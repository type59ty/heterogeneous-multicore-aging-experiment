// Verilog
// c5315
// Ninputs 178
// Noutputs 123
// NtotalGates 2307
// BUFF1 313
// AND2 319
// NOT1 581
// NAND2 454
// AND4 27
// OR2 95
// AND3 359
// OR3 50
// OR4 61
// NOR2 19
// AND5 11
// OR5 8
// NOR3 6
// NOR4 2
// AND9 2

module c5315d (N11,N14,N111,N114,N117,N120,N123,N124,N125,N126,
               N127,N131,N134,N137,N140,N143,N146,N149,N152,N153,
               N154,N161,N164,N167,N170,N173,N176,N179,N180,N181,
               N182,N183,N186,N187,N188,N191,N194,N197,N1100,N1103,
               N1106,N1109,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,
               N1120,N1121,N1122,N1123,N1126,N1127,N1128,N1129,N1130,N1131,
               N1132,N1135,N1136,N1137,N1140,N1141,N1145,N1146,N1149,N1152,
               N1155,N1158,N1161,N1164,N1167,N1170,N1173,N1176,N1179,N1182,
               N1185,N1188,N1191,N1194,N1197,N1200,N1203,N1206,N1209,N1210,
               N1217,N1218,N1225,N1226,N1233,N1234,N1241,N1242,N1245,N1248,
               N1251,N1254,N1257,N1264,N1265,N1272,N1273,N1280,N1281,N1288,
               N1289,N1292,N1293,N1299,N1302,N1307,N1308,N1315,N1316,N1323,
               N1324,N1331,N1332,N1335,N1338,N1341,N1348,N1351,N1358,N1361,
               N1366,N1369,N1372,N1373,N1374,N1386,N1389,N1400,N1411,N1422,
               N1435,N1446,N1457,N1468,N1479,N1490,N1503,N1514,N1523,N1534,
               N1545,N1549,N1552,N1556,N1559,N1562,N1566,N1571,N1574,N1577,
               N1580,N1583,N1588,N1591,N1592,N1595,N1596,N1597,N1598,N1599,
               N1603,N1607,N1610,N1613,N1616,N1619,N1625,N1631,N1709,N1816,
               N11066,N11137,N11138,N11139,N11140,N11141,N11142,N11143,N11144,N11145,
               N11147,N11152,N11153,N11154,N11155,N11972,N12054,N12060,N12061,N12139,
               N12142,N12309,N12387,N12527,N12584,N12590,N12623,N13357,N13358,N13359,
               N13360,N13604,N13613,N14272,N14275,N14278,N14279,N14737,N14738,N14739,
               N14740,N15240,N15388,N16641,N16643,N16646,N16648,N16716,N16877,N16924,
               N16925,N16926,N16927,N17015,N17363,N17365,N17432,N17449,N17465,N17466,
               N17467,N17469,N17470,N17471,N17472,N17473,N17474,N17476,N17503,N17504,
               N17506,N17511,N17515,N17516,N17517,N17518,N17519,N17520,N17521,N17522,
               N17600,N17601,N17602,N17603,N17604,N17605,N17606,N17607,N17626,N17698,
               N17699,N17700,N17701,N17702,N17703,N17704,N17705,N17706,N17707,N17735,
               N17736,N17737,N17738,N17739,N17740,N17741,N17742,N17754,N17755,N17756,
               N17757,N17758,N17759,N17760,N17761,N18075,N18076,N18123,N18124,N18127,
               N18128,
               N21,N24,N211,N214,N217,N220,N223,N224,N225,N226,
               N227,N231,N234,N237,N240,N243,N246,N249,N252,N253,
               N254,N261,N264,N267,N270,N273,N276,N279,N280,N281,
               N282,N283,N286,N287,N288,N291,N294,N297,N2100,N2103,
               N2106,N2109,N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,
               N2120,N2121,N2122,N2123,N2126,N2127,N2128,N2129,N2130,N2131,
               N2132,N2135,N2136,N2137,N2140,N2141,N2145,N2146,N2149,N2152,
               N2155,N2158,N2161,N2164,N2167,N2170,N2173,N2176,N2179,N2182,
               N2185,N2188,N2191,N2194,N2197,N2200,N2203,N2206,N2209,N2210,
               N2217,N2218,N2225,N2226,N2233,N2234,N2241,N2242,N2245,N2248,
               N2251,N2254,N2257,N2264,N2265,N2272,N2273,N2280,N2281,N2288,
               N2289,N2292,N2293,N2299,N2302,N2307,N2308,N2315,N2316,N2323,
               N2324,N2331,N2332,N2335,N2338,N2341,N2348,N2351,N2358,N2361,
               N2366,N2369,N2372,N2373,N2374,N2386,N2389,N2400,N2411,N2422,
               N2435,N2446,N2457,N2468,N2479,N2490,N2503,N2514,N2523,N2534,
               N2545,N2549,N2552,N2556,N2559,N2562,N2566,N2571,N2574,N2577,
               N2580,N2583,N2588,N2591,N2592,N2595,N2596,N2597,N2598,N2599,
               N2603,N2607,N2610,N2613,N2616,N2619,N2625,N2631,N2709,N2816,
               N21066,N21137,N21138,N21139,N21140,N21141,N21142,N21143,N21144,N21145,
               N21147,N21152,N21153,N21154,N21155,N21972,N22054,N22060,N22061,N22139,
               N22142,N22309,N22387,N22527,N22584,N22590,N22623,N23357,N23358,N23359,
               N23360,N23604,N23613,N24272,N24275,N24278,N24279,N24737,N24738,N24739,
               N24740,N25240,N25388,N26641,N26643,N26646,N26648,N26716,N26877,N26924,
               N26925,N26926,N26927,N27015,N27363,N27365,N27432,N27449,N27465,N27466,
               N27467,N27469,N27470,N27471,N27472,N27473,N27474,N27476,N27503,N27504,
               N27506,N27511,N27515,N27516,N27517,N27518,N27519,N27520,N27521,N27522,
               N27600,N27601,N27602,N27603,N27604,N27605,N27606,N27607,N27626,N27698,
               N27699,N27700,N27701,N27702,N27703,N27704,N27705,N27706,N27707,N27735,
               N27736,N27737,N27738,N27739,N27740,N27741,N27742,N27754,N27755,N27756,
               N27757,N27758,N27759,N27760,N27761,N28075,N28076,N28123,N28124,N28127,
               N28128);

input N11,N14,N111,N114,N117,N120,N123,N124,N125,N126,
      N127,N131,N134,N137,N140,N143,N146,N149,N152,N153,
      N154,N161,N164,N167,N170,N173,N176,N179,N180,N181,
      N182,N183,N186,N187,N188,N191,N194,N197,N1100,N1103,
      N1106,N1109,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,
      N1120,N1121,N1122,N1123,N1126,N1127,N1128,N1129,N1130,N1131,
      N1132,N1135,N1136,N1137,N1140,N1141,N1145,N1146,N1149,N1152,
      N1155,N1158,N1161,N1164,N1167,N1170,N1173,N1176,N1179,N1182,
      N1185,N1188,N1191,N1194,N1197,N1200,N1203,N1206,N1209,N1210,
      N1217,N1218,N1225,N1226,N1233,N1234,N1241,N1242,N1245,N1248,
      N1251,N1254,N1257,N1264,N1265,N1272,N1273,N1280,N1281,N1288,
      N1289,N1292,N1293,N1299,N1302,N1307,N1308,N1315,N1316,N1323,
      N1324,N1331,N1332,N1335,N1338,N1341,N1348,N1351,N1358,N1361,
      N1366,N1369,N1372,N1373,N1374,N1386,N1389,N1400,N1411,N1422,
      N1435,N1446,N1457,N1468,N1479,N1490,N1503,N1514,N1523,N1534,
      N1545,N1549,N1552,N1556,N1559,N1562,N1566,N1571,N1574,N1577,
      N1580,N1583,N1588,N1591,N1592,N1595,N1596,N1597,N1598,N1599,
      N1603,N1607,N1610,N1613,N1616,N1619,N1625,N1631,
      N21,N24,N211,N214,N217,N220,N223,N224,N225,N226,
      N227,N231,N234,N237,N240,N243,N246,N249,N252,N253,
      N254,N261,N264,N267,N270,N273,N276,N279,N280,N281,
      N282,N283,N286,N287,N288,N291,N294,N297,N2100,N2103,
      N2106,N2109,N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,
      N2120,N2121,N2122,N2123,N2126,N2127,N2128,N2129,N2130,N2131,
      N2132,N2135,N2136,N2137,N2140,N2141,N2145,N2146,N2149,N2152,
      N2155,N2158,N2161,N2164,N2167,N2170,N2173,N2176,N2179,N2182,
      N2185,N2188,N2191,N2194,N2197,N2200,N2203,N2206,N2209,N2210,
      N2217,N2218,N2225,N2226,N2233,N2234,N2241,N2242,N2245,N2248,
      N2251,N2254,N2257,N2264,N2265,N2272,N2273,N2280,N2281,N2288,
      N2289,N2292,N2293,N2299,N2302,N2307,N2308,N2315,N2316,N2323,
      N2324,N2331,N2332,N2335,N2338,N2341,N2348,N2351,N2358,N2361,
      N2366,N2369,N2372,N2373,N2374,N2386,N2389,N2400,N2411,N2422,
      N2435,N2446,N2457,N2468,N2479,N2490,N2503,N2514,N2523,N2534,
      N2545,N2549,N2552,N2556,N2559,N2562,N2566,N2571,N2574,N2577,
      N2580,N2583,N2588,N2591,N2592,N2595,N2596,N2597,N2598,N2599,
      N2603,N2607,N2610,N2613,N2616,N2619,N2625,N2631;

output N1709,N1816,N11066,N11137,N11138,N11139,N11140,N11141,N11142,N11143,
       N11144,N11145,N11147,N11152,N11153,N11154,N11155,N11972,N12054,N12060,
       N12061,N12139,N12142,N12309,N12387,N12527,N12584,N12590,N12623,N13357,
       N13358,N13359,N13360,N13604,N13613,N14272,N14275,N14278,N14279,N14737,
       N14738,N14739,N14740,N15240,N15388,N16641,N16643,N16646,N16648,N16716,
       N16877,N16924,N16925,N16926,N16927,N17015,N17363,N17365,N17432,N17449,
       N17465,N17466,N17467,N17469,N17470,N17471,N17472,N17473,N17474,N17476,
       N17503,N17504,N17506,N17511,N17515,N17516,N17517,N17518,N17519,N17520,
       N17521,N17522,N17600,N17601,N17602,N17603,N17604,N17605,N17606,N17607,
       N17626,N17698,N17699,N17700,N17701,N17702,N17703,N17704,N17705,N17706,
       N17707,N17735,N17736,N17737,N17738,N17739,N17740,N17741,N17742,N17754,
       N17755,N17756,N17757,N17758,N17759,N17760,N17761,N18075,N18076,N18123,
       N18124,N18127,N18128,
       N2709,N2816,N21066,N21137,N21138,N21139,N21140,N21141,N21142,N21143,
       N21144,N21145,N21147,N21152,N21153,N21154,N21155,N21972,N22054,N22060,
       N22061,N22139,N22142,N22309,N22387,N22527,N22584,N22590,N22623,N23357,
       N23358,N23359,N23360,N23604,N23613,N24272,N24275,N24278,N24279,N24737,
       N24738,N24739,N24740,N25240,N25388,N26641,N26643,N26646,N26648,N26716,
       N26877,N26924,N26925,N26926,N26927,N27015,N27363,N27365,N27432,N27449,
       N27465,N27466,N27467,N27469,N27470,N27471,N27472,N27473,N27474,N27476,
       N27503,N27504,N27506,N27511,N27515,N27516,N27517,N27518,N27519,N27520,
       N27521,N27522,N27600,N27601,N27602,N27603,N27604,N27605,N27606,N27607,
       N27626,N27698,N27699,N27700,N27701,N27702,N27703,N27704,N27705,N27706,
       N27707,N27735,N27736,N27737,N27738,N27739,N27740,N27741,N27742,N27754,
       N27755,N27756,N27757,N27758,N27759,N27760,N27761,N28075,N28076,N28123,
       N28124,N28127,N28128;

wire N11042,N11043,N11067,N11080,N11092,N11104,N11146,N11148,N11149,N11150,
     N11151,N11156,N11157,N11161,N11173,N11185,N11197,N11209,N11213,N11216,
     N11219,N11223,N11235,N11247,N11259,N11271,N11280,N11292,N11303,N11315,
     N11327,N11339,N11351,N11363,N11375,N11378,N11381,N11384,N11387,N11390,
     N11393,N11396,N11415,N11418,N11421,N11424,N11427,N11430,N11433,N11436,
     N11455,N11462,N11469,N11475,N11479,N11482,N11492,N11495,N11498,N11501,
     N11504,N11507,N11510,N11513,N11516,N11519,N11522,N11525,N11542,N11545,
     N11548,N11551,N11554,N11557,N11560,N11563,N11566,N11573,N11580,N11583,
     N11588,N11594,N11597,N11600,N11603,N11606,N11609,N11612,N11615,N11618,
     N11621,N11624,N11627,N11630,N11633,N11636,N11639,N11642,N11645,N11648,
     N11651,N11654,N11657,N11660,N11663,N11675,N11685,N11697,N11709,N11721,
     N11727,N11731,N11743,N11755,N11758,N11761,N11769,N11777,N11785,N11793,
     N11800,N11807,N11814,N11821,N11824,N11827,N11830,N11833,N11836,N11839,
     N11842,N11845,N11848,N11851,N11854,N11857,N11860,N11863,N11866,N11869,
     N11872,N11875,N11878,N11881,N11884,N11887,N11890,N11893,N11896,N11899,
     N11902,N11905,N11908,N11911,N11914,N11917,N11920,N11923,N11926,N11929,
     N11932,N11935,N11938,N11941,N11944,N11947,N11950,N11953,N11956,N11959,
     N11962,N11965,N11968,N12349,N12350,N12585,N12586,N12587,N12588,N12589,
     N12591,N12592,N12593,N12594,N12595,N12596,N12597,N12598,N12599,N12600,
     N12601,N12602,N12603,N12604,N12605,N12606,N12607,N12608,N12609,N12610,
     N12611,N12612,N12613,N12614,N12615,N12616,N12617,N12618,N12619,N12620,
     N12621,N12622,N12624,N12625,N12626,N12627,N12628,N12629,N12630,N12631,
     N12632,N12633,N12634,N12635,N12636,N12637,N12638,N12639,N12640,N12641,
     N12642,N12643,N12644,N12645,N12646,N12647,N12653,N12664,N12675,N12681,
     N12692,N12703,N12704,N12709,N12710,N12711,N12712,N12713,N12714,N12715,
     N12716,N12717,N12718,N12719,N12720,N12721,N12722,N12728,N12739,N12750,
     N12756,N12767,N12778,N12779,N12790,N12801,N12812,N12823,N12824,N12825,
     N12826,N12827,N12828,N12829,N12830,N12831,N12832,N12833,N12834,N12835,
     N12836,N12837,N12838,N12839,N12840,N12841,N12842,N12843,N12844,N12845,
     N12846,N12847,N12848,N12849,N12850,N12851,N12852,N12853,N12854,N12855,
     N12861,N12867,N12868,N12869,N12870,N12871,N12872,N12873,N12874,N12875,
     N12876,N12877,N12882,N12891,N12901,N12902,N12903,N12904,N12905,N12906,
     N12907,N12908,N12909,N12910,N12911,N12912,N12913,N12914,N12915,N12916,
     N12917,N12918,N12919,N12920,N12921,N12922,N12923,N12924,N12925,N12926,
     N12927,N12928,N12929,N12930,N12931,N12932,N12933,N12934,N12935,N12936,
     N12937,N12938,N12939,N12940,N12941,N12942,N12948,N12954,N12955,N12956,
     N12957,N12958,N12959,N12960,N12961,N12962,N12963,N12964,N12969,N12970,
     N12971,N12972,N12973,N12974,N12975,N12976,N12977,N12978,N12979,N12980,
     N12981,N12982,N12983,N12984,N12985,N12986,N12987,N12988,N12989,N12990,
     N12991,N12992,N12993,N12994,N12995,N12996,N12997,N12998,N12999,N13000,
     N13003,N13006,N13007,N13010,N13013,N13014,N13015,N13016,N13017,N13018,
     N13019,N13020,N13021,N13022,N13023,N13024,N13025,N13026,N13027,N13028,
     N13029,N13030,N13031,N13032,N13033,N13034,N13035,N13038,N13041,N13052,
     N13063,N13068,N13071,N13072,N13073,N13074,N13075,N13086,N13097,N13108,
     N13119,N13130,N13141,N13142,N13143,N13144,N13145,N13146,N13147,N13158,
     N13169,N13180,N13191,N13194,N13195,N13196,N13197,N13198,N13199,N13200,
     N13203,N13401,N13402,N13403,N13404,N13405,N13406,N13407,N13408,N13409,
     N13410,N13411,N13412,N13413,N13414,N13415,N13416,N13444,N13445,N13446,
     N13447,N13448,N13449,N13450,N13451,N13452,N13453,N13454,N13455,N13456,
     N13459,N13460,N13461,N13462,N13463,N13464,N13465,N13466,N13481,N13482,
     N13483,N13484,N13485,N13486,N13487,N13488,N13489,N13490,N13491,N13492,
     N13493,N13502,N13503,N13504,N13505,N13506,N13507,N13508,N13509,N13510,
     N13511,N13512,N13513,N13514,N13515,N13558,N13559,N13560,N13561,N13562,
     N13563,N13605,N13606,N13607,N13608,N13609,N13610,N13614,N13615,N13616,
     N13617,N13618,N13619,N13620,N13621,N13622,N13623,N13624,N13625,N13626,
     N13627,N13628,N13629,N13630,N13631,N13632,N13633,N13634,N13635,N13636,
     N13637,N13638,N13639,N13640,N13641,N13642,N13643,N13644,N13645,N13646,
     N13647,N13648,N13649,N13650,N13651,N13652,N13653,N13654,N13655,N13656,
     N13657,N13658,N13659,N13660,N13661,N13662,N13663,N13664,N13665,N13666,
     N13667,N13668,N13669,N13670,N13671,N13672,N13673,N13674,N13675,N13676,
     N13677,N13678,N13679,N13680,N13681,N13682,N13683,N13684,N13685,N13686,
     N13687,N13688,N13689,N13691,N13700,N13701,N13702,N13703,N13704,N13705,
     N13708,N13709,N13710,N13711,N13712,N13713,N13715,N13716,N13717,N13718,
     N13719,N13720,N13721,N13722,N13723,N13724,N13725,N13726,N13727,N13728,
     N13729,N13730,N13731,N13732,N13738,N13739,N13740,N13741,N13742,N13743,
     N13744,N13745,N13746,N13747,N13748,N13749,N13750,N13751,N13752,N13753,
     N13754,N13755,N13756,N13757,N13758,N13759,N13760,N13761,N13762,N13763,
     N13764,N13765,N13766,N13767,N13768,N13769,N13770,N13771,N13775,N13779,
     N13780,N13781,N13782,N13783,N13784,N13785,N13786,N13787,N13788,N13789,
     N13793,N13797,N13800,N13801,N13802,N13803,N13804,N13805,N13806,N13807,
     N13808,N13809,N13810,N13813,N13816,N13819,N13822,N13823,N13824,N13827,
     N13828,N13829,N13830,N13831,N13834,N13835,N13836,N13837,N13838,N13839,
     N13840,N13841,N13842,N13849,N13855,N13861,N13867,N13873,N13881,N13887,
     N13893,N13908,N13909,N13911,N13914,N13915,N13916,N13917,N13918,N13919,
     N13920,N13921,N13927,N13933,N13942,N13948,N13956,N13962,N13968,N13975,
     N13976,N13977,N13978,N13979,N13980,N13981,N13982,N13983,N13984,N13987,
     N13988,N13989,N13990,N13991,N13998,N14008,N14011,N14021,N14024,N14027,
     N14031,N14032,N14033,N14034,N14035,N14036,N14037,N14038,N14039,N14040,
     N14041,N14042,N14067,N14080,N14088,N14091,N14094,N14097,N14100,N14103,
     N14106,N14109,N14144,N14147,N14150,N14153,N14156,N14159,N14183,N14184,
     N14185,N14186,N14188,N14191,N14196,N14197,N14198,N14199,N14200,N14203,
     N14206,N14209,N14212,N14215,N14219,N14223,N14224,N14225,N14228,N14231,
     N14234,N14237,N14240,N14243,N14246,N14249,N14252,N14255,N14258,N14263,
     N14264,N14267,N14268,N14269,N14270,N14271,N14273,N14274,N14276,N14277,
     N14280,N14284,N14290,N14297,N14298,N14301,N14305,N14310,N14316,N14320,
     N14325,N14331,N14332,N14336,N14342,N14349,N14357,N14364,N14375,N14379,
     N14385,N14392,N14396,N14400,N14405,N14412,N14418,N14425,N14436,N14440,
     N14445,N14451,N14456,N14462,N14469,N14477,N14512,N14515,N14516,N14521,
     N14523,N14524,N14532,N14547,N14548,N14551,N14554,N14557,N14560,N14563,
     N14566,N14569,N14572,N14575,N14578,N14581,N14584,N14587,N14590,N14593,
     N14596,N14599,N14602,N14605,N14608,N14611,N14614,N14617,N14621,N14624,
     N14627,N14630,N14633,N14637,N14640,N14643,N14646,N14649,N14652,N14655,
     N14658,N14662,N14665,N14668,N14671,N14674,N14677,N14680,N14683,N14686,
     N14689,N14692,N14695,N14698,N14701,N14702,N14720,N14721,N14724,N14725,
     N14726,N14727,N14728,N14729,N14730,N14731,N14732,N14733,N14734,N14735,
     N14736,N14741,N14855,N14856,N14908,N14909,N14939,N14942,N14947,N14953,
     N14954,N14955,N14956,N14957,N14958,N14959,N14960,N14961,N14965,N14966,
     N14967,N14968,N14972,N14973,N14974,N14975,N14976,N14977,N14978,N14979,
     N14980,N14981,N14982,N14983,N14984,N14985,N14986,N14987,N15049,N15052,
     N15053,N15054,N15055,N15056,N15057,N15058,N15059,N15060,N15061,N15062,
     N15063,N15065,N15066,N15067,N15068,N15069,N15070,N15071,N15072,N15073,
     N15074,N15075,N15076,N15077,N15078,N15079,N15080,N15081,N15082,N15083,
     N15084,N15085,N15086,N15087,N15088,N15089,N15090,N15091,N15092,N15093,
     N15094,N15095,N15096,N15097,N15098,N15099,N15100,N15101,N15102,N15103,
     N15104,N15105,N15106,N15107,N15108,N15109,N15110,N15111,N15112,N15113,
     N15114,N15115,N15116,N15117,N15118,N15119,N15120,N15121,N15122,N15123,
     N15124,N15125,N15126,N15127,N15128,N15129,N15130,N15131,N15132,N15133,
     N15135,N15136,N15137,N15138,N15139,N15140,N15141,N15142,N15143,N15144,
     N15145,N15146,N15147,N15148,N15150,N15153,N15154,N15155,N15156,N15157,
     N15160,N15161,N15162,N15163,N15164,N15165,N15166,N15169,N15172,N15173,
     N15176,N15177,N15180,N15183,N15186,N15189,N15192,N15195,N15198,N15199,
     N15202,N15205,N15208,N15211,N15214,N15217,N15220,N15223,N15224,N15225,
     N15226,N15227,N15228,N15229,N15230,N15232,N15233,N15234,N15235,N15236,
     N15239,N15241,N15242,N15243,N15244,N15245,N15246,N15247,N15248,N15249,
     N15250,N15252,N15253,N15254,N15255,N15256,N15257,N15258,N15259,N15260,
     N15261,N15262,N15263,N15264,N15274,N15275,N15282,N15283,N15284,N15298,
     N15299,N15300,N15303,N15304,N15305,N15306,N15307,N15308,N15309,N15310,
     N15311,N15312,N15315,N15319,N15324,N15328,N15331,N15332,N15346,N15363,
     N15364,N15365,N15366,N15367,N15368,N15369,N15370,N15371,N15374,N15377,
     N15382,N15385,N15389,N15396,N15407,N15418,N15424,N15431,N15441,N15452,
     N15462,N15469,N15470,N15477,N15488,N15498,N15506,N15520,N15536,N15549,
     N15555,N15562,N15573,N15579,N15595,N15606,N15616,N15617,N15618,N15619,
     N15620,N15621,N15622,N15624,N15634,N15655,N15671,N15684,N15690,N15691,
     N15692,N15696,N15700,N15703,N15707,N15711,N15726,N15727,N15728,N15730,
     N15731,N15732,N15733,N15734,N15735,N15736,N15739,N15742,N15745,N15755,
     N15756,N15954,N15955,N15956,N16005,N16006,N16023,N16024,N16025,N16028,
     N16031,N16034,N16037,N16040,N16044,N16045,N16048,N16051,N16054,N16065,
     N16066,N16067,N16068,N16069,N16071,N16072,N16073,N16074,N16075,N16076,
     N16077,N16078,N16079,N16080,N16083,N16084,N16085,N16086,N16087,N16088,
     N16089,N16090,N16091,N16094,N16095,N16096,N16097,N16098,N16099,N16100,
     N16101,N16102,N16103,N16104,N16105,N16106,N16107,N16108,N16111,N16112,
     N16113,N16114,N16115,N16116,N16117,N16120,N16121,N16122,N16123,N16124,
     N16125,N16126,N16127,N16128,N16129,N16130,N16131,N16132,N16133,N16134,
     N16135,N16136,N16137,N16138,N16139,N16140,N16143,N16144,N16145,N16146,
     N16147,N16148,N16149,N16152,N16153,N16154,N16155,N16156,N16157,N16158,
     N16159,N16160,N16161,N16162,N16163,N16164,N16168,N16171,N16172,N16173,
     N16174,N16175,N16178,N16179,N16180,N16181,N16182,N16183,N16184,N16185,
     N16186,N16187,N16188,N16189,N16190,N16191,N16192,N16193,N16194,N16197,
     N16200,N16203,N16206,N16209,N16212,N16215,N16218,N16221,N16234,N16235,
     N16238,N16241,N16244,N16247,N16250,N16253,N16256,N16259,N16262,N16265,
     N16268,N16271,N16274,N16277,N16280,N16283,N16286,N16289,N16292,N16295,
     N16298,N16301,N16304,N16307,N16310,N16313,N16316,N16319,N16322,N16325,
     N16328,N16331,N16335,N16338,N16341,N16344,N16347,N16350,N16353,N16356,
     N16359,N16364,N16367,N16370,N16373,N16374,N16375,N16376,N16377,N16378,
     N16382,N16386,N16388,N16392,N16397,N16411,N16415,N16419,N16427,N16434,
     N16437,N16441,N16445,N16448,N16449,N16466,N16469,N16470,N16471,N16472,
     N16473,N16474,N16475,N16476,N16477,N16478,N16482,N16486,N16490,N16494,
     N16500,N16504,N16508,N16512,N16516,N16526,N16536,N16539,N16553,N16556,
     N16566,N16569,N16572,N16575,N16580,N16584,N16587,N16592,N16599,N16606,
     N16609,N16619,N16622,N16630,N16631,N16632,N16633,N16634,N16637,N16640,
     N16650,N16651,N16653,N16655,N16657,N16659,N16660,N16661,N16662,N16663,
     N16664,N16666,N16668,N16670,N16672,N16675,N16680,N16681,N16682,N16683,
     N16689,N16690,N16691,N16692,N16693,N16695,N16698,N16699,N16700,N16703,
     N16708,N16709,N16710,N16711,N16712,N16713,N16714,N16715,N16718,N16719,
     N16720,N16721,N16722,N16724,N16739,N16740,N16741,N16744,N16745,N16746,
     N16751,N16752,N16753,N16754,N16755,N16760,N16761,N16762,N16772,N16773,
     N16776,N16777,N16782,N16783,N16784,N16785,N16790,N16791,N16792,N16795,
     N16801,N16802,N16803,N16804,N16805,N16806,N16807,N16808,N16809,N16810,
     N16811,N16812,N16813,N16814,N16815,N16816,N16817,N16823,N16824,N16825,
     N16826,N16827,N16828,N16829,N16830,N16831,N16834,N16835,N16836,N16837,
     N16838,N16839,N16840,N16841,N16842,N16843,N16844,N16850,N16851,N16852,
     N16853,N16854,N16855,N16856,N16857,N16860,N16861,N16862,N16863,N16866,
     N16872,N16873,N16874,N16875,N16876,N16879,N16880,N16881,N16884,N16885,
     N16888,N16889,N16890,N16891,N16894,N16895,N16896,N16897,N16900,N16901,
     N16904,N16905,N16908,N16909,N16912,N16913,N16914,N16915,N16916,N16919,
     N16922,N16923,N16930,N16932,N16935,N16936,N16937,N16938,N16939,N16940,
     N16946,N16947,N16948,N16949,N16953,N16954,N16955,N16956,N16957,N16958,
     N16964,N16965,N16966,N16967,N16973,N16974,N16975,N16976,N16977,N16978,
     N16979,N16987,N16990,N16999,N17002,N17003,N17006,N17011,N17012,N17013,
     N17016,N17018,N17019,N17020,N17021,N17022,N17023,N17028,N17031,N17034,
     N17037,N17040,N17041,N17044,N17045,N17046,N17047,N17048,N17049,N17054,
     N17057,N17060,N17064,N17065,N17072,N17073,N17074,N17075,N17076,N17079,
     N17080,N17083,N17084,N17085,N17086,N17087,N17088,N17089,N17090,N17093,
     N17094,N17097,N17101,N17105,N17110,N17114,N17115,N17116,N17125,N17126,
     N17127,N17130,N17131,N17139,N17140,N17141,N17146,N17147,N17149,N17150,
     N17151,N17152,N17153,N17158,N17159,N17160,N17166,N17167,N17168,N17169,
     N17170,N17171,N17172,N17173,N17174,N17175,N17176,N17177,N17178,N17179,
     N17180,N17181,N17182,N17183,N17184,N17185,N17186,N17187,N17188,N17189,
     N17190,N17196,N17197,N17198,N17204,N17205,N17206,N17207,N17208,N17209,
     N17212,N17215,N17216,N17217,N17218,N17219,N17222,N17225,N17228,N17229,
     N17236,N17239,N17242,N17245,N17250,N17257,N17260,N17263,N17268,N17269,
     N17270,N17276,N17282,N17288,N17294,N17300,N17301,N17304,N17310,N17320,
     N17321,N17328,N17338,N17339,N17340,N17341,N17342,N17349,N17357,N17364,
     N17394,N17397,N17402,N17405,N17406,N17407,N17408,N17409,N17412,N17415,
     N17416,N17417,N17418,N17419,N17420,N17421,N17424,N17425,N17426,N17427,
     N17428,N17429,N17430,N17431,N17433,N17434,N17435,N17436,N17437,N17438,
     N17439,N17440,N17441,N17442,N17443,N17444,N17445,N17446,N17447,N17448,
     N17450,N17451,N17452,N17453,N17454,N17455,N17456,N17457,N17458,N17459,
     N17460,N17461,N17462,N17463,N17464,N17468,N17479,N17481,N17482,N17483,
     N17484,N17485,N17486,N17487,N17488,N17489,N17492,N17493,N17498,N17499,
     N17500,N17505,N17507,N17508,N17509,N17510,N17512,N17513,N17514,N17525,
     N17526,N17527,N17528,N17529,N17530,N17531,N17537,N17543,N17549,N17555,
     N17561,N17567,N17573,N17579,N17582,N17585,N17586,N17587,N17588,N17589,
     N17592,N17595,N17598,N17599,N17624,N17625,N17631,N17636,N17657,N17658,
     N17665,N17666,N17667,N17668,N17669,N17670,N17671,N17672,N17673,N17674,
     N17675,N17676,N17677,N17678,N17679,N17680,N17681,N17682,N17683,N17684,
     N17685,N17686,N17687,N17688,N17689,N17690,N17691,N17692,N17693,N17694,
     N17695,N17696,N17697,N17708,N17709,N17710,N17711,N17712,N17715,N17718,
     N17719,N17720,N17721,N17722,N17723,N17724,N17727,N17728,N17729,N17730,
     N17731,N17732,N17733,N17734,N17743,N17744,N17749,N17750,N17751,N17762,
     N17765,N17768,N17769,N17770,N17771,N17772,N17775,N17778,N17781,N17782,
     N17787,N17788,N17795,N17796,N17797,N17798,N17799,N17800,N17803,N17806,
     N17807,N17808,N17809,N17810,N17811,N17812,N17815,N17816,N17821,N17822,
     N17823,N17826,N17829,N17832,N17833,N17834,N17835,N17836,N17839,N17842,
     N17845,N17846,N17851,N17852,N17859,N17860,N17861,N17862,N17863,N17864,
     N17867,N17870,N17871,N17872,N17873,N17874,N17875,N17876,N17879,N17880,
     N17885,N17886,N17887,N17890,N17893,N17896,N17897,N17898,N17899,N17900,
     N17903,N17906,N17909,N17910,N17917,N17918,N17923,N17924,N17925,N17926,
     N17927,N17928,N17929,N17930,N17931,N17932,N17935,N17938,N17939,N17940,
     N17943,N17944,N17945,N17946,N17951,N17954,N17957,N17960,N17963,N17966,
     N17967,N17968,N17969,N17970,N17973,N17974,N17984,N17985,N17987,N17988,
     N17989,N17990,N17991,N17992,N17993,N17994,N17995,N17996,N17997,N17998,
     N18001,N18004,N18009,N18013,N18017,N18020,N18021,N18022,N18023,N18025,
     N18026,N18027,N18031,N18032,N18033,N18034,N18035,N18036,N18037,N18038,
     N18039,N18040,N18041,N18042,N18043,N18044,N18045,N18048,N18055,N18056,
     N18057,N18058,N18059,N18060,N18061,N18064,N18071,N18072,N18073,N18074,
     N18077,N18078,N18079,N18082,N18089,N18090,N18091,N18092,N18093,N18096,
     N18099,N18102,N18113,N18114,N18115,N18116,N18117,N18118,N18119,N18120,
     N18121,N18122,N18125,N18126,

     N21042,N21043,N21067,N21080,N21092,N21104,N21146,N21148,N21149,N21150,
     N21151,N21156,N21157,N21161,N21173,N21185,N21197,N21209,N21213,N21216,
     N21219,N21223,N21235,N21247,N21259,N21271,N21280,N21292,N21303,N21315,
     N21327,N21339,N21351,N21363,N21375,N21378,N21381,N21384,N21387,N21390,
     N21393,N21396,N21415,N21418,N21421,N21424,N21427,N21430,N21433,N21436,
     N21455,N21462,N21469,N21475,N21479,N21482,N21492,N21495,N21498,N21501,
     N21504,N21507,N21510,N21513,N21516,N21519,N21522,N21525,N21542,N21545,
     N21548,N21551,N21554,N21557,N21560,N21563,N21566,N21573,N21580,N21583,
     N21588,N21594,N21597,N21600,N21603,N21606,N21609,N21612,N21615,N21618,
     N21621,N21624,N21627,N21630,N21633,N21636,N21639,N21642,N21645,N21648,
     N21651,N21654,N21657,N21660,N21663,N21675,N21685,N21697,N21709,N21721,
     N21727,N21731,N21743,N21755,N21758,N21761,N21769,N21777,N21785,N21793,
     N21800,N21807,N21814,N21821,N21824,N21827,N21830,N21833,N21836,N21839,
     N21842,N21845,N21848,N21851,N21854,N21857,N21860,N21863,N21866,N21869,
     N21872,N21875,N21878,N21881,N21884,N21887,N21890,N21893,N21896,N21899,
     N21902,N21905,N21908,N21911,N21914,N21917,N21920,N21923,N21926,N21929,
     N21932,N21935,N21938,N21941,N21944,N21947,N21950,N21953,N21956,N21959,
     N21962,N21965,N21968,N22349,N22350,N22585,N22586,N22587,N22588,N22589,
     N22591,N22592,N22593,N22594,N22595,N22596,N22597,N22598,N22599,N22600,
     N22601,N22602,N22603,N22604,N22605,N22606,N22607,N22608,N22609,N22610,
     N22611,N22612,N22613,N22614,N22615,N22616,N22617,N22618,N22619,N22620,
     N22621,N22622,N22624,N22625,N22626,N22627,N22628,N22629,N22630,N22631,
     N22632,N22633,N22634,N22635,N22636,N22637,N22638,N22639,N22640,N22641,
     N22642,N22643,N22644,N22645,N22646,N22647,N22653,N22664,N22675,N22681,
     N22692,N22703,N22704,N22709,N22710,N22711,N22712,N22713,N22714,N22715,
     N22716,N22717,N22718,N22719,N22720,N22721,N22722,N22728,N22739,N22750,
     N22756,N22767,N22778,N22779,N22790,N22801,N22812,N22823,N22824,N22825,
     N22826,N22827,N22828,N22829,N22830,N22831,N22832,N22833,N22834,N22835,
     N22836,N22837,N22838,N22839,N22840,N22841,N22842,N22843,N22844,N22845,
     N22846,N22847,N22848,N22849,N22850,N22851,N22852,N22853,N22854,N22855,
     N22861,N22867,N22868,N22869,N22870,N22871,N22872,N22873,N22874,N22875,
     N22876,N22877,N22882,N22891,N22901,N22902,N22903,N22904,N22905,N22906,
     N22907,N22908,N22909,N22910,N22911,N22912,N22913,N22914,N22915,N22916,
     N22917,N22918,N22919,N22920,N22921,N22922,N22923,N22924,N22925,N22926,
     N22927,N22928,N22929,N22930,N22931,N22932,N22933,N22934,N22935,N22936,
     N22937,N22938,N22939,N22940,N22941,N22942,N22948,N22954,N22955,N22956,
     N22957,N22958,N22959,N22960,N22961,N22962,N22963,N22964,N22969,N22970,
     N22971,N22972,N22973,N22974,N22975,N22976,N22977,N22978,N22979,N22980,
     N22981,N22982,N22983,N22984,N22985,N22986,N22987,N22988,N22989,N22990,
     N22991,N22992,N22993,N22994,N22995,N22996,N22997,N22998,N22999,N23000,
     N23003,N23006,N23007,N23010,N23013,N23014,N23015,N23016,N23017,N23018,
     N23019,N23020,N23021,N23022,N23023,N23024,N23025,N23026,N23027,N23028,
     N23029,N23030,N23031,N23032,N23033,N23034,N23035,N23038,N23041,N23052,
     N23063,N23068,N23071,N23072,N23073,N23074,N23075,N23086,N23097,N23108,
     N23119,N23130,N23141,N23142,N23143,N23144,N23145,N23146,N23147,N23158,
     N23169,N23180,N23191,N23194,N23195,N23196,N23197,N23198,N23199,N23200,
     N23203,N23401,N23402,N23403,N23404,N23405,N23406,N23407,N23408,N23409,
     N23410,N23411,N23412,N23413,N23414,N23415,N23416,N23444,N23445,N23446,
     N23447,N23448,N23449,N23450,N23451,N23452,N23453,N23454,N23455,N23456,
     N23459,N23460,N23461,N23462,N23463,N23464,N23465,N23466,N23481,N23482,
     N23483,N23484,N23485,N23486,N23487,N23488,N23489,N23490,N23491,N23492,
     N23493,N23502,N23503,N23504,N23505,N23506,N23507,N23508,N23509,N23510,
     N23511,N23512,N23513,N23514,N23515,N23558,N23559,N23560,N23561,N23562,
     N23563,N23605,N23606,N23607,N23608,N23609,N23610,N23614,N23615,N23616,
     N23617,N23618,N23619,N23620,N23621,N23622,N23623,N23624,N23625,N23626,
     N23627,N23628,N23629,N23630,N23631,N23632,N23633,N23634,N23635,N23636,
     N23637,N23638,N23639,N23640,N23641,N23642,N23643,N23644,N23645,N23646,
     N23647,N23648,N23649,N23650,N23651,N23652,N23653,N23654,N23655,N23656,
     N23657,N23658,N23659,N23660,N23661,N23662,N23663,N23664,N23665,N23666,
     N23667,N23668,N23669,N23670,N23671,N23672,N23673,N23674,N23675,N23676,
     N23677,N23678,N23679,N23680,N23681,N23682,N23683,N23684,N23685,N23686,
     N23687,N23688,N23689,N23691,N23700,N23701,N23702,N23703,N23704,N23705,
     N23708,N23709,N23710,N23711,N23712,N23713,N23715,N23716,N23717,N23718,
     N23719,N23720,N23721,N23722,N23723,N23724,N23725,N23726,N23727,N23728,
     N23729,N23730,N23731,N23732,N23738,N23739,N23740,N23741,N23742,N23743,
     N23744,N23745,N23746,N23747,N23748,N23749,N23750,N23751,N23752,N23753,
     N23754,N23755,N23756,N23757,N23758,N23759,N23760,N23761,N23762,N23763,
     N23764,N23765,N23766,N23767,N23768,N23769,N23770,N23771,N23775,N23779,
     N23780,N23781,N23782,N23783,N23784,N23785,N23786,N23787,N23788,N23789,
     N23793,N23797,N23800,N23801,N23802,N23803,N23804,N23805,N23806,N23807,
     N23808,N23809,N23810,N23813,N23816,N23819,N23822,N23823,N23824,N23827,
     N23828,N23829,N23830,N23831,N23834,N23835,N23836,N23837,N23838,N23839,
     N23840,N23841,N23842,N23849,N23855,N23861,N23867,N23873,N23881,N23887,
     N23893,N23908,N23909,N23911,N23914,N23915,N23916,N23917,N23918,N23919,
     N23920,N23921,N23927,N23933,N23942,N23948,N23956,N23962,N23968,N23975,
     N23976,N23977,N23978,N23979,N23980,N23981,N23982,N23983,N23984,N23987,
     N23988,N23989,N23990,N23991,N23998,N24008,N24011,N24021,N24024,N24027,
     N24031,N24032,N24033,N24034,N24035,N24036,N24037,N24038,N24039,N24040,
     N24041,N24042,N24067,N24080,N24088,N24091,N24094,N24097,N24100,N24103,
     N24106,N24109,N24144,N24147,N24150,N24153,N24156,N24159,N24183,N24184,
     N24185,N24186,N24188,N24191,N24196,N24197,N24198,N24199,N24200,N24203,
     N24206,N24209,N24212,N24215,N24219,N24223,N24224,N24225,N24228,N24231,
     N24234,N24237,N24240,N24243,N24246,N24249,N24252,N24255,N24258,N24263,
     N24264,N24267,N24268,N24269,N24270,N24271,N24273,N24274,N24276,N24277,
     N24280,N24284,N24290,N24297,N24298,N24301,N24305,N24310,N24316,N24320,
     N24325,N24331,N24332,N24336,N24342,N24349,N24357,N24364,N24375,N24379,
     N24385,N24392,N24396,N24400,N24405,N24412,N24418,N24425,N24436,N24440,
     N24445,N24451,N24456,N24462,N24469,N24477,N24512,N24515,N24516,N24521,
     N24523,N24524,N24532,N24547,N24548,N24551,N24554,N24557,N24560,N24563,
     N24566,N24569,N24572,N24575,N24578,N24581,N24584,N24587,N24590,N24593,
     N24596,N24599,N24602,N24605,N24608,N24611,N24614,N24617,N24621,N24624,
     N24627,N24630,N24633,N24637,N24640,N24643,N24646,N24649,N24652,N24655,
     N24658,N24662,N24665,N24668,N24671,N24674,N24677,N24680,N24683,N24686,
     N24689,N24692,N24695,N24698,N24701,N24702,N24720,N24721,N24724,N24725,
     N24726,N24727,N24728,N24729,N24730,N24731,N24732,N24733,N24734,N24735,
     N24736,N24741,N24855,N24856,N24908,N24909,N24939,N24942,N24947,N24953,
     N24954,N24955,N24956,N24957,N24958,N24959,N24960,N24961,N24965,N24966,
     N24967,N24968,N24972,N24973,N24974,N24975,N24976,N24977,N24978,N24979,
     N24980,N24981,N24982,N24983,N24984,N24985,N24986,N24987,N25049,N25052,
     N25053,N25054,N25055,N25056,N25057,N25058,N25059,N25060,N25061,N25062,
     N25063,N25065,N25066,N25067,N25068,N25069,N25070,N25071,N25072,N25073,
     N25074,N25075,N25076,N25077,N25078,N25079,N25080,N25081,N25082,N25083,
     N25084,N25085,N25086,N25087,N25088,N25089,N25090,N25091,N25092,N25093,
     N25094,N25095,N25096,N25097,N25098,N25099,N25100,N25101,N25102,N25103,
     N25104,N25105,N25106,N25107,N25108,N25109,N25110,N25111,N25112,N25113,
     N25114,N25115,N25116,N25117,N25118,N25119,N25120,N25121,N25122,N25123,
     N25124,N25125,N25126,N25127,N25128,N25129,N25130,N25131,N25132,N25133,
     N25135,N25136,N25137,N25138,N25139,N25140,N25141,N25142,N25143,N25144,
     N25145,N25146,N25147,N25148,N25150,N25153,N25154,N25155,N25156,N25157,
     N25160,N25161,N25162,N25163,N25164,N25165,N25166,N25169,N25172,N25173,
     N25176,N25177,N25180,N25183,N25186,N25189,N25192,N25195,N25198,N25199,
     N25202,N25205,N25208,N25211,N25214,N25217,N25220,N25223,N25224,N25225,
     N25226,N25227,N25228,N25229,N25230,N25232,N25233,N25234,N25235,N25236,
     N25239,N25241,N25242,N25243,N25244,N25245,N25246,N25247,N25248,N25249,
     N25250,N25252,N25253,N25254,N25255,N25256,N25257,N25258,N25259,N25260,
     N25261,N25262,N25263,N25264,N25274,N25275,N25282,N25283,N25284,N25298,
     N25299,N25300,N25303,N25304,N25305,N25306,N25307,N25308,N25309,N25310,
     N25311,N25312,N25315,N25319,N25324,N25328,N25331,N25332,N25346,N25363,
     N25364,N25365,N25366,N25367,N25368,N25369,N25370,N25371,N25374,N25377,
     N25382,N25385,N25389,N25396,N25407,N25418,N25424,N25431,N25441,N25452,
     N25462,N25469,N25470,N25477,N25488,N25498,N25506,N25520,N25536,N25549,
     N25555,N25562,N25573,N25579,N25595,N25606,N25616,N25617,N25618,N25619,
     N25620,N25621,N25622,N25624,N25634,N25655,N25671,N25684,N25690,N25691,
     N25692,N25696,N25700,N25703,N25707,N25711,N25726,N25727,N25728,N25730,
     N25731,N25732,N25733,N25734,N25735,N25736,N25739,N25742,N25745,N25755,
     N25756,N25954,N25955,N25956,N26005,N26006,N26023,N26024,N26025,N26028,
     N26031,N26034,N26037,N26040,N26044,N26045,N26048,N26051,N26054,N26065,
     N26066,N26067,N26068,N26069,N26071,N26072,N26073,N26074,N26075,N26076,
     N26077,N26078,N26079,N26080,N26083,N26084,N26085,N26086,N26087,N26088,
     N26089,N26090,N26091,N26094,N26095,N26096,N26097,N26098,N26099,N26100,
     N26101,N26102,N26103,N26104,N26105,N26106,N26107,N26108,N26111,N26112,
     N26113,N26114,N26115,N26116,N26117,N26120,N26121,N26122,N26123,N26124,
     N26125,N26126,N26127,N26128,N26129,N26130,N26131,N26132,N26133,N26134,
     N26135,N26136,N26137,N26138,N26139,N26140,N26143,N26144,N26145,N26146,
     N26147,N26148,N26149,N26152,N26153,N26154,N26155,N26156,N26157,N26158,
     N26159,N26160,N26161,N26162,N26163,N26164,N26168,N26171,N26172,N26173,
     N26174,N26175,N26178,N26179,N26180,N26181,N26182,N26183,N26184,N26185,
     N26186,N26187,N26188,N26189,N26190,N26191,N26192,N26193,N26194,N26197,
     N26200,N26203,N26206,N26209,N26212,N26215,N26218,N26221,N26234,N26235,
     N26238,N26241,N26244,N26247,N26250,N26253,N26256,N26259,N26262,N26265,
     N26268,N26271,N26274,N26277,N26280,N26283,N26286,N26289,N26292,N26295,
     N26298,N26301,N26304,N26307,N26310,N26313,N26316,N26319,N26322,N26325,
     N26328,N26331,N26335,N26338,N26341,N26344,N26347,N26350,N26353,N26356,
     N26359,N26364,N26367,N26370,N26373,N26374,N26375,N26376,N26377,N26378,
     N26382,N26386,N26388,N26392,N26397,N26411,N26415,N26419,N26427,N26434,
     N26437,N26441,N26445,N26448,N26449,N26466,N26469,N26470,N26471,N26472,
     N26473,N26474,N26475,N26476,N26477,N26478,N26482,N26486,N26490,N26494,
     N26500,N26504,N26508,N26512,N26516,N26526,N26536,N26539,N26553,N26556,
     N26566,N26569,N26572,N26575,N26580,N26584,N26587,N26592,N26599,N26606,
     N26609,N26619,N26622,N26630,N26631,N26632,N26633,N26634,N26637,N26640,
     N26650,N26651,N26653,N26655,N26657,N26659,N26660,N26661,N26662,N26663,
     N26664,N26666,N26668,N26670,N26672,N26675,N26680,N26681,N26682,N26683,
     N26689,N26690,N26691,N26692,N26693,N26695,N26698,N26699,N26700,N26703,
     N26708,N26709,N26710,N26711,N26712,N26713,N26714,N26715,N26718,N26719,
     N26720,N26721,N26722,N26724,N26739,N26740,N26741,N26744,N26745,N26746,
     N26751,N26752,N26753,N26754,N26755,N26760,N26761,N26762,N26772,N26773,
     N26776,N26777,N26782,N26783,N26784,N26785,N26790,N26791,N26792,N26795,
     N26801,N26802,N26803,N26804,N26805,N26806,N26807,N26808,N26809,N26810,
     N26811,N26812,N26813,N26814,N26815,N26816,N26817,N26823,N26824,N26825,
     N26826,N26827,N26828,N26829,N26830,N26831,N26834,N26835,N26836,N26837,
     N26838,N26839,N26840,N26841,N26842,N26843,N26844,N26850,N26851,N26852,
     N26853,N26854,N26855,N26856,N26857,N26860,N26861,N26862,N26863,N26866,
     N26872,N26873,N26874,N26875,N26876,N26879,N26880,N26881,N26884,N26885,
     N26888,N26889,N26890,N26891,N26894,N26895,N26896,N26897,N26900,N26901,
     N26904,N26905,N26908,N26909,N26912,N26913,N26914,N26915,N26916,N26919,
     N26922,N26923,N26930,N26932,N26935,N26936,N26937,N26938,N26939,N26940,
     N26946,N26947,N26948,N26949,N26953,N26954,N26955,N26956,N26957,N26958,
     N26964,N26965,N26966,N26967,N26973,N26974,N26975,N26976,N26977,N26978,
     N26979,N26987,N26990,N26999,N27002,N27003,N27006,N27011,N27012,N27013,
     N27016,N27018,N27019,N27020,N27021,N27022,N27023,N27028,N27031,N27034,
     N27037,N27040,N27041,N27044,N27045,N27046,N27047,N27048,N27049,N27054,
     N27057,N27060,N27064,N27065,N27072,N27073,N27074,N27075,N27076,N27079,
     N27080,N27083,N27084,N27085,N27086,N27087,N27088,N27089,N27090,N27093,
     N27094,N27097,N27101,N27105,N27110,N27114,N27115,N27116,N27125,N27126,
     N27127,N27130,N27131,N27139,N27140,N27141,N27146,N27147,N27149,N27150,
     N27151,N27152,N27153,N27158,N27159,N27160,N27166,N27167,N27168,N27169,
     N27170,N27171,N27172,N27173,N27174,N27175,N27176,N27177,N27178,N27179,
     N27180,N27181,N27182,N27183,N27184,N27185,N27186,N27187,N27188,N27189,
     N27190,N27196,N27197,N27198,N27204,N27205,N27206,N27207,N27208,N27209,
     N27212,N27215,N27216,N27217,N27218,N27219,N27222,N27225,N27228,N27229,
     N27236,N27239,N27242,N27245,N27250,N27257,N27260,N27263,N27268,N27269,
     N27270,N27276,N27282,N27288,N27294,N27300,N27301,N27304,N27310,N27320,
     N27321,N27328,N27338,N27339,N27340,N27341,N27342,N27349,N27357,N27364,
     N27394,N27397,N27402,N27405,N27406,N27407,N27408,N27409,N27412,N27415,
     N27416,N27417,N27418,N27419,N27420,N27421,N27424,N27425,N27426,N27427,
     N27428,N27429,N27430,N27431,N27433,N27434,N27435,N27436,N27437,N27438,
     N27439,N27440,N27441,N27442,N27443,N27444,N27445,N27446,N27447,N27448,
     N27450,N27451,N27452,N27453,N27454,N27455,N27456,N27457,N27458,N27459,
     N27460,N27461,N27462,N27463,N27464,N27468,N27479,N27481,N27482,N27483,
     N27484,N27485,N27486,N27487,N27488,N27489,N27492,N27493,N27498,N27499,
     N27500,N27505,N27507,N27508,N27509,N27510,N27512,N27513,N27514,N27525,
     N27526,N27527,N27528,N27529,N27530,N27531,N27537,N27543,N27549,N27555,
     N27561,N27567,N27573,N27579,N27582,N27585,N27586,N27587,N27588,N27589,
     N27592,N27595,N27598,N27599,N27624,N27625,N27631,N27636,N27657,N27658,
     N27665,N27666,N27667,N27668,N27669,N27670,N27671,N27672,N27673,N27674,
     N27675,N27676,N27677,N27678,N27679,N27680,N27681,N27682,N27683,N27684,
     N27685,N27686,N27687,N27688,N27689,N27690,N27691,N27692,N27693,N27694,
     N27695,N27696,N27697,N27708,N27709,N27710,N27711,N27712,N27715,N27718,
     N27719,N27720,N27721,N27722,N27723,N27724,N27727,N27728,N27729,N27730,
     N27731,N27732,N27733,N27734,N27743,N27744,N27749,N27750,N27751,N27762,
     N27765,N27768,N27769,N27770,N27771,N27772,N27775,N27778,N27781,N27782,
     N27787,N27788,N27795,N27796,N27797,N27798,N27799,N27800,N27803,N27806,
     N27807,N27808,N27809,N27810,N27811,N27812,N27815,N27816,N27821,N27822,
     N27823,N27826,N27829,N27832,N27833,N27834,N27835,N27836,N27839,N27842,
     N27845,N27846,N27851,N27852,N27859,N27860,N27861,N27862,N27863,N27864,
     N27867,N27870,N27871,N27872,N27873,N27874,N27875,N27876,N27879,N27880,
     N27885,N27886,N27887,N27890,N27893,N27896,N27897,N27898,N27899,N27900,
     N27903,N27906,N27909,N27910,N27917,N27918,N27923,N27924,N27925,N27926,
     N27927,N27928,N27929,N27930,N27931,N27932,N27935,N27938,N27939,N27940,
     N27943,N27944,N27945,N27946,N27951,N27954,N27957,N27960,N27963,N27966,
     N27967,N27968,N27969,N27970,N27973,N27974,N27984,N27985,N27987,N27988,
     N27989,N27990,N27991,N27992,N27993,N27994,N27995,N27996,N27997,N27998,
     N28001,N28004,N28009,N28013,N28017,N28020,N28021,N28022,N28023,N28025,
     N28026,N28027,N28031,N28032,N28033,N28034,N28035,N28036,N28037,N28038,
     N28039,N28040,N28041,N28042,N28043,N28044,N28045,N28048,N28055,N28056,
     N28057,N28058,N28059,N28060,N28061,N28064,N28071,N28072,N28073,N28074,
     N28077,N28078,N28079,N28082,N28089,N28090,N28091,N28092,N28093,N28096,
     N28099,N28102,N28113,N28114,N28115,N28116,N28117,N28118,N28119,N28120,
     N28121,N28122,N28125,N28126;

buf BUFF1_11 (N1709, N1141);
buf BUFF1_12 (N1816, N1293);
and AND2_13 (N11042, N1135, N1631);
not NOT1_14 (N11043, N1591);
buf BUFF1_15 (N11066, N1592);
not NOT1_16 (N11067, N1595);
not NOT1_17 (N11080, N1596);
not NOT1_18 (N11092, N1597);
not NOT1_19 (N11104, N1598);
not NOT1_110 (N11137, N1545);
not NOT1_111 (N11138, N1348);
not NOT1_112 (N11139, N1366);
and AND2_113 (N11140, N1552, N1562);
not NOT1_114 (N11141, N1549);
not NOT1_115 (N11142, N1545);
not NOT1_116 (N11143, N1545);
not NOT1_117 (N11144, N1338);
not NOT1_118 (N11145, N1358);
nand NAND2_119 (N11146, N1373, N11);
and AND2_120 (N11147, N1141, N1145);
not NOT1_121 (N11148, N1592);
not NOT1_122 (N11149, N11042);
and AND2_123 (N11150, N11043, N127);
and AND2_124 (N11151, N1386, N1556);
not NOT1_125 (N11152, N1245);
not NOT1_126 (N11153, N1552);
not NOT1_127 (N11154, N1562);
not NOT1_128 (N11155, N1559);
and AND4_129 (N11156, N1386, N1559, N1556, N1552);
not NOT1_130 (N11157, N1566);
buf BUFF1_131 (N11161, N1571);
buf BUFF1_132 (N11173, N1574);
buf BUFF1_133 (N11185, N1571);
buf BUFF1_134 (N11197, N1574);
buf BUFF1_135 (N11209, N1137);
buf BUFF1_136 (N11213, N1137);
buf BUFF1_137 (N11216, N1141);
not NOT1_138 (N11219, N1583);
buf BUFF1_139 (N11223, N1577);
buf BUFF1_140 (N11235, N1580);
buf BUFF1_141 (N11247, N1577);
buf BUFF1_142 (N11259, N1580);
buf BUFF1_143 (N11271, N1254);
buf BUFF1_144 (N11280, N1251);
buf BUFF1_145 (N11292, N1251);
buf BUFF1_146 (N11303, N1248);
buf BUFF1_147 (N11315, N1248);
buf BUFF1_148 (N11327, N1610);
buf BUFF1_149 (N11339, N1607);
buf BUFF1_150 (N11351, N1613);
buf BUFF1_151 (N11363, N1616);
buf BUFF1_152 (N11375, N1210);
buf BUFF1_153 (N11378, N1210);
buf BUFF1_154 (N11381, N1218);
buf BUFF1_155 (N11384, N1218);
buf BUFF1_156 (N11387, N1226);
buf BUFF1_157 (N11390, N1226);
buf BUFF1_158 (N11393, N1234);
buf BUFF1_159 (N11396, N1234);
buf BUFF1_160 (N11415, N1257);
buf BUFF1_161 (N11418, N1257);
buf BUFF1_162 (N11421, N1265);
buf BUFF1_163 (N11424, N1265);
buf BUFF1_164 (N11427, N1273);
buf BUFF1_165 (N11430, N1273);
buf BUFF1_166 (N11433, N1281);
buf BUFF1_167 (N11436, N1281);
buf BUFF1_168 (N11455, N1335);
buf BUFF1_169 (N11462, N1335);
buf BUFF1_170 (N11469, N1206);
and AND2_171 (N11475, N127, N131);
buf BUFF1_172 (N11479, N11);
buf BUFF1_173 (N11482, N1588);
buf BUFF1_174 (N11492, N1293);
buf BUFF1_175 (N11495, N1302);
buf BUFF1_176 (N11498, N1308);
buf BUFF1_177 (N11501, N1308);
buf BUFF1_178 (N11504, N1316);
buf BUFF1_179 (N11507, N1316);
buf BUFF1_180 (N11510, N1324);
buf BUFF1_181 (N11513, N1324);
buf BUFF1_182 (N11516, N1341);
buf BUFF1_183 (N11519, N1341);
buf BUFF1_184 (N11522, N1351);
buf BUFF1_185 (N11525, N1351);
buf BUFF1_186 (N11542, N1257);
buf BUFF1_187 (N11545, N1257);
buf BUFF1_188 (N11548, N1265);
buf BUFF1_189 (N11551, N1265);
buf BUFF1_190 (N11554, N1273);
buf BUFF1_191 (N11557, N1273);
buf BUFF1_192 (N11560, N1281);
buf BUFF1_193 (N11563, N1281);
buf BUFF1_194 (N11566, N1332);
buf BUFF1_195 (N11573, N1332);
buf BUFF1_196 (N11580, N1549);
and AND2_197 (N11583, N131, N127);
not NOT1_198 (N11588, N1588);
buf BUFF1_199 (N11594, N1324);
buf BUFF1_1100 (N11597, N1324);
buf BUFF1_1101 (N11600, N1341);
buf BUFF1_1102 (N11603, N1341);
buf BUFF1_1103 (N11606, N1351);
buf BUFF1_1104 (N11609, N1351);
buf BUFF1_1105 (N11612, N1293);
buf BUFF1_1106 (N11615, N1302);
buf BUFF1_1107 (N11618, N1308);
buf BUFF1_1108 (N11621, N1308);
buf BUFF1_1109 (N11624, N1316);
buf BUFF1_1110 (N11627, N1316);
buf BUFF1_1111 (N11630, N1361);
buf BUFF1_1112 (N11633, N1361);
buf BUFF1_1113 (N11636, N1210);
buf BUFF1_1114 (N11639, N1210);
buf BUFF1_1115 (N11642, N1218);
buf BUFF1_1116 (N11645, N1218);
buf BUFF1_1117 (N11648, N1226);
buf BUFF1_1118 (N11651, N1226);
buf BUFF1_1119 (N11654, N1234);
buf BUFF1_1120 (N11657, N1234);
not NOT1_1121 (N11660, N1324);
buf BUFF1_1122 (N11663, N1242);
buf BUFF1_1123 (N11675, N1242);
buf BUFF1_1124 (N11685, N1254);
buf BUFF1_1125 (N11697, N1610);
buf BUFF1_1126 (N11709, N1607);
buf BUFF1_1127 (N11721, N1625);
buf BUFF1_1128 (N11727, N1619);
buf BUFF1_1129 (N11731, N1613);
buf BUFF1_1130 (N11743, N1616);
not NOT1_1131 (N11755, N1599);
not NOT1_1132 (N11758, N1603);
buf BUFF1_1133 (N11761, N1619);
buf BUFF1_1134 (N11769, N1625);
buf BUFF1_1135 (N11777, N1619);
buf BUFF1_1136 (N11785, N1625);
buf BUFF1_1137 (N11793, N1619);
buf BUFF1_1138 (N11800, N1625);
buf BUFF1_1139 (N11807, N1619);
buf BUFF1_1140 (N11814, N1625);
buf BUFF1_1141 (N11821, N1299);
buf BUFF1_1142 (N11824, N1446);
buf BUFF1_1143 (N11827, N1457);
buf BUFF1_1144 (N11830, N1468);
buf BUFF1_1145 (N11833, N1422);
buf BUFF1_1146 (N11836, N1435);
buf BUFF1_1147 (N11839, N1389);
buf BUFF1_1148 (N11842, N1400);
buf BUFF1_1149 (N11845, N1411);
buf BUFF1_1150 (N11848, N1374);
buf BUFF1_1151 (N11851, N14);
buf BUFF1_1152 (N11854, N1446);
buf BUFF1_1153 (N11857, N1457);
buf BUFF1_1154 (N11860, N1468);
buf BUFF1_1155 (N11863, N1435);
buf BUFF1_1156 (N11866, N1389);
buf BUFF1_1157 (N11869, N1400);
buf BUFF1_1158 (N11872, N1411);
buf BUFF1_1159 (N11875, N1422);
buf BUFF1_1160 (N11878, N1374);
buf BUFF1_1161 (N11881, N1479);
buf BUFF1_1162 (N11884, N1490);
buf BUFF1_1163 (N11887, N1503);
buf BUFF1_1164 (N11890, N1514);
buf BUFF1_1165 (N11893, N1523);
buf BUFF1_1166 (N11896, N1534);
buf BUFF1_1167 (N11899, N154);
buf BUFF1_1168 (N11902, N1479);
buf BUFF1_1169 (N11905, N1503);
buf BUFF1_1170 (N11908, N1514);
buf BUFF1_1171 (N11911, N1523);
buf BUFF1_1172 (N11914, N1534);
buf BUFF1_1173 (N11917, N1490);
buf BUFF1_1174 (N11920, N1361);
buf BUFF1_1175 (N11923, N1369);
buf BUFF1_1176 (N11926, N1341);
buf BUFF1_1177 (N11929, N1351);
buf BUFF1_1178 (N11932, N1308);
buf BUFF1_1179 (N11935, N1316);
buf BUFF1_1180 (N11938, N1293);
buf BUFF1_1181 (N11941, N1302);
buf BUFF1_1182 (N11944, N1281);
buf BUFF1_1183 (N11947, N1289);
buf BUFF1_1184 (N11950, N1265);
buf BUFF1_1185 (N11953, N1273);
buf BUFF1_1186 (N11956, N1234);
buf BUFF1_1187 (N11959, N1257);
buf BUFF1_1188 (N11962, N1218);
buf BUFF1_1189 (N11965, N1226);
buf BUFF1_1190 (N11968, N1210);
not NOT1_1191 (N11972, N11146);
and AND2_1192 (N12054, N1136, N11148);
not NOT1_1193 (N12060, N11150);
not NOT1_1194 (N12061, N11151);
buf BUFF1_1195 (N12139, N11209);
buf BUFF1_1196 (N12142, N11216);
buf BUFF1_1197 (N12309, N11479);
and AND2_1198 (N12349, N11104, N1514);
or OR2_1199 (N12350, N11067, N1514);
buf BUFF1_1200 (N12387, N11580);
buf BUFF1_1201 (N12527, N11821);
not NOT1_1202 (N12584, N11580);
and AND3_1203 (N12585, N1170, N11161, N11173);
and AND3_1204 (N12586, N1173, N11161, N11173);
and AND3_1205 (N12587, N1167, N11161, N11173);
and AND3_1206 (N12588, N1164, N11161, N11173);
and AND3_1207 (N12589, N1161, N11161, N11173);
nand NAND2_1208 (N12590, N11475, N1140);
and AND3_1209 (N12591, N1185, N11185, N11197);
and AND3_1210 (N12592, N1158, N11185, N11197);
and AND3_1211 (N12593, N1152, N11185, N11197);
and AND3_1212 (N12594, N1146, N11185, N11197);
and AND3_1213 (N12595, N1170, N11223, N11235);
and AND3_1214 (N12596, N1173, N11223, N11235);
and AND3_1215 (N12597, N1167, N11223, N11235);
and AND3_1216 (N12598, N1164, N11223, N11235);
and AND3_1217 (N12599, N1161, N11223, N11235);
and AND3_1218 (N12600, N1185, N11247, N11259);
and AND3_1219 (N12601, N1158, N11247, N11259);
and AND3_1220 (N12602, N1152, N11247, N11259);
and AND3_1221 (N12603, N1146, N11247, N11259);
and AND3_1222 (N12604, N1106, N11731, N11743);
and AND3_1223 (N12605, N161, N11327, N11339);
and AND3_1224 (N12606, N1106, N11697, N11709);
and AND3_1225 (N12607, N149, N11697, N11709);
and AND3_1226 (N12608, N1103, N11697, N11709);
and AND3_1227 (N12609, N140, N11697, N11709);
and AND3_1228 (N12610, N137, N11697, N11709);
and AND3_1229 (N12611, N120, N11327, N11339);
and AND3_1230 (N12612, N117, N11327, N11339);
and AND3_1231 (N12613, N170, N11327, N11339);
and AND3_1232 (N12614, N164, N11327, N11339);
and AND3_1233 (N12615, N149, N11731, N11743);
and AND3_1234 (N12616, N1103, N11731, N11743);
and AND3_1235 (N12617, N140, N11731, N11743);
and AND3_1236 (N12618, N137, N11731, N11743);
and AND3_1237 (N12619, N120, N11351, N11363);
and AND3_1238 (N12620, N117, N11351, N11363);
and AND3_1239 (N12621, N170, N11351, N11363);
and AND3_1240 (N12622, N164, N11351, N11363);
not NOT1_1241 (N12623, N11475);
and AND3_1242 (N12624, N1123, N11758, N1599);
and AND2_1243 (N12625, N11777, N11785);
and AND3_1244 (N12626, N161, N11351, N11363);
and AND2_1245 (N12627, N11761, N11769);
not NOT1_1246 (N12628, N11824);
not NOT1_1247 (N12629, N11827);
not NOT1_1248 (N12630, N11830);
not NOT1_1249 (N12631, N11833);
not NOT1_1250 (N12632, N11836);
not NOT1_1251 (N12633, N11839);
not NOT1_1252 (N12634, N11842);
not NOT1_1253 (N12635, N11845);
not NOT1_1254 (N12636, N11848);
not NOT1_1255 (N12637, N11851);
not NOT1_1256 (N12638, N11854);
not NOT1_1257 (N12639, N11857);
not NOT1_1258 (N12640, N11860);
not NOT1_1259 (N12641, N11863);
not NOT1_1260 (N12642, N11866);
not NOT1_1261 (N12643, N11869);
not NOT1_1262 (N12644, N11872);
not NOT1_1263 (N12645, N11875);
not NOT1_1264 (N12646, N11878);
buf BUFF1_1265 (N12647, N11209);
not NOT1_1266 (N12653, N11161);
not NOT1_1267 (N12664, N11173);
buf BUFF1_1268 (N12675, N11209);
not NOT1_1269 (N12681, N11185);
not NOT1_1270 (N12692, N11197);
and AND3_1271 (N12703, N1179, N11185, N11197);
buf BUFF1_1272 (N12704, N11479);
not NOT1_1273 (N12709, N11881);
not NOT1_1274 (N12710, N11884);
not NOT1_1275 (N12711, N11887);
not NOT1_1276 (N12712, N11890);
not NOT1_1277 (N12713, N11893);
not NOT1_1278 (N12714, N11896);
not NOT1_1279 (N12715, N11899);
not NOT1_1280 (N12716, N11902);
not NOT1_1281 (N12717, N11905);
not NOT1_1282 (N12718, N11908);
not NOT1_1283 (N12719, N11911);
not NOT1_1284 (N12720, N11914);
not NOT1_1285 (N12721, N11917);
buf BUFF1_1286 (N12722, N11213);
not NOT1_1287 (N12728, N11223);
not NOT1_1288 (N12739, N11235);
buf BUFF1_1289 (N12750, N11213);
not NOT1_1290 (N12756, N11247);
not NOT1_1291 (N12767, N11259);
and AND3_1292 (N12778, N1179, N11247, N11259);
not NOT1_1293 (N12779, N11327);
not NOT1_1294 (N12790, N11339);
not NOT1_1295 (N12801, N11351);
not NOT1_1296 (N12812, N11363);
not NOT1_1297 (N12823, N11375);
not NOT1_1298 (N12824, N11378);
not NOT1_1299 (N12825, N11381);
not NOT1_1300 (N12826, N11384);
not NOT1_1301 (N12827, N11387);
not NOT1_1302 (N12828, N11390);
not NOT1_1303 (N12829, N11393);
not NOT1_1304 (N12830, N11396);
and AND3_1305 (N12831, N11104, N1457, N11378);
and AND3_1306 (N12832, N11104, N1468, N11384);
and AND3_1307 (N12833, N11104, N1422, N11390);
and AND3_1308 (N12834, N11104, N1435, N11396);
and AND2_1309 (N12835, N11067, N11375);
and AND2_1310 (N12836, N11067, N11381);
and AND2_1311 (N12837, N11067, N11387);
and AND2_1312 (N12838, N11067, N11393);
not NOT1_1313 (N12839, N11415);
not NOT1_1314 (N12840, N11418);
not NOT1_1315 (N12841, N11421);
not NOT1_1316 (N12842, N11424);
not NOT1_1317 (N12843, N11427);
not NOT1_1318 (N12844, N11430);
not NOT1_1319 (N12845, N11433);
not NOT1_1320 (N12846, N11436);
and AND3_1321 (N12847, N11104, N1389, N11418);
and AND3_1322 (N12848, N11104, N1400, N11424);
and AND3_1323 (N12849, N11104, N1411, N11430);
and AND3_1324 (N12850, N11104, N1374, N11436);
and AND2_1325 (N12851, N11067, N11415);
and AND2_1326 (N12852, N11067, N11421);
and AND2_1327 (N12853, N11067, N11427);
and AND2_1328 (N12854, N11067, N11433);
not NOT1_1329 (N12855, N11455);
not NOT1_1330 (N12861, N11462);
and AND2_1331 (N12867, N1292, N11455);
and AND2_1332 (N12868, N1288, N11455);
and AND2_1333 (N12869, N1280, N11455);
and AND2_1334 (N12870, N1272, N11455);
and AND2_1335 (N12871, N1264, N11455);
and AND2_1336 (N12872, N1241, N11462);
and AND2_1337 (N12873, N1233, N11462);
and AND2_1338 (N12874, N1225, N11462);
and AND2_1339 (N12875, N1217, N11462);
and AND2_1340 (N12876, N1209, N11462);
buf BUFF1_1341 (N12877, N11216);
not NOT1_1342 (N12882, N11482);
not NOT1_1343 (N12891, N11475);
not NOT1_1344 (N12901, N11492);
not NOT1_1345 (N12902, N11495);
not NOT1_1346 (N12903, N11498);
not NOT1_1347 (N12904, N11501);
not NOT1_1348 (N12905, N11504);
not NOT1_1349 (N12906, N11507);
and AND2_1350 (N12907, N11303, N11495);
and AND3_1351 (N12908, N11303, N1479, N11501);
and AND3_1352 (N12909, N11303, N1490, N11507);
and AND2_1353 (N12910, N11663, N11492);
and AND2_1354 (N12911, N11663, N11498);
and AND2_1355 (N12912, N11663, N11504);
not NOT1_1356 (N12913, N11510);
not NOT1_1357 (N12914, N11513);
not NOT1_1358 (N12915, N11516);
not NOT1_1359 (N12916, N11519);
not NOT1_1360 (N12917, N11522);
not NOT1_1361 (N12918, N11525);
and AND3_1362 (N12919, N11104, N1503, N11513);
not NOT1_1363 (N12920, N12349);
and AND3_1364 (N12921, N11104, N1523, N11519);
and AND3_1365 (N12922, N11104, N1534, N11525);
and AND2_1366 (N12923, N11067, N11510);
and AND2_1367 (N12924, N11067, N11516);
and AND2_1368 (N12925, N11067, N11522);
not NOT1_1369 (N12926, N11542);
not NOT1_1370 (N12927, N11545);
not NOT1_1371 (N12928, N11548);
not NOT1_1372 (N12929, N11551);
not NOT1_1373 (N12930, N11554);
not NOT1_1374 (N12931, N11557);
not NOT1_1375 (N12932, N11560);
not NOT1_1376 (N12933, N11563);
and AND3_1377 (N12934, N11303, N1389, N11545);
and AND3_1378 (N12935, N11303, N1400, N11551);
and AND3_1379 (N12936, N11303, N1411, N11557);
and AND3_1380 (N12937, N11303, N1374, N11563);
and AND2_1381 (N12938, N11663, N11542);
and AND2_1382 (N12939, N11663, N11548);
and AND2_1383 (N12940, N11663, N11554);
and AND2_1384 (N12941, N11663, N11560);
not NOT1_1385 (N12942, N11566);
not NOT1_1386 (N12948, N11573);
and AND2_1387 (N12954, N1372, N11566);
and AND2_1388 (N12955, N1366, N11566);
and AND2_1389 (N12956, N1358, N11566);
and AND2_1390 (N12957, N1348, N11566);
and AND2_1391 (N12958, N1338, N11566);
and AND2_1392 (N12959, N1331, N11573);
and AND2_1393 (N12960, N1323, N11573);
and AND2_1394 (N12961, N1315, N11573);
and AND2_1395 (N12962, N1307, N11573);
and AND2_1396 (N12963, N1299, N11573);
not NOT1_1397 (N12964, N11588);
and AND2_1398 (N12969, N183, N11588);
and AND2_1399 (N12970, N186, N11588);
and AND2_1400 (N12971, N188, N11588);
and AND2_1401 (N12972, N188, N11588);
not NOT1_1402 (N12973, N11594);
not NOT1_1403 (N12974, N11597);
not NOT1_1404 (N12975, N11600);
not NOT1_1405 (N12976, N11603);
not NOT1_1406 (N12977, N11606);
not NOT1_1407 (N12978, N11609);
and AND3_1408 (N12979, N11315, N1503, N11597);
and AND2_1409 (N12980, N11315, N1514);
and AND3_1410 (N12981, N11315, N1523, N11603);
and AND3_1411 (N12982, N11315, N1534, N11609);
and AND2_1412 (N12983, N11675, N11594);
or OR2_1413 (N12984, N11675, N1514);
and AND2_1414 (N12985, N11675, N11600);
and AND2_1415 (N12986, N11675, N11606);
not NOT1_1416 (N12987, N11612);
not NOT1_1417 (N12988, N11615);
not NOT1_1418 (N12989, N11618);
not NOT1_1419 (N12990, N11621);
not NOT1_1420 (N12991, N11624);
not NOT1_1421 (N12992, N11627);
and AND2_1422 (N12993, N11315, N11615);
and AND3_1423 (N12994, N11315, N1479, N11621);
and AND3_1424 (N12995, N11315, N1490, N11627);
and AND2_1425 (N12996, N11675, N11612);
and AND2_1426 (N12997, N11675, N11618);
and AND2_1427 (N12998, N11675, N11624);
not NOT1_1428 (N12999, N11630);
buf BUFF1_1429 (N13000, N11469);
buf BUFF1_1430 (N13003, N11469);
not NOT1_1431 (N13006, N11633);
buf BUFF1_1432 (N13007, N11469);
buf BUFF1_1433 (N13010, N11469);
and AND2_1434 (N13013, N11315, N11630);
and AND2_1435 (N13014, N11315, N11633);
not NOT1_1436 (N13015, N11636);
not NOT1_1437 (N13016, N11639);
not NOT1_1438 (N13017, N11642);
not NOT1_1439 (N13018, N11645);
not NOT1_1440 (N13019, N11648);
not NOT1_1441 (N13020, N11651);
not NOT1_1442 (N13021, N11654);
not NOT1_1443 (N13022, N11657);
and AND3_1444 (N13023, N11303, N1457, N11639);
and AND3_1445 (N13024, N11303, N1468, N11645);
and AND3_1446 (N13025, N11303, N1422, N11651);
and AND3_1447 (N13026, N11303, N1435, N11657);
and AND2_1448 (N13027, N11663, N11636);
and AND2_1449 (N13028, N11663, N11642);
and AND2_1450 (N13029, N11663, N11648);
and AND2_1451 (N13030, N11663, N11654);
not NOT1_1452 (N13031, N11920);
not NOT1_1453 (N13032, N11923);
not NOT1_1454 (N13033, N11926);
not NOT1_1455 (N13034, N11929);
buf BUFF1_1456 (N13035, N11660);
buf BUFF1_1457 (N13038, N11660);
not NOT1_1458 (N13041, N11697);
not NOT1_1459 (N13052, N11709);
not NOT1_1460 (N13063, N11721);
not NOT1_1461 (N13068, N11727);
and AND2_1462 (N13071, N197, N11721);
and AND2_1463 (N13072, N194, N11721);
and AND2_1464 (N13073, N197, N11721);
and AND2_1465 (N13074, N194, N11721);
not NOT1_1466 (N13075, N11731);
not NOT1_1467 (N13086, N11743);
not NOT1_1468 (N13097, N11761);
not NOT1_1469 (N13108, N11769);
not NOT1_1470 (N13119, N11777);
not NOT1_1471 (N13130, N11785);
not NOT1_1472 (N13141, N11944);
not NOT1_1473 (N13142, N11947);
not NOT1_1474 (N13143, N11950);
not NOT1_1475 (N13144, N11953);
not NOT1_1476 (N13145, N11956);
not NOT1_1477 (N13146, N11959);
not NOT1_1478 (N13147, N11793);
not NOT1_1479 (N13158, N11800);
not NOT1_1480 (N13169, N11807);
not NOT1_1481 (N13180, N11814);
buf BUFF1_1482 (N13191, N11821);
not NOT1_1483 (N13194, N11932);
not NOT1_1484 (N13195, N11935);
not NOT1_1485 (N13196, N11938);
not NOT1_1486 (N13197, N11941);
not NOT1_1487 (N13198, N11962);
not NOT1_1488 (N13199, N11965);
buf BUFF1_1489 (N13200, N11469);
not NOT1_1490 (N13203, N11968);
buf BUFF1_1491 (N13357, N12704);
buf BUFF1_1492 (N13358, N12704);
buf BUFF1_1493 (N13359, N12704);
buf BUFF1_1494 (N13360, N12704);
and AND3_1495 (N13401, N1457, N11092, N12824);
and AND3_1496 (N13402, N1468, N11092, N12826);
and AND3_1497 (N13403, N1422, N11092, N12828);
and AND3_1498 (N13404, N1435, N11092, N12830);
and AND2_1499 (N13405, N11080, N12823);
and AND2_1500 (N13406, N11080, N12825);
and AND2_1501 (N13407, N11080, N12827);
and AND2_1502 (N13408, N11080, N12829);
and AND3_1503 (N13409, N1389, N11092, N12840);
and AND3_1504 (N13410, N1400, N11092, N12842);
and AND3_1505 (N13411, N1411, N11092, N12844);
and AND3_1506 (N13412, N1374, N11092, N12846);
and AND2_1507 (N13413, N11080, N12839);
and AND2_1508 (N13414, N11080, N12841);
and AND2_1509 (N13415, N11080, N12843);
and AND2_1510 (N13416, N11080, N12845);
and AND2_1511 (N13444, N11280, N12902);
and AND3_1512 (N13445, N1479, N11280, N12904);
and AND3_1513 (N13446, N1490, N11280, N12906);
and AND2_1514 (N13447, N11685, N12901);
and AND2_1515 (N13448, N11685, N12903);
and AND2_1516 (N13449, N11685, N12905);
and AND3_1517 (N13450, N1503, N11092, N12914);
and AND3_1518 (N13451, N1523, N11092, N12916);
and AND3_1519 (N13452, N1534, N11092, N12918);
and AND2_1520 (N13453, N11080, N12913);
and AND2_1521 (N13454, N11080, N12915);
and AND2_1522 (N13455, N11080, N12917);
and AND2_1523 (N13456, N12920, N12350);
and AND3_1524 (N13459, N1389, N11280, N12927);
and AND3_1525 (N13460, N1400, N11280, N12929);
and AND3_1526 (N13461, N1411, N11280, N12931);
and AND3_1527 (N13462, N1374, N11280, N12933);
and AND2_1528 (N13463, N11685, N12926);
and AND2_1529 (N13464, N11685, N12928);
and AND2_1530 (N13465, N11685, N12930);
and AND2_1531 (N13466, N11685, N12932);
and AND3_1532 (N13481, N1503, N11292, N12974);
not NOT1_1533 (N13482, N12980);
and AND3_1534 (N13483, N1523, N11292, N12976);
and AND3_1535 (N13484, N1534, N11292, N12978);
and AND2_1536 (N13485, N11271, N12973);
and AND2_1537 (N13486, N11271, N12975);
and AND2_1538 (N13487, N11271, N12977);
and AND2_1539 (N13488, N11292, N12988);
and AND3_1540 (N13489, N1479, N11292, N12990);
and AND3_1541 (N13490, N1490, N11292, N12992);
and AND2_1542 (N13491, N11271, N12987);
and AND2_1543 (N13492, N11271, N12989);
and AND2_1544 (N13493, N11271, N12991);
and AND2_1545 (N13502, N11292, N12999);
and AND2_1546 (N13503, N11292, N13006);
and AND3_1547 (N13504, N1457, N11280, N13016);
and AND3_1548 (N13505, N1468, N11280, N13018);
and AND3_1549 (N13506, N1422, N11280, N13020);
and AND3_1550 (N13507, N1435, N11280, N13022);
and AND2_1551 (N13508, N11685, N13015);
and AND2_1552 (N13509, N11685, N13017);
and AND2_1553 (N13510, N11685, N13019);
and AND2_1554 (N13511, N11685, N13021);
nand NAND2_1555 (N13512, N11923, N13031);
nand NAND2_1556 (N13513, N11920, N13032);
nand NAND2_1557 (N13514, N11929, N13033);
nand NAND2_1558 (N13515, N11926, N13034);
nand NAND2_1559 (N13558, N11947, N13141);
nand NAND2_1560 (N13559, N11944, N13142);
nand NAND2_1561 (N13560, N11953, N13143);
nand NAND2_1562 (N13561, N11950, N13144);
nand NAND2_1563 (N13562, N11959, N13145);
nand NAND2_1564 (N13563, N11956, N13146);
buf BUFF1_1565 (N13604, N13191);
nand NAND2_1566 (N13605, N11935, N13194);
nand NAND2_1567 (N13606, N11932, N13195);
nand NAND2_1568 (N13607, N11941, N13196);
nand NAND2_1569 (N13608, N11938, N13197);
nand NAND2_1570 (N13609, N11965, N13198);
nand NAND2_1571 (N13610, N11962, N13199);
not NOT1_1572 (N13613, N13191);
and AND2_1573 (N13614, N12882, N12891);
and AND2_1574 (N13615, N11482, N12891);
and AND3_1575 (N13616, N1200, N12653, N11173);
and AND3_1576 (N13617, N1203, N12653, N11173);
and AND3_1577 (N13618, N1197, N12653, N11173);
and AND3_1578 (N13619, N1194, N12653, N11173);
and AND3_1579 (N13620, N1191, N12653, N11173);
and AND3_1580 (N13621, N1182, N12681, N11197);
and AND3_1581 (N13622, N1188, N12681, N11197);
and AND3_1582 (N13623, N1155, N12681, N11197);
and AND3_1583 (N13624, N1149, N12681, N11197);
and AND2_1584 (N13625, N12882, N12891);
and AND2_1585 (N13626, N11482, N12891);
and AND3_1586 (N13627, N1200, N12728, N11235);
and AND3_1587 (N13628, N1203, N12728, N11235);
and AND3_1588 (N13629, N1197, N12728, N11235);
and AND3_1589 (N13630, N1194, N12728, N11235);
and AND3_1590 (N13631, N1191, N12728, N11235);
and AND3_1591 (N13632, N1182, N12756, N11259);
and AND3_1592 (N13633, N1188, N12756, N11259);
and AND3_1593 (N13634, N1155, N12756, N11259);
and AND3_1594 (N13635, N1149, N12756, N11259);
and AND2_1595 (N13636, N12882, N12891);
and AND2_1596 (N13637, N11482, N12891);
and AND3_1597 (N13638, N1109, N13075, N11743);
and AND2_1598 (N13639, N12882, N12891);
and AND2_1599 (N13640, N11482, N12891);
and AND3_1600 (N13641, N111, N12779, N11339);
and AND3_1601 (N13642, N1109, N13041, N11709);
and AND3_1602 (N13643, N146, N13041, N11709);
and AND3_1603 (N13644, N1100, N13041, N11709);
and AND3_1604 (N13645, N191, N13041, N11709);
and AND3_1605 (N13646, N143, N13041, N11709);
and AND3_1606 (N13647, N176, N12779, N11339);
and AND3_1607 (N13648, N173, N12779, N11339);
and AND3_1608 (N13649, N167, N12779, N11339);
and AND3_1609 (N13650, N114, N12779, N11339);
and AND3_1610 (N13651, N146, N13075, N11743);
and AND3_1611 (N13652, N1100, N13075, N11743);
and AND3_1612 (N13653, N191, N13075, N11743);
and AND3_1613 (N13654, N143, N13075, N11743);
and AND3_1614 (N13655, N176, N12801, N11363);
and AND3_1615 (N13656, N173, N12801, N11363);
and AND3_1616 (N13657, N167, N12801, N11363);
and AND3_1617 (N13658, N114, N12801, N11363);
and AND3_1618 (N13659, N1120, N13119, N11785);
and AND3_1619 (N13660, N111, N12801, N11363);
and AND3_1620 (N13661, N1118, N13097, N11769);
and AND3_1621 (N13662, N1176, N12681, N11197);
and AND3_1622 (N13663, N1176, N12756, N11259);
or OR2_1623 (N13664, N12831, N13401);
or OR2_1624 (N13665, N12832, N13402);
or OR2_1625 (N13666, N12833, N13403);
or OR2_1626 (N13667, N12834, N13404);
or OR3_1627 (N13668, N12835, N13405, N1457);
or OR3_1628 (N13669, N12836, N13406, N1468);
or OR3_1629 (N13670, N12837, N13407, N1422);
or OR3_1630 (N13671, N12838, N13408, N1435);
or OR2_1631 (N13672, N12847, N13409);
or OR2_1632 (N13673, N12848, N13410);
or OR2_1633 (N13674, N12849, N13411);
or OR2_1634 (N13675, N12850, N13412);
or OR3_1635 (N13676, N12851, N13413, N1389);
or OR3_1636 (N13677, N12852, N13414, N1400);
or OR3_1637 (N13678, N12853, N13415, N1411);
or OR3_1638 (N13679, N12854, N13416, N1374);
and AND2_1639 (N13680, N1289, N12855);
and AND2_1640 (N13681, N1281, N12855);
and AND2_1641 (N13682, N1273, N12855);
and AND2_1642 (N13683, N1265, N12855);
and AND2_1643 (N13684, N1257, N12855);
and AND2_1644 (N13685, N1234, N12861);
and AND2_1645 (N13686, N1226, N12861);
and AND2_1646 (N13687, N1218, N12861);
and AND2_1647 (N13688, N1210, N12861);
and AND2_1648 (N13689, N1206, N12861);
not NOT1_1649 (N13691, N12891);
or OR2_1650 (N13700, N12907, N13444);
or OR2_1651 (N13701, N12908, N13445);
or OR2_1652 (N13702, N12909, N13446);
or OR3_1653 (N13703, N12911, N13448, N1479);
or OR3_1654 (N13704, N12912, N13449, N1490);
or OR2_1655 (N13705, N12910, N13447);
or OR2_1656 (N13708, N12919, N13450);
or OR2_1657 (N13709, N12921, N13451);
or OR2_1658 (N13710, N12922, N13452);
or OR3_1659 (N13711, N12923, N13453, N1503);
or OR3_1660 (N13712, N12924, N13454, N1523);
or OR3_1661 (N13713, N12925, N13455, N1534);
or OR2_1662 (N13715, N12934, N13459);
or OR2_1663 (N13716, N12935, N13460);
or OR2_1664 (N13717, N12936, N13461);
or OR2_1665 (N13718, N12937, N13462);
or OR3_1666 (N13719, N12938, N13463, N1389);
or OR3_1667 (N13720, N12939, N13464, N1400);
or OR3_1668 (N13721, N12940, N13465, N1411);
or OR3_1669 (N13722, N12941, N13466, N1374);
and AND2_1670 (N13723, N1369, N12942);
and AND2_1671 (N13724, N1361, N12942);
and AND2_1672 (N13725, N1351, N12942);
and AND2_1673 (N13726, N1341, N12942);
and AND2_1674 (N13727, N1324, N12948);
and AND2_1675 (N13728, N1316, N12948);
and AND2_1676 (N13729, N1308, N12948);
and AND2_1677 (N13730, N1302, N12948);
and AND2_1678 (N13731, N1293, N12948);
or OR2_1679 (N13732, N12942, N12958);
and AND2_1680 (N13738, N183, N12964);
and AND2_1681 (N13739, N187, N12964);
and AND2_1682 (N13740, N134, N12964);
and AND2_1683 (N13741, N134, N12964);
or OR2_1684 (N13742, N12979, N13481);
or OR2_1685 (N13743, N12981, N13483);
or OR2_1686 (N13744, N12982, N13484);
or OR3_1687 (N13745, N12983, N13485, N1503);
or OR3_1688 (N13746, N12985, N13486, N1523);
or OR3_1689 (N13747, N12986, N13487, N1534);
or OR2_1690 (N13748, N12993, N13488);
or OR2_1691 (N13749, N12994, N13489);
or OR2_1692 (N13750, N12995, N13490);
or OR3_1693 (N13751, N12997, N13492, N1479);
or OR3_1694 (N13752, N12998, N13493, N1490);
not NOT1_1695 (N13753, N13000);
not NOT1_1696 (N13754, N13003);
not NOT1_1697 (N13755, N13007);
not NOT1_1698 (N13756, N13010);
or OR2_1699 (N13757, N13013, N13502);
and AND3_1700 (N13758, N11315, N1446, N13003);
or OR2_1701 (N13759, N13014, N13503);
and AND3_1702 (N13760, N11315, N1446, N13010);
and AND2_1703 (N13761, N11675, N13000);
and AND2_1704 (N13762, N11675, N13007);
or OR2_1705 (N13763, N13023, N13504);
or OR2_1706 (N13764, N13024, N13505);
or OR2_1707 (N13765, N13025, N13506);
or OR2_1708 (N13766, N13026, N13507);
or OR3_1709 (N13767, N13027, N13508, N1457);
or OR3_1710 (N13768, N13028, N13509, N1468);
or OR3_1711 (N13769, N13029, N13510, N1422);
or OR3_1712 (N13770, N13030, N13511, N1435);
nand NAND2_1713 (N13771, N13512, N13513);
nand NAND2_1714 (N13775, N13514, N13515);
not NOT1_1715 (N13779, N13035);
not NOT1_1716 (N13780, N13038);
and AND3_1717 (N13781, N1117, N13097, N11769);
and AND3_1718 (N13782, N1126, N13097, N11769);
and AND3_1719 (N13783, N1127, N13097, N11769);
and AND3_1720 (N13784, N1128, N13097, N11769);
and AND3_1721 (N13785, N1131, N13119, N11785);
and AND3_1722 (N13786, N1129, N13119, N11785);
and AND3_1723 (N13787, N1119, N13119, N11785);
and AND3_1724 (N13788, N1130, N13119, N11785);
nand NAND2_1725 (N13789, N13558, N13559);
nand NAND2_1726 (N13793, N13560, N13561);
nand NAND2_1727 (N13797, N13562, N13563);
and AND3_1728 (N13800, N1122, N13147, N11800);
and AND3_1729 (N13801, N1113, N13147, N11800);
and AND3_1730 (N13802, N153, N13147, N11800);
and AND3_1731 (N13803, N1114, N13147, N11800);
and AND3_1732 (N13804, N1115, N13147, N11800);
and AND3_1733 (N13805, N152, N13169, N11814);
and AND3_1734 (N13806, N1112, N13169, N11814);
and AND3_1735 (N13807, N1116, N13169, N11814);
and AND3_1736 (N13808, N1121, N13169, N11814);
and AND3_1737 (N13809, N1123, N13169, N11814);
nand NAND2_1738 (N13810, N13607, N13608);
nand NAND2_1739 (N13813, N13605, N13606);
and AND2_1740 (N13816, N13482, N12984);
or OR2_1741 (N13819, N12996, N13491);
not NOT1_1742 (N13822, N13200);
nand NAND2_1743 (N13823, N13200, N13203);
nand NAND2_1744 (N13824, N13609, N13610);
not NOT1_1745 (N13827, N13456);
or OR2_1746 (N13828, N13739, N12970);
or OR2_1747 (N13829, N13740, N12971);
or OR2_1748 (N13830, N13741, N12972);
or OR2_1749 (N13831, N13738, N12969);
not NOT1_1750 (N13834, N13664);
not NOT1_1751 (N13835, N13665);
not NOT1_1752 (N13836, N13666);
not NOT1_1753 (N13837, N13667);
not NOT1_1754 (N13838, N13672);
not NOT1_1755 (N13839, N13673);
not NOT1_1756 (N13840, N13674);
not NOT1_1757 (N13841, N13675);
or OR2_1758 (N13842, N13681, N12868);
or OR2_1759 (N13849, N13682, N12869);
or OR2_1760 (N13855, N13683, N12870);
or OR2_1761 (N13861, N13684, N12871);
or OR2_1762 (N13867, N13685, N12872);
or OR2_1763 (N13873, N13686, N12873);
or OR2_1764 (N13881, N13687, N12874);
or OR2_1765 (N13887, N13688, N12875);
or OR2_1766 (N13893, N13689, N12876);
not NOT1_1767 (N13908, N13701);
not NOT1_1768 (N13909, N13702);
not NOT1_1769 (N13911, N13700);
not NOT1_1770 (N13914, N13708);
not NOT1_1771 (N13915, N13709);
not NOT1_1772 (N13916, N13710);
not NOT1_1773 (N13917, N13715);
not NOT1_1774 (N13918, N13716);
not NOT1_1775 (N13919, N13717);
not NOT1_1776 (N13920, N13718);
or OR2_1777 (N13921, N13724, N12955);
or OR2_1778 (N13927, N13725, N12956);
or OR2_1779 (N13933, N13726, N12957);
or OR2_1780 (N13942, N13727, N12959);
or OR2_1781 (N13948, N13728, N12960);
or OR2_1782 (N13956, N13729, N12961);
or OR2_1783 (N13962, N13730, N12962);
or OR2_1784 (N13968, N13731, N12963);
not NOT1_1785 (N13975, N13742);
not NOT1_1786 (N13976, N13743);
not NOT1_1787 (N13977, N13744);
not NOT1_1788 (N13978, N13749);
not NOT1_1789 (N13979, N13750);
and AND3_1790 (N13980, N1446, N11292, N13754);
and AND3_1791 (N13981, N1446, N11292, N13756);
and AND2_1792 (N13982, N11271, N13753);
and AND2_1793 (N13983, N11271, N13755);
not NOT1_1794 (N13984, N13757);
not NOT1_1795 (N13987, N13759);
not NOT1_1796 (N13988, N13763);
not NOT1_1797 (N13989, N13764);
not NOT1_1798 (N13990, N13765);
not NOT1_1799 (N13991, N13766);
and AND3_1800 (N13998, N13456, N13119, N13130);
or OR2_1801 (N14008, N13723, N12954);
or OR2_1802 (N14011, N13680, N12867);
not NOT1_1803 (N14021, N13748);
nand NAND2_1804 (N14024, N11968, N13822);
not NOT1_1805 (N14027, N13705);
and AND2_1806 (N14031, N13828, N11583);
and AND3_1807 (N14032, N124, N12882, N13691);
and AND3_1808 (N14033, N125, N11482, N13691);
and AND3_1809 (N14034, N126, N12882, N13691);
and AND3_1810 (N14035, N181, N11482, N13691);
and AND2_1811 (N14036, N13829, N11583);
and AND3_1812 (N14037, N179, N12882, N13691);
and AND3_1813 (N14038, N123, N11482, N13691);
and AND3_1814 (N14039, N182, N12882, N13691);
and AND3_1815 (N14040, N180, N11482, N13691);
and AND2_1816 (N14041, N13830, N11583);
and AND2_1817 (N14042, N13831, N11583);
and AND2_1818 (N14067, N13732, N1514);
and AND2_1819 (N14080, N1514, N13732);
and AND2_1820 (N14088, N13834, N13668);
and AND2_1821 (N14091, N13835, N13669);
and AND2_1822 (N14094, N13836, N13670);
and AND2_1823 (N14097, N13837, N13671);
and AND2_1824 (N14100, N13838, N13676);
and AND2_1825 (N14103, N13839, N13677);
and AND2_1826 (N14106, N13840, N13678);
and AND2_1827 (N14109, N13841, N13679);
and AND2_1828 (N14144, N13908, N13703);
and AND2_1829 (N14147, N13909, N13704);
buf BUFF1_1830 (N14150, N13705);
and AND2_1831 (N14153, N13914, N13711);
and AND2_1832 (N14156, N13915, N13712);
and AND2_1833 (N14159, N13916, N13713);
or OR2_1834 (N14183, N13758, N13980);
or OR2_1835 (N14184, N13760, N13981);
or OR3_1836 (N14185, N13761, N13982, N1446);
or OR3_1837 (N14186, N13762, N13983, N1446);
not NOT1_1838 (N14188, N13771);
not NOT1_1839 (N14191, N13775);
and AND3_1840 (N14196, N13775, N13771, N13035);
and AND3_1841 (N14197, N13987, N13119, N13130);
and AND2_1842 (N14198, N13920, N13722);
not NOT1_1843 (N14199, N13816);
not NOT1_1844 (N14200, N13789);
not NOT1_1845 (N14203, N13793);
buf BUFF1_1846 (N14206, N13797);
buf BUFF1_1847 (N14209, N13797);
buf BUFF1_1848 (N14212, N13732);
buf BUFF1_1849 (N14215, N13732);
buf BUFF1_1850 (N14219, N13732);
not NOT1_1851 (N14223, N13810);
not NOT1_1852 (N14224, N13813);
and AND2_1853 (N14225, N13918, N13720);
and AND2_1854 (N14228, N13919, N13721);
and AND2_1855 (N14231, N13991, N13770);
and AND2_1856 (N14234, N13917, N13719);
and AND2_1857 (N14237, N13989, N13768);
and AND2_1858 (N14240, N13990, N13769);
and AND2_1859 (N14243, N13988, N13767);
and AND2_1860 (N14246, N13976, N13746);
and AND2_1861 (N14249, N13977, N13747);
and AND2_1862 (N14252, N13975, N13745);
and AND2_1863 (N14255, N13978, N13751);
and AND2_1864 (N14258, N13979, N13752);
not NOT1_1865 (N14263, N13819);
nand NAND2_1866 (N14264, N14024, N13823);
not NOT1_1867 (N14267, N13824);
and AND2_1868 (N14268, N1446, N13893);
not NOT1_1869 (N14269, N13911);
not NOT1_1870 (N14270, N13984);
and AND2_1871 (N14271, N13893, N1446);
not NOT1_1872 (N14272, N14031);
or OR4_1873 (N14273, N14032, N14033, N13614, N13615);
or OR4_1874 (N14274, N14034, N14035, N13625, N13626);
not NOT1_1875 (N14275, N14036);
or OR4_1876 (N14276, N14037, N14038, N13636, N13637);
or OR4_1877 (N14277, N14039, N14040, N13639, N13640);
not NOT1_1878 (N14278, N14041);
not NOT1_1879 (N14279, N14042);
and AND2_1880 (N14280, N13887, N1457);
and AND2_1881 (N14284, N13881, N1468);
and AND2_1882 (N14290, N1422, N13873);
and AND2_1883 (N14297, N13867, N1435);
and AND2_1884 (N14298, N13861, N1389);
and AND2_1885 (N14301, N13855, N1400);
and AND2_1886 (N14305, N13849, N1411);
and AND2_1887 (N14310, N13842, N1374);
and AND2_1888 (N14316, N1457, N13887);
and AND2_1889 (N14320, N1468, N13881);
and AND2_1890 (N14325, N1422, N13873);
and AND2_1891 (N14331, N1435, N13867);
and AND2_1892 (N14332, N1389, N13861);
and AND2_1893 (N14336, N1400, N13855);
and AND2_1894 (N14342, N1411, N13849);
and AND2_1895 (N14349, N1374, N13842);
not NOT1_1896 (N14357, N13968);
not NOT1_1897 (N14364, N13962);
buf BUFF1_1898 (N14375, N13962);
and AND2_1899 (N14379, N13956, N1479);
and AND2_1900 (N14385, N1490, N13948);
and AND2_1901 (N14392, N13942, N1503);
and AND2_1902 (N14396, N13933, N1523);
and AND2_1903 (N14400, N13927, N1534);
not NOT1_1904 (N14405, N13921);
buf BUFF1_1905 (N14412, N13921);
not NOT1_1906 (N14418, N13968);
not NOT1_1907 (N14425, N13962);
buf BUFF1_1908 (N14436, N13962);
and AND2_1909 (N14440, N1479, N13956);
and AND2_1910 (N14445, N1490, N13948);
and AND2_1911 (N14451, N1503, N13942);
and AND2_1912 (N14456, N1523, N13933);
and AND2_1913 (N14462, N1534, N13927);
buf BUFF1_1914 (N14469, N13921);
not NOT1_1915 (N14477, N13921);
buf BUFF1_1916 (N14512, N13968);
not NOT1_1917 (N14515, N14183);
not NOT1_1918 (N14516, N14184);
not NOT1_1919 (N14521, N14008);
not NOT1_1920 (N14523, N14011);
not NOT1_1921 (N14524, N14198);
not NOT1_1922 (N14532, N13984);
and AND3_1923 (N14547, N13911, N13169, N13180);
buf BUFF1_1924 (N14548, N13893);
buf BUFF1_1925 (N14551, N13887);
buf BUFF1_1926 (N14554, N13881);
buf BUFF1_1927 (N14557, N13873);
buf BUFF1_1928 (N14560, N13867);
buf BUFF1_1929 (N14563, N13861);
buf BUFF1_1930 (N14566, N13855);
buf BUFF1_1931 (N14569, N13849);
buf BUFF1_1932 (N14572, N13842);
nor N1OR2_1933 (N14575, N1422, N13873);
buf BUFF1_1934 (N14578, N13893);
buf BUFF1_1935 (N14581, N13887);
buf BUFF1_1936 (N14584, N13881);
buf BUFF1_1937 (N14587, N13867);
buf BUFF1_1938 (N14590, N13861);
buf BUFF1_1939 (N14593, N13855);
buf BUFF1_1940 (N14596, N13849);
buf BUFF1_1941 (N14599, N13873);
buf BUFF1_1942 (N14602, N13842);
nor N1OR2_1943 (N14605, N1422, N13873);
nor N1OR2_1944 (N14608, N1374, N13842);
buf BUFF1_1945 (N14611, N13956);
buf BUFF1_1946 (N14614, N13948);
buf BUFF1_1947 (N14617, N13942);
buf BUFF1_1948 (N14621, N13933);
buf BUFF1_1949 (N14624, N13927);
nor N1OR2_1950 (N14627, N1490, N13948);
buf BUFF1_1951 (N14630, N13956);
buf BUFF1_1952 (N14633, N13942);
buf BUFF1_1953 (N14637, N13933);
buf BUFF1_1954 (N14640, N13927);
buf BUFF1_1955 (N14643, N13948);
nor N1OR2_1956 (N14646, N1490, N13948);
buf BUFF1_1957 (N14649, N13927);
buf BUFF1_1958 (N14652, N13933);
buf BUFF1_1959 (N14655, N13921);
buf BUFF1_1960 (N14658, N13942);
buf BUFF1_1961 (N14662, N13956);
buf BUFF1_1962 (N14665, N13948);
buf BUFF1_1963 (N14668, N13968);
buf BUFF1_1964 (N14671, N13962);
buf BUFF1_1965 (N14674, N13873);
buf BUFF1_1966 (N14677, N13867);
buf BUFF1_1967 (N14680, N13887);
buf BUFF1_1968 (N14683, N13881);
buf BUFF1_1969 (N14686, N13893);
buf BUFF1_1970 (N14689, N13849);
buf BUFF1_1971 (N14692, N13842);
buf BUFF1_1972 (N14695, N13861);
buf BUFF1_1973 (N14698, N13855);
nand NAND2_1974 (N14701, N13813, N14223);
nand NAND2_1975 (N14702, N13810, N14224);
not NOT1_1976 (N14720, N14021);
nand NAND2_1977 (N14721, N14021, N14263);
not NOT1_1978 (N14724, N14147);
not NOT1_1979 (N14725, N14144);
not NOT1_1980 (N14726, N14159);
not NOT1_1981 (N14727, N14156);
not NOT1_1982 (N14728, N14153);
not NOT1_1983 (N14729, N14097);
not NOT1_1984 (N14730, N14094);
not NOT1_1985 (N14731, N14091);
not NOT1_1986 (N14732, N14088);
not NOT1_1987 (N14733, N14109);
not NOT1_1988 (N14734, N14106);
not NOT1_1989 (N14735, N14103);
not NOT1_1990 (N14736, N14100);
and AND2_1991 (N14737, N14273, N12877);
and AND2_1992 (N14738, N14274, N12877);
and AND2_1993 (N14739, N14276, N12877);
and AND2_1994 (N14740, N14277, N12877);
and AND3_1995 (N14741, N14150, N11758, N11755);
not NOT1_1996 (N14855, N14212);
nand NAND2_1997 (N14856, N14212, N12712);
nand NAND2_1998 (N14908, N14215, N12718);
not NOT1_1999 (N14909, N14215);
and AND2_11000 (N14939, N14515, N14185);
and AND2_11001 (N14942, N14516, N14186);
not NOT1_11002 (N14947, N14219);
and AND3_11003 (N14953, N14188, N13775, N13779);
and AND3_11004 (N14954, N13771, N14191, N13780);
and AND3_11005 (N14955, N14191, N14188, N13038);
and AND3_11006 (N14956, N14109, N13097, N13108);
and AND3_11007 (N14957, N14106, N13097, N13108);
and AND3_11008 (N14958, N14103, N13097, N13108);
and AND3_11009 (N14959, N14100, N13097, N13108);
and AND3_11010 (N14960, N14159, N13119, N13130);
and AND3_11011 (N14961, N14156, N13119, N13130);
not NOT1_11012 (N14965, N14225);
not NOT1_11013 (N14966, N14228);
not NOT1_11014 (N14967, N14231);
not NOT1_11015 (N14968, N14234);
not NOT1_11016 (N14972, N14246);
not NOT1_11017 (N14973, N14249);
not NOT1_11018 (N14974, N14252);
nand NAND2_11019 (N14975, N14252, N14199);
not NOT1_11020 (N14976, N14206);
not NOT1_11021 (N14977, N14209);
and AND3_11022 (N14978, N13793, N13789, N14206);
and AND3_11023 (N14979, N14203, N14200, N14209);
and AND3_11024 (N14980, N14097, N13147, N13158);
and AND3_11025 (N14981, N14094, N13147, N13158);
and AND3_11026 (N14982, N14091, N13147, N13158);
and AND3_11027 (N14983, N14088, N13147, N13158);
and AND3_11028 (N14984, N14153, N13169, N13180);
and AND3_11029 (N14985, N14147, N13169, N13180);
and AND3_11030 (N14986, N14144, N13169, N13180);
and AND3_11031 (N14987, N14150, N13169, N13180);
nand NAND2_11032 (N15049, N14701, N14702);
not NOT1_11033 (N15052, N14237);
not NOT1_11034 (N15053, N14240);
not NOT1_11035 (N15054, N14243);
not NOT1_11036 (N15055, N14255);
not NOT1_11037 (N15056, N14258);
nand NAND2_11038 (N15057, N13819, N14720);
not NOT1_11039 (N15058, N14264);
nand NAND2_11040 (N15059, N14264, N14267);
and AND4_11041 (N15060, N14724, N14725, N14269, N14027);
and AND4_11042 (N15061, N14726, N14727, N13827, N14728);
and AND4_11043 (N15062, N14729, N14730, N14731, N14732);
and AND4_11044 (N15063, N14733, N14734, N14735, N14736);
and AND2_11045 (N15065, N14357, N14375);
and AND3_11046 (N15066, N14364, N14357, N14379);
and AND2_11047 (N15067, N14418, N14436);
and AND3_11048 (N15068, N14425, N14418, N14440);
not NOT1_11049 (N15069, N14548);
nand NAND2_11050 (N15070, N14548, N12628);
not NOT1_11051 (N15071, N14551);
nand NAND2_11052 (N15072, N14551, N12629);
not NOT1_11053 (N15073, N14554);
nand NAND2_11054 (N15074, N14554, N12630);
not NOT1_11055 (N15075, N14557);
nand NAND2_11056 (N15076, N14557, N12631);
not NOT1_11057 (N15077, N14560);
nand NAND2_11058 (N15078, N14560, N12632);
not NOT1_11059 (N15079, N14563);
nand NAND2_11060 (N15080, N14563, N12633);
not NOT1_11061 (N15081, N14566);
nand NAND2_11062 (N15082, N14566, N12634);
not NOT1_11063 (N15083, N14569);
nand NAND2_11064 (N15084, N14569, N12635);
not NOT1_11065 (N15085, N14572);
nand NAND2_11066 (N15086, N14572, N12636);
not NOT1_11067 (N15087, N14575);
nand NAND2_11068 (N15088, N14578, N12638);
not NOT1_11069 (N15089, N14578);
nand NAND2_11070 (N15090, N14581, N12639);
not NOT1_11071 (N15091, N14581);
nand NAND2_11072 (N15092, N14584, N12640);
not NOT1_11073 (N15093, N14584);
nand NAND2_11074 (N15094, N14587, N12641);
not NOT1_11075 (N15095, N14587);
nand NAND2_11076 (N15096, N14590, N12642);
not NOT1_11077 (N15097, N14590);
nand NAND2_11078 (N15098, N14593, N12643);
not NOT1_11079 (N15099, N14593);
nand NAND2_11080 (N15100, N14596, N12644);
not NOT1_11081 (N15101, N14596);
nand NAND2_11082 (N15102, N14599, N12645);
not NOT1_11083 (N15103, N14599);
nand NAND2_11084 (N15104, N14602, N12646);
not NOT1_11085 (N15105, N14602);
not NOT1_11086 (N15106, N14611);
nand NAND2_11087 (N15107, N14611, N12709);
not NOT1_11088 (N15108, N14614);
nand NAND2_11089 (N15109, N14614, N12710);
not NOT1_11090 (N15110, N14617);
nand NAND2_11091 (N15111, N14617, N12711);
nand NAND2_11092 (N15112, N11890, N14855);
not NOT1_11093 (N15113, N14621);
nand NAND2_11094 (N15114, N14621, N12713);
not NOT1_11095 (N15115, N14624);
nand NAND2_11096 (N15116, N14624, N12714);
and AND2_11097 (N15117, N14364, N14379);
and AND2_11098 (N15118, N14364, N14379);
and AND2_11099 (N15119, N154, N14405);
not NOT1_11100 (N15120, N14627);
nand NAND2_11101 (N15121, N14630, N12716);
not NOT1_11102 (N15122, N14630);
nand NAND2_11103 (N15123, N14633, N12717);
not NOT1_11104 (N15124, N14633);
nand NAND2_11105 (N15125, N11908, N14909);
nand NAND2_11106 (N15126, N14637, N12719);
not NOT1_11107 (N15127, N14637);
nand NAND2_11108 (N15128, N14640, N12720);
not NOT1_11109 (N15129, N14640);
nand NAND2_11110 (N15130, N14643, N12721);
not NOT1_11111 (N15131, N14643);
and AND2_11112 (N15132, N14425, N14440);
and AND2_11113 (N15133, N14425, N14440);
not NOT1_11114 (N15135, N14649);
not NOT1_11115 (N15136, N14652);
nand NAND2_11116 (N15137, N14655, N14521);
not NOT1_11117 (N15138, N14655);
not NOT1_11118 (N15139, N14658);
nand NAND2_11119 (N15140, N14658, N14947);
not NOT1_11120 (N15141, N14674);
not NOT1_11121 (N15142, N14677);
not NOT1_11122 (N15143, N14680);
not NOT1_11123 (N15144, N14683);
nand NAND2_11124 (N15145, N14686, N14523);
not NOT1_11125 (N15146, N14686);
nor N1OR2_11126 (N15147, N14953, N14196);
nor N1OR2_11127 (N15148, N14954, N14955);
not NOT1_11128 (N15150, N14524);
nand NAND2_11129 (N15153, N14228, N14965);
nand NAND2_11130 (N15154, N14225, N14966);
nand NAND2_11131 (N15155, N14234, N14967);
nand NAND2_11132 (N15156, N14231, N14968);
not NOT1_11133 (N15157, N14532);
nand NAND2_11134 (N15160, N14249, N14972);
nand NAND2_11135 (N15161, N14246, N14973);
nand NAND2_11136 (N15162, N13816, N14974);
and AND3_11137 (N15163, N14200, N13793, N14976);
and AND3_11138 (N15164, N13789, N14203, N14977);
and AND3_11139 (N15165, N14942, N13147, N13158);
not NOT1_11140 (N15166, N14512);
buf BUFF1_11141 (N15169, N14290);
not NOT1_11142 (N15172, N14605);
buf BUFF1_11143 (N15173, N14325);
not NOT1_11144 (N15176, N14608);
buf BUFF1_11145 (N15177, N14349);
buf BUFF1_11146 (N15180, N14405);
buf BUFF1_11147 (N15183, N14357);
buf BUFF1_11148 (N15186, N14357);
buf BUFF1_11149 (N15189, N14364);
buf BUFF1_11150 (N15192, N14364);
buf BUFF1_11151 (N15195, N14385);
not NOT1_11152 (N15198, N14646);
buf BUFF1_11153 (N15199, N14418);
buf BUFF1_11154 (N15202, N14425);
buf BUFF1_11155 (N15205, N14445);
buf BUFF1_11156 (N15208, N14418);
buf BUFF1_11157 (N15211, N14425);
buf BUFF1_11158 (N15214, N14477);
buf BUFF1_11159 (N15217, N14469);
buf BUFF1_11160 (N15220, N14477);
not NOT1_11161 (N15223, N14662);
not NOT1_11162 (N15224, N14665);
not NOT1_11163 (N15225, N14668);
not NOT1_11164 (N15226, N14671);
not NOT1_11165 (N15227, N14689);
not NOT1_11166 (N15228, N14692);
not NOT1_11167 (N15229, N14695);
not NOT1_11168 (N15230, N14698);
nand NAND2_11169 (N15232, N14240, N15052);
nand NAND2_11170 (N15233, N14237, N15053);
nand NAND2_11171 (N15234, N14258, N15055);
nand NAND2_11172 (N15235, N14255, N15056);
nand NAND2_11173 (N15236, N14721, N15057);
nand NAND2_11174 (N15239, N13824, N15058);
and AND3_11175 (N15240, N15060, N15061, N14270);
not NOT1_11176 (N15241, N14939);
nand NAND2_11177 (N15242, N11824, N15069);
nand NAND2_11178 (N15243, N11827, N15071);
nand NAND2_11179 (N15244, N11830, N15073);
nand NAND2_11180 (N15245, N11833, N15075);
nand NAND2_11181 (N15246, N11836, N15077);
nand NAND2_11182 (N15247, N11839, N15079);
nand NAND2_11183 (N15248, N11842, N15081);
nand NAND2_11184 (N15249, N11845, N15083);
nand NAND2_11185 (N15250, N11848, N15085);
nand NAND2_11186 (N15252, N11854, N15089);
nand NAND2_11187 (N15253, N11857, N15091);
nand NAND2_11188 (N15254, N11860, N15093);
nand NAND2_11189 (N15255, N11863, N15095);
nand NAND2_11190 (N15256, N11866, N15097);
nand NAND2_11191 (N15257, N11869, N15099);
nand NAND2_11192 (N15258, N11872, N15101);
nand NAND2_11193 (N15259, N11875, N15103);
nand NAND2_11194 (N15260, N11878, N15105);
nand NAND2_11195 (N15261, N11881, N15106);
nand NAND2_11196 (N15262, N11884, N15108);
nand NAND2_11197 (N15263, N11887, N15110);
nand NAND2_11198 (N15264, N15112, N14856);
nand NAND2_11199 (N15274, N11893, N15113);
nand NAND2_11200 (N15275, N11896, N15115);
nand NAND2_11201 (N15282, N11902, N15122);
nand NAND2_11202 (N15283, N11905, N15124);
nand NAND2_11203 (N15284, N14908, N15125);
nand NAND2_11204 (N15298, N11911, N15127);
nand NAND2_11205 (N15299, N11914, N15129);
nand NAND2_11206 (N15300, N11917, N15131);
nand NAND2_11207 (N15303, N14652, N15135);
nand NAND2_11208 (N15304, N14649, N15136);
nand NAND2_11209 (N15305, N14008, N15138);
nand NAND2_11210 (N15306, N14219, N15139);
nand NAND2_11211 (N15307, N14677, N15141);
nand NAND2_11212 (N15308, N14674, N15142);
nand NAND2_11213 (N15309, N14683, N15143);
nand NAND2_11214 (N15310, N14680, N15144);
nand NAND2_11215 (N15311, N14011, N15146);
not NOT1_11216 (N15312, N15049);
nand NAND2_11217 (N15315, N15153, N15154);
nand NAND2_11218 (N15319, N15155, N15156);
nand NAND2_11219 (N15324, N15160, N15161);
nand NAND2_11220 (N15328, N15162, N14975);
nor N1OR2_11221 (N15331, N15163, N14978);
nor N1OR2_11222 (N15332, N15164, N14979);
or OR2_11223 (N15346, N14412, N15119);
nand NAND2_11224 (N15363, N14665, N15223);
nand NAND2_11225 (N15364, N14662, N15224);
nand NAND2_11226 (N15365, N14671, N15225);
nand NAND2_11227 (N15366, N14668, N15226);
nand NAND2_11228 (N15367, N14692, N15227);
nand NAND2_11229 (N15368, N14689, N15228);
nand NAND2_11230 (N15369, N14698, N15229);
nand NAND2_11231 (N15370, N14695, N15230);
nand NAND2_11232 (N15371, N15148, N15147);
buf BUFF1_11233 (N15374, N14939);
nand NAND2_11234 (N15377, N15232, N15233);
nand NAND2_11235 (N15382, N15234, N15235);
nand NAND2_11236 (N15385, N15239, N15059);
and AND3_11237 (N15388, N15062, N15063, N15241);
nand NAND2_11238 (N15389, N15242, N15070);
nand NAND2_11239 (N15396, N15243, N15072);
nand NAND2_11240 (N15407, N15244, N15074);
nand NAND2_11241 (N15418, N15245, N15076);
nand NAND2_11242 (N15424, N15246, N15078);
nand NAND2_11243 (N15431, N15247, N15080);
nand NAND2_11244 (N15441, N15248, N15082);
nand NAND2_11245 (N15452, N15249, N15084);
nand NAND2_11246 (N15462, N15250, N15086);
not NOT1_11247 (N15469, N15169);
nand NAND2_11248 (N15470, N15088, N15252);
nand NAND2_11249 (N15477, N15090, N15253);
nand NAND2_11250 (N15488, N15092, N15254);
nand NAND2_11251 (N15498, N15094, N15255);
nand NAND2_11252 (N15506, N15096, N15256);
nand NAND2_11253 (N15520, N15098, N15257);
nand NAND2_11254 (N15536, N15100, N15258);
nand NAND2_11255 (N15549, N15102, N15259);
nand NAND2_11256 (N15555, N15104, N15260);
nand NAND2_11257 (N15562, N15261, N15107);
nand NAND2_11258 (N15573, N15262, N15109);
nand NAND2_11259 (N15579, N15263, N15111);
nand NAND2_11260 (N15595, N15274, N15114);
nand NAND2_11261 (N15606, N15275, N15116);
nand NAND2_11262 (N15616, N15180, N12715);
not NOT1_11263 (N15617, N15180);
not NOT1_11264 (N15618, N15183);
not NOT1_11265 (N15619, N15186);
not NOT1_11266 (N15620, N15189);
not NOT1_11267 (N15621, N15192);
not NOT1_11268 (N15622, N15195);
nand NAND2_11269 (N15624, N15121, N15282);
nand NAND2_11270 (N15634, N15123, N15283);
nand NAND2_11271 (N15655, N15126, N15298);
nand NAND2_11272 (N15671, N15128, N15299);
nand NAND2_11273 (N15684, N15130, N15300);
not NOT1_11274 (N15690, N15202);
not NOT1_11275 (N15691, N15211);
nand NAND2_11276 (N15692, N15303, N15304);
nand NAND2_11277 (N15696, N15137, N15305);
nand NAND2_11278 (N15700, N15306, N15140);
nand NAND2_11279 (N15703, N15307, N15308);
nand NAND2_11280 (N15707, N15309, N15310);
nand NAND2_11281 (N15711, N15145, N15311);
and AND2_11282 (N15726, N15166, N14512);
not NOT1_11283 (N15727, N15173);
not NOT1_11284 (N15728, N15177);
not NOT1_11285 (N15730, N15199);
not NOT1_11286 (N15731, N15205);
not NOT1_11287 (N15732, N15208);
not NOT1_11288 (N15733, N15214);
not NOT1_11289 (N15734, N15217);
not NOT1_11290 (N15735, N15220);
nand NAND2_11291 (N15736, N15365, N15366);
nand NAND2_11292 (N15739, N15363, N15364);
nand NAND2_11293 (N15742, N15369, N15370);
nand NAND2_11294 (N15745, N15367, N15368);
not NOT1_11295 (N15755, N15236);
nand NAND2_11296 (N15756, N15332, N15331);
and AND2_11297 (N15954, N15264, N14396);
nand NAND2_11298 (N15955, N11899, N15617);
not NOT1_11299 (N15956, N15346);
and AND2_11300 (N16005, N15284, N14456);
and AND2_11301 (N16006, N15284, N14456);
not NOT1_11302 (N16023, N15371);
nand NAND2_11303 (N16024, N15371, N15312);
not NOT1_11304 (N16025, N15315);
not NOT1_11305 (N16028, N15324);
buf BUFF1_11306 (N16031, N15319);
buf BUFF1_11307 (N16034, N15319);
buf BUFF1_11308 (N16037, N15328);
buf BUFF1_11309 (N16040, N15328);
not NOT1_11310 (N16044, N15385);
or OR2_11311 (N16045, N15166, N15726);
buf BUFF1_11312 (N16048, N15264);
buf BUFF1_11313 (N16051, N15284);
buf BUFF1_11314 (N16054, N15284);
not NOT1_11315 (N16065, N15374);
nand NAND2_11316 (N16066, N15374, N15054);
not NOT1_11317 (N16067, N15377);
not NOT1_11318 (N16068, N15382);
nand NAND2_11319 (N16069, N15382, N15755);
and AND2_11320 (N16071, N15470, N14316);
and AND3_11321 (N16072, N15477, N15470, N14320);
and AND4_11322 (N16073, N15488, N15470, N14325, N15477);
and AND4_11323 (N16074, N15562, N14357, N14385, N14364);
and AND2_11324 (N16075, N15389, N14280);
and AND3_11325 (N16076, N15396, N15389, N14284);
and AND4_11326 (N16077, N15407, N15389, N14290, N15396);
and AND4_11327 (N16078, N15624, N14418, N14445, N14425);
not NOT1_11328 (N16079, N15418);
and AND4_11329 (N16080, N15396, N15418, N15407, N15389);
and AND2_11330 (N16083, N15396, N14284);
and AND3_11331 (N16084, N15407, N14290, N15396);
and AND3_11332 (N16085, N15418, N15407, N15396);
and AND2_11333 (N16086, N15396, N14284);
and AND3_11334 (N16087, N14290, N15407, N15396);
and AND2_11335 (N16088, N15407, N14290);
and AND2_11336 (N16089, N15418, N15407);
and AND2_11337 (N16090, N15407, N14290);
and AND5_11338 (N16091, N15431, N15462, N15441, N15424, N15452);
and AND2_11339 (N16094, N15424, N14298);
and AND3_11340 (N16095, N15431, N15424, N14301);
and AND4_11341 (N16096, N15441, N15424, N14305, N15431);
and AND5_11342 (N16097, N15452, N15441, N15424, N14310, N15431);
and AND2_11343 (N16098, N15431, N14301);
and AND3_11344 (N16099, N15441, N14305, N15431);
and AND4_11345 (N16100, N15452, N15441, N14310, N15431);
and AND5_11346 (N16101, N14, N15462, N15441, N15452, N15431);
and AND2_11347 (N16102, N14305, N15441);
and AND3_11348 (N16103, N15452, N15441, N14310);
and AND4_11349 (N16104, N14, N15462, N15441, N15452);
and AND2_11350 (N16105, N15452, N14310);
and AND3_11351 (N16106, N14, N15462, N15452);
and AND2_11352 (N16107, N14, N15462);
and AND4_11353 (N16108, N15549, N15488, N15477, N15470);
and AND2_11354 (N16111, N15477, N14320);
and AND3_11355 (N16112, N15488, N14325, N15477);
and AND3_11356 (N16113, N15549, N15488, N15477);
and AND2_11357 (N16114, N15477, N14320);
and AND3_11358 (N16115, N15488, N14325, N15477);
and AND2_11359 (N16116, N15488, N14325);
and AND5_11360 (N16117, N15555, N15536, N15520, N15506, N15498);
and AND2_11361 (N16120, N15498, N14332);
and AND3_11362 (N16121, N15506, N15498, N14336);
and AND4_11363 (N16122, N15520, N15498, N14342, N15506);
and AND5_11364 (N16123, N15536, N15520, N15498, N14349, N15506);
and AND2_11365 (N16124, N15506, N14336);
and AND3_11366 (N16125, N15520, N14342, N15506);
and AND4_11367 (N16126, N15536, N15520, N14349, N15506);
and AND4_11368 (N16127, N15555, N15520, N15506, N15536);
and AND2_11369 (N16128, N15506, N14336);
and AND3_11370 (N16129, N15520, N14342, N15506);
and AND4_11371 (N16130, N15536, N15520, N14349, N15506);
and AND2_11372 (N16131, N15520, N14342);
and AND3_11373 (N16132, N15536, N15520, N14349);
and AND3_11374 (N16133, N15555, N15520, N15536);
and AND2_11375 (N16134, N15520, N14342);
and AND3_11376 (N16135, N15536, N15520, N14349);
and AND2_11377 (N16136, N15536, N14349);
and AND2_11378 (N16137, N15549, N15488);
and AND2_11379 (N16138, N15555, N15536);
not NOT1_11380 (N16139, N15573);
and AND4_11381 (N16140, N14364, N15573, N15562, N14357);
and AND3_11382 (N16143, N15562, N14385, N14364);
and AND3_11383 (N16144, N15573, N15562, N14364);
and AND3_11384 (N16145, N14385, N15562, N14364);
and AND2_11385 (N16146, N15562, N14385);
and AND2_11386 (N16147, N15573, N15562);
and AND2_11387 (N16148, N15562, N14385);
and AND5_11388 (N16149, N15264, N14405, N15595, N15579, N15606);
and AND2_11389 (N16152, N15579, N14067);
and AND3_11390 (N16153, N15264, N15579, N14396);
and AND4_11391 (N16154, N15595, N15579, N14400, N15264);
and AND5_11392 (N16155, N15606, N15595, N15579, N14412, N15264);
and AND3_11393 (N16156, N15595, N14400, N15264);
and AND4_11394 (N16157, N15606, N15595, N14412, N15264);
and AND5_11395 (N16158, N154, N14405, N15595, N15606, N15264);
and AND2_11396 (N16159, N14400, N15595);
and AND3_11397 (N16160, N15606, N15595, N14412);
and AND4_11398 (N16161, N154, N14405, N15595, N15606);
and AND2_11399 (N16162, N15606, N14412);
and AND3_11400 (N16163, N154, N14405, N15606);
nand NAND2_11401 (N16164, N15616, N15955);
and AND4_11402 (N16168, N15684, N15624, N14425, N14418);
and AND3_11403 (N16171, N15624, N14445, N14425);
and AND3_11404 (N16172, N15684, N15624, N14425);
and AND3_11405 (N16173, N15624, N14445, N14425);
and AND2_11406 (N16174, N15624, N14445);
and AND5_11407 (N16175, N14477, N15671, N15655, N15284, N15634);
and AND2_11408 (N16178, N15634, N14080);
and AND3_11409 (N16179, N15284, N15634, N14456);
and AND4_11410 (N16180, N15655, N15634, N14462, N15284);
and AND5_11411 (N16181, N15671, N15655, N15634, N14469, N15284);
and AND3_11412 (N16182, N15655, N14462, N15284);
and AND4_11413 (N16183, N15671, N15655, N14469, N15284);
and AND4_11414 (N16184, N14477, N15655, N15284, N15671);
and AND3_11415 (N16185, N15655, N14462, N15284);
and AND4_11416 (N16186, N15671, N15655, N14469, N15284);
and AND2_11417 (N16187, N15655, N14462);
and AND3_11418 (N16188, N15671, N15655, N14469);
and AND3_11419 (N16189, N14477, N15655, N15671);
and AND2_11420 (N16190, N15655, N14462);
and AND3_11421 (N16191, N15671, N15655, N14469);
and AND2_11422 (N16192, N15671, N14469);
and AND2_11423 (N16193, N15684, N15624);
and AND2_11424 (N16194, N14477, N15671);
not NOT1_11425 (N16197, N15692);
not NOT1_11426 (N16200, N15696);
not NOT1_11427 (N16203, N15703);
not NOT1_11428 (N16206, N15707);
buf BUFF1_11429 (N16209, N15700);
buf BUFF1_11430 (N16212, N15700);
buf BUFF1_11431 (N16215, N15711);
buf BUFF1_11432 (N16218, N15711);
nand NAND2_11433 (N16221, N15049, N16023);
not NOT1_11434 (N16234, N15756);
nand NAND2_11435 (N16235, N15756, N16044);
buf BUFF1_11436 (N16238, N15462);
buf BUFF1_11437 (N16241, N15389);
buf BUFF1_11438 (N16244, N15389);
buf BUFF1_11439 (N16247, N15396);
buf BUFF1_11440 (N16250, N15396);
buf BUFF1_11441 (N16253, N15407);
buf BUFF1_11442 (N16256, N15407);
buf BUFF1_11443 (N16259, N15424);
buf BUFF1_11444 (N16262, N15431);
buf BUFF1_11445 (N16265, N15441);
buf BUFF1_11446 (N16268, N15452);
buf BUFF1_11447 (N16271, N15549);
buf BUFF1_11448 (N16274, N15488);
buf BUFF1_11449 (N16277, N15470);
buf BUFF1_11450 (N16280, N15477);
buf BUFF1_11451 (N16283, N15549);
buf BUFF1_11452 (N16286, N15488);
buf BUFF1_11453 (N16289, N15470);
buf BUFF1_11454 (N16292, N15477);
buf BUFF1_11455 (N16295, N15555);
buf BUFF1_11456 (N16298, N15536);
buf BUFF1_11457 (N16301, N15498);
buf BUFF1_11458 (N16304, N15520);
buf BUFF1_11459 (N16307, N15506);
buf BUFF1_11460 (N16310, N15506);
buf BUFF1_11461 (N16313, N15555);
buf BUFF1_11462 (N16316, N15536);
buf BUFF1_11463 (N16319, N15498);
buf BUFF1_11464 (N16322, N15520);
buf BUFF1_11465 (N16325, N15562);
buf BUFF1_11466 (N16328, N15562);
buf BUFF1_11467 (N16331, N15579);
buf BUFF1_11468 (N16335, N15595);
buf BUFF1_11469 (N16338, N15606);
buf BUFF1_11470 (N16341, N15684);
buf BUFF1_11471 (N16344, N15624);
buf BUFF1_11472 (N16347, N15684);
buf BUFF1_11473 (N16350, N15624);
buf BUFF1_11474 (N16353, N15671);
buf BUFF1_11475 (N16356, N15634);
buf BUFF1_11476 (N16359, N15655);
buf BUFF1_11477 (N16364, N15671);
buf BUFF1_11478 (N16367, N15634);
buf BUFF1_11479 (N16370, N15655);
not NOT1_11480 (N16373, N15736);
not NOT1_11481 (N16374, N15739);
not NOT1_11482 (N16375, N15742);
not NOT1_11483 (N16376, N15745);
nand NAND2_11484 (N16377, N14243, N16065);
nand NAND2_11485 (N16378, N15236, N16068);
or OR4_11486 (N16382, N14268, N16071, N16072, N16073);
or OR4_11487 (N16386, N13968, N15065, N15066, N16074);
or OR4_11488 (N16388, N14271, N16075, N16076, N16077);
or OR4_11489 (N16392, N13968, N15067, N15068, N16078);
or OR5_11490 (N16397, N14297, N16094, N16095, N16096, N16097);
or OR2_11491 (N16411, N14320, N16116);
or OR5_11492 (N16415, N14331, N16120, N16121, N16122, N16123);
or OR2_11493 (N16419, N14342, N16136);
or OR5_11494 (N16427, N14392, N16152, N16153, N16154, N16155);
not NOT1_11495 (N16434, N16048);
or OR2_11496 (N16437, N14440, N16174);
or OR5_11497 (N16441, N14451, N16178, N16179, N16180, N16181);
or OR2_11498 (N16445, N14462, N16192);
not NOT1_11499 (N16448, N16051);
not NOT1_11500 (N16449, N16054);
nand NAND2_11501 (N16466, N16221, N16024);
not NOT1_11502 (N16469, N16031);
not NOT1_11503 (N16470, N16034);
not NOT1_11504 (N16471, N16037);
not NOT1_11505 (N16472, N16040);
and AND3_11506 (N16473, N15315, N14524, N16031);
and AND3_11507 (N16474, N16025, N15150, N16034);
and AND3_11508 (N16475, N15324, N14532, N16037);
and AND3_11509 (N16476, N16028, N15157, N16040);
nand NAND2_11510 (N16477, N15385, N16234);
nand NAND2_11511 (N16478, N16045, N1132);
or OR4_11512 (N16482, N14280, N16083, N16084, N16085);
nor N1OR3_11513 (N16486, N14280, N16086, N16087);
or OR3_11514 (N16490, N14284, N16088, N16089);
nor N1OR2_11515 (N16494, N14284, N16090);
or OR5_11516 (N16500, N14298, N16098, N16099, N16100, N16101);
or OR4_11517 (N16504, N14301, N16102, N16103, N16104);
or OR3_11518 (N16508, N14305, N16105, N16106);
or OR2_11519 (N16512, N14310, N16107);
or OR4_11520 (N16516, N14316, N16111, N16112, N16113);
nor N1OR3_11521 (N16526, N14316, N16114, N16115);
or OR4_11522 (N16536, N14336, N16131, N16132, N16133);
or OR5_11523 (N16539, N14332, N16124, N16125, N16126, N16127);
nor N1OR3_11524 (N16553, N14336, N16134, N16135);
nor N1OR4_11525 (N16556, N14332, N16128, N16129, N16130);
or OR4_11526 (N16566, N14375, N15117, N16143, N16144);
nor N1OR3_11527 (N16569, N14375, N15118, N16145);
or OR3_11528 (N16572, N14379, N16146, N16147);
nor N1OR2_11529 (N16575, N14379, N16148);
or OR5_11530 (N16580, N14067, N15954, N16156, N16157, N16158);
or OR4_11531 (N16584, N14396, N16159, N16160, N16161);
or OR3_11532 (N16587, N14400, N16162, N16163);
or OR4_11533 (N16592, N14436, N15132, N16171, N16172);
nor N1OR3_11534 (N16599, N14436, N15133, N16173);
or OR4_11535 (N16606, N14456, N16187, N16188, N16189);
or OR5_11536 (N16609, N14080, N16005, N16182, N16183, N16184);
nor N1OR3_11537 (N16619, N14456, N16190, N16191);
nor N1OR4_11538 (N16622, N14080, N16006, N16185, N16186);
nand NAND2_11539 (N16630, N15739, N16373);
nand NAND2_11540 (N16631, N15736, N16374);
nand NAND2_11541 (N16632, N15745, N16375);
nand NAND2_11542 (N16633, N15742, N16376);
nand NAND2_11543 (N16634, N16377, N16066);
nand NAND2_11544 (N16637, N16069, N16378);
not NOT1_11545 (N16640, N16164);
and AND2_11546 (N16641, N16108, N16117);
and AND2_11547 (N16643, N16140, N16149);
and AND2_11548 (N16646, N16168, N16175);
and AND2_11549 (N16648, N16080, N16091);
nand NAND2_11550 (N16650, N16238, N12637);
not NOT1_11551 (N16651, N16238);
not NOT1_11552 (N16653, N16241);
not NOT1_11553 (N16655, N16244);
not NOT1_11554 (N16657, N16247);
not NOT1_11555 (N16659, N16250);
nand NAND2_11556 (N16660, N16253, N15087);
not NOT1_11557 (N16661, N16253);
nand NAND2_11558 (N16662, N16256, N15469);
not NOT1_11559 (N16663, N16256);
and AND2_11560 (N16664, N16091, N14);
not NOT1_11561 (N16666, N16259);
not NOT1_11562 (N16668, N16262);
not NOT1_11563 (N16670, N16265);
not NOT1_11564 (N16672, N16268);
not NOT1_11565 (N16675, N16117);
not NOT1_11566 (N16680, N16280);
not NOT1_11567 (N16681, N16292);
not NOT1_11568 (N16682, N16307);
not NOT1_11569 (N16683, N16310);
nand NAND2_11570 (N16689, N16325, N15120);
not NOT1_11571 (N16690, N16325);
nand NAND2_11572 (N16691, N16328, N15622);
not NOT1_11573 (N16692, N16328);
and AND2_11574 (N16693, N16149, N154);
not NOT1_11575 (N16695, N16331);
not NOT1_11576 (N16698, N16335);
nand NAND2_11577 (N16699, N16338, N15956);
not NOT1_11578 (N16700, N16338);
not NOT1_11579 (N16703, N16175);
not NOT1_11580 (N16708, N16209);
not NOT1_11581 (N16709, N16212);
not NOT1_11582 (N16710, N16215);
not NOT1_11583 (N16711, N16218);
and AND3_11584 (N16712, N15696, N15692, N16209);
and AND3_11585 (N16713, N16200, N16197, N16212);
and AND3_11586 (N16714, N15707, N15703, N16215);
and AND3_11587 (N16715, N16206, N16203, N16218);
buf BUFF1_11588 (N16716, N16466);
and AND3_11589 (N16718, N16164, N11777, N13130);
and AND3_11590 (N16719, N15150, N15315, N16469);
and AND3_11591 (N16720, N14524, N16025, N16470);
and AND3_11592 (N16721, N15157, N15324, N16471);
and AND3_11593 (N16722, N14532, N16028, N16472);
nand NAND2_11594 (N16724, N16477, N16235);
not NOT1_11595 (N16739, N16271);
not NOT1_11596 (N16740, N16274);
not NOT1_11597 (N16741, N16277);
not NOT1_11598 (N16744, N16283);
not NOT1_11599 (N16745, N16286);
not NOT1_11600 (N16746, N16289);
not NOT1_11601 (N16751, N16295);
not NOT1_11602 (N16752, N16298);
not NOT1_11603 (N16753, N16301);
not NOT1_11604 (N16754, N16304);
not NOT1_11605 (N16755, N16322);
not NOT1_11606 (N16760, N16313);
not NOT1_11607 (N16761, N16316);
not NOT1_11608 (N16762, N16319);
not NOT1_11609 (N16772, N16341);
not NOT1_11610 (N16773, N16344);
not NOT1_11611 (N16776, N16347);
not NOT1_11612 (N16777, N16350);
not NOT1_11613 (N16782, N16353);
not NOT1_11614 (N16783, N16356);
not NOT1_11615 (N16784, N16359);
not NOT1_11616 (N16785, N16370);
not NOT1_11617 (N16790, N16364);
not NOT1_11618 (N16791, N16367);
nand NAND2_11619 (N16792, N16630, N16631);
nand NAND2_11620 (N16795, N16632, N16633);
and AND2_11621 (N16801, N16108, N16415);
and AND2_11622 (N16802, N16427, N16140);
and AND2_11623 (N16803, N16397, N16080);
and AND2_11624 (N16804, N16168, N16441);
not NOT1_11625 (N16805, N16466);
nand NAND2_11626 (N16806, N11851, N16651);
not NOT1_11627 (N16807, N16482);
nand NAND2_11628 (N16808, N16482, N16653);
not NOT1_11629 (N16809, N16486);
nand NAND2_11630 (N16810, N16486, N16655);
not NOT1_11631 (N16811, N16490);
nand NAND2_11632 (N16812, N16490, N16657);
not NOT1_11633 (N16813, N16494);
nand NAND2_11634 (N16814, N16494, N16659);
nand NAND2_11635 (N16815, N14575, N16661);
nand NAND2_11636 (N16816, N15169, N16663);
or OR2_11637 (N16817, N16397, N16664);
not NOT1_11638 (N16823, N16500);
nand NAND2_11639 (N16824, N16500, N16666);
not NOT1_11640 (N16825, N16504);
nand NAND2_11641 (N16826, N16504, N16668);
not NOT1_11642 (N16827, N16508);
nand NAND2_11643 (N16828, N16508, N16670);
not NOT1_11644 (N16829, N16512);
nand NAND2_11645 (N16830, N16512, N16672);
not NOT1_11646 (N16831, N16415);
not NOT1_11647 (N16834, N16566);
nand NAND2_11648 (N16835, N16566, N15618);
not NOT1_11649 (N16836, N16569);
nand NAND2_11650 (N16837, N16569, N15619);
not NOT1_11651 (N16838, N16572);
nand NAND2_11652 (N16839, N16572, N15620);
not NOT1_11653 (N16840, N16575);
nand NAND2_11654 (N16841, N16575, N15621);
nand NAND2_11655 (N16842, N14627, N16690);
nand NAND2_11656 (N16843, N15195, N16692);
or OR2_11657 (N16844, N16427, N16693);
not NOT1_11658 (N16850, N16580);
nand NAND2_11659 (N16851, N16580, N16695);
not NOT1_11660 (N16852, N16584);
nand NAND2_11661 (N16853, N16584, N16434);
not NOT1_11662 (N16854, N16587);
nand NAND2_11663 (N16855, N16587, N16698);
nand NAND2_11664 (N16856, N15346, N16700);
not NOT1_11665 (N16857, N16441);
and AND3_11666 (N16860, N16197, N15696, N16708);
and AND3_11667 (N16861, N15692, N16200, N16709);
and AND3_11668 (N16862, N16203, N15707, N16710);
and AND3_11669 (N16863, N15703, N16206, N16711);
or OR3_11670 (N16866, N14197, N16718, N13785);
nor N1OR2_11671 (N16872, N16719, N16473);
nor N1OR2_11672 (N16873, N16720, N16474);
nor N1OR2_11673 (N16874, N16721, N16475);
nor N1OR2_11674 (N16875, N16722, N16476);
not NOT1_11675 (N16876, N16637);
buf BUFF1_11676 (N16877, N16724);
and AND2_11677 (N16879, N16045, N16478);
and AND2_11678 (N16880, N16478, N1132);
or OR2_11679 (N16881, N16411, N16137);
not NOT1_11680 (N16884, N16516);
not NOT1_11681 (N16885, N16411);
not NOT1_11682 (N16888, N16526);
not NOT1_11683 (N16889, N16536);
nand NAND2_11684 (N16890, N16536, N15176);
or OR2_11685 (N16891, N16419, N16138);
not NOT1_11686 (N16894, N16539);
not NOT1_11687 (N16895, N16553);
nand NAND2_11688 (N16896, N16553, N15728);
not NOT1_11689 (N16897, N16419);
not NOT1_11690 (N16900, N16556);
or OR2_11691 (N16901, N16437, N16193);
not NOT1_11692 (N16904, N16592);
not NOT1_11693 (N16905, N16437);
not NOT1_11694 (N16908, N16599);
or OR2_11695 (N16909, N16445, N16194);
not NOT1_11696 (N16912, N16606);
not NOT1_11697 (N16913, N16609);
not NOT1_11698 (N16914, N16619);
nand NAND2_11699 (N16915, N16619, N15734);
not NOT1_11700 (N16916, N16445);
not NOT1_11701 (N16919, N16622);
not NOT1_11702 (N16922, N16634);
nand NAND2_11703 (N16923, N16634, N16067);
or OR2_11704 (N16924, N16382, N16801);
or OR2_11705 (N16925, N16386, N16802);
or OR2_11706 (N16926, N16388, N16803);
or OR2_11707 (N16927, N16392, N16804);
not NOT1_11708 (N16930, N16724);
nand NAND2_11709 (N16932, N16650, N16806);
nand NAND2_11710 (N16935, N16241, N16807);
nand NAND2_11711 (N16936, N16244, N16809);
nand NAND2_11712 (N16937, N16247, N16811);
nand NAND2_11713 (N16938, N16250, N16813);
nand NAND2_11714 (N16939, N16660, N16815);
nand NAND2_11715 (N16940, N16662, N16816);
nand NAND2_11716 (N16946, N16259, N16823);
nand NAND2_11717 (N16947, N16262, N16825);
nand NAND2_11718 (N16948, N16265, N16827);
nand NAND2_11719 (N16949, N16268, N16829);
nand NAND2_11720 (N16953, N15183, N16834);
nand NAND2_11721 (N16954, N15186, N16836);
nand NAND2_11722 (N16955, N15189, N16838);
nand NAND2_11723 (N16956, N15192, N16840);
nand NAND2_11724 (N16957, N16689, N16842);
nand NAND2_11725 (N16958, N16691, N16843);
nand NAND2_11726 (N16964, N16331, N16850);
nand NAND2_11727 (N16965, N16048, N16852);
nand NAND2_11728 (N16966, N16335, N16854);
nand NAND2_11729 (N16967, N16699, N16856);
nor N1OR2_11730 (N16973, N16860, N16712);
nor N1OR2_11731 (N16974, N16861, N16713);
nor N1OR2_11732 (N16975, N16862, N16714);
nor N1OR2_11733 (N16976, N16863, N16715);
not NOT1_11734 (N16977, N16792);
not NOT1_11735 (N16978, N16795);
or OR2_11736 (N16979, N16879, N16880);
nand NAND2_11737 (N16987, N14608, N16889);
nand NAND2_11738 (N16990, N15177, N16895);
nand NAND2_11739 (N16999, N15217, N16914);
nand NAND2_11740 (N17002, N15377, N16922);
nand NAND2_11741 (N17003, N16873, N16872);
nand NAND2_11742 (N17006, N16875, N16874);
and AND3_11743 (N17011, N16866, N12681, N12692);
and AND3_11744 (N17012, N16866, N12756, N12767);
and AND3_11745 (N17013, N16866, N12779, N12790);
not NOT1_11746 (N17015, N16866);
and AND3_11747 (N17016, N16866, N12801, N12812);
nand NAND2_11748 (N17018, N16935, N16808);
nand NAND2_11749 (N17019, N16936, N16810);
nand NAND2_11750 (N17020, N16937, N16812);
nand NAND2_11751 (N17021, N16938, N16814);
not NOT1_11752 (N17022, N16939);
not NOT1_11753 (N17023, N16817);
nand NAND2_11754 (N17028, N16946, N16824);
nand NAND2_11755 (N17031, N16947, N16826);
nand NAND2_11756 (N17034, N16948, N16828);
nand NAND2_11757 (N17037, N16949, N16830);
and AND2_11758 (N17040, N16817, N16079);
and AND2_11759 (N17041, N16831, N16675);
nand NAND2_11760 (N17044, N16953, N16835);
nand NAND2_11761 (N17045, N16954, N16837);
nand NAND2_11762 (N17046, N16955, N16839);
nand NAND2_11763 (N17047, N16956, N16841);
not NOT1_11764 (N17048, N16957);
not NOT1_11765 (N17049, N16844);
nand NAND2_11766 (N17054, N16964, N16851);
nand NAND2_11767 (N17057, N16965, N16853);
nand NAND2_11768 (N17060, N16966, N16855);
and AND2_11769 (N17064, N16844, N16139);
and AND2_11770 (N17065, N16857, N16703);
not NOT1_11771 (N17072, N16881);
nand NAND2_11772 (N17073, N16881, N15172);
not NOT1_11773 (N17074, N16885);
nand NAND2_11774 (N17075, N16885, N15727);
nand NAND2_11775 (N17076, N16890, N16987);
not NOT1_11776 (N17079, N16891);
nand NAND2_11777 (N17080, N16896, N16990);
not NOT1_11778 (N17083, N16897);
not NOT1_11779 (N17084, N16901);
nand NAND2_11780 (N17085, N16901, N15198);
not NOT1_11781 (N17086, N16905);
nand NAND2_11782 (N17087, N16905, N15731);
not NOT1_11783 (N17088, N16909);
nand NAND2_11784 (N17089, N16909, N16912);
nand NAND2_11785 (N17090, N16915, N16999);
not NOT1_11786 (N17093, N16916);
nand NAND2_11787 (N17094, N16974, N16973);
nand NAND2_11788 (N17097, N16976, N16975);
nand NAND2_11789 (N17101, N17002, N16923);
not NOT1_11790 (N17105, N16932);
not NOT1_11791 (N17110, N16967);
and AND3_11792 (N17114, N16979, N1603, N11755);
not NOT1_11793 (N17115, N17019);
not NOT1_11794 (N17116, N17021);
and AND2_11795 (N17125, N16817, N17018);
and AND2_11796 (N17126, N16817, N17020);
and AND2_11797 (N17127, N16817, N17022);
not NOT1_11798 (N17130, N17045);
not NOT1_11799 (N17131, N17047);
and AND2_11800 (N17139, N16844, N17044);
and AND2_11801 (N17140, N16844, N17046);
and AND2_11802 (N17141, N16844, N17048);
and AND3_11803 (N17146, N16932, N11761, N13108);
and AND3_11804 (N17147, N16967, N11777, N13130);
not NOT1_11805 (N17149, N17003);
not NOT1_11806 (N17150, N17006);
nand NAND2_11807 (N17151, N17006, N16876);
nand NAND2_11808 (N17152, N14605, N17072);
nand NAND2_11809 (N17153, N15173, N17074);
nand NAND2_11810 (N17158, N14646, N17084);
nand NAND2_11811 (N17159, N15205, N17086);
nand NAND2_11812 (N17160, N16606, N17088);
not NOT1_11813 (N17166, N17037);
not NOT1_11814 (N17167, N17034);
not NOT1_11815 (N17168, N17031);
not NOT1_11816 (N17169, N17028);
not NOT1_11817 (N17170, N17060);
not NOT1_11818 (N17171, N17057);
not NOT1_11819 (N17172, N17054);
and AND2_11820 (N17173, N17115, N17023);
and AND2_11821 (N17174, N17116, N17023);
and AND2_11822 (N17175, N16940, N17023);
and AND2_11823 (N17176, N15418, N17023);
not NOT1_11824 (N17177, N17041);
and AND2_11825 (N17178, N17130, N17049);
and AND2_11826 (N17179, N17131, N17049);
and AND2_11827 (N17180, N16958, N17049);
and AND2_11828 (N17181, N15573, N17049);
not NOT1_11829 (N17182, N17065);
not NOT1_11830 (N17183, N17094);
nand NAND2_11831 (N17184, N17094, N16977);
not NOT1_11832 (N17185, N17097);
nand NAND2_11833 (N17186, N17097, N16978);
and AND3_11834 (N17187, N17037, N11761, N13108);
and AND3_11835 (N17188, N17034, N11761, N13108);
and AND3_11836 (N17189, N17031, N11761, N13108);
or OR3_11837 (N17190, N14956, N17146, N13781);
and AND3_11838 (N17196, N17060, N11777, N13130);
and AND3_11839 (N17197, N17057, N11777, N13130);
or OR3_11840 (N17198, N14960, N17147, N13786);
nand NAND2_11841 (N17204, N17101, N17149);
not NOT1_11842 (N17205, N17101);
nand NAND2_11843 (N17206, N16637, N17150);
and AND3_11844 (N17207, N17028, N11793, N13158);
and AND3_11845 (N17208, N17054, N11807, N13180);
nand NAND2_11846 (N17209, N17073, N17152);
nand NAND2_11847 (N17212, N17075, N17153);
not NOT1_11848 (N17215, N17076);
nand NAND2_11849 (N17216, N17076, N17079);
not NOT1_11850 (N17217, N17080);
nand NAND2_11851 (N17218, N17080, N17083);
nand NAND2_11852 (N17219, N17085, N17158);
nand NAND2_11853 (N17222, N17087, N17159);
nand NAND2_11854 (N17225, N17089, N17160);
not NOT1_11855 (N17228, N17090);
nand NAND2_11856 (N17229, N17090, N17093);
or OR2_11857 (N17236, N17173, N17125);
or OR2_11858 (N17239, N17174, N17126);
or OR2_11859 (N17242, N17175, N17127);
or OR2_11860 (N17245, N17176, N17040);
or OR2_11861 (N17250, N17178, N17139);
or OR2_11862 (N17257, N17179, N17140);
or OR2_11863 (N17260, N17180, N17141);
or OR2_11864 (N17263, N17181, N17064);
nand NAND2_11865 (N17268, N16792, N17183);
nand NAND2_11866 (N17269, N16795, N17185);
or OR3_11867 (N17270, N14957, N17187, N13782);
or OR3_11868 (N17276, N14958, N17188, N13783);
or OR3_11869 (N17282, N14959, N17189, N13784);
or OR3_11870 (N17288, N14961, N17196, N13787);
or OR3_11871 (N17294, N13998, N17197, N13788);
nand NAND2_11872 (N17300, N17003, N17205);
nand NAND2_11873 (N17301, N17206, N17151);
or OR3_11874 (N17304, N14980, N17207, N13800);
or OR3_11875 (N17310, N14984, N17208, N13805);
nand NAND2_11876 (N17320, N16891, N17215);
nand NAND2_11877 (N17321, N16897, N17217);
nand NAND2_11878 (N17328, N16916, N17228);
and AND3_11879 (N17338, N17190, N11185, N12692);
and AND3_11880 (N17339, N17198, N12681, N12692);
and AND3_11881 (N17340, N17190, N11247, N12767);
and AND3_11882 (N17341, N17198, N12756, N12767);
and AND3_11883 (N17342, N17190, N11327, N12790);
and AND3_11884 (N17349, N17198, N12779, N12790);
and AND3_11885 (N17357, N17198, N12801, N12812);
not NOT1_11886 (N17363, N17198);
and AND3_11887 (N17364, N17190, N11351, N12812);
not NOT1_11888 (N17365, N17190);
nand NAND2_11889 (N17394, N17268, N17184);
nand NAND2_11890 (N17397, N17269, N17186);
nand NAND2_11891 (N17402, N17204, N17300);
not NOT1_11892 (N17405, N17209);
nand NAND2_11893 (N17406, N17209, N16884);
not NOT1_11894 (N17407, N17212);
nand NAND2_11895 (N17408, N17212, N16888);
nand NAND2_11896 (N17409, N17320, N17216);
nand NAND2_11897 (N17412, N17321, N17218);
not NOT1_11898 (N17415, N17219);
nand NAND2_11899 (N17416, N17219, N16904);
not NOT1_11900 (N17417, N17222);
nand NAND2_11901 (N17418, N17222, N16908);
not NOT1_11902 (N17419, N17225);
nand NAND2_11903 (N17420, N17225, N16913);
nand NAND2_11904 (N17421, N17328, N17229);
not NOT1_11905 (N17424, N17245);
not NOT1_11906 (N17425, N17242);
not NOT1_11907 (N17426, N17239);
not NOT1_11908 (N17427, N17236);
not NOT1_11909 (N17428, N17263);
not NOT1_11910 (N17429, N17260);
not NOT1_11911 (N17430, N17257);
not NOT1_11912 (N17431, N17250);
not NOT1_11913 (N17432, N17250);
and AND3_11914 (N17433, N17310, N12653, N12664);
and AND3_11915 (N17434, N17304, N11161, N12664);
or OR4_11916 (N17435, N17011, N17338, N13621, N12591);
and AND3_11917 (N17436, N17270, N11185, N12692);
and AND3_11918 (N17437, N17288, N12681, N12692);
and AND3_11919 (N17438, N17276, N11185, N12692);
and AND3_11920 (N17439, N17294, N12681, N12692);
and AND3_11921 (N17440, N17282, N11185, N12692);
and AND3_11922 (N17441, N17310, N12728, N12739);
and AND3_11923 (N17442, N17304, N11223, N12739);
or OR4_11924 (N17443, N17012, N17340, N13632, N12600);
and AND3_11925 (N17444, N17270, N11247, N12767);
and AND3_11926 (N17445, N17288, N12756, N12767);
and AND3_11927 (N17446, N17276, N11247, N12767);
and AND3_11928 (N17447, N17294, N12756, N12767);
and AND3_11929 (N17448, N17282, N11247, N12767);
or OR4_11930 (N17449, N17013, N17342, N13641, N12605);
and AND3_11931 (N17450, N17310, N13041, N13052);
and AND3_11932 (N17451, N17304, N11697, N13052);
and AND3_11933 (N17452, N17294, N12779, N12790);
and AND3_11934 (N17453, N17282, N11327, N12790);
and AND3_11935 (N17454, N17288, N12779, N12790);
and AND3_11936 (N17455, N17276, N11327, N12790);
and AND3_11937 (N17456, N17270, N11327, N12790);
and AND3_11938 (N17457, N17310, N13075, N13086);
and AND3_11939 (N17458, N17304, N11731, N13086);
and AND3_11940 (N17459, N17294, N12801, N12812);
and AND3_11941 (N17460, N17282, N11351, N12812);
and AND3_11942 (N17461, N17288, N12801, N12812);
and AND3_11943 (N17462, N17276, N11351, N12812);
and AND3_11944 (N17463, N17270, N11351, N12812);
and AND3_11945 (N17464, N17250, N1603, N1599);
not NOT1_11946 (N17465, N17310);
not NOT1_11947 (N17466, N17294);
not NOT1_11948 (N17467, N17288);
not NOT1_11949 (N17468, N17301);
or OR4_11950 (N17469, N17016, N17364, N13660, N12626);
not NOT1_11951 (N17470, N17304);
not NOT1_11952 (N17471, N17282);
not NOT1_11953 (N17472, N17276);
not NOT1_11954 (N17473, N17270);
buf BUFF1_11955 (N17474, N17394);
buf BUFF1_11956 (N17476, N17397);
and AND2_11957 (N17479, N17301, N13068);
and AND3_11958 (N17481, N17245, N11793, N13158);
and AND3_11959 (N17482, N17242, N11793, N13158);
and AND3_11960 (N17483, N17239, N11793, N13158);
and AND3_11961 (N17484, N17236, N11793, N13158);
and AND3_11962 (N17485, N17263, N11807, N13180);
and AND3_11963 (N17486, N17260, N11807, N13180);
and AND3_11964 (N17487, N17257, N11807, N13180);
and AND3_11965 (N17488, N17250, N11807, N13180);
nand NAND2_11966 (N17489, N16979, N17250);
nand NAND2_11967 (N17492, N16516, N17405);
nand NAND2_11968 (N17493, N16526, N17407);
nand NAND2_11969 (N17498, N16592, N17415);
nand NAND2_11970 (N17499, N16599, N17417);
nand NAND2_11971 (N17500, N16609, N17419);
and AND9_11972 (N17503, N17105, N17166, N17167, N17168, N17169, N17424, N17425, N17426, N17427);
and AND9_11973 (N17504, N16640, N17110, N17170, N17171, N17172, N17428, N17429, N17430, N17431);
or OR4_11974 (N17505, N17433, N17434, N13616, N12585);
and AND2_11975 (N17506, N17435, N12675);
or OR4_11976 (N17507, N17339, N17436, N13622, N12592);
or OR4_11977 (N17508, N17437, N17438, N13623, N12593);
or OR4_11978 (N17509, N17439, N17440, N13624, N12594);
or OR4_11979 (N17510, N17441, N17442, N13627, N12595);
and AND2_11980 (N17511, N17443, N12750);
or OR4_11981 (N17512, N17341, N17444, N13633, N12601);
or OR4_11982 (N17513, N17445, N17446, N13634, N12602);
or OR4_11983 (N17514, N17447, N17448, N13635, N12603);
or OR4_11984 (N17515, N17450, N17451, N13646, N12610);
or OR4_11985 (N17516, N17452, N17453, N13647, N12611);
or OR4_11986 (N17517, N17454, N17455, N13648, N12612);
or OR4_11987 (N17518, N17349, N17456, N13649, N12613);
or OR4_11988 (N17519, N17457, N17458, N13654, N12618);
or OR4_11989 (N17520, N17459, N17460, N13655, N12619);
or OR4_11990 (N17521, N17461, N17462, N13656, N12620);
or OR4_11991 (N17522, N17357, N17463, N13657, N12621);
or OR4_11992 (N17525, N14741, N17114, N12624, N17464);
and AND3_11993 (N17526, N17468, N13119, N13130);
not NOT1_11994 (N17527, N17394);
not NOT1_11995 (N17528, N17397);
not NOT1_11996 (N17529, N17402);
and AND2_11997 (N17530, N17402, N13068);
or OR3_11998 (N17531, N14981, N17481, N13801);
or OR3_11999 (N17537, N14982, N17482, N13802);
or OR3_12000 (N17543, N14983, N17483, N13803);
or OR3_12001 (N17549, N15165, N17484, N13804);
or OR3_12002 (N17555, N14985, N17485, N13806);
or OR3_12003 (N17561, N14986, N17486, N13807);
or OR3_12004 (N17567, N14547, N17487, N13808);
or OR3_12005 (N17573, N14987, N17488, N13809);
nand NAND2_12006 (N17579, N17492, N17406);
nand NAND2_12007 (N17582, N17493, N17408);
not NOT1_12008 (N17585, N17409);
nand NAND2_12009 (N17586, N17409, N16894);
not NOT1_12010 (N17587, N17412);
nand NAND2_12011 (N17588, N17412, N16900);
nand NAND2_12012 (N17589, N17498, N17416);
nand NAND2_12013 (N17592, N17499, N17418);
nand NAND2_12014 (N17595, N17500, N17420);
not NOT1_12015 (N17598, N17421);
nand NAND2_12016 (N17599, N17421, N16919);
and AND2_12017 (N17600, N17505, N12647);
and AND2_12018 (N17601, N17507, N12675);
and AND2_12019 (N17602, N17508, N12675);
and AND2_12020 (N17603, N17509, N12675);
and AND2_12021 (N17604, N17510, N12722);
and AND2_12022 (N17605, N17512, N12750);
and AND2_12023 (N17606, N17513, N12750);
and AND2_12024 (N17607, N17514, N12750);
and AND2_12025 (N17624, N16979, N17489);
and AND2_12026 (N17625, N17489, N17250);
and AND2_12027 (N17626, N11149, N17525);
and AND5_12028 (N17631, N1562, N17527, N17528, N16805, N16930);
and AND3_12029 (N17636, N17529, N13097, N13108);
nand NAND2_12030 (N17657, N16539, N17585);
nand NAND2_12031 (N17658, N16556, N17587);
nand NAND2_12032 (N17665, N16622, N17598);
and AND3_12033 (N17666, N17555, N12653, N12664);
and AND3_12034 (N17667, N17531, N11161, N12664);
and AND3_12035 (N17668, N17561, N12653, N12664);
and AND3_12036 (N17669, N17537, N11161, N12664);
and AND3_12037 (N17670, N17567, N12653, N12664);
and AND3_12038 (N17671, N17543, N11161, N12664);
and AND3_12039 (N17672, N17573, N12653, N12664);
and AND3_12040 (N17673, N17549, N11161, N12664);
and AND3_12041 (N17674, N17555, N12728, N12739);
and AND3_12042 (N17675, N17531, N11223, N12739);
and AND3_12043 (N17676, N17561, N12728, N12739);
and AND3_12044 (N17677, N17537, N11223, N12739);
and AND3_12045 (N17678, N17567, N12728, N12739);
and AND3_12046 (N17679, N17543, N11223, N12739);
and AND3_12047 (N17680, N17573, N12728, N12739);
and AND3_12048 (N17681, N17549, N11223, N12739);
and AND3_12049 (N17682, N17573, N13075, N13086);
and AND3_12050 (N17683, N17549, N11731, N13086);
and AND3_12051 (N17684, N17573, N13041, N13052);
and AND3_12052 (N17685, N17549, N11697, N13052);
and AND3_12053 (N17686, N17567, N13041, N13052);
and AND3_12054 (N17687, N17543, N11697, N13052);
and AND3_12055 (N17688, N17561, N13041, N13052);
and AND3_12056 (N17689, N17537, N11697, N13052);
and AND3_12057 (N17690, N17555, N13041, N13052);
and AND3_12058 (N17691, N17531, N11697, N13052);
and AND3_12059 (N17692, N17567, N13075, N13086);
and AND3_12060 (N17693, N17543, N11731, N13086);
and AND3_12061 (N17694, N17561, N13075, N13086);
and AND3_12062 (N17695, N17537, N11731, N13086);
and AND3_12063 (N17696, N17555, N13075, N13086);
and AND3_12064 (N17697, N17531, N11731, N13086);
or OR2_12065 (N17698, N17624, N17625);
not NOT1_12066 (N17699, N17573);
not NOT1_12067 (N17700, N17567);
not NOT1_12068 (N17701, N17561);
not NOT1_12069 (N17702, N17555);
and AND3_12070 (N17703, N11156, N17631, N1245);
not NOT1_12071 (N17704, N17549);
not NOT1_12072 (N17705, N17543);
not NOT1_12073 (N17706, N17537);
not NOT1_12074 (N17707, N17531);
not NOT1_12075 (N17708, N17579);
nand NAND2_12076 (N17709, N17579, N16739);
not NOT1_12077 (N17710, N17582);
nand NAND2_12078 (N17711, N17582, N16744);
nand NAND2_12079 (N17712, N17657, N17586);
nand NAND2_12080 (N17715, N17658, N17588);
not NOT1_12081 (N17718, N17589);
nand NAND2_12082 (N17719, N17589, N16772);
not NOT1_12083 (N17720, N17592);
nand NAND2_12084 (N17721, N17592, N16776);
not NOT1_12085 (N17722, N17595);
nand NAND2_12086 (N17723, N17595, N15733);
nand NAND2_12087 (N17724, N17665, N17599);
or OR4_12088 (N17727, N17666, N17667, N13617, N12586);
or OR4_12089 (N17728, N17668, N17669, N13618, N12587);
or OR4_12090 (N17729, N17670, N17671, N13619, N12588);
or OR4_12091 (N17730, N17672, N17673, N13620, N12589);
or OR4_12092 (N17731, N17674, N17675, N13628, N12596);
or OR4_12093 (N17732, N17676, N17677, N13629, N12597);
or OR4_12094 (N17733, N17678, N17679, N13630, N12598);
or OR4_12095 (N17734, N17680, N17681, N13631, N12599);
or OR4_12096 (N17735, N17682, N17683, N13638, N12604);
or OR4_12097 (N17736, N17684, N17685, N13642, N12606);
or OR4_12098 (N17737, N17686, N17687, N13643, N12607);
or OR4_12099 (N17738, N17688, N17689, N13644, N12608);
or OR4_12100 (N17739, N17690, N17691, N13645, N12609);
or OR4_12101 (N17740, N17692, N17693, N13651, N12615);
or OR4_12102 (N17741, N17694, N17695, N13652, N12616);
or OR4_12103 (N17742, N17696, N17697, N13653, N12617);
nand NAND2_12104 (N17743, N16271, N17708);
nand NAND2_12105 (N17744, N16283, N17710);
nand NAND2_12106 (N17749, N16341, N17718);
nand NAND2_12107 (N17750, N16347, N17720);
nand NAND2_12108 (N17751, N15214, N17722);
and AND2_12109 (N17754, N17727, N12647);
and AND2_12110 (N17755, N17728, N12647);
and AND2_12111 (N17756, N17729, N12647);
and AND2_12112 (N17757, N17730, N12647);
and AND2_12113 (N17758, N17731, N12722);
and AND2_12114 (N17759, N17732, N12722);
and AND2_12115 (N17760, N17733, N12722);
and AND2_12116 (N17761, N17734, N12722);
nand NAND2_12117 (N17762, N17743, N17709);
nand NAND2_12118 (N17765, N17744, N17711);
not NOT1_12119 (N17768, N17712);
nand NAND2_12120 (N17769, N17712, N16751);
not NOT1_12121 (N17770, N17715);
nand NAND2_12122 (N17771, N17715, N16760);
nand NAND2_12123 (N17772, N17749, N17719);
nand NAND2_12124 (N17775, N17750, N17721);
nand NAND2_12125 (N17778, N17751, N17723);
not NOT1_12126 (N17781, N17724);
nand NAND2_12127 (N17782, N17724, N15735);
nand NAND2_12128 (N17787, N16295, N17768);
nand NAND2_12129 (N17788, N16313, N17770);
nand NAND2_12130 (N17795, N15220, N17781);
not NOT1_12131 (N17796, N17762);
nand NAND2_12132 (N17797, N17762, N16740);
not NOT1_12133 (N17798, N17765);
nand NAND2_12134 (N17799, N17765, N16745);
nand NAND2_12135 (N17800, N17787, N17769);
nand NAND2_12136 (N17803, N17788, N17771);
not NOT1_12137 (N17806, N17772);
nand NAND2_12138 (N17807, N17772, N16773);
not NOT1_12139 (N17808, N17775);
nand NAND2_12140 (N17809, N17775, N16777);
not NOT1_12141 (N17810, N17778);
nand NAND2_12142 (N17811, N17778, N16782);
nand NAND2_12143 (N17812, N17795, N17782);
nand NAND2_12144 (N17815, N16274, N17796);
nand NAND2_12145 (N17816, N16286, N17798);
nand NAND2_12146 (N17821, N16344, N17806);
nand NAND2_12147 (N17822, N16350, N17808);
nand NAND2_12148 (N17823, N16353, N17810);
nand NAND2_12149 (N17826, N17815, N17797);
nand NAND2_12150 (N17829, N17816, N17799);
not NOT1_12151 (N17832, N17800);
nand NAND2_12152 (N17833, N17800, N16752);
not NOT1_12153 (N17834, N17803);
nand NAND2_12154 (N17835, N17803, N16761);
nand NAND2_12155 (N17836, N17821, N17807);
nand NAND2_12156 (N17839, N17822, N17809);
nand NAND2_12157 (N17842, N17823, N17811);
not NOT1_12158 (N17845, N17812);
nand NAND2_12159 (N17846, N17812, N16790);
nand NAND2_12160 (N17851, N16298, N17832);
nand NAND2_12161 (N17852, N16316, N17834);
nand NAND2_12162 (N17859, N16364, N17845);
not NOT1_12163 (N17860, N17826);
nand NAND2_12164 (N17861, N17826, N16741);
not NOT1_12165 (N17862, N17829);
nand NAND2_12166 (N17863, N17829, N16746);
nand NAND2_12167 (N17864, N17851, N17833);
nand NAND2_12168 (N17867, N17852, N17835);
not NOT1_12169 (N17870, N17836);
nand NAND2_12170 (N17871, N17836, N15730);
not NOT1_12171 (N17872, N17839);
nand NAND2_12172 (N17873, N17839, N15732);
not NOT1_12173 (N17874, N17842);
nand NAND2_12174 (N17875, N17842, N16783);
nand NAND2_12175 (N17876, N17859, N17846);
nand NAND2_12176 (N17879, N16277, N17860);
nand NAND2_12177 (N17880, N16289, N17862);
nand NAND2_12178 (N17885, N15199, N17870);
nand NAND2_12179 (N17886, N15208, N17872);
nand NAND2_12180 (N17887, N16356, N17874);
nand NAND2_12181 (N17890, N17879, N17861);
nand NAND2_12182 (N17893, N17880, N17863);
not NOT1_12183 (N17896, N17864);
nand NAND2_12184 (N17897, N17864, N16753);
not NOT1_12185 (N17898, N17867);
nand NAND2_12186 (N17899, N17867, N16762);
nand NAND2_12187 (N17900, N17885, N17871);
nand NAND2_12188 (N17903, N17886, N17873);
nand NAND2_12189 (N17906, N17887, N17875);
not NOT1_12190 (N17909, N17876);
nand NAND2_12191 (N17910, N17876, N16791);
nand NAND2_12192 (N17917, N16301, N17896);
nand NAND2_12193 (N17918, N16319, N17898);
nand NAND2_12194 (N17923, N16367, N17909);
not NOT1_12195 (N17924, N17890);
nand NAND2_12196 (N17925, N17890, N16680);
not NOT1_12197 (N17926, N17893);
nand NAND2_12198 (N17927, N17893, N16681);
not NOT1_12199 (N17928, N17900);
nand NAND2_12200 (N17929, N17900, N15690);
not NOT1_12201 (N17930, N17903);
nand NAND2_12202 (N17931, N17903, N15691);
nand NAND2_12203 (N17932, N17917, N17897);
nand NAND2_12204 (N17935, N17918, N17899);
not NOT1_12205 (N17938, N17906);
nand NAND2_12206 (N17939, N17906, N16784);
nand NAND2_12207 (N17940, N17923, N17910);
nand NAND2_12208 (N17943, N16280, N17924);
nand NAND2_12209 (N17944, N16292, N17926);
nand NAND2_12210 (N17945, N15202, N17928);
nand NAND2_12211 (N17946, N15211, N17930);
nand NAND2_12212 (N17951, N16359, N17938);
nand NAND2_12213 (N17954, N17943, N17925);
nand NAND2_12214 (N17957, N17944, N17927);
nand NAND2_12215 (N17960, N17945, N17929);
nand NAND2_12216 (N17963, N17946, N17931);
not NOT1_12217 (N17966, N17932);
nand NAND2_12218 (N17967, N17932, N16754);
not NOT1_12219 (N17968, N17935);
nand NAND2_12220 (N17969, N17935, N16755);
nand NAND2_12221 (N17970, N17951, N17939);
not NOT1_12222 (N17973, N17940);
nand NAND2_12223 (N17974, N17940, N16785);
nand NAND2_12224 (N17984, N16304, N17966);
nand NAND2_12225 (N17985, N16322, N17968);
nand NAND2_12226 (N17987, N16370, N17973);
and AND3_12227 (N17988, N17957, N16831, N11157);
and AND3_12228 (N17989, N17954, N16415, N11157);
and AND3_12229 (N17990, N17957, N17041, N1566);
and AND3_12230 (N17991, N17954, N17177, N1566);
not NOT1_12231 (N17992, N17970);
nand NAND2_12232 (N17993, N17970, N16448);
and AND3_12233 (N17994, N17963, N16857, N11219);
and AND3_12234 (N17995, N17960, N16441, N11219);
and AND3_12235 (N17996, N17963, N17065, N1583);
and AND3_12236 (N17997, N17960, N17182, N1583);
nand NAND2_12237 (N17998, N17984, N17967);
nand NAND2_12238 (N18001, N17985, N17969);
nand NAND2_12239 (N18004, N17987, N17974);
nand NAND2_12240 (N18009, N16051, N17992);
or OR4_12241 (N18013, N17988, N17989, N17990, N17991);
or OR4_12242 (N18017, N17994, N17995, N17996, N17997);
not NOT1_12243 (N18020, N17998);
nand NAND2_12244 (N18021, N17998, N16682);
not NOT1_12245 (N18022, N18001);
nand NAND2_12246 (N18023, N18001, N16683);
nand NAND2_12247 (N18025, N18009, N17993);
not NOT1_12248 (N18026, N18004);
nand NAND2_12249 (N18027, N18004, N16449);
nand NAND2_12250 (N18031, N16307, N18020);
nand NAND2_12251 (N18032, N16310, N18022);
not NOT1_12252 (N18033, N18013);
nand NAND2_12253 (N18034, N16054, N18026);
and AND2_12254 (N18035, N1583, N18025);
not NOT1_12255 (N18036, N18017);
nand NAND2_12256 (N18037, N18031, N18021);
nand NAND2_12257 (N18038, N18032, N18023);
nand NAND2_12258 (N18039, N18034, N18027);
not NOT1_12259 (N18040, N18038);
and AND2_12260 (N18041, N1566, N18037);
not NOT1_12261 (N18042, N18039);
and AND2_12262 (N18043, N18040, N11157);
and AND2_12263 (N18044, N18042, N11219);
or OR2_12264 (N18045, N18043, N18041);
or OR2_12265 (N18048, N18044, N18035);
nand NAND2_12266 (N18055, N18045, N18033);
not NOT1_12267 (N18056, N18045);
nand NAND2_12268 (N18057, N18048, N18036);
not NOT1_12269 (N18058, N18048);
nand NAND2_12270 (N18059, N18013, N18056);
nand NAND2_12271 (N18060, N18017, N18058);
nand NAND2_12272 (N18061, N18055, N18059);
nand NAND2_12273 (N18064, N18057, N18060);
and AND3_12274 (N18071, N18064, N11777, N13130);
and AND3_12275 (N18072, N18061, N11761, N13108);
not NOT1_12276 (N18073, N18061);
not NOT1_12277 (N18074, N18064);
or OR4_12278 (N18075, N17526, N18071, N13659, N12625);
or OR4_12279 (N18076, N17636, N18072, N13661, N12627);
and AND2_12280 (N18077, N18073, N11727);
and AND2_12281 (N18078, N18074, N11727);
or OR2_12282 (N18079, N17530, N18077);
or OR2_12283 (N18082, N17479, N18078);
and AND2_12284 (N18089, N18079, N13063);
and AND2_12285 (N18090, N18082, N13063);
and AND2_12286 (N18091, N18079, N13063);
and AND2_12287 (N18092, N18082, N13063);
or OR2_12288 (N18093, N18089, N13071);
or OR2_12289 (N18096, N18090, N13072);
or OR2_12290 (N18099, N18091, N13073);
or OR2_12291 (N18102, N18092, N13074);
and AND3_12292 (N18113, N18102, N12779, N12790);
and AND3_12293 (N18114, N18099, N11327, N12790);
and AND3_12294 (N18115, N18102, N12801, N12812);
and AND3_12295 (N18116, N18099, N11351, N12812);
and AND3_12296 (N18117, N18096, N12681, N12692);
and AND3_12297 (N18118, N18093, N11185, N12692);
and AND3_12298 (N18119, N18096, N12756, N12767);
and AND3_12299 (N18120, N18093, N11247, N12767);
or OR4_12300 (N18121, N18117, N18118, N13662, N12703);
or OR4_12301 (N18122, N18119, N18120, N13663, N12778);
or OR4_12302 (N18123, N18113, N18114, N13650, N12614);
or OR4_12303 (N18124, N18115, N18116, N13658, N12622);
and AND2_12304 (N18125, N18121, N12675);
and AND2_12305 (N18126, N18122, N12750);
not NOT1_12306 (N18127, N18125);
not NOT1_12307 (N18128, N18126);

buf BUFF1_21 (N2709, N2141);
buf BUFF1_22 (N2816, N2293);
and AND2_23 (N21042, N2135, N2631);
not NOT1_24 (N21043, N2591);
buf BUFF1_25 (N21066, N2592);
not NOT1_26 (N21067, N2595);
not NOT1_27 (N21080, N2596);
not NOT1_28 (N21092, N2597);
not NOT1_29 (N21104, N2598);
not NOT1_210 (N21137, N2545);
not NOT1_211 (N21138, N2348);
not NOT1_212 (N21139, N2366);
and AND2_213 (N21140, N2552, N2562);
not NOT1_214 (N21141, N2549);
not NOT1_215 (N21142, N2545);
not NOT1_216 (N21143, N2545);
not NOT1_217 (N21144, N2338);
not NOT1_218 (N21145, N2358);
nand NAND2_219 (N21146, N2373, N21);
and AND2_220 (N21147, N2141, N2145);
not NOT1_221 (N21148, N2592);
not NOT1_222 (N21149, N21042);
and AND2_223 (N21150, N21043, N227);
and AND2_224 (N21151, N2386, N2556);
not NOT1_225 (N21152, N2245);
not NOT1_226 (N21153, N2552);
not NOT1_227 (N21154, N2562);
not NOT1_228 (N21155, N2559);
and AND4_229 (N21156, N2386, N2559, N2556, N2552);
not NOT1_230 (N21157, N2566);
buf BUFF1_231 (N21161, N2571);
buf BUFF1_232 (N21173, N2574);
buf BUFF1_233 (N21185, N2571);
buf BUFF1_234 (N21197, N2574);
buf BUFF1_235 (N21209, N2137);
buf BUFF1_236 (N21213, N2137);
buf BUFF1_237 (N21216, N2141);
not NOT1_238 (N21219, N2583);
buf BUFF1_239 (N21223, N2577);
buf BUFF1_240 (N21235, N2580);
buf BUFF1_241 (N21247, N2577);
buf BUFF1_242 (N21259, N2580);
buf BUFF1_243 (N21271, N2254);
buf BUFF1_244 (N21280, N2251);
buf BUFF1_245 (N21292, N2251);
buf BUFF1_246 (N21303, N2248);
buf BUFF1_247 (N21315, N2248);
buf BUFF1_248 (N21327, N2610);
buf BUFF1_249 (N21339, N2607);
buf BUFF1_250 (N21351, N2613);
buf BUFF1_251 (N21363, N2616);
buf BUFF1_252 (N21375, N2210);
buf BUFF1_253 (N21378, N2210);
buf BUFF1_254 (N21381, N2218);
buf BUFF1_255 (N21384, N2218);
buf BUFF1_256 (N21387, N2226);
buf BUFF1_257 (N21390, N2226);
buf BUFF1_258 (N21393, N2234);
buf BUFF1_259 (N21396, N2234);
buf BUFF1_260 (N21415, N2257);
buf BUFF1_261 (N21418, N2257);
buf BUFF1_262 (N21421, N2265);
buf BUFF1_263 (N21424, N2265);
buf BUFF1_264 (N21427, N2273);
buf BUFF1_265 (N21430, N2273);
buf BUFF1_266 (N21433, N2281);
buf BUFF1_267 (N21436, N2281);
buf BUFF1_268 (N21455, N2335);
buf BUFF1_269 (N21462, N2335);
buf BUFF1_270 (N21469, N2206);
and AND2_271 (N21475, N227, N231);
buf BUFF1_272 (N21479, N21);
buf BUFF1_273 (N21482, N2588);
buf BUFF1_274 (N21492, N2293);
buf BUFF1_275 (N21495, N2302);
buf BUFF1_276 (N21498, N2308);
buf BUFF1_277 (N21501, N2308);
buf BUFF1_278 (N21504, N2316);
buf BUFF1_279 (N21507, N2316);
buf BUFF1_280 (N21510, N2324);
buf BUFF1_281 (N21513, N2324);
buf BUFF1_282 (N21516, N2341);
buf BUFF1_283 (N21519, N2341);
buf BUFF1_284 (N21522, N2351);
buf BUFF1_285 (N21525, N2351);
buf BUFF1_286 (N21542, N2257);
buf BUFF1_287 (N21545, N2257);
buf BUFF1_288 (N21548, N2265);
buf BUFF1_289 (N21551, N2265);
buf BUFF1_290 (N21554, N2273);
buf BUFF1_291 (N21557, N2273);
buf BUFF1_292 (N21560, N2281);
buf BUFF1_293 (N21563, N2281);
buf BUFF1_294 (N21566, N2332);
buf BUFF1_295 (N21573, N2332);
buf BUFF1_296 (N21580, N2549);
and AND2_297 (N21583, N231, N227);
not NOT1_298 (N21588, N2588);
buf BUFF1_299 (N21594, N2324);
buf BUFF1_2100 (N21597, N2324);
buf BUFF1_2101 (N21600, N2341);
buf BUFF1_2102 (N21603, N2341);
buf BUFF1_2103 (N21606, N2351);
buf BUFF1_2104 (N21609, N2351);
buf BUFF1_2105 (N21612, N2293);
buf BUFF1_2106 (N21615, N2302);
buf BUFF1_2107 (N21618, N2308);
buf BUFF1_2108 (N21621, N2308);
buf BUFF1_2109 (N21624, N2316);
buf BUFF1_2110 (N21627, N2316);
buf BUFF1_2111 (N21630, N2361);
buf BUFF1_2112 (N21633, N2361);
buf BUFF1_2113 (N21636, N2210);
buf BUFF1_2114 (N21639, N2210);
buf BUFF1_2115 (N21642, N2218);
buf BUFF1_2116 (N21645, N2218);
buf BUFF1_2117 (N21648, N2226);
buf BUFF1_2118 (N21651, N2226);
buf BUFF1_2119 (N21654, N2234);
buf BUFF1_2120 (N21657, N2234);
not NOT1_2121 (N21660, N2324);
buf BUFF1_2122 (N21663, N2242);
buf BUFF1_2123 (N21675, N2242);
buf BUFF1_2124 (N21685, N2254);
buf BUFF1_2125 (N21697, N2610);
buf BUFF1_2126 (N21709, N2607);
buf BUFF1_2127 (N21721, N2625);
buf BUFF1_2128 (N21727, N2619);
buf BUFF1_2129 (N21731, N2613);
buf BUFF1_2130 (N21743, N2616);
not NOT1_2131 (N21755, N2599);
not NOT1_2132 (N21758, N2603);
buf BUFF1_2133 (N21761, N2619);
buf BUFF1_2134 (N21769, N2625);
buf BUFF1_2135 (N21777, N2619);
buf BUFF1_2136 (N21785, N2625);
buf BUFF1_2137 (N21793, N2619);
buf BUFF1_2138 (N21800, N2625);
buf BUFF1_2139 (N21807, N2619);
buf BUFF1_2140 (N21814, N2625);
buf BUFF1_2141 (N21821, N2299);
buf BUFF1_2142 (N21824, N2446);
buf BUFF1_2143 (N21827, N2457);
buf BUFF1_2144 (N21830, N2468);
buf BUFF1_2145 (N21833, N2422);
buf BUFF1_2146 (N21836, N2435);
buf BUFF1_2147 (N21839, N2389);
buf BUFF1_2148 (N21842, N2400);
buf BUFF1_2149 (N21845, N2411);
buf BUFF1_2150 (N21848, N2374);
buf BUFF1_2151 (N21851, N24);
buf BUFF1_2152 (N21854, N2446);
buf BUFF1_2153 (N21857, N2457);
buf BUFF1_2154 (N21860, N2468);
buf BUFF1_2155 (N21863, N2435);
buf BUFF1_2156 (N21866, N2389);
buf BUFF1_2157 (N21869, N2400);
buf BUFF1_2158 (N21872, N2411);
buf BUFF1_2159 (N21875, N2422);
buf BUFF1_2160 (N21878, N2374);
buf BUFF1_2161 (N21881, N2479);
buf BUFF1_2162 (N21884, N2490);
buf BUFF1_2163 (N21887, N2503);
buf BUFF1_2164 (N21890, N2514);
buf BUFF1_2165 (N21893, N2523);
buf BUFF1_2166 (N21896, N2534);
buf BUFF1_2167 (N21899, N254);
buf BUFF1_2168 (N21902, N2479);
buf BUFF1_2169 (N21905, N2503);
buf BUFF1_2170 (N21908, N2514);
buf BUFF1_2171 (N21911, N2523);
buf BUFF1_2172 (N21914, N2534);
buf BUFF1_2173 (N21917, N2490);
buf BUFF1_2174 (N21920, N2361);
buf BUFF1_2175 (N21923, N2369);
buf BUFF1_2176 (N21926, N2341);
buf BUFF1_2177 (N21929, N2351);
buf BUFF1_2178 (N21932, N2308);
buf BUFF1_2179 (N21935, N2316);
buf BUFF1_2180 (N21938, N2293);
buf BUFF1_2181 (N21941, N2302);
buf BUFF1_2182 (N21944, N2281);
buf BUFF1_2183 (N21947, N2289);
buf BUFF1_2184 (N21950, N2265);
buf BUFF1_2185 (N21953, N2273);
buf BUFF1_2186 (N21956, N2234);
buf BUFF1_2187 (N21959, N2257);
buf BUFF1_2188 (N21962, N2218);
buf BUFF1_2189 (N21965, N2226);
buf BUFF1_2190 (N21968, N2210);
not NOT1_2191 (N21972, N21146);
and AND2_2192 (N22054, N2136, N21148);
not NOT1_2193 (N22060, N21150);
not NOT1_2194 (N22061, N21151);
buf BUFF1_2195 (N22139, N21209);
buf BUFF1_2196 (N22142, N21216);
buf BUFF1_2197 (N22309, N21479);
and AND2_2198 (N22349, N21104, N2514);
or OR2_2199 (N22350, N21067, N2514);
buf BUFF1_2200 (N22387, N21580);
buf BUFF1_2201 (N22527, N21821);
not NOT1_2202 (N22584, N21580);
and AND3_2203 (N22585, N2170, N21161, N21173);
and AND3_2204 (N22586, N2173, N21161, N21173);
and AND3_2205 (N22587, N2167, N21161, N21173);
and AND3_2206 (N22588, N2164, N21161, N21173);
and AND3_2207 (N22589, N2161, N21161, N21173);
nand NAND2_2208 (N22590, N21475, N2140);
and AND3_2209 (N22591, N2185, N21185, N21197);
and AND3_2210 (N22592, N2158, N21185, N21197);
and AND3_2211 (N22593, N2152, N21185, N21197);
and AND3_2212 (N22594, N2146, N21185, N21197);
and AND3_2213 (N22595, N2170, N21223, N21235);
and AND3_2214 (N22596, N2173, N21223, N21235);
and AND3_2215 (N22597, N2167, N21223, N21235);
and AND3_2216 (N22598, N2164, N21223, N21235);
and AND3_2217 (N22599, N2161, N21223, N21235);
and AND3_2218 (N22600, N2185, N21247, N21259);
and AND3_2219 (N22601, N2158, N21247, N21259);
and AND3_2220 (N22602, N2152, N21247, N21259);
and AND3_2221 (N22603, N2146, N21247, N21259);
and AND3_2222 (N22604, N2106, N21731, N21743);
and AND3_2223 (N22605, N261, N21327, N21339);
and AND3_2224 (N22606, N2106, N21697, N21709);
and AND3_2225 (N22607, N249, N21697, N21709);
and AND3_2226 (N22608, N2103, N21697, N21709);
and AND3_2227 (N22609, N240, N21697, N21709);
and AND3_2228 (N22610, N237, N21697, N21709);
and AND3_2229 (N22611, N220, N21327, N21339);
and AND3_2230 (N22612, N217, N21327, N21339);
and AND3_2231 (N22613, N270, N21327, N21339);
and AND3_2232 (N22614, N264, N21327, N21339);
and AND3_2233 (N22615, N249, N21731, N21743);
and AND3_2234 (N22616, N2103, N21731, N21743);
and AND3_2235 (N22617, N240, N21731, N21743);
and AND3_2236 (N22618, N237, N21731, N21743);
and AND3_2237 (N22619, N220, N21351, N21363);
and AND3_2238 (N22620, N217, N21351, N21363);
and AND3_2239 (N22621, N270, N21351, N21363);
and AND3_2240 (N22622, N264, N21351, N21363);
not NOT1_2241 (N22623, N21475);
and AND3_2242 (N22624, N2123, N21758, N2599);
and AND2_2243 (N22625, N21777, N21785);
and AND3_2244 (N22626, N261, N21351, N21363);
and AND2_2245 (N22627, N21761, N21769);
not NOT1_2246 (N22628, N21824);
not NOT1_2247 (N22629, N21827);
not NOT1_2248 (N22630, N21830);
not NOT1_2249 (N22631, N21833);
not NOT1_2250 (N22632, N21836);
not NOT1_2251 (N22633, N21839);
not NOT1_2252 (N22634, N21842);
not NOT1_2253 (N22635, N21845);
not NOT1_2254 (N22636, N21848);
not NOT1_2255 (N22637, N21851);
not NOT1_2256 (N22638, N21854);
not NOT1_2257 (N22639, N21857);
not NOT1_2258 (N22640, N21860);
not NOT1_2259 (N22641, N21863);
not NOT1_2260 (N22642, N21866);
not NOT1_2261 (N22643, N21869);
not NOT1_2262 (N22644, N21872);
not NOT1_2263 (N22645, N21875);
not NOT1_2264 (N22646, N21878);
buf BUFF1_2265 (N22647, N21209);
not NOT1_2266 (N22653, N21161);
not NOT1_2267 (N22664, N21173);
buf BUFF1_2268 (N22675, N21209);
not NOT1_2269 (N22681, N21185);
not NOT1_2270 (N22692, N21197);
and AND3_2271 (N22703, N2179, N21185, N21197);
buf BUFF1_2272 (N22704, N21479);
not NOT1_2273 (N22709, N21881);
not NOT1_2274 (N22710, N21884);
not NOT1_2275 (N22711, N21887);
not NOT1_2276 (N22712, N21890);
not NOT1_2277 (N22713, N21893);
not NOT1_2278 (N22714, N21896);
not NOT1_2279 (N22715, N21899);
not NOT1_2280 (N22716, N21902);
not NOT1_2281 (N22717, N21905);
not NOT1_2282 (N22718, N21908);
not NOT1_2283 (N22719, N21911);
not NOT1_2284 (N22720, N21914);
not NOT1_2285 (N22721, N21917);
buf BUFF1_2286 (N22722, N21213);
not NOT1_2287 (N22728, N21223);
not NOT1_2288 (N22739, N21235);
buf BUFF1_2289 (N22750, N21213);
not NOT1_2290 (N22756, N21247);
not NOT1_2291 (N22767, N21259);
and AND3_2292 (N22778, N2179, N21247, N21259);
not NOT1_2293 (N22779, N21327);
not NOT1_2294 (N22790, N21339);
not NOT1_2295 (N22801, N21351);
not NOT1_2296 (N22812, N21363);
not NOT1_2297 (N22823, N21375);
not NOT1_2298 (N22824, N21378);
not NOT1_2299 (N22825, N21381);
not NOT1_2300 (N22826, N21384);
not NOT1_2301 (N22827, N21387);
not NOT1_2302 (N22828, N21390);
not NOT1_2303 (N22829, N21393);
not NOT1_2304 (N22830, N21396);
and AND3_2305 (N22831, N21104, N2457, N21378);
and AND3_2306 (N22832, N21104, N2468, N21384);
and AND3_2307 (N22833, N21104, N2422, N21390);
and AND3_2308 (N22834, N21104, N2435, N21396);
and AND2_2309 (N22835, N21067, N21375);
and AND2_2310 (N22836, N21067, N21381);
and AND2_2311 (N22837, N21067, N21387);
and AND2_2312 (N22838, N21067, N21393);
not NOT1_2313 (N22839, N21415);
not NOT1_2314 (N22840, N21418);
not NOT1_2315 (N22841, N21421);
not NOT1_2316 (N22842, N21424);
not NOT1_2317 (N22843, N21427);
not NOT1_2318 (N22844, N21430);
not NOT1_2319 (N22845, N21433);
not NOT1_2320 (N22846, N21436);
and AND3_2321 (N22847, N21104, N2389, N21418);
and AND3_2322 (N22848, N21104, N2400, N21424);
and AND3_2323 (N22849, N21104, N2411, N21430);
and AND3_2324 (N22850, N21104, N2374, N21436);
and AND2_2325 (N22851, N21067, N21415);
and AND2_2326 (N22852, N21067, N21421);
and AND2_2327 (N22853, N21067, N21427);
and AND2_2328 (N22854, N21067, N21433);
not NOT1_2329 (N22855, N21455);
not NOT1_2330 (N22861, N21462);
and AND2_2331 (N22867, N2292, N21455);
and AND2_2332 (N22868, N2288, N21455);
and AND2_2333 (N22869, N2280, N21455);
and AND2_2334 (N22870, N2272, N21455);
and AND2_2335 (N22871, N2264, N21455);
and AND2_2336 (N22872, N2241, N21462);
and AND2_2337 (N22873, N2233, N21462);
and AND2_2338 (N22874, N2225, N21462);
and AND2_2339 (N22875, N2217, N21462);
and AND2_2340 (N22876, N2209, N21462);
buf BUFF1_2341 (N22877, N21216);
not NOT1_2342 (N22882, N21482);
not NOT1_2343 (N22891, N21475);
not NOT1_2344 (N22901, N21492);
not NOT1_2345 (N22902, N21495);
not NOT1_2346 (N22903, N21498);
not NOT1_2347 (N22904, N21501);
not NOT1_2348 (N22905, N21504);
not NOT1_2349 (N22906, N21507);
and AND2_2350 (N22907, N21303, N21495);
and AND3_2351 (N22908, N21303, N2479, N21501);
and AND3_2352 (N22909, N21303, N2490, N21507);
and AND2_2353 (N22910, N21663, N21492);
and AND2_2354 (N22911, N21663, N21498);
and AND2_2355 (N22912, N21663, N21504);
not NOT1_2356 (N22913, N21510);
not NOT1_2357 (N22914, N21513);
not NOT1_2358 (N22915, N21516);
not NOT1_2359 (N22916, N21519);
not NOT1_2360 (N22917, N21522);
not NOT1_2361 (N22918, N21525);
and AND3_2362 (N22919, N21104, N2503, N21513);
not NOT1_2363 (N22920, N22349);
and AND3_2364 (N22921, N21104, N2523, N21519);
and AND3_2365 (N22922, N21104, N2534, N21525);
and AND2_2366 (N22923, N21067, N21510);
and AND2_2367 (N22924, N21067, N21516);
and AND2_2368 (N22925, N21067, N21522);
not NOT1_2369 (N22926, N21542);
not NOT1_2370 (N22927, N21545);
not NOT1_2371 (N22928, N21548);
not NOT1_2372 (N22929, N21551);
not NOT1_2373 (N22930, N21554);
not NOT1_2374 (N22931, N21557);
not NOT1_2375 (N22932, N21560);
not NOT1_2376 (N22933, N21563);
and AND3_2377 (N22934, N21303, N2389, N21545);
and AND3_2378 (N22935, N21303, N2400, N21551);
and AND3_2379 (N22936, N21303, N2411, N21557);
and AND3_2380 (N22937, N21303, N2374, N21563);
and AND2_2381 (N22938, N21663, N21542);
and AND2_2382 (N22939, N21663, N21548);
and AND2_2383 (N22940, N21663, N21554);
and AND2_2384 (N22941, N21663, N21560);
not NOT1_2385 (N22942, N21566);
not NOT1_2386 (N22948, N21573);
and AND2_2387 (N22954, N2372, N21566);
and AND2_2388 (N22955, N2366, N21566);
and AND2_2389 (N22956, N2358, N21566);
and AND2_2390 (N22957, N2348, N21566);
and AND2_2391 (N22958, N2338, N21566);
and AND2_2392 (N22959, N2331, N21573);
and AND2_2393 (N22960, N2323, N21573);
and AND2_2394 (N22961, N2315, N21573);
and AND2_2395 (N22962, N2307, N21573);
and AND2_2396 (N22963, N2299, N21573);
not NOT1_2397 (N22964, N21588);
and AND2_2398 (N22969, N283, N21588);
and AND2_2399 (N22970, N286, N21588);
and AND2_2400 (N22971, N288, N21588);
and AND2_2401 (N22972, N288, N21588);
not NOT1_2402 (N22973, N21594);
not NOT1_2403 (N22974, N21597);
not NOT1_2404 (N22975, N21600);
not NOT1_2405 (N22976, N21603);
not NOT1_2406 (N22977, N21606);
not NOT1_2407 (N22978, N21609);
and AND3_2408 (N22979, N21315, N2503, N21597);
and AND2_2409 (N22980, N21315, N2514);
and AND3_2410 (N22981, N21315, N2523, N21603);
and AND3_2411 (N22982, N21315, N2534, N21609);
and AND2_2412 (N22983, N21675, N21594);
or OR2_2413 (N22984, N21675, N2514);
and AND2_2414 (N22985, N21675, N21600);
and AND2_2415 (N22986, N21675, N21606);
not NOT1_2416 (N22987, N21612);
not NOT1_2417 (N22988, N21615);
not NOT1_2418 (N22989, N21618);
not NOT1_2419 (N22990, N21621);
not NOT1_2420 (N22991, N21624);
not NOT1_2421 (N22992, N21627);
and AND2_2422 (N22993, N21315, N21615);
and AND3_2423 (N22994, N21315, N2479, N21621);
and AND3_2424 (N22995, N21315, N2490, N21627);
and AND2_2425 (N22996, N21675, N21612);
and AND2_2426 (N22997, N21675, N21618);
and AND2_2427 (N22998, N21675, N21624);
not NOT1_2428 (N22999, N21630);
buf BUFF1_2429 (N23000, N21469);
buf BUFF1_2430 (N23003, N21469);
not NOT1_2431 (N23006, N21633);
buf BUFF1_2432 (N23007, N21469);
buf BUFF1_2433 (N23010, N21469);
and AND2_2434 (N23013, N21315, N21630);
and AND2_2435 (N23014, N21315, N21633);
not NOT1_2436 (N23015, N21636);
not NOT1_2437 (N23016, N21639);
not NOT1_2438 (N23017, N21642);
not NOT1_2439 (N23018, N21645);
not NOT1_2440 (N23019, N21648);
not NOT1_2441 (N23020, N21651);
not NOT1_2442 (N23021, N21654);
not NOT1_2443 (N23022, N21657);
and AND3_2444 (N23023, N21303, N2457, N21639);
and AND3_2445 (N23024, N21303, N2468, N21645);
and AND3_2446 (N23025, N21303, N2422, N21651);
and AND3_2447 (N23026, N21303, N2435, N21657);
and AND2_2448 (N23027, N21663, N21636);
and AND2_2449 (N23028, N21663, N21642);
and AND2_2450 (N23029, N21663, N21648);
and AND2_2451 (N23030, N21663, N21654);
not NOT1_2452 (N23031, N21920);
not NOT1_2453 (N23032, N21923);
not NOT1_2454 (N23033, N21926);
not NOT1_2455 (N23034, N21929);
buf BUFF1_2456 (N23035, N21660);
buf BUFF1_2457 (N23038, N21660);
not NOT1_2458 (N23041, N21697);
not NOT1_2459 (N23052, N21709);
not NOT1_2460 (N23063, N21721);
not NOT1_2461 (N23068, N21727);
and AND2_2462 (N23071, N297, N21721);
and AND2_2463 (N23072, N294, N21721);
and AND2_2464 (N23073, N297, N21721);
and AND2_2465 (N23074, N294, N21721);
not NOT1_2466 (N23075, N21731);
not NOT1_2467 (N23086, N21743);
not NOT1_2468 (N23097, N21761);
not NOT1_2469 (N23108, N21769);
not NOT1_2470 (N23119, N21777);
not NOT1_2471 (N23130, N21785);
not NOT1_2472 (N23141, N21944);
not NOT1_2473 (N23142, N21947);
not NOT1_2474 (N23143, N21950);
not NOT1_2475 (N23144, N21953);
not NOT1_2476 (N23145, N21956);
not NOT1_2477 (N23146, N21959);
not NOT1_2478 (N23147, N21793);
not NOT1_2479 (N23158, N21800);
not NOT1_2480 (N23169, N21807);
not NOT1_2481 (N23180, N21814);
buf BUFF1_2482 (N23191, N21821);
not NOT1_2483 (N23194, N21932);
not NOT1_2484 (N23195, N21935);
not NOT1_2485 (N23196, N21938);
not NOT1_2486 (N23197, N21941);
not NOT1_2487 (N23198, N21962);
not NOT1_2488 (N23199, N21965);
buf BUFF1_2489 (N23200, N21469);
not NOT1_2490 (N23203, N21968);
buf BUFF1_2491 (N23357, N22704);
buf BUFF1_2492 (N23358, N22704);
buf BUFF1_2493 (N23359, N22704);
buf BUFF1_2494 (N23360, N22704);
and AND3_2495 (N23401, N2457, N21092, N22824);
and AND3_2496 (N23402, N2468, N21092, N22826);
and AND3_2497 (N23403, N2422, N21092, N22828);
and AND3_2498 (N23404, N2435, N21092, N22830);
and AND2_2499 (N23405, N21080, N22823);
and AND2_2500 (N23406, N21080, N22825);
and AND2_2501 (N23407, N21080, N22827);
and AND2_2502 (N23408, N21080, N22829);
and AND3_2503 (N23409, N2389, N21092, N22840);
and AND3_2504 (N23410, N2400, N21092, N22842);
and AND3_2505 (N23411, N2411, N21092, N22844);
and AND3_2506 (N23412, N2374, N21092, N22846);
and AND2_2507 (N23413, N21080, N22839);
and AND2_2508 (N23414, N21080, N22841);
and AND2_2509 (N23415, N21080, N22843);
and AND2_2510 (N23416, N21080, N22845);
and AND2_2511 (N23444, N21280, N22902);
and AND3_2512 (N23445, N2479, N21280, N22904);
and AND3_2513 (N23446, N2490, N21280, N22906);
and AND2_2514 (N23447, N21685, N22901);
and AND2_2515 (N23448, N21685, N22903);
and AND2_2516 (N23449, N21685, N22905);
and AND3_2517 (N23450, N2503, N21092, N22914);
and AND3_2518 (N23451, N2523, N21092, N22916);
and AND3_2519 (N23452, N2534, N21092, N22918);
and AND2_2520 (N23453, N21080, N22913);
and AND2_2521 (N23454, N21080, N22915);
and AND2_2522 (N23455, N21080, N22917);
and AND2_2523 (N23456, N22920, N22350);
and AND3_2524 (N23459, N2389, N21280, N22927);
and AND3_2525 (N23460, N2400, N21280, N22929);
and AND3_2526 (N23461, N2411, N21280, N22931);
and AND3_2527 (N23462, N2374, N21280, N22933);
and AND2_2528 (N23463, N21685, N22926);
and AND2_2529 (N23464, N21685, N22928);
and AND2_2530 (N23465, N21685, N22930);
and AND2_2531 (N23466, N21685, N22932);
and AND3_2532 (N23481, N2503, N21292, N22974);
not NOT1_2533 (N23482, N22980);
and AND3_2534 (N23483, N2523, N21292, N22976);
and AND3_2535 (N23484, N2534, N21292, N22978);
and AND2_2536 (N23485, N21271, N22973);
and AND2_2537 (N23486, N21271, N22975);
and AND2_2538 (N23487, N21271, N22977);
and AND2_2539 (N23488, N21292, N22988);
and AND3_2540 (N23489, N2479, N21292, N22990);
and AND3_2541 (N23490, N2490, N21292, N22992);
and AND2_2542 (N23491, N21271, N22987);
and AND2_2543 (N23492, N21271, N22989);
and AND2_2544 (N23493, N21271, N22991);
and AND2_2545 (N23502, N21292, N22999);
and AND2_2546 (N23503, N21292, N23006);
and AND3_2547 (N23504, N2457, N21280, N23016);
and AND3_2548 (N23505, N2468, N21280, N23018);
and AND3_2549 (N23506, N2422, N21280, N23020);
and AND3_2550 (N23507, N2435, N21280, N23022);
and AND2_2551 (N23508, N21685, N23015);
and AND2_2552 (N23509, N21685, N23017);
and AND2_2553 (N23510, N21685, N23019);
and AND2_2554 (N23511, N21685, N23021);
nand NAND2_2555 (N23512, N21923, N23031);
nand NAND2_2556 (N23513, N21920, N23032);
nand NAND2_2557 (N23514, N21929, N23033);
nand NAND2_2558 (N23515, N21926, N23034);
nand NAND2_2559 (N23558, N21947, N23141);
nand NAND2_2560 (N23559, N21944, N23142);
nand NAND2_2561 (N23560, N21953, N23143);
nand NAND2_2562 (N23561, N21950, N23144);
nand NAND2_2563 (N23562, N21959, N23145);
nand NAND2_2564 (N23563, N21956, N23146);
buf BUFF1_2565 (N23604, N23191);
nand NAND2_2566 (N23605, N21935, N23194);
nand NAND2_2567 (N23606, N21932, N23195);
nand NAND2_2568 (N23607, N21941, N23196);
nand NAND2_2569 (N23608, N21938, N23197);
nand NAND2_2570 (N23609, N21965, N23198);
nand NAND2_2571 (N23610, N21962, N23199);
not NOT1_2572 (N23613, N23191);
and AND2_2573 (N23614, N22882, N22891);
and AND2_2574 (N23615, N21482, N22891);
and AND3_2575 (N23616, N2200, N22653, N21173);
and AND3_2576 (N23617, N2203, N22653, N21173);
and AND3_2577 (N23618, N2197, N22653, N21173);
and AND3_2578 (N23619, N2194, N22653, N21173);
and AND3_2579 (N23620, N2191, N22653, N21173);
and AND3_2580 (N23621, N2182, N22681, N21197);
and AND3_2581 (N23622, N2188, N22681, N21197);
and AND3_2582 (N23623, N2155, N22681, N21197);
and AND3_2583 (N23624, N2149, N22681, N21197);
and AND2_2584 (N23625, N22882, N22891);
and AND2_2585 (N23626, N21482, N22891);
and AND3_2586 (N23627, N2200, N22728, N21235);
and AND3_2587 (N23628, N2203, N22728, N21235);
and AND3_2588 (N23629, N2197, N22728, N21235);
and AND3_2589 (N23630, N2194, N22728, N21235);
and AND3_2590 (N23631, N2191, N22728, N21235);
and AND3_2591 (N23632, N2182, N22756, N21259);
and AND3_2592 (N23633, N2188, N22756, N21259);
and AND3_2593 (N23634, N2155, N22756, N21259);
and AND3_2594 (N23635, N2149, N22756, N21259);
and AND2_2595 (N23636, N22882, N22891);
and AND2_2596 (N23637, N21482, N22891);
and AND3_2597 (N23638, N2109, N23075, N21743);
and AND2_2598 (N23639, N22882, N22891);
and AND2_2599 (N23640, N21482, N22891);
and AND3_2600 (N23641, N211, N22779, N21339);
and AND3_2601 (N23642, N2109, N23041, N21709);
and AND3_2602 (N23643, N246, N23041, N21709);
and AND3_2603 (N23644, N2100, N23041, N21709);
and AND3_2604 (N23645, N291, N23041, N21709);
and AND3_2605 (N23646, N243, N23041, N21709);
and AND3_2606 (N23647, N276, N22779, N21339);
and AND3_2607 (N23648, N273, N22779, N21339);
and AND3_2608 (N23649, N267, N22779, N21339);
and AND3_2609 (N23650, N214, N22779, N21339);
and AND3_2610 (N23651, N246, N23075, N21743);
and AND3_2611 (N23652, N2100, N23075, N21743);
and AND3_2612 (N23653, N291, N23075, N21743);
and AND3_2613 (N23654, N243, N23075, N21743);
and AND3_2614 (N23655, N276, N22801, N21363);
and AND3_2615 (N23656, N273, N22801, N21363);
and AND3_2616 (N23657, N267, N22801, N21363);
and AND3_2617 (N23658, N214, N22801, N21363);
and AND3_2618 (N23659, N2120, N23119, N21785);
and AND3_2619 (N23660, N211, N22801, N21363);
and AND3_2620 (N23661, N2118, N23097, N21769);
and AND3_2621 (N23662, N2176, N22681, N21197);
and AND3_2622 (N23663, N2176, N22756, N21259);
or OR2_2623 (N23664, N22831, N23401);
or OR2_2624 (N23665, N22832, N23402);
or OR2_2625 (N23666, N22833, N23403);
or OR2_2626 (N23667, N22834, N23404);
or OR3_2627 (N23668, N22835, N23405, N2457);
or OR3_2628 (N23669, N22836, N23406, N2468);
or OR3_2629 (N23670, N22837, N23407, N2422);
or OR3_2630 (N23671, N22838, N23408, N2435);
or OR2_2631 (N23672, N22847, N23409);
or OR2_2632 (N23673, N22848, N23410);
or OR2_2633 (N23674, N22849, N23411);
or OR2_2634 (N23675, N22850, N23412);
or OR3_2635 (N23676, N22851, N23413, N2389);
or OR3_2636 (N23677, N22852, N23414, N2400);
or OR3_2637 (N23678, N22853, N23415, N2411);
or OR3_2638 (N23679, N22854, N23416, N2374);
and AND2_2639 (N23680, N2289, N22855);
and AND2_2640 (N23681, N2281, N22855);
and AND2_2641 (N23682, N2273, N22855);
and AND2_2642 (N23683, N2265, N22855);
and AND2_2643 (N23684, N2257, N22855);
and AND2_2644 (N23685, N2234, N22861);
and AND2_2645 (N23686, N2226, N22861);
and AND2_2646 (N23687, N2218, N22861);
and AND2_2647 (N23688, N2210, N22861);
and AND2_2648 (N23689, N2206, N22861);
not NOT1_2649 (N23691, N22891);
or OR2_2650 (N23700, N22907, N23444);
or OR2_2651 (N23701, N22908, N23445);
or OR2_2652 (N23702, N22909, N23446);
or OR3_2653 (N23703, N22911, N23448, N2479);
or OR3_2654 (N23704, N22912, N23449, N2490);
or OR2_2655 (N23705, N22910, N23447);
or OR2_2656 (N23708, N22919, N23450);
or OR2_2657 (N23709, N22921, N23451);
or OR2_2658 (N23710, N22922, N23452);
or OR3_2659 (N23711, N22923, N23453, N2503);
or OR3_2660 (N23712, N22924, N23454, N2523);
or OR3_2661 (N23713, N22925, N23455, N2534);
or OR2_2662 (N23715, N22934, N23459);
or OR2_2663 (N23716, N22935, N23460);
or OR2_2664 (N23717, N22936, N23461);
or OR2_2665 (N23718, N22937, N23462);
or OR3_2666 (N23719, N22938, N23463, N2389);
or OR3_2667 (N23720, N22939, N23464, N2400);
or OR3_2668 (N23721, N22940, N23465, N2411);
or OR3_2669 (N23722, N22941, N23466, N2374);
and AND2_2670 (N23723, N2369, N22942);
and AND2_2671 (N23724, N2361, N22942);
and AND2_2672 (N23725, N2351, N22942);
and AND2_2673 (N23726, N2341, N22942);
and AND2_2674 (N23727, N2324, N22948);
and AND2_2675 (N23728, N2316, N22948);
and AND2_2676 (N23729, N2308, N22948);
and AND2_2677 (N23730, N2302, N22948);
and AND2_2678 (N23731, N2293, N22948);
or OR2_2679 (N23732, N22942, N22958);
and AND2_2680 (N23738, N283, N22964);
and AND2_2681 (N23739, N287, N22964);
and AND2_2682 (N23740, N234, N22964);
and AND2_2683 (N23741, N234, N22964);
or OR2_2684 (N23742, N22979, N23481);
or OR2_2685 (N23743, N22981, N23483);
or OR2_2686 (N23744, N22982, N23484);
or OR3_2687 (N23745, N22983, N23485, N2503);
or OR3_2688 (N23746, N22985, N23486, N2523);
or OR3_2689 (N23747, N22986, N23487, N2534);
or OR2_2690 (N23748, N22993, N23488);
or OR2_2691 (N23749, N22994, N23489);
or OR2_2692 (N23750, N22995, N23490);
or OR3_2693 (N23751, N22997, N23492, N2479);
or OR3_2694 (N23752, N22998, N23493, N2490);
not NOT1_2695 (N23753, N23000);
not NOT1_2696 (N23754, N23003);
not NOT1_2697 (N23755, N23007);
not NOT1_2698 (N23756, N23010);
or OR2_2699 (N23757, N23013, N23502);
and AND3_2700 (N23758, N21315, N2446, N23003);
or OR2_2701 (N23759, N23014, N23503);
and AND3_2702 (N23760, N21315, N2446, N23010);
and AND2_2703 (N23761, N21675, N23000);
and AND2_2704 (N23762, N21675, N23007);
or OR2_2705 (N23763, N23023, N23504);
or OR2_2706 (N23764, N23024, N23505);
or OR2_2707 (N23765, N23025, N23506);
or OR2_2708 (N23766, N23026, N23507);
or OR3_2709 (N23767, N23027, N23508, N2457);
or OR3_2710 (N23768, N23028, N23509, N2468);
or OR3_2711 (N23769, N23029, N23510, N2422);
or OR3_2712 (N23770, N23030, N23511, N2435);
nand NAND2_2713 (N23771, N23512, N23513);
nand NAND2_2714 (N23775, N23514, N23515);
not NOT1_2715 (N23779, N23035);
not NOT1_2716 (N23780, N23038);
and AND3_2717 (N23781, N2117, N23097, N21769);
and AND3_2718 (N23782, N2126, N23097, N21769);
and AND3_2719 (N23783, N2127, N23097, N21769);
and AND3_2720 (N23784, N2128, N23097, N21769);
and AND3_2721 (N23785, N2131, N23119, N21785);
and AND3_2722 (N23786, N2129, N23119, N21785);
and AND3_2723 (N23787, N2119, N23119, N21785);
and AND3_2724 (N23788, N2130, N23119, N21785);
nand NAND2_2725 (N23789, N23558, N23559);
nand NAND2_2726 (N23793, N23560, N23561);
nand NAND2_2727 (N23797, N23562, N23563);
and AND3_2728 (N23800, N2122, N23147, N21800);
and AND3_2729 (N23801, N2113, N23147, N21800);
and AND3_2730 (N23802, N253, N23147, N21800);
and AND3_2731 (N23803, N2114, N23147, N21800);
and AND3_2732 (N23804, N2115, N23147, N21800);
and AND3_2733 (N23805, N252, N23169, N21814);
and AND3_2734 (N23806, N2112, N23169, N21814);
and AND3_2735 (N23807, N2116, N23169, N21814);
and AND3_2736 (N23808, N2121, N23169, N21814);
and AND3_2737 (N23809, N2123, N23169, N21814);
nand NAND2_2738 (N23810, N23607, N23608);
nand NAND2_2739 (N23813, N23605, N23606);
and AND2_2740 (N23816, N23482, N22984);
or OR2_2741 (N23819, N22996, N23491);
not NOT1_2742 (N23822, N23200);
nand NAND2_2743 (N23823, N23200, N23203);
nand NAND2_2744 (N23824, N23609, N23610);
not NOT1_2745 (N23827, N23456);
or OR2_2746 (N23828, N23739, N22970);
or OR2_2747 (N23829, N23740, N22971);
or OR2_2748 (N23830, N23741, N22972);
or OR2_2749 (N23831, N23738, N22969);
not NOT1_2750 (N23834, N23664);
not NOT1_2751 (N23835, N23665);
not NOT1_2752 (N23836, N23666);
not NOT1_2753 (N23837, N23667);
not NOT1_2754 (N23838, N23672);
not NOT1_2755 (N23839, N23673);
not NOT1_2756 (N23840, N23674);
not NOT1_2757 (N23841, N23675);
or OR2_2758 (N23842, N23681, N22868);
or OR2_2759 (N23849, N23682, N22869);
or OR2_2760 (N23855, N23683, N22870);
or OR2_2761 (N23861, N23684, N22871);
or OR2_2762 (N23867, N23685, N22872);
or OR2_2763 (N23873, N23686, N22873);
or OR2_2764 (N23881, N23687, N22874);
or OR2_2765 (N23887, N23688, N22875);
or OR2_2766 (N23893, N23689, N22876);
not NOT1_2767 (N23908, N23701);
not NOT1_2768 (N23909, N23702);
not NOT1_2769 (N23911, N23700);
not NOT1_2770 (N23914, N23708);
not NOT1_2771 (N23915, N23709);
not NOT1_2772 (N23916, N23710);
not NOT1_2773 (N23917, N23715);
not NOT1_2774 (N23918, N23716);
not NOT1_2775 (N23919, N23717);
not NOT1_2776 (N23920, N23718);
or OR2_2777 (N23921, N23724, N22955);
or OR2_2778 (N23927, N23725, N22956);
or OR2_2779 (N23933, N23726, N22957);
or OR2_2780 (N23942, N23727, N22959);
or OR2_2781 (N23948, N23728, N22960);
or OR2_2782 (N23956, N23729, N22961);
or OR2_2783 (N23962, N23730, N22962);
or OR2_2784 (N23968, N23731, N22963);
not NOT1_2785 (N23975, N23742);
not NOT1_2786 (N23976, N23743);
not NOT1_2787 (N23977, N23744);
not NOT1_2788 (N23978, N23749);
not NOT1_2789 (N23979, N23750);
and AND3_2790 (N23980, N2446, N21292, N23754);
and AND3_2791 (N23981, N2446, N21292, N23756);
and AND2_2792 (N23982, N21271, N23753);
and AND2_2793 (N23983, N21271, N23755);
not NOT1_2794 (N23984, N23757);
not NOT1_2795 (N23987, N23759);
not NOT1_2796 (N23988, N23763);
not NOT1_2797 (N23989, N23764);
not NOT1_2798 (N23990, N23765);
not NOT1_2799 (N23991, N23766);
and AND3_2800 (N23998, N23456, N23119, N23130);
or OR2_2801 (N24008, N23723, N22954);
or OR2_2802 (N24011, N23680, N22867);
not NOT1_2803 (N24021, N23748);
nand NAND2_2804 (N24024, N21968, N23822);
not NOT1_2805 (N24027, N23705);
and AND2_2806 (N24031, N23828, N21583);
and AND3_2807 (N24032, N224, N22882, N23691);
and AND3_2808 (N24033, N225, N21482, N23691);
and AND3_2809 (N24034, N226, N22882, N23691);
and AND3_2810 (N24035, N281, N21482, N23691);
and AND2_2811 (N24036, N23829, N21583);
and AND3_2812 (N24037, N279, N22882, N23691);
and AND3_2813 (N24038, N223, N21482, N23691);
and AND3_2814 (N24039, N282, N22882, N23691);
and AND3_2815 (N24040, N280, N21482, N23691);
and AND2_2816 (N24041, N23830, N21583);
and AND2_2817 (N24042, N23831, N21583);
and AND2_2818 (N24067, N23732, N2514);
and AND2_2819 (N24080, N2514, N23732);
and AND2_2820 (N24088, N23834, N23668);
and AND2_2821 (N24091, N23835, N23669);
and AND2_2822 (N24094, N23836, N23670);
and AND2_2823 (N24097, N23837, N23671);
and AND2_2824 (N24100, N23838, N23676);
and AND2_2825 (N24103, N23839, N23677);
and AND2_2826 (N24106, N23840, N23678);
and AND2_2827 (N24109, N23841, N23679);
and AND2_2828 (N24144, N23908, N23703);
and AND2_2829 (N24147, N23909, N23704);
buf BUFF1_2830 (N24150, N23705);
and AND2_2831 (N24153, N23914, N23711);
and AND2_2832 (N24156, N23915, N23712);
and AND2_2833 (N24159, N23916, N23713);
or OR2_2834 (N24183, N23758, N23980);
or OR2_2835 (N24184, N23760, N23981);
or OR3_2836 (N24185, N23761, N23982, N2446);
or OR3_2837 (N24186, N23762, N23983, N2446);
not NOT1_2838 (N24188, N23771);
not NOT1_2839 (N24191, N23775);
and AND3_2840 (N24196, N23775, N23771, N23035);
and AND3_2841 (N24197, N23987, N23119, N23130);
and AND2_2842 (N24198, N23920, N23722);
not NOT1_2843 (N24199, N23816);
not NOT1_2844 (N24200, N23789);
not NOT1_2845 (N24203, N23793);
buf BUFF1_2846 (N24206, N23797);
buf BUFF1_2847 (N24209, N23797);
buf BUFF1_2848 (N24212, N23732);
buf BUFF1_2849 (N24215, N23732);
buf BUFF1_2850 (N24219, N23732);
not NOT1_2851 (N24223, N23810);
not NOT1_2852 (N24224, N23813);
and AND2_2853 (N24225, N23918, N23720);
and AND2_2854 (N24228, N23919, N23721);
and AND2_2855 (N24231, N23991, N23770);
and AND2_2856 (N24234, N23917, N23719);
and AND2_2857 (N24237, N23989, N23768);
and AND2_2858 (N24240, N23990, N23769);
and AND2_2859 (N24243, N23988, N23767);
and AND2_2860 (N24246, N23976, N23746);
and AND2_2861 (N24249, N23977, N23747);
and AND2_2862 (N24252, N23975, N23745);
and AND2_2863 (N24255, N23978, N23751);
and AND2_2864 (N24258, N23979, N23752);
not NOT1_2865 (N24263, N23819);
nand NAND2_2866 (N24264, N24024, N23823);
not NOT1_2867 (N24267, N23824);
and AND2_2868 (N24268, N2446, N23893);
not NOT1_2869 (N24269, N23911);
not NOT1_2870 (N24270, N23984);
and AND2_2871 (N24271, N23893, N2446);
not NOT1_2872 (N24272, N24031);
or OR4_2873 (N24273, N24032, N24033, N23614, N23615);
or OR4_2874 (N24274, N24034, N24035, N23625, N23626);
not NOT1_2875 (N24275, N24036);
or OR4_2876 (N24276, N24037, N24038, N23636, N23637);
or OR4_2877 (N24277, N24039, N24040, N23639, N23640);
not NOT1_2878 (N24278, N24041);
not NOT1_2879 (N24279, N24042);
and AND2_2880 (N24280, N23887, N2457);
and AND2_2881 (N24284, N23881, N2468);
and AND2_2882 (N24290, N2422, N23873);
and AND2_2883 (N24297, N23867, N2435);
and AND2_2884 (N24298, N23861, N2389);
and AND2_2885 (N24301, N23855, N2400);
and AND2_2886 (N24305, N23849, N2411);
and AND2_2887 (N24310, N23842, N2374);
and AND2_2888 (N24316, N2457, N23887);
and AND2_2889 (N24320, N2468, N23881);
and AND2_2890 (N24325, N2422, N23873);
and AND2_2891 (N24331, N2435, N23867);
and AND2_2892 (N24332, N2389, N23861);
and AND2_2893 (N24336, N2400, N23855);
and AND2_2894 (N24342, N2411, N23849);
and AND2_2895 (N24349, N2374, N23842);
not NOT1_2896 (N24357, N23968);
not NOT1_2897 (N24364, N23962);
buf BUFF1_2898 (N24375, N23962);
and AND2_2899 (N24379, N23956, N2479);
and AND2_2900 (N24385, N2490, N23948);
and AND2_2901 (N24392, N23942, N2503);
and AND2_2902 (N24396, N23933, N2523);
and AND2_2903 (N24400, N23927, N2534);
not NOT1_2904 (N24405, N23921);
buf BUFF1_2905 (N24412, N23921);
not NOT1_2906 (N24418, N23968);
not NOT1_2907 (N24425, N23962);
buf BUFF1_2908 (N24436, N23962);
and AND2_2909 (N24440, N2479, N23956);
and AND2_2910 (N24445, N2490, N23948);
and AND2_2911 (N24451, N2503, N23942);
and AND2_2912 (N24456, N2523, N23933);
and AND2_2913 (N24462, N2534, N23927);
buf BUFF1_2914 (N24469, N23921);
not NOT1_2915 (N24477, N23921);
buf BUFF1_2916 (N24512, N23968);
not NOT1_2917 (N24515, N24183);
not NOT1_2918 (N24516, N24184);
not NOT1_2919 (N24521, N24008);
not NOT1_2920 (N24523, N24011);
not NOT1_2921 (N24524, N24198);
not NOT1_2922 (N24532, N23984);
and AND3_2923 (N24547, N23911, N23169, N23180);
buf BUFF1_2924 (N24548, N23893);
buf BUFF1_2925 (N24551, N23887);
buf BUFF1_2926 (N24554, N23881);
buf BUFF1_2927 (N24557, N23873);
buf BUFF1_2928 (N24560, N23867);
buf BUFF1_2929 (N24563, N23861);
buf BUFF1_2930 (N24566, N23855);
buf BUFF1_2931 (N24569, N23849);
buf BUFF1_2932 (N24572, N23842);
nor N2OR2_2933 (N24575, N2422, N23873);
buf BUFF1_2934 (N24578, N23893);
buf BUFF1_2935 (N24581, N23887);
buf BUFF1_2936 (N24584, N23881);
buf BUFF1_2937 (N24587, N23867);
buf BUFF1_2938 (N24590, N23861);
buf BUFF1_2939 (N24593, N23855);
buf BUFF1_2940 (N24596, N23849);
buf BUFF1_2941 (N24599, N23873);
buf BUFF1_2942 (N24602, N23842);
nor N2OR2_2943 (N24605, N2422, N23873);
nor N2OR2_2944 (N24608, N2374, N23842);
buf BUFF1_2945 (N24611, N23956);
buf BUFF1_2946 (N24614, N23948);
buf BUFF1_2947 (N24617, N23942);
buf BUFF1_2948 (N24621, N23933);
buf BUFF1_2949 (N24624, N23927);
nor N2OR2_2950 (N24627, N2490, N23948);
buf BUFF1_2951 (N24630, N23956);
buf BUFF1_2952 (N24633, N23942);
buf BUFF1_2953 (N24637, N23933);
buf BUFF1_2954 (N24640, N23927);
buf BUFF1_2955 (N24643, N23948);
nor N2OR2_2956 (N24646, N2490, N23948);
buf BUFF1_2957 (N24649, N23927);
buf BUFF1_2958 (N24652, N23933);
buf BUFF1_2959 (N24655, N23921);
buf BUFF1_2960 (N24658, N23942);
buf BUFF1_2961 (N24662, N23956);
buf BUFF1_2962 (N24665, N23948);
buf BUFF1_2963 (N24668, N23968);
buf BUFF1_2964 (N24671, N23962);
buf BUFF1_2965 (N24674, N23873);
buf BUFF1_2966 (N24677, N23867);
buf BUFF1_2967 (N24680, N23887);
buf BUFF1_2968 (N24683, N23881);
buf BUFF1_2969 (N24686, N23893);
buf BUFF1_2970 (N24689, N23849);
buf BUFF1_2971 (N24692, N23842);
buf BUFF1_2972 (N24695, N23861);
buf BUFF1_2973 (N24698, N23855);
nand NAND2_2974 (N24701, N23813, N24223);
nand NAND2_2975 (N24702, N23810, N24224);
not NOT1_2976 (N24720, N24021);
nand NAND2_2977 (N24721, N24021, N24263);
not NOT1_2978 (N24724, N24147);
not NOT1_2979 (N24725, N24144);
not NOT1_2980 (N24726, N24159);
not NOT1_2981 (N24727, N24156);
not NOT1_2982 (N24728, N24153);
not NOT1_2983 (N24729, N24097);
not NOT1_2984 (N24730, N24094);
not NOT1_2985 (N24731, N24091);
not NOT1_2986 (N24732, N24088);
not NOT1_2987 (N24733, N24109);
not NOT1_2988 (N24734, N24106);
not NOT1_2989 (N24735, N24103);
not NOT1_2990 (N24736, N24100);
and AND2_2991 (N24737, N24273, N22877);
and AND2_2992 (N24738, N24274, N22877);
and AND2_2993 (N24739, N24276, N22877);
and AND2_2994 (N24740, N24277, N22877);
and AND3_2995 (N24741, N24150, N21758, N21755);
not NOT1_2996 (N24855, N24212);
nand NAND2_2997 (N24856, N24212, N22712);
nand NAND2_2998 (N24908, N24215, N22718);
not NOT1_2999 (N24909, N24215);
and AND2_21000 (N24939, N24515, N24185);
and AND2_21001 (N24942, N24516, N24186);
not NOT1_21002 (N24947, N24219);
and AND3_21003 (N24953, N24188, N23775, N23779);
and AND3_21004 (N24954, N23771, N24191, N23780);
and AND3_21005 (N24955, N24191, N24188, N23038);
and AND3_21006 (N24956, N24109, N23097, N23108);
and AND3_21007 (N24957, N24106, N23097, N23108);
and AND3_21008 (N24958, N24103, N23097, N23108);
and AND3_21009 (N24959, N24100, N23097, N23108);
and AND3_21010 (N24960, N24159, N23119, N23130);
and AND3_21011 (N24961, N24156, N23119, N23130);
not NOT1_21012 (N24965, N24225);
not NOT1_21013 (N24966, N24228);
not NOT1_21014 (N24967, N24231);
not NOT1_21015 (N24968, N24234);
not NOT1_21016 (N24972, N24246);
not NOT1_21017 (N24973, N24249);
not NOT1_21018 (N24974, N24252);
nand NAND2_21019 (N24975, N24252, N24199);
not NOT1_21020 (N24976, N24206);
not NOT1_21021 (N24977, N24209);
and AND3_21022 (N24978, N23793, N23789, N24206);
and AND3_21023 (N24979, N24203, N24200, N24209);
and AND3_21024 (N24980, N24097, N23147, N23158);
and AND3_21025 (N24981, N24094, N23147, N23158);
and AND3_21026 (N24982, N24091, N23147, N23158);
and AND3_21027 (N24983, N24088, N23147, N23158);
and AND3_21028 (N24984, N24153, N23169, N23180);
and AND3_21029 (N24985, N24147, N23169, N23180);
and AND3_21030 (N24986, N24144, N23169, N23180);
and AND3_21031 (N24987, N24150, N23169, N23180);
nand NAND2_21032 (N25049, N24701, N24702);
not NOT1_21033 (N25052, N24237);
not NOT1_21034 (N25053, N24240);
not NOT1_21035 (N25054, N24243);
not NOT1_21036 (N25055, N24255);
not NOT1_21037 (N25056, N24258);
nand NAND2_21038 (N25057, N23819, N24720);
not NOT1_21039 (N25058, N24264);
nand NAND2_21040 (N25059, N24264, N24267);
and AND4_21041 (N25060, N24724, N24725, N24269, N24027);
and AND4_21042 (N25061, N24726, N24727, N23827, N24728);
and AND4_21043 (N25062, N24729, N24730, N24731, N24732);
and AND4_21044 (N25063, N24733, N24734, N24735, N24736);
and AND2_21045 (N25065, N24357, N24375);
and AND3_21046 (N25066, N24364, N24357, N24379);
and AND2_21047 (N25067, N24418, N24436);
and AND3_21048 (N25068, N24425, N24418, N24440);
not NOT1_21049 (N25069, N24548);
nand NAND2_21050 (N25070, N24548, N22628);
not NOT1_21051 (N25071, N24551);
nand NAND2_21052 (N25072, N24551, N22629);
not NOT1_21053 (N25073, N24554);
nand NAND2_21054 (N25074, N24554, N22630);
not NOT1_21055 (N25075, N24557);
nand NAND2_21056 (N25076, N24557, N22631);
not NOT1_21057 (N25077, N24560);
nand NAND2_21058 (N25078, N24560, N22632);
not NOT1_21059 (N25079, N24563);
nand NAND2_21060 (N25080, N24563, N22633);
not NOT1_21061 (N25081, N24566);
nand NAND2_21062 (N25082, N24566, N22634);
not NOT1_21063 (N25083, N24569);
nand NAND2_21064 (N25084, N24569, N22635);
not NOT1_21065 (N25085, N24572);
nand NAND2_21066 (N25086, N24572, N22636);
not NOT1_21067 (N25087, N24575);
nand NAND2_21068 (N25088, N24578, N22638);
not NOT1_21069 (N25089, N24578);
nand NAND2_21070 (N25090, N24581, N22639);
not NOT1_21071 (N25091, N24581);
nand NAND2_21072 (N25092, N24584, N22640);
not NOT1_21073 (N25093, N24584);
nand NAND2_21074 (N25094, N24587, N22641);
not NOT1_21075 (N25095, N24587);
nand NAND2_21076 (N25096, N24590, N22642);
not NOT1_21077 (N25097, N24590);
nand NAND2_21078 (N25098, N24593, N22643);
not NOT1_21079 (N25099, N24593);
nand NAND2_21080 (N25100, N24596, N22644);
not NOT1_21081 (N25101, N24596);
nand NAND2_21082 (N25102, N24599, N22645);
not NOT1_21083 (N25103, N24599);
nand NAND2_21084 (N25104, N24602, N22646);
not NOT1_21085 (N25105, N24602);
not NOT1_21086 (N25106, N24611);
nand NAND2_21087 (N25107, N24611, N22709);
not NOT1_21088 (N25108, N24614);
nand NAND2_21089 (N25109, N24614, N22710);
not NOT1_21090 (N25110, N24617);
nand NAND2_21091 (N25111, N24617, N22711);
nand NAND2_21092 (N25112, N21890, N24855);
not NOT1_21093 (N25113, N24621);
nand NAND2_21094 (N25114, N24621, N22713);
not NOT1_21095 (N25115, N24624);
nand NAND2_21096 (N25116, N24624, N22714);
and AND2_21097 (N25117, N24364, N24379);
and AND2_21098 (N25118, N24364, N24379);
and AND2_21099 (N25119, N254, N24405);
not NOT1_21100 (N25120, N24627);
nand NAND2_21101 (N25121, N24630, N22716);
not NOT1_21102 (N25122, N24630);
nand NAND2_21103 (N25123, N24633, N22717);
not NOT1_21104 (N25124, N24633);
nand NAND2_21105 (N25125, N21908, N24909);
nand NAND2_21106 (N25126, N24637, N22719);
not NOT1_21107 (N25127, N24637);
nand NAND2_21108 (N25128, N24640, N22720);
not NOT1_21109 (N25129, N24640);
nand NAND2_21110 (N25130, N24643, N22721);
not NOT1_21111 (N25131, N24643);
and AND2_21112 (N25132, N24425, N24440);
and AND2_21113 (N25133, N24425, N24440);
not NOT1_21114 (N25135, N24649);
not NOT1_21115 (N25136, N24652);
nand NAND2_21116 (N25137, N24655, N24521);
not NOT1_21117 (N25138, N24655);
not NOT1_21118 (N25139, N24658);
nand NAND2_21119 (N25140, N24658, N24947);
not NOT1_21120 (N25141, N24674);
not NOT1_21121 (N25142, N24677);
not NOT1_21122 (N25143, N24680);
not NOT1_21123 (N25144, N24683);
nand NAND2_21124 (N25145, N24686, N24523);
not NOT1_21125 (N25146, N24686);
nor N2OR2_21126 (N25147, N24953, N24196);
nor N2OR2_21127 (N25148, N24954, N24955);
not NOT1_21128 (N25150, N24524);
nand NAND2_21129 (N25153, N24228, N24965);
nand NAND2_21130 (N25154, N24225, N24966);
nand NAND2_21131 (N25155, N24234, N24967);
nand NAND2_21132 (N25156, N24231, N24968);
not NOT1_21133 (N25157, N24532);
nand NAND2_21134 (N25160, N24249, N24972);
nand NAND2_21135 (N25161, N24246, N24973);
nand NAND2_21136 (N25162, N23816, N24974);
and AND3_21137 (N25163, N24200, N23793, N24976);
and AND3_21138 (N25164, N23789, N24203, N24977);
and AND3_21139 (N25165, N24942, N23147, N23158);
not NOT1_21140 (N25166, N24512);
buf BUFF1_21141 (N25169, N24290);
not NOT1_21142 (N25172, N24605);
buf BUFF1_21143 (N25173, N24325);
not NOT1_21144 (N25176, N24608);
buf BUFF1_21145 (N25177, N24349);
buf BUFF1_21146 (N25180, N24405);
buf BUFF1_21147 (N25183, N24357);
buf BUFF1_21148 (N25186, N24357);
buf BUFF1_21149 (N25189, N24364);
buf BUFF1_21150 (N25192, N24364);
buf BUFF1_21151 (N25195, N24385);
not NOT1_21152 (N25198, N24646);
buf BUFF1_21153 (N25199, N24418);
buf BUFF1_21154 (N25202, N24425);
buf BUFF1_21155 (N25205, N24445);
buf BUFF1_21156 (N25208, N24418);
buf BUFF1_21157 (N25211, N24425);
buf BUFF1_21158 (N25214, N24477);
buf BUFF1_21159 (N25217, N24469);
buf BUFF1_21160 (N25220, N24477);
not NOT1_21161 (N25223, N24662);
not NOT1_21162 (N25224, N24665);
not NOT1_21163 (N25225, N24668);
not NOT1_21164 (N25226, N24671);
not NOT1_21165 (N25227, N24689);
not NOT1_21166 (N25228, N24692);
not NOT1_21167 (N25229, N24695);
not NOT1_21168 (N25230, N24698);
nand NAND2_21169 (N25232, N24240, N25052);
nand NAND2_21170 (N25233, N24237, N25053);
nand NAND2_21171 (N25234, N24258, N25055);
nand NAND2_21172 (N25235, N24255, N25056);
nand NAND2_21173 (N25236, N24721, N25057);
nand NAND2_21174 (N25239, N23824, N25058);
and AND3_21175 (N25240, N25060, N25061, N24270);
not NOT1_21176 (N25241, N24939);
nand NAND2_21177 (N25242, N21824, N25069);
nand NAND2_21178 (N25243, N21827, N25071);
nand NAND2_21179 (N25244, N21830, N25073);
nand NAND2_21180 (N25245, N21833, N25075);
nand NAND2_21181 (N25246, N21836, N25077);
nand NAND2_21182 (N25247, N21839, N25079);
nand NAND2_21183 (N25248, N21842, N25081);
nand NAND2_21184 (N25249, N21845, N25083);
nand NAND2_21185 (N25250, N21848, N25085);
nand NAND2_21186 (N25252, N21854, N25089);
nand NAND2_21187 (N25253, N21857, N25091);
nand NAND2_21188 (N25254, N21860, N25093);
nand NAND2_21189 (N25255, N21863, N25095);
nand NAND2_21190 (N25256, N21866, N25097);
nand NAND2_21191 (N25257, N21869, N25099);
nand NAND2_21192 (N25258, N21872, N25101);
nand NAND2_21193 (N25259, N21875, N25103);
nand NAND2_21194 (N25260, N21878, N25105);
nand NAND2_21195 (N25261, N21881, N25106);
nand NAND2_21196 (N25262, N21884, N25108);
nand NAND2_21197 (N25263, N21887, N25110);
nand NAND2_21198 (N25264, N25112, N24856);
nand NAND2_21199 (N25274, N21893, N25113);
nand NAND2_21200 (N25275, N21896, N25115);
nand NAND2_21201 (N25282, N21902, N25122);
nand NAND2_21202 (N25283, N21905, N25124);
nand NAND2_21203 (N25284, N24908, N25125);
nand NAND2_21204 (N25298, N21911, N25127);
nand NAND2_21205 (N25299, N21914, N25129);
nand NAND2_21206 (N25300, N21917, N25131);
nand NAND2_21207 (N25303, N24652, N25135);
nand NAND2_21208 (N25304, N24649, N25136);
nand NAND2_21209 (N25305, N24008, N25138);
nand NAND2_21210 (N25306, N24219, N25139);
nand NAND2_21211 (N25307, N24677, N25141);
nand NAND2_21212 (N25308, N24674, N25142);
nand NAND2_21213 (N25309, N24683, N25143);
nand NAND2_21214 (N25310, N24680, N25144);
nand NAND2_21215 (N25311, N24011, N25146);
not NOT1_21216 (N25312, N25049);
nand NAND2_21217 (N25315, N25153, N25154);
nand NAND2_21218 (N25319, N25155, N25156);
nand NAND2_21219 (N25324, N25160, N25161);
nand NAND2_21220 (N25328, N25162, N24975);
nor N2OR2_21221 (N25331, N25163, N24978);
nor N2OR2_21222 (N25332, N25164, N24979);
or OR2_21223 (N25346, N24412, N25119);
nand NAND2_21224 (N25363, N24665, N25223);
nand NAND2_21225 (N25364, N24662, N25224);
nand NAND2_21226 (N25365, N24671, N25225);
nand NAND2_21227 (N25366, N24668, N25226);
nand NAND2_21228 (N25367, N24692, N25227);
nand NAND2_21229 (N25368, N24689, N25228);
nand NAND2_21230 (N25369, N24698, N25229);
nand NAND2_21231 (N25370, N24695, N25230);
nand NAND2_21232 (N25371, N25148, N25147);
buf BUFF1_21233 (N25374, N24939);
nand NAND2_21234 (N25377, N25232, N25233);
nand NAND2_21235 (N25382, N25234, N25235);
nand NAND2_21236 (N25385, N25239, N25059);
and AND3_21237 (N25388, N25062, N25063, N25241);
nand NAND2_21238 (N25389, N25242, N25070);
nand NAND2_21239 (N25396, N25243, N25072);
nand NAND2_21240 (N25407, N25244, N25074);
nand NAND2_21241 (N25418, N25245, N25076);
nand NAND2_21242 (N25424, N25246, N25078);
nand NAND2_21243 (N25431, N25247, N25080);
nand NAND2_21244 (N25441, N25248, N25082);
nand NAND2_21245 (N25452, N25249, N25084);
nand NAND2_21246 (N25462, N25250, N25086);
not NOT1_21247 (N25469, N25169);
nand NAND2_21248 (N25470, N25088, N25252);
nand NAND2_21249 (N25477, N25090, N25253);
nand NAND2_21250 (N25488, N25092, N25254);
nand NAND2_21251 (N25498, N25094, N25255);
nand NAND2_21252 (N25506, N25096, N25256);
nand NAND2_21253 (N25520, N25098, N25257);
nand NAND2_21254 (N25536, N25100, N25258);
nand NAND2_21255 (N25549, N25102, N25259);
nand NAND2_21256 (N25555, N25104, N25260);
nand NAND2_21257 (N25562, N25261, N25107);
nand NAND2_21258 (N25573, N25262, N25109);
nand NAND2_21259 (N25579, N25263, N25111);
nand NAND2_21260 (N25595, N25274, N25114);
nand NAND2_21261 (N25606, N25275, N25116);
nand NAND2_21262 (N25616, N25180, N22715);
not NOT1_21263 (N25617, N25180);
not NOT1_21264 (N25618, N25183);
not NOT1_21265 (N25619, N25186);
not NOT1_21266 (N25620, N25189);
not NOT1_21267 (N25621, N25192);
not NOT1_21268 (N25622, N25195);
nand NAND2_21269 (N25624, N25121, N25282);
nand NAND2_21270 (N25634, N25123, N25283);
nand NAND2_21271 (N25655, N25126, N25298);
nand NAND2_21272 (N25671, N25128, N25299);
nand NAND2_21273 (N25684, N25130, N25300);
not NOT1_21274 (N25690, N25202);
not NOT1_21275 (N25691, N25211);
nand NAND2_21276 (N25692, N25303, N25304);
nand NAND2_21277 (N25696, N25137, N25305);
nand NAND2_21278 (N25700, N25306, N25140);
nand NAND2_21279 (N25703, N25307, N25308);
nand NAND2_21280 (N25707, N25309, N25310);
nand NAND2_21281 (N25711, N25145, N25311);
and AND2_21282 (N25726, N25166, N24512);
not NOT1_21283 (N25727, N25173);
not NOT1_21284 (N25728, N25177);
not NOT1_21285 (N25730, N25199);
not NOT1_21286 (N25731, N25205);
not NOT1_21287 (N25732, N25208);
not NOT1_21288 (N25733, N25214);
not NOT1_21289 (N25734, N25217);
not NOT1_21290 (N25735, N25220);
nand NAND2_21291 (N25736, N25365, N25366);
nand NAND2_21292 (N25739, N25363, N25364);
nand NAND2_21293 (N25742, N25369, N25370);
nand NAND2_21294 (N25745, N25367, N25368);
not NOT1_21295 (N25755, N25236);
nand NAND2_21296 (N25756, N25332, N25331);
and AND2_21297 (N25954, N25264, N24396);
nand NAND2_21298 (N25955, N21899, N25617);
not NOT1_21299 (N25956, N25346);
and AND2_21300 (N26005, N25284, N24456);
and AND2_21301 (N26006, N25284, N24456);
not NOT1_21302 (N26023, N25371);
nand NAND2_21303 (N26024, N25371, N25312);
not NOT1_21304 (N26025, N25315);
not NOT1_21305 (N26028, N25324);
buf BUFF1_21306 (N26031, N25319);
buf BUFF1_21307 (N26034, N25319);
buf BUFF1_21308 (N26037, N25328);
buf BUFF1_21309 (N26040, N25328);
not NOT1_21310 (N26044, N25385);
or OR2_21311 (N26045, N25166, N25726);
buf BUFF1_21312 (N26048, N25264);
buf BUFF1_21313 (N26051, N25284);
buf BUFF1_21314 (N26054, N25284);
not NOT1_21315 (N26065, N25374);
nand NAND2_21316 (N26066, N25374, N25054);
not NOT1_21317 (N26067, N25377);
not NOT1_21318 (N26068, N25382);
nand NAND2_21319 (N26069, N25382, N25755);
and AND2_21320 (N26071, N25470, N24316);
and AND3_21321 (N26072, N25477, N25470, N24320);
and AND4_21322 (N26073, N25488, N25470, N24325, N25477);
and AND4_21323 (N26074, N25562, N24357, N24385, N24364);
and AND2_21324 (N26075, N25389, N24280);
and AND3_21325 (N26076, N25396, N25389, N24284);
and AND4_21326 (N26077, N25407, N25389, N24290, N25396);
and AND4_21327 (N26078, N25624, N24418, N24445, N24425);
not NOT1_21328 (N26079, N25418);
and AND4_21329 (N26080, N25396, N25418, N25407, N25389);
and AND2_21330 (N26083, N25396, N24284);
and AND3_21331 (N26084, N25407, N24290, N25396);
and AND3_21332 (N26085, N25418, N25407, N25396);
and AND2_21333 (N26086, N25396, N24284);
and AND3_21334 (N26087, N24290, N25407, N25396);
and AND2_21335 (N26088, N25407, N24290);
and AND2_21336 (N26089, N25418, N25407);
and AND2_21337 (N26090, N25407, N24290);
and AND5_21338 (N26091, N25431, N25462, N25441, N25424, N25452);
and AND2_21339 (N26094, N25424, N24298);
and AND3_21340 (N26095, N25431, N25424, N24301);
and AND4_21341 (N26096, N25441, N25424, N24305, N25431);
and AND5_21342 (N26097, N25452, N25441, N25424, N24310, N25431);
and AND2_21343 (N26098, N25431, N24301);
and AND3_21344 (N26099, N25441, N24305, N25431);
and AND4_21345 (N26100, N25452, N25441, N24310, N25431);
and AND5_21346 (N26101, N24, N25462, N25441, N25452, N25431);
and AND2_21347 (N26102, N24305, N25441);
and AND3_21348 (N26103, N25452, N25441, N24310);
and AND4_21349 (N26104, N24, N25462, N25441, N25452);
and AND2_21350 (N26105, N25452, N24310);
and AND3_21351 (N26106, N24, N25462, N25452);
and AND2_21352 (N26107, N24, N25462);
and AND4_21353 (N26108, N25549, N25488, N25477, N25470);
and AND2_21354 (N26111, N25477, N24320);
and AND3_21355 (N26112, N25488, N24325, N25477);
and AND3_21356 (N26113, N25549, N25488, N25477);
and AND2_21357 (N26114, N25477, N24320);
and AND3_21358 (N26115, N25488, N24325, N25477);
and AND2_21359 (N26116, N25488, N24325);
and AND5_21360 (N26117, N25555, N25536, N25520, N25506, N25498);
and AND2_21361 (N26120, N25498, N24332);
and AND3_21362 (N26121, N25506, N25498, N24336);
and AND4_21363 (N26122, N25520, N25498, N24342, N25506);
and AND5_21364 (N26123, N25536, N25520, N25498, N24349, N25506);
and AND2_21365 (N26124, N25506, N24336);
and AND3_21366 (N26125, N25520, N24342, N25506);
and AND4_21367 (N26126, N25536, N25520, N24349, N25506);
and AND4_21368 (N26127, N25555, N25520, N25506, N25536);
and AND2_21369 (N26128, N25506, N24336);
and AND3_21370 (N26129, N25520, N24342, N25506);
and AND4_21371 (N26130, N25536, N25520, N24349, N25506);
and AND2_21372 (N26131, N25520, N24342);
and AND3_21373 (N26132, N25536, N25520, N24349);
and AND3_21374 (N26133, N25555, N25520, N25536);
and AND2_21375 (N26134, N25520, N24342);
and AND3_21376 (N26135, N25536, N25520, N24349);
and AND2_21377 (N26136, N25536, N24349);
and AND2_21378 (N26137, N25549, N25488);
and AND2_21379 (N26138, N25555, N25536);
not NOT1_21380 (N26139, N25573);
and AND4_21381 (N26140, N24364, N25573, N25562, N24357);
and AND3_21382 (N26143, N25562, N24385, N24364);
and AND3_21383 (N26144, N25573, N25562, N24364);
and AND3_21384 (N26145, N24385, N25562, N24364);
and AND2_21385 (N26146, N25562, N24385);
and AND2_21386 (N26147, N25573, N25562);
and AND2_21387 (N26148, N25562, N24385);
and AND5_21388 (N26149, N25264, N24405, N25595, N25579, N25606);
and AND2_21389 (N26152, N25579, N24067);
and AND3_21390 (N26153, N25264, N25579, N24396);
and AND4_21391 (N26154, N25595, N25579, N24400, N25264);
and AND5_21392 (N26155, N25606, N25595, N25579, N24412, N25264);
and AND3_21393 (N26156, N25595, N24400, N25264);
and AND4_21394 (N26157, N25606, N25595, N24412, N25264);
and AND5_21395 (N26158, N254, N24405, N25595, N25606, N25264);
and AND2_21396 (N26159, N24400, N25595);
and AND3_21397 (N26160, N25606, N25595, N24412);
and AND4_21398 (N26161, N254, N24405, N25595, N25606);
and AND2_21399 (N26162, N25606, N24412);
and AND3_21400 (N26163, N254, N24405, N25606);
nand NAND2_21401 (N26164, N25616, N25955);
and AND4_21402 (N26168, N25684, N25624, N24425, N24418);
and AND3_21403 (N26171, N25624, N24445, N24425);
and AND3_21404 (N26172, N25684, N25624, N24425);
and AND3_21405 (N26173, N25624, N24445, N24425);
and AND2_21406 (N26174, N25624, N24445);
and AND5_21407 (N26175, N24477, N25671, N25655, N25284, N25634);
and AND2_21408 (N26178, N25634, N24080);
and AND3_21409 (N26179, N25284, N25634, N24456);
and AND4_21410 (N26180, N25655, N25634, N24462, N25284);
and AND5_21411 (N26181, N25671, N25655, N25634, N24469, N25284);
and AND3_21412 (N26182, N25655, N24462, N25284);
and AND4_21413 (N26183, N25671, N25655, N24469, N25284);
and AND4_21414 (N26184, N24477, N25655, N25284, N25671);
and AND3_21415 (N26185, N25655, N24462, N25284);
and AND4_21416 (N26186, N25671, N25655, N24469, N25284);
and AND2_21417 (N26187, N25655, N24462);
and AND3_21418 (N26188, N25671, N25655, N24469);
and AND3_21419 (N26189, N24477, N25655, N25671);
and AND2_21420 (N26190, N25655, N24462);
and AND3_21421 (N26191, N25671, N25655, N24469);
and AND2_21422 (N26192, N25671, N24469);
and AND2_21423 (N26193, N25684, N25624);
and AND2_21424 (N26194, N24477, N25671);
not NOT1_21425 (N26197, N25692);
not NOT1_21426 (N26200, N25696);
not NOT1_21427 (N26203, N25703);
not NOT1_21428 (N26206, N25707);
buf BUFF1_21429 (N26209, N25700);
buf BUFF1_21430 (N26212, N25700);
buf BUFF1_21431 (N26215, N25711);
buf BUFF1_21432 (N26218, N25711);
nand NAND2_21433 (N26221, N25049, N26023);
not NOT1_21434 (N26234, N25756);
nand NAND2_21435 (N26235, N25756, N26044);
buf BUFF1_21436 (N26238, N25462);
buf BUFF1_21437 (N26241, N25389);
buf BUFF1_21438 (N26244, N25389);
buf BUFF1_21439 (N26247, N25396);
buf BUFF1_21440 (N26250, N25396);
buf BUFF1_21441 (N26253, N25407);
buf BUFF1_21442 (N26256, N25407);
buf BUFF1_21443 (N26259, N25424);
buf BUFF1_21444 (N26262, N25431);
buf BUFF1_21445 (N26265, N25441);
buf BUFF1_21446 (N26268, N25452);
buf BUFF1_21447 (N26271, N25549);
buf BUFF1_21448 (N26274, N25488);
buf BUFF1_21449 (N26277, N25470);
buf BUFF1_21450 (N26280, N25477);
buf BUFF1_21451 (N26283, N25549);
buf BUFF1_21452 (N26286, N25488);
buf BUFF1_21453 (N26289, N25470);
buf BUFF1_21454 (N26292, N25477);
buf BUFF1_21455 (N26295, N25555);
buf BUFF1_21456 (N26298, N25536);
buf BUFF1_21457 (N26301, N25498);
buf BUFF1_21458 (N26304, N25520);
buf BUFF1_21459 (N26307, N25506);
buf BUFF1_21460 (N26310, N25506);
buf BUFF1_21461 (N26313, N25555);
buf BUFF1_21462 (N26316, N25536);
buf BUFF1_21463 (N26319, N25498);
buf BUFF1_21464 (N26322, N25520);
buf BUFF1_21465 (N26325, N25562);
buf BUFF1_21466 (N26328, N25562);
buf BUFF1_21467 (N26331, N25579);
buf BUFF1_21468 (N26335, N25595);
buf BUFF1_21469 (N26338, N25606);
buf BUFF1_21470 (N26341, N25684);
buf BUFF1_21471 (N26344, N25624);
buf BUFF1_21472 (N26347, N25684);
buf BUFF1_21473 (N26350, N25624);
buf BUFF1_21474 (N26353, N25671);
buf BUFF1_21475 (N26356, N25634);
buf BUFF1_21476 (N26359, N25655);
buf BUFF1_21477 (N26364, N25671);
buf BUFF1_21478 (N26367, N25634);
buf BUFF1_21479 (N26370, N25655);
not NOT1_21480 (N26373, N25736);
not NOT1_21481 (N26374, N25739);
not NOT1_21482 (N26375, N25742);
not NOT1_21483 (N26376, N25745);
nand NAND2_21484 (N26377, N24243, N26065);
nand NAND2_21485 (N26378, N25236, N26068);
or OR4_21486 (N26382, N24268, N26071, N26072, N26073);
or OR4_21487 (N26386, N23968, N25065, N25066, N26074);
or OR4_21488 (N26388, N24271, N26075, N26076, N26077);
or OR4_21489 (N26392, N23968, N25067, N25068, N26078);
or OR5_21490 (N26397, N24297, N26094, N26095, N26096, N26097);
or OR2_21491 (N26411, N24320, N26116);
or OR5_21492 (N26415, N24331, N26120, N26121, N26122, N26123);
or OR2_21493 (N26419, N24342, N26136);
or OR5_21494 (N26427, N24392, N26152, N26153, N26154, N26155);
not NOT1_21495 (N26434, N26048);
or OR2_21496 (N26437, N24440, N26174);
or OR5_21497 (N26441, N24451, N26178, N26179, N26180, N26181);
or OR2_21498 (N26445, N24462, N26192);
not NOT1_21499 (N26448, N26051);
not NOT1_21500 (N26449, N26054);
nand NAND2_21501 (N26466, N26221, N26024);
not NOT1_21502 (N26469, N26031);
not NOT1_21503 (N26470, N26034);
not NOT1_21504 (N26471, N26037);
not NOT1_21505 (N26472, N26040);
and AND3_21506 (N26473, N25315, N24524, N26031);
and AND3_21507 (N26474, N26025, N25150, N26034);
and AND3_21508 (N26475, N25324, N24532, N26037);
and AND3_21509 (N26476, N26028, N25157, N26040);
nand NAND2_21510 (N26477, N25385, N26234);
nand NAND2_21511 (N26478, N26045, N2132);
or OR4_21512 (N26482, N24280, N26083, N26084, N26085);
nor N2OR3_21513 (N26486, N24280, N26086, N26087);
or OR3_21514 (N26490, N24284, N26088, N26089);
nor N2OR2_21515 (N26494, N24284, N26090);
or OR5_21516 (N26500, N24298, N26098, N26099, N26100, N26101);
or OR4_21517 (N26504, N24301, N26102, N26103, N26104);
or OR3_21518 (N26508, N24305, N26105, N26106);
or OR2_21519 (N26512, N24310, N26107);
or OR4_21520 (N26516, N24316, N26111, N26112, N26113);
nor N2OR3_21521 (N26526, N24316, N26114, N26115);
or OR4_21522 (N26536, N24336, N26131, N26132, N26133);
or OR5_21523 (N26539, N24332, N26124, N26125, N26126, N26127);
nor N2OR3_21524 (N26553, N24336, N26134, N26135);
nor N2OR4_21525 (N26556, N24332, N26128, N26129, N26130);
or OR4_21526 (N26566, N24375, N25117, N26143, N26144);
nor N2OR3_21527 (N26569, N24375, N25118, N26145);
or OR3_21528 (N26572, N24379, N26146, N26147);
nor N2OR2_21529 (N26575, N24379, N26148);
or OR5_21530 (N26580, N24067, N25954, N26156, N26157, N26158);
or OR4_21531 (N26584, N24396, N26159, N26160, N26161);
or OR3_21532 (N26587, N24400, N26162, N26163);
or OR4_21533 (N26592, N24436, N25132, N26171, N26172);
nor N2OR3_21534 (N26599, N24436, N25133, N26173);
or OR4_21535 (N26606, N24456, N26187, N26188, N26189);
or OR5_21536 (N26609, N24080, N26005, N26182, N26183, N26184);
nor N2OR3_21537 (N26619, N24456, N26190, N26191);
nor N2OR4_21538 (N26622, N24080, N26006, N26185, N26186);
nand NAND2_21539 (N26630, N25739, N26373);
nand NAND2_21540 (N26631, N25736, N26374);
nand NAND2_21541 (N26632, N25745, N26375);
nand NAND2_21542 (N26633, N25742, N26376);
nand NAND2_21543 (N26634, N26377, N26066);
nand NAND2_21544 (N26637, N26069, N26378);
not NOT1_21545 (N26640, N26164);
and AND2_21546 (N26641, N26108, N26117);
and AND2_21547 (N26643, N26140, N26149);
and AND2_21548 (N26646, N26168, N26175);
and AND2_21549 (N26648, N26080, N26091);
nand NAND2_21550 (N26650, N26238, N22637);
not NOT1_21551 (N26651, N26238);
not NOT1_21552 (N26653, N26241);
not NOT1_21553 (N26655, N26244);
not NOT1_21554 (N26657, N26247);
not NOT1_21555 (N26659, N26250);
nand NAND2_21556 (N26660, N26253, N25087);
not NOT1_21557 (N26661, N26253);
nand NAND2_21558 (N26662, N26256, N25469);
not NOT1_21559 (N26663, N26256);
and AND2_21560 (N26664, N26091, N24);
not NOT1_21561 (N26666, N26259);
not NOT1_21562 (N26668, N26262);
not NOT1_21563 (N26670, N26265);
not NOT1_21564 (N26672, N26268);
not NOT1_21565 (N26675, N26117);
not NOT1_21566 (N26680, N26280);
not NOT1_21567 (N26681, N26292);
not NOT1_21568 (N26682, N26307);
not NOT1_21569 (N26683, N26310);
nand NAND2_21570 (N26689, N26325, N25120);
not NOT1_21571 (N26690, N26325);
nand NAND2_21572 (N26691, N26328, N25622);
not NOT1_21573 (N26692, N26328);
and AND2_21574 (N26693, N26149, N254);
not NOT1_21575 (N26695, N26331);
not NOT1_21576 (N26698, N26335);
nand NAND2_21577 (N26699, N26338, N25956);
not NOT1_21578 (N26700, N26338);
not NOT1_21579 (N26703, N26175);
not NOT1_21580 (N26708, N26209);
not NOT1_21581 (N26709, N26212);
not NOT1_21582 (N26710, N26215);
not NOT1_21583 (N26711, N26218);
and AND3_21584 (N26712, N25696, N25692, N26209);
and AND3_21585 (N26713, N26200, N26197, N26212);
and AND3_21586 (N26714, N25707, N25703, N26215);
and AND3_21587 (N26715, N26206, N26203, N26218);
buf BUFF1_21588 (N26716, N26466);
and AND3_21589 (N26718, N26164, N21777, N23130);
and AND3_21590 (N26719, N25150, N25315, N26469);
and AND3_21591 (N26720, N24524, N26025, N26470);
and AND3_21592 (N26721, N25157, N25324, N26471);
and AND3_21593 (N26722, N24532, N26028, N26472);
nand NAND2_21594 (N26724, N26477, N26235);
not NOT1_21595 (N26739, N26271);
not NOT1_21596 (N26740, N26274);
not NOT1_21597 (N26741, N26277);
not NOT1_21598 (N26744, N26283);
not NOT1_21599 (N26745, N26286);
not NOT1_21600 (N26746, N26289);
not NOT1_21601 (N26751, N26295);
not NOT1_21602 (N26752, N26298);
not NOT1_21603 (N26753, N26301);
not NOT1_21604 (N26754, N26304);
not NOT1_21605 (N26755, N26322);
not NOT1_21606 (N26760, N26313);
not NOT1_21607 (N26761, N26316);
not NOT1_21608 (N26762, N26319);
not NOT1_21609 (N26772, N26341);
not NOT1_21610 (N26773, N26344);
not NOT1_21611 (N26776, N26347);
not NOT1_21612 (N26777, N26350);
not NOT1_21613 (N26782, N26353);
not NOT1_21614 (N26783, N26356);
not NOT1_21615 (N26784, N26359);
not NOT1_21616 (N26785, N26370);
not NOT1_21617 (N26790, N26364);
not NOT1_21618 (N26791, N26367);
nand NAND2_21619 (N26792, N26630, N26631);
nand NAND2_21620 (N26795, N26632, N26633);
and AND2_21621 (N26801, N26108, N26415);
and AND2_21622 (N26802, N26427, N26140);
and AND2_21623 (N26803, N26397, N26080);
and AND2_21624 (N26804, N26168, N26441);
not NOT1_21625 (N26805, N26466);
nand NAND2_21626 (N26806, N21851, N26651);
not NOT1_21627 (N26807, N26482);
nand NAND2_21628 (N26808, N26482, N26653);
not NOT1_21629 (N26809, N26486);
nand NAND2_21630 (N26810, N26486, N26655);
not NOT1_21631 (N26811, N26490);
nand NAND2_21632 (N26812, N26490, N26657);
not NOT1_21633 (N26813, N26494);
nand NAND2_21634 (N26814, N26494, N26659);
nand NAND2_21635 (N26815, N24575, N26661);
nand NAND2_21636 (N26816, N25169, N26663);
or OR2_21637 (N26817, N26397, N26664);
not NOT1_21638 (N26823, N26500);
nand NAND2_21639 (N26824, N26500, N26666);
not NOT1_21640 (N26825, N26504);
nand NAND2_21641 (N26826, N26504, N26668);
not NOT1_21642 (N26827, N26508);
nand NAND2_21643 (N26828, N26508, N26670);
not NOT1_21644 (N26829, N26512);
nand NAND2_21645 (N26830, N26512, N26672);
not NOT1_21646 (N26831, N26415);
not NOT1_21647 (N26834, N26566);
nand NAND2_21648 (N26835, N26566, N25618);
not NOT1_21649 (N26836, N26569);
nand NAND2_21650 (N26837, N26569, N25619);
not NOT1_21651 (N26838, N26572);
nand NAND2_21652 (N26839, N26572, N25620);
not NOT1_21653 (N26840, N26575);
nand NAND2_21654 (N26841, N26575, N25621);
nand NAND2_21655 (N26842, N24627, N26690);
nand NAND2_21656 (N26843, N25195, N26692);
or OR2_21657 (N26844, N26427, N26693);
not NOT1_21658 (N26850, N26580);
nand NAND2_21659 (N26851, N26580, N26695);
not NOT1_21660 (N26852, N26584);
nand NAND2_21661 (N26853, N26584, N26434);
not NOT1_21662 (N26854, N26587);
nand NAND2_21663 (N26855, N26587, N26698);
nand NAND2_21664 (N26856, N25346, N26700);
not NOT1_21665 (N26857, N26441);
and AND3_21666 (N26860, N26197, N25696, N26708);
and AND3_21667 (N26861, N25692, N26200, N26709);
and AND3_21668 (N26862, N26203, N25707, N26710);
and AND3_21669 (N26863, N25703, N26206, N26711);
or OR3_21670 (N26866, N24197, N26718, N23785);
nor N2OR2_21671 (N26872, N26719, N26473);
nor N2OR2_21672 (N26873, N26720, N26474);
nor N2OR2_21673 (N26874, N26721, N26475);
nor N2OR2_21674 (N26875, N26722, N26476);
not NOT1_21675 (N26876, N26637);
buf BUFF1_21676 (N26877, N26724);
and AND2_21677 (N26879, N26045, N26478);
and AND2_21678 (N26880, N26478, N2132);
or OR2_21679 (N26881, N26411, N26137);
not NOT1_21680 (N26884, N26516);
not NOT1_21681 (N26885, N26411);
not NOT1_21682 (N26888, N26526);
not NOT1_21683 (N26889, N26536);
nand NAND2_21684 (N26890, N26536, N25176);
or OR2_21685 (N26891, N26419, N26138);
not NOT1_21686 (N26894, N26539);
not NOT1_21687 (N26895, N26553);
nand NAND2_21688 (N26896, N26553, N25728);
not NOT1_21689 (N26897, N26419);
not NOT1_21690 (N26900, N26556);
or OR2_21691 (N26901, N26437, N26193);
not NOT1_21692 (N26904, N26592);
not NOT1_21693 (N26905, N26437);
not NOT1_21694 (N26908, N26599);
or OR2_21695 (N26909, N26445, N26194);
not NOT1_21696 (N26912, N26606);
not NOT1_21697 (N26913, N26609);
not NOT1_21698 (N26914, N26619);
nand NAND2_21699 (N26915, N26619, N25734);
not NOT1_21700 (N26916, N26445);
not NOT1_21701 (N26919, N26622);
not NOT1_21702 (N26922, N26634);
nand NAND2_21703 (N26923, N26634, N26067);
or OR2_21704 (N26924, N26382, N26801);
or OR2_21705 (N26925, N26386, N26802);
or OR2_21706 (N26926, N26388, N26803);
or OR2_21707 (N26927, N26392, N26804);
not NOT1_21708 (N26930, N26724);
nand NAND2_21709 (N26932, N26650, N26806);
nand NAND2_21710 (N26935, N26241, N26807);
nand NAND2_21711 (N26936, N26244, N26809);
nand NAND2_21712 (N26937, N26247, N26811);
nand NAND2_21713 (N26938, N26250, N26813);
nand NAND2_21714 (N26939, N26660, N26815);
nand NAND2_21715 (N26940, N26662, N26816);
nand NAND2_21716 (N26946, N26259, N26823);
nand NAND2_21717 (N26947, N26262, N26825);
nand NAND2_21718 (N26948, N26265, N26827);
nand NAND2_21719 (N26949, N26268, N26829);
nand NAND2_21720 (N26953, N25183, N26834);
nand NAND2_21721 (N26954, N25186, N26836);
nand NAND2_21722 (N26955, N25189, N26838);
nand NAND2_21723 (N26956, N25192, N26840);
nand NAND2_21724 (N26957, N26689, N26842);
nand NAND2_21725 (N26958, N26691, N26843);
nand NAND2_21726 (N26964, N26331, N26850);
nand NAND2_21727 (N26965, N26048, N26852);
nand NAND2_21728 (N26966, N26335, N26854);
nand NAND2_21729 (N26967, N26699, N26856);
nor N2OR2_21730 (N26973, N26860, N26712);
nor N2OR2_21731 (N26974, N26861, N26713);
nor N2OR2_21732 (N26975, N26862, N26714);
nor N2OR2_21733 (N26976, N26863, N26715);
not NOT1_21734 (N26977, N26792);
not NOT1_21735 (N26978, N26795);
or OR2_21736 (N26979, N26879, N26880);
nand NAND2_21737 (N26987, N24608, N26889);
nand NAND2_21738 (N26990, N25177, N26895);
nand NAND2_21739 (N26999, N25217, N26914);
nand NAND2_21740 (N27002, N25377, N26922);
nand NAND2_21741 (N27003, N26873, N26872);
nand NAND2_21742 (N27006, N26875, N26874);
and AND3_21743 (N27011, N26866, N22681, N22692);
and AND3_21744 (N27012, N26866, N22756, N22767);
and AND3_21745 (N27013, N26866, N22779, N22790);
not NOT1_21746 (N27015, N26866);
and AND3_21747 (N27016, N26866, N22801, N22812);
nand NAND2_21748 (N27018, N26935, N26808);
nand NAND2_21749 (N27019, N26936, N26810);
nand NAND2_21750 (N27020, N26937, N26812);
nand NAND2_21751 (N27021, N26938, N26814);
not NOT1_21752 (N27022, N26939);
not NOT1_21753 (N27023, N26817);
nand NAND2_21754 (N27028, N26946, N26824);
nand NAND2_21755 (N27031, N26947, N26826);
nand NAND2_21756 (N27034, N26948, N26828);
nand NAND2_21757 (N27037, N26949, N26830);
and AND2_21758 (N27040, N26817, N26079);
and AND2_21759 (N27041, N26831, N26675);
nand NAND2_21760 (N27044, N26953, N26835);
nand NAND2_21761 (N27045, N26954, N26837);
nand NAND2_21762 (N27046, N26955, N26839);
nand NAND2_21763 (N27047, N26956, N26841);
not NOT1_21764 (N27048, N26957);
not NOT1_21765 (N27049, N26844);
nand NAND2_21766 (N27054, N26964, N26851);
nand NAND2_21767 (N27057, N26965, N26853);
nand NAND2_21768 (N27060, N26966, N26855);
and AND2_21769 (N27064, N26844, N26139);
and AND2_21770 (N27065, N26857, N26703);
not NOT1_21771 (N27072, N26881);
nand NAND2_21772 (N27073, N26881, N25172);
not NOT1_21773 (N27074, N26885);
nand NAND2_21774 (N27075, N26885, N25727);
nand NAND2_21775 (N27076, N26890, N26987);
not NOT1_21776 (N27079, N26891);
nand NAND2_21777 (N27080, N26896, N26990);
not NOT1_21778 (N27083, N26897);
not NOT1_21779 (N27084, N26901);
nand NAND2_21780 (N27085, N26901, N25198);
not NOT1_21781 (N27086, N26905);
nand NAND2_21782 (N27087, N26905, N25731);
not NOT1_21783 (N27088, N26909);
nand NAND2_21784 (N27089, N26909, N26912);
nand NAND2_21785 (N27090, N26915, N26999);
not NOT1_21786 (N27093, N26916);
nand NAND2_21787 (N27094, N26974, N26973);
nand NAND2_21788 (N27097, N26976, N26975);
nand NAND2_21789 (N27101, N27002, N26923);
not NOT1_21790 (N27105, N26932);
not NOT1_21791 (N27110, N26967);
and AND3_21792 (N27114, N26979, N2603, N21755);
not NOT1_21793 (N27115, N27019);
not NOT1_21794 (N27116, N27021);
and AND2_21795 (N27125, N26817, N27018);
and AND2_21796 (N27126, N26817, N27020);
and AND2_21797 (N27127, N26817, N27022);
not NOT1_21798 (N27130, N27045);
not NOT1_21799 (N27131, N27047);
and AND2_21800 (N27139, N26844, N27044);
and AND2_21801 (N27140, N26844, N27046);
and AND2_21802 (N27141, N26844, N27048);
and AND3_21803 (N27146, N26932, N21761, N23108);
and AND3_21804 (N27147, N26967, N21777, N23130);
not NOT1_21805 (N27149, N27003);
not NOT1_21806 (N27150, N27006);
nand NAND2_21807 (N27151, N27006, N26876);
nand NAND2_21808 (N27152, N24605, N27072);
nand NAND2_21809 (N27153, N25173, N27074);
nand NAND2_21810 (N27158, N24646, N27084);
nand NAND2_21811 (N27159, N25205, N27086);
nand NAND2_21812 (N27160, N26606, N27088);
not NOT1_21813 (N27166, N27037);
not NOT1_21814 (N27167, N27034);
not NOT1_21815 (N27168, N27031);
not NOT1_21816 (N27169, N27028);
not NOT1_21817 (N27170, N27060);
not NOT1_21818 (N27171, N27057);
not NOT1_21819 (N27172, N27054);
and AND2_21820 (N27173, N27115, N27023);
and AND2_21821 (N27174, N27116, N27023);
and AND2_21822 (N27175, N26940, N27023);
and AND2_21823 (N27176, N25418, N27023);
not NOT1_21824 (N27177, N27041);
and AND2_21825 (N27178, N27130, N27049);
and AND2_21826 (N27179, N27131, N27049);
and AND2_21827 (N27180, N26958, N27049);
and AND2_21828 (N27181, N25573, N27049);
not NOT1_21829 (N27182, N27065);
not NOT1_21830 (N27183, N27094);
nand NAND2_21831 (N27184, N27094, N26977);
not NOT1_21832 (N27185, N27097);
nand NAND2_21833 (N27186, N27097, N26978);
and AND3_21834 (N27187, N27037, N21761, N23108);
and AND3_21835 (N27188, N27034, N21761, N23108);
and AND3_21836 (N27189, N27031, N21761, N23108);
or OR3_21837 (N27190, N24956, N27146, N23781);
and AND3_21838 (N27196, N27060, N21777, N23130);
and AND3_21839 (N27197, N27057, N21777, N23130);
or OR3_21840 (N27198, N24960, N27147, N23786);
nand NAND2_21841 (N27204, N27101, N27149);
not NOT1_21842 (N27205, N27101);
nand NAND2_21843 (N27206, N26637, N27150);
and AND3_21844 (N27207, N27028, N21793, N23158);
and AND3_21845 (N27208, N27054, N21807, N23180);
nand NAND2_21846 (N27209, N27073, N27152);
nand NAND2_21847 (N27212, N27075, N27153);
not NOT1_21848 (N27215, N27076);
nand NAND2_21849 (N27216, N27076, N27079);
not NOT1_21850 (N27217, N27080);
nand NAND2_21851 (N27218, N27080, N27083);
nand NAND2_21852 (N27219, N27085, N27158);
nand NAND2_21853 (N27222, N27087, N27159);
nand NAND2_21854 (N27225, N27089, N27160);
not NOT1_21855 (N27228, N27090);
nand NAND2_21856 (N27229, N27090, N27093);
or OR2_21857 (N27236, N27173, N27125);
or OR2_21858 (N27239, N27174, N27126);
or OR2_21859 (N27242, N27175, N27127);
or OR2_21860 (N27245, N27176, N27040);
or OR2_21861 (N27250, N27178, N27139);
or OR2_21862 (N27257, N27179, N27140);
or OR2_21863 (N27260, N27180, N27141);
or OR2_21864 (N27263, N27181, N27064);
nand NAND2_21865 (N27268, N26792, N27183);
nand NAND2_21866 (N27269, N26795, N27185);
or OR3_21867 (N27270, N24957, N27187, N23782);
or OR3_21868 (N27276, N24958, N27188, N23783);
or OR3_21869 (N27282, N24959, N27189, N23784);
or OR3_21870 (N27288, N24961, N27196, N23787);
or OR3_21871 (N27294, N23998, N27197, N23788);
nand NAND2_21872 (N27300, N27003, N27205);
nand NAND2_21873 (N27301, N27206, N27151);
or OR3_21874 (N27304, N24980, N27207, N23800);
or OR3_21875 (N27310, N24984, N27208, N23805);
nand NAND2_21876 (N27320, N26891, N27215);
nand NAND2_21877 (N27321, N26897, N27217);
nand NAND2_21878 (N27328, N26916, N27228);
and AND3_21879 (N27338, N27190, N21185, N22692);
and AND3_21880 (N27339, N27198, N22681, N22692);
and AND3_21881 (N27340, N27190, N21247, N22767);
and AND3_21882 (N27341, N27198, N22756, N22767);
and AND3_21883 (N27342, N27190, N21327, N22790);
and AND3_21884 (N27349, N27198, N22779, N22790);
and AND3_21885 (N27357, N27198, N22801, N22812);
not NOT1_21886 (N27363, N27198);
and AND3_21887 (N27364, N27190, N21351, N22812);
not NOT1_21888 (N27365, N27190);
nand NAND2_21889 (N27394, N27268, N27184);
nand NAND2_21890 (N27397, N27269, N27186);
nand NAND2_21891 (N27402, N27204, N27300);
not NOT1_21892 (N27405, N27209);
nand NAND2_21893 (N27406, N27209, N26884);
not NOT1_21894 (N27407, N27212);
nand NAND2_21895 (N27408, N27212, N26888);
nand NAND2_21896 (N27409, N27320, N27216);
nand NAND2_21897 (N27412, N27321, N27218);
not NOT1_21898 (N27415, N27219);
nand NAND2_21899 (N27416, N27219, N26904);
not NOT1_21900 (N27417, N27222);
nand NAND2_21901 (N27418, N27222, N26908);
not NOT1_21902 (N27419, N27225);
nand NAND2_21903 (N27420, N27225, N26913);
nand NAND2_21904 (N27421, N27328, N27229);
not NOT1_21905 (N27424, N27245);
not NOT1_21906 (N27425, N27242);
not NOT1_21907 (N27426, N27239);
not NOT1_21908 (N27427, N27236);
not NOT1_21909 (N27428, N27263);
not NOT1_21910 (N27429, N27260);
not NOT1_21911 (N27430, N27257);
not NOT1_21912 (N27431, N27250);
not NOT1_21913 (N27432, N27250);
and AND3_21914 (N27433, N27310, N22653, N22664);
and AND3_21915 (N27434, N27304, N21161, N22664);
or OR4_21916 (N27435, N27011, N27338, N23621, N22591);
and AND3_21917 (N27436, N27270, N21185, N22692);
and AND3_21918 (N27437, N27288, N22681, N22692);
and AND3_21919 (N27438, N27276, N21185, N22692);
and AND3_21920 (N27439, N27294, N22681, N22692);
and AND3_21921 (N27440, N27282, N21185, N22692);
and AND3_21922 (N27441, N27310, N22728, N22739);
and AND3_21923 (N27442, N27304, N21223, N22739);
or OR4_21924 (N27443, N27012, N27340, N23632, N22600);
and AND3_21925 (N27444, N27270, N21247, N22767);
and AND3_21926 (N27445, N27288, N22756, N22767);
and AND3_21927 (N27446, N27276, N21247, N22767);
and AND3_21928 (N27447, N27294, N22756, N22767);
and AND3_21929 (N27448, N27282, N21247, N22767);
or OR4_21930 (N27449, N27013, N27342, N23641, N22605);
and AND3_21931 (N27450, N27310, N23041, N23052);
and AND3_21932 (N27451, N27304, N21697, N23052);
and AND3_21933 (N27452, N27294, N22779, N22790);
and AND3_21934 (N27453, N27282, N21327, N22790);
and AND3_21935 (N27454, N27288, N22779, N22790);
and AND3_21936 (N27455, N27276, N21327, N22790);
and AND3_21937 (N27456, N27270, N21327, N22790);
and AND3_21938 (N27457, N27310, N23075, N23086);
and AND3_21939 (N27458, N27304, N21731, N23086);
and AND3_21940 (N27459, N27294, N22801, N22812);
and AND3_21941 (N27460, N27282, N21351, N22812);
and AND3_21942 (N27461, N27288, N22801, N22812);
and AND3_21943 (N27462, N27276, N21351, N22812);
and AND3_21944 (N27463, N27270, N21351, N22812);
and AND3_21945 (N27464, N27250, N2603, N2599);
not NOT1_21946 (N27465, N27310);
not NOT1_21947 (N27466, N27294);
not NOT1_21948 (N27467, N27288);
not NOT1_21949 (N27468, N27301);
or OR4_21950 (N27469, N27016, N27364, N23660, N22626);
not NOT1_21951 (N27470, N27304);
not NOT1_21952 (N27471, N27282);
not NOT1_21953 (N27472, N27276);
not NOT1_21954 (N27473, N27270);
buf BUFF1_21955 (N27474, N27394);
buf BUFF1_21956 (N27476, N27397);
and AND2_21957 (N27479, N27301, N23068);
and AND3_21958 (N27481, N27245, N21793, N23158);
and AND3_21959 (N27482, N27242, N21793, N23158);
and AND3_21960 (N27483, N27239, N21793, N23158);
and AND3_21961 (N27484, N27236, N21793, N23158);
and AND3_21962 (N27485, N27263, N21807, N23180);
and AND3_21963 (N27486, N27260, N21807, N23180);
and AND3_21964 (N27487, N27257, N21807, N23180);
and AND3_21965 (N27488, N27250, N21807, N23180);
nand NAND2_21966 (N27489, N26979, N27250);
nand NAND2_21967 (N27492, N26516, N27405);
nand NAND2_21968 (N27493, N26526, N27407);
nand NAND2_21969 (N27498, N26592, N27415);
nand NAND2_21970 (N27499, N26599, N27417);
nand NAND2_21971 (N27500, N26609, N27419);
and AND9_21972 (N27503, N27105, N27166, N27167, N27168, N27169, N27424, N27425, N27426, N27427);
and AND9_21973 (N27504, N26640, N27110, N27170, N27171, N27172, N27428, N27429, N27430, N27431);
or OR4_21974 (N27505, N27433, N27434, N23616, N22585);
and AND2_21975 (N27506, N27435, N22675);
or OR4_21976 (N27507, N27339, N27436, N23622, N22592);
or OR4_21977 (N27508, N27437, N27438, N23623, N22593);
or OR4_21978 (N27509, N27439, N27440, N23624, N22594);
or OR4_21979 (N27510, N27441, N27442, N23627, N22595);
and AND2_21980 (N27511, N27443, N22750);
or OR4_21981 (N27512, N27341, N27444, N23633, N22601);
or OR4_21982 (N27513, N27445, N27446, N23634, N22602);
or OR4_21983 (N27514, N27447, N27448, N23635, N22603);
or OR4_21984 (N27515, N27450, N27451, N23646, N22610);
or OR4_21985 (N27516, N27452, N27453, N23647, N22611);
or OR4_21986 (N27517, N27454, N27455, N23648, N22612);
or OR4_21987 (N27518, N27349, N27456, N23649, N22613);
or OR4_21988 (N27519, N27457, N27458, N23654, N22618);
or OR4_21989 (N27520, N27459, N27460, N23655, N22619);
or OR4_21990 (N27521, N27461, N27462, N23656, N22620);
or OR4_21991 (N27522, N27357, N27463, N23657, N22621);
or OR4_21992 (N27525, N24741, N27114, N22624, N27464);
and AND3_21993 (N27526, N27468, N23119, N23130);
not NOT1_21994 (N27527, N27394);
not NOT1_21995 (N27528, N27397);
not NOT1_21996 (N27529, N27402);
and AND2_21997 (N27530, N27402, N23068);
or OR3_21998 (N27531, N24981, N27481, N23801);
or OR3_21999 (N27537, N24982, N27482, N23802);
or OR3_22000 (N27543, N24983, N27483, N23803);
or OR3_22001 (N27549, N25165, N27484, N23804);
or OR3_22002 (N27555, N24985, N27485, N23806);
or OR3_22003 (N27561, N24986, N27486, N23807);
or OR3_22004 (N27567, N24547, N27487, N23808);
or OR3_22005 (N27573, N24987, N27488, N23809);
nand NAND2_22006 (N27579, N27492, N27406);
nand NAND2_22007 (N27582, N27493, N27408);
not NOT1_22008 (N27585, N27409);
nand NAND2_22009 (N27586, N27409, N26894);
not NOT1_22010 (N27587, N27412);
nand NAND2_22011 (N27588, N27412, N26900);
nand NAND2_22012 (N27589, N27498, N27416);
nand NAND2_22013 (N27592, N27499, N27418);
nand NAND2_22014 (N27595, N27500, N27420);
not NOT1_22015 (N27598, N27421);
nand NAND2_22016 (N27599, N27421, N26919);
and AND2_22017 (N27600, N27505, N22647);
and AND2_22018 (N27601, N27507, N22675);
and AND2_22019 (N27602, N27508, N22675);
and AND2_22020 (N27603, N27509, N22675);
and AND2_22021 (N27604, N27510, N22722);
and AND2_22022 (N27605, N27512, N22750);
and AND2_22023 (N27606, N27513, N22750);
and AND2_22024 (N27607, N27514, N22750);
and AND2_22025 (N27624, N26979, N27489);
and AND2_22026 (N27625, N27489, N27250);
and AND2_22027 (N27626, N21149, N27525);
and AND5_22028 (N27631, N2562, N27527, N27528, N26805, N26930);
and AND3_22029 (N27636, N27529, N23097, N23108);
nand NAND2_22030 (N27657, N26539, N27585);
nand NAND2_22031 (N27658, N26556, N27587);
nand NAND2_22032 (N27665, N26622, N27598);
and AND3_22033 (N27666, N27555, N22653, N22664);
and AND3_22034 (N27667, N27531, N21161, N22664);
and AND3_22035 (N27668, N27561, N22653, N22664);
and AND3_22036 (N27669, N27537, N21161, N22664);
and AND3_22037 (N27670, N27567, N22653, N22664);
and AND3_22038 (N27671, N27543, N21161, N22664);
and AND3_22039 (N27672, N27573, N22653, N22664);
and AND3_22040 (N27673, N27549, N21161, N22664);
and AND3_22041 (N27674, N27555, N22728, N22739);
and AND3_22042 (N27675, N27531, N21223, N22739);
and AND3_22043 (N27676, N27561, N22728, N22739);
and AND3_22044 (N27677, N27537, N21223, N22739);
and AND3_22045 (N27678, N27567, N22728, N22739);
and AND3_22046 (N27679, N27543, N21223, N22739);
and AND3_22047 (N27680, N27573, N22728, N22739);
and AND3_22048 (N27681, N27549, N21223, N22739);
and AND3_22049 (N27682, N27573, N23075, N23086);
and AND3_22050 (N27683, N27549, N21731, N23086);
and AND3_22051 (N27684, N27573, N23041, N23052);
and AND3_22052 (N27685, N27549, N21697, N23052);
and AND3_22053 (N27686, N27567, N23041, N23052);
and AND3_22054 (N27687, N27543, N21697, N23052);
and AND3_22055 (N27688, N27561, N23041, N23052);
and AND3_22056 (N27689, N27537, N21697, N23052);
and AND3_22057 (N27690, N27555, N23041, N23052);
and AND3_22058 (N27691, N27531, N21697, N23052);
and AND3_22059 (N27692, N27567, N23075, N23086);
and AND3_22060 (N27693, N27543, N21731, N23086);
and AND3_22061 (N27694, N27561, N23075, N23086);
and AND3_22062 (N27695, N27537, N21731, N23086);
and AND3_22063 (N27696, N27555, N23075, N23086);
and AND3_22064 (N27697, N27531, N21731, N23086);
or OR2_22065 (N27698, N27624, N27625);
not NOT1_22066 (N27699, N27573);
not NOT1_22067 (N27700, N27567);
not NOT1_22068 (N27701, N27561);
not NOT1_22069 (N27702, N27555);
and AND3_22070 (N27703, N21156, N27631, N2245);
not NOT1_22071 (N27704, N27549);
not NOT1_22072 (N27705, N27543);
not NOT1_22073 (N27706, N27537);
not NOT1_22074 (N27707, N27531);
not NOT1_22075 (N27708, N27579);
nand NAND2_22076 (N27709, N27579, N26739);
not NOT1_22077 (N27710, N27582);
nand NAND2_22078 (N27711, N27582, N26744);
nand NAND2_22079 (N27712, N27657, N27586);
nand NAND2_22080 (N27715, N27658, N27588);
not NOT1_22081 (N27718, N27589);
nand NAND2_22082 (N27719, N27589, N26772);
not NOT1_22083 (N27720, N27592);
nand NAND2_22084 (N27721, N27592, N26776);
not NOT1_22085 (N27722, N27595);
nand NAND2_22086 (N27723, N27595, N25733);
nand NAND2_22087 (N27724, N27665, N27599);
or OR4_22088 (N27727, N27666, N27667, N23617, N22586);
or OR4_22089 (N27728, N27668, N27669, N23618, N22587);
or OR4_22090 (N27729, N27670, N27671, N23619, N22588);
or OR4_22091 (N27730, N27672, N27673, N23620, N22589);
or OR4_22092 (N27731, N27674, N27675, N23628, N22596);
or OR4_22093 (N27732, N27676, N27677, N23629, N22597);
or OR4_22094 (N27733, N27678, N27679, N23630, N22598);
or OR4_22095 (N27734, N27680, N27681, N23631, N22599);
or OR4_22096 (N27735, N27682, N27683, N23638, N22604);
or OR4_22097 (N27736, N27684, N27685, N23642, N22606);
or OR4_22098 (N27737, N27686, N27687, N23643, N22607);
or OR4_22099 (N27738, N27688, N27689, N23644, N22608);
or OR4_22100 (N27739, N27690, N27691, N23645, N22609);
or OR4_22101 (N27740, N27692, N27693, N23651, N22615);
or OR4_22102 (N27741, N27694, N27695, N23652, N22616);
or OR4_22103 (N27742, N27696, N27697, N23653, N22617);
nand NAND2_22104 (N27743, N26271, N27708);
nand NAND2_22105 (N27744, N26283, N27710);
nand NAND2_22106 (N27749, N26341, N27718);
nand NAND2_22107 (N27750, N26347, N27720);
nand NAND2_22108 (N27751, N25214, N27722);
and AND2_22109 (N27754, N27727, N22647);
and AND2_22110 (N27755, N27728, N22647);
and AND2_22111 (N27756, N27729, N22647);
and AND2_22112 (N27757, N27730, N22647);
and AND2_22113 (N27758, N27731, N22722);
and AND2_22114 (N27759, N27732, N22722);
and AND2_22115 (N27760, N27733, N22722);
and AND2_22116 (N27761, N27734, N22722);
nand NAND2_22117 (N27762, N27743, N27709);
nand NAND2_22118 (N27765, N27744, N27711);
not NOT1_22119 (N27768, N27712);
nand NAND2_22120 (N27769, N27712, N26751);
not NOT1_22121 (N27770, N27715);
nand NAND2_22122 (N27771, N27715, N26760);
nand NAND2_22123 (N27772, N27749, N27719);
nand NAND2_22124 (N27775, N27750, N27721);
nand NAND2_22125 (N27778, N27751, N27723);
not NOT1_22126 (N27781, N27724);
nand NAND2_22127 (N27782, N27724, N25735);
nand NAND2_22128 (N27787, N26295, N27768);
nand NAND2_22129 (N27788, N26313, N27770);
nand NAND2_22130 (N27795, N25220, N27781);
not NOT1_22131 (N27796, N27762);
nand NAND2_22132 (N27797, N27762, N26740);
not NOT1_22133 (N27798, N27765);
nand NAND2_22134 (N27799, N27765, N26745);
nand NAND2_22135 (N27800, N27787, N27769);
nand NAND2_22136 (N27803, N27788, N27771);
not NOT1_22137 (N27806, N27772);
nand NAND2_22138 (N27807, N27772, N26773);
not NOT1_22139 (N27808, N27775);
nand NAND2_22140 (N27809, N27775, N26777);
not NOT1_22141 (N27810, N27778);
nand NAND2_22142 (N27811, N27778, N26782);
nand NAND2_22143 (N27812, N27795, N27782);
nand NAND2_22144 (N27815, N26274, N27796);
nand NAND2_22145 (N27816, N26286, N27798);
nand NAND2_22146 (N27821, N26344, N27806);
nand NAND2_22147 (N27822, N26350, N27808);
nand NAND2_22148 (N27823, N26353, N27810);
nand NAND2_22149 (N27826, N27815, N27797);
nand NAND2_22150 (N27829, N27816, N27799);
not NOT1_22151 (N27832, N27800);
nand NAND2_22152 (N27833, N27800, N26752);
not NOT1_22153 (N27834, N27803);
nand NAND2_22154 (N27835, N27803, N26761);
nand NAND2_22155 (N27836, N27821, N27807);
nand NAND2_22156 (N27839, N27822, N27809);
nand NAND2_22157 (N27842, N27823, N27811);
not NOT1_22158 (N27845, N27812);
nand NAND2_22159 (N27846, N27812, N26790);
nand NAND2_22160 (N27851, N26298, N27832);
nand NAND2_22161 (N27852, N26316, N27834);
nand NAND2_22162 (N27859, N26364, N27845);
not NOT1_22163 (N27860, N27826);
nand NAND2_22164 (N27861, N27826, N26741);
not NOT1_22165 (N27862, N27829);
nand NAND2_22166 (N27863, N27829, N26746);
nand NAND2_22167 (N27864, N27851, N27833);
nand NAND2_22168 (N27867, N27852, N27835);
not NOT1_22169 (N27870, N27836);
nand NAND2_22170 (N27871, N27836, N25730);
not NOT1_22171 (N27872, N27839);
nand NAND2_22172 (N27873, N27839, N25732);
not NOT1_22173 (N27874, N27842);
nand NAND2_22174 (N27875, N27842, N26783);
nand NAND2_22175 (N27876, N27859, N27846);
nand NAND2_22176 (N27879, N26277, N27860);
nand NAND2_22177 (N27880, N26289, N27862);
nand NAND2_22178 (N27885, N25199, N27870);
nand NAND2_22179 (N27886, N25208, N27872);
nand NAND2_22180 (N27887, N26356, N27874);
nand NAND2_22181 (N27890, N27879, N27861);
nand NAND2_22182 (N27893, N27880, N27863);
not NOT1_22183 (N27896, N27864);
nand NAND2_22184 (N27897, N27864, N26753);
not NOT1_22185 (N27898, N27867);
nand NAND2_22186 (N27899, N27867, N26762);
nand NAND2_22187 (N27900, N27885, N27871);
nand NAND2_22188 (N27903, N27886, N27873);
nand NAND2_22189 (N27906, N27887, N27875);
not NOT1_22190 (N27909, N27876);
nand NAND2_22191 (N27910, N27876, N26791);
nand NAND2_22192 (N27917, N26301, N27896);
nand NAND2_22193 (N27918, N26319, N27898);
nand NAND2_22194 (N27923, N26367, N27909);
not NOT1_22195 (N27924, N27890);
nand NAND2_22196 (N27925, N27890, N26680);
not NOT1_22197 (N27926, N27893);
nand NAND2_22198 (N27927, N27893, N26681);
not NOT1_22199 (N27928, N27900);
nand NAND2_22200 (N27929, N27900, N25690);
not NOT1_22201 (N27930, N27903);
nand NAND2_22202 (N27931, N27903, N25691);
nand NAND2_22203 (N27932, N27917, N27897);
nand NAND2_22204 (N27935, N27918, N27899);
not NOT1_22205 (N27938, N27906);
nand NAND2_22206 (N27939, N27906, N26784);
nand NAND2_22207 (N27940, N27923, N27910);
nand NAND2_22208 (N27943, N26280, N27924);
nand NAND2_22209 (N27944, N26292, N27926);
nand NAND2_22210 (N27945, N25202, N27928);
nand NAND2_22211 (N27946, N25211, N27930);
nand NAND2_22212 (N27951, N26359, N27938);
nand NAND2_22213 (N27954, N27943, N27925);
nand NAND2_22214 (N27957, N27944, N27927);
nand NAND2_22215 (N27960, N27945, N27929);
nand NAND2_22216 (N27963, N27946, N27931);
not NOT1_22217 (N27966, N27932);
nand NAND2_22218 (N27967, N27932, N26754);
not NOT1_22219 (N27968, N27935);
nand NAND2_22220 (N27969, N27935, N26755);
nand NAND2_22221 (N27970, N27951, N27939);
not NOT1_22222 (N27973, N27940);
nand NAND2_22223 (N27974, N27940, N26785);
nand NAND2_22224 (N27984, N26304, N27966);
nand NAND2_22225 (N27985, N26322, N27968);
nand NAND2_22226 (N27987, N26370, N27973);
and AND3_22227 (N27988, N27957, N26831, N21157);
and AND3_22228 (N27989, N27954, N26415, N21157);
and AND3_22229 (N27990, N27957, N27041, N2566);
and AND3_22230 (N27991, N27954, N27177, N2566);
not NOT1_22231 (N27992, N27970);
nand NAND2_22232 (N27993, N27970, N26448);
and AND3_22233 (N27994, N27963, N26857, N21219);
and AND3_22234 (N27995, N27960, N26441, N21219);
and AND3_22235 (N27996, N27963, N27065, N2583);
and AND3_22236 (N27997, N27960, N27182, N2583);
nand NAND2_22237 (N27998, N27984, N27967);
nand NAND2_22238 (N28001, N27985, N27969);
nand NAND2_22239 (N28004, N27987, N27974);
nand NAND2_22240 (N28009, N26051, N27992);
or OR4_22241 (N28013, N27988, N27989, N27990, N27991);
or OR4_22242 (N28017, N27994, N27995, N27996, N27997);
not NOT1_22243 (N28020, N27998);
nand NAND2_22244 (N28021, N27998, N26682);
not NOT1_22245 (N28022, N28001);
nand NAND2_22246 (N28023, N28001, N26683);
nand NAND2_22247 (N28025, N28009, N27993);
not NOT1_22248 (N28026, N28004);
nand NAND2_22249 (N28027, N28004, N26449);
nand NAND2_22250 (N28031, N26307, N28020);
nand NAND2_22251 (N28032, N26310, N28022);
not NOT1_22252 (N28033, N28013);
nand NAND2_22253 (N28034, N26054, N28026);
and AND2_22254 (N28035, N2583, N28025);
not NOT1_22255 (N28036, N28017);
nand NAND2_22256 (N28037, N28031, N28021);
nand NAND2_22257 (N28038, N28032, N28023);
nand NAND2_22258 (N28039, N28034, N28027);
not NOT1_22259 (N28040, N28038);
and AND2_22260 (N28041, N2566, N28037);
not NOT1_22261 (N28042, N28039);
and AND2_22262 (N28043, N28040, N21157);
and AND2_22263 (N28044, N28042, N21219);
or OR2_22264 (N28045, N28043, N28041);
or OR2_22265 (N28048, N28044, N28035);
nand NAND2_22266 (N28055, N28045, N28033);
not NOT1_22267 (N28056, N28045);
nand NAND2_22268 (N28057, N28048, N28036);
not NOT1_22269 (N28058, N28048);
nand NAND2_22270 (N28059, N28013, N28056);
nand NAND2_22271 (N28060, N28017, N28058);
nand NAND2_22272 (N28061, N28055, N28059);
nand NAND2_22273 (N28064, N28057, N28060);
and AND3_22274 (N28071, N28064, N21777, N23130);
and AND3_22275 (N28072, N28061, N21761, N23108);
not NOT1_22276 (N28073, N28061);
not NOT1_22277 (N28074, N28064);
or OR4_22278 (N28075, N27526, N28071, N23659, N22625);
or OR4_22279 (N28076, N27636, N28072, N23661, N22627);
and AND2_22280 (N28077, N28073, N21727);
and AND2_22281 (N28078, N28074, N21727);
or OR2_22282 (N28079, N27530, N28077);
or OR2_22283 (N28082, N27479, N28078);
and AND2_22284 (N28089, N28079, N23063);
and AND2_22285 (N28090, N28082, N23063);
and AND2_22286 (N28091, N28079, N23063);
and AND2_22287 (N28092, N28082, N23063);
or OR2_22288 (N28093, N28089, N23071);
or OR2_22289 (N28096, N28090, N23072);
or OR2_22290 (N28099, N28091, N23073);
or OR2_22291 (N28102, N28092, N23074);
and AND3_22292 (N28113, N28102, N22779, N22790);
and AND3_22293 (N28114, N28099, N21327, N22790);
and AND3_22294 (N28115, N28102, N22801, N22812);
and AND3_22295 (N28116, N28099, N21351, N22812);
and AND3_22296 (N28117, N28096, N22681, N22692);
and AND3_22297 (N28118, N28093, N21185, N22692);
and AND3_22298 (N28119, N28096, N22756, N22767);
and AND3_22299 (N28120, N28093, N21247, N22767);
or OR4_22300 (N28121, N28117, N28118, N23662, N22703);
or OR4_22301 (N28122, N28119, N28120, N23663, N22778);
or OR4_22302 (N28123, N28113, N28114, N23650, N22614);
or OR4_22303 (N28124, N28115, N28116, N23658, N22622);
and AND2_22304 (N28125, N28121, N22675);
and AND2_22305 (N28126, N28122, N22750);
not NOT1_22306 (N28127, N28125);
not NOT1_22307 (N28128, N28126);

endmodule
