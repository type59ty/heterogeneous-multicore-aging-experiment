`timescale 1ns/10ps

`define cycle 10.0
`define terminate_cycle 400000//200000 // Modify your terminate ycle here

module b22_ras_testfixture;

`define in_file "b22_ras/rand_input_vector_b22_ras_0.out"
`define out_file "b22_ras/rand_output_vector_b22_ras_0.out"

parameter vec_width = 767;
parameter vec_length = 7;

reg clk = 0;


reg [vec_width-1:0] input_vec_mem [0:vec_length-1];
reg [vec_width-1:0] vec;

wire sub_1596_u4, sub_1596_u62, sub_1596_u63, sub_1596_u64, sub_1596_u65, sub_1596_u66, sub_1596_u67, sub_1596_u68, sub_1596_u69, sub_1596_u70, sub_1596_u54, sub_1596_u55, sub_1596_u56, sub_1596_u57, sub_1596_u58, sub_1596_u59, sub_1596_u60, sub_1596_u61, sub_1596_u5, sub_1596_u53, u29, u28, p1_u3355, p1_u3354, p1_u3353, p1_u3352, p1_u3351, p1_u3350, p1_u3349, p1_u3348, p1_u3347, p1_u3346, p1_u3345, p1_u3344, p1_u3343, p1_u3342, p1_u3341, p1_u3340, p1_u3339, p1_u3338, p1_u3337, p1_u3336, p1_u3335, p1_u3334, p1_u3333, p1_u3332, p1_u3331, p1_u3330, p1_u3329, p1_u3328, p1_u3327, p1_u3326, p1_u3325, p1_u3324, p1_u3445, p1_u3446, p1_u3323, p1_u3322, p1_u3321, p1_u3320, p1_u3319, p1_u3318, p1_u3317, p1_u3316, p1_u3315, p1_u3314, p1_u3313, p1_u3312, p1_u3311, p1_u3310, p1_u3309, p1_u3308, p1_u3307, p1_u3306, p1_u3305, p1_u3304, p1_u3303, p1_u3302, p1_u3301, p1_u3300, p1_u3299, p1_u3298, p1_u3297, p1_u3296, p1_u3295, p1_u3294, p1_u3459, p1_u3462, p1_u3465, p1_u3468, p1_u3471, p1_u3474, p1_u3477, p1_u3480, p1_u3483, p1_u3486, p1_u3489, p1_u3492, p1_u3495, p1_u3498, p1_u3501, p1_u3504, p1_u3507, p1_u3510, p1_u3513, p1_u3515, p1_u3516, p1_u3517, p1_u3518, p1_u3519, p1_u3520, p1_u3521, p1_u3522, p1_u3523, p1_u3524, p1_u3525, p1_u3526, p1_u3527, p1_u3528, p1_u3529, p1_u3530, p1_u3531, p1_u3532, p1_u3533, p1_u3534, p1_u3535, p1_u3536, p1_u3537, p1_u3538, p1_u3539, p1_u3540, p1_u3541, p1_u3542, p1_u3543, p1_u3544, p1_u3545, p1_u3546, p1_u3547, p1_u3548, p1_u3549, p1_u3550, p1_u3551, p1_u3552, p1_u3553, p1_u3554, p1_u3555, p1_u3556, p1_u3557, p1_u3558, p1_u3559, p1_u3293, p1_u3292, p1_u3291, p1_u3290, p1_u3289, p1_u3288, p1_u3287, p1_u3286, p1_u3285, p1_u3284, p1_u3283, p1_u3282, p1_u3281, p1_u3280, p1_u3279, p1_u3278, p1_u3277, p1_u3276, p1_u3275, p1_u3274, p1_u3273, p1_u3272, p1_u3271, p1_u3270, p1_u3269, p1_u3268, p1_u3267, p1_u3266, p1_u3265, p1_u3356, p1_u3264, p1_u3263, p1_u3262, p1_u3261, p1_u3260, p1_u3259, p1_u3258, p1_u3257, p1_u3256, p1_u3255, p1_u3254, p1_u3253, p1_u3252, p1_u3251, p1_u3250, p1_u3249, p1_u3248, p1_u3247, p1_u3246, p1_u3245, p1_u3244, p1_u3243, p1_u3560, p1_u3561, p1_u3562, p1_u3563, p1_u3564, p1_u3565, p1_u3566, p1_u3567, p1_u3568, p1_u3569, p1_u3570, p1_u3571, p1_u3572, p1_u3573, p1_u3574, p1_u3575, p1_u3576, p1_u3577, p1_u3578, p1_u3579, p1_u3580, p1_u3581, p1_u3582, p1_u3583, p1_u3584, p1_u3585, p1_u3586, p1_u3587, p1_u3588, p1_u3589, p1_u3590, p1_u3591, p1_u3242, p1_u3241, p1_u3240, p1_u3239, p1_u3238, p1_u3237, p1_u3236, p1_u3235, p1_u3234, p1_u3233, p1_u3232, p1_u3231, p1_u3230, p1_u3229, p1_u3228, p1_u3227, p1_u3226, p1_u3225, p1_u3224, p1_u3223, p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218, p1_u3217, p1_u3216, p1_u3215, p1_u3214, p1_u3213, p1_u3086, p1_u3085, p1_u4016, p2_u3327, p2_u3326, p2_u3325, p2_u3324, p2_u3323, p2_u3322, p2_u3321, p2_u3320, p2_u3319, p2_u3318, p2_u3317, p2_u3316, p2_u3315, p2_u3314, p2_u3313, p2_u3312, p2_u3311, p2_u3310, p2_u3309, p2_u3308, p2_u3307, p2_u3306, p2_u3305, p2_u3304, p2_u3303, p2_u3302, p2_u3301, p2_u3300, p2_u3299, p2_u3298, p2_u3297, p2_u3296, p2_u3416, p2_u3417, p2_u3295, p2_u3294, p2_u3293, p2_u3292, p2_u3291, p2_u3290, p2_u3289, p2_u3288, p2_u3287, p2_u3286, p2_u3285, p2_u3284, p2_u3283, p2_u3282, p2_u3281, p2_u3280, p2_u3279, p2_u3278, p2_u3277, p2_u3276, p2_u3275, p2_u3274, p2_u3273, p2_u3272, p2_u3271, p2_u3270, p2_u3269, p2_u3268, p2_u3267, p2_u3266, p2_u3430, p2_u3433, p2_u3436, p2_u3439, p2_u3442, p2_u3445, p2_u3448, p2_u3451, p2_u3454, p2_u3457, p2_u3460, p2_u3463, p2_u3466, p2_u3469, p2_u3472, p2_u3475, p2_u3478, p2_u3481, p2_u3484, p2_u3486, p2_u3487, p2_u3488, p2_u3489, p2_u3490, p2_u3491, p2_u3492, p2_u3493, p2_u3494, p2_u3495, p2_u3496, p2_u3497, p2_u3498, p2_u3499, p2_u3500, p2_u3501, p2_u3502, p2_u3503, p2_u3504, p2_u3505, p2_u3506, p2_u3507, p2_u3508, p2_u3509, p2_u3510, p2_u3511, p2_u3512, p2_u3513, p2_u3514, p2_u3515, p2_u3516, p2_u3517, p2_u3518, p2_u3519, p2_u3520, p2_u3521, p2_u3522, p2_u3523, p2_u3524, p2_u3525, p2_u3526, p2_u3527, p2_u3528, p2_u3529, p2_u3530, p2_u3265, p2_u3264, p2_u3263, p2_u3262, p2_u3261, p2_u3260, p2_u3259, p2_u3258, p2_u3257, p2_u3256, p2_u3255, p2_u3254, p2_u3253, p2_u3252, p2_u3251, p2_u3250, p2_u3249, p2_u3248, p2_u3247, p2_u3246, p2_u3245, p2_u3244, p2_u3243, p2_u3242, p2_u3241, p2_u3240, p2_u3239, p2_u3238, p2_u3237, p2_u3236, p2_u3235, p2_u3234, p2_u3233, p2_u3232, p2_u3231, p2_u3230, p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225, p2_u3224, p2_u3223, p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218, p2_u3217, p2_u3216, p2_u3215, p2_u3214, p2_u3531, p2_u3532, p2_u3533, p2_u3534, p2_u3535, p2_u3536, p2_u3537, p2_u3538, p2_u3539, p2_u3540, p2_u3541, p2_u3542, p2_u3543, p2_u3544, p2_u3545, p2_u3546, p2_u3547, p2_u3548, p2_u3549, p2_u3550, p2_u3551, p2_u3552, p2_u3553, p2_u3554, p2_u3555, p2_u3556, p2_u3557, p2_u3558, p2_u3559, p2_u3560, p2_u3561, p2_u3562, p2_u3328, p2_u3213, p2_u3212, p2_u3211, p2_u3210, p2_u3209, p2_u3208, p2_u3207, p2_u3206, p2_u3205, p2_u3204, p2_u3203, p2_u3202, p2_u3201, p2_u3200, p2_u3199, p2_u3198, p2_u3197, p2_u3196, p2_u3195, p2_u3194, p2_u3193, p2_u3192, p2_u3191, p2_u3190, p2_u3189, p2_u3188, p2_u3187, p2_u3186, p2_u3185, p2_u3088, p2_u3087, p2_u3947, p3_u3295, p3_u3294, p3_u3293, p3_u3292, p3_u3291, p3_u3290, p3_u3289, p3_u3288, p3_u3287, p3_u3286, p3_u3285, p3_u3284, p3_u3283, p3_u3282, p3_u3281, p3_u3280, p3_u3279, p3_u3278, p3_u3277, p3_u3276, p3_u3275, p3_u3274, p3_u3273, p3_u3272, p3_u3271, p3_u3270, p3_u3269, p3_u3268, p3_u3267, p3_u3266, p3_u3265, p3_u3264, p3_u3376, p3_u3377, p3_u3263, p3_u3262, p3_u3261, p3_u3260, p3_u3259, p3_u3258, p3_u3257, p3_u3256, p3_u3255, p3_u3254, p3_u3253, p3_u3252, p3_u3251, p3_u3250, p3_u3249, p3_u3248, p3_u3247, p3_u3246, p3_u3245, p3_u3244, p3_u3243, p3_u3242, p3_u3241, p3_u3240, p3_u3239, p3_u3238, p3_u3237, p3_u3236, p3_u3235, p3_u3234, p3_u3390, p3_u3393, p3_u3396, p3_u3399, p3_u3402, p3_u3405, p3_u3408, p3_u3411, p3_u3414, p3_u3417, p3_u3420, p3_u3423, p3_u3426, p3_u3429, p3_u3432, p3_u3435, p3_u3438, p3_u3441, p3_u3444, p3_u3446, p3_u3447, p3_u3448, p3_u3449, p3_u3450, p3_u3451, p3_u3452, p3_u3453, p3_u3454, p3_u3455, p3_u3456, p3_u3457, p3_u3458, p3_u3459, p3_u3460, p3_u3461, p3_u3462, p3_u3463, p3_u3464, p3_u3465, p3_u3466, p3_u3467, p3_u3468, p3_u3469, p3_u3470, p3_u3471, p3_u3472, p3_u3473, p3_u3474, p3_u3475, p3_u3476, p3_u3477, p3_u3478, p3_u3479, p3_u3480, p3_u3481, p3_u3482, p3_u3483, p3_u3484, p3_u3485, p3_u3486, p3_u3487, p3_u3488, p3_u3489, p3_u3490, p3_u3233, p3_u3232, p3_u3231, p3_u3230, p3_u3229, p3_u3228, p3_u3227, p3_u3226, p3_u3225, p3_u3224, p3_u3223, p3_u3222, p3_u3221, p3_u3220, p3_u3219, p3_u3218, p3_u3217, p3_u3216, p3_u3215, p3_u3214, p3_u3213, p3_u3212, p3_u3211, p3_u3210, p3_u3209, p3_u3208, p3_u3207, p3_u3206, p3_u3205, p3_u3204, p3_u3203, p3_u3202, p3_u3201, p3_u3200, p3_u3199, p3_u3198, p3_u3197, p3_u3196, p3_u3195, p3_u3194, p3_u3193, p3_u3192, p3_u3191, p3_u3190, p3_u3189, p3_u3188, p3_u3187, p3_u3186, p3_u3185, p3_u3184, p3_u3183, p3_u3182, p3_u3491, p3_u3492, p3_u3493, p3_u3494, p3_u3495, p3_u3496, p3_u3497, p3_u3498, p3_u3499, p3_u3500, p3_u3501, p3_u3502, p3_u3503, p3_u3504, p3_u3505, p3_u3506, p3_u3507, p3_u3508, p3_u3509, p3_u3510, p3_u3511, p3_u3512, p3_u3513, p3_u3514, p3_u3515, p3_u3516, p3_u3517, p3_u3518, p3_u3519, p3_u3520, p3_u3521, p3_u3522, p3_u3296, p3_u3181, p3_u3180, p3_u3179, p3_u3178, p3_u3177, p3_u3176, p3_u3175, p3_u3174, p3_u3173, p3_u3172, p3_u3171, p3_u3170, p3_u3169, p3_u3168, p3_u3167, p3_u3166, p3_u3165, p3_u3164, p3_u3163, p3_u3162, p3_u3161, p3_u3160, p3_u3159, p3_u3158, p3_u3157, p3_u3156, p3_u3155, p3_u3154, p3_u3153, p3_u3151, p3_u3150, p3_u3897;
initial begin
	$readmemb(`in_file, input_vec_mem );
end

always #(`cycle/2) clk = ~clk;

b22_ras cc (.SI_31_(vec[766]), .SI_30_(vec[765]), .SI_29_(vec[764]), .SI_28_(vec[763]), .SI_27_(vec[762]), .SI_26_(vec[761]), .SI_25_(vec[760]), .SI_24_(vec[759]), .SI_23_(vec[758]), .SI_22_(vec[757]), .SI_21_(vec[756]), .SI_20_(vec[755]), .SI_19_(vec[754]), .SI_18_(vec[753]), .SI_17_(vec[752]), .SI_16_(vec[751]), .SI_15_(vec[750]), .SI_14_(vec[749]), .SI_13_(vec[748]), .SI_12_(vec[747]), .SI_11_(vec[746]), .SI_10_(vec[745]), .SI_9_(vec[744]), .SI_8_(vec[743]), .SI_7_(vec[742]), .SI_6_(vec[741]), .SI_5_(vec[740]), .SI_4_(vec[739]), .SI_3_(vec[738]), .SI_2_(vec[737]), .SI_1_(vec[736]), .SI_0_(vec[735]), .P1_IR_REG_0_(vec[734]), .P1_IR_REG_1_(vec[733]), .P1_IR_REG_2_(vec[732]), .P1_IR_REG_3_(vec[731]), .P1_IR_REG_4_(vec[730]), .P1_IR_REG_5_(vec[729]), .P1_IR_REG_6_(vec[728]), .P1_IR_REG_7_(vec[727]), .P1_IR_REG_8_(vec[726]), .P1_IR_REG_9_(vec[725]), .P1_IR_REG_10_(vec[724]), .P1_IR_REG_11_(vec[723]), .P1_IR_REG_12_(vec[722]), .P1_IR_REG_13_(vec[721]), .P1_IR_REG_14_(vec[720]), .P1_IR_REG_15_(vec[719]), .P1_IR_REG_16_(vec[718]), .P1_IR_REG_17_(vec[717]), .P1_IR_REG_18_(vec[716]), .P1_IR_REG_19_(vec[715]), .P1_IR_REG_20_(vec[714]), .P1_IR_REG_21_(vec[713]), .P1_IR_REG_22_(vec[712]), .P1_IR_REG_23_(vec[711]), .P1_IR_REG_24_(vec[710]), .P1_IR_REG_25_(vec[709]), .P1_IR_REG_26_(vec[708]), .P1_IR_REG_27_(vec[707]), .P1_IR_REG_28_(vec[706]), .P1_IR_REG_29_(vec[705]), .P1_IR_REG_30_(vec[704]), .P1_IR_REG_31_(vec[703]), .P1_D_REG_0_(vec[702]), .P1_D_REG_1_(vec[701]), .P1_D_REG_2_(vec[700]), .P1_D_REG_3_(vec[699]), .P1_D_REG_4_(vec[698]), .P1_D_REG_5_(vec[697]), .P1_D_REG_6_(vec[696]), .P1_D_REG_7_(vec[695]), .P1_D_REG_8_(vec[694]), .P1_D_REG_9_(vec[693]), .P1_D_REG_10_(vec[692]), .P1_D_REG_11_(vec[691]), .P1_D_REG_12_(vec[690]), .P1_D_REG_13_(vec[689]), .P1_D_REG_14_(vec[688]), .P1_D_REG_15_(vec[687]), .P1_D_REG_16_(vec[686]), .P1_D_REG_17_(vec[685]), .P1_D_REG_18_(vec[684]), .P1_D_REG_19_(vec[683]), .P1_D_REG_20_(vec[682]), .P1_D_REG_21_(vec[681]), .P1_D_REG_22_(vec[680]), .P1_D_REG_23_(vec[679]), .P1_D_REG_24_(vec[678]), .P1_D_REG_25_(vec[677]), .P1_D_REG_26_(vec[676]), .P1_D_REG_27_(vec[675]), .P1_D_REG_28_(vec[674]), .P1_D_REG_29_(vec[673]), .P1_D_REG_30_(vec[672]), .P1_D_REG_31_(vec[671]), .P1_REG0_REG_0_(vec[670]), .P1_REG0_REG_1_(vec[669]), .P1_REG0_REG_2_(vec[668]), .P1_REG0_REG_3_(vec[667]), .P1_REG0_REG_4_(vec[666]), .P1_REG0_REG_5_(vec[665]), .P1_REG0_REG_6_(vec[664]), .P1_REG0_REG_7_(vec[663]), .P1_REG0_REG_8_(vec[662]), .P1_REG0_REG_9_(vec[661]), .P1_REG0_REG_10_(vec[660]), .P1_REG0_REG_11_(vec[659]), .P1_REG0_REG_12_(vec[658]), .P1_REG0_REG_13_(vec[657]), .P1_REG0_REG_14_(vec[656]), .P1_REG0_REG_15_(vec[655]), .P1_REG0_REG_16_(vec[654]), .P1_REG0_REG_17_(vec[653]), .P1_REG0_REG_18_(vec[652]), .P1_REG0_REG_19_(vec[651]), .P1_REG0_REG_20_(vec[650]), .P1_REG0_REG_21_(vec[649]), .P1_REG0_REG_22_(vec[648]), .P1_REG0_REG_23_(vec[647]), .P1_REG0_REG_24_(vec[646]), .P1_REG0_REG_25_(vec[645]), .P1_REG0_REG_26_(vec[644]), .P1_REG0_REG_27_(vec[643]), .P1_REG0_REG_28_(vec[642]), .P1_REG0_REG_29_(vec[641]), .P1_REG0_REG_30_(vec[640]), .P1_REG0_REG_31_(vec[639]), .P1_REG1_REG_0_(vec[638]), .P1_REG1_REG_1_(vec[637]), .P1_REG1_REG_2_(vec[636]), .P1_REG1_REG_3_(vec[635]), .P1_REG1_REG_4_(vec[634]), .P1_REG1_REG_5_(vec[633]), .P1_REG1_REG_6_(vec[632]), .P1_REG1_REG_7_(vec[631]), .P1_REG1_REG_8_(vec[630]), .P1_REG1_REG_9_(vec[629]), .P1_REG1_REG_10_(vec[628]), .P1_REG1_REG_11_(vec[627]), .P1_REG1_REG_12_(vec[626]), .P1_REG1_REG_13_(vec[625]), .P1_REG1_REG_14_(vec[624]), .P1_REG1_REG_15_(vec[623]), .P1_REG1_REG_16_(vec[622]), .P1_REG1_REG_17_(vec[621]), .P1_REG1_REG_18_(vec[620]), .P1_REG1_REG_19_(vec[619]), .P1_REG1_REG_20_(vec[618]), .P1_REG1_REG_21_(vec[617]), .P1_REG1_REG_22_(vec[616]), .P1_REG1_REG_23_(vec[615]), .P1_REG1_REG_24_(vec[614]), .P1_REG1_REG_25_(vec[613]), .P1_REG1_REG_26_(vec[612]), .P1_REG1_REG_27_(vec[611]), .P1_REG1_REG_28_(vec[610]), .P1_REG1_REG_29_(vec[609]), .P1_REG1_REG_30_(vec[608]), .P1_REG1_REG_31_(vec[607]), .P1_REG2_REG_0_(vec[606]), .P1_REG2_REG_1_(vec[605]), .P1_REG2_REG_2_(vec[604]), .P1_REG2_REG_3_(vec[603]), .P1_REG2_REG_4_(vec[602]), .P1_REG2_REG_5_(vec[601]), .P1_REG2_REG_6_(vec[600]), .P1_REG2_REG_7_(vec[599]), .P1_REG2_REG_8_(vec[598]), .P1_REG2_REG_9_(vec[597]), .P1_REG2_REG_10_(vec[596]), .P1_REG2_REG_11_(vec[595]), .P1_REG2_REG_12_(vec[594]), .P1_REG2_REG_13_(vec[593]), .P1_REG2_REG_14_(vec[592]), .P1_REG2_REG_15_(vec[591]), .P1_REG2_REG_16_(vec[590]), .P1_REG2_REG_17_(vec[589]), .P1_REG2_REG_18_(vec[588]), .P1_REG2_REG_19_(vec[587]), .P1_REG2_REG_20_(vec[586]), .P1_REG2_REG_21_(vec[585]), .P1_REG2_REG_22_(vec[584]), .P1_REG2_REG_23_(vec[583]), .P1_REG2_REG_24_(vec[582]), .P1_REG2_REG_25_(vec[581]), .P1_REG2_REG_26_(vec[580]), .P1_REG2_REG_27_(vec[579]), .P1_REG2_REG_28_(vec[578]), .P1_REG2_REG_29_(vec[577]), .P1_REG2_REG_30_(vec[576]), .P1_REG2_REG_31_(vec[575]), .P1_ADDR_REG_19_(vec[574]), .P1_ADDR_REG_18_(vec[573]), .P1_ADDR_REG_17_(vec[572]), .P1_ADDR_REG_16_(vec[571]), .P1_ADDR_REG_15_(vec[570]), .P1_ADDR_REG_14_(vec[569]), .P1_ADDR_REG_13_(vec[568]), .P1_ADDR_REG_12_(vec[567]), .P1_ADDR_REG_11_(vec[566]), .P1_ADDR_REG_10_(vec[565]), .P1_ADDR_REG_9_(vec[564]), .P1_ADDR_REG_8_(vec[563]), .P1_ADDR_REG_7_(vec[562]), .P1_ADDR_REG_6_(vec[561]), .P1_ADDR_REG_5_(vec[560]), .P1_ADDR_REG_4_(vec[559]), .P1_ADDR_REG_3_(vec[558]), .P1_ADDR_REG_2_(vec[557]), .P1_ADDR_REG_1_(vec[556]), .P1_ADDR_REG_0_(vec[555]), .P1_DATAO_REG_0_(vec[554]), .P1_DATAO_REG_1_(vec[553]), .P1_DATAO_REG_2_(vec[552]), .P1_DATAO_REG_3_(vec[551]), .P1_DATAO_REG_4_(vec[550]), .P1_DATAO_REG_5_(vec[549]), .P1_DATAO_REG_6_(vec[548]), .P1_DATAO_REG_7_(vec[547]), .P1_DATAO_REG_8_(vec[546]), .P1_DATAO_REG_9_(vec[545]), .P1_DATAO_REG_10_(vec[544]), .P1_DATAO_REG_11_(vec[543]), .P1_DATAO_REG_12_(vec[542]), .P1_DATAO_REG_13_(vec[541]), .P1_DATAO_REG_14_(vec[540]), .P1_DATAO_REG_15_(vec[539]), .P1_DATAO_REG_16_(vec[538]), .P1_DATAO_REG_17_(vec[537]), .P1_DATAO_REG_18_(vec[536]), .P1_DATAO_REG_19_(vec[535]), .P1_DATAO_REG_20_(vec[534]), .P1_DATAO_REG_21_(vec[533]), .P1_DATAO_REG_22_(vec[532]), .P1_DATAO_REG_23_(vec[531]), .P1_DATAO_REG_24_(vec[530]), .P1_DATAO_REG_25_(vec[529]), .P1_DATAO_REG_26_(vec[528]), .P1_DATAO_REG_27_(vec[527]), .P1_DATAO_REG_28_(vec[526]), .P1_DATAO_REG_29_(vec[525]), .P1_DATAO_REG_30_(vec[524]), .P1_DATAO_REG_31_(vec[523]), .P1_B_REG(vec[522]), .P1_REG3_REG_15_(vec[521]), .P1_REG3_REG_26_(vec[520]), .P1_REG3_REG_6_(vec[519]), .P1_REG3_REG_18_(vec[518]), .P1_REG3_REG_2_(vec[517]), .P1_REG3_REG_11_(vec[516]), .P1_REG3_REG_22_(vec[515]), .P1_REG3_REG_13_(vec[514]), .P1_REG3_REG_20_(vec[513]), .P1_REG3_REG_0_(vec[512]), .P1_REG3_REG_9_(vec[511]), .P1_REG3_REG_4_(vec[510]), .P1_REG3_REG_24_(vec[509]), .P1_REG3_REG_17_(vec[508]), .P1_REG3_REG_5_(vec[507]), .P1_REG3_REG_16_(vec[506]), .P1_REG3_REG_25_(vec[505]), .P1_REG3_REG_12_(vec[504]), .P1_REG3_REG_21_(vec[503]), .P1_REG3_REG_1_(vec[502]), .P1_REG3_REG_8_(vec[501]), .P1_REG3_REG_28_(vec[500]), .P1_REG3_REG_19_(vec[499]), .P1_REG3_REG_3_(vec[498]), .P1_REG3_REG_10_(vec[497]), .P1_REG3_REG_23_(vec[496]), .P1_REG3_REG_14_(vec[495]), .P1_REG3_REG_27_(vec[494]), .P1_REG3_REG_7_(vec[493]), .P1_STATE_REG(vec[492]), .P1_RD_REG(vec[491]), .P1_WR_REG(vec[490]), .P2_IR_REG_0_(vec[489]), .P2_IR_REG_1_(vec[488]), .P2_IR_REG_2_(vec[487]), .P2_IR_REG_3_(vec[486]), .P2_IR_REG_4_(vec[485]), .P2_IR_REG_5_(vec[484]), .P2_IR_REG_6_(vec[483]), .P2_IR_REG_7_(vec[482]), .P2_IR_REG_8_(vec[481]), .P2_IR_REG_9_(vec[480]), .P2_IR_REG_10_(vec[479]), .P2_IR_REG_11_(vec[478]), .P2_IR_REG_12_(vec[477]), .P2_IR_REG_13_(vec[476]), .P2_IR_REG_14_(vec[475]), .P2_IR_REG_15_(vec[474]), .P2_IR_REG_16_(vec[473]), .P2_IR_REG_17_(vec[472]), .P2_IR_REG_18_(vec[471]), .P2_IR_REG_19_(vec[470]), .P2_IR_REG_20_(vec[469]), .P2_IR_REG_21_(vec[468]), .P2_IR_REG_22_(vec[467]), .P2_IR_REG_23_(vec[466]), .P2_IR_REG_24_(vec[465]), .P2_IR_REG_25_(vec[464]), .P2_IR_REG_26_(vec[463]), .P2_IR_REG_27_(vec[462]), .P2_IR_REG_28_(vec[461]), .P2_IR_REG_29_(vec[460]), .P2_IR_REG_30_(vec[459]), .P2_IR_REG_31_(vec[458]), .P2_D_REG_0_(vec[457]), .P2_D_REG_1_(vec[456]), .P2_D_REG_2_(vec[455]), .P2_D_REG_3_(vec[454]), .P2_D_REG_4_(vec[453]), .P2_D_REG_5_(vec[452]), .P2_D_REG_6_(vec[451]), .P2_D_REG_7_(vec[450]), .P2_D_REG_8_(vec[449]), .P2_D_REG_9_(vec[448]), .P2_D_REG_10_(vec[447]), .P2_D_REG_11_(vec[446]), .P2_D_REG_12_(vec[445]), .P2_D_REG_13_(vec[444]), .P2_D_REG_14_(vec[443]), .P2_D_REG_15_(vec[442]), .P2_D_REG_16_(vec[441]), .P2_D_REG_17_(vec[440]), .P2_D_REG_18_(vec[439]), .P2_D_REG_19_(vec[438]), .P2_D_REG_20_(vec[437]), .P2_D_REG_21_(vec[436]), .P2_D_REG_22_(vec[435]), .P2_D_REG_23_(vec[434]), .P2_D_REG_24_(vec[433]), .P2_D_REG_25_(vec[432]), .P2_D_REG_26_(vec[431]), .P2_D_REG_27_(vec[430]), .P2_D_REG_28_(vec[429]), .P2_D_REG_29_(vec[428]), .P2_D_REG_30_(vec[427]), .P2_D_REG_31_(vec[426]), .P2_REG0_REG_0_(vec[425]), .P2_REG0_REG_1_(vec[424]), .P2_REG0_REG_2_(vec[423]), .P2_REG0_REG_3_(vec[422]), .P2_REG0_REG_4_(vec[421]), .P2_REG0_REG_5_(vec[420]), .P2_REG0_REG_6_(vec[419]), .P2_REG0_REG_7_(vec[418]), .P2_REG0_REG_8_(vec[417]), .P2_REG0_REG_9_(vec[416]), .P2_REG0_REG_10_(vec[415]), .P2_REG0_REG_11_(vec[414]), .P2_REG0_REG_12_(vec[413]), .P2_REG0_REG_13_(vec[412]), .P2_REG0_REG_14_(vec[411]), .P2_REG0_REG_15_(vec[410]), .P2_REG0_REG_16_(vec[409]), .P2_REG0_REG_17_(vec[408]), .P2_REG0_REG_18_(vec[407]), .P2_REG0_REG_19_(vec[406]), .P2_REG0_REG_20_(vec[405]), .P2_REG0_REG_21_(vec[404]), .P2_REG0_REG_22_(vec[403]), .P2_REG0_REG_23_(vec[402]), .P2_REG0_REG_24_(vec[401]), .P2_REG0_REG_25_(vec[400]), .P2_REG0_REG_26_(vec[399]), .P2_REG0_REG_27_(vec[398]), .P2_REG0_REG_28_(vec[397]), .P2_REG0_REG_29_(vec[396]), .P2_REG0_REG_30_(vec[395]), .P2_REG0_REG_31_(vec[394]), .P2_REG1_REG_0_(vec[393]), .P2_REG1_REG_1_(vec[392]), .P2_REG1_REG_2_(vec[391]), .P2_REG1_REG_3_(vec[390]), .P2_REG1_REG_4_(vec[389]), .P2_REG1_REG_5_(vec[388]), .P2_REG1_REG_6_(vec[387]), .P2_REG1_REG_7_(vec[386]), .P2_REG1_REG_8_(vec[385]), .P2_REG1_REG_9_(vec[384]), .P2_REG1_REG_10_(vec[383]), .P2_REG1_REG_11_(vec[382]), .P2_REG1_REG_12_(vec[381]), .P2_REG1_REG_13_(vec[380]), .P2_REG1_REG_14_(vec[379]), .P2_REG1_REG_15_(vec[378]), .P2_REG1_REG_16_(vec[377]), .P2_REG1_REG_17_(vec[376]), .P2_REG1_REG_18_(vec[375]), .P2_REG1_REG_19_(vec[374]), .P2_REG1_REG_20_(vec[373]), .P2_REG1_REG_21_(vec[372]), .P2_REG1_REG_22_(vec[371]), .P2_REG1_REG_23_(vec[370]), .P2_REG1_REG_24_(vec[369]), .P2_REG1_REG_25_(vec[368]), .P2_REG1_REG_26_(vec[367]), .P2_REG1_REG_27_(vec[366]), .P2_REG1_REG_28_(vec[365]), .P2_REG1_REG_29_(vec[364]), .P2_REG1_REG_30_(vec[363]), .P2_REG1_REG_31_(vec[362]), .P2_REG2_REG_0_(vec[361]), .P2_REG2_REG_1_(vec[360]), .P2_REG2_REG_2_(vec[359]), .P2_REG2_REG_3_(vec[358]), .P2_REG2_REG_4_(vec[357]), .P2_REG2_REG_5_(vec[356]), .P2_REG2_REG_6_(vec[355]), .P2_REG2_REG_7_(vec[354]), .P2_REG2_REG_8_(vec[353]), .P2_REG2_REG_9_(vec[352]), .P2_REG2_REG_10_(vec[351]), .P2_REG2_REG_11_(vec[350]), .P2_REG2_REG_12_(vec[349]), .P2_REG2_REG_13_(vec[348]), .P2_REG2_REG_14_(vec[347]), .P2_REG2_REG_15_(vec[346]), .P2_REG2_REG_16_(vec[345]), .P2_REG2_REG_17_(vec[344]), .P2_REG2_REG_18_(vec[343]), .P2_REG2_REG_19_(vec[342]), .P2_REG2_REG_20_(vec[341]), .P2_REG2_REG_21_(vec[340]), .P2_REG2_REG_22_(vec[339]), .P2_REG2_REG_23_(vec[338]), .P2_REG2_REG_24_(vec[337]), .P2_REG2_REG_25_(vec[336]), .P2_REG2_REG_26_(vec[335]), .P2_REG2_REG_27_(vec[334]), .P2_REG2_REG_28_(vec[333]), .P2_REG2_REG_29_(vec[332]), .P2_REG2_REG_30_(vec[331]), .P2_REG2_REG_31_(vec[330]), .P2_ADDR_REG_19_(vec[329]), .P2_ADDR_REG_18_(vec[328]), .P2_ADDR_REG_17_(vec[327]), .P2_ADDR_REG_16_(vec[326]), .P2_ADDR_REG_15_(vec[325]), .P2_ADDR_REG_14_(vec[324]), .P2_ADDR_REG_13_(vec[323]), .P2_ADDR_REG_12_(vec[322]), .P2_ADDR_REG_11_(vec[321]), .P2_ADDR_REG_10_(vec[320]), .P2_ADDR_REG_9_(vec[319]), .P2_ADDR_REG_8_(vec[318]), .P2_ADDR_REG_7_(vec[317]), .P2_ADDR_REG_6_(vec[316]), .P2_ADDR_REG_5_(vec[315]), .P2_ADDR_REG_4_(vec[314]), .P2_ADDR_REG_3_(vec[313]), .P2_ADDR_REG_2_(vec[312]), .P2_ADDR_REG_1_(vec[311]), .P2_ADDR_REG_0_(vec[310]), .P2_DATAO_REG_0_(vec[309]), .P2_DATAO_REG_1_(vec[308]), .P2_DATAO_REG_2_(vec[307]), .P2_DATAO_REG_3_(vec[306]), .P2_DATAO_REG_4_(vec[305]), .P2_DATAO_REG_5_(vec[304]), .P2_DATAO_REG_6_(vec[303]), .P2_DATAO_REG_7_(vec[302]), .P2_DATAO_REG_8_(vec[301]), .P2_DATAO_REG_9_(vec[300]), .P2_DATAO_REG_10_(vec[299]), .P2_DATAO_REG_11_(vec[298]), .P2_DATAO_REG_12_(vec[297]), .P2_DATAO_REG_13_(vec[296]), .P2_DATAO_REG_14_(vec[295]), .P2_DATAO_REG_15_(vec[294]), .P2_DATAO_REG_16_(vec[293]), .P2_DATAO_REG_17_(vec[292]), .P2_DATAO_REG_18_(vec[291]), .P2_DATAO_REG_19_(vec[290]), .P2_DATAO_REG_20_(vec[289]), .P2_DATAO_REG_21_(vec[288]), .P2_DATAO_REG_22_(vec[287]), .P2_DATAO_REG_23_(vec[286]), .P2_DATAO_REG_24_(vec[285]), .P2_DATAO_REG_25_(vec[284]), .P2_DATAO_REG_26_(vec[283]), .P2_DATAO_REG_27_(vec[282]), .P2_DATAO_REG_28_(vec[281]), .P2_DATAO_REG_29_(vec[280]), .P2_DATAO_REG_30_(vec[279]), .P2_DATAO_REG_31_(vec[278]), .P2_B_REG(vec[277]), .P2_REG3_REG_15_(vec[276]), .P2_REG3_REG_26_(vec[275]), .P2_REG3_REG_6_(vec[274]), .P2_REG3_REG_18_(vec[273]), .P2_REG3_REG_2_(vec[272]), .P2_REG3_REG_11_(vec[271]), .P2_REG3_REG_22_(vec[270]), .P2_REG3_REG_13_(vec[269]), .P2_REG3_REG_20_(vec[268]), .P2_REG3_REG_0_(vec[267]), .P2_REG3_REG_9_(vec[266]), .P2_REG3_REG_4_(vec[265]), .P2_REG3_REG_24_(vec[264]), .P2_REG3_REG_17_(vec[263]), .P2_REG3_REG_5_(vec[262]), .P2_REG3_REG_16_(vec[261]), .P2_REG3_REG_25_(vec[260]), .P2_REG3_REG_12_(vec[259]), .P2_REG3_REG_21_(vec[258]), .P2_REG3_REG_1_(vec[257]), .P2_REG3_REG_8_(vec[256]), .P2_REG3_REG_28_(vec[255]), .P2_REG3_REG_19_(vec[254]), .P2_REG3_REG_3_(vec[253]), .P2_REG3_REG_10_(vec[252]), .P2_REG3_REG_23_(vec[251]), .P2_REG3_REG_14_(vec[250]), .P2_REG3_REG_27_(vec[249]), .P2_REG3_REG_7_(vec[248]), .P2_STATE_REG(vec[247]), .P2_RD_REG(vec[246]), .P2_WR_REG(vec[245]), .P3_IR_REG_0_(vec[244]), .P3_IR_REG_1_(vec[243]), .P3_IR_REG_2_(vec[242]), .P3_IR_REG_3_(vec[241]), .P3_IR_REG_4_(vec[240]), .P3_IR_REG_5_(vec[239]), .P3_IR_REG_6_(vec[238]), .P3_IR_REG_7_(vec[237]), .P3_IR_REG_8_(vec[236]), .P3_IR_REG_9_(vec[235]), .P3_IR_REG_10_(vec[234]), .P3_IR_REG_11_(vec[233]), .P3_IR_REG_12_(vec[232]), .P3_IR_REG_13_(vec[231]), .P3_IR_REG_14_(vec[230]), .P3_IR_REG_15_(vec[229]), .P3_IR_REG_16_(vec[228]), .P3_IR_REG_17_(vec[227]), .P3_IR_REG_18_(vec[226]), .P3_IR_REG_19_(vec[225]), .P3_IR_REG_20_(vec[224]), .P3_IR_REG_21_(vec[223]), .P3_IR_REG_22_(vec[222]), .P3_IR_REG_23_(vec[221]), .P3_IR_REG_24_(vec[220]), .P3_IR_REG_25_(vec[219]), .P3_IR_REG_26_(vec[218]), .P3_IR_REG_27_(vec[217]), .P3_IR_REG_28_(vec[216]), .P3_IR_REG_29_(vec[215]), .P3_IR_REG_30_(vec[214]), .P3_IR_REG_31_(vec[213]), .P3_D_REG_0_(vec[212]), .P3_D_REG_1_(vec[211]), .P3_D_REG_2_(vec[210]), .P3_D_REG_3_(vec[209]), .P3_D_REG_4_(vec[208]), .P3_D_REG_5_(vec[207]), .P3_D_REG_6_(vec[206]), .P3_D_REG_7_(vec[205]), .P3_D_REG_8_(vec[204]), .P3_D_REG_9_(vec[203]), .P3_D_REG_10_(vec[202]), .P3_D_REG_11_(vec[201]), .P3_D_REG_12_(vec[200]), .P3_D_REG_13_(vec[199]), .P3_D_REG_14_(vec[198]), .P3_D_REG_15_(vec[197]), .P3_D_REG_16_(vec[196]), .P3_D_REG_17_(vec[195]), .P3_D_REG_18_(vec[194]), .P3_D_REG_19_(vec[193]), .P3_D_REG_20_(vec[192]), .P3_D_REG_21_(vec[191]), .P3_D_REG_22_(vec[190]), .P3_D_REG_23_(vec[189]), .P3_D_REG_24_(vec[188]), .P3_D_REG_25_(vec[187]), .P3_D_REG_26_(vec[186]), .P3_D_REG_27_(vec[185]), .P3_D_REG_28_(vec[184]), .P3_D_REG_29_(vec[183]), .P3_D_REG_30_(vec[182]), .P3_D_REG_31_(vec[181]), .P3_REG0_REG_0_(vec[180]), .P3_REG0_REG_1_(vec[179]), .P3_REG0_REG_2_(vec[178]), .P3_REG0_REG_3_(vec[177]), .P3_REG0_REG_4_(vec[176]), .P3_REG0_REG_5_(vec[175]), .P3_REG0_REG_6_(vec[174]), .P3_REG0_REG_7_(vec[173]), .P3_REG0_REG_8_(vec[172]), .P3_REG0_REG_9_(vec[171]), .P3_REG0_REG_10_(vec[170]), .P3_REG0_REG_11_(vec[169]), .P3_REG0_REG_12_(vec[168]), .P3_REG0_REG_13_(vec[167]), .P3_REG0_REG_14_(vec[166]), .P3_REG0_REG_15_(vec[165]), .P3_REG0_REG_16_(vec[164]), .P3_REG0_REG_17_(vec[163]), .P3_REG0_REG_18_(vec[162]), .P3_REG0_REG_19_(vec[161]), .P3_REG0_REG_20_(vec[160]), .P3_REG0_REG_21_(vec[159]), .P3_REG0_REG_22_(vec[158]), .P3_REG0_REG_23_(vec[157]), .P3_REG0_REG_24_(vec[156]), .P3_REG0_REG_25_(vec[155]), .P3_REG0_REG_26_(vec[154]), .P3_REG0_REG_27_(vec[153]), .P3_REG0_REG_28_(vec[152]), .P3_REG0_REG_29_(vec[151]), .P3_REG0_REG_30_(vec[150]), .P3_REG0_REG_31_(vec[149]), .P3_REG1_REG_0_(vec[148]), .P3_REG1_REG_1_(vec[147]), .P3_REG1_REG_2_(vec[146]), .P3_REG1_REG_3_(vec[145]), .P3_REG1_REG_4_(vec[144]), .P3_REG1_REG_5_(vec[143]), .P3_REG1_REG_6_(vec[142]), .P3_REG1_REG_7_(vec[141]), .P3_REG1_REG_8_(vec[140]), .P3_REG1_REG_9_(vec[139]), .P3_REG1_REG_10_(vec[138]), .P3_REG1_REG_11_(vec[137]), .P3_REG1_REG_12_(vec[136]), .P3_REG1_REG_13_(vec[135]), .P3_REG1_REG_14_(vec[134]), .P3_REG1_REG_15_(vec[133]), .P3_REG1_REG_16_(vec[132]), .P3_REG1_REG_17_(vec[131]), .P3_REG1_REG_18_(vec[130]), .P3_REG1_REG_19_(vec[129]), .P3_REG1_REG_20_(vec[128]), .P3_REG1_REG_21_(vec[127]), .P3_REG1_REG_22_(vec[126]), .P3_REG1_REG_23_(vec[125]), .P3_REG1_REG_24_(vec[124]), .P3_REG1_REG_25_(vec[123]), .P3_REG1_REG_26_(vec[122]), .P3_REG1_REG_27_(vec[121]), .P3_REG1_REG_28_(vec[120]), .P3_REG1_REG_29_(vec[119]), .P3_REG1_REG_30_(vec[118]), .P3_REG1_REG_31_(vec[117]), .P3_REG2_REG_0_(vec[116]), .P3_REG2_REG_1_(vec[115]), .P3_REG2_REG_2_(vec[114]), .P3_REG2_REG_3_(vec[113]), .P3_REG2_REG_4_(vec[112]), .P3_REG2_REG_5_(vec[111]), .P3_REG2_REG_6_(vec[110]), .P3_REG2_REG_7_(vec[109]), .P3_REG2_REG_8_(vec[108]), .P3_REG2_REG_9_(vec[107]), .P3_REG2_REG_10_(vec[106]), .P3_REG2_REG_11_(vec[105]), .P3_REG2_REG_12_(vec[104]), .P3_REG2_REG_13_(vec[103]), .P3_REG2_REG_14_(vec[102]), .P3_REG2_REG_15_(vec[101]), .P3_REG2_REG_16_(vec[100]), .P3_REG2_REG_17_(vec[99]), .P3_REG2_REG_18_(vec[98]), .P3_REG2_REG_19_(vec[97]), .P3_REG2_REG_20_(vec[96]), .P3_REG2_REG_21_(vec[95]), .P3_REG2_REG_22_(vec[94]), .P3_REG2_REG_23_(vec[93]), .P3_REG2_REG_24_(vec[92]), .P3_REG2_REG_25_(vec[91]), .P3_REG2_REG_26_(vec[90]), .P3_REG2_REG_27_(vec[89]), .P3_REG2_REG_28_(vec[88]), .P3_REG2_REG_29_(vec[87]), .P3_REG2_REG_30_(vec[86]), .P3_REG2_REG_31_(vec[85]), .P3_ADDR_REG_19_(vec[84]), .P3_ADDR_REG_18_(vec[83]), .P3_ADDR_REG_17_(vec[82]), .P3_ADDR_REG_16_(vec[81]), .P3_ADDR_REG_15_(vec[80]), .P3_ADDR_REG_14_(vec[79]), .P3_ADDR_REG_13_(vec[78]), .P3_ADDR_REG_12_(vec[77]), .P3_ADDR_REG_11_(vec[76]), .P3_ADDR_REG_10_(vec[75]), .P3_ADDR_REG_9_(vec[74]), .P3_ADDR_REG_8_(vec[73]), .P3_ADDR_REG_7_(vec[72]), .P3_ADDR_REG_6_(vec[71]), .P3_ADDR_REG_5_(vec[70]), .P3_ADDR_REG_4_(vec[69]), .P3_ADDR_REG_3_(vec[68]), .P3_ADDR_REG_2_(vec[67]), .P3_ADDR_REG_1_(vec[66]), .P3_ADDR_REG_0_(vec[65]), .P3_DATAO_REG_0_(vec[64]), .P3_DATAO_REG_1_(vec[63]), .P3_DATAO_REG_2_(vec[62]), .P3_DATAO_REG_3_(vec[61]), .P3_DATAO_REG_4_(vec[60]), .P3_DATAO_REG_5_(vec[59]), .P3_DATAO_REG_6_(vec[58]), .P3_DATAO_REG_7_(vec[57]), .P3_DATAO_REG_8_(vec[56]), .P3_DATAO_REG_9_(vec[55]), .P3_DATAO_REG_10_(vec[54]), .P3_DATAO_REG_11_(vec[53]), .P3_DATAO_REG_12_(vec[52]), .P3_DATAO_REG_13_(vec[51]), .P3_DATAO_REG_14_(vec[50]), .P3_DATAO_REG_15_(vec[49]), .P3_DATAO_REG_16_(vec[48]), .P3_DATAO_REG_17_(vec[47]), .P3_DATAO_REG_18_(vec[46]), .P3_DATAO_REG_19_(vec[45]), .P3_DATAO_REG_20_(vec[44]), .P3_DATAO_REG_21_(vec[43]), .P3_DATAO_REG_22_(vec[42]), .P3_DATAO_REG_23_(vec[41]), .P3_DATAO_REG_24_(vec[40]), .P3_DATAO_REG_25_(vec[39]), .P3_DATAO_REG_26_(vec[38]), .P3_DATAO_REG_27_(vec[37]), .P3_DATAO_REG_28_(vec[36]), .P3_DATAO_REG_29_(vec[35]), .P3_DATAO_REG_30_(vec[34]), .P3_DATAO_REG_31_(vec[33]), .P3_B_REG(vec[32]), .P3_REG3_REG_15_(vec[31]), .P3_REG3_REG_26_(vec[30]), .P3_REG3_REG_6_(vec[29]), .P3_REG3_REG_18_(vec[28]), .P3_REG3_REG_2_(vec[27]), .P3_REG3_REG_11_(vec[26]), .P3_REG3_REG_22_(vec[25]), .P3_REG3_REG_13_(vec[24]), .P3_REG3_REG_20_(vec[23]), .P3_REG3_REG_0_(vec[22]), .P3_REG3_REG_9_(vec[21]), .P3_REG3_REG_4_(vec[20]), .P3_REG3_REG_24_(vec[19]), .P3_REG3_REG_17_(vec[18]), .P3_REG3_REG_5_(vec[17]), .P3_REG3_REG_16_(vec[16]), .P3_REG3_REG_25_(vec[15]), .P3_REG3_REG_12_(vec[14]), .P3_REG3_REG_21_(vec[13]), .P3_REG3_REG_1_(vec[12]), .P3_REG3_REG_8_(vec[11]), .P3_REG3_REG_28_(vec[10]), .P3_REG3_REG_19_(vec[9]), .P3_REG3_REG_3_(vec[8]), .P3_REG3_REG_10_(vec[7]), .P3_REG3_REG_23_(vec[6]), .P3_REG3_REG_14_(vec[5]), .P3_REG3_REG_27_(vec[4]), .P3_REG3_REG_7_(vec[3]), .P3_STATE_REG(vec[2]), .P3_RD_REG(vec[1]), .P3_WR_REG(vec[0]), .SUB_1596_U4(sub_1596_u4), .SUB_1596_U62(sub_1596_u62), .SUB_1596_U63(sub_1596_u63), .SUB_1596_U64(sub_1596_u64), .SUB_1596_U65(sub_1596_u65), .SUB_1596_U66(sub_1596_u66), .SUB_1596_U67(sub_1596_u67), .SUB_1596_U68(sub_1596_u68), .SUB_1596_U69(sub_1596_u69), .SUB_1596_U70(sub_1596_u70), .SUB_1596_U54(sub_1596_u54), .SUB_1596_U55(sub_1596_u55), .SUB_1596_U56(sub_1596_u56), .SUB_1596_U57(sub_1596_u57), .SUB_1596_U58(sub_1596_u58), .SUB_1596_U59(sub_1596_u59), .SUB_1596_U60(sub_1596_u60), .SUB_1596_U61(sub_1596_u61), .SUB_1596_U5(sub_1596_u5), .SUB_1596_U53(sub_1596_u53), .U29(u29), .U28(u28), .P1_U3355(p1_u3355), .P1_U3354(p1_u3354), .P1_U3353(p1_u3353), .P1_U3352(p1_u3352), .P1_U3351(p1_u3351), .P1_U3350(p1_u3350), .P1_U3349(p1_u3349), .P1_U3348(p1_u3348), .P1_U3347(p1_u3347), .P1_U3346(p1_u3346), .P1_U3345(p1_u3345), .P1_U3344(p1_u3344), .P1_U3343(p1_u3343), .P1_U3342(p1_u3342), .P1_U3341(p1_u3341), .P1_U3340(p1_u3340), .P1_U3339(p1_u3339), .P1_U3338(p1_u3338), .P1_U3337(p1_u3337), .P1_U3336(p1_u3336), .P1_U3335(p1_u3335), .P1_U3334(p1_u3334), .P1_U3333(p1_u3333), .P1_U3332(p1_u3332), .P1_U3331(p1_u3331), .P1_U3330(p1_u3330), .P1_U3329(p1_u3329), .P1_U3328(p1_u3328), .P1_U3327(p1_u3327), .P1_U3326(p1_u3326), .P1_U3325(p1_u3325), .P1_U3324(p1_u3324), .P1_U3445(p1_u3445), .P1_U3446(p1_u3446), .P1_U3323(p1_u3323), .P1_U3322(p1_u3322), .P1_U3321(p1_u3321), .P1_U3320(p1_u3320), .P1_U3319(p1_u3319), .P1_U3318(p1_u3318), .P1_U3317(p1_u3317), .P1_U3316(p1_u3316), .P1_U3315(p1_u3315), .P1_U3314(p1_u3314), .P1_U3313(p1_u3313), .P1_U3312(p1_u3312), .P1_U3311(p1_u3311), .P1_U3310(p1_u3310), .P1_U3309(p1_u3309), .P1_U3308(p1_u3308), .P1_U3307(p1_u3307), .P1_U3306(p1_u3306), .P1_U3305(p1_u3305), .P1_U3304(p1_u3304), .P1_U3303(p1_u3303), .P1_U3302(p1_u3302), .P1_U3301(p1_u3301), .P1_U3300(p1_u3300), .P1_U3299(p1_u3299), .P1_U3298(p1_u3298), .P1_U3297(p1_u3297), .P1_U3296(p1_u3296), .P1_U3295(p1_u3295), .P1_U3294(p1_u3294), .P1_U3459(p1_u3459), .P1_U3462(p1_u3462), .P1_U3465(p1_u3465), .P1_U3468(p1_u3468), .P1_U3471(p1_u3471), .P1_U3474(p1_u3474), .P1_U3477(p1_u3477), .P1_U3480(p1_u3480), .P1_U3483(p1_u3483), .P1_U3486(p1_u3486), .P1_U3489(p1_u3489), .P1_U3492(p1_u3492), .P1_U3495(p1_u3495), .P1_U3498(p1_u3498), .P1_U3501(p1_u3501), .P1_U3504(p1_u3504), .P1_U3507(p1_u3507), .P1_U3510(p1_u3510), .P1_U3513(p1_u3513), .P1_U3515(p1_u3515), .P1_U3516(p1_u3516), .P1_U3517(p1_u3517), .P1_U3518(p1_u3518), .P1_U3519(p1_u3519), .P1_U3520(p1_u3520), .P1_U3521(p1_u3521), .P1_U3522(p1_u3522), .P1_U3523(p1_u3523), .P1_U3524(p1_u3524), .P1_U3525(p1_u3525), .P1_U3526(p1_u3526), .P1_U3527(p1_u3527), .P1_U3528(p1_u3528), .P1_U3529(p1_u3529), .P1_U3530(p1_u3530), .P1_U3531(p1_u3531), .P1_U3532(p1_u3532), .P1_U3533(p1_u3533), .P1_U3534(p1_u3534), .P1_U3535(p1_u3535), .P1_U3536(p1_u3536), .P1_U3537(p1_u3537), .P1_U3538(p1_u3538), .P1_U3539(p1_u3539), .P1_U3540(p1_u3540), .P1_U3541(p1_u3541), .P1_U3542(p1_u3542), .P1_U3543(p1_u3543), .P1_U3544(p1_u3544), .P1_U3545(p1_u3545), .P1_U3546(p1_u3546), .P1_U3547(p1_u3547), .P1_U3548(p1_u3548), .P1_U3549(p1_u3549), .P1_U3550(p1_u3550), .P1_U3551(p1_u3551), .P1_U3552(p1_u3552), .P1_U3553(p1_u3553), .P1_U3554(p1_u3554), .P1_U3555(p1_u3555), .P1_U3556(p1_u3556), .P1_U3557(p1_u3557), .P1_U3558(p1_u3558), .P1_U3559(p1_u3559), .P1_U3293(p1_u3293), .P1_U3292(p1_u3292), .P1_U3291(p1_u3291), .P1_U3290(p1_u3290), .P1_U3289(p1_u3289), .P1_U3288(p1_u3288), .P1_U3287(p1_u3287), .P1_U3286(p1_u3286), .P1_U3285(p1_u3285), .P1_U3284(p1_u3284), .P1_U3283(p1_u3283), .P1_U3282(p1_u3282), .P1_U3281(p1_u3281), .P1_U3280(p1_u3280), .P1_U3279(p1_u3279), .P1_U3278(p1_u3278), .P1_U3277(p1_u3277), .P1_U3276(p1_u3276), .P1_U3275(p1_u3275), .P1_U3274(p1_u3274), .P1_U3273(p1_u3273), .P1_U3272(p1_u3272), .P1_U3271(p1_u3271), .P1_U3270(p1_u3270), .P1_U3269(p1_u3269), .P1_U3268(p1_u3268), .P1_U3267(p1_u3267), .P1_U3266(p1_u3266), .P1_U3265(p1_u3265), .P1_U3356(p1_u3356), .P1_U3264(p1_u3264), .P1_U3263(p1_u3263), .P1_U3262(p1_u3262), .P1_U3261(p1_u3261), .P1_U3260(p1_u3260), .P1_U3259(p1_u3259), .P1_U3258(p1_u3258), .P1_U3257(p1_u3257), .P1_U3256(p1_u3256), .P1_U3255(p1_u3255), .P1_U3254(p1_u3254), .P1_U3253(p1_u3253), .P1_U3252(p1_u3252), .P1_U3251(p1_u3251), .P1_U3250(p1_u3250), .P1_U3249(p1_u3249), .P1_U3248(p1_u3248), .P1_U3247(p1_u3247), .P1_U3246(p1_u3246), .P1_U3245(p1_u3245), .P1_U3244(p1_u3244), .P1_U3243(p1_u3243), .P1_U3560(p1_u3560), .P1_U3561(p1_u3561), .P1_U3562(p1_u3562), .P1_U3563(p1_u3563), .P1_U3564(p1_u3564), .P1_U3565(p1_u3565), .P1_U3566(p1_u3566), .P1_U3567(p1_u3567), .P1_U3568(p1_u3568), .P1_U3569(p1_u3569), .P1_U3570(p1_u3570), .P1_U3571(p1_u3571), .P1_U3572(p1_u3572), .P1_U3573(p1_u3573), .P1_U3574(p1_u3574), .P1_U3575(p1_u3575), .P1_U3576(p1_u3576), .P1_U3577(p1_u3577), .P1_U3578(p1_u3578), .P1_U3579(p1_u3579), .P1_U3580(p1_u3580), .P1_U3581(p1_u3581), .P1_U3582(p1_u3582), .P1_U3583(p1_u3583), .P1_U3584(p1_u3584), .P1_U3585(p1_u3585), .P1_U3586(p1_u3586), .P1_U3587(p1_u3587), .P1_U3588(p1_u3588), .P1_U3589(p1_u3589), .P1_U3590(p1_u3590), .P1_U3591(p1_u3591), .P1_U3242(p1_u3242), .P1_U3241(p1_u3241), .P1_U3240(p1_u3240), .P1_U3239(p1_u3239), .P1_U3238(p1_u3238), .P1_U3237(p1_u3237), .P1_U3236(p1_u3236), .P1_U3235(p1_u3235), .P1_U3234(p1_u3234), .P1_U3233(p1_u3233), .P1_U3232(p1_u3232), .P1_U3231(p1_u3231), .P1_U3230(p1_u3230), .P1_U3229(p1_u3229), .P1_U3228(p1_u3228), .P1_U3227(p1_u3227), .P1_U3226(p1_u3226), .P1_U3225(p1_u3225), .P1_U3224(p1_u3224), .P1_U3223(p1_u3223), .P1_U3222(p1_u3222), .P1_U3221(p1_u3221), .P1_U3220(p1_u3220), .P1_U3219(p1_u3219), .P1_U3218(p1_u3218), .P1_U3217(p1_u3217), .P1_U3216(p1_u3216), .P1_U3215(p1_u3215), .P1_U3214(p1_u3214), .P1_U3213(p1_u3213), .P1_U3086(p1_u3086), .P1_U3085(p1_u3085), .P1_U4016(p1_u4016), .P2_U3327(p2_u3327), .P2_U3326(p2_u3326), .P2_U3325(p2_u3325), .P2_U3324(p2_u3324), .P2_U3323(p2_u3323), .P2_U3322(p2_u3322), .P2_U3321(p2_u3321), .P2_U3320(p2_u3320), .P2_U3319(p2_u3319), .P2_U3318(p2_u3318), .P2_U3317(p2_u3317), .P2_U3316(p2_u3316), .P2_U3315(p2_u3315), .P2_U3314(p2_u3314), .P2_U3313(p2_u3313), .P2_U3312(p2_u3312), .P2_U3311(p2_u3311), .P2_U3310(p2_u3310), .P2_U3309(p2_u3309), .P2_U3308(p2_u3308), .P2_U3307(p2_u3307), .P2_U3306(p2_u3306), .P2_U3305(p2_u3305), .P2_U3304(p2_u3304), .P2_U3303(p2_u3303), .P2_U3302(p2_u3302), .P2_U3301(p2_u3301), .P2_U3300(p2_u3300), .P2_U3299(p2_u3299), .P2_U3298(p2_u3298), .P2_U3297(p2_u3297), .P2_U3296(p2_u3296), .P2_U3416(p2_u3416), .P2_U3417(p2_u3417), .P2_U3295(p2_u3295), .P2_U3294(p2_u3294), .P2_U3293(p2_u3293), .P2_U3292(p2_u3292), .P2_U3291(p2_u3291), .P2_U3290(p2_u3290), .P2_U3289(p2_u3289), .P2_U3288(p2_u3288), .P2_U3287(p2_u3287), .P2_U3286(p2_u3286), .P2_U3285(p2_u3285), .P2_U3284(p2_u3284), .P2_U3283(p2_u3283), .P2_U3282(p2_u3282), .P2_U3281(p2_u3281), .P2_U3280(p2_u3280), .P2_U3279(p2_u3279), .P2_U3278(p2_u3278), .P2_U3277(p2_u3277), .P2_U3276(p2_u3276), .P2_U3275(p2_u3275), .P2_U3274(p2_u3274), .P2_U3273(p2_u3273), .P2_U3272(p2_u3272), .P2_U3271(p2_u3271), .P2_U3270(p2_u3270), .P2_U3269(p2_u3269), .P2_U3268(p2_u3268), .P2_U3267(p2_u3267), .P2_U3266(p2_u3266), .P2_U3430(p2_u3430), .P2_U3433(p2_u3433), .P2_U3436(p2_u3436), .P2_U3439(p2_u3439), .P2_U3442(p2_u3442), .P2_U3445(p2_u3445), .P2_U3448(p2_u3448), .P2_U3451(p2_u3451), .P2_U3454(p2_u3454), .P2_U3457(p2_u3457), .P2_U3460(p2_u3460), .P2_U3463(p2_u3463), .P2_U3466(p2_u3466), .P2_U3469(p2_u3469), .P2_U3472(p2_u3472), .P2_U3475(p2_u3475), .P2_U3478(p2_u3478), .P2_U3481(p2_u3481), .P2_U3484(p2_u3484), .P2_U3486(p2_u3486), .P2_U3487(p2_u3487), .P2_U3488(p2_u3488), .P2_U3489(p2_u3489), .P2_U3490(p2_u3490), .P2_U3491(p2_u3491), .P2_U3492(p2_u3492), .P2_U3493(p2_u3493), .P2_U3494(p2_u3494), .P2_U3495(p2_u3495), .P2_U3496(p2_u3496), .P2_U3497(p2_u3497), .P2_U3498(p2_u3498), .P2_U3499(p2_u3499), .P2_U3500(p2_u3500), .P2_U3501(p2_u3501), .P2_U3502(p2_u3502), .P2_U3503(p2_u3503), .P2_U3504(p2_u3504), .P2_U3505(p2_u3505), .P2_U3506(p2_u3506), .P2_U3507(p2_u3507), .P2_U3508(p2_u3508), .P2_U3509(p2_u3509), .P2_U3510(p2_u3510), .P2_U3511(p2_u3511), .P2_U3512(p2_u3512), .P2_U3513(p2_u3513), .P2_U3514(p2_u3514), .P2_U3515(p2_u3515), .P2_U3516(p2_u3516), .P2_U3517(p2_u3517), .P2_U3518(p2_u3518), .P2_U3519(p2_u3519), .P2_U3520(p2_u3520), .P2_U3521(p2_u3521), .P2_U3522(p2_u3522), .P2_U3523(p2_u3523), .P2_U3524(p2_u3524), .P2_U3525(p2_u3525), .P2_U3526(p2_u3526), .P2_U3527(p2_u3527), .P2_U3528(p2_u3528), .P2_U3529(p2_u3529), .P2_U3530(p2_u3530), .P2_U3265(p2_u3265), .P2_U3264(p2_u3264), .P2_U3263(p2_u3263), .P2_U3262(p2_u3262), .P2_U3261(p2_u3261), .P2_U3260(p2_u3260), .P2_U3259(p2_u3259), .P2_U3258(p2_u3258), .P2_U3257(p2_u3257), .P2_U3256(p2_u3256), .P2_U3255(p2_u3255), .P2_U3254(p2_u3254), .P2_U3253(p2_u3253), .P2_U3252(p2_u3252), .P2_U3251(p2_u3251), .P2_U3250(p2_u3250), .P2_U3249(p2_u3249), .P2_U3248(p2_u3248), .P2_U3247(p2_u3247), .P2_U3246(p2_u3246), .P2_U3245(p2_u3245), .P2_U3244(p2_u3244), .P2_U3243(p2_u3243), .P2_U3242(p2_u3242), .P2_U3241(p2_u3241), .P2_U3240(p2_u3240), .P2_U3239(p2_u3239), .P2_U3238(p2_u3238), .P2_U3237(p2_u3237), .P2_U3236(p2_u3236), .P2_U3235(p2_u3235), .P2_U3234(p2_u3234), .P2_U3233(p2_u3233), .P2_U3232(p2_u3232), .P2_U3231(p2_u3231), .P2_U3230(p2_u3230), .P2_U3229(p2_u3229), .P2_U3228(p2_u3228), .P2_U3227(p2_u3227), .P2_U3226(p2_u3226), .P2_U3225(p2_u3225), .P2_U3224(p2_u3224), .P2_U3223(p2_u3223), .P2_U3222(p2_u3222), .P2_U3221(p2_u3221), .P2_U3220(p2_u3220), .P2_U3219(p2_u3219), .P2_U3218(p2_u3218), .P2_U3217(p2_u3217), .P2_U3216(p2_u3216), .P2_U3215(p2_u3215), .P2_U3214(p2_u3214), .P2_U3531(p2_u3531), .P2_U3532(p2_u3532), .P2_U3533(p2_u3533), .P2_U3534(p2_u3534), .P2_U3535(p2_u3535), .P2_U3536(p2_u3536), .P2_U3537(p2_u3537), .P2_U3538(p2_u3538), .P2_U3539(p2_u3539), .P2_U3540(p2_u3540), .P2_U3541(p2_u3541), .P2_U3542(p2_u3542), .P2_U3543(p2_u3543), .P2_U3544(p2_u3544), .P2_U3545(p2_u3545), .P2_U3546(p2_u3546), .P2_U3547(p2_u3547), .P2_U3548(p2_u3548), .P2_U3549(p2_u3549), .P2_U3550(p2_u3550), .P2_U3551(p2_u3551), .P2_U3552(p2_u3552), .P2_U3553(p2_u3553), .P2_U3554(p2_u3554), .P2_U3555(p2_u3555), .P2_U3556(p2_u3556), .P2_U3557(p2_u3557), .P2_U3558(p2_u3558), .P2_U3559(p2_u3559), .P2_U3560(p2_u3560), .P2_U3561(p2_u3561), .P2_U3562(p2_u3562), .P2_U3328(p2_u3328), .P2_U3213(p2_u3213), .P2_U3212(p2_u3212), .P2_U3211(p2_u3211), .P2_U3210(p2_u3210), .P2_U3209(p2_u3209), .P2_U3208(p2_u3208), .P2_U3207(p2_u3207), .P2_U3206(p2_u3206), .P2_U3205(p2_u3205), .P2_U3204(p2_u3204), .P2_U3203(p2_u3203), .P2_U3202(p2_u3202), .P2_U3201(p2_u3201), .P2_U3200(p2_u3200), .P2_U3199(p2_u3199), .P2_U3198(p2_u3198), .P2_U3197(p2_u3197), .P2_U3196(p2_u3196), .P2_U3195(p2_u3195), .P2_U3194(p2_u3194), .P2_U3193(p2_u3193), .P2_U3192(p2_u3192), .P2_U3191(p2_u3191), .P2_U3190(p2_u3190), .P2_U3189(p2_u3189), .P2_U3188(p2_u3188), .P2_U3187(p2_u3187), .P2_U3186(p2_u3186), .P2_U3185(p2_u3185), .P2_U3088(p2_u3088), .P2_U3087(p2_u3087), .P2_U3947(p2_u3947), .P3_U3295(p3_u3295), .P3_U3294(p3_u3294), .P3_U3293(p3_u3293), .P3_U3292(p3_u3292), .P3_U3291(p3_u3291), .P3_U3290(p3_u3290), .P3_U3289(p3_u3289), .P3_U3288(p3_u3288), .P3_U3287(p3_u3287), .P3_U3286(p3_u3286), .P3_U3285(p3_u3285), .P3_U3284(p3_u3284), .P3_U3283(p3_u3283), .P3_U3282(p3_u3282), .P3_U3281(p3_u3281), .P3_U3280(p3_u3280), .P3_U3279(p3_u3279), .P3_U3278(p3_u3278), .P3_U3277(p3_u3277), .P3_U3276(p3_u3276), .P3_U3275(p3_u3275), .P3_U3274(p3_u3274), .P3_U3273(p3_u3273), .P3_U3272(p3_u3272), .P3_U3271(p3_u3271), .P3_U3270(p3_u3270), .P3_U3269(p3_u3269), .P3_U3268(p3_u3268), .P3_U3267(p3_u3267), .P3_U3266(p3_u3266), .P3_U3265(p3_u3265), .P3_U3264(p3_u3264), .P3_U3376(p3_u3376), .P3_U3377(p3_u3377), .P3_U3263(p3_u3263), .P3_U3262(p3_u3262), .P3_U3261(p3_u3261), .P3_U3260(p3_u3260), .P3_U3259(p3_u3259), .P3_U3258(p3_u3258), .P3_U3257(p3_u3257), .P3_U3256(p3_u3256), .P3_U3255(p3_u3255), .P3_U3254(p3_u3254), .P3_U3253(p3_u3253), .P3_U3252(p3_u3252), .P3_U3251(p3_u3251), .P3_U3250(p3_u3250), .P3_U3249(p3_u3249), .P3_U3248(p3_u3248), .P3_U3247(p3_u3247), .P3_U3246(p3_u3246), .P3_U3245(p3_u3245), .P3_U3244(p3_u3244), .P3_U3243(p3_u3243), .P3_U3242(p3_u3242), .P3_U3241(p3_u3241), .P3_U3240(p3_u3240), .P3_U3239(p3_u3239), .P3_U3238(p3_u3238), .P3_U3237(p3_u3237), .P3_U3236(p3_u3236), .P3_U3235(p3_u3235), .P3_U3234(p3_u3234), .P3_U3390(p3_u3390), .P3_U3393(p3_u3393), .P3_U3396(p3_u3396), .P3_U3399(p3_u3399), .P3_U3402(p3_u3402), .P3_U3405(p3_u3405), .P3_U3408(p3_u3408), .P3_U3411(p3_u3411), .P3_U3414(p3_u3414), .P3_U3417(p3_u3417), .P3_U3420(p3_u3420), .P3_U3423(p3_u3423), .P3_U3426(p3_u3426), .P3_U3429(p3_u3429), .P3_U3432(p3_u3432), .P3_U3435(p3_u3435), .P3_U3438(p3_u3438), .P3_U3441(p3_u3441), .P3_U3444(p3_u3444), .P3_U3446(p3_u3446), .P3_U3447(p3_u3447), .P3_U3448(p3_u3448), .P3_U3449(p3_u3449), .P3_U3450(p3_u3450), .P3_U3451(p3_u3451), .P3_U3452(p3_u3452), .P3_U3453(p3_u3453), .P3_U3454(p3_u3454), .P3_U3455(p3_u3455), .P3_U3456(p3_u3456), .P3_U3457(p3_u3457), .P3_U3458(p3_u3458), .P3_U3459(p3_u3459), .P3_U3460(p3_u3460), .P3_U3461(p3_u3461), .P3_U3462(p3_u3462), .P3_U3463(p3_u3463), .P3_U3464(p3_u3464), .P3_U3465(p3_u3465), .P3_U3466(p3_u3466), .P3_U3467(p3_u3467), .P3_U3468(p3_u3468), .P3_U3469(p3_u3469), .P3_U3470(p3_u3470), .P3_U3471(p3_u3471), .P3_U3472(p3_u3472), .P3_U3473(p3_u3473), .P3_U3474(p3_u3474), .P3_U3475(p3_u3475), .P3_U3476(p3_u3476), .P3_U3477(p3_u3477), .P3_U3478(p3_u3478), .P3_U3479(p3_u3479), .P3_U3480(p3_u3480), .P3_U3481(p3_u3481), .P3_U3482(p3_u3482), .P3_U3483(p3_u3483), .P3_U3484(p3_u3484), .P3_U3485(p3_u3485), .P3_U3486(p3_u3486), .P3_U3487(p3_u3487), .P3_U3488(p3_u3488), .P3_U3489(p3_u3489), .P3_U3490(p3_u3490), .P3_U3233(p3_u3233), .P3_U3232(p3_u3232), .P3_U3231(p3_u3231), .P3_U3230(p3_u3230), .P3_U3229(p3_u3229), .P3_U3228(p3_u3228), .P3_U3227(p3_u3227), .P3_U3226(p3_u3226), .P3_U3225(p3_u3225), .P3_U3224(p3_u3224), .P3_U3223(p3_u3223), .P3_U3222(p3_u3222), .P3_U3221(p3_u3221), .P3_U3220(p3_u3220), .P3_U3219(p3_u3219), .P3_U3218(p3_u3218), .P3_U3217(p3_u3217), .P3_U3216(p3_u3216), .P3_U3215(p3_u3215), .P3_U3214(p3_u3214), .P3_U3213(p3_u3213), .P3_U3212(p3_u3212), .P3_U3211(p3_u3211), .P3_U3210(p3_u3210), .P3_U3209(p3_u3209), .P3_U3208(p3_u3208), .P3_U3207(p3_u3207), .P3_U3206(p3_u3206), .P3_U3205(p3_u3205), .P3_U3204(p3_u3204), .P3_U3203(p3_u3203), .P3_U3202(p3_u3202), .P3_U3201(p3_u3201), .P3_U3200(p3_u3200), .P3_U3199(p3_u3199), .P3_U3198(p3_u3198), .P3_U3197(p3_u3197), .P3_U3196(p3_u3196), .P3_U3195(p3_u3195), .P3_U3194(p3_u3194), .P3_U3193(p3_u3193), .P3_U3192(p3_u3192), .P3_U3191(p3_u3191), .P3_U3190(p3_u3190), .P3_U3189(p3_u3189), .P3_U3188(p3_u3188), .P3_U3187(p3_u3187), .P3_U3186(p3_u3186), .P3_U3185(p3_u3185), .P3_U3184(p3_u3184), .P3_U3183(p3_u3183), .P3_U3182(p3_u3182), .P3_U3491(p3_u3491), .P3_U3492(p3_u3492), .P3_U3493(p3_u3493), .P3_U3494(p3_u3494), .P3_U3495(p3_u3495), .P3_U3496(p3_u3496), .P3_U3497(p3_u3497), .P3_U3498(p3_u3498), .P3_U3499(p3_u3499), .P3_U3500(p3_u3500), .P3_U3501(p3_u3501), .P3_U3502(p3_u3502), .P3_U3503(p3_u3503), .P3_U3504(p3_u3504), .P3_U3505(p3_u3505), .P3_U3506(p3_u3506), .P3_U3507(p3_u3507), .P3_U3508(p3_u3508), .P3_U3509(p3_u3509), .P3_U3510(p3_u3510), .P3_U3511(p3_u3511), .P3_U3512(p3_u3512), .P3_U3513(p3_u3513), .P3_U3514(p3_u3514), .P3_U3515(p3_u3515), .P3_U3516(p3_u3516), .P3_U3517(p3_u3517), .P3_U3518(p3_u3518), .P3_U3519(p3_u3519), .P3_U3520(p3_u3520), .P3_U3521(p3_u3521), .P3_U3522(p3_u3522), .P3_U3296(p3_u3296), .P3_U3181(p3_u3181), .P3_U3180(p3_u3180), .P3_U3179(p3_u3179), .P3_U3178(p3_u3178), .P3_U3177(p3_u3177), .P3_U3176(p3_u3176), .P3_U3175(p3_u3175), .P3_U3174(p3_u3174), .P3_U3173(p3_u3173), .P3_U3172(p3_u3172), .P3_U3171(p3_u3171), .P3_U3170(p3_u3170), .P3_U3169(p3_u3169), .P3_U3168(p3_u3168), .P3_U3167(p3_u3167), .P3_U3166(p3_u3166), .P3_U3165(p3_u3165), .P3_U3164(p3_u3164), .P3_U3163(p3_u3163), .P3_U3162(p3_u3162), .P3_U3161(p3_u3161), .P3_U3160(p3_u3160), .P3_U3159(p3_u3159), .P3_U3158(p3_u3158), .P3_U3157(p3_u3157), .P3_U3156(p3_u3156), .P3_U3155(p3_u3155), .P3_U3154(p3_u3154), .P3_U3153(p3_u3153), .P3_U3151(p3_u3151), .P3_U3150(p3_u3150), .P3_U3897(p3_u3897));

integer i=0;
always @ (posedge clk) begin
	vec = input_vec_mem[i];
	$monitor(vec);
	i = i + 1;

end

always @ (negedge clk)begin
	$fdisplay ( fh_w, sub_1596_u4, sub_1596_u62, sub_1596_u63, sub_1596_u64, sub_1596_u65, sub_1596_u66, sub_1596_u67, sub_1596_u68, sub_1596_u69, sub_1596_u70, sub_1596_u54, sub_1596_u55, sub_1596_u56, sub_1596_u57, sub_1596_u58, sub_1596_u59, sub_1596_u60, sub_1596_u61, sub_1596_u5, sub_1596_u53, u29, u28, p1_u3355, p1_u3354, p1_u3353, p1_u3352, p1_u3351, p1_u3350, p1_u3349, p1_u3348, p1_u3347, p1_u3346, p1_u3345, p1_u3344, p1_u3343, p1_u3342, p1_u3341, p1_u3340, p1_u3339, p1_u3338, p1_u3337, p1_u3336, p1_u3335, p1_u3334, p1_u3333, p1_u3332, p1_u3331, p1_u3330, p1_u3329, p1_u3328, p1_u3327, p1_u3326, p1_u3325, p1_u3324, p1_u3445, p1_u3446, p1_u3323, p1_u3322, p1_u3321, p1_u3320, p1_u3319, p1_u3318, p1_u3317, p1_u3316, p1_u3315, p1_u3314, p1_u3313, p1_u3312, p1_u3311, p1_u3310, p1_u3309, p1_u3308, p1_u3307, p1_u3306, p1_u3305, p1_u3304, p1_u3303, p1_u3302, p1_u3301, p1_u3300, p1_u3299, p1_u3298, p1_u3297, p1_u3296, p1_u3295, p1_u3294, p1_u3459, p1_u3462, p1_u3465, p1_u3468, p1_u3471, p1_u3474, p1_u3477, p1_u3480, p1_u3483, p1_u3486, p1_u3489, p1_u3492, p1_u3495, p1_u3498, p1_u3501, p1_u3504, p1_u3507, p1_u3510, p1_u3513, p1_u3515, p1_u3516, p1_u3517, p1_u3518, p1_u3519, p1_u3520, p1_u3521, p1_u3522, p1_u3523, p1_u3524, p1_u3525, p1_u3526, p1_u3527, p1_u3528, p1_u3529, p1_u3530, p1_u3531, p1_u3532, p1_u3533, p1_u3534, p1_u3535, p1_u3536, p1_u3537, p1_u3538, p1_u3539, p1_u3540, p1_u3541, p1_u3542, p1_u3543, p1_u3544, p1_u3545, p1_u3546, p1_u3547, p1_u3548, p1_u3549, p1_u3550, p1_u3551, p1_u3552, p1_u3553, p1_u3554, p1_u3555, p1_u3556, p1_u3557, p1_u3558, p1_u3559, p1_u3293, p1_u3292, p1_u3291, p1_u3290, p1_u3289, p1_u3288, p1_u3287, p1_u3286, p1_u3285, p1_u3284, p1_u3283, p1_u3282, p1_u3281, p1_u3280, p1_u3279, p1_u3278, p1_u3277, p1_u3276, p1_u3275, p1_u3274, p1_u3273, p1_u3272, p1_u3271, p1_u3270, p1_u3269, p1_u3268, p1_u3267, p1_u3266, p1_u3265, p1_u3356, p1_u3264, p1_u3263, p1_u3262, p1_u3261, p1_u3260, p1_u3259, p1_u3258, p1_u3257, p1_u3256, p1_u3255, p1_u3254, p1_u3253, p1_u3252, p1_u3251, p1_u3250, p1_u3249, p1_u3248, p1_u3247, p1_u3246, p1_u3245, p1_u3244, p1_u3243, p1_u3560, p1_u3561, p1_u3562, p1_u3563, p1_u3564, p1_u3565, p1_u3566, p1_u3567, p1_u3568, p1_u3569, p1_u3570, p1_u3571, p1_u3572, p1_u3573, p1_u3574, p1_u3575, p1_u3576, p1_u3577, p1_u3578, p1_u3579, p1_u3580, p1_u3581, p1_u3582, p1_u3583, p1_u3584, p1_u3585, p1_u3586, p1_u3587, p1_u3588, p1_u3589, p1_u3590, p1_u3591, p1_u3242, p1_u3241, p1_u3240, p1_u3239, p1_u3238, p1_u3237, p1_u3236, p1_u3235, p1_u3234, p1_u3233, p1_u3232, p1_u3231, p1_u3230, p1_u3229, p1_u3228, p1_u3227, p1_u3226, p1_u3225, p1_u3224, p1_u3223, p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218, p1_u3217, p1_u3216, p1_u3215, p1_u3214, p1_u3213, p1_u3086, p1_u3085, p1_u4016, p2_u3327, p2_u3326, p2_u3325, p2_u3324, p2_u3323, p2_u3322, p2_u3321, p2_u3320, p2_u3319, p2_u3318, p2_u3317, p2_u3316, p2_u3315, p2_u3314, p2_u3313, p2_u3312, p2_u3311, p2_u3310, p2_u3309, p2_u3308, p2_u3307, p2_u3306, p2_u3305, p2_u3304, p2_u3303, p2_u3302, p2_u3301, p2_u3300, p2_u3299, p2_u3298, p2_u3297, p2_u3296, p2_u3416, p2_u3417, p2_u3295, p2_u3294, p2_u3293, p2_u3292, p2_u3291, p2_u3290, p2_u3289, p2_u3288, p2_u3287, p2_u3286, p2_u3285, p2_u3284, p2_u3283, p2_u3282, p2_u3281, p2_u3280, p2_u3279, p2_u3278, p2_u3277, p2_u3276, p2_u3275, p2_u3274, p2_u3273, p2_u3272, p2_u3271, p2_u3270, p2_u3269, p2_u3268, p2_u3267, p2_u3266, p2_u3430, p2_u3433, p2_u3436, p2_u3439, p2_u3442, p2_u3445, p2_u3448, p2_u3451, p2_u3454, p2_u3457, p2_u3460, p2_u3463, p2_u3466, p2_u3469, p2_u3472, p2_u3475, p2_u3478, p2_u3481, p2_u3484, p2_u3486, p2_u3487, p2_u3488, p2_u3489, p2_u3490, p2_u3491, p2_u3492, p2_u3493, p2_u3494, p2_u3495, p2_u3496, p2_u3497, p2_u3498, p2_u3499, p2_u3500, p2_u3501, p2_u3502, p2_u3503, p2_u3504, p2_u3505, p2_u3506, p2_u3507, p2_u3508, p2_u3509, p2_u3510, p2_u3511, p2_u3512, p2_u3513, p2_u3514, p2_u3515, p2_u3516, p2_u3517, p2_u3518, p2_u3519, p2_u3520, p2_u3521, p2_u3522, p2_u3523, p2_u3524, p2_u3525, p2_u3526, p2_u3527, p2_u3528, p2_u3529, p2_u3530, p2_u3265, p2_u3264, p2_u3263, p2_u3262, p2_u3261, p2_u3260, p2_u3259, p2_u3258, p2_u3257, p2_u3256, p2_u3255, p2_u3254, p2_u3253, p2_u3252, p2_u3251, p2_u3250, p2_u3249, p2_u3248, p2_u3247, p2_u3246, p2_u3245, p2_u3244, p2_u3243, p2_u3242, p2_u3241, p2_u3240, p2_u3239, p2_u3238, p2_u3237, p2_u3236, p2_u3235, p2_u3234, p2_u3233, p2_u3232, p2_u3231, p2_u3230, p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225, p2_u3224, p2_u3223, p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218, p2_u3217, p2_u3216, p2_u3215, p2_u3214, p2_u3531, p2_u3532, p2_u3533, p2_u3534, p2_u3535, p2_u3536, p2_u3537, p2_u3538, p2_u3539, p2_u3540, p2_u3541, p2_u3542, p2_u3543, p2_u3544, p2_u3545, p2_u3546, p2_u3547, p2_u3548, p2_u3549, p2_u3550, p2_u3551, p2_u3552, p2_u3553, p2_u3554, p2_u3555, p2_u3556, p2_u3557, p2_u3558, p2_u3559, p2_u3560, p2_u3561, p2_u3562, p2_u3328, p2_u3213, p2_u3212, p2_u3211, p2_u3210, p2_u3209, p2_u3208, p2_u3207, p2_u3206, p2_u3205, p2_u3204, p2_u3203, p2_u3202, p2_u3201, p2_u3200, p2_u3199, p2_u3198, p2_u3197, p2_u3196, p2_u3195, p2_u3194, p2_u3193, p2_u3192, p2_u3191, p2_u3190, p2_u3189, p2_u3188, p2_u3187, p2_u3186, p2_u3185, p2_u3088, p2_u3087, p2_u3947, p3_u3295, p3_u3294, p3_u3293, p3_u3292, p3_u3291, p3_u3290, p3_u3289, p3_u3288, p3_u3287, p3_u3286, p3_u3285, p3_u3284, p3_u3283, p3_u3282, p3_u3281, p3_u3280, p3_u3279, p3_u3278, p3_u3277, p3_u3276, p3_u3275, p3_u3274, p3_u3273, p3_u3272, p3_u3271, p3_u3270, p3_u3269, p3_u3268, p3_u3267, p3_u3266, p3_u3265, p3_u3264, p3_u3376, p3_u3377, p3_u3263, p3_u3262, p3_u3261, p3_u3260, p3_u3259, p3_u3258, p3_u3257, p3_u3256, p3_u3255, p3_u3254, p3_u3253, p3_u3252, p3_u3251, p3_u3250, p3_u3249, p3_u3248, p3_u3247, p3_u3246, p3_u3245, p3_u3244, p3_u3243, p3_u3242, p3_u3241, p3_u3240, p3_u3239, p3_u3238, p3_u3237, p3_u3236, p3_u3235, p3_u3234, p3_u3390, p3_u3393, p3_u3396, p3_u3399, p3_u3402, p3_u3405, p3_u3408, p3_u3411, p3_u3414, p3_u3417, p3_u3420, p3_u3423, p3_u3426, p3_u3429, p3_u3432, p3_u3435, p3_u3438, p3_u3441, p3_u3444, p3_u3446, p3_u3447, p3_u3448, p3_u3449, p3_u3450, p3_u3451, p3_u3452, p3_u3453, p3_u3454, p3_u3455, p3_u3456, p3_u3457, p3_u3458, p3_u3459, p3_u3460, p3_u3461, p3_u3462, p3_u3463, p3_u3464, p3_u3465, p3_u3466, p3_u3467, p3_u3468, p3_u3469, p3_u3470, p3_u3471, p3_u3472, p3_u3473, p3_u3474, p3_u3475, p3_u3476, p3_u3477, p3_u3478, p3_u3479, p3_u3480, p3_u3481, p3_u3482, p3_u3483, p3_u3484, p3_u3485, p3_u3486, p3_u3487, p3_u3488, p3_u3489, p3_u3490, p3_u3233, p3_u3232, p3_u3231, p3_u3230, p3_u3229, p3_u3228, p3_u3227, p3_u3226, p3_u3225, p3_u3224, p3_u3223, p3_u3222, p3_u3221, p3_u3220, p3_u3219, p3_u3218, p3_u3217, p3_u3216, p3_u3215, p3_u3214, p3_u3213, p3_u3212, p3_u3211, p3_u3210, p3_u3209, p3_u3208, p3_u3207, p3_u3206, p3_u3205, p3_u3204, p3_u3203, p3_u3202, p3_u3201, p3_u3200, p3_u3199, p3_u3198, p3_u3197, p3_u3196, p3_u3195, p3_u3194, p3_u3193, p3_u3192, p3_u3191, p3_u3190, p3_u3189, p3_u3188, p3_u3187, p3_u3186, p3_u3185, p3_u3184, p3_u3183, p3_u3182, p3_u3491, p3_u3492, p3_u3493, p3_u3494, p3_u3495, p3_u3496, p3_u3497, p3_u3498, p3_u3499, p3_u3500, p3_u3501, p3_u3502, p3_u3503, p3_u3504, p3_u3505, p3_u3506, p3_u3507, p3_u3508, p3_u3509, p3_u3510, p3_u3511, p3_u3512, p3_u3513, p3_u3514, p3_u3515, p3_u3516, p3_u3517, p3_u3518, p3_u3519, p3_u3520, p3_u3521, p3_u3522, p3_u3296, p3_u3181, p3_u3180, p3_u3179, p3_u3178, p3_u3177, p3_u3176, p3_u3175, p3_u3174, p3_u3173, p3_u3172, p3_u3171, p3_u3170, p3_u3169, p3_u3168, p3_u3167, p3_u3166, p3_u3165, p3_u3164, p3_u3163, p3_u3162, p3_u3161, p3_u3160, p3_u3159, p3_u3158, p3_u3157, p3_u3156, p3_u3155, p3_u3154, p3_u3153, p3_u3151, p3_u3150, p3_u3897);
	if(i == vec_length)begin
		$finish;
	end
end

integer fh_w;
initial begin
	fh_w = $fopen(`out_file, "w");
end
 
initial begin
	//$fsdbDumpfile("SET.fsdb");
	//$fsdbDumpvars;
	//$fsdbDumpMDA;
	$dumpfile("test_result.vcd");
    $dumpvars;

end
endmodule
