// b21
// 522 inputs  (32 PIs + 490 PPIs)
// 512 outputs (22 POs + 490 PPOs)
// 20027 gates (16938 gates + 3089 inverters + 0 buffers )
// ( 2196 AND + 542 OR + 14073 NAND + 127 NOR )
// Time: Wed Mar 25 17:47:25 2009
// All copyrigh from NCKU EE TestLAB, Taiwan. [2008.12. WCL]

module b21_ras ( P1_U3353 , P1_U3352 , P1_U3351 , P1_U3350 , P1_U3349 , P1_U3348 ,
             P1_U3347 , P1_U3346 , P1_U3345 , P1_U3344 , P1_U3343 , P1_U3342 ,
             P1_U3341 , P1_U3340 , P1_U3339 , P1_U3338 , P1_U3337 , P1_U3336 ,
             P1_U3335 , P1_U3334 , P1_U3333 , P1_U3332 , P1_U3331 , P1_U3330 ,
             P1_U3329 , P1_U3328 , P1_U3327 , P1_U3326 , P1_U3325 , P1_U3324 ,
             P1_U3323 , P1_U3322 , P1_U3440 , P1_U3441 , P1_U3321 , P1_U3320 ,
             P1_U3319 , P1_U3318 , P1_U3317 , P1_U3316 , P1_U3315 , P1_U3314 ,
             P1_U3313 , P1_U3312 , P1_U3311 , P1_U3310 , P1_U3309 , P1_U3308 ,
             P1_U3307 , P1_U3306 , P1_U3305 , P1_U3304 , P1_U3303 , P1_U3302 ,
             P1_U3301 , P1_U3300 , P1_U3299 , P1_U3298 , P1_U3297 , P1_U3296 ,
             P1_U3295 , P1_U3294 , P1_U3293 , P1_U3292 , P1_U3454 , P1_U3457 ,
             P1_U3460 , P1_U3463 , P1_U3466 , P1_U3469 , P1_U3472 , P1_U3475 ,
             P1_U3478 , P1_U3481 , P1_U3484 , P1_U3487 , P1_U3490 , P1_U3493 ,
             P1_U3496 , P1_U3499 , P1_U3502 , P1_U3505 , P1_U3508 , P1_U3510 ,
             P1_U3511 , P1_U3512 , P1_U3513 , P1_U3514 , P1_U3515 , P1_U3516 ,
             P1_U3517 , P1_U3518 , P1_U3519 , P1_U3520 , P1_U3521 , P1_U3522 ,
             P1_U3523 , P1_U3524 , P1_U3525 , P1_U3526 , P1_U3527 , P1_U3528 ,
             P1_U3529 , P1_U3530 , P1_U3531 , P1_U3532 , P1_U3533 , P1_U3534 ,
             P1_U3535 , P1_U3536 , P1_U3537 , P1_U3538 , P1_U3539 , P1_U3540 ,
             P1_U3541 , P1_U3542 , P1_U3543 , P1_U3544 , P1_U3545 , P1_U3546 ,
             P1_U3547 , P1_U3548 , P1_U3549 , P1_U3550 , P1_U3551 , P1_U3552 ,
             P1_U3553 , P1_U3554 , P1_U3291 , P1_U3290 , P1_U3289 , P1_U3288 ,
             P1_U3287 , P1_U3286 , P1_U3285 , P1_U3284 , P1_U3283 , P1_U3282 ,
             P1_U3281 , P1_U3280 , P1_U3279 , P1_U3278 , P1_U3277 , P1_U3276 ,
             P1_U3275 , P1_U3274 , P1_U3273 , P1_U3272 , P1_U3271 , P1_U3270 ,
             P1_U3269 , P1_U3268 , P1_U3267 , P1_U3266 , P1_U3265 , P1_U3264 ,
             P1_U3263 , P1_U3355 , P1_U3262 , P1_U3261 , P1_U3260 , P1_U3259 ,
             P1_U3258 , P1_U3257 , P1_U3256 , P1_U3255 , P1_U3254 , P1_U3253 ,
             P1_U3252 , P1_U3251 , P1_U3250 , P1_U3249 , P1_U3248 , P1_U3247 ,
             P1_U3246 , P1_U3245 , P1_U3244 , P1_U3243 , P1_U3242 , P1_U3241 ,
             P1_U3555 , P1_U3556 , P1_U3557 , P1_U3558 , P1_U3559 , P1_U3560 ,
             P1_U3561 , P1_U3562 , P1_U3563 , P1_U3564 , P1_U3565 , P1_U3566 ,
             P1_U3567 , P1_U3568 , P1_U3569 , P1_U3570 , P1_U3571 , P1_U3572 ,
             P1_U3573 , P1_U3574 , P1_U3575 , P1_U3576 , P1_U3577 , P1_U3578 ,
             P1_U3579 , P1_U3580 , P1_U3581 , P1_U3582 , P1_U3583 , P1_U3584 ,
             P1_U3585 , P1_U3586 , P1_U3240 , P1_U3239 , P1_U3238 , P1_U3237 ,
             P1_U3236 , P1_U3235 , P1_U3234 , P1_U3233 , P1_U3232 , P1_U3231 ,
             P1_U3230 , P1_U3229 , P1_U3228 , P1_U3227 , P1_U3226 , P1_U3225 ,
             P1_U3224 , P1_U3223 , P1_U3222 , P1_U3221 , P1_U3220 , P1_U3219 ,
             P1_U3218 , P1_U3217 , P1_U3216 , P1_U3215 , P1_U3214 , P1_U3213 ,
             P1_U3212 , P1_U3211 , P1_U3084 , P1_U3083 , P1_U4006 , P2_U3358 ,
             P2_U3357 , P2_U3356 , P2_U3355 , P2_U3354 , P2_U3353 , P2_U3352 ,
             P2_U3351 , P2_U3350 , P2_U3349 , P2_U3348 , P2_U3347 , P2_U3346 ,
             P2_U3345 , P2_U3344 , P2_U3343 , P2_U3342 , P2_U3341 , P2_U3340 ,
             P2_U3339 , P2_U3338 , P2_U3337 , P2_U3336 , P2_U3335 , P2_U3334 ,
             P2_U3333 , P2_U3332 , P2_U3331 , P2_U3330 , P2_U3329 , P2_U3328 ,
             P2_U3327 , P2_U3437 , P2_U3438 , P2_U3326 , P2_U3325 , P2_U3324 ,
             P2_U3323 , P2_U3322 , P2_U3321 , P2_U3320 , P2_U3319 , P2_U3318 ,
             P2_U3317 , P2_U3316 , P2_U3315 , P2_U3314 , P2_U3313 , P2_U3312 ,
             P2_U3311 , P2_U3310 , P2_U3309 , P2_U3308 , P2_U3307 , P2_U3306 ,
             P2_U3305 , P2_U3304 , P2_U3303 , P2_U3302 , P2_U3301 , P2_U3300 ,
             P2_U3299 , P2_U3298 , P2_U3297 , P2_U3451 , P2_U3454 , P2_U3457 ,
             P2_U3460 , P2_U3463 , P2_U3466 , P2_U3469 , P2_U3472 , P2_U3475 ,
             P2_U3478 , P2_U3481 , P2_U3484 , P2_U3487 , P2_U3490 , P2_U3493 ,
             P2_U3496 , P2_U3499 , P2_U3502 , P2_U3505 , P2_U3507 , P2_U3508 ,
             P2_U3509 , P2_U3510 , P2_U3511 , P2_U3512 , P2_U3513 , P2_U3514 ,
             P2_U3515 , P2_U3516 , P2_U3517 , P2_U3518 , P2_U3519 , P2_U3520 ,
             P2_U3521 , P2_U3522 , P2_U3523 , P2_U3524 , P2_U3525 , P2_U3526 ,
             P2_U3527 , P2_U3528 , P2_U3529 , P2_U3530 , P2_U3531 , P2_U3532 ,
             P2_U3533 , P2_U3534 , P2_U3535 , P2_U3536 , P2_U3537 , P2_U3538 ,
             P2_U3539 , P2_U3540 , P2_U3541 , P2_U3542 , P2_U3543 , P2_U3544 ,
             P2_U3545 , P2_U3546 , P2_U3547 , P2_U3548 , P2_U3549 , P2_U3550 ,
             P2_U3551 , P2_U3296 , P2_U3295 , P2_U3294 , P2_U3293 , P2_U3292 ,
             P2_U3291 , P2_U3290 , P2_U3289 , P2_U3288 , P2_U3287 , P2_U3286 ,
             P2_U3285 , P2_U3284 , P2_U3283 , P2_U3282 , P2_U3281 , P2_U3280 ,
             P2_U3279 , P2_U3278 , P2_U3277 , P2_U3276 , P2_U3275 , P2_U3274 ,
             P2_U3273 , P2_U3272 , P2_U3271 , P2_U3270 , P2_U3269 , P2_U3268 ,
             P2_U3267 , P2_U3266 , P2_U3265 , P2_U3264 , P2_U3263 , P2_U3262 ,
             P2_U3261 , P2_U3260 , P2_U3259 , P2_U3258 , P2_U3257 , P2_U3256 ,
             P2_U3255 , P2_U3254 , P2_U3253 , P2_U3252 , P2_U3251 , P2_U3250 ,
             P2_U3249 , P2_U3248 , P2_U3247 , P2_U3246 , P2_U3245 , P2_U3552 ,
             P2_U3553 , P2_U3554 , P2_U3555 , P2_U3556 , P2_U3557 , P2_U3558 ,
             P2_U3559 , P2_U3560 , P2_U3561 , P2_U3562 , P2_U3563 , P2_U3564 ,
             P2_U3565 , P2_U3566 , P2_U3567 , P2_U3568 , P2_U3569 , P2_U3570 ,
             P2_U3571 , P2_U3572 , P2_U3573 , P2_U3574 , P2_U3575 , P2_U3576 ,
             P2_U3577 , P2_U3578 , P2_U3579 , P2_U3580 , P2_U3581 , P2_U3582 ,
             P2_U3583 , P2_U3244 , P2_U3243 , P2_U3242 , P2_U3241 , P2_U3240 ,
             P2_U3239 , P2_U3238 , P2_U3237 , P2_U3236 , P2_U3235 , P2_U3234 ,
             P2_U3233 , P2_U3232 , P2_U3231 , P2_U3230 , P2_U3229 , P2_U3228 ,
             P2_U3227 , P2_U3226 , P2_U3225 , P2_U3224 , P2_U3223 , P2_U3222 ,
             P2_U3221 , P2_U3220 , P2_U3219 , P2_U3218 , P2_U3217 , P2_U3216 ,
             P2_U3215 , P2_U3152 , P2_U3151 , P2_U3966 , ADD_1071_U4 , ADD_1071_U55 ,
             ADD_1071_U56 , ADD_1071_U57 , ADD_1071_U58 , ADD_1071_U59 , ADD_1071_U60 , ADD_1071_U61 ,
             ADD_1071_U62 , ADD_1071_U63 , ADD_1071_U47 , ADD_1071_U48 , ADD_1071_U49 , ADD_1071_U50 ,
             ADD_1071_U51 , ADD_1071_U52 , ADD_1071_U53 , ADD_1071_U54 , ADD_1071_U5 , ADD_1071_U46 ,
             U126 , U123 ,
             P1_IR_REG_0_ , P1_IR_REG_1_ , P1_IR_REG_2_ , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ ,
             P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_10_ , P1_IR_REG_11_ ,
             P1_IR_REG_12_ , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_ ,
             P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_20_ , P1_IR_REG_21_ , P1_IR_REG_22_ , P1_IR_REG_23_ ,
             P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ , P1_IR_REG_27_ , P1_IR_REG_28_ , P1_IR_REG_29_ ,
             P1_IR_REG_30_ , P1_IR_REG_31_ , P1_D_REG_0_ , P1_D_REG_1_ , P1_D_REG_2_ , P1_D_REG_3_ ,
             P1_D_REG_4_ , P1_D_REG_5_ , P1_D_REG_6_ , P1_D_REG_7_ , P1_D_REG_8_ , P1_D_REG_9_ ,
             P1_D_REG_10_ , P1_D_REG_11_ , P1_D_REG_12_ , P1_D_REG_13_ , P1_D_REG_14_ , P1_D_REG_15_ ,
             P1_D_REG_16_ , P1_D_REG_17_ , P1_D_REG_18_ , P1_D_REG_19_ , P1_D_REG_20_ , P1_D_REG_21_ ,
             P1_D_REG_22_ , P1_D_REG_23_ , P1_D_REG_24_ , P1_D_REG_25_ , P1_D_REG_26_ , P1_D_REG_27_ ,
             P1_D_REG_28_ , P1_D_REG_29_ , P1_D_REG_30_ , P1_D_REG_31_ , P1_REG0_REG_0_ , P1_REG0_REG_1_ ,
             P1_REG0_REG_2_ , P1_REG0_REG_3_ , P1_REG0_REG_4_ , P1_REG0_REG_5_ , P1_REG0_REG_6_ , P1_REG0_REG_7_ ,
             P1_REG0_REG_8_ , P1_REG0_REG_9_ , P1_REG0_REG_10_ , P1_REG0_REG_11_ , P1_REG0_REG_12_ , P1_REG0_REG_13_ ,
             P1_REG0_REG_14_ , P1_REG0_REG_15_ , P1_REG0_REG_16_ , P1_REG0_REG_17_ , P1_REG0_REG_18_ , P1_REG0_REG_19_ ,
             P1_REG0_REG_20_ , P1_REG0_REG_21_ , P1_REG0_REG_22_ , P1_REG0_REG_23_ , P1_REG0_REG_24_ , P1_REG0_REG_25_ ,
             P1_REG0_REG_26_ , P1_REG0_REG_27_ , P1_REG0_REG_28_ , P1_REG0_REG_29_ , P1_REG0_REG_30_ , P1_REG0_REG_31_ ,
             P1_REG1_REG_0_ , P1_REG1_REG_1_ , P1_REG1_REG_2_ , P1_REG1_REG_3_ , P1_REG1_REG_4_ , P1_REG1_REG_5_ ,
             P1_REG1_REG_6_ , P1_REG1_REG_7_ , P1_REG1_REG_8_ , P1_REG1_REG_9_ , P1_REG1_REG_10_ , P1_REG1_REG_11_ ,
             P1_REG1_REG_12_ , P1_REG1_REG_13_ , P1_REG1_REG_14_ , P1_REG1_REG_15_ , P1_REG1_REG_16_ , P1_REG1_REG_17_ ,
             P1_REG1_REG_18_ , P1_REG1_REG_19_ , P1_REG1_REG_20_ , P1_REG1_REG_21_ , P1_REG1_REG_22_ , P1_REG1_REG_23_ ,
             P1_REG1_REG_24_ , P1_REG1_REG_25_ , P1_REG1_REG_26_ , P1_REG1_REG_27_ , P1_REG1_REG_28_ , P1_REG1_REG_29_ ,
             P1_REG1_REG_30_ , P1_REG1_REG_31_ , P1_REG2_REG_0_ , P1_REG2_REG_1_ , P1_REG2_REG_2_ , P1_REG2_REG_3_ ,
             P1_REG2_REG_4_ , P1_REG2_REG_5_ , P1_REG2_REG_6_ , P1_REG2_REG_7_ , P1_REG2_REG_8_ , P1_REG2_REG_9_ ,
             P1_REG2_REG_10_ , P1_REG2_REG_11_ , P1_REG2_REG_12_ , P1_REG2_REG_13_ , P1_REG2_REG_14_ , P1_REG2_REG_15_ ,
             P1_REG2_REG_16_ , P1_REG2_REG_17_ , P1_REG2_REG_18_ , P1_REG2_REG_19_ , P1_REG2_REG_20_ , P1_REG2_REG_21_ ,
             P1_REG2_REG_22_ , P1_REG2_REG_23_ , P1_REG2_REG_24_ , P1_REG2_REG_25_ , P1_REG2_REG_26_ , P1_REG2_REG_27_ ,
             P1_REG2_REG_28_ , P1_REG2_REG_29_ , P1_REG2_REG_30_ , P1_REG2_REG_31_ , P1_ADDR_REG_19_ , P1_ADDR_REG_18_ ,
             P1_ADDR_REG_17_ , P1_ADDR_REG_16_ , P1_ADDR_REG_15_ , P1_ADDR_REG_14_ , P1_ADDR_REG_13_ , P1_ADDR_REG_12_ ,
             P1_ADDR_REG_11_ , P1_ADDR_REG_10_ , P1_ADDR_REG_9_ , P1_ADDR_REG_8_ , P1_ADDR_REG_7_ , P1_ADDR_REG_6_ ,
             P1_ADDR_REG_5_ , P1_ADDR_REG_4_ , P1_ADDR_REG_3_ , P1_ADDR_REG_2_ , P1_ADDR_REG_1_ , P1_ADDR_REG_0_ ,
             P1_DATAO_REG_0_ , P1_DATAO_REG_1_ , P1_DATAO_REG_2_ , P1_DATAO_REG_3_ , P1_DATAO_REG_4_ , P1_DATAO_REG_5_ ,
             P1_DATAO_REG_6_ , P1_DATAO_REG_7_ , P1_DATAO_REG_8_ , P1_DATAO_REG_9_ , P1_DATAO_REG_10_ , P1_DATAO_REG_11_ ,
             P1_DATAO_REG_12_ , P1_DATAO_REG_13_ , P1_DATAO_REG_14_ , P1_DATAO_REG_15_ , P1_DATAO_REG_16_ , P1_DATAO_REG_17_ ,
             P1_DATAO_REG_18_ , P1_DATAO_REG_19_ , P1_DATAO_REG_20_ , P1_DATAO_REG_21_ , P1_DATAO_REG_22_ , P1_DATAO_REG_23_ ,
             P1_DATAO_REG_24_ , P1_DATAO_REG_25_ , P1_DATAO_REG_26_ , P1_DATAO_REG_27_ , P1_DATAO_REG_28_ , P1_DATAO_REG_29_ ,
             P1_DATAO_REG_30_ , P1_DATAO_REG_31_ , P1_B_REG , P1_REG3_REG_15_ , P1_REG3_REG_26_ , P1_REG3_REG_6_ ,
             P1_REG3_REG_18_ , P1_REG3_REG_2_ , P1_REG3_REG_11_ , P1_REG3_REG_22_ , P1_REG3_REG_13_ , P1_REG3_REG_20_ ,
             P1_REG3_REG_0_ , P1_REG3_REG_9_ , P1_REG3_REG_4_ , P1_REG3_REG_24_ , P1_REG3_REG_17_ , P1_REG3_REG_5_ ,
             P1_REG3_REG_16_ , P1_REG3_REG_25_ , P1_REG3_REG_12_ , P1_REG3_REG_21_ , P1_REG3_REG_1_ , P1_REG3_REG_8_ ,
             P1_REG3_REG_28_ , P1_REG3_REG_19_ , P1_REG3_REG_3_ , P1_REG3_REG_10_ , P1_REG3_REG_23_ , P1_REG3_REG_14_ ,
             P1_REG3_REG_27_ , P1_REG3_REG_7_ , P1_STATE_REG , P1_RD_REG , P1_WR_REG , P2_IR_REG_0_ ,
             P2_IR_REG_1_ , P2_IR_REG_2_ , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ , P2_IR_REG_6_ ,
             P2_IR_REG_7_ , P2_IR_REG_8_ , P2_IR_REG_9_ , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_ ,
             P2_IR_REG_13_ , P2_IR_REG_14_ , P2_IR_REG_15_ , P2_IR_REG_16_ , P2_IR_REG_17_ , P2_IR_REG_18_ ,
             P2_IR_REG_19_ , P2_IR_REG_20_ , P2_IR_REG_21_ , P2_IR_REG_22_ , P2_IR_REG_23_ , P2_IR_REG_24_ ,
             P2_IR_REG_25_ , P2_IR_REG_26_ , P2_IR_REG_27_ , P2_IR_REG_28_ , P2_IR_REG_29_ , P2_IR_REG_30_ ,
             P2_IR_REG_31_ , P2_D_REG_0_ , P2_D_REG_1_ , P2_D_REG_2_ , P2_D_REG_3_ , P2_D_REG_4_ ,
             P2_D_REG_5_ , P2_D_REG_6_ , P2_D_REG_7_ , P2_D_REG_8_ , P2_D_REG_9_ , P2_D_REG_10_ ,
             P2_D_REG_11_ , P2_D_REG_12_ , P2_D_REG_13_ , P2_D_REG_14_ , P2_D_REG_15_ , P2_D_REG_16_ ,
             P2_D_REG_17_ , P2_D_REG_18_ , P2_D_REG_19_ , P2_D_REG_20_ , P2_D_REG_21_ , P2_D_REG_22_ ,
             P2_D_REG_23_ , P2_D_REG_24_ , P2_D_REG_25_ , P2_D_REG_26_ , P2_D_REG_27_ , P2_D_REG_28_ ,
             P2_D_REG_29_ , P2_D_REG_30_ , P2_D_REG_31_ , P2_REG0_REG_0_ , P2_REG0_REG_1_ , P2_REG0_REG_2_ ,
             P2_REG0_REG_3_ , P2_REG0_REG_4_ , P2_REG0_REG_5_ , P2_REG0_REG_6_ , P2_REG0_REG_7_ , P2_REG0_REG_8_ ,
             P2_REG0_REG_9_ , P2_REG0_REG_10_ , P2_REG0_REG_11_ , P2_REG0_REG_12_ , P2_REG0_REG_13_ , P2_REG0_REG_14_ ,
             P2_REG0_REG_15_ , P2_REG0_REG_16_ , P2_REG0_REG_17_ , P2_REG0_REG_18_ , P2_REG0_REG_19_ , P2_REG0_REG_20_ ,
             P2_REG0_REG_21_ , P2_REG0_REG_22_ , P2_REG0_REG_23_ , P2_REG0_REG_24_ , P2_REG0_REG_25_ , P2_REG0_REG_26_ ,
             P2_REG0_REG_27_ , P2_REG0_REG_28_ , P2_REG0_REG_29_ , P2_REG0_REG_30_ , P2_REG0_REG_31_ , P2_REG1_REG_0_ ,
             P2_REG1_REG_1_ , P2_REG1_REG_2_ , P2_REG1_REG_3_ , P2_REG1_REG_4_ , P2_REG1_REG_5_ , P2_REG1_REG_6_ ,
             P2_REG1_REG_7_ , P2_REG1_REG_8_ , P2_REG1_REG_9_ , P2_REG1_REG_10_ , P2_REG1_REG_11_ , P2_REG1_REG_12_ ,
             P2_REG1_REG_13_ , P2_REG1_REG_14_ , P2_REG1_REG_15_ , P2_REG1_REG_16_ , P2_REG1_REG_17_ , P2_REG1_REG_18_ ,
             P2_REG1_REG_19_ , P2_REG1_REG_20_ , P2_REG1_REG_21_ , P2_REG1_REG_22_ , P2_REG1_REG_23_ , P2_REG1_REG_24_ ,
             P2_REG1_REG_25_ , P2_REG1_REG_26_ , P2_REG1_REG_27_ , P2_REG1_REG_28_ , P2_REG1_REG_29_ , P2_REG1_REG_30_ ,
             P2_REG1_REG_31_ , P2_REG2_REG_0_ , P2_REG2_REG_1_ , P2_REG2_REG_2_ , P2_REG2_REG_3_ , P2_REG2_REG_4_ ,
             P2_REG2_REG_5_ , P2_REG2_REG_6_ , P2_REG2_REG_7_ , P2_REG2_REG_8_ , P2_REG2_REG_9_ , P2_REG2_REG_10_ ,
             P2_REG2_REG_11_ , P2_REG2_REG_12_ , P2_REG2_REG_13_ , P2_REG2_REG_14_ , P2_REG2_REG_15_ , P2_REG2_REG_16_ ,
             P2_REG2_REG_17_ , P2_REG2_REG_18_ , P2_REG2_REG_19_ , P2_REG2_REG_20_ , P2_REG2_REG_21_ , P2_REG2_REG_22_ ,
             P2_REG2_REG_23_ , P2_REG2_REG_24_ , P2_REG2_REG_25_ , P2_REG2_REG_26_ , P2_REG2_REG_27_ , P2_REG2_REG_28_ ,
             P2_REG2_REG_29_ , P2_REG2_REG_30_ , P2_REG2_REG_31_ , P2_ADDR_REG_19_ , P2_ADDR_REG_18_ , P2_ADDR_REG_17_ ,
             P2_ADDR_REG_16_ , P2_ADDR_REG_15_ , P2_ADDR_REG_14_ , P2_ADDR_REG_13_ , P2_ADDR_REG_12_ , P2_ADDR_REG_11_ ,
             P2_ADDR_REG_10_ , P2_ADDR_REG_9_ , P2_ADDR_REG_8_ , P2_ADDR_REG_7_ , P2_ADDR_REG_6_ , P2_ADDR_REG_5_ ,
             P2_ADDR_REG_4_ , P2_ADDR_REG_3_ , P2_ADDR_REG_2_ , P2_ADDR_REG_1_ , P2_ADDR_REG_0_ , P2_DATAO_REG_0_ ,
             P2_DATAO_REG_1_ , P2_DATAO_REG_2_ , P2_DATAO_REG_3_ , P2_DATAO_REG_4_ , P2_DATAO_REG_5_ , P2_DATAO_REG_6_ ,
             P2_DATAO_REG_7_ , P2_DATAO_REG_8_ , P2_DATAO_REG_9_ , P2_DATAO_REG_10_ , P2_DATAO_REG_11_ , P2_DATAO_REG_12_ ,
             P2_DATAO_REG_13_ , P2_DATAO_REG_14_ , P2_DATAO_REG_15_ , P2_DATAO_REG_16_ , P2_DATAO_REG_17_ , P2_DATAO_REG_18_ ,
             P2_DATAO_REG_19_ , P2_DATAO_REG_20_ , P2_DATAO_REG_21_ , P2_DATAO_REG_22_ , P2_DATAO_REG_23_ , P2_DATAO_REG_24_ ,
             P2_DATAO_REG_25_ , P2_DATAO_REG_26_ , P2_DATAO_REG_27_ , P2_DATAO_REG_28_ , P2_DATAO_REG_29_ , P2_DATAO_REG_30_ ,
             P2_DATAO_REG_31_ , P2_B_REG , P2_REG3_REG_15_ , P2_REG3_REG_26_ , P2_REG3_REG_6_ , P2_REG3_REG_18_ ,
             P2_REG3_REG_2_ , P2_REG3_REG_11_ , P2_REG3_REG_22_ , P2_REG3_REG_13_ , P2_REG3_REG_20_ , P2_REG3_REG_0_ ,
             P2_REG3_REG_9_ , P2_REG3_REG_4_ , P2_REG3_REG_24_ , P2_REG3_REG_17_ , P2_REG3_REG_5_ , P2_REG3_REG_16_ ,
             P2_REG3_REG_25_ , P2_REG3_REG_12_ , P2_REG3_REG_21_ , P2_REG3_REG_1_ , P2_REG3_REG_8_ , P2_REG3_REG_28_ ,
             P2_REG3_REG_19_ , P2_REG3_REG_3_ , P2_REG3_REG_10_ , P2_REG3_REG_23_ , P2_REG3_REG_14_ , P2_REG3_REG_27_ ,
             P2_REG3_REG_7_ , P2_STATE_REG , P2_RD_REG , P2_WR_REG , SI_31_ , SI_30_ ,
             SI_29_ , SI_28_ , SI_27_ , SI_26_ , SI_25_ , SI_24_ ,
             SI_23_ , SI_22_ , SI_21_ , SI_20_ , SI_19_ , SI_18_ ,
             SI_17_ , SI_16_ , SI_15_ , SI_14_ , SI_13_ , SI_12_ ,
             SI_11_ , SI_10_ , SI_9_ , SI_8_ , SI_7_ , SI_6_ ,
             SI_5_ , SI_4_ , SI_3_ , SI_2_ , SI_1_ , SI_0_ );

output ADD_1071_U4 , ADD_1071_U55 , ADD_1071_U56 , ADD_1071_U57 , ADD_1071_U58 , ADD_1071_U59;
output ADD_1071_U60 , ADD_1071_U61 , ADD_1071_U62 , ADD_1071_U63 , ADD_1071_U47 , ADD_1071_U48;
output ADD_1071_U49 , ADD_1071_U50 , ADD_1071_U51 , ADD_1071_U52 , ADD_1071_U53 , ADD_1071_U54;
output ADD_1071_U5 , ADD_1071_U46 , U126 , U123;
output P1_U3353 , P1_U3352 , P1_U3351 , P1_U3350 , P1_U3349 , P1_U3348 , P1_U3347;
output P1_U3346 , P1_U3345 , P1_U3344 , P1_U3343 , P1_U3342 , P1_U3341 , P1_U3340;
output P1_U3339 , P1_U3338 , P1_U3337 , P1_U3336 , P1_U3335 , P1_U3334 , P1_U3333;
output P1_U3332 , P1_U3331 , P1_U3330 , P1_U3329 , P1_U3328 , P1_U3327 , P1_U3326;
output P1_U3325 , P1_U3324 , P1_U3323 , P1_U3322 , P1_U3440 , P1_U3441 , P1_U3321;
output P1_U3320 , P1_U3319 , P1_U3318 , P1_U3317 , P1_U3316 , P1_U3315 , P1_U3314;
output P1_U3313 , P1_U3312 , P1_U3311 , P1_U3310 , P1_U3309 , P1_U3308 , P1_U3307;
output P1_U3306 , P1_U3305 , P1_U3304 , P1_U3303 , P1_U3302 , P1_U3301 , P1_U3300;
output P1_U3299 , P1_U3298 , P1_U3297 , P1_U3296 , P1_U3295 , P1_U3294 , P1_U3293;
output P1_U3292 , P1_U3454 , P1_U3457 , P1_U3460 , P1_U3463 , P1_U3466 , P1_U3469;
output P1_U3472 , P1_U3475 , P1_U3478 , P1_U3481 , P1_U3484 , P1_U3487 , P1_U3490;
output P1_U3493 , P1_U3496 , P1_U3499 , P1_U3502 , P1_U3505 , P1_U3508 , P1_U3510;
output P1_U3511 , P1_U3512 , P1_U3513 , P1_U3514 , P1_U3515 , P1_U3516 , P1_U3517;
output P1_U3518 , P1_U3519 , P1_U3520 , P1_U3521 , P1_U3522 , P1_U3523 , P1_U3524;
output P1_U3525 , P1_U3526 , P1_U3527 , P1_U3528 , P1_U3529 , P1_U3530 , P1_U3531;
output P1_U3532 , P1_U3533 , P1_U3534 , P1_U3535 , P1_U3536 , P1_U3537 , P1_U3538;
output P1_U3539 , P1_U3540 , P1_U3541 , P1_U3542 , P1_U3543 , P1_U3544 , P1_U3545;
output P1_U3546 , P1_U3547 , P1_U3548 , P1_U3549 , P1_U3550 , P1_U3551 , P1_U3552;
output P1_U3553 , P1_U3554 , P1_U3291 , P1_U3290 , P1_U3289 , P1_U3288 , P1_U3287;
output P1_U3286 , P1_U3285 , P1_U3284 , P1_U3283 , P1_U3282 , P1_U3281 , P1_U3280;
output P1_U3279 , P1_U3278 , P1_U3277 , P1_U3276 , P1_U3275 , P1_U3274 , P1_U3273;
output P1_U3272 , P1_U3271 , P1_U3270 , P1_U3269 , P1_U3268 , P1_U3267 , P1_U3266;
output P1_U3265 , P1_U3264 , P1_U3263 , P1_U3355 , P1_U3262 , P1_U3261 , P1_U3260;
output P1_U3259 , P1_U3258 , P1_U3257 , P1_U3256 , P1_U3255 , P1_U3254 , P1_U3253;
output P1_U3252 , P1_U3251 , P1_U3250 , P1_U3249 , P1_U3248 , P1_U3247 , P1_U3246;
output P1_U3245 , P1_U3244 , P1_U3243 , P1_U3242 , P1_U3241 , P1_U3555 , P1_U3556;
output P1_U3557 , P1_U3558 , P1_U3559 , P1_U3560 , P1_U3561 , P1_U3562 , P1_U3563;
output P1_U3564 , P1_U3565 , P1_U3566 , P1_U3567 , P1_U3568 , P1_U3569 , P1_U3570;
output P1_U3571 , P1_U3572 , P1_U3573 , P1_U3574 , P1_U3575 , P1_U3576 , P1_U3577;
output P1_U3578 , P1_U3579 , P1_U3580 , P1_U3581 , P1_U3582 , P1_U3583 , P1_U3584;
output P1_U3585 , P1_U3586 , P1_U3240 , P1_U3239 , P1_U3238 , P1_U3237 , P1_U3236;
output P1_U3235 , P1_U3234 , P1_U3233 , P1_U3232 , P1_U3231 , P1_U3230 , P1_U3229;
output P1_U3228 , P1_U3227 , P1_U3226 , P1_U3225 , P1_U3224 , P1_U3223 , P1_U3222;
output P1_U3221 , P1_U3220 , P1_U3219 , P1_U3218 , P1_U3217 , P1_U3216 , P1_U3215;
output P1_U3214 , P1_U3213 , P1_U3212 , P1_U3211 , P1_U3084 , P1_U3083 , P1_U4006;
output P2_U3358 , P2_U3357 , P2_U3356 , P2_U3355 , P2_U3354 , P2_U3353 , P2_U3352;
output P2_U3351 , P2_U3350 , P2_U3349 , P2_U3348 , P2_U3347 , P2_U3346 , P2_U3345;
output P2_U3344 , P2_U3343 , P2_U3342 , P2_U3341 , P2_U3340 , P2_U3339 , P2_U3338;
output P2_U3337 , P2_U3336 , P2_U3335 , P2_U3334 , P2_U3333 , P2_U3332 , P2_U3331;
output P2_U3330 , P2_U3329 , P2_U3328 , P2_U3327 , P2_U3437 , P2_U3438 , P2_U3326;
output P2_U3325 , P2_U3324 , P2_U3323 , P2_U3322 , P2_U3321 , P2_U3320 , P2_U3319;
output P2_U3318 , P2_U3317 , P2_U3316 , P2_U3315 , P2_U3314 , P2_U3313 , P2_U3312;
output P2_U3311 , P2_U3310 , P2_U3309 , P2_U3308 , P2_U3307 , P2_U3306 , P2_U3305;
output P2_U3304 , P2_U3303 , P2_U3302 , P2_U3301 , P2_U3300 , P2_U3299 , P2_U3298;
output P2_U3297 , P2_U3451 , P2_U3454 , P2_U3457 , P2_U3460 , P2_U3463 , P2_U3466;
output P2_U3469 , P2_U3472 , P2_U3475 , P2_U3478 , P2_U3481 , P2_U3484 , P2_U3487;
output P2_U3490 , P2_U3493 , P2_U3496 , P2_U3499 , P2_U3502 , P2_U3505 , P2_U3507;
output P2_U3508 , P2_U3509 , P2_U3510 , P2_U3511 , P2_U3512 , P2_U3513 , P2_U3514;
output P2_U3515 , P2_U3516 , P2_U3517 , P2_U3518 , P2_U3519 , P2_U3520 , P2_U3521;
output P2_U3522 , P2_U3523 , P2_U3524 , P2_U3525 , P2_U3526 , P2_U3527 , P2_U3528;
output P2_U3529 , P2_U3530 , P2_U3531 , P2_U3532 , P2_U3533 , P2_U3534 , P2_U3535;
output P2_U3536 , P2_U3537 , P2_U3538 , P2_U3539 , P2_U3540 , P2_U3541 , P2_U3542;
output P2_U3543 , P2_U3544 , P2_U3545 , P2_U3546 , P2_U3547 , P2_U3548 , P2_U3549;
output P2_U3550 , P2_U3551 , P2_U3296 , P2_U3295 , P2_U3294 , P2_U3293 , P2_U3292;
output P2_U3291 , P2_U3290 , P2_U3289 , P2_U3288 , P2_U3287 , P2_U3286 , P2_U3285;
output P2_U3284 , P2_U3283 , P2_U3282 , P2_U3281 , P2_U3280 , P2_U3279 , P2_U3278;
output P2_U3277 , P2_U3276 , P2_U3275 , P2_U3274 , P2_U3273 , P2_U3272 , P2_U3271;
output P2_U3270 , P2_U3269 , P2_U3268 , P2_U3267 , P2_U3266 , P2_U3265 , P2_U3264;
output P2_U3263 , P2_U3262 , P2_U3261 , P2_U3260 , P2_U3259 , P2_U3258 , P2_U3257;
output P2_U3256 , P2_U3255 , P2_U3254 , P2_U3253 , P2_U3252 , P2_U3251 , P2_U3250;
output P2_U3249 , P2_U3248 , P2_U3247 , P2_U3246 , P2_U3245 , P2_U3552 , P2_U3553;
output P2_U3554 , P2_U3555 , P2_U3556 , P2_U3557 , P2_U3558 , P2_U3559 , P2_U3560;
output P2_U3561 , P2_U3562 , P2_U3563 , P2_U3564 , P2_U3565 , P2_U3566 , P2_U3567;
output P2_U3568 , P2_U3569 , P2_U3570 , P2_U3571 , P2_U3572 , P2_U3573 , P2_U3574;
output P2_U3575 , P2_U3576 , P2_U3577 , P2_U3578 , P2_U3579 , P2_U3580 , P2_U3581;
output P2_U3582 , P2_U3583 , P2_U3244 , P2_U3243 , P2_U3242 , P2_U3241 , P2_U3240;
output P2_U3239 , P2_U3238 , P2_U3237 , P2_U3236 , P2_U3235 , P2_U3234 , P2_U3233;
output P2_U3232 , P2_U3231 , P2_U3230 , P2_U3229 , P2_U3228 , P2_U3227 , P2_U3226;
output P2_U3225 , P2_U3224 , P2_U3223 , P2_U3222 , P2_U3221 , P2_U3220 , P2_U3219;
output P2_U3218 , P2_U3217 , P2_U3216 , P2_U3215 , P2_U3152 , P2_U3151 , P2_U3966;

input SI_31_ , SI_30_ , SI_29_ , SI_28_ , SI_27_ , SI_26_;
input SI_25_ , SI_24_ , SI_23_ , SI_22_ , SI_21_ , SI_20_;
input SI_19_ , SI_18_ , SI_17_ , SI_16_ , SI_15_ , SI_14_;
input SI_13_ , SI_12_ , SI_11_ , SI_10_ , SI_9_ , SI_8_;
input SI_7_ , SI_6_ , SI_5_ , SI_4_ , SI_3_ , SI_2_;
input SI_1_ , SI_0_;
input P1_IR_REG_0_ , P1_IR_REG_1_ , P1_IR_REG_2_ , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_;
input P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_10_ , P1_IR_REG_11_;
input P1_IR_REG_12_ , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_;
input P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_20_ , P1_IR_REG_21_ , P1_IR_REG_22_ , P1_IR_REG_23_;
input P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ , P1_IR_REG_27_ , P1_IR_REG_28_ , P1_IR_REG_29_;
input P1_IR_REG_30_ , P1_IR_REG_31_ , P1_D_REG_0_ , P1_D_REG_1_ , P1_D_REG_2_ , P1_D_REG_3_;
input P1_D_REG_4_ , P1_D_REG_5_ , P1_D_REG_6_ , P1_D_REG_7_ , P1_D_REG_8_ , P1_D_REG_9_;
input P1_D_REG_10_ , P1_D_REG_11_ , P1_D_REG_12_ , P1_D_REG_13_ , P1_D_REG_14_ , P1_D_REG_15_;
input P1_D_REG_16_ , P1_D_REG_17_ , P1_D_REG_18_ , P1_D_REG_19_ , P1_D_REG_20_ , P1_D_REG_21_;
input P1_D_REG_22_ , P1_D_REG_23_ , P1_D_REG_24_ , P1_D_REG_25_ , P1_D_REG_26_ , P1_D_REG_27_;
input P1_D_REG_28_ , P1_D_REG_29_ , P1_D_REG_30_ , P1_D_REG_31_ , P1_REG0_REG_0_ , P1_REG0_REG_1_;
input P1_REG0_REG_2_ , P1_REG0_REG_3_ , P1_REG0_REG_4_ , P1_REG0_REG_5_ , P1_REG0_REG_6_ , P1_REG0_REG_7_;
input P1_REG0_REG_8_ , P1_REG0_REG_9_ , P1_REG0_REG_10_ , P1_REG0_REG_11_ , P1_REG0_REG_12_ , P1_REG0_REG_13_;
input P1_REG0_REG_14_ , P1_REG0_REG_15_ , P1_REG0_REG_16_ , P1_REG0_REG_17_ , P1_REG0_REG_18_ , P1_REG0_REG_19_;
input P1_REG0_REG_20_ , P1_REG0_REG_21_ , P1_REG0_REG_22_ , P1_REG0_REG_23_ , P1_REG0_REG_24_ , P1_REG0_REG_25_;
input P1_REG0_REG_26_ , P1_REG0_REG_27_ , P1_REG0_REG_28_ , P1_REG0_REG_29_ , P1_REG0_REG_30_ , P1_REG0_REG_31_;
input P1_REG1_REG_0_ , P1_REG1_REG_1_ , P1_REG1_REG_2_ , P1_REG1_REG_3_ , P1_REG1_REG_4_ , P1_REG1_REG_5_;
input P1_REG1_REG_6_ , P1_REG1_REG_7_ , P1_REG1_REG_8_ , P1_REG1_REG_9_ , P1_REG1_REG_10_ , P1_REG1_REG_11_;
input P1_REG1_REG_12_ , P1_REG1_REG_13_ , P1_REG1_REG_14_ , P1_REG1_REG_15_ , P1_REG1_REG_16_ , P1_REG1_REG_17_;
input P1_REG1_REG_18_ , P1_REG1_REG_19_ , P1_REG1_REG_20_ , P1_REG1_REG_21_ , P1_REG1_REG_22_ , P1_REG1_REG_23_;
input P1_REG1_REG_24_ , P1_REG1_REG_25_ , P1_REG1_REG_26_ , P1_REG1_REG_27_ , P1_REG1_REG_28_ , P1_REG1_REG_29_;
input P1_REG1_REG_30_ , P1_REG1_REG_31_ , P1_REG2_REG_0_ , P1_REG2_REG_1_ , P1_REG2_REG_2_ , P1_REG2_REG_3_;
input P1_REG2_REG_4_ , P1_REG2_REG_5_ , P1_REG2_REG_6_ , P1_REG2_REG_7_ , P1_REG2_REG_8_ , P1_REG2_REG_9_;
input P1_REG2_REG_10_ , P1_REG2_REG_11_ , P1_REG2_REG_12_ , P1_REG2_REG_13_ , P1_REG2_REG_14_ , P1_REG2_REG_15_;
input P1_REG2_REG_16_ , P1_REG2_REG_17_ , P1_REG2_REG_18_ , P1_REG2_REG_19_ , P1_REG2_REG_20_ , P1_REG2_REG_21_;
input P1_REG2_REG_22_ , P1_REG2_REG_23_ , P1_REG2_REG_24_ , P1_REG2_REG_25_ , P1_REG2_REG_26_ , P1_REG2_REG_27_;
input P1_REG2_REG_28_ , P1_REG2_REG_29_ , P1_REG2_REG_30_ , P1_REG2_REG_31_ , P1_ADDR_REG_19_ , P1_ADDR_REG_18_;
input P1_ADDR_REG_17_ , P1_ADDR_REG_16_ , P1_ADDR_REG_15_ , P1_ADDR_REG_14_ , P1_ADDR_REG_13_ , P1_ADDR_REG_12_;
input P1_ADDR_REG_11_ , P1_ADDR_REG_10_ , P1_ADDR_REG_9_ , P1_ADDR_REG_8_ , P1_ADDR_REG_7_ , P1_ADDR_REG_6_;
input P1_ADDR_REG_5_ , P1_ADDR_REG_4_ , P1_ADDR_REG_3_ , P1_ADDR_REG_2_ , P1_ADDR_REG_1_ , P1_ADDR_REG_0_;
input P1_DATAO_REG_0_ , P1_DATAO_REG_1_ , P1_DATAO_REG_2_ , P1_DATAO_REG_3_ , P1_DATAO_REG_4_ , P1_DATAO_REG_5_;
input P1_DATAO_REG_6_ , P1_DATAO_REG_7_ , P1_DATAO_REG_8_ , P1_DATAO_REG_9_ , P1_DATAO_REG_10_ , P1_DATAO_REG_11_;
input P1_DATAO_REG_12_ , P1_DATAO_REG_13_ , P1_DATAO_REG_14_ , P1_DATAO_REG_15_ , P1_DATAO_REG_16_ , P1_DATAO_REG_17_;
input P1_DATAO_REG_18_ , P1_DATAO_REG_19_ , P1_DATAO_REG_20_ , P1_DATAO_REG_21_ , P1_DATAO_REG_22_ , P1_DATAO_REG_23_;
input P1_DATAO_REG_24_ , P1_DATAO_REG_25_ , P1_DATAO_REG_26_ , P1_DATAO_REG_27_ , P1_DATAO_REG_28_ , P1_DATAO_REG_29_;
input P1_DATAO_REG_30_ , P1_DATAO_REG_31_ , P1_B_REG , P1_REG3_REG_15_ , P1_REG3_REG_26_ , P1_REG3_REG_6_;
input P1_REG3_REG_18_ , P1_REG3_REG_2_ , P1_REG3_REG_11_ , P1_REG3_REG_22_ , P1_REG3_REG_13_ , P1_REG3_REG_20_;
input P1_REG3_REG_0_ , P1_REG3_REG_9_ , P1_REG3_REG_4_ , P1_REG3_REG_24_ , P1_REG3_REG_17_ , P1_REG3_REG_5_;
input P1_REG3_REG_16_ , P1_REG3_REG_25_ , P1_REG3_REG_12_ , P1_REG3_REG_21_ , P1_REG3_REG_1_ , P1_REG3_REG_8_;
input P1_REG3_REG_28_ , P1_REG3_REG_19_ , P1_REG3_REG_3_ , P1_REG3_REG_10_ , P1_REG3_REG_23_ , P1_REG3_REG_14_;
input P1_REG3_REG_27_ , P1_REG3_REG_7_ , P1_STATE_REG , P1_RD_REG , P1_WR_REG , P2_IR_REG_0_;
input P2_IR_REG_1_ , P2_IR_REG_2_ , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ , P2_IR_REG_6_;
input P2_IR_REG_7_ , P2_IR_REG_8_ , P2_IR_REG_9_ , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_;
input P2_IR_REG_13_ , P2_IR_REG_14_ , P2_IR_REG_15_ , P2_IR_REG_16_ , P2_IR_REG_17_ , P2_IR_REG_18_;
input P2_IR_REG_19_ , P2_IR_REG_20_ , P2_IR_REG_21_ , P2_IR_REG_22_ , P2_IR_REG_23_ , P2_IR_REG_24_;
input P2_IR_REG_25_ , P2_IR_REG_26_ , P2_IR_REG_27_ , P2_IR_REG_28_ , P2_IR_REG_29_ , P2_IR_REG_30_;
input P2_IR_REG_31_ , P2_D_REG_0_ , P2_D_REG_1_ , P2_D_REG_2_ , P2_D_REG_3_ , P2_D_REG_4_;
input P2_D_REG_5_ , P2_D_REG_6_ , P2_D_REG_7_ , P2_D_REG_8_ , P2_D_REG_9_ , P2_D_REG_10_;
input P2_D_REG_11_ , P2_D_REG_12_ , P2_D_REG_13_ , P2_D_REG_14_ , P2_D_REG_15_ , P2_D_REG_16_;
input P2_D_REG_17_ , P2_D_REG_18_ , P2_D_REG_19_ , P2_D_REG_20_ , P2_D_REG_21_ , P2_D_REG_22_;
input P2_D_REG_23_ , P2_D_REG_24_ , P2_D_REG_25_ , P2_D_REG_26_ , P2_D_REG_27_ , P2_D_REG_28_;
input P2_D_REG_29_ , P2_D_REG_30_ , P2_D_REG_31_ , P2_REG0_REG_0_ , P2_REG0_REG_1_ , P2_REG0_REG_2_;
input P2_REG0_REG_3_ , P2_REG0_REG_4_ , P2_REG0_REG_5_ , P2_REG0_REG_6_ , P2_REG0_REG_7_ , P2_REG0_REG_8_;
input P2_REG0_REG_9_ , P2_REG0_REG_10_ , P2_REG0_REG_11_ , P2_REG0_REG_12_ , P2_REG0_REG_13_ , P2_REG0_REG_14_;
input P2_REG0_REG_15_ , P2_REG0_REG_16_ , P2_REG0_REG_17_ , P2_REG0_REG_18_ , P2_REG0_REG_19_ , P2_REG0_REG_20_;
input P2_REG0_REG_21_ , P2_REG0_REG_22_ , P2_REG0_REG_23_ , P2_REG0_REG_24_ , P2_REG0_REG_25_ , P2_REG0_REG_26_;
input P2_REG0_REG_27_ , P2_REG0_REG_28_ , P2_REG0_REG_29_ , P2_REG0_REG_30_ , P2_REG0_REG_31_ , P2_REG1_REG_0_;
input P2_REG1_REG_1_ , P2_REG1_REG_2_ , P2_REG1_REG_3_ , P2_REG1_REG_4_ , P2_REG1_REG_5_ , P2_REG1_REG_6_;
input P2_REG1_REG_7_ , P2_REG1_REG_8_ , P2_REG1_REG_9_ , P2_REG1_REG_10_ , P2_REG1_REG_11_ , P2_REG1_REG_12_;
input P2_REG1_REG_13_ , P2_REG1_REG_14_ , P2_REG1_REG_15_ , P2_REG1_REG_16_ , P2_REG1_REG_17_ , P2_REG1_REG_18_;
input P2_REG1_REG_19_ , P2_REG1_REG_20_ , P2_REG1_REG_21_ , P2_REG1_REG_22_ , P2_REG1_REG_23_ , P2_REG1_REG_24_;
input P2_REG1_REG_25_ , P2_REG1_REG_26_ , P2_REG1_REG_27_ , P2_REG1_REG_28_ , P2_REG1_REG_29_ , P2_REG1_REG_30_;
input P2_REG1_REG_31_ , P2_REG2_REG_0_ , P2_REG2_REG_1_ , P2_REG2_REG_2_ , P2_REG2_REG_3_ , P2_REG2_REG_4_;
input P2_REG2_REG_5_ , P2_REG2_REG_6_ , P2_REG2_REG_7_ , P2_REG2_REG_8_ , P2_REG2_REG_9_ , P2_REG2_REG_10_;
input P2_REG2_REG_11_ , P2_REG2_REG_12_ , P2_REG2_REG_13_ , P2_REG2_REG_14_ , P2_REG2_REG_15_ , P2_REG2_REG_16_;
input P2_REG2_REG_17_ , P2_REG2_REG_18_ , P2_REG2_REG_19_ , P2_REG2_REG_20_ , P2_REG2_REG_21_ , P2_REG2_REG_22_;
input P2_REG2_REG_23_ , P2_REG2_REG_24_ , P2_REG2_REG_25_ , P2_REG2_REG_26_ , P2_REG2_REG_27_ , P2_REG2_REG_28_;
input P2_REG2_REG_29_ , P2_REG2_REG_30_ , P2_REG2_REG_31_ , P2_ADDR_REG_19_ , P2_ADDR_REG_18_ , P2_ADDR_REG_17_;
input P2_ADDR_REG_16_ , P2_ADDR_REG_15_ , P2_ADDR_REG_14_ , P2_ADDR_REG_13_ , P2_ADDR_REG_12_ , P2_ADDR_REG_11_;
input P2_ADDR_REG_10_ , P2_ADDR_REG_9_ , P2_ADDR_REG_8_ , P2_ADDR_REG_7_ , P2_ADDR_REG_6_ , P2_ADDR_REG_5_;
input P2_ADDR_REG_4_ , P2_ADDR_REG_3_ , P2_ADDR_REG_2_ , P2_ADDR_REG_1_ , P2_ADDR_REG_0_ , P2_DATAO_REG_0_;
input P2_DATAO_REG_1_ , P2_DATAO_REG_2_ , P2_DATAO_REG_3_ , P2_DATAO_REG_4_ , P2_DATAO_REG_5_ , P2_DATAO_REG_6_;
input P2_DATAO_REG_7_ , P2_DATAO_REG_8_ , P2_DATAO_REG_9_ , P2_DATAO_REG_10_ , P2_DATAO_REG_11_ , P2_DATAO_REG_12_;
input P2_DATAO_REG_13_ , P2_DATAO_REG_14_ , P2_DATAO_REG_15_ , P2_DATAO_REG_16_ , P2_DATAO_REG_17_ , P2_DATAO_REG_18_;
input P2_DATAO_REG_19_ , P2_DATAO_REG_20_ , P2_DATAO_REG_21_ , P2_DATAO_REG_22_ , P2_DATAO_REG_23_ , P2_DATAO_REG_24_;
input P2_DATAO_REG_25_ , P2_DATAO_REG_26_ , P2_DATAO_REG_27_ , P2_DATAO_REG_28_ , P2_DATAO_REG_29_ , P2_DATAO_REG_30_;
input P2_DATAO_REG_31_ , P2_B_REG , P2_REG3_REG_15_ , P2_REG3_REG_26_ , P2_REG3_REG_6_ , P2_REG3_REG_18_;
input P2_REG3_REG_2_ , P2_REG3_REG_11_ , P2_REG3_REG_22_ , P2_REG3_REG_13_ , P2_REG3_REG_20_ , P2_REG3_REG_0_;
input P2_REG3_REG_9_ , P2_REG3_REG_4_ , P2_REG3_REG_24_ , P2_REG3_REG_17_ , P2_REG3_REG_5_ , P2_REG3_REG_16_;
input P2_REG3_REG_25_ , P2_REG3_REG_12_ , P2_REG3_REG_21_ , P2_REG3_REG_1_ , P2_REG3_REG_8_ , P2_REG3_REG_28_;
input P2_REG3_REG_19_ , P2_REG3_REG_3_ , P2_REG3_REG_10_ , P2_REG3_REG_23_ , P2_REG3_REG_14_ , P2_REG3_REG_27_;
input P2_REG3_REG_7_ , P2_STATE_REG , P2_RD_REG , P2_WR_REG;

wire P2_R1113_U477 , P2_R1113_U476 , P2_R1113_U475 , U25 , U26 , U27 , U28 , U29 , U30 , U31;
wire U32 , U33 , U34 , U35 , U36 , U37 , U38 , U39 , U40 , U41;
wire U42 , U43 , U44 , U45 , U46 , U47 , U48 , U49 , U50 , U51;
wire U52 , U53 , U54 , U55 , U56 , U57 , U58 , U59 , U60 , U61;
wire U62 , U63 , U64 , U65 , U66 , U67 , U68 , U69 , U70 , U71;
wire U72 , U73 , U74 , U75 , U76 , U77 , U78 , U79 , U80 , U81;
wire U82 , U83 , U84 , U85 , U86 , U87 , U88 , U89 , U90 , U91;
wire U92 , U93 , U94 , U95 , U96 , U97 , U98 , U99 , U100 , U101;
wire U102 , U103 , U104 , U105 , U106 , U107 , U108 , U109 , U110 , U111;
wire U112 , U113 , U114 , U115 , U116 , U117 , U118 , U119 , U120 , U121;
wire U122 , U124 , U125 , U127 , U128 , U129 , U130 , U131 , U132 , U133;
wire U134 , U135 , U136 , U137 , U138 , U139 , U140 , U141 , U142 , U143;
wire U144 , U145 , U146 , U147 , U148 , U149 , U150 , U151 , U152 , U153;
wire U154 , U155 , U156 , U157 , U158 , U159 , U160 , U161 , U162 , U163;
wire U164 , U165 , U166 , U167 , U168 , U169 , U170 , U171 , U172 , U173;
wire U174 , U175 , U176 , U177 , U178 , U179 , U180 , U181 , U182 , U183;
wire U184 , U185 , U186 , U187 , U188 , U189 , U190 , U191 , U192 , U193;
wire U194 , U195 , U196 , U197 , U198 , U199 , U200 , U201 , U202 , U203;
wire U204 , U205 , U206 , U207 , U208 , U209 , U210 , U211 , U212 , U213;
wire U214 , U215 , U216 , U217 , U218 , U219 , U220 , U221 , U222 , U223;
wire U224 , U225 , U226 , U227 , U228 , U229 , U230 , U231 , U232 , U233;
wire U234 , U235 , U236 , U237 , U238 , U239 , U240 , U241 , U242 , U243;
wire U244 , U245 , U246 , U247 , U248 , U249 , U250 , U251 , U252 , U253;
wire U254 , U255 , U256 , U257 , U258 , U259 , U260 , U261 , U262 , U263;
wire U264 , U265 , U266 , U267 , U268 , U269 , U270 , U271 , U272 , U273;
wire U274 , U275 , U276 , U277 , U278 , U279 , U280 , U281 , U282 , U283;
wire U284 , U285 , U286 , U287 , U288 , U289 , U290 , U291 , U292 , U293;
wire U294 , U295 , U296 , U297 , U298 , U299 , U300 , U301 , U302 , U303;
wire U304 , U305 , U306 , U307 , U308 , U309 , U310 , U311 , U312 , U313;
wire U314 , U315 , U316 , U317 , U318 , U319 , U320 , U321 , U322 , U323;
wire U324 , U325 , U326 , P2_R1113_U474 , P2_R1113_U473 , P2_R1113_U472 , P2_R1113_U471 , P2_R1113_U470 , P2_R1113_U469 , P2_R1113_U468;
wire P2_R1113_U467 , P2_R1113_U466 , P2_R1113_U465 , P2_R1113_U464 , P2_R1113_U463 , P1_U3014 , P1_U3015 , P1_U3016 , P1_U3017 , P1_U3018;
wire P1_U3019 , P1_U3020 , P1_U3021 , P1_U3022 , P1_U3023 , P1_U3024 , P1_U3025 , P1_U3026 , P1_U3027 , P1_U3028;
wire P1_U3029 , P1_U3030 , P1_U3031 , P1_U3032 , P1_U3033 , P1_U3034 , P1_U3035 , P1_U3036 , P1_U3037 , P1_U3038;
wire P1_U3039 , P1_U3040 , P1_U3041 , P1_U3042 , P1_U3043 , P1_U3044 , P1_U3045 , P1_U3046 , P1_U3047 , P1_U3048;
wire P1_U3049 , P1_U3050 , P1_U3051 , P1_U3052 , P1_U3053 , P1_U3054 , P1_U3055 , P1_U3056 , P1_U3057 , P1_U3058;
wire P1_U3059 , P1_U3060 , P1_U3061 , P1_U3062 , P1_U3063 , P1_U3064 , P1_U3065 , P1_U3066 , P1_U3067 , P1_U3068;
wire P1_U3069 , P1_U3070 , P1_U3071 , P1_U3072 , P1_U3073 , P1_U3074 , P1_U3075 , P1_U3076 , P1_U3077 , P1_U3078;
wire P1_U3079 , P1_U3080 , P1_U3081 , P1_U3082 , P1_U3085 , P1_U3086 , P1_U3087 , P1_U3088 , P1_U3089 , P1_U3090;
wire P1_U3091 , P1_U3092 , P1_U3093 , P1_U3094 , P1_U3095 , P1_U3096 , P1_U3097 , P1_U3098 , P1_U3099 , P1_U3100;
wire P1_U3101 , P1_U3102 , P1_U3103 , P1_U3104 , P1_U3105 , P1_U3106 , P1_U3107 , P1_U3108 , P1_U3109 , P1_U3110;
wire P1_U3111 , P1_U3112 , P1_U3113 , P1_U3114 , P1_U3115 , P1_U3116 , P1_U3117 , P1_U3118 , P1_U3119 , P1_U3120;
wire P1_U3121 , P1_U3122 , P1_U3123 , P1_U3124 , P1_U3125 , P1_U3126 , P1_U3127 , P1_U3128 , P1_U3129 , P1_U3130;
wire P1_U3131 , P1_U3132 , P1_U3133 , P1_U3134 , P1_U3135 , P1_U3136 , P1_U3137 , P1_U3138 , P1_U3139 , P1_U3140;
wire P1_U3141 , P1_U3142 , P1_U3143 , P1_U3144 , P1_U3145 , P1_U3146 , P1_U3147 , P1_U3148 , P1_U3149 , P1_U3150;
wire P1_U3151 , P1_U3152 , P1_U3153 , P1_U3154 , P1_U3155 , P1_U3156 , P1_U3157 , P1_U3158 , P1_U3159 , P1_U3160;
wire P1_U3161 , P1_U3162 , P1_U3163 , P1_U3164 , P1_U3165 , P1_U3166 , P1_U3167 , P1_U3168 , P1_U3169 , P1_U3170;
wire P1_U3171 , P1_U3172 , P1_U3173 , P1_U3174 , P1_U3175 , P1_U3176 , P1_U3177 , P1_U3178 , P1_U3179 , P1_U3180;
wire P1_U3181 , P1_U3182 , P1_U3183 , P1_U3184 , P1_U3185 , P1_U3186 , P1_U3187 , P1_U3188 , P1_U3189 , P1_U3190;
wire P1_U3191 , P1_U3192 , P1_U3193 , P1_U3194 , P1_U3195 , P1_U3196 , P1_U3197 , P1_U3198 , P1_U3199 , P1_U3200;
wire P1_U3201 , P1_U3202 , P1_U3203 , P1_U3204 , P1_U3205 , P1_U3206 , P1_U3207 , P1_U3208 , P1_U3209 , P1_U3210;
wire P1_U3354 , P1_U3356 , P1_U3357 , P1_U3358 , P1_U3359 , P1_U3360 , P1_U3361 , P1_U3362 , P1_U3363 , P1_U3364;
wire P1_U3365 , P1_U3366 , P1_U3367 , P1_U3368 , P1_U3369 , P1_U3370 , P1_U3371 , P1_U3372 , P1_U3373 , P1_U3374;
wire P1_U3375 , P1_U3376 , P1_U3377 , P1_U3378 , P1_U3379 , P1_U3380 , P1_U3381 , P1_U3382 , P1_U3383 , P1_U3384;
wire P1_U3385 , P1_U3386 , P1_U3387 , P1_U3388 , P1_U3389 , P1_U3390 , P1_U3391 , P1_U3392 , P1_U3393 , P1_U3394;
wire P1_U3395 , P1_U3396 , P1_U3397 , P1_U3398 , P1_U3399 , P1_U3400 , P1_U3401 , P1_U3402 , P1_U3403 , P1_U3404;
wire P1_U3405 , P1_U3406 , P1_U3407 , P1_U3408 , P1_U3409 , P1_U3410 , P1_U3411 , P1_U3412 , P1_U3413 , P1_U3414;
wire P1_U3415 , P1_U3416 , P1_U3417 , P1_U3418 , P1_U3419 , P1_U3420 , P1_U3421 , P1_U3422 , P1_U3423 , P1_U3424;
wire P1_U3425 , P1_U3426 , P1_U3427 , P1_U3428 , P1_U3429 , P1_U3430 , P1_U3431 , P1_U3432 , P1_U3433 , P1_U3434;
wire P1_U3435 , P1_U3436 , P1_U3437 , P1_U3438 , P1_U3439 , P1_U3442 , P1_U3443 , P1_U3444 , P1_U3445 , P1_U3446;
wire P1_U3447 , P1_U3448 , P1_U3449 , P1_U3450 , P1_U3451 , P1_U3452 , P1_U3453 , P1_U3455 , P1_U3456 , P1_U3458;
wire P1_U3459 , P1_U3461 , P1_U3462 , P1_U3464 , P1_U3465 , P1_U3467 , P1_U3468 , P1_U3470 , P1_U3471 , P1_U3473;
wire P1_U3474 , P1_U3476 , P1_U3477 , P1_U3479 , P1_U3480 , P1_U3482 , P1_U3483 , P1_U3485 , P1_U3486 , P1_U3488;
wire P1_U3489 , P1_U3491 , P1_U3492 , P1_U3494 , P1_U3495 , P1_U3497 , P1_U3498 , P1_U3500 , P1_U3501 , P1_U3503;
wire P1_U3504 , P1_U3506 , P1_U3507 , P1_U3509 , P1_U3587 , P1_U3588 , P1_U3589 , P1_U3590 , P1_U3591 , P1_U3592;
wire P1_U3593 , P1_U3594 , P1_U3595 , P1_U3596 , P1_U3597 , P1_U3598 , P1_U3599 , P1_U3600 , P1_U3601 , P1_U3602;
wire P1_U3603 , P1_U3604 , P1_U3605 , P1_U3606 , P1_U3607 , P1_U3608 , P1_U3609 , P1_U3610 , P1_U3611 , P1_U3612;
wire P1_U3613 , P1_U3614 , P1_U3615 , P1_U3616 , P1_U3617 , P1_U3618 , P1_U3619 , P1_U3620 , P1_U3621 , P1_U3622;
wire P1_U3623 , P1_U3624 , P1_U3625 , P1_U3626 , P1_U3627 , P1_U3628 , P1_U3629 , P1_U3630 , P1_U3631 , P1_U3632;
wire P1_U3633 , P1_U3634 , P1_U3635 , P1_U3636 , P1_U3637 , P1_U3638 , P1_U3639 , P1_U3640 , P1_U3641 , P1_U3642;
wire P1_U3643 , P1_U3644 , P1_U3645 , P1_U3646 , P1_U3647 , P1_U3648 , P1_U3649 , P1_U3650 , P1_U3651 , P1_U3652;
wire P1_U3653 , P1_U3654 , P1_U3655 , P1_U3656 , P1_U3657 , P1_U3658 , P1_U3659 , P1_U3660 , P1_U3661 , P1_U3662;
wire P1_U3663 , P1_U3664 , P1_U3665 , P1_U3666 , P1_U3667 , P1_U3668 , P1_U3669 , P1_U3670 , P1_U3671 , P1_U3672;
wire P1_U3673 , P1_U3674 , P1_U3675 , P1_U3676 , P1_U3677 , P1_U3678 , P1_U3679 , P1_U3680 , P1_U3681 , P1_U3682;
wire P1_U3683 , P1_U3684 , P1_U3685 , P1_U3686 , P1_U3687 , P1_U3688 , P1_U3689 , P1_U3690 , P1_U3691 , P1_U3692;
wire P1_U3693 , P1_U3694 , P1_U3695 , P1_U3696 , P1_U3697 , P1_U3698 , P1_U3699 , P1_U3700 , P1_U3701 , P1_U3702;
wire P1_U3703 , P1_U3704 , P1_U3705 , P1_U3706 , P1_U3707 , P1_U3708 , P1_U3709 , P1_U3710 , P1_U3711 , P1_U3712;
wire P1_U3713 , P1_U3714 , P1_U3715 , P1_U3716 , P1_U3717 , P1_U3718 , P1_U3719 , P1_U3720 , P1_U3721 , P1_U3722;
wire P1_U3723 , P1_U3724 , P1_U3725 , P1_U3726 , P1_U3727 , P1_U3728 , P1_U3729 , P1_U3730 , P1_U3731 , P1_U3732;
wire P1_U3733 , P1_U3734 , P1_U3735 , P1_U3736 , P1_U3737 , P1_U3738 , P1_U3739 , P1_U3740 , P1_U3741 , P1_U3742;
wire P1_U3743 , P1_U3744 , P1_U3745 , P1_U3746 , P1_U3747 , P1_U3748 , P1_U3749 , P1_U3750 , P1_U3751 , P1_U3752;
wire P1_U3753 , P1_U3754 , P1_U3755 , P1_U3756 , P1_U3757 , P1_U3758 , P1_U3759 , P1_U3760 , P1_U3761 , P1_U3762;
wire P1_U3763 , P1_U3764 , P1_U3765 , P1_U3766 , P1_U3767 , P1_U3768 , P1_U3769 , P1_U3770 , P1_U3771 , P1_U3772;
wire P1_U3773 , P1_U3774 , P1_U3775 , P1_U3776 , P1_U3777 , P1_U3778 , P1_U3779 , P1_U3780 , P1_U3781 , P1_U3782;
wire P1_U3783 , P1_U3784 , P1_U3785 , P1_U3786 , P1_U3787 , P1_U3788 , P1_U3789 , P1_U3790 , P1_U3791 , P1_U3792;
wire P1_U3793 , P1_U3794 , P1_U3795 , P1_U3796 , P1_U3797 , P1_U3798 , P1_U3799 , P1_U3800 , P1_U3801 , P1_U3802;
wire P1_U3803 , P1_U3804 , P1_U3805 , P1_U3806 , P1_U3807 , P1_U3808 , P1_U3809 , P1_U3810 , P1_U3811 , P1_U3812;
wire P1_U3813 , P1_U3814 , P1_U3815 , P1_U3816 , P1_U3817 , P1_U3818 , P1_U3819 , P1_U3820 , P1_U3821 , P1_U3822;
wire P1_U3823 , P1_U3824 , P1_U3825 , P1_U3826 , P1_U3827 , P1_U3828 , P1_U3829 , P1_U3830 , P1_U3831 , P1_U3832;
wire P1_U3833 , P1_U3834 , P1_U3835 , P1_U3836 , P1_U3837 , P1_U3838 , P1_U3839 , P1_U3840 , P1_U3841 , P1_U3842;
wire P1_U3843 , P1_U3844 , P1_U3845 , P1_U3846 , P1_U3847 , P1_U3848 , P1_U3849 , P1_U3850 , P1_U3851 , P1_U3852;
wire P1_U3853 , P1_U3854 , P1_U3855 , P1_U3856 , P1_U3857 , P1_U3858 , P1_U3859 , P1_U3860 , P1_U3861 , P1_U3862;
wire P1_U3863 , P1_U3864 , P1_U3865 , P1_U3866 , P1_U3867 , P1_U3868 , P1_U3869 , P1_U3870 , P1_U3871 , P1_U3872;
wire P1_U3873 , P1_U3874 , P1_U3875 , P1_U3876 , P1_U3877 , P1_U3878 , P1_U3879 , P1_U3880 , P1_U3881 , P1_U3882;
wire P1_U3883 , P1_U3884 , P1_U3885 , P1_U3886 , P1_U3887 , P1_U3888 , P1_U3889 , P1_U3890 , P1_U3891 , P1_U3892;
wire P1_U3893 , P1_U3894 , P1_U3895 , P1_U3896 , P1_U3897 , P1_U3898 , P1_U3899 , P1_U3900 , P1_U3901 , P1_U3902;
wire P1_U3903 , P1_U3904 , P1_U3905 , P1_U3906 , P1_U3907 , P1_U3908 , P1_U3909 , P1_U3910 , P1_U3911 , P1_U3912;
wire P1_U3913 , P1_U3914 , P1_U3915 , P1_U3916 , P1_U3917 , P1_U3918 , P1_U3919 , P1_U3920 , P1_U3921 , P1_U3922;
wire P1_U3923 , P1_U3924 , P1_U3925 , P1_U3926 , P1_U3927 , P1_U3928 , P1_U3929 , P1_U3930 , P1_U3931 , P1_U3932;
wire P1_U3933 , P1_U3934 , P1_U3935 , P1_U3936 , P1_U3937 , P1_U3938 , P1_U3939 , P1_U3940 , P1_U3941 , P1_U3942;
wire P1_U3943 , P1_U3944 , P1_U3945 , P1_U3946 , P1_U3947 , P1_U3948 , P1_U3949 , P1_U3950 , P1_U3951 , P1_U3952;
wire P1_U3953 , P1_U3954 , P1_U3955 , P1_U3956 , P1_U3957 , P1_U3958 , P1_U3959 , P1_U3960 , P1_U3961 , P1_U3962;
wire P1_U3963 , P1_U3964 , P1_U3965 , P1_U3966 , P1_U3967 , P1_U3968 , P1_U3969 , P1_U3970 , P1_U3971 , P1_U3972;
wire P1_U3973 , P1_U3974 , P1_U3975 , P1_U3976 , P1_U3977 , P1_U3978 , P1_U3979 , P1_U3980 , P1_U3981 , P1_U3982;
wire P1_U3983 , P1_U3984 , P1_U3985 , P1_U3986 , P1_U3987 , P1_U3988 , P1_U3989 , P1_U3990 , P1_U3991 , P1_U3992;
wire P1_U3993 , P1_U3994 , P1_U3995 , P1_U3996 , P1_U3997 , P1_U3998 , P1_U3999 , P1_U4000 , P1_U4001 , P1_U4002;
wire P1_U4003 , P1_U4004 , P1_U4005 , P1_U4007 , P1_U4008 , P1_U4009 , P1_U4010 , P1_U4011 , P1_U4012 , P1_U4013;
wire P1_U4014 , P1_U4015 , P1_U4016 , P1_U4017 , P1_U4018 , P1_U4019 , P1_U4020 , P1_U4021 , P1_U4022 , P1_U4023;
wire P1_U4024 , P1_U4025 , P1_U4026 , P1_U4027 , P1_U4028 , P1_U4029 , P1_U4030 , P1_U4031 , P1_U4032 , P1_U4033;
wire P1_U4034 , P1_U4035 , P1_U4036 , P1_U4037 , P1_U4038 , P1_U4039 , P1_U4040 , P1_U4041 , P1_U4042 , P1_U4043;
wire P1_U4044 , P1_U4045 , P1_U4046 , P1_U4047 , P1_U4048 , P1_U4049 , P1_U4050 , P1_U4051 , P1_U4052 , P1_U4053;
wire P1_U4054 , P1_U4055 , P1_U4056 , P1_U4057 , P1_U4058 , P1_U4059 , P1_U4060 , P1_U4061 , P1_U4062 , P1_U4063;
wire P1_U4064 , P1_U4065 , P1_U4066 , P1_U4067 , P1_U4068 , P1_U4069 , P1_U4070 , P1_U4071 , P1_U4072 , P1_U4073;
wire P1_U4074 , P1_U4075 , P1_U4076 , P1_U4077 , P1_U4078 , P1_U4079 , P1_U4080 , P1_U4081 , P1_U4082 , P1_U4083;
wire P1_U4084 , P1_U4085 , P1_U4086 , P1_U4087 , P1_U4088 , P1_U4089 , P1_U4090 , P1_U4091 , P1_U4092 , P1_U4093;
wire P1_U4094 , P1_U4095 , P1_U4096 , P1_U4097 , P1_U4098 , P1_U4099 , P1_U4100 , P1_U4101 , P1_U4102 , P1_U4103;
wire P1_U4104 , P1_U4105 , P1_U4106 , P1_U4107 , P1_U4108 , P1_U4109 , P1_U4110 , P1_U4111 , P1_U4112 , P1_U4113;
wire P1_U4114 , P1_U4115 , P1_U4116 , P1_U4117 , P1_U4118 , P1_U4119 , P1_U4120 , P1_U4121 , P1_U4122 , P1_U4123;
wire P1_U4124 , P1_U4125 , P1_U4126 , P1_U4127 , P1_U4128 , P1_U4129 , P1_U4130 , P1_U4131 , P1_U4132 , P1_U4133;
wire P1_U4134 , P1_U4135 , P1_U4136 , P1_U4137 , P1_U4138 , P1_U4139 , P1_U4140 , P1_U4141 , P1_U4142 , P1_U4143;
wire P1_U4144 , P1_U4145 , P1_U4146 , P1_U4147 , P1_U4148 , P1_U4149 , P1_U4150 , P1_U4151 , P1_U4152 , P1_U4153;
wire P1_U4154 , P1_U4155 , P1_U4156 , P1_U4157 , P1_U4158 , P1_U4159 , P1_U4160 , P1_U4161 , P1_U4162 , P1_U4163;
wire P1_U4164 , P1_U4165 , P1_U4166 , P1_U4167 , P1_U4168 , P1_U4169 , P1_U4170 , P1_U4171 , P1_U4172 , P1_U4173;
wire P1_U4174 , P1_U4175 , P1_U4176 , P1_U4177 , P1_U4178 , P1_U4179 , P1_U4180 , P1_U4181 , P1_U4182 , P1_U4183;
wire P1_U4184 , P1_U4185 , P1_U4186 , P1_U4187 , P1_U4188 , P1_U4189 , P1_U4190 , P1_U4191 , P1_U4192 , P1_U4193;
wire P1_U4194 , P1_U4195 , P1_U4196 , P1_U4197 , P1_U4198 , P1_U4199 , P1_U4200 , P1_U4201 , P1_U4202 , P1_U4203;
wire P1_U4204 , P1_U4205 , P1_U4206 , P1_U4207 , P1_U4208 , P1_U4209 , P1_U4210 , P1_U4211 , P1_U4212 , P1_U4213;
wire P1_U4214 , P1_U4215 , P1_U4216 , P1_U4217 , P1_U4218 , P1_U4219 , P1_U4220 , P1_U4221 , P1_U4222 , P1_U4223;
wire P1_U4224 , P1_U4225 , P1_U4226 , P1_U4227 , P1_U4228 , P1_U4229 , P1_U4230 , P1_U4231 , P1_U4232 , P1_U4233;
wire P1_U4234 , P1_U4235 , P1_U4236 , P1_U4237 , P1_U4238 , P1_U4239 , P1_U4240 , P1_U4241 , P1_U4242 , P1_U4243;
wire P1_U4244 , P1_U4245 , P1_U4246 , P1_U4247 , P1_U4248 , P1_U4249 , P1_U4250 , P1_U4251 , P1_U4252 , P1_U4253;
wire P1_U4254 , P1_U4255 , P1_U4256 , P1_U4257 , P1_U4258 , P1_U4259 , P1_U4260 , P1_U4261 , P1_U4262 , P1_U4263;
wire P1_U4264 , P1_U4265 , P1_U4266 , P1_U4267 , P1_U4268 , P1_U4269 , P1_U4270 , P1_U4271 , P1_U4272 , P1_U4273;
wire P1_U4274 , P1_U4275 , P1_U4276 , P1_U4277 , P1_U4278 , P1_U4279 , P1_U4280 , P1_U4281 , P1_U4282 , P1_U4283;
wire P1_U4284 , P1_U4285 , P1_U4286 , P1_U4287 , P1_U4288 , P1_U4289 , P1_U4290 , P1_U4291 , P1_U4292 , P1_U4293;
wire P1_U4294 , P1_U4295 , P1_U4296 , P1_U4297 , P1_U4298 , P1_U4299 , P1_U4300 , P1_U4301 , P1_U4302 , P1_U4303;
wire P1_U4304 , P1_U4305 , P1_U4306 , P1_U4307 , P1_U4308 , P1_U4309 , P1_U4310 , P1_U4311 , P1_U4312 , P1_U4313;
wire P1_U4314 , P1_U4315 , P1_U4316 , P1_U4317 , P1_U4318 , P1_U4319 , P1_U4320 , P1_U4321 , P1_U4322 , P1_U4323;
wire P1_U4324 , P1_U4325 , P1_U4326 , P1_U4327 , P1_U4328 , P1_U4329 , P1_U4330 , P1_U4331 , P1_U4332 , P1_U4333;
wire P1_U4334 , P1_U4335 , P1_U4336 , P1_U4337 , P1_U4338 , P1_U4339 , P1_U4340 , P1_U4341 , P1_U4342 , P1_U4343;
wire P1_U4344 , P1_U4345 , P1_U4346 , P1_U4347 , P1_U4348 , P1_U4349 , P1_U4350 , P1_U4351 , P1_U4352 , P1_U4353;
wire P1_U4354 , P1_U4355 , P1_U4356 , P1_U4357 , P1_U4358 , P1_U4359 , P1_U4360 , P1_U4361 , P1_U4362 , P1_U4363;
wire P1_U4364 , P1_U4365 , P1_U4366 , P1_U4367 , P1_U4368 , P1_U4369 , P1_U4370 , P1_U4371 , P1_U4372 , P1_U4373;
wire P1_U4374 , P1_U4375 , P1_U4376 , P1_U4377 , P1_U4378 , P1_U4379 , P1_U4380 , P1_U4381 , P1_U4382 , P1_U4383;
wire P1_U4384 , P1_U4385 , P1_U4386 , P1_U4387 , P1_U4388 , P1_U4389 , P1_U4390 , P1_U4391 , P1_U4392 , P1_U4393;
wire P1_U4394 , P1_U4395 , P1_U4396 , P1_U4397 , P1_U4398 , P1_U4399 , P1_U4400 , P1_U4401 , P1_U4402 , P1_U4403;
wire P1_U4404 , P1_U4405 , P1_U4406 , P1_U4407 , P1_U4408 , P1_U4409 , P1_U4410 , P1_U4411 , P1_U4412 , P1_U4413;
wire P1_U4414 , P1_U4415 , P1_U4416 , P1_U4417 , P1_U4418 , P1_U4419 , P1_U4420 , P1_U4421 , P1_U4422 , P1_U4423;
wire P1_U4424 , P1_U4425 , P1_U4426 , P1_U4427 , P1_U4428 , P1_U4429 , P1_U4430 , P1_U4431 , P1_U4432 , P1_U4433;
wire P1_U4434 , P1_U4435 , P1_U4436 , P1_U4437 , P1_U4438 , P1_U4439 , P1_U4440 , P1_U4441 , P1_U4442 , P1_U4443;
wire P1_U4444 , P1_U4445 , P1_U4446 , P1_U4447 , P1_U4448 , P1_U4449 , P1_U4450 , P1_U4451 , P1_U4452 , P1_U4453;
wire P1_U4454 , P1_U4455 , P1_U4456 , P1_U4457 , P1_U4458 , P1_U4459 , P1_U4460 , P1_U4461 , P1_U4462 , P1_U4463;
wire P1_U4464 , P1_U4465 , P1_U4466 , P1_U4467 , P1_U4468 , P1_U4469 , P1_U4470 , P1_U4471 , P1_U4472 , P1_U4473;
wire P1_U4474 , P1_U4475 , P1_U4476 , P1_U4477 , P1_U4478 , P1_U4479 , P1_U4480 , P1_U4481 , P1_U4482 , P1_U4483;
wire P1_U4484 , P1_U4485 , P1_U4486 , P1_U4487 , P1_U4488 , P1_U4489 , P1_U4490 , P1_U4491 , P1_U4492 , P1_U4493;
wire P1_U4494 , P1_U4495 , P1_U4496 , P1_U4497 , P1_U4498 , P1_U4499 , P1_U4500 , P1_U4501 , P1_U4502 , P1_U4503;
wire P1_U4504 , P1_U4505 , P1_U4506 , P1_U4507 , P1_U4508 , P1_U4509 , P1_U4510 , P1_U4511 , P1_U4512 , P1_U4513;
wire P1_U4514 , P1_U4515 , P1_U4516 , P1_U4517 , P1_U4518 , P1_U4519 , P1_U4520 , P1_U4521 , P1_U4522 , P1_U4523;
wire P1_U4524 , P1_U4525 , P1_U4526 , P1_U4527 , P1_U4528 , P1_U4529 , P1_U4530 , P1_U4531 , P1_U4532 , P1_U4533;
wire P1_U4534 , P1_U4535 , P1_U4536 , P1_U4537 , P1_U4538 , P1_U4539 , P1_U4540 , P1_U4541 , P1_U4542 , P1_U4543;
wire P1_U4544 , P1_U4545 , P1_U4546 , P1_U4547 , P1_U4548 , P1_U4549 , P1_U4550 , P1_U4551 , P1_U4552 , P1_U4553;
wire P1_U4554 , P1_U4555 , P1_U4556 , P1_U4557 , P1_U4558 , P1_U4559 , P1_U4560 , P1_U4561 , P1_U4562 , P1_U4563;
wire P1_U4564 , P1_U4565 , P1_U4566 , P1_U4567 , P1_U4568 , P1_U4569 , P1_U4570 , P1_U4571 , P1_U4572 , P1_U4573;
wire P1_U4574 , P1_U4575 , P1_U4576 , P1_U4577 , P1_U4578 , P1_U4579 , P1_U4580 , P1_U4581 , P1_U4582 , P1_U4583;
wire P1_U4584 , P1_U4585 , P1_U4586 , P1_U4587 , P1_U4588 , P1_U4589 , P1_U4590 , P1_U4591 , P1_U4592 , P1_U4593;
wire P1_U4594 , P1_U4595 , P1_U4596 , P1_U4597 , P1_U4598 , P1_U4599 , P1_U4600 , P1_U4601 , P1_U4602 , P1_U4603;
wire P1_U4604 , P1_U4605 , P1_U4606 , P1_U4607 , P1_U4608 , P1_U4609 , P1_U4610 , P1_U4611 , P1_U4612 , P1_U4613;
wire P1_U4614 , P1_U4615 , P1_U4616 , P1_U4617 , P1_U4618 , P1_U4619 , P1_U4620 , P1_U4621 , P1_U4622 , P1_U4623;
wire P1_U4624 , P1_U4625 , P1_U4626 , P1_U4627 , P1_U4628 , P1_U4629 , P1_U4630 , P1_U4631 , P1_U4632 , P1_U4633;
wire P1_U4634 , P1_U4635 , P1_U4636 , P1_U4637 , P1_U4638 , P1_U4639 , P1_U4640 , P1_U4641 , P1_U4642 , P1_U4643;
wire P1_U4644 , P1_U4645 , P1_U4646 , P1_U4647 , P1_U4648 , P1_U4649 , P1_U4650 , P1_U4651 , P1_U4652 , P1_U4653;
wire P1_U4654 , P1_U4655 , P1_U4656 , P1_U4657 , P1_U4658 , P1_U4659 , P1_U4660 , P1_U4661 , P1_U4662 , P1_U4663;
wire P1_U4664 , P1_U4665 , P1_U4666 , P1_U4667 , P1_U4668 , P1_U4669 , P1_U4670 , P1_U4671 , P1_U4672 , P1_U4673;
wire P1_U4674 , P1_U4675 , P1_U4676 , P1_U4677 , P1_U4678 , P1_U4679 , P1_U4680 , P1_U4681 , P1_U4682 , P1_U4683;
wire P1_U4684 , P1_U4685 , P1_U4686 , P1_U4687 , P1_U4688 , P1_U4689 , P1_U4690 , P1_U4691 , P1_U4692 , P1_U4693;
wire P1_U4694 , P1_U4695 , P1_U4696 , P1_U4697 , P1_U4698 , P1_U4699 , P1_U4700 , P1_U4701 , P1_U4702 , P1_U4703;
wire P1_U4704 , P1_U4705 , P1_U4706 , P1_U4707 , P1_U4708 , P1_U4709 , P1_U4710 , P1_U4711 , P1_U4712 , P1_U4713;
wire P1_U4714 , P1_U4715 , P1_U4716 , P1_U4717 , P1_U4718 , P1_U4719 , P1_U4720 , P1_U4721 , P1_U4722 , P1_U4723;
wire P1_U4724 , P1_U4725 , P1_U4726 , P1_U4727 , P1_U4728 , P1_U4729 , P1_U4730 , P1_U4731 , P1_U4732 , P1_U4733;
wire P1_U4734 , P1_U4735 , P1_U4736 , P1_U4737 , P1_U4738 , P1_U4739 , P1_U4740 , P1_U4741 , P1_U4742 , P1_U4743;
wire P1_U4744 , P1_U4745 , P1_U4746 , P1_U4747 , P1_U4748 , P1_U4749 , P1_U4750 , P1_U4751 , P1_U4752 , P1_U4753;
wire P1_U4754 , P1_U4755 , P1_U4756 , P1_U4757 , P1_U4758 , P1_U4759 , P1_U4760 , P1_U4761 , P1_U4762 , P1_U4763;
wire P1_U4764 , P1_U4765 , P1_U4766 , P1_U4767 , P1_U4768 , P1_U4769 , P1_U4770 , P1_U4771 , P1_U4772 , P1_U4773;
wire P1_U4774 , P1_U4775 , P1_U4776 , P1_U4777 , P1_U4778 , P1_U4779 , P1_U4780 , P1_U4781 , P1_U4782 , P1_U4783;
wire P1_U4784 , P1_U4785 , P1_U4786 , P1_U4787 , P1_U4788 , P1_U4789 , P1_U4790 , P1_U4791 , P1_U4792 , P1_U4793;
wire P1_U4794 , P1_U4795 , P1_U4796 , P1_U4797 , P1_U4798 , P1_U4799 , P1_U4800 , P1_U4801 , P1_U4802 , P1_U4803;
wire P1_U4804 , P1_U4805 , P1_U4806 , P1_U4807 , P1_U4808 , P1_U4809 , P1_U4810 , P1_U4811 , P1_U4812 , P1_U4813;
wire P1_U4814 , P1_U4815 , P1_U4816 , P1_U4817 , P1_U4818 , P1_U4819 , P1_U4820 , P1_U4821 , P1_U4822 , P1_U4823;
wire P1_U4824 , P1_U4825 , P1_U4826 , P1_U4827 , P1_U4828 , P1_U4829 , P1_U4830 , P1_U4831 , P1_U4832 , P1_U4833;
wire P1_U4834 , P1_U4835 , P1_U4836 , P1_U4837 , P1_U4838 , P1_U4839 , P1_U4840 , P1_U4841 , P1_U4842 , P1_U4843;
wire P1_U4844 , P1_U4845 , P1_U4846 , P1_U4847 , P1_U4848 , P1_U4849 , P1_U4850 , P1_U4851 , P1_U4852 , P1_U4853;
wire P1_U4854 , P1_U4855 , P1_U4856 , P1_U4857 , P1_U4858 , P1_U4859 , P1_U4860 , P1_U4861 , P1_U4862 , P1_U4863;
wire P1_U4864 , P1_U4865 , P1_U4866 , P1_U4867 , P1_U4868 , P1_U4869 , P1_U4870 , P1_U4871 , P1_U4872 , P1_U4873;
wire P1_U4874 , P1_U4875 , P1_U4876 , P1_U4877 , P1_U4878 , P1_U4879 , P1_U4880 , P1_U4881 , P1_U4882 , P1_U4883;
wire P1_U4884 , P1_U4885 , P1_U4886 , P1_U4887 , P1_U4888 , P1_U4889 , P1_U4890 , P1_U4891 , P1_U4892 , P1_U4893;
wire P1_U4894 , P1_U4895 , P1_U4896 , P1_U4897 , P1_U4898 , P1_U4899 , P1_U4900 , P1_U4901 , P1_U4902 , P1_U4903;
wire P1_U4904 , P1_U4905 , P1_U4906 , P1_U4907 , P1_U4908 , P1_U4909 , P1_U4910 , P1_U4911 , P1_U4912 , P1_U4913;
wire P1_U4914 , P1_U4915 , P1_U4916 , P1_U4917 , P1_U4918 , P1_U4919 , P1_U4920 , P1_U4921 , P1_U4922 , P1_U4923;
wire P1_U4924 , P1_U4925 , P1_U4926 , P1_U4927 , P1_U4928 , P1_U4929 , P1_U4930 , P1_U4931 , P1_U4932 , P1_U4933;
wire P1_U4934 , P1_U4935 , P1_U4936 , P1_U4937 , P1_U4938 , P1_U4939 , P1_U4940 , P1_U4941 , P1_U4942 , P1_U4943;
wire P1_U4944 , P1_U4945 , P1_U4946 , P1_U4947 , P1_U4948 , P1_U4949 , P1_U4950 , P1_U4951 , P1_U4952 , P1_U4953;
wire P1_U4954 , P1_U4955 , P1_U4956 , P1_U4957 , P1_U4958 , P1_U4959 , P1_U4960 , P1_U4961 , P1_U4962 , P1_U4963;
wire P1_U4964 , P1_U4965 , P1_U4966 , P1_U4967 , P1_U4968 , P1_U4969 , P1_U4970 , P1_U4971 , P1_U4972 , P1_U4973;
wire P1_U4974 , P1_U4975 , P1_U4976 , P1_U4977 , P1_U4978 , P1_U4979 , P1_U4980 , P1_U4981 , P1_U4982 , P1_U4983;
wire P1_U4984 , P1_U4985 , P1_U4986 , P1_U4987 , P1_U4988 , P1_U4989 , P1_U4990 , P1_U4991 , P1_U4992 , P1_U4993;
wire P1_U4994 , P1_U4995 , P1_U4996 , P1_U4997 , P1_U4998 , P1_U4999 , P1_U5000 , P1_U5001 , P1_U5002 , P1_U5003;
wire P1_U5004 , P1_U5005 , P1_U5006 , P1_U5007 , P1_U5008 , P1_U5009 , P1_U5010 , P1_U5011 , P1_U5012 , P1_U5013;
wire P1_U5014 , P1_U5015 , P1_U5016 , P1_U5017 , P1_U5018 , P1_U5019 , P1_U5020 , P1_U5021 , P1_U5022 , P1_U5023;
wire P1_U5024 , P1_U5025 , P1_U5026 , P1_U5027 , P1_U5028 , P1_U5029 , P1_U5030 , P1_U5031 , P1_U5032 , P1_U5033;
wire P1_U5034 , P1_U5035 , P1_U5036 , P1_U5037 , P1_U5038 , P1_U5039 , P1_U5040 , P1_U5041 , P1_U5042 , P1_U5043;
wire P1_U5044 , P1_U5045 , P1_U5046 , P1_U5047 , P1_U5048 , P1_U5049 , P1_U5050 , P1_U5051 , P1_U5052 , P1_U5053;
wire P1_U5054 , P1_U5055 , P1_U5056 , P1_U5057 , P1_U5058 , P1_U5059 , P1_U5060 , P1_U5061 , P1_U5062 , P1_U5063;
wire P1_U5064 , P1_U5065 , P1_U5066 , P1_U5067 , P1_U5068 , P1_U5069 , P1_U5070 , P1_U5071 , P1_U5072 , P1_U5073;
wire P1_U5074 , P1_U5075 , P1_U5076 , P1_U5077 , P1_U5078 , P1_U5079 , P1_U5080 , P1_U5081 , P1_U5082 , P1_U5083;
wire P1_U5084 , P1_U5085 , P1_U5086 , P1_U5087 , P1_U5088 , P1_U5089 , P1_U5090 , P1_U5091 , P1_U5092 , P1_U5093;
wire P1_U5094 , P1_U5095 , P1_U5096 , P1_U5097 , P1_U5098 , P1_U5099 , P1_U5100 , P1_U5101 , P1_U5102 , P1_U5103;
wire P1_U5104 , P1_U5105 , P1_U5106 , P1_U5107 , P1_U5108 , P1_U5109 , P1_U5110 , P1_U5111 , P1_U5112 , P1_U5113;
wire P1_U5114 , P1_U5115 , P1_U5116 , P1_U5117 , P1_U5118 , P1_U5119 , P1_U5120 , P1_U5121 , P1_U5122 , P1_U5123;
wire P1_U5124 , P1_U5125 , P1_U5126 , P1_U5127 , P1_U5128 , P1_U5129 , P1_U5130 , P1_U5131 , P1_U5132 , P1_U5133;
wire P1_U5134 , P1_U5135 , P1_U5136 , P1_U5137 , P1_U5138 , P1_U5139 , P1_U5140 , P1_U5141 , P1_U5142 , P1_U5143;
wire P1_U5144 , P1_U5145 , P1_U5146 , P1_U5147 , P1_U5148 , P1_U5149 , P1_U5150 , P1_U5151 , P1_U5152 , P1_U5153;
wire P1_U5154 , P1_U5155 , P1_U5156 , P1_U5157 , P1_U5158 , P1_U5159 , P1_U5160 , P1_U5161 , P1_U5162 , P1_U5163;
wire P1_U5164 , P1_U5165 , P1_U5166 , P1_U5167 , P1_U5168 , P1_U5169 , P1_U5170 , P1_U5171 , P1_U5172 , P1_U5173;
wire P1_U5174 , P1_U5175 , P1_U5176 , P1_U5177 , P1_U5178 , P1_U5179 , P1_U5180 , P1_U5181 , P1_U5182 , P1_U5183;
wire P1_U5184 , P1_U5185 , P1_U5186 , P1_U5187 , P1_U5188 , P1_U5189 , P1_U5190 , P1_U5191 , P1_U5192 , P1_U5193;
wire P1_U5194 , P1_U5195 , P1_U5196 , P1_U5197 , P1_U5198 , P1_U5199 , P1_U5200 , P1_U5201 , P1_U5202 , P1_U5203;
wire P1_U5204 , P1_U5205 , P1_U5206 , P1_U5207 , P1_U5208 , P1_U5209 , P1_U5210 , P1_U5211 , P1_U5212 , P1_U5213;
wire P1_U5214 , P1_U5215 , P1_U5216 , P1_U5217 , P1_U5218 , P1_U5219 , P1_U5220 , P1_U5221 , P1_U5222 , P1_U5223;
wire P1_U5224 , P1_U5225 , P1_U5226 , P1_U5227 , P1_U5228 , P1_U5229 , P1_U5230 , P1_U5231 , P1_U5232 , P1_U5233;
wire P1_U5234 , P1_U5235 , P1_U5236 , P1_U5237 , P1_U5238 , P1_U5239 , P1_U5240 , P1_U5241 , P1_U5242 , P1_U5243;
wire P1_U5244 , P1_U5245 , P1_U5246 , P1_U5247 , P1_U5248 , P1_U5249 , P1_U5250 , P1_U5251 , P1_U5252 , P1_U5253;
wire P1_U5254 , P1_U5255 , P1_U5256 , P1_U5257 , P1_U5258 , P1_U5259 , P1_U5260 , P1_U5261 , P1_U5262 , P1_U5263;
wire P1_U5264 , P1_U5265 , P1_U5266 , P1_U5267 , P1_U5268 , P1_U5269 , P1_U5270 , P1_U5271 , P1_U5272 , P1_U5273;
wire P1_U5274 , P1_U5275 , P1_U5276 , P1_U5277 , P1_U5278 , P1_U5279 , P1_U5280 , P1_U5281 , P1_U5282 , P1_U5283;
wire P1_U5284 , P1_U5285 , P1_U5286 , P1_U5287 , P1_U5288 , P1_U5289 , P1_U5290 , P1_U5291 , P1_U5292 , P1_U5293;
wire P1_U5294 , P1_U5295 , P1_U5296 , P1_U5297 , P1_U5298 , P1_U5299 , P1_U5300 , P1_U5301 , P1_U5302 , P1_U5303;
wire P1_U5304 , P1_U5305 , P1_U5306 , P1_U5307 , P1_U5308 , P1_U5309 , P1_U5310 , P1_U5311 , P1_U5312 , P1_U5313;
wire P1_U5314 , P1_U5315 , P1_U5316 , P1_U5317 , P1_U5318 , P1_U5319 , P1_U5320 , P1_U5321 , P1_U5322 , P1_U5323;
wire P1_U5324 , P1_U5325 , P1_U5326 , P1_U5327 , P1_U5328 , P1_U5329 , P1_U5330 , P1_U5331 , P1_U5332 , P1_U5333;
wire P1_U5334 , P1_U5335 , P1_U5336 , P1_U5337 , P1_U5338 , P1_U5339 , P1_U5340 , P1_U5341 , P1_U5342 , P1_U5343;
wire P1_U5344 , P1_U5345 , P1_U5346 , P1_U5347 , P1_U5348 , P1_U5349 , P1_U5350 , P1_U5351 , P1_U5352 , P1_U5353;
wire P1_U5354 , P1_U5355 , P1_U5356 , P1_U5357 , P1_U5358 , P1_U5359 , P1_U5360 , P1_U5361 , P1_U5362 , P1_U5363;
wire P1_U5364 , P1_U5365 , P1_U5366 , P1_U5367 , P1_U5368 , P1_U5369 , P1_U5370 , P1_U5371 , P1_U5372 , P1_U5373;
wire P1_U5374 , P1_U5375 , P1_U5376 , P1_U5377 , P1_U5378 , P1_U5379 , P1_U5380 , P1_U5381 , P1_U5382 , P1_U5383;
wire P1_U5384 , P1_U5385 , P1_U5386 , P1_U5387 , P1_U5388 , P1_U5389 , P1_U5390 , P1_U5391 , P1_U5392 , P1_U5393;
wire P1_U5394 , P1_U5395 , P1_U5396 , P1_U5397 , P1_U5398 , P1_U5399 , P1_U5400 , P1_U5401 , P1_U5402 , P1_U5403;
wire P1_U5404 , P1_U5405 , P1_U5406 , P1_U5407 , P1_U5408 , P1_U5409 , P1_U5410 , P1_U5411 , P1_U5412 , P1_U5413;
wire P1_U5414 , P1_U5415 , P1_U5416 , P1_U5417 , P1_U5418 , P1_U5419 , P1_U5420 , P1_U5421 , P1_U5422 , P1_U5423;
wire P1_U5424 , P1_U5425 , P1_U5426 , P1_U5427 , P1_U5428 , P1_U5429 , P1_U5430 , P1_U5431 , P1_U5432 , P1_U5433;
wire P1_U5434 , P1_U5435 , P1_U5436 , P1_U5437 , P1_U5438 , P1_U5439 , P1_U5440 , P1_U5441 , P1_U5442 , P1_U5443;
wire P1_U5444 , P1_U5445 , P1_U5446 , P1_U5447 , P1_U5448 , P1_U5449 , P1_U5450 , P1_U5451 , P1_U5452 , P1_U5453;
wire P1_U5454 , P1_U5455 , P1_U5456 , P1_U5457 , P1_U5458 , P1_U5459 , P1_U5460 , P1_U5461 , P1_U5462 , P1_U5463;
wire P1_U5464 , P1_U5465 , P1_U5466 , P1_U5467 , P1_U5468 , P1_U5469 , P1_U5470 , P1_U5471 , P1_U5472 , P1_U5473;
wire P1_U5474 , P1_U5475 , P1_U5476 , P1_U5477 , P1_U5478 , P1_U5479 , P1_U5480 , P1_U5481 , P1_U5482 , P1_U5483;
wire P1_U5484 , P1_U5485 , P1_U5486 , P1_U5487 , P1_U5488 , P1_U5489 , P1_U5490 , P1_U5491 , P1_U5492 , P1_U5493;
wire P1_U5494 , P1_U5495 , P1_U5496 , P1_U5497 , P1_U5498 , P1_U5499 , P1_U5500 , P1_U5501 , P1_U5502 , P1_U5503;
wire P1_U5504 , P1_U5505 , P1_U5506 , P1_U5507 , P1_U5508 , P1_U5509 , P1_U5510 , P1_U5511 , P1_U5512 , P1_U5513;
wire P1_U5514 , P1_U5515 , P1_U5516 , P1_U5517 , P1_U5518 , P1_U5519 , P1_U5520 , P1_U5521 , P1_U5522 , P1_U5523;
wire P1_U5524 , P1_U5525 , P1_U5526 , P1_U5527 , P1_U5528 , P1_U5529 , P1_U5530 , P1_U5531 , P1_U5532 , P1_U5533;
wire P1_U5534 , P1_U5535 , P1_U5536 , P1_U5537 , P1_U5538 , P1_U5539 , P1_U5540 , P1_U5541 , P1_U5542 , P1_U5543;
wire P1_U5544 , P1_U5545 , P1_U5546 , P1_U5547 , P1_U5548 , P1_U5549 , P1_U5550 , P1_U5551 , P1_U5552 , P1_U5553;
wire P1_U5554 , P1_U5555 , P1_U5556 , P1_U5557 , P1_U5558 , P1_U5559 , P1_U5560 , P1_U5561 , P1_U5562 , P1_U5563;
wire P1_U5564 , P1_U5565 , P1_U5566 , P1_U5567 , P1_U5568 , P1_U5569 , P1_U5570 , P1_U5571 , P1_U5572 , P1_U5573;
wire P1_U5574 , P1_U5575 , P1_U5576 , P1_U5577 , P1_U5578 , P1_U5579 , P1_U5580 , P1_U5581 , P1_U5582 , P1_U5583;
wire P1_U5584 , P1_U5585 , P1_U5586 , P1_U5587 , P1_U5588 , P1_U5589 , P1_U5590 , P1_U5591 , P1_U5592 , P1_U5593;
wire P1_U5594 , P1_U5595 , P1_U5596 , P1_U5597 , P1_U5598 , P1_U5599 , P1_U5600 , P1_U5601 , P1_U5602 , P1_U5603;
wire P1_U5604 , P1_U5605 , P1_U5606 , P1_U5607 , P1_U5608 , P1_U5609 , P1_U5610 , P1_U5611 , P1_U5612 , P1_U5613;
wire P1_U5614 , P1_U5615 , P1_U5616 , P1_U5617 , P1_U5618 , P1_U5619 , P1_U5620 , P1_U5621 , P1_U5622 , P1_U5623;
wire P1_U5624 , P1_U5625 , P1_U5626 , P1_U5627 , P1_U5628 , P1_U5629 , P1_U5630 , P1_U5631 , P1_U5632 , P1_U5633;
wire P1_U5634 , P1_U5635 , P1_U5636 , P1_U5637 , P1_U5638 , P1_U5639 , P1_U5640 , P1_U5641 , P1_U5642 , P1_U5643;
wire P1_U5644 , P1_U5645 , P1_U5646 , P1_U5647 , P1_U5648 , P1_U5649 , P1_U5650 , P1_U5651 , P1_U5652 , P1_U5653;
wire P1_U5654 , P1_U5655 , P1_U5656 , P1_U5657 , P1_U5658 , P1_U5659 , P1_U5660 , P1_U5661 , P1_U5662 , P1_U5663;
wire P1_U5664 , P1_U5665 , P1_U5666 , P1_U5667 , P1_U5668 , P1_U5669 , P1_U5670 , P1_U5671 , P1_U5672 , P1_U5673;
wire P1_U5674 , P1_U5675 , P1_U5676 , P1_U5677 , P1_U5678 , P1_U5679 , P1_U5680 , P1_U5681 , P1_U5682 , P1_U5683;
wire P1_U5684 , P1_U5685 , P1_U5686 , P1_U5687 , P1_U5688 , P1_U5689 , P1_U5690 , P1_U5691 , P1_U5692 , P1_U5693;
wire P1_U5694 , P1_U5695 , P1_U5696 , P1_U5697 , P1_U5698 , P1_U5699 , P1_U5700 , P1_U5701 , P1_U5702 , P1_U5703;
wire P1_U5704 , P1_U5705 , P1_U5706 , P1_U5707 , P1_U5708 , P1_U5709 , P1_U5710 , P1_U5711 , P1_U5712 , P1_U5713;
wire P1_U5714 , P1_U5715 , P1_U5716 , P1_U5717 , P1_U5718 , P1_U5719 , P1_U5720 , P1_U5721 , P1_U5722 , P1_U5723;
wire P1_U5724 , P1_U5725 , P1_U5726 , P1_U5727 , P1_U5728 , P1_U5729 , P1_U5730 , P1_U5731 , P1_U5732 , P1_U5733;
wire P1_U5734 , P1_U5735 , P1_U5736 , P1_U5737 , P1_U5738 , P1_U5739 , P1_U5740 , P1_U5741 , P1_U5742 , P1_U5743;
wire P1_U5744 , P1_U5745 , P1_U5746 , P1_U5747 , P1_U5748 , P1_U5749 , P1_U5750 , P1_U5751 , P1_U5752 , P1_U5753;
wire P1_U5754 , P1_U5755 , P1_U5756 , P1_U5757 , P1_U5758 , P1_U5759 , P1_U5760 , P1_U5761 , P1_U5762 , P1_U5763;
wire P1_U5764 , P1_U5765 , P1_U5766 , P1_U5767 , P1_U5768 , P1_U5769 , P1_U5770 , P1_U5771 , P1_U5772 , P1_U5773;
wire P1_U5774 , P1_U5775 , P1_U5776 , P1_U5777 , P1_U5778 , P1_U5779 , P1_U5780 , P1_U5781 , P1_U5782 , P1_U5783;
wire P1_U5784 , P1_U5785 , P1_U5786 , P1_U5787 , P1_U5788 , P1_U5789 , P1_U5790 , P1_U5791 , P1_U5792 , P1_U5793;
wire P1_U5794 , P1_U5795 , P1_U5796 , P1_U5797 , P1_U5798 , P1_U5799 , P1_U5800 , P1_U5801 , P1_U5802 , P1_U5803;
wire P1_U5804 , P1_U5805 , P1_U5806 , P1_U5807 , P1_U5808 , P1_U5809 , P1_U5810 , P1_U5811 , P1_U5812 , P1_U5813;
wire P1_U5814 , P1_U5815 , P1_U5816 , P1_U5817 , P1_U5818 , P1_U5819 , P1_U5820 , P1_U5821 , P1_U5822 , P1_U5823;
wire P1_U5824 , P1_U5825 , P1_U5826 , P1_U5827 , P1_U5828 , P1_U5829 , P1_U5830 , P1_U5831 , P1_U5832 , P1_U5833;
wire P1_U5834 , P1_U5835 , P1_U5836 , P1_U5837 , P1_U5838 , P1_U5839 , P1_U5840 , P1_U5841 , P1_U5842 , P1_U5843;
wire P1_U5844 , P1_U5845 , P1_U5846 , P1_U5847 , P1_U5848 , P1_U5849 , P1_U5850 , P1_U5851 , P1_U5852 , P1_U5853;
wire P1_U5854 , P1_U5855 , P1_U5856 , P1_U5857 , P1_U5858 , P1_U5859 , P1_U5860 , P1_U5861 , P1_U5862 , P1_U5863;
wire P1_U5864 , P1_U5865 , P1_U5866 , P1_U5867 , P1_U5868 , P1_U5869 , P1_U5870 , P1_U5871 , P1_U5872 , P1_U5873;
wire P1_U5874 , P1_U5875 , P1_U5876 , P1_U5877 , P1_U5878 , P1_U5879 , P1_U5880 , P1_U5881 , P1_U5882 , P1_U5883;
wire P1_U5884 , P1_U5885 , P1_U5886 , P1_U5887 , P1_U5888 , P1_U5889 , P1_U5890 , P1_U5891 , P1_U5892 , P1_U5893;
wire P1_U5894 , P1_U5895 , P1_U5896 , P1_U5897 , P1_U5898 , P1_U5899 , P1_U5900 , P1_U5901 , P1_U5902 , P1_U5903;
wire P1_U5904 , P1_U5905 , P1_U5906 , P1_U5907 , P1_U5908 , P1_U5909 , P1_U5910 , P1_U5911 , P1_U5912 , P1_U5913;
wire P1_U5914 , P1_U5915 , P1_U5916 , P1_U5917 , P1_U5918 , P1_U5919 , P1_U5920 , P1_U5921 , P1_U5922 , P1_U5923;
wire P1_U5924 , P1_U5925 , P1_U5926 , P1_U5927 , P1_U5928 , P1_U5929 , P1_U5930 , P1_U5931 , P1_U5932 , P1_U5933;
wire P1_U5934 , P1_U5935 , P1_U5936 , P1_U5937 , P1_U5938 , P1_U5939 , P1_U5940 , P1_U5941 , P1_U5942 , P1_U5943;
wire P1_U5944 , P1_U5945 , P1_U5946 , P1_U5947 , P1_U5948 , P1_U5949 , P1_U5950 , P1_U5951 , P1_U5952 , P1_U5953;
wire P1_U5954 , P1_U5955 , P1_U5956 , P1_U5957 , P1_U5958 , P1_U5959 , P1_U5960 , P1_U5961 , P1_U5962 , P1_U5963;
wire P1_U5964 , P1_U5965 , P1_U5966 , P1_U5967 , P1_U5968 , P1_U5969 , P1_U5970 , P1_U5971 , P1_U5972 , P1_U5973;
wire P1_U5974 , P1_U5975 , P1_U5976 , P1_U5977 , P1_U5978 , P1_U5979 , P1_U5980 , P1_U5981 , P1_U5982 , P1_U5983;
wire P1_U5984 , P1_U5985 , P1_U5986 , P1_U5987 , P1_U5988 , P1_U5989 , P1_U5990 , P1_U5991 , P1_U5992 , P1_U5993;
wire P1_U5994 , P1_U5995 , P1_U5996 , P1_U5997 , P1_U5998 , P1_U5999 , P1_U6000 , P1_U6001 , P1_U6002 , P1_U6003;
wire P1_U6004 , P1_U6005 , P1_U6006 , P1_U6007 , P1_U6008 , P1_U6009 , P1_U6010 , P1_U6011 , P1_U6012 , P1_U6013;
wire P1_U6014 , P1_U6015 , P1_U6016 , P1_U6017 , P1_U6018 , P1_U6019 , P1_U6020 , P1_U6021 , P1_U6022 , P1_U6023;
wire P1_U6024 , P1_U6025 , P1_U6026 , P1_U6027 , P1_U6028 , P1_U6029 , P1_U6030 , P1_U6031 , P1_U6032 , P1_U6033;
wire P1_U6034 , P1_U6035 , P1_U6036 , P1_U6037 , P1_U6038 , P1_U6039 , P1_U6040 , P1_U6041 , P1_U6042 , P1_U6043;
wire P1_U6044 , P1_U6045 , P1_U6046 , P1_U6047 , P1_U6048 , P1_U6049 , P1_U6050 , P1_U6051 , P1_U6052 , P1_U6053;
wire P1_U6054 , P1_U6055 , P1_U6056 , P1_U6057 , P1_U6058 , P1_U6059 , P1_U6060 , P1_U6061 , P1_U6062 , P1_U6063;
wire P1_U6064 , P1_U6065 , P1_U6066 , P1_U6067 , P1_U6068 , P1_U6069 , P1_U6070 , P1_U6071 , P1_U6072 , P1_U6073;
wire P1_U6074 , P1_U6075 , P1_U6076 , P1_U6077 , P1_U6078 , P1_U6079 , P1_U6080 , P1_U6081 , P1_U6082 , P1_U6083;
wire P1_U6084 , P1_U6085 , P1_U6086 , P1_U6087 , P1_U6088 , P1_U6089 , P1_U6090 , P1_U6091 , P1_U6092 , P1_U6093;
wire P1_U6094 , P1_U6095 , P1_U6096 , P1_U6097 , P1_U6098 , P1_U6099 , P1_U6100 , P1_U6101 , P1_U6102 , P1_U6103;
wire P1_U6104 , P1_U6105 , P1_U6106 , P1_U6107 , P1_U6108 , P1_U6109 , P1_U6110 , P1_U6111 , P1_U6112 , P1_U6113;
wire P1_U6114 , P1_U6115 , P1_U6116 , P1_U6117 , P1_U6118 , P1_U6119 , P1_U6120 , P1_U6121 , P1_U6122 , P1_U6123;
wire P1_U6124 , P1_U6125 , P1_U6126 , P1_U6127 , P1_U6128 , P1_U6129 , P1_U6130 , P1_U6131 , P1_U6132 , P1_U6133;
wire P1_U6134 , P1_U6135 , P1_U6136 , P1_U6137 , P1_U6138 , P1_U6139 , P1_U6140 , P1_U6141 , P1_U6142 , P1_U6143;
wire P1_U6144 , P1_U6145 , P1_U6146 , P1_U6147 , P1_U6148 , P1_U6149 , P1_U6150 , P1_U6151 , P1_U6152 , P1_U6153;
wire P1_U6154 , P1_U6155 , P1_U6156 , P1_U6157 , P1_U6158 , P1_U6159 , P1_U6160 , P1_U6161 , P1_U6162 , P1_U6163;
wire P1_U6164 , P1_U6165 , P1_U6166 , P1_U6167 , P1_U6168 , P1_U6169 , P1_U6170 , P1_U6171 , P1_U6172 , P1_U6173;
wire P1_U6174 , P1_U6175 , P1_U6176 , P1_U6177 , P1_U6178 , P1_U6179 , P1_U6180 , P1_U6181 , P1_U6182 , P1_U6183;
wire P1_U6184 , P1_U6185 , P1_U6186 , P1_U6187 , P1_U6188 , P1_U6189 , P1_U6190 , P1_U6191 , P1_U6192 , P1_U6193;
wire P1_U6194 , P1_U6195 , P1_U6196 , P1_U6197 , P1_U6198 , P1_U6199 , P1_U6200 , P1_U6201 , P1_U6202 , P1_U6203;
wire P1_U6204 , P1_U6205 , P1_U6206 , P1_U6207 , P1_U6208 , P1_U6209 , P1_U6210 , P1_U6211 , P1_U6212 , P1_U6213;
wire P1_U6214 , P1_U6215 , P1_U6216 , P1_U6217 , P1_U6218 , P1_U6219 , P1_U6220 , P1_U6221 , P1_U6222 , P1_U6223;
wire P1_U6224 , P1_U6225 , P1_U6226 , P1_U6227 , P1_U6228 , P1_U6229 , P1_U6230 , P1_U6231 , P1_U6232 , P1_U6233;
wire P1_U6234 , P1_U6235 , P1_U6236 , P1_U6237 , P1_U6238 , P1_U6239 , P1_U6240 , P1_U6241 , P1_U6242 , P1_U6243;
wire P1_U6244 , P1_U6245 , P1_U6246 , P1_U6247 , P1_U6248 , P1_U6249 , P1_U6250 , P1_U6251 , P1_U6252 , P1_U6253;
wire P1_U6254 , P1_U6255 , P1_U6256 , P1_U6257 , P1_U6258 , P1_U6259 , P1_U6260 , P1_U6261 , P1_U6262 , P1_U6263;
wire P1_U6264 , P1_U6265 , P1_U6266 , P2_R1113_U462 , P2_R1113_U461 , P2_R1113_U460 , P2_R1113_U459 , P2_R1113_U458 , P2_R1113_U457 , P2_R1113_U456;
wire P2_R1113_U455 , P2_R1113_U454 , P2_R1113_U453 , P2_R1113_U452 , P2_R1113_U451 , P2_R1113_U450 , P2_R1113_U449 , P2_R1113_U448 , P2_R1113_U447 , P2_R1113_U446;
wire P2_R1113_U445 , P2_R1113_U444 , P2_R1113_U443 , P2_R1113_U442 , P2_R1113_U441 , P2_R1113_U440 , P2_R1113_U439 , P2_U3014 , P2_U3015 , P2_U3016;
wire P2_U3017 , P2_U3018 , P2_U3019 , P2_U3020 , P2_U3021 , P2_U3022 , P2_U3023 , P2_U3024 , P2_U3025 , P2_U3026;
wire P2_U3027 , P2_U3028 , P2_U3029 , P2_U3030 , P2_U3031 , P2_U3032 , P2_U3033 , P2_U3034 , P2_U3035 , P2_U3036;
wire P2_U3037 , P2_U3038 , P2_U3039 , P2_U3040 , P2_U3041 , P2_U3042 , P2_U3043 , P2_U3044 , P2_U3045 , P2_U3046;
wire P2_U3047 , P2_U3048 , P2_U3049 , P2_U3050 , P2_U3051 , P2_U3052 , P2_U3053 , P2_U3054 , P2_U3055 , P2_U3056;
wire P2_U3057 , P2_U3058 , P2_U3059 , P2_U3060 , P2_U3061 , P2_U3062 , P2_U3063 , P2_U3064 , P2_U3065 , P2_U3066;
wire P2_U3067 , P2_U3068 , P2_U3069 , P2_U3070 , P2_U3071 , P2_U3072 , P2_U3073 , P2_U3074 , P2_U3075 , P2_U3076;
wire P2_U3077 , P2_U3078 , P2_U3079 , P2_U3080 , P2_U3081 , P2_U3082 , P2_U3083 , P2_U3084 , P2_U3085 , P2_U3086;
wire P2_U3087 , P2_U3088 , P2_U3089 , P2_U3090 , P2_U3091 , P2_U3092 , P2_U3093 , P2_U3094 , P2_U3095 , P2_U3096;
wire P2_U3097 , P2_U3098 , P2_U3099 , P2_U3100 , P2_U3101 , P2_U3102 , P2_U3103 , P2_U3104 , P2_U3105 , P2_U3106;
wire P2_U3107 , P2_U3108 , P2_U3109 , P2_U3110 , P2_U3111 , P2_U3112 , P2_U3113 , P2_U3114 , P2_U3115 , P2_U3116;
wire P2_U3117 , P2_U3118 , P2_U3119 , P2_U3120 , P2_U3121 , P2_U3122 , P2_U3123 , P2_U3124 , P2_U3125 , P2_U3126;
wire P2_U3127 , P2_U3128 , P2_U3129 , P2_U3130 , P2_U3131 , P2_U3132 , P2_U3133 , P2_U3134 , P2_U3135 , P2_U3136;
wire P2_U3137 , P2_U3138 , P2_U3139 , P2_U3140 , P2_U3141 , P2_U3142 , P2_U3143 , P2_U3144 , P2_U3145 , P2_U3146;
wire P2_U3147 , P2_U3148 , P2_U3149 , P2_U3150 , P2_U3153 , P2_U3154 , P2_U3155 , P2_U3156 , P2_U3157 , P2_U3158;
wire P2_U3159 , P2_U3160 , P2_U3161 , P2_U3162 , P2_U3163 , P2_U3164 , P2_U3165 , P2_U3166 , P2_U3167 , P2_U3168;
wire P2_U3169 , P2_U3170 , P2_U3171 , P2_U3172 , P2_U3173 , P2_U3174 , P2_U3175 , P2_U3176 , P2_U3177 , P2_U3178;
wire P2_U3179 , P2_U3180 , P2_U3181 , P2_U3182 , P2_U3183 , P2_U3184 , P2_U3185 , P2_U3186 , P2_U3187 , P2_U3188;
wire P2_U3189 , P2_U3190 , P2_U3191 , P2_U3192 , P2_U3193 , P2_U3194 , P2_U3195 , P2_U3196 , P2_U3197 , P2_U3198;
wire P2_U3199 , P2_U3200 , P2_U3201 , P2_U3202 , P2_U3203 , P2_U3204 , P2_U3205 , P2_U3206 , P2_U3207 , P2_U3208;
wire P2_U3209 , P2_U3210 , P2_U3211 , P2_U3212 , P2_U3213 , P2_U3214 , P2_U3359 , P2_U3360 , P2_U3361 , P2_U3362;
wire P2_U3363 , P2_U3364 , P2_U3365 , P2_U3366 , P2_U3367 , P2_U3368 , P2_U3369 , P2_U3370 , P2_U3371 , P2_U3372;
wire P2_U3373 , P2_U3374 , P2_U3375 , P2_U3376 , P2_U3377 , P2_U3378 , P2_U3379 , P2_U3380 , P2_U3381 , P2_U3382;
wire P2_U3383 , P2_U3384 , P2_U3385 , P2_U3386 , P2_U3387 , P2_U3388 , P2_U3389 , P2_U3390 , P2_U3391 , P2_U3392;
wire P2_U3393 , P2_U3394 , P2_U3395 , P2_U3396 , P2_U3397 , P2_U3398 , P2_U3399 , P2_U3400 , P2_U3401 , P2_U3402;
wire P2_U3403 , P2_U3404 , P2_U3405 , P2_U3406 , P2_U3407 , P2_U3408 , P2_U3409 , P2_U3410 , P2_U3411 , P2_U3412;
wire P2_U3413 , P2_U3414 , P2_U3415 , P2_U3416 , P2_U3417 , P2_U3418 , P2_U3419 , P2_U3420 , P2_U3421 , P2_U3422;
wire P2_U3423 , P2_U3424 , P2_U3425 , P2_U3426 , P2_U3427 , P2_U3428 , P2_U3429 , P2_U3430 , P2_U3431 , P2_U3432;
wire P2_U3433 , P2_U3434 , P2_U3435 , P2_U3436 , P2_U3439 , P2_U3440 , P2_U3441 , P2_U3442 , P2_U3443 , P2_U3444;
wire P2_U3445 , P2_U3446 , P2_U3447 , P2_U3448 , P2_U3449 , P2_U3450 , P2_U3452 , P2_U3453 , P2_U3455 , P2_U3456;
wire P2_U3458 , P2_U3459 , P2_U3461 , P2_U3462 , P2_U3464 , P2_U3465 , P2_U3467 , P2_U3468 , P2_U3470 , P2_U3471;
wire P2_U3473 , P2_U3474 , P2_U3476 , P2_U3477 , P2_U3479 , P2_U3480 , P2_U3482 , P2_U3483 , P2_U3485 , P2_U3486;
wire P2_U3488 , P2_U3489 , P2_U3491 , P2_U3492 , P2_U3494 , P2_U3495 , P2_U3497 , P2_U3498 , P2_U3500 , P2_U3501;
wire P2_U3503 , P2_U3504 , P2_U3506 , P2_U3584 , P2_U3585 , P2_U3586 , P2_U3587 , P2_U3588 , P2_U3589 , P2_U3590;
wire P2_U3591 , P2_U3592 , P2_U3593 , P2_U3594 , P2_U3595 , P2_U3596 , P2_U3597 , P2_U3598 , P2_U3599 , P2_U3600;
wire P2_U3601 , P2_U3602 , P2_U3603 , P2_U3604 , P2_U3605 , P2_U3606 , P2_U3607 , P2_U3608 , P2_U3609 , P2_U3610;
wire P2_U3611 , P2_U3612 , P2_U3613 , P2_U3614 , P2_U3615 , P2_U3616 , P2_U3617 , P2_U3618 , P2_U3619 , P2_U3620;
wire P2_U3621 , P2_U3622 , P2_U3623 , P2_U3624 , P2_U3625 , P2_U3626 , P2_U3627 , P2_U3628 , P2_U3629 , P2_U3630;
wire P2_U3631 , P2_U3632 , P2_U3633 , P2_U3634 , P2_U3635 , P2_U3636 , P2_U3637 , P2_U3638 , P2_U3639 , P2_U3640;
wire P2_U3641 , P2_U3642 , P2_U3643 , P2_U3644 , P2_U3645 , P2_U3646 , P2_U3647 , P2_U3648 , P2_U3649 , P2_U3650;
wire P2_U3651 , P2_U3652 , P2_U3653 , P2_U3654 , P2_U3655 , P2_U3656 , P2_U3657 , P2_U3658 , P2_U3659 , P2_U3660;
wire P2_U3661 , P2_U3662 , P2_U3663 , P2_U3664 , P2_U3665 , P2_U3666 , P2_U3667 , P2_U3668 , P2_U3669 , P2_U3670;
wire P2_U3671 , P2_U3672 , P2_U3673 , P2_U3674 , P2_U3675 , P2_U3676 , P2_U3677 , P2_U3678 , P2_U3679 , P2_U3680;
wire P2_U3681 , P2_U3682 , P2_U3683 , P2_U3684 , P2_U3685 , P2_U3686 , P2_U3687 , P2_U3688 , P2_U3689 , P2_U3690;
wire P2_U3691 , P2_U3692 , P2_U3693 , P2_U3694 , P2_U3695 , P2_U3696 , P2_U3697 , P2_U3698 , P2_U3699 , P2_U3700;
wire P2_U3701 , P2_U3702 , P2_U3703 , P2_U3704 , P2_U3705 , P2_U3706 , P2_U3707 , P2_U3708 , P2_U3709 , P2_U3710;
wire P2_U3711 , P2_U3712 , P2_U3713 , P2_U3714 , P2_U3715 , P2_U3716 , P2_U3717 , P2_U3718 , P2_U3719 , P2_U3720;
wire P2_U3721 , P2_U3722 , P2_U3723 , P2_U3724 , P2_U3725 , P2_U3726 , P2_U3727 , P2_U3728 , P2_U3729 , P2_U3730;
wire P2_U3731 , P2_U3732 , P2_U3733 , P2_U3734 , P2_U3735 , P2_U3736 , P2_U3737 , P2_U3738 , P2_U3739 , P2_U3740;
wire P2_U3741 , P2_U3742 , P2_U3743 , P2_U3744 , P2_U3745 , P2_U3746 , P2_U3747 , P2_U3748 , P2_U3749 , P2_U3750;
wire P2_U3751 , P2_U3752 , P2_U3753 , P2_U3754 , P2_U3755 , P2_U3756 , P2_U3757 , P2_U3758 , P2_U3759 , P2_U3760;
wire P2_U3761 , P2_U3762 , P2_U3763 , P2_U3764 , P2_U3765 , P2_U3766 , P2_U3767 , P2_U3768 , P2_U3769 , P2_U3770;
wire P2_U3771 , P2_U3772 , P2_U3773 , P2_U3774 , P2_U3775 , P2_U3776 , P2_U3777 , P2_U3778 , P2_U3779 , P2_U3780;
wire P2_U3781 , P2_U3782 , P2_U3783 , P2_U3784 , P2_U3785 , P2_U3786 , P2_U3787 , P2_U3788 , P2_U3789 , P2_U3790;
wire P2_U3791 , P2_U3792 , P2_U3793 , P2_U3794 , P2_U3795 , P2_U3796 , P2_U3797 , P2_U3798 , P2_U3799 , P2_U3800;
wire P2_U3801 , P2_U3802 , P2_U3803 , P2_U3804 , P2_U3805 , P2_U3806 , P2_U3807 , P2_U3808 , P2_U3809 , P2_U3810;
wire P2_U3811 , P2_U3812 , P2_U3813 , P2_U3814 , P2_U3815 , P2_U3816 , P2_U3817 , P2_U3818 , P2_U3819 , P2_U3820;
wire P2_U3821 , P2_U3822 , P2_U3823 , P2_U3824 , P2_U3825 , P2_U3826 , P2_U3827 , P2_U3828 , P2_U3829 , P2_U3830;
wire P2_U3831 , P2_U3832 , P2_U3833 , P2_U3834 , P2_U3835 , P2_U3836 , P2_U3837 , P2_U3838 , P2_U3839 , P2_U3840;
wire P2_U3841 , P2_U3842 , P2_U3843 , P2_U3844 , P2_U3845 , P2_U3846 , P2_U3847 , P2_U3848 , P2_U3849 , P2_U3850;
wire P2_U3851 , P2_U3852 , P2_U3853 , P2_U3854 , P2_U3855 , P2_U3856 , P2_U3857 , P2_U3858 , P2_U3859 , P2_U3860;
wire P2_U3861 , P2_U3862 , P2_U3863 , P2_U3864 , P2_U3865 , P2_U3866 , P2_U3867 , P2_U3868 , P2_U3869 , P2_U3870;
wire P2_U3871 , P2_U3872 , P2_U3873 , P2_U3874 , P2_U3875 , P2_U3876 , P2_U3877 , P2_U3878 , P2_U3879 , P2_U3880;
wire P2_U3881 , P2_U3882 , P2_U3883 , P2_U3884 , P2_U3885 , P2_U3886 , P2_U3887 , P2_U3888 , P2_U3889 , P2_U3890;
wire P2_U3891 , P2_U3892 , P2_U3893 , P2_U3894 , P2_U3895 , P2_U3896 , P2_U3897 , P2_U3898 , P2_U3899 , P2_U3900;
wire P2_U3901 , P2_U3902 , P2_U3903 , P2_U3904 , P2_U3905 , P2_U3906 , P2_U3907 , P2_U3908 , P2_U3909 , P2_U3910;
wire P2_U3911 , P2_U3912 , P2_U3913 , P2_U3914 , P2_U3915 , P2_U3916 , P2_U3917 , P2_U3918 , P2_U3919 , P2_U3920;
wire P2_U3921 , P2_U3922 , P2_U3923 , P2_U3924 , P2_U3925 , P2_U3926 , P2_U3927 , P2_U3928 , P2_U3929 , P2_U3930;
wire P2_U3931 , P2_U3932 , P2_U3933 , P2_U3934 , P2_U3935 , P2_U3936 , P2_U3937 , P2_U3938 , P2_U3939 , P2_U3940;
wire P2_U3941 , P2_U3942 , P2_U3943 , P2_U3944 , P2_U3945 , P2_U3946 , P2_U3947 , P2_U3948 , P2_U3949 , P2_U3950;
wire P2_U3951 , P2_U3952 , P2_U3953 , P2_U3954 , P2_U3955 , P2_U3956 , P2_U3957 , P2_U3958 , P2_U3959 , P2_U3960;
wire P2_U3961 , P2_U3962 , P2_U3963 , P2_U3964 , P2_U3965 , P2_U3967 , P2_U3968 , P2_U3969 , P2_U3970 , P2_U3971;
wire P2_U3972 , P2_U3973 , P2_U3974 , P2_U3975 , P2_U3976 , P2_U3977 , P2_U3978 , P2_U3979 , P2_U3980 , P2_U3981;
wire P2_U3982 , P2_U3983 , P2_U3984 , P2_U3985 , P2_U3986 , P2_U3987 , P2_U3988 , P2_U3989 , P2_U3990 , P2_U3991;
wire P2_U3992 , P2_U3993 , P2_U3994 , P2_U3995 , P2_U3996 , P2_U3997 , P2_U3998 , P2_U3999 , P2_U4000 , P2_U4001;
wire P2_U4002 , P2_U4003 , P2_U4004 , P2_U4005 , P2_U4006 , P2_U4007 , P2_U4008 , P2_U4009 , P2_U4010 , P2_U4011;
wire P2_U4012 , P2_U4013 , P2_U4014 , P2_U4015 , P2_U4016 , P2_U4017 , P2_U4018 , P2_U4019 , P2_U4020 , P2_U4021;
wire P2_U4022 , P2_U4023 , P2_U4024 , P2_U4025 , P2_U4026 , P2_U4027 , P2_U4028 , P2_U4029 , P2_U4030 , P2_U4031;
wire P2_U4032 , P2_U4033 , P2_U4034 , P2_U4035 , P2_U4036 , P2_U4037 , P2_U4038 , P2_U4039 , P2_U4040 , P2_U4041;
wire P2_U4042 , P2_U4043 , P2_U4044 , P2_U4045 , P2_U4046 , P2_U4047 , P2_U4048 , P2_U4049 , P2_U4050 , P2_U4051;
wire P2_U4052 , P2_U4053 , P2_U4054 , P2_U4055 , P2_U4056 , P2_U4057 , P2_U4058 , P2_U4059 , P2_U4060 , P2_U4061;
wire P2_U4062 , P2_U4063 , P2_U4064 , P2_U4065 , P2_U4066 , P2_U4067 , P2_U4068 , P2_U4069 , P2_U4070 , P2_U4071;
wire P2_U4072 , P2_U4073 , P2_U4074 , P2_U4075 , P2_U4076 , P2_U4077 , P2_U4078 , P2_U4079 , P2_U4080 , P2_U4081;
wire P2_U4082 , P2_U4083 , P2_U4084 , P2_U4085 , P2_U4086 , P2_U4087 , P2_U4088 , P2_U4089 , P2_U4090 , P2_U4091;
wire P2_U4092 , P2_U4093 , P2_U4094 , P2_U4095 , P2_U4096 , P2_U4097 , P2_U4098 , P2_U4099 , P2_U4100 , P2_U4101;
wire P2_U4102 , P2_U4103 , P2_U4104 , P2_U4105 , P2_U4106 , P2_U4107 , P2_U4108 , P2_U4109 , P2_U4110 , P2_U4111;
wire P2_U4112 , P2_U4113 , P2_U4114 , P2_U4115 , P2_U4116 , P2_U4117 , P2_U4118 , P2_U4119 , P2_U4120 , P2_U4121;
wire P2_U4122 , P2_U4123 , P2_U4124 , P2_U4125 , P2_U4126 , P2_U4127 , P2_U4128 , P2_U4129 , P2_U4130 , P2_U4131;
wire P2_U4132 , P2_U4133 , P2_U4134 , P2_U4135 , P2_U4136 , P2_U4137 , P2_U4138 , P2_U4139 , P2_U4140 , P2_U4141;
wire P2_U4142 , P2_U4143 , P2_U4144 , P2_U4145 , P2_U4146 , P2_U4147 , P2_U4148 , P2_U4149 , P2_U4150 , P2_U4151;
wire P2_U4152 , P2_U4153 , P2_U4154 , P2_U4155 , P2_U4156 , P2_U4157 , P2_U4158 , P2_U4159 , P2_U4160 , P2_U4161;
wire P2_U4162 , P2_U4163 , P2_U4164 , P2_U4165 , P2_U4166 , P2_U4167 , P2_U4168 , P2_U4169 , P2_U4170 , P2_U4171;
wire P2_U4172 , P2_U4173 , P2_U4174 , P2_U4175 , P2_U4176 , P2_U4177 , P2_U4178 , P2_U4179 , P2_U4180 , P2_U4181;
wire P2_U4182 , P2_U4183 , P2_U4184 , P2_U4185 , P2_U4186 , P2_U4187 , P2_U4188 , P2_U4189 , P2_U4190 , P2_U4191;
wire P2_U4192 , P2_U4193 , P2_U4194 , P2_U4195 , P2_U4196 , P2_U4197 , P2_U4198 , P2_U4199 , P2_U4200 , P2_U4201;
wire P2_U4202 , P2_U4203 , P2_U4204 , P2_U4205 , P2_U4206 , P2_U4207 , P2_U4208 , P2_U4209 , P2_U4210 , P2_U4211;
wire P2_U4212 , P2_U4213 , P2_U4214 , P2_U4215 , P2_U4216 , P2_U4217 , P2_U4218 , P2_U4219 , P2_U4220 , P2_U4221;
wire P2_U4222 , P2_U4223 , P2_U4224 , P2_U4225 , P2_U4226 , P2_U4227 , P2_U4228 , P2_U4229 , P2_U4230 , P2_U4231;
wire P2_U4232 , P2_U4233 , P2_U4234 , P2_U4235 , P2_U4236 , P2_U4237 , P2_U4238 , P2_U4239 , P2_U4240 , P2_U4241;
wire P2_U4242 , P2_U4243 , P2_U4244 , P2_U4245 , P2_U4246 , P2_U4247 , P2_U4248 , P2_U4249 , P2_U4250 , P2_U4251;
wire P2_U4252 , P2_U4253 , P2_U4254 , P2_U4255 , P2_U4256 , P2_U4257 , P2_U4258 , P2_U4259 , P2_U4260 , P2_U4261;
wire P2_U4262 , P2_U4263 , P2_U4264 , P2_U4265 , P2_U4266 , P2_U4267 , P2_U4268 , P2_U4269 , P2_U4270 , P2_U4271;
wire P2_U4272 , P2_U4273 , P2_U4274 , P2_U4275 , P2_U4276 , P2_U4277 , P2_U4278 , P2_U4279 , P2_U4280 , P2_U4281;
wire P2_U4282 , P2_U4283 , P2_U4284 , P2_U4285 , P2_U4286 , P2_U4287 , P2_U4288 , P2_U4289 , P2_U4290 , P2_U4291;
wire P2_U4292 , P2_U4293 , P2_U4294 , P2_U4295 , P2_U4296 , P2_U4297 , P2_U4298 , P2_U4299 , P2_U4300 , P2_U4301;
wire P2_U4302 , P2_U4303 , P2_U4304 , P2_U4305 , P2_U4306 , P2_U4307 , P2_U4308 , P2_U4309 , P2_U4310 , P2_U4311;
wire P2_U4312 , P2_U4313 , P2_U4314 , P2_U4315 , P2_U4316 , P2_U4317 , P2_U4318 , P2_U4319 , P2_U4320 , P2_U4321;
wire P2_U4322 , P2_U4323 , P2_U4324 , P2_U4325 , P2_U4326 , P2_U4327 , P2_U4328 , P2_U4329 , P2_U4330 , P2_U4331;
wire P2_U4332 , P2_U4333 , P2_U4334 , P2_U4335 , P2_U4336 , P2_U4337 , P2_U4338 , P2_U4339 , P2_U4340 , P2_U4341;
wire P2_U4342 , P2_U4343 , P2_U4344 , P2_U4345 , P2_U4346 , P2_U4347 , P2_U4348 , P2_U4349 , P2_U4350 , P2_U4351;
wire P2_U4352 , P2_U4353 , P2_U4354 , P2_U4355 , P2_U4356 , P2_U4357 , P2_U4358 , P2_U4359 , P2_U4360 , P2_U4361;
wire P2_U4362 , P2_U4363 , P2_U4364 , P2_U4365 , P2_U4366 , P2_U4367 , P2_U4368 , P2_U4369 , P2_U4370 , P2_U4371;
wire P2_U4372 , P2_U4373 , P2_U4374 , P2_U4375 , P2_U4376 , P2_U4377 , P2_U4378 , P2_U4379 , P2_U4380 , P2_U4381;
wire P2_U4382 , P2_U4383 , P2_U4384 , P2_U4385 , P2_U4386 , P2_U4387 , P2_U4388 , P2_U4389 , P2_U4390 , P2_U4391;
wire P2_U4392 , P2_U4393 , P2_U4394 , P2_U4395 , P2_U4396 , P2_U4397 , P2_U4398 , P2_U4399 , P2_U4400 , P2_U4401;
wire P2_U4402 , P2_U4403 , P2_U4404 , P2_U4405 , P2_U4406 , P2_U4407 , P2_U4408 , P2_U4409 , P2_U4410 , P2_U4411;
wire P2_U4412 , P2_U4413 , P2_U4414 , P2_U4415 , P2_U4416 , P2_U4417 , P2_U4418 , P2_U4419 , P2_U4420 , P2_U4421;
wire P2_U4422 , P2_U4423 , P2_U4424 , P2_U4425 , P2_U4426 , P2_U4427 , P2_U4428 , P2_U4429 , P2_U4430 , P2_U4431;
wire P2_U4432 , P2_U4433 , P2_U4434 , P2_U4435 , P2_U4436 , P2_U4437 , P2_U4438 , P2_U4439 , P2_U4440 , P2_U4441;
wire P2_U4442 , P2_U4443 , P2_U4444 , P2_U4445 , P2_U4446 , P2_U4447 , P2_U4448 , P2_U4449 , P2_U4450 , P2_U4451;
wire P2_U4452 , P2_U4453 , P2_U4454 , P2_U4455 , P2_U4456 , P2_U4457 , P2_U4458 , P2_U4459 , P2_U4460 , P2_U4461;
wire P2_U4462 , P2_U4463 , P2_U4464 , P2_U4465 , P2_U4466 , P2_U4467 , P2_U4468 , P2_U4469 , P2_U4470 , P2_U4471;
wire P2_U4472 , P2_U4473 , P2_U4474 , P2_U4475 , P2_U4476 , P2_U4477 , P2_U4478 , P2_U4479 , P2_U4480 , P2_U4481;
wire P2_U4482 , P2_U4483 , P2_U4484 , P2_U4485 , P2_U4486 , P2_U4487 , P2_U4488 , P2_U4489 , P2_U4490 , P2_U4491;
wire P2_U4492 , P2_U4493 , P2_U4494 , P2_U4495 , P2_U4496 , P2_U4497 , P2_U4498 , P2_U4499 , P2_U4500 , P2_U4501;
wire P2_U4502 , P2_U4503 , P2_U4504 , P2_U4505 , P2_U4506 , P2_U4507 , P2_U4508 , P2_U4509 , P2_U4510 , P2_U4511;
wire P2_U4512 , P2_U4513 , P2_U4514 , P2_U4515 , P2_U4516 , P2_U4517 , P2_U4518 , P2_U4519 , P2_U4520 , P2_U4521;
wire P2_U4522 , P2_U4523 , P2_U4524 , P2_U4525 , P2_U4526 , P2_U4527 , P2_U4528 , P2_U4529 , P2_U4530 , P2_U4531;
wire P2_U4532 , P2_U4533 , P2_U4534 , P2_U4535 , P2_U4536 , P2_U4537 , P2_U4538 , P2_U4539 , P2_U4540 , P2_U4541;
wire P2_U4542 , P2_U4543 , P2_U4544 , P2_U4545 , P2_U4546 , P2_U4547 , P2_U4548 , P2_U4549 , P2_U4550 , P2_U4551;
wire P2_U4552 , P2_U4553 , P2_U4554 , P2_U4555 , P2_U4556 , P2_U4557 , P2_U4558 , P2_U4559 , P2_U4560 , P2_U4561;
wire P2_U4562 , P2_U4563 , P2_U4564 , P2_U4565 , P2_U4566 , P2_U4567 , P2_U4568 , P2_U4569 , P2_U4570 , P2_U4571;
wire P2_U4572 , P2_U4573 , P2_U4574 , P2_U4575 , P2_U4576 , P2_U4577 , P2_U4578 , P2_U4579 , P2_U4580 , P2_U4581;
wire P2_U4582 , P2_U4583 , P2_U4584 , P2_U4585 , P2_U4586 , P2_U4587 , P2_U4588 , P2_U4589 , P2_U4590 , P2_U4591;
wire P2_U4592 , P2_U4593 , P2_U4594 , P2_U4595 , P2_U4596 , P2_U4597 , P2_U4598 , P2_U4599 , P2_U4600 , P2_U4601;
wire P2_U4602 , P2_U4603 , P2_U4604 , P2_U4605 , P2_U4606 , P2_U4607 , P2_U4608 , P2_U4609 , P2_U4610 , P2_U4611;
wire P2_U4612 , P2_U4613 , P2_U4614 , P2_U4615 , P2_U4616 , P2_U4617 , P2_U4618 , P2_U4619 , P2_U4620 , P2_U4621;
wire P2_U4622 , P2_U4623 , P2_U4624 , P2_U4625 , P2_U4626 , P2_U4627 , P2_U4628 , P2_U4629 , P2_U4630 , P2_U4631;
wire P2_U4632 , P2_U4633 , P2_U4634 , P2_U4635 , P2_U4636 , P2_U4637 , P2_U4638 , P2_U4639 , P2_U4640 , P2_U4641;
wire P2_U4642 , P2_U4643 , P2_U4644 , P2_U4645 , P2_U4646 , P2_U4647 , P2_U4648 , P2_U4649 , P2_U4650 , P2_U4651;
wire P2_U4652 , P2_U4653 , P2_U4654 , P2_U4655 , P2_U4656 , P2_U4657 , P2_U4658 , P2_U4659 , P2_U4660 , P2_U4661;
wire P2_U4662 , P2_U4663 , P2_U4664 , P2_U4665 , P2_U4666 , P2_U4667 , P2_U4668 , P2_U4669 , P2_U4670 , P2_U4671;
wire P2_U4672 , P2_U4673 , P2_U4674 , P2_U4675 , P2_U4676 , P2_U4677 , P2_U4678 , P2_U4679 , P2_U4680 , P2_U4681;
wire P2_U4682 , P2_U4683 , P2_U4684 , P2_U4685 , P2_U4686 , P2_U4687 , P2_U4688 , P2_U4689 , P2_U4690 , P2_U4691;
wire P2_U4692 , P2_U4693 , P2_U4694 , P2_U4695 , P2_U4696 , P2_U4697 , P2_U4698 , P2_U4699 , P2_U4700 , P2_U4701;
wire P2_U4702 , P2_U4703 , P2_U4704 , P2_U4705 , P2_U4706 , P2_U4707 , P2_U4708 , P2_U4709 , P2_U4710 , P2_U4711;
wire P2_U4712 , P2_U4713 , P2_U4714 , P2_U4715 , P2_U4716 , P2_U4717 , P2_U4718 , P2_U4719 , P2_U4720 , P2_U4721;
wire P2_U4722 , P2_U4723 , P2_U4724 , P2_U4725 , P2_U4726 , P2_U4727 , P2_U4728 , P2_U4729 , P2_U4730 , P2_U4731;
wire P2_U4732 , P2_U4733 , P2_U4734 , P2_U4735 , P2_U4736 , P2_U4737 , P2_U4738 , P2_U4739 , P2_U4740 , P2_U4741;
wire P2_U4742 , P2_U4743 , P2_U4744 , P2_U4745 , P2_U4746 , P2_U4747 , P2_U4748 , P2_U4749 , P2_U4750 , P2_U4751;
wire P2_U4752 , P2_U4753 , P2_U4754 , P2_U4755 , P2_U4756 , P2_U4757 , P2_U4758 , P2_U4759 , P2_U4760 , P2_U4761;
wire P2_U4762 , P2_U4763 , P2_U4764 , P2_U4765 , P2_U4766 , P2_U4767 , P2_U4768 , P2_U4769 , P2_U4770 , P2_U4771;
wire P2_U4772 , P2_U4773 , P2_U4774 , P2_U4775 , P2_U4776 , P2_U4777 , P2_U4778 , P2_U4779 , P2_U4780 , P2_U4781;
wire P2_U4782 , P2_U4783 , P2_U4784 , P2_U4785 , P2_U4786 , P2_U4787 , P2_U4788 , P2_U4789 , P2_U4790 , P2_U4791;
wire P2_U4792 , P2_U4793 , P2_U4794 , P2_U4795 , P2_U4796 , P2_U4797 , P2_U4798 , P2_U4799 , P2_U4800 , P2_U4801;
wire P2_U4802 , P2_U4803 , P2_U4804 , P2_U4805 , P2_U4806 , P2_U4807 , P2_U4808 , P2_U4809 , P2_U4810 , P2_U4811;
wire P2_U4812 , P2_U4813 , P2_U4814 , P2_U4815 , P2_U4816 , P2_U4817 , P2_U4818 , P2_U4819 , P2_U4820 , P2_U4821;
wire P2_U4822 , P2_U4823 , P2_U4824 , P2_U4825 , P2_U4826 , P2_U4827 , P2_U4828 , P2_U4829 , P2_U4830 , P2_U4831;
wire P2_U4832 , P2_U4833 , P2_U4834 , P2_U4835 , P2_U4836 , P2_U4837 , P2_U4838 , P2_U4839 , P2_U4840 , P2_U4841;
wire P2_U4842 , P2_U4843 , P2_U4844 , P2_U4845 , P2_U4846 , P2_U4847 , P2_U4848 , P2_U4849 , P2_U4850 , P2_U4851;
wire P2_U4852 , P2_U4853 , P2_U4854 , P2_U4855 , P2_U4856 , P2_U4857 , P2_U4858 , P2_U4859 , P2_U4860 , P2_U4861;
wire P2_U4862 , P2_U4863 , P2_U4864 , P2_U4865 , P2_U4866 , P2_U4867 , P2_U4868 , P2_U4869 , P2_U4870 , P2_U4871;
wire P2_U4872 , P2_U4873 , P2_U4874 , P2_U4875 , P2_U4876 , P2_U4877 , P2_U4878 , P2_U4879 , P2_U4880 , P2_U4881;
wire P2_U4882 , P2_U4883 , P2_U4884 , P2_U4885 , P2_U4886 , P2_U4887 , P2_U4888 , P2_U4889 , P2_U4890 , P2_U4891;
wire P2_U4892 , P2_U4893 , P2_U4894 , P2_U4895 , P2_U4896 , P2_U4897 , P2_U4898 , P2_U4899 , P2_U4900 , P2_U4901;
wire P2_U4902 , P2_U4903 , P2_U4904 , P2_U4905 , P2_U4906 , P2_U4907 , P2_U4908 , P2_U4909 , P2_U4910 , P2_U4911;
wire P2_U4912 , P2_U4913 , P2_U4914 , P2_U4915 , P2_U4916 , P2_U4917 , P2_U4918 , P2_U4919 , P2_U4920 , P2_U4921;
wire P2_U4922 , P2_U4923 , P2_U4924 , P2_U4925 , P2_U4926 , P2_U4927 , P2_U4928 , P2_U4929 , P2_U4930 , P2_U4931;
wire P2_U4932 , P2_U4933 , P2_U4934 , P2_U4935 , P2_U4936 , P2_U4937 , P2_U4938 , P2_U4939 , P2_U4940 , P2_U4941;
wire P2_U4942 , P2_U4943 , P2_U4944 , P2_U4945 , P2_U4946 , P2_U4947 , P2_U4948 , P2_U4949 , P2_U4950 , P2_U4951;
wire P2_U4952 , P2_U4953 , P2_U4954 , P2_U4955 , P2_U4956 , P2_U4957 , P2_U4958 , P2_U4959 , P2_U4960 , P2_U4961;
wire P2_U4962 , P2_U4963 , P2_U4964 , P2_U4965 , P2_U4966 , P2_U4967 , P2_U4968 , P2_U4969 , P2_U4970 , P2_U4971;
wire P2_U4972 , P2_U4973 , P2_U4974 , P2_U4975 , P2_U4976 , P2_U4977 , P2_U4978 , P2_U4979 , P2_U4980 , P2_U4981;
wire P2_U4982 , P2_U4983 , P2_U4984 , P2_U4985 , P2_U4986 , P2_U4987 , P2_U4988 , P2_U4989 , P2_U4990 , P2_U4991;
wire P2_U4992 , P2_U4993 , P2_U4994 , P2_U4995 , P2_U4996 , P2_U4997 , P2_U4998 , P2_U4999 , P2_U5000 , P2_U5001;
wire P2_U5002 , P2_U5003 , P2_U5004 , P2_U5005 , P2_U5006 , P2_U5007 , P2_U5008 , P2_U5009 , P2_U5010 , P2_U5011;
wire P2_U5012 , P2_U5013 , P2_U5014 , P2_U5015 , P2_U5016 , P2_U5017 , P2_U5018 , P2_U5019 , P2_U5020 , P2_U5021;
wire P2_U5022 , P2_U5023 , P2_U5024 , P2_U5025 , P2_U5026 , P2_U5027 , P2_U5028 , P2_U5029 , P2_U5030 , P2_U5031;
wire P2_U5032 , P2_U5033 , P2_U5034 , P2_U5035 , P2_U5036 , P2_U5037 , P2_U5038 , P2_U5039 , P2_U5040 , P2_U5041;
wire P2_U5042 , P2_U5043 , P2_U5044 , P2_U5045 , P2_U5046 , P2_U5047 , P2_U5048 , P2_U5049 , P2_U5050 , P2_U5051;
wire P2_U5052 , P2_U5053 , P2_U5054 , P2_U5055 , P2_U5056 , P2_U5057 , P2_U5058 , P2_U5059 , P2_U5060 , P2_U5061;
wire P2_U5062 , P2_U5063 , P2_U5064 , P2_U5065 , P2_U5066 , P2_U5067 , P2_U5068 , P2_U5069 , P2_U5070 , P2_U5071;
wire P2_U5072 , P2_U5073 , P2_U5074 , P2_U5075 , P2_U5076 , P2_U5077 , P2_U5078 , P2_U5079 , P2_U5080 , P2_U5081;
wire P2_U5082 , P2_U5083 , P2_U5084 , P2_U5085 , P2_U5086 , P2_U5087 , P2_U5088 , P2_U5089 , P2_U5090 , P2_U5091;
wire P2_U5092 , P2_U5093 , P2_U5094 , P2_U5095 , P2_U5096 , P2_U5097 , P2_U5098 , P2_U5099 , P2_U5100 , P2_U5101;
wire P2_U5102 , P2_U5103 , P2_U5104 , P2_U5105 , P2_U5106 , P2_U5107 , P2_U5108 , P2_U5109 , P2_U5110 , P2_U5111;
wire P2_U5112 , P2_U5113 , P2_U5114 , P2_U5115 , P2_U5116 , P2_U5117 , P2_U5118 , P2_U5119 , P2_U5120 , P2_U5121;
wire P2_U5122 , P2_U5123 , P2_U5124 , P2_U5125 , P2_U5126 , P2_U5127 , P2_U5128 , P2_U5129 , P2_U5130 , P2_U5131;
wire P2_U5132 , P2_U5133 , P2_U5134 , P2_U5135 , P2_U5136 , P2_U5137 , P2_U5138 , P2_U5139 , P2_U5140 , P2_U5141;
wire P2_U5142 , P2_U5143 , P2_U5144 , P2_U5145 , P2_U5146 , P2_U5147 , P2_U5148 , P2_U5149 , P2_U5150 , P2_U5151;
wire P2_U5152 , P2_U5153 , P2_U5154 , P2_U5155 , P2_U5156 , P2_U5157 , P2_U5158 , P2_U5159 , P2_U5160 , P2_U5161;
wire P2_U5162 , P2_U5163 , P2_U5164 , P2_U5165 , P2_U5166 , P2_U5167 , P2_U5168 , P2_U5169 , P2_U5170 , P2_U5171;
wire P2_U5172 , P2_U5173 , P2_U5174 , P2_U5175 , P2_U5176 , P2_U5177 , P2_U5178 , P2_U5179 , P2_U5180 , P2_U5181;
wire P2_U5182 , P2_U5183 , P2_U5184 , P2_U5185 , P2_U5186 , P2_U5187 , P2_U5188 , P2_U5189 , P2_U5190 , P2_U5191;
wire P2_U5192 , P2_U5193 , P2_U5194 , P2_U5195 , P2_U5196 , P2_U5197 , P2_U5198 , P2_U5199 , P2_U5200 , P2_U5201;
wire P2_U5202 , P2_U5203 , P2_U5204 , P2_U5205 , P2_U5206 , P2_U5207 , P2_U5208 , P2_U5209 , P2_U5210 , P2_U5211;
wire P2_U5212 , P2_U5213 , P2_U5214 , P2_U5215 , P2_U5216 , P2_U5217 , P2_U5218 , P2_U5219 , P2_U5220 , P2_U5221;
wire P2_U5222 , P2_U5223 , P2_U5224 , P2_U5225 , P2_U5226 , P2_U5227 , P2_U5228 , P2_U5229 , P2_U5230 , P2_U5231;
wire P2_U5232 , P2_U5233 , P2_U5234 , P2_U5235 , P2_U5236 , P2_U5237 , P2_U5238 , P2_U5239 , P2_U5240 , P2_U5241;
wire P2_U5242 , P2_U5243 , P2_U5244 , P2_U5245 , P2_U5246 , P2_U5247 , P2_U5248 , P2_U5249 , P2_U5250 , P2_U5251;
wire P2_U5252 , P2_U5253 , P2_U5254 , P2_U5255 , P2_U5256 , P2_U5257 , P2_U5258 , P2_U5259 , P2_U5260 , P2_U5261;
wire P2_U5262 , P2_U5263 , P2_U5264 , P2_U5265 , P2_U5266 , P2_U5267 , P2_U5268 , P2_U5269 , P2_U5270 , P2_U5271;
wire P2_U5272 , P2_U5273 , P2_U5274 , P2_U5275 , P2_U5276 , P2_U5277 , P2_U5278 , P2_U5279 , P2_U5280 , P2_U5281;
wire P2_U5282 , P2_U5283 , P2_U5284 , P2_U5285 , P2_U5286 , P2_U5287 , P2_U5288 , P2_U5289 , P2_U5290 , P2_U5291;
wire P2_U5292 , P2_U5293 , P2_U5294 , P2_U5295 , P2_U5296 , P2_U5297 , P2_U5298 , P2_U5299 , P2_U5300 , P2_U5301;
wire P2_U5302 , P2_U5303 , P2_U5304 , P2_U5305 , P2_U5306 , P2_U5307 , P2_U5308 , P2_U5309 , P2_U5310 , P2_U5311;
wire P2_U5312 , P2_U5313 , P2_U5314 , P2_U5315 , P2_U5316 , P2_U5317 , P2_U5318 , P2_U5319 , P2_U5320 , P2_U5321;
wire P2_U5322 , P2_U5323 , P2_U5324 , P2_U5325 , P2_U5326 , P2_U5327 , P2_U5328 , P2_U5329 , P2_U5330 , P2_U5331;
wire P2_U5332 , P2_U5333 , P2_U5334 , P2_U5335 , P2_U5336 , P2_U5337 , P2_U5338 , P2_U5339 , P2_U5340 , P2_U5341;
wire P2_U5342 , P2_U5343 , P2_U5344 , P2_U5345 , P2_U5346 , P2_U5347 , P2_U5348 , P2_U5349 , P2_U5350 , P2_U5351;
wire P2_U5352 , P2_U5353 , P2_U5354 , P2_U5355 , P2_U5356 , P2_U5357 , P2_U5358 , P2_U5359 , P2_U5360 , P2_U5361;
wire P2_U5362 , P2_U5363 , P2_U5364 , P2_U5365 , P2_U5366 , P2_U5367 , P2_U5368 , P2_U5369 , P2_U5370 , P2_U5371;
wire P2_U5372 , P2_U5373 , P2_U5374 , P2_U5375 , P2_U5376 , P2_U5377 , P2_U5378 , P2_U5379 , P2_U5380 , P2_U5381;
wire P2_U5382 , P2_U5383 , P2_U5384 , P2_U5385 , P2_U5386 , P2_U5387 , P2_U5388 , P2_U5389 , P2_U5390 , P2_U5391;
wire P2_U5392 , P2_U5393 , P2_U5394 , P2_U5395 , P2_U5396 , P2_U5397 , P2_U5398 , P2_U5399 , P2_U5400 , P2_U5401;
wire P2_U5402 , P2_U5403 , P2_U5404 , P2_U5405 , P2_U5406 , P2_U5407 , P2_U5408 , P2_U5409 , P2_U5410 , P2_U5411;
wire P2_U5412 , P2_U5413 , P2_U5414 , P2_U5415 , P2_U5416 , P2_U5417 , P2_U5418 , P2_U5419 , P2_U5420 , P2_U5421;
wire P2_U5422 , P2_U5423 , P2_U5424 , P2_U5425 , P2_U5426 , P2_U5427 , P2_U5428 , P2_U5429 , P2_U5430 , P2_U5431;
wire P2_U5432 , P2_U5433 , P2_U5434 , P2_U5435 , P2_U5436 , P2_U5437 , P2_U5438 , P2_U5439 , P2_U5440 , P2_U5441;
wire P2_U5442 , P2_U5443 , P2_U5444 , P2_U5445 , P2_U5446 , P2_U5447 , P2_U5448 , P2_U5449 , P2_U5450 , P2_U5451;
wire P2_U5452 , P2_U5453 , P2_U5454 , P2_U5455 , P2_U5456 , P2_U5457 , P2_U5458 , P2_U5459 , P2_U5460 , P2_U5461;
wire P2_U5462 , P2_U5463 , P2_U5464 , P2_U5465 , P2_U5466 , P2_U5467 , P2_U5468 , P2_U5469 , P2_U5470 , P2_U5471;
wire P2_U5472 , P2_U5473 , P2_U5474 , P2_U5475 , P2_U5476 , P2_U5477 , P2_U5478 , P2_U5479 , P2_U5480 , P2_U5481;
wire P2_U5482 , P2_U5483 , P2_U5484 , P2_U5485 , P2_U5486 , P2_U5487 , P2_U5488 , P2_U5489 , P2_U5490 , P2_U5491;
wire P2_U5492 , P2_U5493 , P2_U5494 , P2_U5495 , P2_U5496 , P2_U5497 , P2_U5498 , P2_U5499 , P2_U5500 , P2_U5501;
wire P2_U5502 , P2_U5503 , P2_U5504 , P2_U5505 , P2_U5506 , P2_U5507 , P2_U5508 , P2_U5509 , P2_U5510 , P2_U5511;
wire P2_U5512 , P2_U5513 , P2_U5514 , P2_U5515 , P2_U5516 , P2_U5517 , P2_U5518 , P2_U5519 , P2_U5520 , P2_U5521;
wire P2_U5522 , P2_U5523 , P2_U5524 , P2_U5525 , P2_U5526 , P2_U5527 , P2_U5528 , P2_U5529 , P2_U5530 , P2_U5531;
wire P2_U5532 , P2_U5533 , P2_U5534 , P2_U5535 , P2_U5536 , P2_U5537 , P2_U5538 , P2_U5539 , P2_U5540 , P2_U5541;
wire P2_U5542 , P2_U5543 , P2_U5544 , P2_U5545 , P2_U5546 , P2_U5547 , P2_U5548 , P2_U5549 , P2_U5550 , P2_U5551;
wire P2_U5552 , P2_U5553 , P2_U5554 , P2_U5555 , P2_U5556 , P2_U5557 , P2_U5558 , P2_U5559 , P2_U5560 , P2_U5561;
wire P2_U5562 , P2_U5563 , P2_U5564 , P2_U5565 , P2_U5566 , P2_U5567 , P2_U5568 , P2_U5569 , P2_U5570 , P2_U5571;
wire P2_U5572 , P2_U5573 , P2_U5574 , P2_U5575 , P2_U5576 , P2_U5577 , P2_U5578 , P2_U5579 , P2_U5580 , P2_U5581;
wire P2_U5582 , P2_U5583 , P2_U5584 , P2_U5585 , P2_U5586 , P2_U5587 , P2_U5588 , P2_U5589 , P2_U5590 , P2_U5591;
wire P2_U5592 , P2_U5593 , P2_U5594 , P2_U5595 , P2_U5596 , P2_U5597 , P2_U5598 , P2_U5599 , P2_U5600 , P2_U5601;
wire P2_U5602 , P2_U5603 , P2_U5604 , P2_U5605 , P2_U5606 , P2_U5607 , P2_U5608 , P2_U5609 , P2_U5610 , P2_U5611;
wire P2_U5612 , P2_U5613 , P2_U5614 , P2_U5615 , P2_U5616 , P2_U5617 , P2_U5618 , P2_U5619 , P2_U5620 , P2_U5621;
wire P2_U5622 , P2_U5623 , P2_U5624 , P2_U5625 , P2_U5626 , P2_U5627 , P2_U5628 , P2_U5629 , P2_U5630 , P2_U5631;
wire P2_U5632 , P2_U5633 , P2_U5634 , P2_U5635 , P2_U5636 , P2_U5637 , P2_U5638 , P2_U5639 , P2_U5640 , P2_U5641;
wire P2_U5642 , P2_U5643 , P2_U5644 , P2_U5645 , P2_U5646 , P2_U5647 , P2_U5648 , P2_U5649 , P2_U5650 , P2_U5651;
wire P2_U5652 , P2_U5653 , P2_U5654 , P2_U5655 , P2_U5656 , P2_U5657 , P2_U5658 , P2_U5659 , P2_U5660 , P2_U5661;
wire P2_U5662 , P2_U5663 , P2_U5664 , P2_U5665 , P2_U5666 , P2_U5667 , P2_U5668 , P2_U5669 , P2_U5670 , P2_U5671;
wire P2_U5672 , P2_U5673 , P2_U5674 , P2_U5675 , P2_U5676 , P2_U5677 , P2_U5678 , P2_U5679 , P2_U5680 , P2_U5681;
wire P2_U5682 , P2_U5683 , P2_U5684 , P2_U5685 , P2_U5686 , P2_U5687 , P2_U5688 , P2_U5689 , P2_U5690 , P2_U5691;
wire P2_U5692 , P2_U5693 , P2_U5694 , P2_U5695 , P2_U5696 , P2_U5697 , P2_U5698 , P2_U5699 , P2_U5700 , P2_U5701;
wire P2_U5702 , P2_U5703 , P2_U5704 , P2_U5705 , P2_U5706 , P2_U5707 , P2_U5708 , P2_U5709 , P2_U5710 , P2_U5711;
wire P2_U5712 , P2_U5713 , P2_U5714 , P2_U5715 , P2_U5716 , P2_U5717 , P2_U5718 , P2_U5719 , P2_U5720 , P2_U5721;
wire P2_U5722 , P2_U5723 , P2_U5724 , P2_U5725 , P2_U5726 , P2_U5727 , P2_U5728 , P2_U5729 , P2_U5730 , P2_U5731;
wire P2_U5732 , P2_U5733 , P2_U5734 , P2_U5735 , P2_U5736 , P2_U5737 , P2_U5738 , P2_U5739 , P2_U5740 , P2_U5741;
wire P2_U5742 , P2_U5743 , P2_U5744 , P2_U5745 , P2_U5746 , P2_U5747 , P2_U5748 , P2_U5749 , P2_U5750 , P2_U5751;
wire P2_U5752 , P2_U5753 , P2_U5754 , P2_U5755 , P2_U5756 , P2_U5757 , P2_U5758 , P2_U5759 , P2_U5760 , P2_U5761;
wire P2_U5762 , P2_U5763 , P2_U5764 , P2_U5765 , P2_U5766 , P2_U5767 , P2_U5768 , P2_U5769 , P2_U5770 , P2_U5771;
wire P2_U5772 , P2_U5773 , P2_U5774 , P2_U5775 , P2_U5776 , P2_U5777 , P2_U5778 , P2_U5779 , P2_U5780 , P2_U5781;
wire P2_U5782 , P2_U5783 , P2_U5784 , P2_U5785 , P2_U5786 , P2_U5787 , P2_U5788 , P2_U5789 , P2_U5790 , P2_U5791;
wire P2_U5792 , P2_U5793 , P2_U5794 , P2_U5795 , P2_U5796 , P2_U5797 , P2_U5798 , P2_U5799 , P2_U5800 , P2_U5801;
wire P2_U5802 , P2_U5803 , P2_U5804 , P2_U5805 , P2_U5806 , P2_U5807 , P2_U5808 , P2_U5809 , P2_U5810 , P2_U5811;
wire P2_U5812 , P2_U5813 , P2_U5814 , P2_U5815 , P2_U5816 , P2_U5817 , P2_U5818 , P2_U5819 , P2_U5820 , P2_U5821;
wire P2_U5822 , P2_U5823 , P2_U5824 , P2_U5825 , P2_U5826 , P2_U5827 , P2_U5828 , P2_U5829 , P2_U5830 , P2_U5831;
wire P2_U5832 , P2_U5833 , P2_U5834 , P2_U5835 , P2_U5836 , P2_U5837 , P2_U5838 , P2_U5839 , P2_U5840 , P2_U5841;
wire P2_U5842 , P2_U5843 , P2_U5844 , P2_U5845 , P2_U5846 , P2_U5847 , P2_U5848 , P2_U5849 , P2_U5850 , P2_U5851;
wire P2_U5852 , P2_U5853 , P2_U5854 , P2_U5855 , P2_U5856 , P2_U5857 , P2_U5858 , P2_U5859 , P2_U5860 , P2_U5861;
wire P2_U5862 , P2_U5863 , P2_U5864 , P2_U5865 , P2_U5866 , P2_U5867 , P2_U5868 , P2_U5869 , P2_U5870 , P2_U5871;
wire P2_U5872 , P2_U5873 , P2_U5874 , P2_U5875 , P2_U5876 , P2_U5877 , P2_U5878 , P2_U5879 , P2_U5880 , P2_U5881;
wire P2_U5882 , P2_U5883 , P2_U5884 , P2_U5885 , P2_U5886 , P2_U5887 , P2_U5888 , P2_U5889 , P2_U5890 , P2_U5891;
wire P2_U5892 , P2_U5893 , P2_U5894 , P2_U5895 , P2_U5896 , P2_U5897 , P2_U5898 , P2_U5899 , P2_U5900 , P2_U5901;
wire P2_U5902 , P2_U5903 , P2_U5904 , P2_U5905 , P2_U5906 , P2_U5907 , P2_U5908 , P2_U5909 , P2_U5910 , P2_U5911;
wire P2_U5912 , P2_U5913 , P2_U5914 , P2_U5915 , P2_U5916 , P2_U5917 , P2_U5918 , P2_U5919 , P2_U5920 , P2_U5921;
wire P2_U5922 , P2_U5923 , P2_U5924 , P2_U5925 , P2_U5926 , P2_U5927 , P2_U5928 , P2_U5929 , P2_U5930 , P2_U5931;
wire P2_U5932 , P2_U5933 , P2_U5934 , P2_U5935 , P2_U5936 , P2_U5937 , P2_U5938 , P2_U5939 , P2_U5940 , P2_U5941;
wire P2_U5942 , P2_U5943 , P2_U5944 , P2_U5945 , P2_U5946 , P2_U5947 , P2_U5948 , P2_U5949 , P2_U5950 , P2_U5951;
wire P2_U5952 , P2_U5953 , P2_U5954 , P2_U5955 , P2_U5956 , P2_U5957 , P2_U5958 , P2_U5959 , P2_U5960 , P2_U5961;
wire P2_U5962 , P2_U5963 , P2_U5964 , P2_U5965 , P2_U5966 , P2_U5967 , P2_U5968 , P2_U5969 , P2_U5970 , P2_U5971;
wire P2_U5972 , P2_U5973 , P2_U5974 , P2_U5975 , P2_U5976 , P2_U5977 , P2_U5978 , P2_U5979 , P2_U5980 , P2_U5981;
wire P2_U5982 , P2_U5983 , P2_U5984 , P2_U5985 , P2_U5986 , P2_U5987 , P2_U5988 , P2_U5989 , P2_U5990 , P2_U5991;
wire P2_U5992 , P2_U5993 , P2_U5994 , P2_U5995 , P2_U5996 , P2_U5997 , P2_U5998 , P2_U5999 , P2_U6000 , P2_U6001;
wire P2_U6002 , P2_U6003 , P2_U6004 , P2_U6005 , P2_U6006 , P2_U6007 , P2_U6008 , P2_U6009 , P2_U6010 , P2_U6011;
wire P2_U6012 , P2_U6013 , P2_U6014 , P2_U6015 , P2_U6016 , P2_U6017 , P2_U6018 , P2_U6019 , P2_U6020 , P2_U6021;
wire P2_U6022 , P2_U6023 , P2_U6024 , P2_U6025 , P2_U6026 , P2_U6027 , P2_U6028 , P2_U6029 , P2_U6030 , P2_U6031;
wire P2_U6032 , P2_U6033 , P2_U6034 , P2_U6035 , P2_U6036 , P2_U6037 , P2_U6038 , P2_U6039 , P2_U6040 , P2_U6041;
wire P2_U6042 , P2_U6043 , P2_U6044 , P2_U6045 , P2_U6046 , P2_U6047 , P2_U6048 , P2_U6049 , P2_U6050 , P2_U6051;
wire P2_U6052 , P2_U6053 , P2_U6054 , P2_U6055 , P2_U6056 , P2_U6057 , P2_U6058 , P2_U6059 , P2_U6060 , P2_U6061;
wire P2_U6062 , P2_U6063 , P2_U6064 , P2_U6065 , P2_U6066 , P2_U6067 , P2_U6068 , P2_U6069 , P2_U6070 , P2_U6071;
wire P2_U6072 , P2_U6073 , P2_U6074 , P2_U6075 , P2_U6076 , P2_U6077 , P2_U6078 , P2_U6079 , P2_U6080 , P2_U6081;
wire P2_U6082 , P2_U6083 , P2_U6084 , P2_U6085 , P2_U6086 , P2_U6087 , P2_U6088 , P2_U6089 , P2_U6090 , P2_U6091;
wire P2_U6092 , P2_U6093 , P2_U6094 , P2_U6095 , P2_U6096 , P2_U6097 , P2_U6098 , P2_U6099 , P2_U6100 , P2_U6101;
wire P2_U6102 , P2_U6103 , P2_U6104 , P2_U6105 , P2_U6106 , P2_U6107 , P2_U6108 , P2_U6109 , P2_U6110 , P2_U6111;
wire P2_U6112 , P2_U6113 , P2_U6114 , P2_U6115 , P2_U6116 , P2_U6117 , P2_U6118 , P2_U6119 , P2_U6120 , P2_U6121;
wire P2_U6122 , P2_U6123 , P2_U6124 , P2_U6125 , P2_U6126 , P2_U6127 , P2_U6128 , P2_U6129 , P2_U6130 , P2_U6131;
wire P2_U6132 , P2_U6133 , P2_U6134 , P2_U6135 , P2_U6136 , P2_U6137 , P2_U6138 , P2_U6139 , P2_U6140 , P2_U6141;
wire P2_U6142 , P2_U6143 , P2_U6144 , P2_U6145 , P2_U6146 , P2_U6147 , P2_U6148 , P2_U6149 , P2_U6150 , P2_U6151;
wire P2_U6152 , P2_U6153 , P2_U6154 , P2_U6155 , P2_U6156 , P2_U6157 , P2_U6158 , P2_U6159 , P2_U6160 , P2_U6161;
wire P2_U6162 , P2_U6163 , P2_U6164 , P2_U6165 , P2_U6166 , P2_U6167 , P2_U6168 , P2_U6169 , P2_U6170 , P2_U6171;
wire P2_U6172 , P2_U6173 , P2_U6174 , P2_U6175 , P2_U6176 , P2_U6177 , P2_U6178 , P2_U6179 , P2_U6180 , P2_U6181;
wire P2_U6182 , P2_U6183 , P2_U6184 , P2_U6185 , P2_U6186 , P2_U6187 , P2_U6188 , P2_U6189 , P2_U6190 , P2_U6191;
wire P2_U6192 , P2_U6193 , P2_U6194 , P2_U6195 , P2_U6196 , P2_U6197 , P2_U6198 , P2_U6199 , P2_U6200 , P2_U6201;
wire P2_U6202 , P2_U6203 , P2_U6204 , P2_U6205 , P2_U6206 , P2_U6207 , P2_U6208 , P2_U6209 , P2_U6210 , P2_U6211;
wire P2_U6212 , P2_U6213 , P2_U6214 , P2_U6215 , P2_U6216 , P2_U6217 , P2_U6218 , P2_U6219 , P2_U6220 , P2_U6221;
wire P2_U6222 , P2_U6223 , P2_U6224 , P2_U6225 , P2_U6226 , P2_U6227 , P2_U6228 , P2_U6229 , P2_U6230 , P2_U6231;
wire P2_U6232 , P2_U6233 , P2_U6234 , P2_U6235 , P2_U6236 , P2_U6237 , P2_U6238 , P2_U6239 , P2_U6240 , P2_U6241;
wire P2_U6242 , P2_U6243 , P2_U6244 , P2_U6245 , P2_U6246 , P2_U6247 , P2_U6248 , P2_U6249 , P2_U6250 , P2_U6251;
wire P2_U6252 , P2_U6253 , P2_U6254 , P2_U6255 , P2_U6256 , P2_U6257 , P2_U6258 , P2_U6259 , P2_U6260 , P2_U6261;
wire P2_U6262 , P2_U6263 , P2_U6264 , P2_U6265 , P2_U6266 , P2_U6267 , P2_U6268 , P2_U6269 , P2_U6270 , P2_R1113_U438;
wire P2_R1113_U437 , P2_R1113_U436 , P2_R1113_U435 , P2_R1113_U434 , P2_R1113_U433 , P2_R1113_U432 , P2_R1113_U431 , P2_R1113_U430 , P2_R1113_U429 , P2_R1113_U428;
wire P2_R1113_U427 , P2_R1113_U426 , P2_R1113_U425 , P2_R1113_U424 , P2_R1113_U423 , P2_R1113_U422 , P2_R1113_U421 , P2_R1113_U420 , P2_R1113_U419 , LT_1079_U6;
wire ADD_1071_U6 , ADD_1071_U7 , ADD_1071_U8 , ADD_1071_U9 , ADD_1071_U10 , ADD_1071_U11 , ADD_1071_U12 , ADD_1071_U13 , ADD_1071_U14 , ADD_1071_U15;
wire ADD_1071_U16 , ADD_1071_U17 , ADD_1071_U18 , ADD_1071_U19 , ADD_1071_U20 , ADD_1071_U21 , ADD_1071_U22 , ADD_1071_U23 , ADD_1071_U24 , ADD_1071_U25;
wire ADD_1071_U26 , ADD_1071_U27 , ADD_1071_U28 , ADD_1071_U29 , ADD_1071_U30 , ADD_1071_U31 , ADD_1071_U32 , ADD_1071_U33 , ADD_1071_U34 , ADD_1071_U35;
wire ADD_1071_U36 , ADD_1071_U37 , ADD_1071_U38 , ADD_1071_U39 , ADD_1071_U40 , ADD_1071_U41 , ADD_1071_U42 , ADD_1071_U43 , ADD_1071_U44 , ADD_1071_U45;
wire ADD_1071_U64 , ADD_1071_U65 , ADD_1071_U66 , ADD_1071_U67 , ADD_1071_U68 , ADD_1071_U69 , ADD_1071_U70 , ADD_1071_U71 , ADD_1071_U72 , ADD_1071_U73;
wire ADD_1071_U74 , ADD_1071_U75 , ADD_1071_U76 , ADD_1071_U77 , ADD_1071_U78 , ADD_1071_U79 , ADD_1071_U80 , ADD_1071_U81 , ADD_1071_U82 , ADD_1071_U83;
wire ADD_1071_U84 , ADD_1071_U85 , ADD_1071_U86 , ADD_1071_U87 , ADD_1071_U88 , ADD_1071_U89 , ADD_1071_U90 , ADD_1071_U91 , ADD_1071_U92 , ADD_1071_U93;
wire ADD_1071_U94 , ADD_1071_U95 , ADD_1071_U96 , ADD_1071_U97 , ADD_1071_U98 , ADD_1071_U99 , ADD_1071_U100 , ADD_1071_U101 , ADD_1071_U102 , ADD_1071_U103;
wire ADD_1071_U104 , ADD_1071_U105 , ADD_1071_U106 , ADD_1071_U107 , ADD_1071_U108 , ADD_1071_U109 , ADD_1071_U110 , ADD_1071_U111 , ADD_1071_U112 , ADD_1071_U113;
wire ADD_1071_U114 , ADD_1071_U115 , ADD_1071_U116 , ADD_1071_U117 , ADD_1071_U118 , ADD_1071_U119 , ADD_1071_U120 , ADD_1071_U121 , ADD_1071_U122 , ADD_1071_U123;
wire ADD_1071_U124 , ADD_1071_U125 , ADD_1071_U126 , ADD_1071_U127 , ADD_1071_U128 , ADD_1071_U129 , ADD_1071_U130 , ADD_1071_U131 , ADD_1071_U132 , ADD_1071_U133;
wire ADD_1071_U134 , ADD_1071_U135 , ADD_1071_U136 , ADD_1071_U137 , ADD_1071_U138 , ADD_1071_U139 , ADD_1071_U140 , ADD_1071_U141 , ADD_1071_U142 , ADD_1071_U143;
wire ADD_1071_U144 , ADD_1071_U145 , ADD_1071_U146 , ADD_1071_U147 , ADD_1071_U148 , ADD_1071_U149 , ADD_1071_U150 , ADD_1071_U151 , ADD_1071_U152 , ADD_1071_U153;
wire ADD_1071_U154 , ADD_1071_U155 , ADD_1071_U156 , ADD_1071_U157 , ADD_1071_U158 , ADD_1071_U159 , ADD_1071_U160 , ADD_1071_U161 , ADD_1071_U162 , ADD_1071_U163;
wire ADD_1071_U164 , ADD_1071_U165 , ADD_1071_U166 , ADD_1071_U167 , ADD_1071_U168 , ADD_1071_U169 , ADD_1071_U170 , ADD_1071_U171 , ADD_1071_U172 , ADD_1071_U173;
wire ADD_1071_U174 , ADD_1071_U175 , ADD_1071_U176 , ADD_1071_U177 , ADD_1071_U178 , ADD_1071_U179 , ADD_1071_U180 , ADD_1071_U181 , ADD_1071_U182 , ADD_1071_U183;
wire ADD_1071_U184 , ADD_1071_U185 , ADD_1071_U186 , ADD_1071_U187 , ADD_1071_U188 , ADD_1071_U189 , ADD_1071_U190 , ADD_1071_U191 , ADD_1071_U192 , ADD_1071_U193;
wire ADD_1071_U194 , ADD_1071_U195 , ADD_1071_U196 , ADD_1071_U197 , ADD_1071_U198 , ADD_1071_U199 , ADD_1071_U200 , ADD_1071_U201 , ADD_1071_U202 , ADD_1071_U203;
wire ADD_1071_U204 , ADD_1071_U205 , ADD_1071_U206 , ADD_1071_U207 , ADD_1071_U208 , ADD_1071_U209 , ADD_1071_U210 , ADD_1071_U211 , ADD_1071_U212 , ADD_1071_U213;
wire ADD_1071_U214 , ADD_1071_U215 , ADD_1071_U216 , ADD_1071_U217 , ADD_1071_U218 , ADD_1071_U219 , ADD_1071_U220 , ADD_1071_U221 , ADD_1071_U222 , ADD_1071_U223;
wire ADD_1071_U224 , ADD_1071_U225 , ADD_1071_U226 , ADD_1071_U227 , ADD_1071_U228 , ADD_1071_U229 , ADD_1071_U230 , ADD_1071_U231 , ADD_1071_U232 , ADD_1071_U233;
wire ADD_1071_U234 , ADD_1071_U235 , ADD_1071_U236 , ADD_1071_U237 , ADD_1071_U238 , ADD_1071_U239 , ADD_1071_U240 , ADD_1071_U241 , ADD_1071_U242 , ADD_1071_U243;
wire ADD_1071_U244 , ADD_1071_U245 , ADD_1071_U246 , ADD_1071_U247 , ADD_1071_U248 , ADD_1071_U249 , ADD_1071_U250 , ADD_1071_U251 , ADD_1071_U252 , ADD_1071_U253;
wire ADD_1071_U254 , ADD_1071_U255 , ADD_1071_U256 , ADD_1071_U257 , ADD_1071_U258 , ADD_1071_U259 , ADD_1071_U260 , ADD_1071_U261 , ADD_1071_U262 , ADD_1071_U263;
wire ADD_1071_U264 , ADD_1071_U265 , ADD_1071_U266 , ADD_1071_U267 , ADD_1071_U268 , ADD_1071_U269 , ADD_1071_U270 , ADD_1071_U271 , ADD_1071_U272 , ADD_1071_U273;
wire ADD_1071_U274 , ADD_1071_U275 , ADD_1071_U276 , ADD_1071_U277 , ADD_1071_U278 , ADD_1071_U279 , ADD_1071_U280 , ADD_1071_U281 , ADD_1071_U282 , ADD_1071_U283;
wire ADD_1071_U284 , ADD_1071_U285 , ADD_1071_U286 , ADD_1071_U287 , ADD_1071_U288 , ADD_1071_U289 , ADD_1071_U290 , ADD_1071_U291 , R140_U4 , R140_U5;
wire R140_U6 , R140_U7 , R140_U8 , R140_U9 , R140_U10 , R140_U11 , R140_U12 , R140_U13 , R140_U14 , R140_U15;
wire R140_U16 , R140_U17 , R140_U18 , R140_U19 , R140_U20 , R140_U21 , R140_U22 , R140_U23 , R140_U24 , R140_U25;
wire R140_U26 , R140_U27 , R140_U28 , R140_U29 , R140_U30 , R140_U31 , R140_U32 , R140_U33 , R140_U34 , R140_U35;
wire R140_U36 , R140_U37 , R140_U38 , R140_U39 , R140_U40 , R140_U41 , R140_U42 , R140_U43 , R140_U44 , R140_U45;
wire R140_U46 , R140_U47 , R140_U48 , R140_U49 , R140_U50 , R140_U51 , R140_U52 , R140_U53 , R140_U54 , R140_U55;
wire R140_U56 , R140_U57 , R140_U58 , R140_U59 , R140_U60 , R140_U61 , R140_U62 , R140_U63 , R140_U64 , R140_U65;
wire R140_U66 , R140_U67 , R140_U68 , R140_U69 , R140_U70 , R140_U71 , R140_U72 , R140_U73 , R140_U74 , R140_U75;
wire R140_U76 , R140_U77 , R140_U78 , R140_U79 , R140_U80 , R140_U81 , R140_U82 , R140_U83 , R140_U84 , R140_U85;
wire R140_U86 , R140_U87 , R140_U88 , R140_U89 , R140_U90 , R140_U91 , R140_U92 , R140_U93 , R140_U94 , R140_U95;
wire R140_U96 , R140_U97 , R140_U98 , R140_U99 , R140_U100 , R140_U101 , R140_U102 , R140_U103 , R140_U104 , R140_U105;
wire R140_U106 , R140_U107 , R140_U108 , R140_U109 , R140_U110 , R140_U111 , R140_U112 , R140_U113 , R140_U114 , R140_U115;
wire R140_U116 , R140_U117 , R140_U118 , R140_U119 , R140_U120 , R140_U121 , R140_U122 , R140_U123 , R140_U124 , R140_U125;
wire R140_U126 , R140_U127 , R140_U128 , R140_U129 , R140_U130 , R140_U131 , R140_U132 , R140_U133 , R140_U134 , R140_U135;
wire R140_U136 , R140_U137 , R140_U138 , R140_U139 , R140_U140 , R140_U141 , R140_U142 , R140_U143 , R140_U144 , R140_U145;
wire R140_U146 , R140_U147 , R140_U148 , R140_U149 , R140_U150 , R140_U151 , R140_U152 , R140_U153 , R140_U154 , R140_U155;
wire R140_U156 , R140_U157 , R140_U158 , R140_U159 , R140_U160 , R140_U161 , R140_U162 , R140_U163 , R140_U164 , R140_U165;
wire R140_U166 , R140_U167 , R140_U168 , R140_U169 , R140_U170 , R140_U171 , R140_U172 , R140_U173 , R140_U174 , R140_U175;
wire R140_U176 , R140_U177 , R140_U178 , R140_U179 , R140_U180 , R140_U181 , R140_U182 , R140_U183 , R140_U184 , R140_U185;
wire R140_U186 , R140_U187 , R140_U188 , R140_U189 , R140_U190 , R140_U191 , R140_U192 , R140_U193 , R140_U194 , R140_U195;
wire R140_U196 , R140_U197 , R140_U198 , R140_U199 , R140_U200 , R140_U201 , R140_U202 , R140_U203 , R140_U204 , R140_U205;
wire R140_U206 , R140_U207 , R140_U208 , R140_U209 , R140_U210 , R140_U211 , R140_U212 , R140_U213 , R140_U214 , R140_U215;
wire R140_U216 , R140_U217 , R140_U218 , R140_U219 , R140_U220 , R140_U221 , R140_U222 , R140_U223 , R140_U224 , R140_U225;
wire R140_U226 , R140_U227 , R140_U228 , R140_U229 , R140_U230 , R140_U231 , R140_U232 , R140_U233 , R140_U234 , R140_U235;
wire R140_U236 , R140_U237 , R140_U238 , R140_U239 , R140_U240 , R140_U241 , R140_U242 , R140_U243 , R140_U244 , R140_U245;
wire R140_U246 , R140_U247 , R140_U248 , R140_U249 , R140_U250 , R140_U251 , R140_U252 , R140_U253 , R140_U254 , R140_U255;
wire R140_U256 , R140_U257 , R140_U258 , R140_U259 , R140_U260 , R140_U261 , R140_U262 , R140_U263 , R140_U264 , R140_U265;
wire R140_U266 , R140_U267 , R140_U268 , R140_U269 , R140_U270 , R140_U271 , R140_U272 , R140_U273 , R140_U274 , R140_U275;
wire R140_U276 , R140_U277 , R140_U278 , R140_U279 , R140_U280 , R140_U281 , R140_U282 , R140_U283 , R140_U284 , R140_U285;
wire R140_U286 , R140_U287 , R140_U288 , R140_U289 , R140_U290 , R140_U291 , R140_U292 , R140_U293 , R140_U294 , R140_U295;
wire R140_U296 , R140_U297 , R140_U298 , R140_U299 , R140_U300 , R140_U301 , R140_U302 , R140_U303 , R140_U304 , R140_U305;
wire R140_U306 , R140_U307 , R140_U308 , R140_U309 , R140_U310 , R140_U311 , R140_U312 , R140_U313 , R140_U314 , R140_U315;
wire R140_U316 , R140_U317 , R140_U318 , R140_U319 , R140_U320 , R140_U321 , R140_U322 , R140_U323 , R140_U324 , R140_U325;
wire R140_U326 , R140_U327 , R140_U328 , R140_U329 , R140_U330 , R140_U331 , R140_U332 , R140_U333 , R140_U334 , R140_U335;
wire R140_U336 , R140_U337 , R140_U338 , R140_U339 , R140_U340 , R140_U341 , R140_U342 , R140_U343 , R140_U344 , R140_U345;
wire R140_U346 , R140_U347 , R140_U348 , R140_U349 , R140_U350 , R140_U351 , R140_U352 , R140_U353 , R140_U354 , R140_U355;
wire R140_U356 , R140_U357 , R140_U358 , R140_U359 , R140_U360 , R140_U361 , R140_U362 , R140_U363 , R140_U364 , R140_U365;
wire R140_U366 , R140_U367 , R140_U368 , R140_U369 , R140_U370 , R140_U371 , R140_U372 , R140_U373 , R140_U374 , R140_U375;
wire R140_U376 , R140_U377 , R140_U378 , R140_U379 , R140_U380 , R140_U381 , R140_U382 , R140_U383 , R140_U384 , R140_U385;
wire R140_U386 , R140_U387 , R140_U388 , R140_U389 , R140_U390 , R140_U391 , R140_U392 , R140_U393 , R140_U394 , R140_U395;
wire R140_U396 , R140_U397 , R140_U398 , R140_U399 , R140_U400 , R140_U401 , R140_U402 , R140_U403 , R140_U404 , R140_U405;
wire R140_U406 , R140_U407 , R140_U408 , R140_U409 , R140_U410 , R140_U411 , R140_U412 , R140_U413 , R140_U414 , R140_U415;
wire R140_U416 , R140_U417 , R140_U418 , R140_U419 , R140_U420 , R140_U421 , R140_U422 , R140_U423 , R140_U424 , R140_U425;
wire R140_U426 , R140_U427 , R140_U428 , R140_U429 , R140_U430 , R140_U431 , R140_U432 , R140_U433 , R140_U434 , R140_U435;
wire R140_U436 , R140_U437 , R140_U438 , R140_U439 , R140_U440 , R140_U441 , R140_U442 , R140_U443 , R140_U444 , R140_U445;
wire R140_U446 , R140_U447 , R140_U448 , R140_U449 , R140_U450 , R140_U451 , R140_U452 , R140_U453 , R140_U454 , R140_U455;
wire R140_U456 , R140_U457 , R140_U458 , R140_U459 , R140_U460 , R140_U461 , R140_U462 , R140_U463 , R140_U464 , R140_U465;
wire R140_U466 , R140_U467 , R140_U468 , R140_U469 , R140_U470 , R140_U471 , R140_U472 , R140_U473 , R140_U474 , R140_U475;
wire R140_U476 , R140_U477 , R140_U478 , R140_U479 , R140_U480 , R140_U481 , R140_U482 , R140_U483 , R140_U484 , R140_U485;
wire R140_U486 , R140_U487 , R140_U488 , R140_U489 , R140_U490 , R140_U491 , R140_U492 , R140_U493 , R140_U494 , R140_U495;
wire R140_U496 , R140_U497 , R140_U498 , R140_U499 , R140_U500 , R140_U501 , R140_U502 , R140_U503 , R140_U504 , R140_U505;
wire R140_U506 , R140_U507 , R140_U508 , R140_U509 , R140_U510 , R140_U511 , R140_U512 , R140_U513 , R140_U514 , R140_U515;
wire R140_U516 , R140_U517 , R140_U518 , R140_U519 , R140_U520 , R140_U521 , R140_U522 , R140_U523 , R140_U524 , R140_U525;
wire R140_U526 , R140_U527 , R140_U528 , R140_U529 , R140_U530 , R140_U531 , R140_U532 , R140_U533 , R140_U534 , R140_U535;
wire R140_U536 , R140_U537 , R140_U538 , R140_U539 , R140_U540 , R140_U541 , LT_1079_19_U6 , P1_ADD_99_U4 , P1_ADD_99_U5 , P1_ADD_99_U6;
wire P1_ADD_99_U7 , P1_ADD_99_U8 , P1_ADD_99_U9 , P1_ADD_99_U10 , P1_ADD_99_U11 , P1_ADD_99_U12 , P1_ADD_99_U13 , P1_ADD_99_U14 , P1_ADD_99_U15 , P1_ADD_99_U16;
wire P1_ADD_99_U17 , P1_ADD_99_U18 , P1_ADD_99_U19 , P1_ADD_99_U20 , P1_ADD_99_U21 , P1_ADD_99_U22 , P1_ADD_99_U23 , P1_ADD_99_U24 , P1_ADD_99_U25 , P1_ADD_99_U26;
wire P1_ADD_99_U27 , P1_ADD_99_U28 , P1_ADD_99_U29 , P1_ADD_99_U30 , P1_ADD_99_U31 , P1_ADD_99_U32 , P1_ADD_99_U33 , P1_ADD_99_U34 , P1_ADD_99_U35 , P1_ADD_99_U36;
wire P1_ADD_99_U37 , P1_ADD_99_U38 , P1_ADD_99_U39 , P1_ADD_99_U40 , P1_ADD_99_U41 , P1_ADD_99_U42 , P1_ADD_99_U43 , P1_ADD_99_U44 , P1_ADD_99_U45 , P1_ADD_99_U46;
wire P1_ADD_99_U47 , P1_ADD_99_U48 , P1_ADD_99_U49 , P1_ADD_99_U50 , P1_ADD_99_U51 , P1_ADD_99_U52 , P1_ADD_99_U53 , P1_ADD_99_U54 , P1_ADD_99_U55 , P1_ADD_99_U56;
wire P1_ADD_99_U57 , P1_ADD_99_U58 , P1_ADD_99_U59 , P1_ADD_99_U60 , P1_ADD_99_U61 , P1_ADD_99_U62 , P1_ADD_99_U63 , P1_ADD_99_U64 , P1_ADD_99_U65 , P1_ADD_99_U66;
wire P1_ADD_99_U67 , P1_ADD_99_U68 , P1_ADD_99_U69 , P1_ADD_99_U70 , P1_ADD_99_U71 , P1_ADD_99_U72 , P1_ADD_99_U73 , P1_ADD_99_U74 , P1_ADD_99_U75 , P1_ADD_99_U76;
wire P1_ADD_99_U77 , P1_ADD_99_U78 , P1_ADD_99_U79 , P1_ADD_99_U80 , P1_ADD_99_U81 , P1_ADD_99_U82 , P1_ADD_99_U83 , P1_ADD_99_U84 , P1_ADD_99_U85 , P1_ADD_99_U86;
wire P1_ADD_99_U87 , P1_ADD_99_U88 , P1_ADD_99_U89 , P1_ADD_99_U90 , P1_ADD_99_U91 , P1_ADD_99_U92 , P1_ADD_99_U93 , P1_ADD_99_U94 , P1_ADD_99_U95 , P1_ADD_99_U96;
wire P1_ADD_99_U97 , P1_ADD_99_U98 , P1_ADD_99_U99 , P1_ADD_99_U100 , P1_ADD_99_U101 , P1_ADD_99_U102 , P1_ADD_99_U103 , P1_ADD_99_U104 , P1_ADD_99_U105 , P1_ADD_99_U106;
wire P1_ADD_99_U107 , P1_ADD_99_U108 , P1_ADD_99_U109 , P1_ADD_99_U110 , P1_ADD_99_U111 , P1_ADD_99_U112 , P1_ADD_99_U113 , P1_ADD_99_U114 , P1_ADD_99_U115 , P1_ADD_99_U116;
wire P1_ADD_99_U117 , P1_ADD_99_U118 , P1_ADD_99_U119 , P1_ADD_99_U120 , P1_ADD_99_U121 , P1_ADD_99_U122 , P1_ADD_99_U123 , P1_ADD_99_U124 , P1_ADD_99_U125 , P1_ADD_99_U126;
wire P1_ADD_99_U127 , P1_ADD_99_U128 , P1_ADD_99_U129 , P1_ADD_99_U130 , P1_ADD_99_U131 , P1_ADD_99_U132 , P1_ADD_99_U133 , P1_ADD_99_U134 , P1_ADD_99_U135 , P1_ADD_99_U136;
wire P1_ADD_99_U137 , P1_ADD_99_U138 , P1_ADD_99_U139 , P1_ADD_99_U140 , P1_ADD_99_U141 , P1_ADD_99_U142 , P1_ADD_99_U143 , P1_ADD_99_U144 , P1_ADD_99_U145 , P1_ADD_99_U146;
wire P1_ADD_99_U147 , P1_ADD_99_U148 , P1_ADD_99_U149 , P1_ADD_99_U150 , P1_ADD_99_U151 , P1_ADD_99_U152 , P1_ADD_99_U153 , P1_R1105_U4 , P1_R1105_U5 , P1_R1105_U6;
wire P1_R1105_U7 , P1_R1105_U8 , P1_R1105_U9 , P1_R1105_U10 , P1_R1105_U11 , P1_R1105_U12 , P1_R1105_U13 , P1_R1105_U14 , P1_R1105_U15 , P1_R1105_U16;
wire P1_R1105_U17 , P1_R1105_U18 , P1_R1105_U19 , P1_R1105_U20 , P1_R1105_U21 , P1_R1105_U22 , P1_R1105_U23 , P1_R1105_U24 , P1_R1105_U25 , P1_R1105_U26;
wire P1_R1105_U27 , P1_R1105_U28 , P1_R1105_U29 , P1_R1105_U30 , P1_R1105_U31 , P1_R1105_U32 , P1_R1105_U33 , P1_R1105_U34 , P1_R1105_U35 , P1_R1105_U36;
wire P1_R1105_U37 , P1_R1105_U38 , P1_R1105_U39 , P1_R1105_U40 , P1_R1105_U41 , P1_R1105_U42 , P1_R1105_U43 , P1_R1105_U44 , P1_R1105_U45 , P1_R1105_U46;
wire P1_R1105_U47 , P1_R1105_U48 , P1_R1105_U49 , P1_R1105_U50 , P1_R1105_U51 , P1_R1105_U52 , P1_R1105_U53 , P1_R1105_U54 , P1_R1105_U55 , P1_R1105_U56;
wire P1_R1105_U57 , P1_R1105_U58 , P1_R1105_U59 , P1_R1105_U60 , P1_R1105_U61 , P1_R1105_U62 , P1_R1105_U63 , P1_R1105_U64 , P1_R1105_U65 , P1_R1105_U66;
wire P1_R1105_U67 , P1_R1105_U68 , P1_R1105_U69 , P1_R1105_U70 , P1_R1105_U71 , P1_R1105_U72 , P1_R1105_U73 , P1_R1105_U74 , P1_R1105_U75 , P1_R1105_U76;
wire P1_R1105_U77 , P1_R1105_U78 , P1_R1105_U79 , P1_R1105_U80 , P1_R1105_U81 , P1_R1105_U82 , P1_R1105_U83 , P1_R1105_U84 , P1_R1105_U85 , P1_R1105_U86;
wire P1_R1105_U87 , P1_R1105_U88 , P1_R1105_U89 , P1_R1105_U90 , P1_R1105_U91 , P1_R1105_U92 , P1_R1105_U93 , P1_R1105_U94 , P1_R1105_U95 , P1_R1105_U96;
wire P1_R1105_U97 , P1_R1105_U98 , P1_R1105_U99 , P1_R1105_U100 , P1_R1105_U101 , P1_R1105_U102 , P1_R1105_U103 , P1_R1105_U104 , P1_R1105_U105 , P1_R1105_U106;
wire P1_R1105_U107 , P1_R1105_U108 , P1_R1105_U109 , P1_R1105_U110 , P1_R1105_U111 , P1_R1105_U112 , P1_R1105_U113 , P1_R1105_U114 , P1_R1105_U115 , P1_R1105_U116;
wire P1_R1105_U117 , P1_R1105_U118 , P1_R1105_U119 , P1_R1105_U120 , P1_R1105_U121 , P1_R1105_U122 , P1_R1105_U123 , P1_R1105_U124 , P1_R1105_U125 , P1_R1105_U126;
wire P1_R1105_U127 , P1_R1105_U128 , P1_R1105_U129 , P1_R1105_U130 , P1_R1105_U131 , P1_R1105_U132 , P1_R1105_U133 , P1_R1105_U134 , P1_R1105_U135 , P1_R1105_U136;
wire P1_R1105_U137 , P1_R1105_U138 , P1_R1105_U139 , P1_R1105_U140 , P1_R1105_U141 , P1_R1105_U142 , P1_R1105_U143 , P1_R1105_U144 , P1_R1105_U145 , P1_R1105_U146;
wire P1_R1105_U147 , P1_R1105_U148 , P1_R1105_U149 , P1_R1105_U150 , P1_R1105_U151 , P1_R1105_U152 , P1_R1105_U153 , P1_R1105_U154 , P1_R1105_U155 , P1_R1105_U156;
wire P1_R1105_U157 , P1_R1105_U158 , P1_R1105_U159 , P1_R1105_U160 , P1_R1105_U161 , P1_R1105_U162 , P1_R1105_U163 , P1_R1105_U164 , P1_R1105_U165 , P1_R1105_U166;
wire P1_R1105_U167 , P1_R1105_U168 , P1_R1105_U169 , P1_R1105_U170 , P1_R1105_U171 , P1_R1105_U172 , P1_R1105_U173 , P1_R1105_U174 , P1_R1105_U175 , P1_R1105_U176;
wire P1_R1105_U177 , P1_R1105_U178 , P1_R1105_U179 , P1_R1105_U180 , P1_R1105_U181 , P1_R1105_U182 , P1_R1105_U183 , P1_R1105_U184 , P1_R1105_U185 , P1_R1105_U186;
wire P1_R1105_U187 , P1_R1105_U188 , P1_R1105_U189 , P1_R1105_U190 , P1_R1105_U191 , P1_R1105_U192 , P1_R1105_U193 , P1_R1105_U194 , P1_R1105_U195 , P1_R1105_U196;
wire P1_R1105_U197 , P1_R1105_U198 , P1_R1105_U199 , P1_R1105_U200 , P1_R1105_U201 , P1_R1105_U202 , P1_R1105_U203 , P1_R1105_U204 , P1_R1105_U205 , P1_R1105_U206;
wire P1_R1105_U207 , P1_R1105_U208 , P1_R1105_U209 , P1_R1105_U210 , P1_R1105_U211 , P1_R1105_U212 , P1_R1105_U213 , P1_R1105_U214 , P1_R1105_U215 , P1_R1105_U216;
wire P1_R1105_U217 , P1_R1105_U218 , P1_R1105_U219 , P1_R1105_U220 , P1_R1105_U221 , P1_R1105_U222 , P1_R1105_U223 , P1_R1105_U224 , P1_R1105_U225 , P1_R1105_U226;
wire P1_R1105_U227 , P1_R1105_U228 , P1_R1105_U229 , P1_R1105_U230 , P1_R1105_U231 , P1_R1105_U232 , P1_R1105_U233 , P1_R1105_U234 , P1_R1105_U235 , P1_R1105_U236;
wire P1_R1105_U237 , P1_R1105_U238 , P1_R1105_U239 , P1_R1105_U240 , P1_R1105_U241 , P1_R1105_U242 , P1_R1105_U243 , P1_R1105_U244 , P1_R1105_U245 , P1_R1105_U246;
wire P1_R1105_U247 , P1_R1105_U248 , P1_R1105_U249 , P1_R1105_U250 , P1_R1105_U251 , P1_R1105_U252 , P1_R1105_U253 , P1_R1105_U254 , P1_R1105_U255 , P1_R1105_U256;
wire P1_R1105_U257 , P1_R1105_U258 , P1_R1105_U259 , P1_R1105_U260 , P1_R1105_U261 , P1_R1105_U262 , P1_R1105_U263 , P1_R1105_U264 , P1_R1105_U265 , P1_R1105_U266;
wire P1_R1105_U267 , P1_R1105_U268 , P1_R1105_U269 , P1_R1105_U270 , P1_R1105_U271 , P1_R1105_U272 , P1_R1105_U273 , P1_R1105_U274 , P1_R1105_U275 , P1_R1105_U276;
wire P1_R1105_U277 , P1_R1105_U278 , P1_R1105_U279 , P1_R1105_U280 , P1_R1105_U281 , P1_R1105_U282 , P1_R1105_U283 , P1_R1105_U284 , P1_R1105_U285 , P1_R1105_U286;
wire P1_R1105_U287 , P1_R1105_U288 , P1_R1105_U289 , P1_R1105_U290 , P1_R1105_U291 , P1_R1105_U292 , P1_R1105_U293 , P1_R1105_U294 , P1_R1105_U295 , P1_R1105_U296;
wire P1_R1105_U297 , P1_R1105_U298 , P1_R1105_U299 , P1_R1105_U300 , P1_R1105_U301 , P1_R1105_U302 , P1_R1105_U303 , P1_R1105_U304 , P1_R1105_U305 , P1_R1105_U306;
wire P1_R1105_U307 , P1_R1105_U308 , P1_SUB_88_U6 , P1_SUB_88_U7 , P1_SUB_88_U8 , P1_SUB_88_U9 , P1_SUB_88_U10 , P1_SUB_88_U11 , P1_SUB_88_U12 , P1_SUB_88_U13;
wire P1_SUB_88_U14 , P1_SUB_88_U15 , P1_SUB_88_U16 , P1_SUB_88_U17 , P1_SUB_88_U18 , P1_SUB_88_U19 , P1_SUB_88_U20 , P1_SUB_88_U21 , P1_SUB_88_U22 , P1_SUB_88_U23;
wire P1_SUB_88_U24 , P1_SUB_88_U25 , P1_SUB_88_U26 , P1_SUB_88_U27 , P1_SUB_88_U28 , P1_SUB_88_U29 , P1_SUB_88_U30 , P1_SUB_88_U31 , P1_SUB_88_U32 , P1_SUB_88_U33;
wire P1_SUB_88_U34 , P1_SUB_88_U35 , P1_SUB_88_U36 , P1_SUB_88_U37 , P1_SUB_88_U38 , P1_SUB_88_U39 , P1_SUB_88_U40 , P1_SUB_88_U41 , P1_SUB_88_U42 , P1_SUB_88_U43;
wire P1_SUB_88_U44 , P1_SUB_88_U45 , P1_SUB_88_U46 , P1_SUB_88_U47 , P1_SUB_88_U48 , P1_SUB_88_U49 , P1_SUB_88_U50 , P1_SUB_88_U51 , P1_SUB_88_U52 , P1_SUB_88_U53;
wire P1_SUB_88_U54 , P1_SUB_88_U55 , P1_SUB_88_U56 , P1_SUB_88_U57 , P1_SUB_88_U58 , P1_SUB_88_U59 , P1_SUB_88_U60 , P1_SUB_88_U61 , P1_SUB_88_U62 , P1_SUB_88_U63;
wire P1_SUB_88_U64 , P1_SUB_88_U65 , P1_SUB_88_U66 , P1_SUB_88_U67 , P1_SUB_88_U68 , P1_SUB_88_U69 , P1_SUB_88_U70 , P1_SUB_88_U71 , P1_SUB_88_U72 , P1_SUB_88_U73;
wire P1_SUB_88_U74 , P1_SUB_88_U75 , P1_SUB_88_U76 , P1_SUB_88_U77 , P1_SUB_88_U78 , P1_SUB_88_U79 , P1_SUB_88_U80 , P1_SUB_88_U81 , P1_SUB_88_U82 , P1_SUB_88_U83;
wire P1_SUB_88_U84 , P1_SUB_88_U85 , P1_SUB_88_U86 , P1_SUB_88_U87 , P1_SUB_88_U88 , P1_SUB_88_U89 , P1_SUB_88_U90 , P1_SUB_88_U91 , P1_SUB_88_U92 , P1_SUB_88_U93;
wire P1_SUB_88_U94 , P1_SUB_88_U95 , P1_SUB_88_U96 , P1_SUB_88_U97 , P1_SUB_88_U98 , P1_SUB_88_U99 , P1_SUB_88_U100 , P1_SUB_88_U101 , P1_SUB_88_U102 , P1_SUB_88_U103;
wire P1_SUB_88_U104 , P1_SUB_88_U105 , P1_SUB_88_U106 , P1_SUB_88_U107 , P1_SUB_88_U108 , P1_SUB_88_U109 , P1_SUB_88_U110 , P1_SUB_88_U111 , P1_SUB_88_U112 , P1_SUB_88_U113;
wire P1_SUB_88_U114 , P1_SUB_88_U115 , P1_SUB_88_U116 , P1_SUB_88_U117 , P1_SUB_88_U118 , P1_SUB_88_U119 , P1_SUB_88_U120 , P1_SUB_88_U121 , P1_SUB_88_U122 , P1_SUB_88_U123;
wire P1_SUB_88_U124 , P1_SUB_88_U125 , P1_SUB_88_U126 , P1_SUB_88_U127 , P1_SUB_88_U128 , P1_SUB_88_U129 , P1_SUB_88_U130 , P1_SUB_88_U131 , P1_SUB_88_U132 , P1_SUB_88_U133;
wire P1_SUB_88_U134 , P1_SUB_88_U135 , P1_SUB_88_U136 , P1_SUB_88_U137 , P1_SUB_88_U138 , P1_SUB_88_U139 , P1_SUB_88_U140 , P1_SUB_88_U141 , P1_SUB_88_U142 , P1_SUB_88_U143;
wire P1_SUB_88_U144 , P1_SUB_88_U145 , P1_SUB_88_U146 , P1_SUB_88_U147 , P1_SUB_88_U148 , P1_SUB_88_U149 , P1_SUB_88_U150 , P1_SUB_88_U151 , P1_SUB_88_U152 , P1_SUB_88_U153;
wire P1_SUB_88_U154 , P1_SUB_88_U155 , P1_SUB_88_U156 , P1_SUB_88_U157 , P1_SUB_88_U158 , P1_SUB_88_U159 , P1_SUB_88_U160 , P1_SUB_88_U161 , P1_SUB_88_U162 , P1_SUB_88_U163;
wire P1_SUB_88_U164 , P1_SUB_88_U165 , P1_SUB_88_U166 , P1_SUB_88_U167 , P1_SUB_88_U168 , P1_SUB_88_U169 , P1_SUB_88_U170 , P1_SUB_88_U171 , P1_SUB_88_U172 , P1_SUB_88_U173;
wire P1_SUB_88_U174 , P1_SUB_88_U175 , P1_SUB_88_U176 , P1_SUB_88_U177 , P1_SUB_88_U178 , P1_SUB_88_U179 , P1_SUB_88_U180 , P1_SUB_88_U181 , P1_SUB_88_U182 , P1_SUB_88_U183;
wire P1_SUB_88_U184 , P1_SUB_88_U185 , P1_SUB_88_U186 , P1_SUB_88_U187 , P1_SUB_88_U188 , P1_SUB_88_U189 , P1_SUB_88_U190 , P1_SUB_88_U191 , P1_SUB_88_U192 , P1_SUB_88_U193;
wire P1_SUB_88_U194 , P1_SUB_88_U195 , P1_SUB_88_U196 , P1_SUB_88_U197 , P1_SUB_88_U198 , P1_SUB_88_U199 , P1_SUB_88_U200 , P1_SUB_88_U201 , P1_SUB_88_U202 , P1_SUB_88_U203;
wire P1_SUB_88_U204 , P1_SUB_88_U205 , P1_SUB_88_U206 , P1_SUB_88_U207 , P1_SUB_88_U208 , P1_SUB_88_U209 , P1_SUB_88_U210 , P1_SUB_88_U211 , P1_SUB_88_U212 , P1_SUB_88_U213;
wire P1_SUB_88_U214 , P1_SUB_88_U215 , P1_SUB_88_U216 , P1_SUB_88_U217 , P1_SUB_88_U218 , P1_SUB_88_U219 , P1_SUB_88_U220 , P1_SUB_88_U221 , P1_SUB_88_U222 , P1_SUB_88_U223;
wire P1_SUB_88_U224 , P1_SUB_88_U225 , P1_SUB_88_U226 , P1_SUB_88_U227 , P1_SUB_88_U228 , P1_SUB_88_U229 , P1_SUB_88_U230 , P1_SUB_88_U231 , P1_SUB_88_U232 , P1_SUB_88_U233;
wire P1_SUB_88_U234 , P1_SUB_88_U235 , P1_SUB_88_U236 , P1_SUB_88_U237 , P1_SUB_88_U238 , P1_SUB_88_U239 , P1_SUB_88_U240 , P1_SUB_88_U241 , P1_SUB_88_U242 , P1_SUB_88_U243;
wire P1_SUB_88_U244 , P1_SUB_88_U245 , P1_SUB_88_U246 , P1_SUB_88_U247 , P1_SUB_88_U248 , P1_SUB_88_U249 , P1_SUB_88_U250 , P1_SUB_88_U251 , P1_R1309_U6 , P1_R1309_U7;
wire P1_R1309_U8 , P1_R1309_U9 , P1_R1309_U10 , P1_R1282_U6 , P1_R1282_U7 , P1_R1282_U8 , P1_R1282_U9 , P1_R1282_U10 , P1_R1282_U11 , P1_R1282_U12;
wire P1_R1282_U13 , P1_R1282_U14 , P1_R1282_U15 , P1_R1282_U16 , P1_R1282_U17 , P1_R1282_U18 , P1_R1282_U19 , P1_R1282_U20 , P1_R1282_U21 , P1_R1282_U22;
wire P1_R1282_U23 , P1_R1282_U24 , P1_R1282_U25 , P1_R1282_U26 , P1_R1282_U27 , P1_R1282_U28 , P1_R1282_U29 , P1_R1282_U30 , P1_R1282_U31 , P1_R1282_U32;
wire P1_R1282_U33 , P1_R1282_U34 , P1_R1282_U35 , P1_R1282_U36 , P1_R1282_U37 , P1_R1282_U38 , P1_R1282_U39 , P1_R1282_U40 , P1_R1282_U41 , P1_R1282_U42;
wire P1_R1282_U43 , P1_R1282_U44 , P1_R1282_U45 , P1_R1282_U46 , P1_R1282_U47 , P1_R1282_U48 , P1_R1282_U49 , P1_R1282_U50 , P1_R1282_U51 , P1_R1282_U52;
wire P1_R1282_U53 , P1_R1282_U54 , P1_R1282_U55 , P1_R1282_U56 , P1_R1282_U57 , P1_R1282_U58 , P1_R1282_U59 , P1_R1282_U60 , P1_R1282_U61 , P1_R1282_U62;
wire P1_R1282_U63 , P1_R1282_U64 , P1_R1282_U65 , P1_R1282_U66 , P1_R1282_U67 , P1_R1282_U68 , P1_R1282_U69 , P1_R1282_U70 , P1_R1282_U71 , P1_R1282_U72;
wire P1_R1282_U73 , P1_R1282_U74 , P1_R1282_U75 , P1_R1282_U76 , P1_R1282_U77 , P1_R1282_U78 , P1_R1282_U79 , P1_R1282_U80 , P1_R1282_U81 , P1_R1282_U82;
wire P1_R1282_U83 , P1_R1282_U84 , P1_R1282_U85 , P1_R1282_U86 , P1_R1282_U87 , P1_R1282_U88 , P1_R1282_U89 , P1_R1282_U90 , P1_R1282_U91 , P1_R1282_U92;
wire P1_R1282_U93 , P1_R1282_U94 , P1_R1282_U95 , P1_R1282_U96 , P1_R1282_U97 , P1_R1282_U98 , P1_R1282_U99 , P1_R1282_U100 , P1_R1282_U101 , P1_R1282_U102;
wire P1_R1282_U103 , P1_R1282_U104 , P1_R1282_U105 , P1_R1282_U106 , P1_R1282_U107 , P1_R1282_U108 , P1_R1282_U109 , P1_R1282_U110 , P1_R1282_U111 , P1_R1282_U112;
wire P1_R1282_U113 , P1_R1282_U114 , P1_R1282_U115 , P1_R1282_U116 , P1_R1282_U117 , P1_R1282_U118 , P1_R1282_U119 , P1_R1282_U120 , P1_R1282_U121 , P1_R1282_U122;
wire P1_R1282_U123 , P1_R1282_U124 , P1_R1282_U125 , P1_R1282_U126 , P1_R1282_U127 , P1_R1282_U128 , P1_R1282_U129 , P1_R1282_U130 , P1_R1282_U131 , P1_R1282_U132;
wire P1_R1282_U133 , P1_R1282_U134 , P1_R1282_U135 , P1_R1282_U136 , P1_R1282_U137 , P1_R1282_U138 , P1_R1282_U139 , P1_R1282_U140 , P1_R1282_U141 , P1_R1282_U142;
wire P1_R1282_U143 , P1_R1282_U144 , P1_R1282_U145 , P1_R1282_U146 , P1_R1282_U147 , P1_R1282_U148 , P1_R1282_U149 , P1_R1282_U150 , P1_R1282_U151 , P1_R1282_U152;
wire P1_R1282_U153 , P1_R1282_U154 , P1_R1282_U155 , P1_R1282_U156 , P1_R1282_U157 , P1_R1282_U158 , P1_R1282_U159 , P1_R1240_U4 , P1_R1240_U5 , P1_R1240_U6;
wire P1_R1240_U7 , P1_R1240_U8 , P1_R1240_U9 , P1_R1240_U10 , P1_R1240_U11 , P1_R1240_U12 , P1_R1240_U13 , P1_R1240_U14 , P1_R1240_U15 , P1_R1240_U16;
wire P1_R1240_U17 , P1_R1240_U18 , P1_R1240_U19 , P1_R1240_U20 , P1_R1240_U21 , P1_R1240_U22 , P1_R1240_U23 , P1_R1240_U24 , P1_R1240_U25 , P1_R1240_U26;
wire P1_R1240_U27 , P1_R1240_U28 , P1_R1240_U29 , P1_R1240_U30 , P1_R1240_U31 , P1_R1240_U32 , P1_R1240_U33 , P1_R1240_U34 , P1_R1240_U35 , P1_R1240_U36;
wire P1_R1240_U37 , P1_R1240_U38 , P1_R1240_U39 , P1_R1240_U40 , P1_R1240_U41 , P1_R1240_U42 , P1_R1240_U43 , P1_R1240_U44 , P1_R1240_U45 , P1_R1240_U46;
wire P1_R1240_U47 , P1_R1240_U48 , P1_R1240_U49 , P1_R1240_U50 , P1_R1240_U51 , P1_R1240_U52 , P1_R1240_U53 , P1_R1240_U54 , P1_R1240_U55 , P1_R1240_U56;
wire P1_R1240_U57 , P1_R1240_U58 , P1_R1240_U59 , P1_R1240_U60 , P1_R1240_U61 , P1_R1240_U62 , P1_R1240_U63 , P1_R1240_U64 , P1_R1240_U65 , P1_R1240_U66;
wire P1_R1240_U67 , P1_R1240_U68 , P1_R1240_U69 , P1_R1240_U70 , P1_R1240_U71 , P1_R1240_U72 , P1_R1240_U73 , P1_R1240_U74 , P1_R1240_U75 , P1_R1240_U76;
wire P1_R1240_U77 , P1_R1240_U78 , P1_R1240_U79 , P1_R1240_U80 , P1_R1240_U81 , P1_R1240_U82 , P1_R1240_U83 , P1_R1240_U84 , P1_R1240_U85 , P1_R1240_U86;
wire P1_R1240_U87 , P1_R1240_U88 , P1_R1240_U89 , P1_R1240_U90 , P1_R1240_U91 , P1_R1240_U92 , P1_R1240_U93 , P1_R1240_U94 , P1_R1240_U95 , P1_R1240_U96;
wire P1_R1240_U97 , P1_R1240_U98 , P1_R1240_U99 , P1_R1240_U100 , P1_R1240_U101 , P1_R1240_U102 , P1_R1240_U103 , P1_R1240_U104 , P1_R1240_U105 , P1_R1240_U106;
wire P1_R1240_U107 , P1_R1240_U108 , P1_R1240_U109 , P1_R1240_U110 , P1_R1240_U111 , P1_R1240_U112 , P1_R1240_U113 , P1_R1240_U114 , P1_R1240_U115 , P1_R1240_U116;
wire P1_R1240_U117 , P1_R1240_U118 , P1_R1240_U119 , P1_R1240_U120 , P1_R1240_U121 , P1_R1240_U122 , P1_R1240_U123 , P1_R1240_U124 , P1_R1240_U125 , P1_R1240_U126;
wire P1_R1240_U127 , P1_R1240_U128 , P1_R1240_U129 , P1_R1240_U130 , P1_R1240_U131 , P1_R1240_U132 , P1_R1240_U133 , P1_R1240_U134 , P1_R1240_U135 , P1_R1240_U136;
wire P1_R1240_U137 , P1_R1240_U138 , P1_R1240_U139 , P1_R1240_U140 , P1_R1240_U141 , P1_R1240_U142 , P1_R1240_U143 , P1_R1240_U144 , P1_R1240_U145 , P1_R1240_U146;
wire P1_R1240_U147 , P1_R1240_U148 , P1_R1240_U149 , P1_R1240_U150 , P1_R1240_U151 , P1_R1240_U152 , P1_R1240_U153 , P1_R1240_U154 , P1_R1240_U155 , P1_R1240_U156;
wire P1_R1240_U157 , P1_R1240_U158 , P1_R1240_U159 , P1_R1240_U160 , P1_R1240_U161 , P1_R1240_U162 , P1_R1240_U163 , P1_R1240_U164 , P1_R1240_U165 , P1_R1240_U166;
wire P1_R1240_U167 , P1_R1240_U168 , P1_R1240_U169 , P1_R1240_U170 , P1_R1240_U171 , P1_R1240_U172 , P1_R1240_U173 , P1_R1240_U174 , P1_R1240_U175 , P1_R1240_U176;
wire P1_R1240_U177 , P1_R1240_U178 , P1_R1240_U179 , P1_R1240_U180 , P1_R1240_U181 , P1_R1240_U182 , P1_R1240_U183 , P1_R1240_U184 , P1_R1240_U185 , P1_R1240_U186;
wire P1_R1240_U187 , P1_R1240_U188 , P1_R1240_U189 , P1_R1240_U190 , P1_R1240_U191 , P1_R1240_U192 , P1_R1240_U193 , P1_R1240_U194 , P1_R1240_U195 , P1_R1240_U196;
wire P1_R1240_U197 , P1_R1240_U198 , P1_R1240_U199 , P1_R1240_U200 , P1_R1240_U201 , P1_R1240_U202 , P1_R1240_U203 , P1_R1240_U204 , P1_R1240_U205 , P1_R1240_U206;
wire P1_R1240_U207 , P1_R1240_U208 , P1_R1240_U209 , P1_R1240_U210 , P1_R1240_U211 , P1_R1240_U212 , P1_R1240_U213 , P1_R1240_U214 , P1_R1240_U215 , P1_R1240_U216;
wire P1_R1240_U217 , P1_R1240_U218 , P1_R1240_U219 , P1_R1240_U220 , P1_R1240_U221 , P1_R1240_U222 , P1_R1240_U223 , P1_R1240_U224 , P1_R1240_U225 , P1_R1240_U226;
wire P1_R1240_U227 , P1_R1240_U228 , P1_R1240_U229 , P1_R1240_U230 , P1_R1240_U231 , P1_R1240_U232 , P1_R1240_U233 , P1_R1240_U234 , P1_R1240_U235 , P1_R1240_U236;
wire P1_R1240_U237 , P1_R1240_U238 , P1_R1240_U239 , P1_R1240_U240 , P1_R1240_U241 , P1_R1240_U242 , P1_R1240_U243 , P1_R1240_U244 , P1_R1240_U245 , P1_R1240_U246;
wire P1_R1240_U247 , P1_R1240_U248 , P1_R1240_U249 , P1_R1240_U250 , P1_R1240_U251 , P1_R1240_U252 , P1_R1240_U253 , P1_R1240_U254 , P1_R1240_U255 , P1_R1240_U256;
wire P1_R1240_U257 , P1_R1240_U258 , P1_R1240_U259 , P1_R1240_U260 , P1_R1240_U261 , P1_R1240_U262 , P1_R1240_U263 , P1_R1240_U264 , P1_R1240_U265 , P1_R1240_U266;
wire P1_R1240_U267 , P1_R1240_U268 , P1_R1240_U269 , P1_R1240_U270 , P1_R1240_U271 , P1_R1240_U272 , P1_R1240_U273 , P1_R1240_U274 , P1_R1240_U275 , P1_R1240_U276;
wire P1_R1240_U277 , P1_R1240_U278 , P1_R1240_U279 , P1_R1240_U280 , P1_R1240_U281 , P1_R1240_U282 , P1_R1240_U283 , P1_R1240_U284 , P1_R1240_U285 , P1_R1240_U286;
wire P1_R1240_U287 , P1_R1240_U288 , P1_R1240_U289 , P1_R1240_U290 , P1_R1240_U291 , P1_R1240_U292 , P1_R1240_U293 , P1_R1240_U294 , P1_R1240_U295 , P1_R1240_U296;
wire P1_R1240_U297 , P1_R1240_U298 , P1_R1240_U299 , P1_R1240_U300 , P1_R1240_U301 , P1_R1240_U302 , P1_R1240_U303 , P1_R1240_U304 , P1_R1240_U305 , P1_R1240_U306;
wire P1_R1240_U307 , P1_R1240_U308 , P1_R1240_U309 , P1_R1240_U310 , P1_R1240_U311 , P1_R1240_U312 , P1_R1240_U313 , P1_R1240_U314 , P1_R1240_U315 , P1_R1240_U316;
wire P1_R1240_U317 , P1_R1240_U318 , P1_R1240_U319 , P1_R1240_U320 , P1_R1240_U321 , P1_R1240_U322 , P1_R1240_U323 , P1_R1240_U324 , P1_R1240_U325 , P1_R1240_U326;
wire P1_R1240_U327 , P1_R1240_U328 , P1_R1240_U329 , P1_R1240_U330 , P1_R1240_U331 , P1_R1240_U332 , P1_R1240_U333 , P1_R1240_U334 , P1_R1240_U335 , P1_R1240_U336;
wire P1_R1240_U337 , P1_R1240_U338 , P1_R1240_U339 , P1_R1240_U340 , P1_R1240_U341 , P1_R1240_U342 , P1_R1240_U343 , P1_R1240_U344 , P1_R1240_U345 , P1_R1240_U346;
wire P1_R1240_U347 , P1_R1240_U348 , P1_R1240_U349 , P1_R1240_U350 , P1_R1240_U351 , P1_R1240_U352 , P1_R1240_U353 , P1_R1240_U354 , P1_R1240_U355 , P1_R1240_U356;
wire P1_R1240_U357 , P1_R1240_U358 , P1_R1240_U359 , P1_R1240_U360 , P1_R1240_U361 , P1_R1240_U362 , P1_R1240_U363 , P1_R1240_U364 , P1_R1240_U365 , P1_R1240_U366;
wire P1_R1240_U367 , P1_R1240_U368 , P1_R1240_U369 , P1_R1240_U370 , P1_R1240_U371 , P1_R1240_U372 , P1_R1240_U373 , P1_R1240_U374 , P1_R1240_U375 , P1_R1240_U376;
wire P1_R1240_U377 , P1_R1240_U378 , P1_R1240_U379 , P1_R1240_U380 , P1_R1240_U381 , P1_R1240_U382 , P1_R1240_U383 , P1_R1240_U384 , P1_R1240_U385 , P1_R1240_U386;
wire P1_R1240_U387 , P1_R1240_U388 , P1_R1240_U389 , P1_R1240_U390 , P1_R1240_U391 , P1_R1240_U392 , P1_R1240_U393 , P1_R1240_U394 , P1_R1240_U395 , P1_R1240_U396;
wire P1_R1240_U397 , P1_R1240_U398 , P1_R1240_U399 , P1_R1240_U400 , P1_R1240_U401 , P1_R1240_U402 , P1_R1240_U403 , P1_R1240_U404 , P1_R1240_U405 , P1_R1240_U406;
wire P1_R1240_U407 , P1_R1240_U408 , P1_R1240_U409 , P1_R1240_U410 , P1_R1240_U411 , P1_R1240_U412 , P1_R1240_U413 , P1_R1240_U414 , P1_R1240_U415 , P1_R1240_U416;
wire P1_R1240_U417 , P1_R1240_U418 , P1_R1240_U419 , P1_R1240_U420 , P1_R1240_U421 , P1_R1240_U422 , P1_R1240_U423 , P1_R1240_U424 , P1_R1240_U425 , P1_R1240_U426;
wire P1_R1240_U427 , P1_R1240_U428 , P1_R1240_U429 , P1_R1240_U430 , P1_R1240_U431 , P1_R1240_U432 , P1_R1240_U433 , P1_R1240_U434 , P1_R1240_U435 , P1_R1240_U436;
wire P1_R1240_U437 , P1_R1240_U438 , P1_R1240_U439 , P1_R1240_U440 , P1_R1240_U441 , P1_R1240_U442 , P1_R1240_U443 , P1_R1240_U444 , P1_R1240_U445 , P1_R1240_U446;
wire P1_R1240_U447 , P1_R1240_U448 , P1_R1240_U449 , P1_R1240_U450 , P1_R1240_U451 , P1_R1240_U452 , P1_R1240_U453 , P1_R1240_U454 , P1_R1240_U455 , P1_R1240_U456;
wire P1_R1240_U457 , P1_R1240_U458 , P1_R1240_U459 , P1_R1240_U460 , P1_R1240_U461 , P1_R1240_U462 , P1_R1240_U463 , P1_R1240_U464 , P1_R1240_U465 , P1_R1240_U466;
wire P1_R1240_U467 , P1_R1240_U468 , P1_R1240_U469 , P1_R1240_U470 , P1_R1240_U471 , P1_R1240_U472 , P1_R1240_U473 , P1_R1240_U474 , P1_R1240_U475 , P1_R1240_U476;
wire P1_R1240_U477 , P1_R1240_U478 , P1_R1240_U479 , P1_R1240_U480 , P1_R1240_U481 , P1_R1240_U482 , P1_R1240_U483 , P1_R1240_U484 , P1_R1240_U485 , P1_R1240_U486;
wire P1_R1240_U487 , P1_R1240_U488 , P1_R1240_U489 , P1_R1240_U490 , P1_R1240_U491 , P1_R1240_U492 , P1_R1240_U493 , P1_R1240_U494 , P1_R1240_U495 , P1_R1240_U496;
wire P1_R1240_U497 , P1_R1240_U498 , P1_R1240_U499 , P1_R1240_U500 , P1_R1240_U501 , P1_R1162_U4 , P1_R1162_U5 , P1_R1162_U6 , P1_R1162_U7 , P1_R1162_U8;
wire P1_R1162_U9 , P1_R1162_U10 , P1_R1162_U11 , P1_R1162_U12 , P1_R1162_U13 , P1_R1162_U14 , P1_R1162_U15 , P1_R1162_U16 , P1_R1162_U17 , P1_R1162_U18;
wire P1_R1162_U19 , P1_R1162_U20 , P1_R1162_U21 , P1_R1162_U22 , P1_R1162_U23 , P1_R1162_U24 , P1_R1162_U25 , P1_R1162_U26 , P1_R1162_U27 , P1_R1162_U28;
wire P1_R1162_U29 , P1_R1162_U30 , P1_R1162_U31 , P1_R1162_U32 , P1_R1162_U33 , P1_R1162_U34 , P1_R1162_U35 , P1_R1162_U36 , P1_R1162_U37 , P1_R1162_U38;
wire P1_R1162_U39 , P1_R1162_U40 , P1_R1162_U41 , P1_R1162_U42 , P1_R1162_U43 , P1_R1162_U44 , P1_R1162_U45 , P1_R1162_U46 , P1_R1162_U47 , P1_R1162_U48;
wire P1_R1162_U49 , P1_R1162_U50 , P1_R1162_U51 , P1_R1162_U52 , P1_R1162_U53 , P1_R1162_U54 , P1_R1162_U55 , P1_R1162_U56 , P1_R1162_U57 , P1_R1162_U58;
wire P1_R1162_U59 , P1_R1162_U60 , P1_R1162_U61 , P1_R1162_U62 , P1_R1162_U63 , P1_R1162_U64 , P1_R1162_U65 , P1_R1162_U66 , P1_R1162_U67 , P1_R1162_U68;
wire P1_R1162_U69 , P1_R1162_U70 , P1_R1162_U71 , P1_R1162_U72 , P1_R1162_U73 , P1_R1162_U74 , P1_R1162_U75 , P1_R1162_U76 , P1_R1162_U77 , P1_R1162_U78;
wire P1_R1162_U79 , P1_R1162_U80 , P1_R1162_U81 , P1_R1162_U82 , P1_R1162_U83 , P1_R1162_U84 , P1_R1162_U85 , P1_R1162_U86 , P1_R1162_U87 , P1_R1162_U88;
wire P1_R1162_U89 , P1_R1162_U90 , P1_R1162_U91 , P1_R1162_U92 , P1_R1162_U93 , P1_R1162_U94 , P1_R1162_U95 , P1_R1162_U96 , P1_R1162_U97 , P1_R1162_U98;
wire P1_R1162_U99 , P1_R1162_U100 , P1_R1162_U101 , P1_R1162_U102 , P1_R1162_U103 , P1_R1162_U104 , P1_R1162_U105 , P1_R1162_U106 , P1_R1162_U107 , P1_R1162_U108;
wire P1_R1162_U109 , P1_R1162_U110 , P1_R1162_U111 , P1_R1162_U112 , P1_R1162_U113 , P1_R1162_U114 , P1_R1162_U115 , P1_R1162_U116 , P1_R1162_U117 , P1_R1162_U118;
wire P1_R1162_U119 , P1_R1162_U120 , P1_R1162_U121 , P1_R1162_U122 , P1_R1162_U123 , P1_R1162_U124 , P1_R1162_U125 , P1_R1162_U126 , P1_R1162_U127 , P1_R1162_U128;
wire P1_R1162_U129 , P1_R1162_U130 , P1_R1162_U131 , P1_R1162_U132 , P1_R1162_U133 , P1_R1162_U134 , P1_R1162_U135 , P1_R1162_U136 , P1_R1162_U137 , P1_R1162_U138;
wire P1_R1162_U139 , P1_R1162_U140 , P1_R1162_U141 , P1_R1162_U142 , P1_R1162_U143 , P1_R1162_U144 , P1_R1162_U145 , P1_R1162_U146 , P1_R1162_U147 , P1_R1162_U148;
wire P1_R1162_U149 , P1_R1162_U150 , P1_R1162_U151 , P1_R1162_U152 , P1_R1162_U153 , P1_R1162_U154 , P1_R1162_U155 , P1_R1162_U156 , P1_R1162_U157 , P1_R1162_U158;
wire P1_R1162_U159 , P1_R1162_U160 , P1_R1162_U161 , P1_R1162_U162 , P1_R1162_U163 , P1_R1162_U164 , P1_R1162_U165 , P1_R1162_U166 , P1_R1162_U167 , P1_R1162_U168;
wire P1_R1162_U169 , P1_R1162_U170 , P1_R1162_U171 , P1_R1162_U172 , P1_R1162_U173 , P1_R1162_U174 , P1_R1162_U175 , P1_R1162_U176 , P1_R1162_U177 , P1_R1162_U178;
wire P1_R1162_U179 , P1_R1162_U180 , P1_R1162_U181 , P1_R1162_U182 , P1_R1162_U183 , P1_R1162_U184 , P1_R1162_U185 , P1_R1162_U186 , P1_R1162_U187 , P1_R1162_U188;
wire P1_R1162_U189 , P1_R1162_U190 , P1_R1162_U191 , P1_R1162_U192 , P1_R1162_U193 , P1_R1162_U194 , P1_R1162_U195 , P1_R1162_U196 , P1_R1162_U197 , P1_R1162_U198;
wire P1_R1162_U199 , P1_R1162_U200 , P1_R1162_U201 , P1_R1162_U202 , P1_R1162_U203 , P1_R1162_U204 , P1_R1162_U205 , P1_R1162_U206 , P1_R1162_U207 , P1_R1162_U208;
wire P1_R1162_U209 , P1_R1162_U210 , P1_R1162_U211 , P1_R1162_U212 , P1_R1162_U213 , P1_R1162_U214 , P1_R1162_U215 , P1_R1162_U216 , P1_R1162_U217 , P1_R1162_U218;
wire P1_R1162_U219 , P1_R1162_U220 , P1_R1162_U221 , P1_R1162_U222 , P1_R1162_U223 , P1_R1162_U224 , P1_R1162_U225 , P1_R1162_U226 , P1_R1162_U227 , P1_R1162_U228;
wire P1_R1162_U229 , P1_R1162_U230 , P1_R1162_U231 , P1_R1162_U232 , P1_R1162_U233 , P1_R1162_U234 , P1_R1162_U235 , P1_R1162_U236 , P1_R1162_U237 , P1_R1162_U238;
wire P1_R1162_U239 , P1_R1162_U240 , P1_R1162_U241 , P1_R1162_U242 , P1_R1162_U243 , P1_R1162_U244 , P1_R1162_U245 , P1_R1162_U246 , P1_R1162_U247 , P1_R1162_U248;
wire P1_R1162_U249 , P1_R1162_U250 , P1_R1162_U251 , P1_R1162_U252 , P1_R1162_U253 , P1_R1162_U254 , P1_R1162_U255 , P1_R1162_U256 , P1_R1162_U257 , P1_R1162_U258;
wire P1_R1162_U259 , P1_R1162_U260 , P1_R1162_U261 , P1_R1162_U262 , P1_R1162_U263 , P1_R1162_U264 , P1_R1162_U265 , P1_R1162_U266 , P1_R1162_U267 , P1_R1162_U268;
wire P1_R1162_U269 , P1_R1162_U270 , P1_R1162_U271 , P1_R1162_U272 , P1_R1162_U273 , P1_R1162_U274 , P1_R1162_U275 , P1_R1162_U276 , P1_R1162_U277 , P1_R1162_U278;
wire P1_R1162_U279 , P1_R1162_U280 , P1_R1162_U281 , P1_R1162_U282 , P1_R1162_U283 , P1_R1162_U284 , P1_R1162_U285 , P1_R1162_U286 , P1_R1162_U287 , P1_R1162_U288;
wire P1_R1162_U289 , P1_R1162_U290 , P1_R1162_U291 , P1_R1162_U292 , P1_R1162_U293 , P1_R1162_U294 , P1_R1162_U295 , P1_R1162_U296 , P1_R1162_U297 , P1_R1162_U298;
wire P1_R1162_U299 , P1_R1162_U300 , P1_R1162_U301 , P1_R1162_U302 , P1_R1162_U303 , P1_R1162_U304 , P1_R1162_U305 , P1_R1162_U306 , P1_R1162_U307 , P1_R1162_U308;
wire P1_R1117_U6 , P1_R1117_U7 , P1_R1117_U8 , P1_R1117_U9 , P1_R1117_U10 , P1_R1117_U11 , P1_R1117_U12 , P1_R1117_U13 , P1_R1117_U14 , P1_R1117_U15;
wire P1_R1117_U16 , P1_R1117_U17 , P1_R1117_U18 , P1_R1117_U19 , P1_R1117_U20 , P1_R1117_U21 , P1_R1117_U22 , P1_R1117_U23 , P1_R1117_U24 , P1_R1117_U25;
wire P1_R1117_U26 , P1_R1117_U27 , P1_R1117_U28 , P1_R1117_U29 , P1_R1117_U30 , P1_R1117_U31 , P1_R1117_U32 , P1_R1117_U33 , P1_R1117_U34 , P1_R1117_U35;
wire P1_R1117_U36 , P1_R1117_U37 , P1_R1117_U38 , P1_R1117_U39 , P1_R1117_U40 , P1_R1117_U41 , P1_R1117_U42 , P1_R1117_U43 , P1_R1117_U44 , P1_R1117_U45;
wire P1_R1117_U46 , P1_R1117_U47 , P1_R1117_U48 , P1_R1117_U49 , P1_R1117_U50 , P1_R1117_U51 , P1_R1117_U52 , P1_R1117_U53 , P1_R1117_U54 , P1_R1117_U55;
wire P1_R1117_U56 , P1_R1117_U57 , P1_R1117_U58 , P1_R1117_U59 , P1_R1117_U60 , P1_R1117_U61 , P1_R1117_U62 , P1_R1117_U63 , P1_R1117_U64 , P1_R1117_U65;
wire P1_R1117_U66 , P1_R1117_U67 , P1_R1117_U68 , P1_R1117_U69 , P1_R1117_U70 , P1_R1117_U71 , P1_R1117_U72 , P1_R1117_U73 , P1_R1117_U74 , P1_R1117_U75;
wire P1_R1117_U76 , P1_R1117_U77 , P1_R1117_U78 , P1_R1117_U79 , P1_R1117_U80 , P1_R1117_U81 , P1_R1117_U82 , P1_R1117_U83 , P1_R1117_U84 , P1_R1117_U85;
wire P1_R1117_U86 , P1_R1117_U87 , P1_R1117_U88 , P1_R1117_U89 , P1_R1117_U90 , P1_R1117_U91 , P1_R1117_U92 , P1_R1117_U93 , P1_R1117_U94 , P1_R1117_U95;
wire P1_R1117_U96 , P1_R1117_U97 , P1_R1117_U98 , P1_R1117_U99 , P1_R1117_U100 , P1_R1117_U101 , P1_R1117_U102 , P1_R1117_U103 , P1_R1117_U104 , P1_R1117_U105;
wire P1_R1117_U106 , P1_R1117_U107 , P1_R1117_U108 , P1_R1117_U109 , P1_R1117_U110 , P1_R1117_U111 , P1_R1117_U112 , P1_R1117_U113 , P1_R1117_U114 , P1_R1117_U115;
wire P1_R1117_U116 , P1_R1117_U117 , P1_R1117_U118 , P1_R1117_U119 , P1_R1117_U120 , P1_R1117_U121 , P1_R1117_U122 , P1_R1117_U123 , P1_R1117_U124 , P1_R1117_U125;
wire P1_R1117_U126 , P1_R1117_U127 , P1_R1117_U128 , P1_R1117_U129 , P1_R1117_U130 , P1_R1117_U131 , P1_R1117_U132 , P1_R1117_U133 , P1_R1117_U134 , P1_R1117_U135;
wire P1_R1117_U136 , P1_R1117_U137 , P1_R1117_U138 , P1_R1117_U139 , P1_R1117_U140 , P1_R1117_U141 , P1_R1117_U142 , P1_R1117_U143 , P1_R1117_U144 , P1_R1117_U145;
wire P1_R1117_U146 , P1_R1117_U147 , P1_R1117_U148 , P1_R1117_U149 , P1_R1117_U150 , P1_R1117_U151 , P1_R1117_U152 , P1_R1117_U153 , P1_R1117_U154 , P1_R1117_U155;
wire P1_R1117_U156 , P1_R1117_U157 , P1_R1117_U158 , P1_R1117_U159 , P1_R1117_U160 , P1_R1117_U161 , P1_R1117_U162 , P1_R1117_U163 , P1_R1117_U164 , P1_R1117_U165;
wire P1_R1117_U166 , P1_R1117_U167 , P1_R1117_U168 , P1_R1117_U169 , P1_R1117_U170 , P1_R1117_U171 , P1_R1117_U172 , P1_R1117_U173 , P1_R1117_U174 , P1_R1117_U175;
wire P1_R1117_U176 , P1_R1117_U177 , P1_R1117_U178 , P1_R1117_U179 , P1_R1117_U180 , P1_R1117_U181 , P1_R1117_U182 , P1_R1117_U183 , P1_R1117_U184 , P1_R1117_U185;
wire P1_R1117_U186 , P1_R1117_U187 , P1_R1117_U188 , P1_R1117_U189 , P1_R1117_U190 , P1_R1117_U191 , P1_R1117_U192 , P1_R1117_U193 , P1_R1117_U194 , P1_R1117_U195;
wire P1_R1117_U196 , P1_R1117_U197 , P1_R1117_U198 , P1_R1117_U199 , P1_R1117_U200 , P1_R1117_U201 , P1_R1117_U202 , P1_R1117_U203 , P1_R1117_U204 , P1_R1117_U205;
wire P1_R1117_U206 , P1_R1117_U207 , P1_R1117_U208 , P1_R1117_U209 , P1_R1117_U210 , P1_R1117_U211 , P1_R1117_U212 , P1_R1117_U213 , P1_R1117_U214 , P1_R1117_U215;
wire P1_R1117_U216 , P1_R1117_U217 , P1_R1117_U218 , P1_R1117_U219 , P1_R1117_U220 , P1_R1117_U221 , P1_R1117_U222 , P1_R1117_U223 , P1_R1117_U224 , P1_R1117_U225;
wire P1_R1117_U226 , P1_R1117_U227 , P1_R1117_U228 , P1_R1117_U229 , P1_R1117_U230 , P1_R1117_U231 , P1_R1117_U232 , P1_R1117_U233 , P1_R1117_U234 , P1_R1117_U235;
wire P1_R1117_U236 , P1_R1117_U237 , P1_R1117_U238 , P1_R1117_U239 , P1_R1117_U240 , P1_R1117_U241 , P1_R1117_U242 , P1_R1117_U243 , P1_R1117_U244 , P1_R1117_U245;
wire P1_R1117_U246 , P1_R1117_U247 , P1_R1117_U248 , P1_R1117_U249 , P1_R1117_U250 , P1_R1117_U251 , P1_R1117_U252 , P1_R1117_U253 , P1_R1117_U254 , P1_R1117_U255;
wire P1_R1117_U256 , P1_R1117_U257 , P1_R1117_U258 , P1_R1117_U259 , P1_R1117_U260 , P1_R1117_U261 , P1_R1117_U262 , P1_R1117_U263 , P1_R1117_U264 , P1_R1117_U265;
wire P1_R1117_U266 , P1_R1117_U267 , P1_R1117_U268 , P1_R1117_U269 , P1_R1117_U270 , P1_R1117_U271 , P1_R1117_U272 , P1_R1117_U273 , P1_R1117_U274 , P1_R1117_U275;
wire P1_R1117_U276 , P1_R1117_U277 , P1_R1117_U278 , P1_R1117_U279 , P1_R1117_U280 , P1_R1117_U281 , P1_R1117_U282 , P1_R1117_U283 , P1_R1117_U284 , P1_R1117_U285;
wire P1_R1117_U286 , P1_R1117_U287 , P1_R1117_U288 , P1_R1117_U289 , P1_R1117_U290 , P1_R1117_U291 , P1_R1117_U292 , P1_R1117_U293 , P1_R1117_U294 , P1_R1117_U295;
wire P1_R1117_U296 , P1_R1117_U297 , P1_R1117_U298 , P1_R1117_U299 , P1_R1117_U300 , P1_R1117_U301 , P1_R1117_U302 , P1_R1117_U303 , P1_R1117_U304 , P1_R1117_U305;
wire P1_R1117_U306 , P1_R1117_U307 , P1_R1117_U308 , P1_R1117_U309 , P1_R1117_U310 , P1_R1117_U311 , P1_R1117_U312 , P1_R1117_U313 , P1_R1117_U314 , P1_R1117_U315;
wire P1_R1117_U316 , P1_R1117_U317 , P1_R1117_U318 , P1_R1117_U319 , P1_R1117_U320 , P1_R1117_U321 , P1_R1117_U322 , P1_R1117_U323 , P1_R1117_U324 , P1_R1117_U325;
wire P1_R1117_U326 , P1_R1117_U327 , P1_R1117_U328 , P1_R1117_U329 , P1_R1117_U330 , P1_R1117_U331 , P1_R1117_U332 , P1_R1117_U333 , P1_R1117_U334 , P1_R1117_U335;
wire P1_R1117_U336 , P1_R1117_U337 , P1_R1117_U338 , P1_R1117_U339 , P1_R1117_U340 , P1_R1117_U341 , P1_R1117_U342 , P1_R1117_U343 , P1_R1117_U344 , P1_R1117_U345;
wire P1_R1117_U346 , P1_R1117_U347 , P1_R1117_U348 , P1_R1117_U349 , P1_R1117_U350 , P1_R1117_U351 , P1_R1117_U352 , P1_R1117_U353 , P1_R1117_U354 , P1_R1117_U355;
wire P1_R1117_U356 , P1_R1117_U357 , P1_R1117_U358 , P1_R1117_U359 , P1_R1117_U360 , P1_R1117_U361 , P1_R1117_U362 , P1_R1117_U363 , P1_R1117_U364 , P1_R1117_U365;
wire P1_R1117_U366 , P1_R1117_U367 , P1_R1117_U368 , P1_R1117_U369 , P1_R1117_U370 , P1_R1117_U371 , P1_R1117_U372 , P1_R1117_U373 , P1_R1117_U374 , P1_R1117_U375;
wire P1_R1117_U376 , P1_R1117_U377 , P1_R1117_U378 , P1_R1117_U379 , P1_R1117_U380 , P1_R1117_U381 , P1_R1117_U382 , P1_R1117_U383 , P1_R1117_U384 , P1_R1117_U385;
wire P1_R1117_U386 , P1_R1117_U387 , P1_R1117_U388 , P1_R1117_U389 , P1_R1117_U390 , P1_R1117_U391 , P1_R1117_U392 , P1_R1117_U393 , P1_R1117_U394 , P1_R1117_U395;
wire P1_R1117_U396 , P1_R1117_U397 , P1_R1117_U398 , P1_R1117_U399 , P1_R1117_U400 , P1_R1117_U401 , P1_R1117_U402 , P1_R1117_U403 , P1_R1117_U404 , P1_R1117_U405;
wire P1_R1117_U406 , P1_R1117_U407 , P1_R1117_U408 , P1_R1117_U409 , P1_R1117_U410 , P1_R1117_U411 , P1_R1117_U412 , P1_R1117_U413 , P1_R1117_U414 , P1_R1117_U415;
wire P1_R1117_U416 , P1_R1117_U417 , P1_R1117_U418 , P1_R1117_U419 , P1_R1117_U420 , P1_R1117_U421 , P1_R1117_U422 , P1_R1117_U423 , P1_R1117_U424 , P1_R1117_U425;
wire P1_R1117_U426 , P1_R1117_U427 , P1_R1117_U428 , P1_R1117_U429 , P1_R1117_U430 , P1_R1117_U431 , P1_R1117_U432 , P1_R1117_U433 , P1_R1117_U434 , P1_R1117_U435;
wire P1_R1117_U436 , P1_R1117_U437 , P1_R1117_U438 , P1_R1117_U439 , P1_R1117_U440 , P1_R1117_U441 , P1_R1117_U442 , P1_R1117_U443 , P1_R1117_U444 , P1_R1117_U445;
wire P1_R1117_U446 , P1_R1117_U447 , P1_R1117_U448 , P1_R1117_U449 , P1_R1117_U450 , P1_R1117_U451 , P1_R1117_U452 , P1_R1117_U453 , P1_R1117_U454 , P1_R1117_U455;
wire P1_R1117_U456 , P1_R1117_U457 , P1_R1117_U458 , P1_R1117_U459 , P1_R1117_U460 , P1_R1117_U461 , P1_R1117_U462 , P1_R1117_U463 , P1_R1117_U464 , P1_R1117_U465;
wire P1_R1117_U466 , P1_R1117_U467 , P1_R1117_U468 , P1_R1117_U469 , P1_R1117_U470 , P1_R1117_U471 , P1_R1117_U472 , P1_R1117_U473 , P1_R1117_U474 , P1_R1117_U475;
wire P1_R1117_U476 , P1_R1375_U6 , P1_R1375_U7 , P1_R1375_U8 , P1_R1375_U9 , P1_R1375_U10 , P1_R1375_U11 , P1_R1375_U12 , P1_R1375_U13 , P1_R1375_U14;
wire P1_R1375_U15 , P1_R1375_U16 , P1_R1375_U17 , P1_R1375_U18 , P1_R1375_U19 , P1_R1375_U20 , P1_R1375_U21 , P1_R1375_U22 , P1_R1375_U23 , P1_R1375_U24;
wire P1_R1375_U25 , P1_R1375_U26 , P1_R1375_U27 , P1_R1375_U28 , P1_R1375_U29 , P1_R1375_U30 , P1_R1375_U31 , P1_R1375_U32 , P1_R1375_U33 , P1_R1375_U34;
wire P1_R1375_U35 , P1_R1375_U36 , P1_R1375_U37 , P1_R1375_U38 , P1_R1375_U39 , P1_R1375_U40 , P1_R1375_U41 , P1_R1375_U42 , P1_R1375_U43 , P1_R1375_U44;
wire P1_R1375_U45 , P1_R1375_U46 , P1_R1375_U47 , P1_R1375_U48 , P1_R1375_U49 , P1_R1375_U50 , P1_R1375_U51 , P1_R1375_U52 , P1_R1375_U53 , P1_R1375_U54;
wire P1_R1375_U55 , P1_R1375_U56 , P1_R1375_U57 , P1_R1375_U58 , P1_R1375_U59 , P1_R1375_U60 , P1_R1375_U61 , P1_R1375_U62 , P1_R1375_U63 , P1_R1375_U64;
wire P1_R1375_U65 , P1_R1375_U66 , P1_R1375_U67 , P1_R1375_U68 , P1_R1375_U69 , P1_R1375_U70 , P1_R1375_U71 , P1_R1375_U72 , P1_R1375_U73 , P1_R1375_U74;
wire P1_R1375_U75 , P1_R1375_U76 , P1_R1375_U77 , P1_R1375_U78 , P1_R1375_U79 , P1_R1375_U80 , P1_R1375_U81 , P1_R1375_U82 , P1_R1375_U83 , P1_R1375_U84;
wire P1_R1375_U85 , P1_R1375_U86 , P1_R1375_U87 , P1_R1375_U88 , P1_R1375_U89 , P1_R1375_U90 , P1_R1375_U91 , P1_R1375_U92 , P1_R1375_U93 , P1_R1375_U94;
wire P1_R1375_U95 , P1_R1375_U96 , P1_R1375_U97 , P1_R1375_U98 , P1_R1375_U99 , P1_R1375_U100 , P1_R1375_U101 , P1_R1375_U102 , P1_R1375_U103 , P1_R1375_U104;
wire P1_R1375_U105 , P1_R1375_U106 , P1_R1375_U107 , P1_R1375_U108 , P1_R1375_U109 , P1_R1375_U110 , P1_R1375_U111 , P1_R1375_U112 , P1_R1375_U113 , P1_R1375_U114;
wire P1_R1375_U115 , P1_R1375_U116 , P1_R1375_U117 , P1_R1375_U118 , P1_R1375_U119 , P1_R1375_U120 , P1_R1375_U121 , P1_R1375_U122 , P1_R1375_U123 , P1_R1375_U124;
wire P1_R1375_U125 , P1_R1375_U126 , P1_R1375_U127 , P1_R1375_U128 , P1_R1375_U129 , P1_R1375_U130 , P1_R1375_U131 , P1_R1375_U132 , P1_R1375_U133 , P1_R1375_U134;
wire P1_R1375_U135 , P1_R1375_U136 , P1_R1375_U137 , P1_R1375_U138 , P1_R1375_U139 , P1_R1375_U140 , P1_R1375_U141 , P1_R1375_U142 , P1_R1375_U143 , P1_R1375_U144;
wire P1_R1375_U145 , P1_R1375_U146 , P1_R1375_U147 , P1_R1375_U148 , P1_R1375_U149 , P1_R1375_U150 , P1_R1375_U151 , P1_R1375_U152 , P1_R1375_U153 , P1_R1375_U154;
wire P1_R1375_U155 , P1_R1375_U156 , P1_R1375_U157 , P1_R1375_U158 , P1_R1375_U159 , P1_R1375_U160 , P1_R1375_U161 , P1_R1375_U162 , P1_R1375_U163 , P1_R1375_U164;
wire P1_R1375_U165 , P1_R1375_U166 , P1_R1375_U167 , P1_R1375_U168 , P1_R1375_U169 , P1_R1375_U170 , P1_R1375_U171 , P1_R1375_U172 , P1_R1375_U173 , P1_R1375_U174;
wire P1_R1375_U175 , P1_R1375_U176 , P1_R1375_U177 , P1_R1375_U178 , P1_R1375_U179 , P1_R1375_U180 , P1_R1375_U181 , P1_R1375_U182 , P1_R1375_U183 , P1_R1375_U184;
wire P1_R1375_U185 , P1_R1375_U186 , P1_R1375_U187 , P1_R1375_U188 , P1_R1375_U189 , P1_R1375_U190 , P1_R1375_U191 , P1_R1375_U192 , P1_R1375_U193 , P1_R1375_U194;
wire P1_R1375_U195 , P1_R1375_U196 , P1_R1375_U197 , P1_R1375_U198 , P1_R1375_U199 , P1_R1375_U200 , P1_R1375_U201 , P1_R1375_U202 , P1_R1375_U203 , P1_R1375_U204;
wire P1_R1375_U205 , P1_R1375_U206 , P1_R1375_U207 , P1_R1352_U6 , P1_R1352_U7 , P1_R1207_U6 , P1_R1207_U7 , P1_R1207_U8 , P1_R1207_U9 , P1_R1207_U10;
wire P1_R1207_U11 , P1_R1207_U12 , P1_R1207_U13 , P1_R1207_U14 , P1_R1207_U15 , P1_R1207_U16 , P1_R1207_U17 , P1_R1207_U18 , P1_R1207_U19 , P1_R1207_U20;
wire P1_R1207_U21 , P1_R1207_U22 , P1_R1207_U23 , P1_R1207_U24 , P1_R1207_U25 , P1_R1207_U26 , P1_R1207_U27 , P1_R1207_U28 , P1_R1207_U29 , P1_R1207_U30;
wire P1_R1207_U31 , P1_R1207_U32 , P1_R1207_U33 , P1_R1207_U34 , P1_R1207_U35 , P1_R1207_U36 , P1_R1207_U37 , P1_R1207_U38 , P1_R1207_U39 , P1_R1207_U40;
wire P1_R1207_U41 , P1_R1207_U42 , P1_R1207_U43 , P1_R1207_U44 , P1_R1207_U45 , P1_R1207_U46 , P1_R1207_U47 , P1_R1207_U48 , P1_R1207_U49 , P1_R1207_U50;
wire P1_R1207_U51 , P1_R1207_U52 , P1_R1207_U53 , P1_R1207_U54 , P1_R1207_U55 , P1_R1207_U56 , P1_R1207_U57 , P1_R1207_U58 , P1_R1207_U59 , P1_R1207_U60;
wire P1_R1207_U61 , P1_R1207_U62 , P1_R1207_U63 , P1_R1207_U64 , P1_R1207_U65 , P1_R1207_U66 , P1_R1207_U67 , P1_R1207_U68 , P1_R1207_U69 , P1_R1207_U70;
wire P1_R1207_U71 , P1_R1207_U72 , P1_R1207_U73 , P1_R1207_U74 , P1_R1207_U75 , P1_R1207_U76 , P1_R1207_U77 , P1_R1207_U78 , P1_R1207_U79 , P1_R1207_U80;
wire P1_R1207_U81 , P1_R1207_U82 , P1_R1207_U83 , P1_R1207_U84 , P1_R1207_U85 , P1_R1207_U86 , P1_R1207_U87 , P1_R1207_U88 , P1_R1207_U89 , P1_R1207_U90;
wire P1_R1207_U91 , P1_R1207_U92 , P1_R1207_U93 , P1_R1207_U94 , P1_R1207_U95 , P1_R1207_U96 , P1_R1207_U97 , P1_R1207_U98 , P1_R1207_U99 , P1_R1207_U100;
wire P1_R1207_U101 , P1_R1207_U102 , P1_R1207_U103 , P1_R1207_U104 , P1_R1207_U105 , P1_R1207_U106 , P1_R1207_U107 , P1_R1207_U108 , P1_R1207_U109 , P1_R1207_U110;
wire P1_R1207_U111 , P1_R1207_U112 , P1_R1207_U113 , P1_R1207_U114 , P1_R1207_U115 , P1_R1207_U116 , P1_R1207_U117 , P1_R1207_U118 , P1_R1207_U119 , P1_R1207_U120;
wire P1_R1207_U121 , P1_R1207_U122 , P1_R1207_U123 , P1_R1207_U124 , P1_R1207_U125 , P1_R1207_U126 , P1_R1207_U127 , P1_R1207_U128 , P1_R1207_U129 , P1_R1207_U130;
wire P1_R1207_U131 , P1_R1207_U132 , P1_R1207_U133 , P1_R1207_U134 , P1_R1207_U135 , P1_R1207_U136 , P1_R1207_U137 , P1_R1207_U138 , P1_R1207_U139 , P1_R1207_U140;
wire P1_R1207_U141 , P1_R1207_U142 , P1_R1207_U143 , P1_R1207_U144 , P1_R1207_U145 , P1_R1207_U146 , P1_R1207_U147 , P1_R1207_U148 , P1_R1207_U149 , P1_R1207_U150;
wire P1_R1207_U151 , P1_R1207_U152 , P1_R1207_U153 , P1_R1207_U154 , P1_R1207_U155 , P1_R1207_U156 , P1_R1207_U157 , P1_R1207_U158 , P1_R1207_U159 , P1_R1207_U160;
wire P1_R1207_U161 , P1_R1207_U162 , P1_R1207_U163 , P1_R1207_U164 , P1_R1207_U165 , P1_R1207_U166 , P1_R1207_U167 , P1_R1207_U168 , P1_R1207_U169 , P1_R1207_U170;
wire P1_R1207_U171 , P1_R1207_U172 , P1_R1207_U173 , P1_R1207_U174 , P1_R1207_U175 , P1_R1207_U176 , P1_R1207_U177 , P1_R1207_U178 , P1_R1207_U179 , P1_R1207_U180;
wire P1_R1207_U181 , P1_R1207_U182 , P1_R1207_U183 , P1_R1207_U184 , P1_R1207_U185 , P1_R1207_U186 , P1_R1207_U187 , P1_R1207_U188 , P1_R1207_U189 , P1_R1207_U190;
wire P1_R1207_U191 , P1_R1207_U192 , P1_R1207_U193 , P1_R1207_U194 , P1_R1207_U195 , P1_R1207_U196 , P1_R1207_U197 , P1_R1207_U198 , P1_R1207_U199 , P1_R1207_U200;
wire P1_R1207_U201 , P1_R1207_U202 , P1_R1207_U203 , P1_R1207_U204 , P1_R1207_U205 , P1_R1207_U206 , P1_R1207_U207 , P1_R1207_U208 , P1_R1207_U209 , P1_R1207_U210;
wire P1_R1207_U211 , P1_R1207_U212 , P1_R1207_U213 , P1_R1207_U214 , P1_R1207_U215 , P1_R1207_U216 , P1_R1207_U217 , P1_R1207_U218 , P1_R1207_U219 , P1_R1207_U220;
wire P1_R1207_U221 , P1_R1207_U222 , P1_R1207_U223 , P1_R1207_U224 , P1_R1207_U225 , P1_R1207_U226 , P1_R1207_U227 , P1_R1207_U228 , P1_R1207_U229 , P1_R1207_U230;
wire P1_R1207_U231 , P1_R1207_U232 , P1_R1207_U233 , P1_R1207_U234 , P1_R1207_U235 , P1_R1207_U236 , P1_R1207_U237 , P1_R1207_U238 , P1_R1207_U239 , P1_R1207_U240;
wire P1_R1207_U241 , P1_R1207_U242 , P1_R1207_U243 , P1_R1207_U244 , P1_R1207_U245 , P1_R1207_U246 , P1_R1207_U247 , P1_R1207_U248 , P1_R1207_U249 , P1_R1207_U250;
wire P1_R1207_U251 , P1_R1207_U252 , P1_R1207_U253 , P1_R1207_U254 , P1_R1207_U255 , P1_R1207_U256 , P1_R1207_U257 , P1_R1207_U258 , P1_R1207_U259 , P1_R1207_U260;
wire P1_R1207_U261 , P1_R1207_U262 , P1_R1207_U263 , P1_R1207_U264 , P1_R1207_U265 , P1_R1207_U266 , P1_R1207_U267 , P1_R1207_U268 , P1_R1207_U269 , P1_R1207_U270;
wire P1_R1207_U271 , P1_R1207_U272 , P1_R1207_U273 , P1_R1207_U274 , P1_R1207_U275 , P1_R1207_U276 , P1_R1207_U277 , P1_R1207_U278 , P1_R1207_U279 , P1_R1207_U280;
wire P1_R1207_U281 , P1_R1207_U282 , P1_R1207_U283 , P1_R1207_U284 , P1_R1207_U285 , P1_R1207_U286 , P1_R1207_U287 , P1_R1207_U288 , P1_R1207_U289 , P1_R1207_U290;
wire P1_R1207_U291 , P1_R1207_U292 , P1_R1207_U293 , P1_R1207_U294 , P1_R1207_U295 , P1_R1207_U296 , P1_R1207_U297 , P1_R1207_U298 , P1_R1207_U299 , P1_R1207_U300;
wire P1_R1207_U301 , P1_R1207_U302 , P1_R1207_U303 , P1_R1207_U304 , P1_R1207_U305 , P1_R1207_U306 , P1_R1207_U307 , P1_R1207_U308 , P1_R1207_U309 , P1_R1207_U310;
wire P1_R1207_U311 , P1_R1207_U312 , P1_R1207_U313 , P1_R1207_U314 , P1_R1207_U315 , P1_R1207_U316 , P1_R1207_U317 , P1_R1207_U318 , P1_R1207_U319 , P1_R1207_U320;
wire P1_R1207_U321 , P1_R1207_U322 , P1_R1207_U323 , P1_R1207_U324 , P1_R1207_U325 , P1_R1207_U326 , P1_R1207_U327 , P1_R1207_U328 , P1_R1207_U329 , P1_R1207_U330;
wire P1_R1207_U331 , P1_R1207_U332 , P1_R1207_U333 , P1_R1207_U334 , P1_R1207_U335 , P1_R1207_U336 , P1_R1207_U337 , P1_R1207_U338 , P1_R1207_U339 , P1_R1207_U340;
wire P1_R1207_U341 , P1_R1207_U342 , P1_R1207_U343 , P1_R1207_U344 , P1_R1207_U345 , P1_R1207_U346 , P1_R1207_U347 , P1_R1207_U348 , P1_R1207_U349 , P1_R1207_U350;
wire P1_R1207_U351 , P1_R1207_U352 , P1_R1207_U353 , P1_R1207_U354 , P1_R1207_U355 , P1_R1207_U356 , P1_R1207_U357 , P1_R1207_U358 , P1_R1207_U359 , P1_R1207_U360;
wire P1_R1207_U361 , P1_R1207_U362 , P1_R1207_U363 , P1_R1207_U364 , P1_R1207_U365 , P1_R1207_U366 , P1_R1207_U367 , P1_R1207_U368 , P1_R1207_U369 , P1_R1207_U370;
wire P1_R1207_U371 , P1_R1207_U372 , P1_R1207_U373 , P1_R1207_U374 , P1_R1207_U375 , P1_R1207_U376 , P1_R1207_U377 , P1_R1207_U378 , P1_R1207_U379 , P1_R1207_U380;
wire P1_R1207_U381 , P1_R1207_U382 , P1_R1207_U383 , P1_R1207_U384 , P1_R1207_U385 , P1_R1207_U386 , P1_R1207_U387 , P1_R1207_U388 , P1_R1207_U389 , P1_R1207_U390;
wire P1_R1207_U391 , P1_R1207_U392 , P1_R1207_U393 , P1_R1207_U394 , P1_R1207_U395 , P1_R1207_U396 , P1_R1207_U397 , P1_R1207_U398 , P1_R1207_U399 , P1_R1207_U400;
wire P1_R1207_U401 , P1_R1207_U402 , P1_R1207_U403 , P1_R1207_U404 , P1_R1207_U405 , P1_R1207_U406 , P1_R1207_U407 , P1_R1207_U408 , P1_R1207_U409 , P1_R1207_U410;
wire P1_R1207_U411 , P1_R1207_U412 , P1_R1207_U413 , P1_R1207_U414 , P1_R1207_U415 , P1_R1207_U416 , P1_R1207_U417 , P1_R1207_U418 , P1_R1207_U419 , P1_R1207_U420;
wire P1_R1207_U421 , P1_R1207_U422 , P1_R1207_U423 , P1_R1207_U424 , P1_R1207_U425 , P1_R1207_U426 , P1_R1207_U427 , P1_R1207_U428 , P1_R1207_U429 , P1_R1207_U430;
wire P1_R1207_U431 , P1_R1207_U432 , P1_R1207_U433 , P1_R1207_U434 , P1_R1207_U435 , P1_R1207_U436 , P1_R1207_U437 , P1_R1207_U438 , P1_R1207_U439 , P1_R1207_U440;
wire P1_R1207_U441 , P1_R1207_U442 , P1_R1207_U443 , P1_R1207_U444 , P1_R1207_U445 , P1_R1207_U446 , P1_R1207_U447 , P1_R1207_U448 , P1_R1207_U449 , P1_R1207_U450;
wire P1_R1207_U451 , P1_R1207_U452 , P1_R1207_U453 , P1_R1207_U454 , P1_R1207_U455 , P1_R1207_U456 , P1_R1207_U457 , P1_R1207_U458 , P1_R1207_U459 , P1_R1207_U460;
wire P1_R1207_U461 , P1_R1207_U462 , P1_R1207_U463 , P1_R1207_U464 , P1_R1207_U465 , P1_R1207_U466 , P1_R1207_U467 , P1_R1207_U468 , P1_R1207_U469 , P1_R1207_U470;
wire P1_R1207_U471 , P1_R1207_U472 , P1_R1207_U473 , P1_R1207_U474 , P1_R1207_U475 , P1_R1207_U476 , P1_R1165_U4 , P1_R1165_U5 , P1_R1165_U6 , P1_R1165_U7;
wire P1_R1165_U8 , P1_R1165_U9 , P1_R1165_U10 , P1_R1165_U11 , P1_R1165_U12 , P1_R1165_U13 , P1_R1165_U14 , P1_R1165_U15 , P1_R1165_U16 , P1_R1165_U17;
wire P1_R1165_U18 , P1_R1165_U19 , P1_R1165_U20 , P1_R1165_U21 , P1_R1165_U22 , P1_R1165_U23 , P1_R1165_U24 , P1_R1165_U25 , P1_R1165_U26 , P1_R1165_U27;
wire P1_R1165_U28 , P1_R1165_U29 , P1_R1165_U30 , P1_R1165_U31 , P1_R1165_U32 , P1_R1165_U33 , P1_R1165_U34 , P1_R1165_U35 , P1_R1165_U36 , P1_R1165_U37;
wire P1_R1165_U38 , P1_R1165_U39 , P1_R1165_U40 , P1_R1165_U41 , P1_R1165_U42 , P1_R1165_U43 , P1_R1165_U44 , P1_R1165_U45 , P1_R1165_U46 , P1_R1165_U47;
wire P1_R1165_U48 , P1_R1165_U49 , P1_R1165_U50 , P1_R1165_U51 , P1_R1165_U52 , P1_R1165_U53 , P1_R1165_U54 , P1_R1165_U55 , P1_R1165_U56 , P1_R1165_U57;
wire P1_R1165_U58 , P1_R1165_U59 , P1_R1165_U60 , P1_R1165_U61 , P1_R1165_U62 , P1_R1165_U63 , P1_R1165_U64 , P1_R1165_U65 , P1_R1165_U66 , P1_R1165_U67;
wire P1_R1165_U68 , P1_R1165_U69 , P1_R1165_U70 , P1_R1165_U71 , P1_R1165_U72 , P1_R1165_U73 , P1_R1165_U74 , P1_R1165_U75 , P1_R1165_U76 , P1_R1165_U77;
wire P1_R1165_U78 , P1_R1165_U79 , P1_R1165_U80 , P1_R1165_U81 , P1_R1165_U82 , P1_R1165_U83 , P1_R1165_U84 , P1_R1165_U85 , P1_R1165_U86 , P1_R1165_U87;
wire P1_R1165_U88 , P1_R1165_U89 , P1_R1165_U90 , P1_R1165_U91 , P1_R1165_U92 , P1_R1165_U93 , P1_R1165_U94 , P1_R1165_U95 , P1_R1165_U96 , P1_R1165_U97;
wire P1_R1165_U98 , P1_R1165_U99 , P1_R1165_U100 , P1_R1165_U101 , P1_R1165_U102 , P1_R1165_U103 , P1_R1165_U104 , P1_R1165_U105 , P1_R1165_U106 , P1_R1165_U107;
wire P1_R1165_U108 , P1_R1165_U109 , P1_R1165_U110 , P1_R1165_U111 , P1_R1165_U112 , P1_R1165_U113 , P1_R1165_U114 , P1_R1165_U115 , P1_R1165_U116 , P1_R1165_U117;
wire P1_R1165_U118 , P1_R1165_U119 , P1_R1165_U120 , P1_R1165_U121 , P1_R1165_U122 , P1_R1165_U123 , P1_R1165_U124 , P1_R1165_U125 , P1_R1165_U126 , P1_R1165_U127;
wire P1_R1165_U128 , P1_R1165_U129 , P1_R1165_U130 , P1_R1165_U131 , P1_R1165_U132 , P1_R1165_U133 , P1_R1165_U134 , P1_R1165_U135 , P1_R1165_U136 , P1_R1165_U137;
wire P1_R1165_U138 , P1_R1165_U139 , P1_R1165_U140 , P1_R1165_U141 , P1_R1165_U142 , P1_R1165_U143 , P1_R1165_U144 , P1_R1165_U145 , P1_R1165_U146 , P1_R1165_U147;
wire P1_R1165_U148 , P1_R1165_U149 , P1_R1165_U150 , P1_R1165_U151 , P1_R1165_U152 , P1_R1165_U153 , P1_R1165_U154 , P1_R1165_U155 , P1_R1165_U156 , P1_R1165_U157;
wire P1_R1165_U158 , P1_R1165_U159 , P1_R1165_U160 , P1_R1165_U161 , P1_R1165_U162 , P1_R1165_U163 , P1_R1165_U164 , P1_R1165_U165 , P1_R1165_U166 , P1_R1165_U167;
wire P1_R1165_U168 , P1_R1165_U169 , P1_R1165_U170 , P1_R1165_U171 , P1_R1165_U172 , P1_R1165_U173 , P1_R1165_U174 , P1_R1165_U175 , P1_R1165_U176 , P1_R1165_U177;
wire P1_R1165_U178 , P1_R1165_U179 , P1_R1165_U180 , P1_R1165_U181 , P1_R1165_U182 , P1_R1165_U183 , P1_R1165_U184 , P1_R1165_U185 , P1_R1165_U186 , P1_R1165_U187;
wire P1_R1165_U188 , P1_R1165_U189 , P1_R1165_U190 , P1_R1165_U191 , P1_R1165_U192 , P1_R1165_U193 , P1_R1165_U194 , P1_R1165_U195 , P1_R1165_U196 , P1_R1165_U197;
wire P1_R1165_U198 , P1_R1165_U199 , P1_R1165_U200 , P1_R1165_U201 , P1_R1165_U202 , P1_R1165_U203 , P1_R1165_U204 , P1_R1165_U205 , P1_R1165_U206 , P1_R1165_U207;
wire P1_R1165_U208 , P1_R1165_U209 , P1_R1165_U210 , P1_R1165_U211 , P1_R1165_U212 , P1_R1165_U213 , P1_R1165_U214 , P1_R1165_U215 , P1_R1165_U216 , P1_R1165_U217;
wire P1_R1165_U218 , P1_R1165_U219 , P1_R1165_U220 , P1_R1165_U221 , P1_R1165_U222 , P1_R1165_U223 , P1_R1165_U224 , P1_R1165_U225 , P1_R1165_U226 , P1_R1165_U227;
wire P1_R1165_U228 , P1_R1165_U229 , P1_R1165_U230 , P1_R1165_U231 , P1_R1165_U232 , P1_R1165_U233 , P1_R1165_U234 , P1_R1165_U235 , P1_R1165_U236 , P1_R1165_U237;
wire P1_R1165_U238 , P1_R1165_U239 , P1_R1165_U240 , P1_R1165_U241 , P1_R1165_U242 , P1_R1165_U243 , P1_R1165_U244 , P1_R1165_U245 , P1_R1165_U246 , P1_R1165_U247;
wire P1_R1165_U248 , P1_R1165_U249 , P1_R1165_U250 , P1_R1165_U251 , P1_R1165_U252 , P1_R1165_U253 , P1_R1165_U254 , P1_R1165_U255 , P1_R1165_U256 , P1_R1165_U257;
wire P1_R1165_U258 , P1_R1165_U259 , P1_R1165_U260 , P1_R1165_U261 , P1_R1165_U262 , P1_R1165_U263 , P1_R1165_U264 , P1_R1165_U265 , P1_R1165_U266 , P1_R1165_U267;
wire P1_R1165_U268 , P1_R1165_U269 , P1_R1165_U270 , P1_R1165_U271 , P1_R1165_U272 , P1_R1165_U273 , P1_R1165_U274 , P1_R1165_U275 , P1_R1165_U276 , P1_R1165_U277;
wire P1_R1165_U278 , P1_R1165_U279 , P1_R1165_U280 , P1_R1165_U281 , P1_R1165_U282 , P1_R1165_U283 , P1_R1165_U284 , P1_R1165_U285 , P1_R1165_U286 , P1_R1165_U287;
wire P1_R1165_U288 , P1_R1165_U289 , P1_R1165_U290 , P1_R1165_U291 , P1_R1165_U292 , P1_R1165_U293 , P1_R1165_U294 , P1_R1165_U295 , P1_R1165_U296 , P1_R1165_U297;
wire P1_R1165_U298 , P1_R1165_U299 , P1_R1165_U300 , P1_R1165_U301 , P1_R1165_U302 , P1_R1165_U303 , P1_R1165_U304 , P1_R1165_U305 , P1_R1165_U306 , P1_R1165_U307;
wire P1_R1165_U308 , P1_R1165_U309 , P1_R1165_U310 , P1_R1165_U311 , P1_R1165_U312 , P1_R1165_U313 , P1_R1165_U314 , P1_R1165_U315 , P1_R1165_U316 , P1_R1165_U317;
wire P1_R1165_U318 , P1_R1165_U319 , P1_R1165_U320 , P1_R1165_U321 , P1_R1165_U322 , P1_R1165_U323 , P1_R1165_U324 , P1_R1165_U325 , P1_R1165_U326 , P1_R1165_U327;
wire P1_R1165_U328 , P1_R1165_U329 , P1_R1165_U330 , P1_R1165_U331 , P1_R1165_U332 , P1_R1165_U333 , P1_R1165_U334 , P1_R1165_U335 , P1_R1165_U336 , P1_R1165_U337;
wire P1_R1165_U338 , P1_R1165_U339 , P1_R1165_U340 , P1_R1165_U341 , P1_R1165_U342 , P1_R1165_U343 , P1_R1165_U344 , P1_R1165_U345 , P1_R1165_U346 , P1_R1165_U347;
wire P1_R1165_U348 , P1_R1165_U349 , P1_R1165_U350 , P1_R1165_U351 , P1_R1165_U352 , P1_R1165_U353 , P1_R1165_U354 , P1_R1165_U355 , P1_R1165_U356 , P1_R1165_U357;
wire P1_R1165_U358 , P1_R1165_U359 , P1_R1165_U360 , P1_R1165_U361 , P1_R1165_U362 , P1_R1165_U363 , P1_R1165_U364 , P1_R1165_U365 , P1_R1165_U366 , P1_R1165_U367;
wire P1_R1165_U368 , P1_R1165_U369 , P1_R1165_U370 , P1_R1165_U371 , P1_R1165_U372 , P1_R1165_U373 , P1_R1165_U374 , P1_R1165_U375 , P1_R1165_U376 , P1_R1165_U377;
wire P1_R1165_U378 , P1_R1165_U379 , P1_R1165_U380 , P1_R1165_U381 , P1_R1165_U382 , P1_R1165_U383 , P1_R1165_U384 , P1_R1165_U385 , P1_R1165_U386 , P1_R1165_U387;
wire P1_R1165_U388 , P1_R1165_U389 , P1_R1165_U390 , P1_R1165_U391 , P1_R1165_U392 , P1_R1165_U393 , P1_R1165_U394 , P1_R1165_U395 , P1_R1165_U396 , P1_R1165_U397;
wire P1_R1165_U398 , P1_R1165_U399 , P1_R1165_U400 , P1_R1165_U401 , P1_R1165_U402 , P1_R1165_U403 , P1_R1165_U404 , P1_R1165_U405 , P1_R1165_U406 , P1_R1165_U407;
wire P1_R1165_U408 , P1_R1165_U409 , P1_R1165_U410 , P1_R1165_U411 , P1_R1165_U412 , P1_R1165_U413 , P1_R1165_U414 , P1_R1165_U415 , P1_R1165_U416 , P1_R1165_U417;
wire P1_R1165_U418 , P1_R1165_U419 , P1_R1165_U420 , P1_R1165_U421 , P1_R1165_U422 , P1_R1165_U423 , P1_R1165_U424 , P1_R1165_U425 , P1_R1165_U426 , P1_R1165_U427;
wire P1_R1165_U428 , P1_R1165_U429 , P1_R1165_U430 , P1_R1165_U431 , P1_R1165_U432 , P1_R1165_U433 , P1_R1165_U434 , P1_R1165_U435 , P1_R1165_U436 , P1_R1165_U437;
wire P1_R1165_U438 , P1_R1165_U439 , P1_R1165_U440 , P1_R1165_U441 , P1_R1165_U442 , P1_R1165_U443 , P1_R1165_U444 , P1_R1165_U445 , P1_R1165_U446 , P1_R1165_U447;
wire P1_R1165_U448 , P1_R1165_U449 , P1_R1165_U450 , P1_R1165_U451 , P1_R1165_U452 , P1_R1165_U453 , P1_R1165_U454 , P1_R1165_U455 , P1_R1165_U456 , P1_R1165_U457;
wire P1_R1165_U458 , P1_R1165_U459 , P1_R1165_U460 , P1_R1165_U461 , P1_R1165_U462 , P1_R1165_U463 , P1_R1165_U464 , P1_R1165_U465 , P1_R1165_U466 , P1_R1165_U467;
wire P1_R1165_U468 , P1_R1165_U469 , P1_R1165_U470 , P1_R1165_U471 , P1_R1165_U472 , P1_R1165_U473 , P1_R1165_U474 , P1_R1165_U475 , P1_R1165_U476 , P1_R1165_U477;
wire P1_R1165_U478 , P1_R1165_U479 , P1_R1165_U480 , P1_R1165_U481 , P1_R1165_U482 , P1_R1165_U483 , P1_R1165_U484 , P1_R1165_U485 , P1_R1165_U486 , P1_R1165_U487;
wire P1_R1165_U488 , P1_R1165_U489 , P1_R1165_U490 , P1_R1165_U491 , P1_R1165_U492 , P1_R1165_U493 , P1_R1165_U494 , P1_R1165_U495 , P1_R1165_U496 , P1_R1165_U497;
wire P1_R1165_U498 , P1_R1165_U499 , P1_R1165_U500 , P1_R1165_U501 , P1_R1165_U502 , P1_R1165_U503 , P1_R1165_U504 , P1_R1165_U505 , P1_R1165_U506 , P1_R1165_U507;
wire P1_R1165_U508 , P1_R1165_U509 , P1_R1165_U510 , P1_R1165_U511 , P1_R1165_U512 , P1_R1165_U513 , P1_R1165_U514 , P1_R1165_U515 , P1_R1165_U516 , P1_R1165_U517;
wire P1_R1165_U518 , P1_R1165_U519 , P1_R1165_U520 , P1_R1165_U521 , P1_R1165_U522 , P1_R1165_U523 , P1_R1165_U524 , P1_R1165_U525 , P1_R1165_U526 , P1_R1165_U527;
wire P1_R1165_U528 , P1_R1165_U529 , P1_R1165_U530 , P1_R1165_U531 , P1_R1165_U532 , P1_R1165_U533 , P1_R1165_U534 , P1_R1165_U535 , P1_R1165_U536 , P1_R1165_U537;
wire P1_R1165_U538 , P1_R1165_U539 , P1_R1165_U540 , P1_R1165_U541 , P1_R1165_U542 , P1_R1165_U543 , P1_R1165_U544 , P1_R1165_U545 , P1_R1165_U546 , P1_R1165_U547;
wire P1_R1165_U548 , P1_R1165_U549 , P1_R1165_U550 , P1_R1165_U551 , P1_R1165_U552 , P1_R1165_U553 , P1_R1165_U554 , P1_R1165_U555 , P1_R1165_U556 , P1_R1165_U557;
wire P1_R1165_U558 , P1_R1165_U559 , P1_R1165_U560 , P1_R1165_U561 , P1_R1165_U562 , P1_R1165_U563 , P1_R1165_U564 , P1_R1165_U565 , P1_R1165_U566 , P1_R1165_U567;
wire P1_R1165_U568 , P1_R1165_U569 , P1_R1165_U570 , P1_R1165_U571 , P1_R1165_U572 , P1_R1165_U573 , P1_R1165_U574 , P1_R1165_U575 , P1_R1165_U576 , P1_R1165_U577;
wire P1_R1165_U578 , P1_R1165_U579 , P1_R1165_U580 , P1_R1165_U581 , P1_R1165_U582 , P1_R1165_U583 , P1_R1165_U584 , P1_R1165_U585 , P1_R1165_U586 , P1_R1165_U587;
wire P1_R1165_U588 , P1_R1165_U589 , P1_R1165_U590 , P1_R1165_U591 , P1_R1165_U592 , P1_R1165_U593 , P1_R1165_U594 , P1_R1165_U595 , P1_R1165_U596 , P1_R1165_U597;
wire P1_R1165_U598 , P1_R1165_U599 , P1_R1165_U600 , P1_R1165_U601 , P1_R1165_U602 , P1_R1150_U6 , P1_R1150_U7 , P1_R1150_U8 , P1_R1150_U9 , P1_R1150_U10;
wire P1_R1150_U11 , P1_R1150_U12 , P1_R1150_U13 , P1_R1150_U14 , P1_R1150_U15 , P1_R1150_U16 , P1_R1150_U17 , P1_R1150_U18 , P1_R1150_U19 , P1_R1150_U20;
wire P1_R1150_U21 , P1_R1150_U22 , P1_R1150_U23 , P1_R1150_U24 , P1_R1150_U25 , P1_R1150_U26 , P1_R1150_U27 , P1_R1150_U28 , P1_R1150_U29 , P1_R1150_U30;
wire P1_R1150_U31 , P1_R1150_U32 , P1_R1150_U33 , P1_R1150_U34 , P1_R1150_U35 , P1_R1150_U36 , P1_R1150_U37 , P1_R1150_U38 , P1_R1150_U39 , P1_R1150_U40;
wire P1_R1150_U41 , P1_R1150_U42 , P1_R1150_U43 , P1_R1150_U44 , P1_R1150_U45 , P1_R1150_U46 , P1_R1150_U47 , P1_R1150_U48 , P1_R1150_U49 , P1_R1150_U50;
wire P1_R1150_U51 , P1_R1150_U52 , P1_R1150_U53 , P1_R1150_U54 , P1_R1150_U55 , P1_R1150_U56 , P1_R1150_U57 , P1_R1150_U58 , P1_R1150_U59 , P1_R1150_U60;
wire P1_R1150_U61 , P1_R1150_U62 , P1_R1150_U63 , P1_R1150_U64 , P1_R1150_U65 , P1_R1150_U66 , P1_R1150_U67 , P1_R1150_U68 , P1_R1150_U69 , P1_R1150_U70;
wire P1_R1150_U71 , P1_R1150_U72 , P1_R1150_U73 , P1_R1150_U74 , P1_R1150_U75 , P1_R1150_U76 , P1_R1150_U77 , P1_R1150_U78 , P1_R1150_U79 , P1_R1150_U80;
wire P1_R1150_U81 , P1_R1150_U82 , P1_R1150_U83 , P1_R1150_U84 , P1_R1150_U85 , P1_R1150_U86 , P1_R1150_U87 , P1_R1150_U88 , P1_R1150_U89 , P1_R1150_U90;
wire P1_R1150_U91 , P1_R1150_U92 , P1_R1150_U93 , P1_R1150_U94 , P1_R1150_U95 , P1_R1150_U96 , P1_R1150_U97 , P1_R1150_U98 , P1_R1150_U99 , P1_R1150_U100;
wire P1_R1150_U101 , P1_R1150_U102 , P1_R1150_U103 , P1_R1150_U104 , P1_R1150_U105 , P1_R1150_U106 , P1_R1150_U107 , P1_R1150_U108 , P1_R1150_U109 , P1_R1150_U110;
wire P1_R1150_U111 , P1_R1150_U112 , P1_R1150_U113 , P1_R1150_U114 , P1_R1150_U115 , P1_R1150_U116 , P1_R1150_U117 , P1_R1150_U118 , P1_R1150_U119 , P1_R1150_U120;
wire P1_R1150_U121 , P1_R1150_U122 , P1_R1150_U123 , P1_R1150_U124 , P1_R1150_U125 , P1_R1150_U126 , P1_R1150_U127 , P1_R1150_U128 , P1_R1150_U129 , P1_R1150_U130;
wire P1_R1150_U131 , P1_R1150_U132 , P1_R1150_U133 , P1_R1150_U134 , P1_R1150_U135 , P1_R1150_U136 , P1_R1150_U137 , P1_R1150_U138 , P1_R1150_U139 , P1_R1150_U140;
wire P1_R1150_U141 , P1_R1150_U142 , P1_R1150_U143 , P1_R1150_U144 , P1_R1150_U145 , P1_R1150_U146 , P1_R1150_U147 , P1_R1150_U148 , P1_R1150_U149 , P1_R1150_U150;
wire P1_R1150_U151 , P1_R1150_U152 , P1_R1150_U153 , P1_R1150_U154 , P1_R1150_U155 , P1_R1150_U156 , P1_R1150_U157 , P1_R1150_U158 , P1_R1150_U159 , P1_R1150_U160;
wire P1_R1150_U161 , P1_R1150_U162 , P1_R1150_U163 , P1_R1150_U164 , P1_R1150_U165 , P1_R1150_U166 , P1_R1150_U167 , P1_R1150_U168 , P1_R1150_U169 , P1_R1150_U170;
wire P1_R1150_U171 , P1_R1150_U172 , P1_R1150_U173 , P1_R1150_U174 , P1_R1150_U175 , P1_R1150_U176 , P1_R1150_U177 , P1_R1150_U178 , P1_R1150_U179 , P1_R1150_U180;
wire P1_R1150_U181 , P1_R1150_U182 , P1_R1150_U183 , P1_R1150_U184 , P1_R1150_U185 , P1_R1150_U186 , P1_R1150_U187 , P1_R1150_U188 , P1_R1150_U189 , P1_R1150_U190;
wire P1_R1150_U191 , P1_R1150_U192 , P1_R1150_U193 , P1_R1150_U194 , P1_R1150_U195 , P1_R1150_U196 , P1_R1150_U197 , P1_R1150_U198 , P1_R1150_U199 , P1_R1150_U200;
wire P1_R1150_U201 , P1_R1150_U202 , P1_R1150_U203 , P1_R1150_U204 , P1_R1150_U205 , P1_R1150_U206 , P1_R1150_U207 , P1_R1150_U208 , P1_R1150_U209 , P1_R1150_U210;
wire P1_R1150_U211 , P1_R1150_U212 , P1_R1150_U213 , P1_R1150_U214 , P1_R1150_U215 , P1_R1150_U216 , P1_R1150_U217 , P1_R1150_U218 , P1_R1150_U219 , P1_R1150_U220;
wire P1_R1150_U221 , P1_R1150_U222 , P1_R1150_U223 , P1_R1150_U224 , P1_R1150_U225 , P1_R1150_U226 , P1_R1150_U227 , P1_R1150_U228 , P1_R1150_U229 , P1_R1150_U230;
wire P1_R1150_U231 , P1_R1150_U232 , P1_R1150_U233 , P1_R1150_U234 , P1_R1150_U235 , P1_R1150_U236 , P1_R1150_U237 , P1_R1150_U238 , P1_R1150_U239 , P1_R1150_U240;
wire P1_R1150_U241 , P1_R1150_U242 , P1_R1150_U243 , P1_R1150_U244 , P1_R1150_U245 , P1_R1150_U246 , P1_R1150_U247 , P1_R1150_U248 , P1_R1150_U249 , P1_R1150_U250;
wire P1_R1150_U251 , P1_R1150_U252 , P1_R1150_U253 , P1_R1150_U254 , P1_R1150_U255 , P1_R1150_U256 , P1_R1150_U257 , P1_R1150_U258 , P1_R1150_U259 , P1_R1150_U260;
wire P1_R1150_U261 , P1_R1150_U262 , P1_R1150_U263 , P1_R1150_U264 , P1_R1150_U265 , P1_R1150_U266 , P1_R1150_U267 , P1_R1150_U268 , P1_R1150_U269 , P1_R1150_U270;
wire P1_R1150_U271 , P1_R1150_U272 , P1_R1150_U273 , P1_R1150_U274 , P1_R1150_U275 , P1_R1150_U276 , P1_R1150_U277 , P1_R1150_U278 , P1_R1150_U279 , P1_R1150_U280;
wire P1_R1150_U281 , P1_R1150_U282 , P1_R1150_U283 , P1_R1150_U284 , P1_R1150_U285 , P1_R1150_U286 , P1_R1150_U287 , P1_R1150_U288 , P1_R1150_U289 , P1_R1150_U290;
wire P1_R1150_U291 , P1_R1150_U292 , P1_R1150_U293 , P1_R1150_U294 , P1_R1150_U295 , P1_R1150_U296 , P1_R1150_U297 , P1_R1150_U298 , P1_R1150_U299 , P1_R1150_U300;
wire P1_R1150_U301 , P1_R1150_U302 , P1_R1150_U303 , P1_R1150_U304 , P1_R1150_U305 , P1_R1150_U306 , P1_R1150_U307 , P1_R1150_U308 , P1_R1150_U309 , P1_R1150_U310;
wire P1_R1150_U311 , P1_R1150_U312 , P1_R1150_U313 , P1_R1150_U314 , P1_R1150_U315 , P1_R1150_U316 , P1_R1150_U317 , P1_R1150_U318 , P1_R1150_U319 , P1_R1150_U320;
wire P1_R1150_U321 , P1_R1150_U322 , P1_R1150_U323 , P1_R1150_U324 , P1_R1150_U325 , P1_R1150_U326 , P1_R1150_U327 , P1_R1150_U328 , P1_R1150_U329 , P1_R1150_U330;
wire P1_R1150_U331 , P1_R1150_U332 , P1_R1150_U333 , P1_R1150_U334 , P1_R1150_U335 , P1_R1150_U336 , P1_R1150_U337 , P1_R1150_U338 , P1_R1150_U339 , P1_R1150_U340;
wire P1_R1150_U341 , P1_R1150_U342 , P1_R1150_U343 , P1_R1150_U344 , P1_R1150_U345 , P1_R1150_U346 , P1_R1150_U347 , P1_R1150_U348 , P1_R1150_U349 , P1_R1150_U350;
wire P1_R1150_U351 , P1_R1150_U352 , P1_R1150_U353 , P1_R1150_U354 , P1_R1150_U355 , P1_R1150_U356 , P1_R1150_U357 , P1_R1150_U358 , P1_R1150_U359 , P1_R1150_U360;
wire P1_R1150_U361 , P1_R1150_U362 , P1_R1150_U363 , P1_R1150_U364 , P1_R1150_U365 , P1_R1150_U366 , P1_R1150_U367 , P1_R1150_U368 , P1_R1150_U369 , P1_R1150_U370;
wire P1_R1150_U371 , P1_R1150_U372 , P1_R1150_U373 , P1_R1150_U374 , P1_R1150_U375 , P1_R1150_U376 , P1_R1150_U377 , P1_R1150_U378 , P1_R1150_U379 , P1_R1150_U380;
wire P1_R1150_U381 , P1_R1150_U382 , P1_R1150_U383 , P1_R1150_U384 , P1_R1150_U385 , P1_R1150_U386 , P1_R1150_U387 , P1_R1150_U388 , P1_R1150_U389 , P1_R1150_U390;
wire P1_R1150_U391 , P1_R1150_U392 , P1_R1150_U393 , P1_R1150_U394 , P1_R1150_U395 , P1_R1150_U396 , P1_R1150_U397 , P1_R1150_U398 , P1_R1150_U399 , P1_R1150_U400;
wire P1_R1150_U401 , P1_R1150_U402 , P1_R1150_U403 , P1_R1150_U404 , P1_R1150_U405 , P1_R1150_U406 , P1_R1150_U407 , P1_R1150_U408 , P1_R1150_U409 , P1_R1150_U410;
wire P1_R1150_U411 , P1_R1150_U412 , P1_R1150_U413 , P1_R1150_U414 , P1_R1150_U415 , P1_R1150_U416 , P1_R1150_U417 , P1_R1150_U418 , P1_R1150_U419 , P1_R1150_U420;
wire P1_R1150_U421 , P1_R1150_U422 , P1_R1150_U423 , P1_R1150_U424 , P1_R1150_U425 , P1_R1150_U426 , P1_R1150_U427 , P1_R1150_U428 , P1_R1150_U429 , P1_R1150_U430;
wire P1_R1150_U431 , P1_R1150_U432 , P1_R1150_U433 , P1_R1150_U434 , P1_R1150_U435 , P1_R1150_U436 , P1_R1150_U437 , P1_R1150_U438 , P1_R1150_U439 , P1_R1150_U440;
wire P1_R1150_U441 , P1_R1150_U442 , P1_R1150_U443 , P1_R1150_U444 , P1_R1150_U445 , P1_R1150_U446 , P1_R1150_U447 , P1_R1150_U448 , P1_R1150_U449 , P1_R1150_U450;
wire P1_R1150_U451 , P1_R1150_U452 , P1_R1150_U453 , P1_R1150_U454 , P1_R1150_U455 , P1_R1150_U456 , P1_R1150_U457 , P1_R1150_U458 , P1_R1150_U459 , P1_R1150_U460;
wire P1_R1150_U461 , P1_R1150_U462 , P1_R1150_U463 , P1_R1150_U464 , P1_R1150_U465 , P1_R1150_U466 , P1_R1150_U467 , P1_R1150_U468 , P1_R1150_U469 , P1_R1150_U470;
wire P1_R1150_U471 , P1_R1150_U472 , P1_R1150_U473 , P1_R1150_U474 , P1_R1150_U475 , P1_R1150_U476 , P1_R1192_U6 , P1_R1192_U7 , P1_R1192_U8 , P1_R1192_U9;
wire P1_R1192_U10 , P1_R1192_U11 , P1_R1192_U12 , P1_R1192_U13 , P1_R1192_U14 , P1_R1192_U15 , P1_R1192_U16 , P1_R1192_U17 , P1_R1192_U18 , P1_R1192_U19;
wire P1_R1192_U20 , P1_R1192_U21 , P1_R1192_U22 , P1_R1192_U23 , P1_R1192_U24 , P1_R1192_U25 , P1_R1192_U26 , P1_R1192_U27 , P1_R1192_U28 , P1_R1192_U29;
wire P1_R1192_U30 , P1_R1192_U31 , P1_R1192_U32 , P1_R1192_U33 , P1_R1192_U34 , P1_R1192_U35 , P1_R1192_U36 , P1_R1192_U37 , P1_R1192_U38 , P1_R1192_U39;
wire P1_R1192_U40 , P1_R1192_U41 , P1_R1192_U42 , P1_R1192_U43 , P1_R1192_U44 , P1_R1192_U45 , P1_R1192_U46 , P1_R1192_U47 , P1_R1192_U48 , P1_R1192_U49;
wire P1_R1192_U50 , P1_R1192_U51 , P1_R1192_U52 , P1_R1192_U53 , P1_R1192_U54 , P1_R1192_U55 , P1_R1192_U56 , P1_R1192_U57 , P1_R1192_U58 , P1_R1192_U59;
wire P1_R1192_U60 , P1_R1192_U61 , P1_R1192_U62 , P1_R1192_U63 , P1_R1192_U64 , P1_R1192_U65 , P1_R1192_U66 , P1_R1192_U67 , P1_R1192_U68 , P1_R1192_U69;
wire P1_R1192_U70 , P1_R1192_U71 , P1_R1192_U72 , P1_R1192_U73 , P1_R1192_U74 , P1_R1192_U75 , P1_R1192_U76 , P1_R1192_U77 , P1_R1192_U78 , P1_R1192_U79;
wire P1_R1192_U80 , P1_R1192_U81 , P1_R1192_U82 , P1_R1192_U83 , P1_R1192_U84 , P1_R1192_U85 , P1_R1192_U86 , P1_R1192_U87 , P1_R1192_U88 , P1_R1192_U89;
wire P1_R1192_U90 , P1_R1192_U91 , P1_R1192_U92 , P1_R1192_U93 , P1_R1192_U94 , P1_R1192_U95 , P1_R1192_U96 , P1_R1192_U97 , P1_R1192_U98 , P1_R1192_U99;
wire P1_R1192_U100 , P1_R1192_U101 , P1_R1192_U102 , P1_R1192_U103 , P1_R1192_U104 , P1_R1192_U105 , P1_R1192_U106 , P1_R1192_U107 , P1_R1192_U108 , P1_R1192_U109;
wire P1_R1192_U110 , P1_R1192_U111 , P1_R1192_U112 , P1_R1192_U113 , P1_R1192_U114 , P1_R1192_U115 , P1_R1192_U116 , P1_R1192_U117 , P1_R1192_U118 , P1_R1192_U119;
wire P1_R1192_U120 , P1_R1192_U121 , P1_R1192_U122 , P1_R1192_U123 , P1_R1192_U124 , P1_R1192_U125 , P1_R1192_U126 , P1_R1192_U127 , P1_R1192_U128 , P1_R1192_U129;
wire P1_R1192_U130 , P1_R1192_U131 , P1_R1192_U132 , P1_R1192_U133 , P1_R1192_U134 , P1_R1192_U135 , P1_R1192_U136 , P1_R1192_U137 , P1_R1192_U138 , P1_R1192_U139;
wire P1_R1192_U140 , P1_R1192_U141 , P1_R1192_U142 , P1_R1192_U143 , P1_R1192_U144 , P1_R1192_U145 , P1_R1192_U146 , P1_R1192_U147 , P1_R1192_U148 , P1_R1192_U149;
wire P1_R1192_U150 , P1_R1192_U151 , P1_R1192_U152 , P1_R1192_U153 , P1_R1192_U154 , P1_R1192_U155 , P1_R1192_U156 , P1_R1192_U157 , P1_R1192_U158 , P1_R1192_U159;
wire P1_R1192_U160 , P1_R1192_U161 , P1_R1192_U162 , P1_R1192_U163 , P1_R1192_U164 , P1_R1192_U165 , P1_R1192_U166 , P1_R1192_U167 , P1_R1192_U168 , P1_R1192_U169;
wire P1_R1192_U170 , P1_R1192_U171 , P1_R1192_U172 , P1_R1192_U173 , P1_R1192_U174 , P1_R1192_U175 , P1_R1192_U176 , P1_R1192_U177 , P1_R1192_U178 , P1_R1192_U179;
wire P1_R1192_U180 , P1_R1192_U181 , P1_R1192_U182 , P1_R1192_U183 , P1_R1192_U184 , P1_R1192_U185 , P1_R1192_U186 , P1_R1192_U187 , P1_R1192_U188 , P1_R1192_U189;
wire P1_R1192_U190 , P1_R1192_U191 , P1_R1192_U192 , P1_R1192_U193 , P1_R1192_U194 , P1_R1192_U195 , P1_R1192_U196 , P1_R1192_U197 , P1_R1192_U198 , P1_R1192_U199;
wire P1_R1192_U200 , P1_R1192_U201 , P1_R1192_U202 , P1_R1192_U203 , P1_R1192_U204 , P1_R1192_U205 , P1_R1192_U206 , P1_R1192_U207 , P1_R1192_U208 , P1_R1192_U209;
wire P1_R1192_U210 , P1_R1192_U211 , P1_R1192_U212 , P1_R1192_U213 , P1_R1192_U214 , P1_R1192_U215 , P1_R1192_U216 , P1_R1192_U217 , P1_R1192_U218 , P1_R1192_U219;
wire P1_R1192_U220 , P1_R1192_U221 , P1_R1192_U222 , P1_R1192_U223 , P1_R1192_U224 , P1_R1192_U225 , P1_R1192_U226 , P1_R1192_U227 , P1_R1192_U228 , P1_R1192_U229;
wire P1_R1192_U230 , P1_R1192_U231 , P1_R1192_U232 , P1_R1192_U233 , P1_R1192_U234 , P1_R1192_U235 , P1_R1192_U236 , P1_R1192_U237 , P1_R1192_U238 , P1_R1192_U239;
wire P1_R1192_U240 , P1_R1192_U241 , P1_R1192_U242 , P1_R1192_U243 , P1_R1192_U244 , P1_R1192_U245 , P1_R1192_U246 , P1_R1192_U247 , P1_R1192_U248 , P1_R1192_U249;
wire P1_R1192_U250 , P1_R1192_U251 , P1_R1192_U252 , P1_R1192_U253 , P1_R1192_U254 , P1_R1192_U255 , P1_R1192_U256 , P1_R1192_U257 , P1_R1192_U258 , P1_R1192_U259;
wire P1_R1192_U260 , P1_R1192_U261 , P1_R1192_U262 , P1_R1192_U263 , P1_R1192_U264 , P1_R1192_U265 , P1_R1192_U266 , P1_R1192_U267 , P1_R1192_U268 , P1_R1192_U269;
wire P1_R1192_U270 , P1_R1192_U271 , P1_R1192_U272 , P1_R1192_U273 , P1_R1192_U274 , P1_R1192_U275 , P1_R1192_U276 , P1_R1192_U277 , P1_R1192_U278 , P1_R1192_U279;
wire P1_R1192_U280 , P1_R1192_U281 , P1_R1192_U282 , P1_R1192_U283 , P1_R1192_U284 , P1_R1192_U285 , P1_R1192_U286 , P1_R1192_U287 , P1_R1192_U288 , P1_R1192_U289;
wire P1_R1192_U290 , P1_R1192_U291 , P1_R1192_U292 , P1_R1192_U293 , P1_R1192_U294 , P1_R1192_U295 , P1_R1192_U296 , P1_R1192_U297 , P1_R1192_U298 , P1_R1192_U299;
wire P1_R1192_U300 , P1_R1192_U301 , P1_R1192_U302 , P1_R1192_U303 , P1_R1192_U304 , P1_R1192_U305 , P1_R1192_U306 , P1_R1192_U307 , P1_R1192_U308 , P1_R1192_U309;
wire P1_R1192_U310 , P1_R1192_U311 , P1_R1192_U312 , P1_R1192_U313 , P1_R1192_U314 , P1_R1192_U315 , P1_R1192_U316 , P1_R1192_U317 , P1_R1192_U318 , P1_R1192_U319;
wire P1_R1192_U320 , P1_R1192_U321 , P1_R1192_U322 , P1_R1192_U323 , P1_R1192_U324 , P1_R1192_U325 , P1_R1192_U326 , P1_R1192_U327 , P1_R1192_U328 , P1_R1192_U329;
wire P1_R1192_U330 , P1_R1192_U331 , P1_R1192_U332 , P1_R1192_U333 , P1_R1192_U334 , P1_R1192_U335 , P1_R1192_U336 , P1_R1192_U337 , P1_R1192_U338 , P1_R1192_U339;
wire P1_R1192_U340 , P1_R1192_U341 , P1_R1192_U342 , P1_R1192_U343 , P1_R1192_U344 , P1_R1192_U345 , P1_R1192_U346 , P1_R1192_U347 , P1_R1192_U348 , P1_R1192_U349;
wire P1_R1192_U350 , P1_R1192_U351 , P1_R1192_U352 , P1_R1192_U353 , P1_R1192_U354 , P1_R1192_U355 , P1_R1192_U356 , P1_R1192_U357 , P1_R1192_U358 , P1_R1192_U359;
wire P1_R1192_U360 , P1_R1192_U361 , P1_R1192_U362 , P1_R1192_U363 , P1_R1192_U364 , P1_R1192_U365 , P1_R1192_U366 , P1_R1192_U367 , P1_R1192_U368 , P1_R1192_U369;
wire P1_R1192_U370 , P1_R1192_U371 , P1_R1192_U372 , P1_R1192_U373 , P1_R1192_U374 , P1_R1192_U375 , P1_R1192_U376 , P1_R1192_U377 , P1_R1192_U378 , P1_R1192_U379;
wire P1_R1192_U380 , P1_R1192_U381 , P1_R1192_U382 , P1_R1192_U383 , P1_R1192_U384 , P1_R1192_U385 , P1_R1192_U386 , P1_R1192_U387 , P1_R1192_U388 , P1_R1192_U389;
wire P1_R1192_U390 , P1_R1192_U391 , P1_R1192_U392 , P1_R1192_U393 , P1_R1192_U394 , P1_R1192_U395 , P1_R1192_U396 , P1_R1192_U397 , P1_R1192_U398 , P1_R1192_U399;
wire P1_R1192_U400 , P1_R1192_U401 , P1_R1192_U402 , P1_R1192_U403 , P1_R1192_U404 , P1_R1192_U405 , P1_R1192_U406 , P1_R1192_U407 , P1_R1192_U408 , P1_R1192_U409;
wire P1_R1192_U410 , P1_R1192_U411 , P1_R1192_U412 , P1_R1192_U413 , P1_R1192_U414 , P1_R1192_U415 , P1_R1192_U416 , P1_R1192_U417 , P1_R1192_U418 , P1_R1192_U419;
wire P1_R1192_U420 , P1_R1192_U421 , P1_R1192_U422 , P1_R1192_U423 , P1_R1192_U424 , P1_R1192_U425 , P1_R1192_U426 , P1_R1192_U427 , P1_R1192_U428 , P1_R1192_U429;
wire P1_R1192_U430 , P1_R1192_U431 , P1_R1192_U432 , P1_R1192_U433 , P1_R1192_U434 , P1_R1192_U435 , P1_R1192_U436 , P1_R1192_U437 , P1_R1192_U438 , P1_R1192_U439;
wire P1_R1192_U440 , P1_R1192_U441 , P1_R1192_U442 , P1_R1192_U443 , P1_R1192_U444 , P1_R1192_U445 , P1_R1192_U446 , P1_R1192_U447 , P1_R1192_U448 , P1_R1192_U449;
wire P1_R1192_U450 , P1_R1192_U451 , P1_R1192_U452 , P1_R1192_U453 , P1_R1192_U454 , P1_R1192_U455 , P1_R1192_U456 , P1_R1192_U457 , P1_R1192_U458 , P1_R1192_U459;
wire P1_R1192_U460 , P1_R1192_U461 , P1_R1192_U462 , P1_R1192_U463 , P1_R1192_U464 , P1_R1192_U465 , P1_R1192_U466 , P1_R1192_U467 , P1_R1192_U468 , P1_R1192_U469;
wire P1_R1192_U470 , P1_R1192_U471 , P1_R1192_U472 , P1_R1192_U473 , P1_R1192_U474 , P1_R1192_U475 , P1_R1192_U476 , P1_LT_201_U6 , P1_LT_201_U7 , P1_LT_201_U8;
wire P1_LT_201_U9 , P1_LT_201_U10 , P1_LT_201_U11 , P1_LT_201_U12 , P1_LT_201_U13 , P1_LT_201_U14 , P1_LT_201_U15 , P1_LT_201_U16 , P1_LT_201_U17 , P1_LT_201_U18;
wire P1_LT_201_U19 , P1_LT_201_U20 , P1_LT_201_U21 , P1_LT_201_U22 , P1_LT_201_U23 , P1_LT_201_U24 , P1_LT_201_U25 , P1_LT_201_U26 , P1_LT_201_U27 , P1_LT_201_U28;
wire P1_LT_201_U29 , P1_LT_201_U30 , P1_LT_201_U31 , P1_LT_201_U32 , P1_LT_201_U33 , P1_LT_201_U34 , P1_LT_201_U35 , P1_LT_201_U36 , P1_LT_201_U37 , P1_LT_201_U38;
wire P1_LT_201_U39 , P1_LT_201_U40 , P1_LT_201_U41 , P1_LT_201_U42 , P1_LT_201_U43 , P1_LT_201_U44 , P1_LT_201_U45 , P1_LT_201_U46 , P1_LT_201_U47 , P1_LT_201_U48;
wire P1_LT_201_U49 , P1_LT_201_U50 , P1_LT_201_U51 , P1_LT_201_U52 , P1_LT_201_U53 , P1_LT_201_U54 , P1_LT_201_U55 , P1_LT_201_U56 , P1_LT_201_U57 , P1_LT_201_U58;
wire P1_LT_201_U59 , P1_LT_201_U60 , P1_LT_201_U61 , P1_LT_201_U62 , P1_LT_201_U63 , P1_LT_201_U64 , P1_LT_201_U65 , P1_LT_201_U66 , P1_LT_201_U67 , P1_LT_201_U68;
wire P1_LT_201_U69 , P1_LT_201_U70 , P1_LT_201_U71 , P1_LT_201_U72 , P1_LT_201_U73 , P1_LT_201_U74 , P1_LT_201_U75 , P1_LT_201_U76 , P1_LT_201_U77 , P1_LT_201_U78;
wire P1_LT_201_U79 , P1_LT_201_U80 , P1_LT_201_U81 , P1_LT_201_U82 , P1_LT_201_U83 , P1_LT_201_U84 , P1_LT_201_U85 , P1_LT_201_U86 , P1_LT_201_U87 , P1_LT_201_U88;
wire P1_LT_201_U89 , P1_LT_201_U90 , P1_LT_201_U91 , P1_LT_201_U92 , P1_LT_201_U93 , P1_LT_201_U94 , P1_LT_201_U95 , P1_LT_201_U96 , P1_LT_201_U97 , P1_LT_201_U98;
wire P1_LT_201_U99 , P1_LT_201_U100 , P1_LT_201_U101 , P1_LT_201_U102 , P1_LT_201_U103 , P1_LT_201_U104 , P1_LT_201_U105 , P1_LT_201_U106 , P1_LT_201_U107 , P1_LT_201_U108;
wire P1_LT_201_U109 , P1_LT_201_U110 , P1_LT_201_U111 , P1_LT_201_U112 , P1_LT_201_U113 , P1_LT_201_U114 , P1_LT_201_U115 , P1_LT_201_U116 , P1_LT_201_U117 , P1_LT_201_U118;
wire P1_LT_201_U119 , P1_LT_201_U120 , P1_LT_201_U121 , P1_LT_201_U122 , P1_LT_201_U123 , P1_LT_201_U124 , P1_LT_201_U125 , P1_LT_201_U126 , P1_LT_201_U127 , P1_LT_201_U128;
wire P1_LT_201_U129 , P1_LT_201_U130 , P1_LT_201_U131 , P1_LT_201_U132 , P1_LT_201_U133 , P1_LT_201_U134 , P1_LT_201_U135 , P1_LT_201_U136 , P1_LT_201_U137 , P1_LT_201_U138;
wire P1_LT_201_U139 , P1_LT_201_U140 , P1_LT_201_U141 , P1_LT_201_U142 , P1_LT_201_U143 , P1_LT_201_U144 , P1_LT_201_U145 , P1_LT_201_U146 , P1_LT_201_U147 , P1_LT_201_U148;
wire P1_LT_201_U149 , P1_LT_201_U150 , P1_LT_201_U151 , P1_LT_201_U152 , P1_LT_201_U153 , P1_LT_201_U154 , P1_LT_201_U155 , P1_LT_201_U156 , P1_LT_201_U157 , P1_LT_201_U158;
wire P1_LT_201_U159 , P1_LT_201_U160 , P1_LT_201_U161 , P1_LT_201_U162 , P1_LT_201_U163 , P1_LT_201_U164 , P1_LT_201_U165 , P1_LT_201_U166 , P1_LT_201_U167 , P1_LT_201_U168;
wire P1_LT_201_U169 , P1_LT_201_U170 , P1_LT_201_U171 , P1_LT_201_U172 , P1_LT_201_U173 , P1_LT_201_U174 , P1_LT_201_U175 , P1_LT_201_U176 , P1_LT_201_U177 , P1_LT_201_U178;
wire P1_LT_201_U179 , P1_LT_201_U180 , P1_LT_201_U181 , P1_LT_201_U182 , P1_LT_201_U183 , P1_LT_201_U184 , P1_LT_201_U185 , P1_LT_201_U186 , P1_LT_201_U187 , P1_LT_201_U188;
wire P1_LT_201_U189 , P1_LT_201_U190 , P1_LT_201_U191 , P1_LT_201_U192 , P1_LT_201_U193 , P1_LT_201_U194 , P1_LT_201_U195 , P1_LT_201_U196 , P1_LT_201_U197 , P1_LT_201_U198;
wire P1_R1360_U6 , P1_R1360_U7 , P1_R1360_U8 , P1_R1360_U9 , P1_R1360_U10 , P1_R1360_U11 , P1_R1360_U12 , P1_R1360_U13 , P1_R1360_U14 , P1_R1360_U15;
wire P1_R1360_U16 , P1_R1360_U17 , P1_R1360_U18 , P1_R1360_U19 , P1_R1360_U20 , P1_R1360_U21 , P1_R1360_U22 , P1_R1360_U23 , P1_R1360_U24 , P1_R1360_U25;
wire P1_R1360_U26 , P1_R1360_U27 , P1_R1360_U28 , P1_R1360_U29 , P1_R1360_U30 , P1_R1360_U31 , P1_R1360_U32 , P1_R1360_U33 , P1_R1360_U34 , P1_R1360_U35;
wire P1_R1360_U36 , P1_R1360_U37 , P1_R1360_U38 , P1_R1360_U39 , P1_R1360_U40 , P1_R1360_U41 , P1_R1360_U42 , P1_R1360_U43 , P1_R1360_U44 , P1_R1360_U45;
wire P1_R1360_U46 , P1_R1360_U47 , P1_R1360_U48 , P1_R1360_U49 , P1_R1360_U50 , P1_R1360_U51 , P1_R1360_U52 , P1_R1360_U53 , P1_R1360_U54 , P1_R1360_U55;
wire P1_R1360_U56 , P1_R1360_U57 , P1_R1360_U58 , P1_R1360_U59 , P1_R1360_U60 , P1_R1360_U61 , P1_R1360_U62 , P1_R1360_U63 , P1_R1360_U64 , P1_R1360_U65;
wire P1_R1360_U66 , P1_R1360_U67 , P1_R1360_U68 , P1_R1360_U69 , P1_R1360_U70 , P1_R1360_U71 , P1_R1360_U72 , P1_R1360_U73 , P1_R1360_U74 , P1_R1360_U75;
wire P1_R1360_U76 , P1_R1360_U77 , P1_R1360_U78 , P1_R1360_U79 , P1_R1360_U80 , P1_R1360_U81 , P1_R1360_U82 , P1_R1360_U83 , P1_R1360_U84 , P1_R1360_U85;
wire P1_R1360_U86 , P1_R1360_U87 , P1_R1360_U88 , P1_R1360_U89 , P1_R1360_U90 , P1_R1360_U91 , P1_R1360_U92 , P1_R1360_U93 , P1_R1360_U94 , P1_R1360_U95;
wire P1_R1360_U96 , P1_R1360_U97 , P1_R1360_U98 , P1_R1360_U99 , P1_R1360_U100 , P1_R1360_U101 , P1_R1360_U102 , P1_R1360_U103 , P1_R1360_U104 , P1_R1360_U105;
wire P1_R1360_U106 , P1_R1360_U107 , P1_R1360_U108 , P1_R1360_U109 , P1_R1360_U110 , P1_R1360_U111 , P1_R1360_U112 , P1_R1360_U113 , P1_R1360_U114 , P1_R1360_U115;
wire P1_R1360_U116 , P1_R1360_U117 , P1_R1360_U118 , P1_R1360_U119 , P1_R1360_U120 , P1_R1360_U121 , P1_R1360_U122 , P1_R1360_U123 , P1_R1360_U124 , P1_R1360_U125;
wire P1_R1360_U126 , P1_R1360_U127 , P1_R1360_U128 , P1_R1360_U129 , P1_R1360_U130 , P1_R1360_U131 , P1_R1360_U132 , P1_R1360_U133 , P1_R1360_U134 , P1_R1360_U135;
wire P1_R1360_U136 , P1_R1360_U137 , P1_R1360_U138 , P1_R1360_U139 , P1_R1360_U140 , P1_R1360_U141 , P1_R1360_U142 , P1_R1360_U143 , P1_R1360_U144 , P1_R1360_U145;
wire P1_R1360_U146 , P1_R1360_U147 , P1_R1360_U148 , P1_R1360_U149 , P1_R1360_U150 , P1_R1360_U151 , P1_R1360_U152 , P1_R1360_U153 , P1_R1360_U154 , P1_R1360_U155;
wire P1_R1360_U156 , P1_R1360_U157 , P1_R1360_U158 , P1_R1360_U159 , P1_R1360_U160 , P1_R1360_U161 , P1_R1360_U162 , P1_R1360_U163 , P1_R1360_U164 , P1_R1360_U165;
wire P1_R1360_U166 , P1_R1360_U167 , P1_R1360_U168 , P1_R1360_U169 , P1_R1360_U170 , P1_R1360_U171 , P1_R1360_U172 , P1_R1360_U173 , P1_R1360_U174 , P1_R1360_U175;
wire P1_R1360_U176 , P1_R1360_U177 , P1_R1360_U178 , P1_R1360_U179 , P1_R1360_U180 , P1_R1360_U181 , P1_R1360_U182 , P1_R1360_U183 , P1_R1360_U184 , P1_R1360_U185;
wire P1_R1360_U186 , P1_R1360_U187 , P1_R1360_U188 , P1_R1360_U189 , P1_R1360_U190 , P1_R1360_U191 , P1_R1360_U192 , P1_R1360_U193 , P1_R1360_U194 , P1_R1360_U195;
wire P1_R1360_U196 , P1_R1360_U197 , P1_R1360_U198 , P1_R1360_U199 , P1_R1360_U200 , P1_R1360_U201 , P1_R1360_U202 , P1_R1360_U203 , P1_R1360_U204 , P1_R1360_U205;
wire P1_R1171_U4 , P1_R1171_U5 , P1_R1171_U6 , P1_R1171_U7 , P1_R1171_U8 , P1_R1171_U9 , P1_R1171_U10 , P1_R1171_U11 , P1_R1171_U12 , P1_R1171_U13;
wire P1_R1171_U14 , P1_R1171_U15 , P1_R1171_U16 , P1_R1171_U17 , P1_R1171_U18 , P1_R1171_U19 , P1_R1171_U20 , P1_R1171_U21 , P1_R1171_U22 , P1_R1171_U23;
wire P1_R1171_U24 , P1_R1171_U25 , P1_R1171_U26 , P1_R1171_U27 , P1_R1171_U28 , P1_R1171_U29 , P1_R1171_U30 , P1_R1171_U31 , P1_R1171_U32 , P1_R1171_U33;
wire P1_R1171_U34 , P1_R1171_U35 , P1_R1171_U36 , P1_R1171_U37 , P1_R1171_U38 , P1_R1171_U39 , P1_R1171_U40 , P1_R1171_U41 , P1_R1171_U42 , P1_R1171_U43;
wire P1_R1171_U44 , P1_R1171_U45 , P1_R1171_U46 , P1_R1171_U47 , P1_R1171_U48 , P1_R1171_U49 , P1_R1171_U50 , P1_R1171_U51 , P1_R1171_U52 , P1_R1171_U53;
wire P1_R1171_U54 , P1_R1171_U55 , P1_R1171_U56 , P1_R1171_U57 , P1_R1171_U58 , P1_R1171_U59 , P1_R1171_U60 , P1_R1171_U61 , P1_R1171_U62 , P1_R1171_U63;
wire P1_R1171_U64 , P1_R1171_U65 , P1_R1171_U66 , P1_R1171_U67 , P1_R1171_U68 , P1_R1171_U69 , P1_R1171_U70 , P1_R1171_U71 , P1_R1171_U72 , P1_R1171_U73;
wire P1_R1171_U74 , P1_R1171_U75 , P1_R1171_U76 , P1_R1171_U77 , P1_R1171_U78 , P1_R1171_U79 , P1_R1171_U80 , P1_R1171_U81 , P1_R1171_U82 , P1_R1171_U83;
wire P1_R1171_U84 , P1_R1171_U85 , P1_R1171_U86 , P1_R1171_U87 , P1_R1171_U88 , P1_R1171_U89 , P1_R1171_U90 , P1_R1171_U91 , P1_R1171_U92 , P1_R1171_U93;
wire P1_R1171_U94 , P1_R1171_U95 , P1_R1171_U96 , P1_R1171_U97 , P1_R1171_U98 , P1_R1171_U99 , P1_R1171_U100 , P1_R1171_U101 , P1_R1171_U102 , P1_R1171_U103;
wire P1_R1171_U104 , P1_R1171_U105 , P1_R1171_U106 , P1_R1171_U107 , P1_R1171_U108 , P1_R1171_U109 , P1_R1171_U110 , P1_R1171_U111 , P1_R1171_U112 , P1_R1171_U113;
wire P1_R1171_U114 , P1_R1171_U115 , P1_R1171_U116 , P1_R1171_U117 , P1_R1171_U118 , P1_R1171_U119 , P1_R1171_U120 , P1_R1171_U121 , P1_R1171_U122 , P1_R1171_U123;
wire P1_R1171_U124 , P1_R1171_U125 , P1_R1171_U126 , P1_R1171_U127 , P1_R1171_U128 , P1_R1171_U129 , P1_R1171_U130 , P1_R1171_U131 , P1_R1171_U132 , P1_R1171_U133;
wire P1_R1171_U134 , P1_R1171_U135 , P1_R1171_U136 , P1_R1171_U137 , P1_R1171_U138 , P1_R1171_U139 , P1_R1171_U140 , P1_R1171_U141 , P1_R1171_U142 , P1_R1171_U143;
wire P1_R1171_U144 , P1_R1171_U145 , P1_R1171_U146 , P1_R1171_U147 , P1_R1171_U148 , P1_R1171_U149 , P1_R1171_U150 , P1_R1171_U151 , P1_R1171_U152 , P1_R1171_U153;
wire P1_R1171_U154 , P1_R1171_U155 , P1_R1171_U156 , P1_R1171_U157 , P1_R1171_U158 , P1_R1171_U159 , P1_R1171_U160 , P1_R1171_U161 , P1_R1171_U162 , P1_R1171_U163;
wire P1_R1171_U164 , P1_R1171_U165 , P1_R1171_U166 , P1_R1171_U167 , P1_R1171_U168 , P1_R1171_U169 , P1_R1171_U170 , P1_R1171_U171 , P1_R1171_U172 , P1_R1171_U173;
wire P1_R1171_U174 , P1_R1171_U175 , P1_R1171_U176 , P1_R1171_U177 , P1_R1171_U178 , P1_R1171_U179 , P1_R1171_U180 , P1_R1171_U181 , P1_R1171_U182 , P1_R1171_U183;
wire P1_R1171_U184 , P1_R1171_U185 , P1_R1171_U186 , P1_R1171_U187 , P1_R1171_U188 , P1_R1171_U189 , P1_R1171_U190 , P1_R1171_U191 , P1_R1171_U192 , P1_R1171_U193;
wire P1_R1171_U194 , P1_R1171_U195 , P1_R1171_U196 , P1_R1171_U197 , P1_R1171_U198 , P1_R1171_U199 , P1_R1171_U200 , P1_R1171_U201 , P1_R1171_U202 , P1_R1171_U203;
wire P1_R1171_U204 , P1_R1171_U205 , P1_R1171_U206 , P1_R1171_U207 , P1_R1171_U208 , P1_R1171_U209 , P1_R1171_U210 , P1_R1171_U211 , P1_R1171_U212 , P1_R1171_U213;
wire P1_R1171_U214 , P1_R1171_U215 , P1_R1171_U216 , P1_R1171_U217 , P1_R1171_U218 , P1_R1171_U219 , P1_R1171_U220 , P1_R1171_U221 , P1_R1171_U222 , P1_R1171_U223;
wire P1_R1171_U224 , P1_R1171_U225 , P1_R1171_U226 , P1_R1171_U227 , P1_R1171_U228 , P1_R1171_U229 , P1_R1171_U230 , P1_R1171_U231 , P1_R1171_U232 , P1_R1171_U233;
wire P1_R1171_U234 , P1_R1171_U235 , P1_R1171_U236 , P1_R1171_U237 , P1_R1171_U238 , P1_R1171_U239 , P1_R1171_U240 , P1_R1171_U241 , P1_R1171_U242 , P1_R1171_U243;
wire P1_R1171_U244 , P1_R1171_U245 , P1_R1171_U246 , P1_R1171_U247 , P1_R1171_U248 , P1_R1171_U249 , P1_R1171_U250 , P1_R1171_U251 , P1_R1171_U252 , P1_R1171_U253;
wire P1_R1171_U254 , P1_R1171_U255 , P1_R1171_U256 , P1_R1171_U257 , P1_R1171_U258 , P1_R1171_U259 , P1_R1171_U260 , P1_R1171_U261 , P1_R1171_U262 , P1_R1171_U263;
wire P1_R1171_U264 , P1_R1171_U265 , P1_R1171_U266 , P1_R1171_U267 , P1_R1171_U268 , P1_R1171_U269 , P1_R1171_U270 , P1_R1171_U271 , P1_R1171_U272 , P1_R1171_U273;
wire P1_R1171_U274 , P1_R1171_U275 , P1_R1171_U276 , P1_R1171_U277 , P1_R1171_U278 , P1_R1171_U279 , P1_R1171_U280 , P1_R1171_U281 , P1_R1171_U282 , P1_R1171_U283;
wire P1_R1171_U284 , P1_R1171_U285 , P1_R1171_U286 , P1_R1171_U287 , P1_R1171_U288 , P1_R1171_U289 , P1_R1171_U290 , P1_R1171_U291 , P1_R1171_U292 , P1_R1171_U293;
wire P1_R1171_U294 , P1_R1171_U295 , P1_R1171_U296 , P1_R1171_U297 , P1_R1171_U298 , P1_R1171_U299 , P1_R1171_U300 , P1_R1171_U301 , P1_R1171_U302 , P1_R1171_U303;
wire P1_R1171_U304 , P1_R1171_U305 , P1_R1171_U306 , P1_R1171_U307 , P1_R1171_U308 , P1_R1171_U309 , P1_R1171_U310 , P1_R1171_U311 , P1_R1171_U312 , P1_R1171_U313;
wire P1_R1171_U314 , P1_R1171_U315 , P1_R1171_U316 , P1_R1171_U317 , P1_R1171_U318 , P1_R1171_U319 , P1_R1171_U320 , P1_R1171_U321 , P1_R1171_U322 , P1_R1171_U323;
wire P1_R1171_U324 , P1_R1171_U325 , P1_R1171_U326 , P1_R1171_U327 , P1_R1171_U328 , P1_R1171_U329 , P1_R1171_U330 , P1_R1171_U331 , P1_R1171_U332 , P1_R1171_U333;
wire P1_R1171_U334 , P1_R1171_U335 , P1_R1171_U336 , P1_R1171_U337 , P1_R1171_U338 , P1_R1171_U339 , P1_R1171_U340 , P1_R1171_U341 , P1_R1171_U342 , P1_R1171_U343;
wire P1_R1171_U344 , P1_R1171_U345 , P1_R1171_U346 , P1_R1171_U347 , P1_R1171_U348 , P1_R1171_U349 , P1_R1171_U350 , P1_R1171_U351 , P1_R1171_U352 , P1_R1171_U353;
wire P1_R1171_U354 , P1_R1171_U355 , P1_R1171_U356 , P1_R1171_U357 , P1_R1171_U358 , P1_R1171_U359 , P1_R1171_U360 , P1_R1171_U361 , P1_R1171_U362 , P1_R1171_U363;
wire P1_R1171_U364 , P1_R1171_U365 , P1_R1171_U366 , P1_R1171_U367 , P1_R1171_U368 , P1_R1171_U369 , P1_R1171_U370 , P1_R1171_U371 , P1_R1171_U372 , P1_R1171_U373;
wire P1_R1171_U374 , P1_R1171_U375 , P1_R1171_U376 , P1_R1171_U377 , P1_R1171_U378 , P1_R1171_U379 , P1_R1171_U380 , P1_R1171_U381 , P1_R1171_U382 , P1_R1171_U383;
wire P1_R1171_U384 , P1_R1171_U385 , P1_R1171_U386 , P1_R1171_U387 , P1_R1171_U388 , P1_R1171_U389 , P1_R1171_U390 , P1_R1171_U391 , P1_R1171_U392 , P1_R1171_U393;
wire P1_R1171_U394 , P1_R1171_U395 , P1_R1171_U396 , P1_R1171_U397 , P1_R1171_U398 , P1_R1171_U399 , P1_R1171_U400 , P1_R1171_U401 , P1_R1171_U402 , P1_R1171_U403;
wire P1_R1171_U404 , P1_R1171_U405 , P1_R1171_U406 , P1_R1171_U407 , P1_R1171_U408 , P1_R1171_U409 , P1_R1171_U410 , P1_R1171_U411 , P1_R1171_U412 , P1_R1171_U413;
wire P1_R1171_U414 , P1_R1171_U415 , P1_R1171_U416 , P1_R1171_U417 , P1_R1171_U418 , P1_R1171_U419 , P1_R1171_U420 , P1_R1171_U421 , P1_R1171_U422 , P1_R1171_U423;
wire P1_R1171_U424 , P1_R1171_U425 , P1_R1171_U426 , P1_R1171_U427 , P1_R1171_U428 , P1_R1171_U429 , P1_R1171_U430 , P1_R1171_U431 , P1_R1171_U432 , P1_R1171_U433;
wire P1_R1171_U434 , P1_R1171_U435 , P1_R1171_U436 , P1_R1171_U437 , P1_R1171_U438 , P1_R1171_U439 , P1_R1171_U440 , P1_R1171_U441 , P1_R1171_U442 , P1_R1171_U443;
wire P1_R1171_U444 , P1_R1171_U445 , P1_R1171_U446 , P1_R1171_U447 , P1_R1171_U448 , P1_R1171_U449 , P1_R1171_U450 , P1_R1171_U451 , P1_R1171_U452 , P1_R1171_U453;
wire P1_R1171_U454 , P1_R1171_U455 , P1_R1171_U456 , P1_R1171_U457 , P1_R1171_U458 , P1_R1171_U459 , P1_R1171_U460 , P1_R1171_U461 , P1_R1171_U462 , P1_R1171_U463;
wire P1_R1171_U464 , P1_R1171_U465 , P1_R1171_U466 , P1_R1171_U467 , P1_R1171_U468 , P1_R1171_U469 , P1_R1171_U470 , P1_R1171_U471 , P1_R1171_U472 , P1_R1171_U473;
wire P1_R1171_U474 , P1_R1171_U475 , P1_R1171_U476 , P1_R1171_U477 , P1_R1171_U478 , P1_R1171_U479 , P1_R1171_U480 , P1_R1171_U481 , P1_R1171_U482 , P1_R1171_U483;
wire P1_R1171_U484 , P1_R1171_U485 , P1_R1171_U486 , P1_R1171_U487 , P1_R1171_U488 , P1_R1171_U489 , P1_R1171_U490 , P1_R1171_U491 , P1_R1171_U492 , P1_R1171_U493;
wire P1_R1171_U494 , P1_R1171_U495 , P1_R1171_U496 , P1_R1171_U497 , P1_R1171_U498 , P1_R1171_U499 , P1_R1171_U500 , P1_R1171_U501 , P1_R1138_U4 , P1_R1138_U5;
wire P1_R1138_U6 , P1_R1138_U7 , P1_R1138_U8 , P1_R1138_U9 , P1_R1138_U10 , P1_R1138_U11 , P1_R1138_U12 , P1_R1138_U13 , P1_R1138_U14 , P1_R1138_U15;
wire P1_R1138_U16 , P1_R1138_U17 , P1_R1138_U18 , P1_R1138_U19 , P1_R1138_U20 , P1_R1138_U21 , P1_R1138_U22 , P1_R1138_U23 , P1_R1138_U24 , P1_R1138_U25;
wire P1_R1138_U26 , P1_R1138_U27 , P1_R1138_U28 , P1_R1138_U29 , P1_R1138_U30 , P1_R1138_U31 , P1_R1138_U32 , P1_R1138_U33 , P1_R1138_U34 , P1_R1138_U35;
wire P1_R1138_U36 , P1_R1138_U37 , P1_R1138_U38 , P1_R1138_U39 , P1_R1138_U40 , P1_R1138_U41 , P1_R1138_U42 , P1_R1138_U43 , P1_R1138_U44 , P1_R1138_U45;
wire P1_R1138_U46 , P1_R1138_U47 , P1_R1138_U48 , P1_R1138_U49 , P1_R1138_U50 , P1_R1138_U51 , P1_R1138_U52 , P1_R1138_U53 , P1_R1138_U54 , P1_R1138_U55;
wire P1_R1138_U56 , P1_R1138_U57 , P1_R1138_U58 , P1_R1138_U59 , P1_R1138_U60 , P1_R1138_U61 , P1_R1138_U62 , P1_R1138_U63 , P1_R1138_U64 , P1_R1138_U65;
wire P1_R1138_U66 , P1_R1138_U67 , P1_R1138_U68 , P1_R1138_U69 , P1_R1138_U70 , P1_R1138_U71 , P1_R1138_U72 , P1_R1138_U73 , P1_R1138_U74 , P1_R1138_U75;
wire P1_R1138_U76 , P1_R1138_U77 , P1_R1138_U78 , P1_R1138_U79 , P1_R1138_U80 , P1_R1138_U81 , P1_R1138_U82 , P1_R1138_U83 , P1_R1138_U84 , P1_R1138_U85;
wire P1_R1138_U86 , P1_R1138_U87 , P1_R1138_U88 , P1_R1138_U89 , P1_R1138_U90 , P1_R1138_U91 , P1_R1138_U92 , P1_R1138_U93 , P1_R1138_U94 , P1_R1138_U95;
wire P1_R1138_U96 , P1_R1138_U97 , P1_R1138_U98 , P1_R1138_U99 , P1_R1138_U100 , P1_R1138_U101 , P1_R1138_U102 , P1_R1138_U103 , P1_R1138_U104 , P1_R1138_U105;
wire P1_R1138_U106 , P1_R1138_U107 , P1_R1138_U108 , P1_R1138_U109 , P1_R1138_U110 , P1_R1138_U111 , P1_R1138_U112 , P1_R1138_U113 , P1_R1138_U114 , P1_R1138_U115;
wire P1_R1138_U116 , P1_R1138_U117 , P1_R1138_U118 , P1_R1138_U119 , P1_R1138_U120 , P1_R1138_U121 , P1_R1138_U122 , P1_R1138_U123 , P1_R1138_U124 , P1_R1138_U125;
wire P1_R1138_U126 , P1_R1138_U127 , P1_R1138_U128 , P1_R1138_U129 , P1_R1138_U130 , P1_R1138_U131 , P1_R1138_U132 , P1_R1138_U133 , P1_R1138_U134 , P1_R1138_U135;
wire P1_R1138_U136 , P1_R1138_U137 , P1_R1138_U138 , P1_R1138_U139 , P1_R1138_U140 , P1_R1138_U141 , P1_R1138_U142 , P1_R1138_U143 , P1_R1138_U144 , P1_R1138_U145;
wire P1_R1138_U146 , P1_R1138_U147 , P1_R1138_U148 , P1_R1138_U149 , P1_R1138_U150 , P1_R1138_U151 , P1_R1138_U152 , P1_R1138_U153 , P1_R1138_U154 , P1_R1138_U155;
wire P1_R1138_U156 , P1_R1138_U157 , P1_R1138_U158 , P1_R1138_U159 , P1_R1138_U160 , P1_R1138_U161 , P1_R1138_U162 , P1_R1138_U163 , P1_R1138_U164 , P1_R1138_U165;
wire P1_R1138_U166 , P1_R1138_U167 , P1_R1138_U168 , P1_R1138_U169 , P1_R1138_U170 , P1_R1138_U171 , P1_R1138_U172 , P1_R1138_U173 , P1_R1138_U174 , P1_R1138_U175;
wire P1_R1138_U176 , P1_R1138_U177 , P1_R1138_U178 , P1_R1138_U179 , P1_R1138_U180 , P1_R1138_U181 , P1_R1138_U182 , P1_R1138_U183 , P1_R1138_U184 , P1_R1138_U185;
wire P1_R1138_U186 , P1_R1138_U187 , P1_R1138_U188 , P1_R1138_U189 , P1_R1138_U190 , P1_R1138_U191 , P1_R1138_U192 , P1_R1138_U193 , P1_R1138_U194 , P1_R1138_U195;
wire P1_R1138_U196 , P1_R1138_U197 , P1_R1138_U198 , P1_R1138_U199 , P1_R1138_U200 , P1_R1138_U201 , P1_R1138_U202 , P1_R1138_U203 , P1_R1138_U204 , P1_R1138_U205;
wire P1_R1138_U206 , P1_R1138_U207 , P1_R1138_U208 , P1_R1138_U209 , P1_R1138_U210 , P1_R1138_U211 , P1_R1138_U212 , P1_R1138_U213 , P1_R1138_U214 , P1_R1138_U215;
wire P1_R1138_U216 , P1_R1138_U217 , P1_R1138_U218 , P1_R1138_U219 , P1_R1138_U220 , P1_R1138_U221 , P1_R1138_U222 , P1_R1138_U223 , P1_R1138_U224 , P1_R1138_U225;
wire P1_R1138_U226 , P1_R1138_U227 , P1_R1138_U228 , P1_R1138_U229 , P1_R1138_U230 , P1_R1138_U231 , P1_R1138_U232 , P1_R1138_U233 , P1_R1138_U234 , P1_R1138_U235;
wire P1_R1138_U236 , P1_R1138_U237 , P1_R1138_U238 , P1_R1138_U239 , P1_R1138_U240 , P1_R1138_U241 , P1_R1138_U242 , P1_R1138_U243 , P1_R1138_U244 , P1_R1138_U245;
wire P1_R1138_U246 , P1_R1138_U247 , P1_R1138_U248 , P1_R1138_U249 , P1_R1138_U250 , P1_R1138_U251 , P1_R1138_U252 , P1_R1138_U253 , P1_R1138_U254 , P1_R1138_U255;
wire P1_R1138_U256 , P1_R1138_U257 , P1_R1138_U258 , P1_R1138_U259 , P1_R1138_U260 , P1_R1138_U261 , P1_R1138_U262 , P1_R1138_U263 , P1_R1138_U264 , P1_R1138_U265;
wire P1_R1138_U266 , P1_R1138_U267 , P1_R1138_U268 , P1_R1138_U269 , P1_R1138_U270 , P1_R1138_U271 , P1_R1138_U272 , P1_R1138_U273 , P1_R1138_U274 , P1_R1138_U275;
wire P1_R1138_U276 , P1_R1138_U277 , P1_R1138_U278 , P1_R1138_U279 , P1_R1138_U280 , P1_R1138_U281 , P1_R1138_U282 , P1_R1138_U283 , P1_R1138_U284 , P1_R1138_U285;
wire P1_R1138_U286 , P1_R1138_U287 , P1_R1138_U288 , P1_R1138_U289 , P1_R1138_U290 , P1_R1138_U291 , P1_R1138_U292 , P1_R1138_U293 , P1_R1138_U294 , P1_R1138_U295;
wire P1_R1138_U296 , P1_R1138_U297 , P1_R1138_U298 , P1_R1138_U299 , P1_R1138_U300 , P1_R1138_U301 , P1_R1138_U302 , P1_R1138_U303 , P1_R1138_U304 , P1_R1138_U305;
wire P1_R1138_U306 , P1_R1138_U307 , P1_R1138_U308 , P1_R1138_U309 , P1_R1138_U310 , P1_R1138_U311 , P1_R1138_U312 , P1_R1138_U313 , P1_R1138_U314 , P1_R1138_U315;
wire P1_R1138_U316 , P1_R1138_U317 , P1_R1138_U318 , P1_R1138_U319 , P1_R1138_U320 , P1_R1138_U321 , P1_R1138_U322 , P1_R1138_U323 , P1_R1138_U324 , P1_R1138_U325;
wire P1_R1138_U326 , P1_R1138_U327 , P1_R1138_U328 , P1_R1138_U329 , P1_R1138_U330 , P1_R1138_U331 , P1_R1138_U332 , P1_R1138_U333 , P1_R1138_U334 , P1_R1138_U335;
wire P1_R1138_U336 , P1_R1138_U337 , P1_R1138_U338 , P1_R1138_U339 , P1_R1138_U340 , P1_R1138_U341 , P1_R1138_U342 , P1_R1138_U343 , P1_R1138_U344 , P1_R1138_U345;
wire P1_R1138_U346 , P1_R1138_U347 , P1_R1138_U348 , P1_R1138_U349 , P1_R1138_U350 , P1_R1138_U351 , P1_R1138_U352 , P1_R1138_U353 , P1_R1138_U354 , P1_R1138_U355;
wire P1_R1138_U356 , P1_R1138_U357 , P1_R1138_U358 , P1_R1138_U359 , P1_R1138_U360 , P1_R1138_U361 , P1_R1138_U362 , P1_R1138_U363 , P1_R1138_U364 , P1_R1138_U365;
wire P1_R1138_U366 , P1_R1138_U367 , P1_R1138_U368 , P1_R1138_U369 , P1_R1138_U370 , P1_R1138_U371 , P1_R1138_U372 , P1_R1138_U373 , P1_R1138_U374 , P1_R1138_U375;
wire P1_R1138_U376 , P1_R1138_U377 , P1_R1138_U378 , P1_R1138_U379 , P1_R1138_U380 , P1_R1138_U381 , P1_R1138_U382 , P1_R1138_U383 , P1_R1138_U384 , P1_R1138_U385;
wire P1_R1138_U386 , P1_R1138_U387 , P1_R1138_U388 , P1_R1138_U389 , P1_R1138_U390 , P1_R1138_U391 , P1_R1138_U392 , P1_R1138_U393 , P1_R1138_U394 , P1_R1138_U395;
wire P1_R1138_U396 , P1_R1138_U397 , P1_R1138_U398 , P1_R1138_U399 , P1_R1138_U400 , P1_R1138_U401 , P1_R1138_U402 , P1_R1138_U403 , P1_R1138_U404 , P1_R1138_U405;
wire P1_R1138_U406 , P1_R1138_U407 , P1_R1138_U408 , P1_R1138_U409 , P1_R1138_U410 , P1_R1138_U411 , P1_R1138_U412 , P1_R1138_U413 , P1_R1138_U414 , P1_R1138_U415;
wire P1_R1138_U416 , P1_R1138_U417 , P1_R1138_U418 , P1_R1138_U419 , P1_R1138_U420 , P1_R1138_U421 , P1_R1138_U422 , P1_R1138_U423 , P1_R1138_U424 , P1_R1138_U425;
wire P1_R1138_U426 , P1_R1138_U427 , P1_R1138_U428 , P1_R1138_U429 , P1_R1138_U430 , P1_R1138_U431 , P1_R1138_U432 , P1_R1138_U433 , P1_R1138_U434 , P1_R1138_U435;
wire P1_R1138_U436 , P1_R1138_U437 , P1_R1138_U438 , P1_R1138_U439 , P1_R1138_U440 , P1_R1138_U441 , P1_R1138_U442 , P1_R1138_U443 , P1_R1138_U444 , P1_R1138_U445;
wire P1_R1138_U446 , P1_R1138_U447 , P1_R1138_U448 , P1_R1138_U449 , P1_R1138_U450 , P1_R1138_U451 , P1_R1138_U452 , P1_R1138_U453 , P1_R1138_U454 , P1_R1138_U455;
wire P1_R1138_U456 , P1_R1138_U457 , P1_R1138_U458 , P1_R1138_U459 , P1_R1138_U460 , P1_R1138_U461 , P1_R1138_U462 , P1_R1138_U463 , P1_R1138_U464 , P1_R1138_U465;
wire P1_R1138_U466 , P1_R1138_U467 , P1_R1138_U468 , P1_R1138_U469 , P1_R1138_U470 , P1_R1138_U471 , P1_R1138_U472 , P1_R1138_U473 , P1_R1138_U474 , P1_R1138_U475;
wire P1_R1138_U476 , P1_R1138_U477 , P1_R1138_U478 , P1_R1138_U479 , P1_R1138_U480 , P1_R1138_U481 , P1_R1138_U482 , P1_R1138_U483 , P1_R1138_U484 , P1_R1138_U485;
wire P1_R1138_U486 , P1_R1138_U487 , P1_R1138_U488 , P1_R1138_U489 , P1_R1138_U490 , P1_R1138_U491 , P1_R1138_U492 , P1_R1138_U493 , P1_R1138_U494 , P1_R1138_U495;
wire P1_R1138_U496 , P1_R1138_U497 , P1_R1138_U498 , P1_R1138_U499 , P1_R1138_U500 , P1_R1138_U501 , P1_R1222_U4 , P1_R1222_U5 , P1_R1222_U6 , P1_R1222_U7;
wire P1_R1222_U8 , P1_R1222_U9 , P1_R1222_U10 , P1_R1222_U11 , P1_R1222_U12 , P1_R1222_U13 , P1_R1222_U14 , P1_R1222_U15 , P1_R1222_U16 , P1_R1222_U17;
wire P1_R1222_U18 , P1_R1222_U19 , P1_R1222_U20 , P1_R1222_U21 , P1_R1222_U22 , P1_R1222_U23 , P1_R1222_U24 , P1_R1222_U25 , P1_R1222_U26 , P1_R1222_U27;
wire P1_R1222_U28 , P1_R1222_U29 , P1_R1222_U30 , P1_R1222_U31 , P1_R1222_U32 , P1_R1222_U33 , P1_R1222_U34 , P1_R1222_U35 , P1_R1222_U36 , P1_R1222_U37;
wire P1_R1222_U38 , P1_R1222_U39 , P1_R1222_U40 , P1_R1222_U41 , P1_R1222_U42 , P1_R1222_U43 , P1_R1222_U44 , P1_R1222_U45 , P1_R1222_U46 , P1_R1222_U47;
wire P1_R1222_U48 , P1_R1222_U49 , P1_R1222_U50 , P1_R1222_U51 , P1_R1222_U52 , P1_R1222_U53 , P1_R1222_U54 , P1_R1222_U55 , P1_R1222_U56 , P1_R1222_U57;
wire P1_R1222_U58 , P1_R1222_U59 , P1_R1222_U60 , P1_R1222_U61 , P1_R1222_U62 , P1_R1222_U63 , P1_R1222_U64 , P1_R1222_U65 , P1_R1222_U66 , P1_R1222_U67;
wire P1_R1222_U68 , P1_R1222_U69 , P1_R1222_U70 , P1_R1222_U71 , P1_R1222_U72 , P1_R1222_U73 , P1_R1222_U74 , P1_R1222_U75 , P1_R1222_U76 , P1_R1222_U77;
wire P1_R1222_U78 , P1_R1222_U79 , P1_R1222_U80 , P1_R1222_U81 , P1_R1222_U82 , P1_R1222_U83 , P1_R1222_U84 , P1_R1222_U85 , P1_R1222_U86 , P1_R1222_U87;
wire P1_R1222_U88 , P1_R1222_U89 , P1_R1222_U90 , P1_R1222_U91 , P1_R1222_U92 , P1_R1222_U93 , P1_R1222_U94 , P1_R1222_U95 , P1_R1222_U96 , P1_R1222_U97;
wire P1_R1222_U98 , P1_R1222_U99 , P1_R1222_U100 , P1_R1222_U101 , P1_R1222_U102 , P1_R1222_U103 , P1_R1222_U104 , P1_R1222_U105 , P1_R1222_U106 , P1_R1222_U107;
wire P1_R1222_U108 , P1_R1222_U109 , P1_R1222_U110 , P1_R1222_U111 , P1_R1222_U112 , P1_R1222_U113 , P1_R1222_U114 , P1_R1222_U115 , P1_R1222_U116 , P1_R1222_U117;
wire P1_R1222_U118 , P1_R1222_U119 , P1_R1222_U120 , P1_R1222_U121 , P1_R1222_U122 , P1_R1222_U123 , P1_R1222_U124 , P1_R1222_U125 , P1_R1222_U126 , P1_R1222_U127;
wire P1_R1222_U128 , P1_R1222_U129 , P1_R1222_U130 , P1_R1222_U131 , P1_R1222_U132 , P1_R1222_U133 , P1_R1222_U134 , P1_R1222_U135 , P1_R1222_U136 , P1_R1222_U137;
wire P1_R1222_U138 , P1_R1222_U139 , P1_R1222_U140 , P1_R1222_U141 , P1_R1222_U142 , P1_R1222_U143 , P1_R1222_U144 , P1_R1222_U145 , P1_R1222_U146 , P1_R1222_U147;
wire P1_R1222_U148 , P1_R1222_U149 , P1_R1222_U150 , P1_R1222_U151 , P1_R1222_U152 , P1_R1222_U153 , P1_R1222_U154 , P1_R1222_U155 , P1_R1222_U156 , P1_R1222_U157;
wire P1_R1222_U158 , P1_R1222_U159 , P1_R1222_U160 , P1_R1222_U161 , P1_R1222_U162 , P1_R1222_U163 , P1_R1222_U164 , P1_R1222_U165 , P1_R1222_U166 , P1_R1222_U167;
wire P1_R1222_U168 , P1_R1222_U169 , P1_R1222_U170 , P1_R1222_U171 , P1_R1222_U172 , P1_R1222_U173 , P1_R1222_U174 , P1_R1222_U175 , P1_R1222_U176 , P1_R1222_U177;
wire P1_R1222_U178 , P1_R1222_U179 , P1_R1222_U180 , P1_R1222_U181 , P1_R1222_U182 , P1_R1222_U183 , P1_R1222_U184 , P1_R1222_U185 , P1_R1222_U186 , P1_R1222_U187;
wire P1_R1222_U188 , P1_R1222_U189 , P1_R1222_U190 , P1_R1222_U191 , P1_R1222_U192 , P1_R1222_U193 , P1_R1222_U194 , P1_R1222_U195 , P1_R1222_U196 , P1_R1222_U197;
wire P1_R1222_U198 , P1_R1222_U199 , P1_R1222_U200 , P1_R1222_U201 , P1_R1222_U202 , P1_R1222_U203 , P1_R1222_U204 , P1_R1222_U205 , P1_R1222_U206 , P1_R1222_U207;
wire P1_R1222_U208 , P1_R1222_U209 , P1_R1222_U210 , P1_R1222_U211 , P1_R1222_U212 , P1_R1222_U213 , P1_R1222_U214 , P1_R1222_U215 , P1_R1222_U216 , P1_R1222_U217;
wire P1_R1222_U218 , P1_R1222_U219 , P1_R1222_U220 , P1_R1222_U221 , P1_R1222_U222 , P1_R1222_U223 , P1_R1222_U224 , P1_R1222_U225 , P1_R1222_U226 , P1_R1222_U227;
wire P1_R1222_U228 , P1_R1222_U229 , P1_R1222_U230 , P1_R1222_U231 , P1_R1222_U232 , P1_R1222_U233 , P1_R1222_U234 , P1_R1222_U235 , P1_R1222_U236 , P1_R1222_U237;
wire P1_R1222_U238 , P1_R1222_U239 , P1_R1222_U240 , P1_R1222_U241 , P1_R1222_U242 , P1_R1222_U243 , P1_R1222_U244 , P1_R1222_U245 , P1_R1222_U246 , P1_R1222_U247;
wire P1_R1222_U248 , P1_R1222_U249 , P1_R1222_U250 , P1_R1222_U251 , P1_R1222_U252 , P1_R1222_U253 , P1_R1222_U254 , P1_R1222_U255 , P1_R1222_U256 , P1_R1222_U257;
wire P1_R1222_U258 , P1_R1222_U259 , P1_R1222_U260 , P1_R1222_U261 , P1_R1222_U262 , P1_R1222_U263 , P1_R1222_U264 , P1_R1222_U265 , P1_R1222_U266 , P1_R1222_U267;
wire P1_R1222_U268 , P1_R1222_U269 , P1_R1222_U270 , P1_R1222_U271 , P1_R1222_U272 , P1_R1222_U273 , P1_R1222_U274 , P1_R1222_U275 , P1_R1222_U276 , P1_R1222_U277;
wire P1_R1222_U278 , P1_R1222_U279 , P1_R1222_U280 , P1_R1222_U281 , P1_R1222_U282 , P1_R1222_U283 , P1_R1222_U284 , P1_R1222_U285 , P1_R1222_U286 , P1_R1222_U287;
wire P1_R1222_U288 , P1_R1222_U289 , P1_R1222_U290 , P1_R1222_U291 , P1_R1222_U292 , P1_R1222_U293 , P1_R1222_U294 , P1_R1222_U295 , P1_R1222_U296 , P1_R1222_U297;
wire P1_R1222_U298 , P1_R1222_U299 , P1_R1222_U300 , P1_R1222_U301 , P1_R1222_U302 , P1_R1222_U303 , P1_R1222_U304 , P1_R1222_U305 , P1_R1222_U306 , P1_R1222_U307;
wire P1_R1222_U308 , P1_R1222_U309 , P1_R1222_U310 , P1_R1222_U311 , P1_R1222_U312 , P1_R1222_U313 , P1_R1222_U314 , P1_R1222_U315 , P1_R1222_U316 , P1_R1222_U317;
wire P1_R1222_U318 , P1_R1222_U319 , P1_R1222_U320 , P1_R1222_U321 , P1_R1222_U322 , P1_R1222_U323 , P1_R1222_U324 , P1_R1222_U325 , P1_R1222_U326 , P1_R1222_U327;
wire P1_R1222_U328 , P1_R1222_U329 , P1_R1222_U330 , P1_R1222_U331 , P1_R1222_U332 , P1_R1222_U333 , P1_R1222_U334 , P1_R1222_U335 , P1_R1222_U336 , P1_R1222_U337;
wire P1_R1222_U338 , P1_R1222_U339 , P1_R1222_U340 , P1_R1222_U341 , P1_R1222_U342 , P1_R1222_U343 , P1_R1222_U344 , P1_R1222_U345 , P1_R1222_U346 , P1_R1222_U347;
wire P1_R1222_U348 , P1_R1222_U349 , P1_R1222_U350 , P1_R1222_U351 , P1_R1222_U352 , P1_R1222_U353 , P1_R1222_U354 , P1_R1222_U355 , P1_R1222_U356 , P1_R1222_U357;
wire P1_R1222_U358 , P1_R1222_U359 , P1_R1222_U360 , P1_R1222_U361 , P1_R1222_U362 , P1_R1222_U363 , P1_R1222_U364 , P1_R1222_U365 , P1_R1222_U366 , P1_R1222_U367;
wire P1_R1222_U368 , P1_R1222_U369 , P1_R1222_U370 , P1_R1222_U371 , P1_R1222_U372 , P1_R1222_U373 , P1_R1222_U374 , P1_R1222_U375 , P1_R1222_U376 , P1_R1222_U377;
wire P1_R1222_U378 , P1_R1222_U379 , P1_R1222_U380 , P1_R1222_U381 , P1_R1222_U382 , P1_R1222_U383 , P1_R1222_U384 , P1_R1222_U385 , P1_R1222_U386 , P1_R1222_U387;
wire P1_R1222_U388 , P1_R1222_U389 , P1_R1222_U390 , P1_R1222_U391 , P1_R1222_U392 , P1_R1222_U393 , P1_R1222_U394 , P1_R1222_U395 , P1_R1222_U396 , P1_R1222_U397;
wire P1_R1222_U398 , P1_R1222_U399 , P1_R1222_U400 , P1_R1222_U401 , P1_R1222_U402 , P1_R1222_U403 , P1_R1222_U404 , P1_R1222_U405 , P1_R1222_U406 , P1_R1222_U407;
wire P1_R1222_U408 , P1_R1222_U409 , P1_R1222_U410 , P1_R1222_U411 , P1_R1222_U412 , P1_R1222_U413 , P1_R1222_U414 , P1_R1222_U415 , P1_R1222_U416 , P1_R1222_U417;
wire P1_R1222_U418 , P1_R1222_U419 , P1_R1222_U420 , P1_R1222_U421 , P1_R1222_U422 , P1_R1222_U423 , P1_R1222_U424 , P1_R1222_U425 , P1_R1222_U426 , P1_R1222_U427;
wire P1_R1222_U428 , P1_R1222_U429 , P1_R1222_U430 , P1_R1222_U431 , P1_R1222_U432 , P1_R1222_U433 , P1_R1222_U434 , P1_R1222_U435 , P1_R1222_U436 , P1_R1222_U437;
wire P1_R1222_U438 , P1_R1222_U439 , P1_R1222_U440 , P1_R1222_U441 , P1_R1222_U442 , P1_R1222_U443 , P1_R1222_U444 , P1_R1222_U445 , P1_R1222_U446 , P1_R1222_U447;
wire P1_R1222_U448 , P1_R1222_U449 , P1_R1222_U450 , P1_R1222_U451 , P1_R1222_U452 , P1_R1222_U453 , P1_R1222_U454 , P1_R1222_U455 , P1_R1222_U456 , P1_R1222_U457;
wire P1_R1222_U458 , P1_R1222_U459 , P1_R1222_U460 , P1_R1222_U461 , P1_R1222_U462 , P1_R1222_U463 , P1_R1222_U464 , P1_R1222_U465 , P1_R1222_U466 , P1_R1222_U467;
wire P1_R1222_U468 , P1_R1222_U469 , P1_R1222_U470 , P1_R1222_U471 , P1_R1222_U472 , P1_R1222_U473 , P1_R1222_U474 , P1_R1222_U475 , P1_R1222_U476 , P1_R1222_U477;
wire P1_R1222_U478 , P1_R1222_U479 , P1_R1222_U480 , P1_R1222_U481 , P1_R1222_U482 , P1_R1222_U483 , P1_R1222_U484 , P1_R1222_U485 , P1_R1222_U486 , P1_R1222_U487;
wire P1_R1222_U488 , P1_R1222_U489 , P1_R1222_U490 , P1_R1222_U491 , P1_R1222_U492 , P1_R1222_U493 , P1_R1222_U494 , P1_R1222_U495 , P1_R1222_U496 , P1_R1222_U497;
wire P1_R1222_U498 , P1_R1222_U499 , P1_R1222_U500 , P1_R1222_U501 , P2_ADD_609_U4 , P2_ADD_609_U5 , P2_ADD_609_U6 , P2_ADD_609_U7 , P2_ADD_609_U8 , P2_ADD_609_U9;
wire P2_ADD_609_U10 , P2_ADD_609_U11 , P2_ADD_609_U12 , P2_ADD_609_U13 , P2_ADD_609_U14 , P2_ADD_609_U15 , P2_ADD_609_U16 , P2_ADD_609_U17 , P2_ADD_609_U18 , P2_ADD_609_U19;
wire P2_ADD_609_U20 , P2_ADD_609_U21 , P2_ADD_609_U22 , P2_ADD_609_U23 , P2_ADD_609_U24 , P2_ADD_609_U25 , P2_ADD_609_U26 , P2_ADD_609_U27 , P2_ADD_609_U28 , P2_ADD_609_U29;
wire P2_ADD_609_U30 , P2_ADD_609_U31 , P2_ADD_609_U32 , P2_ADD_609_U33 , P2_ADD_609_U34 , P2_ADD_609_U35 , P2_ADD_609_U36 , P2_ADD_609_U37 , P2_ADD_609_U38 , P2_ADD_609_U39;
wire P2_ADD_609_U40 , P2_ADD_609_U41 , P2_ADD_609_U42 , P2_ADD_609_U43 , P2_ADD_609_U44 , P2_ADD_609_U45 , P2_ADD_609_U46 , P2_ADD_609_U47 , P2_ADD_609_U48 , P2_ADD_609_U49;
wire P2_ADD_609_U50 , P2_ADD_609_U51 , P2_ADD_609_U52 , P2_ADD_609_U53 , P2_ADD_609_U54 , P2_ADD_609_U55 , P2_ADD_609_U56 , P2_ADD_609_U57 , P2_ADD_609_U58 , P2_ADD_609_U59;
wire P2_ADD_609_U60 , P2_ADD_609_U61 , P2_ADD_609_U62 , P2_ADD_609_U63 , P2_ADD_609_U64 , P2_ADD_609_U65 , P2_ADD_609_U66 , P2_ADD_609_U67 , P2_ADD_609_U68 , P2_ADD_609_U69;
wire P2_ADD_609_U70 , P2_ADD_609_U71 , P2_ADD_609_U72 , P2_ADD_609_U73 , P2_ADD_609_U74 , P2_ADD_609_U75 , P2_ADD_609_U76 , P2_ADD_609_U77 , P2_ADD_609_U78 , P2_ADD_609_U79;
wire P2_ADD_609_U80 , P2_ADD_609_U81 , P2_ADD_609_U82 , P2_ADD_609_U83 , P2_ADD_609_U84 , P2_ADD_609_U85 , P2_ADD_609_U86 , P2_ADD_609_U87 , P2_ADD_609_U88 , P2_ADD_609_U89;
wire P2_ADD_609_U90 , P2_ADD_609_U91 , P2_ADD_609_U92 , P2_ADD_609_U93 , P2_ADD_609_U94 , P2_ADD_609_U95 , P2_ADD_609_U96 , P2_ADD_609_U97 , P2_ADD_609_U98 , P2_ADD_609_U99;
wire P2_ADD_609_U100 , P2_ADD_609_U101 , P2_ADD_609_U102 , P2_ADD_609_U103 , P2_ADD_609_U104 , P2_ADD_609_U105 , P2_ADD_609_U106 , P2_ADD_609_U107 , P2_ADD_609_U108 , P2_ADD_609_U109;
wire P2_ADD_609_U110 , P2_ADD_609_U111 , P2_ADD_609_U112 , P2_ADD_609_U113 , P2_ADD_609_U114 , P2_ADD_609_U115 , P2_ADD_609_U116 , P2_ADD_609_U117 , P2_ADD_609_U118 , P2_ADD_609_U119;
wire P2_ADD_609_U120 , P2_ADD_609_U121 , P2_ADD_609_U122 , P2_ADD_609_U123 , P2_ADD_609_U124 , P2_ADD_609_U125 , P2_ADD_609_U126 , P2_ADD_609_U127 , P2_ADD_609_U128 , P2_ADD_609_U129;
wire P2_ADD_609_U130 , P2_ADD_609_U131 , P2_ADD_609_U132 , P2_ADD_609_U133 , P2_ADD_609_U134 , P2_ADD_609_U135 , P2_ADD_609_U136 , P2_ADD_609_U137 , P2_ADD_609_U138 , P2_ADD_609_U139;
wire P2_ADD_609_U140 , P2_ADD_609_U141 , P2_ADD_609_U142 , P2_ADD_609_U143 , P2_ADD_609_U144 , P2_ADD_609_U145 , P2_ADD_609_U146 , P2_ADD_609_U147 , P2_ADD_609_U148 , P2_ADD_609_U149;
wire P2_ADD_609_U150 , P2_ADD_609_U151 , P2_ADD_609_U152 , P2_ADD_609_U153 , P2_ADD_609_U154 , P2_ADD_609_U155 , P2_ADD_609_U156 , P2_R1340_U6 , P2_R1340_U7 , P2_R1340_U8;
wire P2_R1340_U9 , P2_R1340_U10 , P2_R1340_U11 , P2_R1340_U12 , P2_R1340_U13 , P2_R1340_U14 , P2_R1340_U15 , P2_R1340_U16 , P2_R1340_U17 , P2_R1340_U18;
wire P2_R1340_U19 , P2_R1340_U20 , P2_R1340_U21 , P2_R1340_U22 , P2_R1340_U23 , P2_R1340_U24 , P2_R1340_U25 , P2_R1340_U26 , P2_R1340_U27 , P2_R1340_U28;
wire P2_R1340_U29 , P2_R1340_U30 , P2_R1340_U31 , P2_R1340_U32 , P2_R1340_U33 , P2_R1340_U34 , P2_R1340_U35 , P2_R1340_U36 , P2_R1340_U37 , P2_R1340_U38;
wire P2_R1340_U39 , P2_R1340_U40 , P2_R1340_U41 , P2_R1340_U42 , P2_R1340_U43 , P2_R1340_U44 , P2_R1340_U45 , P2_R1340_U46 , P2_R1340_U47 , P2_R1340_U48;
wire P2_R1340_U49 , P2_R1340_U50 , P2_R1340_U51 , P2_R1340_U52 , P2_R1340_U53 , P2_R1340_U54 , P2_R1340_U55 , P2_R1340_U56 , P2_R1340_U57 , P2_R1340_U58;
wire P2_R1340_U59 , P2_R1340_U60 , P2_R1340_U61 , P2_R1340_U62 , P2_R1340_U63 , P2_R1340_U64 , P2_R1340_U65 , P2_R1340_U66 , P2_R1340_U67 , P2_R1340_U68;
wire P2_R1340_U69 , P2_R1340_U70 , P2_R1340_U71 , P2_R1340_U72 , P2_R1340_U73 , P2_R1340_U74 , P2_R1340_U75 , P2_R1340_U76 , P2_R1340_U77 , P2_R1340_U78;
wire P2_R1340_U79 , P2_R1340_U80 , P2_R1340_U81 , P2_R1340_U82 , P2_R1340_U83 , P2_R1340_U84 , P2_R1340_U85 , P2_R1340_U86 , P2_R1340_U87 , P2_R1340_U88;
wire P2_R1340_U89 , P2_R1340_U90 , P2_R1340_U91 , P2_R1340_U92 , P2_R1340_U93 , P2_R1340_U94 , P2_R1340_U95 , P2_R1340_U96 , P2_R1340_U97 , P2_R1340_U98;
wire P2_R1340_U99 , P2_R1340_U100 , P2_R1340_U101 , P2_R1340_U102 , P2_R1340_U103 , P2_R1340_U104 , P2_R1340_U105 , P2_R1340_U106 , P2_R1340_U107 , P2_R1340_U108;
wire P2_R1340_U109 , P2_R1340_U110 , P2_R1340_U111 , P2_R1340_U112 , P2_R1340_U113 , P2_R1340_U114 , P2_R1340_U115 , P2_R1340_U116 , P2_R1340_U117 , P2_R1340_U118;
wire P2_R1340_U119 , P2_R1340_U120 , P2_R1340_U121 , P2_R1340_U122 , P2_R1340_U123 , P2_R1340_U124 , P2_R1340_U125 , P2_R1340_U126 , P2_R1340_U127 , P2_R1340_U128;
wire P2_R1340_U129 , P2_R1340_U130 , P2_R1340_U131 , P2_R1340_U132 , P2_R1340_U133 , P2_R1340_U134 , P2_R1340_U135 , P2_R1340_U136 , P2_R1340_U137 , P2_R1340_U138;
wire P2_R1340_U139 , P2_R1340_U140 , P2_R1340_U141 , P2_R1340_U142 , P2_R1340_U143 , P2_R1340_U144 , P2_R1340_U145 , P2_R1340_U146 , P2_R1340_U147 , P2_R1340_U148;
wire P2_R1340_U149 , P2_R1340_U150 , P2_R1340_U151 , P2_R1340_U152 , P2_R1340_U153 , P2_R1340_U154 , P2_R1340_U155 , P2_R1340_U156 , P2_R1340_U157 , P2_R1340_U158;
wire P2_R1340_U159 , P2_R1340_U160 , P2_R1340_U161 , P2_R1340_U162 , P2_R1340_U163 , P2_R1340_U164 , P2_R1340_U165 , P2_R1340_U166 , P2_R1340_U167 , P2_R1340_U168;
wire P2_R1340_U169 , P2_R1340_U170 , P2_R1340_U171 , P2_R1340_U172 , P2_R1340_U173 , P2_R1340_U174 , P2_R1340_U175 , P2_R1340_U176 , P2_R1340_U177 , P2_R1340_U178;
wire P2_R1340_U179 , P2_SUB_598_U6 , P2_SUB_598_U7 , P2_SUB_598_U8 , P2_SUB_598_U9 , P2_SUB_598_U10 , P2_SUB_598_U11 , P2_SUB_598_U12 , P2_SUB_598_U13 , P2_SUB_598_U14;
wire P2_SUB_598_U15 , P2_SUB_598_U16 , P2_SUB_598_U17 , P2_SUB_598_U18 , P2_SUB_598_U19 , P2_SUB_598_U20 , P2_SUB_598_U21 , P2_SUB_598_U22 , P2_SUB_598_U23 , P2_SUB_598_U24;
wire P2_SUB_598_U25 , P2_SUB_598_U26 , P2_SUB_598_U27 , P2_SUB_598_U28 , P2_SUB_598_U29 , P2_SUB_598_U30 , P2_SUB_598_U31 , P2_SUB_598_U32 , P2_SUB_598_U33 , P2_SUB_598_U34;
wire P2_SUB_598_U35 , P2_SUB_598_U36 , P2_SUB_598_U37 , P2_SUB_598_U38 , P2_SUB_598_U39 , P2_SUB_598_U40 , P2_SUB_598_U41 , P2_SUB_598_U42 , P2_SUB_598_U43 , P2_SUB_598_U44;
wire P2_SUB_598_U45 , P2_SUB_598_U46 , P2_SUB_598_U47 , P2_SUB_598_U48 , P2_SUB_598_U49 , P2_SUB_598_U50 , P2_SUB_598_U51 , P2_SUB_598_U52 , P2_SUB_598_U53 , P2_SUB_598_U54;
wire P2_SUB_598_U55 , P2_SUB_598_U56 , P2_SUB_598_U57 , P2_SUB_598_U58 , P2_SUB_598_U59 , P2_SUB_598_U60 , P2_SUB_598_U61 , P2_SUB_598_U62 , P2_SUB_598_U63 , P2_SUB_598_U64;
wire P2_SUB_598_U65 , P2_SUB_598_U66 , P2_SUB_598_U67 , P2_SUB_598_U68 , P2_SUB_598_U69 , P2_SUB_598_U70 , P2_SUB_598_U71 , P2_SUB_598_U72 , P2_SUB_598_U73 , P2_SUB_598_U74;
wire P2_SUB_598_U75 , P2_SUB_598_U76 , P2_SUB_598_U77 , P2_SUB_598_U78 , P2_SUB_598_U79 , P2_SUB_598_U80 , P2_SUB_598_U81 , P2_SUB_598_U82 , P2_SUB_598_U83 , P2_SUB_598_U84;
wire P2_SUB_598_U85 , P2_SUB_598_U86 , P2_SUB_598_U87 , P2_SUB_598_U88 , P2_SUB_598_U89 , P2_SUB_598_U90 , P2_SUB_598_U91 , P2_SUB_598_U92 , P2_SUB_598_U93 , P2_SUB_598_U94;
wire P2_SUB_598_U95 , P2_SUB_598_U96 , P2_SUB_598_U97 , P2_SUB_598_U98 , P2_SUB_598_U99 , P2_SUB_598_U100 , P2_SUB_598_U101 , P2_SUB_598_U102 , P2_SUB_598_U103 , P2_SUB_598_U104;
wire P2_SUB_598_U105 , P2_SUB_598_U106 , P2_SUB_598_U107 , P2_SUB_598_U108 , P2_SUB_598_U109 , P2_SUB_598_U110 , P2_SUB_598_U111 , P2_SUB_598_U112 , P2_SUB_598_U113 , P2_SUB_598_U114;
wire P2_SUB_598_U115 , P2_SUB_598_U116 , P2_SUB_598_U117 , P2_SUB_598_U118 , P2_SUB_598_U119 , P2_SUB_598_U120 , P2_SUB_598_U121 , P2_SUB_598_U122 , P2_SUB_598_U123 , P2_SUB_598_U124;
wire P2_SUB_598_U125 , P2_SUB_598_U126 , P2_SUB_598_U127 , P2_SUB_598_U128 , P2_SUB_598_U129 , P2_SUB_598_U130 , P2_SUB_598_U131 , P2_SUB_598_U132 , P2_SUB_598_U133 , P2_SUB_598_U134;
wire P2_SUB_598_U135 , P2_SUB_598_U136 , P2_SUB_598_U137 , P2_SUB_598_U138 , P2_SUB_598_U139 , P2_SUB_598_U140 , P2_SUB_598_U141 , P2_SUB_598_U142 , P2_SUB_598_U143 , P2_SUB_598_U144;
wire P2_SUB_598_U145 , P2_SUB_598_U146 , P2_SUB_598_U147 , P2_SUB_598_U148 , P2_SUB_598_U149 , P2_SUB_598_U150 , P2_SUB_598_U151 , P2_SUB_598_U152 , P2_SUB_598_U153 , P2_SUB_598_U154;
wire P2_SUB_598_U155 , P2_SUB_598_U156 , P2_SUB_598_U157 , P2_SUB_598_U158 , P2_SUB_598_U159 , P2_SUB_598_U160 , P2_SUB_598_U161 , P2_SUB_598_U162 , P2_SUB_598_U163 , P2_SUB_598_U164;
wire P2_SUB_598_U165 , P2_SUB_598_U166 , P2_SUB_598_U167 , P2_SUB_598_U168 , P2_SUB_598_U169 , P2_SUB_598_U170 , P2_SUB_598_U171 , P2_SUB_598_U172 , P2_SUB_598_U173 , P2_R1299_U6;
wire P2_R1299_U7 , P2_R1312_U6 , P2_R1312_U7 , P2_R1312_U8 , P2_R1312_U9 , P2_R1312_U10 , P2_R1312_U11 , P2_R1312_U12 , P2_R1312_U13 , P2_R1312_U14;
wire P2_R1312_U15 , P2_R1312_U16 , P2_R1312_U17 , P2_R1312_U18 , P2_R1312_U19 , P2_R1312_U20 , P2_R1312_U21 , P2_R1312_U22 , P2_R1312_U23 , P2_R1312_U24;
wire P2_R1312_U25 , P2_R1312_U26 , P2_R1312_U27 , P2_R1312_U28 , P2_R1312_U29 , P2_R1312_U30 , P2_R1312_U31 , P2_R1312_U32 , P2_R1312_U33 , P2_R1312_U34;
wire P2_R1312_U35 , P2_R1312_U36 , P2_R1312_U37 , P2_R1312_U38 , P2_R1312_U39 , P2_R1312_U40 , P2_R1312_U41 , P2_R1312_U42 , P2_R1312_U43 , P2_R1312_U44;
wire P2_R1312_U45 , P2_R1312_U46 , P2_R1312_U47 , P2_R1312_U48 , P2_R1312_U49 , P2_R1312_U50 , P2_R1312_U51 , P2_R1312_U52 , P2_R1312_U53 , P2_R1312_U54;
wire P2_R1312_U55 , P2_R1312_U56 , P2_R1312_U57 , P2_R1312_U58 , P2_R1312_U59 , P2_R1312_U60 , P2_R1312_U61 , P2_R1312_U62 , P2_R1312_U63 , P2_R1312_U64;
wire P2_R1312_U65 , P2_R1312_U66 , P2_R1312_U67 , P2_R1312_U68 , P2_R1312_U69 , P2_R1312_U70 , P2_R1312_U71 , P2_R1312_U72 , P2_R1312_U73 , P2_R1312_U74;
wire P2_R1312_U75 , P2_R1312_U76 , P2_R1312_U77 , P2_R1312_U78 , P2_R1312_U79 , P2_R1312_U80 , P2_R1312_U81 , P2_R1312_U82 , P2_R1312_U83 , P2_R1312_U84;
wire P2_R1312_U85 , P2_R1312_U86 , P2_R1312_U87 , P2_R1312_U88 , P2_R1312_U89 , P2_R1312_U90 , P2_R1312_U91 , P2_R1312_U92 , P2_R1312_U93 , P2_R1312_U94;
wire P2_R1312_U95 , P2_R1312_U96 , P2_R1312_U97 , P2_R1312_U98 , P2_R1312_U99 , P2_R1312_U100 , P2_R1312_U101 , P2_R1312_U102 , P2_R1312_U103 , P2_R1312_U104;
wire P2_R1312_U105 , P2_R1312_U106 , P2_R1312_U107 , P2_R1312_U108 , P2_R1312_U109 , P2_R1312_U110 , P2_R1312_U111 , P2_R1312_U112 , P2_R1312_U113 , P2_R1312_U114;
wire P2_R1312_U115 , P2_R1312_U116 , P2_R1312_U117 , P2_R1312_U118 , P2_R1312_U119 , P2_R1312_U120 , P2_R1312_U121 , P2_R1312_U122 , P2_R1312_U123 , P2_R1312_U124;
wire P2_R1312_U125 , P2_R1312_U126 , P2_R1312_U127 , P2_R1312_U128 , P2_R1312_U129 , P2_R1312_U130 , P2_R1312_U131 , P2_R1312_U132 , P2_R1312_U133 , P2_R1312_U134;
wire P2_R1312_U135 , P2_R1312_U136 , P2_R1312_U137 , P2_R1312_U138 , P2_R1312_U139 , P2_R1312_U140 , P2_R1312_U141 , P2_R1312_U142 , P2_R1312_U143 , P2_R1312_U144;
wire P2_R1312_U145 , P2_R1312_U146 , P2_R1312_U147 , P2_R1312_U148 , P2_R1312_U149 , P2_R1312_U150 , P2_R1312_U151 , P2_R1312_U152 , P2_R1312_U153 , P2_R1312_U154;
wire P2_R1312_U155 , P2_R1312_U156 , P2_R1312_U157 , P2_R1312_U158 , P2_R1312_U159 , P2_R1312_U160 , P2_R1312_U161 , P2_R1312_U162 , P2_R1312_U163 , P2_R1312_U164;
wire P2_R1312_U165 , P2_R1312_U166 , P2_R1312_U167 , P2_R1312_U168 , P2_R1312_U169 , P2_R1312_U170 , P2_R1312_U171 , P2_R1312_U172 , P2_R1312_U173 , P2_R1312_U174;
wire P2_R1312_U175 , P2_R1312_U176 , P2_R1312_U177 , P2_R1312_U178 , P2_R1312_U179 , P2_R1312_U180 , P2_R1312_U181 , P2_R1312_U182 , P2_R1312_U183 , P2_R1312_U184;
wire P2_R1312_U185 , P2_R1312_U186 , P2_R1312_U187 , P2_R1312_U188 , P2_R1312_U189 , P2_R1312_U190 , P2_R1312_U191 , P2_R1312_U192 , P2_R1312_U193 , P2_R1312_U194;
wire P2_R1312_U195 , P2_R1312_U196 , P2_R1312_U197 , P2_R1312_U198 , P2_R1312_U199 , P2_R1312_U200 , P2_R1312_U201 , P2_R1312_U202 , P2_R1312_U203 , P2_R1312_U204;
wire P2_R1312_U205 , P2_R1312_U206 , P2_R1312_U207 , P2_R1312_U208 , P2_R1312_U209 , P2_R1335_U6 , P2_R1335_U7 , P2_R1335_U8 , P2_R1335_U9 , P2_R1335_U10;
wire P2_R1209_U4 , P2_R1209_U5 , P2_R1209_U6 , P2_R1209_U7 , P2_R1209_U8 , P2_R1209_U9 , P2_R1209_U10 , P2_R1209_U11 , P2_R1209_U12 , P2_R1209_U13;
wire P2_R1209_U14 , P2_R1209_U15 , P2_R1209_U16 , P2_R1209_U17 , P2_R1209_U18 , P2_R1209_U19 , P2_R1209_U20 , P2_R1209_U21 , P2_R1209_U22 , P2_R1209_U23;
wire P2_R1209_U24 , P2_R1209_U25 , P2_R1209_U26 , P2_R1209_U27 , P2_R1209_U28 , P2_R1209_U29 , P2_R1209_U30 , P2_R1209_U31 , P2_R1209_U32 , P2_R1209_U33;
wire P2_R1209_U34 , P2_R1209_U35 , P2_R1209_U36 , P2_R1209_U37 , P2_R1209_U38 , P2_R1209_U39 , P2_R1209_U40 , P2_R1209_U41 , P2_R1209_U42 , P2_R1209_U43;
wire P2_R1209_U44 , P2_R1209_U45 , P2_R1209_U46 , P2_R1209_U47 , P2_R1209_U48 , P2_R1209_U49 , P2_R1209_U50 , P2_R1209_U51 , P2_R1209_U52 , P2_R1209_U53;
wire P2_R1209_U54 , P2_R1209_U55 , P2_R1209_U56 , P2_R1209_U57 , P2_R1209_U58 , P2_R1209_U59 , P2_R1209_U60 , P2_R1209_U61 , P2_R1209_U62 , P2_R1209_U63;
wire P2_R1209_U64 , P2_R1209_U65 , P2_R1209_U66 , P2_R1209_U67 , P2_R1209_U68 , P2_R1209_U69 , P2_R1209_U70 , P2_R1209_U71 , P2_R1209_U72 , P2_R1209_U73;
wire P2_R1209_U74 , P2_R1209_U75 , P2_R1209_U76 , P2_R1209_U77 , P2_R1209_U78 , P2_R1209_U79 , P2_R1209_U80 , P2_R1209_U81 , P2_R1209_U82 , P2_R1209_U83;
wire P2_R1209_U84 , P2_R1209_U85 , P2_R1209_U86 , P2_R1209_U87 , P2_R1209_U88 , P2_R1209_U89 , P2_R1209_U90 , P2_R1209_U91 , P2_R1209_U92 , P2_R1209_U93;
wire P2_R1209_U94 , P2_R1209_U95 , P2_R1209_U96 , P2_R1209_U97 , P2_R1209_U98 , P2_R1209_U99 , P2_R1209_U100 , P2_R1209_U101 , P2_R1209_U102 , P2_R1209_U103;
wire P2_R1209_U104 , P2_R1209_U105 , P2_R1209_U106 , P2_R1209_U107 , P2_R1209_U108 , P2_R1209_U109 , P2_R1209_U110 , P2_R1209_U111 , P2_R1209_U112 , P2_R1209_U113;
wire P2_R1209_U114 , P2_R1209_U115 , P2_R1209_U116 , P2_R1209_U117 , P2_R1209_U118 , P2_R1209_U119 , P2_R1209_U120 , P2_R1209_U121 , P2_R1209_U122 , P2_R1209_U123;
wire P2_R1209_U124 , P2_R1209_U125 , P2_R1209_U126 , P2_R1209_U127 , P2_R1209_U128 , P2_R1209_U129 , P2_R1209_U130 , P2_R1209_U131 , P2_R1209_U132 , P2_R1209_U133;
wire P2_R1209_U134 , P2_R1209_U135 , P2_R1209_U136 , P2_R1209_U137 , P2_R1209_U138 , P2_R1209_U139 , P2_R1209_U140 , P2_R1209_U141 , P2_R1209_U142 , P2_R1209_U143;
wire P2_R1209_U144 , P2_R1209_U145 , P2_R1209_U146 , P2_R1209_U147 , P2_R1209_U148 , P2_R1209_U149 , P2_R1209_U150 , P2_R1209_U151 , P2_R1209_U152 , P2_R1209_U153;
wire P2_R1209_U154 , P2_R1209_U155 , P2_R1209_U156 , P2_R1209_U157 , P2_R1209_U158 , P2_R1209_U159 , P2_R1209_U160 , P2_R1209_U161 , P2_R1209_U162 , P2_R1209_U163;
wire P2_R1209_U164 , P2_R1209_U165 , P2_R1209_U166 , P2_R1209_U167 , P2_R1209_U168 , P2_R1209_U169 , P2_R1209_U170 , P2_R1209_U171 , P2_R1209_U172 , P2_R1209_U173;
wire P2_R1209_U174 , P2_R1209_U175 , P2_R1209_U176 , P2_R1209_U177 , P2_R1209_U178 , P2_R1209_U179 , P2_R1209_U180 , P2_R1209_U181 , P2_R1209_U182 , P2_R1209_U183;
wire P2_R1209_U184 , P2_R1209_U185 , P2_R1209_U186 , P2_R1209_U187 , P2_R1209_U188 , P2_R1209_U189 , P2_R1209_U190 , P2_R1209_U191 , P2_R1209_U192 , P2_R1209_U193;
wire P2_R1209_U194 , P2_R1209_U195 , P2_R1209_U196 , P2_R1209_U197 , P2_R1209_U198 , P2_R1209_U199 , P2_R1209_U200 , P2_R1209_U201 , P2_R1209_U202 , P2_R1209_U203;
wire P2_R1209_U204 , P2_R1209_U205 , P2_R1209_U206 , P2_R1209_U207 , P2_R1209_U208 , P2_R1209_U209 , P2_R1209_U210 , P2_R1209_U211 , P2_R1209_U212 , P2_R1209_U213;
wire P2_R1209_U214 , P2_R1209_U215 , P2_R1209_U216 , P2_R1209_U217 , P2_R1209_U218 , P2_R1209_U219 , P2_R1209_U220 , P2_R1209_U221 , P2_R1209_U222 , P2_R1209_U223;
wire P2_R1209_U224 , P2_R1209_U225 , P2_R1209_U226 , P2_R1209_U227 , P2_R1209_U228 , P2_R1209_U229 , P2_R1209_U230 , P2_R1209_U231 , P2_R1209_U232 , P2_R1209_U233;
wire P2_R1209_U234 , P2_R1209_U235 , P2_R1209_U236 , P2_R1209_U237 , P2_R1209_U238 , P2_R1209_U239 , P2_R1209_U240 , P2_R1209_U241 , P2_R1209_U242 , P2_R1209_U243;
wire P2_R1209_U244 , P2_R1209_U245 , P2_R1209_U246 , P2_R1209_U247 , P2_R1209_U248 , P2_R1209_U249 , P2_R1209_U250 , P2_R1209_U251 , P2_R1209_U252 , P2_R1209_U253;
wire P2_R1209_U254 , P2_R1209_U255 , P2_R1209_U256 , P2_R1209_U257 , P2_R1209_U258 , P2_R1209_U259 , P2_R1209_U260 , P2_R1209_U261 , P2_R1209_U262 , P2_R1209_U263;
wire P2_R1209_U264 , P2_R1209_U265 , P2_R1209_U266 , P2_R1209_U267 , P2_R1209_U268 , P2_R1209_U269 , P2_R1209_U270 , P2_R1209_U271 , P2_R1209_U272 , P2_R1209_U273;
wire P2_R1209_U274 , P2_R1209_U275 , P2_R1209_U276 , P2_R1209_U277 , P2_R1209_U278 , P2_R1209_U279 , P2_R1209_U280 , P2_R1209_U281 , P2_R1209_U282 , P2_R1209_U283;
wire P2_R1209_U284 , P2_R1209_U285 , P2_R1209_U286 , P2_R1209_U287 , P2_R1209_U288 , P2_R1209_U289 , P2_R1209_U290 , P2_R1209_U291 , P2_R1209_U292 , P2_R1209_U293;
wire P2_R1209_U294 , P2_R1209_U295 , P2_R1209_U296 , P2_R1209_U297 , P2_R1209_U298 , P2_R1209_U299 , P2_R1209_U300 , P2_R1209_U301 , P2_R1209_U302 , P2_R1209_U303;
wire P2_R1209_U304 , P2_R1209_U305 , P2_R1209_U306 , P2_R1209_U307 , P2_R1209_U308 , P2_R1170_U4 , P2_R1170_U5 , P2_R1170_U6 , P2_R1170_U7 , P2_R1170_U8;
wire P2_R1170_U9 , P2_R1170_U10 , P2_R1170_U11 , P2_R1170_U12 , P2_R1170_U13 , P2_R1170_U14 , P2_R1170_U15 , P2_R1170_U16 , P2_R1170_U17 , P2_R1170_U18;
wire P2_R1170_U19 , P2_R1170_U20 , P2_R1170_U21 , P2_R1170_U22 , P2_R1170_U23 , P2_R1170_U24 , P2_R1170_U25 , P2_R1170_U26 , P2_R1170_U27 , P2_R1170_U28;
wire P2_R1170_U29 , P2_R1170_U30 , P2_R1170_U31 , P2_R1170_U32 , P2_R1170_U33 , P2_R1170_U34 , P2_R1170_U35 , P2_R1170_U36 , P2_R1170_U37 , P2_R1170_U38;
wire P2_R1170_U39 , P2_R1170_U40 , P2_R1170_U41 , P2_R1170_U42 , P2_R1170_U43 , P2_R1170_U44 , P2_R1170_U45 , P2_R1170_U46 , P2_R1170_U47 , P2_R1170_U48;
wire P2_R1170_U49 , P2_R1170_U50 , P2_R1170_U51 , P2_R1170_U52 , P2_R1170_U53 , P2_R1170_U54 , P2_R1170_U55 , P2_R1170_U56 , P2_R1170_U57 , P2_R1170_U58;
wire P2_R1170_U59 , P2_R1170_U60 , P2_R1170_U61 , P2_R1170_U62 , P2_R1170_U63 , P2_R1170_U64 , P2_R1170_U65 , P2_R1170_U66 , P2_R1170_U67 , P2_R1170_U68;
wire P2_R1170_U69 , P2_R1170_U70 , P2_R1170_U71 , P2_R1170_U72 , P2_R1170_U73 , P2_R1170_U74 , P2_R1170_U75 , P2_R1170_U76 , P2_R1170_U77 , P2_R1170_U78;
wire P2_R1170_U79 , P2_R1170_U80 , P2_R1170_U81 , P2_R1170_U82 , P2_R1170_U83 , P2_R1170_U84 , P2_R1170_U85 , P2_R1170_U86 , P2_R1170_U87 , P2_R1170_U88;
wire P2_R1170_U89 , P2_R1170_U90 , P2_R1170_U91 , P2_R1170_U92 , P2_R1170_U93 , P2_R1170_U94 , P2_R1170_U95 , P2_R1170_U96 , P2_R1170_U97 , P2_R1170_U98;
wire P2_R1170_U99 , P2_R1170_U100 , P2_R1170_U101 , P2_R1170_U102 , P2_R1170_U103 , P2_R1170_U104 , P2_R1170_U105 , P2_R1170_U106 , P2_R1170_U107 , P2_R1170_U108;
wire P2_R1170_U109 , P2_R1170_U110 , P2_R1170_U111 , P2_R1170_U112 , P2_R1170_U113 , P2_R1170_U114 , P2_R1170_U115 , P2_R1170_U116 , P2_R1170_U117 , P2_R1170_U118;
wire P2_R1170_U119 , P2_R1170_U120 , P2_R1170_U121 , P2_R1170_U122 , P2_R1170_U123 , P2_R1170_U124 , P2_R1170_U125 , P2_R1170_U126 , P2_R1170_U127 , P2_R1170_U128;
wire P2_R1170_U129 , P2_R1170_U130 , P2_R1170_U131 , P2_R1170_U132 , P2_R1170_U133 , P2_R1170_U134 , P2_R1170_U135 , P2_R1170_U136 , P2_R1170_U137 , P2_R1170_U138;
wire P2_R1170_U139 , P2_R1170_U140 , P2_R1170_U141 , P2_R1170_U142 , P2_R1170_U143 , P2_R1170_U144 , P2_R1170_U145 , P2_R1170_U146 , P2_R1170_U147 , P2_R1170_U148;
wire P2_R1170_U149 , P2_R1170_U150 , P2_R1170_U151 , P2_R1170_U152 , P2_R1170_U153 , P2_R1170_U154 , P2_R1170_U155 , P2_R1170_U156 , P2_R1170_U157 , P2_R1170_U158;
wire P2_R1170_U159 , P2_R1170_U160 , P2_R1170_U161 , P2_R1170_U162 , P2_R1170_U163 , P2_R1170_U164 , P2_R1170_U165 , P2_R1170_U166 , P2_R1170_U167 , P2_R1170_U168;
wire P2_R1170_U169 , P2_R1170_U170 , P2_R1170_U171 , P2_R1170_U172 , P2_R1170_U173 , P2_R1170_U174 , P2_R1170_U175 , P2_R1170_U176 , P2_R1170_U177 , P2_R1170_U178;
wire P2_R1170_U179 , P2_R1170_U180 , P2_R1170_U181 , P2_R1170_U182 , P2_R1170_U183 , P2_R1170_U184 , P2_R1170_U185 , P2_R1170_U186 , P2_R1170_U187 , P2_R1170_U188;
wire P2_R1170_U189 , P2_R1170_U190 , P2_R1170_U191 , P2_R1170_U192 , P2_R1170_U193 , P2_R1170_U194 , P2_R1170_U195 , P2_R1170_U196 , P2_R1170_U197 , P2_R1170_U198;
wire P2_R1170_U199 , P2_R1170_U200 , P2_R1170_U201 , P2_R1170_U202 , P2_R1170_U203 , P2_R1170_U204 , P2_R1170_U205 , P2_R1170_U206 , P2_R1170_U207 , P2_R1170_U208;
wire P2_R1170_U209 , P2_R1170_U210 , P2_R1170_U211 , P2_R1170_U212 , P2_R1170_U213 , P2_R1170_U214 , P2_R1170_U215 , P2_R1170_U216 , P2_R1170_U217 , P2_R1170_U218;
wire P2_R1170_U219 , P2_R1170_U220 , P2_R1170_U221 , P2_R1170_U222 , P2_R1170_U223 , P2_R1170_U224 , P2_R1170_U225 , P2_R1170_U226 , P2_R1170_U227 , P2_R1170_U228;
wire P2_R1170_U229 , P2_R1170_U230 , P2_R1170_U231 , P2_R1170_U232 , P2_R1170_U233 , P2_R1170_U234 , P2_R1170_U235 , P2_R1170_U236 , P2_R1170_U237 , P2_R1170_U238;
wire P2_R1170_U239 , P2_R1170_U240 , P2_R1170_U241 , P2_R1170_U242 , P2_R1170_U243 , P2_R1170_U244 , P2_R1170_U245 , P2_R1170_U246 , P2_R1170_U247 , P2_R1170_U248;
wire P2_R1170_U249 , P2_R1170_U250 , P2_R1170_U251 , P2_R1170_U252 , P2_R1170_U253 , P2_R1170_U254 , P2_R1170_U255 , P2_R1170_U256 , P2_R1170_U257 , P2_R1170_U258;
wire P2_R1170_U259 , P2_R1170_U260 , P2_R1170_U261 , P2_R1170_U262 , P2_R1170_U263 , P2_R1170_U264 , P2_R1170_U265 , P2_R1170_U266 , P2_R1170_U267 , P2_R1170_U268;
wire P2_R1170_U269 , P2_R1170_U270 , P2_R1170_U271 , P2_R1170_U272 , P2_R1170_U273 , P2_R1170_U274 , P2_R1170_U275 , P2_R1170_U276 , P2_R1170_U277 , P2_R1170_U278;
wire P2_R1170_U279 , P2_R1170_U280 , P2_R1170_U281 , P2_R1170_U282 , P2_R1170_U283 , P2_R1170_U284 , P2_R1170_U285 , P2_R1170_U286 , P2_R1170_U287 , P2_R1170_U288;
wire P2_R1170_U289 , P2_R1170_U290 , P2_R1170_U291 , P2_R1170_U292 , P2_R1170_U293 , P2_R1170_U294 , P2_R1170_U295 , P2_R1170_U296 , P2_R1170_U297 , P2_R1170_U298;
wire P2_R1170_U299 , P2_R1170_U300 , P2_R1170_U301 , P2_R1170_U302 , P2_R1170_U303 , P2_R1170_U304 , P2_R1170_U305 , P2_R1170_U306 , P2_R1170_U307 , P2_R1170_U308;
wire P2_R1275_U6 , P2_R1275_U7 , P2_R1275_U8 , P2_R1275_U9 , P2_R1275_U10 , P2_R1275_U11 , P2_R1275_U12 , P2_R1275_U13 , P2_R1275_U14 , P2_R1275_U15;
wire P2_R1275_U16 , P2_R1275_U17 , P2_R1275_U18 , P2_R1275_U19 , P2_R1275_U20 , P2_R1275_U21 , P2_R1275_U22 , P2_R1275_U23 , P2_R1275_U24 , P2_R1275_U25;
wire P2_R1275_U26 , P2_R1275_U27 , P2_R1275_U28 , P2_R1275_U29 , P2_R1275_U30 , P2_R1275_U31 , P2_R1275_U32 , P2_R1275_U33 , P2_R1275_U34 , P2_R1275_U35;
wire P2_R1275_U36 , P2_R1275_U37 , P2_R1275_U38 , P2_R1275_U39 , P2_R1275_U40 , P2_R1275_U41 , P2_R1275_U42 , P2_R1275_U43 , P2_R1275_U44 , P2_R1275_U45;
wire P2_R1275_U46 , P2_R1275_U47 , P2_R1275_U48 , P2_R1275_U49 , P2_R1275_U50 , P2_R1275_U51 , P2_R1275_U52 , P2_R1275_U53 , P2_R1275_U54 , P2_R1275_U55;
wire P2_R1275_U56 , P2_R1275_U57 , P2_R1275_U58 , P2_R1275_U59 , P2_R1275_U60 , P2_R1275_U61 , P2_R1275_U62 , P2_R1275_U63 , P2_R1275_U64 , P2_R1275_U65;
wire P2_R1275_U66 , P2_R1275_U67 , P2_R1275_U68 , P2_R1275_U69 , P2_R1275_U70 , P2_R1275_U71 , P2_R1275_U72 , P2_R1275_U73 , P2_R1275_U74 , P2_R1275_U75;
wire P2_R1275_U76 , P2_R1275_U77 , P2_R1275_U78 , P2_R1275_U79 , P2_R1275_U80 , P2_R1275_U81 , P2_R1275_U82 , P2_R1275_U83 , P2_R1275_U84 , P2_R1275_U85;
wire P2_R1275_U86 , P2_R1275_U87 , P2_R1275_U88 , P2_R1275_U89 , P2_R1275_U90 , P2_R1275_U91 , P2_R1275_U92 , P2_R1275_U93 , P2_R1275_U94 , P2_R1275_U95;
wire P2_R1275_U96 , P2_R1275_U97 , P2_R1275_U98 , P2_R1275_U99 , P2_R1275_U100 , P2_R1275_U101 , P2_R1275_U102 , P2_R1275_U103 , P2_R1275_U104 , P2_R1275_U105;
wire P2_R1275_U106 , P2_R1275_U107 , P2_R1275_U108 , P2_R1275_U109 , P2_R1275_U110 , P2_R1275_U111 , P2_R1275_U112 , P2_R1275_U113 , P2_R1275_U114 , P2_R1275_U115;
wire P2_R1275_U116 , P2_R1275_U117 , P2_R1275_U118 , P2_R1275_U119 , P2_R1275_U120 , P2_R1275_U121 , P2_R1275_U122 , P2_R1275_U123 , P2_R1275_U124 , P2_R1275_U125;
wire P2_R1275_U126 , P2_R1275_U127 , P2_R1275_U128 , P2_R1275_U129 , P2_R1275_U130 , P2_R1275_U131 , P2_R1275_U132 , P2_R1275_U133 , P2_R1275_U134 , P2_R1275_U135;
wire P2_R1275_U136 , P2_R1275_U137 , P2_R1275_U138 , P2_R1275_U139 , P2_R1275_U140 , P2_R1275_U141 , P2_R1275_U142 , P2_R1275_U143 , P2_R1275_U144 , P2_R1275_U145;
wire P2_R1275_U146 , P2_R1275_U147 , P2_R1275_U148 , P2_R1275_U149 , P2_R1275_U150 , P2_R1275_U151 , P2_R1275_U152 , P2_R1275_U153 , P2_R1275_U154 , P2_R1275_U155;
wire P2_R1275_U156 , P2_R1275_U157 , P2_R1275_U158 , P2_R1275_U159 , P2_LT_719_U6 , P2_LT_719_U7 , P2_LT_719_U8 , P2_LT_719_U9 , P2_LT_719_U10 , P2_LT_719_U11;
wire P2_LT_719_U12 , P2_LT_719_U13 , P2_LT_719_U14 , P2_LT_719_U15 , P2_LT_719_U16 , P2_LT_719_U17 , P2_LT_719_U18 , P2_LT_719_U19 , P2_LT_719_U20 , P2_LT_719_U21;
wire P2_LT_719_U22 , P2_LT_719_U23 , P2_LT_719_U24 , P2_LT_719_U25 , P2_LT_719_U26 , P2_LT_719_U27 , P2_LT_719_U28 , P2_LT_719_U29 , P2_LT_719_U30 , P2_LT_719_U31;
wire P2_LT_719_U32 , P2_LT_719_U33 , P2_LT_719_U34 , P2_LT_719_U35 , P2_LT_719_U36 , P2_LT_719_U37 , P2_LT_719_U38 , P2_LT_719_U39 , P2_LT_719_U40 , P2_LT_719_U41;
wire P2_LT_719_U42 , P2_LT_719_U43 , P2_LT_719_U44 , P2_LT_719_U45 , P2_LT_719_U46 , P2_LT_719_U47 , P2_LT_719_U48 , P2_LT_719_U49 , P2_LT_719_U50 , P2_LT_719_U51;
wire P2_LT_719_U52 , P2_LT_719_U53 , P2_LT_719_U54 , P2_LT_719_U55 , P2_LT_719_U56 , P2_LT_719_U57 , P2_LT_719_U58 , P2_LT_719_U59 , P2_LT_719_U60 , P2_LT_719_U61;
wire P2_LT_719_U62 , P2_LT_719_U63 , P2_LT_719_U64 , P2_LT_719_U65 , P2_LT_719_U66 , P2_LT_719_U67 , P2_LT_719_U68 , P2_LT_719_U69 , P2_LT_719_U70 , P2_LT_719_U71;
wire P2_LT_719_U72 , P2_LT_719_U73 , P2_LT_719_U74 , P2_LT_719_U75 , P2_LT_719_U76 , P2_LT_719_U77 , P2_LT_719_U78 , P2_LT_719_U79 , P2_LT_719_U80 , P2_LT_719_U81;
wire P2_LT_719_U82 , P2_LT_719_U83 , P2_LT_719_U84 , P2_LT_719_U85 , P2_LT_719_U86 , P2_LT_719_U87 , P2_LT_719_U88 , P2_LT_719_U89 , P2_LT_719_U90 , P2_LT_719_U91;
wire P2_LT_719_U92 , P2_LT_719_U93 , P2_LT_719_U94 , P2_LT_719_U95 , P2_LT_719_U96 , P2_LT_719_U97 , P2_LT_719_U98 , P2_LT_719_U99 , P2_LT_719_U100 , P2_LT_719_U101;
wire P2_LT_719_U102 , P2_LT_719_U103 , P2_LT_719_U104 , P2_LT_719_U105 , P2_LT_719_U106 , P2_LT_719_U107 , P2_LT_719_U108 , P2_LT_719_U109 , P2_LT_719_U110 , P2_LT_719_U111;
wire P2_LT_719_U112 , P2_LT_719_U113 , P2_LT_719_U114 , P2_LT_719_U115 , P2_LT_719_U116 , P2_LT_719_U117 , P2_LT_719_U118 , P2_LT_719_U119 , P2_LT_719_U120 , P2_LT_719_U121;
wire P2_LT_719_U122 , P2_LT_719_U123 , P2_LT_719_U124 , P2_LT_719_U125 , P2_LT_719_U126 , P2_LT_719_U127 , P2_LT_719_U128 , P2_LT_719_U129 , P2_LT_719_U130 , P2_LT_719_U131;
wire P2_LT_719_U132 , P2_LT_719_U133 , P2_LT_719_U134 , P2_LT_719_U135 , P2_LT_719_U136 , P2_LT_719_U137 , P2_LT_719_U138 , P2_LT_719_U139 , P2_LT_719_U140 , P2_LT_719_U141;
wire P2_LT_719_U142 , P2_LT_719_U143 , P2_LT_719_U144 , P2_LT_719_U145 , P2_LT_719_U146 , P2_LT_719_U147 , P2_LT_719_U148 , P2_LT_719_U149 , P2_LT_719_U150 , P2_LT_719_U151;
wire P2_LT_719_U152 , P2_LT_719_U153 , P2_LT_719_U154 , P2_LT_719_U155 , P2_LT_719_U156 , P2_LT_719_U157 , P2_LT_719_U158 , P2_LT_719_U159 , P2_LT_719_U160 , P2_LT_719_U161;
wire P2_LT_719_U162 , P2_LT_719_U163 , P2_LT_719_U164 , P2_LT_719_U165 , P2_LT_719_U166 , P2_LT_719_U167 , P2_LT_719_U168 , P2_LT_719_U169 , P2_LT_719_U170 , P2_LT_719_U171;
wire P2_LT_719_U172 , P2_LT_719_U173 , P2_LT_719_U174 , P2_LT_719_U175 , P2_LT_719_U176 , P2_LT_719_U177 , P2_LT_719_U178 , P2_LT_719_U179 , P2_LT_719_U180 , P2_LT_719_U181;
wire P2_LT_719_U182 , P2_LT_719_U183 , P2_LT_719_U184 , P2_LT_719_U185 , P2_LT_719_U186 , P2_LT_719_U187 , P2_LT_719_U188 , P2_LT_719_U189 , P2_LT_719_U190 , P2_LT_719_U191;
wire P2_LT_719_U192 , P2_LT_719_U193 , P2_LT_719_U194 , P2_R1179_U6 , P2_R1179_U7 , P2_R1179_U8 , P2_R1179_U9 , P2_R1179_U10 , P2_R1179_U11 , P2_R1179_U12;
wire P2_R1179_U13 , P2_R1179_U14 , P2_R1179_U15 , P2_R1179_U16 , P2_R1179_U17 , P2_R1179_U18 , P2_R1179_U19 , P2_R1179_U20 , P2_R1179_U21 , P2_R1179_U22;
wire P2_R1179_U23 , P2_R1179_U24 , P2_R1179_U25 , P2_R1179_U26 , P2_R1179_U27 , P2_R1179_U28 , P2_R1179_U29 , P2_R1179_U30 , P2_R1179_U31 , P2_R1179_U32;
wire P2_R1179_U33 , P2_R1179_U34 , P2_R1179_U35 , P2_R1179_U36 , P2_R1179_U37 , P2_R1179_U38 , P2_R1179_U39 , P2_R1179_U40 , P2_R1179_U41 , P2_R1179_U42;
wire P2_R1179_U43 , P2_R1179_U44 , P2_R1179_U45 , P2_R1179_U46 , P2_R1179_U47 , P2_R1179_U48 , P2_R1179_U49 , P2_R1179_U50 , P2_R1179_U51 , P2_R1179_U52;
wire P2_R1179_U53 , P2_R1179_U54 , P2_R1179_U55 , P2_R1179_U56 , P2_R1179_U57 , P2_R1179_U58 , P2_R1179_U59 , P2_R1179_U60 , P2_R1179_U61 , P2_R1179_U62;
wire P2_R1179_U63 , P2_R1179_U64 , P2_R1179_U65 , P2_R1179_U66 , P2_R1179_U67 , P2_R1179_U68 , P2_R1179_U69 , P2_R1179_U70 , P2_R1179_U71 , P2_R1179_U72;
wire P2_R1179_U73 , P2_R1179_U74 , P2_R1179_U75 , P2_R1179_U76 , P2_R1179_U77 , P2_R1179_U78 , P2_R1179_U79 , P2_R1179_U80 , P2_R1179_U81 , P2_R1179_U82;
wire P2_R1179_U83 , P2_R1179_U84 , P2_R1179_U85 , P2_R1179_U86 , P2_R1179_U87 , P2_R1179_U88 , P2_R1179_U89 , P2_R1179_U90 , P2_R1179_U91 , P2_R1179_U92;
wire P2_R1179_U93 , P2_R1179_U94 , P2_R1179_U95 , P2_R1179_U96 , P2_R1179_U97 , P2_R1179_U98 , P2_R1179_U99 , P2_R1179_U100 , P2_R1179_U101 , P2_R1179_U102;
wire P2_R1179_U103 , P2_R1179_U104 , P2_R1179_U105 , P2_R1179_U106 , P2_R1179_U107 , P2_R1179_U108 , P2_R1179_U109 , P2_R1179_U110 , P2_R1179_U111 , P2_R1179_U112;
wire P2_R1179_U113 , P2_R1179_U114 , P2_R1179_U115 , P2_R1179_U116 , P2_R1179_U117 , P2_R1179_U118 , P2_R1179_U119 , P2_R1179_U120 , P2_R1179_U121 , P2_R1179_U122;
wire P2_R1179_U123 , P2_R1179_U124 , P2_R1179_U125 , P2_R1179_U126 , P2_R1179_U127 , P2_R1179_U128 , P2_R1179_U129 , P2_R1179_U130 , P2_R1179_U131 , P2_R1179_U132;
wire P2_R1179_U133 , P2_R1179_U134 , P2_R1179_U135 , P2_R1179_U136 , P2_R1179_U137 , P2_R1179_U138 , P2_R1179_U139 , P2_R1179_U140 , P2_R1179_U141 , P2_R1179_U142;
wire P2_R1179_U143 , P2_R1179_U144 , P2_R1179_U145 , P2_R1179_U146 , P2_R1179_U147 , P2_R1179_U148 , P2_R1179_U149 , P2_R1179_U150 , P2_R1179_U151 , P2_R1179_U152;
wire P2_R1179_U153 , P2_R1179_U154 , P2_R1179_U155 , P2_R1179_U156 , P2_R1179_U157 , P2_R1179_U158 , P2_R1179_U159 , P2_R1179_U160 , P2_R1179_U161 , P2_R1179_U162;
wire P2_R1179_U163 , P2_R1179_U164 , P2_R1179_U165 , P2_R1179_U166 , P2_R1179_U167 , P2_R1179_U168 , P2_R1179_U169 , P2_R1179_U170 , P2_R1179_U171 , P2_R1179_U172;
wire P2_R1179_U173 , P2_R1179_U174 , P2_R1179_U175 , P2_R1179_U176 , P2_R1179_U177 , P2_R1179_U178 , P2_R1179_U179 , P2_R1179_U180 , P2_R1179_U181 , P2_R1179_U182;
wire P2_R1179_U183 , P2_R1179_U184 , P2_R1179_U185 , P2_R1179_U186 , P2_R1179_U187 , P2_R1179_U188 , P2_R1179_U189 , P2_R1179_U190 , P2_R1179_U191 , P2_R1179_U192;
wire P2_R1179_U193 , P2_R1179_U194 , P2_R1179_U195 , P2_R1179_U196 , P2_R1179_U197 , P2_R1179_U198 , P2_R1179_U199 , P2_R1179_U200 , P2_R1179_U201 , P2_R1179_U202;
wire P2_R1179_U203 , P2_R1179_U204 , P2_R1179_U205 , P2_R1179_U206 , P2_R1179_U207 , P2_R1179_U208 , P2_R1179_U209 , P2_R1179_U210 , P2_R1179_U211 , P2_R1179_U212;
wire P2_R1179_U213 , P2_R1179_U214 , P2_R1179_U215 , P2_R1179_U216 , P2_R1179_U217 , P2_R1179_U218 , P2_R1179_U219 , P2_R1179_U220 , P2_R1179_U221 , P2_R1179_U222;
wire P2_R1179_U223 , P2_R1179_U224 , P2_R1179_U225 , P2_R1179_U226 , P2_R1179_U227 , P2_R1179_U228 , P2_R1179_U229 , P2_R1179_U230 , P2_R1179_U231 , P2_R1179_U232;
wire P2_R1179_U233 , P2_R1179_U234 , P2_R1179_U235 , P2_R1179_U236 , P2_R1179_U237 , P2_R1179_U238 , P2_R1179_U239 , P2_R1179_U240 , P2_R1179_U241 , P2_R1179_U242;
wire P2_R1179_U243 , P2_R1179_U244 , P2_R1179_U245 , P2_R1179_U246 , P2_R1179_U247 , P2_R1179_U248 , P2_R1179_U249 , P2_R1179_U250 , P2_R1179_U251 , P2_R1179_U252;
wire P2_R1179_U253 , P2_R1179_U254 , P2_R1179_U255 , P2_R1179_U256 , P2_R1179_U257 , P2_R1179_U258 , P2_R1179_U259 , P2_R1179_U260 , P2_R1179_U261 , P2_R1179_U262;
wire P2_R1179_U263 , P2_R1179_U264 , P2_R1179_U265 , P2_R1179_U266 , P2_R1179_U267 , P2_R1179_U268 , P2_R1179_U269 , P2_R1179_U270 , P2_R1179_U271 , P2_R1179_U272;
wire P2_R1179_U273 , P2_R1179_U274 , P2_R1179_U275 , P2_R1179_U276 , P2_R1179_U277 , P2_R1179_U278 , P2_R1179_U279 , P2_R1179_U280 , P2_R1179_U281 , P2_R1179_U282;
wire P2_R1179_U283 , P2_R1179_U284 , P2_R1179_U285 , P2_R1179_U286 , P2_R1179_U287 , P2_R1179_U288 , P2_R1179_U289 , P2_R1179_U290 , P2_R1179_U291 , P2_R1179_U292;
wire P2_R1179_U293 , P2_R1179_U294 , P2_R1179_U295 , P2_R1179_U296 , P2_R1179_U297 , P2_R1179_U298 , P2_R1179_U299 , P2_R1179_U300 , P2_R1179_U301 , P2_R1179_U302;
wire P2_R1179_U303 , P2_R1179_U304 , P2_R1179_U305 , P2_R1179_U306 , P2_R1179_U307 , P2_R1179_U308 , P2_R1179_U309 , P2_R1179_U310 , P2_R1179_U311 , P2_R1179_U312;
wire P2_R1179_U313 , P2_R1179_U314 , P2_R1179_U315 , P2_R1179_U316 , P2_R1179_U317 , P2_R1179_U318 , P2_R1179_U319 , P2_R1179_U320 , P2_R1179_U321 , P2_R1179_U322;
wire P2_R1179_U323 , P2_R1179_U324 , P2_R1179_U325 , P2_R1179_U326 , P2_R1179_U327 , P2_R1179_U328 , P2_R1179_U329 , P2_R1179_U330 , P2_R1179_U331 , P2_R1179_U332;
wire P2_R1179_U333 , P2_R1179_U334 , P2_R1179_U335 , P2_R1179_U336 , P2_R1179_U337 , P2_R1179_U338 , P2_R1179_U339 , P2_R1179_U340 , P2_R1179_U341 , P2_R1179_U342;
wire P2_R1179_U343 , P2_R1179_U344 , P2_R1179_U345 , P2_R1179_U346 , P2_R1179_U347 , P2_R1179_U348 , P2_R1179_U349 , P2_R1179_U350 , P2_R1179_U351 , P2_R1179_U352;
wire P2_R1179_U353 , P2_R1179_U354 , P2_R1179_U355 , P2_R1179_U356 , P2_R1179_U357 , P2_R1179_U358 , P2_R1179_U359 , P2_R1179_U360 , P2_R1179_U361 , P2_R1179_U362;
wire P2_R1179_U363 , P2_R1179_U364 , P2_R1179_U365 , P2_R1179_U366 , P2_R1179_U367 , P2_R1179_U368 , P2_R1179_U369 , P2_R1179_U370 , P2_R1179_U371 , P2_R1179_U372;
wire P2_R1179_U373 , P2_R1179_U374 , P2_R1179_U375 , P2_R1179_U376 , P2_R1179_U377 , P2_R1179_U378 , P2_R1179_U379 , P2_R1179_U380 , P2_R1179_U381 , P2_R1179_U382;
wire P2_R1179_U383 , P2_R1179_U384 , P2_R1179_U385 , P2_R1179_U386 , P2_R1179_U387 , P2_R1179_U388 , P2_R1179_U389 , P2_R1179_U390 , P2_R1179_U391 , P2_R1179_U392;
wire P2_R1179_U393 , P2_R1179_U394 , P2_R1179_U395 , P2_R1179_U396 , P2_R1179_U397 , P2_R1179_U398 , P2_R1179_U399 , P2_R1179_U400 , P2_R1179_U401 , P2_R1179_U402;
wire P2_R1179_U403 , P2_R1179_U404 , P2_R1179_U405 , P2_R1179_U406 , P2_R1179_U407 , P2_R1179_U408 , P2_R1179_U409 , P2_R1179_U410 , P2_R1179_U411 , P2_R1179_U412;
wire P2_R1179_U413 , P2_R1179_U414 , P2_R1179_U415 , P2_R1179_U416 , P2_R1179_U417 , P2_R1179_U418 , P2_R1179_U419 , P2_R1179_U420 , P2_R1179_U421 , P2_R1179_U422;
wire P2_R1179_U423 , P2_R1179_U424 , P2_R1179_U425 , P2_R1179_U426 , P2_R1179_U427 , P2_R1179_U428 , P2_R1179_U429 , P2_R1179_U430 , P2_R1179_U431 , P2_R1179_U432;
wire P2_R1179_U433 , P2_R1179_U434 , P2_R1179_U435 , P2_R1179_U436 , P2_R1179_U437 , P2_R1179_U438 , P2_R1179_U439 , P2_R1179_U440 , P2_R1179_U441 , P2_R1179_U442;
wire P2_R1179_U443 , P2_R1179_U444 , P2_R1179_U445 , P2_R1179_U446 , P2_R1179_U447 , P2_R1179_U448 , P2_R1179_U449 , P2_R1179_U450 , P2_R1179_U451 , P2_R1179_U452;
wire P2_R1179_U453 , P2_R1179_U454 , P2_R1179_U455 , P2_R1179_U456 , P2_R1179_U457 , P2_R1179_U458 , P2_R1179_U459 , P2_R1179_U460 , P2_R1179_U461 , P2_R1179_U462;
wire P2_R1179_U463 , P2_R1179_U464 , P2_R1179_U465 , P2_R1179_U466 , P2_R1179_U467 , P2_R1179_U468 , P2_R1179_U469 , P2_R1179_U470 , P2_R1179_U471 , P2_R1179_U472;
wire P2_R1179_U473 , P2_R1179_U474 , P2_R1179_U475 , P2_R1179_U476 , P2_R1179_U477 , P2_R1215_U4 , P2_R1215_U5 , P2_R1215_U6 , P2_R1215_U7 , P2_R1215_U8;
wire P2_R1215_U9 , P2_R1215_U10 , P2_R1215_U11 , P2_R1215_U12 , P2_R1215_U13 , P2_R1215_U14 , P2_R1215_U15 , P2_R1215_U16 , P2_R1215_U17 , P2_R1215_U18;
wire P2_R1215_U19 , P2_R1215_U20 , P2_R1215_U21 , P2_R1215_U22 , P2_R1215_U23 , P2_R1215_U24 , P2_R1215_U25 , P2_R1215_U26 , P2_R1215_U27 , P2_R1215_U28;
wire P2_R1215_U29 , P2_R1215_U30 , P2_R1215_U31 , P2_R1215_U32 , P2_R1215_U33 , P2_R1215_U34 , P2_R1215_U35 , P2_R1215_U36 , P2_R1215_U37 , P2_R1215_U38;
wire P2_R1215_U39 , P2_R1215_U40 , P2_R1215_U41 , P2_R1215_U42 , P2_R1215_U43 , P2_R1215_U44 , P2_R1215_U45 , P2_R1215_U46 , P2_R1215_U47 , P2_R1215_U48;
wire P2_R1215_U49 , P2_R1215_U50 , P2_R1215_U51 , P2_R1215_U52 , P2_R1215_U53 , P2_R1215_U54 , P2_R1215_U55 , P2_R1215_U56 , P2_R1215_U57 , P2_R1215_U58;
wire P2_R1215_U59 , P2_R1215_U60 , P2_R1215_U61 , P2_R1215_U62 , P2_R1215_U63 , P2_R1215_U64 , P2_R1215_U65 , P2_R1215_U66 , P2_R1215_U67 , P2_R1215_U68;
wire P2_R1215_U69 , P2_R1215_U70 , P2_R1215_U71 , P2_R1215_U72 , P2_R1215_U73 , P2_R1215_U74 , P2_R1215_U75 , P2_R1215_U76 , P2_R1215_U77 , P2_R1215_U78;
wire P2_R1215_U79 , P2_R1215_U80 , P2_R1215_U81 , P2_R1215_U82 , P2_R1215_U83 , P2_R1215_U84 , P2_R1215_U85 , P2_R1215_U86 , P2_R1215_U87 , P2_R1215_U88;
wire P2_R1215_U89 , P2_R1215_U90 , P2_R1215_U91 , P2_R1215_U92 , P2_R1215_U93 , P2_R1215_U94 , P2_R1215_U95 , P2_R1215_U96 , P2_R1215_U97 , P2_R1215_U98;
wire P2_R1215_U99 , P2_R1215_U100 , P2_R1215_U101 , P2_R1215_U102 , P2_R1215_U103 , P2_R1215_U104 , P2_R1215_U105 , P2_R1215_U106 , P2_R1215_U107 , P2_R1215_U108;
wire P2_R1215_U109 , P2_R1215_U110 , P2_R1215_U111 , P2_R1215_U112 , P2_R1215_U113 , P2_R1215_U114 , P2_R1215_U115 , P2_R1215_U116 , P2_R1215_U117 , P2_R1215_U118;
wire P2_R1215_U119 , P2_R1215_U120 , P2_R1215_U121 , P2_R1215_U122 , P2_R1215_U123 , P2_R1215_U124 , P2_R1215_U125 , P2_R1215_U126 , P2_R1215_U127 , P2_R1215_U128;
wire P2_R1215_U129 , P2_R1215_U130 , P2_R1215_U131 , P2_R1215_U132 , P2_R1215_U133 , P2_R1215_U134 , P2_R1215_U135 , P2_R1215_U136 , P2_R1215_U137 , P2_R1215_U138;
wire P2_R1215_U139 , P2_R1215_U140 , P2_R1215_U141 , P2_R1215_U142 , P2_R1215_U143 , P2_R1215_U144 , P2_R1215_U145 , P2_R1215_U146 , P2_R1215_U147 , P2_R1215_U148;
wire P2_R1215_U149 , P2_R1215_U150 , P2_R1215_U151 , P2_R1215_U152 , P2_R1215_U153 , P2_R1215_U154 , P2_R1215_U155 , P2_R1215_U156 , P2_R1215_U157 , P2_R1215_U158;
wire P2_R1215_U159 , P2_R1215_U160 , P2_R1215_U161 , P2_R1215_U162 , P2_R1215_U163 , P2_R1215_U164 , P2_R1215_U165 , P2_R1215_U166 , P2_R1215_U167 , P2_R1215_U168;
wire P2_R1215_U169 , P2_R1215_U170 , P2_R1215_U171 , P2_R1215_U172 , P2_R1215_U173 , P2_R1215_U174 , P2_R1215_U175 , P2_R1215_U176 , P2_R1215_U177 , P2_R1215_U178;
wire P2_R1215_U179 , P2_R1215_U180 , P2_R1215_U181 , P2_R1215_U182 , P2_R1215_U183 , P2_R1215_U184 , P2_R1215_U185 , P2_R1215_U186 , P2_R1215_U187 , P2_R1215_U188;
wire P2_R1215_U189 , P2_R1215_U190 , P2_R1215_U191 , P2_R1215_U192 , P2_R1215_U193 , P2_R1215_U194 , P2_R1215_U195 , P2_R1215_U196 , P2_R1215_U197 , P2_R1215_U198;
wire P2_R1215_U199 , P2_R1215_U200 , P2_R1215_U201 , P2_R1215_U202 , P2_R1215_U203 , P2_R1215_U204 , P2_R1215_U205 , P2_R1215_U206 , P2_R1215_U207 , P2_R1215_U208;
wire P2_R1215_U209 , P2_R1215_U210 , P2_R1215_U211 , P2_R1215_U212 , P2_R1215_U213 , P2_R1215_U214 , P2_R1215_U215 , P2_R1215_U216 , P2_R1215_U217 , P2_R1215_U218;
wire P2_R1215_U219 , P2_R1215_U220 , P2_R1215_U221 , P2_R1215_U222 , P2_R1215_U223 , P2_R1215_U224 , P2_R1215_U225 , P2_R1215_U226 , P2_R1215_U227 , P2_R1215_U228;
wire P2_R1215_U229 , P2_R1215_U230 , P2_R1215_U231 , P2_R1215_U232 , P2_R1215_U233 , P2_R1215_U234 , P2_R1215_U235 , P2_R1215_U236 , P2_R1215_U237 , P2_R1215_U238;
wire P2_R1215_U239 , P2_R1215_U240 , P2_R1215_U241 , P2_R1215_U242 , P2_R1215_U243 , P2_R1215_U244 , P2_R1215_U245 , P2_R1215_U246 , P2_R1215_U247 , P2_R1215_U248;
wire P2_R1215_U249 , P2_R1215_U250 , P2_R1215_U251 , P2_R1215_U252 , P2_R1215_U253 , P2_R1215_U254 , P2_R1215_U255 , P2_R1215_U256 , P2_R1215_U257 , P2_R1215_U258;
wire P2_R1215_U259 , P2_R1215_U260 , P2_R1215_U261 , P2_R1215_U262 , P2_R1215_U263 , P2_R1215_U264 , P2_R1215_U265 , P2_R1215_U266 , P2_R1215_U267 , P2_R1215_U268;
wire P2_R1215_U269 , P2_R1215_U270 , P2_R1215_U271 , P2_R1215_U272 , P2_R1215_U273 , P2_R1215_U274 , P2_R1215_U275 , P2_R1215_U276 , P2_R1215_U277 , P2_R1215_U278;
wire P2_R1215_U279 , P2_R1215_U280 , P2_R1215_U281 , P2_R1215_U282 , P2_R1215_U283 , P2_R1215_U284 , P2_R1215_U285 , P2_R1215_U286 , P2_R1215_U287 , P2_R1215_U288;
wire P2_R1215_U289 , P2_R1215_U290 , P2_R1215_U291 , P2_R1215_U292 , P2_R1215_U293 , P2_R1215_U294 , P2_R1215_U295 , P2_R1215_U296 , P2_R1215_U297 , P2_R1215_U298;
wire P2_R1215_U299 , P2_R1215_U300 , P2_R1215_U301 , P2_R1215_U302 , P2_R1215_U303 , P2_R1215_U304 , P2_R1215_U305 , P2_R1215_U306 , P2_R1215_U307 , P2_R1215_U308;
wire P2_R1215_U309 , P2_R1215_U310 , P2_R1215_U311 , P2_R1215_U312 , P2_R1215_U313 , P2_R1215_U314 , P2_R1215_U315 , P2_R1215_U316 , P2_R1215_U317 , P2_R1215_U318;
wire P2_R1215_U319 , P2_R1215_U320 , P2_R1215_U321 , P2_R1215_U322 , P2_R1215_U323 , P2_R1215_U324 , P2_R1215_U325 , P2_R1215_U326 , P2_R1215_U327 , P2_R1215_U328;
wire P2_R1215_U329 , P2_R1215_U330 , P2_R1215_U331 , P2_R1215_U332 , P2_R1215_U333 , P2_R1215_U334 , P2_R1215_U335 , P2_R1215_U336 , P2_R1215_U337 , P2_R1215_U338;
wire P2_R1215_U339 , P2_R1215_U340 , P2_R1215_U341 , P2_R1215_U342 , P2_R1215_U343 , P2_R1215_U344 , P2_R1215_U345 , P2_R1215_U346 , P2_R1215_U347 , P2_R1215_U348;
wire P2_R1215_U349 , P2_R1215_U350 , P2_R1215_U351 , P2_R1215_U352 , P2_R1215_U353 , P2_R1215_U354 , P2_R1215_U355 , P2_R1215_U356 , P2_R1215_U357 , P2_R1215_U358;
wire P2_R1215_U359 , P2_R1215_U360 , P2_R1215_U361 , P2_R1215_U362 , P2_R1215_U363 , P2_R1215_U364 , P2_R1215_U365 , P2_R1215_U366 , P2_R1215_U367 , P2_R1215_U368;
wire P2_R1215_U369 , P2_R1215_U370 , P2_R1215_U371 , P2_R1215_U372 , P2_R1215_U373 , P2_R1215_U374 , P2_R1215_U375 , P2_R1215_U376 , P2_R1215_U377 , P2_R1215_U378;
wire P2_R1215_U379 , P2_R1215_U380 , P2_R1215_U381 , P2_R1215_U382 , P2_R1215_U383 , P2_R1215_U384 , P2_R1215_U385 , P2_R1215_U386 , P2_R1215_U387 , P2_R1215_U388;
wire P2_R1215_U389 , P2_R1215_U390 , P2_R1215_U391 , P2_R1215_U392 , P2_R1215_U393 , P2_R1215_U394 , P2_R1215_U395 , P2_R1215_U396 , P2_R1215_U397 , P2_R1215_U398;
wire P2_R1215_U399 , P2_R1215_U400 , P2_R1215_U401 , P2_R1215_U402 , P2_R1215_U403 , P2_R1215_U404 , P2_R1215_U405 , P2_R1215_U406 , P2_R1215_U407 , P2_R1215_U408;
wire P2_R1215_U409 , P2_R1215_U410 , P2_R1215_U411 , P2_R1215_U412 , P2_R1215_U413 , P2_R1215_U414 , P2_R1215_U415 , P2_R1215_U416 , P2_R1215_U417 , P2_R1215_U418;
wire P2_R1215_U419 , P2_R1215_U420 , P2_R1215_U421 , P2_R1215_U422 , P2_R1215_U423 , P2_R1215_U424 , P2_R1215_U425 , P2_R1215_U426 , P2_R1215_U427 , P2_R1215_U428;
wire P2_R1215_U429 , P2_R1215_U430 , P2_R1215_U431 , P2_R1215_U432 , P2_R1215_U433 , P2_R1215_U434 , P2_R1215_U435 , P2_R1215_U436 , P2_R1215_U437 , P2_R1215_U438;
wire P2_R1215_U439 , P2_R1215_U440 , P2_R1215_U441 , P2_R1215_U442 , P2_R1215_U443 , P2_R1215_U444 , P2_R1215_U445 , P2_R1215_U446 , P2_R1215_U447 , P2_R1215_U448;
wire P2_R1215_U449 , P2_R1215_U450 , P2_R1215_U451 , P2_R1215_U452 , P2_R1215_U453 , P2_R1215_U454 , P2_R1215_U455 , P2_R1215_U456 , P2_R1215_U457 , P2_R1215_U458;
wire P2_R1215_U459 , P2_R1215_U460 , P2_R1215_U461 , P2_R1215_U462 , P2_R1215_U463 , P2_R1215_U464 , P2_R1215_U465 , P2_R1215_U466 , P2_R1215_U467 , P2_R1215_U468;
wire P2_R1215_U469 , P2_R1215_U470 , P2_R1215_U471 , P2_R1215_U472 , P2_R1215_U473 , P2_R1215_U474 , P2_R1215_U475 , P2_R1215_U476 , P2_R1215_U477 , P2_R1215_U478;
wire P2_R1215_U479 , P2_R1215_U480 , P2_R1215_U481 , P2_R1215_U482 , P2_R1215_U483 , P2_R1215_U484 , P2_R1215_U485 , P2_R1215_U486 , P2_R1215_U487 , P2_R1215_U488;
wire P2_R1215_U489 , P2_R1215_U490 , P2_R1215_U491 , P2_R1215_U492 , P2_R1215_U493 , P2_R1215_U494 , P2_R1215_U495 , P2_R1215_U496 , P2_R1215_U497 , P2_R1215_U498;
wire P2_R1215_U499 , P2_R1215_U500 , P2_R1215_U501 , P2_R1215_U502 , P2_R1215_U503 , P2_R1215_U504 , P2_R1164_U4 , P2_R1164_U5 , P2_R1164_U6 , P2_R1164_U7;
wire P2_R1164_U8 , P2_R1164_U9 , P2_R1164_U10 , P2_R1164_U11 , P2_R1164_U12 , P2_R1164_U13 , P2_R1164_U14 , P2_R1164_U15 , P2_R1164_U16 , P2_R1164_U17;
wire P2_R1164_U18 , P2_R1164_U19 , P2_R1164_U20 , P2_R1164_U21 , P2_R1164_U22 , P2_R1164_U23 , P2_R1164_U24 , P2_R1164_U25 , P2_R1164_U26 , P2_R1164_U27;
wire P2_R1164_U28 , P2_R1164_U29 , P2_R1164_U30 , P2_R1164_U31 , P2_R1164_U32 , P2_R1164_U33 , P2_R1164_U34 , P2_R1164_U35 , P2_R1164_U36 , P2_R1164_U37;
wire P2_R1164_U38 , P2_R1164_U39 , P2_R1164_U40 , P2_R1164_U41 , P2_R1164_U42 , P2_R1164_U43 , P2_R1164_U44 , P2_R1164_U45 , P2_R1164_U46 , P2_R1164_U47;
wire P2_R1164_U48 , P2_R1164_U49 , P2_R1164_U50 , P2_R1164_U51 , P2_R1164_U52 , P2_R1164_U53 , P2_R1164_U54 , P2_R1164_U55 , P2_R1164_U56 , P2_R1164_U57;
wire P2_R1164_U58 , P2_R1164_U59 , P2_R1164_U60 , P2_R1164_U61 , P2_R1164_U62 , P2_R1164_U63 , P2_R1164_U64 , P2_R1164_U65 , P2_R1164_U66 , P2_R1164_U67;
wire P2_R1164_U68 , P2_R1164_U69 , P2_R1164_U70 , P2_R1164_U71 , P2_R1164_U72 , P2_R1164_U73 , P2_R1164_U74 , P2_R1164_U75 , P2_R1164_U76 , P2_R1164_U77;
wire P2_R1164_U78 , P2_R1164_U79 , P2_R1164_U80 , P2_R1164_U81 , P2_R1164_U82 , P2_R1164_U83 , P2_R1164_U84 , P2_R1164_U85 , P2_R1164_U86 , P2_R1164_U87;
wire P2_R1164_U88 , P2_R1164_U89 , P2_R1164_U90 , P2_R1164_U91 , P2_R1164_U92 , P2_R1164_U93 , P2_R1164_U94 , P2_R1164_U95 , P2_R1164_U96 , P2_R1164_U97;
wire P2_R1164_U98 , P2_R1164_U99 , P2_R1164_U100 , P2_R1164_U101 , P2_R1164_U102 , P2_R1164_U103 , P2_R1164_U104 , P2_R1164_U105 , P2_R1164_U106 , P2_R1164_U107;
wire P2_R1164_U108 , P2_R1164_U109 , P2_R1164_U110 , P2_R1164_U111 , P2_R1164_U112 , P2_R1164_U113 , P2_R1164_U114 , P2_R1164_U115 , P2_R1164_U116 , P2_R1164_U117;
wire P2_R1164_U118 , P2_R1164_U119 , P2_R1164_U120 , P2_R1164_U121 , P2_R1164_U122 , P2_R1164_U123 , P2_R1164_U124 , P2_R1164_U125 , P2_R1164_U126 , P2_R1164_U127;
wire P2_R1164_U128 , P2_R1164_U129 , P2_R1164_U130 , P2_R1164_U131 , P2_R1164_U132 , P2_R1164_U133 , P2_R1164_U134 , P2_R1164_U135 , P2_R1164_U136 , P2_R1164_U137;
wire P2_R1164_U138 , P2_R1164_U139 , P2_R1164_U140 , P2_R1164_U141 , P2_R1164_U142 , P2_R1164_U143 , P2_R1164_U144 , P2_R1164_U145 , P2_R1164_U146 , P2_R1164_U147;
wire P2_R1164_U148 , P2_R1164_U149 , P2_R1164_U150 , P2_R1164_U151 , P2_R1164_U152 , P2_R1164_U153 , P2_R1164_U154 , P2_R1164_U155 , P2_R1164_U156 , P2_R1164_U157;
wire P2_R1164_U158 , P2_R1164_U159 , P2_R1164_U160 , P2_R1164_U161 , P2_R1164_U162 , P2_R1164_U163 , P2_R1164_U164 , P2_R1164_U165 , P2_R1164_U166 , P2_R1164_U167;
wire P2_R1164_U168 , P2_R1164_U169 , P2_R1164_U170 , P2_R1164_U171 , P2_R1164_U172 , P2_R1164_U173 , P2_R1164_U174 , P2_R1164_U175 , P2_R1164_U176 , P2_R1164_U177;
wire P2_R1164_U178 , P2_R1164_U179 , P2_R1164_U180 , P2_R1164_U181 , P2_R1164_U182 , P2_R1164_U183 , P2_R1164_U184 , P2_R1164_U185 , P2_R1164_U186 , P2_R1164_U187;
wire P2_R1164_U188 , P2_R1164_U189 , P2_R1164_U190 , P2_R1164_U191 , P2_R1164_U192 , P2_R1164_U193 , P2_R1164_U194 , P2_R1164_U195 , P2_R1164_U196 , P2_R1164_U197;
wire P2_R1164_U198 , P2_R1164_U199 , P2_R1164_U200 , P2_R1164_U201 , P2_R1164_U202 , P2_R1164_U203 , P2_R1164_U204 , P2_R1164_U205 , P2_R1164_U206 , P2_R1164_U207;
wire P2_R1164_U208 , P2_R1164_U209 , P2_R1164_U210 , P2_R1164_U211 , P2_R1164_U212 , P2_R1164_U213 , P2_R1164_U214 , P2_R1164_U215 , P2_R1164_U216 , P2_R1164_U217;
wire P2_R1164_U218 , P2_R1164_U219 , P2_R1164_U220 , P2_R1164_U221 , P2_R1164_U222 , P2_R1164_U223 , P2_R1164_U224 , P2_R1164_U225 , P2_R1164_U226 , P2_R1164_U227;
wire P2_R1164_U228 , P2_R1164_U229 , P2_R1164_U230 , P2_R1164_U231 , P2_R1164_U232 , P2_R1164_U233 , P2_R1164_U234 , P2_R1164_U235 , P2_R1164_U236 , P2_R1164_U237;
wire P2_R1164_U238 , P2_R1164_U239 , P2_R1164_U240 , P2_R1164_U241 , P2_R1164_U242 , P2_R1164_U243 , P2_R1164_U244 , P2_R1164_U245 , P2_R1164_U246 , P2_R1164_U247;
wire P2_R1164_U248 , P2_R1164_U249 , P2_R1164_U250 , P2_R1164_U251 , P2_R1164_U252 , P2_R1164_U253 , P2_R1164_U254 , P2_R1164_U255 , P2_R1164_U256 , P2_R1164_U257;
wire P2_R1164_U258 , P2_R1164_U259 , P2_R1164_U260 , P2_R1164_U261 , P2_R1164_U262 , P2_R1164_U263 , P2_R1164_U264 , P2_R1164_U265 , P2_R1164_U266 , P2_R1164_U267;
wire P2_R1164_U268 , P2_R1164_U269 , P2_R1164_U270 , P2_R1164_U271 , P2_R1164_U272 , P2_R1164_U273 , P2_R1164_U274 , P2_R1164_U275 , P2_R1164_U276 , P2_R1164_U277;
wire P2_R1164_U278 , P2_R1164_U279 , P2_R1164_U280 , P2_R1164_U281 , P2_R1164_U282 , P2_R1164_U283 , P2_R1164_U284 , P2_R1164_U285 , P2_R1164_U286 , P2_R1164_U287;
wire P2_R1164_U288 , P2_R1164_U289 , P2_R1164_U290 , P2_R1164_U291 , P2_R1164_U292 , P2_R1164_U293 , P2_R1164_U294 , P2_R1164_U295 , P2_R1164_U296 , P2_R1164_U297;
wire P2_R1164_U298 , P2_R1164_U299 , P2_R1164_U300 , P2_R1164_U301 , P2_R1164_U302 , P2_R1164_U303 , P2_R1164_U304 , P2_R1164_U305 , P2_R1164_U306 , P2_R1164_U307;
wire P2_R1164_U308 , P2_R1164_U309 , P2_R1164_U310 , P2_R1164_U311 , P2_R1164_U312 , P2_R1164_U313 , P2_R1164_U314 , P2_R1164_U315 , P2_R1164_U316 , P2_R1164_U317;
wire P2_R1164_U318 , P2_R1164_U319 , P2_R1164_U320 , P2_R1164_U321 , P2_R1164_U322 , P2_R1164_U323 , P2_R1164_U324 , P2_R1164_U325 , P2_R1164_U326 , P2_R1164_U327;
wire P2_R1164_U328 , P2_R1164_U329 , P2_R1164_U330 , P2_R1164_U331 , P2_R1164_U332 , P2_R1164_U333 , P2_R1164_U334 , P2_R1164_U335 , P2_R1164_U336 , P2_R1164_U337;
wire P2_R1164_U338 , P2_R1164_U339 , P2_R1164_U340 , P2_R1164_U341 , P2_R1164_U342 , P2_R1164_U343 , P2_R1164_U344 , P2_R1164_U345 , P2_R1164_U346 , P2_R1164_U347;
wire P2_R1164_U348 , P2_R1164_U349 , P2_R1164_U350 , P2_R1164_U351 , P2_R1164_U352 , P2_R1164_U353 , P2_R1164_U354 , P2_R1164_U355 , P2_R1164_U356 , P2_R1164_U357;
wire P2_R1164_U358 , P2_R1164_U359 , P2_R1164_U360 , P2_R1164_U361 , P2_R1164_U362 , P2_R1164_U363 , P2_R1164_U364 , P2_R1164_U365 , P2_R1164_U366 , P2_R1164_U367;
wire P2_R1164_U368 , P2_R1164_U369 , P2_R1164_U370 , P2_R1164_U371 , P2_R1164_U372 , P2_R1164_U373 , P2_R1164_U374 , P2_R1164_U375 , P2_R1164_U376 , P2_R1164_U377;
wire P2_R1164_U378 , P2_R1164_U379 , P2_R1164_U380 , P2_R1164_U381 , P2_R1164_U382 , P2_R1164_U383 , P2_R1164_U384 , P2_R1164_U385 , P2_R1164_U386 , P2_R1164_U387;
wire P2_R1164_U388 , P2_R1164_U389 , P2_R1164_U390 , P2_R1164_U391 , P2_R1164_U392 , P2_R1164_U393 , P2_R1164_U394 , P2_R1164_U395 , P2_R1164_U396 , P2_R1164_U397;
wire P2_R1164_U398 , P2_R1164_U399 , P2_R1164_U400 , P2_R1164_U401 , P2_R1164_U402 , P2_R1164_U403 , P2_R1164_U404 , P2_R1164_U405 , P2_R1164_U406 , P2_R1164_U407;
wire P2_R1164_U408 , P2_R1164_U409 , P2_R1164_U410 , P2_R1164_U411 , P2_R1164_U412 , P2_R1164_U413 , P2_R1164_U414 , P2_R1164_U415 , P2_R1164_U416 , P2_R1164_U417;
wire P2_R1164_U418 , P2_R1164_U419 , P2_R1164_U420 , P2_R1164_U421 , P2_R1164_U422 , P2_R1164_U423 , P2_R1164_U424 , P2_R1164_U425 , P2_R1164_U426 , P2_R1164_U427;
wire P2_R1164_U428 , P2_R1164_U429 , P2_R1164_U430 , P2_R1164_U431 , P2_R1164_U432 , P2_R1164_U433 , P2_R1164_U434 , P2_R1164_U435 , P2_R1164_U436 , P2_R1164_U437;
wire P2_R1164_U438 , P2_R1164_U439 , P2_R1164_U440 , P2_R1164_U441 , P2_R1164_U442 , P2_R1164_U443 , P2_R1164_U444 , P2_R1164_U445 , P2_R1164_U446 , P2_R1164_U447;
wire P2_R1164_U448 , P2_R1164_U449 , P2_R1164_U450 , P2_R1164_U451 , P2_R1164_U452 , P2_R1164_U453 , P2_R1164_U454 , P2_R1164_U455 , P2_R1164_U456 , P2_R1164_U457;
wire P2_R1164_U458 , P2_R1164_U459 , P2_R1164_U460 , P2_R1164_U461 , P2_R1164_U462 , P2_R1164_U463 , P2_R1164_U464 , P2_R1164_U465 , P2_R1164_U466 , P2_R1164_U467;
wire P2_R1164_U468 , P2_R1164_U469 , P2_R1164_U470 , P2_R1164_U471 , P2_R1164_U472 , P2_R1164_U473 , P2_R1164_U474 , P2_R1164_U475 , P2_R1164_U476 , P2_R1164_U477;
wire P2_R1164_U478 , P2_R1164_U479 , P2_R1164_U480 , P2_R1164_U481 , P2_R1164_U482 , P2_R1164_U483 , P2_R1164_U484 , P2_R1164_U485 , P2_R1164_U486 , P2_R1164_U487;
wire P2_R1164_U488 , P2_R1164_U489 , P2_R1164_U490 , P2_R1164_U491 , P2_R1164_U492 , P2_R1164_U493 , P2_R1164_U494 , P2_R1164_U495 , P2_R1164_U496 , P2_R1164_U497;
wire P2_R1164_U498 , P2_R1164_U499 , P2_R1164_U500 , P2_R1164_U501 , P2_R1164_U502 , P2_R1164_U503 , P2_R1164_U504 , P2_R1233_U4 , P2_R1233_U5 , P2_R1233_U6;
wire P2_R1233_U7 , P2_R1233_U8 , P2_R1233_U9 , P2_R1233_U10 , P2_R1233_U11 , P2_R1233_U12 , P2_R1233_U13 , P2_R1233_U14 , P2_R1233_U15 , P2_R1233_U16;
wire P2_R1233_U17 , P2_R1233_U18 , P2_R1233_U19 , P2_R1233_U20 , P2_R1233_U21 , P2_R1233_U22 , P2_R1233_U23 , P2_R1233_U24 , P2_R1233_U25 , P2_R1233_U26;
wire P2_R1233_U27 , P2_R1233_U28 , P2_R1233_U29 , P2_R1233_U30 , P2_R1233_U31 , P2_R1233_U32 , P2_R1233_U33 , P2_R1233_U34 , P2_R1233_U35 , P2_R1233_U36;
wire P2_R1233_U37 , P2_R1233_U38 , P2_R1233_U39 , P2_R1233_U40 , P2_R1233_U41 , P2_R1233_U42 , P2_R1233_U43 , P2_R1233_U44 , P2_R1233_U45 , P2_R1233_U46;
wire P2_R1233_U47 , P2_R1233_U48 , P2_R1233_U49 , P2_R1233_U50 , P2_R1233_U51 , P2_R1233_U52 , P2_R1233_U53 , P2_R1233_U54 , P2_R1233_U55 , P2_R1233_U56;
wire P2_R1233_U57 , P2_R1233_U58 , P2_R1233_U59 , P2_R1233_U60 , P2_R1233_U61 , P2_R1233_U62 , P2_R1233_U63 , P2_R1233_U64 , P2_R1233_U65 , P2_R1233_U66;
wire P2_R1233_U67 , P2_R1233_U68 , P2_R1233_U69 , P2_R1233_U70 , P2_R1233_U71 , P2_R1233_U72 , P2_R1233_U73 , P2_R1233_U74 , P2_R1233_U75 , P2_R1233_U76;
wire P2_R1233_U77 , P2_R1233_U78 , P2_R1233_U79 , P2_R1233_U80 , P2_R1233_U81 , P2_R1233_U82 , P2_R1233_U83 , P2_R1233_U84 , P2_R1233_U85 , P2_R1233_U86;
wire P2_R1233_U87 , P2_R1233_U88 , P2_R1233_U89 , P2_R1233_U90 , P2_R1233_U91 , P2_R1233_U92 , P2_R1233_U93 , P2_R1233_U94 , P2_R1233_U95 , P2_R1233_U96;
wire P2_R1233_U97 , P2_R1233_U98 , P2_R1233_U99 , P2_R1233_U100 , P2_R1233_U101 , P2_R1233_U102 , P2_R1233_U103 , P2_R1233_U104 , P2_R1233_U105 , P2_R1233_U106;
wire P2_R1233_U107 , P2_R1233_U108 , P2_R1233_U109 , P2_R1233_U110 , P2_R1233_U111 , P2_R1233_U112 , P2_R1233_U113 , P2_R1233_U114 , P2_R1233_U115 , P2_R1233_U116;
wire P2_R1233_U117 , P2_R1233_U118 , P2_R1233_U119 , P2_R1233_U120 , P2_R1233_U121 , P2_R1233_U122 , P2_R1233_U123 , P2_R1233_U124 , P2_R1233_U125 , P2_R1233_U126;
wire P2_R1233_U127 , P2_R1233_U128 , P2_R1233_U129 , P2_R1233_U130 , P2_R1233_U131 , P2_R1233_U132 , P2_R1233_U133 , P2_R1233_U134 , P2_R1233_U135 , P2_R1233_U136;
wire P2_R1233_U137 , P2_R1233_U138 , P2_R1233_U139 , P2_R1233_U140 , P2_R1233_U141 , P2_R1233_U142 , P2_R1233_U143 , P2_R1233_U144 , P2_R1233_U145 , P2_R1233_U146;
wire P2_R1233_U147 , P2_R1233_U148 , P2_R1233_U149 , P2_R1233_U150 , P2_R1233_U151 , P2_R1233_U152 , P2_R1233_U153 , P2_R1233_U154 , P2_R1233_U155 , P2_R1233_U156;
wire P2_R1233_U157 , P2_R1233_U158 , P2_R1233_U159 , P2_R1233_U160 , P2_R1233_U161 , P2_R1233_U162 , P2_R1233_U163 , P2_R1233_U164 , P2_R1233_U165 , P2_R1233_U166;
wire P2_R1233_U167 , P2_R1233_U168 , P2_R1233_U169 , P2_R1233_U170 , P2_R1233_U171 , P2_R1233_U172 , P2_R1233_U173 , P2_R1233_U174 , P2_R1233_U175 , P2_R1233_U176;
wire P2_R1233_U177 , P2_R1233_U178 , P2_R1233_U179 , P2_R1233_U180 , P2_R1233_U181 , P2_R1233_U182 , P2_R1233_U183 , P2_R1233_U184 , P2_R1233_U185 , P2_R1233_U186;
wire P2_R1233_U187 , P2_R1233_U188 , P2_R1233_U189 , P2_R1233_U190 , P2_R1233_U191 , P2_R1233_U192 , P2_R1233_U193 , P2_R1233_U194 , P2_R1233_U195 , P2_R1233_U196;
wire P2_R1233_U197 , P2_R1233_U198 , P2_R1233_U199 , P2_R1233_U200 , P2_R1233_U201 , P2_R1233_U202 , P2_R1233_U203 , P2_R1233_U204 , P2_R1233_U205 , P2_R1233_U206;
wire P2_R1233_U207 , P2_R1233_U208 , P2_R1233_U209 , P2_R1233_U210 , P2_R1233_U211 , P2_R1233_U212 , P2_R1233_U213 , P2_R1233_U214 , P2_R1233_U215 , P2_R1233_U216;
wire P2_R1233_U217 , P2_R1233_U218 , P2_R1233_U219 , P2_R1233_U220 , P2_R1233_U221 , P2_R1233_U222 , P2_R1233_U223 , P2_R1233_U224 , P2_R1233_U225 , P2_R1233_U226;
wire P2_R1233_U227 , P2_R1233_U228 , P2_R1233_U229 , P2_R1233_U230 , P2_R1233_U231 , P2_R1233_U232 , P2_R1233_U233 , P2_R1233_U234 , P2_R1233_U235 , P2_R1233_U236;
wire P2_R1233_U237 , P2_R1233_U238 , P2_R1233_U239 , P2_R1233_U240 , P2_R1233_U241 , P2_R1233_U242 , P2_R1233_U243 , P2_R1233_U244 , P2_R1233_U245 , P2_R1233_U246;
wire P2_R1233_U247 , P2_R1233_U248 , P2_R1233_U249 , P2_R1233_U250 , P2_R1233_U251 , P2_R1233_U252 , P2_R1233_U253 , P2_R1233_U254 , P2_R1233_U255 , P2_R1233_U256;
wire P2_R1233_U257 , P2_R1233_U258 , P2_R1233_U259 , P2_R1233_U260 , P2_R1233_U261 , P2_R1233_U262 , P2_R1233_U263 , P2_R1233_U264 , P2_R1233_U265 , P2_R1233_U266;
wire P2_R1233_U267 , P2_R1233_U268 , P2_R1233_U269 , P2_R1233_U270 , P2_R1233_U271 , P2_R1233_U272 , P2_R1233_U273 , P2_R1233_U274 , P2_R1233_U275 , P2_R1233_U276;
wire P2_R1233_U277 , P2_R1233_U278 , P2_R1233_U279 , P2_R1233_U280 , P2_R1233_U281 , P2_R1233_U282 , P2_R1233_U283 , P2_R1233_U284 , P2_R1233_U285 , P2_R1233_U286;
wire P2_R1233_U287 , P2_R1233_U288 , P2_R1233_U289 , P2_R1233_U290 , P2_R1233_U291 , P2_R1233_U292 , P2_R1233_U293 , P2_R1233_U294 , P2_R1233_U295 , P2_R1233_U296;
wire P2_R1233_U297 , P2_R1233_U298 , P2_R1233_U299 , P2_R1233_U300 , P2_R1233_U301 , P2_R1233_U302 , P2_R1233_U303 , P2_R1233_U304 , P2_R1233_U305 , P2_R1233_U306;
wire P2_R1233_U307 , P2_R1233_U308 , P2_R1233_U309 , P2_R1233_U310 , P2_R1233_U311 , P2_R1233_U312 , P2_R1233_U313 , P2_R1233_U314 , P2_R1233_U315 , P2_R1233_U316;
wire P2_R1233_U317 , P2_R1233_U318 , P2_R1233_U319 , P2_R1233_U320 , P2_R1233_U321 , P2_R1233_U322 , P2_R1233_U323 , P2_R1233_U324 , P2_R1233_U325 , P2_R1233_U326;
wire P2_R1233_U327 , P2_R1233_U328 , P2_R1233_U329 , P2_R1233_U330 , P2_R1233_U331 , P2_R1233_U332 , P2_R1233_U333 , P2_R1233_U334 , P2_R1233_U335 , P2_R1233_U336;
wire P2_R1233_U337 , P2_R1233_U338 , P2_R1233_U339 , P2_R1233_U340 , P2_R1233_U341 , P2_R1233_U342 , P2_R1233_U343 , P2_R1233_U344 , P2_R1233_U345 , P2_R1233_U346;
wire P2_R1233_U347 , P2_R1233_U348 , P2_R1233_U349 , P2_R1233_U350 , P2_R1233_U351 , P2_R1233_U352 , P2_R1233_U353 , P2_R1233_U354 , P2_R1233_U355 , P2_R1233_U356;
wire P2_R1233_U357 , P2_R1233_U358 , P2_R1233_U359 , P2_R1233_U360 , P2_R1233_U361 , P2_R1233_U362 , P2_R1233_U363 , P2_R1233_U364 , P2_R1233_U365 , P2_R1233_U366;
wire P2_R1233_U367 , P2_R1233_U368 , P2_R1233_U369 , P2_R1233_U370 , P2_R1233_U371 , P2_R1233_U372 , P2_R1233_U373 , P2_R1233_U374 , P2_R1233_U375 , P2_R1233_U376;
wire P2_R1233_U377 , P2_R1233_U378 , P2_R1233_U379 , P2_R1233_U380 , P2_R1233_U381 , P2_R1233_U382 , P2_R1233_U383 , P2_R1233_U384 , P2_R1233_U385 , P2_R1233_U386;
wire P2_R1233_U387 , P2_R1233_U388 , P2_R1233_U389 , P2_R1233_U390 , P2_R1233_U391 , P2_R1233_U392 , P2_R1233_U393 , P2_R1233_U394 , P2_R1233_U395 , P2_R1233_U396;
wire P2_R1233_U397 , P2_R1233_U398 , P2_R1233_U399 , P2_R1233_U400 , P2_R1233_U401 , P2_R1233_U402 , P2_R1233_U403 , P2_R1233_U404 , P2_R1233_U405 , P2_R1233_U406;
wire P2_R1233_U407 , P2_R1233_U408 , P2_R1233_U409 , P2_R1233_U410 , P2_R1233_U411 , P2_R1233_U412 , P2_R1233_U413 , P2_R1233_U414 , P2_R1233_U415 , P2_R1233_U416;
wire P2_R1233_U417 , P2_R1233_U418 , P2_R1233_U419 , P2_R1233_U420 , P2_R1233_U421 , P2_R1233_U422 , P2_R1233_U423 , P2_R1233_U424 , P2_R1233_U425 , P2_R1233_U426;
wire P2_R1233_U427 , P2_R1233_U428 , P2_R1233_U429 , P2_R1233_U430 , P2_R1233_U431 , P2_R1233_U432 , P2_R1233_U433 , P2_R1233_U434 , P2_R1233_U435 , P2_R1233_U436;
wire P2_R1233_U437 , P2_R1233_U438 , P2_R1233_U439 , P2_R1233_U440 , P2_R1233_U441 , P2_R1233_U442 , P2_R1233_U443 , P2_R1233_U444 , P2_R1233_U445 , P2_R1233_U446;
wire P2_R1233_U447 , P2_R1233_U448 , P2_R1233_U449 , P2_R1233_U450 , P2_R1233_U451 , P2_R1233_U452 , P2_R1233_U453 , P2_R1233_U454 , P2_R1233_U455 , P2_R1233_U456;
wire P2_R1233_U457 , P2_R1233_U458 , P2_R1233_U459 , P2_R1233_U460 , P2_R1233_U461 , P2_R1233_U462 , P2_R1233_U463 , P2_R1233_U464 , P2_R1233_U465 , P2_R1233_U466;
wire P2_R1233_U467 , P2_R1233_U468 , P2_R1233_U469 , P2_R1233_U470 , P2_R1233_U471 , P2_R1233_U472 , P2_R1233_U473 , P2_R1233_U474 , P2_R1233_U475 , P2_R1233_U476;
wire P2_R1233_U477 , P2_R1233_U478 , P2_R1233_U479 , P2_R1233_U480 , P2_R1233_U481 , P2_R1233_U482 , P2_R1233_U483 , P2_R1233_U484 , P2_R1233_U485 , P2_R1233_U486;
wire P2_R1233_U487 , P2_R1233_U488 , P2_R1233_U489 , P2_R1233_U490 , P2_R1233_U491 , P2_R1233_U492 , P2_R1233_U493 , P2_R1233_U494 , P2_R1233_U495 , P2_R1233_U496;
wire P2_R1233_U497 , P2_R1233_U498 , P2_R1233_U499 , P2_R1233_U500 , P2_R1233_U501 , P2_R1233_U502 , P2_R1233_U503 , P2_R1233_U504 , P2_R1176_U4 , P2_R1176_U5;
wire P2_R1176_U6 , P2_R1176_U7 , P2_R1176_U8 , P2_R1176_U9 , P2_R1176_U10 , P2_R1176_U11 , P2_R1176_U12 , P2_R1176_U13 , P2_R1176_U14 , P2_R1176_U15;
wire P2_R1176_U16 , P2_R1176_U17 , P2_R1176_U18 , P2_R1176_U19 , P2_R1176_U20 , P2_R1176_U21 , P2_R1176_U22 , P2_R1176_U23 , P2_R1176_U24 , P2_R1176_U25;
wire P2_R1176_U26 , P2_R1176_U27 , P2_R1176_U28 , P2_R1176_U29 , P2_R1176_U30 , P2_R1176_U31 , P2_R1176_U32 , P2_R1176_U33 , P2_R1176_U34 , P2_R1176_U35;
wire P2_R1176_U36 , P2_R1176_U37 , P2_R1176_U38 , P2_R1176_U39 , P2_R1176_U40 , P2_R1176_U41 , P2_R1176_U42 , P2_R1176_U43 , P2_R1176_U44 , P2_R1176_U45;
wire P2_R1176_U46 , P2_R1176_U47 , P2_R1176_U48 , P2_R1176_U49 , P2_R1176_U50 , P2_R1176_U51 , P2_R1176_U52 , P2_R1176_U53 , P2_R1176_U54 , P2_R1176_U55;
wire P2_R1176_U56 , P2_R1176_U57 , P2_R1176_U58 , P2_R1176_U59 , P2_R1176_U60 , P2_R1176_U61 , P2_R1176_U62 , P2_R1176_U63 , P2_R1176_U64 , P2_R1176_U65;
wire P2_R1176_U66 , P2_R1176_U67 , P2_R1176_U68 , P2_R1176_U69 , P2_R1176_U70 , P2_R1176_U71 , P2_R1176_U72 , P2_R1176_U73 , P2_R1176_U74 , P2_R1176_U75;
wire P2_R1176_U76 , P2_R1176_U77 , P2_R1176_U78 , P2_R1176_U79 , P2_R1176_U80 , P2_R1176_U81 , P2_R1176_U82 , P2_R1176_U83 , P2_R1176_U84 , P2_R1176_U85;
wire P2_R1176_U86 , P2_R1176_U87 , P2_R1176_U88 , P2_R1176_U89 , P2_R1176_U90 , P2_R1176_U91 , P2_R1176_U92 , P2_R1176_U93 , P2_R1176_U94 , P2_R1176_U95;
wire P2_R1176_U96 , P2_R1176_U97 , P2_R1176_U98 , P2_R1176_U99 , P2_R1176_U100 , P2_R1176_U101 , P2_R1176_U102 , P2_R1176_U103 , P2_R1176_U104 , P2_R1176_U105;
wire P2_R1176_U106 , P2_R1176_U107 , P2_R1176_U108 , P2_R1176_U109 , P2_R1176_U110 , P2_R1176_U111 , P2_R1176_U112 , P2_R1176_U113 , P2_R1176_U114 , P2_R1176_U115;
wire P2_R1176_U116 , P2_R1176_U117 , P2_R1176_U118 , P2_R1176_U119 , P2_R1176_U120 , P2_R1176_U121 , P2_R1176_U122 , P2_R1176_U123 , P2_R1176_U124 , P2_R1176_U125;
wire P2_R1176_U126 , P2_R1176_U127 , P2_R1176_U128 , P2_R1176_U129 , P2_R1176_U130 , P2_R1176_U131 , P2_R1176_U132 , P2_R1176_U133 , P2_R1176_U134 , P2_R1176_U135;
wire P2_R1176_U136 , P2_R1176_U137 , P2_R1176_U138 , P2_R1176_U139 , P2_R1176_U140 , P2_R1176_U141 , P2_R1176_U142 , P2_R1176_U143 , P2_R1176_U144 , P2_R1176_U145;
wire P2_R1176_U146 , P2_R1176_U147 , P2_R1176_U148 , P2_R1176_U149 , P2_R1176_U150 , P2_R1176_U151 , P2_R1176_U152 , P2_R1176_U153 , P2_R1176_U154 , P2_R1176_U155;
wire P2_R1176_U156 , P2_R1176_U157 , P2_R1176_U158 , P2_R1176_U159 , P2_R1176_U160 , P2_R1176_U161 , P2_R1176_U162 , P2_R1176_U163 , P2_R1176_U164 , P2_R1176_U165;
wire P2_R1176_U166 , P2_R1176_U167 , P2_R1176_U168 , P2_R1176_U169 , P2_R1176_U170 , P2_R1176_U171 , P2_R1176_U172 , P2_R1176_U173 , P2_R1176_U174 , P2_R1176_U175;
wire P2_R1176_U176 , P2_R1176_U177 , P2_R1176_U178 , P2_R1176_U179 , P2_R1176_U180 , P2_R1176_U181 , P2_R1176_U182 , P2_R1176_U183 , P2_R1176_U184 , P2_R1176_U185;
wire P2_R1176_U186 , P2_R1176_U187 , P2_R1176_U188 , P2_R1176_U189 , P2_R1176_U190 , P2_R1176_U191 , P2_R1176_U192 , P2_R1176_U193 , P2_R1176_U194 , P2_R1176_U195;
wire P2_R1176_U196 , P2_R1176_U197 , P2_R1176_U198 , P2_R1176_U199 , P2_R1176_U200 , P2_R1176_U201 , P2_R1176_U202 , P2_R1176_U203 , P2_R1176_U204 , P2_R1176_U205;
wire P2_R1176_U206 , P2_R1176_U207 , P2_R1176_U208 , P2_R1176_U209 , P2_R1176_U210 , P2_R1176_U211 , P2_R1176_U212 , P2_R1176_U213 , P2_R1176_U214 , P2_R1176_U215;
wire P2_R1176_U216 , P2_R1176_U217 , P2_R1176_U218 , P2_R1176_U219 , P2_R1176_U220 , P2_R1176_U221 , P2_R1176_U222 , P2_R1176_U223 , P2_R1176_U224 , P2_R1176_U225;
wire P2_R1176_U226 , P2_R1176_U227 , P2_R1176_U228 , P2_R1176_U229 , P2_R1176_U230 , P2_R1176_U231 , P2_R1176_U232 , P2_R1176_U233 , P2_R1176_U234 , P2_R1176_U235;
wire P2_R1176_U236 , P2_R1176_U237 , P2_R1176_U238 , P2_R1176_U239 , P2_R1176_U240 , P2_R1176_U241 , P2_R1176_U242 , P2_R1176_U243 , P2_R1176_U244 , P2_R1176_U245;
wire P2_R1176_U246 , P2_R1176_U247 , P2_R1176_U248 , P2_R1176_U249 , P2_R1176_U250 , P2_R1176_U251 , P2_R1176_U252 , P2_R1176_U253 , P2_R1176_U254 , P2_R1176_U255;
wire P2_R1176_U256 , P2_R1176_U257 , P2_R1176_U258 , P2_R1176_U259 , P2_R1176_U260 , P2_R1176_U261 , P2_R1176_U262 , P2_R1176_U263 , P2_R1176_U264 , P2_R1176_U265;
wire P2_R1176_U266 , P2_R1176_U267 , P2_R1176_U268 , P2_R1176_U269 , P2_R1176_U270 , P2_R1176_U271 , P2_R1176_U272 , P2_R1176_U273 , P2_R1176_U274 , P2_R1176_U275;
wire P2_R1176_U276 , P2_R1176_U277 , P2_R1176_U278 , P2_R1176_U279 , P2_R1176_U280 , P2_R1176_U281 , P2_R1176_U282 , P2_R1176_U283 , P2_R1176_U284 , P2_R1176_U285;
wire P2_R1176_U286 , P2_R1176_U287 , P2_R1176_U288 , P2_R1176_U289 , P2_R1176_U290 , P2_R1176_U291 , P2_R1176_U292 , P2_R1176_U293 , P2_R1176_U294 , P2_R1176_U295;
wire P2_R1176_U296 , P2_R1176_U297 , P2_R1176_U298 , P2_R1176_U299 , P2_R1176_U300 , P2_R1176_U301 , P2_R1176_U302 , P2_R1176_U303 , P2_R1176_U304 , P2_R1176_U305;
wire P2_R1176_U306 , P2_R1176_U307 , P2_R1176_U308 , P2_R1176_U309 , P2_R1176_U310 , P2_R1176_U311 , P2_R1176_U312 , P2_R1176_U313 , P2_R1176_U314 , P2_R1176_U315;
wire P2_R1176_U316 , P2_R1176_U317 , P2_R1176_U318 , P2_R1176_U319 , P2_R1176_U320 , P2_R1176_U321 , P2_R1176_U322 , P2_R1176_U323 , P2_R1176_U324 , P2_R1176_U325;
wire P2_R1176_U326 , P2_R1176_U327 , P2_R1176_U328 , P2_R1176_U329 , P2_R1176_U330 , P2_R1176_U331 , P2_R1176_U332 , P2_R1176_U333 , P2_R1176_U334 , P2_R1176_U335;
wire P2_R1176_U336 , P2_R1176_U337 , P2_R1176_U338 , P2_R1176_U339 , P2_R1176_U340 , P2_R1176_U341 , P2_R1176_U342 , P2_R1176_U343 , P2_R1176_U344 , P2_R1176_U345;
wire P2_R1176_U346 , P2_R1176_U347 , P2_R1176_U348 , P2_R1176_U349 , P2_R1176_U350 , P2_R1176_U351 , P2_R1176_U352 , P2_R1176_U353 , P2_R1176_U354 , P2_R1176_U355;
wire P2_R1176_U356 , P2_R1176_U357 , P2_R1176_U358 , P2_R1176_U359 , P2_R1176_U360 , P2_R1176_U361 , P2_R1176_U362 , P2_R1176_U363 , P2_R1176_U364 , P2_R1176_U365;
wire P2_R1176_U366 , P2_R1176_U367 , P2_R1176_U368 , P2_R1176_U369 , P2_R1176_U370 , P2_R1176_U371 , P2_R1176_U372 , P2_R1176_U373 , P2_R1176_U374 , P2_R1176_U375;
wire P2_R1176_U376 , P2_R1176_U377 , P2_R1176_U378 , P2_R1176_U379 , P2_R1176_U380 , P2_R1176_U381 , P2_R1176_U382 , P2_R1176_U383 , P2_R1176_U384 , P2_R1176_U385;
wire P2_R1176_U386 , P2_R1176_U387 , P2_R1176_U388 , P2_R1176_U389 , P2_R1176_U390 , P2_R1176_U391 , P2_R1176_U392 , P2_R1176_U393 , P2_R1176_U394 , P2_R1176_U395;
wire P2_R1176_U396 , P2_R1176_U397 , P2_R1176_U398 , P2_R1176_U399 , P2_R1176_U400 , P2_R1176_U401 , P2_R1176_U402 , P2_R1176_U403 , P2_R1176_U404 , P2_R1176_U405;
wire P2_R1176_U406 , P2_R1176_U407 , P2_R1176_U408 , P2_R1176_U409 , P2_R1176_U410 , P2_R1176_U411 , P2_R1176_U412 , P2_R1176_U413 , P2_R1176_U414 , P2_R1176_U415;
wire P2_R1176_U416 , P2_R1176_U417 , P2_R1176_U418 , P2_R1176_U419 , P2_R1176_U420 , P2_R1176_U421 , P2_R1176_U422 , P2_R1176_U423 , P2_R1176_U424 , P2_R1176_U425;
wire P2_R1176_U426 , P2_R1176_U427 , P2_R1176_U428 , P2_R1176_U429 , P2_R1176_U430 , P2_R1176_U431 , P2_R1176_U432 , P2_R1176_U433 , P2_R1176_U434 , P2_R1176_U435;
wire P2_R1176_U436 , P2_R1176_U437 , P2_R1176_U438 , P2_R1176_U439 , P2_R1176_U440 , P2_R1176_U441 , P2_R1176_U442 , P2_R1176_U443 , P2_R1176_U444 , P2_R1176_U445;
wire P2_R1176_U446 , P2_R1176_U447 , P2_R1176_U448 , P2_R1176_U449 , P2_R1176_U450 , P2_R1176_U451 , P2_R1176_U452 , P2_R1176_U453 , P2_R1176_U454 , P2_R1176_U455;
wire P2_R1176_U456 , P2_R1176_U457 , P2_R1176_U458 , P2_R1176_U459 , P2_R1176_U460 , P2_R1176_U461 , P2_R1176_U462 , P2_R1176_U463 , P2_R1176_U464 , P2_R1176_U465;
wire P2_R1176_U466 , P2_R1176_U467 , P2_R1176_U468 , P2_R1176_U469 , P2_R1176_U470 , P2_R1176_U471 , P2_R1176_U472 , P2_R1176_U473 , P2_R1176_U474 , P2_R1176_U475;
wire P2_R1176_U476 , P2_R1176_U477 , P2_R1176_U478 , P2_R1176_U479 , P2_R1176_U480 , P2_R1176_U481 , P2_R1176_U482 , P2_R1176_U483 , P2_R1176_U484 , P2_R1176_U485;
wire P2_R1176_U486 , P2_R1176_U487 , P2_R1176_U488 , P2_R1176_U489 , P2_R1176_U490 , P2_R1176_U491 , P2_R1176_U492 , P2_R1176_U493 , P2_R1176_U494 , P2_R1176_U495;
wire P2_R1176_U496 , P2_R1176_U497 , P2_R1176_U498 , P2_R1176_U499 , P2_R1176_U500 , P2_R1176_U501 , P2_R1176_U502 , P2_R1176_U503 , P2_R1176_U504 , P2_R1176_U505;
wire P2_R1176_U506 , P2_R1176_U507 , P2_R1176_U508 , P2_R1176_U509 , P2_R1176_U510 , P2_R1176_U511 , P2_R1176_U512 , P2_R1176_U513 , P2_R1176_U514 , P2_R1176_U515;
wire P2_R1176_U516 , P2_R1176_U517 , P2_R1176_U518 , P2_R1176_U519 , P2_R1176_U520 , P2_R1176_U521 , P2_R1176_U522 , P2_R1176_U523 , P2_R1176_U524 , P2_R1176_U525;
wire P2_R1176_U526 , P2_R1176_U527 , P2_R1176_U528 , P2_R1176_U529 , P2_R1176_U530 , P2_R1176_U531 , P2_R1176_U532 , P2_R1176_U533 , P2_R1176_U534 , P2_R1176_U535;
wire P2_R1176_U536 , P2_R1176_U537 , P2_R1176_U538 , P2_R1176_U539 , P2_R1176_U540 , P2_R1176_U541 , P2_R1176_U542 , P2_R1176_U543 , P2_R1176_U544 , P2_R1176_U545;
wire P2_R1176_U546 , P2_R1176_U547 , P2_R1176_U548 , P2_R1176_U549 , P2_R1176_U550 , P2_R1176_U551 , P2_R1176_U552 , P2_R1176_U553 , P2_R1176_U554 , P2_R1176_U555;
wire P2_R1176_U556 , P2_R1176_U557 , P2_R1176_U558 , P2_R1176_U559 , P2_R1176_U560 , P2_R1176_U561 , P2_R1176_U562 , P2_R1176_U563 , P2_R1176_U564 , P2_R1176_U565;
wire P2_R1176_U566 , P2_R1176_U567 , P2_R1176_U568 , P2_R1176_U569 , P2_R1176_U570 , P2_R1176_U571 , P2_R1176_U572 , P2_R1176_U573 , P2_R1176_U574 , P2_R1176_U575;
wire P2_R1176_U576 , P2_R1176_U577 , P2_R1176_U578 , P2_R1176_U579 , P2_R1176_U580 , P2_R1176_U581 , P2_R1176_U582 , P2_R1176_U583 , P2_R1176_U584 , P2_R1176_U585;
wire P2_R1176_U586 , P2_R1176_U587 , P2_R1176_U588 , P2_R1176_U589 , P2_R1176_U590 , P2_R1176_U591 , P2_R1176_U592 , P2_R1176_U593 , P2_R1176_U594 , P2_R1176_U595;
wire P2_R1176_U596 , P2_R1176_U597 , P2_R1176_U598 , P2_R1176_U599 , P2_R1176_U600 , P2_R1176_U601 , P2_R1176_U602 , P2_R1131_U4 , P2_R1131_U5 , P2_R1131_U6;
wire P2_R1131_U7 , P2_R1131_U8 , P2_R1131_U9 , P2_R1131_U10 , P2_R1131_U11 , P2_R1131_U12 , P2_R1131_U13 , P2_R1131_U14 , P2_R1131_U15 , P2_R1131_U16;
wire P2_R1131_U17 , P2_R1131_U18 , P2_R1131_U19 , P2_R1131_U20 , P2_R1131_U21 , P2_R1131_U22 , P2_R1131_U23 , P2_R1131_U24 , P2_R1131_U25 , P2_R1131_U26;
wire P2_R1131_U27 , P2_R1131_U28 , P2_R1131_U29 , P2_R1131_U30 , P2_R1131_U31 , P2_R1131_U32 , P2_R1131_U33 , P2_R1131_U34 , P2_R1131_U35 , P2_R1131_U36;
wire P2_R1131_U37 , P2_R1131_U38 , P2_R1131_U39 , P2_R1131_U40 , P2_R1131_U41 , P2_R1131_U42 , P2_R1131_U43 , P2_R1131_U44 , P2_R1131_U45 , P2_R1131_U46;
wire P2_R1131_U47 , P2_R1131_U48 , P2_R1131_U49 , P2_R1131_U50 , P2_R1131_U51 , P2_R1131_U52 , P2_R1131_U53 , P2_R1131_U54 , P2_R1131_U55 , P2_R1131_U56;
wire P2_R1131_U57 , P2_R1131_U58 , P2_R1131_U59 , P2_R1131_U60 , P2_R1131_U61 , P2_R1131_U62 , P2_R1131_U63 , P2_R1131_U64 , P2_R1131_U65 , P2_R1131_U66;
wire P2_R1131_U67 , P2_R1131_U68 , P2_R1131_U69 , P2_R1131_U70 , P2_R1131_U71 , P2_R1131_U72 , P2_R1131_U73 , P2_R1131_U74 , P2_R1131_U75 , P2_R1131_U76;
wire P2_R1131_U77 , P2_R1131_U78 , P2_R1131_U79 , P2_R1131_U80 , P2_R1131_U81 , P2_R1131_U82 , P2_R1131_U83 , P2_R1131_U84 , P2_R1131_U85 , P2_R1131_U86;
wire P2_R1131_U87 , P2_R1131_U88 , P2_R1131_U89 , P2_R1131_U90 , P2_R1131_U91 , P2_R1131_U92 , P2_R1131_U93 , P2_R1131_U94 , P2_R1131_U95 , P2_R1131_U96;
wire P2_R1131_U97 , P2_R1131_U98 , P2_R1131_U99 , P2_R1131_U100 , P2_R1131_U101 , P2_R1131_U102 , P2_R1131_U103 , P2_R1131_U104 , P2_R1131_U105 , P2_R1131_U106;
wire P2_R1131_U107 , P2_R1131_U108 , P2_R1131_U109 , P2_R1131_U110 , P2_R1131_U111 , P2_R1131_U112 , P2_R1131_U113 , P2_R1131_U114 , P2_R1131_U115 , P2_R1131_U116;
wire P2_R1131_U117 , P2_R1131_U118 , P2_R1131_U119 , P2_R1131_U120 , P2_R1131_U121 , P2_R1131_U122 , P2_R1131_U123 , P2_R1131_U124 , P2_R1131_U125 , P2_R1131_U126;
wire P2_R1131_U127 , P2_R1131_U128 , P2_R1131_U129 , P2_R1131_U130 , P2_R1131_U131 , P2_R1131_U132 , P2_R1131_U133 , P2_R1131_U134 , P2_R1131_U135 , P2_R1131_U136;
wire P2_R1131_U137 , P2_R1131_U138 , P2_R1131_U139 , P2_R1131_U140 , P2_R1131_U141 , P2_R1131_U142 , P2_R1131_U143 , P2_R1131_U144 , P2_R1131_U145 , P2_R1131_U146;
wire P2_R1131_U147 , P2_R1131_U148 , P2_R1131_U149 , P2_R1131_U150 , P2_R1131_U151 , P2_R1131_U152 , P2_R1131_U153 , P2_R1131_U154 , P2_R1131_U155 , P2_R1131_U156;
wire P2_R1131_U157 , P2_R1131_U158 , P2_R1131_U159 , P2_R1131_U160 , P2_R1131_U161 , P2_R1131_U162 , P2_R1131_U163 , P2_R1131_U164 , P2_R1131_U165 , P2_R1131_U166;
wire P2_R1131_U167 , P2_R1131_U168 , P2_R1131_U169 , P2_R1131_U170 , P2_R1131_U171 , P2_R1131_U172 , P2_R1131_U173 , P2_R1131_U174 , P2_R1131_U175 , P2_R1131_U176;
wire P2_R1131_U177 , P2_R1131_U178 , P2_R1131_U179 , P2_R1131_U180 , P2_R1131_U181 , P2_R1131_U182 , P2_R1131_U183 , P2_R1131_U184 , P2_R1131_U185 , P2_R1131_U186;
wire P2_R1131_U187 , P2_R1131_U188 , P2_R1131_U189 , P2_R1131_U190 , P2_R1131_U191 , P2_R1131_U192 , P2_R1131_U193 , P2_R1131_U194 , P2_R1131_U195 , P2_R1131_U196;
wire P2_R1131_U197 , P2_R1131_U198 , P2_R1131_U199 , P2_R1131_U200 , P2_R1131_U201 , P2_R1131_U202 , P2_R1131_U203 , P2_R1131_U204 , P2_R1131_U205 , P2_R1131_U206;
wire P2_R1131_U207 , P2_R1131_U208 , P2_R1131_U209 , P2_R1131_U210 , P2_R1131_U211 , P2_R1131_U212 , P2_R1131_U213 , P2_R1131_U214 , P2_R1131_U215 , P2_R1131_U216;
wire P2_R1131_U217 , P2_R1131_U218 , P2_R1131_U219 , P2_R1131_U220 , P2_R1131_U221 , P2_R1131_U222 , P2_R1131_U223 , P2_R1131_U224 , P2_R1131_U225 , P2_R1131_U226;
wire P2_R1131_U227 , P2_R1131_U228 , P2_R1131_U229 , P2_R1131_U230 , P2_R1131_U231 , P2_R1131_U232 , P2_R1131_U233 , P2_R1131_U234 , P2_R1131_U235 , P2_R1131_U236;
wire P2_R1131_U237 , P2_R1131_U238 , P2_R1131_U239 , P2_R1131_U240 , P2_R1131_U241 , P2_R1131_U242 , P2_R1131_U243 , P2_R1131_U244 , P2_R1131_U245 , P2_R1131_U246;
wire P2_R1131_U247 , P2_R1131_U248 , P2_R1131_U249 , P2_R1131_U250 , P2_R1131_U251 , P2_R1131_U252 , P2_R1131_U253 , P2_R1131_U254 , P2_R1131_U255 , P2_R1131_U256;
wire P2_R1131_U257 , P2_R1131_U258 , P2_R1131_U259 , P2_R1131_U260 , P2_R1131_U261 , P2_R1131_U262 , P2_R1131_U263 , P2_R1131_U264 , P2_R1131_U265 , P2_R1131_U266;
wire P2_R1131_U267 , P2_R1131_U268 , P2_R1131_U269 , P2_R1131_U270 , P2_R1131_U271 , P2_R1131_U272 , P2_R1131_U273 , P2_R1131_U274 , P2_R1131_U275 , P2_R1131_U276;
wire P2_R1131_U277 , P2_R1131_U278 , P2_R1131_U279 , P2_R1131_U280 , P2_R1131_U281 , P2_R1131_U282 , P2_R1131_U283 , P2_R1131_U284 , P2_R1131_U285 , P2_R1131_U286;
wire P2_R1131_U287 , P2_R1131_U288 , P2_R1131_U289 , P2_R1131_U290 , P2_R1131_U291 , P2_R1131_U292 , P2_R1131_U293 , P2_R1131_U294 , P2_R1131_U295 , P2_R1131_U296;
wire P2_R1131_U297 , P2_R1131_U298 , P2_R1131_U299 , P2_R1131_U300 , P2_R1131_U301 , P2_R1131_U302 , P2_R1131_U303 , P2_R1131_U304 , P2_R1131_U305 , P2_R1131_U306;
wire P2_R1131_U307 , P2_R1131_U308 , P2_R1131_U309 , P2_R1131_U310 , P2_R1131_U311 , P2_R1131_U312 , P2_R1131_U313 , P2_R1131_U314 , P2_R1131_U315 , P2_R1131_U316;
wire P2_R1131_U317 , P2_R1131_U318 , P2_R1131_U319 , P2_R1131_U320 , P2_R1131_U321 , P2_R1131_U322 , P2_R1131_U323 , P2_R1131_U324 , P2_R1131_U325 , P2_R1131_U326;
wire P2_R1131_U327 , P2_R1131_U328 , P2_R1131_U329 , P2_R1131_U330 , P2_R1131_U331 , P2_R1131_U332 , P2_R1131_U333 , P2_R1131_U334 , P2_R1131_U335 , P2_R1131_U336;
wire P2_R1131_U337 , P2_R1131_U338 , P2_R1131_U339 , P2_R1131_U340 , P2_R1131_U341 , P2_R1131_U342 , P2_R1131_U343 , P2_R1131_U344 , P2_R1131_U345 , P2_R1131_U346;
wire P2_R1131_U347 , P2_R1131_U348 , P2_R1131_U349 , P2_R1131_U350 , P2_R1131_U351 , P2_R1131_U352 , P2_R1131_U353 , P2_R1131_U354 , P2_R1131_U355 , P2_R1131_U356;
wire P2_R1131_U357 , P2_R1131_U358 , P2_R1131_U359 , P2_R1131_U360 , P2_R1131_U361 , P2_R1131_U362 , P2_R1131_U363 , P2_R1131_U364 , P2_R1131_U365 , P2_R1131_U366;
wire P2_R1131_U367 , P2_R1131_U368 , P2_R1131_U369 , P2_R1131_U370 , P2_R1131_U371 , P2_R1131_U372 , P2_R1131_U373 , P2_R1131_U374 , P2_R1131_U375 , P2_R1131_U376;
wire P2_R1131_U377 , P2_R1131_U378 , P2_R1131_U379 , P2_R1131_U380 , P2_R1131_U381 , P2_R1131_U382 , P2_R1131_U383 , P2_R1131_U384 , P2_R1131_U385 , P2_R1131_U386;
wire P2_R1131_U387 , P2_R1131_U388 , P2_R1131_U389 , P2_R1131_U390 , P2_R1131_U391 , P2_R1131_U392 , P2_R1131_U393 , P2_R1131_U394 , P2_R1131_U395 , P2_R1131_U396;
wire P2_R1131_U397 , P2_R1131_U398 , P2_R1131_U399 , P2_R1131_U400 , P2_R1131_U401 , P2_R1131_U402 , P2_R1131_U403 , P2_R1131_U404 , P2_R1131_U405 , P2_R1131_U406;
wire P2_R1131_U407 , P2_R1131_U408 , P2_R1131_U409 , P2_R1131_U410 , P2_R1131_U411 , P2_R1131_U412 , P2_R1131_U413 , P2_R1131_U414 , P2_R1131_U415 , P2_R1131_U416;
wire P2_R1131_U417 , P2_R1131_U418 , P2_R1131_U419 , P2_R1131_U420 , P2_R1131_U421 , P2_R1131_U422 , P2_R1131_U423 , P2_R1131_U424 , P2_R1131_U425 , P2_R1131_U426;
wire P2_R1131_U427 , P2_R1131_U428 , P2_R1131_U429 , P2_R1131_U430 , P2_R1131_U431 , P2_R1131_U432 , P2_R1131_U433 , P2_R1131_U434 , P2_R1131_U435 , P2_R1131_U436;
wire P2_R1131_U437 , P2_R1131_U438 , P2_R1131_U439 , P2_R1131_U440 , P2_R1131_U441 , P2_R1131_U442 , P2_R1131_U443 , P2_R1131_U444 , P2_R1131_U445 , P2_R1131_U446;
wire P2_R1131_U447 , P2_R1131_U448 , P2_R1131_U449 , P2_R1131_U450 , P2_R1131_U451 , P2_R1131_U452 , P2_R1131_U453 , P2_R1131_U454 , P2_R1131_U455 , P2_R1131_U456;
wire P2_R1131_U457 , P2_R1131_U458 , P2_R1131_U459 , P2_R1131_U460 , P2_R1131_U461 , P2_R1131_U462 , P2_R1131_U463 , P2_R1131_U464 , P2_R1131_U465 , P2_R1131_U466;
wire P2_R1131_U467 , P2_R1131_U468 , P2_R1131_U469 , P2_R1131_U470 , P2_R1131_U471 , P2_R1131_U472 , P2_R1131_U473 , P2_R1131_U474 , P2_R1131_U475 , P2_R1131_U476;
wire P2_R1131_U477 , P2_R1131_U478 , P2_R1131_U479 , P2_R1131_U480 , P2_R1131_U481 , P2_R1131_U482 , P2_R1131_U483 , P2_R1131_U484 , P2_R1131_U485 , P2_R1131_U486;
wire P2_R1131_U487 , P2_R1131_U488 , P2_R1131_U489 , P2_R1131_U490 , P2_R1131_U491 , P2_R1131_U492 , P2_R1131_U493 , P2_R1131_U494 , P2_R1131_U495 , P2_R1131_U496;
wire P2_R1131_U497 , P2_R1131_U498 , P2_R1131_U499 , P2_R1131_U500 , P2_R1131_U501 , P2_R1131_U502 , P2_R1131_U503 , P2_R1131_U504 , P2_R1146_U6 , P2_R1146_U7;
wire P2_R1146_U8 , P2_R1146_U9 , P2_R1146_U10 , P2_R1146_U11 , P2_R1146_U12 , P2_R1146_U13 , P2_R1146_U14 , P2_R1146_U15 , P2_R1146_U16 , P2_R1146_U17;
wire P2_R1146_U18 , P2_R1146_U19 , P2_R1146_U20 , P2_R1146_U21 , P2_R1146_U22 , P2_R1146_U23 , P2_R1146_U24 , P2_R1146_U25 , P2_R1146_U26 , P2_R1146_U27;
wire P2_R1146_U28 , P2_R1146_U29 , P2_R1146_U30 , P2_R1146_U31 , P2_R1146_U32 , P2_R1146_U33 , P2_R1146_U34 , P2_R1146_U35 , P2_R1146_U36 , P2_R1146_U37;
wire P2_R1146_U38 , P2_R1146_U39 , P2_R1146_U40 , P2_R1146_U41 , P2_R1146_U42 , P2_R1146_U43 , P2_R1146_U44 , P2_R1146_U45 , P2_R1146_U46 , P2_R1146_U47;
wire P2_R1146_U48 , P2_R1146_U49 , P2_R1146_U50 , P2_R1146_U51 , P2_R1146_U52 , P2_R1146_U53 , P2_R1146_U54 , P2_R1146_U55 , P2_R1146_U56 , P2_R1146_U57;
wire P2_R1146_U58 , P2_R1146_U59 , P2_R1146_U60 , P2_R1146_U61 , P2_R1146_U62 , P2_R1146_U63 , P2_R1146_U64 , P2_R1146_U65 , P2_R1146_U66 , P2_R1146_U67;
wire P2_R1146_U68 , P2_R1146_U69 , P2_R1146_U70 , P2_R1146_U71 , P2_R1146_U72 , P2_R1146_U73 , P2_R1146_U74 , P2_R1146_U75 , P2_R1146_U76 , P2_R1146_U77;
wire P2_R1146_U78 , P2_R1146_U79 , P2_R1146_U80 , P2_R1146_U81 , P2_R1146_U82 , P2_R1146_U83 , P2_R1146_U84 , P2_R1146_U85 , P2_R1146_U86 , P2_R1146_U87;
wire P2_R1146_U88 , P2_R1146_U89 , P2_R1146_U90 , P2_R1146_U91 , P2_R1146_U92 , P2_R1146_U93 , P2_R1146_U94 , P2_R1146_U95 , P2_R1146_U96 , P2_R1146_U97;
wire P2_R1146_U98 , P2_R1146_U99 , P2_R1146_U100 , P2_R1146_U101 , P2_R1146_U102 , P2_R1146_U103 , P2_R1146_U104 , P2_R1146_U105 , P2_R1146_U106 , P2_R1146_U107;
wire P2_R1146_U108 , P2_R1146_U109 , P2_R1146_U110 , P2_R1146_U111 , P2_R1146_U112 , P2_R1146_U113 , P2_R1146_U114 , P2_R1146_U115 , P2_R1146_U116 , P2_R1146_U117;
wire P2_R1146_U118 , P2_R1146_U119 , P2_R1146_U120 , P2_R1146_U121 , P2_R1146_U122 , P2_R1146_U123 , P2_R1146_U124 , P2_R1146_U125 , P2_R1146_U126 , P2_R1146_U127;
wire P2_R1146_U128 , P2_R1146_U129 , P2_R1146_U130 , P2_R1146_U131 , P2_R1146_U132 , P2_R1146_U133 , P2_R1146_U134 , P2_R1146_U135 , P2_R1146_U136 , P2_R1146_U137;
wire P2_R1146_U138 , P2_R1146_U139 , P2_R1146_U140 , P2_R1146_U141 , P2_R1146_U142 , P2_R1146_U143 , P2_R1146_U144 , P2_R1146_U145 , P2_R1146_U146 , P2_R1146_U147;
wire P2_R1146_U148 , P2_R1146_U149 , P2_R1146_U150 , P2_R1146_U151 , P2_R1146_U152 , P2_R1146_U153 , P2_R1146_U154 , P2_R1146_U155 , P2_R1146_U156 , P2_R1146_U157;
wire P2_R1146_U158 , P2_R1146_U159 , P2_R1146_U160 , P2_R1146_U161 , P2_R1146_U162 , P2_R1146_U163 , P2_R1146_U164 , P2_R1146_U165 , P2_R1146_U166 , P2_R1146_U167;
wire P2_R1146_U168 , P2_R1146_U169 , P2_R1146_U170 , P2_R1146_U171 , P2_R1146_U172 , P2_R1146_U173 , P2_R1146_U174 , P2_R1146_U175 , P2_R1146_U176 , P2_R1146_U177;
wire P2_R1146_U178 , P2_R1146_U179 , P2_R1146_U180 , P2_R1146_U181 , P2_R1146_U182 , P2_R1146_U183 , P2_R1146_U184 , P2_R1146_U185 , P2_R1146_U186 , P2_R1146_U187;
wire P2_R1146_U188 , P2_R1146_U189 , P2_R1146_U190 , P2_R1146_U191 , P2_R1146_U192 , P2_R1146_U193 , P2_R1146_U194 , P2_R1146_U195 , P2_R1146_U196 , P2_R1146_U197;
wire P2_R1146_U198 , P2_R1146_U199 , P2_R1146_U200 , P2_R1146_U201 , P2_R1146_U202 , P2_R1146_U203 , P2_R1146_U204 , P2_R1146_U205 , P2_R1146_U206 , P2_R1146_U207;
wire P2_R1146_U208 , P2_R1146_U209 , P2_R1146_U210 , P2_R1146_U211 , P2_R1146_U212 , P2_R1146_U213 , P2_R1146_U214 , P2_R1146_U215 , P2_R1146_U216 , P2_R1146_U217;
wire P2_R1146_U218 , P2_R1146_U219 , P2_R1146_U220 , P2_R1146_U221 , P2_R1146_U222 , P2_R1146_U223 , P2_R1146_U224 , P2_R1146_U225 , P2_R1146_U226 , P2_R1146_U227;
wire P2_R1146_U228 , P2_R1146_U229 , P2_R1146_U230 , P2_R1146_U231 , P2_R1146_U232 , P2_R1146_U233 , P2_R1146_U234 , P2_R1146_U235 , P2_R1146_U236 , P2_R1146_U237;
wire P2_R1146_U238 , P2_R1146_U239 , P2_R1146_U240 , P2_R1146_U241 , P2_R1146_U242 , P2_R1146_U243 , P2_R1146_U244 , P2_R1146_U245 , P2_R1146_U246 , P2_R1146_U247;
wire P2_R1146_U248 , P2_R1146_U249 , P2_R1146_U250 , P2_R1146_U251 , P2_R1146_U252 , P2_R1146_U253 , P2_R1146_U254 , P2_R1146_U255 , P2_R1146_U256 , P2_R1146_U257;
wire P2_R1146_U258 , P2_R1146_U259 , P2_R1146_U260 , P2_R1146_U261 , P2_R1146_U262 , P2_R1146_U263 , P2_R1146_U264 , P2_R1146_U265 , P2_R1146_U266 , P2_R1146_U267;
wire P2_R1146_U268 , P2_R1146_U269 , P2_R1146_U270 , P2_R1146_U271 , P2_R1146_U272 , P2_R1146_U273 , P2_R1146_U274 , P2_R1146_U275 , P2_R1146_U276 , P2_R1146_U277;
wire P2_R1146_U278 , P2_R1146_U279 , P2_R1146_U280 , P2_R1146_U281 , P2_R1146_U282 , P2_R1146_U283 , P2_R1146_U284 , P2_R1146_U285 , P2_R1146_U286 , P2_R1146_U287;
wire P2_R1146_U288 , P2_R1146_U289 , P2_R1146_U290 , P2_R1146_U291 , P2_R1146_U292 , P2_R1146_U293 , P2_R1146_U294 , P2_R1146_U295 , P2_R1146_U296 , P2_R1146_U297;
wire P2_R1146_U298 , P2_R1146_U299 , P2_R1146_U300 , P2_R1146_U301 , P2_R1146_U302 , P2_R1146_U303 , P2_R1146_U304 , P2_R1146_U305 , P2_R1146_U306 , P2_R1146_U307;
wire P2_R1146_U308 , P2_R1146_U309 , P2_R1146_U310 , P2_R1146_U311 , P2_R1146_U312 , P2_R1146_U313 , P2_R1146_U314 , P2_R1146_U315 , P2_R1146_U316 , P2_R1146_U317;
wire P2_R1146_U318 , P2_R1146_U319 , P2_R1146_U320 , P2_R1146_U321 , P2_R1146_U322 , P2_R1146_U323 , P2_R1146_U324 , P2_R1146_U325 , P2_R1146_U326 , P2_R1146_U327;
wire P2_R1146_U328 , P2_R1146_U329 , P2_R1146_U330 , P2_R1146_U331 , P2_R1146_U332 , P2_R1146_U333 , P2_R1146_U334 , P2_R1146_U335 , P2_R1146_U336 , P2_R1146_U337;
wire P2_R1146_U338 , P2_R1146_U339 , P2_R1146_U340 , P2_R1146_U341 , P2_R1146_U342 , P2_R1146_U343 , P2_R1146_U344 , P2_R1146_U345 , P2_R1146_U346 , P2_R1146_U347;
wire P2_R1146_U348 , P2_R1146_U349 , P2_R1146_U350 , P2_R1146_U351 , P2_R1146_U352 , P2_R1146_U353 , P2_R1146_U354 , P2_R1146_U355 , P2_R1146_U356 , P2_R1146_U357;
wire P2_R1146_U358 , P2_R1146_U359 , P2_R1146_U360 , P2_R1146_U361 , P2_R1146_U362 , P2_R1146_U363 , P2_R1146_U364 , P2_R1146_U365 , P2_R1146_U366 , P2_R1146_U367;
wire P2_R1146_U368 , P2_R1146_U369 , P2_R1146_U370 , P2_R1146_U371 , P2_R1146_U372 , P2_R1146_U373 , P2_R1146_U374 , P2_R1146_U375 , P2_R1146_U376 , P2_R1146_U377;
wire P2_R1146_U378 , P2_R1146_U379 , P2_R1146_U380 , P2_R1146_U381 , P2_R1146_U382 , P2_R1146_U383 , P2_R1146_U384 , P2_R1146_U385 , P2_R1146_U386 , P2_R1146_U387;
wire P2_R1146_U388 , P2_R1146_U389 , P2_R1146_U390 , P2_R1146_U391 , P2_R1146_U392 , P2_R1146_U393 , P2_R1146_U394 , P2_R1146_U395 , P2_R1146_U396 , P2_R1146_U397;
wire P2_R1146_U398 , P2_R1146_U399 , P2_R1146_U400 , P2_R1146_U401 , P2_R1146_U402 , P2_R1146_U403 , P2_R1146_U404 , P2_R1146_U405 , P2_R1146_U406 , P2_R1146_U407;
wire P2_R1146_U408 , P2_R1146_U409 , P2_R1146_U410 , P2_R1146_U411 , P2_R1146_U412 , P2_R1146_U413 , P2_R1146_U414 , P2_R1146_U415 , P2_R1146_U416 , P2_R1146_U417;
wire P2_R1146_U418 , P2_R1146_U419 , P2_R1146_U420 , P2_R1146_U421 , P2_R1146_U422 , P2_R1146_U423 , P2_R1146_U424 , P2_R1146_U425 , P2_R1146_U426 , P2_R1146_U427;
wire P2_R1146_U428 , P2_R1146_U429 , P2_R1146_U430 , P2_R1146_U431 , P2_R1146_U432 , P2_R1146_U433 , P2_R1146_U434 , P2_R1146_U435 , P2_R1146_U436 , P2_R1146_U437;
wire P2_R1146_U438 , P2_R1146_U439 , P2_R1146_U440 , P2_R1146_U441 , P2_R1146_U442 , P2_R1146_U443 , P2_R1146_U444 , P2_R1146_U445 , P2_R1146_U446 , P2_R1146_U447;
wire P2_R1146_U448 , P2_R1146_U449 , P2_R1146_U450 , P2_R1146_U451 , P2_R1146_U452 , P2_R1146_U453 , P2_R1146_U454 , P2_R1146_U455 , P2_R1146_U456 , P2_R1146_U457;
wire P2_R1146_U458 , P2_R1146_U459 , P2_R1146_U460 , P2_R1146_U461 , P2_R1146_U462 , P2_R1146_U463 , P2_R1146_U464 , P2_R1146_U465 , P2_R1146_U466 , P2_R1146_U467;
wire P2_R1146_U468 , P2_R1146_U469 , P2_R1146_U470 , P2_R1146_U471 , P2_R1146_U472 , P2_R1146_U473 , P2_R1146_U474 , P2_R1146_U475 , P2_R1146_U476 , P2_R1146_U477;
wire P2_R1203_U6 , P2_R1203_U7 , P2_R1203_U8 , P2_R1203_U9 , P2_R1203_U10 , P2_R1203_U11 , P2_R1203_U12 , P2_R1203_U13 , P2_R1203_U14 , P2_R1203_U15;
wire P2_R1203_U16 , P2_R1203_U17 , P2_R1203_U18 , P2_R1203_U19 , P2_R1203_U20 , P2_R1203_U21 , P2_R1203_U22 , P2_R1203_U23 , P2_R1203_U24 , P2_R1203_U25;
wire P2_R1203_U26 , P2_R1203_U27 , P2_R1203_U28 , P2_R1203_U29 , P2_R1203_U30 , P2_R1203_U31 , P2_R1203_U32 , P2_R1203_U33 , P2_R1203_U34 , P2_R1203_U35;
wire P2_R1203_U36 , P2_R1203_U37 , P2_R1203_U38 , P2_R1203_U39 , P2_R1203_U40 , P2_R1203_U41 , P2_R1203_U42 , P2_R1203_U43 , P2_R1203_U44 , P2_R1203_U45;
wire P2_R1203_U46 , P2_R1203_U47 , P2_R1203_U48 , P2_R1203_U49 , P2_R1203_U50 , P2_R1203_U51 , P2_R1203_U52 , P2_R1203_U53 , P2_R1203_U54 , P2_R1203_U55;
wire P2_R1203_U56 , P2_R1203_U57 , P2_R1203_U58 , P2_R1203_U59 , P2_R1203_U60 , P2_R1203_U61 , P2_R1203_U62 , P2_R1203_U63 , P2_R1203_U64 , P2_R1203_U65;
wire P2_R1203_U66 , P2_R1203_U67 , P2_R1203_U68 , P2_R1203_U69 , P2_R1203_U70 , P2_R1203_U71 , P2_R1203_U72 , P2_R1203_U73 , P2_R1203_U74 , P2_R1203_U75;
wire P2_R1203_U76 , P2_R1203_U77 , P2_R1203_U78 , P2_R1203_U79 , P2_R1203_U80 , P2_R1203_U81 , P2_R1203_U82 , P2_R1203_U83 , P2_R1203_U84 , P2_R1203_U85;
wire P2_R1203_U86 , P2_R1203_U87 , P2_R1203_U88 , P2_R1203_U89 , P2_R1203_U90 , P2_R1203_U91 , P2_R1203_U92 , P2_R1203_U93 , P2_R1203_U94 , P2_R1203_U95;
wire P2_R1203_U96 , P2_R1203_U97 , P2_R1203_U98 , P2_R1203_U99 , P2_R1203_U100 , P2_R1203_U101 , P2_R1203_U102 , P2_R1203_U103 , P2_R1203_U104 , P2_R1203_U105;
wire P2_R1203_U106 , P2_R1203_U107 , P2_R1203_U108 , P2_R1203_U109 , P2_R1203_U110 , P2_R1203_U111 , P2_R1203_U112 , P2_R1203_U113 , P2_R1203_U114 , P2_R1203_U115;
wire P2_R1203_U116 , P2_R1203_U117 , P2_R1203_U118 , P2_R1203_U119 , P2_R1203_U120 , P2_R1203_U121 , P2_R1203_U122 , P2_R1203_U123 , P2_R1203_U124 , P2_R1203_U125;
wire P2_R1203_U126 , P2_R1203_U127 , P2_R1203_U128 , P2_R1203_U129 , P2_R1203_U130 , P2_R1203_U131 , P2_R1203_U132 , P2_R1203_U133 , P2_R1203_U134 , P2_R1203_U135;
wire P2_R1203_U136 , P2_R1203_U137 , P2_R1203_U138 , P2_R1203_U139 , P2_R1203_U140 , P2_R1203_U141 , P2_R1203_U142 , P2_R1203_U143 , P2_R1203_U144 , P2_R1203_U145;
wire P2_R1203_U146 , P2_R1203_U147 , P2_R1203_U148 , P2_R1203_U149 , P2_R1203_U150 , P2_R1203_U151 , P2_R1203_U152 , P2_R1203_U153 , P2_R1203_U154 , P2_R1203_U155;
wire P2_R1203_U156 , P2_R1203_U157 , P2_R1203_U158 , P2_R1203_U159 , P2_R1203_U160 , P2_R1203_U161 , P2_R1203_U162 , P2_R1203_U163 , P2_R1203_U164 , P2_R1203_U165;
wire P2_R1203_U166 , P2_R1203_U167 , P2_R1203_U168 , P2_R1203_U169 , P2_R1203_U170 , P2_R1203_U171 , P2_R1203_U172 , P2_R1203_U173 , P2_R1203_U174 , P2_R1203_U175;
wire P2_R1203_U176 , P2_R1203_U177 , P2_R1203_U178 , P2_R1203_U179 , P2_R1203_U180 , P2_R1203_U181 , P2_R1203_U182 , P2_R1203_U183 , P2_R1203_U184 , P2_R1203_U185;
wire P2_R1203_U186 , P2_R1203_U187 , P2_R1203_U188 , P2_R1203_U189 , P2_R1203_U190 , P2_R1203_U191 , P2_R1203_U192 , P2_R1203_U193 , P2_R1203_U194 , P2_R1203_U195;
wire P2_R1203_U196 , P2_R1203_U197 , P2_R1203_U198 , P2_R1203_U199 , P2_R1203_U200 , P2_R1203_U201 , P2_R1203_U202 , P2_R1203_U203 , P2_R1203_U204 , P2_R1203_U205;
wire P2_R1203_U206 , P2_R1203_U207 , P2_R1203_U208 , P2_R1203_U209 , P2_R1203_U210 , P2_R1203_U211 , P2_R1203_U212 , P2_R1203_U213 , P2_R1203_U214 , P2_R1203_U215;
wire P2_R1203_U216 , P2_R1203_U217 , P2_R1203_U218 , P2_R1203_U219 , P2_R1203_U220 , P2_R1203_U221 , P2_R1203_U222 , P2_R1203_U223 , P2_R1203_U224 , P2_R1203_U225;
wire P2_R1203_U226 , P2_R1203_U227 , P2_R1203_U228 , P2_R1203_U229 , P2_R1203_U230 , P2_R1203_U231 , P2_R1203_U232 , P2_R1203_U233 , P2_R1203_U234 , P2_R1203_U235;
wire P2_R1203_U236 , P2_R1203_U237 , P2_R1203_U238 , P2_R1203_U239 , P2_R1203_U240 , P2_R1203_U241 , P2_R1203_U242 , P2_R1203_U243 , P2_R1203_U244 , P2_R1203_U245;
wire P2_R1203_U246 , P2_R1203_U247 , P2_R1203_U248 , P2_R1203_U249 , P2_R1203_U250 , P2_R1203_U251 , P2_R1203_U252 , P2_R1203_U253 , P2_R1203_U254 , P2_R1203_U255;
wire P2_R1203_U256 , P2_R1203_U257 , P2_R1203_U258 , P2_R1203_U259 , P2_R1203_U260 , P2_R1203_U261 , P2_R1203_U262 , P2_R1203_U263 , P2_R1203_U264 , P2_R1203_U265;
wire P2_R1203_U266 , P2_R1203_U267 , P2_R1203_U268 , P2_R1203_U269 , P2_R1203_U270 , P2_R1203_U271 , P2_R1203_U272 , P2_R1203_U273 , P2_R1203_U274 , P2_R1203_U275;
wire P2_R1203_U276 , P2_R1203_U277 , P2_R1203_U278 , P2_R1203_U279 , P2_R1203_U280 , P2_R1203_U281 , P2_R1203_U282 , P2_R1203_U283 , P2_R1203_U284 , P2_R1203_U285;
wire P2_R1203_U286 , P2_R1203_U287 , P2_R1203_U288 , P2_R1203_U289 , P2_R1203_U290 , P2_R1203_U291 , P2_R1203_U292 , P2_R1203_U293 , P2_R1203_U294 , P2_R1203_U295;
wire P2_R1203_U296 , P2_R1203_U297 , P2_R1203_U298 , P2_R1203_U299 , P2_R1203_U300 , P2_R1203_U301 , P2_R1203_U302 , P2_R1203_U303 , P2_R1203_U304 , P2_R1203_U305;
wire P2_R1203_U306 , P2_R1203_U307 , P2_R1203_U308 , P2_R1203_U309 , P2_R1203_U310 , P2_R1203_U311 , P2_R1203_U312 , P2_R1203_U313 , P2_R1203_U314 , P2_R1203_U315;
wire P2_R1203_U316 , P2_R1203_U317 , P2_R1203_U318 , P2_R1203_U319 , P2_R1203_U320 , P2_R1203_U321 , P2_R1203_U322 , P2_R1203_U323 , P2_R1203_U324 , P2_R1203_U325;
wire P2_R1203_U326 , P2_R1203_U327 , P2_R1203_U328 , P2_R1203_U329 , P2_R1203_U330 , P2_R1203_U331 , P2_R1203_U332 , P2_R1203_U333 , P2_R1203_U334 , P2_R1203_U335;
wire P2_R1203_U336 , P2_R1203_U337 , P2_R1203_U338 , P2_R1203_U339 , P2_R1203_U340 , P2_R1203_U341 , P2_R1203_U342 , P2_R1203_U343 , P2_R1203_U344 , P2_R1203_U345;
wire P2_R1203_U346 , P2_R1203_U347 , P2_R1203_U348 , P2_R1203_U349 , P2_R1203_U350 , P2_R1203_U351 , P2_R1203_U352 , P2_R1203_U353 , P2_R1203_U354 , P2_R1203_U355;
wire P2_R1203_U356 , P2_R1203_U357 , P2_R1203_U358 , P2_R1203_U359 , P2_R1203_U360 , P2_R1203_U361 , P2_R1203_U362 , P2_R1203_U363 , P2_R1203_U364 , P2_R1203_U365;
wire P2_R1203_U366 , P2_R1203_U367 , P2_R1203_U368 , P2_R1203_U369 , P2_R1203_U370 , P2_R1203_U371 , P2_R1203_U372 , P2_R1203_U373 , P2_R1203_U374 , P2_R1203_U375;
wire P2_R1203_U376 , P2_R1203_U377 , P2_R1203_U378 , P2_R1203_U379 , P2_R1203_U380 , P2_R1203_U381 , P2_R1203_U382 , P2_R1203_U383 , P2_R1203_U384 , P2_R1203_U385;
wire P2_R1203_U386 , P2_R1203_U387 , P2_R1203_U388 , P2_R1203_U389 , P2_R1203_U390 , P2_R1203_U391 , P2_R1203_U392 , P2_R1203_U393 , P2_R1203_U394 , P2_R1203_U395;
wire P2_R1203_U396 , P2_R1203_U397 , P2_R1203_U398 , P2_R1203_U399 , P2_R1203_U400 , P2_R1203_U401 , P2_R1203_U402 , P2_R1203_U403 , P2_R1203_U404 , P2_R1203_U405;
wire P2_R1203_U406 , P2_R1203_U407 , P2_R1203_U408 , P2_R1203_U409 , P2_R1203_U410 , P2_R1203_U411 , P2_R1203_U412 , P2_R1203_U413 , P2_R1203_U414 , P2_R1203_U415;
wire P2_R1203_U416 , P2_R1203_U417 , P2_R1203_U418 , P2_R1203_U419 , P2_R1203_U420 , P2_R1203_U421 , P2_R1203_U422 , P2_R1203_U423 , P2_R1203_U424 , P2_R1203_U425;
wire P2_R1203_U426 , P2_R1203_U427 , P2_R1203_U428 , P2_R1203_U429 , P2_R1203_U430 , P2_R1203_U431 , P2_R1203_U432 , P2_R1203_U433 , P2_R1203_U434 , P2_R1203_U435;
wire P2_R1203_U436 , P2_R1203_U437 , P2_R1203_U438 , P2_R1203_U439 , P2_R1203_U440 , P2_R1203_U441 , P2_R1203_U442 , P2_R1203_U443 , P2_R1203_U444 , P2_R1203_U445;
wire P2_R1203_U446 , P2_R1203_U447 , P2_R1203_U448 , P2_R1203_U449 , P2_R1203_U450 , P2_R1203_U451 , P2_R1203_U452 , P2_R1203_U453 , P2_R1203_U454 , P2_R1203_U455;
wire P2_R1203_U456 , P2_R1203_U457 , P2_R1203_U458 , P2_R1203_U459 , P2_R1203_U460 , P2_R1203_U461 , P2_R1203_U462 , P2_R1203_U463 , P2_R1203_U464 , P2_R1203_U465;
wire P2_R1203_U466 , P2_R1203_U467 , P2_R1203_U468 , P2_R1203_U469 , P2_R1203_U470 , P2_R1203_U471 , P2_R1203_U472 , P2_R1203_U473 , P2_R1203_U474 , P2_R1203_U475;
wire P2_R1203_U476 , P2_R1203_U477 , P2_R1113_U6 , P2_R1113_U7 , P2_R1113_U8 , P2_R1113_U9 , P2_R1113_U10 , P2_R1113_U11 , P2_R1113_U12 , P2_R1113_U13;
wire P2_R1113_U14 , P2_R1113_U15 , P2_R1113_U16 , P2_R1113_U17 , P2_R1113_U18 , P2_R1113_U19 , P2_R1113_U20 , P2_R1113_U21 , P2_R1113_U22 , P2_R1113_U23;
wire P2_R1113_U24 , P2_R1113_U25 , P2_R1113_U26 , P2_R1113_U27 , P2_R1113_U28 , P2_R1113_U29 , P2_R1113_U30 , P2_R1113_U31 , P2_R1113_U32 , P2_R1113_U33;
wire P2_R1113_U34 , P2_R1113_U35 , P2_R1113_U36 , P2_R1113_U37 , P2_R1113_U38 , P2_R1113_U39 , P2_R1113_U40 , P2_R1113_U41 , P2_R1113_U42 , P2_R1113_U43;
wire P2_R1113_U44 , P2_R1113_U45 , P2_R1113_U46 , P2_R1113_U47 , P2_R1113_U48 , P2_R1113_U49 , P2_R1113_U50 , P2_R1113_U51 , P2_R1113_U52 , P2_R1113_U53;
wire P2_R1113_U54 , P2_R1113_U55 , P2_R1113_U56 , P2_R1113_U57 , P2_R1113_U58 , P2_R1113_U59 , P2_R1113_U60 , P2_R1113_U61 , P2_R1113_U62 , P2_R1113_U63;
wire P2_R1113_U64 , P2_R1113_U65 , P2_R1113_U66 , P2_R1113_U67 , P2_R1113_U68 , P2_R1113_U69 , P2_R1113_U70 , P2_R1113_U71 , P2_R1113_U72 , P2_R1113_U73;
wire P2_R1113_U74 , P2_R1113_U75 , P2_R1113_U76 , P2_R1113_U77 , P2_R1113_U78 , P2_R1113_U79 , P2_R1113_U80 , P2_R1113_U81 , P2_R1113_U82 , P2_R1113_U83;
wire P2_R1113_U84 , P2_R1113_U85 , P2_R1113_U86 , P2_R1113_U87 , P2_R1113_U88 , P2_R1113_U89 , P2_R1113_U90 , P2_R1113_U91 , P2_R1113_U92 , P2_R1113_U93;
wire P2_R1113_U94 , P2_R1113_U95 , P2_R1113_U96 , P2_R1113_U97 , P2_R1113_U98 , P2_R1113_U99 , P2_R1113_U100 , P2_R1113_U101 , P2_R1113_U102 , P2_R1113_U103;
wire P2_R1113_U104 , P2_R1113_U105 , P2_R1113_U106 , P2_R1113_U107 , P2_R1113_U108 , P2_R1113_U109 , P2_R1113_U110 , P2_R1113_U111 , P2_R1113_U112 , P2_R1113_U113;
wire P2_R1113_U114 , P2_R1113_U115 , P2_R1113_U116 , P2_R1113_U117 , P2_R1113_U118 , P2_R1113_U119 , P2_R1113_U120 , P2_R1113_U121 , P2_R1113_U122 , P2_R1113_U123;
wire P2_R1113_U124 , P2_R1113_U125 , P2_R1113_U126 , P2_R1113_U127 , P2_R1113_U128 , P2_R1113_U129 , P2_R1113_U130 , P2_R1113_U131 , P2_R1113_U132 , P2_R1113_U133;
wire P2_R1113_U134 , P2_R1113_U135 , P2_R1113_U136 , P2_R1113_U137 , P2_R1113_U138 , P2_R1113_U139 , P2_R1113_U140 , P2_R1113_U141 , P2_R1113_U142 , P2_R1113_U143;
wire P2_R1113_U144 , P2_R1113_U145 , P2_R1113_U146 , P2_R1113_U147 , P2_R1113_U148 , P2_R1113_U149 , P2_R1113_U150 , P2_R1113_U151 , P2_R1113_U152 , P2_R1113_U153;
wire P2_R1113_U154 , P2_R1113_U155 , P2_R1113_U156 , P2_R1113_U157 , P2_R1113_U158 , P2_R1113_U159 , P2_R1113_U160 , P2_R1113_U161 , P2_R1113_U162 , P2_R1113_U163;
wire P2_R1113_U164 , P2_R1113_U165 , P2_R1113_U166 , P2_R1113_U167 , P2_R1113_U168 , P2_R1113_U169 , P2_R1113_U170 , P2_R1113_U171 , P2_R1113_U172 , P2_R1113_U173;
wire P2_R1113_U174 , P2_R1113_U175 , P2_R1113_U176 , P2_R1113_U177 , P2_R1113_U178 , P2_R1113_U179 , P2_R1113_U180 , P2_R1113_U181 , P2_R1113_U182 , P2_R1113_U183;
wire P2_R1113_U184 , P2_R1113_U185 , P2_R1113_U186 , P2_R1113_U187 , P2_R1113_U188 , P2_R1113_U189 , P2_R1113_U190 , P2_R1113_U191 , P2_R1113_U192 , P2_R1113_U193;
wire P2_R1113_U194 , P2_R1113_U195 , P2_R1113_U196 , P2_R1113_U197 , P2_R1113_U198 , P2_R1113_U199 , P2_R1113_U200 , P2_R1113_U201 , P2_R1113_U202 , P2_R1113_U203;
wire P2_R1113_U204 , P2_R1113_U205 , P2_R1113_U206 , P2_R1113_U207 , P2_R1113_U208 , P2_R1113_U209 , P2_R1113_U210 , P2_R1113_U211 , P2_R1113_U212 , P2_R1113_U213;
wire P2_R1113_U214 , P2_R1113_U215 , P2_R1113_U216 , P2_R1113_U217 , P2_R1113_U218 , P2_R1113_U219 , P2_R1113_U220 , P2_R1113_U221 , P2_R1113_U222 , P2_R1113_U223;
wire P2_R1113_U224 , P2_R1113_U225 , P2_R1113_U226 , P2_R1113_U227 , P2_R1113_U228 , P2_R1113_U229 , P2_R1113_U230 , P2_R1113_U231 , P2_R1113_U232 , P2_R1113_U233;
wire P2_R1113_U234 , P2_R1113_U235 , P2_R1113_U236 , P2_R1113_U237 , P2_R1113_U238 , P2_R1113_U239 , P2_R1113_U240 , P2_R1113_U241 , P2_R1113_U242 , P2_R1113_U243;
wire P2_R1113_U244 , P2_R1113_U245 , P2_R1113_U246 , P2_R1113_U247 , P2_R1113_U248 , P2_R1113_U249 , P2_R1113_U250 , P2_R1113_U251 , P2_R1113_U252 , P2_R1113_U253;
wire P2_R1113_U254 , P2_R1113_U255 , P2_R1113_U256 , P2_R1113_U257 , P2_R1113_U258 , P2_R1113_U259 , P2_R1113_U260 , P2_R1113_U261 , P2_R1113_U262 , P2_R1113_U263;
wire P2_R1113_U264 , P2_R1113_U265 , P2_R1113_U266 , P2_R1113_U267 , P2_R1113_U268 , P2_R1113_U269 , P2_R1113_U270 , P2_R1113_U271 , P2_R1113_U272 , P2_R1113_U273;
wire P2_R1113_U274 , P2_R1113_U275 , P2_R1113_U276 , P2_R1113_U277 , P2_R1113_U278 , P2_R1113_U279 , P2_R1113_U280 , P2_R1113_U281 , P2_R1113_U282 , P2_R1113_U283;
wire P2_R1113_U284 , P2_R1113_U285 , P2_R1113_U286 , P2_R1113_U287 , P2_R1113_U288 , P2_R1113_U289 , P2_R1113_U290 , P2_R1113_U291 , P2_R1113_U292 , P2_R1113_U293;
wire P2_R1113_U294 , P2_R1113_U295 , P2_R1113_U296 , P2_R1113_U297 , P2_R1113_U298 , P2_R1113_U299 , P2_R1113_U300 , P2_R1113_U301 , P2_R1113_U302 , P2_R1113_U303;
wire P2_R1113_U304 , P2_R1113_U305 , P2_R1113_U306 , P2_R1113_U307 , P2_R1113_U308 , P2_R1113_U309 , P2_R1113_U310 , P2_R1113_U311 , P2_R1113_U312 , P2_R1113_U313;
wire P2_R1113_U314 , P2_R1113_U315 , P2_R1113_U316 , P2_R1113_U317 , P2_R1113_U318 , P2_R1113_U319 , P2_R1113_U320 , P2_R1113_U321 , P2_R1113_U322 , P2_R1113_U323;
wire P2_R1113_U324 , P2_R1113_U325 , P2_R1113_U326 , P2_R1113_U327 , P2_R1113_U328 , P2_R1113_U329 , P2_R1113_U330 , P2_R1113_U331 , P2_R1113_U332 , P2_R1113_U333;
wire P2_R1113_U334 , P2_R1113_U335 , P2_R1113_U336 , P2_R1113_U337 , P2_R1113_U338 , P2_R1113_U339 , P2_R1113_U340 , P2_R1113_U341 , P2_R1113_U342 , P2_R1113_U343;
wire P2_R1113_U344 , P2_R1113_U345 , P2_R1113_U346 , P2_R1113_U347 , P2_R1113_U348 , P2_R1113_U349 , P2_R1113_U350 , P2_R1113_U351 , P2_R1113_U352 , P2_R1113_U353;
wire P2_R1113_U354 , P2_R1113_U355 , P2_R1113_U356 , P2_R1113_U357 , P2_R1113_U358 , P2_R1113_U359 , P2_R1113_U360 , P2_R1113_U361 , P2_R1113_U362 , P2_R1113_U363;
wire P2_R1113_U364 , P2_R1113_U365 , P2_R1113_U366 , P2_R1113_U367 , P2_R1113_U368 , P2_R1113_U369 , P2_R1113_U370 , P2_R1113_U371 , P2_R1113_U372 , P2_R1113_U373;
wire P2_R1113_U374 , P2_R1113_U375 , P2_R1113_U376 , P2_R1113_U377 , P2_R1113_U378 , P2_R1113_U379 , P2_R1113_U380 , P2_R1113_U381 , P2_R1113_U382 , P2_R1113_U383;
wire P2_R1113_U384 , P2_R1113_U385 , P2_R1113_U386 , P2_R1113_U387 , P2_R1113_U388 , P2_R1113_U389 , P2_R1113_U390 , P2_R1113_U391 , P2_R1113_U392 , P2_R1113_U393;
wire P2_R1113_U394 , P2_R1113_U395 , P2_R1113_U396 , P2_R1113_U397 , P2_R1113_U398 , P2_R1113_U399 , P2_R1113_U400 , P2_R1113_U401 , P2_R1113_U402 , P2_R1113_U403;
wire P2_R1113_U404 , P2_R1113_U405 , P2_R1113_U406 , P2_R1113_U407 , P2_R1113_U408 , P2_R1113_U409 , P2_R1113_U410 , P2_R1113_U411 , P2_R1113_U412 , P2_R1113_U413;
wire P2_R1113_U414 , P2_R1113_U415 , P2_R1113_U416 , P2_R1113_U417 , P2_R1113_U418;


nand NAND2_1 ( P2_R1113_U477 , P2_R1113_U176 , P2_R1113_U337 );
nand NAND2_2 ( P2_R1113_U476 , P2_R1113_U345 , P2_R1113_U88 );
nand NAND2_3 ( P2_R1113_U475 , P2_U3062 , P2_R1113_U47 );
nand NAND2_4 ( U25 , U136 , U135 );
nand NAND2_5 ( U26 , U138 , U137 );
nand NAND2_6 ( U27 , U140 , U139 );
nand NAND2_7 ( U28 , U142 , U141 );
nand NAND2_8 ( U29 , U144 , U143 );
nand NAND2_9 ( U30 , U146 , U145 );
nand NAND2_10 ( U31 , U148 , U147 );
nand NAND2_11 ( U32 , U150 , U149 );
nand NAND2_12 ( U33 , U152 , U151 );
nand NAND2_13 ( U34 , U154 , U153 );
nand NAND2_14 ( U35 , U156 , U155 );
nand NAND2_15 ( U36 , U158 , U157 );
nand NAND2_16 ( U37 , U160 , U159 );
nand NAND2_17 ( U38 , U162 , U161 );
nand NAND2_18 ( U39 , U164 , U163 );
nand NAND2_19 ( U40 , U166 , U165 );
nand NAND2_20 ( U41 , U168 , U167 );
nand NAND2_21 ( U42 , U170 , U169 );
nand NAND2_22 ( U43 , U172 , U171 );
nand NAND2_23 ( U44 , U174 , U173 );
nand NAND2_24 ( U45 , U176 , U175 );
nand NAND2_25 ( U46 , U178 , U177 );
nand NAND2_26 ( U47 , U180 , U179 );
nand NAND2_27 ( U48 , U182 , U181 );
nand NAND2_28 ( U49 , U184 , U183 );
nand NAND2_29 ( U50 , U186 , U185 );
nand NAND2_30 ( U51 , U188 , U187 );
nand NAND2_31 ( U52 , U190 , U189 );
nand NAND2_32 ( U53 , U192 , U191 );
nand NAND2_33 ( U54 , U194 , U193 );
nand NAND2_34 ( U55 , U196 , U195 );
nand NAND2_35 ( U56 , U198 , U197 );
nand NAND2_36 ( U57 , U200 , U199 );
nand NAND2_37 ( U58 , U202 , U201 );
nand NAND2_38 ( U59 , U204 , U203 );
nand NAND2_39 ( U60 , U206 , U205 );
nand NAND2_40 ( U61 , U208 , U207 );
nand NAND2_41 ( U62 , U210 , U209 );
nand NAND2_42 ( U63 , U212 , U211 );
nand NAND2_43 ( U64 , U214 , U213 );
nand NAND2_44 ( U65 , U216 , U215 );
nand NAND2_45 ( U66 , U218 , U217 );
nand NAND2_46 ( U67 , U220 , U219 );
nand NAND2_47 ( U68 , U222 , U221 );
nand NAND2_48 ( U69 , U224 , U223 );
nand NAND2_49 ( U70 , U226 , U225 );
nand NAND2_50 ( U71 , U228 , U227 );
nand NAND2_51 ( U72 , U230 , U229 );
nand NAND2_52 ( U73 , U232 , U231 );
nand NAND2_53 ( U74 , U234 , U233 );
nand NAND2_54 ( U75 , U236 , U235 );
nand NAND2_55 ( U76 , U238 , U237 );
nand NAND2_56 ( U77 , U240 , U239 );
nand NAND2_57 ( U78 , U242 , U241 );
nand NAND2_58 ( U79 , U244 , U243 );
nand NAND2_59 ( U80 , U246 , U245 );
nand NAND2_60 ( U81 , U248 , U247 );
nand NAND2_61 ( U82 , U250 , U249 );
nand NAND2_62 ( U83 , U252 , U251 );
nand NAND2_63 ( U84 , U254 , U253 );
nand NAND2_64 ( U85 , U256 , U255 );
nand NAND2_65 ( U86 , U258 , U257 );
nand NAND2_66 ( U87 , U260 , U259 );
nand NAND2_67 ( U88 , U262 , U261 );
nand NAND2_68 ( U89 , U264 , U263 );
nand NAND2_69 ( U90 , U266 , U265 );
nand NAND2_70 ( U91 , U268 , U267 );
nand NAND2_71 ( U92 , U270 , U269 );
nand NAND2_72 ( U93 , U272 , U271 );
nand NAND2_73 ( U94 , U274 , U273 );
nand NAND2_74 ( U95 , U276 , U275 );
nand NAND2_75 ( U96 , U278 , U277 );
nand NAND2_76 ( U97 , U280 , U279 );
nand NAND2_77 ( U98 , U282 , U281 );
nand NAND2_78 ( U99 , U284 , U283 );
nand NAND2_79 ( U100 , U286 , U285 );
nand NAND2_80 ( U101 , U288 , U287 );
nand NAND2_81 ( U102 , U290 , U289 );
nand NAND2_82 ( U103 , U292 , U291 );
nand NAND2_83 ( U104 , U294 , U293 );
nand NAND2_84 ( U105 , U296 , U295 );
nand NAND2_85 ( U106 , U298 , U297 );
nand NAND2_86 ( U107 , U300 , U299 );
nand NAND2_87 ( U108 , U302 , U301 );
nand NAND2_88 ( U109 , U304 , U303 );
nand NAND2_89 ( U110 , U306 , U305 );
nand NAND2_90 ( U111 , U308 , U307 );
nand NAND2_91 ( U112 , U310 , U309 );
nand NAND2_92 ( U113 , U312 , U311 );
nand NAND2_93 ( U114 , U314 , U313 );
nand NAND2_94 ( U115 , U316 , U315 );
nand NAND2_95 ( U116 , U318 , U317 );
nand NAND2_96 ( U117 , U320 , U319 );
nand NAND2_97 ( U118 , U322 , U321 );
nand NAND2_98 ( U119 , U324 , U323 );
nand NAND2_99 ( U120 , U326 , U325 );
not NOT1_100 ( U121 , P2_WR_REG );
not NOT1_101 ( U122 , P1_WR_REG );
and AND2_102 ( U123 , U132 , U131 );
not NOT1_103 ( U124 , P2_RD_REG );
not NOT1_104 ( U125 , P1_RD_REG );
and AND2_105 ( U126 , U134 , U133 );
nand NAND2_106 ( U127 , U129 , U128 );
nand NAND3_107 ( U128 , LT_1079_U6 , U125 , LT_1079_19_U6 );
nand NAND3_108 ( U129 , P1_ADDR_REG_19_ , U124 , P2_ADDR_REG_19_ );
not NOT1_109 ( U130 , U127 );
nand NAND2_110 ( U131 , P2_WR_REG , U122 );
nand NAND2_111 ( U132 , P1_WR_REG , U121 );
nand NAND2_112 ( U133 , P2_RD_REG , U125 );
nand NAND2_113 ( U134 , P1_RD_REG , U124 );
nand NAND2_114 ( U135 , P1_DATAO_REG_9_ , U127 );
nand NAND2_115 ( U136 , R140_U84 , U130 );
nand NAND2_116 ( U137 , P1_DATAO_REG_8_ , U127 );
nand NAND2_117 ( U138 , R140_U85 , U130 );
nand NAND2_118 ( U139 , P1_DATAO_REG_7_ , U127 );
nand NAND2_119 ( U140 , R140_U86 , U130 );
nand NAND2_120 ( U141 , P1_DATAO_REG_6_ , U127 );
nand NAND2_121 ( U142 , R140_U87 , U130 );
nand NAND2_122 ( U143 , P1_DATAO_REG_5_ , U127 );
nand NAND2_123 ( U144 , R140_U88 , U130 );
nand NAND2_124 ( U145 , P1_DATAO_REG_4_ , U127 );
nand NAND2_125 ( U146 , R140_U89 , U130 );
nand NAND2_126 ( U147 , P1_DATAO_REG_3_ , U127 );
nand NAND2_127 ( U148 , R140_U90 , U130 );
nand NAND2_128 ( U149 , P1_DATAO_REG_31_ , U127 );
nand NAND2_129 ( U150 , R140_U11 , U130 );
nand NAND2_130 ( U151 , P1_DATAO_REG_30_ , U127 );
nand NAND2_131 ( U152 , R140_U91 , U130 );
nand NAND2_132 ( U153 , P1_DATAO_REG_2_ , U127 );
nand NAND2_133 ( U154 , R140_U92 , U130 );
nand NAND2_134 ( U155 , P1_DATAO_REG_29_ , U127 );
nand NAND2_135 ( U156 , R140_U93 , U130 );
nand NAND2_136 ( U157 , P1_DATAO_REG_28_ , U127 );
nand NAND2_137 ( U158 , R140_U94 , U130 );
nand NAND2_138 ( U159 , P1_DATAO_REG_27_ , U127 );
nand NAND2_139 ( U160 , R140_U95 , U130 );
nand NAND2_140 ( U161 , P1_DATAO_REG_26_ , U127 );
nand NAND2_141 ( U162 , R140_U96 , U130 );
nand NAND2_142 ( U163 , P1_DATAO_REG_25_ , U127 );
nand NAND2_143 ( U164 , R140_U97 , U130 );
nand NAND2_144 ( U165 , P1_DATAO_REG_24_ , U127 );
nand NAND2_145 ( U166 , R140_U98 , U130 );
nand NAND2_146 ( U167 , P1_DATAO_REG_23_ , U127 );
nand NAND2_147 ( U168 , R140_U99 , U130 );
nand NAND2_148 ( U169 , P1_DATAO_REG_22_ , U127 );
nand NAND2_149 ( U170 , R140_U100 , U130 );
nand NAND2_150 ( U171 , P1_DATAO_REG_21_ , U127 );
nand NAND2_151 ( U172 , R140_U101 , U130 );
nand NAND2_152 ( U173 , P1_DATAO_REG_20_ , U127 );
nand NAND2_153 ( U174 , R140_U102 , U130 );
nand NAND2_154 ( U175 , P1_DATAO_REG_1_ , U127 );
nand NAND2_155 ( U176 , R140_U10 , U130 );
nand NAND2_156 ( U177 , P1_DATAO_REG_19_ , U127 );
nand NAND2_157 ( U178 , R140_U103 , U130 );
nand NAND2_158 ( U179 , P1_DATAO_REG_18_ , U127 );
nand NAND2_159 ( U180 , R140_U104 , U130 );
nand NAND2_160 ( U181 , P1_DATAO_REG_17_ , U127 );
nand NAND2_161 ( U182 , R140_U105 , U130 );
nand NAND2_162 ( U183 , P1_DATAO_REG_16_ , U127 );
nand NAND2_163 ( U184 , R140_U106 , U130 );
nand NAND2_164 ( U185 , P1_DATAO_REG_15_ , U127 );
nand NAND2_165 ( U186 , R140_U107 , U130 );
nand NAND2_166 ( U187 , P1_DATAO_REG_14_ , U127 );
nand NAND2_167 ( U188 , R140_U108 , U130 );
nand NAND2_168 ( U189 , P1_DATAO_REG_13_ , U127 );
nand NAND2_169 ( U190 , R140_U109 , U130 );
nand NAND2_170 ( U191 , P1_DATAO_REG_12_ , U127 );
nand NAND2_171 ( U192 , R140_U110 , U130 );
nand NAND2_172 ( U193 , P1_DATAO_REG_11_ , U127 );
nand NAND2_173 ( U194 , R140_U111 , U130 );
nand NAND2_174 ( U195 , P1_DATAO_REG_10_ , U127 );
nand NAND2_175 ( U196 , R140_U112 , U130 );
nand NAND2_176 ( U197 , P1_DATAO_REG_0_ , U127 );
nand NAND2_177 ( U198 , R140_U83 , U130 );
nand NAND2_178 ( U199 , R140_U84 , U127 );
nand NAND2_179 ( U200 , P2_DATAO_REG_9_ , U130 );
nand NAND2_180 ( U201 , R140_U85 , U127 );
nand NAND2_181 ( U202 , P2_DATAO_REG_8_ , U130 );
nand NAND2_182 ( U203 , R140_U86 , U127 );
nand NAND2_183 ( U204 , P2_DATAO_REG_7_ , U130 );
nand NAND2_184 ( U205 , R140_U87 , U127 );
nand NAND2_185 ( U206 , P2_DATAO_REG_6_ , U130 );
nand NAND2_186 ( U207 , R140_U88 , U127 );
nand NAND2_187 ( U208 , P2_DATAO_REG_5_ , U130 );
nand NAND2_188 ( U209 , R140_U89 , U127 );
nand NAND2_189 ( U210 , P2_DATAO_REG_4_ , U130 );
nand NAND2_190 ( U211 , R140_U90 , U127 );
nand NAND2_191 ( U212 , P2_DATAO_REG_3_ , U130 );
nand NAND2_192 ( U213 , R140_U11 , U127 );
nand NAND2_193 ( U214 , P2_DATAO_REG_31_ , U130 );
nand NAND2_194 ( U215 , R140_U91 , U127 );
nand NAND2_195 ( U216 , P2_DATAO_REG_30_ , U130 );
nand NAND2_196 ( U217 , R140_U92 , U127 );
nand NAND2_197 ( U218 , P2_DATAO_REG_2_ , U130 );
nand NAND2_198 ( U219 , R140_U93 , U127 );
nand NAND2_199 ( U220 , P2_DATAO_REG_29_ , U130 );
nand NAND2_200 ( U221 , R140_U94 , U127 );
nand NAND2_201 ( U222 , P2_DATAO_REG_28_ , U130 );
nand NAND2_202 ( U223 , R140_U95 , U127 );
nand NAND2_203 ( U224 , P2_DATAO_REG_27_ , U130 );
nand NAND2_204 ( U225 , R140_U96 , U127 );
nand NAND2_205 ( U226 , P2_DATAO_REG_26_ , U130 );
nand NAND2_206 ( U227 , R140_U97 , U127 );
nand NAND2_207 ( U228 , P2_DATAO_REG_25_ , U130 );
nand NAND2_208 ( U229 , R140_U98 , U127 );
nand NAND2_209 ( U230 , P2_DATAO_REG_24_ , U130 );
nand NAND2_210 ( U231 , R140_U99 , U127 );
nand NAND2_211 ( U232 , P2_DATAO_REG_23_ , U130 );
nand NAND2_212 ( U233 , R140_U100 , U127 );
nand NAND2_213 ( U234 , P2_DATAO_REG_22_ , U130 );
nand NAND2_214 ( U235 , R140_U101 , U127 );
nand NAND2_215 ( U236 , P2_DATAO_REG_21_ , U130 );
nand NAND2_216 ( U237 , R140_U102 , U127 );
nand NAND2_217 ( U238 , P2_DATAO_REG_20_ , U130 );
nand NAND2_218 ( U239 , R140_U10 , U127 );
nand NAND2_219 ( U240 , P2_DATAO_REG_1_ , U130 );
nand NAND2_220 ( U241 , R140_U103 , U127 );
nand NAND2_221 ( U242 , P2_DATAO_REG_19_ , U130 );
nand NAND2_222 ( U243 , R140_U104 , U127 );
nand NAND2_223 ( U244 , P2_DATAO_REG_18_ , U130 );
nand NAND2_224 ( U245 , R140_U105 , U127 );
nand NAND2_225 ( U246 , P2_DATAO_REG_17_ , U130 );
nand NAND2_226 ( U247 , R140_U106 , U127 );
nand NAND2_227 ( U248 , P2_DATAO_REG_16_ , U130 );
nand NAND2_228 ( U249 , R140_U107 , U127 );
nand NAND2_229 ( U250 , P2_DATAO_REG_15_ , U130 );
nand NAND2_230 ( U251 , R140_U108 , U127 );
nand NAND2_231 ( U252 , P2_DATAO_REG_14_ , U130 );
nand NAND2_232 ( U253 , R140_U109 , U127 );
nand NAND2_233 ( U254 , P2_DATAO_REG_13_ , U130 );
nand NAND2_234 ( U255 , R140_U110 , U127 );
nand NAND2_235 ( U256 , P2_DATAO_REG_12_ , U130 );
nand NAND2_236 ( U257 , R140_U111 , U127 );
nand NAND2_237 ( U258 , P2_DATAO_REG_11_ , U130 );
nand NAND2_238 ( U259 , R140_U112 , U127 );
nand NAND2_239 ( U260 , P2_DATAO_REG_10_ , U130 );
nand NAND2_240 ( U261 , R140_U83 , U127 );
nand NAND2_241 ( U262 , P2_DATAO_REG_0_ , U130 );
nand NAND2_242 ( U263 , P2_DATAO_REG_9_ , U127 );
nand NAND2_243 ( U264 , U130 , P1_DATAO_REG_9_ );
nand NAND2_244 ( U265 , P2_DATAO_REG_8_ , U127 );
nand NAND2_245 ( U266 , P1_DATAO_REG_8_ , U130 );
nand NAND2_246 ( U267 , P2_DATAO_REG_7_ , U127 );
nand NAND2_247 ( U268 , P1_DATAO_REG_7_ , U130 );
nand NAND2_248 ( U269 , P2_DATAO_REG_6_ , U127 );
nand NAND2_249 ( U270 , P1_DATAO_REG_6_ , U130 );
nand NAND2_250 ( U271 , P2_DATAO_REG_5_ , U127 );
nand NAND2_251 ( U272 , P1_DATAO_REG_5_ , U130 );
nand NAND2_252 ( U273 , P2_DATAO_REG_4_ , U127 );
nand NAND2_253 ( U274 , P1_DATAO_REG_4_ , U130 );
nand NAND2_254 ( U275 , P2_DATAO_REG_31_ , U127 );
nand NAND2_255 ( U276 , P1_DATAO_REG_31_ , U130 );
nand NAND2_256 ( U277 , P2_DATAO_REG_30_ , U127 );
nand NAND2_257 ( U278 , P1_DATAO_REG_30_ , U130 );
nand NAND2_258 ( U279 , P2_DATAO_REG_3_ , U127 );
nand NAND2_259 ( U280 , P1_DATAO_REG_3_ , U130 );
nand NAND2_260 ( U281 , P2_DATAO_REG_29_ , U127 );
nand NAND2_261 ( U282 , P1_DATAO_REG_29_ , U130 );
nand NAND2_262 ( U283 , P2_DATAO_REG_28_ , U127 );
nand NAND2_263 ( U284 , P1_DATAO_REG_28_ , U130 );
nand NAND2_264 ( U285 , P2_DATAO_REG_27_ , U127 );
nand NAND2_265 ( U286 , P1_DATAO_REG_27_ , U130 );
nand NAND2_266 ( U287 , P2_DATAO_REG_26_ , U127 );
nand NAND2_267 ( U288 , P1_DATAO_REG_26_ , U130 );
nand NAND2_268 ( U289 , P2_DATAO_REG_25_ , U127 );
nand NAND2_269 ( U290 , P1_DATAO_REG_25_ , U130 );
nand NAND2_270 ( U291 , P2_DATAO_REG_24_ , U127 );
nand NAND2_271 ( U292 , P1_DATAO_REG_24_ , U130 );
nand NAND2_272 ( U293 , P2_DATAO_REG_23_ , U127 );
nand NAND2_273 ( U294 , P1_DATAO_REG_23_ , U130 );
nand NAND2_274 ( U295 , P2_DATAO_REG_22_ , U127 );
nand NAND2_275 ( U296 , P1_DATAO_REG_22_ , U130 );
nand NAND2_276 ( U297 , P2_DATAO_REG_21_ , U127 );
nand NAND2_277 ( U298 , P1_DATAO_REG_21_ , U130 );
nand NAND2_278 ( U299 , P2_DATAO_REG_20_ , U127 );
nand NAND2_279 ( U300 , P1_DATAO_REG_20_ , U130 );
nand NAND2_280 ( U301 , P2_DATAO_REG_2_ , U127 );
nand NAND2_281 ( U302 , P1_DATAO_REG_2_ , U130 );
nand NAND2_282 ( U303 , P2_DATAO_REG_19_ , U127 );
nand NAND2_283 ( U304 , P1_DATAO_REG_19_ , U130 );
nand NAND2_284 ( U305 , P2_DATAO_REG_18_ , U127 );
nand NAND2_285 ( U306 , P1_DATAO_REG_18_ , U130 );
nand NAND2_286 ( U307 , P2_DATAO_REG_17_ , U127 );
nand NAND2_287 ( U308 , P1_DATAO_REG_17_ , U130 );
nand NAND2_288 ( U309 , P2_DATAO_REG_16_ , U127 );
nand NAND2_289 ( U310 , P1_DATAO_REG_16_ , U130 );
nand NAND2_290 ( U311 , P2_DATAO_REG_15_ , U127 );
nand NAND2_291 ( U312 , P1_DATAO_REG_15_ , U130 );
nand NAND2_292 ( U313 , P2_DATAO_REG_14_ , U127 );
nand NAND2_293 ( U314 , P1_DATAO_REG_14_ , U130 );
nand NAND2_294 ( U315 , P2_DATAO_REG_13_ , U127 );
nand NAND2_295 ( U316 , P1_DATAO_REG_13_ , U130 );
nand NAND2_296 ( U317 , P2_DATAO_REG_12_ , U127 );
nand NAND2_297 ( U318 , P1_DATAO_REG_12_ , U130 );
nand NAND2_298 ( U319 , P2_DATAO_REG_11_ , U127 );
nand NAND2_299 ( U320 , P1_DATAO_REG_11_ , U130 );
nand NAND2_300 ( U321 , P2_DATAO_REG_10_ , U127 );
nand NAND2_301 ( U322 , P1_DATAO_REG_10_ , U130 );
nand NAND2_302 ( U323 , P2_DATAO_REG_1_ , U127 );
nand NAND2_303 ( U324 , P1_DATAO_REG_1_ , U130 );
nand NAND2_304 ( U325 , P2_DATAO_REG_0_ , U127 );
nand NAND2_305 ( U326 , P1_DATAO_REG_0_ , U130 );
nand NAND2_306 ( P2_R1113_U474 , P2_U3480 , P2_R1113_U50 );
nand NAND2_307 ( P2_R1113_U473 , P2_R1113_U472 , P2_R1113_U471 );
nand NAND2_308 ( P2_R1113_U472 , P2_U3063 , P2_R1113_U48 );
nand NAND2_309 ( P2_R1113_U471 , P2_U3483 , P2_R1113_U49 );
nand NAND2_310 ( P2_R1113_U470 , P2_R1113_U144 , P2_R1113_U175 );
nand NAND2_311 ( P2_R1113_U469 , P2_R1113_U250 , P2_R1113_U468 );
not NOT1_312 ( P2_R1113_U468 , P2_R1113_U144 );
nand NAND2_313 ( P2_R1113_U467 , P2_U3072 , P2_R1113_U52 );
nand NAND2_314 ( P2_R1113_U466 , P2_U3486 , P2_R1113_U53 );
nand NAND2_315 ( P2_R1113_U465 , P2_R1113_U143 , P2_R1113_U174 );
nand NAND2_316 ( P2_R1113_U464 , P2_R1113_U254 , P2_R1113_U463 );
not NOT1_317 ( P2_R1113_U463 , P2_R1113_U143 );
and AND2_318 ( P1_U3014 , P1_U3989 , P1_U3444 );
and AND2_319 ( P1_U3015 , P1_U3450 , P1_U3447 );
and AND2_320 ( P1_U3016 , P1_U3632 , P1_U3627 );
and AND2_321 ( P1_U3017 , P1_U3445 , P1_U3446 );
and AND2_322 ( P1_U3018 , P1_U5725 , P1_U3445 );
and AND2_323 ( P1_U3019 , P1_U5722 , P1_U3446 );
and AND2_324 ( P1_U3020 , P1_U5722 , P1_U5725 );
and AND2_325 ( P1_U3021 , P1_U5400 , P1_U3421 );
and AND2_326 ( P1_U3022 , P1_U3046 , P1_STATE_REG );
and AND2_327 ( P1_U3023 , P1_U3049 , P1_U5716 );
and AND2_328 ( P1_U3024 , P1_U3817 , P1_U3423 );
and AND2_329 ( P1_U3025 , P1_U4020 , P1_U5728 );
and AND2_330 ( P1_U3026 , P1_U3986 , P1_U5716 );
and AND2_331 ( P1_U3027 , P1_U3880 , P1_U4005 );
and AND2_332 ( P1_U3028 , P1_U3356 , P1_STATE_REG );
and AND2_333 ( P1_U3029 , P1_U3997 , P1_U4022 );
and AND2_334 ( P1_U3030 , P1_U4022 , P1_U3422 );
and AND2_335 ( P1_U3031 , P1_U3990 , P1_U4022 );
and AND2_336 ( P1_U3032 , P1_U3998 , P1_U4022 );
and AND2_337 ( P1_U3033 , P1_U4020 , P1_U3447 );
and AND2_338 ( P1_U3034 , P1_U4005 , P1_U5728 );
and AND2_339 ( P1_U3035 , P1_U4022 , P1_U3025 );
and AND2_340 ( P1_U3036 , P1_U4005 , P1_U3447 );
and AND2_341 ( P1_U3037 , P1_U5734 , P1_U4913 );
and AND2_342 ( P1_U3038 , P1_U3024 , P1_U5734 );
and AND2_343 ( P1_U3039 , P1_U5728 , P1_U4913 );
and AND2_344 ( P1_U3040 , P1_U3024 , P1_U5728 );
and AND2_345 ( P1_U3041 , P1_U3015 , P1_U4913 );
and AND2_346 ( P1_U3042 , P1_U3024 , P1_U3015 );
and AND2_347 ( P1_U3043 , P1_U3022 , P1_U3423 );
and AND2_348 ( P1_U3044 , P1_U5145 , P1_STATE_REG );
and AND2_349 ( P1_U3045 , P1_U3022 , P1_U5147 );
and AND2_350 ( P1_U3046 , P1_U5703 , P1_U3421 );
and AND2_351 ( P1_U3047 , P1_U3633 , P1_U3016 );
and AND2_352 ( P1_U3048 , P1_U5716 , P1_U3443 );
and AND2_353 ( P1_U3049 , P1_U5710 , P1_U5719 );
and AND2_354 ( P1_U3050 , P1_U3436 , P1_U3438 );
nand NAND4_355 ( P1_U3051 , P1_U4670 , P1_U4671 , P1_U4669 , P1_U4672 );
nand NAND4_356 ( P1_U3052 , P1_U4689 , P1_U4690 , P1_U4688 , P1_U4691 );
nand NAND4_357 ( P1_U3053 , P1_U4710 , P1_U4709 , P1_U4708 , P1_U4707 );
nand NAND3_358 ( P1_U3054 , P1_U4747 , P1_U4748 , P1_U4746 );
nand NAND4_359 ( P1_U3055 , P1_U4651 , P1_U4652 , P1_U4650 , P1_U4653 );
nand NAND4_360 ( P1_U3056 , P1_U4632 , P1_U4633 , P1_U4631 , P1_U4634 );
nand NAND3_361 ( P1_U3057 , P1_U4727 , P1_U4728 , P1_U4726 );
nand NAND4_362 ( P1_U3058 , P1_U4235 , P1_U4234 , P1_U4233 , P1_U4232 );
nand NAND4_363 ( P1_U3059 , P1_U4575 , P1_U4576 , P1_U4574 , P1_U4577 );
nand NAND4_364 ( P1_U3060 , P1_U4347 , P1_U4348 , P1_U4346 , P1_U4349 );
nand NAND4_365 ( P1_U3061 , P1_U4366 , P1_U4367 , P1_U4365 , P1_U4368 );
nand NAND4_366 ( P1_U3062 , P1_U4216 , P1_U4215 , P1_U4214 , P1_U4213 );
nand NAND4_367 ( P1_U3063 , P1_U4613 , P1_U4614 , P1_U4612 , P1_U4615 );
nand NAND4_368 ( P1_U3064 , P1_U4594 , P1_U4595 , P1_U4593 , P1_U4596 );
nand NAND4_369 ( P1_U3065 , P1_U4254 , P1_U4253 , P1_U4252 , P1_U4251 );
nand NAND4_370 ( P1_U3066 , P1_U4192 , P1_U4191 , P1_U4190 , P1_U4189 );
nand NAND4_371 ( P1_U3067 , P1_U4480 , P1_U4481 , P1_U4479 , P1_U4482 );
nand NAND4_372 ( P1_U3068 , P1_U4292 , P1_U4291 , P1_U4290 , P1_U4289 );
nand NAND4_373 ( P1_U3069 , P1_U4273 , P1_U4272 , P1_U4271 , P1_U4270 );
nand NAND4_374 ( P1_U3070 , P1_U4385 , P1_U4386 , P1_U4384 , P1_U4387 );
nand NAND4_375 ( P1_U3071 , P1_U4461 , P1_U4462 , P1_U4460 , P1_U4463 );
nand NAND4_376 ( P1_U3072 , P1_U4442 , P1_U4443 , P1_U4441 , P1_U4444 );
nand NAND4_377 ( P1_U3073 , P1_U4556 , P1_U4557 , P1_U4555 , P1_U4558 );
nand NAND4_378 ( P1_U3074 , P1_U4537 , P1_U4538 , P1_U4536 , P1_U4539 );
nand NAND4_379 ( P1_U3075 , P1_U4197 , P1_U4196 , P1_U4195 , P1_U4194 );
nand NAND4_380 ( P1_U3076 , P1_U4173 , P1_U4172 , P1_U4171 , P1_U4170 );
nand NAND4_381 ( P1_U3077 , P1_U4423 , P1_U4424 , P1_U4422 , P1_U4425 );
nand NAND4_382 ( P1_U3078 , P1_U4404 , P1_U4405 , P1_U4403 , P1_U4406 );
nand NAND4_383 ( P1_U3079 , P1_U4518 , P1_U4519 , P1_U4517 , P1_U4520 );
nand NAND4_384 ( P1_U3080 , P1_U4499 , P1_U4500 , P1_U4498 , P1_U4501 );
nand NAND4_385 ( P1_U3081 , P1_U4328 , P1_U4329 , P1_U4327 , P1_U4330 );
nand NAND4_386 ( P1_U3082 , P1_U4311 , P1_U4310 , P1_U4309 , P1_U4308 );
nand NAND2_387 ( P1_U3083 , P1_U4920 , P1_STATE_REG );
not NOT1_388 ( P1_U3084 , P1_STATE_REG );
nand NAND2_389 ( P1_U3085 , P1_U5608 , P1_U5607 );
nand NAND2_390 ( P1_U3086 , P1_U5610 , P1_U5609 );
nand NAND3_391 ( P1_U3087 , P1_U5615 , P1_U5614 , P1_U5616 );
nand NAND2_392 ( P1_U3088 , P1_U3923 , P1_U5618 );
nand NAND2_393 ( P1_U3089 , P1_U3924 , P1_U5621 );
nand NAND2_394 ( P1_U3090 , P1_U3925 , P1_U5624 );
nand NAND2_395 ( P1_U3091 , P1_U3926 , P1_U5627 );
nand NAND2_396 ( P1_U3092 , P1_U3927 , P1_U5630 );
nand NAND2_397 ( P1_U3093 , P1_U3928 , P1_U5633 );
nand NAND2_398 ( P1_U3094 , P1_U3929 , P1_U5636 );
nand NAND2_399 ( P1_U3095 , P1_U3930 , P1_U5639 );
nand NAND2_400 ( P1_U3096 , P1_U3931 , P1_U5642 );
nand NAND2_401 ( P1_U3097 , P1_U3933 , P1_U5648 );
nand NAND2_402 ( P1_U3098 , P1_U3934 , P1_U5651 );
nand NAND2_403 ( P1_U3099 , P1_U3935 , P1_U5654 );
nand NAND2_404 ( P1_U3100 , P1_U3936 , P1_U5657 );
nand NAND2_405 ( P1_U3101 , P1_U3937 , P1_U5660 );
nand NAND2_406 ( P1_U3102 , P1_U3938 , P1_U5663 );
nand NAND2_407 ( P1_U3103 , P1_U3939 , P1_U5666 );
nand NAND2_408 ( P1_U3104 , P1_U3940 , P1_U5669 );
nand NAND2_409 ( P1_U3105 , P1_U3941 , P1_U5672 );
nand NAND2_410 ( P1_U3106 , P1_U3942 , P1_U5675 );
nand NAND3_411 ( P1_U3107 , P1_U5590 , P1_U5591 , P1_U5589 );
nand NAND3_412 ( P1_U3108 , P1_U5593 , P1_U5594 , P1_U5592 );
nand NAND3_413 ( P1_U3109 , P1_U5596 , P1_U5597 , P1_U5595 );
nand NAND3_414 ( P1_U3110 , P1_U5599 , P1_U5600 , P1_U5598 );
nand NAND3_415 ( P1_U3111 , P1_U5602 , P1_U5603 , P1_U5601 );
nand NAND2_416 ( P1_U3112 , P1_U3921 , P1_U5605 );
nand NAND2_417 ( P1_U3113 , P1_U3922 , P1_U5612 );
nand NAND2_418 ( P1_U3114 , P1_U3932 , P1_U5645 );
nand NAND2_419 ( P1_U3115 , P1_U3943 , P1_U5678 );
nand NAND2_420 ( P1_U3116 , P1_U5681 , P1_U5680 );
nand NAND2_421 ( P1_U3117 , P1_U5538 , P1_U5537 );
nand NAND2_422 ( P1_U3118 , P1_U5540 , P1_U5539 );
nand NAND2_423 ( P1_U3119 , P1_U3898 , P1_U5543 );
nand NAND2_424 ( P1_U3120 , P1_U3899 , P1_U5545 );
nand NAND2_425 ( P1_U3121 , P1_U3900 , P1_U5547 );
nand NAND2_426 ( P1_U3122 , P1_U3901 , P1_U5549 );
nand NAND2_427 ( P1_U3123 , P1_U3902 , P1_U5551 );
nand NAND2_428 ( P1_U3124 , P1_U3903 , P1_U5553 );
nand NAND2_429 ( P1_U3125 , P1_U3904 , P1_U5555 );
nand NAND2_430 ( P1_U3126 , P1_U3905 , P1_U5557 );
nand NAND2_431 ( P1_U3127 , P1_U3906 , P1_U5559 );
nand NAND2_432 ( P1_U3128 , P1_U3907 , P1_U5561 );
nand NAND2_433 ( P1_U3129 , P1_U3909 , P1_U5566 );
nand NAND2_434 ( P1_U3130 , P1_U3910 , P1_U5568 );
nand NAND2_435 ( P1_U3131 , P1_U3911 , P1_U5570 );
nand NAND2_436 ( P1_U3132 , P1_U3912 , P1_U5572 );
nand NAND2_437 ( P1_U3133 , P1_U3913 , P1_U5574 );
nand NAND2_438 ( P1_U3134 , P1_U3914 , P1_U5576 );
nand NAND2_439 ( P1_U3135 , P1_U3915 , P1_U5578 );
nand NAND2_440 ( P1_U3136 , P1_U3916 , P1_U5580 );
nand NAND2_441 ( P1_U3137 , P1_U3917 , P1_U5582 );
nand NAND2_442 ( P1_U3138 , P1_U3918 , P1_U5584 );
nand NAND3_443 ( P1_U3139 , P1_U5526 , P1_U3439 , P1_U5525 );
nand NAND3_444 ( P1_U3140 , P1_U5528 , P1_U3439 , P1_U5527 );
nand NAND3_445 ( P1_U3141 , P1_U5530 , P1_U3439 , P1_U5529 );
nand NAND3_446 ( P1_U3142 , P1_U5532 , P1_U3439 , P1_U5531 );
nand NAND3_447 ( P1_U3143 , P1_U5534 , P1_U3439 , P1_U5533 );
nand NAND2_448 ( P1_U3144 , P1_U3896 , P1_U5536 );
nand NAND2_449 ( P1_U3145 , P1_U3897 , P1_U5542 );
nand NAND2_450 ( P1_U3146 , P1_U3908 , P1_U5564 );
nand NAND2_451 ( P1_U3147 , P1_U3919 , P1_U5586 );
nand NAND2_452 ( P1_U3148 , P1_U3920 , P1_U5588 );
nand NAND2_453 ( P1_U3149 , P1_U3986 , P1_U3439 );
nand NAND2_454 ( P1_U3150 , P1_U5703 , P1_U3371 );
nand NAND2_455 ( P1_U3151 , P1_U5480 , P1_U5479 );
nand NAND2_456 ( P1_U3152 , P1_U5482 , P1_U5481 );
nand NAND2_457 ( P1_U3153 , P1_U5484 , P1_U5483 );
nand NAND2_458 ( P1_U3154 , P1_U5486 , P1_U5485 );
nand NAND2_459 ( P1_U3155 , P1_U5488 , P1_U5487 );
nand NAND2_460 ( P1_U3156 , P1_U5490 , P1_U5489 );
nand NAND2_461 ( P1_U3157 , P1_U5492 , P1_U5491 );
nand NAND2_462 ( P1_U3158 , P1_U5494 , P1_U5493 );
nand NAND2_463 ( P1_U3159 , P1_U5496 , P1_U5495 );
nand NAND2_464 ( P1_U3160 , P1_U5500 , P1_U5499 );
nand NAND2_465 ( P1_U3161 , P1_U5502 , P1_U5501 );
nand NAND2_466 ( P1_U3162 , P1_U5504 , P1_U5503 );
nand NAND2_467 ( P1_U3163 , P1_U5506 , P1_U5505 );
nand NAND2_468 ( P1_U3164 , P1_U5508 , P1_U5507 );
nand NAND2_469 ( P1_U3165 , P1_U5510 , P1_U5509 );
nand NAND2_470 ( P1_U3166 , P1_U5512 , P1_U5511 );
nand NAND2_471 ( P1_U3167 , P1_U5514 , P1_U5513 );
nand NAND2_472 ( P1_U3168 , P1_U5516 , P1_U5515 );
nand NAND2_473 ( P1_U3169 , P1_U5518 , P1_U5517 );
nand NAND2_474 ( P1_U3170 , P1_U5466 , P1_U5465 );
nand NAND2_475 ( P1_U3171 , P1_U5468 , P1_U5467 );
nand NAND2_476 ( P1_U3172 , P1_U5470 , P1_U5469 );
nand NAND2_477 ( P1_U3173 , P1_U5472 , P1_U5471 );
nand NAND2_478 ( P1_U3174 , P1_U5474 , P1_U5473 );
nand NAND2_479 ( P1_U3175 , P1_U5476 , P1_U5475 );
nand NAND2_480 ( P1_U3176 , P1_U5478 , P1_U5477 );
nand NAND2_481 ( P1_U3177 , P1_U5498 , P1_U5497 );
nand NAND2_482 ( P1_U3178 , P1_U5520 , P1_U5519 );
nand NAND2_483 ( P1_U3179 , P1_U3895 , P1_U5522 );
nand NAND2_484 ( P1_U3180 , P1_U5421 , P1_U5420 );
nand NAND2_485 ( P1_U3181 , P1_U5423 , P1_U5422 );
nand NAND2_486 ( P1_U3182 , P1_U5425 , P1_U5424 );
nand NAND2_487 ( P1_U3183 , P1_U5427 , P1_U5426 );
nand NAND2_488 ( P1_U3184 , P1_U5429 , P1_U5428 );
nand NAND2_489 ( P1_U3185 , P1_U5431 , P1_U5430 );
nand NAND2_490 ( P1_U3186 , P1_U5433 , P1_U5432 );
nand NAND2_491 ( P1_U3187 , P1_U5435 , P1_U5434 );
nand NAND2_492 ( P1_U3188 , P1_U5437 , P1_U5436 );
nand NAND2_493 ( P1_U3189 , P1_U5441 , P1_U5440 );
nand NAND2_494 ( P1_U3190 , P1_U5443 , P1_U5442 );
nand NAND2_495 ( P1_U3191 , P1_U5445 , P1_U5444 );
nand NAND2_496 ( P1_U3192 , P1_U5447 , P1_U5446 );
nand NAND2_497 ( P1_U3193 , P1_U5449 , P1_U5448 );
nand NAND2_498 ( P1_U3194 , P1_U5451 , P1_U5450 );
nand NAND2_499 ( P1_U3195 , P1_U5453 , P1_U5452 );
nand NAND2_500 ( P1_U3196 , P1_U5455 , P1_U5454 );
nand NAND2_501 ( P1_U3197 , P1_U5457 , P1_U5456 );
nand NAND2_502 ( P1_U3198 , P1_U5459 , P1_U5458 );
nand NAND2_503 ( P1_U3199 , P1_U5407 , P1_U5406 );
nand NAND2_504 ( P1_U3200 , P1_U5409 , P1_U5408 );
nand NAND2_505 ( P1_U3201 , P1_U5411 , P1_U5410 );
nand NAND2_506 ( P1_U3202 , P1_U5413 , P1_U5412 );
nand NAND2_507 ( P1_U3203 , P1_U5415 , P1_U5414 );
nand NAND2_508 ( P1_U3204 , P1_U5417 , P1_U5416 );
nand NAND2_509 ( P1_U3205 , P1_U5419 , P1_U5418 );
nand NAND2_510 ( P1_U3206 , P1_U5439 , P1_U5438 );
nand NAND2_511 ( P1_U3207 , P1_U5461 , P1_U5460 );
nand NAND2_512 ( P1_U3208 , P1_U3894 , P1_U5462 );
and AND2_513 ( P1_U3209 , P1_U5399 , P1_U3421 );
nand NAND3_514 ( P1_U3210 , P1_U6266 , P1_U6265 , P1_U5397 );
nand NAND5_515 ( P1_U3211 , P1_U5391 , P1_U5390 , P1_U5394 , P1_U5392 , P1_U5393 );
nand NAND5_516 ( P1_U3212 , P1_U5382 , P1_U5381 , P1_U5385 , P1_U5383 , P1_U5384 );
nand NAND5_517 ( P1_U3213 , P1_U5373 , P1_U5372 , P1_U5376 , P1_U5374 , P1_U5375 );
nand NAND5_518 ( P1_U3214 , P1_U5364 , P1_U5363 , P1_U5367 , P1_U5365 , P1_U5366 );
nand NAND5_519 ( P1_U3215 , P1_U5355 , P1_U5354 , P1_U5358 , P1_U5356 , P1_U5357 );
nand NAND3_520 ( P1_U3216 , P1_U3891 , P1_U5346 , P1_U5347 );
nand NAND5_521 ( P1_U3217 , P1_U5337 , P1_U5336 , P1_U5340 , P1_U5338 , P1_U5339 );
nand NAND5_522 ( P1_U3218 , P1_U5328 , P1_U5327 , P1_U5331 , P1_U5329 , P1_U5330 );
nand NAND5_523 ( P1_U3219 , P1_U5319 , P1_U5318 , P1_U5322 , P1_U5320 , P1_U5321 );
nand NAND3_524 ( P1_U3220 , P1_U3889 , P1_U5310 , P1_U5311 );
nand NAND5_525 ( P1_U3221 , P1_U5301 , P1_U5300 , P1_U5304 , P1_U5302 , P1_U5303 );
nand NAND5_526 ( P1_U3222 , P1_U5292 , P1_U5291 , P1_U5295 , P1_U5293 , P1_U5294 );
nand NAND5_527 ( P1_U3223 , P1_U5283 , P1_U5282 , P1_U5286 , P1_U5284 , P1_U5285 );
nand NAND5_528 ( P1_U3224 , P1_U5274 , P1_U5273 , P1_U5277 , P1_U5275 , P1_U5276 );
nand NAND4_529 ( P1_U3225 , P1_U5265 , P1_U5264 , P1_U5266 , P1_U3888 );
nand NAND5_530 ( P1_U3226 , P1_U5256 , P1_U5255 , P1_U5259 , P1_U5257 , P1_U5258 );
nand NAND5_531 ( P1_U3227 , P1_U5247 , P1_U5246 , P1_U5250 , P1_U5248 , P1_U5249 );
nand NAND3_532 ( P1_U3228 , P1_U3886 , P1_U5238 , P1_U5239 );
nand NAND5_533 ( P1_U3229 , P1_U5229 , P1_U5228 , P1_U5232 , P1_U5230 , P1_U5231 );
nand NAND3_534 ( P1_U3230 , P1_U3885 , P1_U5221 , P1_U3884 );
nand NAND5_535 ( P1_U3231 , P1_U5212 , P1_U5211 , P1_U5215 , P1_U5213 , P1_U5214 );
nand NAND5_536 ( P1_U3232 , P1_U5203 , P1_U5202 , P1_U5206 , P1_U5204 , P1_U5205 );
nand NAND5_537 ( P1_U3233 , P1_U5194 , P1_U5193 , P1_U5197 , P1_U5195 , P1_U5196 );
nand NAND5_538 ( P1_U3234 , P1_U5185 , P1_U5184 , P1_U5188 , P1_U5186 , P1_U5187 );
nand NAND3_539 ( P1_U3235 , P1_U3881 , P1_U5176 , P1_U5177 );
nand NAND5_540 ( P1_U3236 , P1_U5167 , P1_U5166 , P1_U5170 , P1_U5168 , P1_U5169 );
nand NAND5_541 ( P1_U3237 , P1_U5158 , P1_U5157 , P1_U5161 , P1_U5159 , P1_U5160 );
nand NAND5_542 ( P1_U3238 , P1_U5149 , P1_U5148 , P1_U5152 , P1_U5150 , P1_U5151 );
nand NAND5_543 ( P1_U3239 , P1_U5136 , P1_U5135 , P1_U5139 , P1_U5137 , P1_U5138 );
and AND2_544 ( P1_U3240 , P1_U5120 , P1_U5682 );
nand NAND2_545 ( P1_U3241 , P1_U3859 , P1_U3858 );
nand NAND2_546 ( P1_U3242 , P1_U3857 , P1_U3856 );
nand NAND2_547 ( P1_U3243 , P1_U3855 , P1_U3854 );
nand NAND2_548 ( P1_U3244 , P1_U3852 , P1_U3851 );
nand NAND2_549 ( P1_U3245 , P1_U3850 , P1_U3849 );
nand NAND2_550 ( P1_U3246 , P1_U3847 , P1_U3846 );
nand NAND2_551 ( P1_U3247 , P1_U3845 , P1_U3844 );
nand NAND3_552 ( P1_U3248 , P1_U3842 , P1_U3843 , P1_U5043 );
nand NAND3_553 ( P1_U3249 , P1_U3840 , P1_U3841 , P1_U5033 );
nand NAND3_554 ( P1_U3250 , P1_U3838 , P1_U3839 , P1_U5023 );
nand NAND3_555 ( P1_U3251 , P1_U3836 , P1_U3837 , P1_U5013 );
nand NAND3_556 ( P1_U3252 , P1_U3834 , P1_U3835 , P1_U5003 );
nand NAND3_557 ( P1_U3253 , P1_U3832 , P1_U3833 , P1_U4993 );
nand NAND3_558 ( P1_U3254 , P1_U3830 , P1_U3831 , P1_U4983 );
nand NAND3_559 ( P1_U3255 , P1_U3828 , P1_U3829 , P1_U4973 );
nand NAND3_560 ( P1_U3256 , P1_U3826 , P1_U3827 , P1_U4963 );
nand NAND3_561 ( P1_U3257 , P1_U3824 , P1_U3825 , P1_U4953 );
nand NAND3_562 ( P1_U3258 , P1_U3822 , P1_U3823 , P1_U4943 );
nand NAND3_563 ( P1_U3259 , P1_U3820 , P1_U3821 , P1_U4933 );
nand NAND3_564 ( P1_U3260 , P1_U3818 , P1_U3819 , P1_U4923 );
nand NAND3_565 ( P1_U3261 , P1_U3981 , P1_U4911 , P1_U4912 );
nand NAND3_566 ( P1_U3262 , P1_U3980 , P1_U4909 , P1_U4910 );
nand NAND4_567 ( P1_U3263 , P1_U3811 , P1_U3812 , P1_U4902 , P1_U3977 );
nand NAND4_568 ( P1_U3264 , P1_U3809 , P1_U3810 , P1_U4897 , P1_U3976 );
nand NAND4_569 ( P1_U3265 , P1_U3807 , P1_U3808 , P1_U4892 , P1_U3975 );
nand NAND4_570 ( P1_U3266 , P1_U3805 , P1_U3806 , P1_U4887 , P1_U3974 );
nand NAND4_571 ( P1_U3267 , P1_U3803 , P1_U3804 , P1_U4882 , P1_U3973 );
nand NAND4_572 ( P1_U3268 , P1_U3801 , P1_U3802 , P1_U4877 , P1_U3972 );
nand NAND4_573 ( P1_U3269 , P1_U3799 , P1_U3800 , P1_U4872 , P1_U3971 );
nand NAND4_574 ( P1_U3270 , P1_U3797 , P1_U3798 , P1_U4867 , P1_U3970 );
nand NAND4_575 ( P1_U3271 , P1_U3795 , P1_U3796 , P1_U4862 , P1_U3969 );
nand NAND4_576 ( P1_U3272 , P1_U3793 , P1_U3794 , P1_U4857 , P1_U3968 );
nand NAND3_577 ( P1_U3273 , P1_U3792 , P1_U3791 , P1_U3967 );
nand NAND3_578 ( P1_U3274 , P1_U3790 , P1_U3789 , P1_U3966 );
nand NAND4_579 ( P1_U3275 , P1_U3787 , P1_U3788 , P1_U4842 , P1_U3965 );
nand NAND4_580 ( P1_U3276 , P1_U3785 , P1_U3786 , P1_U4837 , P1_U3964 );
nand NAND3_581 ( P1_U3277 , P1_U3784 , P1_U3783 , P1_U3963 );
nand NAND3_582 ( P1_U3278 , P1_U3782 , P1_U3781 , P1_U3962 );
nand NAND3_583 ( P1_U3279 , P1_U3780 , P1_U3779 , P1_U3961 );
nand NAND3_584 ( P1_U3280 , P1_U3778 , P1_U3777 , P1_U3960 );
nand NAND4_585 ( P1_U3281 , P1_U3775 , P1_U3776 , P1_U4812 , P1_U3959 );
nand NAND4_586 ( P1_U3282 , P1_U3773 , P1_U3774 , P1_U4807 , P1_U3958 );
nand NAND3_587 ( P1_U3283 , P1_U3772 , P1_U3771 , P1_U3957 );
nand NAND3_588 ( P1_U3284 , P1_U3770 , P1_U3769 , P1_U3956 );
nand NAND3_589 ( P1_U3285 , P1_U3768 , P1_U3767 , P1_U3955 );
nand NAND3_590 ( P1_U3286 , P1_U3766 , P1_U3765 , P1_U3954 );
nand NAND2_591 ( P1_U3287 , P1_U3764 , P1_U3763 );
nand NAND2_592 ( P1_U3288 , P1_U3762 , P1_U3761 );
nand NAND2_593 ( P1_U3289 , P1_U3760 , P1_U3759 );
nand NAND2_594 ( P1_U3290 , P1_U3758 , P1_U3757 );
nand NAND2_595 ( P1_U3291 , P1_U3756 , P1_U3755 );
and AND2_596 ( P1_U3292 , P1_D_REG_31_ , P1_U3945 );
and AND2_597 ( P1_U3293 , P1_D_REG_30_ , P1_U3945 );
and AND2_598 ( P1_U3294 , P1_D_REG_29_ , P1_U3945 );
and AND2_599 ( P1_U3295 , P1_D_REG_28_ , P1_U3945 );
and AND2_600 ( P1_U3296 , P1_D_REG_27_ , P1_U3945 );
and AND2_601 ( P1_U3297 , P1_D_REG_26_ , P1_U3945 );
and AND2_602 ( P1_U3298 , P1_D_REG_25_ , P1_U3945 );
and AND2_603 ( P1_U3299 , P1_D_REG_24_ , P1_U3945 );
and AND2_604 ( P1_U3300 , P1_D_REG_23_ , P1_U3945 );
and AND2_605 ( P1_U3301 , P1_D_REG_22_ , P1_U3945 );
and AND2_606 ( P1_U3302 , P1_D_REG_21_ , P1_U3945 );
and AND2_607 ( P1_U3303 , P1_D_REG_20_ , P1_U3945 );
and AND2_608 ( P1_U3304 , P1_D_REG_19_ , P1_U3945 );
and AND2_609 ( P1_U3305 , P1_D_REG_18_ , P1_U3945 );
and AND2_610 ( P1_U3306 , P1_D_REG_17_ , P1_U3945 );
and AND2_611 ( P1_U3307 , P1_D_REG_16_ , P1_U3945 );
and AND2_612 ( P1_U3308 , P1_D_REG_15_ , P1_U3945 );
and AND2_613 ( P1_U3309 , P1_D_REG_14_ , P1_U3945 );
and AND2_614 ( P1_U3310 , P1_D_REG_13_ , P1_U3945 );
and AND2_615 ( P1_U3311 , P1_D_REG_12_ , P1_U3945 );
and AND2_616 ( P1_U3312 , P1_D_REG_11_ , P1_U3945 );
and AND2_617 ( P1_U3313 , P1_D_REG_10_ , P1_U3945 );
and AND2_618 ( P1_U3314 , P1_D_REG_9_ , P1_U3945 );
and AND2_619 ( P1_U3315 , P1_D_REG_8_ , P1_U3945 );
and AND2_620 ( P1_U3316 , P1_D_REG_7_ , P1_U3945 );
and AND2_621 ( P1_U3317 , P1_D_REG_6_ , P1_U3945 );
and AND2_622 ( P1_U3318 , P1_D_REG_5_ , P1_U3945 );
and AND2_623 ( P1_U3319 , P1_D_REG_4_ , P1_U3945 );
and AND2_624 ( P1_U3320 , P1_D_REG_3_ , P1_U3945 );
and AND2_625 ( P1_U3321 , P1_D_REG_2_ , P1_U3945 );
nand NAND3_626 ( P1_U3322 , P1_U4132 , P1_U4133 , P1_U4131 );
nand NAND3_627 ( P1_U3323 , P1_U4129 , P1_U4130 , P1_U4128 );
nand NAND3_628 ( P1_U3324 , P1_U4126 , P1_U4127 , P1_U4125 );
nand NAND3_629 ( P1_U3325 , P1_U4123 , P1_U4124 , P1_U4122 );
nand NAND3_630 ( P1_U3326 , P1_U4120 , P1_U4121 , P1_U4119 );
nand NAND3_631 ( P1_U3327 , P1_U4117 , P1_U4118 , P1_U4116 );
nand NAND3_632 ( P1_U3328 , P1_U4114 , P1_U4115 , P1_U4113 );
nand NAND3_633 ( P1_U3329 , P1_U4111 , P1_U4112 , P1_U4110 );
nand NAND3_634 ( P1_U3330 , P1_U4108 , P1_U4109 , P1_U4107 );
nand NAND3_635 ( P1_U3331 , P1_U4105 , P1_U4106 , P1_U4104 );
nand NAND3_636 ( P1_U3332 , P1_U4102 , P1_U4103 , P1_U4101 );
nand NAND3_637 ( P1_U3333 , P1_U4099 , P1_U4100 , P1_U4098 );
nand NAND3_638 ( P1_U3334 , P1_U4096 , P1_U4097 , P1_U4095 );
nand NAND3_639 ( P1_U3335 , P1_U4093 , P1_U4094 , P1_U4092 );
nand NAND3_640 ( P1_U3336 , P1_U4090 , P1_U4091 , P1_U4089 );
nand NAND3_641 ( P1_U3337 , P1_U4087 , P1_U4088 , P1_U4086 );
nand NAND3_642 ( P1_U3338 , P1_U4084 , P1_U4085 , P1_U4083 );
nand NAND3_643 ( P1_U3339 , P1_U4081 , P1_U4082 , P1_U4080 );
nand NAND3_644 ( P1_U3340 , P1_U4078 , P1_U4079 , P1_U4077 );
nand NAND3_645 ( P1_U3341 , P1_U4075 , P1_U4076 , P1_U4074 );
nand NAND3_646 ( P1_U3342 , P1_U4072 , P1_U4073 , P1_U4071 );
nand NAND3_647 ( P1_U3343 , P1_U4069 , P1_U4070 , P1_U4068 );
nand NAND3_648 ( P1_U3344 , P1_U4066 , P1_U4067 , P1_U4065 );
nand NAND3_649 ( P1_U3345 , P1_U4063 , P1_U4064 , P1_U4062 );
nand NAND3_650 ( P1_U3346 , P1_U4060 , P1_U4061 , P1_U4059 );
nand NAND3_651 ( P1_U3347 , P1_U4057 , P1_U4058 , P1_U4056 );
nand NAND3_652 ( P1_U3348 , P1_U4054 , P1_U4055 , P1_U4053 );
nand NAND3_653 ( P1_U3349 , P1_U4051 , P1_U4052 , P1_U4050 );
nand NAND3_654 ( P1_U3350 , P1_U4048 , P1_U4049 , P1_U4047 );
nand NAND3_655 ( P1_U3351 , P1_U4045 , P1_U4046 , P1_U4044 );
nand NAND3_656 ( P1_U3352 , P1_U4042 , P1_U4043 , P1_U4041 );
nand NAND3_657 ( P1_U3353 , P1_U4039 , P1_U4040 , P1_U4038 );
and AND2_658 ( P1_U3354 , P1_U3443 , P1_U3439 );
nand NAND5_659 ( P1_U3355 , P1_U4907 , P1_U4905 , P1_U4908 , P1_U4906 , P1_U3978 );
nand NAND2_660 ( P1_U3356 , P1_STATE_REG , P1_U3944 );
nand NAND2_661 ( P1_U3357 , P1_U3438 , P1_U5695 );
not NOT1_662 ( P1_U3358 , P1_B_REG );
nand NAND3_663 ( P1_U3359 , P1_U5700 , P1_U5699 , P1_U3438 );
nand NAND2_664 ( P1_U3360 , P1_U3048 , P1_U3444 );
nand NAND3_665 ( P1_U3361 , P1_U3442 , P1_U3443 , P1_U3444 );
nand NAND2_666 ( P1_U3362 , P1_U3442 , P1_U5713 );
nand NAND2_667 ( P1_U3363 , P1_U4034 , P1_U3444 );
nand NAND3_668 ( P1_U3364 , P1_U3442 , P1_U3443 , P1_U3448 );
nand NAND2_669 ( P1_U3365 , P1_U4034 , P1_U3448 );
nand NAND2_670 ( P1_U3366 , P1_U5716 , P1_U5713 );
nand NAND2_671 ( P1_U3367 , P1_U4035 , P1_U3444 );
nand NAND2_672 ( P1_U3368 , P1_U3993 , P1_U5719 );
nand NAND2_673 ( P1_U3369 , P1_U4035 , P1_U3448 );
nand NAND2_674 ( P1_U3370 , P1_U3989 , P1_U5710 );
nand NAND2_675 ( P1_U3371 , P1_U5710 , P1_U3443 );
nand NAND2_676 ( P1_U3372 , P1_U3444 , P1_U3448 );
nand NAND5_677 ( P1_U3373 , P1_U4181 , P1_U4180 , P1_U4182 , P1_U3620 , P1_U3619 );
not NOT1_678 ( P1_U3374 , P1_REG2_REG_0_ );
nand NAND4_679 ( P1_U3375 , P1_U4200 , P1_U4199 , P1_U3635 , P1_U3637 );
nand NAND4_680 ( P1_U3376 , P1_U4219 , P1_U4218 , P1_U3639 , P1_U3641 );
nand NAND4_681 ( P1_U3377 , P1_U4238 , P1_U4237 , P1_U3643 , P1_U3645 );
nand NAND4_682 ( P1_U3378 , P1_U4257 , P1_U4256 , P1_U3647 , P1_U3649 );
nand NAND4_683 ( P1_U3379 , P1_U4276 , P1_U4275 , P1_U3651 , P1_U3653 );
nand NAND4_684 ( P1_U3380 , P1_U4295 , P1_U4294 , P1_U3655 , P1_U3657 );
nand NAND4_685 ( P1_U3381 , P1_U4314 , P1_U4313 , P1_U3659 , P1_U3661 );
nand NAND4_686 ( P1_U3382 , P1_U4333 , P1_U4332 , P1_U3663 , P1_U3665 );
nand NAND4_687 ( P1_U3383 , P1_U4352 , P1_U4351 , P1_U3667 , P1_U3669 );
nand NAND4_688 ( P1_U3384 , P1_U4371 , P1_U4370 , P1_U3671 , P1_U3673 );
nand NAND4_689 ( P1_U3385 , P1_U4390 , P1_U4389 , P1_U3675 , P1_U3677 );
nand NAND4_690 ( P1_U3386 , P1_U4409 , P1_U4408 , P1_U3679 , P1_U3681 );
nand NAND4_691 ( P1_U3387 , P1_U4428 , P1_U4427 , P1_U3683 , P1_U3685 );
nand NAND4_692 ( P1_U3388 , P1_U4447 , P1_U4446 , P1_U3687 , P1_U3689 );
nand NAND4_693 ( P1_U3389 , P1_U4466 , P1_U4465 , P1_U3691 , P1_U3693 );
nand NAND4_694 ( P1_U3390 , P1_U4485 , P1_U4484 , P1_U3695 , P1_U3697 );
nand NAND4_695 ( P1_U3391 , P1_U4504 , P1_U4503 , P1_U3699 , P1_U3701 );
nand NAND4_696 ( P1_U3392 , P1_U4523 , P1_U4522 , P1_U3703 , P1_U3705 );
nand NAND4_697 ( P1_U3393 , P1_U4542 , P1_U4541 , P1_U3707 , P1_U3709 );
nand NAND2_698 ( P1_U3394 , U76 , P1_U3946 );
nand NAND4_699 ( P1_U3395 , P1_U4561 , P1_U4560 , P1_U3711 , P1_U3713 );
nand NAND2_700 ( P1_U3396 , U75 , P1_U3946 );
nand NAND4_701 ( P1_U3397 , P1_U4580 , P1_U4579 , P1_U3715 , P1_U3717 );
nand NAND2_702 ( P1_U3398 , U74 , P1_U3946 );
nand NAND4_703 ( P1_U3399 , P1_U4599 , P1_U4598 , P1_U3719 , P1_U3721 );
nand NAND2_704 ( P1_U3400 , U73 , P1_U3946 );
nand NAND4_705 ( P1_U3401 , P1_U4618 , P1_U4617 , P1_U3723 , P1_U3725 );
nand NAND2_706 ( P1_U3402 , U72 , P1_U3946 );
nand NAND4_707 ( P1_U3403 , P1_U4637 , P1_U4636 , P1_U3727 , P1_U3729 );
nand NAND2_708 ( P1_U3404 , U71 , P1_U3946 );
nand NAND4_709 ( P1_U3405 , P1_U4656 , P1_U4655 , P1_U3731 , P1_U3733 );
nand NAND2_710 ( P1_U3406 , U70 , P1_U3946 );
nand NAND4_711 ( P1_U3407 , P1_U4675 , P1_U4674 , P1_U3735 , P1_U3737 );
nand NAND2_712 ( P1_U3408 , U69 , P1_U3946 );
nand NAND4_713 ( P1_U3409 , P1_U4694 , P1_U4693 , P1_U3739 , P1_U3741 );
nand NAND2_714 ( P1_U3410 , U68 , P1_U3946 );
nand NAND4_715 ( P1_U3411 , P1_U4713 , P1_U4712 , P1_U3743 , P1_U3745 );
nand NAND2_716 ( P1_U3412 , U67 , P1_U3946 );
nand NAND2_717 ( P1_U3413 , P1_U3750 , P1_U3748 );
nand NAND2_718 ( P1_U3414 , U65 , P1_U3946 );
nand NAND2_719 ( P1_U3415 , U64 , P1_U3946 );
nand NAND2_720 ( P1_U3416 , P1_U3986 , P1_U5719 );
nand NAND2_721 ( P1_U3417 , P1_U3022 , P1_U4757 );
nand NAND2_722 ( P1_U3418 , P1_U4021 , P1_U5716 );
nand NAND2_723 ( P1_U3419 , P1_U3048 , P1_U3448 );
nand NAND2_724 ( P1_U3420 , P1_U3023 , P1_U5713 );
nand NAND2_725 ( P1_U3421 , P1_U3050 , P1_U3437 );
nand NAND2_726 ( P1_U3422 , P1_U3999 , P1_U4758 );
nand NAND2_727 ( P1_U3423 , P1_U3424 , P1_U4921 );
nand NAND2_728 ( P1_U3424 , P1_U4135 , P1_U5703 );
nand NAND2_729 ( P1_U3425 , P1_U4032 , P1_STATE_REG );
nand NAND2_730 ( P1_U3426 , P1_U3444 , P1_U3439 );
nand NAND2_731 ( P1_U3427 , P1_U3014 , P1_U3015 );
nand NAND2_732 ( P1_U3428 , P1_U3439 , P1_U5713 );
not NOT1_733 ( P1_U3429 , P1_R1375_U14 );
nand NAND2_734 ( P1_U3430 , P1_U3022 , P1_U3422 );
nand NAND2_735 ( P1_U3431 , P1_U3876 , P1_U3016 );
nand NAND2_736 ( P1_U3432 , P1_U3014 , P1_U3022 );
nand NAND2_737 ( P1_U3433 , P1_U3879 , P1_U5133 );
nand NAND2_738 ( P1_U3434 , P1_U3443 , P1_U5719 );
nand NAND2_739 ( P1_U3435 , P1_U5403 , P1_U5402 );
nand NAND2_740 ( P1_U3436 , P1_U5691 , P1_U5690 );
nand NAND2_741 ( P1_U3437 , P1_U5694 , P1_U5693 );
nand NAND2_742 ( P1_U3438 , P1_U5697 , P1_U5696 );
nand NAND2_743 ( P1_U3439 , P1_U5702 , P1_U5701 );
nand NAND2_744 ( P1_U3440 , P1_U5705 , P1_U5704 );
nand NAND2_745 ( P1_U3441 , P1_U5707 , P1_U5706 );
nand NAND2_746 ( P1_U3442 , P1_U5715 , P1_U5714 );
nand NAND2_747 ( P1_U3443 , P1_U5712 , P1_U5711 );
nand NAND2_748 ( P1_U3444 , P1_U5709 , P1_U5708 );
nand NAND2_749 ( P1_U3445 , P1_U5721 , P1_U5720 );
nand NAND2_750 ( P1_U3446 , P1_U5724 , P1_U5723 );
nand NAND2_751 ( P1_U3447 , P1_U5727 , P1_U5726 );
nand NAND2_752 ( P1_U3448 , P1_U5718 , P1_U5717 );
nand NAND2_753 ( P1_U3449 , P1_U5730 , P1_U5729 );
nand NAND2_754 ( P1_U3450 , P1_U5733 , P1_U5732 );
nand NAND2_755 ( P1_U3451 , P1_U5736 , P1_U5735 );
nand NAND2_756 ( P1_U3452 , P1_U5744 , P1_U5743 );
nand NAND2_757 ( P1_U3453 , P1_U5741 , P1_U5740 );
nand NAND2_758 ( P1_U3454 , P1_U5747 , P1_U5746 );
nand NAND2_759 ( P1_U3455 , P1_U5749 , P1_U5748 );
nand NAND2_760 ( P1_U3456 , P1_U5751 , P1_U5750 );
nand NAND2_761 ( P1_U3457 , P1_U5754 , P1_U5753 );
nand NAND2_762 ( P1_U3458 , P1_U5756 , P1_U5755 );
nand NAND2_763 ( P1_U3459 , P1_U5758 , P1_U5757 );
nand NAND2_764 ( P1_U3460 , P1_U5761 , P1_U5760 );
nand NAND2_765 ( P1_U3461 , P1_U5763 , P1_U5762 );
nand NAND2_766 ( P1_U3462 , P1_U5765 , P1_U5764 );
nand NAND2_767 ( P1_U3463 , P1_U5768 , P1_U5767 );
nand NAND2_768 ( P1_U3464 , P1_U5770 , P1_U5769 );
nand NAND2_769 ( P1_U3465 , P1_U5772 , P1_U5771 );
nand NAND2_770 ( P1_U3466 , P1_U5775 , P1_U5774 );
nand NAND2_771 ( P1_U3467 , P1_U5777 , P1_U5776 );
nand NAND2_772 ( P1_U3468 , P1_U5779 , P1_U5778 );
nand NAND2_773 ( P1_U3469 , P1_U5782 , P1_U5781 );
nand NAND2_774 ( P1_U3470 , P1_U5784 , P1_U5783 );
nand NAND2_775 ( P1_U3471 , P1_U5786 , P1_U5785 );
nand NAND2_776 ( P1_U3472 , P1_U5789 , P1_U5788 );
nand NAND2_777 ( P1_U3473 , P1_U5791 , P1_U5790 );
nand NAND2_778 ( P1_U3474 , P1_U5793 , P1_U5792 );
nand NAND2_779 ( P1_U3475 , P1_U5796 , P1_U5795 );
nand NAND2_780 ( P1_U3476 , P1_U5798 , P1_U5797 );
nand NAND2_781 ( P1_U3477 , P1_U5800 , P1_U5799 );
nand NAND2_782 ( P1_U3478 , P1_U5803 , P1_U5802 );
nand NAND2_783 ( P1_U3479 , P1_U5805 , P1_U5804 );
nand NAND2_784 ( P1_U3480 , P1_U5807 , P1_U5806 );
nand NAND2_785 ( P1_U3481 , P1_U5810 , P1_U5809 );
nand NAND2_786 ( P1_U3482 , P1_U5812 , P1_U5811 );
nand NAND2_787 ( P1_U3483 , P1_U5814 , P1_U5813 );
nand NAND2_788 ( P1_U3484 , P1_U5817 , P1_U5816 );
nand NAND2_789 ( P1_U3485 , P1_U5819 , P1_U5818 );
nand NAND2_790 ( P1_U3486 , P1_U5821 , P1_U5820 );
nand NAND2_791 ( P1_U3487 , P1_U5824 , P1_U5823 );
nand NAND2_792 ( P1_U3488 , P1_U5826 , P1_U5825 );
nand NAND2_793 ( P1_U3489 , P1_U5828 , P1_U5827 );
nand NAND2_794 ( P1_U3490 , P1_U5831 , P1_U5830 );
nand NAND2_795 ( P1_U3491 , P1_U5833 , P1_U5832 );
nand NAND2_796 ( P1_U3492 , P1_U5835 , P1_U5834 );
nand NAND2_797 ( P1_U3493 , P1_U5838 , P1_U5837 );
nand NAND2_798 ( P1_U3494 , P1_U5840 , P1_U5839 );
nand NAND2_799 ( P1_U3495 , P1_U5842 , P1_U5841 );
nand NAND2_800 ( P1_U3496 , P1_U5845 , P1_U5844 );
nand NAND2_801 ( P1_U3497 , P1_U5847 , P1_U5846 );
nand NAND2_802 ( P1_U3498 , P1_U5849 , P1_U5848 );
nand NAND2_803 ( P1_U3499 , P1_U5852 , P1_U5851 );
nand NAND2_804 ( P1_U3500 , P1_U5854 , P1_U5853 );
nand NAND2_805 ( P1_U3501 , P1_U5856 , P1_U5855 );
nand NAND2_806 ( P1_U3502 , P1_U5859 , P1_U5858 );
nand NAND2_807 ( P1_U3503 , P1_U5861 , P1_U5860 );
nand NAND2_808 ( P1_U3504 , P1_U5863 , P1_U5862 );
nand NAND2_809 ( P1_U3505 , P1_U5866 , P1_U5865 );
nand NAND2_810 ( P1_U3506 , P1_U5868 , P1_U5867 );
nand NAND2_811 ( P1_U3507 , P1_U5870 , P1_U5869 );
nand NAND2_812 ( P1_U3508 , P1_U5873 , P1_U5872 );
nand NAND2_813 ( P1_U3509 , P1_U5875 , P1_U5874 );
nand NAND2_814 ( P1_U3510 , P1_U5878 , P1_U5877 );
nand NAND2_815 ( P1_U3511 , P1_U5880 , P1_U5879 );
nand NAND2_816 ( P1_U3512 , P1_U5882 , P1_U5881 );
nand NAND2_817 ( P1_U3513 , P1_U5884 , P1_U5883 );
nand NAND2_818 ( P1_U3514 , P1_U5886 , P1_U5885 );
nand NAND2_819 ( P1_U3515 , P1_U5888 , P1_U5887 );
nand NAND2_820 ( P1_U3516 , P1_U5890 , P1_U5889 );
nand NAND2_821 ( P1_U3517 , P1_U5892 , P1_U5891 );
nand NAND2_822 ( P1_U3518 , P1_U5894 , P1_U5893 );
nand NAND2_823 ( P1_U3519 , P1_U5896 , P1_U5895 );
nand NAND2_824 ( P1_U3520 , P1_U5898 , P1_U5897 );
nand NAND2_825 ( P1_U3521 , P1_U5900 , P1_U5899 );
nand NAND2_826 ( P1_U3522 , P1_U5902 , P1_U5901 );
nand NAND2_827 ( P1_U3523 , P1_U5904 , P1_U5903 );
nand NAND2_828 ( P1_U3524 , P1_U5906 , P1_U5905 );
nand NAND2_829 ( P1_U3525 , P1_U5908 , P1_U5907 );
nand NAND2_830 ( P1_U3526 , P1_U5910 , P1_U5909 );
nand NAND2_831 ( P1_U3527 , P1_U5912 , P1_U5911 );
nand NAND2_832 ( P1_U3528 , P1_U5914 , P1_U5913 );
nand NAND2_833 ( P1_U3529 , P1_U5916 , P1_U5915 );
nand NAND2_834 ( P1_U3530 , P1_U5918 , P1_U5917 );
nand NAND2_835 ( P1_U3531 , P1_U5920 , P1_U5919 );
nand NAND2_836 ( P1_U3532 , P1_U5922 , P1_U5921 );
nand NAND2_837 ( P1_U3533 , P1_U5924 , P1_U5923 );
nand NAND2_838 ( P1_U3534 , P1_U5926 , P1_U5925 );
nand NAND2_839 ( P1_U3535 , P1_U5928 , P1_U5927 );
nand NAND2_840 ( P1_U3536 , P1_U5930 , P1_U5929 );
nand NAND2_841 ( P1_U3537 , P1_U5932 , P1_U5931 );
nand NAND2_842 ( P1_U3538 , P1_U5934 , P1_U5933 );
nand NAND2_843 ( P1_U3539 , P1_U5936 , P1_U5935 );
nand NAND2_844 ( P1_U3540 , P1_U5938 , P1_U5937 );
nand NAND2_845 ( P1_U3541 , P1_U5940 , P1_U5939 );
nand NAND2_846 ( P1_U3542 , P1_U5942 , P1_U5941 );
nand NAND2_847 ( P1_U3543 , P1_U5944 , P1_U5943 );
nand NAND2_848 ( P1_U3544 , P1_U5946 , P1_U5945 );
nand NAND2_849 ( P1_U3545 , P1_U5948 , P1_U5947 );
nand NAND2_850 ( P1_U3546 , P1_U5950 , P1_U5949 );
nand NAND2_851 ( P1_U3547 , P1_U5952 , P1_U5951 );
nand NAND2_852 ( P1_U3548 , P1_U5954 , P1_U5953 );
nand NAND2_853 ( P1_U3549 , P1_U5956 , P1_U5955 );
nand NAND2_854 ( P1_U3550 , P1_U5958 , P1_U5957 );
nand NAND2_855 ( P1_U3551 , P1_U5960 , P1_U5959 );
nand NAND2_856 ( P1_U3552 , P1_U5962 , P1_U5961 );
nand NAND2_857 ( P1_U3553 , P1_U5964 , P1_U5963 );
nand NAND2_858 ( P1_U3554 , P1_U5966 , P1_U5965 );
nand NAND2_859 ( P1_U3555 , P1_U6032 , P1_U6031 );
nand NAND2_860 ( P1_U3556 , P1_U6034 , P1_U6033 );
nand NAND2_861 ( P1_U3557 , P1_U6036 , P1_U6035 );
nand NAND2_862 ( P1_U3558 , P1_U6038 , P1_U6037 );
nand NAND2_863 ( P1_U3559 , P1_U6040 , P1_U6039 );
nand NAND2_864 ( P1_U3560 , P1_U6042 , P1_U6041 );
nand NAND2_865 ( P1_U3561 , P1_U6044 , P1_U6043 );
nand NAND2_866 ( P1_U3562 , P1_U6046 , P1_U6045 );
nand NAND2_867 ( P1_U3563 , P1_U6048 , P1_U6047 );
nand NAND2_868 ( P1_U3564 , P1_U6050 , P1_U6049 );
nand NAND2_869 ( P1_U3565 , P1_U6052 , P1_U6051 );
nand NAND2_870 ( P1_U3566 , P1_U6054 , P1_U6053 );
nand NAND2_871 ( P1_U3567 , P1_U6056 , P1_U6055 );
nand NAND2_872 ( P1_U3568 , P1_U6058 , P1_U6057 );
nand NAND2_873 ( P1_U3569 , P1_U6060 , P1_U6059 );
nand NAND2_874 ( P1_U3570 , P1_U6062 , P1_U6061 );
nand NAND2_875 ( P1_U3571 , P1_U6064 , P1_U6063 );
nand NAND2_876 ( P1_U3572 , P1_U6066 , P1_U6065 );
nand NAND2_877 ( P1_U3573 , P1_U6068 , P1_U6067 );
nand NAND2_878 ( P1_U3574 , P1_U6070 , P1_U6069 );
nand NAND2_879 ( P1_U3575 , P1_U6072 , P1_U6071 );
nand NAND2_880 ( P1_U3576 , P1_U6074 , P1_U6073 );
nand NAND2_881 ( P1_U3577 , P1_U6076 , P1_U6075 );
nand NAND2_882 ( P1_U3578 , P1_U6078 , P1_U6077 );
nand NAND2_883 ( P1_U3579 , P1_U6080 , P1_U6079 );
nand NAND2_884 ( P1_U3580 , P1_U6082 , P1_U6081 );
nand NAND2_885 ( P1_U3581 , P1_U6084 , P1_U6083 );
nand NAND2_886 ( P1_U3582 , P1_U6086 , P1_U6085 );
nand NAND2_887 ( P1_U3583 , P1_U6088 , P1_U6087 );
nand NAND2_888 ( P1_U3584 , P1_U6090 , P1_U6089 );
nand NAND2_889 ( P1_U3585 , P1_U6092 , P1_U6091 );
nand NAND2_890 ( P1_U3586 , P1_U6094 , P1_U6093 );
nand NAND2_891 ( P1_U3587 , P1_U6202 , P1_U6201 );
nand NAND2_892 ( P1_U3588 , P1_U6204 , P1_U6203 );
nand NAND2_893 ( P1_U3589 , P1_U6206 , P1_U6205 );
nand NAND2_894 ( P1_U3590 , P1_U6208 , P1_U6207 );
nand NAND2_895 ( P1_U3591 , P1_U6210 , P1_U6209 );
nand NAND2_896 ( P1_U3592 , P1_U6212 , P1_U6211 );
nand NAND2_897 ( P1_U3593 , P1_U6214 , P1_U6213 );
nand NAND2_898 ( P1_U3594 , P1_U6216 , P1_U6215 );
nand NAND2_899 ( P1_U3595 , P1_U6218 , P1_U6217 );
nand NAND2_900 ( P1_U3596 , P1_U6220 , P1_U6219 );
nand NAND2_901 ( P1_U3597 , P1_U6222 , P1_U6221 );
nand NAND2_902 ( P1_U3598 , P1_U6224 , P1_U6223 );
nand NAND2_903 ( P1_U3599 , P1_U6226 , P1_U6225 );
nand NAND2_904 ( P1_U3600 , P1_U6228 , P1_U6227 );
nand NAND2_905 ( P1_U3601 , P1_U6230 , P1_U6229 );
nand NAND2_906 ( P1_U3602 , P1_U6232 , P1_U6231 );
nand NAND2_907 ( P1_U3603 , P1_U6234 , P1_U6233 );
nand NAND2_908 ( P1_U3604 , P1_U6236 , P1_U6235 );
nand NAND2_909 ( P1_U3605 , P1_U6238 , P1_U6237 );
nand NAND2_910 ( P1_U3606 , P1_U6240 , P1_U6239 );
nand NAND2_911 ( P1_U3607 , P1_U6242 , P1_U6241 );
nand NAND2_912 ( P1_U3608 , P1_U6244 , P1_U6243 );
nand NAND2_913 ( P1_U3609 , P1_U6246 , P1_U6245 );
nand NAND2_914 ( P1_U3610 , P1_U6248 , P1_U6247 );
nand NAND2_915 ( P1_U3611 , P1_U6250 , P1_U6249 );
nand NAND2_916 ( P1_U3612 , P1_U6252 , P1_U6251 );
nand NAND2_917 ( P1_U3613 , P1_U6254 , P1_U6253 );
nand NAND2_918 ( P1_U3614 , P1_U6256 , P1_U6255 );
nand NAND2_919 ( P1_U3615 , P1_U6258 , P1_U6257 );
nand NAND2_920 ( P1_U3616 , P1_U6260 , P1_U6259 );
nand NAND2_921 ( P1_U3617 , P1_U6262 , P1_U6261 );
nand NAND2_922 ( P1_U3618 , P1_U6264 , P1_U6263 );
and AND2_923 ( P1_U3619 , P1_U4177 , P1_U4176 );
and AND2_924 ( P1_U3620 , P1_U4179 , P1_U4178 );
and AND2_925 ( P1_U3621 , P1_U4186 , P1_U4184 );
and AND3_926 ( P1_U3622 , P1_U4187 , P1_U4185 , P1_U3621 );
and AND4_927 ( P1_U3623 , P1_U4141 , P1_U4140 , P1_U4139 , P1_U4138 );
and AND4_928 ( P1_U3624 , P1_U4145 , P1_U4144 , P1_U4143 , P1_U4142 );
and AND4_929 ( P1_U3625 , P1_U4149 , P1_U4148 , P1_U4147 , P1_U4146 );
and AND3_930 ( P1_U3626 , P1_U4151 , P1_U4150 , P1_U4152 );
and AND4_931 ( P1_U3627 , P1_U3626 , P1_U3625 , P1_U3624 , P1_U3623 );
and AND4_932 ( P1_U3628 , P1_U4156 , P1_U4155 , P1_U4154 , P1_U4153 );
and AND4_933 ( P1_U3629 , P1_U4160 , P1_U4159 , P1_U4158 , P1_U4157 );
and AND4_934 ( P1_U3630 , P1_U4164 , P1_U4163 , P1_U4162 , P1_U4161 );
and AND3_935 ( P1_U3631 , P1_U4166 , P1_U4165 , P1_U4167 );
and AND4_936 ( P1_U3632 , P1_U3631 , P1_U3630 , P1_U3629 , P1_U3628 );
and AND2_937 ( P1_U3633 , P1_U5742 , P1_U4169 );
and AND2_938 ( P1_U3634 , P1_U5745 , P1_U3022 );
and AND2_939 ( P1_U3635 , P1_U4202 , P1_U4201 );
and AND2_940 ( P1_U3636 , P1_U4204 , P1_U4203 );
and AND3_941 ( P1_U3637 , P1_U4206 , P1_U4205 , P1_U3636 );
and AND4_942 ( P1_U3638 , P1_U4209 , P1_U4210 , P1_U4211 , P1_U4208 );
and AND2_943 ( P1_U3639 , P1_U4221 , P1_U4220 );
and AND2_944 ( P1_U3640 , P1_U4223 , P1_U4222 );
and AND3_945 ( P1_U3641 , P1_U4225 , P1_U4224 , P1_U3640 );
and AND4_946 ( P1_U3642 , P1_U4228 , P1_U4229 , P1_U4230 , P1_U4227 );
and AND2_947 ( P1_U3643 , P1_U4240 , P1_U4239 );
and AND2_948 ( P1_U3644 , P1_U4242 , P1_U4241 );
and AND3_949 ( P1_U3645 , P1_U4244 , P1_U4243 , P1_U3644 );
and AND4_950 ( P1_U3646 , P1_U4247 , P1_U4248 , P1_U4249 , P1_U4246 );
and AND2_951 ( P1_U3647 , P1_U4259 , P1_U4258 );
and AND2_952 ( P1_U3648 , P1_U4261 , P1_U4260 );
and AND3_953 ( P1_U3649 , P1_U4263 , P1_U4262 , P1_U3648 );
and AND4_954 ( P1_U3650 , P1_U4266 , P1_U4267 , P1_U4268 , P1_U4265 );
and AND2_955 ( P1_U3651 , P1_U4278 , P1_U4277 );
and AND2_956 ( P1_U3652 , P1_U4280 , P1_U4279 );
and AND3_957 ( P1_U3653 , P1_U4282 , P1_U4281 , P1_U3652 );
and AND4_958 ( P1_U3654 , P1_U4285 , P1_U4286 , P1_U4287 , P1_U4284 );
and AND2_959 ( P1_U3655 , P1_U4297 , P1_U4296 );
and AND2_960 ( P1_U3656 , P1_U4299 , P1_U4298 );
and AND3_961 ( P1_U3657 , P1_U4301 , P1_U4300 , P1_U3656 );
and AND4_962 ( P1_U3658 , P1_U4304 , P1_U4305 , P1_U4306 , P1_U4303 );
and AND2_963 ( P1_U3659 , P1_U4316 , P1_U4315 );
and AND2_964 ( P1_U3660 , P1_U4318 , P1_U4317 );
and AND3_965 ( P1_U3661 , P1_U4320 , P1_U4319 , P1_U3660 );
and AND4_966 ( P1_U3662 , P1_U4323 , P1_U4324 , P1_U4325 , P1_U4322 );
and AND2_967 ( P1_U3663 , P1_U4335 , P1_U4334 );
and AND2_968 ( P1_U3664 , P1_U4337 , P1_U4336 );
and AND3_969 ( P1_U3665 , P1_U4339 , P1_U4338 , P1_U3664 );
and AND4_970 ( P1_U3666 , P1_U4342 , P1_U4343 , P1_U4344 , P1_U4341 );
and AND2_971 ( P1_U3667 , P1_U4354 , P1_U4353 );
and AND2_972 ( P1_U3668 , P1_U4356 , P1_U4355 );
and AND3_973 ( P1_U3669 , P1_U4358 , P1_U4357 , P1_U3668 );
and AND4_974 ( P1_U3670 , P1_U4361 , P1_U4362 , P1_U4363 , P1_U4360 );
and AND2_975 ( P1_U3671 , P1_U4373 , P1_U4372 );
and AND2_976 ( P1_U3672 , P1_U4375 , P1_U4374 );
and AND3_977 ( P1_U3673 , P1_U4377 , P1_U4376 , P1_U3672 );
and AND4_978 ( P1_U3674 , P1_U4380 , P1_U4381 , P1_U4382 , P1_U4379 );
and AND2_979 ( P1_U3675 , P1_U4392 , P1_U4391 );
and AND2_980 ( P1_U3676 , P1_U4394 , P1_U4393 );
and AND3_981 ( P1_U3677 , P1_U4396 , P1_U4395 , P1_U3676 );
and AND4_982 ( P1_U3678 , P1_U4401 , P1_U4400 , P1_U4399 , P1_U4398 );
and AND2_983 ( P1_U3679 , P1_U4411 , P1_U4410 );
and AND2_984 ( P1_U3680 , P1_U4413 , P1_U4412 );
and AND3_985 ( P1_U3681 , P1_U4415 , P1_U4414 , P1_U3680 );
and AND4_986 ( P1_U3682 , P1_U4420 , P1_U4419 , P1_U4418 , P1_U4417 );
and AND2_987 ( P1_U3683 , P1_U4430 , P1_U4429 );
and AND2_988 ( P1_U3684 , P1_U4432 , P1_U4431 );
and AND3_989 ( P1_U3685 , P1_U4434 , P1_U4433 , P1_U3684 );
and AND4_990 ( P1_U3686 , P1_U4439 , P1_U4438 , P1_U4437 , P1_U4436 );
and AND2_991 ( P1_U3687 , P1_U4449 , P1_U4448 );
and AND2_992 ( P1_U3688 , P1_U4451 , P1_U4450 );
and AND3_993 ( P1_U3689 , P1_U4453 , P1_U4452 , P1_U3688 );
and AND4_994 ( P1_U3690 , P1_U4458 , P1_U4455 , P1_U4456 , P1_U4457 );
and AND2_995 ( P1_U3691 , P1_U4468 , P1_U4467 );
and AND2_996 ( P1_U3692 , P1_U4470 , P1_U4469 );
and AND3_997 ( P1_U3693 , P1_U4472 , P1_U4471 , P1_U3692 );
and AND4_998 ( P1_U3694 , P1_U4475 , P1_U4476 , P1_U4477 , P1_U4474 );
and AND2_999 ( P1_U3695 , P1_U4487 , P1_U4486 );
and AND2_1000 ( P1_U3696 , P1_U4489 , P1_U4488 );
and AND3_1001 ( P1_U3697 , P1_U4491 , P1_U4490 , P1_U3696 );
and AND4_1002 ( P1_U3698 , P1_U4494 , P1_U4495 , P1_U4496 , P1_U4493 );
and AND2_1003 ( P1_U3699 , P1_U4506 , P1_U4505 );
and AND2_1004 ( P1_U3700 , P1_U4508 , P1_U4507 );
and AND3_1005 ( P1_U3701 , P1_U4510 , P1_U4509 , P1_U3700 );
and AND4_1006 ( P1_U3702 , P1_U4515 , P1_U4512 , P1_U4513 , P1_U4514 );
and AND2_1007 ( P1_U3703 , P1_U4525 , P1_U4524 );
and AND2_1008 ( P1_U3704 , P1_U4527 , P1_U4526 );
and AND3_1009 ( P1_U3705 , P1_U4529 , P1_U4528 , P1_U3704 );
and AND4_1010 ( P1_U3706 , P1_U4534 , P1_U4531 , P1_U4532 , P1_U4533 );
and AND2_1011 ( P1_U3707 , P1_U4544 , P1_U4543 );
and AND2_1012 ( P1_U3708 , P1_U4546 , P1_U4545 );
and AND3_1013 ( P1_U3709 , P1_U4548 , P1_U4547 , P1_U3708 );
and AND4_1014 ( P1_U3710 , P1_U4551 , P1_U4552 , P1_U4553 , P1_U4550 );
and AND2_1015 ( P1_U3711 , P1_U4563 , P1_U4562 );
and AND2_1016 ( P1_U3712 , P1_U4565 , P1_U4564 );
and AND3_1017 ( P1_U3713 , P1_U4567 , P1_U4566 , P1_U3712 );
and AND4_1018 ( P1_U3714 , P1_U4570 , P1_U4571 , P1_U4572 , P1_U4569 );
and AND2_1019 ( P1_U3715 , P1_U4582 , P1_U4581 );
and AND2_1020 ( P1_U3716 , P1_U4584 , P1_U4583 );
and AND3_1021 ( P1_U3717 , P1_U4586 , P1_U4585 , P1_U3716 );
and AND4_1022 ( P1_U3718 , P1_U4589 , P1_U4590 , P1_U4591 , P1_U4588 );
and AND2_1023 ( P1_U3719 , P1_U4601 , P1_U4600 );
and AND2_1024 ( P1_U3720 , P1_U4603 , P1_U4602 );
and AND3_1025 ( P1_U3721 , P1_U4605 , P1_U4604 , P1_U3720 );
and AND4_1026 ( P1_U3722 , P1_U4608 , P1_U4609 , P1_U4610 , P1_U4607 );
and AND2_1027 ( P1_U3723 , P1_U4620 , P1_U4619 );
and AND2_1028 ( P1_U3724 , P1_U4622 , P1_U4621 );
and AND3_1029 ( P1_U3725 , P1_U4624 , P1_U4623 , P1_U3724 );
and AND4_1030 ( P1_U3726 , P1_U4627 , P1_U4628 , P1_U4629 , P1_U4626 );
and AND2_1031 ( P1_U3727 , P1_U4639 , P1_U4638 );
and AND2_1032 ( P1_U3728 , P1_U4641 , P1_U4640 );
and AND3_1033 ( P1_U3729 , P1_U4643 , P1_U4642 , P1_U3728 );
and AND4_1034 ( P1_U3730 , P1_U4646 , P1_U4647 , P1_U4648 , P1_U4645 );
and AND2_1035 ( P1_U3731 , P1_U4658 , P1_U4657 );
and AND2_1036 ( P1_U3732 , P1_U4660 , P1_U4659 );
and AND3_1037 ( P1_U3733 , P1_U4662 , P1_U4661 , P1_U3732 );
and AND4_1038 ( P1_U3734 , P1_U4665 , P1_U4666 , P1_U4667 , P1_U4664 );
and AND2_1039 ( P1_U3735 , P1_U4677 , P1_U4676 );
and AND2_1040 ( P1_U3736 , P1_U4679 , P1_U4678 );
and AND3_1041 ( P1_U3737 , P1_U4681 , P1_U4680 , P1_U3736 );
and AND4_1042 ( P1_U3738 , P1_U4684 , P1_U4685 , P1_U4686 , P1_U4683 );
and AND2_1043 ( P1_U3739 , P1_U4696 , P1_U4695 );
and AND2_1044 ( P1_U3740 , P1_U4698 , P1_U4697 );
and AND3_1045 ( P1_U3741 , P1_U4700 , P1_U4699 , P1_U3740 );
and AND4_1046 ( P1_U3742 , P1_U4703 , P1_U4704 , P1_U4705 , P1_U4702 );
and AND2_1047 ( P1_U3743 , P1_U4715 , P1_U4714 );
and AND2_1048 ( P1_U3744 , P1_U4717 , P1_U4716 );
and AND3_1049 ( P1_U3745 , P1_U4719 , P1_U4718 , P1_U3744 );
and AND4_1050 ( P1_U3746 , P1_U4722 , P1_U4723 , P1_U4724 , P1_U4721 );
and AND2_1051 ( P1_U3747 , P1_U4731 , P1_U4020 );
and AND5_1052 ( P1_U3748 , P1_U4733 , P1_U4732 , P1_U4734 , P1_U4735 , P1_U4736 );
and AND2_1053 ( P1_U3749 , P1_U4738 , P1_U4737 );
and AND3_1054 ( P1_U3750 , P1_U4740 , P1_U4739 , P1_U3749 );
and AND3_1055 ( P1_U3751 , P1_U4743 , P1_U4744 , P1_U4742 );
and AND2_1056 ( P1_U3752 , P1_U4020 , P1_U4731 );
and AND2_1057 ( P1_U3753 , P1_U3022 , P1_U3452 );
and AND3_1058 ( P1_U3754 , P1_U5745 , P1_U4002 , P1_U3453 );
and AND3_1059 ( P1_U3755 , P1_U4761 , P1_U4760 , P1_U4762 );
and AND3_1060 ( P1_U3756 , P1_U4764 , P1_U4763 , P1_U3949 );
and AND3_1061 ( P1_U3757 , P1_U4766 , P1_U4765 , P1_U4767 );
and AND3_1062 ( P1_U3758 , P1_U4769 , P1_U4768 , P1_U3950 );
and AND3_1063 ( P1_U3759 , P1_U4771 , P1_U4770 , P1_U4772 );
and AND3_1064 ( P1_U3760 , P1_U4774 , P1_U4773 , P1_U3951 );
and AND3_1065 ( P1_U3761 , P1_U4776 , P1_U4775 , P1_U4777 );
and AND3_1066 ( P1_U3762 , P1_U4779 , P1_U4778 , P1_U3952 );
and AND3_1067 ( P1_U3763 , P1_U4781 , P1_U4780 , P1_U4782 );
and AND3_1068 ( P1_U3764 , P1_U4784 , P1_U4783 , P1_U3953 );
and AND3_1069 ( P1_U3765 , P1_U4786 , P1_U4785 , P1_U4787 );
and AND2_1070 ( P1_U3766 , P1_U4789 , P1_U4788 );
and AND3_1071 ( P1_U3767 , P1_U4791 , P1_U4790 , P1_U4792 );
and AND2_1072 ( P1_U3768 , P1_U4794 , P1_U4793 );
and AND3_1073 ( P1_U3769 , P1_U4796 , P1_U4795 , P1_U4797 );
and AND2_1074 ( P1_U3770 , P1_U4799 , P1_U4798 );
and AND3_1075 ( P1_U3771 , P1_U4801 , P1_U4800 , P1_U4802 );
and AND2_1076 ( P1_U3772 , P1_U4804 , P1_U4803 );
and AND2_1077 ( P1_U3773 , P1_U4806 , P1_U4805 );
and AND2_1078 ( P1_U3774 , P1_U4809 , P1_U4808 );
and AND2_1079 ( P1_U3775 , P1_U4811 , P1_U4810 );
and AND2_1080 ( P1_U3776 , P1_U4814 , P1_U4813 );
and AND3_1081 ( P1_U3777 , P1_U4816 , P1_U4815 , P1_U4817 );
and AND2_1082 ( P1_U3778 , P1_U4819 , P1_U4818 );
and AND3_1083 ( P1_U3779 , P1_U4821 , P1_U4820 , P1_U4822 );
and AND2_1084 ( P1_U3780 , P1_U4824 , P1_U4823 );
and AND3_1085 ( P1_U3781 , P1_U4826 , P1_U4825 , P1_U4827 );
and AND2_1086 ( P1_U3782 , P1_U4829 , P1_U4828 );
and AND3_1087 ( P1_U3783 , P1_U4831 , P1_U4830 , P1_U4832 );
and AND2_1088 ( P1_U3784 , P1_U4834 , P1_U4833 );
and AND2_1089 ( P1_U3785 , P1_U4836 , P1_U4835 );
and AND2_1090 ( P1_U3786 , P1_U4839 , P1_U4838 );
and AND2_1091 ( P1_U3787 , P1_U4841 , P1_U4840 );
and AND2_1092 ( P1_U3788 , P1_U4844 , P1_U4843 );
and AND3_1093 ( P1_U3789 , P1_U4846 , P1_U4845 , P1_U4847 );
and AND2_1094 ( P1_U3790 , P1_U4849 , P1_U4848 );
and AND3_1095 ( P1_U3791 , P1_U4851 , P1_U4850 , P1_U4852 );
and AND2_1096 ( P1_U3792 , P1_U4854 , P1_U4853 );
and AND2_1097 ( P1_U3793 , P1_U4856 , P1_U4855 );
and AND2_1098 ( P1_U3794 , P1_U4859 , P1_U4858 );
and AND2_1099 ( P1_U3795 , P1_U4861 , P1_U4860 );
and AND2_1100 ( P1_U3796 , P1_U4864 , P1_U4863 );
and AND2_1101 ( P1_U3797 , P1_U4866 , P1_U4865 );
and AND2_1102 ( P1_U3798 , P1_U4869 , P1_U4868 );
and AND2_1103 ( P1_U3799 , P1_U4871 , P1_U4870 );
and AND2_1104 ( P1_U3800 , P1_U4874 , P1_U4873 );
and AND2_1105 ( P1_U3801 , P1_U4876 , P1_U4875 );
and AND2_1106 ( P1_U3802 , P1_U4879 , P1_U4878 );
and AND2_1107 ( P1_U3803 , P1_U4881 , P1_U4880 );
and AND2_1108 ( P1_U3804 , P1_U4884 , P1_U4883 );
and AND2_1109 ( P1_U3805 , P1_U4886 , P1_U4885 );
and AND2_1110 ( P1_U3806 , P1_U4889 , P1_U4888 );
and AND2_1111 ( P1_U3807 , P1_U4891 , P1_U4890 );
and AND2_1112 ( P1_U3808 , P1_U4894 , P1_U4893 );
and AND2_1113 ( P1_U3809 , P1_U4896 , P1_U4895 );
and AND2_1114 ( P1_U3810 , P1_U4899 , P1_U4898 );
and AND2_1115 ( P1_U3811 , P1_U4901 , P1_U4900 );
and AND2_1116 ( P1_U3812 , P1_U4904 , P1_U4903 );
and AND3_1117 ( P1_U3813 , P1_U3419 , P1_U3369 , P1_U3365 );
and AND3_1118 ( P1_U3814 , P1_U3367 , P1_U3364 , P1_U3360 );
and AND2_1119 ( P1_U3815 , P1_U3361 , P1_U3363 );
and AND2_1120 ( P1_U3816 , P1_U3815 , P1_U3420 );
and AND2_1121 ( P1_U3817 , P1_U3439 , P1_STATE_REG );
and AND2_1122 ( P1_U3818 , P1_U4924 , P1_U4925 );
and AND3_1123 ( P1_U3819 , P1_U4928 , P1_U4926 , P1_U4927 );
and AND2_1124 ( P1_U3820 , P1_U4934 , P1_U4935 );
and AND3_1125 ( P1_U3821 , P1_U4938 , P1_U4936 , P1_U4937 );
and AND2_1126 ( P1_U3822 , P1_U4944 , P1_U4945 );
and AND3_1127 ( P1_U3823 , P1_U4948 , P1_U4946 , P1_U4947 );
and AND2_1128 ( P1_U3824 , P1_U4954 , P1_U4955 );
and AND3_1129 ( P1_U3825 , P1_U4958 , P1_U4956 , P1_U4957 );
and AND2_1130 ( P1_U3826 , P1_U4964 , P1_U4965 );
and AND3_1131 ( P1_U3827 , P1_U4968 , P1_U4966 , P1_U4967 );
and AND2_1132 ( P1_U3828 , P1_U4974 , P1_U4975 );
and AND3_1133 ( P1_U3829 , P1_U4978 , P1_U4976 , P1_U4977 );
and AND2_1134 ( P1_U3830 , P1_U4984 , P1_U4985 );
and AND3_1135 ( P1_U3831 , P1_U4988 , P1_U4986 , P1_U4987 );
and AND2_1136 ( P1_U3832 , P1_U4994 , P1_U4995 );
and AND3_1137 ( P1_U3833 , P1_U4998 , P1_U4996 , P1_U4997 );
and AND2_1138 ( P1_U3834 , P1_U5004 , P1_U5005 );
and AND3_1139 ( P1_U3835 , P1_U5008 , P1_U5006 , P1_U5007 );
and AND2_1140 ( P1_U3836 , P1_U5014 , P1_U5015 );
and AND3_1141 ( P1_U3837 , P1_U5018 , P1_U5016 , P1_U5017 );
and AND2_1142 ( P1_U3838 , P1_U5024 , P1_U5025 );
and AND3_1143 ( P1_U3839 , P1_U5028 , P1_U5026 , P1_U5027 );
and AND2_1144 ( P1_U3840 , P1_U5034 , P1_U5035 );
and AND3_1145 ( P1_U3841 , P1_U5038 , P1_U5036 , P1_U5037 );
and AND2_1146 ( P1_U3842 , P1_U5044 , P1_U5045 );
and AND3_1147 ( P1_U3843 , P1_U5047 , P1_U5046 , P1_U5048 );
and AND3_1148 ( P1_U3844 , P1_U5054 , P1_U5055 , P1_U5053 );
and AND3_1149 ( P1_U3845 , P1_U5057 , P1_U5056 , P1_U5058 );
and AND3_1150 ( P1_U3846 , P1_U5064 , P1_U5065 , P1_U5063 );
and AND3_1151 ( P1_U3847 , P1_U5067 , P1_U5066 , P1_U5068 );
and AND2_1152 ( P1_U3848 , P1_U5073 , P1_U4031 );
and AND3_1153 ( P1_U3849 , P1_U5075 , P1_U5074 , P1_U3848 );
and AND3_1154 ( P1_U3850 , P1_U5077 , P1_U5076 , P1_U5078 );
and AND3_1155 ( P1_U3851 , P1_U5084 , P1_U5085 , P1_U5083 );
and AND3_1156 ( P1_U3852 , P1_U5087 , P1_U5086 , P1_U5088 );
and AND2_1157 ( P1_U3853 , P1_U5093 , P1_U4031 );
and AND3_1158 ( P1_U3854 , P1_U5095 , P1_U5094 , P1_U3853 );
and AND3_1159 ( P1_U3855 , P1_U5097 , P1_U5096 , P1_U5098 );
and AND3_1160 ( P1_U3856 , P1_U5104 , P1_U5105 , P1_U5103 );
and AND3_1161 ( P1_U3857 , P1_U5107 , P1_U5106 , P1_U5108 );
and AND3_1162 ( P1_U3858 , P1_U5114 , P1_U5115 , P1_U5113 );
and AND3_1163 ( P1_U3859 , P1_U5117 , P1_U5116 , P1_U5118 );
and AND2_1164 ( P1_U3860 , P1_STATE_REG , P1_U3426 );
and AND2_1165 ( P1_U3861 , P1_U3860 , P1_U3424 );
and AND3_1166 ( P1_U3862 , P1_U6127 , P1_U6124 , P1_U6130 );
and AND3_1167 ( P1_U3863 , P1_U3864 , P1_U3862 , P1_U6142 );
and AND3_1168 ( P1_U3864 , P1_U6139 , P1_U6136 , P1_U6133 );
and AND3_1169 ( P1_U3865 , P1_U6151 , P1_U6148 , P1_U6154 );
and AND3_1170 ( P1_U3866 , P1_U6160 , P1_U6157 , P1_U6163 );
and AND3_1171 ( P1_U3867 , P1_U3866 , P1_U3865 , P1_U6145 );
and AND4_1172 ( P1_U3868 , P1_U3867 , P1_U3863 , P1_U6121 , P1_U6166 );
and AND2_1173 ( P1_U3869 , P1_U6190 , P1_U6187 );
and AND5_1174 ( P1_U3870 , P1_U6181 , P1_U6178 , P1_U6175 , P1_U6172 , P1_U6184 );
and AND2_1175 ( P1_U3871 , P1_U3870 , P1_U6169 );
and AND4_1176 ( P1_U3872 , P1_U6112 , P1_U6109 , P1_U6106 , P1_U6103 );
and AND2_1177 ( P1_U3873 , P1_U6118 , P1_U6115 );
and AND4_1178 ( P1_U3874 , P1_U3873 , P1_U3872 , P1_U6100 , P1_U6097 );
and AND4_1179 ( P1_U3875 , P1_U5689 , P1_U5123 , P1_U3984 , P1_U5687 );
and AND2_1180 ( P1_U3876 , P1_U3452 , P1_U3453 );
and AND3_1181 ( P1_U3877 , P1_U3370 , P1_U3368 , P1_U3420 );
and AND2_1182 ( P1_U3878 , P1_U5703 , P1_U4002 );
and AND2_1183 ( P1_U3879 , P1_U3424 , P1_U3878 );
and AND2_1184 ( P1_U3880 , P1_U3022 , P1_U5132 );
and AND2_1185 ( P1_U3881 , P1_U3882 , P1_U5175 );
and AND2_1186 ( P1_U3882 , P1_U5179 , P1_U5178 );
and AND2_1187 ( P1_U3883 , P1_U4027 , P1_U3076 );
and AND2_1188 ( P1_U3884 , P1_U5220 , P1_U5219 );
and AND2_1189 ( P1_U3885 , P1_U5223 , P1_U5222 );
and AND2_1190 ( P1_U3886 , P1_U3887 , P1_U5237 );
and AND2_1191 ( P1_U3887 , P1_U5241 , P1_U5240 );
and AND2_1192 ( P1_U3888 , P1_U5268 , P1_U5267 );
and AND2_1193 ( P1_U3889 , P1_U3890 , P1_U5309 );
and AND2_1194 ( P1_U3890 , P1_U5313 , P1_U5312 );
and AND2_1195 ( P1_U3891 , P1_U3892 , P1_U5345 );
and AND2_1196 ( P1_U3892 , P1_U5349 , P1_U5348 );
and AND2_1197 ( P1_U3893 , P1_U3434 , P1_U5398 );
and AND2_1198 ( P1_U3894 , P1_U5463 , P1_U5464 );
and AND2_1199 ( P1_U3895 , P1_U5523 , P1_U5521 );
and AND2_1200 ( P1_U3896 , P1_U3439 , P1_U5535 );
and AND2_1201 ( P1_U3897 , P1_U3439 , P1_U5541 );
and AND2_1202 ( P1_U3898 , P1_U5544 , P1_U3439 );
and AND2_1203 ( P1_U3899 , P1_U5546 , P1_U3439 );
and AND2_1204 ( P1_U3900 , P1_U5548 , P1_U3439 );
and AND2_1205 ( P1_U3901 , P1_U5550 , P1_U3439 );
and AND2_1206 ( P1_U3902 , P1_U5552 , P1_U3439 );
and AND2_1207 ( P1_U3903 , P1_U5554 , P1_U3439 );
and AND2_1208 ( P1_U3904 , P1_U5556 , P1_U3439 );
and AND2_1209 ( P1_U3905 , P1_U5558 , P1_U3439 );
and AND2_1210 ( P1_U3906 , P1_U5560 , P1_U3439 );
and AND2_1211 ( P1_U3907 , P1_U5562 , P1_U3439 );
and AND2_1212 ( P1_U3908 , P1_U3439 , P1_U5563 );
and AND2_1213 ( P1_U3909 , P1_U3439 , P1_U5565 );
and AND2_1214 ( P1_U3910 , P1_U3439 , P1_U5567 );
and AND2_1215 ( P1_U3911 , P1_U3439 , P1_U5569 );
and AND2_1216 ( P1_U3912 , P1_U3439 , P1_U5571 );
and AND2_1217 ( P1_U3913 , P1_U3439 , P1_U5573 );
and AND2_1218 ( P1_U3914 , P1_U3439 , P1_U5575 );
and AND2_1219 ( P1_U3915 , P1_U3439 , P1_U5577 );
and AND2_1220 ( P1_U3916 , P1_U3439 , P1_U5579 );
and AND2_1221 ( P1_U3917 , P1_U3439 , P1_U5581 );
and AND2_1222 ( P1_U3918 , P1_U3439 , P1_U5583 );
and AND2_1223 ( P1_U3919 , P1_U3439 , P1_U5585 );
and AND2_1224 ( P1_U3920 , P1_U3439 , P1_U5587 );
and AND2_1225 ( P1_U3921 , P1_U5606 , P1_U5604 );
and AND2_1226 ( P1_U3922 , P1_U5613 , P1_U5611 );
and AND2_1227 ( P1_U3923 , P1_U5619 , P1_U5617 );
and AND2_1228 ( P1_U3924 , P1_U5622 , P1_U5620 );
and AND2_1229 ( P1_U3925 , P1_U5625 , P1_U5623 );
and AND2_1230 ( P1_U3926 , P1_U5628 , P1_U5626 );
and AND2_1231 ( P1_U3927 , P1_U5631 , P1_U5629 );
and AND2_1232 ( P1_U3928 , P1_U5634 , P1_U5632 );
and AND2_1233 ( P1_U3929 , P1_U5637 , P1_U5635 );
and AND2_1234 ( P1_U3930 , P1_U5640 , P1_U5638 );
and AND2_1235 ( P1_U3931 , P1_U5643 , P1_U5641 );
and AND2_1236 ( P1_U3932 , P1_U5646 , P1_U5644 );
and AND2_1237 ( P1_U3933 , P1_U5649 , P1_U5647 );
and AND2_1238 ( P1_U3934 , P1_U5652 , P1_U5650 );
and AND2_1239 ( P1_U3935 , P1_U5655 , P1_U5653 );
and AND2_1240 ( P1_U3936 , P1_U5658 , P1_U5656 );
and AND2_1241 ( P1_U3937 , P1_U5661 , P1_U5659 );
and AND2_1242 ( P1_U3938 , P1_U5664 , P1_U5662 );
and AND2_1243 ( P1_U3939 , P1_U5667 , P1_U5665 );
and AND2_1244 ( P1_U3940 , P1_U5670 , P1_U5668 );
and AND2_1245 ( P1_U3941 , P1_U5673 , P1_U5671 );
and AND2_1246 ( P1_U3942 , P1_U5676 , P1_U5674 );
and AND2_1247 ( P1_U3943 , P1_U5679 , P1_U5677 );
not NOT1_1248 ( P1_U3944 , P1_IR_REG_31_ );
nand NAND2_1249 ( P1_U3945 , P1_U3022 , P1_U3359 );
nand NAND2_1250 ( P1_U3946 , P1_U5734 , P1_U5728 );
nand NAND2_1251 ( P1_U3947 , P1_U3634 , P1_U3047 );
nand NAND2_1252 ( P1_U3948 , P1_U3753 , P1_U3047 );
and AND2_1253 ( P1_U3949 , P1_U5968 , P1_U5967 );
and AND2_1254 ( P1_U3950 , P1_U5970 , P1_U5969 );
and AND2_1255 ( P1_U3951 , P1_U5972 , P1_U5971 );
and AND2_1256 ( P1_U3952 , P1_U5974 , P1_U5973 );
and AND2_1257 ( P1_U3953 , P1_U5976 , P1_U5975 );
and AND2_1258 ( P1_U3954 , P1_U5978 , P1_U5977 );
and AND2_1259 ( P1_U3955 , P1_U5980 , P1_U5979 );
and AND2_1260 ( P1_U3956 , P1_U5982 , P1_U5981 );
and AND2_1261 ( P1_U3957 , P1_U5984 , P1_U5983 );
and AND2_1262 ( P1_U3958 , P1_U5986 , P1_U5985 );
and AND2_1263 ( P1_U3959 , P1_U5988 , P1_U5987 );
and AND2_1264 ( P1_U3960 , P1_U5990 , P1_U5989 );
and AND2_1265 ( P1_U3961 , P1_U5992 , P1_U5991 );
and AND2_1266 ( P1_U3962 , P1_U5994 , P1_U5993 );
and AND2_1267 ( P1_U3963 , P1_U5996 , P1_U5995 );
and AND2_1268 ( P1_U3964 , P1_U5998 , P1_U5997 );
and AND2_1269 ( P1_U3965 , P1_U6000 , P1_U5999 );
and AND2_1270 ( P1_U3966 , P1_U6002 , P1_U6001 );
and AND2_1271 ( P1_U3967 , P1_U6004 , P1_U6003 );
and AND2_1272 ( P1_U3968 , P1_U6006 , P1_U6005 );
and AND2_1273 ( P1_U3969 , P1_U6008 , P1_U6007 );
and AND2_1274 ( P1_U3970 , P1_U6010 , P1_U6009 );
and AND2_1275 ( P1_U3971 , P1_U6012 , P1_U6011 );
and AND2_1276 ( P1_U3972 , P1_U6014 , P1_U6013 );
and AND2_1277 ( P1_U3973 , P1_U6016 , P1_U6015 );
and AND2_1278 ( P1_U3974 , P1_U6018 , P1_U6017 );
and AND2_1279 ( P1_U3975 , P1_U6020 , P1_U6019 );
and AND2_1280 ( P1_U3976 , P1_U6022 , P1_U6021 );
and AND2_1281 ( P1_U3977 , P1_U6024 , P1_U6023 );
and AND2_1282 ( P1_U3978 , P1_U6026 , P1_U6025 );
nand NAND2_1283 ( P1_U3979 , P1_U3752 , P1_U3054 );
and AND2_1284 ( P1_U3980 , P1_U6028 , P1_U6027 );
and AND2_1285 ( P1_U3981 , P1_U6030 , P1_U6029 );
nand NAND4_1286 ( P1_U3982 , P1_U3871 , P1_U3868 , P1_U3869 , P1_U3874 );
not NOT1_1287 ( P1_U3983 , P1_R1360_U14 );
and AND2_1288 ( P1_U3984 , P1_U6200 , P1_U6199 );
not NOT1_1289 ( P1_U3985 , P1_R1352_U6 );
not NOT1_1290 ( P1_U3986 , P1_U3371 );
not NOT1_1291 ( P1_U3987 , P1_U3428 );
not NOT1_1292 ( P1_U3988 , P1_U3426 );
not NOT1_1293 ( P1_U3989 , P1_U3369 );
not NOT1_1294 ( P1_U3990 , P1_U3419 );
not NOT1_1295 ( P1_U3991 , P1_U3365 );
not NOT1_1296 ( P1_U3992 , P1_U3364 );
not NOT1_1297 ( P1_U3993 , P1_U3367 );
not NOT1_1298 ( P1_U3994 , P1_U3360 );
not NOT1_1299 ( P1_U3995 , P1_U3363 );
not NOT1_1300 ( P1_U3996 , P1_U3361 );
not NOT1_1301 ( P1_U3997 , P1_U3420 );
not NOT1_1302 ( P1_U3998 , P1_U3418 );
nand NAND2_1303 ( P1_U3999 , P1_U3049 , P1_U4034 );
not NOT1_1304 ( P1_U4000 , P1_U3370 );
not NOT1_1305 ( P1_U4001 , P1_U3368 );
nand NAND2_1306 ( P1_U4002 , P1_U4020 , P1_U3366 );
nand NAND2_1307 ( P1_U4003 , P1_U3049 , P1_U3421 );
not NOT1_1308 ( P1_U4004 , P1_U3946 );
not NOT1_1309 ( P1_U4005 , P1_U3431 );
not NOT1_1310 ( P1_U4006 , P1_U3425 );
not NOT1_1311 ( P1_U4007 , P1_U3410 );
not NOT1_1312 ( P1_U4008 , P1_U3408 );
not NOT1_1313 ( P1_U4009 , P1_U3406 );
not NOT1_1314 ( P1_U4010 , P1_U3404 );
not NOT1_1315 ( P1_U4011 , P1_U3402 );
not NOT1_1316 ( P1_U4012 , P1_U3400 );
not NOT1_1317 ( P1_U4013 , P1_U3398 );
not NOT1_1318 ( P1_U4014 , P1_U3396 );
not NOT1_1319 ( P1_U4015 , P1_U3394 );
not NOT1_1320 ( P1_U4016 , P1_U3415 );
not NOT1_1321 ( P1_U4017 , P1_U3414 );
not NOT1_1322 ( P1_U4018 , P1_U3412 );
not NOT1_1323 ( P1_U4019 , P1_U3427 );
not NOT1_1324 ( P1_U4020 , P1_U3372 );
not NOT1_1325 ( P1_U4021 , P1_U3416 );
not NOT1_1326 ( P1_U4022 , P1_U3417 );
not NOT1_1327 ( P1_U4023 , P1_U3948 );
not NOT1_1328 ( P1_U4024 , P1_U3947 );
not NOT1_1329 ( P1_U4025 , P1_U3945 );
not NOT1_1330 ( P1_U4026 , P1_U3979 );
not NOT1_1331 ( P1_U4027 , P1_U3432 );
nand NAND2_1332 ( P1_U4028 , P1_U3433 , P1_STATE_REG );
nand NAND2_1333 ( P1_U4029 , P1_U3998 , P1_U3022 );
not NOT1_1334 ( P1_U4030 , P1_U3430 );
nand NAND2_1335 ( P1_U4031 , P1_U4006 , P1_U3210 );
not NOT1_1336 ( P1_U4032 , P1_U3424 );
not NOT1_1337 ( P1_U4033 , P1_U3434 );
not NOT1_1338 ( P1_U4034 , P1_U3362 );
not NOT1_1339 ( P1_U4035 , P1_U3366 );
not NOT1_1340 ( P1_U4036 , P1_U3357 );
not NOT1_1341 ( P1_U4037 , P1_U3356 );
nand NAND2_1342 ( P1_U4038 , U88 , P1_U3084 );
nand NAND2_1343 ( P1_U4039 , P1_IR_REG_0_ , P1_U3028 );
nand NAND2_1344 ( P1_U4040 , P1_IR_REG_0_ , P1_U4037 );
nand NAND2_1345 ( P1_U4041 , U77 , P1_U3084 );
nand NAND2_1346 ( P1_U4042 , P1_SUB_88_U40 , P1_U3028 );
nand NAND2_1347 ( P1_U4043 , P1_IR_REG_1_ , P1_U4037 );
nand NAND2_1348 ( P1_U4044 , U66 , P1_U3084 );
nand NAND2_1349 ( P1_U4045 , P1_SUB_88_U21 , P1_U3028 );
nand NAND2_1350 ( P1_U4046 , P1_IR_REG_2_ , P1_U4037 );
nand NAND2_1351 ( P1_U4047 , U63 , P1_U3084 );
nand NAND2_1352 ( P1_U4048 , P1_SUB_88_U22 , P1_U3028 );
nand NAND2_1353 ( P1_U4049 , P1_IR_REG_3_ , P1_U4037 );
nand NAND2_1354 ( P1_U4050 , U62 , P1_U3084 );
nand NAND2_1355 ( P1_U4051 , P1_SUB_88_U23 , P1_U3028 );
nand NAND2_1356 ( P1_U4052 , P1_IR_REG_4_ , P1_U4037 );
nand NAND2_1357 ( P1_U4053 , U61 , P1_U3084 );
nand NAND2_1358 ( P1_U4054 , P1_SUB_88_U162 , P1_U3028 );
nand NAND2_1359 ( P1_U4055 , P1_IR_REG_5_ , P1_U4037 );
nand NAND2_1360 ( P1_U4056 , U60 , P1_U3084 );
nand NAND2_1361 ( P1_U4057 , P1_SUB_88_U24 , P1_U3028 );
nand NAND2_1362 ( P1_U4058 , P1_IR_REG_6_ , P1_U4037 );
nand NAND2_1363 ( P1_U4059 , U59 , P1_U3084 );
nand NAND2_1364 ( P1_U4060 , P1_SUB_88_U25 , P1_U3028 );
nand NAND2_1365 ( P1_U4061 , P1_IR_REG_7_ , P1_U4037 );
nand NAND2_1366 ( P1_U4062 , U58 , P1_U3084 );
nand NAND2_1367 ( P1_U4063 , P1_SUB_88_U26 , P1_U3028 );
nand NAND2_1368 ( P1_U4064 , P1_IR_REG_8_ , P1_U4037 );
nand NAND2_1369 ( P1_U4065 , U57 , P1_U3084 );
nand NAND2_1370 ( P1_U4066 , P1_SUB_88_U160 , P1_U3028 );
nand NAND2_1371 ( P1_U4067 , P1_IR_REG_9_ , P1_U4037 );
nand NAND2_1372 ( P1_U4068 , U87 , P1_U3084 );
nand NAND2_1373 ( P1_U4069 , P1_SUB_88_U6 , P1_U3028 );
nand NAND2_1374 ( P1_U4070 , P1_IR_REG_10_ , P1_U4037 );
nand NAND2_1375 ( P1_U4071 , U86 , P1_U3084 );
nand NAND2_1376 ( P1_U4072 , P1_SUB_88_U7 , P1_U3028 );
nand NAND2_1377 ( P1_U4073 , P1_IR_REG_11_ , P1_U4037 );
nand NAND2_1378 ( P1_U4074 , U85 , P1_U3084 );
nand NAND2_1379 ( P1_U4075 , P1_SUB_88_U8 , P1_U3028 );
nand NAND2_1380 ( P1_U4076 , P1_IR_REG_12_ , P1_U4037 );
nand NAND2_1381 ( P1_U4077 , U84 , P1_U3084 );
nand NAND2_1382 ( P1_U4078 , P1_SUB_88_U179 , P1_U3028 );
nand NAND2_1383 ( P1_U4079 , P1_IR_REG_13_ , P1_U4037 );
nand NAND2_1384 ( P1_U4080 , U83 , P1_U3084 );
nand NAND2_1385 ( P1_U4081 , P1_SUB_88_U9 , P1_U3028 );
nand NAND2_1386 ( P1_U4082 , P1_IR_REG_14_ , P1_U4037 );
nand NAND2_1387 ( P1_U4083 , U82 , P1_U3084 );
nand NAND2_1388 ( P1_U4084 , P1_SUB_88_U10 , P1_U3028 );
nand NAND2_1389 ( P1_U4085 , P1_IR_REG_15_ , P1_U4037 );
nand NAND2_1390 ( P1_U4086 , U81 , P1_U3084 );
nand NAND2_1391 ( P1_U4087 , P1_SUB_88_U11 , P1_U3028 );
nand NAND2_1392 ( P1_U4088 , P1_IR_REG_16_ , P1_U4037 );
nand NAND2_1393 ( P1_U4089 , U80 , P1_U3084 );
nand NAND2_1394 ( P1_U4090 , P1_SUB_88_U177 , P1_U3028 );
nand NAND2_1395 ( P1_U4091 , P1_IR_REG_17_ , P1_U4037 );
nand NAND2_1396 ( P1_U4092 , U79 , P1_U3084 );
nand NAND2_1397 ( P1_U4093 , P1_SUB_88_U12 , P1_U3028 );
nand NAND2_1398 ( P1_U4094 , P1_IR_REG_18_ , P1_U4037 );
nand NAND2_1399 ( P1_U4095 , U78 , P1_U3084 );
nand NAND2_1400 ( P1_U4096 , P1_SUB_88_U13 , P1_U3028 );
nand NAND2_1401 ( P1_U4097 , P1_IR_REG_19_ , P1_U4037 );
nand NAND2_1402 ( P1_U4098 , U76 , P1_U3084 );
nand NAND2_1403 ( P1_U4099 , P1_SUB_88_U14 , P1_U3028 );
nand NAND2_1404 ( P1_U4100 , P1_IR_REG_20_ , P1_U4037 );
nand NAND2_1405 ( P1_U4101 , U75 , P1_U3084 );
nand NAND2_1406 ( P1_U4102 , P1_SUB_88_U173 , P1_U3028 );
nand NAND2_1407 ( P1_U4103 , P1_IR_REG_21_ , P1_U4037 );
nand NAND2_1408 ( P1_U4104 , U74 , P1_U3084 );
nand NAND2_1409 ( P1_U4105 , P1_SUB_88_U15 , P1_U3028 );
nand NAND2_1410 ( P1_U4106 , P1_IR_REG_22_ , P1_U4037 );
nand NAND2_1411 ( P1_U4107 , U73 , P1_U3084 );
nand NAND2_1412 ( P1_U4108 , P1_SUB_88_U16 , P1_U3028 );
nand NAND2_1413 ( P1_U4109 , P1_IR_REG_23_ , P1_U4037 );
nand NAND2_1414 ( P1_U4110 , U72 , P1_U3084 );
nand NAND2_1415 ( P1_U4111 , P1_SUB_88_U17 , P1_U3028 );
nand NAND2_1416 ( P1_U4112 , P1_IR_REG_24_ , P1_U4037 );
nand NAND2_1417 ( P1_U4113 , U71 , P1_U3084 );
nand NAND2_1418 ( P1_U4114 , P1_SUB_88_U170 , P1_U3028 );
nand NAND2_1419 ( P1_U4115 , P1_IR_REG_25_ , P1_U4037 );
nand NAND2_1420 ( P1_U4116 , U70 , P1_U3084 );
nand NAND2_1421 ( P1_U4117 , P1_SUB_88_U18 , P1_U3028 );
nand NAND2_1422 ( P1_U4118 , P1_IR_REG_26_ , P1_U4037 );
nand NAND2_1423 ( P1_U4119 , U69 , P1_U3084 );
nand NAND2_1424 ( P1_U4120 , P1_SUB_88_U42 , P1_U3028 );
nand NAND2_1425 ( P1_U4121 , P1_IR_REG_27_ , P1_U4037 );
nand NAND2_1426 ( P1_U4122 , U68 , P1_U3084 );
nand NAND2_1427 ( P1_U4123 , P1_SUB_88_U19 , P1_U3028 );
nand NAND2_1428 ( P1_U4124 , P1_IR_REG_28_ , P1_U4037 );
nand NAND2_1429 ( P1_U4125 , U67 , P1_U3084 );
nand NAND2_1430 ( P1_U4126 , P1_SUB_88_U20 , P1_U3028 );
nand NAND2_1431 ( P1_U4127 , P1_IR_REG_29_ , P1_U4037 );
nand NAND2_1432 ( P1_U4128 , U65 , P1_U3084 );
nand NAND2_1433 ( P1_U4129 , P1_SUB_88_U165 , P1_U3028 );
nand NAND2_1434 ( P1_U4130 , P1_IR_REG_30_ , P1_U4037 );
nand NAND2_1435 ( P1_U4131 , U64 , P1_U3084 );
nand NAND2_1436 ( P1_U4132 , P1_SUB_88_U41 , P1_U3028 );
nand NAND2_1437 ( P1_U4133 , P1_IR_REG_31_ , P1_U4037 );
not NOT1_1438 ( P1_U4134 , P1_U3359 );
not NOT1_1439 ( P1_U4135 , P1_U3421 );
nand NAND2_1440 ( P1_U4136 , P1_U3357 , P1_U5692 );
nand NAND2_1441 ( P1_U4137 , P1_U3357 , P1_U5695 );
nand NAND2_1442 ( P1_U4138 , P1_U4134 , P1_D_REG_10_ );
nand NAND2_1443 ( P1_U4139 , P1_U4134 , P1_D_REG_11_ );
nand NAND2_1444 ( P1_U4140 , P1_U4134 , P1_D_REG_12_ );
nand NAND2_1445 ( P1_U4141 , P1_U4134 , P1_D_REG_13_ );
nand NAND2_1446 ( P1_U4142 , P1_U4134 , P1_D_REG_14_ );
nand NAND2_1447 ( P1_U4143 , P1_U4134 , P1_D_REG_15_ );
nand NAND2_1448 ( P1_U4144 , P1_U4134 , P1_D_REG_16_ );
nand NAND2_1449 ( P1_U4145 , P1_U4134 , P1_D_REG_17_ );
nand NAND2_1450 ( P1_U4146 , P1_U4134 , P1_D_REG_18_ );
nand NAND2_1451 ( P1_U4147 , P1_U4134 , P1_D_REG_19_ );
nand NAND2_1452 ( P1_U4148 , P1_U4134 , P1_D_REG_20_ );
nand NAND2_1453 ( P1_U4149 , P1_U4134 , P1_D_REG_21_ );
nand NAND2_1454 ( P1_U4150 , P1_U4134 , P1_D_REG_22_ );
nand NAND2_1455 ( P1_U4151 , P1_U4134 , P1_D_REG_23_ );
nand NAND2_1456 ( P1_U4152 , P1_U4134 , P1_D_REG_24_ );
nand NAND2_1457 ( P1_U4153 , P1_U4134 , P1_D_REG_25_ );
nand NAND2_1458 ( P1_U4154 , P1_U4134 , P1_D_REG_26_ );
nand NAND2_1459 ( P1_U4155 , P1_U4134 , P1_D_REG_27_ );
nand NAND2_1460 ( P1_U4156 , P1_U4134 , P1_D_REG_28_ );
nand NAND2_1461 ( P1_U4157 , P1_U4134 , P1_D_REG_29_ );
nand NAND2_1462 ( P1_U4158 , P1_U4134 , P1_D_REG_2_ );
nand NAND2_1463 ( P1_U4159 , P1_U4134 , P1_D_REG_30_ );
nand NAND2_1464 ( P1_U4160 , P1_U4134 , P1_D_REG_31_ );
nand NAND2_1465 ( P1_U4161 , P1_U4134 , P1_D_REG_3_ );
nand NAND2_1466 ( P1_U4162 , P1_U4134 , P1_D_REG_4_ );
nand NAND2_1467 ( P1_U4163 , P1_U4134 , P1_D_REG_5_ );
nand NAND2_1468 ( P1_U4164 , P1_U4134 , P1_D_REG_6_ );
nand NAND2_1469 ( P1_U4165 , P1_U4134 , P1_D_REG_7_ );
nand NAND2_1470 ( P1_U4166 , P1_U4134 , P1_D_REG_8_ );
nand NAND2_1471 ( P1_U4167 , P1_U4134 , P1_D_REG_9_ );
nand NAND2_1472 ( P1_U4168 , P1_U5716 , P1_U5719 );
nand NAND3_1473 ( P1_U4169 , P1_U5739 , P1_U5738 , P1_U3366 );
nand NAND2_1474 ( P1_U4170 , P1_U3018 , P1_REG2_REG_1_ );
nand NAND2_1475 ( P1_U4171 , P1_U3019 , P1_REG1_REG_1_ );
nand NAND2_1476 ( P1_U4172 , P1_U3020 , P1_REG0_REG_1_ );
nand NAND2_1477 ( P1_U4173 , P1_REG3_REG_1_ , P1_U3017 );
not NOT1_1478 ( P1_U4174 , P1_U3076 );
nand NAND2_1479 ( P1_U4175 , P1_U3999 , P1_U3416 );
nand NAND2_1480 ( P1_U4176 , P1_U3994 , P1_R1150_U21 );
nand NAND2_1481 ( P1_U4177 , P1_U3996 , P1_R1117_U21 );
nand NAND2_1482 ( P1_U4178 , P1_U3995 , P1_R1138_U96 );
nand NAND2_1483 ( P1_U4179 , P1_U3992 , P1_R1192_U21 );
nand NAND2_1484 ( P1_U4180 , P1_U3991 , P1_R1207_U21 );
nand NAND2_1485 ( P1_U4181 , P1_U4001 , P1_R1171_U96 );
nand NAND2_1486 ( P1_U4182 , P1_U4000 , P1_R1240_U96 );
not NOT1_1487 ( P1_U4183 , P1_U3373 );
nand NAND2_1488 ( P1_U4184 , P1_R1222_U96 , P1_U3026 );
nand NAND2_1489 ( P1_U4185 , P1_U3025 , P1_U3076 );
nand NAND2_1490 ( P1_U4186 , P1_U3451 , P1_U3023 );
nand NAND2_1491 ( P1_U4187 , P1_U3451 , P1_U4175 );
nand NAND2_1492 ( P1_U4188 , P1_U3622 , P1_U4183 );
nand NAND2_1493 ( P1_U4189 , P1_REG2_REG_2_ , P1_U3018 );
nand NAND2_1494 ( P1_U4190 , P1_REG1_REG_2_ , P1_U3019 );
nand NAND2_1495 ( P1_U4191 , P1_REG0_REG_2_ , P1_U3020 );
nand NAND2_1496 ( P1_U4192 , P1_REG3_REG_2_ , P1_U3017 );
not NOT1_1497 ( P1_U4193 , P1_U3066 );
nand NAND2_1498 ( P1_U4194 , P1_REG0_REG_0_ , P1_U3020 );
nand NAND2_1499 ( P1_U4195 , P1_REG1_REG_0_ , P1_U3019 );
nand NAND2_1500 ( P1_U4196 , P1_REG2_REG_0_ , P1_U3018 );
nand NAND2_1501 ( P1_U4197 , P1_REG3_REG_0_ , P1_U3017 );
not NOT1_1502 ( P1_U4198 , P1_U3075 );
nand NAND2_1503 ( P1_U4199 , P1_U3033 , P1_U3075 );
nand NAND2_1504 ( P1_U4200 , P1_R1150_U98 , P1_U3994 );
nand NAND2_1505 ( P1_U4201 , P1_R1117_U98 , P1_U3996 );
nand NAND2_1506 ( P1_U4202 , P1_R1138_U95 , P1_U3995 );
nand NAND2_1507 ( P1_U4203 , P1_R1192_U98 , P1_U3992 );
nand NAND2_1508 ( P1_U4204 , P1_R1207_U98 , P1_U3991 );
nand NAND2_1509 ( P1_U4205 , P1_R1171_U95 , P1_U4001 );
nand NAND2_1510 ( P1_U4206 , P1_R1240_U95 , P1_U4000 );
not NOT1_1511 ( P1_U4207 , P1_U3375 );
nand NAND2_1512 ( P1_U4208 , P1_R1222_U95 , P1_U3026 );
nand NAND2_1513 ( P1_U4209 , P1_U3025 , P1_U3066 );
nand NAND2_1514 ( P1_U4210 , P1_R1282_U57 , P1_U3023 );
nand NAND2_1515 ( P1_U4211 , P1_U3456 , P1_U4175 );
nand NAND2_1516 ( P1_U4212 , P1_U3638 , P1_U4207 );
nand NAND2_1517 ( P1_U4213 , P1_REG2_REG_3_ , P1_U3018 );
nand NAND2_1518 ( P1_U4214 , P1_REG1_REG_3_ , P1_U3019 );
nand NAND2_1519 ( P1_U4215 , P1_REG0_REG_3_ , P1_U3020 );
nand NAND2_1520 ( P1_U4216 , P1_ADD_99_U4 , P1_U3017 );
not NOT1_1521 ( P1_U4217 , P1_U3062 );
nand NAND2_1522 ( P1_U4218 , P1_U3033 , P1_U3076 );
nand NAND2_1523 ( P1_U4219 , P1_R1150_U108 , P1_U3994 );
nand NAND2_1524 ( P1_U4220 , P1_R1117_U108 , P1_U3996 );
nand NAND2_1525 ( P1_U4221 , P1_R1138_U17 , P1_U3995 );
nand NAND2_1526 ( P1_U4222 , P1_R1192_U108 , P1_U3992 );
nand NAND2_1527 ( P1_U4223 , P1_R1207_U108 , P1_U3991 );
nand NAND2_1528 ( P1_U4224 , P1_R1171_U17 , P1_U4001 );
nand NAND2_1529 ( P1_U4225 , P1_R1240_U17 , P1_U4000 );
not NOT1_1530 ( P1_U4226 , P1_U3376 );
nand NAND2_1531 ( P1_U4227 , P1_R1222_U17 , P1_U3026 );
nand NAND2_1532 ( P1_U4228 , P1_U3025 , P1_U3062 );
nand NAND2_1533 ( P1_U4229 , P1_R1282_U18 , P1_U3023 );
nand NAND2_1534 ( P1_U4230 , P1_U3459 , P1_U4175 );
nand NAND2_1535 ( P1_U4231 , P1_U3642 , P1_U4226 );
nand NAND2_1536 ( P1_U4232 , P1_REG2_REG_4_ , P1_U3018 );
nand NAND2_1537 ( P1_U4233 , P1_REG1_REG_4_ , P1_U3019 );
nand NAND2_1538 ( P1_U4234 , P1_REG0_REG_4_ , P1_U3020 );
nand NAND2_1539 ( P1_U4235 , P1_ADD_99_U59 , P1_U3017 );
not NOT1_1540 ( P1_U4236 , P1_U3058 );
nand NAND2_1541 ( P1_U4237 , P1_U3033 , P1_U3066 );
nand NAND2_1542 ( P1_U4238 , P1_R1150_U18 , P1_U3994 );
nand NAND2_1543 ( P1_U4239 , P1_R1117_U18 , P1_U3996 );
nand NAND2_1544 ( P1_U4240 , P1_R1138_U101 , P1_U3995 );
nand NAND2_1545 ( P1_U4241 , P1_R1192_U18 , P1_U3992 );
nand NAND2_1546 ( P1_U4242 , P1_R1207_U18 , P1_U3991 );
nand NAND2_1547 ( P1_U4243 , P1_R1171_U101 , P1_U4001 );
nand NAND2_1548 ( P1_U4244 , P1_R1240_U101 , P1_U4000 );
not NOT1_1549 ( P1_U4245 , P1_U3377 );
nand NAND2_1550 ( P1_U4246 , P1_R1222_U101 , P1_U3026 );
nand NAND2_1551 ( P1_U4247 , P1_U3025 , P1_U3058 );
nand NAND2_1552 ( P1_U4248 , P1_R1282_U20 , P1_U3023 );
nand NAND2_1553 ( P1_U4249 , P1_U3462 , P1_U4175 );
nand NAND2_1554 ( P1_U4250 , P1_U3646 , P1_U4245 );
nand NAND2_1555 ( P1_U4251 , P1_REG2_REG_5_ , P1_U3018 );
nand NAND2_1556 ( P1_U4252 , P1_REG1_REG_5_ , P1_U3019 );
nand NAND2_1557 ( P1_U4253 , P1_REG0_REG_5_ , P1_U3020 );
nand NAND2_1558 ( P1_U4254 , P1_ADD_99_U58 , P1_U3017 );
not NOT1_1559 ( P1_U4255 , P1_U3065 );
nand NAND2_1560 ( P1_U4256 , P1_U3033 , P1_U3062 );
nand NAND2_1561 ( P1_U4257 , P1_R1150_U107 , P1_U3994 );
nand NAND2_1562 ( P1_U4258 , P1_R1117_U107 , P1_U3996 );
nand NAND2_1563 ( P1_U4259 , P1_R1138_U100 , P1_U3995 );
nand NAND2_1564 ( P1_U4260 , P1_R1192_U107 , P1_U3992 );
nand NAND2_1565 ( P1_U4261 , P1_R1207_U107 , P1_U3991 );
nand NAND2_1566 ( P1_U4262 , P1_R1171_U100 , P1_U4001 );
nand NAND2_1567 ( P1_U4263 , P1_R1240_U100 , P1_U4000 );
not NOT1_1568 ( P1_U4264 , P1_U3378 );
nand NAND2_1569 ( P1_U4265 , P1_R1222_U100 , P1_U3026 );
nand NAND2_1570 ( P1_U4266 , P1_U3025 , P1_U3065 );
nand NAND2_1571 ( P1_U4267 , P1_R1282_U21 , P1_U3023 );
nand NAND2_1572 ( P1_U4268 , P1_U3465 , P1_U4175 );
nand NAND2_1573 ( P1_U4269 , P1_U3650 , P1_U4264 );
nand NAND2_1574 ( P1_U4270 , P1_REG2_REG_6_ , P1_U3018 );
nand NAND2_1575 ( P1_U4271 , P1_REG1_REG_6_ , P1_U3019 );
nand NAND2_1576 ( P1_U4272 , P1_REG0_REG_6_ , P1_U3020 );
nand NAND2_1577 ( P1_U4273 , P1_ADD_99_U57 , P1_U3017 );
not NOT1_1578 ( P1_U4274 , P1_U3069 );
nand NAND2_1579 ( P1_U4275 , P1_U3033 , P1_U3058 );
nand NAND2_1580 ( P1_U4276 , P1_R1150_U106 , P1_U3994 );
nand NAND2_1581 ( P1_U4277 , P1_R1117_U106 , P1_U3996 );
nand NAND2_1582 ( P1_U4278 , P1_R1138_U18 , P1_U3995 );
nand NAND2_1583 ( P1_U4279 , P1_R1192_U106 , P1_U3992 );
nand NAND2_1584 ( P1_U4280 , P1_R1207_U106 , P1_U3991 );
nand NAND2_1585 ( P1_U4281 , P1_R1171_U18 , P1_U4001 );
nand NAND2_1586 ( P1_U4282 , P1_R1240_U18 , P1_U4000 );
not NOT1_1587 ( P1_U4283 , P1_U3379 );
nand NAND2_1588 ( P1_U4284 , P1_R1222_U18 , P1_U3026 );
nand NAND2_1589 ( P1_U4285 , P1_U3025 , P1_U3069 );
nand NAND2_1590 ( P1_U4286 , P1_R1282_U65 , P1_U3023 );
nand NAND2_1591 ( P1_U4287 , P1_U3468 , P1_U4175 );
nand NAND2_1592 ( P1_U4288 , P1_U3654 , P1_U4283 );
nand NAND2_1593 ( P1_U4289 , P1_REG2_REG_7_ , P1_U3018 );
nand NAND2_1594 ( P1_U4290 , P1_REG1_REG_7_ , P1_U3019 );
nand NAND2_1595 ( P1_U4291 , P1_REG0_REG_7_ , P1_U3020 );
nand NAND2_1596 ( P1_U4292 , P1_ADD_99_U56 , P1_U3017 );
not NOT1_1597 ( P1_U4293 , P1_U3068 );
nand NAND2_1598 ( P1_U4294 , P1_U3033 , P1_U3065 );
nand NAND2_1599 ( P1_U4295 , P1_R1150_U19 , P1_U3994 );
nand NAND2_1600 ( P1_U4296 , P1_R1117_U19 , P1_U3996 );
nand NAND2_1601 ( P1_U4297 , P1_R1138_U99 , P1_U3995 );
nand NAND2_1602 ( P1_U4298 , P1_R1192_U19 , P1_U3992 );
nand NAND2_1603 ( P1_U4299 , P1_R1207_U19 , P1_U3991 );
nand NAND2_1604 ( P1_U4300 , P1_R1171_U99 , P1_U4001 );
nand NAND2_1605 ( P1_U4301 , P1_R1240_U99 , P1_U4000 );
not NOT1_1606 ( P1_U4302 , P1_U3380 );
nand NAND2_1607 ( P1_U4303 , P1_R1222_U99 , P1_U3026 );
nand NAND2_1608 ( P1_U4304 , P1_U3025 , P1_U3068 );
nand NAND2_1609 ( P1_U4305 , P1_R1282_U22 , P1_U3023 );
nand NAND2_1610 ( P1_U4306 , P1_U3471 , P1_U4175 );
nand NAND2_1611 ( P1_U4307 , P1_U3658 , P1_U4302 );
nand NAND2_1612 ( P1_U4308 , P1_REG2_REG_8_ , P1_U3018 );
nand NAND2_1613 ( P1_U4309 , P1_REG1_REG_8_ , P1_U3019 );
nand NAND2_1614 ( P1_U4310 , P1_REG0_REG_8_ , P1_U3020 );
nand NAND2_1615 ( P1_U4311 , P1_ADD_99_U55 , P1_U3017 );
not NOT1_1616 ( P1_U4312 , P1_U3082 );
nand NAND2_1617 ( P1_U4313 , P1_U3033 , P1_U3069 );
nand NAND2_1618 ( P1_U4314 , P1_R1150_U105 , P1_U3994 );
nand NAND2_1619 ( P1_U4315 , P1_R1117_U105 , P1_U3996 );
nand NAND2_1620 ( P1_U4316 , P1_R1138_U19 , P1_U3995 );
nand NAND2_1621 ( P1_U4317 , P1_R1192_U105 , P1_U3992 );
nand NAND2_1622 ( P1_U4318 , P1_R1207_U105 , P1_U3991 );
nand NAND2_1623 ( P1_U4319 , P1_R1171_U19 , P1_U4001 );
nand NAND2_1624 ( P1_U4320 , P1_R1240_U19 , P1_U4000 );
not NOT1_1625 ( P1_U4321 , P1_U3381 );
nand NAND2_1626 ( P1_U4322 , P1_R1222_U19 , P1_U3026 );
nand NAND2_1627 ( P1_U4323 , P1_U3025 , P1_U3082 );
nand NAND2_1628 ( P1_U4324 , P1_R1282_U23 , P1_U3023 );
nand NAND2_1629 ( P1_U4325 , P1_U3474 , P1_U4175 );
nand NAND2_1630 ( P1_U4326 , P1_U3662 , P1_U4321 );
nand NAND2_1631 ( P1_U4327 , P1_REG2_REG_9_ , P1_U3018 );
nand NAND2_1632 ( P1_U4328 , P1_REG1_REG_9_ , P1_U3019 );
nand NAND2_1633 ( P1_U4329 , P1_REG0_REG_9_ , P1_U3020 );
nand NAND2_1634 ( P1_U4330 , P1_ADD_99_U54 , P1_U3017 );
not NOT1_1635 ( P1_U4331 , P1_U3081 );
nand NAND2_1636 ( P1_U4332 , P1_U3033 , P1_U3068 );
nand NAND2_1637 ( P1_U4333 , P1_R1150_U20 , P1_U3994 );
nand NAND2_1638 ( P1_U4334 , P1_R1117_U20 , P1_U3996 );
nand NAND2_1639 ( P1_U4335 , P1_R1138_U98 , P1_U3995 );
nand NAND2_1640 ( P1_U4336 , P1_R1192_U20 , P1_U3992 );
nand NAND2_1641 ( P1_U4337 , P1_R1207_U20 , P1_U3991 );
nand NAND2_1642 ( P1_U4338 , P1_R1171_U98 , P1_U4001 );
nand NAND2_1643 ( P1_U4339 , P1_R1240_U98 , P1_U4000 );
not NOT1_1644 ( P1_U4340 , P1_U3382 );
nand NAND2_1645 ( P1_U4341 , P1_R1222_U98 , P1_U3026 );
nand NAND2_1646 ( P1_U4342 , P1_U3025 , P1_U3081 );
nand NAND2_1647 ( P1_U4343 , P1_R1282_U24 , P1_U3023 );
nand NAND2_1648 ( P1_U4344 , P1_U3477 , P1_U4175 );
nand NAND2_1649 ( P1_U4345 , P1_U3666 , P1_U4340 );
nand NAND2_1650 ( P1_U4346 , P1_REG2_REG_10_ , P1_U3018 );
nand NAND2_1651 ( P1_U4347 , P1_REG1_REG_10_ , P1_U3019 );
nand NAND2_1652 ( P1_U4348 , P1_REG0_REG_10_ , P1_U3020 );
nand NAND2_1653 ( P1_U4349 , P1_ADD_99_U78 , P1_U3017 );
not NOT1_1654 ( P1_U4350 , P1_U3060 );
nand NAND2_1655 ( P1_U4351 , P1_U3033 , P1_U3082 );
nand NAND2_1656 ( P1_U4352 , P1_R1150_U104 , P1_U3994 );
nand NAND2_1657 ( P1_U4353 , P1_R1117_U104 , P1_U3996 );
nand NAND2_1658 ( P1_U4354 , P1_R1138_U97 , P1_U3995 );
nand NAND2_1659 ( P1_U4355 , P1_R1192_U104 , P1_U3992 );
nand NAND2_1660 ( P1_U4356 , P1_R1207_U104 , P1_U3991 );
nand NAND2_1661 ( P1_U4357 , P1_R1171_U97 , P1_U4001 );
nand NAND2_1662 ( P1_U4358 , P1_R1240_U97 , P1_U4000 );
not NOT1_1663 ( P1_U4359 , P1_U3383 );
nand NAND2_1664 ( P1_U4360 , P1_R1222_U97 , P1_U3026 );
nand NAND2_1665 ( P1_U4361 , P1_U3025 , P1_U3060 );
nand NAND2_1666 ( P1_U4362 , P1_R1282_U63 , P1_U3023 );
nand NAND2_1667 ( P1_U4363 , P1_U3480 , P1_U4175 );
nand NAND2_1668 ( P1_U4364 , P1_U3670 , P1_U4359 );
nand NAND2_1669 ( P1_U4365 , P1_REG2_REG_11_ , P1_U3018 );
nand NAND2_1670 ( P1_U4366 , P1_REG1_REG_11_ , P1_U3019 );
nand NAND2_1671 ( P1_U4367 , P1_REG0_REG_11_ , P1_U3020 );
nand NAND2_1672 ( P1_U4368 , P1_ADD_99_U77 , P1_U3017 );
not NOT1_1673 ( P1_U4369 , P1_U3061 );
nand NAND2_1674 ( P1_U4370 , P1_U3033 , P1_U3081 );
nand NAND2_1675 ( P1_U4371 , P1_R1150_U114 , P1_U3994 );
nand NAND2_1676 ( P1_U4372 , P1_R1117_U114 , P1_U3996 );
nand NAND2_1677 ( P1_U4373 , P1_R1138_U11 , P1_U3995 );
nand NAND2_1678 ( P1_U4374 , P1_R1192_U114 , P1_U3992 );
nand NAND2_1679 ( P1_U4375 , P1_R1207_U114 , P1_U3991 );
nand NAND2_1680 ( P1_U4376 , P1_R1171_U11 , P1_U4001 );
nand NAND2_1681 ( P1_U4377 , P1_R1240_U11 , P1_U4000 );
not NOT1_1682 ( P1_U4378 , P1_U3384 );
nand NAND2_1683 ( P1_U4379 , P1_R1222_U11 , P1_U3026 );
nand NAND2_1684 ( P1_U4380 , P1_U3025 , P1_U3061 );
nand NAND2_1685 ( P1_U4381 , P1_R1282_U6 , P1_U3023 );
nand NAND2_1686 ( P1_U4382 , P1_U3483 , P1_U4175 );
nand NAND2_1687 ( P1_U4383 , P1_U3674 , P1_U4378 );
nand NAND2_1688 ( P1_U4384 , P1_REG2_REG_12_ , P1_U3018 );
nand NAND2_1689 ( P1_U4385 , P1_REG1_REG_12_ , P1_U3019 );
nand NAND2_1690 ( P1_U4386 , P1_REG0_REG_12_ , P1_U3020 );
nand NAND2_1691 ( P1_U4387 , P1_ADD_99_U76 , P1_U3017 );
not NOT1_1692 ( P1_U4388 , P1_U3070 );
nand NAND2_1693 ( P1_U4389 , P1_U3033 , P1_U3060 );
nand NAND2_1694 ( P1_U4390 , P1_R1150_U13 , P1_U3994 );
nand NAND2_1695 ( P1_U4391 , P1_R1117_U13 , P1_U3996 );
nand NAND2_1696 ( P1_U4392 , P1_R1138_U115 , P1_U3995 );
nand NAND2_1697 ( P1_U4393 , P1_R1192_U13 , P1_U3992 );
nand NAND2_1698 ( P1_U4394 , P1_R1207_U13 , P1_U3991 );
nand NAND2_1699 ( P1_U4395 , P1_R1171_U115 , P1_U4001 );
nand NAND2_1700 ( P1_U4396 , P1_R1240_U115 , P1_U4000 );
not NOT1_1701 ( P1_U4397 , P1_U3385 );
nand NAND2_1702 ( P1_U4398 , P1_R1222_U115 , P1_U3026 );
nand NAND2_1703 ( P1_U4399 , P1_U3025 , P1_U3070 );
nand NAND2_1704 ( P1_U4400 , P1_R1282_U7 , P1_U3023 );
nand NAND2_1705 ( P1_U4401 , P1_U3486 , P1_U4175 );
nand NAND2_1706 ( P1_U4402 , P1_U3678 , P1_U4397 );
nand NAND2_1707 ( P1_U4403 , P1_REG2_REG_13_ , P1_U3018 );
nand NAND2_1708 ( P1_U4404 , P1_REG1_REG_13_ , P1_U3019 );
nand NAND2_1709 ( P1_U4405 , P1_REG0_REG_13_ , P1_U3020 );
nand NAND2_1710 ( P1_U4406 , P1_ADD_99_U75 , P1_U3017 );
not NOT1_1711 ( P1_U4407 , P1_U3078 );
nand NAND2_1712 ( P1_U4408 , P1_U3033 , P1_U3061 );
nand NAND2_1713 ( P1_U4409 , P1_R1150_U103 , P1_U3994 );
nand NAND2_1714 ( P1_U4410 , P1_R1117_U103 , P1_U3996 );
nand NAND2_1715 ( P1_U4411 , P1_R1138_U114 , P1_U3995 );
nand NAND2_1716 ( P1_U4412 , P1_R1192_U103 , P1_U3992 );
nand NAND2_1717 ( P1_U4413 , P1_R1207_U103 , P1_U3991 );
nand NAND2_1718 ( P1_U4414 , P1_R1171_U114 , P1_U4001 );
nand NAND2_1719 ( P1_U4415 , P1_R1240_U114 , P1_U4000 );
not NOT1_1720 ( P1_U4416 , P1_U3386 );
nand NAND2_1721 ( P1_U4417 , P1_R1222_U114 , P1_U3026 );
nand NAND2_1722 ( P1_U4418 , P1_U3025 , P1_U3078 );
nand NAND2_1723 ( P1_U4419 , P1_R1282_U8 , P1_U3023 );
nand NAND2_1724 ( P1_U4420 , P1_U3489 , P1_U4175 );
nand NAND2_1725 ( P1_U4421 , P1_U3682 , P1_U4416 );
nand NAND2_1726 ( P1_U4422 , P1_REG2_REG_14_ , P1_U3018 );
nand NAND2_1727 ( P1_U4423 , P1_REG1_REG_14_ , P1_U3019 );
nand NAND2_1728 ( P1_U4424 , P1_REG0_REG_14_ , P1_U3020 );
nand NAND2_1729 ( P1_U4425 , P1_ADD_99_U74 , P1_U3017 );
not NOT1_1730 ( P1_U4426 , P1_U3077 );
nand NAND2_1731 ( P1_U4427 , P1_U3033 , P1_U3070 );
nand NAND2_1732 ( P1_U4428 , P1_R1150_U102 , P1_U3994 );
nand NAND2_1733 ( P1_U4429 , P1_R1117_U102 , P1_U3996 );
nand NAND2_1734 ( P1_U4430 , P1_R1138_U12 , P1_U3995 );
nand NAND2_1735 ( P1_U4431 , P1_R1192_U102 , P1_U3992 );
nand NAND2_1736 ( P1_U4432 , P1_R1207_U102 , P1_U3991 );
nand NAND2_1737 ( P1_U4433 , P1_R1171_U12 , P1_U4001 );
nand NAND2_1738 ( P1_U4434 , P1_R1240_U12 , P1_U4000 );
not NOT1_1739 ( P1_U4435 , P1_U3387 );
nand NAND2_1740 ( P1_U4436 , P1_R1222_U12 , P1_U3026 );
nand NAND2_1741 ( P1_U4437 , P1_U3025 , P1_U3077 );
nand NAND2_1742 ( P1_U4438 , P1_R1282_U86 , P1_U3023 );
nand NAND2_1743 ( P1_U4439 , P1_U3492 , P1_U4175 );
nand NAND2_1744 ( P1_U4440 , P1_U3686 , P1_U4435 );
nand NAND2_1745 ( P1_U4441 , P1_REG2_REG_15_ , P1_U3018 );
nand NAND2_1746 ( P1_U4442 , P1_REG1_REG_15_ , P1_U3019 );
nand NAND2_1747 ( P1_U4443 , P1_REG0_REG_15_ , P1_U3020 );
nand NAND2_1748 ( P1_U4444 , P1_ADD_99_U73 , P1_U3017 );
not NOT1_1749 ( P1_U4445 , P1_U3072 );
nand NAND2_1750 ( P1_U4446 , P1_U3033 , P1_U3078 );
nand NAND2_1751 ( P1_U4447 , P1_R1150_U113 , P1_U3994 );
nand NAND2_1752 ( P1_U4448 , P1_R1117_U113 , P1_U3996 );
nand NAND2_1753 ( P1_U4449 , P1_R1138_U113 , P1_U3995 );
nand NAND2_1754 ( P1_U4450 , P1_R1192_U113 , P1_U3992 );
nand NAND2_1755 ( P1_U4451 , P1_R1207_U113 , P1_U3991 );
nand NAND2_1756 ( P1_U4452 , P1_R1171_U113 , P1_U4001 );
nand NAND2_1757 ( P1_U4453 , P1_R1240_U113 , P1_U4000 );
not NOT1_1758 ( P1_U4454 , P1_U3388 );
nand NAND2_1759 ( P1_U4455 , P1_R1222_U113 , P1_U3026 );
nand NAND2_1760 ( P1_U4456 , P1_U3025 , P1_U3072 );
nand NAND2_1761 ( P1_U4457 , P1_R1282_U9 , P1_U3023 );
nand NAND2_1762 ( P1_U4458 , P1_U3495 , P1_U4175 );
nand NAND2_1763 ( P1_U4459 , P1_U3690 , P1_U4454 );
nand NAND2_1764 ( P1_U4460 , P1_REG2_REG_16_ , P1_U3018 );
nand NAND2_1765 ( P1_U4461 , P1_REG1_REG_16_ , P1_U3019 );
nand NAND2_1766 ( P1_U4462 , P1_REG0_REG_16_ , P1_U3020 );
nand NAND2_1767 ( P1_U4463 , P1_ADD_99_U72 , P1_U3017 );
not NOT1_1768 ( P1_U4464 , P1_U3071 );
nand NAND2_1769 ( P1_U4465 , P1_U3033 , P1_U3077 );
nand NAND2_1770 ( P1_U4466 , P1_R1150_U112 , P1_U3994 );
nand NAND2_1771 ( P1_U4467 , P1_R1117_U112 , P1_U3996 );
nand NAND2_1772 ( P1_U4468 , P1_R1138_U112 , P1_U3995 );
nand NAND2_1773 ( P1_U4469 , P1_R1192_U112 , P1_U3992 );
nand NAND2_1774 ( P1_U4470 , P1_R1207_U112 , P1_U3991 );
nand NAND2_1775 ( P1_U4471 , P1_R1171_U112 , P1_U4001 );
nand NAND2_1776 ( P1_U4472 , P1_R1240_U112 , P1_U4000 );
not NOT1_1777 ( P1_U4473 , P1_U3389 );
nand NAND2_1778 ( P1_U4474 , P1_R1222_U112 , P1_U3026 );
nand NAND2_1779 ( P1_U4475 , P1_U3025 , P1_U3071 );
nand NAND2_1780 ( P1_U4476 , P1_R1282_U10 , P1_U3023 );
nand NAND2_1781 ( P1_U4477 , P1_U3498 , P1_U4175 );
nand NAND2_1782 ( P1_U4478 , P1_U3694 , P1_U4473 );
nand NAND2_1783 ( P1_U4479 , P1_REG2_REG_17_ , P1_U3018 );
nand NAND2_1784 ( P1_U4480 , P1_REG1_REG_17_ , P1_U3019 );
nand NAND2_1785 ( P1_U4481 , P1_REG0_REG_17_ , P1_U3020 );
nand NAND2_1786 ( P1_U4482 , P1_ADD_99_U71 , P1_U3017 );
not NOT1_1787 ( P1_U4483 , P1_U3067 );
nand NAND2_1788 ( P1_U4484 , P1_U3033 , P1_U3072 );
nand NAND2_1789 ( P1_U4485 , P1_R1150_U14 , P1_U3994 );
nand NAND2_1790 ( P1_U4486 , P1_R1117_U14 , P1_U3996 );
nand NAND2_1791 ( P1_U4487 , P1_R1138_U111 , P1_U3995 );
nand NAND2_1792 ( P1_U4488 , P1_R1192_U14 , P1_U3992 );
nand NAND2_1793 ( P1_U4489 , P1_R1207_U14 , P1_U3991 );
nand NAND2_1794 ( P1_U4490 , P1_R1171_U111 , P1_U4001 );
nand NAND2_1795 ( P1_U4491 , P1_R1240_U111 , P1_U4000 );
not NOT1_1796 ( P1_U4492 , P1_U3390 );
nand NAND2_1797 ( P1_U4493 , P1_R1222_U111 , P1_U3026 );
nand NAND2_1798 ( P1_U4494 , P1_U3025 , P1_U3067 );
nand NAND2_1799 ( P1_U4495 , P1_R1282_U11 , P1_U3023 );
nand NAND2_1800 ( P1_U4496 , P1_U3501 , P1_U4175 );
nand NAND2_1801 ( P1_U4497 , P1_U3698 , P1_U4492 );
nand NAND2_1802 ( P1_U4498 , P1_REG2_REG_18_ , P1_U3018 );
nand NAND2_1803 ( P1_U4499 , P1_REG1_REG_18_ , P1_U3019 );
nand NAND2_1804 ( P1_U4500 , P1_REG0_REG_18_ , P1_U3020 );
nand NAND2_1805 ( P1_U4501 , P1_ADD_99_U70 , P1_U3017 );
not NOT1_1806 ( P1_U4502 , P1_U3080 );
nand NAND2_1807 ( P1_U4503 , P1_U3033 , P1_U3071 );
nand NAND2_1808 ( P1_U4504 , P1_R1150_U101 , P1_U3994 );
nand NAND2_1809 ( P1_U4505 , P1_R1117_U101 , P1_U3996 );
nand NAND2_1810 ( P1_U4506 , P1_R1138_U13 , P1_U3995 );
nand NAND2_1811 ( P1_U4507 , P1_R1192_U101 , P1_U3992 );
nand NAND2_1812 ( P1_U4508 , P1_R1207_U101 , P1_U3991 );
nand NAND2_1813 ( P1_U4509 , P1_R1171_U13 , P1_U4001 );
nand NAND2_1814 ( P1_U4510 , P1_R1240_U13 , P1_U4000 );
not NOT1_1815 ( P1_U4511 , P1_U3391 );
nand NAND2_1816 ( P1_U4512 , P1_R1222_U13 , P1_U3026 );
nand NAND2_1817 ( P1_U4513 , P1_U3025 , P1_U3080 );
nand NAND2_1818 ( P1_U4514 , P1_R1282_U84 , P1_U3023 );
nand NAND2_1819 ( P1_U4515 , P1_U3504 , P1_U4175 );
nand NAND2_1820 ( P1_U4516 , P1_U3702 , P1_U4511 );
nand NAND2_1821 ( P1_U4517 , P1_REG2_REG_19_ , P1_U3018 );
nand NAND2_1822 ( P1_U4518 , P1_REG1_REG_19_ , P1_U3019 );
nand NAND2_1823 ( P1_U4519 , P1_REG0_REG_19_ , P1_U3020 );
nand NAND2_1824 ( P1_U4520 , P1_ADD_99_U69 , P1_U3017 );
not NOT1_1825 ( P1_U4521 , P1_U3079 );
nand NAND2_1826 ( P1_U4522 , P1_U3033 , P1_U3067 );
nand NAND2_1827 ( P1_U4523 , P1_R1150_U100 , P1_U3994 );
nand NAND2_1828 ( P1_U4524 , P1_R1117_U100 , P1_U3996 );
nand NAND2_1829 ( P1_U4525 , P1_R1138_U110 , P1_U3995 );
nand NAND2_1830 ( P1_U4526 , P1_R1192_U100 , P1_U3992 );
nand NAND2_1831 ( P1_U4527 , P1_R1207_U100 , P1_U3991 );
nand NAND2_1832 ( P1_U4528 , P1_R1171_U110 , P1_U4001 );
nand NAND2_1833 ( P1_U4529 , P1_R1240_U110 , P1_U4000 );
not NOT1_1834 ( P1_U4530 , P1_U3392 );
nand NAND2_1835 ( P1_U4531 , P1_R1222_U110 , P1_U3026 );
nand NAND2_1836 ( P1_U4532 , P1_U3025 , P1_U3079 );
nand NAND2_1837 ( P1_U4533 , P1_R1282_U12 , P1_U3023 );
nand NAND2_1838 ( P1_U4534 , P1_U3507 , P1_U4175 );
nand NAND2_1839 ( P1_U4535 , P1_U3706 , P1_U4530 );
nand NAND2_1840 ( P1_U4536 , P1_REG2_REG_20_ , P1_U3018 );
nand NAND2_1841 ( P1_U4537 , P1_REG1_REG_20_ , P1_U3019 );
nand NAND2_1842 ( P1_U4538 , P1_REG0_REG_20_ , P1_U3020 );
nand NAND2_1843 ( P1_U4539 , P1_ADD_99_U68 , P1_U3017 );
not NOT1_1844 ( P1_U4540 , P1_U3074 );
nand NAND2_1845 ( P1_U4541 , P1_U3033 , P1_U3080 );
nand NAND2_1846 ( P1_U4542 , P1_R1150_U99 , P1_U3994 );
nand NAND2_1847 ( P1_U4543 , P1_R1117_U99 , P1_U3996 );
nand NAND2_1848 ( P1_U4544 , P1_R1138_U109 , P1_U3995 );
nand NAND2_1849 ( P1_U4545 , P1_R1192_U99 , P1_U3992 );
nand NAND2_1850 ( P1_U4546 , P1_R1207_U99 , P1_U3991 );
nand NAND2_1851 ( P1_U4547 , P1_R1171_U109 , P1_U4001 );
nand NAND2_1852 ( P1_U4548 , P1_R1240_U109 , P1_U4000 );
not NOT1_1853 ( P1_U4549 , P1_U3393 );
nand NAND2_1854 ( P1_U4550 , P1_R1222_U109 , P1_U3026 );
nand NAND2_1855 ( P1_U4551 , P1_U3025 , P1_U3074 );
nand NAND2_1856 ( P1_U4552 , P1_R1282_U82 , P1_U3023 );
nand NAND2_1857 ( P1_U4553 , P1_U3509 , P1_U4175 );
nand NAND2_1858 ( P1_U4554 , P1_U3710 , P1_U4549 );
nand NAND2_1859 ( P1_U4555 , P1_REG2_REG_21_ , P1_U3018 );
nand NAND2_1860 ( P1_U4556 , P1_REG1_REG_21_ , P1_U3019 );
nand NAND2_1861 ( P1_U4557 , P1_REG0_REG_21_ , P1_U3020 );
nand NAND2_1862 ( P1_U4558 , P1_ADD_99_U67 , P1_U3017 );
not NOT1_1863 ( P1_U4559 , P1_U3073 );
nand NAND2_1864 ( P1_U4560 , P1_U3033 , P1_U3079 );
nand NAND2_1865 ( P1_U4561 , P1_R1150_U97 , P1_U3994 );
nand NAND2_1866 ( P1_U4562 , P1_R1117_U97 , P1_U3996 );
nand NAND2_1867 ( P1_U4563 , P1_R1138_U14 , P1_U3995 );
nand NAND2_1868 ( P1_U4564 , P1_R1192_U97 , P1_U3992 );
nand NAND2_1869 ( P1_U4565 , P1_R1207_U97 , P1_U3991 );
nand NAND2_1870 ( P1_U4566 , P1_R1171_U14 , P1_U4001 );
nand NAND2_1871 ( P1_U4567 , P1_R1240_U14 , P1_U4000 );
not NOT1_1872 ( P1_U4568 , P1_U3395 );
nand NAND2_1873 ( P1_U4569 , P1_R1222_U14 , P1_U3026 );
nand NAND2_1874 ( P1_U4570 , P1_U3025 , P1_U3073 );
nand NAND2_1875 ( P1_U4571 , P1_R1282_U13 , P1_U3023 );
nand NAND2_1876 ( P1_U4572 , P1_U4015 , P1_U4175 );
nand NAND2_1877 ( P1_U4573 , P1_U3714 , P1_U4568 );
nand NAND2_1878 ( P1_U4574 , P1_REG2_REG_22_ , P1_U3018 );
nand NAND2_1879 ( P1_U4575 , P1_REG1_REG_22_ , P1_U3019 );
nand NAND2_1880 ( P1_U4576 , P1_REG0_REG_22_ , P1_U3020 );
nand NAND2_1881 ( P1_U4577 , P1_ADD_99_U66 , P1_U3017 );
not NOT1_1882 ( P1_U4578 , P1_U3059 );
nand NAND2_1883 ( P1_U4579 , P1_U3033 , P1_U3074 );
nand NAND2_1884 ( P1_U4580 , P1_R1150_U111 , P1_U3994 );
nand NAND2_1885 ( P1_U4581 , P1_R1117_U111 , P1_U3996 );
nand NAND2_1886 ( P1_U4582 , P1_R1138_U15 , P1_U3995 );
nand NAND2_1887 ( P1_U4583 , P1_R1192_U111 , P1_U3992 );
nand NAND2_1888 ( P1_U4584 , P1_R1207_U111 , P1_U3991 );
nand NAND2_1889 ( P1_U4585 , P1_R1171_U15 , P1_U4001 );
nand NAND2_1890 ( P1_U4586 , P1_R1240_U15 , P1_U4000 );
not NOT1_1891 ( P1_U4587 , P1_U3397 );
nand NAND2_1892 ( P1_U4588 , P1_R1222_U15 , P1_U3026 );
nand NAND2_1893 ( P1_U4589 , P1_U3025 , P1_U3059 );
nand NAND2_1894 ( P1_U4590 , P1_R1282_U78 , P1_U3023 );
nand NAND2_1895 ( P1_U4591 , P1_U4014 , P1_U4175 );
nand NAND2_1896 ( P1_U4592 , P1_U3718 , P1_U4587 );
nand NAND2_1897 ( P1_U4593 , P1_REG2_REG_23_ , P1_U3018 );
nand NAND2_1898 ( P1_U4594 , P1_REG1_REG_23_ , P1_U3019 );
nand NAND2_1899 ( P1_U4595 , P1_REG0_REG_23_ , P1_U3020 );
nand NAND2_1900 ( P1_U4596 , P1_ADD_99_U65 , P1_U3017 );
not NOT1_1901 ( P1_U4597 , P1_U3064 );
nand NAND2_1902 ( P1_U4598 , P1_U3033 , P1_U3073 );
nand NAND2_1903 ( P1_U4599 , P1_R1150_U110 , P1_U3994 );
nand NAND2_1904 ( P1_U4600 , P1_R1117_U110 , P1_U3996 );
nand NAND2_1905 ( P1_U4601 , P1_R1138_U108 , P1_U3995 );
nand NAND2_1906 ( P1_U4602 , P1_R1192_U110 , P1_U3992 );
nand NAND2_1907 ( P1_U4603 , P1_R1207_U110 , P1_U3991 );
nand NAND2_1908 ( P1_U4604 , P1_R1171_U108 , P1_U4001 );
nand NAND2_1909 ( P1_U4605 , P1_R1240_U108 , P1_U4000 );
not NOT1_1910 ( P1_U4606 , P1_U3399 );
nand NAND2_1911 ( P1_U4607 , P1_R1222_U108 , P1_U3026 );
nand NAND2_1912 ( P1_U4608 , P1_U3025 , P1_U3064 );
nand NAND2_1913 ( P1_U4609 , P1_R1282_U14 , P1_U3023 );
nand NAND2_1914 ( P1_U4610 , P1_U4013 , P1_U4175 );
nand NAND2_1915 ( P1_U4611 , P1_U3722 , P1_U4606 );
nand NAND2_1916 ( P1_U4612 , P1_REG2_REG_24_ , P1_U3018 );
nand NAND2_1917 ( P1_U4613 , P1_REG1_REG_24_ , P1_U3019 );
nand NAND2_1918 ( P1_U4614 , P1_REG0_REG_24_ , P1_U3020 );
nand NAND2_1919 ( P1_U4615 , P1_ADD_99_U64 , P1_U3017 );
not NOT1_1920 ( P1_U4616 , P1_U3063 );
nand NAND2_1921 ( P1_U4617 , P1_U3033 , P1_U3059 );
nand NAND2_1922 ( P1_U4618 , P1_R1150_U15 , P1_U3994 );
nand NAND2_1923 ( P1_U4619 , P1_R1117_U15 , P1_U3996 );
nand NAND2_1924 ( P1_U4620 , P1_R1138_U107 , P1_U3995 );
nand NAND2_1925 ( P1_U4621 , P1_R1192_U15 , P1_U3992 );
nand NAND2_1926 ( P1_U4622 , P1_R1207_U15 , P1_U3991 );
nand NAND2_1927 ( P1_U4623 , P1_R1171_U107 , P1_U4001 );
nand NAND2_1928 ( P1_U4624 , P1_R1240_U107 , P1_U4000 );
not NOT1_1929 ( P1_U4625 , P1_U3401 );
nand NAND2_1930 ( P1_U4626 , P1_R1222_U107 , P1_U3026 );
nand NAND2_1931 ( P1_U4627 , P1_U3025 , P1_U3063 );
nand NAND2_1932 ( P1_U4628 , P1_R1282_U76 , P1_U3023 );
nand NAND2_1933 ( P1_U4629 , P1_U4012 , P1_U4175 );
nand NAND2_1934 ( P1_U4630 , P1_U3726 , P1_U4625 );
nand NAND2_1935 ( P1_U4631 , P1_REG2_REG_25_ , P1_U3018 );
nand NAND2_1936 ( P1_U4632 , P1_REG1_REG_25_ , P1_U3019 );
nand NAND2_1937 ( P1_U4633 , P1_REG0_REG_25_ , P1_U3020 );
nand NAND2_1938 ( P1_U4634 , P1_ADD_99_U63 , P1_U3017 );
not NOT1_1939 ( P1_U4635 , P1_U3056 );
nand NAND2_1940 ( P1_U4636 , P1_U3033 , P1_U3064 );
nand NAND2_1941 ( P1_U4637 , P1_R1150_U96 , P1_U3994 );
nand NAND2_1942 ( P1_U4638 , P1_R1117_U96 , P1_U3996 );
nand NAND2_1943 ( P1_U4639 , P1_R1138_U106 , P1_U3995 );
nand NAND2_1944 ( P1_U4640 , P1_R1192_U96 , P1_U3992 );
nand NAND2_1945 ( P1_U4641 , P1_R1207_U96 , P1_U3991 );
nand NAND2_1946 ( P1_U4642 , P1_R1171_U106 , P1_U4001 );
nand NAND2_1947 ( P1_U4643 , P1_R1240_U106 , P1_U4000 );
not NOT1_1948 ( P1_U4644 , P1_U3403 );
nand NAND2_1949 ( P1_U4645 , P1_R1222_U106 , P1_U3026 );
nand NAND2_1950 ( P1_U4646 , P1_U3025 , P1_U3056 );
nand NAND2_1951 ( P1_U4647 , P1_R1282_U15 , P1_U3023 );
nand NAND2_1952 ( P1_U4648 , P1_U4011 , P1_U4175 );
nand NAND2_1953 ( P1_U4649 , P1_U3730 , P1_U4644 );
nand NAND2_1954 ( P1_U4650 , P1_REG2_REG_26_ , P1_U3018 );
nand NAND2_1955 ( P1_U4651 , P1_REG1_REG_26_ , P1_U3019 );
nand NAND2_1956 ( P1_U4652 , P1_REG0_REG_26_ , P1_U3020 );
nand NAND2_1957 ( P1_U4653 , P1_ADD_99_U62 , P1_U3017 );
not NOT1_1958 ( P1_U4654 , P1_U3055 );
nand NAND2_1959 ( P1_U4655 , P1_U3033 , P1_U3063 );
nand NAND2_1960 ( P1_U4656 , P1_R1150_U95 , P1_U3994 );
nand NAND2_1961 ( P1_U4657 , P1_R1117_U95 , P1_U3996 );
nand NAND2_1962 ( P1_U4658 , P1_R1138_U105 , P1_U3995 );
nand NAND2_1963 ( P1_U4659 , P1_R1192_U95 , P1_U3992 );
nand NAND2_1964 ( P1_U4660 , P1_R1207_U95 , P1_U3991 );
nand NAND2_1965 ( P1_U4661 , P1_R1171_U105 , P1_U4001 );
nand NAND2_1966 ( P1_U4662 , P1_R1240_U105 , P1_U4000 );
not NOT1_1967 ( P1_U4663 , P1_U3405 );
nand NAND2_1968 ( P1_U4664 , P1_R1222_U105 , P1_U3026 );
nand NAND2_1969 ( P1_U4665 , P1_U3025 , P1_U3055 );
nand NAND2_1970 ( P1_U4666 , P1_R1282_U74 , P1_U3023 );
nand NAND2_1971 ( P1_U4667 , P1_U4010 , P1_U4175 );
nand NAND2_1972 ( P1_U4668 , P1_U3734 , P1_U4663 );
nand NAND2_1973 ( P1_U4669 , P1_REG2_REG_27_ , P1_U3018 );
nand NAND2_1974 ( P1_U4670 , P1_REG1_REG_27_ , P1_U3019 );
nand NAND2_1975 ( P1_U4671 , P1_REG0_REG_27_ , P1_U3020 );
nand NAND2_1976 ( P1_U4672 , P1_ADD_99_U61 , P1_U3017 );
not NOT1_1977 ( P1_U4673 , P1_U3051 );
nand NAND2_1978 ( P1_U4674 , P1_U3033 , P1_U3056 );
nand NAND2_1979 ( P1_U4675 , P1_R1150_U109 , P1_U3994 );
nand NAND2_1980 ( P1_U4676 , P1_R1117_U109 , P1_U3996 );
nand NAND2_1981 ( P1_U4677 , P1_R1138_U16 , P1_U3995 );
nand NAND2_1982 ( P1_U4678 , P1_R1192_U109 , P1_U3992 );
nand NAND2_1983 ( P1_U4679 , P1_R1207_U109 , P1_U3991 );
nand NAND2_1984 ( P1_U4680 , P1_R1171_U16 , P1_U4001 );
nand NAND2_1985 ( P1_U4681 , P1_R1240_U16 , P1_U4000 );
not NOT1_1986 ( P1_U4682 , P1_U3407 );
nand NAND2_1987 ( P1_U4683 , P1_R1222_U16 , P1_U3026 );
nand NAND2_1988 ( P1_U4684 , P1_U3025 , P1_U3051 );
nand NAND2_1989 ( P1_U4685 , P1_R1282_U16 , P1_U3023 );
nand NAND2_1990 ( P1_U4686 , P1_U4009 , P1_U4175 );
nand NAND2_1991 ( P1_U4687 , P1_U3738 , P1_U4682 );
nand NAND2_1992 ( P1_U4688 , P1_REG2_REG_28_ , P1_U3018 );
nand NAND2_1993 ( P1_U4689 , P1_REG1_REG_28_ , P1_U3019 );
nand NAND2_1994 ( P1_U4690 , P1_REG0_REG_28_ , P1_U3020 );
nand NAND2_1995 ( P1_U4691 , P1_ADD_99_U60 , P1_U3017 );
not NOT1_1996 ( P1_U4692 , P1_U3052 );
nand NAND2_1997 ( P1_U4693 , P1_U3033 , P1_U3055 );
nand NAND2_1998 ( P1_U4694 , P1_R1150_U16 , P1_U3994 );
nand NAND2_1999 ( P1_U4695 , P1_R1117_U16 , P1_U3996 );
nand NAND2_2000 ( P1_U4696 , P1_R1138_U104 , P1_U3995 );
nand NAND2_2001 ( P1_U4697 , P1_R1192_U16 , P1_U3992 );
nand NAND2_2002 ( P1_U4698 , P1_R1207_U16 , P1_U3991 );
nand NAND2_2003 ( P1_U4699 , P1_R1171_U104 , P1_U4001 );
nand NAND2_2004 ( P1_U4700 , P1_R1240_U104 , P1_U4000 );
not NOT1_2005 ( P1_U4701 , P1_U3409 );
nand NAND2_2006 ( P1_U4702 , P1_R1222_U104 , P1_U3026 );
nand NAND2_2007 ( P1_U4703 , P1_U3025 , P1_U3052 );
nand NAND2_2008 ( P1_U4704 , P1_R1282_U72 , P1_U3023 );
nand NAND2_2009 ( P1_U4705 , P1_U4008 , P1_U4175 );
nand NAND2_2010 ( P1_U4706 , P1_U3742 , P1_U4701 );
nand NAND2_2011 ( P1_U4707 , P1_ADD_99_U5 , P1_U3017 );
nand NAND2_2012 ( P1_U4708 , P1_REG2_REG_29_ , P1_U3018 );
nand NAND2_2013 ( P1_U4709 , P1_REG1_REG_29_ , P1_U3019 );
nand NAND2_2014 ( P1_U4710 , P1_REG0_REG_29_ , P1_U3020 );
not NOT1_2015 ( P1_U4711 , P1_U3053 );
nand NAND2_2016 ( P1_U4712 , P1_U3033 , P1_U3051 );
nand NAND2_2017 ( P1_U4713 , P1_R1150_U94 , P1_U3994 );
nand NAND2_2018 ( P1_U4714 , P1_R1117_U94 , P1_U3996 );
nand NAND2_2019 ( P1_U4715 , P1_R1138_U103 , P1_U3995 );
nand NAND2_2020 ( P1_U4716 , P1_R1192_U94 , P1_U3992 );
nand NAND2_2021 ( P1_U4717 , P1_R1207_U94 , P1_U3991 );
nand NAND2_2022 ( P1_U4718 , P1_R1171_U103 , P1_U4001 );
nand NAND2_2023 ( P1_U4719 , P1_R1240_U103 , P1_U4000 );
not NOT1_2024 ( P1_U4720 , P1_U3411 );
nand NAND2_2025 ( P1_U4721 , P1_R1222_U103 , P1_U3026 );
nand NAND2_2026 ( P1_U4722 , P1_U3025 , P1_U3053 );
nand NAND2_2027 ( P1_U4723 , P1_R1282_U17 , P1_U3023 );
nand NAND2_2028 ( P1_U4724 , P1_U4007 , P1_U4175 );
nand NAND2_2029 ( P1_U4725 , P1_U3746 , P1_U4720 );
nand NAND2_2030 ( P1_U4726 , P1_REG2_REG_30_ , P1_U3018 );
nand NAND2_2031 ( P1_U4727 , P1_REG1_REG_30_ , P1_U3019 );
nand NAND2_2032 ( P1_U4728 , P1_REG0_REG_30_ , P1_U3020 );
not NOT1_2033 ( P1_U4729 , P1_U3057 );
nand NAND2_2034 ( P1_U4730 , P1_U5728 , P1_U3358 );
nand NAND2_2035 ( P1_U4731 , P1_U3946 , P1_U4730 );
nand NAND2_2036 ( P1_U4732 , P1_U3747 , P1_U3057 );
nand NAND2_2037 ( P1_U4733 , P1_U3033 , P1_U3052 );
nand NAND2_2038 ( P1_U4734 , P1_R1150_U17 , P1_U3994 );
nand NAND2_2039 ( P1_U4735 , P1_R1117_U17 , P1_U3996 );
nand NAND2_2040 ( P1_U4736 , P1_R1138_U102 , P1_U3995 );
nand NAND2_2041 ( P1_U4737 , P1_R1192_U17 , P1_U3992 );
nand NAND2_2042 ( P1_U4738 , P1_R1207_U17 , P1_U3991 );
nand NAND2_2043 ( P1_U4739 , P1_R1171_U102 , P1_U4001 );
nand NAND2_2044 ( P1_U4740 , P1_R1240_U102 , P1_U4000 );
not NOT1_2045 ( P1_U4741 , P1_U3413 );
nand NAND2_2046 ( P1_U4742 , P1_R1222_U102 , P1_U3026 );
nand NAND2_2047 ( P1_U4743 , P1_R1282_U70 , P1_U3023 );
nand NAND2_2048 ( P1_U4744 , P1_U4018 , P1_U4175 );
nand NAND2_2049 ( P1_U4745 , P1_U3751 , P1_U4741 );
nand NAND2_2050 ( P1_U4746 , P1_REG2_REG_31_ , P1_U3018 );
nand NAND2_2051 ( P1_U4747 , P1_REG1_REG_31_ , P1_U3019 );
nand NAND2_2052 ( P1_U4748 , P1_REG0_REG_31_ , P1_U3020 );
not NOT1_2053 ( P1_U4749 , P1_U3054 );
nand NAND2_2054 ( P1_U4750 , P1_R1282_U19 , P1_U3023 );
nand NAND2_2055 ( P1_U4751 , P1_U4017 , P1_U4175 );
nand NAND3_2056 ( P1_U4752 , P1_U4751 , P1_U3979 , P1_U4750 );
nand NAND2_2057 ( P1_U4753 , P1_R1282_U68 , P1_U3023 );
nand NAND2_2058 ( P1_U4754 , P1_U4016 , P1_U4175 );
nand NAND3_2059 ( P1_U4755 , P1_U4754 , P1_U3979 , P1_U4753 );
nand NAND2_2060 ( P1_U4756 , P1_U3754 , P1_U3016 );
nand NAND2_2061 ( P1_U4757 , P1_U3418 , P1_U4756 );
nand NAND2_2062 ( P1_U4758 , P1_U4021 , P1_U3442 );
not NOT1_2063 ( P1_U4759 , P1_U3422 );
nand NAND2_2064 ( P1_U4760 , P1_U3035 , P1_U3076 );
nand NAND2_2065 ( P1_U4761 , P1_U3032 , P1_REG3_REG_0_ );
nand NAND2_2066 ( P1_U4762 , P1_U3031 , P1_R1222_U96 );
nand NAND2_2067 ( P1_U4763 , P1_U3030 , P1_U3451 );
nand NAND2_2068 ( P1_U4764 , P1_U3029 , P1_U3451 );
nand NAND2_2069 ( P1_U4765 , P1_U3035 , P1_U3066 );
nand NAND2_2070 ( P1_U4766 , P1_U3032 , P1_REG3_REG_1_ );
nand NAND2_2071 ( P1_U4767 , P1_U3031 , P1_R1222_U95 );
nand NAND2_2072 ( P1_U4768 , P1_U3030 , P1_U3456 );
nand NAND2_2073 ( P1_U4769 , P1_U3029 , P1_R1282_U57 );
nand NAND2_2074 ( P1_U4770 , P1_U3035 , P1_U3062 );
nand NAND2_2075 ( P1_U4771 , P1_U3032 , P1_REG3_REG_2_ );
nand NAND2_2076 ( P1_U4772 , P1_U3031 , P1_R1222_U17 );
nand NAND2_2077 ( P1_U4773 , P1_U3030 , P1_U3459 );
nand NAND2_2078 ( P1_U4774 , P1_U3029 , P1_R1282_U18 );
nand NAND2_2079 ( P1_U4775 , P1_U3035 , P1_U3058 );
nand NAND2_2080 ( P1_U4776 , P1_U3032 , P1_ADD_99_U4 );
nand NAND2_2081 ( P1_U4777 , P1_U3031 , P1_R1222_U101 );
nand NAND2_2082 ( P1_U4778 , P1_U3030 , P1_U3462 );
nand NAND2_2083 ( P1_U4779 , P1_U3029 , P1_R1282_U20 );
nand NAND2_2084 ( P1_U4780 , P1_U3035 , P1_U3065 );
nand NAND2_2085 ( P1_U4781 , P1_U3032 , P1_ADD_99_U59 );
nand NAND2_2086 ( P1_U4782 , P1_U3031 , P1_R1222_U100 );
nand NAND2_2087 ( P1_U4783 , P1_U3030 , P1_U3465 );
nand NAND2_2088 ( P1_U4784 , P1_U3029 , P1_R1282_U21 );
nand NAND2_2089 ( P1_U4785 , P1_U3035 , P1_U3069 );
nand NAND2_2090 ( P1_U4786 , P1_U3032 , P1_ADD_99_U58 );
nand NAND2_2091 ( P1_U4787 , P1_U3031 , P1_R1222_U18 );
nand NAND2_2092 ( P1_U4788 , P1_U3030 , P1_U3468 );
nand NAND2_2093 ( P1_U4789 , P1_U3029 , P1_R1282_U65 );
nand NAND2_2094 ( P1_U4790 , P1_U3035 , P1_U3068 );
nand NAND2_2095 ( P1_U4791 , P1_U3032 , P1_ADD_99_U57 );
nand NAND2_2096 ( P1_U4792 , P1_U3031 , P1_R1222_U99 );
nand NAND2_2097 ( P1_U4793 , P1_U3030 , P1_U3471 );
nand NAND2_2098 ( P1_U4794 , P1_U3029 , P1_R1282_U22 );
nand NAND2_2099 ( P1_U4795 , P1_U3035 , P1_U3082 );
nand NAND2_2100 ( P1_U4796 , P1_U3032 , P1_ADD_99_U56 );
nand NAND2_2101 ( P1_U4797 , P1_U3031 , P1_R1222_U19 );
nand NAND2_2102 ( P1_U4798 , P1_U3030 , P1_U3474 );
nand NAND2_2103 ( P1_U4799 , P1_U3029 , P1_R1282_U23 );
nand NAND2_2104 ( P1_U4800 , P1_U3035 , P1_U3081 );
nand NAND2_2105 ( P1_U4801 , P1_U3032 , P1_ADD_99_U55 );
nand NAND2_2106 ( P1_U4802 , P1_U3031 , P1_R1222_U98 );
nand NAND2_2107 ( P1_U4803 , P1_U3030 , P1_U3477 );
nand NAND2_2108 ( P1_U4804 , P1_U3029 , P1_R1282_U24 );
nand NAND2_2109 ( P1_U4805 , P1_U3035 , P1_U3060 );
nand NAND2_2110 ( P1_U4806 , P1_U3032 , P1_ADD_99_U54 );
nand NAND2_2111 ( P1_U4807 , P1_U3031 , P1_R1222_U97 );
nand NAND2_2112 ( P1_U4808 , P1_U3030 , P1_U3480 );
nand NAND2_2113 ( P1_U4809 , P1_U3029 , P1_R1282_U63 );
nand NAND2_2114 ( P1_U4810 , P1_U3035 , P1_U3061 );
nand NAND2_2115 ( P1_U4811 , P1_U3032 , P1_ADD_99_U78 );
nand NAND2_2116 ( P1_U4812 , P1_U3031 , P1_R1222_U11 );
nand NAND2_2117 ( P1_U4813 , P1_U3030 , P1_U3483 );
nand NAND2_2118 ( P1_U4814 , P1_U3029 , P1_R1282_U6 );
nand NAND2_2119 ( P1_U4815 , P1_U3035 , P1_U3070 );
nand NAND2_2120 ( P1_U4816 , P1_U3032 , P1_ADD_99_U77 );
nand NAND2_2121 ( P1_U4817 , P1_U3031 , P1_R1222_U115 );
nand NAND2_2122 ( P1_U4818 , P1_U3030 , P1_U3486 );
nand NAND2_2123 ( P1_U4819 , P1_U3029 , P1_R1282_U7 );
nand NAND2_2124 ( P1_U4820 , P1_U3035 , P1_U3078 );
nand NAND2_2125 ( P1_U4821 , P1_U3032 , P1_ADD_99_U76 );
nand NAND2_2126 ( P1_U4822 , P1_U3031 , P1_R1222_U114 );
nand NAND2_2127 ( P1_U4823 , P1_U3030 , P1_U3489 );
nand NAND2_2128 ( P1_U4824 , P1_U3029 , P1_R1282_U8 );
nand NAND2_2129 ( P1_U4825 , P1_U3035 , P1_U3077 );
nand NAND2_2130 ( P1_U4826 , P1_U3032 , P1_ADD_99_U75 );
nand NAND2_2131 ( P1_U4827 , P1_U3031 , P1_R1222_U12 );
nand NAND2_2132 ( P1_U4828 , P1_U3030 , P1_U3492 );
nand NAND2_2133 ( P1_U4829 , P1_U3029 , P1_R1282_U86 );
nand NAND2_2134 ( P1_U4830 , P1_U3035 , P1_U3072 );
nand NAND2_2135 ( P1_U4831 , P1_U3032 , P1_ADD_99_U74 );
nand NAND2_2136 ( P1_U4832 , P1_U3031 , P1_R1222_U113 );
nand NAND2_2137 ( P1_U4833 , P1_U3030 , P1_U3495 );
nand NAND2_2138 ( P1_U4834 , P1_U3029 , P1_R1282_U9 );
nand NAND2_2139 ( P1_U4835 , P1_U3035 , P1_U3071 );
nand NAND2_2140 ( P1_U4836 , P1_U3032 , P1_ADD_99_U73 );
nand NAND2_2141 ( P1_U4837 , P1_U3031 , P1_R1222_U112 );
nand NAND2_2142 ( P1_U4838 , P1_U3030 , P1_U3498 );
nand NAND2_2143 ( P1_U4839 , P1_U3029 , P1_R1282_U10 );
nand NAND2_2144 ( P1_U4840 , P1_U3035 , P1_U3067 );
nand NAND2_2145 ( P1_U4841 , P1_U3032 , P1_ADD_99_U72 );
nand NAND2_2146 ( P1_U4842 , P1_U3031 , P1_R1222_U111 );
nand NAND2_2147 ( P1_U4843 , P1_U3030 , P1_U3501 );
nand NAND2_2148 ( P1_U4844 , P1_U3029 , P1_R1282_U11 );
nand NAND2_2149 ( P1_U4845 , P1_U3035 , P1_U3080 );
nand NAND2_2150 ( P1_U4846 , P1_U3032 , P1_ADD_99_U71 );
nand NAND2_2151 ( P1_U4847 , P1_U3031 , P1_R1222_U13 );
nand NAND2_2152 ( P1_U4848 , P1_U3030 , P1_U3504 );
nand NAND2_2153 ( P1_U4849 , P1_U3029 , P1_R1282_U84 );
nand NAND2_2154 ( P1_U4850 , P1_U3035 , P1_U3079 );
nand NAND2_2155 ( P1_U4851 , P1_U3032 , P1_ADD_99_U70 );
nand NAND2_2156 ( P1_U4852 , P1_U3031 , P1_R1222_U110 );
nand NAND2_2157 ( P1_U4853 , P1_U3030 , P1_U3507 );
nand NAND2_2158 ( P1_U4854 , P1_U3029 , P1_R1282_U12 );
nand NAND2_2159 ( P1_U4855 , P1_U3035 , P1_U3074 );
nand NAND2_2160 ( P1_U4856 , P1_U3032 , P1_ADD_99_U69 );
nand NAND2_2161 ( P1_U4857 , P1_U3031 , P1_R1222_U109 );
nand NAND2_2162 ( P1_U4858 , P1_U3030 , P1_U3509 );
nand NAND2_2163 ( P1_U4859 , P1_U3029 , P1_R1282_U82 );
nand NAND2_2164 ( P1_U4860 , P1_U3035 , P1_U3073 );
nand NAND2_2165 ( P1_U4861 , P1_U3032 , P1_ADD_99_U68 );
nand NAND2_2166 ( P1_U4862 , P1_U3031 , P1_R1222_U14 );
nand NAND2_2167 ( P1_U4863 , P1_U3030 , P1_U4015 );
nand NAND2_2168 ( P1_U4864 , P1_U3029 , P1_R1282_U13 );
nand NAND2_2169 ( P1_U4865 , P1_U3035 , P1_U3059 );
nand NAND2_2170 ( P1_U4866 , P1_U3032 , P1_ADD_99_U67 );
nand NAND2_2171 ( P1_U4867 , P1_U3031 , P1_R1222_U15 );
nand NAND2_2172 ( P1_U4868 , P1_U3030 , P1_U4014 );
nand NAND2_2173 ( P1_U4869 , P1_U3029 , P1_R1282_U78 );
nand NAND2_2174 ( P1_U4870 , P1_U3035 , P1_U3064 );
nand NAND2_2175 ( P1_U4871 , P1_U3032 , P1_ADD_99_U66 );
nand NAND2_2176 ( P1_U4872 , P1_U3031 , P1_R1222_U108 );
nand NAND2_2177 ( P1_U4873 , P1_U3030 , P1_U4013 );
nand NAND2_2178 ( P1_U4874 , P1_U3029 , P1_R1282_U14 );
nand NAND2_2179 ( P1_U4875 , P1_U3035 , P1_U3063 );
nand NAND2_2180 ( P1_U4876 , P1_U3032 , P1_ADD_99_U65 );
nand NAND2_2181 ( P1_U4877 , P1_U3031 , P1_R1222_U107 );
nand NAND2_2182 ( P1_U4878 , P1_U3030 , P1_U4012 );
nand NAND2_2183 ( P1_U4879 , P1_U3029 , P1_R1282_U76 );
nand NAND2_2184 ( P1_U4880 , P1_U3035 , P1_U3056 );
nand NAND2_2185 ( P1_U4881 , P1_U3032 , P1_ADD_99_U64 );
nand NAND2_2186 ( P1_U4882 , P1_U3031 , P1_R1222_U106 );
nand NAND2_2187 ( P1_U4883 , P1_U3030 , P1_U4011 );
nand NAND2_2188 ( P1_U4884 , P1_U3029 , P1_R1282_U15 );
nand NAND2_2189 ( P1_U4885 , P1_U3035 , P1_U3055 );
nand NAND2_2190 ( P1_U4886 , P1_U3032 , P1_ADD_99_U63 );
nand NAND2_2191 ( P1_U4887 , P1_U3031 , P1_R1222_U105 );
nand NAND2_2192 ( P1_U4888 , P1_U3030 , P1_U4010 );
nand NAND2_2193 ( P1_U4889 , P1_U3029 , P1_R1282_U74 );
nand NAND2_2194 ( P1_U4890 , P1_U3035 , P1_U3051 );
nand NAND2_2195 ( P1_U4891 , P1_U3032 , P1_ADD_99_U62 );
nand NAND2_2196 ( P1_U4892 , P1_U3031 , P1_R1222_U16 );
nand NAND2_2197 ( P1_U4893 , P1_U3030 , P1_U4009 );
nand NAND2_2198 ( P1_U4894 , P1_U3029 , P1_R1282_U16 );
nand NAND2_2199 ( P1_U4895 , P1_U3035 , P1_U3052 );
nand NAND2_2200 ( P1_U4896 , P1_U3032 , P1_ADD_99_U61 );
nand NAND2_2201 ( P1_U4897 , P1_U3031 , P1_R1222_U104 );
nand NAND2_2202 ( P1_U4898 , P1_U3030 , P1_U4008 );
nand NAND2_2203 ( P1_U4899 , P1_U3029 , P1_R1282_U72 );
nand NAND2_2204 ( P1_U4900 , P1_U3035 , P1_U3053 );
nand NAND2_2205 ( P1_U4901 , P1_U3032 , P1_ADD_99_U60 );
nand NAND2_2206 ( P1_U4902 , P1_U3031 , P1_R1222_U103 );
nand NAND2_2207 ( P1_U4903 , P1_U3030 , P1_U4007 );
nand NAND2_2208 ( P1_U4904 , P1_U3029 , P1_R1282_U17 );
nand NAND2_2209 ( P1_U4905 , P1_U3032 , P1_ADD_99_U5 );
nand NAND2_2210 ( P1_U4906 , P1_U3031 , P1_R1222_U102 );
nand NAND2_2211 ( P1_U4907 , P1_U3030 , P1_U4018 );
nand NAND2_2212 ( P1_U4908 , P1_U3029 , P1_R1282_U70 );
nand NAND2_2213 ( P1_U4909 , P1_U3030 , P1_U4017 );
nand NAND2_2214 ( P1_U4910 , P1_U3029 , P1_R1282_U19 );
nand NAND2_2215 ( P1_U4911 , P1_U3030 , P1_U4016 );
nand NAND2_2216 ( P1_U4912 , P1_U3029 , P1_R1282_U68 );
nand NAND5_2217 ( P1_U4913 , P1_U3814 , P1_U3813 , P1_U3816 , P1_U4759 , P1_U3418 );
nand NAND2_2218 ( P1_U4914 , P1_R1105_U13 , P1_U3041 );
nand NAND2_2219 ( P1_U4915 , P1_U3039 , P1_U3443 );
nand NAND2_2220 ( P1_U4916 , P1_R1162_U13 , P1_U3037 );
nand NAND3_2221 ( P1_U4917 , P1_U4915 , P1_U4914 , P1_U4916 );
nand NAND2_2222 ( P1_U4918 , P1_U3046 , P1_U3372 );
nand NAND2_2223 ( P1_U4919 , P1_U5703 , P1_U4918 );
nand NAND2_2224 ( P1_U4920 , P1_U4919 , P1_U3946 );
not NOT1_2225 ( P1_U4921 , P1_U3083 );
not NOT1_2226 ( P1_U4922 , P1_U3423 );
nand NAND2_2227 ( P1_U4923 , P1_U3043 , P1_U4917 );
nand NAND2_2228 ( P1_U4924 , P1_U3042 , P1_R1105_U13 );
nand NAND2_2229 ( P1_U4925 , P1_REG3_REG_19_ , P1_U3084 );
nand NAND2_2230 ( P1_U4926 , P1_U3040 , P1_U3443 );
nand NAND2_2231 ( P1_U4927 , P1_U3038 , P1_R1162_U13 );
nand NAND2_2232 ( P1_U4928 , P1_ADDR_REG_19_ , P1_U4922 );
nand NAND2_2233 ( P1_U4929 , P1_R1105_U75 , P1_U3041 );
nand NAND2_2234 ( P1_U4930 , P1_U3039 , P1_U3506 );
nand NAND2_2235 ( P1_U4931 , P1_R1162_U75 , P1_U3037 );
nand NAND3_2236 ( P1_U4932 , P1_U4930 , P1_U4929 , P1_U4931 );
nand NAND2_2237 ( P1_U4933 , P1_U3043 , P1_U4932 );
nand NAND2_2238 ( P1_U4934 , P1_R1105_U75 , P1_U3042 );
nand NAND2_2239 ( P1_U4935 , P1_REG3_REG_18_ , P1_U3084 );
nand NAND2_2240 ( P1_U4936 , P1_U3040 , P1_U3506 );
nand NAND2_2241 ( P1_U4937 , P1_R1162_U75 , P1_U3038 );
nand NAND2_2242 ( P1_U4938 , P1_ADDR_REG_18_ , P1_U4922 );
nand NAND2_2243 ( P1_U4939 , P1_R1105_U12 , P1_U3041 );
nand NAND2_2244 ( P1_U4940 , P1_U3039 , P1_U3503 );
nand NAND2_2245 ( P1_U4941 , P1_R1162_U12 , P1_U3037 );
nand NAND3_2246 ( P1_U4942 , P1_U4940 , P1_U4939 , P1_U4941 );
nand NAND2_2247 ( P1_U4943 , P1_U3043 , P1_U4942 );
nand NAND2_2248 ( P1_U4944 , P1_R1105_U12 , P1_U3042 );
nand NAND2_2249 ( P1_U4945 , P1_REG3_REG_17_ , P1_U3084 );
nand NAND2_2250 ( P1_U4946 , P1_U3040 , P1_U3503 );
nand NAND2_2251 ( P1_U4947 , P1_R1162_U12 , P1_U3038 );
nand NAND2_2252 ( P1_U4948 , P1_ADDR_REG_17_ , P1_U4922 );
nand NAND2_2253 ( P1_U4949 , P1_R1105_U76 , P1_U3041 );
nand NAND2_2254 ( P1_U4950 , P1_U3039 , P1_U3500 );
nand NAND2_2255 ( P1_U4951 , P1_R1162_U76 , P1_U3037 );
nand NAND3_2256 ( P1_U4952 , P1_U4950 , P1_U4949 , P1_U4951 );
nand NAND2_2257 ( P1_U4953 , P1_U3043 , P1_U4952 );
nand NAND2_2258 ( P1_U4954 , P1_R1105_U76 , P1_U3042 );
nand NAND2_2259 ( P1_U4955 , P1_REG3_REG_16_ , P1_U3084 );
nand NAND2_2260 ( P1_U4956 , P1_U3040 , P1_U3500 );
nand NAND2_2261 ( P1_U4957 , P1_R1162_U76 , P1_U3038 );
nand NAND2_2262 ( P1_U4958 , P1_ADDR_REG_16_ , P1_U4922 );
nand NAND2_2263 ( P1_U4959 , P1_R1105_U77 , P1_U3041 );
nand NAND2_2264 ( P1_U4960 , P1_U3039 , P1_U3497 );
nand NAND2_2265 ( P1_U4961 , P1_R1162_U77 , P1_U3037 );
nand NAND3_2266 ( P1_U4962 , P1_U4960 , P1_U4959 , P1_U4961 );
nand NAND2_2267 ( P1_U4963 , P1_U3043 , P1_U4962 );
nand NAND2_2268 ( P1_U4964 , P1_R1105_U77 , P1_U3042 );
nand NAND2_2269 ( P1_U4965 , P1_REG3_REG_15_ , P1_U3084 );
nand NAND2_2270 ( P1_U4966 , P1_U3040 , P1_U3497 );
nand NAND2_2271 ( P1_U4967 , P1_R1162_U77 , P1_U3038 );
nand NAND2_2272 ( P1_U4968 , P1_ADDR_REG_15_ , P1_U4922 );
nand NAND2_2273 ( P1_U4969 , P1_R1105_U78 , P1_U3041 );
nand NAND2_2274 ( P1_U4970 , P1_U3039 , P1_U3494 );
nand NAND2_2275 ( P1_U4971 , P1_R1162_U78 , P1_U3037 );
nand NAND3_2276 ( P1_U4972 , P1_U4970 , P1_U4969 , P1_U4971 );
nand NAND2_2277 ( P1_U4973 , P1_U3043 , P1_U4972 );
nand NAND2_2278 ( P1_U4974 , P1_R1105_U78 , P1_U3042 );
nand NAND2_2279 ( P1_U4975 , P1_REG3_REG_14_ , P1_U3084 );
nand NAND2_2280 ( P1_U4976 , P1_U3040 , P1_U3494 );
nand NAND2_2281 ( P1_U4977 , P1_R1162_U78 , P1_U3038 );
nand NAND2_2282 ( P1_U4978 , P1_ADDR_REG_14_ , P1_U4922 );
nand NAND2_2283 ( P1_U4979 , P1_R1105_U11 , P1_U3041 );
nand NAND2_2284 ( P1_U4980 , P1_U3039 , P1_U3491 );
nand NAND2_2285 ( P1_U4981 , P1_R1162_U11 , P1_U3037 );
nand NAND3_2286 ( P1_U4982 , P1_U4980 , P1_U4979 , P1_U4981 );
nand NAND2_2287 ( P1_U4983 , P1_U3043 , P1_U4982 );
nand NAND2_2288 ( P1_U4984 , P1_R1105_U11 , P1_U3042 );
nand NAND2_2289 ( P1_U4985 , P1_REG3_REG_13_ , P1_U3084 );
nand NAND2_2290 ( P1_U4986 , P1_U3040 , P1_U3491 );
nand NAND2_2291 ( P1_U4987 , P1_R1162_U11 , P1_U3038 );
nand NAND2_2292 ( P1_U4988 , P1_ADDR_REG_13_ , P1_U4922 );
nand NAND2_2293 ( P1_U4989 , P1_R1105_U79 , P1_U3041 );
nand NAND2_2294 ( P1_U4990 , P1_U3039 , P1_U3488 );
nand NAND2_2295 ( P1_U4991 , P1_R1162_U79 , P1_U3037 );
nand NAND3_2296 ( P1_U4992 , P1_U4990 , P1_U4989 , P1_U4991 );
nand NAND2_2297 ( P1_U4993 , P1_U3043 , P1_U4992 );
nand NAND2_2298 ( P1_U4994 , P1_R1105_U79 , P1_U3042 );
nand NAND2_2299 ( P1_U4995 , P1_REG3_REG_12_ , P1_U3084 );
nand NAND2_2300 ( P1_U4996 , P1_U3040 , P1_U3488 );
nand NAND2_2301 ( P1_U4997 , P1_R1162_U79 , P1_U3038 );
nand NAND2_2302 ( P1_U4998 , P1_ADDR_REG_12_ , P1_U4922 );
nand NAND2_2303 ( P1_U4999 , P1_R1105_U80 , P1_U3041 );
nand NAND2_2304 ( P1_U5000 , P1_U3039 , P1_U3485 );
nand NAND2_2305 ( P1_U5001 , P1_R1162_U80 , P1_U3037 );
nand NAND3_2306 ( P1_U5002 , P1_U5000 , P1_U4999 , P1_U5001 );
nand NAND2_2307 ( P1_U5003 , P1_U3043 , P1_U5002 );
nand NAND2_2308 ( P1_U5004 , P1_R1105_U80 , P1_U3042 );
nand NAND2_2309 ( P1_U5005 , P1_REG3_REG_11_ , P1_U3084 );
nand NAND2_2310 ( P1_U5006 , P1_U3040 , P1_U3485 );
nand NAND2_2311 ( P1_U5007 , P1_R1162_U80 , P1_U3038 );
nand NAND2_2312 ( P1_U5008 , P1_ADDR_REG_11_ , P1_U4922 );
nand NAND2_2313 ( P1_U5009 , P1_R1105_U10 , P1_U3041 );
nand NAND2_2314 ( P1_U5010 , P1_U3039 , P1_U3482 );
nand NAND2_2315 ( P1_U5011 , P1_R1162_U10 , P1_U3037 );
nand NAND3_2316 ( P1_U5012 , P1_U5010 , P1_U5009 , P1_U5011 );
nand NAND2_2317 ( P1_U5013 , P1_U3043 , P1_U5012 );
nand NAND2_2318 ( P1_U5014 , P1_R1105_U10 , P1_U3042 );
nand NAND2_2319 ( P1_U5015 , P1_REG3_REG_10_ , P1_U3084 );
nand NAND2_2320 ( P1_U5016 , P1_U3040 , P1_U3482 );
nand NAND2_2321 ( P1_U5017 , P1_R1162_U10 , P1_U3038 );
nand NAND2_2322 ( P1_U5018 , P1_ADDR_REG_10_ , P1_U4922 );
nand NAND2_2323 ( P1_U5019 , P1_R1105_U70 , P1_U3041 );
nand NAND2_2324 ( P1_U5020 , P1_U3039 , P1_U3479 );
nand NAND2_2325 ( P1_U5021 , P1_R1162_U70 , P1_U3037 );
nand NAND3_2326 ( P1_U5022 , P1_U5020 , P1_U5019 , P1_U5021 );
nand NAND2_2327 ( P1_U5023 , P1_U3043 , P1_U5022 );
nand NAND2_2328 ( P1_U5024 , P1_R1105_U70 , P1_U3042 );
nand NAND2_2329 ( P1_U5025 , P1_REG3_REG_9_ , P1_U3084 );
nand NAND2_2330 ( P1_U5026 , P1_U3040 , P1_U3479 );
nand NAND2_2331 ( P1_U5027 , P1_R1162_U70 , P1_U3038 );
nand NAND2_2332 ( P1_U5028 , P1_ADDR_REG_9_ , P1_U4922 );
nand NAND2_2333 ( P1_U5029 , P1_R1105_U71 , P1_U3041 );
nand NAND2_2334 ( P1_U5030 , P1_U3039 , P1_U3476 );
nand NAND2_2335 ( P1_U5031 , P1_R1162_U71 , P1_U3037 );
nand NAND3_2336 ( P1_U5032 , P1_U5030 , P1_U5029 , P1_U5031 );
nand NAND2_2337 ( P1_U5033 , P1_U3043 , P1_U5032 );
nand NAND2_2338 ( P1_U5034 , P1_R1105_U71 , P1_U3042 );
nand NAND2_2339 ( P1_U5035 , P1_REG3_REG_8_ , P1_U3084 );
nand NAND2_2340 ( P1_U5036 , P1_U3040 , P1_U3476 );
nand NAND2_2341 ( P1_U5037 , P1_R1162_U71 , P1_U3038 );
nand NAND2_2342 ( P1_U5038 , P1_ADDR_REG_8_ , P1_U4922 );
nand NAND2_2343 ( P1_U5039 , P1_R1105_U16 , P1_U3041 );
nand NAND2_2344 ( P1_U5040 , P1_U3039 , P1_U3473 );
nand NAND2_2345 ( P1_U5041 , P1_R1162_U16 , P1_U3037 );
nand NAND3_2346 ( P1_U5042 , P1_U5040 , P1_U5039 , P1_U5041 );
nand NAND2_2347 ( P1_U5043 , P1_U3043 , P1_U5042 );
nand NAND2_2348 ( P1_U5044 , P1_R1105_U16 , P1_U3042 );
nand NAND2_2349 ( P1_U5045 , P1_REG3_REG_7_ , P1_U3084 );
nand NAND2_2350 ( P1_U5046 , P1_U3040 , P1_U3473 );
nand NAND2_2351 ( P1_U5047 , P1_R1162_U16 , P1_U3038 );
nand NAND2_2352 ( P1_U5048 , P1_ADDR_REG_7_ , P1_U4922 );
nand NAND2_2353 ( P1_U5049 , P1_R1105_U72 , P1_U3041 );
nand NAND2_2354 ( P1_U5050 , P1_U3039 , P1_U3470 );
nand NAND2_2355 ( P1_U5051 , P1_R1162_U72 , P1_U3037 );
nand NAND3_2356 ( P1_U5052 , P1_U5050 , P1_U5049 , P1_U5051 );
nand NAND2_2357 ( P1_U5053 , P1_U3043 , P1_U5052 );
nand NAND2_2358 ( P1_U5054 , P1_R1105_U72 , P1_U3042 );
nand NAND2_2359 ( P1_U5055 , P1_REG3_REG_6_ , P1_U3084 );
nand NAND2_2360 ( P1_U5056 , P1_U3040 , P1_U3470 );
nand NAND2_2361 ( P1_U5057 , P1_R1162_U72 , P1_U3038 );
nand NAND2_2362 ( P1_U5058 , P1_ADDR_REG_6_ , P1_U4922 );
nand NAND2_2363 ( P1_U5059 , P1_R1105_U15 , P1_U3041 );
nand NAND2_2364 ( P1_U5060 , P1_U3039 , P1_U3467 );
nand NAND2_2365 ( P1_U5061 , P1_R1162_U15 , P1_U3037 );
nand NAND3_2366 ( P1_U5062 , P1_U5060 , P1_U5059 , P1_U5061 );
nand NAND2_2367 ( P1_U5063 , P1_U3043 , P1_U5062 );
nand NAND2_2368 ( P1_U5064 , P1_R1105_U15 , P1_U3042 );
nand NAND2_2369 ( P1_U5065 , P1_REG3_REG_5_ , P1_U3084 );
nand NAND2_2370 ( P1_U5066 , P1_U3040 , P1_U3467 );
nand NAND2_2371 ( P1_U5067 , P1_R1162_U15 , P1_U3038 );
nand NAND2_2372 ( P1_U5068 , P1_ADDR_REG_5_ , P1_U4922 );
nand NAND2_2373 ( P1_U5069 , P1_R1105_U73 , P1_U3041 );
nand NAND2_2374 ( P1_U5070 , P1_U3039 , P1_U3464 );
nand NAND2_2375 ( P1_U5071 , P1_R1162_U73 , P1_U3037 );
nand NAND3_2376 ( P1_U5072 , P1_U5070 , P1_U5069 , P1_U5071 );
nand NAND2_2377 ( P1_U5073 , P1_U3043 , P1_U5072 );
nand NAND2_2378 ( P1_U5074 , P1_R1105_U73 , P1_U3042 );
nand NAND2_2379 ( P1_U5075 , P1_REG3_REG_4_ , P1_U3084 );
nand NAND2_2380 ( P1_U5076 , P1_U3040 , P1_U3464 );
nand NAND2_2381 ( P1_U5077 , P1_R1162_U73 , P1_U3038 );
nand NAND2_2382 ( P1_U5078 , P1_ADDR_REG_4_ , P1_U4922 );
nand NAND2_2383 ( P1_U5079 , P1_R1105_U74 , P1_U3041 );
nand NAND2_2384 ( P1_U5080 , P1_U3039 , P1_U3461 );
nand NAND2_2385 ( P1_U5081 , P1_R1162_U74 , P1_U3037 );
nand NAND3_2386 ( P1_U5082 , P1_U5080 , P1_U5079 , P1_U5081 );
nand NAND2_2387 ( P1_U5083 , P1_U3043 , P1_U5082 );
nand NAND2_2388 ( P1_U5084 , P1_R1105_U74 , P1_U3042 );
nand NAND2_2389 ( P1_U5085 , P1_REG3_REG_3_ , P1_U3084 );
nand NAND2_2390 ( P1_U5086 , P1_U3040 , P1_U3461 );
nand NAND2_2391 ( P1_U5087 , P1_R1162_U74 , P1_U3038 );
nand NAND2_2392 ( P1_U5088 , P1_ADDR_REG_3_ , P1_U4922 );
nand NAND2_2393 ( P1_U5089 , P1_R1105_U14 , P1_U3041 );
nand NAND2_2394 ( P1_U5090 , P1_U3039 , P1_U3458 );
nand NAND2_2395 ( P1_U5091 , P1_R1162_U14 , P1_U3037 );
nand NAND3_2396 ( P1_U5092 , P1_U5090 , P1_U5089 , P1_U5091 );
nand NAND2_2397 ( P1_U5093 , P1_U3043 , P1_U5092 );
nand NAND2_2398 ( P1_U5094 , P1_R1105_U14 , P1_U3042 );
nand NAND2_2399 ( P1_U5095 , P1_REG3_REG_2_ , P1_U3084 );
nand NAND2_2400 ( P1_U5096 , P1_U3040 , P1_U3458 );
nand NAND2_2401 ( P1_U5097 , P1_R1162_U14 , P1_U3038 );
nand NAND2_2402 ( P1_U5098 , P1_ADDR_REG_2_ , P1_U4922 );
nand NAND2_2403 ( P1_U5099 , P1_R1105_U68 , P1_U3041 );
nand NAND2_2404 ( P1_U5100 , P1_U3039 , P1_U3455 );
nand NAND2_2405 ( P1_U5101 , P1_R1162_U68 , P1_U3037 );
nand NAND3_2406 ( P1_U5102 , P1_U5100 , P1_U5099 , P1_U5101 );
nand NAND2_2407 ( P1_U5103 , P1_U3043 , P1_U5102 );
nand NAND2_2408 ( P1_U5104 , P1_R1105_U68 , P1_U3042 );
nand NAND2_2409 ( P1_U5105 , P1_REG3_REG_1_ , P1_U3084 );
nand NAND2_2410 ( P1_U5106 , P1_U3040 , P1_U3455 );
nand NAND2_2411 ( P1_U5107 , P1_R1162_U68 , P1_U3038 );
nand NAND2_2412 ( P1_U5108 , P1_ADDR_REG_1_ , P1_U4922 );
nand NAND2_2413 ( P1_U5109 , P1_R1105_U69 , P1_U3041 );
nand NAND2_2414 ( P1_U5110 , P1_U3039 , P1_U3449 );
nand NAND2_2415 ( P1_U5111 , P1_R1162_U69 , P1_U3037 );
nand NAND3_2416 ( P1_U5112 , P1_U5110 , P1_U5109 , P1_U5111 );
nand NAND2_2417 ( P1_U5113 , P1_U3043 , P1_U5112 );
nand NAND2_2418 ( P1_U5114 , P1_R1105_U69 , P1_U3042 );
nand NAND2_2419 ( P1_U5115 , P1_REG3_REG_0_ , P1_U3084 );
nand NAND2_2420 ( P1_U5116 , P1_U3040 , P1_U3449 );
nand NAND2_2421 ( P1_U5117 , P1_R1162_U69 , P1_U3038 );
nand NAND2_2422 ( P1_U5118 , P1_ADDR_REG_0_ , P1_U4922 );
not NOT1_2423 ( P1_U5119 , P1_U3982 );
nand NAND3_2424 ( P1_U5120 , P1_U6198 , P1_U6197 , P1_U3875 );
nand NAND2_2425 ( P1_U5121 , P1_U5703 , P1_U3427 );
nand NAND2_2426 ( P1_U5122 , P1_U3861 , P1_U5121 );
nand NAND2_2427 ( P1_U5123 , P1_B_REG , P1_U5122 );
nand NAND2_2428 ( P1_U5124 , P1_U3036 , P1_U3077 );
nand NAND2_2429 ( P1_U5125 , P1_U3034 , P1_U3071 );
nand NAND2_2430 ( P1_U5126 , P1_ADD_99_U73 , P1_U3431 );
nand NAND3_2431 ( P1_U5127 , P1_U5126 , P1_U5124 , P1_U5125 );
nand NAND3_2432 ( P1_U5128 , P1_U3363 , P1_U3360 , P1_U3361 );
nand NAND3_2433 ( P1_U5129 , P1_U3365 , P1_U3419 , P1_U3364 );
nand NAND2_2434 ( P1_U5130 , P1_U5710 , P1_U5129 );
nand NAND2_2435 ( P1_U5131 , P1_U5719 , P1_U5128 );
nand NAND3_2436 ( P1_U5132 , P1_U5131 , P1_U5130 , P1_U3877 );
nand NAND2_2437 ( P1_U5133 , P1_U5132 , P1_U3431 );
not NOT1_2438 ( P1_U5134 , P1_U3433 );
nand NAND2_2439 ( P1_U5135 , P1_U3498 , P1_U5686 );
nand NAND2_2440 ( P1_U5136 , P1_ADD_99_U73 , P1_U5685 );
nand NAND2_2441 ( P1_U5137 , P1_U4027 , P1_U5127 );
nand NAND2_2442 ( P1_U5138 , P1_R1165_U104 , P1_U3027 );
nand NAND2_2443 ( P1_U5139 , P1_REG3_REG_15_ , P1_U3084 );
nand NAND2_2444 ( P1_U5140 , P1_U3036 , P1_U3056 );
nand NAND2_2445 ( P1_U5141 , P1_U3034 , P1_U3051 );
nand NAND2_2446 ( P1_U5142 , P1_ADD_99_U62 , P1_U3431 );
nand NAND3_2447 ( P1_U5143 , P1_U5142 , P1_U5140 , P1_U5141 );
nand NAND2_2448 ( P1_U5144 , P1_U3422 , P1_U3431 );
nand NAND2_2449 ( P1_U5145 , P1_U5134 , P1_U5144 );
nand NAND2_2450 ( P1_U5146 , P1_U4005 , P1_U3422 );
nand NAND2_2451 ( P1_U5147 , P1_U3418 , P1_U5146 );
nand NAND2_2452 ( P1_U5148 , P1_U3045 , P1_U4009 );
nand NAND2_2453 ( P1_U5149 , P1_U3044 , P1_ADD_99_U62 );
nand NAND2_2454 ( P1_U5150 , P1_U4027 , P1_U5143 );
nand NAND2_2455 ( P1_U5151 , P1_R1165_U13 , P1_U3027 );
nand NAND2_2456 ( P1_U5152 , P1_REG3_REG_26_ , P1_U3084 );
nand NAND2_2457 ( P1_U5153 , P1_U3036 , P1_U3065 );
nand NAND2_2458 ( P1_U5154 , P1_U3034 , P1_U3068 );
nand NAND2_2459 ( P1_U5155 , P1_ADD_99_U57 , P1_U3431 );
nand NAND3_2460 ( P1_U5156 , P1_U5154 , P1_U5153 , P1_U5155 );
nand NAND2_2461 ( P1_U5157 , P1_U3471 , P1_U5686 );
nand NAND2_2462 ( P1_U5158 , P1_ADD_99_U57 , P1_U5685 );
nand NAND2_2463 ( P1_U5159 , P1_U4027 , P1_U5156 );
nand NAND2_2464 ( P1_U5160 , P1_R1165_U89 , P1_U3027 );
nand NAND2_2465 ( P1_U5161 , P1_REG3_REG_6_ , P1_U3084 );
nand NAND2_2466 ( P1_U5162 , P1_U3036 , P1_U3067 );
nand NAND2_2467 ( P1_U5163 , P1_U3034 , P1_U3079 );
nand NAND2_2468 ( P1_U5164 , P1_ADD_99_U70 , P1_U3431 );
nand NAND3_2469 ( P1_U5165 , P1_U5164 , P1_U5162 , P1_U5163 );
nand NAND2_2470 ( P1_U5166 , P1_U3507 , P1_U5686 );
nand NAND2_2471 ( P1_U5167 , P1_ADD_99_U70 , P1_U5685 );
nand NAND2_2472 ( P1_U5168 , P1_U4027 , P1_U5165 );
nand NAND2_2473 ( P1_U5169 , P1_R1165_U102 , P1_U3027 );
nand NAND2_2474 ( P1_U5170 , P1_REG3_REG_18_ , P1_U3084 );
nand NAND2_2475 ( P1_U5171 , P1_U3036 , P1_U3076 );
nand NAND2_2476 ( P1_U5172 , P1_U3034 , P1_U3062 );
nand NAND2_2477 ( P1_U5173 , P1_REG3_REG_2_ , P1_U3431 );
nand NAND3_2478 ( P1_U5174 , P1_U5172 , P1_U5171 , P1_U5173 );
nand NAND2_2479 ( P1_U5175 , P1_U3459 , P1_U5686 );
nand NAND2_2480 ( P1_U5176 , P1_REG3_REG_2_ , P1_U5685 );
nand NAND2_2481 ( P1_U5177 , P1_U4027 , P1_U5174 );
nand NAND2_2482 ( P1_U5178 , P1_R1165_U92 , P1_U3027 );
nand NAND2_2483 ( P1_U5179 , P1_REG3_REG_2_ , P1_U3084 );
nand NAND2_2484 ( P1_U5180 , P1_U3036 , P1_U3060 );
nand NAND2_2485 ( P1_U5181 , P1_U3034 , P1_U3070 );
nand NAND2_2486 ( P1_U5182 , P1_ADD_99_U77 , P1_U3431 );
nand NAND3_2487 ( P1_U5183 , P1_U5181 , P1_U5180 , P1_U5182 );
nand NAND2_2488 ( P1_U5184 , P1_U3486 , P1_U5686 );
nand NAND2_2489 ( P1_U5185 , P1_ADD_99_U77 , P1_U5685 );
nand NAND2_2490 ( P1_U5186 , P1_U4027 , P1_U5183 );
nand NAND2_2491 ( P1_U5187 , P1_R1165_U107 , P1_U3027 );
nand NAND2_2492 ( P1_U5188 , P1_REG3_REG_11_ , P1_U3084 );
nand NAND2_2493 ( P1_U5189 , P1_U3036 , P1_U3073 );
nand NAND2_2494 ( P1_U5190 , P1_U3034 , P1_U3064 );
nand NAND2_2495 ( P1_U5191 , P1_ADD_99_U66 , P1_U3431 );
nand NAND3_2496 ( P1_U5192 , P1_U5191 , P1_U5189 , P1_U5190 );
nand NAND2_2497 ( P1_U5193 , P1_U3045 , P1_U4013 );
nand NAND2_2498 ( P1_U5194 , P1_U3044 , P1_ADD_99_U66 );
nand NAND2_2499 ( P1_U5195 , P1_U4027 , P1_U5192 );
nand NAND2_2500 ( P1_U5196 , P1_R1165_U98 , P1_U3027 );
nand NAND2_2501 ( P1_U5197 , P1_REG3_REG_22_ , P1_U3084 );
nand NAND2_2502 ( P1_U5198 , P1_U3036 , P1_U3070 );
nand NAND2_2503 ( P1_U5199 , P1_U3034 , P1_U3077 );
nand NAND2_2504 ( P1_U5200 , P1_ADD_99_U75 , P1_U3431 );
nand NAND3_2505 ( P1_U5201 , P1_U5200 , P1_U5198 , P1_U5199 );
nand NAND2_2506 ( P1_U5202 , P1_U3492 , P1_U5686 );
nand NAND2_2507 ( P1_U5203 , P1_ADD_99_U75 , P1_U5685 );
nand NAND2_2508 ( P1_U5204 , P1_U4027 , P1_U5201 );
nand NAND2_2509 ( P1_U5205 , P1_R1165_U10 , P1_U3027 );
nand NAND2_2510 ( P1_U5206 , P1_REG3_REG_13_ , P1_U3084 );
nand NAND2_2511 ( P1_U5207 , P1_U3036 , P1_U3079 );
nand NAND2_2512 ( P1_U5208 , P1_U3034 , P1_U3073 );
nand NAND2_2513 ( P1_U5209 , P1_ADD_99_U68 , P1_U3431 );
nand NAND3_2514 ( P1_U5210 , P1_U5209 , P1_U5207 , P1_U5208 );
nand NAND2_2515 ( P1_U5211 , P1_U3045 , P1_U4015 );
nand NAND2_2516 ( P1_U5212 , P1_U3044 , P1_ADD_99_U68 );
nand NAND2_2517 ( P1_U5213 , P1_U4027 , P1_U5210 );
nand NAND2_2518 ( P1_U5214 , P1_R1165_U99 , P1_U3027 );
nand NAND2_2519 ( P1_U5215 , P1_REG3_REG_20_ , P1_U3084 );
nand NAND2_2520 ( P1_U5216 , P1_U3432 , P1_U3430 );
nand NAND2_2521 ( P1_U5217 , P1_U5216 , P1_U3431 );
nand NAND2_2522 ( P1_U5218 , P1_U4028 , P1_U5217 );
nand NAND2_2523 ( P1_U5219 , P1_U3883 , P1_U3034 );
nand NAND2_2524 ( P1_U5220 , P1_U3451 , P1_U5686 );
nand NAND2_2525 ( P1_U5221 , P1_REG3_REG_0_ , P1_U5218 );
nand NAND2_2526 ( P1_U5222 , P1_R1165_U86 , P1_U3027 );
nand NAND2_2527 ( P1_U5223 , P1_REG3_REG_0_ , P1_U3084 );
nand NAND2_2528 ( P1_U5224 , P1_U3036 , P1_U3082 );
nand NAND2_2529 ( P1_U5225 , P1_U3034 , P1_U3060 );
nand NAND2_2530 ( P1_U5226 , P1_ADD_99_U54 , P1_U3431 );
nand NAND3_2531 ( P1_U5227 , P1_U5225 , P1_U5224 , P1_U5226 );
nand NAND2_2532 ( P1_U5228 , P1_U3480 , P1_U5686 );
nand NAND2_2533 ( P1_U5229 , P1_ADD_99_U54 , P1_U5685 );
nand NAND2_2534 ( P1_U5230 , P1_U4027 , P1_U5227 );
nand NAND2_2535 ( P1_U5231 , P1_R1165_U87 , P1_U3027 );
nand NAND2_2536 ( P1_U5232 , P1_REG3_REG_9_ , P1_U3084 );
nand NAND2_2537 ( P1_U5233 , P1_U3036 , P1_U3062 );
nand NAND2_2538 ( P1_U5234 , P1_U3034 , P1_U3065 );
nand NAND2_2539 ( P1_U5235 , P1_ADD_99_U59 , P1_U3431 );
nand NAND3_2540 ( P1_U5236 , P1_U5234 , P1_U5233 , P1_U5235 );
nand NAND2_2541 ( P1_U5237 , P1_U3465 , P1_U5686 );
nand NAND2_2542 ( P1_U5238 , P1_ADD_99_U59 , P1_U5685 );
nand NAND2_2543 ( P1_U5239 , P1_U4027 , P1_U5236 );
nand NAND2_2544 ( P1_U5240 , P1_R1165_U91 , P1_U3027 );
nand NAND2_2545 ( P1_U5241 , P1_REG3_REG_4_ , P1_U3084 );
nand NAND2_2546 ( P1_U5242 , P1_U3036 , P1_U3064 );
nand NAND2_2547 ( P1_U5243 , P1_U3034 , P1_U3056 );
nand NAND2_2548 ( P1_U5244 , P1_ADD_99_U64 , P1_U3431 );
nand NAND3_2549 ( P1_U5245 , P1_U5244 , P1_U5242 , P1_U5243 );
nand NAND2_2550 ( P1_U5246 , P1_U3045 , P1_U4011 );
nand NAND2_2551 ( P1_U5247 , P1_U3044 , P1_ADD_99_U64 );
nand NAND2_2552 ( P1_U5248 , P1_U4027 , P1_U5245 );
nand NAND2_2553 ( P1_U5249 , P1_R1165_U96 , P1_U3027 );
nand NAND2_2554 ( P1_U5250 , P1_REG3_REG_24_ , P1_U3084 );
nand NAND2_2555 ( P1_U5251 , P1_U3036 , P1_U3071 );
nand NAND2_2556 ( P1_U5252 , P1_U3034 , P1_U3080 );
nand NAND2_2557 ( P1_U5253 , P1_ADD_99_U71 , P1_U3431 );
nand NAND3_2558 ( P1_U5254 , P1_U5253 , P1_U5251 , P1_U5252 );
nand NAND2_2559 ( P1_U5255 , P1_U3504 , P1_U5686 );
nand NAND2_2560 ( P1_U5256 , P1_ADD_99_U71 , P1_U5685 );
nand NAND2_2561 ( P1_U5257 , P1_U4027 , P1_U5254 );
nand NAND2_2562 ( P1_U5258 , P1_R1165_U11 , P1_U3027 );
nand NAND2_2563 ( P1_U5259 , P1_REG3_REG_17_ , P1_U3084 );
nand NAND2_2564 ( P1_U5260 , P1_U3036 , P1_U3058 );
nand NAND2_2565 ( P1_U5261 , P1_U3034 , P1_U3069 );
nand NAND2_2566 ( P1_U5262 , P1_ADD_99_U58 , P1_U3431 );
nand NAND3_2567 ( P1_U5263 , P1_U5261 , P1_U5260 , P1_U5262 );
nand NAND2_2568 ( P1_U5264 , P1_U3468 , P1_U5686 );
nand NAND2_2569 ( P1_U5265 , P1_ADD_99_U58 , P1_U5685 );
nand NAND2_2570 ( P1_U5266 , P1_U4027 , P1_U5263 );
nand NAND2_2571 ( P1_U5267 , P1_R1165_U90 , P1_U3027 );
nand NAND2_2572 ( P1_U5268 , P1_REG3_REG_5_ , P1_U3084 );
nand NAND2_2573 ( P1_U5269 , P1_U3036 , P1_U3072 );
nand NAND2_2574 ( P1_U5270 , P1_U3034 , P1_U3067 );
nand NAND2_2575 ( P1_U5271 , P1_ADD_99_U72 , P1_U3431 );
nand NAND3_2576 ( P1_U5272 , P1_U5271 , P1_U5269 , P1_U5270 );
nand NAND2_2577 ( P1_U5273 , P1_U3501 , P1_U5686 );
nand NAND2_2578 ( P1_U5274 , P1_ADD_99_U72 , P1_U5685 );
nand NAND2_2579 ( P1_U5275 , P1_U4027 , P1_U5272 );
nand NAND2_2580 ( P1_U5276 , P1_R1165_U103 , P1_U3027 );
nand NAND2_2581 ( P1_U5277 , P1_REG3_REG_16_ , P1_U3084 );
nand NAND2_2582 ( P1_U5278 , P1_U3036 , P1_U3063 );
nand NAND2_2583 ( P1_U5279 , P1_U3034 , P1_U3055 );
nand NAND2_2584 ( P1_U5280 , P1_ADD_99_U63 , P1_U3431 );
nand NAND3_2585 ( P1_U5281 , P1_U5280 , P1_U5278 , P1_U5279 );
nand NAND2_2586 ( P1_U5282 , P1_U3045 , P1_U4010 );
nand NAND2_2587 ( P1_U5283 , P1_U3044 , P1_ADD_99_U63 );
nand NAND2_2588 ( P1_U5284 , P1_U4027 , P1_U5281 );
nand NAND2_2589 ( P1_U5285 , P1_R1165_U95 , P1_U3027 );
nand NAND2_2590 ( P1_U5286 , P1_REG3_REG_25_ , P1_U3084 );
nand NAND2_2591 ( P1_U5287 , P1_U3036 , P1_U3061 );
nand NAND2_2592 ( P1_U5288 , P1_U3034 , P1_U3078 );
nand NAND2_2593 ( P1_U5289 , P1_ADD_99_U76 , P1_U3431 );
nand NAND3_2594 ( P1_U5290 , P1_U5289 , P1_U5287 , P1_U5288 );
nand NAND2_2595 ( P1_U5291 , P1_U3489 , P1_U5686 );
nand NAND2_2596 ( P1_U5292 , P1_ADD_99_U76 , P1_U5685 );
nand NAND2_2597 ( P1_U5293 , P1_U4027 , P1_U5290 );
nand NAND2_2598 ( P1_U5294 , P1_R1165_U106 , P1_U3027 );
nand NAND2_2599 ( P1_U5295 , P1_REG3_REG_12_ , P1_U3084 );
nand NAND2_2600 ( P1_U5296 , P1_U3036 , P1_U3074 );
nand NAND2_2601 ( P1_U5297 , P1_U3034 , P1_U3059 );
nand NAND2_2602 ( P1_U5298 , P1_ADD_99_U67 , P1_U3431 );
nand NAND3_2603 ( P1_U5299 , P1_U5298 , P1_U5296 , P1_U5297 );
nand NAND2_2604 ( P1_U5300 , P1_U3045 , P1_U4014 );
nand NAND2_2605 ( P1_U5301 , P1_U3044 , P1_ADD_99_U67 );
nand NAND2_2606 ( P1_U5302 , P1_U4027 , P1_U5299 );
nand NAND2_2607 ( P1_U5303 , P1_R1165_U12 , P1_U3027 );
nand NAND2_2608 ( P1_U5304 , P1_REG3_REG_21_ , P1_U3084 );
nand NAND2_2609 ( P1_U5305 , P1_U3036 , P1_U3075 );
nand NAND2_2610 ( P1_U5306 , P1_U3034 , P1_U3066 );
nand NAND2_2611 ( P1_U5307 , P1_REG3_REG_1_ , P1_U3431 );
nand NAND3_2612 ( P1_U5308 , P1_U5306 , P1_U5305 , P1_U5307 );
nand NAND2_2613 ( P1_U5309 , P1_U3456 , P1_U5686 );
nand NAND2_2614 ( P1_U5310 , P1_REG3_REG_1_ , P1_U5685 );
nand NAND2_2615 ( P1_U5311 , P1_U4027 , P1_U5308 );
nand NAND2_2616 ( P1_U5312 , P1_R1165_U100 , P1_U3027 );
nand NAND2_2617 ( P1_U5313 , P1_REG3_REG_1_ , P1_U3084 );
nand NAND2_2618 ( P1_U5314 , P1_U3036 , P1_U3068 );
nand NAND2_2619 ( P1_U5315 , P1_U3034 , P1_U3081 );
nand NAND2_2620 ( P1_U5316 , P1_ADD_99_U55 , P1_U3431 );
nand NAND3_2621 ( P1_U5317 , P1_U5315 , P1_U5314 , P1_U5316 );
nand NAND2_2622 ( P1_U5318 , P1_U3477 , P1_U5686 );
nand NAND2_2623 ( P1_U5319 , P1_ADD_99_U55 , P1_U5685 );
nand NAND2_2624 ( P1_U5320 , P1_U4027 , P1_U5317 );
nand NAND2_2625 ( P1_U5321 , P1_R1165_U88 , P1_U3027 );
nand NAND2_2626 ( P1_U5322 , P1_REG3_REG_8_ , P1_U3084 );
nand NAND2_2627 ( P1_U5323 , P1_U3036 , P1_U3051 );
nand NAND2_2628 ( P1_U5324 , P1_U3034 , P1_U3053 );
nand NAND2_2629 ( P1_U5325 , P1_ADD_99_U60 , P1_U3431 );
nand NAND3_2630 ( P1_U5326 , P1_U5324 , P1_U5323 , P1_U5325 );
nand NAND2_2631 ( P1_U5327 , P1_U3045 , P1_U4007 );
nand NAND2_2632 ( P1_U5328 , P1_U3044 , P1_ADD_99_U60 );
nand NAND2_2633 ( P1_U5329 , P1_U4027 , P1_U5326 );
nand NAND2_2634 ( P1_U5330 , P1_R1165_U93 , P1_U3027 );
nand NAND2_2635 ( P1_U5331 , P1_REG3_REG_28_ , P1_U3084 );
nand NAND2_2636 ( P1_U5332 , P1_U3036 , P1_U3080 );
nand NAND2_2637 ( P1_U5333 , P1_U3034 , P1_U3074 );
nand NAND2_2638 ( P1_U5334 , P1_ADD_99_U69 , P1_U3431 );
nand NAND3_2639 ( P1_U5335 , P1_U5334 , P1_U5332 , P1_U5333 );
nand NAND2_2640 ( P1_U5336 , P1_U3509 , P1_U5686 );
nand NAND2_2641 ( P1_U5337 , P1_ADD_99_U69 , P1_U5685 );
nand NAND2_2642 ( P1_U5338 , P1_U4027 , P1_U5335 );
nand NAND2_2643 ( P1_U5339 , P1_R1165_U101 , P1_U3027 );
nand NAND2_2644 ( P1_U5340 , P1_REG3_REG_19_ , P1_U3084 );
nand NAND2_2645 ( P1_U5341 , P1_U3036 , P1_U3066 );
nand NAND2_2646 ( P1_U5342 , P1_U3034 , P1_U3058 );
nand NAND2_2647 ( P1_U5343 , P1_ADD_99_U4 , P1_U3431 );
nand NAND3_2648 ( P1_U5344 , P1_U5342 , P1_U5341 , P1_U5343 );
nand NAND2_2649 ( P1_U5345 , P1_U3462 , P1_U5686 );
nand NAND2_2650 ( P1_U5346 , P1_ADD_99_U4 , P1_U5685 );
nand NAND2_2651 ( P1_U5347 , P1_U4027 , P1_U5344 );
nand NAND2_2652 ( P1_U5348 , P1_R1165_U14 , P1_U3027 );
nand NAND2_2653 ( P1_U5349 , P1_REG3_REG_3_ , P1_U3084 );
nand NAND2_2654 ( P1_U5350 , P1_U3036 , P1_U3081 );
nand NAND2_2655 ( P1_U5351 , P1_U3034 , P1_U3061 );
nand NAND2_2656 ( P1_U5352 , P1_ADD_99_U78 , P1_U3431 );
nand NAND3_2657 ( P1_U5353 , P1_U5351 , P1_U5350 , P1_U5352 );
nand NAND2_2658 ( P1_U5354 , P1_U3483 , P1_U5686 );
nand NAND2_2659 ( P1_U5355 , P1_ADD_99_U78 , P1_U5685 );
nand NAND2_2660 ( P1_U5356 , P1_U4027 , P1_U5353 );
nand NAND2_2661 ( P1_U5357 , P1_R1165_U108 , P1_U3027 );
nand NAND2_2662 ( P1_U5358 , P1_REG3_REG_10_ , P1_U3084 );
nand NAND2_2663 ( P1_U5359 , P1_U3036 , P1_U3059 );
nand NAND2_2664 ( P1_U5360 , P1_U3034 , P1_U3063 );
nand NAND2_2665 ( P1_U5361 , P1_ADD_99_U65 , P1_U3431 );
nand NAND3_2666 ( P1_U5362 , P1_U5361 , P1_U5359 , P1_U5360 );
nand NAND2_2667 ( P1_U5363 , P1_U3045 , P1_U4012 );
nand NAND2_2668 ( P1_U5364 , P1_U3044 , P1_ADD_99_U65 );
nand NAND2_2669 ( P1_U5365 , P1_U4027 , P1_U5362 );
nand NAND2_2670 ( P1_U5366 , P1_R1165_U97 , P1_U3027 );
nand NAND2_2671 ( P1_U5367 , P1_REG3_REG_23_ , P1_U3084 );
nand NAND2_2672 ( P1_U5368 , P1_U3036 , P1_U3078 );
nand NAND2_2673 ( P1_U5369 , P1_U3034 , P1_U3072 );
nand NAND2_2674 ( P1_U5370 , P1_ADD_99_U74 , P1_U3431 );
nand NAND3_2675 ( P1_U5371 , P1_U5370 , P1_U5368 , P1_U5369 );
nand NAND2_2676 ( P1_U5372 , P1_U3495 , P1_U5686 );
nand NAND2_2677 ( P1_U5373 , P1_ADD_99_U74 , P1_U5685 );
nand NAND2_2678 ( P1_U5374 , P1_U4027 , P1_U5371 );
nand NAND2_2679 ( P1_U5375 , P1_R1165_U105 , P1_U3027 );
nand NAND2_2680 ( P1_U5376 , P1_REG3_REG_14_ , P1_U3084 );
nand NAND2_2681 ( P1_U5377 , P1_U3036 , P1_U3055 );
nand NAND2_2682 ( P1_U5378 , P1_U3034 , P1_U3052 );
nand NAND2_2683 ( P1_U5379 , P1_ADD_99_U61 , P1_U3431 );
nand NAND3_2684 ( P1_U5380 , P1_U5379 , P1_U5377 , P1_U5378 );
nand NAND2_2685 ( P1_U5381 , P1_U3045 , P1_U4008 );
nand NAND2_2686 ( P1_U5382 , P1_U3044 , P1_ADD_99_U61 );
nand NAND2_2687 ( P1_U5383 , P1_U4027 , P1_U5380 );
nand NAND2_2688 ( P1_U5384 , P1_R1165_U94 , P1_U3027 );
nand NAND2_2689 ( P1_U5385 , P1_REG3_REG_27_ , P1_U3084 );
nand NAND2_2690 ( P1_U5386 , P1_U3036 , P1_U3069 );
nand NAND2_2691 ( P1_U5387 , P1_U3034 , P1_U3082 );
nand NAND2_2692 ( P1_U5388 , P1_ADD_99_U56 , P1_U3431 );
nand NAND3_2693 ( P1_U5389 , P1_U5387 , P1_U5386 , P1_U5388 );
nand NAND2_2694 ( P1_U5390 , P1_U3474 , P1_U5686 );
nand NAND2_2695 ( P1_U5391 , P1_ADD_99_U56 , P1_U5685 );
nand NAND2_2696 ( P1_U5392 , P1_U4027 , P1_U5389 );
nand NAND2_2697 ( P1_U5393 , P1_R1165_U15 , P1_U3027 );
nand NAND2_2698 ( P1_U5394 , P1_REG3_REG_7_ , P1_U3084 );
nand NAND2_2699 ( P1_U5395 , P1_U3450 , P1_U3374 );
nand NAND2_2700 ( P1_U5396 , P1_U3447 , P1_U5395 );
nand NAND3_2701 ( P1_U5397 , P1_U5734 , P1_U3447 , P1_R1165_U86 );
nand NAND2_2702 ( P1_U5398 , P1_U3448 , P1_U3442 );
nand NAND2_2703 ( P1_U5399 , P1_U3893 , P1_U4003 );
nand NAND2_2704 ( P1_U5400 , P1_U3369 , P1_U3419 );
nand NAND3_2705 ( P1_U5401 , P1_U3367 , P1_U3362 , P1_U3364 );
nand NAND2_2706 ( P1_U5402 , P1_U4033 , P1_U3421 );
nand NAND2_2707 ( P1_U5403 , P1_U5401 , P1_U3421 );
not NOT1_2708 ( P1_U5404 , P1_U3435 );
nand NAND2_2709 ( P1_U5405 , P1_U5404 , P1_U4003 );
nand NAND2_2710 ( P1_U5406 , P1_U3480 , P1_U5405 );
nand NAND2_2711 ( P1_U5407 , P1_U3021 , P1_U3081 );
nand NAND2_2712 ( P1_U5408 , P1_U3477 , P1_U5405 );
nand NAND2_2713 ( P1_U5409 , P1_U3021 , P1_U3082 );
nand NAND2_2714 ( P1_U5410 , P1_U3474 , P1_U5405 );
nand NAND2_2715 ( P1_U5411 , P1_U3021 , P1_U3068 );
nand NAND2_2716 ( P1_U5412 , P1_U3471 , P1_U5405 );
nand NAND2_2717 ( P1_U5413 , P1_U3021 , P1_U3069 );
nand NAND2_2718 ( P1_U5414 , P1_U3468 , P1_U5405 );
nand NAND2_2719 ( P1_U5415 , P1_U3021 , P1_U3065 );
nand NAND2_2720 ( P1_U5416 , P1_U3465 , P1_U5405 );
nand NAND2_2721 ( P1_U5417 , P1_U3021 , P1_U3058 );
nand NAND2_2722 ( P1_U5418 , P1_U3462 , P1_U5405 );
nand NAND2_2723 ( P1_U5419 , P1_U3021 , P1_U3062 );
nand NAND2_2724 ( P1_U5420 , P1_U4007 , P1_U5405 );
nand NAND2_2725 ( P1_U5421 , P1_U3021 , P1_U3052 );
nand NAND2_2726 ( P1_U5422 , P1_U4008 , P1_U5405 );
nand NAND2_2727 ( P1_U5423 , P1_U3021 , P1_U3051 );
nand NAND2_2728 ( P1_U5424 , P1_U4009 , P1_U5405 );
nand NAND2_2729 ( P1_U5425 , P1_U3021 , P1_U3055 );
nand NAND2_2730 ( P1_U5426 , P1_U4010 , P1_U5405 );
nand NAND2_2731 ( P1_U5427 , P1_U3021 , P1_U3056 );
nand NAND2_2732 ( P1_U5428 , P1_U4011 , P1_U5405 );
nand NAND2_2733 ( P1_U5429 , P1_U3021 , P1_U3063 );
nand NAND2_2734 ( P1_U5430 , P1_U4012 , P1_U5405 );
nand NAND2_2735 ( P1_U5431 , P1_U3021 , P1_U3064 );
nand NAND2_2736 ( P1_U5432 , P1_U4013 , P1_U5405 );
nand NAND2_2737 ( P1_U5433 , P1_U3021 , P1_U3059 );
nand NAND2_2738 ( P1_U5434 , P1_U4014 , P1_U5405 );
nand NAND2_2739 ( P1_U5435 , P1_U3021 , P1_U3073 );
nand NAND2_2740 ( P1_U5436 , P1_U4015 , P1_U5405 );
nand NAND2_2741 ( P1_U5437 , P1_U3021 , P1_U3074 );
nand NAND2_2742 ( P1_U5438 , P1_U3459 , P1_U5405 );
nand NAND2_2743 ( P1_U5439 , P1_U3021 , P1_U3066 );
nand NAND2_2744 ( P1_U5440 , P1_U3509 , P1_U5405 );
nand NAND2_2745 ( P1_U5441 , P1_U3021 , P1_U3079 );
nand NAND2_2746 ( P1_U5442 , P1_U3507 , P1_U5405 );
nand NAND2_2747 ( P1_U5443 , P1_U3021 , P1_U3080 );
nand NAND2_2748 ( P1_U5444 , P1_U3504 , P1_U5405 );
nand NAND2_2749 ( P1_U5445 , P1_U3021 , P1_U3067 );
nand NAND2_2750 ( P1_U5446 , P1_U3501 , P1_U5405 );
nand NAND2_2751 ( P1_U5447 , P1_U3021 , P1_U3071 );
nand NAND2_2752 ( P1_U5448 , P1_U3498 , P1_U5405 );
nand NAND2_2753 ( P1_U5449 , P1_U3021 , P1_U3072 );
nand NAND2_2754 ( P1_U5450 , P1_U3495 , P1_U5405 );
nand NAND2_2755 ( P1_U5451 , P1_U3021 , P1_U3077 );
nand NAND2_2756 ( P1_U5452 , P1_U3492 , P1_U5405 );
nand NAND2_2757 ( P1_U5453 , P1_U3021 , P1_U3078 );
nand NAND2_2758 ( P1_U5454 , P1_U3489 , P1_U5405 );
nand NAND2_2759 ( P1_U5455 , P1_U3021 , P1_U3070 );
nand NAND2_2760 ( P1_U5456 , P1_U3486 , P1_U5405 );
nand NAND2_2761 ( P1_U5457 , P1_U3021 , P1_U3061 );
nand NAND2_2762 ( P1_U5458 , P1_U3483 , P1_U5405 );
nand NAND2_2763 ( P1_U5459 , P1_U3021 , P1_U3060 );
nand NAND2_2764 ( P1_U5460 , P1_U3456 , P1_U5405 );
nand NAND2_2765 ( P1_U5461 , P1_U3021 , P1_U3076 );
nand NAND2_2766 ( P1_U5462 , P1_U3451 , P1_U5405 );
nand NAND2_2767 ( P1_U5463 , P1_U3021 , P1_U3075 );
nand NAND2_2768 ( P1_U5464 , P1_U4135 , P1_REG1_REG_0_ );
nand NAND2_2769 ( P1_U5465 , P1_U3021 , P1_U3480 );
nand NAND2_2770 ( P1_U5466 , P1_U3435 , P1_U3081 );
nand NAND2_2771 ( P1_U5467 , P1_U3021 , P1_U3477 );
nand NAND2_2772 ( P1_U5468 , P1_U3435 , P1_U3082 );
nand NAND2_2773 ( P1_U5469 , P1_U3021 , P1_U3474 );
nand NAND2_2774 ( P1_U5470 , P1_U3435 , P1_U3068 );
nand NAND2_2775 ( P1_U5471 , P1_U3021 , P1_U3471 );
nand NAND2_2776 ( P1_U5472 , P1_U3435 , P1_U3069 );
nand NAND2_2777 ( P1_U5473 , P1_U3021 , P1_U3468 );
nand NAND2_2778 ( P1_U5474 , P1_U3435 , P1_U3065 );
nand NAND2_2779 ( P1_U5475 , P1_U3021 , P1_U3465 );
nand NAND2_2780 ( P1_U5476 , P1_U3435 , P1_U3058 );
nand NAND2_2781 ( P1_U5477 , P1_U3021 , P1_U3462 );
nand NAND2_2782 ( P1_U5478 , P1_U3435 , P1_U3062 );
nand NAND2_2783 ( P1_U5479 , P1_U3021 , P1_U4007 );
nand NAND2_2784 ( P1_U5480 , P1_U3435 , P1_U3052 );
nand NAND2_2785 ( P1_U5481 , P1_U3021 , P1_U4008 );
nand NAND2_2786 ( P1_U5482 , P1_U3435 , P1_U3051 );
nand NAND2_2787 ( P1_U5483 , P1_U3021 , P1_U4009 );
nand NAND2_2788 ( P1_U5484 , P1_U3435 , P1_U3055 );
nand NAND2_2789 ( P1_U5485 , P1_U3021 , P1_U4010 );
nand NAND2_2790 ( P1_U5486 , P1_U3435 , P1_U3056 );
nand NAND2_2791 ( P1_U5487 , P1_U3021 , P1_U4011 );
nand NAND2_2792 ( P1_U5488 , P1_U3435 , P1_U3063 );
nand NAND2_2793 ( P1_U5489 , P1_U3021 , P1_U4012 );
nand NAND2_2794 ( P1_U5490 , P1_U3435 , P1_U3064 );
nand NAND2_2795 ( P1_U5491 , P1_U3021 , P1_U4013 );
nand NAND2_2796 ( P1_U5492 , P1_U3435 , P1_U3059 );
nand NAND2_2797 ( P1_U5493 , P1_U3021 , P1_U4014 );
nand NAND2_2798 ( P1_U5494 , P1_U3435 , P1_U3073 );
nand NAND2_2799 ( P1_U5495 , P1_U3021 , P1_U4015 );
nand NAND2_2800 ( P1_U5496 , P1_U3435 , P1_U3074 );
nand NAND2_2801 ( P1_U5497 , P1_U3021 , P1_U3459 );
nand NAND2_2802 ( P1_U5498 , P1_U3435 , P1_U3066 );
nand NAND2_2803 ( P1_U5499 , P1_U3021 , P1_U3509 );
nand NAND2_2804 ( P1_U5500 , P1_U3435 , P1_U3079 );
nand NAND2_2805 ( P1_U5501 , P1_U3021 , P1_U3507 );
nand NAND2_2806 ( P1_U5502 , P1_U3435 , P1_U3080 );
nand NAND2_2807 ( P1_U5503 , P1_U3021 , P1_U3504 );
nand NAND2_2808 ( P1_U5504 , P1_U3435 , P1_U3067 );
nand NAND2_2809 ( P1_U5505 , P1_U3021 , P1_U3501 );
nand NAND2_2810 ( P1_U5506 , P1_U3435 , P1_U3071 );
nand NAND2_2811 ( P1_U5507 , P1_U3021 , P1_U3498 );
nand NAND2_2812 ( P1_U5508 , P1_U3435 , P1_U3072 );
nand NAND2_2813 ( P1_U5509 , P1_U3021 , P1_U3495 );
nand NAND2_2814 ( P1_U5510 , P1_U3435 , P1_U3077 );
nand NAND2_2815 ( P1_U5511 , P1_U3021 , P1_U3492 );
nand NAND2_2816 ( P1_U5512 , P1_U3435 , P1_U3078 );
nand NAND2_2817 ( P1_U5513 , P1_U3021 , P1_U3489 );
nand NAND2_2818 ( P1_U5514 , P1_U3435 , P1_U3070 );
nand NAND2_2819 ( P1_U5515 , P1_U3021 , P1_U3486 );
nand NAND2_2820 ( P1_U5516 , P1_U3435 , P1_U3061 );
nand NAND2_2821 ( P1_U5517 , P1_U3021 , P1_U3483 );
nand NAND2_2822 ( P1_U5518 , P1_U3435 , P1_U3060 );
nand NAND2_2823 ( P1_U5519 , P1_U3021 , P1_U3456 );
nand NAND2_2824 ( P1_U5520 , P1_U3435 , P1_U3076 );
nand NAND2_2825 ( P1_U5521 , P1_U3021 , P1_U3451 );
nand NAND2_2826 ( P1_U5522 , P1_U3435 , P1_U3075 );
nand NAND2_2827 ( P1_U5523 , P1_U4135 , P1_U3449 );
nand NAND2_2828 ( P1_U5524 , P1_U3428 , P1_U3426 );
nand NAND2_2829 ( P1_U5525 , P1_U3986 , P1_U3480 );
nand NAND2_2830 ( P1_U5526 , P1_U3587 , P1_U5524 );
nand NAND2_2831 ( P1_U5527 , P1_U3986 , P1_U3477 );
nand NAND2_2832 ( P1_U5528 , P1_U3588 , P1_U5524 );
nand NAND2_2833 ( P1_U5529 , P1_U3986 , P1_U3474 );
nand NAND2_2834 ( P1_U5530 , P1_U3589 , P1_U5524 );
nand NAND2_2835 ( P1_U5531 , P1_U3986 , P1_U3471 );
nand NAND2_2836 ( P1_U5532 , P1_U3590 , P1_U5524 );
nand NAND2_2837 ( P1_U5533 , P1_U3986 , P1_U3468 );
nand NAND2_2838 ( P1_U5534 , P1_U3591 , P1_U5524 );
nand NAND2_2839 ( P1_U5535 , P1_U3986 , P1_U3465 );
nand NAND2_2840 ( P1_U5536 , P1_U3592 , P1_U5524 );
nand NAND2_2841 ( P1_U5537 , P1_U3594 , P1_U5524 );
nand NAND2_2842 ( P1_U5538 , P1_U4016 , P1_U3986 );
nand NAND2_2843 ( P1_U5539 , P1_U3595 , P1_U5524 );
nand NAND2_2844 ( P1_U5540 , P1_U4017 , P1_U3986 );
nand NAND2_2845 ( P1_U5541 , P1_U3986 , P1_U3462 );
nand NAND2_2846 ( P1_U5542 , P1_U3593 , P1_U5524 );
nand NAND2_2847 ( P1_U5543 , P1_U3597 , P1_U5524 );
nand NAND2_2848 ( P1_U5544 , P1_U4018 , P1_U3986 );
nand NAND2_2849 ( P1_U5545 , P1_U3598 , P1_U5524 );
nand NAND2_2850 ( P1_U5546 , P1_U4007 , P1_U3986 );
nand NAND2_2851 ( P1_U5547 , P1_U3599 , P1_U5524 );
nand NAND2_2852 ( P1_U5548 , P1_U4008 , P1_U3986 );
nand NAND2_2853 ( P1_U5549 , P1_U3600 , P1_U5524 );
nand NAND2_2854 ( P1_U5550 , P1_U4009 , P1_U3986 );
nand NAND2_2855 ( P1_U5551 , P1_U3601 , P1_U5524 );
nand NAND2_2856 ( P1_U5552 , P1_U4010 , P1_U3986 );
nand NAND2_2857 ( P1_U5553 , P1_U3602 , P1_U5524 );
nand NAND2_2858 ( P1_U5554 , P1_U4011 , P1_U3986 );
nand NAND2_2859 ( P1_U5555 , P1_U3603 , P1_U5524 );
nand NAND2_2860 ( P1_U5556 , P1_U4012 , P1_U3986 );
nand NAND2_2861 ( P1_U5557 , P1_U3604 , P1_U5524 );
nand NAND2_2862 ( P1_U5558 , P1_U4013 , P1_U3986 );
nand NAND2_2863 ( P1_U5559 , P1_U3605 , P1_U5524 );
nand NAND2_2864 ( P1_U5560 , P1_U4014 , P1_U3986 );
nand NAND2_2865 ( P1_U5561 , P1_U3606 , P1_U5524 );
nand NAND2_2866 ( P1_U5562 , P1_U4015 , P1_U3986 );
nand NAND2_2867 ( P1_U5563 , P1_U3986 , P1_U3459 );
nand NAND2_2868 ( P1_U5564 , P1_U3596 , P1_U5524 );
nand NAND2_2869 ( P1_U5565 , P1_U3986 , P1_U3509 );
nand NAND2_2870 ( P1_U5566 , P1_U3608 , P1_U5524 );
nand NAND2_2871 ( P1_U5567 , P1_U3986 , P1_U3507 );
nand NAND2_2872 ( P1_U5568 , P1_U3609 , P1_U5524 );
nand NAND2_2873 ( P1_U5569 , P1_U3986 , P1_U3504 );
nand NAND2_2874 ( P1_U5570 , P1_U3610 , P1_U5524 );
nand NAND2_2875 ( P1_U5571 , P1_U3986 , P1_U3501 );
nand NAND2_2876 ( P1_U5572 , P1_U3611 , P1_U5524 );
nand NAND2_2877 ( P1_U5573 , P1_U3986 , P1_U3498 );
nand NAND2_2878 ( P1_U5574 , P1_U3612 , P1_U5524 );
nand NAND2_2879 ( P1_U5575 , P1_U3986 , P1_U3495 );
nand NAND2_2880 ( P1_U5576 , P1_U3613 , P1_U5524 );
nand NAND2_2881 ( P1_U5577 , P1_U3986 , P1_U3492 );
nand NAND2_2882 ( P1_U5578 , P1_U3614 , P1_U5524 );
nand NAND2_2883 ( P1_U5579 , P1_U3986 , P1_U3489 );
nand NAND2_2884 ( P1_U5580 , P1_U3615 , P1_U5524 );
nand NAND2_2885 ( P1_U5581 , P1_U3986 , P1_U3486 );
nand NAND2_2886 ( P1_U5582 , P1_U3616 , P1_U5524 );
nand NAND2_2887 ( P1_U5583 , P1_U3986 , P1_U3483 );
nand NAND2_2888 ( P1_U5584 , P1_U3617 , P1_U5524 );
nand NAND2_2889 ( P1_U5585 , P1_U3986 , P1_U3456 );
nand NAND2_2890 ( P1_U5586 , P1_U3607 , P1_U5524 );
nand NAND2_2891 ( P1_U5587 , P1_U3986 , P1_U3451 );
nand NAND2_2892 ( P1_U5588 , P1_U3618 , P1_U5524 );
nand NAND2_2893 ( P1_U5589 , P1_U3480 , P1_U5524 );
nand NAND2_2894 ( P1_U5590 , P1_U3986 , P1_U3587 );
nand NAND2_2895 ( P1_U5591 , P1_U5703 , P1_U3082 );
nand NAND2_2896 ( P1_U5592 , P1_U3477 , P1_U5524 );
nand NAND2_2897 ( P1_U5593 , P1_U3986 , P1_U3588 );
nand NAND2_2898 ( P1_U5594 , P1_U5703 , P1_U3068 );
nand NAND2_2899 ( P1_U5595 , P1_U3474 , P1_U5524 );
nand NAND2_2900 ( P1_U5596 , P1_U3986 , P1_U3589 );
nand NAND2_2901 ( P1_U5597 , P1_U5703 , P1_U3069 );
nand NAND2_2902 ( P1_U5598 , P1_U3471 , P1_U5524 );
nand NAND2_2903 ( P1_U5599 , P1_U3986 , P1_U3590 );
nand NAND2_2904 ( P1_U5600 , P1_U5703 , P1_U3065 );
nand NAND2_2905 ( P1_U5601 , P1_U3468 , P1_U5524 );
nand NAND2_2906 ( P1_U5602 , P1_U3986 , P1_U3591 );
nand NAND2_2907 ( P1_U5603 , P1_U5703 , P1_U3058 );
nand NAND2_2908 ( P1_U5604 , P1_U3465 , P1_U5524 );
nand NAND2_2909 ( P1_U5605 , P1_U3986 , P1_U3592 );
nand NAND2_2910 ( P1_U5606 , P1_U5703 , P1_U3062 );
nand NAND2_2911 ( P1_U5607 , P1_U4016 , P1_U5524 );
nand NAND2_2912 ( P1_U5608 , P1_U3986 , P1_U3594 );
nand NAND2_2913 ( P1_U5609 , P1_U4017 , P1_U5524 );
nand NAND2_2914 ( P1_U5610 , P1_U3986 , P1_U3595 );
nand NAND2_2915 ( P1_U5611 , P1_U3462 , P1_U5524 );
nand NAND2_2916 ( P1_U5612 , P1_U3986 , P1_U3593 );
nand NAND2_2917 ( P1_U5613 , P1_U5703 , P1_U3066 );
nand NAND2_2918 ( P1_U5614 , P1_U4018 , P1_U5524 );
nand NAND2_2919 ( P1_U5615 , P1_U3986 , P1_U3597 );
nand NAND2_2920 ( P1_U5616 , P1_U5703 , P1_U3052 );
nand NAND2_2921 ( P1_U5617 , P1_U4007 , P1_U5524 );
nand NAND2_2922 ( P1_U5618 , P1_U3986 , P1_U3598 );
nand NAND2_2923 ( P1_U5619 , P1_U5703 , P1_U3051 );
nand NAND2_2924 ( P1_U5620 , P1_U4008 , P1_U5524 );
nand NAND2_2925 ( P1_U5621 , P1_U3986 , P1_U3599 );
nand NAND2_2926 ( P1_U5622 , P1_U5703 , P1_U3055 );
nand NAND2_2927 ( P1_U5623 , P1_U4009 , P1_U5524 );
nand NAND2_2928 ( P1_U5624 , P1_U3986 , P1_U3600 );
nand NAND2_2929 ( P1_U5625 , P1_U5703 , P1_U3056 );
nand NAND2_2930 ( P1_U5626 , P1_U4010 , P1_U5524 );
nand NAND2_2931 ( P1_U5627 , P1_U3986 , P1_U3601 );
nand NAND2_2932 ( P1_U5628 , P1_U5703 , P1_U3063 );
nand NAND2_2933 ( P1_U5629 , P1_U4011 , P1_U5524 );
nand NAND2_2934 ( P1_U5630 , P1_U3986 , P1_U3602 );
nand NAND2_2935 ( P1_U5631 , P1_U5703 , P1_U3064 );
nand NAND2_2936 ( P1_U5632 , P1_U4012 , P1_U5524 );
nand NAND2_2937 ( P1_U5633 , P1_U3986 , P1_U3603 );
nand NAND2_2938 ( P1_U5634 , P1_U5703 , P1_U3059 );
nand NAND2_2939 ( P1_U5635 , P1_U4013 , P1_U5524 );
nand NAND2_2940 ( P1_U5636 , P1_U3986 , P1_U3604 );
nand NAND2_2941 ( P1_U5637 , P1_U5703 , P1_U3073 );
nand NAND2_2942 ( P1_U5638 , P1_U4014 , P1_U5524 );
nand NAND2_2943 ( P1_U5639 , P1_U3986 , P1_U3605 );
nand NAND2_2944 ( P1_U5640 , P1_U5703 , P1_U3074 );
nand NAND2_2945 ( P1_U5641 , P1_U4015 , P1_U5524 );
nand NAND2_2946 ( P1_U5642 , P1_U3986 , P1_U3606 );
nand NAND2_2947 ( P1_U5643 , P1_U5703 , P1_U3079 );
nand NAND2_2948 ( P1_U5644 , P1_U3459 , P1_U5524 );
nand NAND2_2949 ( P1_U5645 , P1_U3986 , P1_U3596 );
nand NAND2_2950 ( P1_U5646 , P1_U5703 , P1_U3076 );
nand NAND2_2951 ( P1_U5647 , P1_U3509 , P1_U5524 );
nand NAND2_2952 ( P1_U5648 , P1_U3986 , P1_U3608 );
nand NAND2_2953 ( P1_U5649 , P1_U5703 , P1_U3080 );
nand NAND2_2954 ( P1_U5650 , P1_U3507 , P1_U5524 );
nand NAND2_2955 ( P1_U5651 , P1_U3986 , P1_U3609 );
nand NAND2_2956 ( P1_U5652 , P1_U5703 , P1_U3067 );
nand NAND2_2957 ( P1_U5653 , P1_U3504 , P1_U5524 );
nand NAND2_2958 ( P1_U5654 , P1_U3986 , P1_U3610 );
nand NAND2_2959 ( P1_U5655 , P1_U5703 , P1_U3071 );
nand NAND2_2960 ( P1_U5656 , P1_U3501 , P1_U5524 );
nand NAND2_2961 ( P1_U5657 , P1_U3986 , P1_U3611 );
nand NAND2_2962 ( P1_U5658 , P1_U5703 , P1_U3072 );
nand NAND2_2963 ( P1_U5659 , P1_U3498 , P1_U5524 );
nand NAND2_2964 ( P1_U5660 , P1_U3986 , P1_U3612 );
nand NAND2_2965 ( P1_U5661 , P1_U5703 , P1_U3077 );
nand NAND2_2966 ( P1_U5662 , P1_U3495 , P1_U5524 );
nand NAND2_2967 ( P1_U5663 , P1_U3986 , P1_U3613 );
nand NAND2_2968 ( P1_U5664 , P1_U5703 , P1_U3078 );
nand NAND2_2969 ( P1_U5665 , P1_U3492 , P1_U5524 );
nand NAND2_2970 ( P1_U5666 , P1_U3986 , P1_U3614 );
nand NAND2_2971 ( P1_U5667 , P1_U5703 , P1_U3070 );
nand NAND2_2972 ( P1_U5668 , P1_U3489 , P1_U5524 );
nand NAND2_2973 ( P1_U5669 , P1_U3986 , P1_U3615 );
nand NAND2_2974 ( P1_U5670 , P1_U5703 , P1_U3061 );
nand NAND2_2975 ( P1_U5671 , P1_U3486 , P1_U5524 );
nand NAND2_2976 ( P1_U5672 , P1_U3986 , P1_U3616 );
nand NAND2_2977 ( P1_U5673 , P1_U5703 , P1_U3060 );
nand NAND2_2978 ( P1_U5674 , P1_U3483 , P1_U5524 );
nand NAND2_2979 ( P1_U5675 , P1_U3986 , P1_U3617 );
nand NAND2_2980 ( P1_U5676 , P1_U5703 , P1_U3081 );
nand NAND2_2981 ( P1_U5677 , P1_U3456 , P1_U5524 );
nand NAND2_2982 ( P1_U5678 , P1_U3986 , P1_U3607 );
nand NAND2_2983 ( P1_U5679 , P1_U5703 , P1_U3075 );
nand NAND2_2984 ( P1_U5680 , P1_U3451 , P1_U5524 );
nand NAND2_2985 ( P1_U5681 , P1_U3986 , P1_U3618 );
nand NAND2_2986 ( P1_U5682 , P1_U5123 , P1_U3084 );
nand NAND2_2987 ( P1_U5683 , P1_U4030 , P1_U3431 );
nand NAND2_2988 ( P1_U5684 , P1_U4005 , P1_U4030 );
nand NAND2_2989 ( P1_U5685 , P1_U5683 , P1_U4028 );
nand NAND2_2990 ( P1_U5686 , P1_U5684 , P1_U4029 );
nand NAND3_2991 ( P1_U5687 , P1_U3439 , P1_U3048 , P1_U3429 );
nand NAND2_2992 ( P1_U5688 , P1_U5692 , P1_U5698 );
nand NAND4_2993 ( P1_U5689 , P1_U4020 , P1_U3442 , P1_U3987 , P1_LT_201_U14 );
nand NAND2_2994 ( P1_U5690 , P1_IR_REG_24_ , P1_U3944 );
nand NAND2_2995 ( P1_U5691 , P1_IR_REG_31_ , P1_SUB_88_U17 );
not NOT1_2996 ( P1_U5692 , P1_U3436 );
nand NAND2_2997 ( P1_U5693 , P1_IR_REG_25_ , P1_U3944 );
nand NAND2_2998 ( P1_U5694 , P1_IR_REG_31_ , P1_SUB_88_U170 );
not NOT1_2999 ( P1_U5695 , P1_U3437 );
nand NAND2_3000 ( P1_U5696 , P1_IR_REG_26_ , P1_U3944 );
nand NAND2_3001 ( P1_U5697 , P1_IR_REG_31_ , P1_SUB_88_U18 );
not NOT1_3002 ( P1_U5698 , P1_U3438 );
nand NAND2_3003 ( P1_U5699 , P1_U3050 , P1_U3358 );
nand NAND3_3004 ( P1_U5700 , P1_U4036 , P1_U5692 , P1_B_REG );
nand NAND2_3005 ( P1_U5701 , P1_IR_REG_23_ , P1_U3944 );
nand NAND2_3006 ( P1_U5702 , P1_IR_REG_31_ , P1_SUB_88_U16 );
not NOT1_3007 ( P1_U5703 , P1_U3439 );
nand NAND2_3008 ( P1_U5704 , P1_D_REG_0_ , P1_U3945 );
nand NAND2_3009 ( P1_U5705 , P1_U4025 , P1_U4136 );
nand NAND2_3010 ( P1_U5706 , P1_D_REG_1_ , P1_U3945 );
nand NAND2_3011 ( P1_U5707 , P1_U4025 , P1_U4137 );
nand NAND2_3012 ( P1_U5708 , P1_IR_REG_22_ , P1_U3944 );
nand NAND2_3013 ( P1_U5709 , P1_IR_REG_31_ , P1_SUB_88_U15 );
not NOT1_3014 ( P1_U5710 , P1_U3444 );
nand NAND2_3015 ( P1_U5711 , P1_IR_REG_19_ , P1_U3944 );
nand NAND2_3016 ( P1_U5712 , P1_IR_REG_31_ , P1_SUB_88_U13 );
not NOT1_3017 ( P1_U5713 , P1_U3443 );
nand NAND2_3018 ( P1_U5714 , P1_IR_REG_20_ , P1_U3944 );
nand NAND2_3019 ( P1_U5715 , P1_IR_REG_31_ , P1_SUB_88_U14 );
not NOT1_3020 ( P1_U5716 , P1_U3442 );
nand NAND2_3021 ( P1_U5717 , P1_IR_REG_21_ , P1_U3944 );
nand NAND2_3022 ( P1_U5718 , P1_IR_REG_31_ , P1_SUB_88_U173 );
not NOT1_3023 ( P1_U5719 , P1_U3448 );
nand NAND2_3024 ( P1_U5720 , P1_IR_REG_30_ , P1_U3944 );
nand NAND2_3025 ( P1_U5721 , P1_IR_REG_31_ , P1_SUB_88_U165 );
not NOT1_3026 ( P1_U5722 , P1_U3445 );
nand NAND2_3027 ( P1_U5723 , P1_IR_REG_29_ , P1_U3944 );
nand NAND2_3028 ( P1_U5724 , P1_IR_REG_31_ , P1_SUB_88_U20 );
not NOT1_3029 ( P1_U5725 , P1_U3446 );
nand NAND2_3030 ( P1_U5726 , P1_IR_REG_28_ , P1_U3944 );
nand NAND2_3031 ( P1_U5727 , P1_IR_REG_31_ , P1_SUB_88_U19 );
not NOT1_3032 ( P1_U5728 , P1_U3447 );
nand NAND2_3033 ( P1_U5729 , P1_IR_REG_0_ , P1_U3944 );
nand NAND2_3034 ( P1_U5730 , P1_IR_REG_31_ , P1_IR_REG_0_ );
not NOT1_3035 ( P1_U5731 , P1_U3449 );
nand NAND2_3036 ( P1_U5732 , P1_IR_REG_27_ , P1_U3944 );
nand NAND2_3037 ( P1_U5733 , P1_IR_REG_31_ , P1_SUB_88_U42 );
not NOT1_3038 ( P1_U5734 , P1_U3450 );
nand NAND2_3039 ( P1_U5735 , U88 , P1_U3946 );
nand NAND2_3040 ( P1_U5736 , P1_U4004 , P1_U3449 );
not NOT1_3041 ( P1_U5737 , P1_U3451 );
nand NAND2_3042 ( P1_U5738 , P1_U3444 , P1_U5719 );
nand NAND2_3043 ( P1_U5739 , P1_U5710 , P1_U4168 );
nand NAND2_3044 ( P1_U5740 , P1_D_REG_1_ , P1_U4134 );
nand NAND2_3045 ( P1_U5741 , P1_U4137 , P1_U3359 );
not NOT1_3046 ( P1_U5742 , P1_U3453 );
nand NAND2_3047 ( P1_U5743 , P1_U5688 , P1_U3359 );
nand NAND2_3048 ( P1_U5744 , P1_D_REG_0_ , P1_U4134 );
not NOT1_3049 ( P1_U5745 , P1_U3452 );
nand NAND2_3050 ( P1_U5746 , P1_REG0_REG_0_ , P1_U3947 );
nand NAND2_3051 ( P1_U5747 , P1_U4024 , P1_U4188 );
nand NAND2_3052 ( P1_U5748 , P1_IR_REG_1_ , P1_U3944 );
nand NAND2_3053 ( P1_U5749 , P1_IR_REG_31_ , P1_SUB_88_U40 );
nand NAND2_3054 ( P1_U5750 , U77 , P1_U3946 );
nand NAND2_3055 ( P1_U5751 , P1_U3455 , P1_U4004 );
not NOT1_3056 ( P1_U5752 , P1_U3456 );
nand NAND2_3057 ( P1_U5753 , P1_REG0_REG_1_ , P1_U3947 );
nand NAND2_3058 ( P1_U5754 , P1_U4024 , P1_U4212 );
nand NAND2_3059 ( P1_U5755 , P1_IR_REG_2_ , P1_U3944 );
nand NAND2_3060 ( P1_U5756 , P1_IR_REG_31_ , P1_SUB_88_U21 );
nand NAND2_3061 ( P1_U5757 , U66 , P1_U3946 );
nand NAND2_3062 ( P1_U5758 , P1_U3458 , P1_U4004 );
not NOT1_3063 ( P1_U5759 , P1_U3459 );
nand NAND2_3064 ( P1_U5760 , P1_REG0_REG_2_ , P1_U3947 );
nand NAND2_3065 ( P1_U5761 , P1_U4024 , P1_U4231 );
nand NAND2_3066 ( P1_U5762 , P1_IR_REG_3_ , P1_U3944 );
nand NAND2_3067 ( P1_U5763 , P1_IR_REG_31_ , P1_SUB_88_U22 );
nand NAND2_3068 ( P1_U5764 , U63 , P1_U3946 );
nand NAND2_3069 ( P1_U5765 , P1_U3461 , P1_U4004 );
not NOT1_3070 ( P1_U5766 , P1_U3462 );
nand NAND2_3071 ( P1_U5767 , P1_REG0_REG_3_ , P1_U3947 );
nand NAND2_3072 ( P1_U5768 , P1_U4024 , P1_U4250 );
nand NAND2_3073 ( P1_U5769 , P1_IR_REG_4_ , P1_U3944 );
nand NAND2_3074 ( P1_U5770 , P1_IR_REG_31_ , P1_SUB_88_U23 );
nand NAND2_3075 ( P1_U5771 , U62 , P1_U3946 );
nand NAND2_3076 ( P1_U5772 , P1_U3464 , P1_U4004 );
not NOT1_3077 ( P1_U5773 , P1_U3465 );
nand NAND2_3078 ( P1_U5774 , P1_REG0_REG_4_ , P1_U3947 );
nand NAND2_3079 ( P1_U5775 , P1_U4024 , P1_U4269 );
nand NAND2_3080 ( P1_U5776 , P1_IR_REG_5_ , P1_U3944 );
nand NAND2_3081 ( P1_U5777 , P1_IR_REG_31_ , P1_SUB_88_U162 );
nand NAND2_3082 ( P1_U5778 , U61 , P1_U3946 );
nand NAND2_3083 ( P1_U5779 , P1_U3467 , P1_U4004 );
not NOT1_3084 ( P1_U5780 , P1_U3468 );
nand NAND2_3085 ( P1_U5781 , P1_REG0_REG_5_ , P1_U3947 );
nand NAND2_3086 ( P1_U5782 , P1_U4024 , P1_U4288 );
nand NAND2_3087 ( P1_U5783 , P1_IR_REG_6_ , P1_U3944 );
nand NAND2_3088 ( P1_U5784 , P1_IR_REG_31_ , P1_SUB_88_U24 );
nand NAND2_3089 ( P1_U5785 , U60 , P1_U3946 );
nand NAND2_3090 ( P1_U5786 , P1_U3470 , P1_U4004 );
not NOT1_3091 ( P1_U5787 , P1_U3471 );
nand NAND2_3092 ( P1_U5788 , P1_REG0_REG_6_ , P1_U3947 );
nand NAND2_3093 ( P1_U5789 , P1_U4024 , P1_U4307 );
nand NAND2_3094 ( P1_U5790 , P1_IR_REG_7_ , P1_U3944 );
nand NAND2_3095 ( P1_U5791 , P1_IR_REG_31_ , P1_SUB_88_U25 );
nand NAND2_3096 ( P1_U5792 , U59 , P1_U3946 );
nand NAND2_3097 ( P1_U5793 , P1_U3473 , P1_U4004 );
not NOT1_3098 ( P1_U5794 , P1_U3474 );
nand NAND2_3099 ( P1_U5795 , P1_REG0_REG_7_ , P1_U3947 );
nand NAND2_3100 ( P1_U5796 , P1_U4024 , P1_U4326 );
nand NAND2_3101 ( P1_U5797 , P1_IR_REG_8_ , P1_U3944 );
nand NAND2_3102 ( P1_U5798 , P1_IR_REG_31_ , P1_SUB_88_U26 );
nand NAND2_3103 ( P1_U5799 , U58 , P1_U3946 );
nand NAND2_3104 ( P1_U5800 , P1_U3476 , P1_U4004 );
not NOT1_3105 ( P1_U5801 , P1_U3477 );
nand NAND2_3106 ( P1_U5802 , P1_REG0_REG_8_ , P1_U3947 );
nand NAND2_3107 ( P1_U5803 , P1_U4024 , P1_U4345 );
nand NAND2_3108 ( P1_U5804 , P1_IR_REG_9_ , P1_U3944 );
nand NAND2_3109 ( P1_U5805 , P1_IR_REG_31_ , P1_SUB_88_U160 );
nand NAND2_3110 ( P1_U5806 , U57 , P1_U3946 );
nand NAND2_3111 ( P1_U5807 , P1_U3479 , P1_U4004 );
not NOT1_3112 ( P1_U5808 , P1_U3480 );
nand NAND2_3113 ( P1_U5809 , P1_REG0_REG_9_ , P1_U3947 );
nand NAND2_3114 ( P1_U5810 , P1_U4024 , P1_U4364 );
nand NAND2_3115 ( P1_U5811 , P1_IR_REG_10_ , P1_U3944 );
nand NAND2_3116 ( P1_U5812 , P1_IR_REG_31_ , P1_SUB_88_U6 );
nand NAND2_3117 ( P1_U5813 , U87 , P1_U3946 );
nand NAND2_3118 ( P1_U5814 , P1_U3482 , P1_U4004 );
not NOT1_3119 ( P1_U5815 , P1_U3483 );
nand NAND2_3120 ( P1_U5816 , P1_REG0_REG_10_ , P1_U3947 );
nand NAND2_3121 ( P1_U5817 , P1_U4024 , P1_U4383 );
nand NAND2_3122 ( P1_U5818 , P1_IR_REG_11_ , P1_U3944 );
nand NAND2_3123 ( P1_U5819 , P1_IR_REG_31_ , P1_SUB_88_U7 );
nand NAND2_3124 ( P1_U5820 , U86 , P1_U3946 );
nand NAND2_3125 ( P1_U5821 , P1_U3485 , P1_U4004 );
not NOT1_3126 ( P1_U5822 , P1_U3486 );
nand NAND2_3127 ( P1_U5823 , P1_REG0_REG_11_ , P1_U3947 );
nand NAND2_3128 ( P1_U5824 , P1_U4024 , P1_U4402 );
nand NAND2_3129 ( P1_U5825 , P1_IR_REG_12_ , P1_U3944 );
nand NAND2_3130 ( P1_U5826 , P1_IR_REG_31_ , P1_SUB_88_U8 );
nand NAND2_3131 ( P1_U5827 , U85 , P1_U3946 );
nand NAND2_3132 ( P1_U5828 , P1_U3488 , P1_U4004 );
not NOT1_3133 ( P1_U5829 , P1_U3489 );
nand NAND2_3134 ( P1_U5830 , P1_REG0_REG_12_ , P1_U3947 );
nand NAND2_3135 ( P1_U5831 , P1_U4024 , P1_U4421 );
nand NAND2_3136 ( P1_U5832 , P1_IR_REG_13_ , P1_U3944 );
nand NAND2_3137 ( P1_U5833 , P1_IR_REG_31_ , P1_SUB_88_U179 );
nand NAND2_3138 ( P1_U5834 , U84 , P1_U3946 );
nand NAND2_3139 ( P1_U5835 , P1_U3491 , P1_U4004 );
not NOT1_3140 ( P1_U5836 , P1_U3492 );
nand NAND2_3141 ( P1_U5837 , P1_REG0_REG_13_ , P1_U3947 );
nand NAND2_3142 ( P1_U5838 , P1_U4024 , P1_U4440 );
nand NAND2_3143 ( P1_U5839 , P1_IR_REG_14_ , P1_U3944 );
nand NAND2_3144 ( P1_U5840 , P1_IR_REG_31_ , P1_SUB_88_U9 );
nand NAND2_3145 ( P1_U5841 , U83 , P1_U3946 );
nand NAND2_3146 ( P1_U5842 , P1_U3494 , P1_U4004 );
not NOT1_3147 ( P1_U5843 , P1_U3495 );
nand NAND2_3148 ( P1_U5844 , P1_REG0_REG_14_ , P1_U3947 );
nand NAND2_3149 ( P1_U5845 , P1_U4024 , P1_U4459 );
nand NAND2_3150 ( P1_U5846 , P1_IR_REG_15_ , P1_U3944 );
nand NAND2_3151 ( P1_U5847 , P1_IR_REG_31_ , P1_SUB_88_U10 );
nand NAND2_3152 ( P1_U5848 , U82 , P1_U3946 );
nand NAND2_3153 ( P1_U5849 , P1_U3497 , P1_U4004 );
not NOT1_3154 ( P1_U5850 , P1_U3498 );
nand NAND2_3155 ( P1_U5851 , P1_REG0_REG_15_ , P1_U3947 );
nand NAND2_3156 ( P1_U5852 , P1_U4024 , P1_U4478 );
nand NAND2_3157 ( P1_U5853 , P1_IR_REG_16_ , P1_U3944 );
nand NAND2_3158 ( P1_U5854 , P1_IR_REG_31_ , P1_SUB_88_U11 );
nand NAND2_3159 ( P1_U5855 , U81 , P1_U3946 );
nand NAND2_3160 ( P1_U5856 , P1_U3500 , P1_U4004 );
not NOT1_3161 ( P1_U5857 , P1_U3501 );
nand NAND2_3162 ( P1_U5858 , P1_REG0_REG_16_ , P1_U3947 );
nand NAND2_3163 ( P1_U5859 , P1_U4024 , P1_U4497 );
nand NAND2_3164 ( P1_U5860 , P1_IR_REG_17_ , P1_U3944 );
nand NAND2_3165 ( P1_U5861 , P1_IR_REG_31_ , P1_SUB_88_U177 );
nand NAND2_3166 ( P1_U5862 , U80 , P1_U3946 );
nand NAND2_3167 ( P1_U5863 , P1_U3503 , P1_U4004 );
not NOT1_3168 ( P1_U5864 , P1_U3504 );
nand NAND2_3169 ( P1_U5865 , P1_REG0_REG_17_ , P1_U3947 );
nand NAND2_3170 ( P1_U5866 , P1_U4024 , P1_U4516 );
nand NAND2_3171 ( P1_U5867 , P1_IR_REG_18_ , P1_U3944 );
nand NAND2_3172 ( P1_U5868 , P1_IR_REG_31_ , P1_SUB_88_U12 );
nand NAND2_3173 ( P1_U5869 , U79 , P1_U3946 );
nand NAND2_3174 ( P1_U5870 , P1_U3506 , P1_U4004 );
not NOT1_3175 ( P1_U5871 , P1_U3507 );
nand NAND2_3176 ( P1_U5872 , P1_REG0_REG_18_ , P1_U3947 );
nand NAND2_3177 ( P1_U5873 , P1_U4024 , P1_U4535 );
nand NAND2_3178 ( P1_U5874 , U78 , P1_U3946 );
nand NAND2_3179 ( P1_U5875 , P1_U4004 , P1_U3443 );
not NOT1_3180 ( P1_U5876 , P1_U3509 );
nand NAND2_3181 ( P1_U5877 , P1_REG0_REG_19_ , P1_U3947 );
nand NAND2_3182 ( P1_U5878 , P1_U4024 , P1_U4554 );
nand NAND2_3183 ( P1_U5879 , P1_REG0_REG_20_ , P1_U3947 );
nand NAND2_3184 ( P1_U5880 , P1_U4024 , P1_U4573 );
nand NAND2_3185 ( P1_U5881 , P1_REG0_REG_21_ , P1_U3947 );
nand NAND2_3186 ( P1_U5882 , P1_U4024 , P1_U4592 );
nand NAND2_3187 ( P1_U5883 , P1_REG0_REG_22_ , P1_U3947 );
nand NAND2_3188 ( P1_U5884 , P1_U4024 , P1_U4611 );
nand NAND2_3189 ( P1_U5885 , P1_REG0_REG_23_ , P1_U3947 );
nand NAND2_3190 ( P1_U5886 , P1_U4024 , P1_U4630 );
nand NAND2_3191 ( P1_U5887 , P1_REG0_REG_24_ , P1_U3947 );
nand NAND2_3192 ( P1_U5888 , P1_U4024 , P1_U4649 );
nand NAND2_3193 ( P1_U5889 , P1_REG0_REG_25_ , P1_U3947 );
nand NAND2_3194 ( P1_U5890 , P1_U4024 , P1_U4668 );
nand NAND2_3195 ( P1_U5891 , P1_REG0_REG_26_ , P1_U3947 );
nand NAND2_3196 ( P1_U5892 , P1_U4024 , P1_U4687 );
nand NAND2_3197 ( P1_U5893 , P1_REG0_REG_27_ , P1_U3947 );
nand NAND2_3198 ( P1_U5894 , P1_U4024 , P1_U4706 );
nand NAND2_3199 ( P1_U5895 , P1_REG0_REG_28_ , P1_U3947 );
nand NAND2_3200 ( P1_U5896 , P1_U4024 , P1_U4725 );
nand NAND2_3201 ( P1_U5897 , P1_REG0_REG_29_ , P1_U3947 );
nand NAND2_3202 ( P1_U5898 , P1_U4024 , P1_U4745 );
nand NAND2_3203 ( P1_U5899 , P1_REG0_REG_30_ , P1_U3947 );
nand NAND2_3204 ( P1_U5900 , P1_U4024 , P1_U4752 );
nand NAND2_3205 ( P1_U5901 , P1_REG0_REG_31_ , P1_U3947 );
nand NAND2_3206 ( P1_U5902 , P1_U4024 , P1_U4755 );
nand NAND2_3207 ( P1_U5903 , P1_REG1_REG_0_ , P1_U3948 );
nand NAND2_3208 ( P1_U5904 , P1_U4023 , P1_U4188 );
nand NAND2_3209 ( P1_U5905 , P1_REG1_REG_1_ , P1_U3948 );
nand NAND2_3210 ( P1_U5906 , P1_U4023 , P1_U4212 );
nand NAND2_3211 ( P1_U5907 , P1_REG1_REG_2_ , P1_U3948 );
nand NAND2_3212 ( P1_U5908 , P1_U4023 , P1_U4231 );
nand NAND2_3213 ( P1_U5909 , P1_REG1_REG_3_ , P1_U3948 );
nand NAND2_3214 ( P1_U5910 , P1_U4023 , P1_U4250 );
nand NAND2_3215 ( P1_U5911 , P1_REG1_REG_4_ , P1_U3948 );
nand NAND2_3216 ( P1_U5912 , P1_U4023 , P1_U4269 );
nand NAND2_3217 ( P1_U5913 , P1_REG1_REG_5_ , P1_U3948 );
nand NAND2_3218 ( P1_U5914 , P1_U4023 , P1_U4288 );
nand NAND2_3219 ( P1_U5915 , P1_REG1_REG_6_ , P1_U3948 );
nand NAND2_3220 ( P1_U5916 , P1_U4023 , P1_U4307 );
nand NAND2_3221 ( P1_U5917 , P1_REG1_REG_7_ , P1_U3948 );
nand NAND2_3222 ( P1_U5918 , P1_U4023 , P1_U4326 );
nand NAND2_3223 ( P1_U5919 , P1_REG1_REG_8_ , P1_U3948 );
nand NAND2_3224 ( P1_U5920 , P1_U4023 , P1_U4345 );
nand NAND2_3225 ( P1_U5921 , P1_REG1_REG_9_ , P1_U3948 );
nand NAND2_3226 ( P1_U5922 , P1_U4023 , P1_U4364 );
nand NAND2_3227 ( P1_U5923 , P1_REG1_REG_10_ , P1_U3948 );
nand NAND2_3228 ( P1_U5924 , P1_U4023 , P1_U4383 );
nand NAND2_3229 ( P1_U5925 , P1_REG1_REG_11_ , P1_U3948 );
nand NAND2_3230 ( P1_U5926 , P1_U4023 , P1_U4402 );
nand NAND2_3231 ( P1_U5927 , P1_REG1_REG_12_ , P1_U3948 );
nand NAND2_3232 ( P1_U5928 , P1_U4023 , P1_U4421 );
nand NAND2_3233 ( P1_U5929 , P1_REG1_REG_13_ , P1_U3948 );
nand NAND2_3234 ( P1_U5930 , P1_U4023 , P1_U4440 );
nand NAND2_3235 ( P1_U5931 , P1_REG1_REG_14_ , P1_U3948 );
nand NAND2_3236 ( P1_U5932 , P1_U4023 , P1_U4459 );
nand NAND2_3237 ( P1_U5933 , P1_REG1_REG_15_ , P1_U3948 );
nand NAND2_3238 ( P1_U5934 , P1_U4023 , P1_U4478 );
nand NAND2_3239 ( P1_U5935 , P1_REG1_REG_16_ , P1_U3948 );
nand NAND2_3240 ( P1_U5936 , P1_U4023 , P1_U4497 );
nand NAND2_3241 ( P1_U5937 , P1_REG1_REG_17_ , P1_U3948 );
nand NAND2_3242 ( P1_U5938 , P1_U4023 , P1_U4516 );
nand NAND2_3243 ( P1_U5939 , P1_REG1_REG_18_ , P1_U3948 );
nand NAND2_3244 ( P1_U5940 , P1_U4023 , P1_U4535 );
nand NAND2_3245 ( P1_U5941 , P1_REG1_REG_19_ , P1_U3948 );
nand NAND2_3246 ( P1_U5942 , P1_U4023 , P1_U4554 );
nand NAND2_3247 ( P1_U5943 , P1_REG1_REG_20_ , P1_U3948 );
nand NAND2_3248 ( P1_U5944 , P1_U4023 , P1_U4573 );
nand NAND2_3249 ( P1_U5945 , P1_REG1_REG_21_ , P1_U3948 );
nand NAND2_3250 ( P1_U5946 , P1_U4023 , P1_U4592 );
nand NAND2_3251 ( P1_U5947 , P1_REG1_REG_22_ , P1_U3948 );
nand NAND2_3252 ( P1_U5948 , P1_U4023 , P1_U4611 );
nand NAND2_3253 ( P1_U5949 , P1_REG1_REG_23_ , P1_U3948 );
nand NAND2_3254 ( P1_U5950 , P1_U4023 , P1_U4630 );
nand NAND2_3255 ( P1_U5951 , P1_REG1_REG_24_ , P1_U3948 );
nand NAND2_3256 ( P1_U5952 , P1_U4023 , P1_U4649 );
nand NAND2_3257 ( P1_U5953 , P1_REG1_REG_25_ , P1_U3948 );
nand NAND2_3258 ( P1_U5954 , P1_U4023 , P1_U4668 );
nand NAND2_3259 ( P1_U5955 , P1_REG1_REG_26_ , P1_U3948 );
nand NAND2_3260 ( P1_U5956 , P1_U4023 , P1_U4687 );
nand NAND2_3261 ( P1_U5957 , P1_REG1_REG_27_ , P1_U3948 );
nand NAND2_3262 ( P1_U5958 , P1_U4023 , P1_U4706 );
nand NAND2_3263 ( P1_U5959 , P1_REG1_REG_28_ , P1_U3948 );
nand NAND2_3264 ( P1_U5960 , P1_U4023 , P1_U4725 );
nand NAND2_3265 ( P1_U5961 , P1_REG1_REG_29_ , P1_U3948 );
nand NAND2_3266 ( P1_U5962 , P1_U4023 , P1_U4745 );
nand NAND2_3267 ( P1_U5963 , P1_REG1_REG_30_ , P1_U3948 );
nand NAND2_3268 ( P1_U5964 , P1_U4023 , P1_U4752 );
nand NAND2_3269 ( P1_U5965 , P1_REG1_REG_31_ , P1_U3948 );
nand NAND2_3270 ( P1_U5966 , P1_U4023 , P1_U4755 );
nand NAND2_3271 ( P1_U5967 , P1_REG2_REG_0_ , P1_U3417 );
nand NAND2_3272 ( P1_U5968 , P1_U4022 , P1_U3373 );
nand NAND2_3273 ( P1_U5969 , P1_REG2_REG_1_ , P1_U3417 );
nand NAND2_3274 ( P1_U5970 , P1_U4022 , P1_U3375 );
nand NAND2_3275 ( P1_U5971 , P1_REG2_REG_2_ , P1_U3417 );
nand NAND2_3276 ( P1_U5972 , P1_U4022 , P1_U3376 );
nand NAND2_3277 ( P1_U5973 , P1_REG2_REG_3_ , P1_U3417 );
nand NAND2_3278 ( P1_U5974 , P1_U4022 , P1_U3377 );
nand NAND2_3279 ( P1_U5975 , P1_REG2_REG_4_ , P1_U3417 );
nand NAND2_3280 ( P1_U5976 , P1_U4022 , P1_U3378 );
nand NAND2_3281 ( P1_U5977 , P1_REG2_REG_5_ , P1_U3417 );
nand NAND2_3282 ( P1_U5978 , P1_U4022 , P1_U3379 );
nand NAND2_3283 ( P1_U5979 , P1_REG2_REG_6_ , P1_U3417 );
nand NAND2_3284 ( P1_U5980 , P1_U4022 , P1_U3380 );
nand NAND2_3285 ( P1_U5981 , P1_REG2_REG_7_ , P1_U3417 );
nand NAND2_3286 ( P1_U5982 , P1_U4022 , P1_U3381 );
nand NAND2_3287 ( P1_U5983 , P1_REG2_REG_8_ , P1_U3417 );
nand NAND2_3288 ( P1_U5984 , P1_U4022 , P1_U3382 );
nand NAND2_3289 ( P1_U5985 , P1_REG2_REG_9_ , P1_U3417 );
nand NAND2_3290 ( P1_U5986 , P1_U4022 , P1_U3383 );
nand NAND2_3291 ( P1_U5987 , P1_REG2_REG_10_ , P1_U3417 );
nand NAND2_3292 ( P1_U5988 , P1_U4022 , P1_U3384 );
nand NAND2_3293 ( P1_U5989 , P1_REG2_REG_11_ , P1_U3417 );
nand NAND2_3294 ( P1_U5990 , P1_U4022 , P1_U3385 );
nand NAND2_3295 ( P1_U5991 , P1_REG2_REG_12_ , P1_U3417 );
nand NAND2_3296 ( P1_U5992 , P1_U4022 , P1_U3386 );
nand NAND2_3297 ( P1_U5993 , P1_REG2_REG_13_ , P1_U3417 );
nand NAND2_3298 ( P1_U5994 , P1_U4022 , P1_U3387 );
nand NAND2_3299 ( P1_U5995 , P1_REG2_REG_14_ , P1_U3417 );
nand NAND2_3300 ( P1_U5996 , P1_U4022 , P1_U3388 );
nand NAND2_3301 ( P1_U5997 , P1_REG2_REG_15_ , P1_U3417 );
nand NAND2_3302 ( P1_U5998 , P1_U4022 , P1_U3389 );
nand NAND2_3303 ( P1_U5999 , P1_REG2_REG_16_ , P1_U3417 );
nand NAND2_3304 ( P1_U6000 , P1_U4022 , P1_U3390 );
nand NAND2_3305 ( P1_U6001 , P1_REG2_REG_17_ , P1_U3417 );
nand NAND2_3306 ( P1_U6002 , P1_U4022 , P1_U3391 );
nand NAND2_3307 ( P1_U6003 , P1_REG2_REG_18_ , P1_U3417 );
nand NAND2_3308 ( P1_U6004 , P1_U4022 , P1_U3392 );
nand NAND2_3309 ( P1_U6005 , P1_REG2_REG_19_ , P1_U3417 );
nand NAND2_3310 ( P1_U6006 , P1_U4022 , P1_U3393 );
nand NAND2_3311 ( P1_U6007 , P1_REG2_REG_20_ , P1_U3417 );
nand NAND2_3312 ( P1_U6008 , P1_U4022 , P1_U3395 );
nand NAND2_3313 ( P1_U6009 , P1_REG2_REG_21_ , P1_U3417 );
nand NAND2_3314 ( P1_U6010 , P1_U4022 , P1_U3397 );
nand NAND2_3315 ( P1_U6011 , P1_REG2_REG_22_ , P1_U3417 );
nand NAND2_3316 ( P1_U6012 , P1_U4022 , P1_U3399 );
nand NAND2_3317 ( P1_U6013 , P1_REG2_REG_23_ , P1_U3417 );
nand NAND2_3318 ( P1_U6014 , P1_U4022 , P1_U3401 );
nand NAND2_3319 ( P1_U6015 , P1_REG2_REG_24_ , P1_U3417 );
nand NAND2_3320 ( P1_U6016 , P1_U4022 , P1_U3403 );
nand NAND2_3321 ( P1_U6017 , P1_REG2_REG_25_ , P1_U3417 );
nand NAND2_3322 ( P1_U6018 , P1_U4022 , P1_U3405 );
nand NAND2_3323 ( P1_U6019 , P1_REG2_REG_26_ , P1_U3417 );
nand NAND2_3324 ( P1_U6020 , P1_U4022 , P1_U3407 );
nand NAND2_3325 ( P1_U6021 , P1_REG2_REG_27_ , P1_U3417 );
nand NAND2_3326 ( P1_U6022 , P1_U4022 , P1_U3409 );
nand NAND2_3327 ( P1_U6023 , P1_REG2_REG_28_ , P1_U3417 );
nand NAND2_3328 ( P1_U6024 , P1_U4022 , P1_U3411 );
nand NAND2_3329 ( P1_U6025 , P1_REG2_REG_29_ , P1_U3417 );
nand NAND2_3330 ( P1_U6026 , P1_U4022 , P1_U3413 );
nand NAND2_3331 ( P1_U6027 , P1_REG2_REG_30_ , P1_U3417 );
nand NAND2_3332 ( P1_U6028 , P1_U4026 , P1_U4022 );
nand NAND2_3333 ( P1_U6029 , P1_REG2_REG_31_ , P1_U3417 );
nand NAND2_3334 ( P1_U6030 , P1_U4026 , P1_U4022 );
nand NAND2_3335 ( P1_U6031 , P1_DATAO_REG_0_ , P1_U3425 );
nand NAND2_3336 ( P1_U6032 , P1_U4006 , P1_U3075 );
nand NAND2_3337 ( P1_U6033 , P1_DATAO_REG_1_ , P1_U3425 );
nand NAND2_3338 ( P1_U6034 , P1_U4006 , P1_U3076 );
nand NAND2_3339 ( P1_U6035 , P1_DATAO_REG_2_ , P1_U3425 );
nand NAND2_3340 ( P1_U6036 , P1_U4006 , P1_U3066 );
nand NAND2_3341 ( P1_U6037 , P1_DATAO_REG_3_ , P1_U3425 );
nand NAND2_3342 ( P1_U6038 , P1_U4006 , P1_U3062 );
nand NAND2_3343 ( P1_U6039 , P1_DATAO_REG_4_ , P1_U3425 );
nand NAND2_3344 ( P1_U6040 , P1_U4006 , P1_U3058 );
nand NAND2_3345 ( P1_U6041 , P1_DATAO_REG_5_ , P1_U3425 );
nand NAND2_3346 ( P1_U6042 , P1_U4006 , P1_U3065 );
nand NAND2_3347 ( P1_U6043 , P1_DATAO_REG_6_ , P1_U3425 );
nand NAND2_3348 ( P1_U6044 , P1_U4006 , P1_U3069 );
nand NAND2_3349 ( P1_U6045 , P1_DATAO_REG_7_ , P1_U3425 );
nand NAND2_3350 ( P1_U6046 , P1_U4006 , P1_U3068 );
nand NAND2_3351 ( P1_U6047 , P1_DATAO_REG_8_ , P1_U3425 );
nand NAND2_3352 ( P1_U6048 , P1_U4006 , P1_U3082 );
nand NAND2_3353 ( P1_U6049 , P1_DATAO_REG_9_ , P1_U3425 );
nand NAND2_3354 ( P1_U6050 , P1_U4006 , P1_U3081 );
nand NAND2_3355 ( P1_U6051 , P1_DATAO_REG_10_ , P1_U3425 );
nand NAND2_3356 ( P1_U6052 , P1_U4006 , P1_U3060 );
nand NAND2_3357 ( P1_U6053 , P1_DATAO_REG_11_ , P1_U3425 );
nand NAND2_3358 ( P1_U6054 , P1_U4006 , P1_U3061 );
nand NAND2_3359 ( P1_U6055 , P1_DATAO_REG_12_ , P1_U3425 );
nand NAND2_3360 ( P1_U6056 , P1_U4006 , P1_U3070 );
nand NAND2_3361 ( P1_U6057 , P1_DATAO_REG_13_ , P1_U3425 );
nand NAND2_3362 ( P1_U6058 , P1_U4006 , P1_U3078 );
nand NAND2_3363 ( P1_U6059 , P1_DATAO_REG_14_ , P1_U3425 );
nand NAND2_3364 ( P1_U6060 , P1_U4006 , P1_U3077 );
nand NAND2_3365 ( P1_U6061 , P1_DATAO_REG_15_ , P1_U3425 );
nand NAND2_3366 ( P1_U6062 , P1_U4006 , P1_U3072 );
nand NAND2_3367 ( P1_U6063 , P1_DATAO_REG_16_ , P1_U3425 );
nand NAND2_3368 ( P1_U6064 , P1_U4006 , P1_U3071 );
nand NAND2_3369 ( P1_U6065 , P1_DATAO_REG_17_ , P1_U3425 );
nand NAND2_3370 ( P1_U6066 , P1_U4006 , P1_U3067 );
nand NAND2_3371 ( P1_U6067 , P1_DATAO_REG_18_ , P1_U3425 );
nand NAND2_3372 ( P1_U6068 , P1_U4006 , P1_U3080 );
nand NAND2_3373 ( P1_U6069 , P1_DATAO_REG_19_ , P1_U3425 );
nand NAND2_3374 ( P1_U6070 , P1_U4006 , P1_U3079 );
nand NAND2_3375 ( P1_U6071 , P1_DATAO_REG_20_ , P1_U3425 );
nand NAND2_3376 ( P1_U6072 , P1_U4006 , P1_U3074 );
nand NAND2_3377 ( P1_U6073 , P1_DATAO_REG_21_ , P1_U3425 );
nand NAND2_3378 ( P1_U6074 , P1_U4006 , P1_U3073 );
nand NAND2_3379 ( P1_U6075 , P1_DATAO_REG_22_ , P1_U3425 );
nand NAND2_3380 ( P1_U6076 , P1_U4006 , P1_U3059 );
nand NAND2_3381 ( P1_U6077 , P1_DATAO_REG_23_ , P1_U3425 );
nand NAND2_3382 ( P1_U6078 , P1_U4006 , P1_U3064 );
nand NAND2_3383 ( P1_U6079 , P1_DATAO_REG_24_ , P1_U3425 );
nand NAND2_3384 ( P1_U6080 , P1_U4006 , P1_U3063 );
nand NAND2_3385 ( P1_U6081 , P1_DATAO_REG_25_ , P1_U3425 );
nand NAND2_3386 ( P1_U6082 , P1_U4006 , P1_U3056 );
nand NAND2_3387 ( P1_U6083 , P1_DATAO_REG_26_ , P1_U3425 );
nand NAND2_3388 ( P1_U6084 , P1_U4006 , P1_U3055 );
nand NAND2_3389 ( P1_U6085 , P1_DATAO_REG_27_ , P1_U3425 );
nand NAND2_3390 ( P1_U6086 , P1_U4006 , P1_U3051 );
nand NAND2_3391 ( P1_U6087 , P1_DATAO_REG_28_ , P1_U3425 );
nand NAND2_3392 ( P1_U6088 , P1_U4006 , P1_U3052 );
nand NAND2_3393 ( P1_U6089 , P1_DATAO_REG_29_ , P1_U3425 );
nand NAND2_3394 ( P1_U6090 , P1_U4006 , P1_U3053 );
nand NAND2_3395 ( P1_U6091 , P1_DATAO_REG_30_ , P1_U3425 );
nand NAND2_3396 ( P1_U6092 , P1_U4006 , P1_U3057 );
nand NAND2_3397 ( P1_U6093 , P1_DATAO_REG_31_ , P1_U3425 );
nand NAND2_3398 ( P1_U6094 , P1_U4006 , P1_U3054 );
nand NAND2_3399 ( P1_U6095 , P1_U4007 , P1_U3052 );
nand NAND2_3400 ( P1_U6096 , P1_U3410 , P1_U4692 );
nand NAND2_3401 ( P1_U6097 , P1_U6096 , P1_U6095 );
nand NAND2_3402 ( P1_U6098 , P1_U4008 , P1_U3051 );
nand NAND2_3403 ( P1_U6099 , P1_U3408 , P1_U4673 );
nand NAND2_3404 ( P1_U6100 , P1_U6099 , P1_U6098 );
nand NAND2_3405 ( P1_U6101 , P1_U4011 , P1_U3063 );
nand NAND2_3406 ( P1_U6102 , P1_U3402 , P1_U4616 );
nand NAND2_3407 ( P1_U6103 , P1_U6102 , P1_U6101 );
nand NAND2_3408 ( P1_U6104 , P1_U4012 , P1_U3064 );
nand NAND2_3409 ( P1_U6105 , P1_U3400 , P1_U4597 );
nand NAND2_3410 ( P1_U6106 , P1_U6105 , P1_U6104 );
nand NAND2_3411 ( P1_U6107 , P1_U4014 , P1_U3073 );
nand NAND2_3412 ( P1_U6108 , P1_U3396 , P1_U4559 );
nand NAND2_3413 ( P1_U6109 , P1_U6108 , P1_U6107 );
nand NAND2_3414 ( P1_U6110 , P1_U4013 , P1_U3059 );
nand NAND2_3415 ( P1_U6111 , P1_U3398 , P1_U4578 );
nand NAND2_3416 ( P1_U6112 , P1_U6111 , P1_U6110 );
nand NAND2_3417 ( P1_U6113 , P1_U4010 , P1_U3056 );
nand NAND2_3418 ( P1_U6114 , P1_U3404 , P1_U4635 );
nand NAND2_3419 ( P1_U6115 , P1_U6114 , P1_U6113 );
nand NAND2_3420 ( P1_U6116 , P1_U4009 , P1_U3055 );
nand NAND2_3421 ( P1_U6117 , P1_U3406 , P1_U4654 );
nand NAND2_3422 ( P1_U6118 , P1_U6117 , P1_U6116 );
nand NAND2_3423 ( P1_U6119 , P1_U5864 , P1_U4483 );
nand NAND2_3424 ( P1_U6120 , P1_U3504 , P1_U3067 );
nand NAND2_3425 ( P1_U6121 , P1_U6120 , P1_U6119 );
nand NAND2_3426 ( P1_U6122 , P1_U5801 , P1_U4312 );
nand NAND2_3427 ( P1_U6123 , P1_U3477 , P1_U3082 );
nand NAND2_3428 ( P1_U6124 , P1_U6123 , P1_U6122 );
nand NAND2_3429 ( P1_U6125 , P1_U5808 , P1_U4331 );
nand NAND2_3430 ( P1_U6126 , P1_U3480 , P1_U3081 );
nand NAND2_3431 ( P1_U6127 , P1_U6126 , P1_U6125 );
nand NAND2_3432 ( P1_U6128 , P1_U5836 , P1_U4407 );
nand NAND2_3433 ( P1_U6129 , P1_U3492 , P1_U3078 );
nand NAND2_3434 ( P1_U6130 , P1_U6129 , P1_U6128 );
nand NAND2_3435 ( P1_U6131 , P1_U5843 , P1_U4426 );
nand NAND2_3436 ( P1_U6132 , P1_U3495 , P1_U3077 );
nand NAND2_3437 ( P1_U6133 , P1_U6132 , P1_U6131 );
nand NAND2_3438 ( P1_U6134 , P1_U5737 , P1_U4198 );
nand NAND2_3439 ( P1_U6135 , P1_U3451 , P1_U3075 );
nand NAND2_3440 ( P1_U6136 , P1_U6135 , P1_U6134 );
nand NAND2_3441 ( P1_U6137 , P1_U5752 , P1_U4174 );
nand NAND2_3442 ( P1_U6138 , P1_U3456 , P1_U3076 );
nand NAND2_3443 ( P1_U6139 , P1_U6138 , P1_U6137 );
nand NAND2_3444 ( P1_U6140 , P1_U5850 , P1_U4445 );
nand NAND2_3445 ( P1_U6141 , P1_U3498 , P1_U3072 );
nand NAND2_3446 ( P1_U6142 , P1_U6141 , P1_U6140 );
nand NAND2_3447 ( P1_U6143 , P1_U5857 , P1_U4464 );
nand NAND2_3448 ( P1_U6144 , P1_U3501 , P1_U3071 );
nand NAND2_3449 ( P1_U6145 , P1_U6144 , P1_U6143 );
nand NAND2_3450 ( P1_U6146 , P1_U5787 , P1_U4274 );
nand NAND2_3451 ( P1_U6147 , P1_U3471 , P1_U3069 );
nand NAND2_3452 ( P1_U6148 , P1_U6147 , P1_U6146 );
nand NAND2_3453 ( P1_U6149 , P1_U5794 , P1_U4293 );
nand NAND2_3454 ( P1_U6150 , P1_U3474 , P1_U3068 );
nand NAND2_3455 ( P1_U6151 , P1_U6150 , P1_U6149 );
nand NAND2_3456 ( P1_U6152 , P1_U5829 , P1_U4388 );
nand NAND2_3457 ( P1_U6153 , P1_U3489 , P1_U3070 );
nand NAND2_3458 ( P1_U6154 , P1_U6153 , P1_U6152 );
nand NAND2_3459 ( P1_U6155 , P1_U5759 , P1_U4193 );
nand NAND2_3460 ( P1_U6156 , P1_U3459 , P1_U3066 );
nand NAND2_3461 ( P1_U6157 , P1_U6156 , P1_U6155 );
nand NAND2_3462 ( P1_U6158 , P1_U5766 , P1_U4217 );
nand NAND2_3463 ( P1_U6159 , P1_U3462 , P1_U3062 );
nand NAND2_3464 ( P1_U6160 , P1_U6159 , P1_U6158 );
nand NAND2_3465 ( P1_U6161 , P1_U5780 , P1_U4255 );
nand NAND2_3466 ( P1_U6162 , P1_U3468 , P1_U3065 );
nand NAND2_3467 ( P1_U6163 , P1_U6162 , P1_U6161 );
nand NAND2_3468 ( P1_U6164 , P1_U5871 , P1_U4502 );
nand NAND2_3469 ( P1_U6165 , P1_U3507 , P1_U3080 );
nand NAND2_3470 ( P1_U6166 , P1_U6165 , P1_U6164 );
nand NAND2_3471 ( P1_U6167 , P1_U4016 , P1_U3054 );
nand NAND2_3472 ( P1_U6168 , P1_U3415 , P1_U4749 );
nand NAND2_3473 ( P1_U6169 , P1_U6168 , P1_U6167 );
nand NAND2_3474 ( P1_U6170 , P1_U5876 , P1_U4521 );
nand NAND2_3475 ( P1_U6171 , P1_U3509 , P1_U3079 );
nand NAND2_3476 ( P1_U6172 , P1_U6171 , P1_U6170 );
nand NAND2_3477 ( P1_U6173 , P1_U5822 , P1_U4369 );
nand NAND2_3478 ( P1_U6174 , P1_U3486 , P1_U3061 );
nand NAND2_3479 ( P1_U6175 , P1_U6174 , P1_U6173 );
nand NAND2_3480 ( P1_U6176 , P1_U5773 , P1_U4236 );
nand NAND2_3481 ( P1_U6177 , P1_U3465 , P1_U3058 );
nand NAND2_3482 ( P1_U6178 , P1_U6177 , P1_U6176 );
nand NAND2_3483 ( P1_U6179 , P1_U5815 , P1_U4350 );
nand NAND2_3484 ( P1_U6180 , P1_U3483 , P1_U3060 );
nand NAND2_3485 ( P1_U6181 , P1_U6180 , P1_U6179 );
nand NAND2_3486 ( P1_U6182 , P1_U4015 , P1_U3074 );
nand NAND2_3487 ( P1_U6183 , P1_U3394 , P1_U4540 );
nand NAND2_3488 ( P1_U6184 , P1_U6183 , P1_U6182 );
nand NAND2_3489 ( P1_U6185 , P1_U4018 , P1_U3053 );
nand NAND2_3490 ( P1_U6186 , P1_U3412 , P1_U4711 );
nand NAND2_3491 ( P1_U6187 , P1_U6186 , P1_U6185 );
nand NAND2_3492 ( P1_U6188 , P1_U4017 , P1_U3057 );
nand NAND2_3493 ( P1_U6189 , P1_U3414 , P1_U4729 );
nand NAND2_3494 ( P1_U6190 , P1_U6189 , P1_U6188 );
nand NAND2_3495 ( P1_U6191 , P1_U5119 , P1_U3987 );
nand NAND2_3496 ( P1_U6192 , P1_U3354 , P1_U3982 );
nand NAND2_3497 ( P1_U6193 , P1_U6192 , P1_U6191 );
nand NAND4_3498 ( P1_U6194 , P1_U3439 , P1_U5710 , P1_U3983 , P1_U3448 );
nand NAND2_3499 ( P1_U6195 , P1_U6193 , P1_U5719 );
nand NAND2_3500 ( P1_U6196 , P1_U6195 , P1_U6194 );
nand NAND3_3501 ( P1_U6197 , P1_R1375_U14 , P1_U3987 , P1_U5716 );
nand NAND2_3502 ( P1_U6198 , P1_U6196 , P1_U3442 );
nand NAND3_3503 ( P1_U6199 , P1_U4019 , P1_U3022 , P1_U3983 );
nand NAND3_3504 ( P1_U6200 , P1_U3988 , P1_U3992 , P1_R1360_U14 );
nand NAND2_3505 ( P1_U6201 , P1_U3081 , P1_R1352_U6 );
nand NAND2_3506 ( P1_U6202 , P1_U3081 , P1_U3985 );
nand NAND2_3507 ( P1_U6203 , P1_U3082 , P1_R1352_U6 );
nand NAND2_3508 ( P1_U6204 , P1_U3082 , P1_U3985 );
nand NAND2_3509 ( P1_U6205 , P1_U3068 , P1_R1352_U6 );
nand NAND2_3510 ( P1_U6206 , P1_U3068 , P1_U3985 );
nand NAND2_3511 ( P1_U6207 , P1_U3069 , P1_R1352_U6 );
nand NAND2_3512 ( P1_U6208 , P1_U3069 , P1_U3985 );
nand NAND2_3513 ( P1_U6209 , P1_U3065 , P1_R1352_U6 );
nand NAND2_3514 ( P1_U6210 , P1_U3065 , P1_U3985 );
nand NAND2_3515 ( P1_U6211 , P1_U3058 , P1_R1352_U6 );
nand NAND2_3516 ( P1_U6212 , P1_U3058 , P1_U3985 );
nand NAND2_3517 ( P1_U6213 , P1_U3062 , P1_R1352_U6 );
nand NAND2_3518 ( P1_U6214 , P1_U3062 , P1_U3985 );
nand NAND2_3519 ( P1_U6215 , P1_R1309_U8 , P1_R1352_U6 );
nand NAND2_3520 ( P1_U6216 , P1_U3054 , P1_U3985 );
nand NAND2_3521 ( P1_U6217 , P1_R1309_U6 , P1_R1352_U6 );
nand NAND2_3522 ( P1_U6218 , P1_U3057 , P1_U3985 );
nand NAND2_3523 ( P1_U6219 , P1_U3066 , P1_R1352_U6 );
nand NAND2_3524 ( P1_U6220 , P1_U3066 , P1_U3985 );
nand NAND2_3525 ( P1_U6221 , P1_U3053 , P1_R1352_U6 );
nand NAND2_3526 ( P1_U6222 , P1_U3053 , P1_U3985 );
nand NAND2_3527 ( P1_U6223 , P1_U3052 , P1_R1352_U6 );
nand NAND2_3528 ( P1_U6224 , P1_U3052 , P1_U3985 );
nand NAND2_3529 ( P1_U6225 , P1_U3051 , P1_R1352_U6 );
nand NAND2_3530 ( P1_U6226 , P1_U3051 , P1_U3985 );
nand NAND2_3531 ( P1_U6227 , P1_U3055 , P1_R1352_U6 );
nand NAND2_3532 ( P1_U6228 , P1_U3055 , P1_U3985 );
nand NAND2_3533 ( P1_U6229 , P1_U3056 , P1_R1352_U6 );
nand NAND2_3534 ( P1_U6230 , P1_U3056 , P1_U3985 );
nand NAND2_3535 ( P1_U6231 , P1_U3063 , P1_R1352_U6 );
nand NAND2_3536 ( P1_U6232 , P1_U3063 , P1_U3985 );
nand NAND2_3537 ( P1_U6233 , P1_U3064 , P1_R1352_U6 );
nand NAND2_3538 ( P1_U6234 , P1_U3064 , P1_U3985 );
nand NAND2_3539 ( P1_U6235 , P1_U3059 , P1_R1352_U6 );
nand NAND2_3540 ( P1_U6236 , P1_U3059 , P1_U3985 );
nand NAND2_3541 ( P1_U6237 , P1_U3073 , P1_R1352_U6 );
nand NAND2_3542 ( P1_U6238 , P1_U3073 , P1_U3985 );
nand NAND2_3543 ( P1_U6239 , P1_U3074 , P1_R1352_U6 );
nand NAND2_3544 ( P1_U6240 , P1_U3074 , P1_U3985 );
nand NAND2_3545 ( P1_U6241 , P1_U3076 , P1_R1352_U6 );
nand NAND2_3546 ( P1_U6242 , P1_U3076 , P1_U3985 );
nand NAND2_3547 ( P1_U6243 , P1_U3079 , P1_R1352_U6 );
nand NAND2_3548 ( P1_U6244 , P1_U3079 , P1_U3985 );
nand NAND2_3549 ( P1_U6245 , P1_U3080 , P1_R1352_U6 );
nand NAND2_3550 ( P1_U6246 , P1_U3080 , P1_U3985 );
nand NAND2_3551 ( P1_U6247 , P1_U3067 , P1_R1352_U6 );
nand NAND2_3552 ( P1_U6248 , P1_U3067 , P1_U3985 );
nand NAND2_3553 ( P1_U6249 , P1_U3071 , P1_R1352_U6 );
nand NAND2_3554 ( P1_U6250 , P1_U3071 , P1_U3985 );
nand NAND2_3555 ( P1_U6251 , P1_U3072 , P1_R1352_U6 );
nand NAND2_3556 ( P1_U6252 , P1_U3072 , P1_U3985 );
nand NAND2_3557 ( P1_U6253 , P1_U3077 , P1_R1352_U6 );
nand NAND2_3558 ( P1_U6254 , P1_U3077 , P1_U3985 );
nand NAND2_3559 ( P1_U6255 , P1_U3078 , P1_R1352_U6 );
nand NAND2_3560 ( P1_U6256 , P1_U3078 , P1_U3985 );
nand NAND2_3561 ( P1_U6257 , P1_U3070 , P1_R1352_U6 );
nand NAND2_3562 ( P1_U6258 , P1_U3070 , P1_U3985 );
nand NAND2_3563 ( P1_U6259 , P1_U3061 , P1_R1352_U6 );
nand NAND2_3564 ( P1_U6260 , P1_U3061 , P1_U3985 );
nand NAND2_3565 ( P1_U6261 , P1_U3060 , P1_R1352_U6 );
nand NAND2_3566 ( P1_U6262 , P1_U3060 , P1_U3985 );
nand NAND2_3567 ( P1_U6263 , P1_U3075 , P1_R1352_U6 );
nand NAND2_3568 ( P1_U6264 , P1_U3075 , P1_U3985 );
nand NAND2_3569 ( P1_U6265 , P1_U3449 , P1_U5396 );
nand NAND3_3570 ( P1_U6266 , P1_U3015 , P1_REG2_REG_0_ , P1_U5731 );
nand NAND2_3571 ( P2_R1113_U462 , P2_U3080 , P2_R1113_U54 );
nand NAND2_3572 ( P2_R1113_U461 , P2_U3489 , P2_R1113_U55 );
nand NAND2_3573 ( P2_R1113_U460 , P2_R1113_U258 , P2_R1113_U172 );
nand NAND2_3574 ( P2_R1113_U459 , P2_R1113_U335 , P2_R1113_U173 );
nand NAND2_3575 ( P2_R1113_U458 , P2_U3079 , P2_R1113_U57 );
nand NAND2_3576 ( P2_R1113_U457 , P2_U3492 , P2_R1113_U60 );
nand NAND2_3577 ( P2_R1113_U456 , P2_R1113_U171 , P2_R1113_U326 );
nand NAND2_3578 ( P2_R1113_U455 , P2_R1113_U334 , P2_R1113_U87 );
nand NAND2_3579 ( P2_R1113_U454 , P2_U3074 , P2_R1113_U46 );
nand NAND2_3580 ( P2_R1113_U453 , P2_U3495 , P2_R1113_U59 );
nand NAND2_3581 ( P2_R1113_U452 , P2_R1113_U451 , P2_R1113_U450 );
nand NAND2_3582 ( P2_R1113_U451 , P2_U3073 , P2_R1113_U56 );
nand NAND2_3583 ( P2_R1113_U450 , P2_U3498 , P2_R1113_U58 );
nand NAND2_3584 ( P2_R1113_U449 , P2_R1113_U140 , P2_R1113_U170 );
nand NAND2_3585 ( P2_R1113_U448 , P2_R1113_U268 , P2_R1113_U447 );
not NOT1_3586 ( P2_R1113_U447 , P2_R1113_U140 );
nand NAND2_3587 ( P2_R1113_U446 , P2_U3069 , P2_R1113_U62 );
nand NAND2_3588 ( P2_R1113_U445 , P2_U3501 , P2_R1113_U63 );
nand NAND2_3589 ( P2_R1113_U444 , P2_R1113_U139 , P2_R1113_U169 );
nand NAND2_3590 ( P2_R1113_U443 , P2_R1113_U272 , P2_R1113_U442 );
not NOT1_3591 ( P2_R1113_U442 , P2_R1113_U139 );
nand NAND2_3592 ( P2_R1113_U441 , P2_U3082 , P2_R1113_U168 );
nand NAND2_3593 ( P2_R1113_U440 , P2_U3504 , P2_R1113_U64 );
nand NAND2_3594 ( P2_R1113_U439 , P2_R1113_U138 , P2_R1113_U167 );
and AND3_3595 ( P2_U3014 , P2_U5711 , P2_U3441 , P2_U3439 );
and AND3_3596 ( P2_U3015 , P2_U3439 , P2_U3441 , P2_U3445 );
and AND2_3597 ( P2_U3016 , P2_U3954 , P2_U5714 );
and AND2_3598 ( P2_U3017 , P2_U3961 , P2_U3440 );
and AND3_3599 ( P2_U3018 , P2_U3439 , P2_U3445 , P2_U3440 );
and AND2_3600 ( P2_U3019 , P2_U5674 , P2_U3439 );
and AND2_3601 ( P2_U3020 , P2_U3629 , P2_U3624 );
and AND2_3602 ( P2_U3021 , P2_U5733 , P2_U3444 );
and AND2_3603 ( P2_U3022 , P2_U3447 , P2_U3444 );
and AND2_3604 ( P2_U3023 , P2_U3442 , P2_U3443 );
and AND2_3605 ( P2_U3024 , P2_U5723 , P2_U3443 );
and AND2_3606 ( P2_U3025 , P2_U5720 , P2_U3442 );
and AND2_3607 ( P2_U3026 , P2_U5723 , P2_U5720 );
and AND2_3608 ( P2_U3027 , P2_U3048 , P2_STATE_REG );
and AND2_3609 ( P2_U3028 , P2_U3050 , P2_U5708 );
and AND2_3610 ( P2_U3029 , P2_U3811 , P2_U3424 );
and AND2_3611 ( P2_U3030 , P2_U3982 , P2_U5728 );
and AND2_3612 ( P2_U3031 , P2_U3949 , P2_U5714 );
and AND2_3613 ( P2_U3032 , P2_U3890 , P2_U3965 );
and AND2_3614 ( P2_U3033 , P2_U3359 , P2_STATE_REG );
and AND2_3615 ( P2_U3034 , P2_U3956 , P2_U3983 );
and AND2_3616 ( P2_U3035 , P2_U3983 , P2_U4713 );
and AND2_3617 ( P2_U3036 , P2_U3957 , P2_U3983 );
and AND2_3618 ( P2_U3037 , P2_U3751 , P2_U3983 );
and AND2_3619 ( P2_U3038 , P2_U3982 , P2_U3444 );
and AND2_3620 ( P2_U3039 , P2_U3965 , P2_U5728 );
and AND2_3621 ( P2_U3040 , P2_U3983 , P2_U3030 );
and AND2_3622 ( P2_U3041 , P2_U3965 , P2_U3444 );
and AND2_3623 ( P2_U3042 , P2_U3029 , P2_U5733 );
and AND2_3624 ( P2_U3043 , P2_U3029 , P2_U5728 );
and AND2_3625 ( P2_U3044 , P2_U3029 , P2_U3022 );
and AND2_3626 ( P2_U3045 , P2_U3027 , P2_U3424 );
and AND2_3627 ( P2_U3046 , P2_U5196 , P2_STATE_REG );
and AND2_3628 ( P2_U3047 , P2_U3027 , P2_U5198 );
and AND2_3629 ( P2_U3048 , P2_U5701 , P2_U3420 );
and AND2_3630 ( P2_U3049 , P2_U3630 , P2_U3020 );
and AND2_3631 ( P2_U3050 , P2_U5714 , P2_U3445 );
and AND2_3632 ( P2_U3051 , P2_U3950 , P2_U4709 );
and AND2_3633 ( P2_U3052 , P2_U3422 , P2_STATE_REG );
nand NAND4_3634 ( P2_U3053 , P2_U4623 , P2_U4624 , P2_U4622 , P2_U4625 );
nand NAND4_3635 ( P2_U3054 , P2_U4642 , P2_U4643 , P2_U4641 , P2_U4644 );
nand NAND4_3636 ( P2_U3055 , P2_U4663 , P2_U4662 , P2_U4661 , P2_U4660 );
nand NAND3_3637 ( P2_U3056 , P2_U4700 , P2_U4701 , P2_U4699 );
nand NAND4_3638 ( P2_U3057 , P2_U4604 , P2_U4605 , P2_U4603 , P2_U4606 );
nand NAND4_3639 ( P2_U3058 , P2_U4585 , P2_U4586 , P2_U4584 , P2_U4587 );
nand NAND3_3640 ( P2_U3059 , P2_U4680 , P2_U4681 , P2_U4679 );
nand NAND4_3641 ( P2_U3060 , P2_U4188 , P2_U4187 , P2_U4186 , P2_U4185 );
nand NAND4_3642 ( P2_U3061 , P2_U4528 , P2_U4529 , P2_U4527 , P2_U4530 );
nand NAND4_3643 ( P2_U3062 , P2_U4302 , P2_U4301 , P2_U4300 , P2_U4299 );
nand NAND4_3644 ( P2_U3063 , P2_U4321 , P2_U4320 , P2_U4319 , P2_U4318 );
nand NAND4_3645 ( P2_U3064 , P2_U4169 , P2_U4168 , P2_U4167 , P2_U4166 );
nand NAND4_3646 ( P2_U3065 , P2_U4566 , P2_U4567 , P2_U4565 , P2_U4568 );
nand NAND4_3647 ( P2_U3066 , P2_U4547 , P2_U4548 , P2_U4546 , P2_U4549 );
nand NAND4_3648 ( P2_U3067 , P2_U4207 , P2_U4206 , P2_U4205 , P2_U4204 );
nand NAND4_3649 ( P2_U3068 , P2_U4147 , P2_U4146 , P2_U5755 , P2_U5754 );
nand NAND4_3650 ( P2_U3069 , P2_U4433 , P2_U4434 , P2_U4432 , P2_U4435 );
nand NAND4_3651 ( P2_U3070 , P2_U4245 , P2_U4244 , P2_U4243 , P2_U4242 );
nand NAND4_3652 ( P2_U3071 , P2_U4226 , P2_U4225 , P2_U4224 , P2_U4223 );
nand NAND4_3653 ( P2_U3072 , P2_U4340 , P2_U4339 , P2_U4338 , P2_U4337 );
nand NAND4_3654 ( P2_U3073 , P2_U4416 , P2_U4415 , P2_U4414 , P2_U4413 );
nand NAND4_3655 ( P2_U3074 , P2_U4397 , P2_U4396 , P2_U4395 , P2_U4394 );
nand NAND4_3656 ( P2_U3075 , P2_U4509 , P2_U4510 , P2_U4508 , P2_U4511 );
nand NAND4_3657 ( P2_U3076 , P2_U4490 , P2_U4491 , P2_U4489 , P2_U4492 );
nand NAND4_3658 ( P2_U3077 , P2_U4150 , P2_U4149 , P2_U5748 , P2_U5747 );
nand NAND4_3659 ( P2_U3078 , P2_U4129 , P2_U4128 , P2_U5725 , P2_U5724 );
nand NAND4_3660 ( P2_U3079 , P2_U4378 , P2_U4377 , P2_U4376 , P2_U4375 );
nand NAND4_3661 ( P2_U3080 , P2_U4359 , P2_U4358 , P2_U4357 , P2_U4356 );
nand NAND4_3662 ( P2_U3081 , P2_U4471 , P2_U4472 , P2_U4470 , P2_U4473 );
nand NAND4_3663 ( P2_U3082 , P2_U4452 , P2_U4453 , P2_U4451 , P2_U4454 );
nand NAND4_3664 ( P2_U3083 , P2_U4283 , P2_U4282 , P2_U4281 , P2_U4280 );
nand NAND4_3665 ( P2_U3084 , P2_U4264 , P2_U4263 , P2_U4262 , P2_U4261 );
nand NAND2_3666 ( P2_U3085 , P2_U5596 , P2_U5595 );
nand NAND2_3667 ( P2_U3086 , P2_U5598 , P2_U5597 );
nand NAND3_3668 ( P2_U3087 , P2_U5603 , P2_U5604 , P2_U5602 );
nand NAND3_3669 ( P2_U3088 , P2_U5606 , P2_U5607 , P2_U5605 );
nand NAND3_3670 ( P2_U3089 , P2_U5609 , P2_U5610 , P2_U5608 );
nand NAND3_3671 ( P2_U3090 , P2_U5612 , P2_U5613 , P2_U5611 );
nand NAND3_3672 ( P2_U3091 , P2_U5615 , P2_U5616 , P2_U5614 );
nand NAND3_3673 ( P2_U3092 , P2_U5618 , P2_U5619 , P2_U5617 );
nand NAND3_3674 ( P2_U3093 , P2_U5621 , P2_U5622 , P2_U5620 );
nand NAND3_3675 ( P2_U3094 , P2_U5624 , P2_U5625 , P2_U5623 );
nand NAND3_3676 ( P2_U3095 , P2_U5627 , P2_U5628 , P2_U5626 );
nand NAND3_3677 ( P2_U3096 , P2_U5630 , P2_U5631 , P2_U5629 );
nand NAND3_3678 ( P2_U3097 , P2_U5636 , P2_U5637 , P2_U5635 );
nand NAND3_3679 ( P2_U3098 , P2_U5639 , P2_U5640 , P2_U5638 );
nand NAND3_3680 ( P2_U3099 , P2_U5642 , P2_U5643 , P2_U5641 );
nand NAND3_3681 ( P2_U3100 , P2_U5645 , P2_U5646 , P2_U5644 );
nand NAND3_3682 ( P2_U3101 , P2_U5648 , P2_U5649 , P2_U5647 );
nand NAND3_3683 ( P2_U3102 , P2_U5651 , P2_U5652 , P2_U5650 );
nand NAND3_3684 ( P2_U3103 , P2_U5654 , P2_U5655 , P2_U5653 );
nand NAND3_3685 ( P2_U3104 , P2_U5657 , P2_U5658 , P2_U5656 );
nand NAND3_3686 ( P2_U3105 , P2_U5660 , P2_U5659 , P2_U5661 );
nand NAND3_3687 ( P2_U3106 , P2_U5663 , P2_U5662 , P2_U5664 );
nand NAND3_3688 ( P2_U3107 , P2_U5578 , P2_U5577 , P2_U5579 );
nand NAND3_3689 ( P2_U3108 , P2_U5581 , P2_U5580 , P2_U5582 );
nand NAND3_3690 ( P2_U3109 , P2_U5584 , P2_U5583 , P2_U5585 );
nand NAND3_3691 ( P2_U3110 , P2_U5587 , P2_U5586 , P2_U5588 );
nand NAND3_3692 ( P2_U3111 , P2_U5590 , P2_U5589 , P2_U5591 );
nand NAND3_3693 ( P2_U3112 , P2_U5593 , P2_U5592 , P2_U5594 );
nand NAND3_3694 ( P2_U3113 , P2_U5601 , P2_U5599 , P2_U5600 );
nand NAND3_3695 ( P2_U3114 , P2_U5633 , P2_U5632 , P2_U5634 );
nand NAND3_3696 ( P2_U3115 , P2_U5666 , P2_U5665 , P2_U5667 );
nand NAND2_3697 ( P2_U3116 , P2_U5669 , P2_U5668 );
nand NAND2_3698 ( P2_U3117 , P2_U5527 , P2_U5526 );
and AND2_3699 ( P2_U3118 , P2_U5673 , P2_U5672 );
nand NAND3_3700 ( P2_U3119 , P2_U3436 , P2_U5531 , P2_U5532 );
nand NAND3_3701 ( P2_U3120 , P2_U3436 , P2_U5533 , P2_U5534 );
nand NAND3_3702 ( P2_U3121 , P2_U3436 , P2_U5535 , P2_U5536 );
nand NAND3_3703 ( P2_U3122 , P2_U3436 , P2_U5537 , P2_U5538 );
nand NAND3_3704 ( P2_U3123 , P2_U3436 , P2_U5539 , P2_U5540 );
nand NAND3_3705 ( P2_U3124 , P2_U3436 , P2_U5541 , P2_U5542 );
nand NAND3_3706 ( P2_U3125 , P2_U3436 , P2_U5543 , P2_U5544 );
nand NAND3_3707 ( P2_U3126 , P2_U3436 , P2_U5545 , P2_U5546 );
nand NAND3_3708 ( P2_U3127 , P2_U3436 , P2_U5547 , P2_U5548 );
nand NAND3_3709 ( P2_U3128 , P2_U3436 , P2_U5549 , P2_U5550 );
nand NAND3_3710 ( P2_U3129 , P2_U5554 , P2_U3436 , P2_U5553 );
nand NAND3_3711 ( P2_U3130 , P2_U5556 , P2_U3436 , P2_U5555 );
nand NAND3_3712 ( P2_U3131 , P2_U5558 , P2_U3436 , P2_U5557 );
nand NAND3_3713 ( P2_U3132 , P2_U5560 , P2_U3436 , P2_U5559 );
nand NAND3_3714 ( P2_U3133 , P2_U5562 , P2_U3436 , P2_U5561 );
nand NAND3_3715 ( P2_U3134 , P2_U5564 , P2_U3436 , P2_U5563 );
nand NAND3_3716 ( P2_U3135 , P2_U5566 , P2_U3436 , P2_U5565 );
nand NAND3_3717 ( P2_U3136 , P2_U5568 , P2_U3436 , P2_U5567 );
nand NAND3_3718 ( P2_U3137 , P2_U3436 , P2_U5569 , P2_U5570 );
nand NAND3_3719 ( P2_U3138 , P2_U3436 , P2_U5571 , P2_U5572 );
nand NAND3_3720 ( P2_U3139 , P2_U3436 , P2_U5514 , P2_U5515 );
nand NAND3_3721 ( P2_U3140 , P2_U3436 , P2_U5516 , P2_U5517 );
nand NAND3_3722 ( P2_U3141 , P2_U3436 , P2_U5518 , P2_U5519 );
nand NAND3_3723 ( P2_U3142 , P2_U3436 , P2_U5520 , P2_U5521 );
nand NAND3_3724 ( P2_U3143 , P2_U3436 , P2_U5522 , P2_U5523 );
nand NAND3_3725 ( P2_U3144 , P2_U3436 , P2_U5524 , P2_U5525 );
nand NAND3_3726 ( P2_U3145 , P2_U3436 , P2_U5529 , P2_U5530 );
nand NAND3_3727 ( P2_U3146 , P2_U3436 , P2_U5551 , P2_U5552 );
nand NAND3_3728 ( P2_U3147 , P2_U3436 , P2_U5573 , P2_U5574 );
nand NAND3_3729 ( P2_U3148 , P2_U3436 , P2_U5575 , P2_U5576 );
nand NAND3_3730 ( P2_U3149 , P2_U3436 , P2_U5511 , P2_U3440 );
nand NAND2_3731 ( P2_U3150 , P2_U3905 , P2_U3982 );
nand NAND2_3732 ( P2_U3151 , P2_U3903 , P2_U5446 );
not NOT1_3733 ( P2_U3152 , P2_STATE_REG );
nand NAND2_3734 ( P2_U3153 , P2_U5463 , P2_U5462 );
nand NAND2_3735 ( P2_U3154 , P2_U5465 , P2_U5464 );
nand NAND2_3736 ( P2_U3155 , P2_U5469 , P2_U5468 );
nand NAND2_3737 ( P2_U3156 , P2_U5471 , P2_U5470 );
nand NAND2_3738 ( P2_U3157 , P2_U5473 , P2_U5472 );
nand NAND2_3739 ( P2_U3158 , P2_U5475 , P2_U5474 );
nand NAND2_3740 ( P2_U3159 , P2_U5477 , P2_U5476 );
nand NAND2_3741 ( P2_U3160 , P2_U5479 , P2_U5478 );
nand NAND2_3742 ( P2_U3161 , P2_U5481 , P2_U5480 );
nand NAND2_3743 ( P2_U3162 , P2_U5483 , P2_U5482 );
nand NAND2_3744 ( P2_U3163 , P2_U5485 , P2_U5484 );
nand NAND2_3745 ( P2_U3164 , P2_U5487 , P2_U5486 );
nand NAND2_3746 ( P2_U3165 , P2_U5490 , P2_U5489 );
nand NAND2_3747 ( P2_U3166 , P2_U5492 , P2_U5491 );
nand NAND2_3748 ( P2_U3167 , P2_U5494 , P2_U5493 );
nand NAND2_3749 ( P2_U3168 , P2_U5496 , P2_U5495 );
nand NAND2_3750 ( P2_U3169 , P2_U5498 , P2_U5497 );
nand NAND2_3751 ( P2_U3170 , P2_U5500 , P2_U5499 );
nand NAND2_3752 ( P2_U3171 , P2_U5502 , P2_U5501 );
nand NAND2_3753 ( P2_U3172 , P2_U5504 , P2_U5503 );
nand NAND2_3754 ( P2_U3173 , P2_U5506 , P2_U5505 );
nand NAND2_3755 ( P2_U3174 , P2_U5508 , P2_U5507 );
nand NAND2_3756 ( P2_U3175 , P2_U5451 , P2_U5450 );
nand NAND2_3757 ( P2_U3176 , P2_U5453 , P2_U5452 );
nand NAND2_3758 ( P2_U3177 , P2_U5455 , P2_U5454 );
nand NAND2_3759 ( P2_U3178 , P2_U5457 , P2_U5456 );
nand NAND2_3760 ( P2_U3179 , P2_U5459 , P2_U5458 );
nand NAND2_3761 ( P2_U3180 , P2_U5461 , P2_U5460 );
nand NAND2_3762 ( P2_U3181 , P2_U5467 , P2_U5466 );
and AND2_3763 ( P2_U3182 , P2_U5683 , P2_U5679 );
and AND2_3764 ( P2_U3183 , P2_U5682 , P2_U5680 );
and AND2_3765 ( P2_U3184 , P2_U5684 , P2_U5681 );
and AND2_3766 ( P2_U3185 , P2_U5448 , P2_U3054 );
and AND2_3767 ( P2_U3186 , P2_U5448 , P2_U3053 );
and AND2_3768 ( P2_U3187 , P2_U5448 , P2_U3057 );
and AND2_3769 ( P2_U3188 , P2_U5448 , P2_U3058 );
and AND2_3770 ( P2_U3189 , P2_U5448 , P2_U3065 );
and AND2_3771 ( P2_U3190 , P2_U5448 , P2_U3066 );
and AND2_3772 ( P2_U3191 , P2_U5448 , P2_U3061 );
and AND2_3773 ( P2_U3192 , P2_U5448 , P2_U3075 );
and AND2_3774 ( P2_U3193 , P2_U5448 , P2_U3076 );
and AND2_3775 ( P2_U3194 , P2_U5448 , P2_U3081 );
and AND2_3776 ( P2_U3195 , P2_U5448 , P2_U3082 );
and AND2_3777 ( P2_U3196 , P2_U5448 , P2_U3069 );
and AND2_3778 ( P2_U3197 , P2_U5448 , P2_U3073 );
and AND2_3779 ( P2_U3198 , P2_U5448 , P2_U3074 );
and AND2_3780 ( P2_U3199 , P2_U5448 , P2_U3079 );
and AND2_3781 ( P2_U3200 , P2_U5448 , P2_U3080 );
and AND2_3782 ( P2_U3201 , P2_U5448 , P2_U3072 );
and AND2_3783 ( P2_U3202 , P2_U5448 , P2_U3063 );
and AND2_3784 ( P2_U3203 , P2_U5448 , P2_U3062 );
and AND2_3785 ( P2_U3204 , P2_U5448 , P2_U3083 );
and AND2_3786 ( P2_U3205 , P2_U5448 , P2_U3084 );
and AND2_3787 ( P2_U3206 , P2_U5448 , P2_U3070 );
and AND2_3788 ( P2_U3207 , P2_U5448 , P2_U3071 );
and AND2_3789 ( P2_U3208 , P2_U5448 , P2_U3067 );
and AND2_3790 ( P2_U3209 , P2_U5448 , P2_U3060 );
and AND2_3791 ( P2_U3210 , P2_U5448 , P2_U3064 );
and AND2_3792 ( P2_U3211 , P2_U5448 , P2_U3068 );
and AND2_3793 ( P2_U3212 , P2_U5448 , P2_U3078 );
and AND2_3794 ( P2_U3213 , P2_U5448 , P2_U3077 );
nand NAND3_3795 ( P2_U3214 , P2_U6270 , P2_U6269 , P2_U3370 );
nand NAND5_3796 ( P2_U3215 , P2_U5442 , P2_U5441 , P2_U5445 , P2_U5443 , P2_U5444 );
nand NAND5_3797 ( P2_U3216 , P2_U5433 , P2_U5434 , P2_U5436 , P2_U5432 , P2_U5435 );
nand NAND5_3798 ( P2_U3217 , P2_U5424 , P2_U5423 , P2_U5427 , P2_U5425 , P2_U5426 );
nand NAND5_3799 ( P2_U3218 , P2_U5415 , P2_U5416 , P2_U5418 , P2_U5414 , P2_U5417 );
nand NAND5_3800 ( P2_U3219 , P2_U5406 , P2_U5405 , P2_U5409 , P2_U5407 , P2_U5408 );
nand NAND3_3801 ( P2_U3220 , P2_U3901 , P2_U5397 , P2_U5398 );
nand NAND4_3802 ( P2_U3221 , P2_U5388 , P2_U5389 , P2_U3900 , P2_U5390 );
nand NAND5_3803 ( P2_U3222 , P2_U5379 , P2_U5380 , P2_U5382 , P2_U5378 , P2_U5381 );
nand NAND5_3804 ( P2_U3223 , P2_U5370 , P2_U5369 , P2_U5373 , P2_U5371 , P2_U5372 );
nand NAND3_3805 ( P2_U3224 , P2_U3898 , P2_U5361 , P2_U5362 );
nand NAND5_3806 ( P2_U3225 , P2_U5352 , P2_U5353 , P2_U5355 , P2_U5351 , P2_U5354 );
nand NAND5_3807 ( P2_U3226 , P2_U5343 , P2_U5342 , P2_U5346 , P2_U5344 , P2_U5345 );
nand NAND5_3808 ( P2_U3227 , P2_U5334 , P2_U5335 , P2_U5337 , P2_U5333 , P2_U5336 );
nand NAND5_3809 ( P2_U3228 , P2_U5325 , P2_U5324 , P2_U5328 , P2_U5326 , P2_U5327 );
nand NAND4_3810 ( P2_U3229 , P2_U5316 , P2_U5315 , P2_U5317 , P2_U3897 );
nand NAND5_3811 ( P2_U3230 , P2_U5307 , P2_U5306 , P2_U5310 , P2_U5308 , P2_U5309 );
nand NAND5_3812 ( P2_U3231 , P2_U5298 , P2_U5299 , P2_U5301 , P2_U5297 , P2_U5300 );
nand NAND4_3813 ( P2_U3232 , P2_U5289 , P2_U5288 , P2_U3896 , P2_U5290 );
nand NAND5_3814 ( P2_U3233 , P2_U5280 , P2_U5279 , P2_U5283 , P2_U5281 , P2_U5282 );
nand NAND3_3815 ( P2_U3234 , P2_U3895 , P2_U5272 , P2_U3894 );
nand NAND5_3816 ( P2_U3235 , P2_U5263 , P2_U5264 , P2_U5266 , P2_U5262 , P2_U5265 );
nand NAND5_3817 ( P2_U3236 , P2_U5254 , P2_U5253 , P2_U5257 , P2_U5255 , P2_U5256 );
nand NAND5_3818 ( P2_U3237 , P2_U5245 , P2_U5246 , P2_U5248 , P2_U5244 , P2_U5247 );
nand NAND5_3819 ( P2_U3238 , P2_U5236 , P2_U5235 , P2_U5239 , P2_U5237 , P2_U5238 );
nand NAND3_3820 ( P2_U3239 , P2_U3891 , P2_U5227 , P2_U5228 );
nand NAND5_3821 ( P2_U3240 , P2_U5218 , P2_U5217 , P2_U5221 , P2_U5219 , P2_U5220 );
nand NAND5_3822 ( P2_U3241 , P2_U5209 , P2_U5208 , P2_U5212 , P2_U5210 , P2_U5211 );
nand NAND5_3823 ( P2_U3242 , P2_U5200 , P2_U5201 , P2_U5203 , P2_U5199 , P2_U5202 );
nand NAND5_3824 ( P2_U3243 , P2_U5187 , P2_U5186 , P2_U5190 , P2_U5188 , P2_U5189 );
and AND2_3825 ( P2_U3244 , P2_U5671 , P2_U5174 );
nand NAND2_3826 ( P2_U3245 , P2_U3872 , P2_U3871 );
nand NAND2_3827 ( P2_U3246 , P2_U3868 , P2_U3867 );
nand NAND2_3828 ( P2_U3247 , P2_U3865 , P2_U3864 );
nand NAND2_3829 ( P2_U3248 , P2_U3862 , P2_U3861 );
nand NAND2_3830 ( P2_U3249 , P2_U3859 , P2_U3858 );
nand NAND2_3831 ( P2_U3250 , P2_U3856 , P2_U3855 );
nand NAND2_3832 ( P2_U3251 , P2_U3853 , P2_U3852 );
nand NAND2_3833 ( P2_U3252 , P2_U3850 , P2_U3849 );
nand NAND2_3834 ( P2_U3253 , P2_U3847 , P2_U3846 );
nand NAND3_3835 ( P2_U3254 , P2_U3843 , P2_U3844 , P2_U3842 );
nand NAND3_3836 ( P2_U3255 , P2_U3840 , P2_U3841 , P2_U3839 );
nand NAND3_3837 ( P2_U3256 , P2_U3837 , P2_U3838 , P2_U3836 );
nand NAND3_3838 ( P2_U3257 , P2_U3834 , P2_U3835 , P2_U3833 );
nand NAND3_3839 ( P2_U3258 , P2_U3831 , P2_U3832 , P2_U3830 );
nand NAND3_3840 ( P2_U3259 , P2_U3828 , P2_U3829 , P2_U3827 );
nand NAND3_3841 ( P2_U3260 , P2_U3825 , P2_U3826 , P2_U3824 );
nand NAND3_3842 ( P2_U3261 , P2_U3822 , P2_U3823 , P2_U3821 );
nand NAND3_3843 ( P2_U3262 , P2_U3819 , P2_U3820 , P2_U3818 );
nand NAND3_3844 ( P2_U3263 , P2_U3816 , P2_U3817 , P2_U3815 );
nand NAND3_3845 ( P2_U3264 , P2_U3813 , P2_U3814 , P2_U3812 );
nand NAND3_3846 ( P2_U3265 , P2_U3944 , P2_U4865 , P2_U4866 );
nand NAND3_3847 ( P2_U3266 , P2_U3943 , P2_U4863 , P2_U4864 );
nand NAND5_3848 ( P2_U3267 , P2_U4860 , P2_U4861 , P2_U4862 , P2_U4859 , P2_U3941 );
nand NAND4_3849 ( P2_U3268 , P2_U3808 , P2_U3809 , P2_U4855 , P2_U3940 );
nand NAND4_3850 ( P2_U3269 , P2_U3806 , P2_U3807 , P2_U4850 , P2_U3939 );
nand NAND4_3851 ( P2_U3270 , P2_U3804 , P2_U3805 , P2_U4845 , P2_U3938 );
nand NAND4_3852 ( P2_U3271 , P2_U3802 , P2_U3803 , P2_U4840 , P2_U3937 );
nand NAND4_3853 ( P2_U3272 , P2_U3800 , P2_U3801 , P2_U4835 , P2_U3936 );
nand NAND4_3854 ( P2_U3273 , P2_U3798 , P2_U3799 , P2_U4830 , P2_U3935 );
nand NAND4_3855 ( P2_U3274 , P2_U3796 , P2_U3797 , P2_U4825 , P2_U3934 );
nand NAND4_3856 ( P2_U3275 , P2_U3794 , P2_U3795 , P2_U4820 , P2_U3933 );
nand NAND4_3857 ( P2_U3276 , P2_U3792 , P2_U3793 , P2_U4815 , P2_U3932 );
nand NAND4_3858 ( P2_U3277 , P2_U3790 , P2_U3791 , P2_U4810 , P2_U3931 );
nand NAND4_3859 ( P2_U3278 , P2_U3788 , P2_U3789 , P2_U4805 , P2_U3930 );
nand NAND4_3860 ( P2_U3279 , P2_U3786 , P2_U3787 , P2_U4800 , P2_U3929 );
nand NAND4_3861 ( P2_U3280 , P2_U3784 , P2_U3785 , P2_U4795 , P2_U3928 );
nand NAND4_3862 ( P2_U3281 , P2_U3782 , P2_U3783 , P2_U4790 , P2_U3927 );
nand NAND4_3863 ( P2_U3282 , P2_U3780 , P2_U3781 , P2_U4785 , P2_U3926 );
nand NAND4_3864 ( P2_U3283 , P2_U3778 , P2_U3779 , P2_U4780 , P2_U3925 );
nand NAND4_3865 ( P2_U3284 , P2_U3776 , P2_U3777 , P2_U4775 , P2_U3924 );
nand NAND3_3866 ( P2_U3285 , P2_U3775 , P2_U3774 , P2_U3923 );
nand NAND4_3867 ( P2_U3286 , P2_U3772 , P2_U3773 , P2_U4765 , P2_U3922 );
nand NAND3_3868 ( P2_U3287 , P2_U3771 , P2_U3770 , P2_U3921 );
nand NAND3_3869 ( P2_U3288 , P2_U3769 , P2_U3768 , P2_U3920 );
nand NAND3_3870 ( P2_U3289 , P2_U3767 , P2_U3766 , P2_U3919 );
nand NAND3_3871 ( P2_U3290 , P2_U3765 , P2_U3764 , P2_U3918 );
nand NAND3_3872 ( P2_U3291 , P2_U3763 , P2_U3762 , P2_U3917 );
nand NAND2_3873 ( P2_U3292 , P2_U3761 , P2_U3760 );
nand NAND2_3874 ( P2_U3293 , P2_U3759 , P2_U3758 );
nand NAND2_3875 ( P2_U3294 , P2_U3757 , P2_U3756 );
nand NAND2_3876 ( P2_U3295 , P2_U3755 , P2_U3754 );
nand NAND2_3877 ( P2_U3296 , P2_U3753 , P2_U3752 );
and AND2_3878 ( P2_U3297 , P2_D_REG_31_ , P2_U3908 );
and AND2_3879 ( P2_U3298 , P2_D_REG_30_ , P2_U3908 );
and AND2_3880 ( P2_U3299 , P2_D_REG_29_ , P2_U3908 );
and AND2_3881 ( P2_U3300 , P2_D_REG_28_ , P2_U3908 );
and AND2_3882 ( P2_U3301 , P2_D_REG_27_ , P2_U3908 );
and AND2_3883 ( P2_U3302 , P2_D_REG_26_ , P2_U3908 );
and AND2_3884 ( P2_U3303 , P2_D_REG_25_ , P2_U3908 );
and AND2_3885 ( P2_U3304 , P2_D_REG_24_ , P2_U3908 );
and AND2_3886 ( P2_U3305 , P2_D_REG_23_ , P2_U3908 );
and AND2_3887 ( P2_U3306 , P2_D_REG_22_ , P2_U3908 );
and AND2_3888 ( P2_U3307 , P2_D_REG_21_ , P2_U3908 );
and AND2_3889 ( P2_U3308 , P2_D_REG_20_ , P2_U3908 );
and AND2_3890 ( P2_U3309 , P2_D_REG_19_ , P2_U3908 );
and AND2_3891 ( P2_U3310 , P2_D_REG_18_ , P2_U3908 );
and AND2_3892 ( P2_U3311 , P2_D_REG_17_ , P2_U3908 );
and AND2_3893 ( P2_U3312 , P2_D_REG_16_ , P2_U3908 );
and AND2_3894 ( P2_U3313 , P2_D_REG_15_ , P2_U3908 );
and AND2_3895 ( P2_U3314 , P2_D_REG_14_ , P2_U3908 );
and AND2_3896 ( P2_U3315 , P2_D_REG_13_ , P2_U3908 );
and AND2_3897 ( P2_U3316 , P2_D_REG_12_ , P2_U3908 );
and AND2_3898 ( P2_U3317 , P2_D_REG_11_ , P2_U3908 );
and AND2_3899 ( P2_U3318 , P2_D_REG_10_ , P2_U3908 );
and AND2_3900 ( P2_U3319 , P2_D_REG_9_ , P2_U3908 );
and AND2_3901 ( P2_U3320 , P2_D_REG_8_ , P2_U3908 );
and AND2_3902 ( P2_U3321 , P2_D_REG_7_ , P2_U3908 );
and AND2_3903 ( P2_U3322 , P2_D_REG_6_ , P2_U3908 );
and AND2_3904 ( P2_U3323 , P2_D_REG_5_ , P2_U3908 );
and AND2_3905 ( P2_U3324 , P2_D_REG_4_ , P2_U3908 );
and AND2_3906 ( P2_U3325 , P2_D_REG_3_ , P2_U3908 );
and AND2_3907 ( P2_U3326 , P2_D_REG_2_ , P2_U3908 );
nand NAND3_3908 ( P2_U3327 , P2_U4091 , P2_U4092 , P2_U4090 );
nand NAND3_3909 ( P2_U3328 , P2_U4088 , P2_U4089 , P2_U4087 );
nand NAND3_3910 ( P2_U3329 , P2_U4085 , P2_U4086 , P2_U4084 );
nand NAND3_3911 ( P2_U3330 , P2_U4082 , P2_U4083 , P2_U4081 );
nand NAND3_3912 ( P2_U3331 , P2_U4079 , P2_U4080 , P2_U4078 );
nand NAND3_3913 ( P2_U3332 , P2_U4076 , P2_U4077 , P2_U4075 );
nand NAND3_3914 ( P2_U3333 , P2_U4073 , P2_U4074 , P2_U4072 );
nand NAND3_3915 ( P2_U3334 , P2_U4070 , P2_U4071 , P2_U4069 );
nand NAND3_3916 ( P2_U3335 , P2_U4067 , P2_U4068 , P2_U4066 );
nand NAND3_3917 ( P2_U3336 , P2_U4064 , P2_U4065 , P2_U4063 );
nand NAND3_3918 ( P2_U3337 , P2_U4061 , P2_U4062 , P2_U4060 );
nand NAND3_3919 ( P2_U3338 , P2_U4058 , P2_U4059 , P2_U4057 );
nand NAND3_3920 ( P2_U3339 , P2_U4055 , P2_U4056 , P2_U4054 );
nand NAND3_3921 ( P2_U3340 , P2_U4052 , P2_U4053 , P2_U4051 );
nand NAND3_3922 ( P2_U3341 , P2_U4049 , P2_U4050 , P2_U4048 );
nand NAND3_3923 ( P2_U3342 , P2_U4046 , P2_U4047 , P2_U4045 );
nand NAND3_3924 ( P2_U3343 , P2_U4043 , P2_U4044 , P2_U4042 );
nand NAND3_3925 ( P2_U3344 , P2_U4040 , P2_U4041 , P2_U4039 );
nand NAND3_3926 ( P2_U3345 , P2_U4037 , P2_U4038 , P2_U4036 );
nand NAND3_3927 ( P2_U3346 , P2_U4034 , P2_U4035 , P2_U4033 );
nand NAND3_3928 ( P2_U3347 , P2_U4031 , P2_U4032 , P2_U4030 );
nand NAND3_3929 ( P2_U3348 , P2_U4028 , P2_U4029 , P2_U4027 );
nand NAND3_3930 ( P2_U3349 , P2_U4025 , P2_U4026 , P2_U4024 );
nand NAND3_3931 ( P2_U3350 , P2_U4022 , P2_U4023 , P2_U4021 );
nand NAND3_3932 ( P2_U3351 , P2_U4019 , P2_U4020 , P2_U4018 );
nand NAND3_3933 ( P2_U3352 , P2_U4016 , P2_U4017 , P2_U4015 );
nand NAND3_3934 ( P2_U3353 , P2_U4013 , P2_U4014 , P2_U4012 );
nand NAND3_3935 ( P2_U3354 , P2_U4010 , P2_U4011 , P2_U4009 );
nand NAND3_3936 ( P2_U3355 , P2_U4007 , P2_U4008 , P2_U4006 );
nand NAND3_3937 ( P2_U3356 , P2_U4004 , P2_U4005 , P2_U4003 );
nand NAND3_3938 ( P2_U3357 , P2_U4001 , P2_U4002 , P2_U4000 );
nand NAND3_3939 ( P2_U3358 , P2_U3998 , P2_U3999 , P2_U3997 );
nand NAND2_3940 ( P2_U3359 , P2_STATE_REG , P2_U3907 );
not NOT1_3941 ( P2_U3360 , P2_B_REG );
nand NAND2_3942 ( P2_U3361 , P2_U3435 , P2_U5692 );
nand NAND2_3943 ( P2_U3362 , P2_U3435 , P2_U4093 );
nand NAND2_3944 ( P2_U3363 , P2_U3050 , P2_U3441 );
nand NAND3_3945 ( P2_U3364 , P2_U5711 , P2_U3439 , P2_U3440 );
nand NAND2_3946 ( P2_U3365 , P2_U5714 , P2_U5711 );
nand NAND2_3947 ( P2_U3366 , P2_U3994 , P2_U3441 );
nand NAND2_3948 ( P2_U3367 , P2_U3961 , P2_U5717 );
nand NAND2_3949 ( P2_U3368 , P2_U5708 , P2_U5711 );
nand NAND2_3950 ( P2_U3369 , P2_U3951 , P2_U3440 );
nand NAND2_3951 ( P2_U3370 , P2_U5708 , P2_U5717 );
nand NAND2_3952 ( P2_U3371 , P2_U3440 , P2_U3441 );
nand NAND3_3953 ( P2_U3372 , P2_U5711 , P2_U3439 , P2_U5717 );
nand NAND5_3954 ( P2_U3373 , P2_U4138 , P2_U4137 , P2_U4139 , P2_U3617 , P2_U3616 );
nand NAND4_3955 ( P2_U3374 , P2_U4153 , P2_U4152 , P2_U3632 , P2_U3634 );
nand NAND4_3956 ( P2_U3375 , P2_U4172 , P2_U4171 , P2_U3636 , P2_U3638 );
nand NAND4_3957 ( P2_U3376 , P2_U4191 , P2_U4190 , P2_U3640 , P2_U3642 );
nand NAND4_3958 ( P2_U3377 , P2_U4210 , P2_U4209 , P2_U3644 , P2_U3646 );
nand NAND4_3959 ( P2_U3378 , P2_U4229 , P2_U4228 , P2_U3648 , P2_U3650 );
nand NAND4_3960 ( P2_U3379 , P2_U4248 , P2_U4247 , P2_U3652 , P2_U3654 );
nand NAND4_3961 ( P2_U3380 , P2_U4267 , P2_U4266 , P2_U3656 , P2_U3658 );
nand NAND4_3962 ( P2_U3381 , P2_U4286 , P2_U4285 , P2_U3660 , P2_U3662 );
nand NAND4_3963 ( P2_U3382 , P2_U4305 , P2_U4304 , P2_U3664 , P2_U3666 );
nand NAND4_3964 ( P2_U3383 , P2_U4324 , P2_U4323 , P2_U3668 , P2_U3670 );
nand NAND4_3965 ( P2_U3384 , P2_U4343 , P2_U4342 , P2_U3672 , P2_U3674 );
nand NAND4_3966 ( P2_U3385 , P2_U4362 , P2_U4361 , P2_U3676 , P2_U3678 );
nand NAND4_3967 ( P2_U3386 , P2_U4381 , P2_U4380 , P2_U3680 , P2_U3682 );
nand NAND4_3968 ( P2_U3387 , P2_U4400 , P2_U4399 , P2_U3684 , P2_U3686 );
nand NAND4_3969 ( P2_U3388 , P2_U4419 , P2_U4418 , P2_U3688 , P2_U3690 );
nand NAND4_3970 ( P2_U3389 , P2_U4438 , P2_U4437 , P2_U3692 , P2_U3694 );
nand NAND4_3971 ( P2_U3390 , P2_U4457 , P2_U4456 , P2_U3696 , P2_U3698 );
nand NAND4_3972 ( P2_U3391 , P2_U4476 , P2_U4475 , P2_U3700 , P2_U3702 );
nand NAND4_3973 ( P2_U3392 , P2_U4495 , P2_U4494 , P2_U3704 , P2_U3706 );
nand NAND2_3974 ( P2_U3393 , U44 , P2_U3909 );
nand NAND4_3975 ( P2_U3394 , P2_U4514 , P2_U4513 , P2_U3708 , P2_U3710 );
nand NAND2_3976 ( P2_U3395 , U43 , P2_U3909 );
nand NAND4_3977 ( P2_U3396 , P2_U4533 , P2_U4532 , P2_U3712 , P2_U3714 );
nand NAND2_3978 ( P2_U3397 , U42 , P2_U3909 );
nand NAND4_3979 ( P2_U3398 , P2_U4552 , P2_U4551 , P2_U3716 , P2_U3718 );
nand NAND2_3980 ( P2_U3399 , U41 , P2_U3909 );
nand NAND4_3981 ( P2_U3400 , P2_U4571 , P2_U4570 , P2_U3720 , P2_U3722 );
nand NAND2_3982 ( P2_U3401 , U40 , P2_U3909 );
nand NAND4_3983 ( P2_U3402 , P2_U4590 , P2_U4589 , P2_U3724 , P2_U3726 );
nand NAND2_3984 ( P2_U3403 , U39 , P2_U3909 );
nand NAND4_3985 ( P2_U3404 , P2_U4609 , P2_U4608 , P2_U3728 , P2_U3730 );
nand NAND2_3986 ( P2_U3405 , U38 , P2_U3909 );
nand NAND4_3987 ( P2_U3406 , P2_U4628 , P2_U4627 , P2_U3732 , P2_U3734 );
nand NAND2_3988 ( P2_U3407 , U37 , P2_U3909 );
nand NAND4_3989 ( P2_U3408 , P2_U4647 , P2_U4646 , P2_U3736 , P2_U3738 );
nand NAND2_3990 ( P2_U3409 , U36 , P2_U3909 );
nand NAND5_3991 ( P2_U3410 , P2_U4666 , P2_U4665 , P2_U4667 , P2_U4668 , P2_U3741 );
nand NAND2_3992 ( P2_U3411 , U35 , P2_U3909 );
nand NAND5_3993 ( P2_U3412 , P2_U4686 , P2_U4685 , P2_U4687 , P2_U3744 , P2_U3746 );
nand NAND2_3994 ( P2_U3413 , U33 , P2_U3909 );
nand NAND2_3995 ( P2_U3414 , U32 , P2_U3909 );
nand NAND2_3996 ( P2_U3415 , P2_U3445 , P2_U5717 );
nand NAND2_3997 ( P2_U3416 , P2_U5674 , P2_U5714 );
nand NAND2_3998 ( P2_U3417 , P2_U3027 , P2_U4711 );
nand NAND2_3999 ( P2_U3418 , P2_U3960 , P2_U5708 );
nand NAND2_4000 ( P2_U3419 , P2_U3031 , P2_U5711 );
nand NAND3_4001 ( P2_U3420 , P2_U3434 , P2_U3435 , P2_U3433 );
nand NAND2_4002 ( P2_U3421 , P2_U3371 , P2_U3909 );
nand NAND2_4003 ( P2_U3422 , P2_U3981 , P2_U5701 );
nand NAND2_4004 ( P2_U3423 , P2_U3995 , P2_STATE_REG );
nand NAND2_4005 ( P2_U3424 , P2_U3810 , P2_U3052 );
nand NAND2_4006 ( P2_U3425 , P2_U3017 , P2_U3022 );
nand NAND2_4007 ( P2_U3426 , P2_U3027 , P2_U4713 );
nand NAND2_4008 ( P2_U3427 , P2_U3887 , P2_U3020 );
nand NAND2_4009 ( P2_U3428 , P2_U5708 , P2_U3440 );
nand NAND2_4010 ( P2_U3429 , P2_U3017 , P2_U3027 );
nand NAND2_4011 ( P2_U3430 , P2_U5184 , P2_U3889 );
nand NAND2_4012 ( P2_U3431 , P2_U3951 , P2_U3369 );
nand NAND2_4013 ( P2_U3432 , P2_U3993 , P2_U3445 );
nand NAND2_4014 ( P2_U3433 , P2_U5688 , P2_U5687 );
nand NAND2_4015 ( P2_U3434 , P2_U5691 , P2_U5690 );
nand NAND2_4016 ( P2_U3435 , P2_U5694 , P2_U5693 );
nand NAND2_4017 ( P2_U3436 , P2_U5700 , P2_U5699 );
nand NAND2_4018 ( P2_U3437 , P2_U5703 , P2_U5702 );
nand NAND2_4019 ( P2_U3438 , P2_U5705 , P2_U5704 );
nand NAND2_4020 ( P2_U3439 , P2_U5713 , P2_U5712 );
nand NAND2_4021 ( P2_U3440 , P2_U5716 , P2_U5715 );
nand NAND2_4022 ( P2_U3441 , P2_U5707 , P2_U5706 );
nand NAND2_4023 ( P2_U3442 , P2_U5722 , P2_U5721 );
nand NAND2_4024 ( P2_U3443 , P2_U5719 , P2_U5718 );
nand NAND2_4025 ( P2_U3444 , P2_U5727 , P2_U5726 );
nand NAND2_4026 ( P2_U3445 , P2_U5710 , P2_U5709 );
nand NAND2_4027 ( P2_U3446 , P2_U5730 , P2_U5729 );
nand NAND2_4028 ( P2_U3447 , P2_U5732 , P2_U5731 );
nand NAND2_4029 ( P2_U3448 , P2_U5735 , P2_U5734 );
nand NAND2_4030 ( P2_U3449 , P2_U5743 , P2_U5742 );
nand NAND2_4031 ( P2_U3450 , P2_U5740 , P2_U5739 );
nand NAND2_4032 ( P2_U3451 , P2_U5746 , P2_U5745 );
nand NAND2_4033 ( P2_U3452 , P2_U5750 , P2_U5749 );
nand NAND2_4034 ( P2_U3453 , P2_U5752 , P2_U5751 );
nand NAND2_4035 ( P2_U3454 , P2_U5757 , P2_U5756 );
nand NAND2_4036 ( P2_U3455 , P2_U5759 , P2_U5758 );
nand NAND2_4037 ( P2_U3456 , P2_U5761 , P2_U5760 );
nand NAND2_4038 ( P2_U3457 , P2_U5764 , P2_U5763 );
nand NAND2_4039 ( P2_U3458 , P2_U5766 , P2_U5765 );
nand NAND2_4040 ( P2_U3459 , P2_U5768 , P2_U5767 );
nand NAND2_4041 ( P2_U3460 , P2_U5771 , P2_U5770 );
nand NAND2_4042 ( P2_U3461 , P2_U5773 , P2_U5772 );
nand NAND2_4043 ( P2_U3462 , P2_U5775 , P2_U5774 );
nand NAND2_4044 ( P2_U3463 , P2_U5778 , P2_U5777 );
nand NAND2_4045 ( P2_U3464 , P2_U5780 , P2_U5779 );
nand NAND2_4046 ( P2_U3465 , P2_U5782 , P2_U5781 );
nand NAND2_4047 ( P2_U3466 , P2_U5785 , P2_U5784 );
nand NAND2_4048 ( P2_U3467 , P2_U5787 , P2_U5786 );
nand NAND2_4049 ( P2_U3468 , P2_U5789 , P2_U5788 );
nand NAND2_4050 ( P2_U3469 , P2_U5792 , P2_U5791 );
nand NAND2_4051 ( P2_U3470 , P2_U5794 , P2_U5793 );
nand NAND2_4052 ( P2_U3471 , P2_U5796 , P2_U5795 );
nand NAND2_4053 ( P2_U3472 , P2_U5799 , P2_U5798 );
nand NAND2_4054 ( P2_U3473 , P2_U5801 , P2_U5800 );
nand NAND2_4055 ( P2_U3474 , P2_U5803 , P2_U5802 );
nand NAND2_4056 ( P2_U3475 , P2_U5806 , P2_U5805 );
nand NAND2_4057 ( P2_U3476 , P2_U5808 , P2_U5807 );
nand NAND2_4058 ( P2_U3477 , P2_U5810 , P2_U5809 );
nand NAND2_4059 ( P2_U3478 , P2_U5813 , P2_U5812 );
nand NAND2_4060 ( P2_U3479 , P2_U5815 , P2_U5814 );
nand NAND2_4061 ( P2_U3480 , P2_U5817 , P2_U5816 );
nand NAND2_4062 ( P2_U3481 , P2_U5820 , P2_U5819 );
nand NAND2_4063 ( P2_U3482 , P2_U5822 , P2_U5821 );
nand NAND2_4064 ( P2_U3483 , P2_U5824 , P2_U5823 );
nand NAND2_4065 ( P2_U3484 , P2_U5827 , P2_U5826 );
nand NAND2_4066 ( P2_U3485 , P2_U5829 , P2_U5828 );
nand NAND2_4067 ( P2_U3486 , P2_U5831 , P2_U5830 );
nand NAND2_4068 ( P2_U3487 , P2_U5834 , P2_U5833 );
nand NAND2_4069 ( P2_U3488 , P2_U5836 , P2_U5835 );
nand NAND2_4070 ( P2_U3489 , P2_U5838 , P2_U5837 );
nand NAND2_4071 ( P2_U3490 , P2_U5841 , P2_U5840 );
nand NAND2_4072 ( P2_U3491 , P2_U5843 , P2_U5842 );
nand NAND2_4073 ( P2_U3492 , P2_U5845 , P2_U5844 );
nand NAND2_4074 ( P2_U3493 , P2_U5848 , P2_U5847 );
nand NAND2_4075 ( P2_U3494 , P2_U5850 , P2_U5849 );
nand NAND2_4076 ( P2_U3495 , P2_U5852 , P2_U5851 );
nand NAND2_4077 ( P2_U3496 , P2_U5855 , P2_U5854 );
nand NAND2_4078 ( P2_U3497 , P2_U5857 , P2_U5856 );
nand NAND2_4079 ( P2_U3498 , P2_U5859 , P2_U5858 );
nand NAND2_4080 ( P2_U3499 , P2_U5862 , P2_U5861 );
nand NAND2_4081 ( P2_U3500 , P2_U5864 , P2_U5863 );
nand NAND2_4082 ( P2_U3501 , P2_U5866 , P2_U5865 );
nand NAND2_4083 ( P2_U3502 , P2_U5869 , P2_U5868 );
nand NAND2_4084 ( P2_U3503 , P2_U5871 , P2_U5870 );
nand NAND2_4085 ( P2_U3504 , P2_U5873 , P2_U5872 );
nand NAND2_4086 ( P2_U3505 , P2_U5876 , P2_U5875 );
nand NAND2_4087 ( P2_U3506 , P2_U5878 , P2_U5877 );
nand NAND2_4088 ( P2_U3507 , P2_U5881 , P2_U5880 );
nand NAND2_4089 ( P2_U3508 , P2_U5883 , P2_U5882 );
nand NAND2_4090 ( P2_U3509 , P2_U5885 , P2_U5884 );
nand NAND2_4091 ( P2_U3510 , P2_U5887 , P2_U5886 );
nand NAND2_4092 ( P2_U3511 , P2_U5889 , P2_U5888 );
nand NAND2_4093 ( P2_U3512 , P2_U5891 , P2_U5890 );
nand NAND2_4094 ( P2_U3513 , P2_U5893 , P2_U5892 );
nand NAND2_4095 ( P2_U3514 , P2_U5895 , P2_U5894 );
nand NAND2_4096 ( P2_U3515 , P2_U5897 , P2_U5896 );
nand NAND2_4097 ( P2_U3516 , P2_U5899 , P2_U5898 );
nand NAND2_4098 ( P2_U3517 , P2_U5901 , P2_U5900 );
nand NAND2_4099 ( P2_U3518 , P2_U5903 , P2_U5902 );
nand NAND2_4100 ( P2_U3519 , P2_U5905 , P2_U5904 );
nand NAND2_4101 ( P2_U3520 , P2_U5907 , P2_U5906 );
nand NAND2_4102 ( P2_U3521 , P2_U5909 , P2_U5908 );
nand NAND2_4103 ( P2_U3522 , P2_U5911 , P2_U5910 );
nand NAND2_4104 ( P2_U3523 , P2_U5913 , P2_U5912 );
nand NAND2_4105 ( P2_U3524 , P2_U5915 , P2_U5914 );
nand NAND2_4106 ( P2_U3525 , P2_U5917 , P2_U5916 );
nand NAND2_4107 ( P2_U3526 , P2_U5919 , P2_U5918 );
nand NAND2_4108 ( P2_U3527 , P2_U5921 , P2_U5920 );
nand NAND2_4109 ( P2_U3528 , P2_U5923 , P2_U5922 );
nand NAND2_4110 ( P2_U3529 , P2_U5925 , P2_U5924 );
nand NAND2_4111 ( P2_U3530 , P2_U5927 , P2_U5926 );
nand NAND2_4112 ( P2_U3531 , P2_U5929 , P2_U5928 );
nand NAND2_4113 ( P2_U3532 , P2_U5931 , P2_U5930 );
nand NAND2_4114 ( P2_U3533 , P2_U5933 , P2_U5932 );
nand NAND2_4115 ( P2_U3534 , P2_U5935 , P2_U5934 );
nand NAND2_4116 ( P2_U3535 , P2_U5937 , P2_U5936 );
nand NAND2_4117 ( P2_U3536 , P2_U5939 , P2_U5938 );
nand NAND2_4118 ( P2_U3537 , P2_U5941 , P2_U5940 );
nand NAND2_4119 ( P2_U3538 , P2_U5943 , P2_U5942 );
nand NAND2_4120 ( P2_U3539 , P2_U5945 , P2_U5944 );
nand NAND2_4121 ( P2_U3540 , P2_U5947 , P2_U5946 );
nand NAND2_4122 ( P2_U3541 , P2_U5949 , P2_U5948 );
nand NAND2_4123 ( P2_U3542 , P2_U5951 , P2_U5950 );
nand NAND2_4124 ( P2_U3543 , P2_U5953 , P2_U5952 );
nand NAND2_4125 ( P2_U3544 , P2_U5955 , P2_U5954 );
nand NAND2_4126 ( P2_U3545 , P2_U5957 , P2_U5956 );
nand NAND2_4127 ( P2_U3546 , P2_U5959 , P2_U5958 );
nand NAND2_4128 ( P2_U3547 , P2_U5961 , P2_U5960 );
nand NAND2_4129 ( P2_U3548 , P2_U5963 , P2_U5962 );
nand NAND2_4130 ( P2_U3549 , P2_U5965 , P2_U5964 );
nand NAND2_4131 ( P2_U3550 , P2_U5967 , P2_U5966 );
nand NAND2_4132 ( P2_U3551 , P2_U5969 , P2_U5968 );
nand NAND2_4133 ( P2_U3552 , P2_U6035 , P2_U6034 );
nand NAND2_4134 ( P2_U3553 , P2_U6037 , P2_U6036 );
nand NAND2_4135 ( P2_U3554 , P2_U6039 , P2_U6038 );
nand NAND2_4136 ( P2_U3555 , P2_U6041 , P2_U6040 );
nand NAND2_4137 ( P2_U3556 , P2_U6043 , P2_U6042 );
nand NAND2_4138 ( P2_U3557 , P2_U6045 , P2_U6044 );
nand NAND2_4139 ( P2_U3558 , P2_U6047 , P2_U6046 );
nand NAND2_4140 ( P2_U3559 , P2_U6049 , P2_U6048 );
nand NAND2_4141 ( P2_U3560 , P2_U6051 , P2_U6050 );
nand NAND2_4142 ( P2_U3561 , P2_U6053 , P2_U6052 );
nand NAND2_4143 ( P2_U3562 , P2_U6055 , P2_U6054 );
nand NAND2_4144 ( P2_U3563 , P2_U6057 , P2_U6056 );
nand NAND2_4145 ( P2_U3564 , P2_U6059 , P2_U6058 );
nand NAND2_4146 ( P2_U3565 , P2_U6061 , P2_U6060 );
nand NAND2_4147 ( P2_U3566 , P2_U6063 , P2_U6062 );
nand NAND2_4148 ( P2_U3567 , P2_U6065 , P2_U6064 );
nand NAND2_4149 ( P2_U3568 , P2_U6067 , P2_U6066 );
nand NAND2_4150 ( P2_U3569 , P2_U6069 , P2_U6068 );
nand NAND2_4151 ( P2_U3570 , P2_U6071 , P2_U6070 );
nand NAND2_4152 ( P2_U3571 , P2_U6073 , P2_U6072 );
nand NAND2_4153 ( P2_U3572 , P2_U6075 , P2_U6074 );
nand NAND2_4154 ( P2_U3573 , P2_U6077 , P2_U6076 );
nand NAND2_4155 ( P2_U3574 , P2_U6079 , P2_U6078 );
nand NAND2_4156 ( P2_U3575 , P2_U6081 , P2_U6080 );
nand NAND2_4157 ( P2_U3576 , P2_U6083 , P2_U6082 );
nand NAND2_4158 ( P2_U3577 , P2_U6085 , P2_U6084 );
nand NAND2_4159 ( P2_U3578 , P2_U6087 , P2_U6086 );
nand NAND2_4160 ( P2_U3579 , P2_U6089 , P2_U6088 );
nand NAND2_4161 ( P2_U3580 , P2_U6091 , P2_U6090 );
nand NAND2_4162 ( P2_U3581 , P2_U6093 , P2_U6092 );
nand NAND2_4163 ( P2_U3582 , P2_U6095 , P2_U6094 );
nand NAND2_4164 ( P2_U3583 , P2_U6097 , P2_U6096 );
nand NAND2_4165 ( P2_U3584 , P2_U6203 , P2_U6202 );
nand NAND2_4166 ( P2_U3585 , P2_U6205 , P2_U6204 );
nand NAND2_4167 ( P2_U3586 , P2_U6207 , P2_U6206 );
nand NAND2_4168 ( P2_U3587 , P2_U6209 , P2_U6208 );
nand NAND2_4169 ( P2_U3588 , P2_U6211 , P2_U6210 );
nand NAND2_4170 ( P2_U3589 , P2_U6213 , P2_U6212 );
nand NAND2_4171 ( P2_U3590 , P2_U6215 , P2_U6214 );
nand NAND2_4172 ( P2_U3591 , P2_U6217 , P2_U6216 );
nand NAND2_4173 ( P2_U3592 , P2_U6219 , P2_U6218 );
nand NAND2_4174 ( P2_U3593 , P2_U6221 , P2_U6220 );
nand NAND2_4175 ( P2_U3594 , P2_U6224 , P2_U6223 );
nand NAND2_4176 ( P2_U3595 , P2_U6226 , P2_U6225 );
nand NAND2_4177 ( P2_U3596 , P2_U6228 , P2_U6227 );
nand NAND2_4178 ( P2_U3597 , P2_U6230 , P2_U6229 );
nand NAND2_4179 ( P2_U3598 , P2_U6232 , P2_U6231 );
nand NAND2_4180 ( P2_U3599 , P2_U6234 , P2_U6233 );
nand NAND2_4181 ( P2_U3600 , P2_U6236 , P2_U6235 );
nand NAND2_4182 ( P2_U3601 , P2_U6238 , P2_U6237 );
nand NAND2_4183 ( P2_U3602 , P2_U6240 , P2_U6239 );
nand NAND2_4184 ( P2_U3603 , P2_U6242 , P2_U6241 );
nand NAND2_4185 ( P2_U3604 , P2_U6244 , P2_U6243 );
nand NAND2_4186 ( P2_U3605 , P2_U6247 , P2_U6246 );
nand NAND2_4187 ( P2_U3606 , P2_U6249 , P2_U6248 );
nand NAND2_4188 ( P2_U3607 , P2_U6251 , P2_U6250 );
nand NAND2_4189 ( P2_U3608 , P2_U6253 , P2_U6252 );
nand NAND2_4190 ( P2_U3609 , P2_U6255 , P2_U6254 );
nand NAND2_4191 ( P2_U3610 , P2_U6257 , P2_U6256 );
nand NAND2_4192 ( P2_U3611 , P2_U6259 , P2_U6258 );
nand NAND2_4193 ( P2_U3612 , P2_U6261 , P2_U6260 );
nand NAND2_4194 ( P2_U3613 , P2_U6263 , P2_U6262 );
nand NAND2_4195 ( P2_U3614 , P2_U6265 , P2_U6264 );
nand NAND2_4196 ( P2_U3615 , P2_U6267 , P2_U6266 );
and AND2_4197 ( P2_U3616 , P2_U4134 , P2_U4133 );
and AND2_4198 ( P2_U3617 , P2_U4136 , P2_U4135 );
and AND2_4199 ( P2_U3618 , P2_U4143 , P2_U4141 );
and AND3_4200 ( P2_U3619 , P2_U4144 , P2_U4142 , P2_U3618 );
and AND4_4201 ( P2_U3620 , P2_U4100 , P2_U4099 , P2_U4098 , P2_U4097 );
and AND4_4202 ( P2_U3621 , P2_U4104 , P2_U4103 , P2_U4102 , P2_U4101 );
and AND4_4203 ( P2_U3622 , P2_U4108 , P2_U4107 , P2_U4106 , P2_U4105 );
and AND3_4204 ( P2_U3623 , P2_U4110 , P2_U4109 , P2_U4111 );
and AND4_4205 ( P2_U3624 , P2_U3623 , P2_U3622 , P2_U3621 , P2_U3620 );
and AND4_4206 ( P2_U3625 , P2_U4115 , P2_U4114 , P2_U4113 , P2_U4112 );
and AND4_4207 ( P2_U3626 , P2_U4119 , P2_U4118 , P2_U4117 , P2_U4116 );
and AND4_4208 ( P2_U3627 , P2_U4123 , P2_U4122 , P2_U4121 , P2_U4120 );
and AND3_4209 ( P2_U3628 , P2_U4125 , P2_U4124 , P2_U4126 );
and AND4_4210 ( P2_U3629 , P2_U3628 , P2_U3627 , P2_U3626 , P2_U3625 );
and AND2_4211 ( P2_U3630 , P2_U5741 , P2_U4127 );
and AND2_4212 ( P2_U3631 , P2_U5744 , P2_U3027 );
and AND2_4213 ( P2_U3632 , P2_U4155 , P2_U4154 );
and AND2_4214 ( P2_U3633 , P2_U4157 , P2_U4156 );
and AND3_4215 ( P2_U3634 , P2_U4159 , P2_U4158 , P2_U3633 );
and AND4_4216 ( P2_U3635 , P2_U4162 , P2_U4161 , P2_U4164 , P2_U4163 );
and AND2_4217 ( P2_U3636 , P2_U4174 , P2_U4173 );
and AND2_4218 ( P2_U3637 , P2_U4176 , P2_U4175 );
and AND3_4219 ( P2_U3638 , P2_U4178 , P2_U4177 , P2_U3637 );
and AND4_4220 ( P2_U3639 , P2_U4181 , P2_U4180 , P2_U4183 , P2_U4182 );
and AND2_4221 ( P2_U3640 , P2_U4193 , P2_U4192 );
and AND2_4222 ( P2_U3641 , P2_U4195 , P2_U4194 );
and AND3_4223 ( P2_U3642 , P2_U4197 , P2_U4196 , P2_U3641 );
and AND4_4224 ( P2_U3643 , P2_U4200 , P2_U4199 , P2_U4202 , P2_U4201 );
and AND2_4225 ( P2_U3644 , P2_U4212 , P2_U4211 );
and AND2_4226 ( P2_U3645 , P2_U4214 , P2_U4213 );
and AND3_4227 ( P2_U3646 , P2_U4216 , P2_U4215 , P2_U3645 );
and AND4_4228 ( P2_U3647 , P2_U4219 , P2_U4218 , P2_U4221 , P2_U4220 );
and AND2_4229 ( P2_U3648 , P2_U4231 , P2_U4230 );
and AND2_4230 ( P2_U3649 , P2_U4233 , P2_U4232 );
and AND3_4231 ( P2_U3650 , P2_U4235 , P2_U4234 , P2_U3649 );
and AND4_4232 ( P2_U3651 , P2_U4238 , P2_U4237 , P2_U4240 , P2_U4239 );
and AND2_4233 ( P2_U3652 , P2_U4250 , P2_U4249 );
and AND2_4234 ( P2_U3653 , P2_U4252 , P2_U4251 );
and AND3_4235 ( P2_U3654 , P2_U4254 , P2_U4253 , P2_U3653 );
and AND4_4236 ( P2_U3655 , P2_U4257 , P2_U4256 , P2_U4259 , P2_U4258 );
and AND2_4237 ( P2_U3656 , P2_U4269 , P2_U4268 );
and AND2_4238 ( P2_U3657 , P2_U4271 , P2_U4270 );
and AND3_4239 ( P2_U3658 , P2_U4273 , P2_U4272 , P2_U3657 );
and AND4_4240 ( P2_U3659 , P2_U4276 , P2_U4275 , P2_U4278 , P2_U4277 );
and AND2_4241 ( P2_U3660 , P2_U4288 , P2_U4287 );
and AND2_4242 ( P2_U3661 , P2_U4290 , P2_U4289 );
and AND3_4243 ( P2_U3662 , P2_U4292 , P2_U4291 , P2_U3661 );
and AND4_4244 ( P2_U3663 , P2_U4295 , P2_U4294 , P2_U4297 , P2_U4296 );
and AND2_4245 ( P2_U3664 , P2_U4307 , P2_U4306 );
and AND2_4246 ( P2_U3665 , P2_U4309 , P2_U4308 );
and AND3_4247 ( P2_U3666 , P2_U4311 , P2_U4310 , P2_U3665 );
and AND4_4248 ( P2_U3667 , P2_U4314 , P2_U4313 , P2_U4316 , P2_U4315 );
and AND2_4249 ( P2_U3668 , P2_U4326 , P2_U4325 );
and AND2_4250 ( P2_U3669 , P2_U4328 , P2_U4327 );
and AND3_4251 ( P2_U3670 , P2_U4330 , P2_U4329 , P2_U3669 );
and AND4_4252 ( P2_U3671 , P2_U4333 , P2_U4332 , P2_U4335 , P2_U4334 );
and AND2_4253 ( P2_U3672 , P2_U4345 , P2_U4344 );
and AND2_4254 ( P2_U3673 , P2_U4347 , P2_U4346 );
and AND3_4255 ( P2_U3674 , P2_U4349 , P2_U4348 , P2_U3673 );
and AND4_4256 ( P2_U3675 , P2_U4352 , P2_U4351 , P2_U4354 , P2_U4353 );
and AND2_4257 ( P2_U3676 , P2_U4364 , P2_U4363 );
and AND2_4258 ( P2_U3677 , P2_U4366 , P2_U4365 );
and AND3_4259 ( P2_U3678 , P2_U4368 , P2_U4367 , P2_U3677 );
and AND4_4260 ( P2_U3679 , P2_U4371 , P2_U4370 , P2_U4373 , P2_U4372 );
and AND2_4261 ( P2_U3680 , P2_U4383 , P2_U4382 );
and AND2_4262 ( P2_U3681 , P2_U4385 , P2_U4384 );
and AND3_4263 ( P2_U3682 , P2_U4387 , P2_U4386 , P2_U3681 );
and AND4_4264 ( P2_U3683 , P2_U4390 , P2_U4389 , P2_U4392 , P2_U4391 );
and AND2_4265 ( P2_U3684 , P2_U4402 , P2_U4401 );
and AND2_4266 ( P2_U3685 , P2_U4404 , P2_U4403 );
and AND3_4267 ( P2_U3686 , P2_U4406 , P2_U4405 , P2_U3685 );
and AND4_4268 ( P2_U3687 , P2_U4409 , P2_U4408 , P2_U4411 , P2_U4410 );
and AND2_4269 ( P2_U3688 , P2_U4421 , P2_U4420 );
and AND2_4270 ( P2_U3689 , P2_U4423 , P2_U4422 );
and AND3_4271 ( P2_U3690 , P2_U4425 , P2_U4424 , P2_U3689 );
and AND4_4272 ( P2_U3691 , P2_U4428 , P2_U4427 , P2_U4430 , P2_U4429 );
and AND2_4273 ( P2_U3692 , P2_U4440 , P2_U4439 );
and AND2_4274 ( P2_U3693 , P2_U4442 , P2_U4441 );
and AND3_4275 ( P2_U3694 , P2_U4444 , P2_U4443 , P2_U3693 );
and AND4_4276 ( P2_U3695 , P2_U4447 , P2_U4446 , P2_U4449 , P2_U4448 );
and AND2_4277 ( P2_U3696 , P2_U4459 , P2_U4458 );
and AND2_4278 ( P2_U3697 , P2_U4461 , P2_U4460 );
and AND3_4279 ( P2_U3698 , P2_U4463 , P2_U4462 , P2_U3697 );
and AND4_4280 ( P2_U3699 , P2_U4466 , P2_U4465 , P2_U4468 , P2_U4467 );
and AND2_4281 ( P2_U3700 , P2_U4478 , P2_U4477 );
and AND2_4282 ( P2_U3701 , P2_U4480 , P2_U4479 );
and AND3_4283 ( P2_U3702 , P2_U4482 , P2_U4481 , P2_U3701 );
and AND4_4284 ( P2_U3703 , P2_U4485 , P2_U4484 , P2_U4487 , P2_U4486 );
and AND2_4285 ( P2_U3704 , P2_U4497 , P2_U4496 );
and AND2_4286 ( P2_U3705 , P2_U4499 , P2_U4498 );
and AND3_4287 ( P2_U3706 , P2_U4501 , P2_U4500 , P2_U3705 );
and AND4_4288 ( P2_U3707 , P2_U4504 , P2_U4503 , P2_U4506 , P2_U4505 );
and AND2_4289 ( P2_U3708 , P2_U4516 , P2_U4515 );
and AND2_4290 ( P2_U3709 , P2_U4518 , P2_U4517 );
and AND3_4291 ( P2_U3710 , P2_U4520 , P2_U4519 , P2_U3709 );
and AND4_4292 ( P2_U3711 , P2_U4523 , P2_U4522 , P2_U4525 , P2_U4524 );
and AND2_4293 ( P2_U3712 , P2_U4535 , P2_U4534 );
and AND2_4294 ( P2_U3713 , P2_U4537 , P2_U4536 );
and AND3_4295 ( P2_U3714 , P2_U4539 , P2_U4538 , P2_U3713 );
and AND4_4296 ( P2_U3715 , P2_U4542 , P2_U4541 , P2_U4544 , P2_U4543 );
and AND2_4297 ( P2_U3716 , P2_U4554 , P2_U4553 );
and AND2_4298 ( P2_U3717 , P2_U4556 , P2_U4555 );
and AND3_4299 ( P2_U3718 , P2_U4558 , P2_U4557 , P2_U3717 );
and AND4_4300 ( P2_U3719 , P2_U4561 , P2_U4560 , P2_U4563 , P2_U4562 );
and AND2_4301 ( P2_U3720 , P2_U4573 , P2_U4572 );
and AND2_4302 ( P2_U3721 , P2_U4575 , P2_U4574 );
and AND3_4303 ( P2_U3722 , P2_U4577 , P2_U4576 , P2_U3721 );
and AND4_4304 ( P2_U3723 , P2_U4580 , P2_U4579 , P2_U4582 , P2_U4581 );
and AND2_4305 ( P2_U3724 , P2_U4592 , P2_U4591 );
and AND2_4306 ( P2_U3725 , P2_U4594 , P2_U4593 );
and AND3_4307 ( P2_U3726 , P2_U4596 , P2_U4595 , P2_U3725 );
and AND4_4308 ( P2_U3727 , P2_U4599 , P2_U4598 , P2_U4601 , P2_U4600 );
and AND2_4309 ( P2_U3728 , P2_U4611 , P2_U4610 );
and AND2_4310 ( P2_U3729 , P2_U4613 , P2_U4612 );
and AND3_4311 ( P2_U3730 , P2_U4615 , P2_U4614 , P2_U3729 );
and AND4_4312 ( P2_U3731 , P2_U4618 , P2_U4617 , P2_U4620 , P2_U4619 );
and AND2_4313 ( P2_U3732 , P2_U4630 , P2_U4629 );
and AND2_4314 ( P2_U3733 , P2_U4632 , P2_U4631 );
and AND3_4315 ( P2_U3734 , P2_U4634 , P2_U4633 , P2_U3733 );
and AND4_4316 ( P2_U3735 , P2_U4637 , P2_U4636 , P2_U4639 , P2_U4638 );
and AND2_4317 ( P2_U3736 , P2_U4649 , P2_U4648 );
and AND2_4318 ( P2_U3737 , P2_U4651 , P2_U4650 );
and AND3_4319 ( P2_U3738 , P2_U4653 , P2_U4652 , P2_U3737 );
and AND4_4320 ( P2_U3739 , P2_U4656 , P2_U4655 , P2_U4658 , P2_U4657 );
and AND2_4321 ( P2_U3740 , P2_U4670 , P2_U4669 );
and AND3_4322 ( P2_U3741 , P2_U4672 , P2_U4671 , P2_U3740 );
and AND4_4323 ( P2_U3742 , P2_U4675 , P2_U4674 , P2_U4677 , P2_U4676 );
and AND2_4324 ( P2_U3743 , P2_U4684 , P2_U3982 );
and AND2_4325 ( P2_U3744 , P2_U4689 , P2_U4688 );
and AND2_4326 ( P2_U3745 , P2_U4691 , P2_U4690 );
and AND3_4327 ( P2_U3746 , P2_U4693 , P2_U4692 , P2_U3745 );
and AND3_4328 ( P2_U3747 , P2_U4697 , P2_U4695 , P2_U4696 );
and AND2_4329 ( P2_U3748 , P2_U3982 , P2_U4684 );
and AND2_4330 ( P2_U3749 , P2_U3027 , P2_U3449 );
and AND3_4331 ( P2_U3750 , P2_U5744 , P2_U3051 , P2_U3450 );
and AND3_4332 ( P2_U3751 , P2_U3445 , P2_U5714 , P2_U3440 );
and AND3_4333 ( P2_U3752 , P2_U4715 , P2_U4714 , P2_U4716 );
and AND3_4334 ( P2_U3753 , P2_U4718 , P2_U4717 , P2_U3912 );
and AND3_4335 ( P2_U3754 , P2_U4720 , P2_U4719 , P2_U4721 );
and AND3_4336 ( P2_U3755 , P2_U4723 , P2_U4722 , P2_U3913 );
and AND3_4337 ( P2_U3756 , P2_U4725 , P2_U4724 , P2_U4726 );
and AND3_4338 ( P2_U3757 , P2_U4728 , P2_U4727 , P2_U3914 );
and AND3_4339 ( P2_U3758 , P2_U4730 , P2_U4729 , P2_U4731 );
and AND3_4340 ( P2_U3759 , P2_U4733 , P2_U4732 , P2_U3915 );
and AND3_4341 ( P2_U3760 , P2_U4735 , P2_U4734 , P2_U4736 );
and AND3_4342 ( P2_U3761 , P2_U4738 , P2_U4737 , P2_U3916 );
and AND3_4343 ( P2_U3762 , P2_U4740 , P2_U4739 , P2_U4741 );
and AND2_4344 ( P2_U3763 , P2_U4743 , P2_U4742 );
and AND3_4345 ( P2_U3764 , P2_U4745 , P2_U4744 , P2_U4746 );
and AND2_4346 ( P2_U3765 , P2_U4748 , P2_U4747 );
and AND3_4347 ( P2_U3766 , P2_U4750 , P2_U4749 , P2_U4751 );
and AND2_4348 ( P2_U3767 , P2_U4753 , P2_U4752 );
and AND3_4349 ( P2_U3768 , P2_U4755 , P2_U4754 , P2_U4756 );
and AND2_4350 ( P2_U3769 , P2_U4758 , P2_U4757 );
and AND3_4351 ( P2_U3770 , P2_U4760 , P2_U4759 , P2_U4761 );
and AND2_4352 ( P2_U3771 , P2_U4763 , P2_U4762 );
and AND2_4353 ( P2_U3772 , P2_U4766 , P2_U4764 );
and AND2_4354 ( P2_U3773 , P2_U4768 , P2_U4767 );
and AND3_4355 ( P2_U3774 , P2_U4770 , P2_U4769 , P2_U4771 );
and AND2_4356 ( P2_U3775 , P2_U4773 , P2_U4772 );
and AND2_4357 ( P2_U3776 , P2_U4776 , P2_U4774 );
and AND2_4358 ( P2_U3777 , P2_U4778 , P2_U4777 );
and AND2_4359 ( P2_U3778 , P2_U4781 , P2_U4779 );
and AND2_4360 ( P2_U3779 , P2_U4783 , P2_U4782 );
and AND2_4361 ( P2_U3780 , P2_U4786 , P2_U4784 );
and AND2_4362 ( P2_U3781 , P2_U4788 , P2_U4787 );
and AND2_4363 ( P2_U3782 , P2_U4791 , P2_U4789 );
and AND2_4364 ( P2_U3783 , P2_U4793 , P2_U4792 );
and AND2_4365 ( P2_U3784 , P2_U4796 , P2_U4794 );
and AND2_4366 ( P2_U3785 , P2_U4798 , P2_U4797 );
and AND2_4367 ( P2_U3786 , P2_U4801 , P2_U4799 );
and AND2_4368 ( P2_U3787 , P2_U4803 , P2_U4802 );
and AND2_4369 ( P2_U3788 , P2_U4806 , P2_U4804 );
and AND2_4370 ( P2_U3789 , P2_U4808 , P2_U4807 );
and AND2_4371 ( P2_U3790 , P2_U4811 , P2_U4809 );
and AND2_4372 ( P2_U3791 , P2_U4813 , P2_U4812 );
and AND2_4373 ( P2_U3792 , P2_U4816 , P2_U4814 );
and AND2_4374 ( P2_U3793 , P2_U4818 , P2_U4817 );
and AND2_4375 ( P2_U3794 , P2_U4821 , P2_U4819 );
and AND2_4376 ( P2_U3795 , P2_U4823 , P2_U4822 );
and AND2_4377 ( P2_U3796 , P2_U4826 , P2_U4824 );
and AND2_4378 ( P2_U3797 , P2_U4828 , P2_U4827 );
and AND2_4379 ( P2_U3798 , P2_U4831 , P2_U4829 );
and AND2_4380 ( P2_U3799 , P2_U4833 , P2_U4832 );
and AND2_4381 ( P2_U3800 , P2_U4836 , P2_U4834 );
and AND2_4382 ( P2_U3801 , P2_U4838 , P2_U4837 );
and AND2_4383 ( P2_U3802 , P2_U4841 , P2_U4839 );
and AND2_4384 ( P2_U3803 , P2_U4843 , P2_U4842 );
and AND2_4385 ( P2_U3804 , P2_U4846 , P2_U4844 );
and AND2_4386 ( P2_U3805 , P2_U4848 , P2_U4847 );
and AND2_4387 ( P2_U3806 , P2_U4851 , P2_U4849 );
and AND2_4388 ( P2_U3807 , P2_U4853 , P2_U4852 );
and AND2_4389 ( P2_U3808 , P2_U4856 , P2_U4854 );
and AND2_4390 ( P2_U3809 , P2_U4858 , P2_U4857 );
and AND2_4391 ( P2_U3810 , P2_U5686 , P2_U3421 );
and AND2_4392 ( P2_U3811 , P2_U3436 , P2_STATE_REG );
and AND2_4393 ( P2_U3812 , P2_U4877 , P2_U4876 );
and AND2_4394 ( P2_U3813 , P2_U4879 , P2_U4878 );
and AND3_4395 ( P2_U3814 , P2_U4882 , P2_U4880 , P2_U4881 );
and AND2_4396 ( P2_U3815 , P2_U4892 , P2_U4891 );
and AND2_4397 ( P2_U3816 , P2_U4894 , P2_U4893 );
and AND3_4398 ( P2_U3817 , P2_U4897 , P2_U4895 , P2_U4896 );
and AND2_4399 ( P2_U3818 , P2_U4907 , P2_U4906 );
and AND2_4400 ( P2_U3819 , P2_U4909 , P2_U4908 );
and AND3_4401 ( P2_U3820 , P2_U4912 , P2_U4910 , P2_U4911 );
and AND2_4402 ( P2_U3821 , P2_U4922 , P2_U4921 );
and AND2_4403 ( P2_U3822 , P2_U4924 , P2_U4923 );
and AND3_4404 ( P2_U3823 , P2_U4927 , P2_U4925 , P2_U4926 );
and AND2_4405 ( P2_U3824 , P2_U4937 , P2_U4936 );
and AND2_4406 ( P2_U3825 , P2_U4939 , P2_U4938 );
and AND3_4407 ( P2_U3826 , P2_U4942 , P2_U4940 , P2_U4941 );
and AND2_4408 ( P2_U3827 , P2_U4952 , P2_U4951 );
and AND2_4409 ( P2_U3828 , P2_U4954 , P2_U4953 );
and AND3_4410 ( P2_U3829 , P2_U4957 , P2_U4955 , P2_U4956 );
and AND2_4411 ( P2_U3830 , P2_U4967 , P2_U4966 );
and AND2_4412 ( P2_U3831 , P2_U4969 , P2_U4968 );
and AND3_4413 ( P2_U3832 , P2_U4972 , P2_U4970 , P2_U4971 );
and AND2_4414 ( P2_U3833 , P2_U4982 , P2_U4981 );
and AND2_4415 ( P2_U3834 , P2_U4984 , P2_U4983 );
and AND3_4416 ( P2_U3835 , P2_U4987 , P2_U4985 , P2_U4986 );
and AND2_4417 ( P2_U3836 , P2_U4997 , P2_U4996 );
and AND2_4418 ( P2_U3837 , P2_U4999 , P2_U4998 );
and AND3_4419 ( P2_U3838 , P2_U5002 , P2_U5000 , P2_U5001 );
and AND2_4420 ( P2_U3839 , P2_U5012 , P2_U5011 );
and AND2_4421 ( P2_U3840 , P2_U5014 , P2_U5013 );
and AND3_4422 ( P2_U3841 , P2_U5017 , P2_U5015 , P2_U5016 );
and AND2_4423 ( P2_U3842 , P2_U5027 , P2_U5026 );
and AND2_4424 ( P2_U3843 , P2_U5029 , P2_U5028 );
and AND3_4425 ( P2_U3844 , P2_U5032 , P2_U5030 , P2_U5031 );
and AND2_4426 ( P2_U3845 , P2_U5042 , P2_U5041 );
and AND3_4427 ( P2_U3846 , P2_U5044 , P2_U5043 , P2_U3845 );
and AND3_4428 ( P2_U3847 , P2_U5046 , P2_U5045 , P2_U5047 );
and AND2_4429 ( P2_U3848 , P2_U5057 , P2_U5056 );
and AND3_4430 ( P2_U3849 , P2_U5059 , P2_U5058 , P2_U3848 );
and AND3_4431 ( P2_U3850 , P2_U5061 , P2_U5060 , P2_U5062 );
and AND2_4432 ( P2_U3851 , P2_U5072 , P2_U5071 );
and AND3_4433 ( P2_U3852 , P2_U5074 , P2_U5073 , P2_U3851 );
and AND3_4434 ( P2_U3853 , P2_U5076 , P2_U5075 , P2_U5077 );
and AND2_4435 ( P2_U3854 , P2_U5087 , P2_U5086 );
and AND3_4436 ( P2_U3855 , P2_U5089 , P2_U5088 , P2_U3854 );
and AND3_4437 ( P2_U3856 , P2_U5091 , P2_U5090 , P2_U5092 );
and AND2_4438 ( P2_U3857 , P2_U5102 , P2_U5101 );
and AND3_4439 ( P2_U3858 , P2_U5104 , P2_U5103 , P2_U3857 );
and AND3_4440 ( P2_U3859 , P2_U5106 , P2_U5105 , P2_U5107 );
and AND2_4441 ( P2_U3860 , P2_U5117 , P2_U5116 );
and AND3_4442 ( P2_U3861 , P2_U5119 , P2_U5118 , P2_U3860 );
and AND3_4443 ( P2_U3862 , P2_U5121 , P2_U5120 , P2_U5122 );
and AND2_4444 ( P2_U3863 , P2_U5132 , P2_U5131 );
and AND3_4445 ( P2_U3864 , P2_U5134 , P2_U5133 , P2_U3863 );
and AND3_4446 ( P2_U3865 , P2_U5136 , P2_U5135 , P2_U5137 );
and AND2_4447 ( P2_U3866 , P2_U5147 , P2_U5146 );
and AND3_4448 ( P2_U3867 , P2_U5149 , P2_U5148 , P2_U3866 );
and AND3_4449 ( P2_U3868 , P2_U5151 , P2_U5150 , P2_U5152 );
and AND2_4450 ( P2_U3869 , P2_U5154 , P2_U5155 );
and AND2_4451 ( P2_U3870 , P2_U5162 , P2_U5161 );
and AND3_4452 ( P2_U3871 , P2_U5164 , P2_U5163 , P2_U3870 );
and AND3_4453 ( P2_U3872 , P2_U5166 , P2_U5165 , P2_U5167 );
and AND3_4454 ( P2_U3873 , P2_U6157 , P2_U6154 , P2_U6160 );
and AND2_4455 ( P2_U3874 , P2_U3873 , P2_U3875 );
and AND4_4456 ( P2_U3875 , P2_U6151 , P2_U6148 , P2_U6145 , P2_U6142 );
and AND3_4457 ( P2_U3876 , P2_U6169 , P2_U6166 , P2_U6172 );
and AND3_4458 ( P2_U3877 , P2_U6178 , P2_U6175 , P2_U6181 );
and AND3_4459 ( P2_U3878 , P2_U3877 , P2_U3876 , P2_U6163 );
and AND5_4460 ( P2_U3879 , P2_U3884 , P2_U3883 , P2_U6112 , P2_U6109 , P2_U6106 );
and AND5_4461 ( P2_U3880 , P2_U6196 , P2_U6193 , P2_U6190 , P2_U6187 , P2_U6199 );
and AND5_4462 ( P2_U3881 , P2_U3878 , P2_U3874 , P2_U6139 , P2_U6184 , P2_U3880 );
and AND2_4463 ( P2_U3882 , P2_U6133 , P2_U3879 );
and AND4_4464 ( P2_U3883 , P2_U6124 , P2_U6121 , P2_U6118 , P2_U6115 );
and AND2_4465 ( P2_U3884 , P2_U6130 , P2_U6127 );
and AND3_4466 ( P2_U3885 , P2_U5173 , P2_U5177 , P2_U5172 );
and AND2_4467 ( P2_U3886 , P2_U5670 , P2_U5176 );
and AND2_4468 ( P2_U3887 , P2_U3449 , P2_U3450 );
and AND2_4469 ( P2_U3888 , P2_U3432 , P2_U3952 );
and AND3_4470 ( P2_U3889 , P2_U5701 , P2_U3051 , P2_U3422 );
and AND2_4471 ( P2_U3890 , P2_U3027 , P2_U5183 );
and AND2_4472 ( P2_U3891 , P2_U3892 , P2_U5226 );
and AND2_4473 ( P2_U3892 , P2_U5230 , P2_U5229 );
and AND2_4474 ( P2_U3893 , P2_U3988 , P2_U3078 );
and AND2_4475 ( P2_U3894 , P2_U5271 , P2_U5270 );
and AND2_4476 ( P2_U3895 , P2_U5274 , P2_U5273 );
and AND2_4477 ( P2_U3896 , P2_U5292 , P2_U5291 );
and AND2_4478 ( P2_U3897 , P2_U5319 , P2_U5318 );
and AND2_4479 ( P2_U3898 , P2_U3899 , P2_U5360 );
and AND2_4480 ( P2_U3899 , P2_U5364 , P2_U5363 );
and AND2_4481 ( P2_U3900 , P2_U5391 , P2_U5387 );
and AND2_4482 ( P2_U3901 , P2_U3902 , P2_U5396 );
and AND2_4483 ( P2_U3902 , P2_U5400 , P2_U5399 );
and AND2_4484 ( P2_U3903 , P2_U5447 , P2_STATE_REG );
and AND2_4485 ( P2_U3904 , P2_U5717 , P2_U3415 );
and AND2_4486 ( P2_U3905 , P2_U5711 , P2_U5701 );
and AND2_4487 ( P2_U3906 , P2_U3440 , P2_U5512 );
not NOT1_4488 ( P2_U3907 , P2_IR_REG_31_ );
nand NAND2_4489 ( P2_U3908 , P2_U3027 , P2_U3362 );
nand NAND2_4490 ( P2_U3909 , P2_U5733 , P2_U5728 );
nand NAND2_4491 ( P2_U3910 , P2_U3631 , P2_U3049 );
nand NAND2_4492 ( P2_U3911 , P2_U3749 , P2_U3049 );
and AND2_4493 ( P2_U3912 , P2_U5971 , P2_U5970 );
and AND2_4494 ( P2_U3913 , P2_U5973 , P2_U5972 );
and AND2_4495 ( P2_U3914 , P2_U5975 , P2_U5974 );
and AND2_4496 ( P2_U3915 , P2_U5977 , P2_U5976 );
and AND2_4497 ( P2_U3916 , P2_U5979 , P2_U5978 );
and AND2_4498 ( P2_U3917 , P2_U5981 , P2_U5980 );
and AND2_4499 ( P2_U3918 , P2_U5983 , P2_U5982 );
and AND2_4500 ( P2_U3919 , P2_U5985 , P2_U5984 );
and AND2_4501 ( P2_U3920 , P2_U5987 , P2_U5986 );
and AND2_4502 ( P2_U3921 , P2_U5989 , P2_U5988 );
and AND2_4503 ( P2_U3922 , P2_U5991 , P2_U5990 );
and AND2_4504 ( P2_U3923 , P2_U5993 , P2_U5992 );
and AND2_4505 ( P2_U3924 , P2_U5995 , P2_U5994 );
and AND2_4506 ( P2_U3925 , P2_U5997 , P2_U5996 );
and AND2_4507 ( P2_U3926 , P2_U5999 , P2_U5998 );
and AND2_4508 ( P2_U3927 , P2_U6001 , P2_U6000 );
and AND2_4509 ( P2_U3928 , P2_U6003 , P2_U6002 );
and AND2_4510 ( P2_U3929 , P2_U6005 , P2_U6004 );
and AND2_4511 ( P2_U3930 , P2_U6007 , P2_U6006 );
and AND2_4512 ( P2_U3931 , P2_U6009 , P2_U6008 );
and AND2_4513 ( P2_U3932 , P2_U6011 , P2_U6010 );
and AND2_4514 ( P2_U3933 , P2_U6013 , P2_U6012 );
and AND2_4515 ( P2_U3934 , P2_U6015 , P2_U6014 );
and AND2_4516 ( P2_U3935 , P2_U6017 , P2_U6016 );
and AND2_4517 ( P2_U3936 , P2_U6019 , P2_U6018 );
and AND2_4518 ( P2_U3937 , P2_U6021 , P2_U6020 );
and AND2_4519 ( P2_U3938 , P2_U6023 , P2_U6022 );
and AND2_4520 ( P2_U3939 , P2_U6025 , P2_U6024 );
and AND2_4521 ( P2_U3940 , P2_U6027 , P2_U6026 );
and AND2_4522 ( P2_U3941 , P2_U6029 , P2_U6028 );
nand NAND2_4523 ( P2_U3942 , P2_U3748 , P2_U3056 );
and AND2_4524 ( P2_U3943 , P2_U6031 , P2_U6030 );
and AND2_4525 ( P2_U3944 , P2_U6033 , P2_U6032 );
not NOT1_4526 ( P2_U3945 , P2_R1312_U21 );
and AND2_4527 ( P2_U3946 , P2_U6103 , P2_U6102 );
nand NAND3_4528 ( P2_U3947 , P2_U3881 , P2_U6136 , P2_U3882 );
not NOT1_4529 ( P2_U3948 , P2_R1299_U6 );
not NOT1_4530 ( P2_U3949 , P2_U3370 );
nand NAND2_4531 ( P2_U3950 , P2_U3982 , P2_U3445 );
not NOT1_4532 ( P2_U3951 , P2_U3368 );
nand NAND2_4533 ( P2_U3952 , P2_U5674 , P2_U3441 );
not NOT1_4534 ( P2_U3953 , P2_U3432 );
not NOT1_4535 ( P2_U3954 , P2_U3369 );
not NOT1_4536 ( P2_U3955 , P2_U3363 );
not NOT1_4537 ( P2_U3956 , P2_U3419 );
not NOT1_4538 ( P2_U3957 , P2_U3418 );
nand NAND2_4539 ( P2_U3958 , P2_U3962 , P2_U5708 );
not NOT1_4540 ( P2_U3959 , P2_U3367 );
not NOT1_4541 ( P2_U3960 , P2_U3416 );
not NOT1_4542 ( P2_U3961 , P2_U3366 );
not NOT1_4543 ( P2_U3962 , P2_U3372 );
not NOT1_4544 ( P2_U3963 , P2_U3364 );
not NOT1_4545 ( P2_U3964 , P2_U3909 );
not NOT1_4546 ( P2_U3965 , P2_U3427 );
not NOT1_4547 ( P2_U3966 , P2_U3423 );
not NOT1_4548 ( P2_U3967 , P2_U3421 );
not NOT1_4549 ( P2_U3968 , P2_U3409 );
not NOT1_4550 ( P2_U3969 , P2_U3407 );
not NOT1_4551 ( P2_U3970 , P2_U3405 );
not NOT1_4552 ( P2_U3971 , P2_U3403 );
not NOT1_4553 ( P2_U3972 , P2_U3401 );
not NOT1_4554 ( P2_U3973 , P2_U3399 );
not NOT1_4555 ( P2_U3974 , P2_U3397 );
not NOT1_4556 ( P2_U3975 , P2_U3395 );
not NOT1_4557 ( P2_U3976 , P2_U3393 );
not NOT1_4558 ( P2_U3977 , P2_U3414 );
not NOT1_4559 ( P2_U3978 , P2_U3413 );
not NOT1_4560 ( P2_U3979 , P2_U3411 );
not NOT1_4561 ( P2_U3980 , P2_U3425 );
not NOT1_4562 ( P2_U3981 , P2_U3420 );
not NOT1_4563 ( P2_U3982 , P2_U3371 );
not NOT1_4564 ( P2_U3983 , P2_U3417 );
not NOT1_4565 ( P2_U3984 , P2_U3911 );
not NOT1_4566 ( P2_U3985 , P2_U3910 );
not NOT1_4567 ( P2_U3986 , P2_U3908 );
not NOT1_4568 ( P2_U3987 , P2_U3942 );
not NOT1_4569 ( P2_U3988 , P2_U3429 );
nand NAND2_4570 ( P2_U3989 , P2_U3430 , P2_STATE_REG );
nand NAND2_4571 ( P2_U3990 , P2_U3957 , P2_U3027 );
not NOT1_4572 ( P2_U3991 , P2_U3426 );
not NOT1_4573 ( P2_U3992 , P2_U3361 );
not NOT1_4574 ( P2_U3993 , P2_U3428 );
not NOT1_4575 ( P2_U3994 , P2_U3365 );
not NOT1_4576 ( P2_U3995 , P2_U3422 );
not NOT1_4577 ( P2_U3996 , P2_U3359 );
nand NAND2_4578 ( P2_U3997 , U56 , P2_U3152 );
nand NAND2_4579 ( P2_U3998 , P2_IR_REG_0_ , P2_U3033 );
nand NAND2_4580 ( P2_U3999 , P2_IR_REG_0_ , P2_U3996 );
nand NAND2_4581 ( P2_U4000 , U45 , P2_U3152 );
nand NAND2_4582 ( P2_U4001 , P2_SUB_598_U49 , P2_U3033 );
nand NAND2_4583 ( P2_U4002 , P2_IR_REG_1_ , P2_U3996 );
nand NAND2_4584 ( P2_U4003 , U34 , P2_U3152 );
nand NAND2_4585 ( P2_U4004 , P2_SUB_598_U24 , P2_U3033 );
nand NAND2_4586 ( P2_U4005 , P2_IR_REG_2_ , P2_U3996 );
nand NAND2_4587 ( P2_U4006 , U31 , P2_U3152 );
nand NAND2_4588 ( P2_U4007 , P2_SUB_598_U25 , P2_U3033 );
nand NAND2_4589 ( P2_U4008 , P2_IR_REG_3_ , P2_U3996 );
nand NAND2_4590 ( P2_U4009 , U30 , P2_U3152 );
nand NAND2_4591 ( P2_U4010 , P2_SUB_598_U26 , P2_U3033 );
nand NAND2_4592 ( P2_U4011 , P2_IR_REG_4_ , P2_U3996 );
nand NAND2_4593 ( P2_U4012 , U29 , P2_U3152 );
nand NAND2_4594 ( P2_U4013 , P2_SUB_598_U74 , P2_U3033 );
nand NAND2_4595 ( P2_U4014 , P2_IR_REG_5_ , P2_U3996 );
nand NAND2_4596 ( P2_U4015 , U28 , P2_U3152 );
nand NAND2_4597 ( P2_U4016 , P2_SUB_598_U27 , P2_U3033 );
nand NAND2_4598 ( P2_U4017 , P2_IR_REG_6_ , P2_U3996 );
nand NAND2_4599 ( P2_U4018 , U27 , P2_U3152 );
nand NAND2_4600 ( P2_U4019 , P2_SUB_598_U28 , P2_U3033 );
nand NAND2_4601 ( P2_U4020 , P2_IR_REG_7_ , P2_U3996 );
nand NAND2_4602 ( P2_U4021 , U26 , P2_U3152 );
nand NAND2_4603 ( P2_U4022 , P2_SUB_598_U29 , P2_U3033 );
nand NAND2_4604 ( P2_U4023 , P2_IR_REG_8_ , P2_U3996 );
nand NAND2_4605 ( P2_U4024 , U25 , P2_U3152 );
nand NAND2_4606 ( P2_U4025 , P2_SUB_598_U72 , P2_U3033 );
nand NAND2_4607 ( P2_U4026 , P2_IR_REG_9_ , P2_U3996 );
nand NAND2_4608 ( P2_U4027 , U55 , P2_U3152 );
nand NAND2_4609 ( P2_U4028 , P2_SUB_598_U11 , P2_U3033 );
nand NAND2_4610 ( P2_U4029 , P2_IR_REG_10_ , P2_U3996 );
nand NAND2_4611 ( P2_U4030 , U54 , P2_U3152 );
nand NAND2_4612 ( P2_U4031 , P2_SUB_598_U12 , P2_U3033 );
nand NAND2_4613 ( P2_U4032 , P2_IR_REG_11_ , P2_U3996 );
nand NAND2_4614 ( P2_U4033 , U53 , P2_U3152 );
nand NAND2_4615 ( P2_U4034 , P2_SUB_598_U13 , P2_U3033 );
nand NAND2_4616 ( P2_U4035 , P2_IR_REG_12_ , P2_U3996 );
nand NAND2_4617 ( P2_U4036 , U52 , P2_U3152 );
nand NAND2_4618 ( P2_U4037 , P2_SUB_598_U99 , P2_U3033 );
nand NAND2_4619 ( P2_U4038 , P2_IR_REG_13_ , P2_U3996 );
nand NAND2_4620 ( P2_U4039 , U51 , P2_U3152 );
nand NAND2_4621 ( P2_U4040 , P2_SUB_598_U14 , P2_U3033 );
nand NAND2_4622 ( P2_U4041 , P2_IR_REG_14_ , P2_U3996 );
nand NAND2_4623 ( P2_U4042 , U50 , P2_U3152 );
nand NAND2_4624 ( P2_U4043 , P2_SUB_598_U15 , P2_U3033 );
nand NAND2_4625 ( P2_U4044 , P2_IR_REG_15_ , P2_U3996 );
nand NAND2_4626 ( P2_U4045 , U49 , P2_U3152 );
nand NAND2_4627 ( P2_U4046 , P2_SUB_598_U16 , P2_U3033 );
nand NAND2_4628 ( P2_U4047 , P2_IR_REG_16_ , P2_U3996 );
nand NAND2_4629 ( P2_U4048 , U48 , P2_U3152 );
nand NAND2_4630 ( P2_U4049 , P2_SUB_598_U97 , P2_U3033 );
nand NAND2_4631 ( P2_U4050 , P2_IR_REG_17_ , P2_U3996 );
nand NAND2_4632 ( P2_U4051 , U47 , P2_U3152 );
nand NAND2_4633 ( P2_U4052 , P2_SUB_598_U17 , P2_U3033 );
nand NAND2_4634 ( P2_U4053 , P2_IR_REG_18_ , P2_U3996 );
nand NAND2_4635 ( P2_U4054 , U46 , P2_U3152 );
nand NAND2_4636 ( P2_U4055 , P2_SUB_598_U18 , P2_U3033 );
nand NAND2_4637 ( P2_U4056 , P2_IR_REG_19_ , P2_U3996 );
nand NAND2_4638 ( P2_U4057 , U44 , P2_U3152 );
nand NAND2_4639 ( P2_U4058 , P2_SUB_598_U19 , P2_U3033 );
nand NAND2_4640 ( P2_U4059 , P2_IR_REG_20_ , P2_U3996 );
nand NAND2_4641 ( P2_U4060 , U43 , P2_U3152 );
nand NAND2_4642 ( P2_U4061 , P2_SUB_598_U92 , P2_U3033 );
nand NAND2_4643 ( P2_U4062 , P2_IR_REG_21_ , P2_U3996 );
nand NAND2_4644 ( P2_U4063 , U42 , P2_U3152 );
nand NAND2_4645 ( P2_U4064 , P2_SUB_598_U20 , P2_U3033 );
nand NAND2_4646 ( P2_U4065 , P2_IR_REG_22_ , P2_U3996 );
nand NAND2_4647 ( P2_U4066 , U41 , P2_U3152 );
nand NAND2_4648 ( P2_U4067 , P2_SUB_598_U21 , P2_U3033 );
nand NAND2_4649 ( P2_U4068 , P2_IR_REG_23_ , P2_U3996 );
nand NAND2_4650 ( P2_U4069 , U40 , P2_U3152 );
nand NAND2_4651 ( P2_U4070 , P2_SUB_598_U90 , P2_U3033 );
nand NAND2_4652 ( P2_U4071 , P2_IR_REG_24_ , P2_U3996 );
nand NAND2_4653 ( P2_U4072 , U39 , P2_U3152 );
nand NAND2_4654 ( P2_U4073 , P2_SUB_598_U22 , P2_U3033 );
nand NAND2_4655 ( P2_U4074 , P2_IR_REG_25_ , P2_U3996 );
nand NAND2_4656 ( P2_U4075 , U38 , P2_U3152 );
nand NAND2_4657 ( P2_U4076 , P2_SUB_598_U23 , P2_U3033 );
nand NAND2_4658 ( P2_U4077 , P2_IR_REG_26_ , P2_U3996 );
nand NAND2_4659 ( P2_U4078 , U37 , P2_U3152 );
nand NAND2_4660 ( P2_U4079 , P2_SUB_598_U87 , P2_U3033 );
nand NAND2_4661 ( P2_U4080 , P2_IR_REG_27_ , P2_U3996 );
nand NAND2_4662 ( P2_U4081 , U36 , P2_U3152 );
nand NAND2_4663 ( P2_U4082 , P2_SUB_598_U84 , P2_U3033 );
nand NAND2_4664 ( P2_U4083 , P2_IR_REG_28_ , P2_U3996 );
nand NAND2_4665 ( P2_U4084 , U35 , P2_U3152 );
nand NAND2_4666 ( P2_U4085 , P2_SUB_598_U81 , P2_U3033 );
nand NAND2_4667 ( P2_U4086 , P2_IR_REG_29_ , P2_U3996 );
nand NAND2_4668 ( P2_U4087 , U33 , P2_U3152 );
nand NAND2_4669 ( P2_U4088 , P2_SUB_598_U79 , P2_U3033 );
nand NAND2_4670 ( P2_U4089 , P2_IR_REG_30_ , P2_U3996 );
nand NAND2_4671 ( P2_U4090 , U32 , P2_U3152 );
nand NAND2_4672 ( P2_U4091 , P2_SUB_598_U77 , P2_U3033 );
nand NAND2_4673 ( P2_U4092 , P2_IR_REG_31_ , P2_U3996 );
nand NAND2_4674 ( P2_U4093 , P2_U3992 , P2_U5698 );
not NOT1_4675 ( P2_U4094 , P2_U3362 );
nand NAND2_4676 ( P2_U4095 , P2_U3361 , P2_U5689 );
nand NAND2_4677 ( P2_U4096 , P2_U3361 , P2_U5692 );
nand NAND2_4678 ( P2_U4097 , P2_U4094 , P2_D_REG_10_ );
nand NAND2_4679 ( P2_U4098 , P2_U4094 , P2_D_REG_11_ );
nand NAND2_4680 ( P2_U4099 , P2_U4094 , P2_D_REG_12_ );
nand NAND2_4681 ( P2_U4100 , P2_U4094 , P2_D_REG_13_ );
nand NAND2_4682 ( P2_U4101 , P2_U4094 , P2_D_REG_14_ );
nand NAND2_4683 ( P2_U4102 , P2_U4094 , P2_D_REG_15_ );
nand NAND2_4684 ( P2_U4103 , P2_U4094 , P2_D_REG_16_ );
nand NAND2_4685 ( P2_U4104 , P2_U4094 , P2_D_REG_17_ );
nand NAND2_4686 ( P2_U4105 , P2_U4094 , P2_D_REG_18_ );
nand NAND2_4687 ( P2_U4106 , P2_U4094 , P2_D_REG_19_ );
nand NAND2_4688 ( P2_U4107 , P2_U4094 , P2_D_REG_20_ );
nand NAND2_4689 ( P2_U4108 , P2_U4094 , P2_D_REG_21_ );
nand NAND2_4690 ( P2_U4109 , P2_U4094 , P2_D_REG_22_ );
nand NAND2_4691 ( P2_U4110 , P2_U4094 , P2_D_REG_23_ );
nand NAND2_4692 ( P2_U4111 , P2_U4094 , P2_D_REG_24_ );
nand NAND2_4693 ( P2_U4112 , P2_U4094 , P2_D_REG_25_ );
nand NAND2_4694 ( P2_U4113 , P2_U4094 , P2_D_REG_26_ );
nand NAND2_4695 ( P2_U4114 , P2_U4094 , P2_D_REG_27_ );
nand NAND2_4696 ( P2_U4115 , P2_U4094 , P2_D_REG_28_ );
nand NAND2_4697 ( P2_U4116 , P2_U4094 , P2_D_REG_29_ );
nand NAND2_4698 ( P2_U4117 , P2_U4094 , P2_D_REG_2_ );
nand NAND2_4699 ( P2_U4118 , P2_U4094 , P2_D_REG_30_ );
nand NAND2_4700 ( P2_U4119 , P2_U4094 , P2_D_REG_31_ );
nand NAND2_4701 ( P2_U4120 , P2_U4094 , P2_D_REG_3_ );
nand NAND2_4702 ( P2_U4121 , P2_U4094 , P2_D_REG_4_ );
nand NAND2_4703 ( P2_U4122 , P2_U4094 , P2_D_REG_5_ );
nand NAND2_4704 ( P2_U4123 , P2_U4094 , P2_D_REG_6_ );
nand NAND2_4705 ( P2_U4124 , P2_U4094 , P2_D_REG_7_ );
nand NAND2_4706 ( P2_U4125 , P2_U4094 , P2_D_REG_8_ );
nand NAND2_4707 ( P2_U4126 , P2_U4094 , P2_D_REG_9_ );
nand NAND4_4708 ( P2_U4127 , P2_U3365 , P2_U3428 , P2_U5738 , P2_U5737 );
nand NAND2_4709 ( P2_U4128 , P2_U3025 , P2_REG1_REG_1_ );
nand NAND2_4710 ( P2_U4129 , P2_U3026 , P2_REG0_REG_1_ );
not NOT1_4711 ( P2_U4130 , P2_U3078 );
nand NAND2_4712 ( P2_U4131 , P2_U3949 , P2_U3445 );
nand NAND2_4713 ( P2_U4132 , P2_U3958 , P2_U4131 );
nand NAND2_4714 ( P2_U4133 , P2_U3955 , P2_R1146_U19 );
nand NAND2_4715 ( P2_U4134 , P2_U3015 , P2_R1113_U19 );
nand NAND2_4716 ( P2_U4135 , P2_U3014 , P2_R1131_U95 );
nand NAND2_4717 ( P2_U4136 , P2_U3018 , P2_R1179_U19 );
nand NAND2_4718 ( P2_U4137 , P2_U3963 , P2_R1203_U19 );
nand NAND2_4719 ( P2_U4138 , P2_U3959 , P2_R1164_U95 );
nand NAND2_4720 ( P2_U4139 , P2_U3016 , P2_R1233_U95 );
not NOT1_4721 ( P2_U4140 , P2_U3373 );
nand NAND2_4722 ( P2_U4141 , P2_U3448 , P2_U3031 );
nand NAND2_4723 ( P2_U4142 , P2_U3030 , P2_U3078 );
nand NAND2_4724 ( P2_U4143 , P2_R1215_U95 , P2_U3028 );
nand NAND2_4725 ( P2_U4144 , P2_U3448 , P2_U4132 );
nand NAND2_4726 ( P2_U4145 , P2_U3619 , P2_U4140 );
nand NAND2_4727 ( P2_U4146 , P2_REG1_REG_2_ , P2_U3025 );
nand NAND2_4728 ( P2_U4147 , P2_REG0_REG_2_ , P2_U3026 );
not NOT1_4729 ( P2_U4148 , P2_U3068 );
nand NAND2_4730 ( P2_U4149 , P2_REG1_REG_0_ , P2_U3025 );
nand NAND2_4731 ( P2_U4150 , P2_REG0_REG_0_ , P2_U3026 );
not NOT1_4732 ( P2_U4151 , P2_U3077 );
nand NAND2_4733 ( P2_U4152 , P2_U3038 , P2_U3077 );
nand NAND2_4734 ( P2_U4153 , P2_R1146_U94 , P2_U3955 );
nand NAND2_4735 ( P2_U4154 , P2_R1113_U94 , P2_U3015 );
nand NAND2_4736 ( P2_U4155 , P2_R1131_U94 , P2_U3014 );
nand NAND2_4737 ( P2_U4156 , P2_R1179_U94 , P2_U3018 );
nand NAND2_4738 ( P2_U4157 , P2_R1203_U94 , P2_U3963 );
nand NAND2_4739 ( P2_U4158 , P2_R1164_U94 , P2_U3959 );
nand NAND2_4740 ( P2_U4159 , P2_R1233_U94 , P2_U3016 );
not NOT1_4741 ( P2_U4160 , P2_U3374 );
nand NAND2_4742 ( P2_U4161 , P2_R1275_U55 , P2_U3031 );
nand NAND2_4743 ( P2_U4162 , P2_U3030 , P2_U3068 );
nand NAND2_4744 ( P2_U4163 , P2_R1215_U94 , P2_U3028 );
nand NAND2_4745 ( P2_U4164 , P2_U3453 , P2_U4132 );
nand NAND2_4746 ( P2_U4165 , P2_U3635 , P2_U4160 );
nand NAND2_4747 ( P2_U4166 , P2_U3024 , P2_REG2_REG_3_ );
nand NAND2_4748 ( P2_U4167 , P2_REG1_REG_3_ , P2_U3025 );
nand NAND2_4749 ( P2_U4168 , P2_REG0_REG_3_ , P2_U3026 );
nand NAND2_4750 ( P2_U4169 , P2_ADD_609_U4 , P2_U3023 );
not NOT1_4751 ( P2_U4170 , P2_U3064 );
nand NAND2_4752 ( P2_U4171 , P2_U3038 , P2_U3078 );
nand NAND2_4753 ( P2_U4172 , P2_R1146_U104 , P2_U3955 );
nand NAND2_4754 ( P2_U4173 , P2_R1113_U104 , P2_U3015 );
nand NAND2_4755 ( P2_U4174 , P2_R1131_U16 , P2_U3014 );
nand NAND2_4756 ( P2_U4175 , P2_R1179_U104 , P2_U3018 );
nand NAND2_4757 ( P2_U4176 , P2_R1203_U104 , P2_U3963 );
nand NAND2_4758 ( P2_U4177 , P2_R1164_U16 , P2_U3959 );
nand NAND2_4759 ( P2_U4178 , P2_R1233_U16 , P2_U3016 );
not NOT1_4760 ( P2_U4179 , P2_U3375 );
nand NAND2_4761 ( P2_U4180 , P2_R1275_U18 , P2_U3031 );
nand NAND2_4762 ( P2_U4181 , P2_U3030 , P2_U3064 );
nand NAND2_4763 ( P2_U4182 , P2_R1215_U16 , P2_U3028 );
nand NAND2_4764 ( P2_U4183 , P2_U3456 , P2_U4132 );
nand NAND2_4765 ( P2_U4184 , P2_U3639 , P2_U4179 );
nand NAND2_4766 ( P2_U4185 , P2_REG2_REG_4_ , P2_U3024 );
nand NAND2_4767 ( P2_U4186 , P2_REG1_REG_4_ , P2_U3025 );
nand NAND2_4768 ( P2_U4187 , P2_REG0_REG_4_ , P2_U3026 );
nand NAND2_4769 ( P2_U4188 , P2_ADD_609_U54 , P2_U3023 );
not NOT1_4770 ( P2_U4189 , P2_U3060 );
nand NAND2_4771 ( P2_U4190 , P2_U3038 , P2_U3068 );
nand NAND2_4772 ( P2_U4191 , P2_R1146_U16 , P2_U3955 );
nand NAND2_4773 ( P2_U4192 , P2_R1113_U16 , P2_U3015 );
nand NAND2_4774 ( P2_U4193 , P2_R1131_U100 , P2_U3014 );
nand NAND2_4775 ( P2_U4194 , P2_R1179_U16 , P2_U3018 );
nand NAND2_4776 ( P2_U4195 , P2_R1203_U16 , P2_U3963 );
nand NAND2_4777 ( P2_U4196 , P2_R1164_U100 , P2_U3959 );
nand NAND2_4778 ( P2_U4197 , P2_R1233_U100 , P2_U3016 );
not NOT1_4779 ( P2_U4198 , P2_U3376 );
nand NAND2_4780 ( P2_U4199 , P2_R1275_U20 , P2_U3031 );
nand NAND2_4781 ( P2_U4200 , P2_U3030 , P2_U3060 );
nand NAND2_4782 ( P2_U4201 , P2_R1215_U100 , P2_U3028 );
nand NAND2_4783 ( P2_U4202 , P2_U3459 , P2_U4132 );
nand NAND2_4784 ( P2_U4203 , P2_U3643 , P2_U4198 );
nand NAND2_4785 ( P2_U4204 , P2_REG2_REG_5_ , P2_U3024 );
nand NAND2_4786 ( P2_U4205 , P2_REG1_REG_5_ , P2_U3025 );
nand NAND2_4787 ( P2_U4206 , P2_REG0_REG_5_ , P2_U3026 );
nand NAND2_4788 ( P2_U4207 , P2_ADD_609_U53 , P2_U3023 );
not NOT1_4789 ( P2_U4208 , P2_U3067 );
nand NAND2_4790 ( P2_U4209 , P2_U3038 , P2_U3064 );
nand NAND2_4791 ( P2_U4210 , P2_R1146_U103 , P2_U3955 );
nand NAND2_4792 ( P2_U4211 , P2_R1113_U103 , P2_U3015 );
nand NAND2_4793 ( P2_U4212 , P2_R1131_U99 , P2_U3014 );
nand NAND2_4794 ( P2_U4213 , P2_R1179_U103 , P2_U3018 );
nand NAND2_4795 ( P2_U4214 , P2_R1203_U103 , P2_U3963 );
nand NAND2_4796 ( P2_U4215 , P2_R1164_U99 , P2_U3959 );
nand NAND2_4797 ( P2_U4216 , P2_R1233_U99 , P2_U3016 );
not NOT1_4798 ( P2_U4217 , P2_U3377 );
nand NAND2_4799 ( P2_U4218 , P2_R1275_U21 , P2_U3031 );
nand NAND2_4800 ( P2_U4219 , P2_U3030 , P2_U3067 );
nand NAND2_4801 ( P2_U4220 , P2_R1215_U99 , P2_U3028 );
nand NAND2_4802 ( P2_U4221 , P2_U3462 , P2_U4132 );
nand NAND2_4803 ( P2_U4222 , P2_U3647 , P2_U4217 );
nand NAND2_4804 ( P2_U4223 , P2_REG2_REG_6_ , P2_U3024 );
nand NAND2_4805 ( P2_U4224 , P2_REG1_REG_6_ , P2_U3025 );
nand NAND2_4806 ( P2_U4225 , P2_REG0_REG_6_ , P2_U3026 );
nand NAND2_4807 ( P2_U4226 , P2_ADD_609_U52 , P2_U3023 );
not NOT1_4808 ( P2_U4227 , P2_U3071 );
nand NAND2_4809 ( P2_U4228 , P2_U3038 , P2_U3060 );
nand NAND2_4810 ( P2_U4229 , P2_R1146_U102 , P2_U3955 );
nand NAND2_4811 ( P2_U4230 , P2_R1113_U102 , P2_U3015 );
nand NAND2_4812 ( P2_U4231 , P2_R1131_U17 , P2_U3014 );
nand NAND2_4813 ( P2_U4232 , P2_R1179_U102 , P2_U3018 );
nand NAND2_4814 ( P2_U4233 , P2_R1203_U102 , P2_U3963 );
nand NAND2_4815 ( P2_U4234 , P2_R1164_U17 , P2_U3959 );
nand NAND2_4816 ( P2_U4235 , P2_R1233_U17 , P2_U3016 );
not NOT1_4817 ( P2_U4236 , P2_U3378 );
nand NAND2_4818 ( P2_U4237 , P2_R1275_U65 , P2_U3031 );
nand NAND2_4819 ( P2_U4238 , P2_U3030 , P2_U3071 );
nand NAND2_4820 ( P2_U4239 , P2_R1215_U17 , P2_U3028 );
nand NAND2_4821 ( P2_U4240 , P2_U3465 , P2_U4132 );
nand NAND2_4822 ( P2_U4241 , P2_U3651 , P2_U4236 );
nand NAND2_4823 ( P2_U4242 , P2_REG2_REG_7_ , P2_U3024 );
nand NAND2_4824 ( P2_U4243 , P2_REG1_REG_7_ , P2_U3025 );
nand NAND2_4825 ( P2_U4244 , P2_REG0_REG_7_ , P2_U3026 );
nand NAND2_4826 ( P2_U4245 , P2_ADD_609_U51 , P2_U3023 );
not NOT1_4827 ( P2_U4246 , P2_U3070 );
nand NAND2_4828 ( P2_U4247 , P2_U3038 , P2_U3067 );
nand NAND2_4829 ( P2_U4248 , P2_R1146_U17 , P2_U3955 );
nand NAND2_4830 ( P2_U4249 , P2_R1113_U17 , P2_U3015 );
nand NAND2_4831 ( P2_U4250 , P2_R1131_U98 , P2_U3014 );
nand NAND2_4832 ( P2_U4251 , P2_R1179_U17 , P2_U3018 );
nand NAND2_4833 ( P2_U4252 , P2_R1203_U17 , P2_U3963 );
nand NAND2_4834 ( P2_U4253 , P2_R1164_U98 , P2_U3959 );
nand NAND2_4835 ( P2_U4254 , P2_R1233_U98 , P2_U3016 );
not NOT1_4836 ( P2_U4255 , P2_U3379 );
nand NAND2_4837 ( P2_U4256 , P2_R1275_U22 , P2_U3031 );
nand NAND2_4838 ( P2_U4257 , P2_U3030 , P2_U3070 );
nand NAND2_4839 ( P2_U4258 , P2_R1215_U98 , P2_U3028 );
nand NAND2_4840 ( P2_U4259 , P2_U3468 , P2_U4132 );
nand NAND2_4841 ( P2_U4260 , P2_U3655 , P2_U4255 );
nand NAND2_4842 ( P2_U4261 , P2_REG2_REG_8_ , P2_U3024 );
nand NAND2_4843 ( P2_U4262 , P2_REG1_REG_8_ , P2_U3025 );
nand NAND2_4844 ( P2_U4263 , P2_REG0_REG_8_ , P2_U3026 );
nand NAND2_4845 ( P2_U4264 , P2_ADD_609_U50 , P2_U3023 );
not NOT1_4846 ( P2_U4265 , P2_U3084 );
nand NAND2_4847 ( P2_U4266 , P2_U3038 , P2_U3071 );
nand NAND2_4848 ( P2_U4267 , P2_R1146_U101 , P2_U3955 );
nand NAND2_4849 ( P2_U4268 , P2_R1113_U101 , P2_U3015 );
nand NAND2_4850 ( P2_U4269 , P2_R1131_U18 , P2_U3014 );
nand NAND2_4851 ( P2_U4270 , P2_R1179_U101 , P2_U3018 );
nand NAND2_4852 ( P2_U4271 , P2_R1203_U101 , P2_U3963 );
nand NAND2_4853 ( P2_U4272 , P2_R1164_U18 , P2_U3959 );
nand NAND2_4854 ( P2_U4273 , P2_R1233_U18 , P2_U3016 );
not NOT1_4855 ( P2_U4274 , P2_U3380 );
nand NAND2_4856 ( P2_U4275 , P2_R1275_U23 , P2_U3031 );
nand NAND2_4857 ( P2_U4276 , P2_U3030 , P2_U3084 );
nand NAND2_4858 ( P2_U4277 , P2_R1215_U18 , P2_U3028 );
nand NAND2_4859 ( P2_U4278 , P2_U3471 , P2_U4132 );
nand NAND2_4860 ( P2_U4279 , P2_U3659 , P2_U4274 );
nand NAND2_4861 ( P2_U4280 , P2_REG2_REG_9_ , P2_U3024 );
nand NAND2_4862 ( P2_U4281 , P2_REG1_REG_9_ , P2_U3025 );
nand NAND2_4863 ( P2_U4282 , P2_REG0_REG_9_ , P2_U3026 );
nand NAND2_4864 ( P2_U4283 , P2_ADD_609_U49 , P2_U3023 );
not NOT1_4865 ( P2_U4284 , P2_U3083 );
nand NAND2_4866 ( P2_U4285 , P2_U3038 , P2_U3070 );
nand NAND2_4867 ( P2_U4286 , P2_R1146_U18 , P2_U3955 );
nand NAND2_4868 ( P2_U4287 , P2_R1113_U18 , P2_U3015 );
nand NAND2_4869 ( P2_U4288 , P2_R1131_U97 , P2_U3014 );
nand NAND2_4870 ( P2_U4289 , P2_R1179_U18 , P2_U3018 );
nand NAND2_4871 ( P2_U4290 , P2_R1203_U18 , P2_U3963 );
nand NAND2_4872 ( P2_U4291 , P2_R1164_U97 , P2_U3959 );
nand NAND2_4873 ( P2_U4292 , P2_R1233_U97 , P2_U3016 );
not NOT1_4874 ( P2_U4293 , P2_U3381 );
nand NAND2_4875 ( P2_U4294 , P2_R1275_U24 , P2_U3031 );
nand NAND2_4876 ( P2_U4295 , P2_U3030 , P2_U3083 );
nand NAND2_4877 ( P2_U4296 , P2_R1215_U97 , P2_U3028 );
nand NAND2_4878 ( P2_U4297 , P2_U3474 , P2_U4132 );
nand NAND2_4879 ( P2_U4298 , P2_U3663 , P2_U4293 );
nand NAND2_4880 ( P2_U4299 , P2_REG2_REG_10_ , P2_U3024 );
nand NAND2_4881 ( P2_U4300 , P2_REG1_REG_10_ , P2_U3025 );
nand NAND2_4882 ( P2_U4301 , P2_REG0_REG_10_ , P2_U3026 );
nand NAND2_4883 ( P2_U4302 , P2_ADD_609_U73 , P2_U3023 );
not NOT1_4884 ( P2_U4303 , P2_U3062 );
nand NAND2_4885 ( P2_U4304 , P2_U3038 , P2_U3084 );
nand NAND2_4886 ( P2_U4305 , P2_R1146_U100 , P2_U3955 );
nand NAND2_4887 ( P2_U4306 , P2_R1113_U100 , P2_U3015 );
nand NAND2_4888 ( P2_U4307 , P2_R1131_U96 , P2_U3014 );
nand NAND2_4889 ( P2_U4308 , P2_R1179_U100 , P2_U3018 );
nand NAND2_4890 ( P2_U4309 , P2_R1203_U100 , P2_U3963 );
nand NAND2_4891 ( P2_U4310 , P2_R1164_U96 , P2_U3959 );
nand NAND2_4892 ( P2_U4311 , P2_R1233_U96 , P2_U3016 );
not NOT1_4893 ( P2_U4312 , P2_U3382 );
nand NAND2_4894 ( P2_U4313 , P2_R1275_U63 , P2_U3031 );
nand NAND2_4895 ( P2_U4314 , P2_U3030 , P2_U3062 );
nand NAND2_4896 ( P2_U4315 , P2_R1215_U96 , P2_U3028 );
nand NAND2_4897 ( P2_U4316 , P2_U3477 , P2_U4132 );
nand NAND2_4898 ( P2_U4317 , P2_U3667 , P2_U4312 );
nand NAND2_4899 ( P2_U4318 , P2_REG2_REG_11_ , P2_U3024 );
nand NAND2_4900 ( P2_U4319 , P2_REG1_REG_11_ , P2_U3025 );
nand NAND2_4901 ( P2_U4320 , P2_REG0_REG_11_ , P2_U3026 );
nand NAND2_4902 ( P2_U4321 , P2_ADD_609_U72 , P2_U3023 );
not NOT1_4903 ( P2_U4322 , P2_U3063 );
nand NAND2_4904 ( P2_U4323 , P2_U3038 , P2_U3083 );
nand NAND2_4905 ( P2_U4324 , P2_R1146_U110 , P2_U3955 );
nand NAND2_4906 ( P2_U4325 , P2_R1113_U110 , P2_U3015 );
nand NAND2_4907 ( P2_U4326 , P2_R1131_U10 , P2_U3014 );
nand NAND2_4908 ( P2_U4327 , P2_R1179_U110 , P2_U3018 );
nand NAND2_4909 ( P2_U4328 , P2_R1203_U110 , P2_U3963 );
nand NAND2_4910 ( P2_U4329 , P2_R1164_U10 , P2_U3959 );
nand NAND2_4911 ( P2_U4330 , P2_R1233_U10 , P2_U3016 );
not NOT1_4912 ( P2_U4331 , P2_U3383 );
nand NAND2_4913 ( P2_U4332 , P2_R1275_U6 , P2_U3031 );
nand NAND2_4914 ( P2_U4333 , P2_U3030 , P2_U3063 );
nand NAND2_4915 ( P2_U4334 , P2_R1215_U10 , P2_U3028 );
nand NAND2_4916 ( P2_U4335 , P2_U3480 , P2_U4132 );
nand NAND2_4917 ( P2_U4336 , P2_U3671 , P2_U4331 );
nand NAND2_4918 ( P2_U4337 , P2_REG2_REG_12_ , P2_U3024 );
nand NAND2_4919 ( P2_U4338 , P2_REG1_REG_12_ , P2_U3025 );
nand NAND2_4920 ( P2_U4339 , P2_REG0_REG_12_ , P2_U3026 );
nand NAND2_4921 ( P2_U4340 , P2_ADD_609_U71 , P2_U3023 );
not NOT1_4922 ( P2_U4341 , P2_U3072 );
nand NAND2_4923 ( P2_U4342 , P2_U3038 , P2_U3062 );
nand NAND2_4924 ( P2_U4343 , P2_R1146_U11 , P2_U3955 );
nand NAND2_4925 ( P2_U4344 , P2_R1113_U11 , P2_U3015 );
nand NAND2_4926 ( P2_U4345 , P2_R1131_U114 , P2_U3014 );
nand NAND2_4927 ( P2_U4346 , P2_R1179_U11 , P2_U3018 );
nand NAND2_4928 ( P2_U4347 , P2_R1203_U11 , P2_U3963 );
nand NAND2_4929 ( P2_U4348 , P2_R1164_U114 , P2_U3959 );
nand NAND2_4930 ( P2_U4349 , P2_R1233_U114 , P2_U3016 );
not NOT1_4931 ( P2_U4350 , P2_U3384 );
nand NAND2_4932 ( P2_U4351 , P2_R1275_U7 , P2_U3031 );
nand NAND2_4933 ( P2_U4352 , P2_U3030 , P2_U3072 );
nand NAND2_4934 ( P2_U4353 , P2_R1215_U114 , P2_U3028 );
nand NAND2_4935 ( P2_U4354 , P2_U3483 , P2_U4132 );
nand NAND2_4936 ( P2_U4355 , P2_U3675 , P2_U4350 );
nand NAND2_4937 ( P2_U4356 , P2_REG2_REG_13_ , P2_U3024 );
nand NAND2_4938 ( P2_U4357 , P2_REG1_REG_13_ , P2_U3025 );
nand NAND2_4939 ( P2_U4358 , P2_REG0_REG_13_ , P2_U3026 );
nand NAND2_4940 ( P2_U4359 , P2_ADD_609_U70 , P2_U3023 );
not NOT1_4941 ( P2_U4360 , P2_U3080 );
nand NAND2_4942 ( P2_U4361 , P2_U3038 , P2_U3063 );
nand NAND2_4943 ( P2_U4362 , P2_R1146_U99 , P2_U3955 );
nand NAND2_4944 ( P2_U4363 , P2_R1113_U99 , P2_U3015 );
nand NAND2_4945 ( P2_U4364 , P2_R1131_U113 , P2_U3014 );
nand NAND2_4946 ( P2_U4365 , P2_R1179_U99 , P2_U3018 );
nand NAND2_4947 ( P2_U4366 , P2_R1203_U99 , P2_U3963 );
nand NAND2_4948 ( P2_U4367 , P2_R1164_U113 , P2_U3959 );
nand NAND2_4949 ( P2_U4368 , P2_R1233_U113 , P2_U3016 );
not NOT1_4950 ( P2_U4369 , P2_U3385 );
nand NAND2_4951 ( P2_U4370 , P2_R1275_U8 , P2_U3031 );
nand NAND2_4952 ( P2_U4371 , P2_U3030 , P2_U3080 );
nand NAND2_4953 ( P2_U4372 , P2_R1215_U113 , P2_U3028 );
nand NAND2_4954 ( P2_U4373 , P2_U3486 , P2_U4132 );
nand NAND2_4955 ( P2_U4374 , P2_U3679 , P2_U4369 );
nand NAND2_4956 ( P2_U4375 , P2_REG2_REG_14_ , P2_U3024 );
nand NAND2_4957 ( P2_U4376 , P2_REG1_REG_14_ , P2_U3025 );
nand NAND2_4958 ( P2_U4377 , P2_REG0_REG_14_ , P2_U3026 );
nand NAND2_4959 ( P2_U4378 , P2_ADD_609_U69 , P2_U3023 );
not NOT1_4960 ( P2_U4379 , P2_U3079 );
nand NAND2_4961 ( P2_U4380 , P2_U3038 , P2_U3072 );
nand NAND2_4962 ( P2_U4381 , P2_R1146_U98 , P2_U3955 );
nand NAND2_4963 ( P2_U4382 , P2_R1113_U98 , P2_U3015 );
nand NAND2_4964 ( P2_U4383 , P2_R1131_U11 , P2_U3014 );
nand NAND2_4965 ( P2_U4384 , P2_R1179_U98 , P2_U3018 );
nand NAND2_4966 ( P2_U4385 , P2_R1203_U98 , P2_U3963 );
nand NAND2_4967 ( P2_U4386 , P2_R1164_U11 , P2_U3959 );
nand NAND2_4968 ( P2_U4387 , P2_R1233_U11 , P2_U3016 );
not NOT1_4969 ( P2_U4388 , P2_U3386 );
nand NAND2_4970 ( P2_U4389 , P2_R1275_U86 , P2_U3031 );
nand NAND2_4971 ( P2_U4390 , P2_U3030 , P2_U3079 );
nand NAND2_4972 ( P2_U4391 , P2_R1215_U11 , P2_U3028 );
nand NAND2_4973 ( P2_U4392 , P2_U3489 , P2_U4132 );
nand NAND2_4974 ( P2_U4393 , P2_U3683 , P2_U4388 );
nand NAND2_4975 ( P2_U4394 , P2_REG2_REG_15_ , P2_U3024 );
nand NAND2_4976 ( P2_U4395 , P2_REG1_REG_15_ , P2_U3025 );
nand NAND2_4977 ( P2_U4396 , P2_REG0_REG_15_ , P2_U3026 );
nand NAND2_4978 ( P2_U4397 , P2_ADD_609_U68 , P2_U3023 );
not NOT1_4979 ( P2_U4398 , P2_U3074 );
nand NAND2_4980 ( P2_U4399 , P2_U3038 , P2_U3080 );
nand NAND2_4981 ( P2_U4400 , P2_R1146_U109 , P2_U3955 );
nand NAND2_4982 ( P2_U4401 , P2_R1113_U109 , P2_U3015 );
nand NAND2_4983 ( P2_U4402 , P2_R1131_U112 , P2_U3014 );
nand NAND2_4984 ( P2_U4403 , P2_R1179_U109 , P2_U3018 );
nand NAND2_4985 ( P2_U4404 , P2_R1203_U109 , P2_U3963 );
nand NAND2_4986 ( P2_U4405 , P2_R1164_U112 , P2_U3959 );
nand NAND2_4987 ( P2_U4406 , P2_R1233_U112 , P2_U3016 );
not NOT1_4988 ( P2_U4407 , P2_U3387 );
nand NAND2_4989 ( P2_U4408 , P2_R1275_U9 , P2_U3031 );
nand NAND2_4990 ( P2_U4409 , P2_U3030 , P2_U3074 );
nand NAND2_4991 ( P2_U4410 , P2_R1215_U112 , P2_U3028 );
nand NAND2_4992 ( P2_U4411 , P2_U3492 , P2_U4132 );
nand NAND2_4993 ( P2_U4412 , P2_U3687 , P2_U4407 );
nand NAND2_4994 ( P2_U4413 , P2_REG2_REG_16_ , P2_U3024 );
nand NAND2_4995 ( P2_U4414 , P2_REG1_REG_16_ , P2_U3025 );
nand NAND2_4996 ( P2_U4415 , P2_REG0_REG_16_ , P2_U3026 );
nand NAND2_4997 ( P2_U4416 , P2_ADD_609_U67 , P2_U3023 );
not NOT1_4998 ( P2_U4417 , P2_U3073 );
nand NAND2_4999 ( P2_U4418 , P2_U3038 , P2_U3079 );
nand NAND2_5000 ( P2_U4419 , P2_R1146_U108 , P2_U3955 );
nand NAND2_5001 ( P2_U4420 , P2_R1113_U108 , P2_U3015 );
nand NAND2_5002 ( P2_U4421 , P2_R1131_U111 , P2_U3014 );
nand NAND2_5003 ( P2_U4422 , P2_R1179_U108 , P2_U3018 );
nand NAND2_5004 ( P2_U4423 , P2_R1203_U108 , P2_U3963 );
nand NAND2_5005 ( P2_U4424 , P2_R1164_U111 , P2_U3959 );
nand NAND2_5006 ( P2_U4425 , P2_R1233_U111 , P2_U3016 );
not NOT1_5007 ( P2_U4426 , P2_U3388 );
nand NAND2_5008 ( P2_U4427 , P2_R1275_U10 , P2_U3031 );
nand NAND2_5009 ( P2_U4428 , P2_U3030 , P2_U3073 );
nand NAND2_5010 ( P2_U4429 , P2_R1215_U111 , P2_U3028 );
nand NAND2_5011 ( P2_U4430 , P2_U3495 , P2_U4132 );
nand NAND2_5012 ( P2_U4431 , P2_U3691 , P2_U4426 );
nand NAND2_5013 ( P2_U4432 , P2_REG2_REG_17_ , P2_U3024 );
nand NAND2_5014 ( P2_U4433 , P2_REG1_REG_17_ , P2_U3025 );
nand NAND2_5015 ( P2_U4434 , P2_REG0_REG_17_ , P2_U3026 );
nand NAND2_5016 ( P2_U4435 , P2_ADD_609_U66 , P2_U3023 );
not NOT1_5017 ( P2_U4436 , P2_U3069 );
nand NAND2_5018 ( P2_U4437 , P2_U3038 , P2_U3074 );
nand NAND2_5019 ( P2_U4438 , P2_R1146_U12 , P2_U3955 );
nand NAND2_5020 ( P2_U4439 , P2_R1113_U12 , P2_U3015 );
nand NAND2_5021 ( P2_U4440 , P2_R1131_U110 , P2_U3014 );
nand NAND2_5022 ( P2_U4441 , P2_R1179_U12 , P2_U3018 );
nand NAND2_5023 ( P2_U4442 , P2_R1203_U12 , P2_U3963 );
nand NAND2_5024 ( P2_U4443 , P2_R1164_U110 , P2_U3959 );
nand NAND2_5025 ( P2_U4444 , P2_R1233_U110 , P2_U3016 );
not NOT1_5026 ( P2_U4445 , P2_U3389 );
nand NAND2_5027 ( P2_U4446 , P2_R1275_U11 , P2_U3031 );
nand NAND2_5028 ( P2_U4447 , P2_U3030 , P2_U3069 );
nand NAND2_5029 ( P2_U4448 , P2_R1215_U110 , P2_U3028 );
nand NAND2_5030 ( P2_U4449 , P2_U3498 , P2_U4132 );
nand NAND2_5031 ( P2_U4450 , P2_U3695 , P2_U4445 );
nand NAND2_5032 ( P2_U4451 , P2_REG2_REG_18_ , P2_U3024 );
nand NAND2_5033 ( P2_U4452 , P2_REG1_REG_18_ , P2_U3025 );
nand NAND2_5034 ( P2_U4453 , P2_REG0_REG_18_ , P2_U3026 );
nand NAND2_5035 ( P2_U4454 , P2_ADD_609_U65 , P2_U3023 );
not NOT1_5036 ( P2_U4455 , P2_U3082 );
nand NAND2_5037 ( P2_U4456 , P2_U3038 , P2_U3073 );
nand NAND2_5038 ( P2_U4457 , P2_R1146_U97 , P2_U3955 );
nand NAND2_5039 ( P2_U4458 , P2_R1113_U97 , P2_U3015 );
nand NAND2_5040 ( P2_U4459 , P2_R1131_U12 , P2_U3014 );
nand NAND2_5041 ( P2_U4460 , P2_R1179_U97 , P2_U3018 );
nand NAND2_5042 ( P2_U4461 , P2_R1203_U97 , P2_U3963 );
nand NAND2_5043 ( P2_U4462 , P2_R1164_U12 , P2_U3959 );
nand NAND2_5044 ( P2_U4463 , P2_R1233_U12 , P2_U3016 );
not NOT1_5045 ( P2_U4464 , P2_U3390 );
nand NAND2_5046 ( P2_U4465 , P2_R1275_U84 , P2_U3031 );
nand NAND2_5047 ( P2_U4466 , P2_U3030 , P2_U3082 );
nand NAND2_5048 ( P2_U4467 , P2_R1215_U12 , P2_U3028 );
nand NAND2_5049 ( P2_U4468 , P2_U3501 , P2_U4132 );
nand NAND2_5050 ( P2_U4469 , P2_U3699 , P2_U4464 );
nand NAND2_5051 ( P2_U4470 , P2_REG2_REG_19_ , P2_U3024 );
nand NAND2_5052 ( P2_U4471 , P2_REG1_REG_19_ , P2_U3025 );
nand NAND2_5053 ( P2_U4472 , P2_REG0_REG_19_ , P2_U3026 );
nand NAND2_5054 ( P2_U4473 , P2_ADD_609_U64 , P2_U3023 );
not NOT1_5055 ( P2_U4474 , P2_U3081 );
nand NAND2_5056 ( P2_U4475 , P2_U3038 , P2_U3069 );
nand NAND2_5057 ( P2_U4476 , P2_R1146_U96 , P2_U3955 );
nand NAND2_5058 ( P2_U4477 , P2_R1113_U96 , P2_U3015 );
nand NAND2_5059 ( P2_U4478 , P2_R1131_U109 , P2_U3014 );
nand NAND2_5060 ( P2_U4479 , P2_R1179_U96 , P2_U3018 );
nand NAND2_5061 ( P2_U4480 , P2_R1203_U96 , P2_U3963 );
nand NAND2_5062 ( P2_U4481 , P2_R1164_U109 , P2_U3959 );
nand NAND2_5063 ( P2_U4482 , P2_R1233_U109 , P2_U3016 );
not NOT1_5064 ( P2_U4483 , P2_U3391 );
nand NAND2_5065 ( P2_U4484 , P2_R1275_U12 , P2_U3031 );
nand NAND2_5066 ( P2_U4485 , P2_U3030 , P2_U3081 );
nand NAND2_5067 ( P2_U4486 , P2_R1215_U109 , P2_U3028 );
nand NAND2_5068 ( P2_U4487 , P2_U3504 , P2_U4132 );
nand NAND2_5069 ( P2_U4488 , P2_U3703 , P2_U4483 );
nand NAND2_5070 ( P2_U4489 , P2_REG2_REG_20_ , P2_U3024 );
nand NAND2_5071 ( P2_U4490 , P2_REG1_REG_20_ , P2_U3025 );
nand NAND2_5072 ( P2_U4491 , P2_REG0_REG_20_ , P2_U3026 );
nand NAND2_5073 ( P2_U4492 , P2_ADD_609_U63 , P2_U3023 );
not NOT1_5074 ( P2_U4493 , P2_U3076 );
nand NAND2_5075 ( P2_U4494 , P2_U3038 , P2_U3082 );
nand NAND2_5076 ( P2_U4495 , P2_R1146_U95 , P2_U3955 );
nand NAND2_5077 ( P2_U4496 , P2_R1113_U95 , P2_U3015 );
nand NAND2_5078 ( P2_U4497 , P2_R1131_U108 , P2_U3014 );
nand NAND2_5079 ( P2_U4498 , P2_R1179_U95 , P2_U3018 );
nand NAND2_5080 ( P2_U4499 , P2_R1203_U95 , P2_U3963 );
nand NAND2_5081 ( P2_U4500 , P2_R1164_U108 , P2_U3959 );
nand NAND2_5082 ( P2_U4501 , P2_R1233_U108 , P2_U3016 );
not NOT1_5083 ( P2_U4502 , P2_U3392 );
nand NAND2_5084 ( P2_U4503 , P2_R1275_U82 , P2_U3031 );
nand NAND2_5085 ( P2_U4504 , P2_U3030 , P2_U3076 );
nand NAND2_5086 ( P2_U4505 , P2_R1215_U108 , P2_U3028 );
nand NAND2_5087 ( P2_U4506 , P2_U3506 , P2_U4132 );
nand NAND2_5088 ( P2_U4507 , P2_U3707 , P2_U4502 );
nand NAND2_5089 ( P2_U4508 , P2_REG2_REG_21_ , P2_U3024 );
nand NAND2_5090 ( P2_U4509 , P2_REG1_REG_21_ , P2_U3025 );
nand NAND2_5091 ( P2_U4510 , P2_REG0_REG_21_ , P2_U3026 );
nand NAND2_5092 ( P2_U4511 , P2_ADD_609_U62 , P2_U3023 );
not NOT1_5093 ( P2_U4512 , P2_U3075 );
nand NAND2_5094 ( P2_U4513 , P2_U3038 , P2_U3081 );
nand NAND2_5095 ( P2_U4514 , P2_R1146_U93 , P2_U3955 );
nand NAND2_5096 ( P2_U4515 , P2_R1113_U93 , P2_U3015 );
nand NAND2_5097 ( P2_U4516 , P2_R1131_U13 , P2_U3014 );
nand NAND2_5098 ( P2_U4517 , P2_R1179_U93 , P2_U3018 );
nand NAND2_5099 ( P2_U4518 , P2_R1203_U93 , P2_U3963 );
nand NAND2_5100 ( P2_U4519 , P2_R1164_U13 , P2_U3959 );
nand NAND2_5101 ( P2_U4520 , P2_R1233_U13 , P2_U3016 );
not NOT1_5102 ( P2_U4521 , P2_U3394 );
nand NAND2_5103 ( P2_U4522 , P2_R1275_U13 , P2_U3031 );
nand NAND2_5104 ( P2_U4523 , P2_U3030 , P2_U3075 );
nand NAND2_5105 ( P2_U4524 , P2_R1215_U13 , P2_U3028 );
nand NAND2_5106 ( P2_U4525 , P2_U3976 , P2_U4132 );
nand NAND2_5107 ( P2_U4526 , P2_U3711 , P2_U4521 );
nand NAND2_5108 ( P2_U4527 , P2_REG2_REG_22_ , P2_U3024 );
nand NAND2_5109 ( P2_U4528 , P2_REG1_REG_22_ , P2_U3025 );
nand NAND2_5110 ( P2_U4529 , P2_REG0_REG_22_ , P2_U3026 );
nand NAND2_5111 ( P2_U4530 , P2_ADD_609_U61 , P2_U3023 );
not NOT1_5112 ( P2_U4531 , P2_U3061 );
nand NAND2_5113 ( P2_U4532 , P2_U3038 , P2_U3076 );
nand NAND2_5114 ( P2_U4533 , P2_R1146_U107 , P2_U3955 );
nand NAND2_5115 ( P2_U4534 , P2_R1113_U107 , P2_U3015 );
nand NAND2_5116 ( P2_U4535 , P2_R1131_U14 , P2_U3014 );
nand NAND2_5117 ( P2_U4536 , P2_R1179_U107 , P2_U3018 );
nand NAND2_5118 ( P2_U4537 , P2_R1203_U107 , P2_U3963 );
nand NAND2_5119 ( P2_U4538 , P2_R1164_U14 , P2_U3959 );
nand NAND2_5120 ( P2_U4539 , P2_R1233_U14 , P2_U3016 );
not NOT1_5121 ( P2_U4540 , P2_U3396 );
nand NAND2_5122 ( P2_U4541 , P2_R1275_U78 , P2_U3031 );
nand NAND2_5123 ( P2_U4542 , P2_U3030 , P2_U3061 );
nand NAND2_5124 ( P2_U4543 , P2_R1215_U14 , P2_U3028 );
nand NAND2_5125 ( P2_U4544 , P2_U3975 , P2_U4132 );
nand NAND2_5126 ( P2_U4545 , P2_U3715 , P2_U4540 );
nand NAND2_5127 ( P2_U4546 , P2_REG2_REG_23_ , P2_U3024 );
nand NAND2_5128 ( P2_U4547 , P2_REG1_REG_23_ , P2_U3025 );
nand NAND2_5129 ( P2_U4548 , P2_REG0_REG_23_ , P2_U3026 );
nand NAND2_5130 ( P2_U4549 , P2_ADD_609_U60 , P2_U3023 );
not NOT1_5131 ( P2_U4550 , P2_U3066 );
nand NAND2_5132 ( P2_U4551 , P2_U3038 , P2_U3075 );
nand NAND2_5133 ( P2_U4552 , P2_R1146_U106 , P2_U3955 );
nand NAND2_5134 ( P2_U4553 , P2_R1113_U106 , P2_U3015 );
nand NAND2_5135 ( P2_U4554 , P2_R1131_U107 , P2_U3014 );
nand NAND2_5136 ( P2_U4555 , P2_R1179_U106 , P2_U3018 );
nand NAND2_5137 ( P2_U4556 , P2_R1203_U106 , P2_U3963 );
nand NAND2_5138 ( P2_U4557 , P2_R1164_U107 , P2_U3959 );
nand NAND2_5139 ( P2_U4558 , P2_R1233_U107 , P2_U3016 );
not NOT1_5140 ( P2_U4559 , P2_U3398 );
nand NAND2_5141 ( P2_U4560 , P2_R1275_U14 , P2_U3031 );
nand NAND2_5142 ( P2_U4561 , P2_U3030 , P2_U3066 );
nand NAND2_5143 ( P2_U4562 , P2_R1215_U107 , P2_U3028 );
nand NAND2_5144 ( P2_U4563 , P2_U3974 , P2_U4132 );
nand NAND2_5145 ( P2_U4564 , P2_U3719 , P2_U4559 );
nand NAND2_5146 ( P2_U4565 , P2_REG2_REG_24_ , P2_U3024 );
nand NAND2_5147 ( P2_U4566 , P2_REG1_REG_24_ , P2_U3025 );
nand NAND2_5148 ( P2_U4567 , P2_REG0_REG_24_ , P2_U3026 );
nand NAND2_5149 ( P2_U4568 , P2_ADD_609_U59 , P2_U3023 );
not NOT1_5150 ( P2_U4569 , P2_U3065 );
nand NAND2_5151 ( P2_U4570 , P2_U3038 , P2_U3061 );
nand NAND2_5152 ( P2_U4571 , P2_R1146_U13 , P2_U3955 );
nand NAND2_5153 ( P2_U4572 , P2_R1113_U13 , P2_U3015 );
nand NAND2_5154 ( P2_U4573 , P2_R1131_U106 , P2_U3014 );
nand NAND2_5155 ( P2_U4574 , P2_R1179_U13 , P2_U3018 );
nand NAND2_5156 ( P2_U4575 , P2_R1203_U13 , P2_U3963 );
nand NAND2_5157 ( P2_U4576 , P2_R1164_U106 , P2_U3959 );
nand NAND2_5158 ( P2_U4577 , P2_R1233_U106 , P2_U3016 );
not NOT1_5159 ( P2_U4578 , P2_U3400 );
nand NAND2_5160 ( P2_U4579 , P2_R1275_U76 , P2_U3031 );
nand NAND2_5161 ( P2_U4580 , P2_U3030 , P2_U3065 );
nand NAND2_5162 ( P2_U4581 , P2_R1215_U106 , P2_U3028 );
nand NAND2_5163 ( P2_U4582 , P2_U3973 , P2_U4132 );
nand NAND2_5164 ( P2_U4583 , P2_U3723 , P2_U4578 );
nand NAND2_5165 ( P2_U4584 , P2_REG2_REG_25_ , P2_U3024 );
nand NAND2_5166 ( P2_U4585 , P2_REG1_REG_25_ , P2_U3025 );
nand NAND2_5167 ( P2_U4586 , P2_REG0_REG_25_ , P2_U3026 );
nand NAND2_5168 ( P2_U4587 , P2_ADD_609_U58 , P2_U3023 );
not NOT1_5169 ( P2_U4588 , P2_U3058 );
nand NAND2_5170 ( P2_U4589 , P2_U3038 , P2_U3066 );
nand NAND2_5171 ( P2_U4590 , P2_R1146_U92 , P2_U3955 );
nand NAND2_5172 ( P2_U4591 , P2_R1113_U92 , P2_U3015 );
nand NAND2_5173 ( P2_U4592 , P2_R1131_U105 , P2_U3014 );
nand NAND2_5174 ( P2_U4593 , P2_R1179_U92 , P2_U3018 );
nand NAND2_5175 ( P2_U4594 , P2_R1203_U92 , P2_U3963 );
nand NAND2_5176 ( P2_U4595 , P2_R1164_U105 , P2_U3959 );
nand NAND2_5177 ( P2_U4596 , P2_R1233_U105 , P2_U3016 );
not NOT1_5178 ( P2_U4597 , P2_U3402 );
nand NAND2_5179 ( P2_U4598 , P2_R1275_U15 , P2_U3031 );
nand NAND2_5180 ( P2_U4599 , P2_U3030 , P2_U3058 );
nand NAND2_5181 ( P2_U4600 , P2_R1215_U105 , P2_U3028 );
nand NAND2_5182 ( P2_U4601 , P2_U3972 , P2_U4132 );
nand NAND2_5183 ( P2_U4602 , P2_U3727 , P2_U4597 );
nand NAND2_5184 ( P2_U4603 , P2_REG2_REG_26_ , P2_U3024 );
nand NAND2_5185 ( P2_U4604 , P2_REG1_REG_26_ , P2_U3025 );
nand NAND2_5186 ( P2_U4605 , P2_REG0_REG_26_ , P2_U3026 );
nand NAND2_5187 ( P2_U4606 , P2_ADD_609_U57 , P2_U3023 );
not NOT1_5188 ( P2_U4607 , P2_U3057 );
nand NAND2_5189 ( P2_U4608 , P2_U3038 , P2_U3065 );
nand NAND2_5190 ( P2_U4609 , P2_R1146_U91 , P2_U3955 );
nand NAND2_5191 ( P2_U4610 , P2_R1113_U91 , P2_U3015 );
nand NAND2_5192 ( P2_U4611 , P2_R1131_U104 , P2_U3014 );
nand NAND2_5193 ( P2_U4612 , P2_R1179_U91 , P2_U3018 );
nand NAND2_5194 ( P2_U4613 , P2_R1203_U91 , P2_U3963 );
nand NAND2_5195 ( P2_U4614 , P2_R1164_U104 , P2_U3959 );
nand NAND2_5196 ( P2_U4615 , P2_R1233_U104 , P2_U3016 );
not NOT1_5197 ( P2_U4616 , P2_U3404 );
nand NAND2_5198 ( P2_U4617 , P2_R1275_U74 , P2_U3031 );
nand NAND2_5199 ( P2_U4618 , P2_U3030 , P2_U3057 );
nand NAND2_5200 ( P2_U4619 , P2_R1215_U104 , P2_U3028 );
nand NAND2_5201 ( P2_U4620 , P2_U3971 , P2_U4132 );
nand NAND2_5202 ( P2_U4621 , P2_U3731 , P2_U4616 );
nand NAND2_5203 ( P2_U4622 , P2_REG2_REG_27_ , P2_U3024 );
nand NAND2_5204 ( P2_U4623 , P2_REG1_REG_27_ , P2_U3025 );
nand NAND2_5205 ( P2_U4624 , P2_REG0_REG_27_ , P2_U3026 );
nand NAND2_5206 ( P2_U4625 , P2_ADD_609_U56 , P2_U3023 );
not NOT1_5207 ( P2_U4626 , P2_U3053 );
nand NAND2_5208 ( P2_U4627 , P2_U3038 , P2_U3058 );
nand NAND2_5209 ( P2_U4628 , P2_R1146_U105 , P2_U3955 );
nand NAND2_5210 ( P2_U4629 , P2_R1113_U105 , P2_U3015 );
nand NAND2_5211 ( P2_U4630 , P2_R1131_U15 , P2_U3014 );
nand NAND2_5212 ( P2_U4631 , P2_R1179_U105 , P2_U3018 );
nand NAND2_5213 ( P2_U4632 , P2_R1203_U105 , P2_U3963 );
nand NAND2_5214 ( P2_U4633 , P2_R1164_U15 , P2_U3959 );
nand NAND2_5215 ( P2_U4634 , P2_R1233_U15 , P2_U3016 );
not NOT1_5216 ( P2_U4635 , P2_U3406 );
nand NAND2_5217 ( P2_U4636 , P2_R1275_U16 , P2_U3031 );
nand NAND2_5218 ( P2_U4637 , P2_U3030 , P2_U3053 );
nand NAND2_5219 ( P2_U4638 , P2_R1215_U15 , P2_U3028 );
nand NAND2_5220 ( P2_U4639 , P2_U3970 , P2_U4132 );
nand NAND2_5221 ( P2_U4640 , P2_U3735 , P2_U4635 );
nand NAND2_5222 ( P2_U4641 , P2_REG2_REG_28_ , P2_U3024 );
nand NAND2_5223 ( P2_U4642 , P2_REG1_REG_28_ , P2_U3025 );
nand NAND2_5224 ( P2_U4643 , P2_REG0_REG_28_ , P2_U3026 );
nand NAND2_5225 ( P2_U4644 , P2_ADD_609_U55 , P2_U3023 );
not NOT1_5226 ( P2_U4645 , P2_U3054 );
nand NAND2_5227 ( P2_U4646 , P2_U3038 , P2_U3057 );
nand NAND2_5228 ( P2_U4647 , P2_R1146_U14 , P2_U3955 );
nand NAND2_5229 ( P2_U4648 , P2_R1113_U14 , P2_U3015 );
nand NAND2_5230 ( P2_U4649 , P2_R1131_U103 , P2_U3014 );
nand NAND2_5231 ( P2_U4650 , P2_R1179_U14 , P2_U3018 );
nand NAND2_5232 ( P2_U4651 , P2_R1203_U14 , P2_U3963 );
nand NAND2_5233 ( P2_U4652 , P2_R1164_U103 , P2_U3959 );
nand NAND2_5234 ( P2_U4653 , P2_R1233_U103 , P2_U3016 );
not NOT1_5235 ( P2_U4654 , P2_U3408 );
nand NAND2_5236 ( P2_U4655 , P2_R1275_U72 , P2_U3031 );
nand NAND2_5237 ( P2_U4656 , P2_U3030 , P2_U3054 );
nand NAND2_5238 ( P2_U4657 , P2_R1215_U103 , P2_U3028 );
nand NAND2_5239 ( P2_U4658 , P2_U3969 , P2_U4132 );
nand NAND2_5240 ( P2_U4659 , P2_U3739 , P2_U4654 );
nand NAND2_5241 ( P2_U4660 , P2_ADD_609_U5 , P2_U3023 );
nand NAND2_5242 ( P2_U4661 , P2_REG2_REG_29_ , P2_U3024 );
nand NAND2_5243 ( P2_U4662 , P2_REG1_REG_29_ , P2_U3025 );
nand NAND2_5244 ( P2_U4663 , P2_REG0_REG_29_ , P2_U3026 );
not NOT1_5245 ( P2_U4664 , P2_U3055 );
nand NAND2_5246 ( P2_U4665 , P2_U3038 , P2_U3053 );
nand NAND2_5247 ( P2_U4666 , P2_R1146_U90 , P2_U3955 );
nand NAND2_5248 ( P2_U4667 , P2_R1113_U90 , P2_U3015 );
nand NAND2_5249 ( P2_U4668 , P2_R1131_U102 , P2_U3014 );
nand NAND2_5250 ( P2_U4669 , P2_R1179_U90 , P2_U3018 );
nand NAND2_5251 ( P2_U4670 , P2_R1203_U90 , P2_U3963 );
nand NAND2_5252 ( P2_U4671 , P2_R1164_U102 , P2_U3959 );
nand NAND2_5253 ( P2_U4672 , P2_R1233_U102 , P2_U3016 );
not NOT1_5254 ( P2_U4673 , P2_U3410 );
nand NAND2_5255 ( P2_U4674 , P2_R1275_U17 , P2_U3031 );
nand NAND2_5256 ( P2_U4675 , P2_U3030 , P2_U3055 );
nand NAND2_5257 ( P2_U4676 , P2_R1215_U102 , P2_U3028 );
nand NAND2_5258 ( P2_U4677 , P2_U3968 , P2_U4132 );
nand NAND2_5259 ( P2_U4678 , P2_U3742 , P2_U4673 );
nand NAND2_5260 ( P2_U4679 , P2_REG2_REG_30_ , P2_U3024 );
nand NAND2_5261 ( P2_U4680 , P2_REG1_REG_30_ , P2_U3025 );
nand NAND2_5262 ( P2_U4681 , P2_REG0_REG_30_ , P2_U3026 );
not NOT1_5263 ( P2_U4682 , P2_U3059 );
nand NAND2_5264 ( P2_U4683 , P2_U5728 , P2_U3360 );
nand NAND2_5265 ( P2_U4684 , P2_U3909 , P2_U4683 );
nand NAND2_5266 ( P2_U4685 , P2_U3743 , P2_U3059 );
nand NAND2_5267 ( P2_U4686 , P2_U3038 , P2_U3054 );
nand NAND2_5268 ( P2_U4687 , P2_R1146_U15 , P2_U3955 );
nand NAND2_5269 ( P2_U4688 , P2_R1113_U15 , P2_U3015 );
nand NAND2_5270 ( P2_U4689 , P2_R1131_U101 , P2_U3014 );
nand NAND2_5271 ( P2_U4690 , P2_R1179_U15 , P2_U3018 );
nand NAND2_5272 ( P2_U4691 , P2_R1203_U15 , P2_U3963 );
nand NAND2_5273 ( P2_U4692 , P2_R1164_U101 , P2_U3959 );
nand NAND2_5274 ( P2_U4693 , P2_R1233_U101 , P2_U3016 );
not NOT1_5275 ( P2_U4694 , P2_U3412 );
nand NAND2_5276 ( P2_U4695 , P2_R1275_U70 , P2_U3031 );
nand NAND2_5277 ( P2_U4696 , P2_R1215_U101 , P2_U3028 );
nand NAND2_5278 ( P2_U4697 , P2_U3979 , P2_U4132 );
nand NAND2_5279 ( P2_U4698 , P2_U3747 , P2_U4694 );
nand NAND2_5280 ( P2_U4699 , P2_REG2_REG_31_ , P2_U3024 );
nand NAND2_5281 ( P2_U4700 , P2_REG1_REG_31_ , P2_U3025 );
nand NAND2_5282 ( P2_U4701 , P2_REG0_REG_31_ , P2_U3026 );
not NOT1_5283 ( P2_U4702 , P2_U3056 );
nand NAND2_5284 ( P2_U4703 , P2_R1275_U19 , P2_U3031 );
nand NAND2_5285 ( P2_U4704 , P2_U3978 , P2_U4132 );
nand NAND3_5286 ( P2_U4705 , P2_U4704 , P2_U3942 , P2_U4703 );
nand NAND2_5287 ( P2_U4706 , P2_R1275_U68 , P2_U3031 );
nand NAND2_5288 ( P2_U4707 , P2_U3977 , P2_U4132 );
nand NAND3_5289 ( P2_U4708 , P2_U4707 , P2_U3942 , P2_U4706 );
nand NAND2_5290 ( P2_U4709 , P2_U3982 , P2_U3439 );
nand NAND2_5291 ( P2_U4710 , P2_U3020 , P2_U3750 );
nand NAND2_5292 ( P2_U4711 , P2_U3418 , P2_U4710 );
nand NAND2_5293 ( P2_U4712 , P2_U3019 , P2_U5708 );
nand NAND2_5294 ( P2_U4713 , P2_U3958 , P2_U4712 );
nand NAND2_5295 ( P2_U4714 , P2_U3040 , P2_U3078 );
nand NAND2_5296 ( P2_U4715 , P2_U3037 , P2_R1215_U95 );
nand NAND2_5297 ( P2_U4716 , P2_U3036 , P2_REG3_REG_0_ );
nand NAND2_5298 ( P2_U4717 , P2_U3035 , P2_U3448 );
nand NAND2_5299 ( P2_U4718 , P2_U3034 , P2_U3448 );
nand NAND2_5300 ( P2_U4719 , P2_U3040 , P2_U3068 );
nand NAND2_5301 ( P2_U4720 , P2_U3037 , P2_R1215_U94 );
nand NAND2_5302 ( P2_U4721 , P2_U3036 , P2_REG3_REG_1_ );
nand NAND2_5303 ( P2_U4722 , P2_U3035 , P2_U3453 );
nand NAND2_5304 ( P2_U4723 , P2_U3034 , P2_R1275_U55 );
nand NAND2_5305 ( P2_U4724 , P2_U3040 , P2_U3064 );
nand NAND2_5306 ( P2_U4725 , P2_U3037 , P2_R1215_U16 );
nand NAND2_5307 ( P2_U4726 , P2_U3036 , P2_REG3_REG_2_ );
nand NAND2_5308 ( P2_U4727 , P2_U3035 , P2_U3456 );
nand NAND2_5309 ( P2_U4728 , P2_U3034 , P2_R1275_U18 );
nand NAND2_5310 ( P2_U4729 , P2_U3040 , P2_U3060 );
nand NAND2_5311 ( P2_U4730 , P2_U3037 , P2_R1215_U100 );
nand NAND2_5312 ( P2_U4731 , P2_U3036 , P2_ADD_609_U4 );
nand NAND2_5313 ( P2_U4732 , P2_U3035 , P2_U3459 );
nand NAND2_5314 ( P2_U4733 , P2_U3034 , P2_R1275_U20 );
nand NAND2_5315 ( P2_U4734 , P2_U3040 , P2_U3067 );
nand NAND2_5316 ( P2_U4735 , P2_U3037 , P2_R1215_U99 );
nand NAND2_5317 ( P2_U4736 , P2_U3036 , P2_ADD_609_U54 );
nand NAND2_5318 ( P2_U4737 , P2_U3035 , P2_U3462 );
nand NAND2_5319 ( P2_U4738 , P2_U3034 , P2_R1275_U21 );
nand NAND2_5320 ( P2_U4739 , P2_U3040 , P2_U3071 );
nand NAND2_5321 ( P2_U4740 , P2_U3037 , P2_R1215_U17 );
nand NAND2_5322 ( P2_U4741 , P2_U3036 , P2_ADD_609_U53 );
nand NAND2_5323 ( P2_U4742 , P2_U3035 , P2_U3465 );
nand NAND2_5324 ( P2_U4743 , P2_U3034 , P2_R1275_U65 );
nand NAND2_5325 ( P2_U4744 , P2_U3040 , P2_U3070 );
nand NAND2_5326 ( P2_U4745 , P2_U3037 , P2_R1215_U98 );
nand NAND2_5327 ( P2_U4746 , P2_U3036 , P2_ADD_609_U52 );
nand NAND2_5328 ( P2_U4747 , P2_U3035 , P2_U3468 );
nand NAND2_5329 ( P2_U4748 , P2_U3034 , P2_R1275_U22 );
nand NAND2_5330 ( P2_U4749 , P2_U3040 , P2_U3084 );
nand NAND2_5331 ( P2_U4750 , P2_U3037 , P2_R1215_U18 );
nand NAND2_5332 ( P2_U4751 , P2_U3036 , P2_ADD_609_U51 );
nand NAND2_5333 ( P2_U4752 , P2_U3035 , P2_U3471 );
nand NAND2_5334 ( P2_U4753 , P2_U3034 , P2_R1275_U23 );
nand NAND2_5335 ( P2_U4754 , P2_U3040 , P2_U3083 );
nand NAND2_5336 ( P2_U4755 , P2_U3037 , P2_R1215_U97 );
nand NAND2_5337 ( P2_U4756 , P2_U3036 , P2_ADD_609_U50 );
nand NAND2_5338 ( P2_U4757 , P2_U3035 , P2_U3474 );
nand NAND2_5339 ( P2_U4758 , P2_U3034 , P2_R1275_U24 );
nand NAND2_5340 ( P2_U4759 , P2_U3040 , P2_U3062 );
nand NAND2_5341 ( P2_U4760 , P2_U3037 , P2_R1215_U96 );
nand NAND2_5342 ( P2_U4761 , P2_U3036 , P2_ADD_609_U49 );
nand NAND2_5343 ( P2_U4762 , P2_U3035 , P2_U3477 );
nand NAND2_5344 ( P2_U4763 , P2_U3034 , P2_R1275_U63 );
nand NAND2_5345 ( P2_U4764 , P2_U3040 , P2_U3063 );
nand NAND2_5346 ( P2_U4765 , P2_U3037 , P2_R1215_U10 );
nand NAND2_5347 ( P2_U4766 , P2_U3036 , P2_ADD_609_U73 );
nand NAND2_5348 ( P2_U4767 , P2_U3035 , P2_U3480 );
nand NAND2_5349 ( P2_U4768 , P2_U3034 , P2_R1275_U6 );
nand NAND2_5350 ( P2_U4769 , P2_U3040 , P2_U3072 );
nand NAND2_5351 ( P2_U4770 , P2_U3037 , P2_R1215_U114 );
nand NAND2_5352 ( P2_U4771 , P2_U3036 , P2_ADD_609_U72 );
nand NAND2_5353 ( P2_U4772 , P2_U3035 , P2_U3483 );
nand NAND2_5354 ( P2_U4773 , P2_U3034 , P2_R1275_U7 );
nand NAND2_5355 ( P2_U4774 , P2_U3040 , P2_U3080 );
nand NAND2_5356 ( P2_U4775 , P2_U3037 , P2_R1215_U113 );
nand NAND2_5357 ( P2_U4776 , P2_U3036 , P2_ADD_609_U71 );
nand NAND2_5358 ( P2_U4777 , P2_U3035 , P2_U3486 );
nand NAND2_5359 ( P2_U4778 , P2_U3034 , P2_R1275_U8 );
nand NAND2_5360 ( P2_U4779 , P2_U3040 , P2_U3079 );
nand NAND2_5361 ( P2_U4780 , P2_U3037 , P2_R1215_U11 );
nand NAND2_5362 ( P2_U4781 , P2_U3036 , P2_ADD_609_U70 );
nand NAND2_5363 ( P2_U4782 , P2_U3035 , P2_U3489 );
nand NAND2_5364 ( P2_U4783 , P2_U3034 , P2_R1275_U86 );
nand NAND2_5365 ( P2_U4784 , P2_U3040 , P2_U3074 );
nand NAND2_5366 ( P2_U4785 , P2_U3037 , P2_R1215_U112 );
nand NAND2_5367 ( P2_U4786 , P2_U3036 , P2_ADD_609_U69 );
nand NAND2_5368 ( P2_U4787 , P2_U3035 , P2_U3492 );
nand NAND2_5369 ( P2_U4788 , P2_U3034 , P2_R1275_U9 );
nand NAND2_5370 ( P2_U4789 , P2_U3040 , P2_U3073 );
nand NAND2_5371 ( P2_U4790 , P2_U3037 , P2_R1215_U111 );
nand NAND2_5372 ( P2_U4791 , P2_U3036 , P2_ADD_609_U68 );
nand NAND2_5373 ( P2_U4792 , P2_U3035 , P2_U3495 );
nand NAND2_5374 ( P2_U4793 , P2_U3034 , P2_R1275_U10 );
nand NAND2_5375 ( P2_U4794 , P2_U3040 , P2_U3069 );
nand NAND2_5376 ( P2_U4795 , P2_U3037 , P2_R1215_U110 );
nand NAND2_5377 ( P2_U4796 , P2_U3036 , P2_ADD_609_U67 );
nand NAND2_5378 ( P2_U4797 , P2_U3035 , P2_U3498 );
nand NAND2_5379 ( P2_U4798 , P2_U3034 , P2_R1275_U11 );
nand NAND2_5380 ( P2_U4799 , P2_U3040 , P2_U3082 );
nand NAND2_5381 ( P2_U4800 , P2_U3037 , P2_R1215_U12 );
nand NAND2_5382 ( P2_U4801 , P2_U3036 , P2_ADD_609_U66 );
nand NAND2_5383 ( P2_U4802 , P2_U3035 , P2_U3501 );
nand NAND2_5384 ( P2_U4803 , P2_U3034 , P2_R1275_U84 );
nand NAND2_5385 ( P2_U4804 , P2_U3040 , P2_U3081 );
nand NAND2_5386 ( P2_U4805 , P2_U3037 , P2_R1215_U109 );
nand NAND2_5387 ( P2_U4806 , P2_U3036 , P2_ADD_609_U65 );
nand NAND2_5388 ( P2_U4807 , P2_U3035 , P2_U3504 );
nand NAND2_5389 ( P2_U4808 , P2_U3034 , P2_R1275_U12 );
nand NAND2_5390 ( P2_U4809 , P2_U3040 , P2_U3076 );
nand NAND2_5391 ( P2_U4810 , P2_U3037 , P2_R1215_U108 );
nand NAND2_5392 ( P2_U4811 , P2_U3036 , P2_ADD_609_U64 );
nand NAND2_5393 ( P2_U4812 , P2_U3035 , P2_U3506 );
nand NAND2_5394 ( P2_U4813 , P2_U3034 , P2_R1275_U82 );
nand NAND2_5395 ( P2_U4814 , P2_U3040 , P2_U3075 );
nand NAND2_5396 ( P2_U4815 , P2_U3037 , P2_R1215_U13 );
nand NAND2_5397 ( P2_U4816 , P2_U3036 , P2_ADD_609_U63 );
nand NAND2_5398 ( P2_U4817 , P2_U3035 , P2_U3976 );
nand NAND2_5399 ( P2_U4818 , P2_U3034 , P2_R1275_U13 );
nand NAND2_5400 ( P2_U4819 , P2_U3040 , P2_U3061 );
nand NAND2_5401 ( P2_U4820 , P2_U3037 , P2_R1215_U14 );
nand NAND2_5402 ( P2_U4821 , P2_U3036 , P2_ADD_609_U62 );
nand NAND2_5403 ( P2_U4822 , P2_U3035 , P2_U3975 );
nand NAND2_5404 ( P2_U4823 , P2_U3034 , P2_R1275_U78 );
nand NAND2_5405 ( P2_U4824 , P2_U3040 , P2_U3066 );
nand NAND2_5406 ( P2_U4825 , P2_U3037 , P2_R1215_U107 );
nand NAND2_5407 ( P2_U4826 , P2_U3036 , P2_ADD_609_U61 );
nand NAND2_5408 ( P2_U4827 , P2_U3035 , P2_U3974 );
nand NAND2_5409 ( P2_U4828 , P2_U3034 , P2_R1275_U14 );
nand NAND2_5410 ( P2_U4829 , P2_U3040 , P2_U3065 );
nand NAND2_5411 ( P2_U4830 , P2_U3037 , P2_R1215_U106 );
nand NAND2_5412 ( P2_U4831 , P2_U3036 , P2_ADD_609_U60 );
nand NAND2_5413 ( P2_U4832 , P2_U3035 , P2_U3973 );
nand NAND2_5414 ( P2_U4833 , P2_U3034 , P2_R1275_U76 );
nand NAND2_5415 ( P2_U4834 , P2_U3040 , P2_U3058 );
nand NAND2_5416 ( P2_U4835 , P2_U3037 , P2_R1215_U105 );
nand NAND2_5417 ( P2_U4836 , P2_U3036 , P2_ADD_609_U59 );
nand NAND2_5418 ( P2_U4837 , P2_U3035 , P2_U3972 );
nand NAND2_5419 ( P2_U4838 , P2_U3034 , P2_R1275_U15 );
nand NAND2_5420 ( P2_U4839 , P2_U3040 , P2_U3057 );
nand NAND2_5421 ( P2_U4840 , P2_U3037 , P2_R1215_U104 );
nand NAND2_5422 ( P2_U4841 , P2_U3036 , P2_ADD_609_U58 );
nand NAND2_5423 ( P2_U4842 , P2_U3035 , P2_U3971 );
nand NAND2_5424 ( P2_U4843 , P2_U3034 , P2_R1275_U74 );
nand NAND2_5425 ( P2_U4844 , P2_U3040 , P2_U3053 );
nand NAND2_5426 ( P2_U4845 , P2_U3037 , P2_R1215_U15 );
nand NAND2_5427 ( P2_U4846 , P2_U3036 , P2_ADD_609_U57 );
nand NAND2_5428 ( P2_U4847 , P2_U3035 , P2_U3970 );
nand NAND2_5429 ( P2_U4848 , P2_U3034 , P2_R1275_U16 );
nand NAND2_5430 ( P2_U4849 , P2_U3040 , P2_U3054 );
nand NAND2_5431 ( P2_U4850 , P2_U3037 , P2_R1215_U103 );
nand NAND2_5432 ( P2_U4851 , P2_U3036 , P2_ADD_609_U56 );
nand NAND2_5433 ( P2_U4852 , P2_U3035 , P2_U3969 );
nand NAND2_5434 ( P2_U4853 , P2_U3034 , P2_R1275_U72 );
nand NAND2_5435 ( P2_U4854 , P2_U3040 , P2_U3055 );
nand NAND2_5436 ( P2_U4855 , P2_U3037 , P2_R1215_U102 );
nand NAND2_5437 ( P2_U4856 , P2_U3036 , P2_ADD_609_U55 );
nand NAND2_5438 ( P2_U4857 , P2_U3035 , P2_U3968 );
nand NAND2_5439 ( P2_U4858 , P2_U3034 , P2_R1275_U17 );
nand NAND2_5440 ( P2_U4859 , P2_U3037 , P2_R1215_U101 );
nand NAND2_5441 ( P2_U4860 , P2_U3036 , P2_ADD_609_U5 );
nand NAND2_5442 ( P2_U4861 , P2_U3035 , P2_U3979 );
nand NAND2_5443 ( P2_U4862 , P2_U3034 , P2_R1275_U70 );
nand NAND2_5444 ( P2_U4863 , P2_U3035 , P2_U3978 );
nand NAND2_5445 ( P2_U4864 , P2_U3034 , P2_R1275_U19 );
nand NAND2_5446 ( P2_U4865 , P2_U3035 , P2_U3977 );
nand NAND2_5447 ( P2_U4866 , P2_U3034 , P2_R1275_U68 );
nand NAND2_5448 ( P2_U4867 , P2_R1170_U13 , P2_U3022 );
nand NAND2_5449 ( P2_U4868 , P2_U5728 , P2_U3445 );
nand NAND2_5450 ( P2_U4869 , P2_R1209_U13 , P2_U5733 );
nand NAND3_5451 ( P2_U4870 , P2_U4868 , P2_U4867 , P2_U4869 );
nand NAND2_5452 ( P2_U4871 , P2_R1170_U13 , P2_U3022 );
nand NAND2_5453 ( P2_U4872 , P2_U3021 , P2_R1209_U13 );
nand NAND2_5454 ( P2_U4873 , P2_U5728 , P2_U3445 );
nand NAND3_5455 ( P2_U4874 , P2_U4872 , P2_U4871 , P2_U4873 );
not NOT1_5456 ( P2_U4875 , P2_U3424 );
nand NAND2_5457 ( P2_U4876 , P2_U3045 , P2_U4870 );
nand NAND2_5458 ( P2_U4877 , P2_U3966 , P2_U4874 );
nand NAND2_5459 ( P2_U4878 , P2_U3044 , P2_R1170_U13 );
nand NAND2_5460 ( P2_U4879 , P2_REG3_REG_19_ , P2_U3152 );
nand NAND2_5461 ( P2_U4880 , P2_U3043 , P2_U3445 );
nand NAND2_5462 ( P2_U4881 , P2_U3042 , P2_R1209_U13 );
nand NAND2_5463 ( P2_U4882 , P2_ADDR_REG_19_ , P2_U4875 );
nand NAND2_5464 ( P2_U4883 , P2_R1170_U75 , P2_U3022 );
nand NAND2_5465 ( P2_U4884 , P2_U5728 , P2_U3503 );
nand NAND2_5466 ( P2_U4885 , P2_R1209_U75 , P2_U5733 );
nand NAND3_5467 ( P2_U4886 , P2_U4884 , P2_U4883 , P2_U4885 );
nand NAND2_5468 ( P2_U4887 , P2_R1170_U75 , P2_U3022 );
nand NAND2_5469 ( P2_U4888 , P2_R1209_U75 , P2_U3021 );
nand NAND2_5470 ( P2_U4889 , P2_U5728 , P2_U3503 );
nand NAND3_5471 ( P2_U4890 , P2_U4888 , P2_U4887 , P2_U4889 );
nand NAND2_5472 ( P2_U4891 , P2_U3045 , P2_U4886 );
nand NAND2_5473 ( P2_U4892 , P2_U3966 , P2_U4890 );
nand NAND2_5474 ( P2_U4893 , P2_R1170_U75 , P2_U3044 );
nand NAND2_5475 ( P2_U4894 , P2_REG3_REG_18_ , P2_U3152 );
nand NAND2_5476 ( P2_U4895 , P2_U3043 , P2_U3503 );
nand NAND2_5477 ( P2_U4896 , P2_R1209_U75 , P2_U3042 );
nand NAND2_5478 ( P2_U4897 , P2_ADDR_REG_18_ , P2_U4875 );
nand NAND2_5479 ( P2_U4898 , P2_R1170_U12 , P2_U3022 );
nand NAND2_5480 ( P2_U4899 , P2_U5728 , P2_U3500 );
nand NAND2_5481 ( P2_U4900 , P2_R1209_U12 , P2_U5733 );
nand NAND3_5482 ( P2_U4901 , P2_U4899 , P2_U4898 , P2_U4900 );
nand NAND2_5483 ( P2_U4902 , P2_R1170_U12 , P2_U3022 );
nand NAND2_5484 ( P2_U4903 , P2_R1209_U12 , P2_U3021 );
nand NAND2_5485 ( P2_U4904 , P2_U5728 , P2_U3500 );
nand NAND3_5486 ( P2_U4905 , P2_U4903 , P2_U4902 , P2_U4904 );
nand NAND2_5487 ( P2_U4906 , P2_U3045 , P2_U4901 );
nand NAND2_5488 ( P2_U4907 , P2_U3966 , P2_U4905 );
nand NAND2_5489 ( P2_U4908 , P2_R1170_U12 , P2_U3044 );
nand NAND2_5490 ( P2_U4909 , P2_REG3_REG_17_ , P2_U3152 );
nand NAND2_5491 ( P2_U4910 , P2_U3043 , P2_U3500 );
nand NAND2_5492 ( P2_U4911 , P2_R1209_U12 , P2_U3042 );
nand NAND2_5493 ( P2_U4912 , P2_ADDR_REG_17_ , P2_U4875 );
nand NAND2_5494 ( P2_U4913 , P2_R1170_U76 , P2_U3022 );
nand NAND2_5495 ( P2_U4914 , P2_U5728 , P2_U3497 );
nand NAND2_5496 ( P2_U4915 , P2_R1209_U76 , P2_U5733 );
nand NAND3_5497 ( P2_U4916 , P2_U4914 , P2_U4913 , P2_U4915 );
nand NAND2_5498 ( P2_U4917 , P2_R1170_U76 , P2_U3022 );
nand NAND2_5499 ( P2_U4918 , P2_R1209_U76 , P2_U3021 );
nand NAND2_5500 ( P2_U4919 , P2_U5728 , P2_U3497 );
nand NAND3_5501 ( P2_U4920 , P2_U4918 , P2_U4917 , P2_U4919 );
nand NAND2_5502 ( P2_U4921 , P2_U3045 , P2_U4916 );
nand NAND2_5503 ( P2_U4922 , P2_U3966 , P2_U4920 );
nand NAND2_5504 ( P2_U4923 , P2_R1170_U76 , P2_U3044 );
nand NAND2_5505 ( P2_U4924 , P2_REG3_REG_16_ , P2_U3152 );
nand NAND2_5506 ( P2_U4925 , P2_U3043 , P2_U3497 );
nand NAND2_5507 ( P2_U4926 , P2_R1209_U76 , P2_U3042 );
nand NAND2_5508 ( P2_U4927 , P2_ADDR_REG_16_ , P2_U4875 );
nand NAND2_5509 ( P2_U4928 , P2_R1170_U77 , P2_U3022 );
nand NAND2_5510 ( P2_U4929 , P2_U5728 , P2_U3494 );
nand NAND2_5511 ( P2_U4930 , P2_R1209_U77 , P2_U5733 );
nand NAND3_5512 ( P2_U4931 , P2_U4929 , P2_U4928 , P2_U4930 );
nand NAND2_5513 ( P2_U4932 , P2_R1170_U77 , P2_U3022 );
nand NAND2_5514 ( P2_U4933 , P2_R1209_U77 , P2_U3021 );
nand NAND2_5515 ( P2_U4934 , P2_U5728 , P2_U3494 );
nand NAND3_5516 ( P2_U4935 , P2_U4933 , P2_U4932 , P2_U4934 );
nand NAND2_5517 ( P2_U4936 , P2_U3045 , P2_U4931 );
nand NAND2_5518 ( P2_U4937 , P2_U3966 , P2_U4935 );
nand NAND2_5519 ( P2_U4938 , P2_R1170_U77 , P2_U3044 );
nand NAND2_5520 ( P2_U4939 , P2_REG3_REG_15_ , P2_U3152 );
nand NAND2_5521 ( P2_U4940 , P2_U3043 , P2_U3494 );
nand NAND2_5522 ( P2_U4941 , P2_R1209_U77 , P2_U3042 );
nand NAND2_5523 ( P2_U4942 , P2_ADDR_REG_15_ , P2_U4875 );
nand NAND2_5524 ( P2_U4943 , P2_R1170_U78 , P2_U3022 );
nand NAND2_5525 ( P2_U4944 , P2_U5728 , P2_U3491 );
nand NAND2_5526 ( P2_U4945 , P2_R1209_U78 , P2_U5733 );
nand NAND3_5527 ( P2_U4946 , P2_U4944 , P2_U4943 , P2_U4945 );
nand NAND2_5528 ( P2_U4947 , P2_R1170_U78 , P2_U3022 );
nand NAND2_5529 ( P2_U4948 , P2_R1209_U78 , P2_U3021 );
nand NAND2_5530 ( P2_U4949 , P2_U5728 , P2_U3491 );
nand NAND3_5531 ( P2_U4950 , P2_U4948 , P2_U4947 , P2_U4949 );
nand NAND2_5532 ( P2_U4951 , P2_U3045 , P2_U4946 );
nand NAND2_5533 ( P2_U4952 , P2_U3966 , P2_U4950 );
nand NAND2_5534 ( P2_U4953 , P2_R1170_U78 , P2_U3044 );
nand NAND2_5535 ( P2_U4954 , P2_REG3_REG_14_ , P2_U3152 );
nand NAND2_5536 ( P2_U4955 , P2_U3043 , P2_U3491 );
nand NAND2_5537 ( P2_U4956 , P2_R1209_U78 , P2_U3042 );
nand NAND2_5538 ( P2_U4957 , P2_ADDR_REG_14_ , P2_U4875 );
nand NAND2_5539 ( P2_U4958 , P2_R1170_U11 , P2_U3022 );
nand NAND2_5540 ( P2_U4959 , P2_U5728 , P2_U3488 );
nand NAND2_5541 ( P2_U4960 , P2_R1209_U11 , P2_U5733 );
nand NAND3_5542 ( P2_U4961 , P2_U4959 , P2_U4958 , P2_U4960 );
nand NAND2_5543 ( P2_U4962 , P2_R1170_U11 , P2_U3022 );
nand NAND2_5544 ( P2_U4963 , P2_R1209_U11 , P2_U3021 );
nand NAND2_5545 ( P2_U4964 , P2_U5728 , P2_U3488 );
nand NAND3_5546 ( P2_U4965 , P2_U4963 , P2_U4962 , P2_U4964 );
nand NAND2_5547 ( P2_U4966 , P2_U3045 , P2_U4961 );
nand NAND2_5548 ( P2_U4967 , P2_U3966 , P2_U4965 );
nand NAND2_5549 ( P2_U4968 , P2_R1170_U11 , P2_U3044 );
nand NAND2_5550 ( P2_U4969 , P2_REG3_REG_13_ , P2_U3152 );
nand NAND2_5551 ( P2_U4970 , P2_U3043 , P2_U3488 );
nand NAND2_5552 ( P2_U4971 , P2_R1209_U11 , P2_U3042 );
nand NAND2_5553 ( P2_U4972 , P2_ADDR_REG_13_ , P2_U4875 );
nand NAND2_5554 ( P2_U4973 , P2_R1170_U79 , P2_U3022 );
nand NAND2_5555 ( P2_U4974 , P2_U5728 , P2_U3485 );
nand NAND2_5556 ( P2_U4975 , P2_R1209_U79 , P2_U5733 );
nand NAND3_5557 ( P2_U4976 , P2_U4974 , P2_U4973 , P2_U4975 );
nand NAND2_5558 ( P2_U4977 , P2_R1170_U79 , P2_U3022 );
nand NAND2_5559 ( P2_U4978 , P2_R1209_U79 , P2_U3021 );
nand NAND2_5560 ( P2_U4979 , P2_U5728 , P2_U3485 );
nand NAND3_5561 ( P2_U4980 , P2_U4978 , P2_U4977 , P2_U4979 );
nand NAND2_5562 ( P2_U4981 , P2_U3045 , P2_U4976 );
nand NAND2_5563 ( P2_U4982 , P2_U3966 , P2_U4980 );
nand NAND2_5564 ( P2_U4983 , P2_R1170_U79 , P2_U3044 );
nand NAND2_5565 ( P2_U4984 , P2_REG3_REG_12_ , P2_U3152 );
nand NAND2_5566 ( P2_U4985 , P2_U3043 , P2_U3485 );
nand NAND2_5567 ( P2_U4986 , P2_R1209_U79 , P2_U3042 );
nand NAND2_5568 ( P2_U4987 , P2_ADDR_REG_12_ , P2_U4875 );
nand NAND2_5569 ( P2_U4988 , P2_R1170_U80 , P2_U3022 );
nand NAND2_5570 ( P2_U4989 , P2_U5728 , P2_U3482 );
nand NAND2_5571 ( P2_U4990 , P2_R1209_U80 , P2_U5733 );
nand NAND3_5572 ( P2_U4991 , P2_U4989 , P2_U4988 , P2_U4990 );
nand NAND2_5573 ( P2_U4992 , P2_R1170_U80 , P2_U3022 );
nand NAND2_5574 ( P2_U4993 , P2_R1209_U80 , P2_U3021 );
nand NAND2_5575 ( P2_U4994 , P2_U5728 , P2_U3482 );
nand NAND3_5576 ( P2_U4995 , P2_U4993 , P2_U4992 , P2_U4994 );
nand NAND2_5577 ( P2_U4996 , P2_U3045 , P2_U4991 );
nand NAND2_5578 ( P2_U4997 , P2_U3966 , P2_U4995 );
nand NAND2_5579 ( P2_U4998 , P2_R1170_U80 , P2_U3044 );
nand NAND2_5580 ( P2_U4999 , P2_REG3_REG_11_ , P2_U3152 );
nand NAND2_5581 ( P2_U5000 , P2_U3043 , P2_U3482 );
nand NAND2_5582 ( P2_U5001 , P2_R1209_U80 , P2_U3042 );
nand NAND2_5583 ( P2_U5002 , P2_ADDR_REG_11_ , P2_U4875 );
nand NAND2_5584 ( P2_U5003 , P2_R1170_U10 , P2_U3022 );
nand NAND2_5585 ( P2_U5004 , P2_U5728 , P2_U3479 );
nand NAND2_5586 ( P2_U5005 , P2_R1209_U10 , P2_U5733 );
nand NAND3_5587 ( P2_U5006 , P2_U5004 , P2_U5003 , P2_U5005 );
nand NAND2_5588 ( P2_U5007 , P2_R1170_U10 , P2_U3022 );
nand NAND2_5589 ( P2_U5008 , P2_R1209_U10 , P2_U3021 );
nand NAND2_5590 ( P2_U5009 , P2_U5728 , P2_U3479 );
nand NAND3_5591 ( P2_U5010 , P2_U5008 , P2_U5007 , P2_U5009 );
nand NAND2_5592 ( P2_U5011 , P2_U3045 , P2_U5006 );
nand NAND2_5593 ( P2_U5012 , P2_U3966 , P2_U5010 );
nand NAND2_5594 ( P2_U5013 , P2_R1170_U10 , P2_U3044 );
nand NAND2_5595 ( P2_U5014 , P2_REG3_REG_10_ , P2_U3152 );
nand NAND2_5596 ( P2_U5015 , P2_U3043 , P2_U3479 );
nand NAND2_5597 ( P2_U5016 , P2_R1209_U10 , P2_U3042 );
nand NAND2_5598 ( P2_U5017 , P2_ADDR_REG_10_ , P2_U4875 );
nand NAND2_5599 ( P2_U5018 , P2_R1170_U70 , P2_U3022 );
nand NAND2_5600 ( P2_U5019 , P2_U5728 , P2_U3476 );
nand NAND2_5601 ( P2_U5020 , P2_R1209_U70 , P2_U5733 );
nand NAND3_5602 ( P2_U5021 , P2_U5019 , P2_U5018 , P2_U5020 );
nand NAND2_5603 ( P2_U5022 , P2_R1170_U70 , P2_U3022 );
nand NAND2_5604 ( P2_U5023 , P2_R1209_U70 , P2_U3021 );
nand NAND2_5605 ( P2_U5024 , P2_U5728 , P2_U3476 );
nand NAND3_5606 ( P2_U5025 , P2_U5023 , P2_U5022 , P2_U5024 );
nand NAND2_5607 ( P2_U5026 , P2_U3045 , P2_U5021 );
nand NAND2_5608 ( P2_U5027 , P2_U3966 , P2_U5025 );
nand NAND2_5609 ( P2_U5028 , P2_R1170_U70 , P2_U3044 );
nand NAND2_5610 ( P2_U5029 , P2_REG3_REG_9_ , P2_U3152 );
nand NAND2_5611 ( P2_U5030 , P2_U3043 , P2_U3476 );
nand NAND2_5612 ( P2_U5031 , P2_R1209_U70 , P2_U3042 );
nand NAND2_5613 ( P2_U5032 , P2_ADDR_REG_9_ , P2_U4875 );
nand NAND2_5614 ( P2_U5033 , P2_R1170_U71 , P2_U3022 );
nand NAND2_5615 ( P2_U5034 , P2_U5728 , P2_U3473 );
nand NAND2_5616 ( P2_U5035 , P2_R1209_U71 , P2_U5733 );
nand NAND3_5617 ( P2_U5036 , P2_U5034 , P2_U5033 , P2_U5035 );
nand NAND2_5618 ( P2_U5037 , P2_R1170_U71 , P2_U3022 );
nand NAND2_5619 ( P2_U5038 , P2_R1209_U71 , P2_U3021 );
nand NAND2_5620 ( P2_U5039 , P2_U5728 , P2_U3473 );
nand NAND3_5621 ( P2_U5040 , P2_U5038 , P2_U5037 , P2_U5039 );
nand NAND2_5622 ( P2_U5041 , P2_U3045 , P2_U5036 );
nand NAND2_5623 ( P2_U5042 , P2_U3966 , P2_U5040 );
nand NAND2_5624 ( P2_U5043 , P2_R1170_U71 , P2_U3044 );
nand NAND2_5625 ( P2_U5044 , P2_REG3_REG_8_ , P2_U3152 );
nand NAND2_5626 ( P2_U5045 , P2_U3043 , P2_U3473 );
nand NAND2_5627 ( P2_U5046 , P2_R1209_U71 , P2_U3042 );
nand NAND2_5628 ( P2_U5047 , P2_ADDR_REG_8_ , P2_U4875 );
nand NAND2_5629 ( P2_U5048 , P2_R1170_U16 , P2_U3022 );
nand NAND2_5630 ( P2_U5049 , P2_U5728 , P2_U3470 );
nand NAND2_5631 ( P2_U5050 , P2_R1209_U16 , P2_U5733 );
nand NAND3_5632 ( P2_U5051 , P2_U5049 , P2_U5048 , P2_U5050 );
nand NAND2_5633 ( P2_U5052 , P2_R1170_U16 , P2_U3022 );
nand NAND2_5634 ( P2_U5053 , P2_R1209_U16 , P2_U3021 );
nand NAND2_5635 ( P2_U5054 , P2_U5728 , P2_U3470 );
nand NAND3_5636 ( P2_U5055 , P2_U5053 , P2_U5052 , P2_U5054 );
nand NAND2_5637 ( P2_U5056 , P2_U3045 , P2_U5051 );
nand NAND2_5638 ( P2_U5057 , P2_U3966 , P2_U5055 );
nand NAND2_5639 ( P2_U5058 , P2_R1170_U16 , P2_U3044 );
nand NAND2_5640 ( P2_U5059 , P2_REG3_REG_7_ , P2_U3152 );
nand NAND2_5641 ( P2_U5060 , P2_U3043 , P2_U3470 );
nand NAND2_5642 ( P2_U5061 , P2_R1209_U16 , P2_U3042 );
nand NAND2_5643 ( P2_U5062 , P2_ADDR_REG_7_ , P2_U4875 );
nand NAND2_5644 ( P2_U5063 , P2_R1170_U72 , P2_U3022 );
nand NAND2_5645 ( P2_U5064 , P2_U5728 , P2_U3467 );
nand NAND2_5646 ( P2_U5065 , P2_R1209_U72 , P2_U5733 );
nand NAND3_5647 ( P2_U5066 , P2_U5064 , P2_U5063 , P2_U5065 );
nand NAND2_5648 ( P2_U5067 , P2_R1170_U72 , P2_U3022 );
nand NAND2_5649 ( P2_U5068 , P2_R1209_U72 , P2_U3021 );
nand NAND2_5650 ( P2_U5069 , P2_U5728 , P2_U3467 );
nand NAND3_5651 ( P2_U5070 , P2_U5068 , P2_U5067 , P2_U5069 );
nand NAND2_5652 ( P2_U5071 , P2_U3045 , P2_U5066 );
nand NAND2_5653 ( P2_U5072 , P2_U3966 , P2_U5070 );
nand NAND2_5654 ( P2_U5073 , P2_R1170_U72 , P2_U3044 );
nand NAND2_5655 ( P2_U5074 , P2_REG3_REG_6_ , P2_U3152 );
nand NAND2_5656 ( P2_U5075 , P2_U3043 , P2_U3467 );
nand NAND2_5657 ( P2_U5076 , P2_R1209_U72 , P2_U3042 );
nand NAND2_5658 ( P2_U5077 , P2_ADDR_REG_6_ , P2_U4875 );
nand NAND2_5659 ( P2_U5078 , P2_R1170_U15 , P2_U3022 );
nand NAND2_5660 ( P2_U5079 , P2_U5728 , P2_U3464 );
nand NAND2_5661 ( P2_U5080 , P2_R1209_U15 , P2_U5733 );
nand NAND3_5662 ( P2_U5081 , P2_U5079 , P2_U5078 , P2_U5080 );
nand NAND2_5663 ( P2_U5082 , P2_R1170_U15 , P2_U3022 );
nand NAND2_5664 ( P2_U5083 , P2_R1209_U15 , P2_U3021 );
nand NAND2_5665 ( P2_U5084 , P2_U5728 , P2_U3464 );
nand NAND3_5666 ( P2_U5085 , P2_U5083 , P2_U5082 , P2_U5084 );
nand NAND2_5667 ( P2_U5086 , P2_U3045 , P2_U5081 );
nand NAND2_5668 ( P2_U5087 , P2_U3966 , P2_U5085 );
nand NAND2_5669 ( P2_U5088 , P2_R1170_U15 , P2_U3044 );
nand NAND2_5670 ( P2_U5089 , P2_REG3_REG_5_ , P2_U3152 );
nand NAND2_5671 ( P2_U5090 , P2_U3043 , P2_U3464 );
nand NAND2_5672 ( P2_U5091 , P2_R1209_U15 , P2_U3042 );
nand NAND2_5673 ( P2_U5092 , P2_ADDR_REG_5_ , P2_U4875 );
nand NAND2_5674 ( P2_U5093 , P2_R1170_U73 , P2_U3022 );
nand NAND2_5675 ( P2_U5094 , P2_U5728 , P2_U3461 );
nand NAND2_5676 ( P2_U5095 , P2_R1209_U73 , P2_U5733 );
nand NAND3_5677 ( P2_U5096 , P2_U5094 , P2_U5093 , P2_U5095 );
nand NAND2_5678 ( P2_U5097 , P2_R1170_U73 , P2_U3022 );
nand NAND2_5679 ( P2_U5098 , P2_R1209_U73 , P2_U3021 );
nand NAND2_5680 ( P2_U5099 , P2_U5728 , P2_U3461 );
nand NAND3_5681 ( P2_U5100 , P2_U5098 , P2_U5097 , P2_U5099 );
nand NAND2_5682 ( P2_U5101 , P2_U3045 , P2_U5096 );
nand NAND2_5683 ( P2_U5102 , P2_U3966 , P2_U5100 );
nand NAND2_5684 ( P2_U5103 , P2_R1170_U73 , P2_U3044 );
nand NAND2_5685 ( P2_U5104 , P2_REG3_REG_4_ , P2_U3152 );
nand NAND2_5686 ( P2_U5105 , P2_U3043 , P2_U3461 );
nand NAND2_5687 ( P2_U5106 , P2_R1209_U73 , P2_U3042 );
nand NAND2_5688 ( P2_U5107 , P2_ADDR_REG_4_ , P2_U4875 );
nand NAND2_5689 ( P2_U5108 , P2_R1170_U74 , P2_U3022 );
nand NAND2_5690 ( P2_U5109 , P2_U5728 , P2_U3458 );
nand NAND2_5691 ( P2_U5110 , P2_R1209_U74 , P2_U5733 );
nand NAND3_5692 ( P2_U5111 , P2_U5109 , P2_U5108 , P2_U5110 );
nand NAND2_5693 ( P2_U5112 , P2_R1170_U74 , P2_U3022 );
nand NAND2_5694 ( P2_U5113 , P2_R1209_U74 , P2_U3021 );
nand NAND2_5695 ( P2_U5114 , P2_U5728 , P2_U3458 );
nand NAND3_5696 ( P2_U5115 , P2_U5113 , P2_U5112 , P2_U5114 );
nand NAND2_5697 ( P2_U5116 , P2_U3045 , P2_U5111 );
nand NAND2_5698 ( P2_U5117 , P2_U3966 , P2_U5115 );
nand NAND2_5699 ( P2_U5118 , P2_R1170_U74 , P2_U3044 );
nand NAND2_5700 ( P2_U5119 , P2_REG3_REG_3_ , P2_U3152 );
nand NAND2_5701 ( P2_U5120 , P2_U3043 , P2_U3458 );
nand NAND2_5702 ( P2_U5121 , P2_R1209_U74 , P2_U3042 );
nand NAND2_5703 ( P2_U5122 , P2_ADDR_REG_3_ , P2_U4875 );
nand NAND2_5704 ( P2_U5123 , P2_R1170_U14 , P2_U3022 );
nand NAND2_5705 ( P2_U5124 , P2_U5728 , P2_U3455 );
nand NAND2_5706 ( P2_U5125 , P2_R1209_U14 , P2_U5733 );
nand NAND3_5707 ( P2_U5126 , P2_U5124 , P2_U5123 , P2_U5125 );
nand NAND2_5708 ( P2_U5127 , P2_R1170_U14 , P2_U3022 );
nand NAND2_5709 ( P2_U5128 , P2_R1209_U14 , P2_U3021 );
nand NAND2_5710 ( P2_U5129 , P2_U5728 , P2_U3455 );
nand NAND3_5711 ( P2_U5130 , P2_U5128 , P2_U5127 , P2_U5129 );
nand NAND2_5712 ( P2_U5131 , P2_U3045 , P2_U5126 );
nand NAND2_5713 ( P2_U5132 , P2_U3966 , P2_U5130 );
nand NAND2_5714 ( P2_U5133 , P2_R1170_U14 , P2_U3044 );
nand NAND2_5715 ( P2_U5134 , P2_REG3_REG_2_ , P2_U3152 );
nand NAND2_5716 ( P2_U5135 , P2_U3043 , P2_U3455 );
nand NAND2_5717 ( P2_U5136 , P2_R1209_U14 , P2_U3042 );
nand NAND2_5718 ( P2_U5137 , P2_ADDR_REG_2_ , P2_U4875 );
nand NAND2_5719 ( P2_U5138 , P2_R1170_U68 , P2_U3022 );
nand NAND2_5720 ( P2_U5139 , P2_U5728 , P2_U3452 );
nand NAND2_5721 ( P2_U5140 , P2_R1209_U68 , P2_U5733 );
nand NAND3_5722 ( P2_U5141 , P2_U5139 , P2_U5138 , P2_U5140 );
nand NAND2_5723 ( P2_U5142 , P2_R1170_U68 , P2_U3022 );
nand NAND2_5724 ( P2_U5143 , P2_R1209_U68 , P2_U3021 );
nand NAND2_5725 ( P2_U5144 , P2_U5728 , P2_U3452 );
nand NAND3_5726 ( P2_U5145 , P2_U5143 , P2_U5142 , P2_U5144 );
nand NAND2_5727 ( P2_U5146 , P2_U3045 , P2_U5141 );
nand NAND2_5728 ( P2_U5147 , P2_U3966 , P2_U5145 );
nand NAND2_5729 ( P2_U5148 , P2_R1170_U68 , P2_U3044 );
nand NAND2_5730 ( P2_U5149 , P2_REG3_REG_1_ , P2_U3152 );
nand NAND2_5731 ( P2_U5150 , P2_U3043 , P2_U3452 );
nand NAND2_5732 ( P2_U5151 , P2_R1209_U68 , P2_U3042 );
nand NAND2_5733 ( P2_U5152 , P2_ADDR_REG_1_ , P2_U4875 );
nand NAND2_5734 ( P2_U5153 , P2_R1170_U69 , P2_U3022 );
nand NAND2_5735 ( P2_U5154 , P2_U5728 , P2_U3446 );
nand NAND2_5736 ( P2_U5155 , P2_R1209_U69 , P2_U5733 );
nand NAND2_5737 ( P2_U5156 , P2_U3869 , P2_U5153 );
nand NAND2_5738 ( P2_U5157 , P2_R1170_U69 , P2_U3022 );
nand NAND2_5739 ( P2_U5158 , P2_R1209_U69 , P2_U3021 );
nand NAND2_5740 ( P2_U5159 , P2_U5728 , P2_U3446 );
nand NAND3_5741 ( P2_U5160 , P2_U5158 , P2_U5157 , P2_U5159 );
nand NAND2_5742 ( P2_U5161 , P2_U3045 , P2_U5156 );
nand NAND2_5743 ( P2_U5162 , P2_U3966 , P2_U5160 );
nand NAND2_5744 ( P2_U5163 , P2_R1170_U69 , P2_U3044 );
nand NAND2_5745 ( P2_U5164 , P2_REG3_REG_0_ , P2_U3152 );
nand NAND2_5746 ( P2_U5165 , P2_U3043 , P2_U3446 );
nand NAND2_5747 ( P2_U5166 , P2_R1209_U69 , P2_U3042 );
nand NAND2_5748 ( P2_U5167 , P2_ADDR_REG_0_ , P2_U4875 );
not NOT1_5749 ( P2_U5168 , P2_U3947 );
nand NAND2_5750 ( P2_U5169 , P2_U3363 , P2_U3416 );
nand NAND2_5751 ( P2_U5170 , P2_U3366 , P2_U3428 );
nand NAND2_5752 ( P2_U5171 , P2_U3419 , P2_U3364 );
nand NAND3_5753 ( P2_U5172 , P2_U6099 , P2_U6098 , P2_U3018 );
nand NAND2_5754 ( P2_U5173 , P2_R1340_U6 , P2_U5171 );
nand NAND4_5755 ( P2_U5174 , P2_U6201 , P2_U6200 , P2_U3946 , P2_U3885 );
nand NAND3_5756 ( P2_U5175 , P2_U6101 , P2_U6100 , P2_U3052 );
nand NAND2_5757 ( P2_U5176 , P2_U3980 , P2_U3027 );
nand NAND2_5758 ( P2_U5177 , P2_B_REG , P2_U5175 );
nand NAND2_5759 ( P2_U5178 , P2_U3041 , P2_U3079 );
nand NAND2_5760 ( P2_U5179 , P2_U3039 , P2_U3073 );
nand NAND2_5761 ( P2_U5180 , P2_ADD_609_U68 , P2_U3427 );
nand NAND3_5762 ( P2_U5181 , P2_U5179 , P2_U5178 , P2_U5180 );
nand NAND2_5763 ( P2_U5182 , P2_U3014 , P2_U5717 );
nand NAND5_5764 ( P2_U5183 , P2_U3369 , P2_U3367 , P2_U5182 , P2_U3888 , P2_U3419 );
nand NAND2_5765 ( P2_U5184 , P2_U5183 , P2_U3427 );
not NOT1_5766 ( P2_U5185 , P2_U3430 );
nand NAND2_5767 ( P2_U5186 , P2_U3495 , P2_U5678 );
nand NAND2_5768 ( P2_U5187 , P2_ADD_609_U68 , P2_U5677 );
nand NAND2_5769 ( P2_U5188 , P2_U3988 , P2_U5181 );
nand NAND2_5770 ( P2_U5189 , P2_R1176_U102 , P2_U3032 );
nand NAND2_5771 ( P2_U5190 , P2_REG3_REG_15_ , P2_U3152 );
nand NAND2_5772 ( P2_U5191 , P2_U3041 , P2_U3058 );
nand NAND2_5773 ( P2_U5192 , P2_U3039 , P2_U3053 );
nand NAND2_5774 ( P2_U5193 , P2_ADD_609_U57 , P2_U3427 );
nand NAND3_5775 ( P2_U5194 , P2_U5193 , P2_U5191 , P2_U5192 );
nand NAND2_5776 ( P2_U5195 , P2_U4713 , P2_U3427 );
nand NAND2_5777 ( P2_U5196 , P2_U5185 , P2_U5195 );
nand NAND2_5778 ( P2_U5197 , P2_U3965 , P2_U4713 );
nand NAND2_5779 ( P2_U5198 , P2_U3418 , P2_U5197 );
nand NAND2_5780 ( P2_U5199 , P2_U3047 , P2_U3970 );
nand NAND2_5781 ( P2_U5200 , P2_U3046 , P2_ADD_609_U57 );
nand NAND2_5782 ( P2_U5201 , P2_U3988 , P2_U5194 );
nand NAND2_5783 ( P2_U5202 , P2_R1176_U12 , P2_U3032 );
nand NAND2_5784 ( P2_U5203 , P2_REG3_REG_26_ , P2_U3152 );
nand NAND2_5785 ( P2_U5204 , P2_U3041 , P2_U3067 );
nand NAND2_5786 ( P2_U5205 , P2_U3039 , P2_U3070 );
nand NAND2_5787 ( P2_U5206 , P2_ADD_609_U52 , P2_U3427 );
nand NAND3_5788 ( P2_U5207 , P2_U5205 , P2_U5204 , P2_U5206 );
nand NAND2_5789 ( P2_U5208 , P2_U3468 , P2_U5678 );
nand NAND2_5790 ( P2_U5209 , P2_ADD_609_U52 , P2_U5677 );
nand NAND2_5791 ( P2_U5210 , P2_U3988 , P2_U5207 );
nand NAND2_5792 ( P2_U5211 , P2_R1176_U87 , P2_U3032 );
nand NAND2_5793 ( P2_U5212 , P2_REG3_REG_6_ , P2_U3152 );
nand NAND2_5794 ( P2_U5213 , P2_U3041 , P2_U3069 );
nand NAND2_5795 ( P2_U5214 , P2_U3039 , P2_U3081 );
nand NAND2_5796 ( P2_U5215 , P2_ADD_609_U65 , P2_U3427 );
nand NAND3_5797 ( P2_U5216 , P2_U5214 , P2_U5213 , P2_U5215 );
nand NAND2_5798 ( P2_U5217 , P2_U3504 , P2_U5678 );
nand NAND2_5799 ( P2_U5218 , P2_ADD_609_U65 , P2_U5677 );
nand NAND2_5800 ( P2_U5219 , P2_U3988 , P2_U5216 );
nand NAND2_5801 ( P2_U5220 , P2_R1176_U100 , P2_U3032 );
nand NAND2_5802 ( P2_U5221 , P2_REG3_REG_18_ , P2_U3152 );
nand NAND2_5803 ( P2_U5222 , P2_U3041 , P2_U3078 );
nand NAND2_5804 ( P2_U5223 , P2_U3039 , P2_U3064 );
nand NAND2_5805 ( P2_U5224 , P2_REG3_REG_2_ , P2_U3427 );
nand NAND3_5806 ( P2_U5225 , P2_U5223 , P2_U5222 , P2_U5224 );
nand NAND2_5807 ( P2_U5226 , P2_U3456 , P2_U5678 );
nand NAND2_5808 ( P2_U5227 , P2_REG3_REG_2_ , P2_U5677 );
nand NAND2_5809 ( P2_U5228 , P2_U3988 , P2_U5225 );
nand NAND2_5810 ( P2_U5229 , P2_R1176_U90 , P2_U3032 );
nand NAND2_5811 ( P2_U5230 , P2_REG3_REG_2_ , P2_U3152 );
nand NAND2_5812 ( P2_U5231 , P2_U3041 , P2_U3062 );
nand NAND2_5813 ( P2_U5232 , P2_U3039 , P2_U3072 );
nand NAND2_5814 ( P2_U5233 , P2_ADD_609_U72 , P2_U3427 );
nand NAND3_5815 ( P2_U5234 , P2_U5232 , P2_U5231 , P2_U5233 );
nand NAND2_5816 ( P2_U5235 , P2_U3483 , P2_U5678 );
nand NAND2_5817 ( P2_U5236 , P2_ADD_609_U72 , P2_U5677 );
nand NAND2_5818 ( P2_U5237 , P2_U3988 , P2_U5234 );
nand NAND2_5819 ( P2_U5238 , P2_R1176_U105 , P2_U3032 );
nand NAND2_5820 ( P2_U5239 , P2_REG3_REG_11_ , P2_U3152 );
nand NAND2_5821 ( P2_U5240 , P2_U3041 , P2_U3075 );
nand NAND2_5822 ( P2_U5241 , P2_U3039 , P2_U3066 );
nand NAND2_5823 ( P2_U5242 , P2_ADD_609_U61 , P2_U3427 );
nand NAND3_5824 ( P2_U5243 , P2_U5242 , P2_U5240 , P2_U5241 );
nand NAND2_5825 ( P2_U5244 , P2_U3047 , P2_U3974 );
nand NAND2_5826 ( P2_U5245 , P2_U3046 , P2_ADD_609_U61 );
nand NAND2_5827 ( P2_U5246 , P2_U3988 , P2_U5243 );
nand NAND2_5828 ( P2_U5247 , P2_R1176_U96 , P2_U3032 );
nand NAND2_5829 ( P2_U5248 , P2_REG3_REG_22_ , P2_U3152 );
nand NAND2_5830 ( P2_U5249 , P2_U3041 , P2_U3072 );
nand NAND2_5831 ( P2_U5250 , P2_U3039 , P2_U3079 );
nand NAND2_5832 ( P2_U5251 , P2_ADD_609_U70 , P2_U3427 );
nand NAND3_5833 ( P2_U5252 , P2_U5250 , P2_U5249 , P2_U5251 );
nand NAND2_5834 ( P2_U5253 , P2_U3489 , P2_U5678 );
nand NAND2_5835 ( P2_U5254 , P2_ADD_609_U70 , P2_U5677 );
nand NAND2_5836 ( P2_U5255 , P2_U3988 , P2_U5252 );
nand NAND2_5837 ( P2_U5256 , P2_R1176_U9 , P2_U3032 );
nand NAND2_5838 ( P2_U5257 , P2_REG3_REG_13_ , P2_U3152 );
nand NAND2_5839 ( P2_U5258 , P2_U3041 , P2_U3081 );
nand NAND2_5840 ( P2_U5259 , P2_U3039 , P2_U3075 );
nand NAND2_5841 ( P2_U5260 , P2_ADD_609_U63 , P2_U3427 );
nand NAND3_5842 ( P2_U5261 , P2_U5259 , P2_U5258 , P2_U5260 );
nand NAND2_5843 ( P2_U5262 , P2_U3047 , P2_U3976 );
nand NAND2_5844 ( P2_U5263 , P2_U3046 , P2_ADD_609_U63 );
nand NAND2_5845 ( P2_U5264 , P2_U3988 , P2_U5261 );
nand NAND2_5846 ( P2_U5265 , P2_R1176_U97 , P2_U3032 );
nand NAND2_5847 ( P2_U5266 , P2_REG3_REG_20_ , P2_U3152 );
nand NAND2_5848 ( P2_U5267 , P2_U3429 , P2_U3426 );
nand NAND2_5849 ( P2_U5268 , P2_U5267 , P2_U3427 );
nand NAND2_5850 ( P2_U5269 , P2_U3989 , P2_U5268 );
nand NAND2_5851 ( P2_U5270 , P2_U3893 , P2_U3039 );
nand NAND2_5852 ( P2_U5271 , P2_U3448 , P2_U5678 );
nand NAND2_5853 ( P2_U5272 , P2_REG3_REG_0_ , P2_U5269 );
nand NAND2_5854 ( P2_U5273 , P2_R1176_U84 , P2_U3032 );
nand NAND2_5855 ( P2_U5274 , P2_REG3_REG_0_ , P2_U3152 );
nand NAND2_5856 ( P2_U5275 , P2_U3041 , P2_U3084 );
nand NAND2_5857 ( P2_U5276 , P2_U3039 , P2_U3062 );
nand NAND2_5858 ( P2_U5277 , P2_ADD_609_U49 , P2_U3427 );
nand NAND3_5859 ( P2_U5278 , P2_U5276 , P2_U5275 , P2_U5277 );
nand NAND2_5860 ( P2_U5279 , P2_U3477 , P2_U5678 );
nand NAND2_5861 ( P2_U5280 , P2_ADD_609_U49 , P2_U5677 );
nand NAND2_5862 ( P2_U5281 , P2_U3988 , P2_U5278 );
nand NAND2_5863 ( P2_U5282 , P2_R1176_U85 , P2_U3032 );
nand NAND2_5864 ( P2_U5283 , P2_REG3_REG_9_ , P2_U3152 );
nand NAND2_5865 ( P2_U5284 , P2_U3041 , P2_U3064 );
nand NAND2_5866 ( P2_U5285 , P2_U3039 , P2_U3067 );
nand NAND2_5867 ( P2_U5286 , P2_ADD_609_U54 , P2_U3427 );
nand NAND3_5868 ( P2_U5287 , P2_U5285 , P2_U5284 , P2_U5286 );
nand NAND2_5869 ( P2_U5288 , P2_U3462 , P2_U5678 );
nand NAND2_5870 ( P2_U5289 , P2_ADD_609_U54 , P2_U5677 );
nand NAND2_5871 ( P2_U5290 , P2_U3988 , P2_U5287 );
nand NAND2_5872 ( P2_U5291 , P2_R1176_U89 , P2_U3032 );
nand NAND2_5873 ( P2_U5292 , P2_REG3_REG_4_ , P2_U3152 );
nand NAND2_5874 ( P2_U5293 , P2_U3041 , P2_U3066 );
nand NAND2_5875 ( P2_U5294 , P2_U3039 , P2_U3058 );
nand NAND2_5876 ( P2_U5295 , P2_ADD_609_U59 , P2_U3427 );
nand NAND3_5877 ( P2_U5296 , P2_U5295 , P2_U5293 , P2_U5294 );
nand NAND2_5878 ( P2_U5297 , P2_U3047 , P2_U3972 );
nand NAND2_5879 ( P2_U5298 , P2_U3046 , P2_ADD_609_U59 );
nand NAND2_5880 ( P2_U5299 , P2_U3988 , P2_U5296 );
nand NAND2_5881 ( P2_U5300 , P2_R1176_U94 , P2_U3032 );
nand NAND2_5882 ( P2_U5301 , P2_REG3_REG_24_ , P2_U3152 );
nand NAND2_5883 ( P2_U5302 , P2_U3041 , P2_U3073 );
nand NAND2_5884 ( P2_U5303 , P2_U3039 , P2_U3082 );
nand NAND2_5885 ( P2_U5304 , P2_ADD_609_U66 , P2_U3427 );
nand NAND3_5886 ( P2_U5305 , P2_U5303 , P2_U5302 , P2_U5304 );
nand NAND2_5887 ( P2_U5306 , P2_U3501 , P2_U5678 );
nand NAND2_5888 ( P2_U5307 , P2_ADD_609_U66 , P2_U5677 );
nand NAND2_5889 ( P2_U5308 , P2_U3988 , P2_U5305 );
nand NAND2_5890 ( P2_U5309 , P2_R1176_U10 , P2_U3032 );
nand NAND2_5891 ( P2_U5310 , P2_REG3_REG_17_ , P2_U3152 );
nand NAND2_5892 ( P2_U5311 , P2_U3041 , P2_U3060 );
nand NAND2_5893 ( P2_U5312 , P2_U3039 , P2_U3071 );
nand NAND2_5894 ( P2_U5313 , P2_ADD_609_U53 , P2_U3427 );
nand NAND3_5895 ( P2_U5314 , P2_U5312 , P2_U5311 , P2_U5313 );
nand NAND2_5896 ( P2_U5315 , P2_U3465 , P2_U5678 );
nand NAND2_5897 ( P2_U5316 , P2_ADD_609_U53 , P2_U5677 );
nand NAND2_5898 ( P2_U5317 , P2_U3988 , P2_U5314 );
nand NAND2_5899 ( P2_U5318 , P2_R1176_U88 , P2_U3032 );
nand NAND2_5900 ( P2_U5319 , P2_REG3_REG_5_ , P2_U3152 );
nand NAND2_5901 ( P2_U5320 , P2_U3041 , P2_U3074 );
nand NAND2_5902 ( P2_U5321 , P2_U3039 , P2_U3069 );
nand NAND2_5903 ( P2_U5322 , P2_ADD_609_U67 , P2_U3427 );
nand NAND3_5904 ( P2_U5323 , P2_U5321 , P2_U5320 , P2_U5322 );
nand NAND2_5905 ( P2_U5324 , P2_U3498 , P2_U5678 );
nand NAND2_5906 ( P2_U5325 , P2_ADD_609_U67 , P2_U5677 );
nand NAND2_5907 ( P2_U5326 , P2_U3988 , P2_U5323 );
nand NAND2_5908 ( P2_U5327 , P2_R1176_U101 , P2_U3032 );
nand NAND2_5909 ( P2_U5328 , P2_REG3_REG_16_ , P2_U3152 );
nand NAND2_5910 ( P2_U5329 , P2_U3041 , P2_U3065 );
nand NAND2_5911 ( P2_U5330 , P2_U3039 , P2_U3057 );
nand NAND2_5912 ( P2_U5331 , P2_ADD_609_U58 , P2_U3427 );
nand NAND3_5913 ( P2_U5332 , P2_U5331 , P2_U5329 , P2_U5330 );
nand NAND2_5914 ( P2_U5333 , P2_U3047 , P2_U3971 );
nand NAND2_5915 ( P2_U5334 , P2_U3046 , P2_ADD_609_U58 );
nand NAND2_5916 ( P2_U5335 , P2_U3988 , P2_U5332 );
nand NAND2_5917 ( P2_U5336 , P2_R1176_U93 , P2_U3032 );
nand NAND2_5918 ( P2_U5337 , P2_REG3_REG_25_ , P2_U3152 );
nand NAND2_5919 ( P2_U5338 , P2_U3041 , P2_U3063 );
nand NAND2_5920 ( P2_U5339 , P2_U3039 , P2_U3080 );
nand NAND2_5921 ( P2_U5340 , P2_ADD_609_U71 , P2_U3427 );
nand NAND3_5922 ( P2_U5341 , P2_U5339 , P2_U5338 , P2_U5340 );
nand NAND2_5923 ( P2_U5342 , P2_U3486 , P2_U5678 );
nand NAND2_5924 ( P2_U5343 , P2_ADD_609_U71 , P2_U5677 );
nand NAND2_5925 ( P2_U5344 , P2_U3988 , P2_U5341 );
nand NAND2_5926 ( P2_U5345 , P2_R1176_U104 , P2_U3032 );
nand NAND2_5927 ( P2_U5346 , P2_REG3_REG_12_ , P2_U3152 );
nand NAND2_5928 ( P2_U5347 , P2_U3041 , P2_U3076 );
nand NAND2_5929 ( P2_U5348 , P2_U3039 , P2_U3061 );
nand NAND2_5930 ( P2_U5349 , P2_ADD_609_U62 , P2_U3427 );
nand NAND3_5931 ( P2_U5350 , P2_U5348 , P2_U5347 , P2_U5349 );
nand NAND2_5932 ( P2_U5351 , P2_U3047 , P2_U3975 );
nand NAND2_5933 ( P2_U5352 , P2_U3046 , P2_ADD_609_U62 );
nand NAND2_5934 ( P2_U5353 , P2_U3988 , P2_U5350 );
nand NAND2_5935 ( P2_U5354 , P2_R1176_U11 , P2_U3032 );
nand NAND2_5936 ( P2_U5355 , P2_REG3_REG_21_ , P2_U3152 );
nand NAND2_5937 ( P2_U5356 , P2_U3041 , P2_U3077 );
nand NAND2_5938 ( P2_U5357 , P2_U3039 , P2_U3068 );
nand NAND2_5939 ( P2_U5358 , P2_REG3_REG_1_ , P2_U3427 );
nand NAND3_5940 ( P2_U5359 , P2_U5357 , P2_U5356 , P2_U5358 );
nand NAND2_5941 ( P2_U5360 , P2_U3453 , P2_U5678 );
nand NAND2_5942 ( P2_U5361 , P2_REG3_REG_1_ , P2_U5677 );
nand NAND2_5943 ( P2_U5362 , P2_U3988 , P2_U5359 );
nand NAND2_5944 ( P2_U5363 , P2_R1176_U98 , P2_U3032 );
nand NAND2_5945 ( P2_U5364 , P2_REG3_REG_1_ , P2_U3152 );
nand NAND2_5946 ( P2_U5365 , P2_U3041 , P2_U3070 );
nand NAND2_5947 ( P2_U5366 , P2_U3039 , P2_U3083 );
nand NAND2_5948 ( P2_U5367 , P2_ADD_609_U50 , P2_U3427 );
nand NAND3_5949 ( P2_U5368 , P2_U5366 , P2_U5365 , P2_U5367 );
nand NAND2_5950 ( P2_U5369 , P2_U3474 , P2_U5678 );
nand NAND2_5951 ( P2_U5370 , P2_ADD_609_U50 , P2_U5677 );
nand NAND2_5952 ( P2_U5371 , P2_U3988 , P2_U5368 );
nand NAND2_5953 ( P2_U5372 , P2_R1176_U86 , P2_U3032 );
nand NAND2_5954 ( P2_U5373 , P2_REG3_REG_8_ , P2_U3152 );
nand NAND2_5955 ( P2_U5374 , P2_U3041 , P2_U3053 );
nand NAND2_5956 ( P2_U5375 , P2_U3039 , P2_U3055 );
nand NAND2_5957 ( P2_U5376 , P2_ADD_609_U55 , P2_U3427 );
nand NAND3_5958 ( P2_U5377 , P2_U5375 , P2_U5376 , P2_U5374 );
nand NAND2_5959 ( P2_U5378 , P2_U3047 , P2_U3968 );
nand NAND2_5960 ( P2_U5379 , P2_U3046 , P2_ADD_609_U55 );
nand NAND2_5961 ( P2_U5380 , P2_U3988 , P2_U5377 );
nand NAND2_5962 ( P2_U5381 , P2_R1176_U91 , P2_U3032 );
nand NAND2_5963 ( P2_U5382 , P2_REG3_REG_28_ , P2_U3152 );
nand NAND2_5964 ( P2_U5383 , P2_U3041 , P2_U3082 );
nand NAND2_5965 ( P2_U5384 , P2_U3039 , P2_U3076 );
nand NAND2_5966 ( P2_U5385 , P2_ADD_609_U64 , P2_U3427 );
nand NAND3_5967 ( P2_U5386 , P2_U5384 , P2_U5383 , P2_U5385 );
nand NAND2_5968 ( P2_U5387 , P2_U3506 , P2_U5678 );
nand NAND2_5969 ( P2_U5388 , P2_ADD_609_U64 , P2_U5677 );
nand NAND2_5970 ( P2_U5389 , P2_U3988 , P2_U5386 );
nand NAND2_5971 ( P2_U5390 , P2_R1176_U99 , P2_U3032 );
nand NAND2_5972 ( P2_U5391 , P2_REG3_REG_19_ , P2_U3152 );
nand NAND2_5973 ( P2_U5392 , P2_U3041 , P2_U3068 );
nand NAND2_5974 ( P2_U5393 , P2_U3039 , P2_U3060 );
nand NAND2_5975 ( P2_U5394 , P2_ADD_609_U4 , P2_U3427 );
nand NAND3_5976 ( P2_U5395 , P2_U5393 , P2_U5392 , P2_U5394 );
nand NAND2_5977 ( P2_U5396 , P2_U3459 , P2_U5678 );
nand NAND2_5978 ( P2_U5397 , P2_ADD_609_U4 , P2_U5677 );
nand NAND2_5979 ( P2_U5398 , P2_U3988 , P2_U5395 );
nand NAND2_5980 ( P2_U5399 , P2_R1176_U13 , P2_U3032 );
nand NAND2_5981 ( P2_U5400 , P2_REG3_REG_3_ , P2_U3152 );
nand NAND2_5982 ( P2_U5401 , P2_U3041 , P2_U3083 );
nand NAND2_5983 ( P2_U5402 , P2_U3039 , P2_U3063 );
nand NAND2_5984 ( P2_U5403 , P2_ADD_609_U73 , P2_U3427 );
nand NAND3_5985 ( P2_U5404 , P2_U5402 , P2_U5401 , P2_U5403 );
nand NAND2_5986 ( P2_U5405 , P2_U3480 , P2_U5678 );
nand NAND2_5987 ( P2_U5406 , P2_ADD_609_U73 , P2_U5677 );
nand NAND2_5988 ( P2_U5407 , P2_U3988 , P2_U5404 );
nand NAND2_5989 ( P2_U5408 , P2_R1176_U106 , P2_U3032 );
nand NAND2_5990 ( P2_U5409 , P2_REG3_REG_10_ , P2_U3152 );
nand NAND2_5991 ( P2_U5410 , P2_U3041 , P2_U3061 );
nand NAND2_5992 ( P2_U5411 , P2_U3039 , P2_U3065 );
nand NAND2_5993 ( P2_U5412 , P2_ADD_609_U60 , P2_U3427 );
nand NAND3_5994 ( P2_U5413 , P2_U5412 , P2_U5410 , P2_U5411 );
nand NAND2_5995 ( P2_U5414 , P2_U3047 , P2_U3973 );
nand NAND2_5996 ( P2_U5415 , P2_U3046 , P2_ADD_609_U60 );
nand NAND2_5997 ( P2_U5416 , P2_U3988 , P2_U5413 );
nand NAND2_5998 ( P2_U5417 , P2_R1176_U95 , P2_U3032 );
nand NAND2_5999 ( P2_U5418 , P2_REG3_REG_23_ , P2_U3152 );
nand NAND2_6000 ( P2_U5419 , P2_U3041 , P2_U3080 );
nand NAND2_6001 ( P2_U5420 , P2_U3039 , P2_U3074 );
nand NAND2_6002 ( P2_U5421 , P2_ADD_609_U69 , P2_U3427 );
nand NAND3_6003 ( P2_U5422 , P2_U5420 , P2_U5419 , P2_U5421 );
nand NAND2_6004 ( P2_U5423 , P2_U3492 , P2_U5678 );
nand NAND2_6005 ( P2_U5424 , P2_ADD_609_U69 , P2_U5677 );
nand NAND2_6006 ( P2_U5425 , P2_U3988 , P2_U5422 );
nand NAND2_6007 ( P2_U5426 , P2_R1176_U103 , P2_U3032 );
nand NAND2_6008 ( P2_U5427 , P2_REG3_REG_14_ , P2_U3152 );
nand NAND2_6009 ( P2_U5428 , P2_U3041 , P2_U3057 );
nand NAND2_6010 ( P2_U5429 , P2_U3039 , P2_U3054 );
nand NAND2_6011 ( P2_U5430 , P2_ADD_609_U56 , P2_U3427 );
nand NAND3_6012 ( P2_U5431 , P2_U5430 , P2_U5428 , P2_U5429 );
nand NAND2_6013 ( P2_U5432 , P2_U3047 , P2_U3969 );
nand NAND2_6014 ( P2_U5433 , P2_U3046 , P2_ADD_609_U56 );
nand NAND2_6015 ( P2_U5434 , P2_U3988 , P2_U5431 );
nand NAND2_6016 ( P2_U5435 , P2_R1176_U92 , P2_U3032 );
nand NAND2_6017 ( P2_U5436 , P2_REG3_REG_27_ , P2_U3152 );
nand NAND2_6018 ( P2_U5437 , P2_U3041 , P2_U3071 );
nand NAND2_6019 ( P2_U5438 , P2_U3039 , P2_U3084 );
nand NAND2_6020 ( P2_U5439 , P2_ADD_609_U51 , P2_U3427 );
nand NAND3_6021 ( P2_U5440 , P2_U5438 , P2_U5437 , P2_U5439 );
nand NAND2_6022 ( P2_U5441 , P2_U3471 , P2_U5678 );
nand NAND2_6023 ( P2_U5442 , P2_ADD_609_U51 , P2_U5677 );
nand NAND2_6024 ( P2_U5443 , P2_U3988 , P2_U5440 );
nand NAND2_6025 ( P2_U5444 , P2_R1176_U14 , P2_U3032 );
nand NAND2_6026 ( P2_U5445 , P2_REG3_REG_7_ , P2_U3152 );
nand NAND2_6027 ( P2_U5446 , P2_U3967 , P2_U3048 );
nand NAND2_6028 ( P2_U5447 , P2_U3436 , P2_U3909 );
nand NAND3_6029 ( P2_U5448 , P2_U3372 , P2_U3366 , P2_U3904 );
not NOT1_6030 ( P2_U5449 , P2_U3431 );
nand NAND2_6031 ( P2_U5450 , P2_U3584 , P2_U3431 );
nand NAND2_6032 ( P2_U5451 , P2_U5717 , P2_U3083 );
nand NAND2_6033 ( P2_U5452 , P2_U3585 , P2_U3431 );
nand NAND2_6034 ( P2_U5453 , P2_U5717 , P2_U3084 );
nand NAND2_6035 ( P2_U5454 , P2_U3586 , P2_U3431 );
nand NAND2_6036 ( P2_U5455 , P2_U5717 , P2_U3070 );
nand NAND2_6037 ( P2_U5456 , P2_U3587 , P2_U3431 );
nand NAND2_6038 ( P2_U5457 , P2_U5717 , P2_U3071 );
nand NAND2_6039 ( P2_U5458 , P2_U3588 , P2_U3431 );
nand NAND2_6040 ( P2_U5459 , P2_U5717 , P2_U3067 );
nand NAND2_6041 ( P2_U5460 , P2_U3589 , P2_U3431 );
nand NAND2_6042 ( P2_U5461 , P2_U5717 , P2_U3060 );
nand NAND2_6043 ( P2_U5462 , P2_U3591 , P2_U3431 );
nand NAND2_6044 ( P2_U5463 , P2_U5717 , P2_U3056 );
nand NAND2_6045 ( P2_U5464 , P2_U3592 , P2_U3431 );
nand NAND2_6046 ( P2_U5465 , P2_U5717 , P2_U3059 );
nand NAND2_6047 ( P2_U5466 , P2_U3590 , P2_U3431 );
nand NAND2_6048 ( P2_U5467 , P2_U5717 , P2_U3064 );
nand NAND2_6049 ( P2_U5468 , P2_U3594 , P2_U3431 );
nand NAND2_6050 ( P2_U5469 , P2_U5717 , P2_U3055 );
nand NAND2_6051 ( P2_U5470 , P2_U3595 , P2_U3431 );
nand NAND2_6052 ( P2_U5471 , P2_U5717 , P2_U3054 );
nand NAND2_6053 ( P2_U5472 , P2_U3596 , P2_U3431 );
nand NAND2_6054 ( P2_U5473 , P2_U5717 , P2_U3053 );
nand NAND2_6055 ( P2_U5474 , P2_U3597 , P2_U3431 );
nand NAND2_6056 ( P2_U5475 , P2_U5717 , P2_U3057 );
nand NAND2_6057 ( P2_U5476 , P2_U3598 , P2_U3431 );
nand NAND2_6058 ( P2_U5477 , P2_U5717 , P2_U3058 );
nand NAND2_6059 ( P2_U5478 , P2_U3599 , P2_U3431 );
nand NAND2_6060 ( P2_U5479 , P2_U5717 , P2_U3065 );
nand NAND2_6061 ( P2_U5480 , P2_U3600 , P2_U3431 );
nand NAND2_6062 ( P2_U5481 , P2_U5717 , P2_U3066 );
nand NAND2_6063 ( P2_U5482 , P2_U3601 , P2_U3431 );
nand NAND2_6064 ( P2_U5483 , P2_U5717 , P2_U3061 );
nand NAND2_6065 ( P2_U5484 , P2_U3602 , P2_U3431 );
nand NAND2_6066 ( P2_U5485 , P2_U5717 , P2_U3075 );
nand NAND2_6067 ( P2_U5486 , P2_U3603 , P2_U3431 );
nand NAND2_6068 ( P2_U5487 , P2_U5717 , P2_U3076 );
nand NAND2_6069 ( P2_U5488 , P2_U5717 , P2_U3068 );
nand NAND2_6070 ( P2_U5489 , P2_U3605 , P2_U3431 );
nand NAND2_6071 ( P2_U5490 , P2_U5717 , P2_U3081 );
nand NAND2_6072 ( P2_U5491 , P2_U3606 , P2_U3431 );
nand NAND2_6073 ( P2_U5492 , P2_U5717 , P2_U3082 );
nand NAND2_6074 ( P2_U5493 , P2_U3607 , P2_U3431 );
nand NAND2_6075 ( P2_U5494 , P2_U5717 , P2_U3069 );
nand NAND2_6076 ( P2_U5495 , P2_U3608 , P2_U3431 );
nand NAND2_6077 ( P2_U5496 , P2_U5717 , P2_U3073 );
nand NAND2_6078 ( P2_U5497 , P2_U3609 , P2_U3431 );
nand NAND2_6079 ( P2_U5498 , P2_U5717 , P2_U3074 );
nand NAND2_6080 ( P2_U5499 , P2_U3610 , P2_U3431 );
nand NAND2_6081 ( P2_U5500 , P2_U5717 , P2_U3079 );
nand NAND2_6082 ( P2_U5501 , P2_U3611 , P2_U3431 );
nand NAND2_6083 ( P2_U5502 , P2_U5717 , P2_U3080 );
nand NAND2_6084 ( P2_U5503 , P2_U3612 , P2_U3431 );
nand NAND2_6085 ( P2_U5504 , P2_U5717 , P2_U3072 );
nand NAND2_6086 ( P2_U5505 , P2_U3613 , P2_U3431 );
nand NAND2_6087 ( P2_U5506 , P2_U5717 , P2_U3063 );
nand NAND2_6088 ( P2_U5507 , P2_U3614 , P2_U3431 );
nand NAND2_6089 ( P2_U5508 , P2_U5717 , P2_U3062 );
nand NAND2_6090 ( P2_U5509 , P2_U5717 , P2_U3078 );
nand NAND2_6091 ( P2_U5510 , P2_U5717 , P2_U3077 );
nand NAND2_6092 ( P2_U5511 , P2_U5708 , P2_U3445 );
nand NAND2_6093 ( P2_U5512 , P2_U3436 , P2_U5711 );
nand NAND3_6094 ( P2_U5513 , P2_U3368 , P2_U3950 , P2_U3906 );
nand NAND2_6095 ( P2_U5514 , P2_U3953 , P2_U3477 );
nand NAND2_6096 ( P2_U5515 , P2_U5513 , P2_U3083 );
nand NAND2_6097 ( P2_U5516 , P2_U3953 , P2_U3474 );
nand NAND2_6098 ( P2_U5517 , P2_U5513 , P2_U3084 );
nand NAND2_6099 ( P2_U5518 , P2_U3953 , P2_U3471 );
nand NAND2_6100 ( P2_U5519 , P2_U5513 , P2_U3070 );
nand NAND2_6101 ( P2_U5520 , P2_U3953 , P2_U3468 );
nand NAND2_6102 ( P2_U5521 , P2_U5513 , P2_U3071 );
nand NAND2_6103 ( P2_U5522 , P2_U3953 , P2_U3465 );
nand NAND2_6104 ( P2_U5523 , P2_U5513 , P2_U3067 );
nand NAND2_6105 ( P2_U5524 , P2_U3953 , P2_U3462 );
nand NAND2_6106 ( P2_U5525 , P2_U5513 , P2_U3060 );
nand NAND2_6107 ( P2_U5526 , P2_U5513 , P2_U3056 );
nand NAND2_6108 ( P2_U5527 , P2_U3953 , P2_U3977 );
nand NAND2_6109 ( P2_U5528 , P2_U5513 , P2_U3059 );
nand NAND2_6110 ( P2_U5529 , P2_U3953 , P2_U3459 );
nand NAND2_6111 ( P2_U5530 , P2_U5513 , P2_U3064 );
nand NAND2_6112 ( P2_U5531 , P2_U5513 , P2_U3055 );
nand NAND2_6113 ( P2_U5532 , P2_U3953 , P2_U3979 );
nand NAND2_6114 ( P2_U5533 , P2_U5513 , P2_U3054 );
nand NAND2_6115 ( P2_U5534 , P2_U3953 , P2_U3968 );
nand NAND2_6116 ( P2_U5535 , P2_U5513 , P2_U3053 );
nand NAND2_6117 ( P2_U5536 , P2_U3953 , P2_U3969 );
nand NAND2_6118 ( P2_U5537 , P2_U5513 , P2_U3057 );
nand NAND2_6119 ( P2_U5538 , P2_U3953 , P2_U3970 );
nand NAND2_6120 ( P2_U5539 , P2_U5513 , P2_U3058 );
nand NAND2_6121 ( P2_U5540 , P2_U3953 , P2_U3971 );
nand NAND2_6122 ( P2_U5541 , P2_U5513 , P2_U3065 );
nand NAND2_6123 ( P2_U5542 , P2_U3953 , P2_U3972 );
nand NAND2_6124 ( P2_U5543 , P2_U5513 , P2_U3066 );
nand NAND2_6125 ( P2_U5544 , P2_U3953 , P2_U3973 );
nand NAND2_6126 ( P2_U5545 , P2_U5513 , P2_U3061 );
nand NAND2_6127 ( P2_U5546 , P2_U3953 , P2_U3974 );
nand NAND2_6128 ( P2_U5547 , P2_U5513 , P2_U3075 );
nand NAND2_6129 ( P2_U5548 , P2_U3953 , P2_U3975 );
nand NAND2_6130 ( P2_U5549 , P2_U5513 , P2_U3076 );
nand NAND2_6131 ( P2_U5550 , P2_U3953 , P2_U3976 );
nand NAND2_6132 ( P2_U5551 , P2_U3953 , P2_U3456 );
nand NAND2_6133 ( P2_U5552 , P2_U5513 , P2_U3068 );
nand NAND2_6134 ( P2_U5553 , P2_U3953 , P2_U3506 );
nand NAND2_6135 ( P2_U5554 , P2_U5513 , P2_U3081 );
nand NAND2_6136 ( P2_U5555 , P2_U3953 , P2_U3504 );
nand NAND2_6137 ( P2_U5556 , P2_U5513 , P2_U3082 );
nand NAND2_6138 ( P2_U5557 , P2_U3953 , P2_U3501 );
nand NAND2_6139 ( P2_U5558 , P2_U5513 , P2_U3069 );
nand NAND2_6140 ( P2_U5559 , P2_U3953 , P2_U3498 );
nand NAND2_6141 ( P2_U5560 , P2_U5513 , P2_U3073 );
nand NAND2_6142 ( P2_U5561 , P2_U3953 , P2_U3495 );
nand NAND2_6143 ( P2_U5562 , P2_U5513 , P2_U3074 );
nand NAND2_6144 ( P2_U5563 , P2_U3953 , P2_U3492 );
nand NAND2_6145 ( P2_U5564 , P2_U5513 , P2_U3079 );
nand NAND2_6146 ( P2_U5565 , P2_U3953 , P2_U3489 );
nand NAND2_6147 ( P2_U5566 , P2_U5513 , P2_U3080 );
nand NAND2_6148 ( P2_U5567 , P2_U3953 , P2_U3486 );
nand NAND2_6149 ( P2_U5568 , P2_U5513 , P2_U3072 );
nand NAND2_6150 ( P2_U5569 , P2_U3953 , P2_U3483 );
nand NAND2_6151 ( P2_U5570 , P2_U5513 , P2_U3063 );
nand NAND2_6152 ( P2_U5571 , P2_U3953 , P2_U3480 );
nand NAND2_6153 ( P2_U5572 , P2_U5513 , P2_U3062 );
nand NAND2_6154 ( P2_U5573 , P2_U3953 , P2_U3453 );
nand NAND2_6155 ( P2_U5574 , P2_U5513 , P2_U3078 );
nand NAND2_6156 ( P2_U5575 , P2_U3953 , P2_U3448 );
nand NAND2_6157 ( P2_U5576 , P2_U5513 , P2_U3077 );
nand NAND2_6158 ( P2_U5577 , P2_U3477 , P2_U5513 );
nand NAND2_6159 ( P2_U5578 , P2_U3953 , P2_U3083 );
nand NAND2_6160 ( P2_U5579 , P2_U5701 , P2_U3084 );
nand NAND2_6161 ( P2_U5580 , P2_U3474 , P2_U5513 );
nand NAND2_6162 ( P2_U5581 , P2_U3953 , P2_U3084 );
nand NAND2_6163 ( P2_U5582 , P2_U5701 , P2_U3070 );
nand NAND2_6164 ( P2_U5583 , P2_U3471 , P2_U5513 );
nand NAND2_6165 ( P2_U5584 , P2_U3953 , P2_U3070 );
nand NAND2_6166 ( P2_U5585 , P2_U5701 , P2_U3071 );
nand NAND2_6167 ( P2_U5586 , P2_U3468 , P2_U5513 );
nand NAND2_6168 ( P2_U5587 , P2_U3953 , P2_U3071 );
nand NAND2_6169 ( P2_U5588 , P2_U5701 , P2_U3067 );
nand NAND2_6170 ( P2_U5589 , P2_U3465 , P2_U5513 );
nand NAND2_6171 ( P2_U5590 , P2_U3953 , P2_U3067 );
nand NAND2_6172 ( P2_U5591 , P2_U5701 , P2_U3060 );
nand NAND2_6173 ( P2_U5592 , P2_U3462 , P2_U5513 );
nand NAND2_6174 ( P2_U5593 , P2_U3953 , P2_U3060 );
nand NAND2_6175 ( P2_U5594 , P2_U5701 , P2_U3064 );
nand NAND2_6176 ( P2_U5595 , P2_U3977 , P2_U5513 );
nand NAND2_6177 ( P2_U5596 , P2_U3953 , P2_U3056 );
nand NAND2_6178 ( P2_U5597 , P2_U3978 , P2_U5513 );
nand NAND2_6179 ( P2_U5598 , P2_U3953 , P2_U3059 );
nand NAND2_6180 ( P2_U5599 , P2_U3459 , P2_U5513 );
nand NAND2_6181 ( P2_U5600 , P2_U3953 , P2_U3064 );
nand NAND2_6182 ( P2_U5601 , P2_U5701 , P2_U3068 );
nand NAND2_6183 ( P2_U5602 , P2_U3979 , P2_U5513 );
nand NAND2_6184 ( P2_U5603 , P2_U3953 , P2_U3055 );
nand NAND2_6185 ( P2_U5604 , P2_U5701 , P2_U3054 );
nand NAND2_6186 ( P2_U5605 , P2_U3968 , P2_U5513 );
nand NAND2_6187 ( P2_U5606 , P2_U3953 , P2_U3054 );
nand NAND2_6188 ( P2_U5607 , P2_U5701 , P2_U3053 );
nand NAND2_6189 ( P2_U5608 , P2_U3969 , P2_U5513 );
nand NAND2_6190 ( P2_U5609 , P2_U3953 , P2_U3053 );
nand NAND2_6191 ( P2_U5610 , P2_U5701 , P2_U3057 );
nand NAND2_6192 ( P2_U5611 , P2_U3970 , P2_U5513 );
nand NAND2_6193 ( P2_U5612 , P2_U3953 , P2_U3057 );
nand NAND2_6194 ( P2_U5613 , P2_U5701 , P2_U3058 );
nand NAND2_6195 ( P2_U5614 , P2_U3971 , P2_U5513 );
nand NAND2_6196 ( P2_U5615 , P2_U3953 , P2_U3058 );
nand NAND2_6197 ( P2_U5616 , P2_U5701 , P2_U3065 );
nand NAND2_6198 ( P2_U5617 , P2_U3972 , P2_U5513 );
nand NAND2_6199 ( P2_U5618 , P2_U3953 , P2_U3065 );
nand NAND2_6200 ( P2_U5619 , P2_U5701 , P2_U3066 );
nand NAND2_6201 ( P2_U5620 , P2_U3973 , P2_U5513 );
nand NAND2_6202 ( P2_U5621 , P2_U3953 , P2_U3066 );
nand NAND2_6203 ( P2_U5622 , P2_U5701 , P2_U3061 );
nand NAND2_6204 ( P2_U5623 , P2_U3974 , P2_U5513 );
nand NAND2_6205 ( P2_U5624 , P2_U3953 , P2_U3061 );
nand NAND2_6206 ( P2_U5625 , P2_U5701 , P2_U3075 );
nand NAND2_6207 ( P2_U5626 , P2_U3975 , P2_U5513 );
nand NAND2_6208 ( P2_U5627 , P2_U3953 , P2_U3075 );
nand NAND2_6209 ( P2_U5628 , P2_U5701 , P2_U3076 );
nand NAND2_6210 ( P2_U5629 , P2_U3976 , P2_U5513 );
nand NAND2_6211 ( P2_U5630 , P2_U3953 , P2_U3076 );
nand NAND2_6212 ( P2_U5631 , P2_U5701 , P2_U3081 );
nand NAND2_6213 ( P2_U5632 , P2_U3456 , P2_U5513 );
nand NAND2_6214 ( P2_U5633 , P2_U3953 , P2_U3068 );
nand NAND2_6215 ( P2_U5634 , P2_U5701 , P2_U3078 );
nand NAND2_6216 ( P2_U5635 , P2_U3506 , P2_U5513 );
nand NAND2_6217 ( P2_U5636 , P2_U3953 , P2_U3081 );
nand NAND2_6218 ( P2_U5637 , P2_U5701 , P2_U3082 );
nand NAND2_6219 ( P2_U5638 , P2_U3504 , P2_U5513 );
nand NAND2_6220 ( P2_U5639 , P2_U3953 , P2_U3082 );
nand NAND2_6221 ( P2_U5640 , P2_U5701 , P2_U3069 );
nand NAND2_6222 ( P2_U5641 , P2_U3501 , P2_U5513 );
nand NAND2_6223 ( P2_U5642 , P2_U3953 , P2_U3069 );
nand NAND2_6224 ( P2_U5643 , P2_U5701 , P2_U3073 );
nand NAND2_6225 ( P2_U5644 , P2_U3498 , P2_U5513 );
nand NAND2_6226 ( P2_U5645 , P2_U3953 , P2_U3073 );
nand NAND2_6227 ( P2_U5646 , P2_U5701 , P2_U3074 );
nand NAND2_6228 ( P2_U5647 , P2_U3495 , P2_U5513 );
nand NAND2_6229 ( P2_U5648 , P2_U3953 , P2_U3074 );
nand NAND2_6230 ( P2_U5649 , P2_U5701 , P2_U3079 );
nand NAND2_6231 ( P2_U5650 , P2_U3492 , P2_U5513 );
nand NAND2_6232 ( P2_U5651 , P2_U3953 , P2_U3079 );
nand NAND2_6233 ( P2_U5652 , P2_U5701 , P2_U3080 );
nand NAND2_6234 ( P2_U5653 , P2_U3489 , P2_U5513 );
nand NAND2_6235 ( P2_U5654 , P2_U3953 , P2_U3080 );
nand NAND2_6236 ( P2_U5655 , P2_U5701 , P2_U3072 );
nand NAND2_6237 ( P2_U5656 , P2_U3486 , P2_U5513 );
nand NAND2_6238 ( P2_U5657 , P2_U3953 , P2_U3072 );
nand NAND2_6239 ( P2_U5658 , P2_U5701 , P2_U3063 );
nand NAND2_6240 ( P2_U5659 , P2_U3483 , P2_U5513 );
nand NAND2_6241 ( P2_U5660 , P2_U3953 , P2_U3063 );
nand NAND2_6242 ( P2_U5661 , P2_U5701 , P2_U3062 );
nand NAND2_6243 ( P2_U5662 , P2_U3480 , P2_U5513 );
nand NAND2_6244 ( P2_U5663 , P2_U3953 , P2_U3062 );
nand NAND2_6245 ( P2_U5664 , P2_U5701 , P2_U3083 );
nand NAND2_6246 ( P2_U5665 , P2_U3453 , P2_U5513 );
nand NAND2_6247 ( P2_U5666 , P2_U3953 , P2_U3078 );
nand NAND2_6248 ( P2_U5667 , P2_U5701 , P2_U3077 );
nand NAND2_6249 ( P2_U5668 , P2_U3448 , P2_U5513 );
nand NAND2_6250 ( P2_U5669 , P2_U3953 , P2_U3077 );
nand NAND2_6251 ( P2_U5670 , P2_U3436 , P2_STATE_REG );
nand NAND2_6252 ( P2_U5671 , P2_U3886 , P2_U5177 );
nand NAND2_6253 ( P2_U5672 , P2_U5528 , P2_U3413 );
nand NAND2_6254 ( P2_U5673 , P2_U3432 , P2_U5528 );
not NOT1_6255 ( P2_U5674 , P2_U3415 );
nand NAND2_6256 ( P2_U5675 , P2_U3991 , P2_U3427 );
nand NAND2_6257 ( P2_U5676 , P2_U3965 , P2_U3991 );
nand NAND2_6258 ( P2_U5677 , P2_U5675 , P2_U3989 );
nand NAND2_6259 ( P2_U5678 , P2_U5676 , P2_U3990 );
nand NAND2_6260 ( P2_U5679 , P2_U6222 , P2_U5488 );
nand NAND2_6261 ( P2_U5680 , P2_U6245 , P2_U5509 );
nand NAND2_6262 ( P2_U5681 , P2_U6268 , P2_U5510 );
nand NAND2_6263 ( P2_U5682 , P2_U5449 , P2_U5509 );
nand NAND2_6264 ( P2_U5683 , P2_U5449 , P2_U5488 );
nand NAND2_6265 ( P2_U5684 , P2_U5449 , P2_U5510 );
nand NAND2_6266 ( P2_U5685 , P2_U5695 , P2_U5689 );
nand NAND2_6267 ( P2_U5686 , P2_U3436 , P2_U3909 );
nand NAND2_6268 ( P2_U5687 , P2_IR_REG_24_ , P2_U3907 );
nand NAND2_6269 ( P2_U5688 , P2_IR_REG_31_ , P2_SUB_598_U90 );
not NOT1_6270 ( P2_U5689 , P2_U3433 );
nand NAND2_6271 ( P2_U5690 , P2_IR_REG_25_ , P2_U3907 );
nand NAND2_6272 ( P2_U5691 , P2_IR_REG_31_ , P2_SUB_598_U22 );
not NOT1_6273 ( P2_U5692 , P2_U3434 );
nand NAND2_6274 ( P2_U5693 , P2_IR_REG_26_ , P2_U3907 );
nand NAND2_6275 ( P2_U5694 , P2_IR_REG_31_ , P2_SUB_598_U23 );
not NOT1_6276 ( P2_U5695 , P2_U3435 );
nand NAND2_6277 ( P2_U5696 , P2_U5689 , P2_B_REG );
nand NAND2_6278 ( P2_U5697 , P2_U3433 , P2_U3360 );
nand NAND2_6279 ( P2_U5698 , P2_U5697 , P2_U5696 );
nand NAND2_6280 ( P2_U5699 , P2_IR_REG_23_ , P2_U3907 );
nand NAND2_6281 ( P2_U5700 , P2_IR_REG_31_ , P2_SUB_598_U21 );
not NOT1_6282 ( P2_U5701 , P2_U3436 );
nand NAND2_6283 ( P2_U5702 , P2_D_REG_0_ , P2_U3908 );
nand NAND2_6284 ( P2_U5703 , P2_U3986 , P2_U4095 );
nand NAND2_6285 ( P2_U5704 , P2_D_REG_1_ , P2_U3908 );
nand NAND2_6286 ( P2_U5705 , P2_U3986 , P2_U4096 );
nand NAND2_6287 ( P2_U5706 , P2_IR_REG_22_ , P2_U3907 );
nand NAND2_6288 ( P2_U5707 , P2_IR_REG_31_ , P2_SUB_598_U20 );
not NOT1_6289 ( P2_U5708 , P2_U3441 );
nand NAND2_6290 ( P2_U5709 , P2_IR_REG_19_ , P2_U3907 );
nand NAND2_6291 ( P2_U5710 , P2_IR_REG_31_ , P2_SUB_598_U18 );
not NOT1_6292 ( P2_U5711 , P2_U3445 );
nand NAND2_6293 ( P2_U5712 , P2_IR_REG_20_ , P2_U3907 );
nand NAND2_6294 ( P2_U5713 , P2_IR_REG_31_ , P2_SUB_598_U19 );
not NOT1_6295 ( P2_U5714 , P2_U3439 );
nand NAND2_6296 ( P2_U5715 , P2_IR_REG_21_ , P2_U3907 );
nand NAND2_6297 ( P2_U5716 , P2_IR_REG_31_ , P2_SUB_598_U92 );
not NOT1_6298 ( P2_U5717 , P2_U3440 );
nand NAND2_6299 ( P2_U5718 , P2_IR_REG_30_ , P2_U3907 );
nand NAND2_6300 ( P2_U5719 , P2_IR_REG_31_ , P2_SUB_598_U79 );
not NOT1_6301 ( P2_U5720 , P2_U3443 );
nand NAND2_6302 ( P2_U5721 , P2_IR_REG_29_ , P2_U3907 );
nand NAND2_6303 ( P2_U5722 , P2_IR_REG_31_ , P2_SUB_598_U81 );
not NOT1_6304 ( P2_U5723 , P2_U3442 );
nand NAND3_6305 ( P2_U5724 , P2_REG2_REG_1_ , P2_U3443 , P2_U5723 );
nand NAND3_6306 ( P2_U5725 , P2_REG3_REG_1_ , P2_U3443 , P2_U3442 );
nand NAND2_6307 ( P2_U5726 , P2_IR_REG_28_ , P2_U3907 );
nand NAND2_6308 ( P2_U5727 , P2_IR_REG_31_ , P2_SUB_598_U84 );
not NOT1_6309 ( P2_U5728 , P2_U3444 );
nand NAND2_6310 ( P2_U5729 , P2_IR_REG_0_ , P2_U3907 );
nand NAND2_6311 ( P2_U5730 , P2_IR_REG_31_ , P2_IR_REG_0_ );
nand NAND2_6312 ( P2_U5731 , P2_IR_REG_27_ , P2_U3907 );
nand NAND2_6313 ( P2_U5732 , P2_IR_REG_31_ , P2_SUB_598_U87 );
not NOT1_6314 ( P2_U5733 , P2_U3447 );
nand NAND2_6315 ( P2_U5734 , U56 , P2_U3909 );
nand NAND2_6316 ( P2_U5735 , P2_U3964 , P2_U3446 );
not NOT1_6317 ( P2_U5736 , P2_U3448 );
nand NAND2_6318 ( P2_U5737 , P2_U3441 , P2_U5717 );
nand NAND2_6319 ( P2_U5738 , P2_U3439 , P2_U5708 );
nand NAND2_6320 ( P2_U5739 , P2_D_REG_1_ , P2_U4094 );
nand NAND2_6321 ( P2_U5740 , P2_U4096 , P2_U3362 );
not NOT1_6322 ( P2_U5741 , P2_U3450 );
nand NAND2_6323 ( P2_U5742 , P2_U5685 , P2_U3362 );
nand NAND2_6324 ( P2_U5743 , P2_D_REG_0_ , P2_U4094 );
not NOT1_6325 ( P2_U5744 , P2_U3449 );
nand NAND2_6326 ( P2_U5745 , P2_REG0_REG_0_ , P2_U3910 );
nand NAND2_6327 ( P2_U5746 , P2_U3985 , P2_U4145 );
nand NAND3_6328 ( P2_U5747 , P2_REG2_REG_0_ , P2_U3443 , P2_U5723 );
nand NAND3_6329 ( P2_U5748 , P2_REG3_REG_0_ , P2_U3443 , P2_U3442 );
nand NAND2_6330 ( P2_U5749 , P2_IR_REG_1_ , P2_U3907 );
nand NAND2_6331 ( P2_U5750 , P2_IR_REG_31_ , P2_SUB_598_U49 );
nand NAND2_6332 ( P2_U5751 , U45 , P2_U3909 );
nand NAND2_6333 ( P2_U5752 , P2_U3452 , P2_U3964 );
not NOT1_6334 ( P2_U5753 , P2_U3453 );
nand NAND3_6335 ( P2_U5754 , P2_REG2_REG_2_ , P2_U3443 , P2_U5723 );
nand NAND3_6336 ( P2_U5755 , P2_REG3_REG_2_ , P2_U3443 , P2_U3442 );
nand NAND2_6337 ( P2_U5756 , P2_REG0_REG_1_ , P2_U3910 );
nand NAND2_6338 ( P2_U5757 , P2_U3985 , P2_U4165 );
nand NAND2_6339 ( P2_U5758 , P2_IR_REG_2_ , P2_U3907 );
nand NAND2_6340 ( P2_U5759 , P2_IR_REG_31_ , P2_SUB_598_U24 );
nand NAND2_6341 ( P2_U5760 , U34 , P2_U3909 );
nand NAND2_6342 ( P2_U5761 , P2_U3455 , P2_U3964 );
not NOT1_6343 ( P2_U5762 , P2_U3456 );
nand NAND2_6344 ( P2_U5763 , P2_REG0_REG_2_ , P2_U3910 );
nand NAND2_6345 ( P2_U5764 , P2_U3985 , P2_U4184 );
nand NAND2_6346 ( P2_U5765 , P2_IR_REG_3_ , P2_U3907 );
nand NAND2_6347 ( P2_U5766 , P2_IR_REG_31_ , P2_SUB_598_U25 );
nand NAND2_6348 ( P2_U5767 , U31 , P2_U3909 );
nand NAND2_6349 ( P2_U5768 , P2_U3458 , P2_U3964 );
not NOT1_6350 ( P2_U5769 , P2_U3459 );
nand NAND2_6351 ( P2_U5770 , P2_REG0_REG_3_ , P2_U3910 );
nand NAND2_6352 ( P2_U5771 , P2_U3985 , P2_U4203 );
nand NAND2_6353 ( P2_U5772 , P2_IR_REG_4_ , P2_U3907 );
nand NAND2_6354 ( P2_U5773 , P2_IR_REG_31_ , P2_SUB_598_U26 );
nand NAND2_6355 ( P2_U5774 , U30 , P2_U3909 );
nand NAND2_6356 ( P2_U5775 , P2_U3461 , P2_U3964 );
not NOT1_6357 ( P2_U5776 , P2_U3462 );
nand NAND2_6358 ( P2_U5777 , P2_REG0_REG_4_ , P2_U3910 );
nand NAND2_6359 ( P2_U5778 , P2_U3985 , P2_U4222 );
nand NAND2_6360 ( P2_U5779 , P2_IR_REG_5_ , P2_U3907 );
nand NAND2_6361 ( P2_U5780 , P2_IR_REG_31_ , P2_SUB_598_U74 );
nand NAND2_6362 ( P2_U5781 , U29 , P2_U3909 );
nand NAND2_6363 ( P2_U5782 , P2_U3464 , P2_U3964 );
not NOT1_6364 ( P2_U5783 , P2_U3465 );
nand NAND2_6365 ( P2_U5784 , P2_REG0_REG_5_ , P2_U3910 );
nand NAND2_6366 ( P2_U5785 , P2_U3985 , P2_U4241 );
nand NAND2_6367 ( P2_U5786 , P2_IR_REG_6_ , P2_U3907 );
nand NAND2_6368 ( P2_U5787 , P2_IR_REG_31_ , P2_SUB_598_U27 );
nand NAND2_6369 ( P2_U5788 , U28 , P2_U3909 );
nand NAND2_6370 ( P2_U5789 , P2_U3467 , P2_U3964 );
not NOT1_6371 ( P2_U5790 , P2_U3468 );
nand NAND2_6372 ( P2_U5791 , P2_REG0_REG_6_ , P2_U3910 );
nand NAND2_6373 ( P2_U5792 , P2_U3985 , P2_U4260 );
nand NAND2_6374 ( P2_U5793 , P2_IR_REG_7_ , P2_U3907 );
nand NAND2_6375 ( P2_U5794 , P2_IR_REG_31_ , P2_SUB_598_U28 );
nand NAND2_6376 ( P2_U5795 , U27 , P2_U3909 );
nand NAND2_6377 ( P2_U5796 , P2_U3470 , P2_U3964 );
not NOT1_6378 ( P2_U5797 , P2_U3471 );
nand NAND2_6379 ( P2_U5798 , P2_REG0_REG_7_ , P2_U3910 );
nand NAND2_6380 ( P2_U5799 , P2_U3985 , P2_U4279 );
nand NAND2_6381 ( P2_U5800 , P2_IR_REG_8_ , P2_U3907 );
nand NAND2_6382 ( P2_U5801 , P2_IR_REG_31_ , P2_SUB_598_U29 );
nand NAND2_6383 ( P2_U5802 , U26 , P2_U3909 );
nand NAND2_6384 ( P2_U5803 , P2_U3473 , P2_U3964 );
not NOT1_6385 ( P2_U5804 , P2_U3474 );
nand NAND2_6386 ( P2_U5805 , P2_REG0_REG_8_ , P2_U3910 );
nand NAND2_6387 ( P2_U5806 , P2_U3985 , P2_U4298 );
nand NAND2_6388 ( P2_U5807 , P2_IR_REG_9_ , P2_U3907 );
nand NAND2_6389 ( P2_U5808 , P2_IR_REG_31_ , P2_SUB_598_U72 );
nand NAND2_6390 ( P2_U5809 , U25 , P2_U3909 );
nand NAND2_6391 ( P2_U5810 , P2_U3476 , P2_U3964 );
not NOT1_6392 ( P2_U5811 , P2_U3477 );
nand NAND2_6393 ( P2_U5812 , P2_REG0_REG_9_ , P2_U3910 );
nand NAND2_6394 ( P2_U5813 , P2_U3985 , P2_U4317 );
nand NAND2_6395 ( P2_U5814 , P2_IR_REG_10_ , P2_U3907 );
nand NAND2_6396 ( P2_U5815 , P2_IR_REG_31_ , P2_SUB_598_U11 );
nand NAND2_6397 ( P2_U5816 , U55 , P2_U3909 );
nand NAND2_6398 ( P2_U5817 , P2_U3479 , P2_U3964 );
not NOT1_6399 ( P2_U5818 , P2_U3480 );
nand NAND2_6400 ( P2_U5819 , P2_REG0_REG_10_ , P2_U3910 );
nand NAND2_6401 ( P2_U5820 , P2_U3985 , P2_U4336 );
nand NAND2_6402 ( P2_U5821 , P2_IR_REG_11_ , P2_U3907 );
nand NAND2_6403 ( P2_U5822 , P2_IR_REG_31_ , P2_SUB_598_U12 );
nand NAND2_6404 ( P2_U5823 , U54 , P2_U3909 );
nand NAND2_6405 ( P2_U5824 , P2_U3482 , P2_U3964 );
not NOT1_6406 ( P2_U5825 , P2_U3483 );
nand NAND2_6407 ( P2_U5826 , P2_REG0_REG_11_ , P2_U3910 );
nand NAND2_6408 ( P2_U5827 , P2_U3985 , P2_U4355 );
nand NAND2_6409 ( P2_U5828 , P2_IR_REG_12_ , P2_U3907 );
nand NAND2_6410 ( P2_U5829 , P2_IR_REG_31_ , P2_SUB_598_U13 );
nand NAND2_6411 ( P2_U5830 , U53 , P2_U3909 );
nand NAND2_6412 ( P2_U5831 , P2_U3485 , P2_U3964 );
not NOT1_6413 ( P2_U5832 , P2_U3486 );
nand NAND2_6414 ( P2_U5833 , P2_REG0_REG_12_ , P2_U3910 );
nand NAND2_6415 ( P2_U5834 , P2_U3985 , P2_U4374 );
nand NAND2_6416 ( P2_U5835 , P2_IR_REG_13_ , P2_U3907 );
nand NAND2_6417 ( P2_U5836 , P2_IR_REG_31_ , P2_SUB_598_U99 );
nand NAND2_6418 ( P2_U5837 , U52 , P2_U3909 );
nand NAND2_6419 ( P2_U5838 , P2_U3488 , P2_U3964 );
not NOT1_6420 ( P2_U5839 , P2_U3489 );
nand NAND2_6421 ( P2_U5840 , P2_REG0_REG_13_ , P2_U3910 );
nand NAND2_6422 ( P2_U5841 , P2_U3985 , P2_U4393 );
nand NAND2_6423 ( P2_U5842 , P2_IR_REG_14_ , P2_U3907 );
nand NAND2_6424 ( P2_U5843 , P2_IR_REG_31_ , P2_SUB_598_U14 );
nand NAND2_6425 ( P2_U5844 , U51 , P2_U3909 );
nand NAND2_6426 ( P2_U5845 , P2_U3491 , P2_U3964 );
not NOT1_6427 ( P2_U5846 , P2_U3492 );
nand NAND2_6428 ( P2_U5847 , P2_REG0_REG_14_ , P2_U3910 );
nand NAND2_6429 ( P2_U5848 , P2_U3985 , P2_U4412 );
nand NAND2_6430 ( P2_U5849 , P2_IR_REG_15_ , P2_U3907 );
nand NAND2_6431 ( P2_U5850 , P2_IR_REG_31_ , P2_SUB_598_U15 );
nand NAND2_6432 ( P2_U5851 , U50 , P2_U3909 );
nand NAND2_6433 ( P2_U5852 , P2_U3494 , P2_U3964 );
not NOT1_6434 ( P2_U5853 , P2_U3495 );
nand NAND2_6435 ( P2_U5854 , P2_REG0_REG_15_ , P2_U3910 );
nand NAND2_6436 ( P2_U5855 , P2_U3985 , P2_U4431 );
nand NAND2_6437 ( P2_U5856 , P2_IR_REG_16_ , P2_U3907 );
nand NAND2_6438 ( P2_U5857 , P2_IR_REG_31_ , P2_SUB_598_U16 );
nand NAND2_6439 ( P2_U5858 , U49 , P2_U3909 );
nand NAND2_6440 ( P2_U5859 , P2_U3497 , P2_U3964 );
not NOT1_6441 ( P2_U5860 , P2_U3498 );
nand NAND2_6442 ( P2_U5861 , P2_REG0_REG_16_ , P2_U3910 );
nand NAND2_6443 ( P2_U5862 , P2_U3985 , P2_U4450 );
nand NAND2_6444 ( P2_U5863 , P2_IR_REG_17_ , P2_U3907 );
nand NAND2_6445 ( P2_U5864 , P2_IR_REG_31_ , P2_SUB_598_U97 );
nand NAND2_6446 ( P2_U5865 , U48 , P2_U3909 );
nand NAND2_6447 ( P2_U5866 , P2_U3500 , P2_U3964 );
not NOT1_6448 ( P2_U5867 , P2_U3501 );
nand NAND2_6449 ( P2_U5868 , P2_REG0_REG_17_ , P2_U3910 );
nand NAND2_6450 ( P2_U5869 , P2_U3985 , P2_U4469 );
nand NAND2_6451 ( P2_U5870 , P2_IR_REG_18_ , P2_U3907 );
nand NAND2_6452 ( P2_U5871 , P2_IR_REG_31_ , P2_SUB_598_U17 );
nand NAND2_6453 ( P2_U5872 , U47 , P2_U3909 );
nand NAND2_6454 ( P2_U5873 , P2_U3503 , P2_U3964 );
not NOT1_6455 ( P2_U5874 , P2_U3504 );
nand NAND2_6456 ( P2_U5875 , P2_REG0_REG_18_ , P2_U3910 );
nand NAND2_6457 ( P2_U5876 , P2_U3985 , P2_U4488 );
nand NAND2_6458 ( P2_U5877 , U46 , P2_U3909 );
nand NAND2_6459 ( P2_U5878 , P2_U3964 , P2_U3445 );
not NOT1_6460 ( P2_U5879 , P2_U3506 );
nand NAND2_6461 ( P2_U5880 , P2_REG0_REG_19_ , P2_U3910 );
nand NAND2_6462 ( P2_U5881 , P2_U3985 , P2_U4507 );
nand NAND2_6463 ( P2_U5882 , P2_REG0_REG_20_ , P2_U3910 );
nand NAND2_6464 ( P2_U5883 , P2_U3985 , P2_U4526 );
nand NAND2_6465 ( P2_U5884 , P2_REG0_REG_21_ , P2_U3910 );
nand NAND2_6466 ( P2_U5885 , P2_U3985 , P2_U4545 );
nand NAND2_6467 ( P2_U5886 , P2_REG0_REG_22_ , P2_U3910 );
nand NAND2_6468 ( P2_U5887 , P2_U3985 , P2_U4564 );
nand NAND2_6469 ( P2_U5888 , P2_REG0_REG_23_ , P2_U3910 );
nand NAND2_6470 ( P2_U5889 , P2_U3985 , P2_U4583 );
nand NAND2_6471 ( P2_U5890 , P2_REG0_REG_24_ , P2_U3910 );
nand NAND2_6472 ( P2_U5891 , P2_U3985 , P2_U4602 );
nand NAND2_6473 ( P2_U5892 , P2_REG0_REG_25_ , P2_U3910 );
nand NAND2_6474 ( P2_U5893 , P2_U3985 , P2_U4621 );
nand NAND2_6475 ( P2_U5894 , P2_REG0_REG_26_ , P2_U3910 );
nand NAND2_6476 ( P2_U5895 , P2_U3985 , P2_U4640 );
nand NAND2_6477 ( P2_U5896 , P2_REG0_REG_27_ , P2_U3910 );
nand NAND2_6478 ( P2_U5897 , P2_U3985 , P2_U4659 );
nand NAND2_6479 ( P2_U5898 , P2_REG0_REG_28_ , P2_U3910 );
nand NAND2_6480 ( P2_U5899 , P2_U3985 , P2_U4678 );
nand NAND2_6481 ( P2_U5900 , P2_REG0_REG_29_ , P2_U3910 );
nand NAND2_6482 ( P2_U5901 , P2_U3985 , P2_U4698 );
nand NAND2_6483 ( P2_U5902 , P2_REG0_REG_30_ , P2_U3910 );
nand NAND2_6484 ( P2_U5903 , P2_U3985 , P2_U4705 );
nand NAND2_6485 ( P2_U5904 , P2_REG0_REG_31_ , P2_U3910 );
nand NAND2_6486 ( P2_U5905 , P2_U3985 , P2_U4708 );
nand NAND2_6487 ( P2_U5906 , P2_REG1_REG_0_ , P2_U3911 );
nand NAND2_6488 ( P2_U5907 , P2_U3984 , P2_U4145 );
nand NAND2_6489 ( P2_U5908 , P2_REG1_REG_1_ , P2_U3911 );
nand NAND2_6490 ( P2_U5909 , P2_U3984 , P2_U4165 );
nand NAND2_6491 ( P2_U5910 , P2_REG1_REG_2_ , P2_U3911 );
nand NAND2_6492 ( P2_U5911 , P2_U3984 , P2_U4184 );
nand NAND2_6493 ( P2_U5912 , P2_REG1_REG_3_ , P2_U3911 );
nand NAND2_6494 ( P2_U5913 , P2_U3984 , P2_U4203 );
nand NAND2_6495 ( P2_U5914 , P2_REG1_REG_4_ , P2_U3911 );
nand NAND2_6496 ( P2_U5915 , P2_U3984 , P2_U4222 );
nand NAND2_6497 ( P2_U5916 , P2_REG1_REG_5_ , P2_U3911 );
nand NAND2_6498 ( P2_U5917 , P2_U3984 , P2_U4241 );
nand NAND2_6499 ( P2_U5918 , P2_REG1_REG_6_ , P2_U3911 );
nand NAND2_6500 ( P2_U5919 , P2_U3984 , P2_U4260 );
nand NAND2_6501 ( P2_U5920 , P2_REG1_REG_7_ , P2_U3911 );
nand NAND2_6502 ( P2_U5921 , P2_U3984 , P2_U4279 );
nand NAND2_6503 ( P2_U5922 , P2_REG1_REG_8_ , P2_U3911 );
nand NAND2_6504 ( P2_U5923 , P2_U3984 , P2_U4298 );
nand NAND2_6505 ( P2_U5924 , P2_REG1_REG_9_ , P2_U3911 );
nand NAND2_6506 ( P2_U5925 , P2_U3984 , P2_U4317 );
nand NAND2_6507 ( P2_U5926 , P2_REG1_REG_10_ , P2_U3911 );
nand NAND2_6508 ( P2_U5927 , P2_U3984 , P2_U4336 );
nand NAND2_6509 ( P2_U5928 , P2_REG1_REG_11_ , P2_U3911 );
nand NAND2_6510 ( P2_U5929 , P2_U3984 , P2_U4355 );
nand NAND2_6511 ( P2_U5930 , P2_REG1_REG_12_ , P2_U3911 );
nand NAND2_6512 ( P2_U5931 , P2_U3984 , P2_U4374 );
nand NAND2_6513 ( P2_U5932 , P2_REG1_REG_13_ , P2_U3911 );
nand NAND2_6514 ( P2_U5933 , P2_U3984 , P2_U4393 );
nand NAND2_6515 ( P2_U5934 , P2_REG1_REG_14_ , P2_U3911 );
nand NAND2_6516 ( P2_U5935 , P2_U3984 , P2_U4412 );
nand NAND2_6517 ( P2_U5936 , P2_REG1_REG_15_ , P2_U3911 );
nand NAND2_6518 ( P2_U5937 , P2_U3984 , P2_U4431 );
nand NAND2_6519 ( P2_U5938 , P2_REG1_REG_16_ , P2_U3911 );
nand NAND2_6520 ( P2_U5939 , P2_U3984 , P2_U4450 );
nand NAND2_6521 ( P2_U5940 , P2_REG1_REG_17_ , P2_U3911 );
nand NAND2_6522 ( P2_U5941 , P2_U3984 , P2_U4469 );
nand NAND2_6523 ( P2_U5942 , P2_REG1_REG_18_ , P2_U3911 );
nand NAND2_6524 ( P2_U5943 , P2_U3984 , P2_U4488 );
nand NAND2_6525 ( P2_U5944 , P2_REG1_REG_19_ , P2_U3911 );
nand NAND2_6526 ( P2_U5945 , P2_U3984 , P2_U4507 );
nand NAND2_6527 ( P2_U5946 , P2_REG1_REG_20_ , P2_U3911 );
nand NAND2_6528 ( P2_U5947 , P2_U3984 , P2_U4526 );
nand NAND2_6529 ( P2_U5948 , P2_REG1_REG_21_ , P2_U3911 );
nand NAND2_6530 ( P2_U5949 , P2_U3984 , P2_U4545 );
nand NAND2_6531 ( P2_U5950 , P2_REG1_REG_22_ , P2_U3911 );
nand NAND2_6532 ( P2_U5951 , P2_U3984 , P2_U4564 );
nand NAND2_6533 ( P2_U5952 , P2_REG1_REG_23_ , P2_U3911 );
nand NAND2_6534 ( P2_U5953 , P2_U3984 , P2_U4583 );
nand NAND2_6535 ( P2_U5954 , P2_REG1_REG_24_ , P2_U3911 );
nand NAND2_6536 ( P2_U5955 , P2_U3984 , P2_U4602 );
nand NAND2_6537 ( P2_U5956 , P2_REG1_REG_25_ , P2_U3911 );
nand NAND2_6538 ( P2_U5957 , P2_U3984 , P2_U4621 );
nand NAND2_6539 ( P2_U5958 , P2_REG1_REG_26_ , P2_U3911 );
nand NAND2_6540 ( P2_U5959 , P2_U3984 , P2_U4640 );
nand NAND2_6541 ( P2_U5960 , P2_REG1_REG_27_ , P2_U3911 );
nand NAND2_6542 ( P2_U5961 , P2_U3984 , P2_U4659 );
nand NAND2_6543 ( P2_U5962 , P2_REG1_REG_28_ , P2_U3911 );
nand NAND2_6544 ( P2_U5963 , P2_U3984 , P2_U4678 );
nand NAND2_6545 ( P2_U5964 , P2_REG1_REG_29_ , P2_U3911 );
nand NAND2_6546 ( P2_U5965 , P2_U3984 , P2_U4698 );
nand NAND2_6547 ( P2_U5966 , P2_REG1_REG_30_ , P2_U3911 );
nand NAND2_6548 ( P2_U5967 , P2_U3984 , P2_U4705 );
nand NAND2_6549 ( P2_U5968 , P2_REG1_REG_31_ , P2_U3911 );
nand NAND2_6550 ( P2_U5969 , P2_U3984 , P2_U4708 );
nand NAND2_6551 ( P2_U5970 , P2_REG2_REG_0_ , P2_U3417 );
nand NAND2_6552 ( P2_U5971 , P2_U3983 , P2_U3373 );
nand NAND2_6553 ( P2_U5972 , P2_REG2_REG_1_ , P2_U3417 );
nand NAND2_6554 ( P2_U5973 , P2_U3983 , P2_U3374 );
nand NAND2_6555 ( P2_U5974 , P2_REG2_REG_2_ , P2_U3417 );
nand NAND2_6556 ( P2_U5975 , P2_U3983 , P2_U3375 );
nand NAND2_6557 ( P2_U5976 , P2_REG2_REG_3_ , P2_U3417 );
nand NAND2_6558 ( P2_U5977 , P2_U3983 , P2_U3376 );
nand NAND2_6559 ( P2_U5978 , P2_REG2_REG_4_ , P2_U3417 );
nand NAND2_6560 ( P2_U5979 , P2_U3983 , P2_U3377 );
nand NAND2_6561 ( P2_U5980 , P2_REG2_REG_5_ , P2_U3417 );
nand NAND2_6562 ( P2_U5981 , P2_U3983 , P2_U3378 );
nand NAND2_6563 ( P2_U5982 , P2_REG2_REG_6_ , P2_U3417 );
nand NAND2_6564 ( P2_U5983 , P2_U3983 , P2_U3379 );
nand NAND2_6565 ( P2_U5984 , P2_REG2_REG_7_ , P2_U3417 );
nand NAND2_6566 ( P2_U5985 , P2_U3983 , P2_U3380 );
nand NAND2_6567 ( P2_U5986 , P2_REG2_REG_8_ , P2_U3417 );
nand NAND2_6568 ( P2_U5987 , P2_U3983 , P2_U3381 );
nand NAND2_6569 ( P2_U5988 , P2_REG2_REG_9_ , P2_U3417 );
nand NAND2_6570 ( P2_U5989 , P2_U3983 , P2_U3382 );
nand NAND2_6571 ( P2_U5990 , P2_REG2_REG_10_ , P2_U3417 );
nand NAND2_6572 ( P2_U5991 , P2_U3983 , P2_U3383 );
nand NAND2_6573 ( P2_U5992 , P2_REG2_REG_11_ , P2_U3417 );
nand NAND2_6574 ( P2_U5993 , P2_U3983 , P2_U3384 );
nand NAND2_6575 ( P2_U5994 , P2_REG2_REG_12_ , P2_U3417 );
nand NAND2_6576 ( P2_U5995 , P2_U3983 , P2_U3385 );
nand NAND2_6577 ( P2_U5996 , P2_REG2_REG_13_ , P2_U3417 );
nand NAND2_6578 ( P2_U5997 , P2_U3983 , P2_U3386 );
nand NAND2_6579 ( P2_U5998 , P2_REG2_REG_14_ , P2_U3417 );
nand NAND2_6580 ( P2_U5999 , P2_U3983 , P2_U3387 );
nand NAND2_6581 ( P2_U6000 , P2_REG2_REG_15_ , P2_U3417 );
nand NAND2_6582 ( P2_U6001 , P2_U3983 , P2_U3388 );
nand NAND2_6583 ( P2_U6002 , P2_REG2_REG_16_ , P2_U3417 );
nand NAND2_6584 ( P2_U6003 , P2_U3983 , P2_U3389 );
nand NAND2_6585 ( P2_U6004 , P2_REG2_REG_17_ , P2_U3417 );
nand NAND2_6586 ( P2_U6005 , P2_U3983 , P2_U3390 );
nand NAND2_6587 ( P2_U6006 , P2_REG2_REG_18_ , P2_U3417 );
nand NAND2_6588 ( P2_U6007 , P2_U3983 , P2_U3391 );
nand NAND2_6589 ( P2_U6008 , P2_REG2_REG_19_ , P2_U3417 );
nand NAND2_6590 ( P2_U6009 , P2_U3983 , P2_U3392 );
nand NAND2_6591 ( P2_U6010 , P2_REG2_REG_20_ , P2_U3417 );
nand NAND2_6592 ( P2_U6011 , P2_U3983 , P2_U3394 );
nand NAND2_6593 ( P2_U6012 , P2_REG2_REG_21_ , P2_U3417 );
nand NAND2_6594 ( P2_U6013 , P2_U3983 , P2_U3396 );
nand NAND2_6595 ( P2_U6014 , P2_REG2_REG_22_ , P2_U3417 );
nand NAND2_6596 ( P2_U6015 , P2_U3983 , P2_U3398 );
nand NAND2_6597 ( P2_U6016 , P2_REG2_REG_23_ , P2_U3417 );
nand NAND2_6598 ( P2_U6017 , P2_U3983 , P2_U3400 );
nand NAND2_6599 ( P2_U6018 , P2_REG2_REG_24_ , P2_U3417 );
nand NAND2_6600 ( P2_U6019 , P2_U3983 , P2_U3402 );
nand NAND2_6601 ( P2_U6020 , P2_REG2_REG_25_ , P2_U3417 );
nand NAND2_6602 ( P2_U6021 , P2_U3983 , P2_U3404 );
nand NAND2_6603 ( P2_U6022 , P2_REG2_REG_26_ , P2_U3417 );
nand NAND2_6604 ( P2_U6023 , P2_U3983 , P2_U3406 );
nand NAND2_6605 ( P2_U6024 , P2_REG2_REG_27_ , P2_U3417 );
nand NAND2_6606 ( P2_U6025 , P2_U3983 , P2_U3408 );
nand NAND2_6607 ( P2_U6026 , P2_REG2_REG_28_ , P2_U3417 );
nand NAND2_6608 ( P2_U6027 , P2_U3983 , P2_U3410 );
nand NAND2_6609 ( P2_U6028 , P2_REG2_REG_29_ , P2_U3417 );
nand NAND2_6610 ( P2_U6029 , P2_U3983 , P2_U3412 );
nand NAND2_6611 ( P2_U6030 , P2_REG2_REG_30_ , P2_U3417 );
nand NAND2_6612 ( P2_U6031 , P2_U3987 , P2_U3983 );
nand NAND2_6613 ( P2_U6032 , P2_REG2_REG_31_ , P2_U3417 );
nand NAND2_6614 ( P2_U6033 , P2_U3987 , P2_U3983 );
nand NAND2_6615 ( P2_U6034 , P2_DATAO_REG_0_ , P2_U3423 );
nand NAND2_6616 ( P2_U6035 , P2_U3966 , P2_U3077 );
nand NAND2_6617 ( P2_U6036 , P2_DATAO_REG_1_ , P2_U3423 );
nand NAND2_6618 ( P2_U6037 , P2_U3966 , P2_U3078 );
nand NAND2_6619 ( P2_U6038 , P2_DATAO_REG_2_ , P2_U3423 );
nand NAND2_6620 ( P2_U6039 , P2_U3966 , P2_U3068 );
nand NAND2_6621 ( P2_U6040 , P2_DATAO_REG_3_ , P2_U3423 );
nand NAND2_6622 ( P2_U6041 , P2_U3966 , P2_U3064 );
nand NAND2_6623 ( P2_U6042 , P2_DATAO_REG_4_ , P2_U3423 );
nand NAND2_6624 ( P2_U6043 , P2_U3966 , P2_U3060 );
nand NAND2_6625 ( P2_U6044 , P2_DATAO_REG_5_ , P2_U3423 );
nand NAND2_6626 ( P2_U6045 , P2_U3966 , P2_U3067 );
nand NAND2_6627 ( P2_U6046 , P2_DATAO_REG_6_ , P2_U3423 );
nand NAND2_6628 ( P2_U6047 , P2_U3966 , P2_U3071 );
nand NAND2_6629 ( P2_U6048 , P2_DATAO_REG_7_ , P2_U3423 );
nand NAND2_6630 ( P2_U6049 , P2_U3966 , P2_U3070 );
nand NAND2_6631 ( P2_U6050 , P2_DATAO_REG_8_ , P2_U3423 );
nand NAND2_6632 ( P2_U6051 , P2_U3966 , P2_U3084 );
nand NAND2_6633 ( P2_U6052 , P2_DATAO_REG_9_ , P2_U3423 );
nand NAND2_6634 ( P2_U6053 , P2_U3966 , P2_U3083 );
nand NAND2_6635 ( P2_U6054 , P2_DATAO_REG_10_ , P2_U3423 );
nand NAND2_6636 ( P2_U6055 , P2_U3966 , P2_U3062 );
nand NAND2_6637 ( P2_U6056 , P2_DATAO_REG_11_ , P2_U3423 );
nand NAND2_6638 ( P2_U6057 , P2_U3966 , P2_U3063 );
nand NAND2_6639 ( P2_U6058 , P2_DATAO_REG_12_ , P2_U3423 );
nand NAND2_6640 ( P2_U6059 , P2_U3966 , P2_U3072 );
nand NAND2_6641 ( P2_U6060 , P2_DATAO_REG_13_ , P2_U3423 );
nand NAND2_6642 ( P2_U6061 , P2_U3966 , P2_U3080 );
nand NAND2_6643 ( P2_U6062 , P2_DATAO_REG_14_ , P2_U3423 );
nand NAND2_6644 ( P2_U6063 , P2_U3966 , P2_U3079 );
nand NAND2_6645 ( P2_U6064 , P2_DATAO_REG_15_ , P2_U3423 );
nand NAND2_6646 ( P2_U6065 , P2_U3966 , P2_U3074 );
nand NAND2_6647 ( P2_U6066 , P2_DATAO_REG_16_ , P2_U3423 );
nand NAND2_6648 ( P2_U6067 , P2_U3966 , P2_U3073 );
nand NAND2_6649 ( P2_U6068 , P2_DATAO_REG_17_ , P2_U3423 );
nand NAND2_6650 ( P2_U6069 , P2_U3966 , P2_U3069 );
nand NAND2_6651 ( P2_U6070 , P2_DATAO_REG_18_ , P2_U3423 );
nand NAND2_6652 ( P2_U6071 , P2_U3966 , P2_U3082 );
nand NAND2_6653 ( P2_U6072 , P2_DATAO_REG_19_ , P2_U3423 );
nand NAND2_6654 ( P2_U6073 , P2_U3966 , P2_U3081 );
nand NAND2_6655 ( P2_U6074 , P2_DATAO_REG_20_ , P2_U3423 );
nand NAND2_6656 ( P2_U6075 , P2_U3966 , P2_U3076 );
nand NAND2_6657 ( P2_U6076 , P2_DATAO_REG_21_ , P2_U3423 );
nand NAND2_6658 ( P2_U6077 , P2_U3966 , P2_U3075 );
nand NAND2_6659 ( P2_U6078 , P2_DATAO_REG_22_ , P2_U3423 );
nand NAND2_6660 ( P2_U6079 , P2_U3966 , P2_U3061 );
nand NAND2_6661 ( P2_U6080 , P2_DATAO_REG_23_ , P2_U3423 );
nand NAND2_6662 ( P2_U6081 , P2_U3966 , P2_U3066 );
nand NAND2_6663 ( P2_U6082 , P2_DATAO_REG_24_ , P2_U3423 );
nand NAND2_6664 ( P2_U6083 , P2_U3966 , P2_U3065 );
nand NAND2_6665 ( P2_U6084 , P2_DATAO_REG_25_ , P2_U3423 );
nand NAND2_6666 ( P2_U6085 , P2_U3966 , P2_U3058 );
nand NAND2_6667 ( P2_U6086 , P2_DATAO_REG_26_ , P2_U3423 );
nand NAND2_6668 ( P2_U6087 , P2_U3966 , P2_U3057 );
nand NAND2_6669 ( P2_U6088 , P2_DATAO_REG_27_ , P2_U3423 );
nand NAND2_6670 ( P2_U6089 , P2_U3966 , P2_U3053 );
nand NAND2_6671 ( P2_U6090 , P2_DATAO_REG_28_ , P2_U3423 );
nand NAND2_6672 ( P2_U6091 , P2_U3966 , P2_U3054 );
nand NAND2_6673 ( P2_U6092 , P2_DATAO_REG_29_ , P2_U3423 );
nand NAND2_6674 ( P2_U6093 , P2_U3966 , P2_U3055 );
nand NAND2_6675 ( P2_U6094 , P2_DATAO_REG_30_ , P2_U3423 );
nand NAND2_6676 ( P2_U6095 , P2_U3966 , P2_U3059 );
nand NAND2_6677 ( P2_U6096 , P2_DATAO_REG_31_ , P2_U3423 );
nand NAND2_6678 ( P2_U6097 , P2_U3966 , P2_U3056 );
nand NAND2_6679 ( P2_U6098 , P2_U5708 , P2_R1340_U6 );
nand NAND2_6680 ( P2_U6099 , P2_LT_719_U11 , P2_U3441 );
nand NAND2_6681 ( P2_U6100 , P2_U5701 , P2_U3425 );
nand NAND2_6682 ( P2_U6101 , P2_U3441 , P2_U3436 );
nand NAND2_6683 ( P2_U6102 , P2_R1312_U21 , P2_U5169 );
nand NAND3_6684 ( P2_U6103 , P2_U5714 , P2_U5170 , P2_U3945 );
nand NAND2_6685 ( P2_U6104 , P2_U3979 , P2_U3055 );
nand NAND2_6686 ( P2_U6105 , P2_U3411 , P2_U4664 );
nand NAND2_6687 ( P2_U6106 , P2_U6105 , P2_U6104 );
nand NAND2_6688 ( P2_U6107 , P2_U3968 , P2_U3054 );
nand NAND2_6689 ( P2_U6108 , P2_U3409 , P2_U4645 );
nand NAND2_6690 ( P2_U6109 , P2_U6108 , P2_U6107 );
nand NAND2_6691 ( P2_U6110 , P2_U3969 , P2_U3053 );
nand NAND2_6692 ( P2_U6111 , P2_U3407 , P2_U4626 );
nand NAND2_6693 ( P2_U6112 , P2_U6111 , P2_U6110 );
nand NAND2_6694 ( P2_U6113 , P2_U3972 , P2_U3065 );
nand NAND2_6695 ( P2_U6114 , P2_U3401 , P2_U4569 );
nand NAND2_6696 ( P2_U6115 , P2_U6114 , P2_U6113 );
nand NAND2_6697 ( P2_U6116 , P2_U3973 , P2_U3066 );
nand NAND2_6698 ( P2_U6117 , P2_U3399 , P2_U4550 );
nand NAND2_6699 ( P2_U6118 , P2_U6117 , P2_U6116 );
nand NAND2_6700 ( P2_U6119 , P2_U3975 , P2_U3075 );
nand NAND2_6701 ( P2_U6120 , P2_U3395 , P2_U4512 );
nand NAND2_6702 ( P2_U6121 , P2_U6120 , P2_U6119 );
nand NAND2_6703 ( P2_U6122 , P2_U3974 , P2_U3061 );
nand NAND2_6704 ( P2_U6123 , P2_U3397 , P2_U4531 );
nand NAND2_6705 ( P2_U6124 , P2_U6123 , P2_U6122 );
nand NAND2_6706 ( P2_U6125 , P2_U3971 , P2_U3058 );
nand NAND2_6707 ( P2_U6126 , P2_U3403 , P2_U4588 );
nand NAND2_6708 ( P2_U6127 , P2_U6126 , P2_U6125 );
nand NAND2_6709 ( P2_U6128 , P2_U3970 , P2_U3057 );
nand NAND2_6710 ( P2_U6129 , P2_U3405 , P2_U4607 );
nand NAND2_6711 ( P2_U6130 , P2_U6129 , P2_U6128 );
nand NAND2_6712 ( P2_U6131 , P2_U3978 , P2_U3059 );
nand NAND2_6713 ( P2_U6132 , P2_U3413 , P2_U4682 );
nand NAND2_6714 ( P2_U6133 , P2_U6132 , P2_U6131 );
nand NAND2_6715 ( P2_U6134 , P2_U3977 , P2_U3056 );
nand NAND2_6716 ( P2_U6135 , P2_U3414 , P2_U4702 );
nand NAND2_6717 ( P2_U6136 , P2_U6135 , P2_U6134 );
nand NAND2_6718 ( P2_U6137 , P2_U5867 , P2_U4436 );
nand NAND2_6719 ( P2_U6138 , P2_U3501 , P2_U3069 );
nand NAND2_6720 ( P2_U6139 , P2_U6138 , P2_U6137 );
nand NAND2_6721 ( P2_U6140 , P2_U5846 , P2_U4379 );
nand NAND2_6722 ( P2_U6141 , P2_U3492 , P2_U3079 );
nand NAND2_6723 ( P2_U6142 , P2_U6141 , P2_U6140 );
nand NAND2_6724 ( P2_U6143 , P2_U5753 , P2_U4130 );
nand NAND2_6725 ( P2_U6144 , P2_U3453 , P2_U3078 );
nand NAND2_6726 ( P2_U6145 , P2_U6144 , P2_U6143 );
nand NAND2_6727 ( P2_U6146 , P2_U5736 , P2_U4151 );
nand NAND2_6728 ( P2_U6147 , P2_U3448 , P2_U3077 );
nand NAND2_6729 ( P2_U6148 , P2_U6147 , P2_U6146 );
nand NAND2_6730 ( P2_U6149 , P2_U5853 , P2_U4398 );
nand NAND2_6731 ( P2_U6150 , P2_U3495 , P2_U3074 );
nand NAND2_6732 ( P2_U6151 , P2_U6150 , P2_U6149 );
nand NAND2_6733 ( P2_U6152 , P2_U5804 , P2_U4265 );
nand NAND2_6734 ( P2_U6153 , P2_U3474 , P2_U3084 );
nand NAND2_6735 ( P2_U6154 , P2_U6153 , P2_U6152 );
nand NAND2_6736 ( P2_U6155 , P2_U5811 , P2_U4284 );
nand NAND2_6737 ( P2_U6156 , P2_U3477 , P2_U3083 );
nand NAND2_6738 ( P2_U6157 , P2_U6156 , P2_U6155 );
nand NAND2_6739 ( P2_U6158 , P2_U5839 , P2_U4360 );
nand NAND2_6740 ( P2_U6159 , P2_U3489 , P2_U3080 );
nand NAND2_6741 ( P2_U6160 , P2_U6159 , P2_U6158 );
nand NAND2_6742 ( P2_U6161 , P2_U5860 , P2_U4417 );
nand NAND2_6743 ( P2_U6162 , P2_U3498 , P2_U3073 );
nand NAND2_6744 ( P2_U6163 , P2_U6162 , P2_U6161 );
nand NAND2_6745 ( P2_U6164 , P2_U5790 , P2_U4227 );
nand NAND2_6746 ( P2_U6165 , P2_U3468 , P2_U3071 );
nand NAND2_6747 ( P2_U6166 , P2_U6165 , P2_U6164 );
nand NAND2_6748 ( P2_U6167 , P2_U5797 , P2_U4246 );
nand NAND2_6749 ( P2_U6168 , P2_U3471 , P2_U3070 );
nand NAND2_6750 ( P2_U6169 , P2_U6168 , P2_U6167 );
nand NAND2_6751 ( P2_U6170 , P2_U5832 , P2_U4341 );
nand NAND2_6752 ( P2_U6171 , P2_U3486 , P2_U3072 );
nand NAND2_6753 ( P2_U6172 , P2_U6171 , P2_U6170 );
nand NAND2_6754 ( P2_U6173 , P2_U5783 , P2_U4208 );
nand NAND2_6755 ( P2_U6174 , P2_U3465 , P2_U3067 );
nand NAND2_6756 ( P2_U6175 , P2_U6174 , P2_U6173 );
nand NAND2_6757 ( P2_U6176 , P2_U5769 , P2_U4170 );
nand NAND2_6758 ( P2_U6177 , P2_U3459 , P2_U3064 );
nand NAND2_6759 ( P2_U6178 , P2_U6177 , P2_U6176 );
nand NAND2_6760 ( P2_U6179 , P2_U5762 , P2_U4148 );
nand NAND2_6761 ( P2_U6180 , P2_U3456 , P2_U3068 );
nand NAND2_6762 ( P2_U6181 , P2_U6180 , P2_U6179 );
nand NAND2_6763 ( P2_U6182 , P2_U5874 , P2_U4455 );
nand NAND2_6764 ( P2_U6183 , P2_U3504 , P2_U3082 );
nand NAND2_6765 ( P2_U6184 , P2_U6183 , P2_U6182 );
nand NAND2_6766 ( P2_U6185 , P2_U5879 , P2_U4474 );
nand NAND2_6767 ( P2_U6186 , P2_U3506 , P2_U3081 );
nand NAND2_6768 ( P2_U6187 , P2_U6186 , P2_U6185 );
nand NAND2_6769 ( P2_U6188 , P2_U5776 , P2_U4189 );
nand NAND2_6770 ( P2_U6189 , P2_U3462 , P2_U3060 );
nand NAND2_6771 ( P2_U6190 , P2_U6189 , P2_U6188 );
nand NAND2_6772 ( P2_U6191 , P2_U5825 , P2_U4322 );
nand NAND2_6773 ( P2_U6192 , P2_U3483 , P2_U3063 );
nand NAND2_6774 ( P2_U6193 , P2_U6192 , P2_U6191 );
nand NAND2_6775 ( P2_U6194 , P2_U5818 , P2_U4303 );
nand NAND2_6776 ( P2_U6195 , P2_U3480 , P2_U3062 );
nand NAND2_6777 ( P2_U6196 , P2_U6195 , P2_U6194 );
nand NAND2_6778 ( P2_U6197 , P2_U3976 , P2_U3076 );
nand NAND2_6779 ( P2_U6198 , P2_U3393 , P2_U4493 );
nand NAND2_6780 ( P2_U6199 , P2_U6198 , P2_U6197 );
nand NAND2_6781 ( P2_U6200 , P2_U3019 , P2_U3947 );
nand NAND2_6782 ( P2_U6201 , P2_U5168 , P2_U3962 );
nand NAND2_6783 ( P2_U6202 , P2_U3083 , P2_R1299_U6 );
nand NAND2_6784 ( P2_U6203 , P2_U3083 , P2_U3948 );
nand NAND2_6785 ( P2_U6204 , P2_U3084 , P2_R1299_U6 );
nand NAND2_6786 ( P2_U6205 , P2_U3084 , P2_U3948 );
nand NAND2_6787 ( P2_U6206 , P2_U3070 , P2_R1299_U6 );
nand NAND2_6788 ( P2_U6207 , P2_U3070 , P2_U3948 );
nand NAND2_6789 ( P2_U6208 , P2_U3071 , P2_R1299_U6 );
nand NAND2_6790 ( P2_U6209 , P2_U3071 , P2_U3948 );
nand NAND2_6791 ( P2_U6210 , P2_U3067 , P2_R1299_U6 );
nand NAND2_6792 ( P2_U6211 , P2_U3067 , P2_U3948 );
nand NAND2_6793 ( P2_U6212 , P2_U3060 , P2_R1299_U6 );
nand NAND2_6794 ( P2_U6213 , P2_U3060 , P2_U3948 );
nand NAND2_6795 ( P2_U6214 , P2_U3064 , P2_R1299_U6 );
nand NAND2_6796 ( P2_U6215 , P2_U3064 , P2_U3948 );
nand NAND2_6797 ( P2_U6216 , P2_R1335_U8 , P2_R1299_U6 );
nand NAND2_6798 ( P2_U6217 , P2_U3056 , P2_U3948 );
nand NAND2_6799 ( P2_U6218 , P2_R1335_U6 , P2_R1299_U6 );
nand NAND2_6800 ( P2_U6219 , P2_U3059 , P2_U3948 );
nand NAND2_6801 ( P2_U6220 , P2_U3068 , P2_R1299_U6 );
nand NAND2_6802 ( P2_U6221 , P2_U3068 , P2_U3948 );
not NOT1_6803 ( P2_U6222 , P2_U3593 );
nand NAND2_6804 ( P2_U6223 , P2_U3055 , P2_R1299_U6 );
nand NAND2_6805 ( P2_U6224 , P2_U3055 , P2_U3948 );
nand NAND2_6806 ( P2_U6225 , P2_U3054 , P2_R1299_U6 );
nand NAND2_6807 ( P2_U6226 , P2_U3054 , P2_U3948 );
nand NAND2_6808 ( P2_U6227 , P2_U3053 , P2_R1299_U6 );
nand NAND2_6809 ( P2_U6228 , P2_U3053 , P2_U3948 );
nand NAND2_6810 ( P2_U6229 , P2_U3057 , P2_R1299_U6 );
nand NAND2_6811 ( P2_U6230 , P2_U3057 , P2_U3948 );
nand NAND2_6812 ( P2_U6231 , P2_U3058 , P2_R1299_U6 );
nand NAND2_6813 ( P2_U6232 , P2_U3058 , P2_U3948 );
nand NAND2_6814 ( P2_U6233 , P2_U3065 , P2_R1299_U6 );
nand NAND2_6815 ( P2_U6234 , P2_U3065 , P2_U3948 );
nand NAND2_6816 ( P2_U6235 , P2_U3066 , P2_R1299_U6 );
nand NAND2_6817 ( P2_U6236 , P2_U3066 , P2_U3948 );
nand NAND2_6818 ( P2_U6237 , P2_U3061 , P2_R1299_U6 );
nand NAND2_6819 ( P2_U6238 , P2_U3061 , P2_U3948 );
nand NAND2_6820 ( P2_U6239 , P2_U3075 , P2_R1299_U6 );
nand NAND2_6821 ( P2_U6240 , P2_U3075 , P2_U3948 );
nand NAND2_6822 ( P2_U6241 , P2_U3076 , P2_R1299_U6 );
nand NAND2_6823 ( P2_U6242 , P2_U3076 , P2_U3948 );
nand NAND2_6824 ( P2_U6243 , P2_U3078 , P2_R1299_U6 );
nand NAND2_6825 ( P2_U6244 , P2_U3078 , P2_U3948 );
not NOT1_6826 ( P2_U6245 , P2_U3604 );
nand NAND2_6827 ( P2_U6246 , P2_U3081 , P2_R1299_U6 );
nand NAND2_6828 ( P2_U6247 , P2_U3081 , P2_U3948 );
nand NAND2_6829 ( P2_U6248 , P2_U3082 , P2_R1299_U6 );
nand NAND2_6830 ( P2_U6249 , P2_U3082 , P2_U3948 );
nand NAND2_6831 ( P2_U6250 , P2_U3069 , P2_R1299_U6 );
nand NAND2_6832 ( P2_U6251 , P2_U3069 , P2_U3948 );
nand NAND2_6833 ( P2_U6252 , P2_U3073 , P2_R1299_U6 );
nand NAND2_6834 ( P2_U6253 , P2_U3073 , P2_U3948 );
nand NAND2_6835 ( P2_U6254 , P2_U3074 , P2_R1299_U6 );
nand NAND2_6836 ( P2_U6255 , P2_U3074 , P2_U3948 );
nand NAND2_6837 ( P2_U6256 , P2_U3079 , P2_R1299_U6 );
nand NAND2_6838 ( P2_U6257 , P2_U3079 , P2_U3948 );
nand NAND2_6839 ( P2_U6258 , P2_U3080 , P2_R1299_U6 );
nand NAND2_6840 ( P2_U6259 , P2_U3080 , P2_U3948 );
nand NAND2_6841 ( P2_U6260 , P2_U3072 , P2_R1299_U6 );
nand NAND2_6842 ( P2_U6261 , P2_U3072 , P2_U3948 );
nand NAND2_6843 ( P2_U6262 , P2_U3063 , P2_R1299_U6 );
nand NAND2_6844 ( P2_U6263 , P2_U3063 , P2_U3948 );
nand NAND2_6845 ( P2_U6264 , P2_U3062 , P2_R1299_U6 );
nand NAND2_6846 ( P2_U6265 , P2_U3062 , P2_U3948 );
nand NAND2_6847 ( P2_U6266 , P2_U3077 , P2_R1299_U6 );
nand NAND2_6848 ( P2_U6267 , P2_U3077 , P2_U3948 );
not NOT1_6849 ( P2_U6268 , P2_U3615 );
nand NAND2_6850 ( P2_U6269 , P2_U3445 , P2_U5717 );
nand NAND2_6851 ( P2_U6270 , P2_U3440 , P2_U3439 );
nand NAND2_6852 ( P2_R1113_U438 , P2_R1113_U274 , P2_R1113_U437 );
not NOT1_6853 ( P2_R1113_U437 , P2_R1113_U138 );
nand NAND2_6854 ( P2_R1113_U436 , P2_U3081 , P2_R1113_U65 );
nand NAND2_6855 ( P2_R1113_U435 , P2_U3506 , P2_R1113_U66 );
nand NAND2_6856 ( P2_R1113_U434 , P2_R1113_U137 , P2_R1113_U166 );
nand NAND2_6857 ( P2_R1113_U433 , P2_R1113_U194 , P2_R1113_U432 );
not NOT1_6858 ( P2_R1113_U432 , P2_R1113_U137 );
nand NAND2_6859 ( P2_R1113_U431 , P2_U3078 , P2_R1113_U165 );
nand NAND2_6860 ( P2_R1113_U430 , P2_U3453 , P2_R1113_U24 );
nand NAND2_6861 ( P2_R1113_U429 , P2_R1113_U136 , P2_R1113_U164 );
nand NAND2_6862 ( P2_R1113_U428 , P2_R1113_U278 , P2_R1113_U427 );
not NOT1_6863 ( P2_R1113_U427 , P2_R1113_U136 );
nand NAND2_6864 ( P2_R1113_U426 , P2_U3076 , P2_R1113_U67 );
nand NAND2_6865 ( P2_R1113_U425 , P2_U3976 , P2_R1113_U68 );
nand NAND2_6866 ( P2_R1113_U424 , P2_R1113_U282 , P2_R1113_U162 );
nand NAND2_6867 ( P2_R1113_U423 , P2_R1113_U324 , P2_R1113_U163 );
nand NAND2_6868 ( P2_R1113_U422 , P2_U3075 , P2_R1113_U70 );
nand NAND2_6869 ( P2_R1113_U421 , P2_U3975 , P2_R1113_U73 );
nand NAND2_6870 ( P2_R1113_U420 , P2_R1113_U161 , P2_R1113_U315 );
nand NAND2_6871 ( P2_R1113_U419 , P2_R1113_U323 , P2_R1113_U86 );
not NOT1_6872 ( LT_1079_U6 , P1_ADDR_REG_19_ );
and AND2_6873 ( ADD_1071_U4 , ADD_1071_U159 , ADD_1071_U155 );
nand NAND3_6874 ( ADD_1071_U5 , ADD_1071_U221 , ADD_1071_U220 , ADD_1071_U160 );
not NOT1_6875 ( ADD_1071_U6 , P1_ADDR_REG_0_ );
not NOT1_6876 ( ADD_1071_U7 , P2_ADDR_REG_0_ );
not NOT1_6877 ( ADD_1071_U8 , P2_ADDR_REG_1_ );
nand NAND2_6878 ( ADD_1071_U9 , P2_ADDR_REG_0_ , P1_ADDR_REG_0_ );
not NOT1_6879 ( ADD_1071_U10 , P1_ADDR_REG_1_ );
not NOT1_6880 ( ADD_1071_U11 , P1_ADDR_REG_2_ );
not NOT1_6881 ( ADD_1071_U12 , P2_ADDR_REG_2_ );
not NOT1_6882 ( ADD_1071_U13 , P1_ADDR_REG_3_ );
not NOT1_6883 ( ADD_1071_U14 , P2_ADDR_REG_3_ );
not NOT1_6884 ( ADD_1071_U15 , P1_ADDR_REG_4_ );
not NOT1_6885 ( ADD_1071_U16 , P2_ADDR_REG_4_ );
not NOT1_6886 ( ADD_1071_U17 , P1_ADDR_REG_5_ );
not NOT1_6887 ( ADD_1071_U18 , P2_ADDR_REG_5_ );
not NOT1_6888 ( ADD_1071_U19 , P1_ADDR_REG_6_ );
not NOT1_6889 ( ADD_1071_U20 , P2_ADDR_REG_6_ );
not NOT1_6890 ( ADD_1071_U21 , P1_ADDR_REG_7_ );
not NOT1_6891 ( ADD_1071_U22 , P2_ADDR_REG_7_ );
not NOT1_6892 ( ADD_1071_U23 , P1_ADDR_REG_8_ );
not NOT1_6893 ( ADD_1071_U24 , P2_ADDR_REG_8_ );
not NOT1_6894 ( ADD_1071_U25 , P2_ADDR_REG_9_ );
not NOT1_6895 ( ADD_1071_U26 , P1_ADDR_REG_9_ );
not NOT1_6896 ( ADD_1071_U27 , P1_ADDR_REG_10_ );
not NOT1_6897 ( ADD_1071_U28 , P2_ADDR_REG_10_ );
not NOT1_6898 ( ADD_1071_U29 , P1_ADDR_REG_11_ );
not NOT1_6899 ( ADD_1071_U30 , P2_ADDR_REG_11_ );
not NOT1_6900 ( ADD_1071_U31 , P1_ADDR_REG_12_ );
not NOT1_6901 ( ADD_1071_U32 , P2_ADDR_REG_12_ );
not NOT1_6902 ( ADD_1071_U33 , P1_ADDR_REG_13_ );
not NOT1_6903 ( ADD_1071_U34 , P2_ADDR_REG_13_ );
not NOT1_6904 ( ADD_1071_U35 , P1_ADDR_REG_14_ );
not NOT1_6905 ( ADD_1071_U36 , P2_ADDR_REG_14_ );
not NOT1_6906 ( ADD_1071_U37 , P1_ADDR_REG_15_ );
not NOT1_6907 ( ADD_1071_U38 , P2_ADDR_REG_15_ );
not NOT1_6908 ( ADD_1071_U39 , P1_ADDR_REG_16_ );
not NOT1_6909 ( ADD_1071_U40 , P2_ADDR_REG_16_ );
not NOT1_6910 ( ADD_1071_U41 , P1_ADDR_REG_17_ );
not NOT1_6911 ( ADD_1071_U42 , P2_ADDR_REG_17_ );
not NOT1_6912 ( ADD_1071_U43 , P1_ADDR_REG_18_ );
not NOT1_6913 ( ADD_1071_U44 , P2_ADDR_REG_18_ );
nand NAND2_6914 ( ADD_1071_U45 , ADD_1071_U150 , ADD_1071_U149 );
nand NAND2_6915 ( ADD_1071_U46 , ADD_1071_U291 , ADD_1071_U290 );
nand NAND2_6916 ( ADD_1071_U47 , ADD_1071_U167 , ADD_1071_U166 );
nand NAND2_6917 ( ADD_1071_U48 , ADD_1071_U174 , ADD_1071_U173 );
nand NAND2_6918 ( ADD_1071_U49 , ADD_1071_U181 , ADD_1071_U180 );
nand NAND2_6919 ( ADD_1071_U50 , ADD_1071_U188 , ADD_1071_U187 );
nand NAND2_6920 ( ADD_1071_U51 , ADD_1071_U195 , ADD_1071_U194 );
nand NAND2_6921 ( ADD_1071_U52 , ADD_1071_U202 , ADD_1071_U201 );
nand NAND2_6922 ( ADD_1071_U53 , ADD_1071_U209 , ADD_1071_U208 );
nand NAND2_6923 ( ADD_1071_U54 , ADD_1071_U216 , ADD_1071_U215 );
nand NAND2_6924 ( ADD_1071_U55 , ADD_1071_U233 , ADD_1071_U232 );
nand NAND2_6925 ( ADD_1071_U56 , ADD_1071_U240 , ADD_1071_U239 );
nand NAND2_6926 ( ADD_1071_U57 , ADD_1071_U247 , ADD_1071_U246 );
nand NAND2_6927 ( ADD_1071_U58 , ADD_1071_U254 , ADD_1071_U253 );
nand NAND2_6928 ( ADD_1071_U59 , ADD_1071_U261 , ADD_1071_U260 );
nand NAND2_6929 ( ADD_1071_U60 , ADD_1071_U268 , ADD_1071_U267 );
nand NAND2_6930 ( ADD_1071_U61 , ADD_1071_U275 , ADD_1071_U274 );
nand NAND2_6931 ( ADD_1071_U62 , ADD_1071_U282 , ADD_1071_U281 );
nand NAND2_6932 ( ADD_1071_U63 , ADD_1071_U289 , ADD_1071_U288 );
nand NAND2_6933 ( ADD_1071_U64 , ADD_1071_U114 , ADD_1071_U113 );
nand NAND2_6934 ( ADD_1071_U65 , ADD_1071_U110 , ADD_1071_U109 );
nand NAND2_6935 ( ADD_1071_U66 , ADD_1071_U106 , ADD_1071_U105 );
nand NAND2_6936 ( ADD_1071_U67 , ADD_1071_U102 , ADD_1071_U101 );
nand NAND2_6937 ( ADD_1071_U68 , ADD_1071_U98 , ADD_1071_U97 );
nand NAND2_6938 ( ADD_1071_U69 , ADD_1071_U94 , ADD_1071_U93 );
nand NAND2_6939 ( ADD_1071_U70 , ADD_1071_U90 , ADD_1071_U89 );
nand NAND2_6940 ( ADD_1071_U71 , ADD_1071_U72 , ADD_1071_U86 );
nand NAND2_6941 ( ADD_1071_U72 , P1_ADDR_REG_1_ , ADD_1071_U84 );
not NOT1_6942 ( ADD_1071_U73 , P2_ADDR_REG_19_ );
not NOT1_6943 ( ADD_1071_U74 , P1_ADDR_REG_19_ );
nand NAND2_6944 ( ADD_1071_U75 , ADD_1071_U146 , ADD_1071_U145 );
nand NAND2_6945 ( ADD_1071_U76 , ADD_1071_U142 , ADD_1071_U141 );
nand NAND2_6946 ( ADD_1071_U77 , ADD_1071_U138 , ADD_1071_U137 );
nand NAND2_6947 ( ADD_1071_U78 , ADD_1071_U134 , ADD_1071_U133 );
nand NAND2_6948 ( ADD_1071_U79 , ADD_1071_U130 , ADD_1071_U129 );
nand NAND2_6949 ( ADD_1071_U80 , ADD_1071_U126 , ADD_1071_U125 );
nand NAND2_6950 ( ADD_1071_U81 , ADD_1071_U122 , ADD_1071_U121 );
nand NAND2_6951 ( ADD_1071_U82 , ADD_1071_U118 , ADD_1071_U117 );
not NOT1_6952 ( ADD_1071_U83 , ADD_1071_U72 );
not NOT1_6953 ( ADD_1071_U84 , ADD_1071_U9 );
nand NAND2_6954 ( ADD_1071_U85 , ADD_1071_U10 , ADD_1071_U9 );
nand NAND2_6955 ( ADD_1071_U86 , P2_ADDR_REG_1_ , ADD_1071_U85 );
not NOT1_6956 ( ADD_1071_U87 , ADD_1071_U71 );
or OR2_6957 ( ADD_1071_U88 , P1_ADDR_REG_2_ , P2_ADDR_REG_2_ );
nand NAND2_6958 ( ADD_1071_U89 , ADD_1071_U88 , ADD_1071_U71 );
nand NAND2_6959 ( ADD_1071_U90 , P2_ADDR_REG_2_ , P1_ADDR_REG_2_ );
not NOT1_6960 ( ADD_1071_U91 , ADD_1071_U70 );
or OR2_6961 ( ADD_1071_U92 , P1_ADDR_REG_3_ , P2_ADDR_REG_3_ );
nand NAND2_6962 ( ADD_1071_U93 , ADD_1071_U92 , ADD_1071_U70 );
nand NAND2_6963 ( ADD_1071_U94 , P2_ADDR_REG_3_ , P1_ADDR_REG_3_ );
not NOT1_6964 ( ADD_1071_U95 , ADD_1071_U69 );
or OR2_6965 ( ADD_1071_U96 , P1_ADDR_REG_4_ , P2_ADDR_REG_4_ );
nand NAND2_6966 ( ADD_1071_U97 , ADD_1071_U96 , ADD_1071_U69 );
nand NAND2_6967 ( ADD_1071_U98 , P2_ADDR_REG_4_ , P1_ADDR_REG_4_ );
not NOT1_6968 ( ADD_1071_U99 , ADD_1071_U68 );
or OR2_6969 ( ADD_1071_U100 , P1_ADDR_REG_5_ , P2_ADDR_REG_5_ );
nand NAND2_6970 ( ADD_1071_U101 , ADD_1071_U100 , ADD_1071_U68 );
nand NAND2_6971 ( ADD_1071_U102 , P2_ADDR_REG_5_ , P1_ADDR_REG_5_ );
not NOT1_6972 ( ADD_1071_U103 , ADD_1071_U67 );
or OR2_6973 ( ADD_1071_U104 , P1_ADDR_REG_6_ , P2_ADDR_REG_6_ );
nand NAND2_6974 ( ADD_1071_U105 , ADD_1071_U104 , ADD_1071_U67 );
nand NAND2_6975 ( ADD_1071_U106 , P2_ADDR_REG_6_ , P1_ADDR_REG_6_ );
not NOT1_6976 ( ADD_1071_U107 , ADD_1071_U66 );
or OR2_6977 ( ADD_1071_U108 , P1_ADDR_REG_7_ , P2_ADDR_REG_7_ );
nand NAND2_6978 ( ADD_1071_U109 , ADD_1071_U108 , ADD_1071_U66 );
nand NAND2_6979 ( ADD_1071_U110 , P2_ADDR_REG_7_ , P1_ADDR_REG_7_ );
not NOT1_6980 ( ADD_1071_U111 , ADD_1071_U65 );
or OR2_6981 ( ADD_1071_U112 , P1_ADDR_REG_8_ , P2_ADDR_REG_8_ );
nand NAND2_6982 ( ADD_1071_U113 , ADD_1071_U112 , ADD_1071_U65 );
nand NAND2_6983 ( ADD_1071_U114 , P2_ADDR_REG_8_ , P1_ADDR_REG_8_ );
not NOT1_6984 ( ADD_1071_U115 , ADD_1071_U64 );
or OR2_6985 ( ADD_1071_U116 , P1_ADDR_REG_9_ , P2_ADDR_REG_9_ );
nand NAND2_6986 ( ADD_1071_U117 , ADD_1071_U116 , ADD_1071_U64 );
nand NAND2_6987 ( ADD_1071_U118 , P1_ADDR_REG_9_ , P2_ADDR_REG_9_ );
not NOT1_6988 ( ADD_1071_U119 , ADD_1071_U82 );
or OR2_6989 ( ADD_1071_U120 , P1_ADDR_REG_10_ , P2_ADDR_REG_10_ );
nand NAND2_6990 ( ADD_1071_U121 , ADD_1071_U120 , ADD_1071_U82 );
nand NAND2_6991 ( ADD_1071_U122 , P2_ADDR_REG_10_ , P1_ADDR_REG_10_ );
not NOT1_6992 ( ADD_1071_U123 , ADD_1071_U81 );
or OR2_6993 ( ADD_1071_U124 , P1_ADDR_REG_11_ , P2_ADDR_REG_11_ );
nand NAND2_6994 ( ADD_1071_U125 , ADD_1071_U124 , ADD_1071_U81 );
nand NAND2_6995 ( ADD_1071_U126 , P2_ADDR_REG_11_ , P1_ADDR_REG_11_ );
not NOT1_6996 ( ADD_1071_U127 , ADD_1071_U80 );
or OR2_6997 ( ADD_1071_U128 , P1_ADDR_REG_12_ , P2_ADDR_REG_12_ );
nand NAND2_6998 ( ADD_1071_U129 , ADD_1071_U128 , ADD_1071_U80 );
nand NAND2_6999 ( ADD_1071_U130 , P2_ADDR_REG_12_ , P1_ADDR_REG_12_ );
not NOT1_7000 ( ADD_1071_U131 , ADD_1071_U79 );
or OR2_7001 ( ADD_1071_U132 , P1_ADDR_REG_13_ , P2_ADDR_REG_13_ );
nand NAND2_7002 ( ADD_1071_U133 , ADD_1071_U132 , ADD_1071_U79 );
nand NAND2_7003 ( ADD_1071_U134 , P2_ADDR_REG_13_ , P1_ADDR_REG_13_ );
not NOT1_7004 ( ADD_1071_U135 , ADD_1071_U78 );
or OR2_7005 ( ADD_1071_U136 , P1_ADDR_REG_14_ , P2_ADDR_REG_14_ );
nand NAND2_7006 ( ADD_1071_U137 , ADD_1071_U136 , ADD_1071_U78 );
nand NAND2_7007 ( ADD_1071_U138 , P2_ADDR_REG_14_ , P1_ADDR_REG_14_ );
not NOT1_7008 ( ADD_1071_U139 , ADD_1071_U77 );
or OR2_7009 ( ADD_1071_U140 , P1_ADDR_REG_15_ , P2_ADDR_REG_15_ );
nand NAND2_7010 ( ADD_1071_U141 , ADD_1071_U140 , ADD_1071_U77 );
nand NAND2_7011 ( ADD_1071_U142 , P2_ADDR_REG_15_ , P1_ADDR_REG_15_ );
not NOT1_7012 ( ADD_1071_U143 , ADD_1071_U76 );
or OR2_7013 ( ADD_1071_U144 , P1_ADDR_REG_16_ , P2_ADDR_REG_16_ );
nand NAND2_7014 ( ADD_1071_U145 , ADD_1071_U144 , ADD_1071_U76 );
nand NAND2_7015 ( ADD_1071_U146 , P2_ADDR_REG_16_ , P1_ADDR_REG_16_ );
not NOT1_7016 ( ADD_1071_U147 , ADD_1071_U75 );
or OR2_7017 ( ADD_1071_U148 , P1_ADDR_REG_17_ , P2_ADDR_REG_17_ );
nand NAND2_7018 ( ADD_1071_U149 , ADD_1071_U148 , ADD_1071_U75 );
nand NAND2_7019 ( ADD_1071_U150 , P2_ADDR_REG_17_ , P1_ADDR_REG_17_ );
not NOT1_7020 ( ADD_1071_U151 , ADD_1071_U45 );
or OR2_7021 ( ADD_1071_U152 , P1_ADDR_REG_18_ , P2_ADDR_REG_18_ );
nand NAND2_7022 ( ADD_1071_U153 , ADD_1071_U152 , ADD_1071_U45 );
nand NAND2_7023 ( ADD_1071_U154 , P2_ADDR_REG_18_ , P1_ADDR_REG_18_ );
nand NAND4_7024 ( ADD_1071_U155 , ADD_1071_U223 , ADD_1071_U222 , ADD_1071_U154 , ADD_1071_U153 );
nand NAND2_7025 ( ADD_1071_U156 , P2_ADDR_REG_18_ , P1_ADDR_REG_18_ );
nand NAND2_7026 ( ADD_1071_U157 , ADD_1071_U151 , ADD_1071_U156 );
or OR2_7027 ( ADD_1071_U158 , P2_ADDR_REG_18_ , P1_ADDR_REG_18_ );
nand NAND3_7028 ( ADD_1071_U159 , ADD_1071_U158 , ADD_1071_U226 , ADD_1071_U157 );
nand NAND2_7029 ( ADD_1071_U160 , ADD_1071_U219 , ADD_1071_U10 );
nand NAND2_7030 ( ADD_1071_U161 , P2_ADDR_REG_9_ , ADD_1071_U26 );
nand NAND2_7031 ( ADD_1071_U162 , P1_ADDR_REG_9_ , ADD_1071_U25 );
nand NAND2_7032 ( ADD_1071_U163 , P2_ADDR_REG_9_ , ADD_1071_U26 );
nand NAND2_7033 ( ADD_1071_U164 , P1_ADDR_REG_9_ , ADD_1071_U25 );
nand NAND2_7034 ( ADD_1071_U165 , ADD_1071_U164 , ADD_1071_U163 );
nand NAND3_7035 ( ADD_1071_U166 , ADD_1071_U162 , ADD_1071_U161 , ADD_1071_U64 );
nand NAND2_7036 ( ADD_1071_U167 , ADD_1071_U115 , ADD_1071_U165 );
nand NAND2_7037 ( ADD_1071_U168 , P2_ADDR_REG_8_ , ADD_1071_U23 );
nand NAND2_7038 ( ADD_1071_U169 , P1_ADDR_REG_8_ , ADD_1071_U24 );
nand NAND2_7039 ( ADD_1071_U170 , P2_ADDR_REG_8_ , ADD_1071_U23 );
nand NAND2_7040 ( ADD_1071_U171 , P1_ADDR_REG_8_ , ADD_1071_U24 );
nand NAND2_7041 ( ADD_1071_U172 , ADD_1071_U171 , ADD_1071_U170 );
nand NAND3_7042 ( ADD_1071_U173 , ADD_1071_U169 , ADD_1071_U168 , ADD_1071_U65 );
nand NAND2_7043 ( ADD_1071_U174 , ADD_1071_U111 , ADD_1071_U172 );
nand NAND2_7044 ( ADD_1071_U175 , P2_ADDR_REG_7_ , ADD_1071_U21 );
nand NAND2_7045 ( ADD_1071_U176 , P1_ADDR_REG_7_ , ADD_1071_U22 );
nand NAND2_7046 ( ADD_1071_U177 , P2_ADDR_REG_7_ , ADD_1071_U21 );
nand NAND2_7047 ( ADD_1071_U178 , P1_ADDR_REG_7_ , ADD_1071_U22 );
nand NAND2_7048 ( ADD_1071_U179 , ADD_1071_U178 , ADD_1071_U177 );
nand NAND3_7049 ( ADD_1071_U180 , ADD_1071_U176 , ADD_1071_U175 , ADD_1071_U66 );
nand NAND2_7050 ( ADD_1071_U181 , ADD_1071_U107 , ADD_1071_U179 );
nand NAND2_7051 ( ADD_1071_U182 , P2_ADDR_REG_6_ , ADD_1071_U19 );
nand NAND2_7052 ( ADD_1071_U183 , P1_ADDR_REG_6_ , ADD_1071_U20 );
nand NAND2_7053 ( ADD_1071_U184 , P2_ADDR_REG_6_ , ADD_1071_U19 );
nand NAND2_7054 ( ADD_1071_U185 , P1_ADDR_REG_6_ , ADD_1071_U20 );
nand NAND2_7055 ( ADD_1071_U186 , ADD_1071_U185 , ADD_1071_U184 );
nand NAND3_7056 ( ADD_1071_U187 , ADD_1071_U183 , ADD_1071_U182 , ADD_1071_U67 );
nand NAND2_7057 ( ADD_1071_U188 , ADD_1071_U103 , ADD_1071_U186 );
nand NAND2_7058 ( ADD_1071_U189 , P2_ADDR_REG_5_ , ADD_1071_U17 );
nand NAND2_7059 ( ADD_1071_U190 , P1_ADDR_REG_5_ , ADD_1071_U18 );
nand NAND2_7060 ( ADD_1071_U191 , P2_ADDR_REG_5_ , ADD_1071_U17 );
nand NAND2_7061 ( ADD_1071_U192 , P1_ADDR_REG_5_ , ADD_1071_U18 );
nand NAND2_7062 ( ADD_1071_U193 , ADD_1071_U192 , ADD_1071_U191 );
nand NAND3_7063 ( ADD_1071_U194 , ADD_1071_U190 , ADD_1071_U189 , ADD_1071_U68 );
nand NAND2_7064 ( ADD_1071_U195 , ADD_1071_U99 , ADD_1071_U193 );
nand NAND2_7065 ( ADD_1071_U196 , P2_ADDR_REG_4_ , ADD_1071_U15 );
nand NAND2_7066 ( ADD_1071_U197 , P1_ADDR_REG_4_ , ADD_1071_U16 );
nand NAND2_7067 ( ADD_1071_U198 , P2_ADDR_REG_4_ , ADD_1071_U15 );
nand NAND2_7068 ( ADD_1071_U199 , P1_ADDR_REG_4_ , ADD_1071_U16 );
nand NAND2_7069 ( ADD_1071_U200 , ADD_1071_U199 , ADD_1071_U198 );
nand NAND3_7070 ( ADD_1071_U201 , ADD_1071_U197 , ADD_1071_U196 , ADD_1071_U69 );
nand NAND2_7071 ( ADD_1071_U202 , ADD_1071_U95 , ADD_1071_U200 );
nand NAND2_7072 ( ADD_1071_U203 , P2_ADDR_REG_3_ , ADD_1071_U13 );
nand NAND2_7073 ( ADD_1071_U204 , P1_ADDR_REG_3_ , ADD_1071_U14 );
nand NAND2_7074 ( ADD_1071_U205 , P2_ADDR_REG_3_ , ADD_1071_U13 );
nand NAND2_7075 ( ADD_1071_U206 , P1_ADDR_REG_3_ , ADD_1071_U14 );
nand NAND2_7076 ( ADD_1071_U207 , ADD_1071_U206 , ADD_1071_U205 );
nand NAND3_7077 ( ADD_1071_U208 , ADD_1071_U204 , ADD_1071_U203 , ADD_1071_U70 );
nand NAND2_7078 ( ADD_1071_U209 , ADD_1071_U91 , ADD_1071_U207 );
nand NAND2_7079 ( ADD_1071_U210 , P2_ADDR_REG_2_ , ADD_1071_U11 );
nand NAND2_7080 ( ADD_1071_U211 , P1_ADDR_REG_2_ , ADD_1071_U12 );
nand NAND2_7081 ( ADD_1071_U212 , P2_ADDR_REG_2_ , ADD_1071_U11 );
nand NAND2_7082 ( ADD_1071_U213 , P1_ADDR_REG_2_ , ADD_1071_U12 );
nand NAND2_7083 ( ADD_1071_U214 , ADD_1071_U213 , ADD_1071_U212 );
nand NAND3_7084 ( ADD_1071_U215 , ADD_1071_U211 , ADD_1071_U210 , ADD_1071_U71 );
nand NAND2_7085 ( ADD_1071_U216 , ADD_1071_U87 , ADD_1071_U214 );
nand NAND2_7086 ( ADD_1071_U217 , P2_ADDR_REG_1_ , ADD_1071_U9 );
nand NAND2_7087 ( ADD_1071_U218 , ADD_1071_U84 , ADD_1071_U8 );
nand NAND2_7088 ( ADD_1071_U219 , ADD_1071_U218 , ADD_1071_U217 );
nand NAND3_7089 ( ADD_1071_U220 , P1_ADDR_REG_1_ , ADD_1071_U9 , ADD_1071_U8 );
nand NAND2_7090 ( ADD_1071_U221 , ADD_1071_U83 , P2_ADDR_REG_1_ );
nand NAND2_7091 ( ADD_1071_U222 , P2_ADDR_REG_19_ , ADD_1071_U74 );
nand NAND2_7092 ( ADD_1071_U223 , P1_ADDR_REG_19_ , ADD_1071_U73 );
nand NAND2_7093 ( ADD_1071_U224 , P2_ADDR_REG_19_ , ADD_1071_U74 );
nand NAND2_7094 ( ADD_1071_U225 , P1_ADDR_REG_19_ , ADD_1071_U73 );
nand NAND2_7095 ( ADD_1071_U226 , ADD_1071_U225 , ADD_1071_U224 );
nand NAND2_7096 ( ADD_1071_U227 , P2_ADDR_REG_18_ , ADD_1071_U43 );
nand NAND2_7097 ( ADD_1071_U228 , P1_ADDR_REG_18_ , ADD_1071_U44 );
nand NAND2_7098 ( ADD_1071_U229 , P2_ADDR_REG_18_ , ADD_1071_U43 );
nand NAND2_7099 ( ADD_1071_U230 , P1_ADDR_REG_18_ , ADD_1071_U44 );
nand NAND2_7100 ( ADD_1071_U231 , ADD_1071_U230 , ADD_1071_U229 );
nand NAND3_7101 ( ADD_1071_U232 , ADD_1071_U228 , ADD_1071_U227 , ADD_1071_U45 );
nand NAND2_7102 ( ADD_1071_U233 , ADD_1071_U231 , ADD_1071_U151 );
nand NAND2_7103 ( ADD_1071_U234 , P2_ADDR_REG_17_ , ADD_1071_U41 );
nand NAND2_7104 ( ADD_1071_U235 , P1_ADDR_REG_17_ , ADD_1071_U42 );
nand NAND2_7105 ( ADD_1071_U236 , P2_ADDR_REG_17_ , ADD_1071_U41 );
nand NAND2_7106 ( ADD_1071_U237 , P1_ADDR_REG_17_ , ADD_1071_U42 );
nand NAND2_7107 ( ADD_1071_U238 , ADD_1071_U237 , ADD_1071_U236 );
nand NAND3_7108 ( ADD_1071_U239 , ADD_1071_U235 , ADD_1071_U234 , ADD_1071_U75 );
nand NAND2_7109 ( ADD_1071_U240 , ADD_1071_U147 , ADD_1071_U238 );
nand NAND2_7110 ( ADD_1071_U241 , P2_ADDR_REG_16_ , ADD_1071_U39 );
nand NAND2_7111 ( ADD_1071_U242 , P1_ADDR_REG_16_ , ADD_1071_U40 );
nand NAND2_7112 ( ADD_1071_U243 , P2_ADDR_REG_16_ , ADD_1071_U39 );
nand NAND2_7113 ( ADD_1071_U244 , P1_ADDR_REG_16_ , ADD_1071_U40 );
nand NAND2_7114 ( ADD_1071_U245 , ADD_1071_U244 , ADD_1071_U243 );
nand NAND3_7115 ( ADD_1071_U246 , ADD_1071_U242 , ADD_1071_U241 , ADD_1071_U76 );
nand NAND2_7116 ( ADD_1071_U247 , ADD_1071_U143 , ADD_1071_U245 );
nand NAND2_7117 ( ADD_1071_U248 , P2_ADDR_REG_15_ , ADD_1071_U37 );
nand NAND2_7118 ( ADD_1071_U249 , P1_ADDR_REG_15_ , ADD_1071_U38 );
nand NAND2_7119 ( ADD_1071_U250 , P2_ADDR_REG_15_ , ADD_1071_U37 );
nand NAND2_7120 ( ADD_1071_U251 , P1_ADDR_REG_15_ , ADD_1071_U38 );
nand NAND2_7121 ( ADD_1071_U252 , ADD_1071_U251 , ADD_1071_U250 );
nand NAND3_7122 ( ADD_1071_U253 , ADD_1071_U249 , ADD_1071_U248 , ADD_1071_U77 );
nand NAND2_7123 ( ADD_1071_U254 , ADD_1071_U139 , ADD_1071_U252 );
nand NAND2_7124 ( ADD_1071_U255 , P2_ADDR_REG_14_ , ADD_1071_U35 );
nand NAND2_7125 ( ADD_1071_U256 , P1_ADDR_REG_14_ , ADD_1071_U36 );
nand NAND2_7126 ( ADD_1071_U257 , P2_ADDR_REG_14_ , ADD_1071_U35 );
nand NAND2_7127 ( ADD_1071_U258 , P1_ADDR_REG_14_ , ADD_1071_U36 );
nand NAND2_7128 ( ADD_1071_U259 , ADD_1071_U258 , ADD_1071_U257 );
nand NAND3_7129 ( ADD_1071_U260 , ADD_1071_U256 , ADD_1071_U255 , ADD_1071_U78 );
nand NAND2_7130 ( ADD_1071_U261 , ADD_1071_U135 , ADD_1071_U259 );
nand NAND2_7131 ( ADD_1071_U262 , P2_ADDR_REG_13_ , ADD_1071_U33 );
nand NAND2_7132 ( ADD_1071_U263 , P1_ADDR_REG_13_ , ADD_1071_U34 );
nand NAND2_7133 ( ADD_1071_U264 , P2_ADDR_REG_13_ , ADD_1071_U33 );
nand NAND2_7134 ( ADD_1071_U265 , P1_ADDR_REG_13_ , ADD_1071_U34 );
nand NAND2_7135 ( ADD_1071_U266 , ADD_1071_U265 , ADD_1071_U264 );
nand NAND3_7136 ( ADD_1071_U267 , ADD_1071_U263 , ADD_1071_U262 , ADD_1071_U79 );
nand NAND2_7137 ( ADD_1071_U268 , ADD_1071_U131 , ADD_1071_U266 );
nand NAND2_7138 ( ADD_1071_U269 , P2_ADDR_REG_12_ , ADD_1071_U31 );
nand NAND2_7139 ( ADD_1071_U270 , P1_ADDR_REG_12_ , ADD_1071_U32 );
nand NAND2_7140 ( ADD_1071_U271 , P2_ADDR_REG_12_ , ADD_1071_U31 );
nand NAND2_7141 ( ADD_1071_U272 , P1_ADDR_REG_12_ , ADD_1071_U32 );
nand NAND2_7142 ( ADD_1071_U273 , ADD_1071_U272 , ADD_1071_U271 );
nand NAND3_7143 ( ADD_1071_U274 , ADD_1071_U270 , ADD_1071_U269 , ADD_1071_U80 );
nand NAND2_7144 ( ADD_1071_U275 , ADD_1071_U127 , ADD_1071_U273 );
nand NAND2_7145 ( ADD_1071_U276 , P2_ADDR_REG_11_ , ADD_1071_U29 );
nand NAND2_7146 ( ADD_1071_U277 , P1_ADDR_REG_11_ , ADD_1071_U30 );
nand NAND2_7147 ( ADD_1071_U278 , P2_ADDR_REG_11_ , ADD_1071_U29 );
nand NAND2_7148 ( ADD_1071_U279 , P1_ADDR_REG_11_ , ADD_1071_U30 );
nand NAND2_7149 ( ADD_1071_U280 , ADD_1071_U279 , ADD_1071_U278 );
nand NAND3_7150 ( ADD_1071_U281 , ADD_1071_U277 , ADD_1071_U276 , ADD_1071_U81 );
nand NAND2_7151 ( ADD_1071_U282 , ADD_1071_U123 , ADD_1071_U280 );
nand NAND2_7152 ( ADD_1071_U283 , P2_ADDR_REG_10_ , ADD_1071_U27 );
nand NAND2_7153 ( ADD_1071_U284 , P1_ADDR_REG_10_ , ADD_1071_U28 );
nand NAND2_7154 ( ADD_1071_U285 , P2_ADDR_REG_10_ , ADD_1071_U27 );
nand NAND2_7155 ( ADD_1071_U286 , P1_ADDR_REG_10_ , ADD_1071_U28 );
nand NAND2_7156 ( ADD_1071_U287 , ADD_1071_U286 , ADD_1071_U285 );
nand NAND3_7157 ( ADD_1071_U288 , ADD_1071_U284 , ADD_1071_U283 , ADD_1071_U82 );
nand NAND2_7158 ( ADD_1071_U289 , ADD_1071_U119 , ADD_1071_U287 );
nand NAND2_7159 ( ADD_1071_U290 , P2_ADDR_REG_0_ , ADD_1071_U6 );
nand NAND2_7160 ( ADD_1071_U291 , P1_ADDR_REG_0_ , ADD_1071_U7 );
and AND2_7161 ( R140_U4 , R140_U197 , R140_U195 );
and AND2_7162 ( R140_U5 , R140_U203 , R140_U201 );
and AND2_7163 ( R140_U6 , R140_U5 , R140_U205 );
and AND2_7164 ( R140_U7 , R140_U213 , R140_U209 );
and AND2_7165 ( R140_U8 , R140_U7 , R140_U216 );
and AND2_7166 ( R140_U9 , R140_U378 , R140_U377 );
nand NAND3_7167 ( R140_U10 , R140_U469 , R140_U468 , R140_U324 );
and AND2_7168 ( R140_U11 , R140_U124 , R140_U323 );
not NOT1_7169 ( R140_U12 , SI_8_ );
not NOT1_7170 ( R140_U13 , U90 );
not NOT1_7171 ( R140_U14 , SI_7_ );
not NOT1_7172 ( R140_U15 , U91 );
nand NAND2_7173 ( R140_U16 , U91 , SI_7_ );
not NOT1_7174 ( R140_U17 , SI_6_ );
not NOT1_7175 ( R140_U18 , U92 );
not NOT1_7176 ( R140_U19 , SI_5_ );
not NOT1_7177 ( R140_U20 , U93 );
not NOT1_7178 ( R140_U21 , SI_4_ );
not NOT1_7179 ( R140_U22 , U94 );
nand NAND2_7180 ( R140_U23 , U94 , SI_4_ );
not NOT1_7181 ( R140_U24 , SI_3_ );
not NOT1_7182 ( R140_U25 , U97 );
not NOT1_7183 ( R140_U26 , SI_2_ );
not NOT1_7184 ( R140_U27 , U108 );
nand NAND2_7185 ( R140_U28 , U108 , SI_2_ );
not NOT1_7186 ( R140_U29 , SI_1_ );
not NOT1_7187 ( R140_U30 , SI_0_ );
not NOT1_7188 ( R140_U31 , U120 );
not NOT1_7189 ( R140_U32 , U119 );
not NOT1_7190 ( R140_U33 , U89 );
not NOT1_7191 ( R140_U34 , SI_9_ );
nand NAND2_7192 ( R140_U35 , R140_U288 , R140_U198 );
not NOT1_7193 ( R140_U36 , SI_14_ );
not NOT1_7194 ( R140_U37 , U114 );
not NOT1_7195 ( R140_U38 , SI_10_ );
not NOT1_7196 ( R140_U39 , U118 );
not NOT1_7197 ( R140_U40 , SI_13_ );
not NOT1_7198 ( R140_U41 , U115 );
not NOT1_7199 ( R140_U42 , SI_12_ );
not NOT1_7200 ( R140_U43 , U116 );
not NOT1_7201 ( R140_U44 , SI_11_ );
not NOT1_7202 ( R140_U45 , U117 );
nand NAND2_7203 ( R140_U46 , U117 , SI_11_ );
not NOT1_7204 ( R140_U47 , SI_15_ );
not NOT1_7205 ( R140_U48 , U113 );
not NOT1_7206 ( R140_U49 , SI_16_ );
not NOT1_7207 ( R140_U50 , U112 );
not NOT1_7208 ( R140_U51 , SI_17_ );
not NOT1_7209 ( R140_U52 , U111 );
not NOT1_7210 ( R140_U53 , SI_18_ );
not NOT1_7211 ( R140_U54 , U110 );
not NOT1_7212 ( R140_U55 , SI_19_ );
not NOT1_7213 ( R140_U56 , U109 );
not NOT1_7214 ( R140_U57 , SI_20_ );
not NOT1_7215 ( R140_U58 , U107 );
not NOT1_7216 ( R140_U59 , SI_21_ );
not NOT1_7217 ( R140_U60 , U106 );
not NOT1_7218 ( R140_U61 , SI_22_ );
not NOT1_7219 ( R140_U62 , U105 );
not NOT1_7220 ( R140_U63 , SI_23_ );
not NOT1_7221 ( R140_U64 , U104 );
not NOT1_7222 ( R140_U65 , SI_24_ );
not NOT1_7223 ( R140_U66 , U103 );
not NOT1_7224 ( R140_U67 , SI_25_ );
not NOT1_7225 ( R140_U68 , U102 );
not NOT1_7226 ( R140_U69 , SI_26_ );
not NOT1_7227 ( R140_U70 , U101 );
not NOT1_7228 ( R140_U71 , SI_27_ );
not NOT1_7229 ( R140_U72 , U100 );
not NOT1_7230 ( R140_U73 , SI_28_ );
not NOT1_7231 ( R140_U74 , U99 );
not NOT1_7232 ( R140_U75 , SI_29_ );
not NOT1_7233 ( R140_U76 , U98 );
not NOT1_7234 ( R140_U77 , SI_30_ );
not NOT1_7235 ( R140_U78 , U96 );
nand NAND3_7236 ( R140_U79 , SI_0_ , SI_1_ , U120 );
nand NAND2_7237 ( R140_U80 , R140_U300 , R140_U217 );
nand NAND2_7238 ( R140_U81 , R140_U297 , R140_U214 );
nand NAND2_7239 ( R140_U82 , R140_U293 , R140_U206 );
nand NAND2_7240 ( R140_U83 , R140_U541 , R140_U540 );
nand NAND2_7241 ( R140_U84 , R140_U331 , R140_U330 );
nand NAND2_7242 ( R140_U85 , R140_U338 , R140_U337 );
nand NAND2_7243 ( R140_U86 , R140_U345 , R140_U344 );
nand NAND2_7244 ( R140_U87 , R140_U352 , R140_U351 );
nand NAND2_7245 ( R140_U88 , R140_U359 , R140_U358 );
nand NAND2_7246 ( R140_U89 , R140_U366 , R140_U365 );
nand NAND2_7247 ( R140_U90 , R140_U373 , R140_U372 );
nand NAND2_7248 ( R140_U91 , R140_U387 , R140_U386 );
nand NAND2_7249 ( R140_U92 , R140_U394 , R140_U393 );
nand NAND2_7250 ( R140_U93 , R140_U401 , R140_U400 );
nand NAND2_7251 ( R140_U94 , R140_U408 , R140_U407 );
nand NAND2_7252 ( R140_U95 , R140_U415 , R140_U414 );
nand NAND2_7253 ( R140_U96 , R140_U422 , R140_U421 );
nand NAND2_7254 ( R140_U97 , R140_U429 , R140_U428 );
nand NAND2_7255 ( R140_U98 , R140_U436 , R140_U435 );
nand NAND2_7256 ( R140_U99 , R140_U443 , R140_U442 );
nand NAND2_7257 ( R140_U100 , R140_U450 , R140_U449 );
nand NAND2_7258 ( R140_U101 , R140_U457 , R140_U456 );
nand NAND2_7259 ( R140_U102 , R140_U464 , R140_U463 );
nand NAND2_7260 ( R140_U103 , R140_U476 , R140_U475 );
nand NAND2_7261 ( R140_U104 , R140_U483 , R140_U482 );
nand NAND2_7262 ( R140_U105 , R140_U490 , R140_U489 );
nand NAND2_7263 ( R140_U106 , R140_U497 , R140_U496 );
nand NAND2_7264 ( R140_U107 , R140_U504 , R140_U503 );
nand NAND2_7265 ( R140_U108 , R140_U511 , R140_U510 );
nand NAND2_7266 ( R140_U109 , R140_U518 , R140_U517 );
nand NAND2_7267 ( R140_U110 , R140_U525 , R140_U524 );
nand NAND2_7268 ( R140_U111 , R140_U532 , R140_U531 );
nand NAND2_7269 ( R140_U112 , R140_U539 , R140_U538 );
and AND2_7270 ( R140_U113 , R140_U189 , R140_U193 );
and AND2_7271 ( R140_U114 , R140_U287 , R140_U194 );
and AND2_7272 ( R140_U115 , R140_U4 , R140_U199 );
and AND2_7273 ( R140_U116 , R140_U290 , R140_U200 );
and AND2_7274 ( R140_U117 , R140_U291 , R140_U204 );
and AND2_7275 ( R140_U118 , R140_U6 , R140_U207 );
and AND2_7276 ( R140_U119 , R140_U295 , R140_U208 );
and AND2_7277 ( R140_U120 , R140_U8 , R140_U219 );
and AND2_7278 ( R140_U121 , R140_U303 , R140_U220 );
and AND3_7279 ( R140_U122 , R140_U9 , R140_U282 , R140_U280 );
and AND2_7280 ( R140_U123 , R140_U283 , R140_U376 );
and AND2_7281 ( R140_U124 , R140_U141 , R140_U284 );
and AND2_7282 ( R140_U125 , R140_U326 , R140_U325 );
nand NAND2_7283 ( R140_U126 , R140_U117 , R140_U309 );
and AND2_7284 ( R140_U127 , R140_U333 , R140_U332 );
nand NAND2_7285 ( R140_U128 , R140_U307 , R140_U16 );
and AND2_7286 ( R140_U129 , R140_U340 , R140_U339 );
nand NAND2_7287 ( R140_U130 , R140_U116 , R140_U319 );
and AND2_7288 ( R140_U131 , R140_U347 , R140_U346 );
nand NAND2_7289 ( R140_U132 , R140_U289 , R140_U317 );
and AND2_7290 ( R140_U133 , R140_U354 , R140_U353 );
nand NAND2_7291 ( R140_U134 , R140_U315 , R140_U23 );
and AND2_7292 ( R140_U135 , R140_U361 , R140_U360 );
nand NAND2_7293 ( R140_U136 , R140_U114 , R140_U321 );
and AND2_7294 ( R140_U137 , R140_U368 , R140_U367 );
nand NAND2_7295 ( R140_U138 , R140_U28 , R140_U190 );
not NOT1_7296 ( R140_U139 , U95 );
not NOT1_7297 ( R140_U140 , SI_31_ );
and AND2_7298 ( R140_U141 , R140_U380 , R140_U379 );
and AND2_7299 ( R140_U142 , R140_U382 , R140_U381 );
nand NAND2_7300 ( R140_U143 , R140_U280 , R140_U279 );
nand NAND3_7301 ( R140_U144 , R140_U286 , R140_U79 , R140_U285 );
and AND2_7302 ( R140_U145 , R140_U396 , R140_U395 );
nand NAND2_7303 ( R140_U146 , R140_U276 , R140_U275 );
and AND2_7304 ( R140_U147 , R140_U403 , R140_U402 );
nand NAND2_7305 ( R140_U148 , R140_U272 , R140_U271 );
and AND2_7306 ( R140_U149 , R140_U410 , R140_U409 );
nand NAND2_7307 ( R140_U150 , R140_U268 , R140_U267 );
and AND2_7308 ( R140_U151 , R140_U417 , R140_U416 );
nand NAND2_7309 ( R140_U152 , R140_U264 , R140_U263 );
and AND2_7310 ( R140_U153 , R140_U424 , R140_U423 );
nand NAND2_7311 ( R140_U154 , R140_U260 , R140_U259 );
and AND2_7312 ( R140_U155 , R140_U431 , R140_U430 );
nand NAND2_7313 ( R140_U156 , R140_U256 , R140_U255 );
and AND2_7314 ( R140_U157 , R140_U438 , R140_U437 );
nand NAND2_7315 ( R140_U158 , R140_U252 , R140_U251 );
and AND2_7316 ( R140_U159 , R140_U445 , R140_U444 );
nand NAND2_7317 ( R140_U160 , R140_U248 , R140_U247 );
and AND2_7318 ( R140_U161 , R140_U452 , R140_U451 );
nand NAND2_7319 ( R140_U162 , R140_U244 , R140_U243 );
and AND2_7320 ( R140_U163 , R140_U459 , R140_U458 );
nand NAND2_7321 ( R140_U164 , R140_U240 , R140_U239 );
nand NAND2_7322 ( R140_U165 , U120 , SI_0_ );
and AND2_7323 ( R140_U166 , R140_U471 , R140_U470 );
nand NAND2_7324 ( R140_U167 , R140_U236 , R140_U235 );
and AND2_7325 ( R140_U168 , R140_U478 , R140_U477 );
nand NAND2_7326 ( R140_U169 , R140_U232 , R140_U231 );
and AND2_7327 ( R140_U170 , R140_U485 , R140_U484 );
nand NAND2_7328 ( R140_U171 , R140_U228 , R140_U227 );
and AND2_7329 ( R140_U172 , R140_U492 , R140_U491 );
nand NAND2_7330 ( R140_U173 , R140_U224 , R140_U223 );
and AND2_7331 ( R140_U174 , R140_U499 , R140_U498 );
nand NAND2_7332 ( R140_U175 , R140_U121 , R140_U302 );
and AND2_7333 ( R140_U176 , R140_U506 , R140_U505 );
nand NAND2_7334 ( R140_U177 , R140_U301 , R140_U299 );
and AND2_7335 ( R140_U178 , R140_U513 , R140_U512 );
nand NAND2_7336 ( R140_U179 , R140_U298 , R140_U296 );
and AND2_7337 ( R140_U180 , R140_U520 , R140_U519 );
nand NAND2_7338 ( R140_U181 , R140_U46 , R140_U210 );
and AND2_7339 ( R140_U182 , R140_U527 , R140_U526 );
nand NAND2_7340 ( R140_U183 , R140_U119 , R140_U313 );
and AND2_7341 ( R140_U184 , R140_U534 , R140_U533 );
nand NAND2_7342 ( R140_U185 , R140_U294 , R140_U311 );
not NOT1_7343 ( R140_U186 , R140_U79 );
not NOT1_7344 ( R140_U187 , R140_U165 );
not NOT1_7345 ( R140_U188 , R140_U144 );
or OR2_7346 ( R140_U189 , SI_2_ , U108 );
nand NAND2_7347 ( R140_U190 , R140_U304 , R140_U189 );
not NOT1_7348 ( R140_U191 , R140_U28 );
not NOT1_7349 ( R140_U192 , R140_U138 );
or OR2_7350 ( R140_U193 , SI_3_ , U97 );
nand NAND2_7351 ( R140_U194 , U97 , SI_3_ );
or OR2_7352 ( R140_U195 , SI_4_ , U94 );
not NOT1_7353 ( R140_U196 , R140_U23 );
or OR2_7354 ( R140_U197 , SI_5_ , U93 );
nand NAND2_7355 ( R140_U198 , U93 , SI_5_ );
or OR2_7356 ( R140_U199 , SI_6_ , U92 );
nand NAND2_7357 ( R140_U200 , U92 , SI_6_ );
or OR2_7358 ( R140_U201 , SI_7_ , U91 );
not NOT1_7359 ( R140_U202 , R140_U16 );
or OR2_7360 ( R140_U203 , SI_8_ , U90 );
nand NAND2_7361 ( R140_U204 , U90 , SI_8_ );
or OR2_7362 ( R140_U205 , SI_9_ , U89 );
nand NAND2_7363 ( R140_U206 , SI_9_ , U89 );
or OR2_7364 ( R140_U207 , SI_10_ , U118 );
nand NAND2_7365 ( R140_U208 , U118 , SI_10_ );
or OR2_7366 ( R140_U209 , SI_11_ , U117 );
nand NAND2_7367 ( R140_U210 , R140_U209 , R140_U183 );
not NOT1_7368 ( R140_U211 , R140_U46 );
not NOT1_7369 ( R140_U212 , R140_U181 );
or OR2_7370 ( R140_U213 , SI_12_ , U116 );
nand NAND2_7371 ( R140_U214 , U116 , SI_12_ );
not NOT1_7372 ( R140_U215 , R140_U179 );
or OR2_7373 ( R140_U216 , SI_13_ , U115 );
nand NAND2_7374 ( R140_U217 , U115 , SI_13_ );
not NOT1_7375 ( R140_U218 , R140_U177 );
or OR2_7376 ( R140_U219 , SI_14_ , U114 );
nand NAND2_7377 ( R140_U220 , U114 , SI_14_ );
not NOT1_7378 ( R140_U221 , R140_U175 );
or OR2_7379 ( R140_U222 , SI_15_ , U113 );
nand NAND2_7380 ( R140_U223 , R140_U222 , R140_U175 );
nand NAND2_7381 ( R140_U224 , U113 , SI_15_ );
not NOT1_7382 ( R140_U225 , R140_U173 );
or OR2_7383 ( R140_U226 , SI_16_ , U112 );
nand NAND2_7384 ( R140_U227 , R140_U226 , R140_U173 );
nand NAND2_7385 ( R140_U228 , U112 , SI_16_ );
not NOT1_7386 ( R140_U229 , R140_U171 );
or OR2_7387 ( R140_U230 , SI_17_ , U111 );
nand NAND2_7388 ( R140_U231 , R140_U230 , R140_U171 );
nand NAND2_7389 ( R140_U232 , U111 , SI_17_ );
not NOT1_7390 ( R140_U233 , R140_U169 );
or OR2_7391 ( R140_U234 , SI_18_ , U110 );
nand NAND2_7392 ( R140_U235 , R140_U234 , R140_U169 );
nand NAND2_7393 ( R140_U236 , U110 , SI_18_ );
not NOT1_7394 ( R140_U237 , R140_U167 );
or OR2_7395 ( R140_U238 , SI_19_ , U109 );
nand NAND2_7396 ( R140_U239 , R140_U238 , R140_U167 );
nand NAND2_7397 ( R140_U240 , U109 , SI_19_ );
not NOT1_7398 ( R140_U241 , R140_U164 );
or OR2_7399 ( R140_U242 , SI_20_ , U107 );
nand NAND2_7400 ( R140_U243 , R140_U242 , R140_U164 );
nand NAND2_7401 ( R140_U244 , U107 , SI_20_ );
not NOT1_7402 ( R140_U245 , R140_U162 );
or OR2_7403 ( R140_U246 , SI_21_ , U106 );
nand NAND2_7404 ( R140_U247 , R140_U246 , R140_U162 );
nand NAND2_7405 ( R140_U248 , U106 , SI_21_ );
not NOT1_7406 ( R140_U249 , R140_U160 );
or OR2_7407 ( R140_U250 , SI_22_ , U105 );
nand NAND2_7408 ( R140_U251 , R140_U250 , R140_U160 );
nand NAND2_7409 ( R140_U252 , U105 , SI_22_ );
not NOT1_7410 ( R140_U253 , R140_U158 );
or OR2_7411 ( R140_U254 , SI_23_ , U104 );
nand NAND2_7412 ( R140_U255 , R140_U254 , R140_U158 );
nand NAND2_7413 ( R140_U256 , U104 , SI_23_ );
not NOT1_7414 ( R140_U257 , R140_U156 );
or OR2_7415 ( R140_U258 , SI_24_ , U103 );
nand NAND2_7416 ( R140_U259 , R140_U258 , R140_U156 );
nand NAND2_7417 ( R140_U260 , U103 , SI_24_ );
not NOT1_7418 ( R140_U261 , R140_U154 );
or OR2_7419 ( R140_U262 , SI_25_ , U102 );
nand NAND2_7420 ( R140_U263 , R140_U262 , R140_U154 );
nand NAND2_7421 ( R140_U264 , U102 , SI_25_ );
not NOT1_7422 ( R140_U265 , R140_U152 );
or OR2_7423 ( R140_U266 , SI_26_ , U101 );
nand NAND2_7424 ( R140_U267 , R140_U266 , R140_U152 );
nand NAND2_7425 ( R140_U268 , U101 , SI_26_ );
not NOT1_7426 ( R140_U269 , R140_U150 );
or OR2_7427 ( R140_U270 , SI_27_ , U100 );
nand NAND2_7428 ( R140_U271 , R140_U270 , R140_U150 );
nand NAND2_7429 ( R140_U272 , U100 , SI_27_ );
not NOT1_7430 ( R140_U273 , R140_U148 );
or OR2_7431 ( R140_U274 , SI_28_ , U99 );
nand NAND2_7432 ( R140_U275 , R140_U274 , R140_U148 );
nand NAND2_7433 ( R140_U276 , U99 , SI_28_ );
not NOT1_7434 ( R140_U277 , R140_U146 );
or OR2_7435 ( R140_U278 , SI_29_ , U98 );
nand NAND2_7436 ( R140_U279 , R140_U278 , R140_U146 );
nand NAND2_7437 ( R140_U280 , U98 , SI_29_ );
not NOT1_7438 ( R140_U281 , R140_U143 );
nand NAND2_7439 ( R140_U282 , U96 , SI_30_ );
or OR2_7440 ( R140_U283 , U96 , SI_30_ );
nand NAND2_7441 ( R140_U284 , R140_U279 , R140_U122 );
nand NAND3_7442 ( R140_U285 , U120 , SI_0_ , U119 );
nand NAND2_7443 ( R140_U286 , U119 , SI_1_ );
nand NAND2_7444 ( R140_U287 , R140_U191 , R140_U193 );
nand NAND2_7445 ( R140_U288 , R140_U196 , R140_U197 );
not NOT1_7446 ( R140_U289 , R140_U35 );
nand NAND2_7447 ( R140_U290 , R140_U35 , R140_U199 );
nand NAND2_7448 ( R140_U291 , R140_U202 , R140_U203 );
nand NAND2_7449 ( R140_U292 , R140_U291 , R140_U204 );
nand NAND2_7450 ( R140_U293 , R140_U292 , R140_U205 );
not NOT1_7451 ( R140_U294 , R140_U82 );
nand NAND2_7452 ( R140_U295 , R140_U82 , R140_U207 );
nand NAND2_7453 ( R140_U296 , R140_U7 , R140_U183 );
nand NAND2_7454 ( R140_U297 , R140_U211 , R140_U213 );
not NOT1_7455 ( R140_U298 , R140_U81 );
nand NAND2_7456 ( R140_U299 , R140_U8 , R140_U183 );
nand NAND2_7457 ( R140_U300 , R140_U81 , R140_U216 );
not NOT1_7458 ( R140_U301 , R140_U80 );
nand NAND2_7459 ( R140_U302 , R140_U120 , R140_U183 );
nand NAND2_7460 ( R140_U303 , R140_U80 , R140_U219 );
nand NAND3_7461 ( R140_U304 , R140_U306 , R140_U286 , R140_U305 );
nand NAND3_7462 ( R140_U305 , U120 , SI_0_ , U119 );
nand NAND3_7463 ( R140_U306 , SI_0_ , SI_1_ , U120 );
nand NAND2_7464 ( R140_U307 , R140_U201 , R140_U130 );
not NOT1_7465 ( R140_U308 , R140_U128 );
nand NAND2_7466 ( R140_U309 , R140_U5 , R140_U130 );
not NOT1_7467 ( R140_U310 , R140_U126 );
nand NAND2_7468 ( R140_U311 , R140_U6 , R140_U130 );
not NOT1_7469 ( R140_U312 , R140_U185 );
nand NAND2_7470 ( R140_U313 , R140_U118 , R140_U130 );
not NOT1_7471 ( R140_U314 , R140_U183 );
nand NAND2_7472 ( R140_U315 , R140_U195 , R140_U136 );
not NOT1_7473 ( R140_U316 , R140_U134 );
nand NAND2_7474 ( R140_U317 , R140_U4 , R140_U136 );
not NOT1_7475 ( R140_U318 , R140_U132 );
nand NAND2_7476 ( R140_U319 , R140_U115 , R140_U136 );
not NOT1_7477 ( R140_U320 , R140_U130 );
nand NAND2_7478 ( R140_U321 , R140_U113 , R140_U144 );
not NOT1_7479 ( R140_U322 , R140_U136 );
nand NAND2_7480 ( R140_U323 , R140_U123 , R140_U143 );
nand NAND2_7481 ( R140_U324 , R140_U186 , U119 );
nand NAND2_7482 ( R140_U325 , U89 , R140_U34 );
nand NAND2_7483 ( R140_U326 , SI_9_ , R140_U33 );
nand NAND2_7484 ( R140_U327 , U89 , R140_U34 );
nand NAND2_7485 ( R140_U328 , SI_9_ , R140_U33 );
nand NAND2_7486 ( R140_U329 , R140_U328 , R140_U327 );
nand NAND2_7487 ( R140_U330 , R140_U125 , R140_U126 );
nand NAND2_7488 ( R140_U331 , R140_U310 , R140_U329 );
nand NAND2_7489 ( R140_U332 , U90 , R140_U12 );
nand NAND2_7490 ( R140_U333 , SI_8_ , R140_U13 );
nand NAND2_7491 ( R140_U334 , U90 , R140_U12 );
nand NAND2_7492 ( R140_U335 , SI_8_ , R140_U13 );
nand NAND2_7493 ( R140_U336 , R140_U335 , R140_U334 );
nand NAND2_7494 ( R140_U337 , R140_U127 , R140_U128 );
nand NAND2_7495 ( R140_U338 , R140_U308 , R140_U336 );
nand NAND2_7496 ( R140_U339 , U91 , R140_U14 );
nand NAND2_7497 ( R140_U340 , SI_7_ , R140_U15 );
nand NAND2_7498 ( R140_U341 , U91 , R140_U14 );
nand NAND2_7499 ( R140_U342 , SI_7_ , R140_U15 );
nand NAND2_7500 ( R140_U343 , R140_U342 , R140_U341 );
nand NAND2_7501 ( R140_U344 , R140_U129 , R140_U130 );
nand NAND2_7502 ( R140_U345 , R140_U320 , R140_U343 );
nand NAND2_7503 ( R140_U346 , U92 , R140_U17 );
nand NAND2_7504 ( R140_U347 , SI_6_ , R140_U18 );
nand NAND2_7505 ( R140_U348 , U92 , R140_U17 );
nand NAND2_7506 ( R140_U349 , SI_6_ , R140_U18 );
nand NAND2_7507 ( R140_U350 , R140_U349 , R140_U348 );
nand NAND2_7508 ( R140_U351 , R140_U131 , R140_U132 );
nand NAND2_7509 ( R140_U352 , R140_U318 , R140_U350 );
nand NAND2_7510 ( R140_U353 , U93 , R140_U19 );
nand NAND2_7511 ( R140_U354 , SI_5_ , R140_U20 );
nand NAND2_7512 ( R140_U355 , U93 , R140_U19 );
nand NAND2_7513 ( R140_U356 , SI_5_ , R140_U20 );
nand NAND2_7514 ( R140_U357 , R140_U356 , R140_U355 );
nand NAND2_7515 ( R140_U358 , R140_U133 , R140_U134 );
nand NAND2_7516 ( R140_U359 , R140_U316 , R140_U357 );
nand NAND2_7517 ( R140_U360 , U94 , R140_U21 );
nand NAND2_7518 ( R140_U361 , SI_4_ , R140_U22 );
nand NAND2_7519 ( R140_U362 , U94 , R140_U21 );
nand NAND2_7520 ( R140_U363 , SI_4_ , R140_U22 );
nand NAND2_7521 ( R140_U364 , R140_U363 , R140_U362 );
nand NAND2_7522 ( R140_U365 , R140_U135 , R140_U136 );
nand NAND2_7523 ( R140_U366 , R140_U322 , R140_U364 );
nand NAND2_7524 ( R140_U367 , U97 , R140_U24 );
nand NAND2_7525 ( R140_U368 , SI_3_ , R140_U25 );
nand NAND2_7526 ( R140_U369 , U97 , R140_U24 );
nand NAND2_7527 ( R140_U370 , SI_3_ , R140_U25 );
nand NAND2_7528 ( R140_U371 , R140_U370 , R140_U369 );
nand NAND2_7529 ( R140_U372 , R140_U137 , R140_U138 );
nand NAND2_7530 ( R140_U373 , R140_U192 , R140_U371 );
nand NAND2_7531 ( R140_U374 , U95 , R140_U140 );
nand NAND2_7532 ( R140_U375 , SI_31_ , R140_U139 );
nand NAND2_7533 ( R140_U376 , R140_U375 , R140_U374 );
nand NAND2_7534 ( R140_U377 , U95 , R140_U140 );
nand NAND2_7535 ( R140_U378 , SI_31_ , R140_U139 );
nand NAND3_7536 ( R140_U379 , R140_U9 , R140_U77 , R140_U78 );
nand NAND3_7537 ( R140_U380 , SI_30_ , R140_U376 , U96 );
nand NAND2_7538 ( R140_U381 , U96 , R140_U77 );
nand NAND2_7539 ( R140_U382 , SI_30_ , R140_U78 );
nand NAND2_7540 ( R140_U383 , U96 , R140_U77 );
nand NAND2_7541 ( R140_U384 , SI_30_ , R140_U78 );
nand NAND2_7542 ( R140_U385 , R140_U384 , R140_U383 );
nand NAND2_7543 ( R140_U386 , R140_U142 , R140_U143 );
nand NAND2_7544 ( R140_U387 , R140_U281 , R140_U385 );
nand NAND2_7545 ( R140_U388 , U108 , R140_U26 );
nand NAND2_7546 ( R140_U389 , SI_2_ , R140_U27 );
nand NAND2_7547 ( R140_U390 , U108 , R140_U26 );
nand NAND2_7548 ( R140_U391 , SI_2_ , R140_U27 );
nand NAND2_7549 ( R140_U392 , R140_U391 , R140_U390 );
nand NAND3_7550 ( R140_U393 , R140_U389 , R140_U388 , R140_U144 );
nand NAND2_7551 ( R140_U394 , R140_U188 , R140_U392 );
nand NAND2_7552 ( R140_U395 , U98 , R140_U75 );
nand NAND2_7553 ( R140_U396 , SI_29_ , R140_U76 );
nand NAND2_7554 ( R140_U397 , U98 , R140_U75 );
nand NAND2_7555 ( R140_U398 , SI_29_ , R140_U76 );
nand NAND2_7556 ( R140_U399 , R140_U398 , R140_U397 );
nand NAND2_7557 ( R140_U400 , R140_U145 , R140_U146 );
nand NAND2_7558 ( R140_U401 , R140_U277 , R140_U399 );
nand NAND2_7559 ( R140_U402 , U99 , R140_U73 );
nand NAND2_7560 ( R140_U403 , SI_28_ , R140_U74 );
nand NAND2_7561 ( R140_U404 , U99 , R140_U73 );
nand NAND2_7562 ( R140_U405 , SI_28_ , R140_U74 );
nand NAND2_7563 ( R140_U406 , R140_U405 , R140_U404 );
nand NAND2_7564 ( R140_U407 , R140_U147 , R140_U148 );
nand NAND2_7565 ( R140_U408 , R140_U273 , R140_U406 );
nand NAND2_7566 ( R140_U409 , U100 , R140_U71 );
nand NAND2_7567 ( R140_U410 , SI_27_ , R140_U72 );
nand NAND2_7568 ( R140_U411 , U100 , R140_U71 );
nand NAND2_7569 ( R140_U412 , SI_27_ , R140_U72 );
nand NAND2_7570 ( R140_U413 , R140_U412 , R140_U411 );
nand NAND2_7571 ( R140_U414 , R140_U149 , R140_U150 );
nand NAND2_7572 ( R140_U415 , R140_U269 , R140_U413 );
nand NAND2_7573 ( R140_U416 , U101 , R140_U69 );
nand NAND2_7574 ( R140_U417 , SI_26_ , R140_U70 );
nand NAND2_7575 ( R140_U418 , U101 , R140_U69 );
nand NAND2_7576 ( R140_U419 , SI_26_ , R140_U70 );
nand NAND2_7577 ( R140_U420 , R140_U419 , R140_U418 );
nand NAND2_7578 ( R140_U421 , R140_U151 , R140_U152 );
nand NAND2_7579 ( R140_U422 , R140_U265 , R140_U420 );
nand NAND2_7580 ( R140_U423 , U102 , R140_U67 );
nand NAND2_7581 ( R140_U424 , SI_25_ , R140_U68 );
nand NAND2_7582 ( R140_U425 , U102 , R140_U67 );
nand NAND2_7583 ( R140_U426 , SI_25_ , R140_U68 );
nand NAND2_7584 ( R140_U427 , R140_U426 , R140_U425 );
nand NAND2_7585 ( R140_U428 , R140_U153 , R140_U154 );
nand NAND2_7586 ( R140_U429 , R140_U261 , R140_U427 );
nand NAND2_7587 ( R140_U430 , U103 , R140_U65 );
nand NAND2_7588 ( R140_U431 , SI_24_ , R140_U66 );
nand NAND2_7589 ( R140_U432 , U103 , R140_U65 );
nand NAND2_7590 ( R140_U433 , SI_24_ , R140_U66 );
nand NAND2_7591 ( R140_U434 , R140_U433 , R140_U432 );
nand NAND2_7592 ( R140_U435 , R140_U155 , R140_U156 );
nand NAND2_7593 ( R140_U436 , R140_U257 , R140_U434 );
nand NAND2_7594 ( R140_U437 , U104 , R140_U63 );
nand NAND2_7595 ( R140_U438 , SI_23_ , R140_U64 );
nand NAND2_7596 ( R140_U439 , U104 , R140_U63 );
nand NAND2_7597 ( R140_U440 , SI_23_ , R140_U64 );
nand NAND2_7598 ( R140_U441 , R140_U440 , R140_U439 );
nand NAND2_7599 ( R140_U442 , R140_U157 , R140_U158 );
nand NAND2_7600 ( R140_U443 , R140_U253 , R140_U441 );
nand NAND2_7601 ( R140_U444 , U105 , R140_U61 );
nand NAND2_7602 ( R140_U445 , SI_22_ , R140_U62 );
nand NAND2_7603 ( R140_U446 , U105 , R140_U61 );
nand NAND2_7604 ( R140_U447 , SI_22_ , R140_U62 );
nand NAND2_7605 ( R140_U448 , R140_U447 , R140_U446 );
nand NAND2_7606 ( R140_U449 , R140_U159 , R140_U160 );
nand NAND2_7607 ( R140_U450 , R140_U249 , R140_U448 );
nand NAND2_7608 ( R140_U451 , U106 , R140_U59 );
nand NAND2_7609 ( R140_U452 , SI_21_ , R140_U60 );
nand NAND2_7610 ( R140_U453 , U106 , R140_U59 );
nand NAND2_7611 ( R140_U454 , SI_21_ , R140_U60 );
nand NAND2_7612 ( R140_U455 , R140_U454 , R140_U453 );
nand NAND2_7613 ( R140_U456 , R140_U161 , R140_U162 );
nand NAND2_7614 ( R140_U457 , R140_U245 , R140_U455 );
nand NAND2_7615 ( R140_U458 , U107 , R140_U57 );
nand NAND2_7616 ( R140_U459 , SI_20_ , R140_U58 );
nand NAND2_7617 ( R140_U460 , U107 , R140_U57 );
nand NAND2_7618 ( R140_U461 , SI_20_ , R140_U58 );
nand NAND2_7619 ( R140_U462 , R140_U461 , R140_U460 );
nand NAND2_7620 ( R140_U463 , R140_U163 , R140_U164 );
nand NAND2_7621 ( R140_U464 , R140_U241 , R140_U462 );
nand NAND2_7622 ( R140_U465 , U119 , R140_U165 );
nand NAND2_7623 ( R140_U466 , R140_U187 , R140_U32 );
nand NAND2_7624 ( R140_U467 , R140_U466 , R140_U465 );
nand NAND3_7625 ( R140_U468 , R140_U165 , R140_U32 , SI_1_ );
nand NAND2_7626 ( R140_U469 , R140_U467 , R140_U29 );
nand NAND2_7627 ( R140_U470 , U109 , R140_U55 );
nand NAND2_7628 ( R140_U471 , SI_19_ , R140_U56 );
nand NAND2_7629 ( R140_U472 , U109 , R140_U55 );
nand NAND2_7630 ( R140_U473 , SI_19_ , R140_U56 );
nand NAND2_7631 ( R140_U474 , R140_U473 , R140_U472 );
nand NAND2_7632 ( R140_U475 , R140_U166 , R140_U167 );
nand NAND2_7633 ( R140_U476 , R140_U237 , R140_U474 );
nand NAND2_7634 ( R140_U477 , U110 , R140_U53 );
nand NAND2_7635 ( R140_U478 , SI_18_ , R140_U54 );
nand NAND2_7636 ( R140_U479 , U110 , R140_U53 );
nand NAND2_7637 ( R140_U480 , SI_18_ , R140_U54 );
nand NAND2_7638 ( R140_U481 , R140_U480 , R140_U479 );
nand NAND2_7639 ( R140_U482 , R140_U168 , R140_U169 );
nand NAND2_7640 ( R140_U483 , R140_U233 , R140_U481 );
nand NAND2_7641 ( R140_U484 , U111 , R140_U51 );
nand NAND2_7642 ( R140_U485 , SI_17_ , R140_U52 );
nand NAND2_7643 ( R140_U486 , U111 , R140_U51 );
nand NAND2_7644 ( R140_U487 , SI_17_ , R140_U52 );
nand NAND2_7645 ( R140_U488 , R140_U487 , R140_U486 );
nand NAND2_7646 ( R140_U489 , R140_U170 , R140_U171 );
nand NAND2_7647 ( R140_U490 , R140_U229 , R140_U488 );
nand NAND2_7648 ( R140_U491 , U112 , R140_U49 );
nand NAND2_7649 ( R140_U492 , SI_16_ , R140_U50 );
nand NAND2_7650 ( R140_U493 , U112 , R140_U49 );
nand NAND2_7651 ( R140_U494 , SI_16_ , R140_U50 );
nand NAND2_7652 ( R140_U495 , R140_U494 , R140_U493 );
nand NAND2_7653 ( R140_U496 , R140_U172 , R140_U173 );
nand NAND2_7654 ( R140_U497 , R140_U225 , R140_U495 );
nand NAND2_7655 ( R140_U498 , U113 , R140_U47 );
nand NAND2_7656 ( R140_U499 , SI_15_ , R140_U48 );
nand NAND2_7657 ( R140_U500 , U113 , R140_U47 );
nand NAND2_7658 ( R140_U501 , SI_15_ , R140_U48 );
nand NAND2_7659 ( R140_U502 , R140_U501 , R140_U500 );
nand NAND2_7660 ( R140_U503 , R140_U174 , R140_U175 );
nand NAND2_7661 ( R140_U504 , R140_U221 , R140_U502 );
nand NAND2_7662 ( R140_U505 , U114 , R140_U36 );
nand NAND2_7663 ( R140_U506 , SI_14_ , R140_U37 );
nand NAND2_7664 ( R140_U507 , U114 , R140_U36 );
nand NAND2_7665 ( R140_U508 , SI_14_ , R140_U37 );
nand NAND2_7666 ( R140_U509 , R140_U508 , R140_U507 );
nand NAND2_7667 ( R140_U510 , R140_U176 , R140_U177 );
nand NAND2_7668 ( R140_U511 , R140_U218 , R140_U509 );
nand NAND2_7669 ( R140_U512 , U115 , R140_U40 );
nand NAND2_7670 ( R140_U513 , SI_13_ , R140_U41 );
nand NAND2_7671 ( R140_U514 , U115 , R140_U40 );
nand NAND2_7672 ( R140_U515 , SI_13_ , R140_U41 );
nand NAND2_7673 ( R140_U516 , R140_U515 , R140_U514 );
nand NAND2_7674 ( R140_U517 , R140_U178 , R140_U179 );
nand NAND2_7675 ( R140_U518 , R140_U215 , R140_U516 );
nand NAND2_7676 ( R140_U519 , U116 , R140_U42 );
nand NAND2_7677 ( R140_U520 , SI_12_ , R140_U43 );
nand NAND2_7678 ( R140_U521 , U116 , R140_U42 );
nand NAND2_7679 ( R140_U522 , SI_12_ , R140_U43 );
nand NAND2_7680 ( R140_U523 , R140_U522 , R140_U521 );
nand NAND2_7681 ( R140_U524 , R140_U180 , R140_U181 );
nand NAND2_7682 ( R140_U525 , R140_U212 , R140_U523 );
nand NAND2_7683 ( R140_U526 , U117 , R140_U44 );
nand NAND2_7684 ( R140_U527 , SI_11_ , R140_U45 );
nand NAND2_7685 ( R140_U528 , U117 , R140_U44 );
nand NAND2_7686 ( R140_U529 , SI_11_ , R140_U45 );
nand NAND2_7687 ( R140_U530 , R140_U529 , R140_U528 );
nand NAND2_7688 ( R140_U531 , R140_U182 , R140_U183 );
nand NAND2_7689 ( R140_U532 , R140_U314 , R140_U530 );
nand NAND2_7690 ( R140_U533 , U118 , R140_U38 );
nand NAND2_7691 ( R140_U534 , SI_10_ , R140_U39 );
nand NAND2_7692 ( R140_U535 , U118 , R140_U38 );
nand NAND2_7693 ( R140_U536 , SI_10_ , R140_U39 );
nand NAND2_7694 ( R140_U537 , R140_U536 , R140_U535 );
nand NAND2_7695 ( R140_U538 , R140_U184 , R140_U185 );
nand NAND2_7696 ( R140_U539 , R140_U312 , R140_U537 );
nand NAND2_7697 ( R140_U540 , U120 , R140_U30 );
nand NAND2_7698 ( R140_U541 , SI_0_ , R140_U31 );
not NOT1_7699 ( LT_1079_19_U6 , P2_ADDR_REG_19_ );
not NOT1_7700 ( P1_ADD_99_U4 , P1_REG3_REG_3_ );
and AND3_7701 ( P1_ADD_99_U5 , P1_REG3_REG_28_ , P1_REG3_REG_27_ , P1_ADD_99_U102 );
not NOT1_7702 ( P1_ADD_99_U6 , P1_REG3_REG_4_ );
nand NAND2_7703 ( P1_ADD_99_U7 , P1_REG3_REG_4_ , P1_REG3_REG_3_ );
not NOT1_7704 ( P1_ADD_99_U8 , P1_REG3_REG_5_ );
nand NAND2_7705 ( P1_ADD_99_U9 , P1_REG3_REG_5_ , P1_ADD_99_U80 );
not NOT1_7706 ( P1_ADD_99_U10 , P1_REG3_REG_6_ );
nand NAND2_7707 ( P1_ADD_99_U11 , P1_REG3_REG_6_ , P1_ADD_99_U81 );
not NOT1_7708 ( P1_ADD_99_U12 , P1_REG3_REG_7_ );
nand NAND2_7709 ( P1_ADD_99_U13 , P1_REG3_REG_7_ , P1_ADD_99_U82 );
not NOT1_7710 ( P1_ADD_99_U14 , P1_REG3_REG_8_ );
not NOT1_7711 ( P1_ADD_99_U15 , P1_REG3_REG_9_ );
nand NAND2_7712 ( P1_ADD_99_U16 , P1_REG3_REG_8_ , P1_ADD_99_U83 );
nand NAND2_7713 ( P1_ADD_99_U17 , P1_ADD_99_U84 , P1_REG3_REG_9_ );
not NOT1_7714 ( P1_ADD_99_U18 , P1_REG3_REG_10_ );
nand NAND2_7715 ( P1_ADD_99_U19 , P1_REG3_REG_10_ , P1_ADD_99_U85 );
not NOT1_7716 ( P1_ADD_99_U20 , P1_REG3_REG_11_ );
nand NAND2_7717 ( P1_ADD_99_U21 , P1_REG3_REG_11_ , P1_ADD_99_U86 );
not NOT1_7718 ( P1_ADD_99_U22 , P1_REG3_REG_12_ );
nand NAND2_7719 ( P1_ADD_99_U23 , P1_REG3_REG_12_ , P1_ADD_99_U87 );
not NOT1_7720 ( P1_ADD_99_U24 , P1_REG3_REG_13_ );
nand NAND2_7721 ( P1_ADD_99_U25 , P1_REG3_REG_13_ , P1_ADD_99_U88 );
not NOT1_7722 ( P1_ADD_99_U26 , P1_REG3_REG_14_ );
nand NAND2_7723 ( P1_ADD_99_U27 , P1_REG3_REG_14_ , P1_ADD_99_U89 );
not NOT1_7724 ( P1_ADD_99_U28 , P1_REG3_REG_15_ );
nand NAND2_7725 ( P1_ADD_99_U29 , P1_REG3_REG_15_ , P1_ADD_99_U90 );
not NOT1_7726 ( P1_ADD_99_U30 , P1_REG3_REG_16_ );
nand NAND2_7727 ( P1_ADD_99_U31 , P1_REG3_REG_16_ , P1_ADD_99_U91 );
not NOT1_7728 ( P1_ADD_99_U32 , P1_REG3_REG_17_ );
nand NAND2_7729 ( P1_ADD_99_U33 , P1_REG3_REG_17_ , P1_ADD_99_U92 );
not NOT1_7730 ( P1_ADD_99_U34 , P1_REG3_REG_18_ );
nand NAND2_7731 ( P1_ADD_99_U35 , P1_REG3_REG_18_ , P1_ADD_99_U93 );
not NOT1_7732 ( P1_ADD_99_U36 , P1_REG3_REG_19_ );
nand NAND2_7733 ( P1_ADD_99_U37 , P1_REG3_REG_19_ , P1_ADD_99_U94 );
not NOT1_7734 ( P1_ADD_99_U38 , P1_REG3_REG_20_ );
nand NAND2_7735 ( P1_ADD_99_U39 , P1_REG3_REG_20_ , P1_ADD_99_U95 );
not NOT1_7736 ( P1_ADD_99_U40 , P1_REG3_REG_21_ );
nand NAND2_7737 ( P1_ADD_99_U41 , P1_REG3_REG_21_ , P1_ADD_99_U96 );
not NOT1_7738 ( P1_ADD_99_U42 , P1_REG3_REG_22_ );
nand NAND2_7739 ( P1_ADD_99_U43 , P1_REG3_REG_22_ , P1_ADD_99_U97 );
not NOT1_7740 ( P1_ADD_99_U44 , P1_REG3_REG_23_ );
nand NAND2_7741 ( P1_ADD_99_U45 , P1_REG3_REG_23_ , P1_ADD_99_U98 );
not NOT1_7742 ( P1_ADD_99_U46 , P1_REG3_REG_24_ );
nand NAND2_7743 ( P1_ADD_99_U47 , P1_REG3_REG_24_ , P1_ADD_99_U99 );
not NOT1_7744 ( P1_ADD_99_U48 , P1_REG3_REG_25_ );
nand NAND2_7745 ( P1_ADD_99_U49 , P1_REG3_REG_25_ , P1_ADD_99_U100 );
not NOT1_7746 ( P1_ADD_99_U50 , P1_REG3_REG_26_ );
nand NAND2_7747 ( P1_ADD_99_U51 , P1_REG3_REG_26_ , P1_ADD_99_U101 );
not NOT1_7748 ( P1_ADD_99_U52 , P1_REG3_REG_28_ );
not NOT1_7749 ( P1_ADD_99_U53 , P1_REG3_REG_27_ );
nand NAND2_7750 ( P1_ADD_99_U54 , P1_ADD_99_U105 , P1_ADD_99_U104 );
nand NAND2_7751 ( P1_ADD_99_U55 , P1_ADD_99_U107 , P1_ADD_99_U106 );
nand NAND2_7752 ( P1_ADD_99_U56 , P1_ADD_99_U109 , P1_ADD_99_U108 );
nand NAND2_7753 ( P1_ADD_99_U57 , P1_ADD_99_U111 , P1_ADD_99_U110 );
nand NAND2_7754 ( P1_ADD_99_U58 , P1_ADD_99_U113 , P1_ADD_99_U112 );
nand NAND2_7755 ( P1_ADD_99_U59 , P1_ADD_99_U115 , P1_ADD_99_U114 );
nand NAND2_7756 ( P1_ADD_99_U60 , P1_ADD_99_U117 , P1_ADD_99_U116 );
nand NAND2_7757 ( P1_ADD_99_U61 , P1_ADD_99_U119 , P1_ADD_99_U118 );
nand NAND2_7758 ( P1_ADD_99_U62 , P1_ADD_99_U121 , P1_ADD_99_U120 );
nand NAND2_7759 ( P1_ADD_99_U63 , P1_ADD_99_U123 , P1_ADD_99_U122 );
nand NAND2_7760 ( P1_ADD_99_U64 , P1_ADD_99_U125 , P1_ADD_99_U124 );
nand NAND2_7761 ( P1_ADD_99_U65 , P1_ADD_99_U127 , P1_ADD_99_U126 );
nand NAND2_7762 ( P1_ADD_99_U66 , P1_ADD_99_U129 , P1_ADD_99_U128 );
nand NAND2_7763 ( P1_ADD_99_U67 , P1_ADD_99_U131 , P1_ADD_99_U130 );
nand NAND2_7764 ( P1_ADD_99_U68 , P1_ADD_99_U133 , P1_ADD_99_U132 );
nand NAND2_7765 ( P1_ADD_99_U69 , P1_ADD_99_U135 , P1_ADD_99_U134 );
nand NAND2_7766 ( P1_ADD_99_U70 , P1_ADD_99_U137 , P1_ADD_99_U136 );
nand NAND2_7767 ( P1_ADD_99_U71 , P1_ADD_99_U139 , P1_ADD_99_U138 );
nand NAND2_7768 ( P1_ADD_99_U72 , P1_ADD_99_U141 , P1_ADD_99_U140 );
nand NAND2_7769 ( P1_ADD_99_U73 , P1_ADD_99_U143 , P1_ADD_99_U142 );
nand NAND2_7770 ( P1_ADD_99_U74 , P1_ADD_99_U145 , P1_ADD_99_U144 );
nand NAND2_7771 ( P1_ADD_99_U75 , P1_ADD_99_U147 , P1_ADD_99_U146 );
nand NAND2_7772 ( P1_ADD_99_U76 , P1_ADD_99_U149 , P1_ADD_99_U148 );
nand NAND2_7773 ( P1_ADD_99_U77 , P1_ADD_99_U151 , P1_ADD_99_U150 );
nand NAND2_7774 ( P1_ADD_99_U78 , P1_ADD_99_U153 , P1_ADD_99_U152 );
nand NAND2_7775 ( P1_ADD_99_U79 , P1_REG3_REG_27_ , P1_ADD_99_U102 );
not NOT1_7776 ( P1_ADD_99_U80 , P1_ADD_99_U7 );
not NOT1_7777 ( P1_ADD_99_U81 , P1_ADD_99_U9 );
not NOT1_7778 ( P1_ADD_99_U82 , P1_ADD_99_U11 );
not NOT1_7779 ( P1_ADD_99_U83 , P1_ADD_99_U13 );
not NOT1_7780 ( P1_ADD_99_U84 , P1_ADD_99_U16 );
not NOT1_7781 ( P1_ADD_99_U85 , P1_ADD_99_U17 );
not NOT1_7782 ( P1_ADD_99_U86 , P1_ADD_99_U19 );
not NOT1_7783 ( P1_ADD_99_U87 , P1_ADD_99_U21 );
not NOT1_7784 ( P1_ADD_99_U88 , P1_ADD_99_U23 );
not NOT1_7785 ( P1_ADD_99_U89 , P1_ADD_99_U25 );
not NOT1_7786 ( P1_ADD_99_U90 , P1_ADD_99_U27 );
not NOT1_7787 ( P1_ADD_99_U91 , P1_ADD_99_U29 );
not NOT1_7788 ( P1_ADD_99_U92 , P1_ADD_99_U31 );
not NOT1_7789 ( P1_ADD_99_U93 , P1_ADD_99_U33 );
not NOT1_7790 ( P1_ADD_99_U94 , P1_ADD_99_U35 );
not NOT1_7791 ( P1_ADD_99_U95 , P1_ADD_99_U37 );
not NOT1_7792 ( P1_ADD_99_U96 , P1_ADD_99_U39 );
not NOT1_7793 ( P1_ADD_99_U97 , P1_ADD_99_U41 );
not NOT1_7794 ( P1_ADD_99_U98 , P1_ADD_99_U43 );
not NOT1_7795 ( P1_ADD_99_U99 , P1_ADD_99_U45 );
not NOT1_7796 ( P1_ADD_99_U100 , P1_ADD_99_U47 );
not NOT1_7797 ( P1_ADD_99_U101 , P1_ADD_99_U49 );
not NOT1_7798 ( P1_ADD_99_U102 , P1_ADD_99_U51 );
not NOT1_7799 ( P1_ADD_99_U103 , P1_ADD_99_U79 );
nand NAND2_7800 ( P1_ADD_99_U104 , P1_REG3_REG_9_ , P1_ADD_99_U16 );
nand NAND2_7801 ( P1_ADD_99_U105 , P1_ADD_99_U84 , P1_ADD_99_U15 );
nand NAND2_7802 ( P1_ADD_99_U106 , P1_REG3_REG_8_ , P1_ADD_99_U13 );
nand NAND2_7803 ( P1_ADD_99_U107 , P1_ADD_99_U83 , P1_ADD_99_U14 );
nand NAND2_7804 ( P1_ADD_99_U108 , P1_REG3_REG_7_ , P1_ADD_99_U11 );
nand NAND2_7805 ( P1_ADD_99_U109 , P1_ADD_99_U82 , P1_ADD_99_U12 );
nand NAND2_7806 ( P1_ADD_99_U110 , P1_REG3_REG_6_ , P1_ADD_99_U9 );
nand NAND2_7807 ( P1_ADD_99_U111 , P1_ADD_99_U81 , P1_ADD_99_U10 );
nand NAND2_7808 ( P1_ADD_99_U112 , P1_REG3_REG_5_ , P1_ADD_99_U7 );
nand NAND2_7809 ( P1_ADD_99_U113 , P1_ADD_99_U80 , P1_ADD_99_U8 );
nand NAND2_7810 ( P1_ADD_99_U114 , P1_REG3_REG_4_ , P1_ADD_99_U4 );
nand NAND2_7811 ( P1_ADD_99_U115 , P1_REG3_REG_3_ , P1_ADD_99_U6 );
nand NAND2_7812 ( P1_ADD_99_U116 , P1_REG3_REG_28_ , P1_ADD_99_U79 );
nand NAND2_7813 ( P1_ADD_99_U117 , P1_ADD_99_U103 , P1_ADD_99_U52 );
nand NAND2_7814 ( P1_ADD_99_U118 , P1_REG3_REG_27_ , P1_ADD_99_U51 );
nand NAND2_7815 ( P1_ADD_99_U119 , P1_ADD_99_U102 , P1_ADD_99_U53 );
nand NAND2_7816 ( P1_ADD_99_U120 , P1_REG3_REG_26_ , P1_ADD_99_U49 );
nand NAND2_7817 ( P1_ADD_99_U121 , P1_ADD_99_U101 , P1_ADD_99_U50 );
nand NAND2_7818 ( P1_ADD_99_U122 , P1_REG3_REG_25_ , P1_ADD_99_U47 );
nand NAND2_7819 ( P1_ADD_99_U123 , P1_ADD_99_U100 , P1_ADD_99_U48 );
nand NAND2_7820 ( P1_ADD_99_U124 , P1_REG3_REG_24_ , P1_ADD_99_U45 );
nand NAND2_7821 ( P1_ADD_99_U125 , P1_ADD_99_U99 , P1_ADD_99_U46 );
nand NAND2_7822 ( P1_ADD_99_U126 , P1_REG3_REG_23_ , P1_ADD_99_U43 );
nand NAND2_7823 ( P1_ADD_99_U127 , P1_ADD_99_U98 , P1_ADD_99_U44 );
nand NAND2_7824 ( P1_ADD_99_U128 , P1_REG3_REG_22_ , P1_ADD_99_U41 );
nand NAND2_7825 ( P1_ADD_99_U129 , P1_ADD_99_U97 , P1_ADD_99_U42 );
nand NAND2_7826 ( P1_ADD_99_U130 , P1_REG3_REG_21_ , P1_ADD_99_U39 );
nand NAND2_7827 ( P1_ADD_99_U131 , P1_ADD_99_U96 , P1_ADD_99_U40 );
nand NAND2_7828 ( P1_ADD_99_U132 , P1_REG3_REG_20_ , P1_ADD_99_U37 );
nand NAND2_7829 ( P1_ADD_99_U133 , P1_ADD_99_U95 , P1_ADD_99_U38 );
nand NAND2_7830 ( P1_ADD_99_U134 , P1_REG3_REG_19_ , P1_ADD_99_U35 );
nand NAND2_7831 ( P1_ADD_99_U135 , P1_ADD_99_U94 , P1_ADD_99_U36 );
nand NAND2_7832 ( P1_ADD_99_U136 , P1_REG3_REG_18_ , P1_ADD_99_U33 );
nand NAND2_7833 ( P1_ADD_99_U137 , P1_ADD_99_U93 , P1_ADD_99_U34 );
nand NAND2_7834 ( P1_ADD_99_U138 , P1_REG3_REG_17_ , P1_ADD_99_U31 );
nand NAND2_7835 ( P1_ADD_99_U139 , P1_ADD_99_U92 , P1_ADD_99_U32 );
nand NAND2_7836 ( P1_ADD_99_U140 , P1_REG3_REG_16_ , P1_ADD_99_U29 );
nand NAND2_7837 ( P1_ADD_99_U141 , P1_ADD_99_U91 , P1_ADD_99_U30 );
nand NAND2_7838 ( P1_ADD_99_U142 , P1_REG3_REG_15_ , P1_ADD_99_U27 );
nand NAND2_7839 ( P1_ADD_99_U143 , P1_ADD_99_U90 , P1_ADD_99_U28 );
nand NAND2_7840 ( P1_ADD_99_U144 , P1_REG3_REG_14_ , P1_ADD_99_U25 );
nand NAND2_7841 ( P1_ADD_99_U145 , P1_ADD_99_U89 , P1_ADD_99_U26 );
nand NAND2_7842 ( P1_ADD_99_U146 , P1_REG3_REG_13_ , P1_ADD_99_U23 );
nand NAND2_7843 ( P1_ADD_99_U147 , P1_ADD_99_U88 , P1_ADD_99_U24 );
nand NAND2_7844 ( P1_ADD_99_U148 , P1_REG3_REG_12_ , P1_ADD_99_U21 );
nand NAND2_7845 ( P1_ADD_99_U149 , P1_ADD_99_U87 , P1_ADD_99_U22 );
nand NAND2_7846 ( P1_ADD_99_U150 , P1_REG3_REG_11_ , P1_ADD_99_U19 );
nand NAND2_7847 ( P1_ADD_99_U151 , P1_ADD_99_U86 , P1_ADD_99_U20 );
nand NAND2_7848 ( P1_ADD_99_U152 , P1_REG3_REG_10_ , P1_ADD_99_U17 );
nand NAND2_7849 ( P1_ADD_99_U153 , P1_ADD_99_U85 , P1_ADD_99_U18 );
and AND2_7850 ( P1_R1105_U4 , P1_R1105_U95 , P1_R1105_U94 );
and AND2_7851 ( P1_R1105_U5 , P1_R1105_U96 , P1_R1105_U97 );
and AND2_7852 ( P1_R1105_U6 , P1_R1105_U113 , P1_R1105_U112 );
and AND2_7853 ( P1_R1105_U7 , P1_R1105_U155 , P1_R1105_U154 );
and AND2_7854 ( P1_R1105_U8 , P1_R1105_U164 , P1_R1105_U163 );
and AND2_7855 ( P1_R1105_U9 , P1_R1105_U182 , P1_R1105_U181 );
and AND2_7856 ( P1_R1105_U10 , P1_R1105_U218 , P1_R1105_U215 );
and AND2_7857 ( P1_R1105_U11 , P1_R1105_U211 , P1_R1105_U208 );
and AND2_7858 ( P1_R1105_U12 , P1_R1105_U202 , P1_R1105_U199 );
and AND2_7859 ( P1_R1105_U13 , P1_R1105_U196 , P1_R1105_U192 );
and AND2_7860 ( P1_R1105_U14 , P1_R1105_U151 , P1_R1105_U148 );
and AND2_7861 ( P1_R1105_U15 , P1_R1105_U143 , P1_R1105_U140 );
and AND2_7862 ( P1_R1105_U16 , P1_R1105_U129 , P1_R1105_U126 );
not NOT1_7863 ( P1_R1105_U17 , P1_REG2_REG_6_ );
not NOT1_7864 ( P1_R1105_U18 , P1_U3470 );
not NOT1_7865 ( P1_R1105_U19 , P1_U3473 );
nand NAND2_7866 ( P1_R1105_U20 , P1_U3470 , P1_REG2_REG_6_ );
not NOT1_7867 ( P1_R1105_U21 , P1_REG2_REG_7_ );
not NOT1_7868 ( P1_R1105_U22 , P1_REG2_REG_4_ );
not NOT1_7869 ( P1_R1105_U23 , P1_U3464 );
not NOT1_7870 ( P1_R1105_U24 , P1_U3467 );
not NOT1_7871 ( P1_R1105_U25 , P1_REG2_REG_2_ );
not NOT1_7872 ( P1_R1105_U26 , P1_U3458 );
not NOT1_7873 ( P1_R1105_U27 , P1_REG2_REG_0_ );
not NOT1_7874 ( P1_R1105_U28 , P1_U3449 );
nand NAND2_7875 ( P1_R1105_U29 , P1_U3449 , P1_REG2_REG_0_ );
not NOT1_7876 ( P1_R1105_U30 , P1_REG2_REG_3_ );
not NOT1_7877 ( P1_R1105_U31 , P1_U3461 );
nand NAND2_7878 ( P1_R1105_U32 , P1_U3464 , P1_REG2_REG_4_ );
not NOT1_7879 ( P1_R1105_U33 , P1_REG2_REG_5_ );
not NOT1_7880 ( P1_R1105_U34 , P1_REG2_REG_8_ );
not NOT1_7881 ( P1_R1105_U35 , P1_U3476 );
not NOT1_7882 ( P1_R1105_U36 , P1_U3479 );
not NOT1_7883 ( P1_R1105_U37 , P1_REG2_REG_9_ );
nand NAND2_7884 ( P1_R1105_U38 , P1_R1105_U49 , P1_R1105_U121 );
nand NAND3_7885 ( P1_R1105_U39 , P1_R1105_U110 , P1_R1105_U108 , P1_R1105_U109 );
nand NAND2_7886 ( P1_R1105_U40 , P1_R1105_U98 , P1_R1105_U99 );
nand NAND2_7887 ( P1_R1105_U41 , P1_REG2_REG_1_ , P1_U3455 );
nand NAND3_7888 ( P1_R1105_U42 , P1_R1105_U136 , P1_R1105_U134 , P1_R1105_U135 );
nand NAND2_7889 ( P1_R1105_U43 , P1_R1105_U132 , P1_R1105_U131 );
not NOT1_7890 ( P1_R1105_U44 , P1_REG2_REG_16_ );
not NOT1_7891 ( P1_R1105_U45 , P1_U3500 );
not NOT1_7892 ( P1_R1105_U46 , P1_U3503 );
nand NAND2_7893 ( P1_R1105_U47 , P1_U3500 , P1_REG2_REG_16_ );
not NOT1_7894 ( P1_R1105_U48 , P1_REG2_REG_17_ );
nand NAND2_7895 ( P1_R1105_U49 , P1_U3476 , P1_REG2_REG_8_ );
not NOT1_7896 ( P1_R1105_U50 , P1_REG2_REG_10_ );
not NOT1_7897 ( P1_R1105_U51 , P1_U3482 );
not NOT1_7898 ( P1_R1105_U52 , P1_REG2_REG_12_ );
not NOT1_7899 ( P1_R1105_U53 , P1_U3488 );
not NOT1_7900 ( P1_R1105_U54 , P1_REG2_REG_11_ );
not NOT1_7901 ( P1_R1105_U55 , P1_U3485 );
nand NAND2_7902 ( P1_R1105_U56 , P1_U3485 , P1_REG2_REG_11_ );
not NOT1_7903 ( P1_R1105_U57 , P1_REG2_REG_13_ );
not NOT1_7904 ( P1_R1105_U58 , P1_U3491 );
not NOT1_7905 ( P1_R1105_U59 , P1_REG2_REG_14_ );
not NOT1_7906 ( P1_R1105_U60 , P1_U3494 );
not NOT1_7907 ( P1_R1105_U61 , P1_REG2_REG_15_ );
not NOT1_7908 ( P1_R1105_U62 , P1_U3497 );
not NOT1_7909 ( P1_R1105_U63 , P1_REG2_REG_18_ );
not NOT1_7910 ( P1_R1105_U64 , P1_U3506 );
nand NAND3_7911 ( P1_R1105_U65 , P1_R1105_U186 , P1_R1105_U185 , P1_R1105_U187 );
nand NAND2_7912 ( P1_R1105_U66 , P1_R1105_U179 , P1_R1105_U178 );
nand NAND2_7913 ( P1_R1105_U67 , P1_R1105_U56 , P1_R1105_U204 );
nand NAND2_7914 ( P1_R1105_U68 , P1_R1105_U259 , P1_R1105_U258 );
nand NAND2_7915 ( P1_R1105_U69 , P1_R1105_U308 , P1_R1105_U307 );
nand NAND2_7916 ( P1_R1105_U70 , P1_R1105_U231 , P1_R1105_U230 );
nand NAND2_7917 ( P1_R1105_U71 , P1_R1105_U236 , P1_R1105_U235 );
nand NAND2_7918 ( P1_R1105_U72 , P1_R1105_U243 , P1_R1105_U242 );
nand NAND2_7919 ( P1_R1105_U73 , P1_R1105_U250 , P1_R1105_U249 );
nand NAND2_7920 ( P1_R1105_U74 , P1_R1105_U255 , P1_R1105_U254 );
nand NAND2_7921 ( P1_R1105_U75 , P1_R1105_U271 , P1_R1105_U270 );
nand NAND2_7922 ( P1_R1105_U76 , P1_R1105_U278 , P1_R1105_U277 );
nand NAND2_7923 ( P1_R1105_U77 , P1_R1105_U285 , P1_R1105_U284 );
nand NAND2_7924 ( P1_R1105_U78 , P1_R1105_U292 , P1_R1105_U291 );
nand NAND2_7925 ( P1_R1105_U79 , P1_R1105_U299 , P1_R1105_U298 );
nand NAND2_7926 ( P1_R1105_U80 , P1_R1105_U304 , P1_R1105_U303 );
nand NAND3_7927 ( P1_R1105_U81 , P1_R1105_U117 , P1_R1105_U116 , P1_R1105_U118 );
nand NAND2_7928 ( P1_R1105_U82 , P1_R1105_U133 , P1_R1105_U145 );
nand NAND2_7929 ( P1_R1105_U83 , P1_R1105_U41 , P1_R1105_U152 );
not NOT1_7930 ( P1_R1105_U84 , P1_U3443 );
not NOT1_7931 ( P1_R1105_U85 , P1_REG2_REG_19_ );
nand NAND2_7932 ( P1_R1105_U86 , P1_R1105_U175 , P1_R1105_U174 );
nand NAND2_7933 ( P1_R1105_U87 , P1_R1105_U171 , P1_R1105_U170 );
nand NAND2_7934 ( P1_R1105_U88 , P1_R1105_U161 , P1_R1105_U160 );
not NOT1_7935 ( P1_R1105_U89 , P1_R1105_U32 );
nand NAND2_7936 ( P1_R1105_U90 , P1_REG2_REG_9_ , P1_U3479 );
nand NAND2_7937 ( P1_R1105_U91 , P1_U3488 , P1_REG2_REG_12_ );
not NOT1_7938 ( P1_R1105_U92 , P1_R1105_U56 );
not NOT1_7939 ( P1_R1105_U93 , P1_R1105_U49 );
or OR2_7940 ( P1_R1105_U94 , P1_U3467 , P1_REG2_REG_5_ );
or OR2_7941 ( P1_R1105_U95 , P1_U3464 , P1_REG2_REG_4_ );
or OR2_7942 ( P1_R1105_U96 , P1_REG2_REG_3_ , P1_U3461 );
or OR2_7943 ( P1_R1105_U97 , P1_REG2_REG_2_ , P1_U3458 );
not NOT1_7944 ( P1_R1105_U98 , P1_R1105_U29 );
or OR2_7945 ( P1_R1105_U99 , P1_REG2_REG_1_ , P1_U3455 );
not NOT1_7946 ( P1_R1105_U100 , P1_R1105_U40 );
not NOT1_7947 ( P1_R1105_U101 , P1_R1105_U41 );
nand NAND2_7948 ( P1_R1105_U102 , P1_R1105_U40 , P1_R1105_U41 );
nand NAND3_7949 ( P1_R1105_U103 , P1_REG2_REG_2_ , P1_U3458 , P1_R1105_U96 );
nand NAND2_7950 ( P1_R1105_U104 , P1_R1105_U5 , P1_R1105_U102 );
nand NAND2_7951 ( P1_R1105_U105 , P1_U3461 , P1_REG2_REG_3_ );
nand NAND3_7952 ( P1_R1105_U106 , P1_R1105_U105 , P1_R1105_U103 , P1_R1105_U104 );
nand NAND2_7953 ( P1_R1105_U107 , P1_R1105_U33 , P1_R1105_U32 );
nand NAND2_7954 ( P1_R1105_U108 , P1_U3467 , P1_R1105_U107 );
nand NAND2_7955 ( P1_R1105_U109 , P1_R1105_U4 , P1_R1105_U106 );
nand NAND2_7956 ( P1_R1105_U110 , P1_REG2_REG_5_ , P1_R1105_U89 );
not NOT1_7957 ( P1_R1105_U111 , P1_R1105_U39 );
or OR2_7958 ( P1_R1105_U112 , P1_U3473 , P1_REG2_REG_7_ );
or OR2_7959 ( P1_R1105_U113 , P1_U3470 , P1_REG2_REG_6_ );
not NOT1_7960 ( P1_R1105_U114 , P1_R1105_U20 );
nand NAND2_7961 ( P1_R1105_U115 , P1_R1105_U21 , P1_R1105_U20 );
nand NAND2_7962 ( P1_R1105_U116 , P1_U3473 , P1_R1105_U115 );
nand NAND2_7963 ( P1_R1105_U117 , P1_REG2_REG_7_ , P1_R1105_U114 );
nand NAND2_7964 ( P1_R1105_U118 , P1_R1105_U6 , P1_R1105_U39 );
not NOT1_7965 ( P1_R1105_U119 , P1_R1105_U81 );
or OR2_7966 ( P1_R1105_U120 , P1_REG2_REG_8_ , P1_U3476 );
nand NAND2_7967 ( P1_R1105_U121 , P1_R1105_U120 , P1_R1105_U81 );
not NOT1_7968 ( P1_R1105_U122 , P1_R1105_U38 );
or OR2_7969 ( P1_R1105_U123 , P1_U3479 , P1_REG2_REG_9_ );
or OR2_7970 ( P1_R1105_U124 , P1_REG2_REG_6_ , P1_U3470 );
nand NAND2_7971 ( P1_R1105_U125 , P1_R1105_U124 , P1_R1105_U39 );
nand NAND4_7972 ( P1_R1105_U126 , P1_R1105_U238 , P1_R1105_U237 , P1_R1105_U20 , P1_R1105_U125 );
nand NAND2_7973 ( P1_R1105_U127 , P1_R1105_U111 , P1_R1105_U20 );
nand NAND2_7974 ( P1_R1105_U128 , P1_REG2_REG_7_ , P1_U3473 );
nand NAND3_7975 ( P1_R1105_U129 , P1_R1105_U128 , P1_R1105_U6 , P1_R1105_U127 );
or OR2_7976 ( P1_R1105_U130 , P1_U3470 , P1_REG2_REG_6_ );
nand NAND2_7977 ( P1_R1105_U131 , P1_R1105_U101 , P1_R1105_U97 );
nand NAND2_7978 ( P1_R1105_U132 , P1_U3458 , P1_REG2_REG_2_ );
not NOT1_7979 ( P1_R1105_U133 , P1_R1105_U43 );
nand NAND2_7980 ( P1_R1105_U134 , P1_R1105_U100 , P1_R1105_U5 );
nand NAND2_7981 ( P1_R1105_U135 , P1_R1105_U43 , P1_R1105_U96 );
nand NAND2_7982 ( P1_R1105_U136 , P1_U3461 , P1_REG2_REG_3_ );
not NOT1_7983 ( P1_R1105_U137 , P1_R1105_U42 );
or OR2_7984 ( P1_R1105_U138 , P1_REG2_REG_4_ , P1_U3464 );
nand NAND2_7985 ( P1_R1105_U139 , P1_R1105_U138 , P1_R1105_U42 );
nand NAND4_7986 ( P1_R1105_U140 , P1_R1105_U245 , P1_R1105_U244 , P1_R1105_U32 , P1_R1105_U139 );
nand NAND2_7987 ( P1_R1105_U141 , P1_R1105_U137 , P1_R1105_U32 );
nand NAND2_7988 ( P1_R1105_U142 , P1_REG2_REG_5_ , P1_U3467 );
nand NAND3_7989 ( P1_R1105_U143 , P1_R1105_U142 , P1_R1105_U4 , P1_R1105_U141 );
or OR2_7990 ( P1_R1105_U144 , P1_U3464 , P1_REG2_REG_4_ );
nand NAND2_7991 ( P1_R1105_U145 , P1_R1105_U100 , P1_R1105_U97 );
not NOT1_7992 ( P1_R1105_U146 , P1_R1105_U82 );
nand NAND2_7993 ( P1_R1105_U147 , P1_U3461 , P1_REG2_REG_3_ );
nand NAND4_7994 ( P1_R1105_U148 , P1_R1105_U41 , P1_R1105_U40 , P1_R1105_U257 , P1_R1105_U256 );
nand NAND2_7995 ( P1_R1105_U149 , P1_R1105_U41 , P1_R1105_U40 );
nand NAND2_7996 ( P1_R1105_U150 , P1_U3458 , P1_REG2_REG_2_ );
nand NAND3_7997 ( P1_R1105_U151 , P1_R1105_U150 , P1_R1105_U97 , P1_R1105_U149 );
or OR2_7998 ( P1_R1105_U152 , P1_REG2_REG_1_ , P1_U3455 );
not NOT1_7999 ( P1_R1105_U153 , P1_R1105_U83 );
or OR2_8000 ( P1_R1105_U154 , P1_U3479 , P1_REG2_REG_9_ );
or OR2_8001 ( P1_R1105_U155 , P1_U3482 , P1_REG2_REG_10_ );
nand NAND2_8002 ( P1_R1105_U156 , P1_R1105_U93 , P1_R1105_U7 );
nand NAND2_8003 ( P1_R1105_U157 , P1_U3482 , P1_REG2_REG_10_ );
nand NAND3_8004 ( P1_R1105_U158 , P1_R1105_U157 , P1_R1105_U90 , P1_R1105_U156 );
or OR2_8005 ( P1_R1105_U159 , P1_REG2_REG_10_ , P1_U3482 );
nand NAND3_8006 ( P1_R1105_U160 , P1_R1105_U120 , P1_R1105_U7 , P1_R1105_U81 );
nand NAND2_8007 ( P1_R1105_U161 , P1_R1105_U159 , P1_R1105_U158 );
not NOT1_8008 ( P1_R1105_U162 , P1_R1105_U88 );
or OR2_8009 ( P1_R1105_U163 , P1_U3491 , P1_REG2_REG_13_ );
or OR2_8010 ( P1_R1105_U164 , P1_U3488 , P1_REG2_REG_12_ );
nand NAND2_8011 ( P1_R1105_U165 , P1_R1105_U92 , P1_R1105_U8 );
nand NAND2_8012 ( P1_R1105_U166 , P1_U3491 , P1_REG2_REG_13_ );
nand NAND3_8013 ( P1_R1105_U167 , P1_R1105_U166 , P1_R1105_U91 , P1_R1105_U165 );
or OR2_8014 ( P1_R1105_U168 , P1_REG2_REG_11_ , P1_U3485 );
or OR2_8015 ( P1_R1105_U169 , P1_REG2_REG_13_ , P1_U3491 );
nand NAND3_8016 ( P1_R1105_U170 , P1_R1105_U168 , P1_R1105_U8 , P1_R1105_U88 );
nand NAND2_8017 ( P1_R1105_U171 , P1_R1105_U169 , P1_R1105_U167 );
not NOT1_8018 ( P1_R1105_U172 , P1_R1105_U87 );
or OR2_8019 ( P1_R1105_U173 , P1_REG2_REG_14_ , P1_U3494 );
nand NAND2_8020 ( P1_R1105_U174 , P1_R1105_U173 , P1_R1105_U87 );
nand NAND2_8021 ( P1_R1105_U175 , P1_U3494 , P1_REG2_REG_14_ );
not NOT1_8022 ( P1_R1105_U176 , P1_R1105_U86 );
or OR2_8023 ( P1_R1105_U177 , P1_REG2_REG_15_ , P1_U3497 );
nand NAND2_8024 ( P1_R1105_U178 , P1_R1105_U177 , P1_R1105_U86 );
nand NAND2_8025 ( P1_R1105_U179 , P1_U3497 , P1_REG2_REG_15_ );
not NOT1_8026 ( P1_R1105_U180 , P1_R1105_U66 );
or OR2_8027 ( P1_R1105_U181 , P1_U3503 , P1_REG2_REG_17_ );
or OR2_8028 ( P1_R1105_U182 , P1_U3500 , P1_REG2_REG_16_ );
not NOT1_8029 ( P1_R1105_U183 , P1_R1105_U47 );
nand NAND2_8030 ( P1_R1105_U184 , P1_R1105_U48 , P1_R1105_U47 );
nand NAND2_8031 ( P1_R1105_U185 , P1_U3503 , P1_R1105_U184 );
nand NAND2_8032 ( P1_R1105_U186 , P1_REG2_REG_17_ , P1_R1105_U183 );
nand NAND2_8033 ( P1_R1105_U187 , P1_R1105_U9 , P1_R1105_U66 );
not NOT1_8034 ( P1_R1105_U188 , P1_R1105_U65 );
or OR2_8035 ( P1_R1105_U189 , P1_REG2_REG_18_ , P1_U3506 );
nand NAND2_8036 ( P1_R1105_U190 , P1_R1105_U189 , P1_R1105_U65 );
nand NAND2_8037 ( P1_R1105_U191 , P1_U3506 , P1_REG2_REG_18_ );
nand NAND4_8038 ( P1_R1105_U192 , P1_R1105_U261 , P1_R1105_U260 , P1_R1105_U191 , P1_R1105_U190 );
nand NAND2_8039 ( P1_R1105_U193 , P1_U3506 , P1_REG2_REG_18_ );
nand NAND2_8040 ( P1_R1105_U194 , P1_R1105_U188 , P1_R1105_U193 );
or OR2_8041 ( P1_R1105_U195 , P1_U3506 , P1_REG2_REG_18_ );
nand NAND3_8042 ( P1_R1105_U196 , P1_R1105_U195 , P1_R1105_U264 , P1_R1105_U194 );
or OR2_8043 ( P1_R1105_U197 , P1_REG2_REG_16_ , P1_U3500 );
nand NAND2_8044 ( P1_R1105_U198 , P1_R1105_U197 , P1_R1105_U66 );
nand NAND4_8045 ( P1_R1105_U199 , P1_R1105_U273 , P1_R1105_U272 , P1_R1105_U47 , P1_R1105_U198 );
nand NAND2_8046 ( P1_R1105_U200 , P1_R1105_U180 , P1_R1105_U47 );
nand NAND2_8047 ( P1_R1105_U201 , P1_REG2_REG_17_ , P1_U3503 );
nand NAND3_8048 ( P1_R1105_U202 , P1_R1105_U201 , P1_R1105_U9 , P1_R1105_U200 );
or OR2_8049 ( P1_R1105_U203 , P1_U3500 , P1_REG2_REG_16_ );
nand NAND2_8050 ( P1_R1105_U204 , P1_R1105_U168 , P1_R1105_U88 );
not NOT1_8051 ( P1_R1105_U205 , P1_R1105_U67 );
or OR2_8052 ( P1_R1105_U206 , P1_REG2_REG_12_ , P1_U3488 );
nand NAND2_8053 ( P1_R1105_U207 , P1_R1105_U206 , P1_R1105_U67 );
nand NAND4_8054 ( P1_R1105_U208 , P1_R1105_U294 , P1_R1105_U293 , P1_R1105_U91 , P1_R1105_U207 );
nand NAND2_8055 ( P1_R1105_U209 , P1_R1105_U205 , P1_R1105_U91 );
nand NAND2_8056 ( P1_R1105_U210 , P1_U3491 , P1_REG2_REG_13_ );
nand NAND3_8057 ( P1_R1105_U211 , P1_R1105_U210 , P1_R1105_U8 , P1_R1105_U209 );
or OR2_8058 ( P1_R1105_U212 , P1_U3488 , P1_REG2_REG_12_ );
or OR2_8059 ( P1_R1105_U213 , P1_REG2_REG_9_ , P1_U3479 );
nand NAND2_8060 ( P1_R1105_U214 , P1_R1105_U213 , P1_R1105_U38 );
nand NAND4_8061 ( P1_R1105_U215 , P1_R1105_U306 , P1_R1105_U305 , P1_R1105_U90 , P1_R1105_U214 );
nand NAND2_8062 ( P1_R1105_U216 , P1_R1105_U122 , P1_R1105_U90 );
nand NAND2_8063 ( P1_R1105_U217 , P1_U3482 , P1_REG2_REG_10_ );
nand NAND3_8064 ( P1_R1105_U218 , P1_R1105_U217 , P1_R1105_U7 , P1_R1105_U216 );
nand NAND2_8065 ( P1_R1105_U219 , P1_R1105_U123 , P1_R1105_U90 );
nand NAND2_8066 ( P1_R1105_U220 , P1_R1105_U120 , P1_R1105_U49 );
nand NAND2_8067 ( P1_R1105_U221 , P1_R1105_U130 , P1_R1105_U20 );
nand NAND2_8068 ( P1_R1105_U222 , P1_R1105_U144 , P1_R1105_U32 );
nand NAND2_8069 ( P1_R1105_U223 , P1_R1105_U147 , P1_R1105_U96 );
nand NAND2_8070 ( P1_R1105_U224 , P1_R1105_U203 , P1_R1105_U47 );
nand NAND2_8071 ( P1_R1105_U225 , P1_R1105_U212 , P1_R1105_U91 );
nand NAND2_8072 ( P1_R1105_U226 , P1_R1105_U168 , P1_R1105_U56 );
nand NAND2_8073 ( P1_R1105_U227 , P1_U3479 , P1_R1105_U37 );
nand NAND2_8074 ( P1_R1105_U228 , P1_REG2_REG_9_ , P1_R1105_U36 );
nand NAND2_8075 ( P1_R1105_U229 , P1_R1105_U228 , P1_R1105_U227 );
nand NAND2_8076 ( P1_R1105_U230 , P1_R1105_U219 , P1_R1105_U38 );
nand NAND2_8077 ( P1_R1105_U231 , P1_R1105_U229 , P1_R1105_U122 );
nand NAND2_8078 ( P1_R1105_U232 , P1_U3476 , P1_R1105_U34 );
nand NAND2_8079 ( P1_R1105_U233 , P1_REG2_REG_8_ , P1_R1105_U35 );
nand NAND2_8080 ( P1_R1105_U234 , P1_R1105_U233 , P1_R1105_U232 );
nand NAND2_8081 ( P1_R1105_U235 , P1_R1105_U220 , P1_R1105_U81 );
nand NAND2_8082 ( P1_R1105_U236 , P1_R1105_U119 , P1_R1105_U234 );
nand NAND2_8083 ( P1_R1105_U237 , P1_U3473 , P1_R1105_U21 );
nand NAND2_8084 ( P1_R1105_U238 , P1_REG2_REG_7_ , P1_R1105_U19 );
nand NAND2_8085 ( P1_R1105_U239 , P1_U3470 , P1_R1105_U17 );
nand NAND2_8086 ( P1_R1105_U240 , P1_REG2_REG_6_ , P1_R1105_U18 );
nand NAND2_8087 ( P1_R1105_U241 , P1_R1105_U240 , P1_R1105_U239 );
nand NAND2_8088 ( P1_R1105_U242 , P1_R1105_U221 , P1_R1105_U39 );
nand NAND2_8089 ( P1_R1105_U243 , P1_R1105_U241 , P1_R1105_U111 );
nand NAND2_8090 ( P1_R1105_U244 , P1_U3467 , P1_R1105_U33 );
nand NAND2_8091 ( P1_R1105_U245 , P1_REG2_REG_5_ , P1_R1105_U24 );
nand NAND2_8092 ( P1_R1105_U246 , P1_U3464 , P1_R1105_U22 );
nand NAND2_8093 ( P1_R1105_U247 , P1_REG2_REG_4_ , P1_R1105_U23 );
nand NAND2_8094 ( P1_R1105_U248 , P1_R1105_U247 , P1_R1105_U246 );
nand NAND2_8095 ( P1_R1105_U249 , P1_R1105_U222 , P1_R1105_U42 );
nand NAND2_8096 ( P1_R1105_U250 , P1_R1105_U248 , P1_R1105_U137 );
nand NAND2_8097 ( P1_R1105_U251 , P1_U3461 , P1_R1105_U30 );
nand NAND2_8098 ( P1_R1105_U252 , P1_REG2_REG_3_ , P1_R1105_U31 );
nand NAND2_8099 ( P1_R1105_U253 , P1_R1105_U252 , P1_R1105_U251 );
nand NAND2_8100 ( P1_R1105_U254 , P1_R1105_U223 , P1_R1105_U82 );
nand NAND2_8101 ( P1_R1105_U255 , P1_R1105_U146 , P1_R1105_U253 );
nand NAND2_8102 ( P1_R1105_U256 , P1_U3458 , P1_R1105_U25 );
nand NAND2_8103 ( P1_R1105_U257 , P1_REG2_REG_2_ , P1_R1105_U26 );
nand NAND2_8104 ( P1_R1105_U258 , P1_R1105_U98 , P1_R1105_U83 );
nand NAND2_8105 ( P1_R1105_U259 , P1_R1105_U153 , P1_R1105_U29 );
nand NAND2_8106 ( P1_R1105_U260 , P1_U3443 , P1_R1105_U85 );
nand NAND2_8107 ( P1_R1105_U261 , P1_REG2_REG_19_ , P1_R1105_U84 );
nand NAND2_8108 ( P1_R1105_U262 , P1_U3443 , P1_R1105_U85 );
nand NAND2_8109 ( P1_R1105_U263 , P1_REG2_REG_19_ , P1_R1105_U84 );
nand NAND2_8110 ( P1_R1105_U264 , P1_R1105_U263 , P1_R1105_U262 );
nand NAND2_8111 ( P1_R1105_U265 , P1_U3506 , P1_R1105_U63 );
nand NAND2_8112 ( P1_R1105_U266 , P1_REG2_REG_18_ , P1_R1105_U64 );
nand NAND2_8113 ( P1_R1105_U267 , P1_U3506 , P1_R1105_U63 );
nand NAND2_8114 ( P1_R1105_U268 , P1_REG2_REG_18_ , P1_R1105_U64 );
nand NAND2_8115 ( P1_R1105_U269 , P1_R1105_U268 , P1_R1105_U267 );
nand NAND3_8116 ( P1_R1105_U270 , P1_R1105_U266 , P1_R1105_U265 , P1_R1105_U65 );
nand NAND2_8117 ( P1_R1105_U271 , P1_R1105_U269 , P1_R1105_U188 );
nand NAND2_8118 ( P1_R1105_U272 , P1_U3503 , P1_R1105_U48 );
nand NAND2_8119 ( P1_R1105_U273 , P1_REG2_REG_17_ , P1_R1105_U46 );
nand NAND2_8120 ( P1_R1105_U274 , P1_U3500 , P1_R1105_U44 );
nand NAND2_8121 ( P1_R1105_U275 , P1_REG2_REG_16_ , P1_R1105_U45 );
nand NAND2_8122 ( P1_R1105_U276 , P1_R1105_U275 , P1_R1105_U274 );
nand NAND2_8123 ( P1_R1105_U277 , P1_R1105_U224 , P1_R1105_U66 );
nand NAND2_8124 ( P1_R1105_U278 , P1_R1105_U276 , P1_R1105_U180 );
nand NAND2_8125 ( P1_R1105_U279 , P1_U3497 , P1_R1105_U61 );
nand NAND2_8126 ( P1_R1105_U280 , P1_REG2_REG_15_ , P1_R1105_U62 );
nand NAND2_8127 ( P1_R1105_U281 , P1_U3497 , P1_R1105_U61 );
nand NAND2_8128 ( P1_R1105_U282 , P1_REG2_REG_15_ , P1_R1105_U62 );
nand NAND2_8129 ( P1_R1105_U283 , P1_R1105_U282 , P1_R1105_U281 );
nand NAND3_8130 ( P1_R1105_U284 , P1_R1105_U280 , P1_R1105_U279 , P1_R1105_U86 );
nand NAND2_8131 ( P1_R1105_U285 , P1_R1105_U176 , P1_R1105_U283 );
nand NAND2_8132 ( P1_R1105_U286 , P1_U3494 , P1_R1105_U59 );
nand NAND2_8133 ( P1_R1105_U287 , P1_REG2_REG_14_ , P1_R1105_U60 );
nand NAND2_8134 ( P1_R1105_U288 , P1_U3494 , P1_R1105_U59 );
nand NAND2_8135 ( P1_R1105_U289 , P1_REG2_REG_14_ , P1_R1105_U60 );
nand NAND2_8136 ( P1_R1105_U290 , P1_R1105_U289 , P1_R1105_U288 );
nand NAND3_8137 ( P1_R1105_U291 , P1_R1105_U287 , P1_R1105_U286 , P1_R1105_U87 );
nand NAND2_8138 ( P1_R1105_U292 , P1_R1105_U172 , P1_R1105_U290 );
nand NAND2_8139 ( P1_R1105_U293 , P1_U3491 , P1_R1105_U57 );
nand NAND2_8140 ( P1_R1105_U294 , P1_REG2_REG_13_ , P1_R1105_U58 );
nand NAND2_8141 ( P1_R1105_U295 , P1_U3488 , P1_R1105_U52 );
nand NAND2_8142 ( P1_R1105_U296 , P1_REG2_REG_12_ , P1_R1105_U53 );
nand NAND2_8143 ( P1_R1105_U297 , P1_R1105_U296 , P1_R1105_U295 );
nand NAND2_8144 ( P1_R1105_U298 , P1_R1105_U225 , P1_R1105_U67 );
nand NAND2_8145 ( P1_R1105_U299 , P1_R1105_U297 , P1_R1105_U205 );
nand NAND2_8146 ( P1_R1105_U300 , P1_U3485 , P1_R1105_U54 );
nand NAND2_8147 ( P1_R1105_U301 , P1_REG2_REG_11_ , P1_R1105_U55 );
nand NAND2_8148 ( P1_R1105_U302 , P1_R1105_U301 , P1_R1105_U300 );
nand NAND2_8149 ( P1_R1105_U303 , P1_R1105_U226 , P1_R1105_U88 );
nand NAND2_8150 ( P1_R1105_U304 , P1_R1105_U162 , P1_R1105_U302 );
nand NAND2_8151 ( P1_R1105_U305 , P1_U3482 , P1_R1105_U50 );
nand NAND2_8152 ( P1_R1105_U306 , P1_REG2_REG_10_ , P1_R1105_U51 );
nand NAND2_8153 ( P1_R1105_U307 , P1_U3449 , P1_R1105_U27 );
nand NAND2_8154 ( P1_R1105_U308 , P1_REG2_REG_0_ , P1_R1105_U28 );
and AND2_8155 ( P1_SUB_88_U6 , P1_SUB_88_U227 , P1_SUB_88_U38 );
and AND2_8156 ( P1_SUB_88_U7 , P1_SUB_88_U225 , P1_SUB_88_U192 );
and AND2_8157 ( P1_SUB_88_U8 , P1_SUB_88_U224 , P1_SUB_88_U35 );
and AND2_8158 ( P1_SUB_88_U9 , P1_SUB_88_U223 , P1_SUB_88_U36 );
and AND2_8159 ( P1_SUB_88_U10 , P1_SUB_88_U221 , P1_SUB_88_U195 );
and AND2_8160 ( P1_SUB_88_U11 , P1_SUB_88_U220 , P1_SUB_88_U34 );
and AND2_8161 ( P1_SUB_88_U12 , P1_SUB_88_U219 , P1_SUB_88_U197 );
and AND2_8162 ( P1_SUB_88_U13 , P1_SUB_88_U217 , P1_SUB_88_U198 );
and AND2_8163 ( P1_SUB_88_U14 , P1_SUB_88_U216 , P1_SUB_88_U172 );
and AND2_8164 ( P1_SUB_88_U15 , P1_SUB_88_U215 , P1_SUB_88_U200 );
and AND2_8165 ( P1_SUB_88_U16 , P1_SUB_88_U213 , P1_SUB_88_U201 );
and AND2_8166 ( P1_SUB_88_U17 , P1_SUB_88_U212 , P1_SUB_88_U169 );
and AND2_8167 ( P1_SUB_88_U18 , P1_SUB_88_U211 , P1_SUB_88_U167 );
and AND2_8168 ( P1_SUB_88_U19 , P1_SUB_88_U209 , P1_SUB_88_U204 );
and AND2_8169 ( P1_SUB_88_U20 , P1_SUB_88_U208 , P1_SUB_88_U33 );
and AND2_8170 ( P1_SUB_88_U21 , P1_SUB_88_U207 , P1_SUB_88_U27 );
and AND2_8171 ( P1_SUB_88_U22 , P1_SUB_88_U190 , P1_SUB_88_U180 );
and AND2_8172 ( P1_SUB_88_U23 , P1_SUB_88_U189 , P1_SUB_88_U29 );
and AND2_8173 ( P1_SUB_88_U24 , P1_SUB_88_U188 , P1_SUB_88_U30 );
and AND2_8174 ( P1_SUB_88_U25 , P1_SUB_88_U186 , P1_SUB_88_U183 );
and AND2_8175 ( P1_SUB_88_U26 , P1_SUB_88_U185 , P1_SUB_88_U28 );
or OR3_8176 ( P1_SUB_88_U27 , P1_IR_REG_1_ , P1_IR_REG_0_ , P1_IR_REG_2_ );
nand NAND3_8177 ( P1_SUB_88_U28 , P1_SUB_88_U44 , P1_SUB_88_U230 , P1_SUB_88_U43 );
nand NAND2_8178 ( P1_SUB_88_U29 , P1_SUB_88_U45 , P1_SUB_88_U230 );
nand NAND2_8179 ( P1_SUB_88_U30 , P1_SUB_88_U46 , P1_SUB_88_U181 );
not NOT1_8180 ( P1_SUB_88_U31 , P1_IR_REG_7_ );
not NOT1_8181 ( P1_SUB_88_U32 , P1_IR_REG_3_ );
nand NAND2_8182 ( P1_SUB_88_U33 , P1_SUB_88_U56 , P1_SUB_88_U51 );
nand NAND4_8183 ( P1_SUB_88_U34 , P1_SUB_88_U130 , P1_SUB_88_U129 , P1_SUB_88_U128 , P1_SUB_88_U127 );
nand NAND2_8184 ( P1_SUB_88_U35 , P1_SUB_88_U156 , P1_SUB_88_U184 );
nand NAND2_8185 ( P1_SUB_88_U36 , P1_SUB_88_U157 , P1_SUB_88_U193 );
not NOT1_8186 ( P1_SUB_88_U37 , P1_IR_REG_15_ );
nand NAND2_8187 ( P1_SUB_88_U38 , P1_SUB_88_U158 , P1_SUB_88_U184 );
not NOT1_8188 ( P1_SUB_88_U39 , P1_IR_REG_11_ );
nand NAND2_8189 ( P1_SUB_88_U40 , P1_SUB_88_U247 , P1_SUB_88_U246 );
nand NAND2_8190 ( P1_SUB_88_U41 , P1_SUB_88_U237 , P1_SUB_88_U236 );
nand NAND2_8191 ( P1_SUB_88_U42 , P1_SUB_88_U241 , P1_SUB_88_U240 );
nor nor_8192 ( P1_SUB_88_U43 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8193 ( P1_SUB_88_U44 , P1_IR_REG_7_ , P1_IR_REG_8_ );
nor nor_8194 ( P1_SUB_88_U45 , P1_IR_REG_3_ , P1_IR_REG_4_ );
nor nor_8195 ( P1_SUB_88_U46 , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8196 ( P1_SUB_88_U47 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_8197 ( P1_SUB_88_U48 , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_8198 ( P1_SUB_88_U49 , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_8199 ( P1_SUB_88_U50 , P1_IR_REG_22_ , P1_IR_REG_20_ , P1_IR_REG_21_ );
and AND4_8200 ( P1_SUB_88_U51 , P1_SUB_88_U50 , P1_SUB_88_U49 , P1_SUB_88_U48 , P1_SUB_88_U47 );
nor nor_8201 ( P1_SUB_88_U52 , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ );
nor nor_8202 ( P1_SUB_88_U53 , P1_IR_REG_27_ , P1_IR_REG_28_ , P1_IR_REG_29_ , P1_IR_REG_2_ );
nor nor_8203 ( P1_SUB_88_U54 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8204 ( P1_SUB_88_U55 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_8205 ( P1_SUB_88_U56 , P1_SUB_88_U55 , P1_SUB_88_U54 , P1_SUB_88_U53 , P1_SUB_88_U52 );
nor nor_8206 ( P1_SUB_88_U57 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_8207 ( P1_SUB_88_U58 , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_8208 ( P1_SUB_88_U59 , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_8209 ( P1_SUB_88_U60 , P1_IR_REG_22_ , P1_IR_REG_20_ , P1_IR_REG_21_ );
and AND4_8210 ( P1_SUB_88_U61 , P1_SUB_88_U60 , P1_SUB_88_U59 , P1_SUB_88_U58 , P1_SUB_88_U57 );
nor nor_8211 ( P1_SUB_88_U62 , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ );
nor nor_8212 ( P1_SUB_88_U63 , P1_IR_REG_2_ , P1_IR_REG_27_ , P1_IR_REG_28_ );
nor nor_8213 ( P1_SUB_88_U64 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8214 ( P1_SUB_88_U65 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_8215 ( P1_SUB_88_U66 , P1_SUB_88_U65 , P1_SUB_88_U64 , P1_SUB_88_U63 , P1_SUB_88_U62 );
nor nor_8216 ( P1_SUB_88_U67 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_8217 ( P1_SUB_88_U68 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_8218 ( P1_SUB_88_U69 , P1_IR_REG_17_ , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
nor nor_8219 ( P1_SUB_88_U70 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
and AND4_8220 ( P1_SUB_88_U71 , P1_SUB_88_U70 , P1_SUB_88_U69 , P1_SUB_88_U68 , P1_SUB_88_U67 );
nor nor_8221 ( P1_SUB_88_U72 , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ );
nor nor_8222 ( P1_SUB_88_U73 , P1_IR_REG_2_ , P1_IR_REG_26_ , P1_IR_REG_27_ );
nor nor_8223 ( P1_SUB_88_U74 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8224 ( P1_SUB_88_U75 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_8225 ( P1_SUB_88_U76 , P1_SUB_88_U75 , P1_SUB_88_U74 , P1_SUB_88_U73 , P1_SUB_88_U72 );
nor nor_8226 ( P1_SUB_88_U77 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_8227 ( P1_SUB_88_U78 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_8228 ( P1_SUB_88_U79 , P1_IR_REG_17_ , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
nor nor_8229 ( P1_SUB_88_U80 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
and AND4_8230 ( P1_SUB_88_U81 , P1_SUB_88_U80 , P1_SUB_88_U79 , P1_SUB_88_U78 , P1_SUB_88_U77 );
nor nor_8231 ( P1_SUB_88_U82 , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ );
nor nor_8232 ( P1_SUB_88_U83 , P1_IR_REG_3_ , P1_IR_REG_26_ , P1_IR_REG_2_ );
nor nor_8233 ( P1_SUB_88_U84 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_8234 ( P1_SUB_88_U85 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_8235 ( P1_SUB_88_U86 , P1_SUB_88_U85 , P1_SUB_88_U84 , P1_SUB_88_U83 , P1_SUB_88_U82 );
nor nor_8236 ( P1_SUB_88_U87 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_8237 ( P1_SUB_88_U88 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_8238 ( P1_SUB_88_U89 , P1_IR_REG_17_ , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
nor nor_8239 ( P1_SUB_88_U90 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
and AND4_8240 ( P1_SUB_88_U91 , P1_SUB_88_U90 , P1_SUB_88_U89 , P1_SUB_88_U88 , P1_SUB_88_U87 );
nor nor_8241 ( P1_SUB_88_U92 , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ );
nor nor_8242 ( P1_SUB_88_U93 , P1_IR_REG_3_ , P1_IR_REG_26_ , P1_IR_REG_2_ );
nor nor_8243 ( P1_SUB_88_U94 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_8244 ( P1_SUB_88_U95 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_8245 ( P1_SUB_88_U96 , P1_SUB_88_U95 , P1_SUB_88_U94 , P1_SUB_88_U93 , P1_SUB_88_U92 );
nor nor_8246 ( P1_SUB_88_U97 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_8247 ( P1_SUB_88_U98 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_8248 ( P1_SUB_88_U99 , P1_IR_REG_19_ , P1_IR_REG_17_ , P1_IR_REG_18_ );
nor nor_8249 ( P1_SUB_88_U100 , P1_IR_REG_20_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
and AND4_8250 ( P1_SUB_88_U101 , P1_SUB_88_U100 , P1_SUB_88_U99 , P1_SUB_88_U98 , P1_SUB_88_U97 );
nor nor_8251 ( P1_SUB_88_U102 , P1_IR_REG_21_ , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ );
nor nor_8252 ( P1_SUB_88_U103 , P1_IR_REG_3_ , P1_IR_REG_25_ , P1_IR_REG_2_ );
nor nor_8253 ( P1_SUB_88_U104 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_8254 ( P1_SUB_88_U105 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_8255 ( P1_SUB_88_U106 , P1_SUB_88_U105 , P1_SUB_88_U104 , P1_SUB_88_U103 , P1_SUB_88_U102 );
nor nor_8256 ( P1_SUB_88_U107 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_8257 ( P1_SUB_88_U108 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_8258 ( P1_SUB_88_U109 , P1_IR_REG_19_ , P1_IR_REG_17_ , P1_IR_REG_18_ );
nor nor_8259 ( P1_SUB_88_U110 , P1_IR_REG_20_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
and AND4_8260 ( P1_SUB_88_U111 , P1_SUB_88_U110 , P1_SUB_88_U109 , P1_SUB_88_U108 , P1_SUB_88_U107 );
nor nor_8261 ( P1_SUB_88_U112 , P1_IR_REG_23_ , P1_IR_REG_21_ , P1_IR_REG_22_ );
nor nor_8262 ( P1_SUB_88_U113 , P1_IR_REG_3_ , P1_IR_REG_24_ , P1_IR_REG_2_ );
nor nor_8263 ( P1_SUB_88_U114 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_8264 ( P1_SUB_88_U115 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_8265 ( P1_SUB_88_U116 , P1_SUB_88_U115 , P1_SUB_88_U114 , P1_SUB_88_U113 , P1_SUB_88_U112 );
nor nor_8266 ( P1_SUB_88_U117 , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8267 ( P1_SUB_88_U118 , P1_IR_REG_15_ , P1_IR_REG_13_ , P1_IR_REG_14_ );
nor nor_8268 ( P1_SUB_88_U119 , P1_IR_REG_18_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_8269 ( P1_SUB_88_U120 , P1_IR_REG_0_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
and AND4_8270 ( P1_SUB_88_U121 , P1_SUB_88_U120 , P1_SUB_88_U119 , P1_SUB_88_U118 , P1_SUB_88_U117 );
nor nor_8271 ( P1_SUB_88_U122 , P1_IR_REG_22_ , P1_IR_REG_20_ , P1_IR_REG_21_ );
nor nor_8272 ( P1_SUB_88_U123 , P1_IR_REG_3_ , P1_IR_REG_23_ , P1_IR_REG_2_ );
nor nor_8273 ( P1_SUB_88_U124 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_8274 ( P1_SUB_88_U125 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_8275 ( P1_SUB_88_U126 , P1_SUB_88_U125 , P1_SUB_88_U124 , P1_SUB_88_U123 , P1_SUB_88_U122 );
nor nor_8276 ( P1_SUB_88_U127 , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8277 ( P1_SUB_88_U128 , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_8278 ( P1_SUB_88_U129 , P1_IR_REG_2_ , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_8279 ( P1_SUB_88_U130 , P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ );
nor nor_8280 ( P1_SUB_88_U131 , P1_IR_REG_17_ , P1_IR_REG_18_ );
nor nor_8281 ( P1_SUB_88_U132 , P1_IR_REG_19_ , P1_IR_REG_20_ );
nor nor_8282 ( P1_SUB_88_U133 , P1_IR_REG_21_ , P1_IR_REG_22_ );
and AND3_8283 ( P1_SUB_88_U134 , P1_SUB_88_U132 , P1_SUB_88_U131 , P1_SUB_88_U133 );
nor nor_8284 ( P1_SUB_88_U135 , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8285 ( P1_SUB_88_U136 , P1_IR_REG_15_ , P1_IR_REG_13_ , P1_IR_REG_14_ );
and AND2_8286 ( P1_SUB_88_U137 , P1_SUB_88_U136 , P1_SUB_88_U135 );
nor nor_8287 ( P1_SUB_88_U138 , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_18_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_8288 ( P1_SUB_88_U139 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
nor nor_8289 ( P1_SUB_88_U140 , P1_IR_REG_4_ , P1_IR_REG_2_ , P1_IR_REG_3_ );
and AND2_8290 ( P1_SUB_88_U141 , P1_SUB_88_U140 , P1_SUB_88_U139 );
nor nor_8291 ( P1_SUB_88_U142 , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8292 ( P1_SUB_88_U143 , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8293 ( P1_SUB_88_U144 , P1_IR_REG_15_ , P1_IR_REG_13_ , P1_IR_REG_14_ );
nor nor_8294 ( P1_SUB_88_U145 , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_18_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_8295 ( P1_SUB_88_U146 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_2_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
nor nor_8296 ( P1_SUB_88_U147 , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8297 ( P1_SUB_88_U148 , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8298 ( P1_SUB_88_U149 , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_17_ , P1_IR_REG_15_ , P1_IR_REG_16_ );
nor nor_8299 ( P1_SUB_88_U150 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_2_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_8300 ( P1_SUB_88_U151 , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8301 ( P1_SUB_88_U152 , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8302 ( P1_SUB_88_U153 , P1_IR_REG_18_ , P1_IR_REG_1_ , P1_IR_REG_17_ , P1_IR_REG_15_ , P1_IR_REG_16_ );
nor nor_8303 ( P1_SUB_88_U154 , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_3_ , P1_IR_REG_0_ , P1_IR_REG_2_ );
nor nor_8304 ( P1_SUB_88_U155 , P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ );
nor nor_8305 ( P1_SUB_88_U156 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_9_ );
nor nor_8306 ( P1_SUB_88_U157 , P1_IR_REG_13_ , P1_IR_REG_14_ );
nor nor_8307 ( P1_SUB_88_U158 , P1_IR_REG_10_ , P1_IR_REG_9_ );
not NOT1_8308 ( P1_SUB_88_U159 , P1_IR_REG_9_ );
and AND2_8309 ( P1_SUB_88_U160 , P1_SUB_88_U233 , P1_SUB_88_U232 );
not NOT1_8310 ( P1_SUB_88_U161 , P1_IR_REG_5_ );
and AND2_8311 ( P1_SUB_88_U162 , P1_SUB_88_U235 , P1_SUB_88_U234 );
not NOT1_8312 ( P1_SUB_88_U163 , P1_IR_REG_31_ );
not NOT1_8313 ( P1_SUB_88_U164 , P1_IR_REG_30_ );
and AND2_8314 ( P1_SUB_88_U165 , P1_SUB_88_U239 , P1_SUB_88_U238 );
not NOT1_8315 ( P1_SUB_88_U166 , P1_IR_REG_27_ );
nand NAND2_8316 ( P1_SUB_88_U167 , P1_SUB_88_U96 , P1_SUB_88_U91 );
not NOT1_8317 ( P1_SUB_88_U168 , P1_IR_REG_25_ );
nand NAND2_8318 ( P1_SUB_88_U169 , P1_SUB_88_U116 , P1_SUB_88_U111 );
and AND2_8319 ( P1_SUB_88_U170 , P1_SUB_88_U243 , P1_SUB_88_U242 );
not NOT1_8320 ( P1_SUB_88_U171 , P1_IR_REG_21_ );
nand NAND5_8321 ( P1_SUB_88_U172 , P1_SUB_88_U144 , P1_SUB_88_U143 , P1_SUB_88_U145 , P1_SUB_88_U147 , P1_SUB_88_U146 );
and AND2_8322 ( P1_SUB_88_U173 , P1_SUB_88_U245 , P1_SUB_88_U244 );
not NOT1_8323 ( P1_SUB_88_U174 , P1_IR_REG_1_ );
not NOT1_8324 ( P1_SUB_88_U175 , P1_IR_REG_0_ );
not NOT1_8325 ( P1_SUB_88_U176 , P1_IR_REG_17_ );
and AND2_8326 ( P1_SUB_88_U177 , P1_SUB_88_U249 , P1_SUB_88_U248 );
not NOT1_8327 ( P1_SUB_88_U178 , P1_IR_REG_13_ );
and AND2_8328 ( P1_SUB_88_U179 , P1_SUB_88_U251 , P1_SUB_88_U250 );
nand NAND2_8329 ( P1_SUB_88_U180 , P1_SUB_88_U230 , P1_SUB_88_U32 );
not NOT1_8330 ( P1_SUB_88_U181 , P1_SUB_88_U29 );
not NOT1_8331 ( P1_SUB_88_U182 , P1_SUB_88_U30 );
nand NAND2_8332 ( P1_SUB_88_U183 , P1_SUB_88_U182 , P1_SUB_88_U31 );
not NOT1_8333 ( P1_SUB_88_U184 , P1_SUB_88_U28 );
nand NAND2_8334 ( P1_SUB_88_U185 , P1_IR_REG_8_ , P1_SUB_88_U183 );
nand NAND2_8335 ( P1_SUB_88_U186 , P1_IR_REG_7_ , P1_SUB_88_U30 );
nand NAND2_8336 ( P1_SUB_88_U187 , P1_SUB_88_U181 , P1_SUB_88_U161 );
nand NAND2_8337 ( P1_SUB_88_U188 , P1_IR_REG_6_ , P1_SUB_88_U187 );
nand NAND2_8338 ( P1_SUB_88_U189 , P1_IR_REG_4_ , P1_SUB_88_U180 );
nand NAND2_8339 ( P1_SUB_88_U190 , P1_IR_REG_3_ , P1_SUB_88_U27 );
not NOT1_8340 ( P1_SUB_88_U191 , P1_SUB_88_U38 );
nand NAND2_8341 ( P1_SUB_88_U192 , P1_SUB_88_U191 , P1_SUB_88_U39 );
not NOT1_8342 ( P1_SUB_88_U193 , P1_SUB_88_U35 );
not NOT1_8343 ( P1_SUB_88_U194 , P1_SUB_88_U36 );
nand NAND2_8344 ( P1_SUB_88_U195 , P1_SUB_88_U194 , P1_SUB_88_U37 );
not NOT1_8345 ( P1_SUB_88_U196 , P1_SUB_88_U34 );
nand NAND4_8346 ( P1_SUB_88_U197 , P1_SUB_88_U155 , P1_SUB_88_U154 , P1_SUB_88_U153 , P1_SUB_88_U152 );
nand NAND4_8347 ( P1_SUB_88_U198 , P1_SUB_88_U151 , P1_SUB_88_U150 , P1_SUB_88_U149 , P1_SUB_88_U148 );
not NOT1_8348 ( P1_SUB_88_U199 , P1_SUB_88_U172 );
nand NAND2_8349 ( P1_SUB_88_U200 , P1_SUB_88_U134 , P1_SUB_88_U196 );
nand NAND2_8350 ( P1_SUB_88_U201 , P1_SUB_88_U126 , P1_SUB_88_U121 );
not NOT1_8351 ( P1_SUB_88_U202 , P1_SUB_88_U169 );
not NOT1_8352 ( P1_SUB_88_U203 , P1_SUB_88_U167 );
nand NAND2_8353 ( P1_SUB_88_U204 , P1_SUB_88_U66 , P1_SUB_88_U61 );
not NOT1_8354 ( P1_SUB_88_U205 , P1_SUB_88_U33 );
or OR2_8355 ( P1_SUB_88_U206 , P1_IR_REG_1_ , P1_IR_REG_0_ );
nand NAND2_8356 ( P1_SUB_88_U207 , P1_IR_REG_2_ , P1_SUB_88_U206 );
nand NAND2_8357 ( P1_SUB_88_U208 , P1_IR_REG_29_ , P1_SUB_88_U204 );
nand NAND2_8358 ( P1_SUB_88_U209 , P1_IR_REG_28_ , P1_SUB_88_U229 );
nand NAND2_8359 ( P1_SUB_88_U210 , P1_SUB_88_U106 , P1_SUB_88_U101 );
nand NAND2_8360 ( P1_SUB_88_U211 , P1_IR_REG_26_ , P1_SUB_88_U210 );
nand NAND2_8361 ( P1_SUB_88_U212 , P1_IR_REG_24_ , P1_SUB_88_U201 );
nand NAND2_8362 ( P1_SUB_88_U213 , P1_IR_REG_23_ , P1_SUB_88_U200 );
nand NAND4_8363 ( P1_SUB_88_U214 , P1_SUB_88_U142 , P1_SUB_88_U141 , P1_SUB_88_U138 , P1_SUB_88_U137 );
nand NAND2_8364 ( P1_SUB_88_U215 , P1_IR_REG_22_ , P1_SUB_88_U214 );
nand NAND2_8365 ( P1_SUB_88_U216 , P1_IR_REG_20_ , P1_SUB_88_U198 );
nand NAND2_8366 ( P1_SUB_88_U217 , P1_IR_REG_19_ , P1_SUB_88_U197 );
nand NAND2_8367 ( P1_SUB_88_U218 , P1_SUB_88_U196 , P1_SUB_88_U176 );
nand NAND2_8368 ( P1_SUB_88_U219 , P1_IR_REG_18_ , P1_SUB_88_U218 );
nand NAND2_8369 ( P1_SUB_88_U220 , P1_IR_REG_16_ , P1_SUB_88_U195 );
nand NAND2_8370 ( P1_SUB_88_U221 , P1_IR_REG_15_ , P1_SUB_88_U36 );
nand NAND2_8371 ( P1_SUB_88_U222 , P1_SUB_88_U193 , P1_SUB_88_U178 );
nand NAND2_8372 ( P1_SUB_88_U223 , P1_IR_REG_14_ , P1_SUB_88_U222 );
nand NAND2_8373 ( P1_SUB_88_U224 , P1_IR_REG_12_ , P1_SUB_88_U192 );
nand NAND2_8374 ( P1_SUB_88_U225 , P1_IR_REG_11_ , P1_SUB_88_U38 );
nand NAND2_8375 ( P1_SUB_88_U226 , P1_SUB_88_U184 , P1_SUB_88_U159 );
nand NAND2_8376 ( P1_SUB_88_U227 , P1_IR_REG_10_ , P1_SUB_88_U226 );
nand NAND2_8377 ( P1_SUB_88_U228 , P1_SUB_88_U205 , P1_SUB_88_U164 );
nand NAND2_8378 ( P1_SUB_88_U229 , P1_SUB_88_U76 , P1_SUB_88_U71 );
not NOT1_8379 ( P1_SUB_88_U230 , P1_SUB_88_U27 );
nand NAND2_8380 ( P1_SUB_88_U231 , P1_SUB_88_U86 , P1_SUB_88_U81 );
nand NAND2_8381 ( P1_SUB_88_U232 , P1_IR_REG_9_ , P1_SUB_88_U28 );
nand NAND2_8382 ( P1_SUB_88_U233 , P1_SUB_88_U184 , P1_SUB_88_U159 );
nand NAND2_8383 ( P1_SUB_88_U234 , P1_IR_REG_5_ , P1_SUB_88_U29 );
nand NAND2_8384 ( P1_SUB_88_U235 , P1_SUB_88_U181 , P1_SUB_88_U161 );
nand NAND2_8385 ( P1_SUB_88_U236 , P1_SUB_88_U228 , P1_SUB_88_U163 );
nand NAND3_8386 ( P1_SUB_88_U237 , P1_SUB_88_U205 , P1_SUB_88_U164 , P1_IR_REG_31_ );
nand NAND2_8387 ( P1_SUB_88_U238 , P1_IR_REG_30_ , P1_SUB_88_U33 );
nand NAND2_8388 ( P1_SUB_88_U239 , P1_SUB_88_U205 , P1_SUB_88_U164 );
nand NAND2_8389 ( P1_SUB_88_U240 , P1_SUB_88_U203 , P1_IR_REG_27_ );
nand NAND2_8390 ( P1_SUB_88_U241 , P1_SUB_88_U231 , P1_SUB_88_U166 );
nand NAND2_8391 ( P1_SUB_88_U242 , P1_IR_REG_25_ , P1_SUB_88_U169 );
nand NAND2_8392 ( P1_SUB_88_U243 , P1_SUB_88_U202 , P1_SUB_88_U168 );
nand NAND2_8393 ( P1_SUB_88_U244 , P1_IR_REG_21_ , P1_SUB_88_U172 );
nand NAND2_8394 ( P1_SUB_88_U245 , P1_SUB_88_U199 , P1_SUB_88_U171 );
nand NAND2_8395 ( P1_SUB_88_U246 , P1_IR_REG_1_ , P1_SUB_88_U175 );
nand NAND2_8396 ( P1_SUB_88_U247 , P1_IR_REG_0_ , P1_SUB_88_U174 );
nand NAND2_8397 ( P1_SUB_88_U248 , P1_IR_REG_17_ , P1_SUB_88_U34 );
nand NAND2_8398 ( P1_SUB_88_U249 , P1_SUB_88_U196 , P1_SUB_88_U176 );
nand NAND2_8399 ( P1_SUB_88_U250 , P1_IR_REG_13_ , P1_SUB_88_U35 );
nand NAND2_8400 ( P1_SUB_88_U251 , P1_SUB_88_U193 , P1_SUB_88_U178 );
not NOT1_8401 ( P1_R1309_U6 , P1_U3057 );
not NOT1_8402 ( P1_R1309_U7 , P1_U3054 );
and AND2_8403 ( P1_R1309_U8 , P1_R1309_U10 , P1_R1309_U9 );
nand NAND2_8404 ( P1_R1309_U9 , P1_U3054 , P1_R1309_U6 );
nand NAND2_8405 ( P1_R1309_U10 , P1_U3057 , P1_R1309_U7 );
and AND2_8406 ( P1_R1282_U6 , P1_R1282_U135 , P1_R1282_U35 );
and AND2_8407 ( P1_R1282_U7 , P1_R1282_U133 , P1_R1282_U36 );
and AND2_8408 ( P1_R1282_U8 , P1_R1282_U132 , P1_R1282_U37 );
and AND2_8409 ( P1_R1282_U9 , P1_R1282_U131 , P1_R1282_U38 );
and AND2_8410 ( P1_R1282_U10 , P1_R1282_U129 , P1_R1282_U39 );
and AND2_8411 ( P1_R1282_U11 , P1_R1282_U128 , P1_R1282_U40 );
and AND2_8412 ( P1_R1282_U12 , P1_R1282_U127 , P1_R1282_U41 );
and AND2_8413 ( P1_R1282_U13 , P1_R1282_U125 , P1_R1282_U42 );
and AND2_8414 ( P1_R1282_U14 , P1_R1282_U123 , P1_R1282_U43 );
and AND2_8415 ( P1_R1282_U15 , P1_R1282_U121 , P1_R1282_U44 );
and AND2_8416 ( P1_R1282_U16 , P1_R1282_U119 , P1_R1282_U45 );
and AND2_8417 ( P1_R1282_U17 , P1_R1282_U117 , P1_R1282_U46 );
and AND2_8418 ( P1_R1282_U18 , P1_R1282_U115 , P1_R1282_U25 );
and AND2_8419 ( P1_R1282_U19 , P1_R1282_U113 , P1_R1282_U67 );
and AND2_8420 ( P1_R1282_U20 , P1_R1282_U98 , P1_R1282_U26 );
and AND2_8421 ( P1_R1282_U21 , P1_R1282_U97 , P1_R1282_U27 );
and AND2_8422 ( P1_R1282_U22 , P1_R1282_U96 , P1_R1282_U28 );
and AND2_8423 ( P1_R1282_U23 , P1_R1282_U94 , P1_R1282_U29 );
and AND2_8424 ( P1_R1282_U24 , P1_R1282_U93 , P1_R1282_U30 );
or OR3_8425 ( P1_R1282_U25 , P1_U3456 , P1_U3451 , P1_U3459 );
nand NAND2_8426 ( P1_R1282_U26 , P1_R1282_U87 , P1_R1282_U34 );
nand NAND2_8427 ( P1_R1282_U27 , P1_R1282_U88 , P1_R1282_U33 );
nand NAND2_8428 ( P1_R1282_U28 , P1_R1282_U58 , P1_R1282_U89 );
nand NAND2_8429 ( P1_R1282_U29 , P1_R1282_U90 , P1_R1282_U32 );
nand NAND2_8430 ( P1_R1282_U30 , P1_R1282_U91 , P1_R1282_U31 );
not NOT1_8431 ( P1_R1282_U31 , P1_U3477 );
not NOT1_8432 ( P1_R1282_U32 , P1_U3474 );
not NOT1_8433 ( P1_R1282_U33 , P1_U3465 );
not NOT1_8434 ( P1_R1282_U34 , P1_U3462 );
nand NAND2_8435 ( P1_R1282_U35 , P1_R1282_U59 , P1_R1282_U92 );
nand NAND2_8436 ( P1_R1282_U36 , P1_R1282_U99 , P1_R1282_U56 );
nand NAND2_8437 ( P1_R1282_U37 , P1_R1282_U100 , P1_R1282_U55 );
nand NAND2_8438 ( P1_R1282_U38 , P1_R1282_U60 , P1_R1282_U101 );
nand NAND2_8439 ( P1_R1282_U39 , P1_R1282_U102 , P1_R1282_U54 );
nand NAND2_8440 ( P1_R1282_U40 , P1_R1282_U103 , P1_R1282_U53 );
nand NAND2_8441 ( P1_R1282_U41 , P1_R1282_U61 , P1_R1282_U104 );
nand NAND3_8442 ( P1_R1282_U42 , P1_R1282_U105 , P1_R1282_U81 , P1_R1282_U52 );
nand NAND3_8443 ( P1_R1282_U43 , P1_R1282_U106 , P1_R1282_U77 , P1_R1282_U51 );
nand NAND3_8444 ( P1_R1282_U44 , P1_R1282_U107 , P1_R1282_U75 , P1_R1282_U50 );
nand NAND3_8445 ( P1_R1282_U45 , P1_R1282_U108 , P1_R1282_U73 , P1_R1282_U49 );
nand NAND3_8446 ( P1_R1282_U46 , P1_R1282_U109 , P1_R1282_U71 , P1_R1282_U48 );
not NOT1_8447 ( P1_R1282_U47 , P1_U4017 );
not NOT1_8448 ( P1_R1282_U48 , P1_U4007 );
not NOT1_8449 ( P1_R1282_U49 , P1_U4009 );
not NOT1_8450 ( P1_R1282_U50 , P1_U4011 );
not NOT1_8451 ( P1_R1282_U51 , P1_U4013 );
not NOT1_8452 ( P1_R1282_U52 , P1_U4015 );
not NOT1_8453 ( P1_R1282_U53 , P1_U3501 );
not NOT1_8454 ( P1_R1282_U54 , P1_U3498 );
not NOT1_8455 ( P1_R1282_U55 , P1_U3489 );
not NOT1_8456 ( P1_R1282_U56 , P1_U3486 );
nand NAND2_8457 ( P1_R1282_U57 , P1_R1282_U153 , P1_R1282_U152 );
nor nor_8458 ( P1_R1282_U58 , P1_U3468 , P1_U3471 );
nor nor_8459 ( P1_R1282_U59 , P1_U3483 , P1_U3480 );
nor nor_8460 ( P1_R1282_U60 , P1_U3492 , P1_U3495 );
nor nor_8461 ( P1_R1282_U61 , P1_U3504 , P1_U3507 );
not NOT1_8462 ( P1_R1282_U62 , P1_U3480 );
and AND2_8463 ( P1_R1282_U63 , P1_R1282_U137 , P1_R1282_U136 );
not NOT1_8464 ( P1_R1282_U64 , P1_U3468 );
and AND2_8465 ( P1_R1282_U65 , P1_R1282_U139 , P1_R1282_U138 );
not NOT1_8466 ( P1_R1282_U66 , P1_U4016 );
nand NAND3_8467 ( P1_R1282_U67 , P1_R1282_U110 , P1_R1282_U69 , P1_R1282_U47 );
and AND2_8468 ( P1_R1282_U68 , P1_R1282_U141 , P1_R1282_U140 );
not NOT1_8469 ( P1_R1282_U69 , P1_U4018 );
and AND2_8470 ( P1_R1282_U70 , P1_R1282_U143 , P1_R1282_U142 );
not NOT1_8471 ( P1_R1282_U71 , P1_U4008 );
and AND2_8472 ( P1_R1282_U72 , P1_R1282_U145 , P1_R1282_U144 );
not NOT1_8473 ( P1_R1282_U73 , P1_U4010 );
and AND2_8474 ( P1_R1282_U74 , P1_R1282_U147 , P1_R1282_U146 );
not NOT1_8475 ( P1_R1282_U75 , P1_U4012 );
and AND2_8476 ( P1_R1282_U76 , P1_R1282_U149 , P1_R1282_U148 );
not NOT1_8477 ( P1_R1282_U77 , P1_U4014 );
and AND2_8478 ( P1_R1282_U78 , P1_R1282_U151 , P1_R1282_U150 );
not NOT1_8479 ( P1_R1282_U79 , P1_U3456 );
not NOT1_8480 ( P1_R1282_U80 , P1_U3451 );
not NOT1_8481 ( P1_R1282_U81 , P1_U3509 );
and AND2_8482 ( P1_R1282_U82 , P1_R1282_U155 , P1_R1282_U154 );
not NOT1_8483 ( P1_R1282_U83 , P1_U3504 );
and AND2_8484 ( P1_R1282_U84 , P1_R1282_U157 , P1_R1282_U156 );
not NOT1_8485 ( P1_R1282_U85 , P1_U3492 );
and AND2_8486 ( P1_R1282_U86 , P1_R1282_U159 , P1_R1282_U158 );
not NOT1_8487 ( P1_R1282_U87 , P1_R1282_U25 );
not NOT1_8488 ( P1_R1282_U88 , P1_R1282_U26 );
not NOT1_8489 ( P1_R1282_U89 , P1_R1282_U27 );
not NOT1_8490 ( P1_R1282_U90 , P1_R1282_U28 );
not NOT1_8491 ( P1_R1282_U91 , P1_R1282_U29 );
not NOT1_8492 ( P1_R1282_U92 , P1_R1282_U30 );
nand NAND2_8493 ( P1_R1282_U93 , P1_U3477 , P1_R1282_U29 );
nand NAND2_8494 ( P1_R1282_U94 , P1_U3474 , P1_R1282_U28 );
nand NAND2_8495 ( P1_R1282_U95 , P1_R1282_U89 , P1_R1282_U64 );
nand NAND2_8496 ( P1_R1282_U96 , P1_U3471 , P1_R1282_U95 );
nand NAND2_8497 ( P1_R1282_U97 , P1_U3465 , P1_R1282_U26 );
nand NAND2_8498 ( P1_R1282_U98 , P1_U3462 , P1_R1282_U25 );
not NOT1_8499 ( P1_R1282_U99 , P1_R1282_U35 );
not NOT1_8500 ( P1_R1282_U100 , P1_R1282_U36 );
not NOT1_8501 ( P1_R1282_U101 , P1_R1282_U37 );
not NOT1_8502 ( P1_R1282_U102 , P1_R1282_U38 );
not NOT1_8503 ( P1_R1282_U103 , P1_R1282_U39 );
not NOT1_8504 ( P1_R1282_U104 , P1_R1282_U40 );
not NOT1_8505 ( P1_R1282_U105 , P1_R1282_U41 );
not NOT1_8506 ( P1_R1282_U106 , P1_R1282_U42 );
not NOT1_8507 ( P1_R1282_U107 , P1_R1282_U43 );
not NOT1_8508 ( P1_R1282_U108 , P1_R1282_U44 );
not NOT1_8509 ( P1_R1282_U109 , P1_R1282_U45 );
not NOT1_8510 ( P1_R1282_U110 , P1_R1282_U46 );
not NOT1_8511 ( P1_R1282_U111 , P1_R1282_U67 );
nand NAND2_8512 ( P1_R1282_U112 , P1_R1282_U110 , P1_R1282_U69 );
nand NAND2_8513 ( P1_R1282_U113 , P1_U4017 , P1_R1282_U112 );
or OR2_8514 ( P1_R1282_U114 , P1_U3456 , P1_U3451 );
nand NAND2_8515 ( P1_R1282_U115 , P1_U3459 , P1_R1282_U114 );
nand NAND2_8516 ( P1_R1282_U116 , P1_R1282_U109 , P1_R1282_U71 );
nand NAND2_8517 ( P1_R1282_U117 , P1_U4007 , P1_R1282_U116 );
nand NAND2_8518 ( P1_R1282_U118 , P1_R1282_U108 , P1_R1282_U73 );
nand NAND2_8519 ( P1_R1282_U119 , P1_U4009 , P1_R1282_U118 );
nand NAND2_8520 ( P1_R1282_U120 , P1_R1282_U107 , P1_R1282_U75 );
nand NAND2_8521 ( P1_R1282_U121 , P1_U4011 , P1_R1282_U120 );
nand NAND2_8522 ( P1_R1282_U122 , P1_R1282_U106 , P1_R1282_U77 );
nand NAND2_8523 ( P1_R1282_U123 , P1_U4013 , P1_R1282_U122 );
nand NAND2_8524 ( P1_R1282_U124 , P1_R1282_U105 , P1_R1282_U81 );
nand NAND2_8525 ( P1_R1282_U125 , P1_U4015 , P1_R1282_U124 );
nand NAND2_8526 ( P1_R1282_U126 , P1_R1282_U104 , P1_R1282_U83 );
nand NAND2_8527 ( P1_R1282_U127 , P1_U3507 , P1_R1282_U126 );
nand NAND2_8528 ( P1_R1282_U128 , P1_U3501 , P1_R1282_U39 );
nand NAND2_8529 ( P1_R1282_U129 , P1_U3498 , P1_R1282_U38 );
nand NAND2_8530 ( P1_R1282_U130 , P1_R1282_U101 , P1_R1282_U85 );
nand NAND2_8531 ( P1_R1282_U131 , P1_U3495 , P1_R1282_U130 );
nand NAND2_8532 ( P1_R1282_U132 , P1_U3489 , P1_R1282_U36 );
nand NAND2_8533 ( P1_R1282_U133 , P1_U3486 , P1_R1282_U35 );
nand NAND2_8534 ( P1_R1282_U134 , P1_R1282_U92 , P1_R1282_U62 );
nand NAND2_8535 ( P1_R1282_U135 , P1_U3483 , P1_R1282_U134 );
nand NAND2_8536 ( P1_R1282_U136 , P1_U3480 , P1_R1282_U30 );
nand NAND2_8537 ( P1_R1282_U137 , P1_R1282_U92 , P1_R1282_U62 );
nand NAND2_8538 ( P1_R1282_U138 , P1_U3468 , P1_R1282_U27 );
nand NAND2_8539 ( P1_R1282_U139 , P1_R1282_U89 , P1_R1282_U64 );
nand NAND2_8540 ( P1_R1282_U140 , P1_U4016 , P1_R1282_U67 );
nand NAND2_8541 ( P1_R1282_U141 , P1_R1282_U111 , P1_R1282_U66 );
nand NAND2_8542 ( P1_R1282_U142 , P1_U4018 , P1_R1282_U46 );
nand NAND2_8543 ( P1_R1282_U143 , P1_R1282_U110 , P1_R1282_U69 );
nand NAND2_8544 ( P1_R1282_U144 , P1_U4008 , P1_R1282_U45 );
nand NAND2_8545 ( P1_R1282_U145 , P1_R1282_U109 , P1_R1282_U71 );
nand NAND2_8546 ( P1_R1282_U146 , P1_U4010 , P1_R1282_U44 );
nand NAND2_8547 ( P1_R1282_U147 , P1_R1282_U108 , P1_R1282_U73 );
nand NAND2_8548 ( P1_R1282_U148 , P1_U4012 , P1_R1282_U43 );
nand NAND2_8549 ( P1_R1282_U149 , P1_R1282_U107 , P1_R1282_U75 );
nand NAND2_8550 ( P1_R1282_U150 , P1_U4014 , P1_R1282_U42 );
nand NAND2_8551 ( P1_R1282_U151 , P1_R1282_U106 , P1_R1282_U77 );
nand NAND2_8552 ( P1_R1282_U152 , P1_U3456 , P1_R1282_U80 );
nand NAND2_8553 ( P1_R1282_U153 , P1_U3451 , P1_R1282_U79 );
nand NAND2_8554 ( P1_R1282_U154 , P1_U3509 , P1_R1282_U41 );
nand NAND2_8555 ( P1_R1282_U155 , P1_R1282_U105 , P1_R1282_U81 );
nand NAND2_8556 ( P1_R1282_U156 , P1_U3504 , P1_R1282_U40 );
nand NAND2_8557 ( P1_R1282_U157 , P1_R1282_U104 , P1_R1282_U83 );
nand NAND2_8558 ( P1_R1282_U158 , P1_U3492 , P1_R1282_U37 );
nand NAND2_8559 ( P1_R1282_U159 , P1_R1282_U101 , P1_R1282_U85 );
and AND2_8560 ( P1_R1240_U4 , P1_R1240_U176 , P1_R1240_U175 );
and AND2_8561 ( P1_R1240_U5 , P1_R1240_U177 , P1_R1240_U178 );
and AND2_8562 ( P1_R1240_U6 , P1_R1240_U194 , P1_R1240_U193 );
and AND2_8563 ( P1_R1240_U7 , P1_R1240_U234 , P1_R1240_U233 );
and AND2_8564 ( P1_R1240_U8 , P1_R1240_U243 , P1_R1240_U242 );
and AND2_8565 ( P1_R1240_U9 , P1_R1240_U261 , P1_R1240_U260 );
and AND2_8566 ( P1_R1240_U10 , P1_R1240_U269 , P1_R1240_U268 );
and AND2_8567 ( P1_R1240_U11 , P1_R1240_U348 , P1_R1240_U345 );
and AND2_8568 ( P1_R1240_U12 , P1_R1240_U341 , P1_R1240_U338 );
and AND2_8569 ( P1_R1240_U13 , P1_R1240_U332 , P1_R1240_U329 );
and AND2_8570 ( P1_R1240_U14 , P1_R1240_U323 , P1_R1240_U320 );
and AND2_8571 ( P1_R1240_U15 , P1_R1240_U317 , P1_R1240_U315 );
and AND2_8572 ( P1_R1240_U16 , P1_R1240_U310 , P1_R1240_U307 );
and AND2_8573 ( P1_R1240_U17 , P1_R1240_U232 , P1_R1240_U229 );
and AND2_8574 ( P1_R1240_U18 , P1_R1240_U224 , P1_R1240_U221 );
and AND2_8575 ( P1_R1240_U19 , P1_R1240_U210 , P1_R1240_U207 );
not NOT1_8576 ( P1_R1240_U20 , P1_U3471 );
not NOT1_8577 ( P1_R1240_U21 , P1_U3069 );
not NOT1_8578 ( P1_R1240_U22 , P1_U3068 );
nand NAND2_8579 ( P1_R1240_U23 , P1_U3069 , P1_U3471 );
not NOT1_8580 ( P1_R1240_U24 , P1_U3474 );
not NOT1_8581 ( P1_R1240_U25 , P1_U3465 );
not NOT1_8582 ( P1_R1240_U26 , P1_U3058 );
not NOT1_8583 ( P1_R1240_U27 , P1_U3065 );
not NOT1_8584 ( P1_R1240_U28 , P1_U3459 );
not NOT1_8585 ( P1_R1240_U29 , P1_U3066 );
not NOT1_8586 ( P1_R1240_U30 , P1_U3451 );
not NOT1_8587 ( P1_R1240_U31 , P1_U3075 );
nand NAND2_8588 ( P1_R1240_U32 , P1_U3075 , P1_U3451 );
not NOT1_8589 ( P1_R1240_U33 , P1_U3462 );
not NOT1_8590 ( P1_R1240_U34 , P1_U3062 );
nand NAND2_8591 ( P1_R1240_U35 , P1_U3058 , P1_U3465 );
not NOT1_8592 ( P1_R1240_U36 , P1_U3468 );
not NOT1_8593 ( P1_R1240_U37 , P1_U3477 );
not NOT1_8594 ( P1_R1240_U38 , P1_U3082 );
not NOT1_8595 ( P1_R1240_U39 , P1_U3081 );
not NOT1_8596 ( P1_R1240_U40 , P1_U3480 );
nand NAND2_8597 ( P1_R1240_U41 , P1_R1240_U62 , P1_R1240_U202 );
nand NAND2_8598 ( P1_R1240_U42 , P1_R1240_U118 , P1_R1240_U190 );
nand NAND2_8599 ( P1_R1240_U43 , P1_R1240_U179 , P1_R1240_U180 );
nand NAND2_8600 ( P1_R1240_U44 , P1_U3456 , P1_U3076 );
nand NAND2_8601 ( P1_R1240_U45 , P1_R1240_U122 , P1_R1240_U216 );
nand NAND2_8602 ( P1_R1240_U46 , P1_R1240_U213 , P1_R1240_U212 );
not NOT1_8603 ( P1_R1240_U47 , P1_U4008 );
not NOT1_8604 ( P1_R1240_U48 , P1_U3051 );
not NOT1_8605 ( P1_R1240_U49 , P1_U3055 );
not NOT1_8606 ( P1_R1240_U50 , P1_U4009 );
not NOT1_8607 ( P1_R1240_U51 , P1_U4010 );
not NOT1_8608 ( P1_R1240_U52 , P1_U3056 );
not NOT1_8609 ( P1_R1240_U53 , P1_U4011 );
not NOT1_8610 ( P1_R1240_U54 , P1_U3063 );
not NOT1_8611 ( P1_R1240_U55 , P1_U4014 );
not NOT1_8612 ( P1_R1240_U56 , P1_U3073 );
not NOT1_8613 ( P1_R1240_U57 , P1_U3501 );
not NOT1_8614 ( P1_R1240_U58 , P1_U3071 );
not NOT1_8615 ( P1_R1240_U59 , P1_U3067 );
nand NAND2_8616 ( P1_R1240_U60 , P1_U3071 , P1_U3501 );
not NOT1_8617 ( P1_R1240_U61 , P1_U3504 );
nand NAND2_8618 ( P1_R1240_U62 , P1_U3082 , P1_U3477 );
not NOT1_8619 ( P1_R1240_U63 , P1_U3483 );
not NOT1_8620 ( P1_R1240_U64 , P1_U3060 );
not NOT1_8621 ( P1_R1240_U65 , P1_U3489 );
not NOT1_8622 ( P1_R1240_U66 , P1_U3070 );
not NOT1_8623 ( P1_R1240_U67 , P1_U3486 );
not NOT1_8624 ( P1_R1240_U68 , P1_U3061 );
nand NAND2_8625 ( P1_R1240_U69 , P1_U3061 , P1_U3486 );
not NOT1_8626 ( P1_R1240_U70 , P1_U3492 );
not NOT1_8627 ( P1_R1240_U71 , P1_U3078 );
not NOT1_8628 ( P1_R1240_U72 , P1_U3495 );
not NOT1_8629 ( P1_R1240_U73 , P1_U3077 );
not NOT1_8630 ( P1_R1240_U74 , P1_U3498 );
not NOT1_8631 ( P1_R1240_U75 , P1_U3072 );
not NOT1_8632 ( P1_R1240_U76 , P1_U3507 );
not NOT1_8633 ( P1_R1240_U77 , P1_U3080 );
nand NAND2_8634 ( P1_R1240_U78 , P1_U3080 , P1_U3507 );
not NOT1_8635 ( P1_R1240_U79 , P1_U3509 );
not NOT1_8636 ( P1_R1240_U80 , P1_U3079 );
nand NAND2_8637 ( P1_R1240_U81 , P1_U3079 , P1_U3509 );
not NOT1_8638 ( P1_R1240_U82 , P1_U4015 );
not NOT1_8639 ( P1_R1240_U83 , P1_U4013 );
not NOT1_8640 ( P1_R1240_U84 , P1_U3059 );
not NOT1_8641 ( P1_R1240_U85 , P1_U4012 );
not NOT1_8642 ( P1_R1240_U86 , P1_U3064 );
nand NAND2_8643 ( P1_R1240_U87 , P1_U4009 , P1_U3055 );
not NOT1_8644 ( P1_R1240_U88 , P1_U3052 );
not NOT1_8645 ( P1_R1240_U89 , P1_U4007 );
nand NAND2_8646 ( P1_R1240_U90 , P1_R1240_U303 , P1_R1240_U173 );
not NOT1_8647 ( P1_R1240_U91 , P1_U3074 );
nand NAND2_8648 ( P1_R1240_U92 , P1_R1240_U78 , P1_R1240_U312 );
nand NAND2_8649 ( P1_R1240_U93 , P1_R1240_U258 , P1_R1240_U257 );
nand NAND2_8650 ( P1_R1240_U94 , P1_R1240_U69 , P1_R1240_U334 );
nand NAND2_8651 ( P1_R1240_U95 , P1_R1240_U454 , P1_R1240_U453 );
nand NAND2_8652 ( P1_R1240_U96 , P1_R1240_U501 , P1_R1240_U500 );
nand NAND2_8653 ( P1_R1240_U97 , P1_R1240_U372 , P1_R1240_U371 );
nand NAND2_8654 ( P1_R1240_U98 , P1_R1240_U377 , P1_R1240_U376 );
nand NAND2_8655 ( P1_R1240_U99 , P1_R1240_U384 , P1_R1240_U383 );
nand NAND2_8656 ( P1_R1240_U100 , P1_R1240_U391 , P1_R1240_U390 );
nand NAND2_8657 ( P1_R1240_U101 , P1_R1240_U396 , P1_R1240_U395 );
nand NAND2_8658 ( P1_R1240_U102 , P1_R1240_U405 , P1_R1240_U404 );
nand NAND2_8659 ( P1_R1240_U103 , P1_R1240_U412 , P1_R1240_U411 );
nand NAND2_8660 ( P1_R1240_U104 , P1_R1240_U419 , P1_R1240_U418 );
nand NAND2_8661 ( P1_R1240_U105 , P1_R1240_U426 , P1_R1240_U425 );
nand NAND2_8662 ( P1_R1240_U106 , P1_R1240_U431 , P1_R1240_U430 );
nand NAND2_8663 ( P1_R1240_U107 , P1_R1240_U438 , P1_R1240_U437 );
nand NAND2_8664 ( P1_R1240_U108 , P1_R1240_U445 , P1_R1240_U444 );
nand NAND2_8665 ( P1_R1240_U109 , P1_R1240_U459 , P1_R1240_U458 );
nand NAND2_8666 ( P1_R1240_U110 , P1_R1240_U464 , P1_R1240_U463 );
nand NAND2_8667 ( P1_R1240_U111 , P1_R1240_U471 , P1_R1240_U470 );
nand NAND2_8668 ( P1_R1240_U112 , P1_R1240_U478 , P1_R1240_U477 );
nand NAND2_8669 ( P1_R1240_U113 , P1_R1240_U485 , P1_R1240_U484 );
nand NAND2_8670 ( P1_R1240_U114 , P1_R1240_U492 , P1_R1240_U491 );
nand NAND2_8671 ( P1_R1240_U115 , P1_R1240_U497 , P1_R1240_U496 );
and AND2_8672 ( P1_R1240_U116 , P1_U3459 , P1_U3066 );
and AND2_8673 ( P1_R1240_U117 , P1_R1240_U186 , P1_R1240_U184 );
and AND2_8674 ( P1_R1240_U118 , P1_R1240_U191 , P1_R1240_U189 );
and AND2_8675 ( P1_R1240_U119 , P1_R1240_U198 , P1_R1240_U197 );
and AND3_8676 ( P1_R1240_U120 , P1_R1240_U379 , P1_R1240_U378 , P1_R1240_U23 );
and AND2_8677 ( P1_R1240_U121 , P1_R1240_U209 , P1_R1240_U6 );
and AND2_8678 ( P1_R1240_U122 , P1_R1240_U217 , P1_R1240_U215 );
and AND3_8679 ( P1_R1240_U123 , P1_R1240_U386 , P1_R1240_U385 , P1_R1240_U35 );
and AND2_8680 ( P1_R1240_U124 , P1_R1240_U223 , P1_R1240_U4 );
and AND2_8681 ( P1_R1240_U125 , P1_R1240_U231 , P1_R1240_U178 );
and AND2_8682 ( P1_R1240_U126 , P1_R1240_U201 , P1_R1240_U7 );
and AND2_8683 ( P1_R1240_U127 , P1_R1240_U236 , P1_R1240_U168 );
and AND2_8684 ( P1_R1240_U128 , P1_R1240_U245 , P1_R1240_U169 );
and AND2_8685 ( P1_R1240_U129 , P1_R1240_U265 , P1_R1240_U264 );
and AND2_8686 ( P1_R1240_U130 , P1_R1240_U10 , P1_R1240_U279 );
and AND2_8687 ( P1_R1240_U131 , P1_R1240_U282 , P1_R1240_U277 );
and AND2_8688 ( P1_R1240_U132 , P1_R1240_U298 , P1_R1240_U295 );
and AND2_8689 ( P1_R1240_U133 , P1_R1240_U365 , P1_R1240_U299 );
and AND2_8690 ( P1_R1240_U134 , P1_R1240_U156 , P1_R1240_U275 );
and AND3_8691 ( P1_R1240_U135 , P1_R1240_U466 , P1_R1240_U465 , P1_R1240_U60 );
and AND3_8692 ( P1_R1240_U136 , P1_R1240_U487 , P1_R1240_U486 , P1_R1240_U169 );
and AND2_8693 ( P1_R1240_U137 , P1_R1240_U340 , P1_R1240_U8 );
and AND3_8694 ( P1_R1240_U138 , P1_R1240_U499 , P1_R1240_U498 , P1_R1240_U168 );
and AND2_8695 ( P1_R1240_U139 , P1_R1240_U347 , P1_R1240_U7 );
nand NAND2_8696 ( P1_R1240_U140 , P1_R1240_U119 , P1_R1240_U199 );
nand NAND2_8697 ( P1_R1240_U141 , P1_R1240_U214 , P1_R1240_U226 );
not NOT1_8698 ( P1_R1240_U142 , P1_U3053 );
not NOT1_8699 ( P1_R1240_U143 , P1_U4018 );
and AND2_8700 ( P1_R1240_U144 , P1_R1240_U400 , P1_R1240_U399 );
nand NAND3_8701 ( P1_R1240_U145 , P1_R1240_U301 , P1_R1240_U166 , P1_R1240_U361 );
and AND2_8702 ( P1_R1240_U146 , P1_R1240_U407 , P1_R1240_U406 );
nand NAND3_8703 ( P1_R1240_U147 , P1_R1240_U367 , P1_R1240_U366 , P1_R1240_U133 );
and AND2_8704 ( P1_R1240_U148 , P1_R1240_U414 , P1_R1240_U413 );
nand NAND3_8705 ( P1_R1240_U149 , P1_R1240_U362 , P1_R1240_U296 , P1_R1240_U87 );
and AND2_8706 ( P1_R1240_U150 , P1_R1240_U421 , P1_R1240_U420 );
nand NAND2_8707 ( P1_R1240_U151 , P1_R1240_U290 , P1_R1240_U289 );
and AND2_8708 ( P1_R1240_U152 , P1_R1240_U433 , P1_R1240_U432 );
nand NAND2_8709 ( P1_R1240_U153 , P1_R1240_U286 , P1_R1240_U285 );
and AND2_8710 ( P1_R1240_U154 , P1_R1240_U440 , P1_R1240_U439 );
nand NAND2_8711 ( P1_R1240_U155 , P1_R1240_U131 , P1_R1240_U281 );
and AND2_8712 ( P1_R1240_U156 , P1_R1240_U447 , P1_R1240_U446 );
and AND2_8713 ( P1_R1240_U157 , P1_R1240_U452 , P1_R1240_U451 );
nand NAND2_8714 ( P1_R1240_U158 , P1_R1240_U44 , P1_R1240_U324 );
nand NAND2_8715 ( P1_R1240_U159 , P1_R1240_U129 , P1_R1240_U266 );
and AND2_8716 ( P1_R1240_U160 , P1_R1240_U473 , P1_R1240_U472 );
nand NAND2_8717 ( P1_R1240_U161 , P1_R1240_U254 , P1_R1240_U253 );
and AND2_8718 ( P1_R1240_U162 , P1_R1240_U480 , P1_R1240_U479 );
nand NAND2_8719 ( P1_R1240_U163 , P1_R1240_U250 , P1_R1240_U249 );
nand NAND2_8720 ( P1_R1240_U164 , P1_R1240_U240 , P1_R1240_U239 );
nand NAND2_8721 ( P1_R1240_U165 , P1_R1240_U364 , P1_R1240_U363 );
nand NAND2_8722 ( P1_R1240_U166 , P1_U3052 , P1_R1240_U147 );
not NOT1_8723 ( P1_R1240_U167 , P1_R1240_U35 );
nand NAND2_8724 ( P1_R1240_U168 , P1_U3480 , P1_U3081 );
nand NAND2_8725 ( P1_R1240_U169 , P1_U3070 , P1_U3489 );
nand NAND2_8726 ( P1_R1240_U170 , P1_U3056 , P1_U4010 );
not NOT1_8727 ( P1_R1240_U171 , P1_R1240_U69 );
not NOT1_8728 ( P1_R1240_U172 , P1_R1240_U78 );
nand NAND2_8729 ( P1_R1240_U173 , P1_U3063 , P1_U4011 );
not NOT1_8730 ( P1_R1240_U174 , P1_R1240_U62 );
or OR2_8731 ( P1_R1240_U175 , P1_U3065 , P1_U3468 );
or OR2_8732 ( P1_R1240_U176 , P1_U3058 , P1_U3465 );
or OR2_8733 ( P1_R1240_U177 , P1_U3462 , P1_U3062 );
or OR2_8734 ( P1_R1240_U178 , P1_U3459 , P1_U3066 );
not NOT1_8735 ( P1_R1240_U179 , P1_R1240_U32 );
or OR2_8736 ( P1_R1240_U180 , P1_U3456 , P1_U3076 );
not NOT1_8737 ( P1_R1240_U181 , P1_R1240_U43 );
not NOT1_8738 ( P1_R1240_U182 , P1_R1240_U44 );
nand NAND2_8739 ( P1_R1240_U183 , P1_R1240_U43 , P1_R1240_U44 );
nand NAND2_8740 ( P1_R1240_U184 , P1_R1240_U116 , P1_R1240_U177 );
nand NAND2_8741 ( P1_R1240_U185 , P1_R1240_U5 , P1_R1240_U183 );
nand NAND2_8742 ( P1_R1240_U186 , P1_U3062 , P1_U3462 );
nand NAND2_8743 ( P1_R1240_U187 , P1_R1240_U117 , P1_R1240_U185 );
nand NAND2_8744 ( P1_R1240_U188 , P1_R1240_U36 , P1_R1240_U35 );
nand NAND2_8745 ( P1_R1240_U189 , P1_U3065 , P1_R1240_U188 );
nand NAND2_8746 ( P1_R1240_U190 , P1_R1240_U4 , P1_R1240_U187 );
nand NAND2_8747 ( P1_R1240_U191 , P1_U3468 , P1_R1240_U167 );
not NOT1_8748 ( P1_R1240_U192 , P1_R1240_U42 );
or OR2_8749 ( P1_R1240_U193 , P1_U3068 , P1_U3474 );
or OR2_8750 ( P1_R1240_U194 , P1_U3069 , P1_U3471 );
not NOT1_8751 ( P1_R1240_U195 , P1_R1240_U23 );
nand NAND2_8752 ( P1_R1240_U196 , P1_R1240_U24 , P1_R1240_U23 );
nand NAND2_8753 ( P1_R1240_U197 , P1_U3068 , P1_R1240_U196 );
nand NAND2_8754 ( P1_R1240_U198 , P1_U3474 , P1_R1240_U195 );
nand NAND2_8755 ( P1_R1240_U199 , P1_R1240_U6 , P1_R1240_U42 );
not NOT1_8756 ( P1_R1240_U200 , P1_R1240_U140 );
or OR2_8757 ( P1_R1240_U201 , P1_U3477 , P1_U3082 );
nand NAND2_8758 ( P1_R1240_U202 , P1_R1240_U201 , P1_R1240_U140 );
not NOT1_8759 ( P1_R1240_U203 , P1_R1240_U41 );
or OR2_8760 ( P1_R1240_U204 , P1_U3081 , P1_U3480 );
or OR2_8761 ( P1_R1240_U205 , P1_U3471 , P1_U3069 );
nand NAND2_8762 ( P1_R1240_U206 , P1_R1240_U205 , P1_R1240_U42 );
nand NAND2_8763 ( P1_R1240_U207 , P1_R1240_U120 , P1_R1240_U206 );
nand NAND2_8764 ( P1_R1240_U208 , P1_R1240_U192 , P1_R1240_U23 );
nand NAND2_8765 ( P1_R1240_U209 , P1_U3474 , P1_U3068 );
nand NAND2_8766 ( P1_R1240_U210 , P1_R1240_U121 , P1_R1240_U208 );
or OR2_8767 ( P1_R1240_U211 , P1_U3069 , P1_U3471 );
nand NAND2_8768 ( P1_R1240_U212 , P1_R1240_U182 , P1_R1240_U178 );
nand NAND2_8769 ( P1_R1240_U213 , P1_U3066 , P1_U3459 );
not NOT1_8770 ( P1_R1240_U214 , P1_R1240_U46 );
nand NAND2_8771 ( P1_R1240_U215 , P1_R1240_U181 , P1_R1240_U5 );
nand NAND2_8772 ( P1_R1240_U216 , P1_R1240_U46 , P1_R1240_U177 );
nand NAND2_8773 ( P1_R1240_U217 , P1_U3062 , P1_U3462 );
not NOT1_8774 ( P1_R1240_U218 , P1_R1240_U45 );
or OR2_8775 ( P1_R1240_U219 , P1_U3465 , P1_U3058 );
nand NAND2_8776 ( P1_R1240_U220 , P1_R1240_U219 , P1_R1240_U45 );
nand NAND2_8777 ( P1_R1240_U221 , P1_R1240_U123 , P1_R1240_U220 );
nand NAND2_8778 ( P1_R1240_U222 , P1_R1240_U218 , P1_R1240_U35 );
nand NAND2_8779 ( P1_R1240_U223 , P1_U3468 , P1_U3065 );
nand NAND2_8780 ( P1_R1240_U224 , P1_R1240_U124 , P1_R1240_U222 );
or OR2_8781 ( P1_R1240_U225 , P1_U3058 , P1_U3465 );
nand NAND2_8782 ( P1_R1240_U226 , P1_R1240_U181 , P1_R1240_U178 );
not NOT1_8783 ( P1_R1240_U227 , P1_R1240_U141 );
nand NAND2_8784 ( P1_R1240_U228 , P1_U3062 , P1_U3462 );
nand NAND4_8785 ( P1_R1240_U229 , P1_R1240_U398 , P1_R1240_U397 , P1_R1240_U44 , P1_R1240_U43 );
nand NAND2_8786 ( P1_R1240_U230 , P1_R1240_U44 , P1_R1240_U43 );
nand NAND2_8787 ( P1_R1240_U231 , P1_U3066 , P1_U3459 );
nand NAND2_8788 ( P1_R1240_U232 , P1_R1240_U125 , P1_R1240_U230 );
or OR2_8789 ( P1_R1240_U233 , P1_U3081 , P1_U3480 );
or OR2_8790 ( P1_R1240_U234 , P1_U3060 , P1_U3483 );
nand NAND2_8791 ( P1_R1240_U235 , P1_R1240_U174 , P1_R1240_U7 );
nand NAND2_8792 ( P1_R1240_U236 , P1_U3060 , P1_U3483 );
nand NAND2_8793 ( P1_R1240_U237 , P1_R1240_U127 , P1_R1240_U235 );
or OR2_8794 ( P1_R1240_U238 , P1_U3483 , P1_U3060 );
nand NAND2_8795 ( P1_R1240_U239 , P1_R1240_U126 , P1_R1240_U140 );
nand NAND2_8796 ( P1_R1240_U240 , P1_R1240_U238 , P1_R1240_U237 );
not NOT1_8797 ( P1_R1240_U241 , P1_R1240_U164 );
or OR2_8798 ( P1_R1240_U242 , P1_U3078 , P1_U3492 );
or OR2_8799 ( P1_R1240_U243 , P1_U3070 , P1_U3489 );
nand NAND2_8800 ( P1_R1240_U244 , P1_R1240_U171 , P1_R1240_U8 );
nand NAND2_8801 ( P1_R1240_U245 , P1_U3078 , P1_U3492 );
nand NAND2_8802 ( P1_R1240_U246 , P1_R1240_U128 , P1_R1240_U244 );
or OR2_8803 ( P1_R1240_U247 , P1_U3486 , P1_U3061 );
or OR2_8804 ( P1_R1240_U248 , P1_U3492 , P1_U3078 );
nand NAND3_8805 ( P1_R1240_U249 , P1_R1240_U247 , P1_R1240_U164 , P1_R1240_U8 );
nand NAND2_8806 ( P1_R1240_U250 , P1_R1240_U248 , P1_R1240_U246 );
not NOT1_8807 ( P1_R1240_U251 , P1_R1240_U163 );
or OR2_8808 ( P1_R1240_U252 , P1_U3495 , P1_U3077 );
nand NAND2_8809 ( P1_R1240_U253 , P1_R1240_U252 , P1_R1240_U163 );
nand NAND2_8810 ( P1_R1240_U254 , P1_U3077 , P1_U3495 );
not NOT1_8811 ( P1_R1240_U255 , P1_R1240_U161 );
or OR2_8812 ( P1_R1240_U256 , P1_U3498 , P1_U3072 );
nand NAND2_8813 ( P1_R1240_U257 , P1_R1240_U256 , P1_R1240_U161 );
nand NAND2_8814 ( P1_R1240_U258 , P1_U3072 , P1_U3498 );
not NOT1_8815 ( P1_R1240_U259 , P1_R1240_U93 );
or OR2_8816 ( P1_R1240_U260 , P1_U3067 , P1_U3504 );
or OR2_8817 ( P1_R1240_U261 , P1_U3071 , P1_U3501 );
not NOT1_8818 ( P1_R1240_U262 , P1_R1240_U60 );
nand NAND2_8819 ( P1_R1240_U263 , P1_R1240_U61 , P1_R1240_U60 );
nand NAND2_8820 ( P1_R1240_U264 , P1_U3067 , P1_R1240_U263 );
nand NAND2_8821 ( P1_R1240_U265 , P1_U3504 , P1_R1240_U262 );
nand NAND2_8822 ( P1_R1240_U266 , P1_R1240_U9 , P1_R1240_U93 );
not NOT1_8823 ( P1_R1240_U267 , P1_R1240_U159 );
or OR2_8824 ( P1_R1240_U268 , P1_U3074 , P1_U4015 );
or OR2_8825 ( P1_R1240_U269 , P1_U3079 , P1_U3509 );
or OR2_8826 ( P1_R1240_U270 , P1_U3073 , P1_U4014 );
not NOT1_8827 ( P1_R1240_U271 , P1_R1240_U81 );
nand NAND2_8828 ( P1_R1240_U272 , P1_U4015 , P1_R1240_U271 );
nand NAND2_8829 ( P1_R1240_U273 , P1_R1240_U272 , P1_R1240_U91 );
nand NAND2_8830 ( P1_R1240_U274 , P1_R1240_U81 , P1_R1240_U82 );
nand NAND2_8831 ( P1_R1240_U275 , P1_R1240_U274 , P1_R1240_U273 );
nand NAND2_8832 ( P1_R1240_U276 , P1_R1240_U172 , P1_R1240_U10 );
nand NAND2_8833 ( P1_R1240_U277 , P1_U3073 , P1_U4014 );
nand NAND2_8834 ( P1_R1240_U278 , P1_R1240_U275 , P1_R1240_U276 );
or OR2_8835 ( P1_R1240_U279 , P1_U3507 , P1_U3080 );
or OR2_8836 ( P1_R1240_U280 , P1_U4014 , P1_U3073 );
nand NAND3_8837 ( P1_R1240_U281 , P1_R1240_U270 , P1_R1240_U159 , P1_R1240_U130 );
nand NAND2_8838 ( P1_R1240_U282 , P1_R1240_U280 , P1_R1240_U278 );
not NOT1_8839 ( P1_R1240_U283 , P1_R1240_U155 );
or OR2_8840 ( P1_R1240_U284 , P1_U4013 , P1_U3059 );
nand NAND2_8841 ( P1_R1240_U285 , P1_R1240_U284 , P1_R1240_U155 );
nand NAND2_8842 ( P1_R1240_U286 , P1_U3059 , P1_U4013 );
not NOT1_8843 ( P1_R1240_U287 , P1_R1240_U153 );
or OR2_8844 ( P1_R1240_U288 , P1_U4012 , P1_U3064 );
nand NAND2_8845 ( P1_R1240_U289 , P1_R1240_U288 , P1_R1240_U153 );
nand NAND2_8846 ( P1_R1240_U290 , P1_U3064 , P1_U4012 );
not NOT1_8847 ( P1_R1240_U291 , P1_R1240_U151 );
or OR2_8848 ( P1_R1240_U292 , P1_U3056 , P1_U4010 );
nand NAND2_8849 ( P1_R1240_U293 , P1_R1240_U173 , P1_R1240_U170 );
not NOT1_8850 ( P1_R1240_U294 , P1_R1240_U87 );
or OR2_8851 ( P1_R1240_U295 , P1_U4011 , P1_U3063 );
nand NAND3_8852 ( P1_R1240_U296 , P1_R1240_U151 , P1_R1240_U295 , P1_R1240_U165 );
not NOT1_8853 ( P1_R1240_U297 , P1_R1240_U149 );
or OR2_8854 ( P1_R1240_U298 , P1_U4008 , P1_U3051 );
nand NAND2_8855 ( P1_R1240_U299 , P1_U3051 , P1_U4008 );
not NOT1_8856 ( P1_R1240_U300 , P1_R1240_U147 );
nand NAND2_8857 ( P1_R1240_U301 , P1_U4007 , P1_R1240_U147 );
not NOT1_8858 ( P1_R1240_U302 , P1_R1240_U145 );
nand NAND2_8859 ( P1_R1240_U303 , P1_R1240_U295 , P1_R1240_U151 );
not NOT1_8860 ( P1_R1240_U304 , P1_R1240_U90 );
or OR2_8861 ( P1_R1240_U305 , P1_U4010 , P1_U3056 );
nand NAND2_8862 ( P1_R1240_U306 , P1_R1240_U305 , P1_R1240_U90 );
nand NAND3_8863 ( P1_R1240_U307 , P1_R1240_U306 , P1_R1240_U170 , P1_R1240_U150 );
nand NAND2_8864 ( P1_R1240_U308 , P1_R1240_U304 , P1_R1240_U170 );
nand NAND2_8865 ( P1_R1240_U309 , P1_U4009 , P1_U3055 );
nand NAND3_8866 ( P1_R1240_U310 , P1_R1240_U308 , P1_R1240_U309 , P1_R1240_U165 );
or OR2_8867 ( P1_R1240_U311 , P1_U3056 , P1_U4010 );
nand NAND2_8868 ( P1_R1240_U312 , P1_R1240_U279 , P1_R1240_U159 );
not NOT1_8869 ( P1_R1240_U313 , P1_R1240_U92 );
nand NAND2_8870 ( P1_R1240_U314 , P1_R1240_U10 , P1_R1240_U92 );
nand NAND2_8871 ( P1_R1240_U315 , P1_R1240_U134 , P1_R1240_U314 );
nand NAND2_8872 ( P1_R1240_U316 , P1_R1240_U314 , P1_R1240_U275 );
nand NAND2_8873 ( P1_R1240_U317 , P1_R1240_U450 , P1_R1240_U316 );
or OR2_8874 ( P1_R1240_U318 , P1_U3509 , P1_U3079 );
nand NAND2_8875 ( P1_R1240_U319 , P1_R1240_U318 , P1_R1240_U92 );
nand NAND3_8876 ( P1_R1240_U320 , P1_R1240_U319 , P1_R1240_U81 , P1_R1240_U157 );
nand NAND2_8877 ( P1_R1240_U321 , P1_R1240_U313 , P1_R1240_U81 );
nand NAND2_8878 ( P1_R1240_U322 , P1_U3074 , P1_U4015 );
nand NAND3_8879 ( P1_R1240_U323 , P1_R1240_U322 , P1_R1240_U321 , P1_R1240_U10 );
or OR2_8880 ( P1_R1240_U324 , P1_U3456 , P1_U3076 );
not NOT1_8881 ( P1_R1240_U325 , P1_R1240_U158 );
or OR2_8882 ( P1_R1240_U326 , P1_U3079 , P1_U3509 );
or OR2_8883 ( P1_R1240_U327 , P1_U3501 , P1_U3071 );
nand NAND2_8884 ( P1_R1240_U328 , P1_R1240_U327 , P1_R1240_U93 );
nand NAND2_8885 ( P1_R1240_U329 , P1_R1240_U135 , P1_R1240_U328 );
nand NAND2_8886 ( P1_R1240_U330 , P1_R1240_U259 , P1_R1240_U60 );
nand NAND2_8887 ( P1_R1240_U331 , P1_U3504 , P1_U3067 );
nand NAND3_8888 ( P1_R1240_U332 , P1_R1240_U331 , P1_R1240_U330 , P1_R1240_U9 );
or OR2_8889 ( P1_R1240_U333 , P1_U3071 , P1_U3501 );
nand NAND2_8890 ( P1_R1240_U334 , P1_R1240_U247 , P1_R1240_U164 );
not NOT1_8891 ( P1_R1240_U335 , P1_R1240_U94 );
or OR2_8892 ( P1_R1240_U336 , P1_U3489 , P1_U3070 );
nand NAND2_8893 ( P1_R1240_U337 , P1_R1240_U336 , P1_R1240_U94 );
nand NAND2_8894 ( P1_R1240_U338 , P1_R1240_U136 , P1_R1240_U337 );
nand NAND2_8895 ( P1_R1240_U339 , P1_R1240_U335 , P1_R1240_U169 );
nand NAND2_8896 ( P1_R1240_U340 , P1_U3078 , P1_U3492 );
nand NAND2_8897 ( P1_R1240_U341 , P1_R1240_U137 , P1_R1240_U339 );
or OR2_8898 ( P1_R1240_U342 , P1_U3070 , P1_U3489 );
or OR2_8899 ( P1_R1240_U343 , P1_U3480 , P1_U3081 );
nand NAND2_8900 ( P1_R1240_U344 , P1_R1240_U343 , P1_R1240_U41 );
nand NAND2_8901 ( P1_R1240_U345 , P1_R1240_U138 , P1_R1240_U344 );
nand NAND2_8902 ( P1_R1240_U346 , P1_R1240_U203 , P1_R1240_U168 );
nand NAND2_8903 ( P1_R1240_U347 , P1_U3060 , P1_U3483 );
nand NAND2_8904 ( P1_R1240_U348 , P1_R1240_U139 , P1_R1240_U346 );
nand NAND2_8905 ( P1_R1240_U349 , P1_R1240_U204 , P1_R1240_U168 );
nand NAND2_8906 ( P1_R1240_U350 , P1_R1240_U201 , P1_R1240_U62 );
nand NAND2_8907 ( P1_R1240_U351 , P1_R1240_U211 , P1_R1240_U23 );
nand NAND2_8908 ( P1_R1240_U352 , P1_R1240_U225 , P1_R1240_U35 );
nand NAND2_8909 ( P1_R1240_U353 , P1_R1240_U228 , P1_R1240_U177 );
nand NAND2_8910 ( P1_R1240_U354 , P1_R1240_U311 , P1_R1240_U170 );
nand NAND2_8911 ( P1_R1240_U355 , P1_R1240_U295 , P1_R1240_U173 );
nand NAND2_8912 ( P1_R1240_U356 , P1_R1240_U326 , P1_R1240_U81 );
nand NAND2_8913 ( P1_R1240_U357 , P1_R1240_U279 , P1_R1240_U78 );
nand NAND2_8914 ( P1_R1240_U358 , P1_R1240_U333 , P1_R1240_U60 );
nand NAND2_8915 ( P1_R1240_U359 , P1_R1240_U342 , P1_R1240_U169 );
nand NAND2_8916 ( P1_R1240_U360 , P1_R1240_U247 , P1_R1240_U69 );
nand NAND2_8917 ( P1_R1240_U361 , P1_U4007 , P1_U3052 );
nand NAND2_8918 ( P1_R1240_U362 , P1_R1240_U293 , P1_R1240_U165 );
nand NAND2_8919 ( P1_R1240_U363 , P1_U3055 , P1_R1240_U292 );
nand NAND2_8920 ( P1_R1240_U364 , P1_U4009 , P1_R1240_U292 );
nand NAND3_8921 ( P1_R1240_U365 , P1_R1240_U293 , P1_R1240_U165 , P1_R1240_U298 );
nand NAND3_8922 ( P1_R1240_U366 , P1_R1240_U151 , P1_R1240_U165 , P1_R1240_U132 );
nand NAND2_8923 ( P1_R1240_U367 , P1_R1240_U294 , P1_R1240_U298 );
nand NAND2_8924 ( P1_R1240_U368 , P1_U3081 , P1_R1240_U40 );
nand NAND2_8925 ( P1_R1240_U369 , P1_U3480 , P1_R1240_U39 );
nand NAND2_8926 ( P1_R1240_U370 , P1_R1240_U369 , P1_R1240_U368 );
nand NAND2_8927 ( P1_R1240_U371 , P1_R1240_U349 , P1_R1240_U41 );
nand NAND2_8928 ( P1_R1240_U372 , P1_R1240_U370 , P1_R1240_U203 );
nand NAND2_8929 ( P1_R1240_U373 , P1_U3082 , P1_R1240_U37 );
nand NAND2_8930 ( P1_R1240_U374 , P1_U3477 , P1_R1240_U38 );
nand NAND2_8931 ( P1_R1240_U375 , P1_R1240_U374 , P1_R1240_U373 );
nand NAND2_8932 ( P1_R1240_U376 , P1_R1240_U350 , P1_R1240_U140 );
nand NAND2_8933 ( P1_R1240_U377 , P1_R1240_U200 , P1_R1240_U375 );
nand NAND2_8934 ( P1_R1240_U378 , P1_U3068 , P1_R1240_U24 );
nand NAND2_8935 ( P1_R1240_U379 , P1_U3474 , P1_R1240_U22 );
nand NAND2_8936 ( P1_R1240_U380 , P1_U3069 , P1_R1240_U20 );
nand NAND2_8937 ( P1_R1240_U381 , P1_U3471 , P1_R1240_U21 );
nand NAND2_8938 ( P1_R1240_U382 , P1_R1240_U381 , P1_R1240_U380 );
nand NAND2_8939 ( P1_R1240_U383 , P1_R1240_U351 , P1_R1240_U42 );
nand NAND2_8940 ( P1_R1240_U384 , P1_R1240_U382 , P1_R1240_U192 );
nand NAND2_8941 ( P1_R1240_U385 , P1_U3065 , P1_R1240_U36 );
nand NAND2_8942 ( P1_R1240_U386 , P1_U3468 , P1_R1240_U27 );
nand NAND2_8943 ( P1_R1240_U387 , P1_U3058 , P1_R1240_U25 );
nand NAND2_8944 ( P1_R1240_U388 , P1_U3465 , P1_R1240_U26 );
nand NAND2_8945 ( P1_R1240_U389 , P1_R1240_U388 , P1_R1240_U387 );
nand NAND2_8946 ( P1_R1240_U390 , P1_R1240_U352 , P1_R1240_U45 );
nand NAND2_8947 ( P1_R1240_U391 , P1_R1240_U389 , P1_R1240_U218 );
nand NAND2_8948 ( P1_R1240_U392 , P1_U3062 , P1_R1240_U33 );
nand NAND2_8949 ( P1_R1240_U393 , P1_U3462 , P1_R1240_U34 );
nand NAND2_8950 ( P1_R1240_U394 , P1_R1240_U393 , P1_R1240_U392 );
nand NAND2_8951 ( P1_R1240_U395 , P1_R1240_U353 , P1_R1240_U141 );
nand NAND2_8952 ( P1_R1240_U396 , P1_R1240_U227 , P1_R1240_U394 );
nand NAND2_8953 ( P1_R1240_U397 , P1_U3066 , P1_R1240_U28 );
nand NAND2_8954 ( P1_R1240_U398 , P1_U3459 , P1_R1240_U29 );
nand NAND2_8955 ( P1_R1240_U399 , P1_U3053 , P1_R1240_U143 );
nand NAND2_8956 ( P1_R1240_U400 , P1_U4018 , P1_R1240_U142 );
nand NAND2_8957 ( P1_R1240_U401 , P1_U3053 , P1_R1240_U143 );
nand NAND2_8958 ( P1_R1240_U402 , P1_U4018 , P1_R1240_U142 );
nand NAND2_8959 ( P1_R1240_U403 , P1_R1240_U402 , P1_R1240_U401 );
nand NAND2_8960 ( P1_R1240_U404 , P1_R1240_U144 , P1_R1240_U145 );
nand NAND2_8961 ( P1_R1240_U405 , P1_R1240_U302 , P1_R1240_U403 );
nand NAND2_8962 ( P1_R1240_U406 , P1_U3052 , P1_R1240_U89 );
nand NAND2_8963 ( P1_R1240_U407 , P1_U4007 , P1_R1240_U88 );
nand NAND2_8964 ( P1_R1240_U408 , P1_U3052 , P1_R1240_U89 );
nand NAND2_8965 ( P1_R1240_U409 , P1_U4007 , P1_R1240_U88 );
nand NAND2_8966 ( P1_R1240_U410 , P1_R1240_U409 , P1_R1240_U408 );
nand NAND2_8967 ( P1_R1240_U411 , P1_R1240_U146 , P1_R1240_U147 );
nand NAND2_8968 ( P1_R1240_U412 , P1_R1240_U300 , P1_R1240_U410 );
nand NAND2_8969 ( P1_R1240_U413 , P1_U3051 , P1_R1240_U47 );
nand NAND2_8970 ( P1_R1240_U414 , P1_U4008 , P1_R1240_U48 );
nand NAND2_8971 ( P1_R1240_U415 , P1_U3051 , P1_R1240_U47 );
nand NAND2_8972 ( P1_R1240_U416 , P1_U4008 , P1_R1240_U48 );
nand NAND2_8973 ( P1_R1240_U417 , P1_R1240_U416 , P1_R1240_U415 );
nand NAND2_8974 ( P1_R1240_U418 , P1_R1240_U148 , P1_R1240_U149 );
nand NAND2_8975 ( P1_R1240_U419 , P1_R1240_U297 , P1_R1240_U417 );
nand NAND2_8976 ( P1_R1240_U420 , P1_U3055 , P1_R1240_U50 );
nand NAND2_8977 ( P1_R1240_U421 , P1_U4009 , P1_R1240_U49 );
nand NAND2_8978 ( P1_R1240_U422 , P1_U3056 , P1_R1240_U51 );
nand NAND2_8979 ( P1_R1240_U423 , P1_U4010 , P1_R1240_U52 );
nand NAND2_8980 ( P1_R1240_U424 , P1_R1240_U423 , P1_R1240_U422 );
nand NAND2_8981 ( P1_R1240_U425 , P1_R1240_U354 , P1_R1240_U90 );
nand NAND2_8982 ( P1_R1240_U426 , P1_R1240_U424 , P1_R1240_U304 );
nand NAND2_8983 ( P1_R1240_U427 , P1_U3063 , P1_R1240_U53 );
nand NAND2_8984 ( P1_R1240_U428 , P1_U4011 , P1_R1240_U54 );
nand NAND2_8985 ( P1_R1240_U429 , P1_R1240_U428 , P1_R1240_U427 );
nand NAND2_8986 ( P1_R1240_U430 , P1_R1240_U355 , P1_R1240_U151 );
nand NAND2_8987 ( P1_R1240_U431 , P1_R1240_U291 , P1_R1240_U429 );
nand NAND2_8988 ( P1_R1240_U432 , P1_U3064 , P1_R1240_U85 );
nand NAND2_8989 ( P1_R1240_U433 , P1_U4012 , P1_R1240_U86 );
nand NAND2_8990 ( P1_R1240_U434 , P1_U3064 , P1_R1240_U85 );
nand NAND2_8991 ( P1_R1240_U435 , P1_U4012 , P1_R1240_U86 );
nand NAND2_8992 ( P1_R1240_U436 , P1_R1240_U435 , P1_R1240_U434 );
nand NAND2_8993 ( P1_R1240_U437 , P1_R1240_U152 , P1_R1240_U153 );
nand NAND2_8994 ( P1_R1240_U438 , P1_R1240_U287 , P1_R1240_U436 );
nand NAND2_8995 ( P1_R1240_U439 , P1_U3059 , P1_R1240_U83 );
nand NAND2_8996 ( P1_R1240_U440 , P1_U4013 , P1_R1240_U84 );
nand NAND2_8997 ( P1_R1240_U441 , P1_U3059 , P1_R1240_U83 );
nand NAND2_8998 ( P1_R1240_U442 , P1_U4013 , P1_R1240_U84 );
nand NAND2_8999 ( P1_R1240_U443 , P1_R1240_U442 , P1_R1240_U441 );
nand NAND2_9000 ( P1_R1240_U444 , P1_R1240_U154 , P1_R1240_U155 );
nand NAND2_9001 ( P1_R1240_U445 , P1_R1240_U283 , P1_R1240_U443 );
nand NAND2_9002 ( P1_R1240_U446 , P1_U3073 , P1_R1240_U55 );
nand NAND2_9003 ( P1_R1240_U447 , P1_U4014 , P1_R1240_U56 );
nand NAND2_9004 ( P1_R1240_U448 , P1_U3073 , P1_R1240_U55 );
nand NAND2_9005 ( P1_R1240_U449 , P1_U4014 , P1_R1240_U56 );
nand NAND2_9006 ( P1_R1240_U450 , P1_R1240_U449 , P1_R1240_U448 );
nand NAND2_9007 ( P1_R1240_U451 , P1_U3074 , P1_R1240_U82 );
nand NAND2_9008 ( P1_R1240_U452 , P1_U4015 , P1_R1240_U91 );
nand NAND2_9009 ( P1_R1240_U453 , P1_R1240_U179 , P1_R1240_U158 );
nand NAND2_9010 ( P1_R1240_U454 , P1_R1240_U325 , P1_R1240_U32 );
nand NAND2_9011 ( P1_R1240_U455 , P1_U3079 , P1_R1240_U79 );
nand NAND2_9012 ( P1_R1240_U456 , P1_U3509 , P1_R1240_U80 );
nand NAND2_9013 ( P1_R1240_U457 , P1_R1240_U456 , P1_R1240_U455 );
nand NAND2_9014 ( P1_R1240_U458 , P1_R1240_U356 , P1_R1240_U92 );
nand NAND2_9015 ( P1_R1240_U459 , P1_R1240_U457 , P1_R1240_U313 );
nand NAND2_9016 ( P1_R1240_U460 , P1_U3080 , P1_R1240_U76 );
nand NAND2_9017 ( P1_R1240_U461 , P1_U3507 , P1_R1240_U77 );
nand NAND2_9018 ( P1_R1240_U462 , P1_R1240_U461 , P1_R1240_U460 );
nand NAND2_9019 ( P1_R1240_U463 , P1_R1240_U357 , P1_R1240_U159 );
nand NAND2_9020 ( P1_R1240_U464 , P1_R1240_U267 , P1_R1240_U462 );
nand NAND2_9021 ( P1_R1240_U465 , P1_U3067 , P1_R1240_U61 );
nand NAND2_9022 ( P1_R1240_U466 , P1_U3504 , P1_R1240_U59 );
nand NAND2_9023 ( P1_R1240_U467 , P1_U3071 , P1_R1240_U57 );
nand NAND2_9024 ( P1_R1240_U468 , P1_U3501 , P1_R1240_U58 );
nand NAND2_9025 ( P1_R1240_U469 , P1_R1240_U468 , P1_R1240_U467 );
nand NAND2_9026 ( P1_R1240_U470 , P1_R1240_U358 , P1_R1240_U93 );
nand NAND2_9027 ( P1_R1240_U471 , P1_R1240_U469 , P1_R1240_U259 );
nand NAND2_9028 ( P1_R1240_U472 , P1_U3072 , P1_R1240_U74 );
nand NAND2_9029 ( P1_R1240_U473 , P1_U3498 , P1_R1240_U75 );
nand NAND2_9030 ( P1_R1240_U474 , P1_U3072 , P1_R1240_U74 );
nand NAND2_9031 ( P1_R1240_U475 , P1_U3498 , P1_R1240_U75 );
nand NAND2_9032 ( P1_R1240_U476 , P1_R1240_U475 , P1_R1240_U474 );
nand NAND2_9033 ( P1_R1240_U477 , P1_R1240_U160 , P1_R1240_U161 );
nand NAND2_9034 ( P1_R1240_U478 , P1_R1240_U255 , P1_R1240_U476 );
nand NAND2_9035 ( P1_R1240_U479 , P1_U3077 , P1_R1240_U72 );
nand NAND2_9036 ( P1_R1240_U480 , P1_U3495 , P1_R1240_U73 );
nand NAND2_9037 ( P1_R1240_U481 , P1_U3077 , P1_R1240_U72 );
nand NAND2_9038 ( P1_R1240_U482 , P1_U3495 , P1_R1240_U73 );
nand NAND2_9039 ( P1_R1240_U483 , P1_R1240_U482 , P1_R1240_U481 );
nand NAND2_9040 ( P1_R1240_U484 , P1_R1240_U162 , P1_R1240_U163 );
nand NAND2_9041 ( P1_R1240_U485 , P1_R1240_U251 , P1_R1240_U483 );
nand NAND2_9042 ( P1_R1240_U486 , P1_U3078 , P1_R1240_U70 );
nand NAND2_9043 ( P1_R1240_U487 , P1_U3492 , P1_R1240_U71 );
nand NAND2_9044 ( P1_R1240_U488 , P1_U3070 , P1_R1240_U65 );
nand NAND2_9045 ( P1_R1240_U489 , P1_U3489 , P1_R1240_U66 );
nand NAND2_9046 ( P1_R1240_U490 , P1_R1240_U489 , P1_R1240_U488 );
nand NAND2_9047 ( P1_R1240_U491 , P1_R1240_U359 , P1_R1240_U94 );
nand NAND2_9048 ( P1_R1240_U492 , P1_R1240_U490 , P1_R1240_U335 );
nand NAND2_9049 ( P1_R1240_U493 , P1_U3061 , P1_R1240_U67 );
nand NAND2_9050 ( P1_R1240_U494 , P1_U3486 , P1_R1240_U68 );
nand NAND2_9051 ( P1_R1240_U495 , P1_R1240_U494 , P1_R1240_U493 );
nand NAND2_9052 ( P1_R1240_U496 , P1_R1240_U360 , P1_R1240_U164 );
nand NAND2_9053 ( P1_R1240_U497 , P1_R1240_U241 , P1_R1240_U495 );
nand NAND2_9054 ( P1_R1240_U498 , P1_U3060 , P1_R1240_U63 );
nand NAND2_9055 ( P1_R1240_U499 , P1_U3483 , P1_R1240_U64 );
nand NAND2_9056 ( P1_R1240_U500 , P1_U3075 , P1_R1240_U30 );
nand NAND2_9057 ( P1_R1240_U501 , P1_U3451 , P1_R1240_U31 );
and AND2_9058 ( P1_R1162_U4 , P1_R1162_U95 , P1_R1162_U94 );
and AND2_9059 ( P1_R1162_U5 , P1_R1162_U96 , P1_R1162_U97 );
and AND2_9060 ( P1_R1162_U6 , P1_R1162_U113 , P1_R1162_U112 );
and AND2_9061 ( P1_R1162_U7 , P1_R1162_U155 , P1_R1162_U154 );
and AND2_9062 ( P1_R1162_U8 , P1_R1162_U164 , P1_R1162_U163 );
and AND2_9063 ( P1_R1162_U9 , P1_R1162_U182 , P1_R1162_U181 );
and AND2_9064 ( P1_R1162_U10 , P1_R1162_U218 , P1_R1162_U215 );
and AND2_9065 ( P1_R1162_U11 , P1_R1162_U211 , P1_R1162_U208 );
and AND2_9066 ( P1_R1162_U12 , P1_R1162_U202 , P1_R1162_U199 );
and AND2_9067 ( P1_R1162_U13 , P1_R1162_U196 , P1_R1162_U192 );
and AND2_9068 ( P1_R1162_U14 , P1_R1162_U151 , P1_R1162_U148 );
and AND2_9069 ( P1_R1162_U15 , P1_R1162_U143 , P1_R1162_U140 );
and AND2_9070 ( P1_R1162_U16 , P1_R1162_U129 , P1_R1162_U126 );
not NOT1_9071 ( P1_R1162_U17 , P1_REG1_REG_6_ );
not NOT1_9072 ( P1_R1162_U18 , P1_U3470 );
not NOT1_9073 ( P1_R1162_U19 , P1_U3473 );
nand NAND2_9074 ( P1_R1162_U20 , P1_U3470 , P1_REG1_REG_6_ );
not NOT1_9075 ( P1_R1162_U21 , P1_REG1_REG_7_ );
not NOT1_9076 ( P1_R1162_U22 , P1_REG1_REG_4_ );
not NOT1_9077 ( P1_R1162_U23 , P1_U3464 );
not NOT1_9078 ( P1_R1162_U24 , P1_U3467 );
not NOT1_9079 ( P1_R1162_U25 , P1_REG1_REG_2_ );
not NOT1_9080 ( P1_R1162_U26 , P1_U3458 );
not NOT1_9081 ( P1_R1162_U27 , P1_REG1_REG_0_ );
not NOT1_9082 ( P1_R1162_U28 , P1_U3449 );
nand NAND2_9083 ( P1_R1162_U29 , P1_U3449 , P1_REG1_REG_0_ );
not NOT1_9084 ( P1_R1162_U30 , P1_REG1_REG_3_ );
not NOT1_9085 ( P1_R1162_U31 , P1_U3461 );
nand NAND2_9086 ( P1_R1162_U32 , P1_U3464 , P1_REG1_REG_4_ );
not NOT1_9087 ( P1_R1162_U33 , P1_REG1_REG_5_ );
not NOT1_9088 ( P1_R1162_U34 , P1_REG1_REG_8_ );
not NOT1_9089 ( P1_R1162_U35 , P1_U3476 );
not NOT1_9090 ( P1_R1162_U36 , P1_U3479 );
not NOT1_9091 ( P1_R1162_U37 , P1_REG1_REG_9_ );
nand NAND2_9092 ( P1_R1162_U38 , P1_R1162_U49 , P1_R1162_U121 );
nand NAND3_9093 ( P1_R1162_U39 , P1_R1162_U110 , P1_R1162_U108 , P1_R1162_U109 );
nand NAND2_9094 ( P1_R1162_U40 , P1_R1162_U98 , P1_R1162_U99 );
nand NAND2_9095 ( P1_R1162_U41 , P1_REG1_REG_1_ , P1_U3455 );
nand NAND3_9096 ( P1_R1162_U42 , P1_R1162_U136 , P1_R1162_U134 , P1_R1162_U135 );
nand NAND2_9097 ( P1_R1162_U43 , P1_R1162_U132 , P1_R1162_U131 );
not NOT1_9098 ( P1_R1162_U44 , P1_REG1_REG_16_ );
not NOT1_9099 ( P1_R1162_U45 , P1_U3500 );
not NOT1_9100 ( P1_R1162_U46 , P1_U3503 );
nand NAND2_9101 ( P1_R1162_U47 , P1_U3500 , P1_REG1_REG_16_ );
not NOT1_9102 ( P1_R1162_U48 , P1_REG1_REG_17_ );
nand NAND2_9103 ( P1_R1162_U49 , P1_U3476 , P1_REG1_REG_8_ );
not NOT1_9104 ( P1_R1162_U50 , P1_REG1_REG_10_ );
not NOT1_9105 ( P1_R1162_U51 , P1_U3482 );
not NOT1_9106 ( P1_R1162_U52 , P1_REG1_REG_12_ );
not NOT1_9107 ( P1_R1162_U53 , P1_U3488 );
not NOT1_9108 ( P1_R1162_U54 , P1_REG1_REG_11_ );
not NOT1_9109 ( P1_R1162_U55 , P1_U3485 );
nand NAND2_9110 ( P1_R1162_U56 , P1_U3485 , P1_REG1_REG_11_ );
not NOT1_9111 ( P1_R1162_U57 , P1_REG1_REG_13_ );
not NOT1_9112 ( P1_R1162_U58 , P1_U3491 );
not NOT1_9113 ( P1_R1162_U59 , P1_REG1_REG_14_ );
not NOT1_9114 ( P1_R1162_U60 , P1_U3494 );
not NOT1_9115 ( P1_R1162_U61 , P1_REG1_REG_15_ );
not NOT1_9116 ( P1_R1162_U62 , P1_U3497 );
not NOT1_9117 ( P1_R1162_U63 , P1_REG1_REG_18_ );
not NOT1_9118 ( P1_R1162_U64 , P1_U3506 );
nand NAND3_9119 ( P1_R1162_U65 , P1_R1162_U186 , P1_R1162_U185 , P1_R1162_U187 );
nand NAND2_9120 ( P1_R1162_U66 , P1_R1162_U179 , P1_R1162_U178 );
nand NAND2_9121 ( P1_R1162_U67 , P1_R1162_U56 , P1_R1162_U204 );
nand NAND2_9122 ( P1_R1162_U68 , P1_R1162_U259 , P1_R1162_U258 );
nand NAND2_9123 ( P1_R1162_U69 , P1_R1162_U308 , P1_R1162_U307 );
nand NAND2_9124 ( P1_R1162_U70 , P1_R1162_U231 , P1_R1162_U230 );
nand NAND2_9125 ( P1_R1162_U71 , P1_R1162_U236 , P1_R1162_U235 );
nand NAND2_9126 ( P1_R1162_U72 , P1_R1162_U243 , P1_R1162_U242 );
nand NAND2_9127 ( P1_R1162_U73 , P1_R1162_U250 , P1_R1162_U249 );
nand NAND2_9128 ( P1_R1162_U74 , P1_R1162_U255 , P1_R1162_U254 );
nand NAND2_9129 ( P1_R1162_U75 , P1_R1162_U271 , P1_R1162_U270 );
nand NAND2_9130 ( P1_R1162_U76 , P1_R1162_U278 , P1_R1162_U277 );
nand NAND2_9131 ( P1_R1162_U77 , P1_R1162_U285 , P1_R1162_U284 );
nand NAND2_9132 ( P1_R1162_U78 , P1_R1162_U292 , P1_R1162_U291 );
nand NAND2_9133 ( P1_R1162_U79 , P1_R1162_U299 , P1_R1162_U298 );
nand NAND2_9134 ( P1_R1162_U80 , P1_R1162_U304 , P1_R1162_U303 );
nand NAND3_9135 ( P1_R1162_U81 , P1_R1162_U117 , P1_R1162_U116 , P1_R1162_U118 );
nand NAND2_9136 ( P1_R1162_U82 , P1_R1162_U133 , P1_R1162_U145 );
nand NAND2_9137 ( P1_R1162_U83 , P1_R1162_U41 , P1_R1162_U152 );
not NOT1_9138 ( P1_R1162_U84 , P1_U3443 );
not NOT1_9139 ( P1_R1162_U85 , P1_REG1_REG_19_ );
nand NAND2_9140 ( P1_R1162_U86 , P1_R1162_U175 , P1_R1162_U174 );
nand NAND2_9141 ( P1_R1162_U87 , P1_R1162_U171 , P1_R1162_U170 );
nand NAND2_9142 ( P1_R1162_U88 , P1_R1162_U161 , P1_R1162_U160 );
not NOT1_9143 ( P1_R1162_U89 , P1_R1162_U32 );
nand NAND2_9144 ( P1_R1162_U90 , P1_REG1_REG_9_ , P1_U3479 );
nand NAND2_9145 ( P1_R1162_U91 , P1_U3488 , P1_REG1_REG_12_ );
not NOT1_9146 ( P1_R1162_U92 , P1_R1162_U56 );
not NOT1_9147 ( P1_R1162_U93 , P1_R1162_U49 );
or OR2_9148 ( P1_R1162_U94 , P1_U3467 , P1_REG1_REG_5_ );
or OR2_9149 ( P1_R1162_U95 , P1_U3464 , P1_REG1_REG_4_ );
or OR2_9150 ( P1_R1162_U96 , P1_REG1_REG_3_ , P1_U3461 );
or OR2_9151 ( P1_R1162_U97 , P1_REG1_REG_2_ , P1_U3458 );
not NOT1_9152 ( P1_R1162_U98 , P1_R1162_U29 );
or OR2_9153 ( P1_R1162_U99 , P1_REG1_REG_1_ , P1_U3455 );
not NOT1_9154 ( P1_R1162_U100 , P1_R1162_U40 );
not NOT1_9155 ( P1_R1162_U101 , P1_R1162_U41 );
nand NAND2_9156 ( P1_R1162_U102 , P1_R1162_U40 , P1_R1162_U41 );
nand NAND3_9157 ( P1_R1162_U103 , P1_REG1_REG_2_ , P1_U3458 , P1_R1162_U96 );
nand NAND2_9158 ( P1_R1162_U104 , P1_R1162_U5 , P1_R1162_U102 );
nand NAND2_9159 ( P1_R1162_U105 , P1_U3461 , P1_REG1_REG_3_ );
nand NAND3_9160 ( P1_R1162_U106 , P1_R1162_U105 , P1_R1162_U103 , P1_R1162_U104 );
nand NAND2_9161 ( P1_R1162_U107 , P1_R1162_U33 , P1_R1162_U32 );
nand NAND2_9162 ( P1_R1162_U108 , P1_U3467 , P1_R1162_U107 );
nand NAND2_9163 ( P1_R1162_U109 , P1_R1162_U4 , P1_R1162_U106 );
nand NAND2_9164 ( P1_R1162_U110 , P1_REG1_REG_5_ , P1_R1162_U89 );
not NOT1_9165 ( P1_R1162_U111 , P1_R1162_U39 );
or OR2_9166 ( P1_R1162_U112 , P1_U3473 , P1_REG1_REG_7_ );
or OR2_9167 ( P1_R1162_U113 , P1_U3470 , P1_REG1_REG_6_ );
not NOT1_9168 ( P1_R1162_U114 , P1_R1162_U20 );
nand NAND2_9169 ( P1_R1162_U115 , P1_R1162_U21 , P1_R1162_U20 );
nand NAND2_9170 ( P1_R1162_U116 , P1_U3473 , P1_R1162_U115 );
nand NAND2_9171 ( P1_R1162_U117 , P1_REG1_REG_7_ , P1_R1162_U114 );
nand NAND2_9172 ( P1_R1162_U118 , P1_R1162_U6 , P1_R1162_U39 );
not NOT1_9173 ( P1_R1162_U119 , P1_R1162_U81 );
or OR2_9174 ( P1_R1162_U120 , P1_REG1_REG_8_ , P1_U3476 );
nand NAND2_9175 ( P1_R1162_U121 , P1_R1162_U120 , P1_R1162_U81 );
not NOT1_9176 ( P1_R1162_U122 , P1_R1162_U38 );
or OR2_9177 ( P1_R1162_U123 , P1_U3479 , P1_REG1_REG_9_ );
or OR2_9178 ( P1_R1162_U124 , P1_REG1_REG_6_ , P1_U3470 );
nand NAND2_9179 ( P1_R1162_U125 , P1_R1162_U124 , P1_R1162_U39 );
nand NAND4_9180 ( P1_R1162_U126 , P1_R1162_U238 , P1_R1162_U237 , P1_R1162_U20 , P1_R1162_U125 );
nand NAND2_9181 ( P1_R1162_U127 , P1_R1162_U111 , P1_R1162_U20 );
nand NAND2_9182 ( P1_R1162_U128 , P1_REG1_REG_7_ , P1_U3473 );
nand NAND3_9183 ( P1_R1162_U129 , P1_R1162_U128 , P1_R1162_U6 , P1_R1162_U127 );
or OR2_9184 ( P1_R1162_U130 , P1_U3470 , P1_REG1_REG_6_ );
nand NAND2_9185 ( P1_R1162_U131 , P1_R1162_U101 , P1_R1162_U97 );
nand NAND2_9186 ( P1_R1162_U132 , P1_U3458 , P1_REG1_REG_2_ );
not NOT1_9187 ( P1_R1162_U133 , P1_R1162_U43 );
nand NAND2_9188 ( P1_R1162_U134 , P1_R1162_U100 , P1_R1162_U5 );
nand NAND2_9189 ( P1_R1162_U135 , P1_R1162_U43 , P1_R1162_U96 );
nand NAND2_9190 ( P1_R1162_U136 , P1_U3461 , P1_REG1_REG_3_ );
not NOT1_9191 ( P1_R1162_U137 , P1_R1162_U42 );
or OR2_9192 ( P1_R1162_U138 , P1_REG1_REG_4_ , P1_U3464 );
nand NAND2_9193 ( P1_R1162_U139 , P1_R1162_U138 , P1_R1162_U42 );
nand NAND4_9194 ( P1_R1162_U140 , P1_R1162_U245 , P1_R1162_U244 , P1_R1162_U32 , P1_R1162_U139 );
nand NAND2_9195 ( P1_R1162_U141 , P1_R1162_U137 , P1_R1162_U32 );
nand NAND2_9196 ( P1_R1162_U142 , P1_REG1_REG_5_ , P1_U3467 );
nand NAND3_9197 ( P1_R1162_U143 , P1_R1162_U142 , P1_R1162_U4 , P1_R1162_U141 );
or OR2_9198 ( P1_R1162_U144 , P1_U3464 , P1_REG1_REG_4_ );
nand NAND2_9199 ( P1_R1162_U145 , P1_R1162_U100 , P1_R1162_U97 );
not NOT1_9200 ( P1_R1162_U146 , P1_R1162_U82 );
nand NAND2_9201 ( P1_R1162_U147 , P1_U3461 , P1_REG1_REG_3_ );
nand NAND4_9202 ( P1_R1162_U148 , P1_R1162_U257 , P1_R1162_U256 , P1_R1162_U41 , P1_R1162_U40 );
nand NAND2_9203 ( P1_R1162_U149 , P1_R1162_U41 , P1_R1162_U40 );
nand NAND2_9204 ( P1_R1162_U150 , P1_U3458 , P1_REG1_REG_2_ );
nand NAND3_9205 ( P1_R1162_U151 , P1_R1162_U150 , P1_R1162_U97 , P1_R1162_U149 );
or OR2_9206 ( P1_R1162_U152 , P1_REG1_REG_1_ , P1_U3455 );
not NOT1_9207 ( P1_R1162_U153 , P1_R1162_U83 );
or OR2_9208 ( P1_R1162_U154 , P1_U3479 , P1_REG1_REG_9_ );
or OR2_9209 ( P1_R1162_U155 , P1_U3482 , P1_REG1_REG_10_ );
nand NAND2_9210 ( P1_R1162_U156 , P1_R1162_U93 , P1_R1162_U7 );
nand NAND2_9211 ( P1_R1162_U157 , P1_U3482 , P1_REG1_REG_10_ );
nand NAND3_9212 ( P1_R1162_U158 , P1_R1162_U157 , P1_R1162_U90 , P1_R1162_U156 );
or OR2_9213 ( P1_R1162_U159 , P1_REG1_REG_10_ , P1_U3482 );
nand NAND3_9214 ( P1_R1162_U160 , P1_R1162_U120 , P1_R1162_U7 , P1_R1162_U81 );
nand NAND2_9215 ( P1_R1162_U161 , P1_R1162_U159 , P1_R1162_U158 );
not NOT1_9216 ( P1_R1162_U162 , P1_R1162_U88 );
or OR2_9217 ( P1_R1162_U163 , P1_U3491 , P1_REG1_REG_13_ );
or OR2_9218 ( P1_R1162_U164 , P1_U3488 , P1_REG1_REG_12_ );
nand NAND2_9219 ( P1_R1162_U165 , P1_R1162_U92 , P1_R1162_U8 );
nand NAND2_9220 ( P1_R1162_U166 , P1_U3491 , P1_REG1_REG_13_ );
nand NAND3_9221 ( P1_R1162_U167 , P1_R1162_U166 , P1_R1162_U91 , P1_R1162_U165 );
or OR2_9222 ( P1_R1162_U168 , P1_REG1_REG_11_ , P1_U3485 );
or OR2_9223 ( P1_R1162_U169 , P1_REG1_REG_13_ , P1_U3491 );
nand NAND3_9224 ( P1_R1162_U170 , P1_R1162_U168 , P1_R1162_U8 , P1_R1162_U88 );
nand NAND2_9225 ( P1_R1162_U171 , P1_R1162_U169 , P1_R1162_U167 );
not NOT1_9226 ( P1_R1162_U172 , P1_R1162_U87 );
or OR2_9227 ( P1_R1162_U173 , P1_REG1_REG_14_ , P1_U3494 );
nand NAND2_9228 ( P1_R1162_U174 , P1_R1162_U173 , P1_R1162_U87 );
nand NAND2_9229 ( P1_R1162_U175 , P1_U3494 , P1_REG1_REG_14_ );
not NOT1_9230 ( P1_R1162_U176 , P1_R1162_U86 );
or OR2_9231 ( P1_R1162_U177 , P1_REG1_REG_15_ , P1_U3497 );
nand NAND2_9232 ( P1_R1162_U178 , P1_R1162_U177 , P1_R1162_U86 );
nand NAND2_9233 ( P1_R1162_U179 , P1_U3497 , P1_REG1_REG_15_ );
not NOT1_9234 ( P1_R1162_U180 , P1_R1162_U66 );
or OR2_9235 ( P1_R1162_U181 , P1_U3503 , P1_REG1_REG_17_ );
or OR2_9236 ( P1_R1162_U182 , P1_U3500 , P1_REG1_REG_16_ );
not NOT1_9237 ( P1_R1162_U183 , P1_R1162_U47 );
nand NAND2_9238 ( P1_R1162_U184 , P1_R1162_U48 , P1_R1162_U47 );
nand NAND2_9239 ( P1_R1162_U185 , P1_U3503 , P1_R1162_U184 );
nand NAND2_9240 ( P1_R1162_U186 , P1_REG1_REG_17_ , P1_R1162_U183 );
nand NAND2_9241 ( P1_R1162_U187 , P1_R1162_U9 , P1_R1162_U66 );
not NOT1_9242 ( P1_R1162_U188 , P1_R1162_U65 );
or OR2_9243 ( P1_R1162_U189 , P1_REG1_REG_18_ , P1_U3506 );
nand NAND2_9244 ( P1_R1162_U190 , P1_R1162_U189 , P1_R1162_U65 );
nand NAND2_9245 ( P1_R1162_U191 , P1_U3506 , P1_REG1_REG_18_ );
nand NAND4_9246 ( P1_R1162_U192 , P1_R1162_U261 , P1_R1162_U260 , P1_R1162_U191 , P1_R1162_U190 );
nand NAND2_9247 ( P1_R1162_U193 , P1_U3506 , P1_REG1_REG_18_ );
nand NAND2_9248 ( P1_R1162_U194 , P1_R1162_U188 , P1_R1162_U193 );
or OR2_9249 ( P1_R1162_U195 , P1_U3506 , P1_REG1_REG_18_ );
nand NAND3_9250 ( P1_R1162_U196 , P1_R1162_U195 , P1_R1162_U264 , P1_R1162_U194 );
or OR2_9251 ( P1_R1162_U197 , P1_REG1_REG_16_ , P1_U3500 );
nand NAND2_9252 ( P1_R1162_U198 , P1_R1162_U197 , P1_R1162_U66 );
nand NAND4_9253 ( P1_R1162_U199 , P1_R1162_U273 , P1_R1162_U272 , P1_R1162_U47 , P1_R1162_U198 );
nand NAND2_9254 ( P1_R1162_U200 , P1_R1162_U180 , P1_R1162_U47 );
nand NAND2_9255 ( P1_R1162_U201 , P1_REG1_REG_17_ , P1_U3503 );
nand NAND3_9256 ( P1_R1162_U202 , P1_R1162_U201 , P1_R1162_U9 , P1_R1162_U200 );
or OR2_9257 ( P1_R1162_U203 , P1_U3500 , P1_REG1_REG_16_ );
nand NAND2_9258 ( P1_R1162_U204 , P1_R1162_U168 , P1_R1162_U88 );
not NOT1_9259 ( P1_R1162_U205 , P1_R1162_U67 );
or OR2_9260 ( P1_R1162_U206 , P1_REG1_REG_12_ , P1_U3488 );
nand NAND2_9261 ( P1_R1162_U207 , P1_R1162_U206 , P1_R1162_U67 );
nand NAND4_9262 ( P1_R1162_U208 , P1_R1162_U294 , P1_R1162_U293 , P1_R1162_U91 , P1_R1162_U207 );
nand NAND2_9263 ( P1_R1162_U209 , P1_R1162_U205 , P1_R1162_U91 );
nand NAND2_9264 ( P1_R1162_U210 , P1_U3491 , P1_REG1_REG_13_ );
nand NAND3_9265 ( P1_R1162_U211 , P1_R1162_U210 , P1_R1162_U8 , P1_R1162_U209 );
or OR2_9266 ( P1_R1162_U212 , P1_U3488 , P1_REG1_REG_12_ );
or OR2_9267 ( P1_R1162_U213 , P1_REG1_REG_9_ , P1_U3479 );
nand NAND2_9268 ( P1_R1162_U214 , P1_R1162_U213 , P1_R1162_U38 );
nand NAND4_9269 ( P1_R1162_U215 , P1_R1162_U306 , P1_R1162_U305 , P1_R1162_U90 , P1_R1162_U214 );
nand NAND2_9270 ( P1_R1162_U216 , P1_R1162_U122 , P1_R1162_U90 );
nand NAND2_9271 ( P1_R1162_U217 , P1_U3482 , P1_REG1_REG_10_ );
nand NAND3_9272 ( P1_R1162_U218 , P1_R1162_U217 , P1_R1162_U7 , P1_R1162_U216 );
nand NAND2_9273 ( P1_R1162_U219 , P1_R1162_U123 , P1_R1162_U90 );
nand NAND2_9274 ( P1_R1162_U220 , P1_R1162_U120 , P1_R1162_U49 );
nand NAND2_9275 ( P1_R1162_U221 , P1_R1162_U130 , P1_R1162_U20 );
nand NAND2_9276 ( P1_R1162_U222 , P1_R1162_U144 , P1_R1162_U32 );
nand NAND2_9277 ( P1_R1162_U223 , P1_R1162_U147 , P1_R1162_U96 );
nand NAND2_9278 ( P1_R1162_U224 , P1_R1162_U203 , P1_R1162_U47 );
nand NAND2_9279 ( P1_R1162_U225 , P1_R1162_U212 , P1_R1162_U91 );
nand NAND2_9280 ( P1_R1162_U226 , P1_R1162_U168 , P1_R1162_U56 );
nand NAND2_9281 ( P1_R1162_U227 , P1_U3479 , P1_R1162_U37 );
nand NAND2_9282 ( P1_R1162_U228 , P1_REG1_REG_9_ , P1_R1162_U36 );
nand NAND2_9283 ( P1_R1162_U229 , P1_R1162_U228 , P1_R1162_U227 );
nand NAND2_9284 ( P1_R1162_U230 , P1_R1162_U219 , P1_R1162_U38 );
nand NAND2_9285 ( P1_R1162_U231 , P1_R1162_U229 , P1_R1162_U122 );
nand NAND2_9286 ( P1_R1162_U232 , P1_U3476 , P1_R1162_U34 );
nand NAND2_9287 ( P1_R1162_U233 , P1_REG1_REG_8_ , P1_R1162_U35 );
nand NAND2_9288 ( P1_R1162_U234 , P1_R1162_U233 , P1_R1162_U232 );
nand NAND2_9289 ( P1_R1162_U235 , P1_R1162_U220 , P1_R1162_U81 );
nand NAND2_9290 ( P1_R1162_U236 , P1_R1162_U119 , P1_R1162_U234 );
nand NAND2_9291 ( P1_R1162_U237 , P1_U3473 , P1_R1162_U21 );
nand NAND2_9292 ( P1_R1162_U238 , P1_REG1_REG_7_ , P1_R1162_U19 );
nand NAND2_9293 ( P1_R1162_U239 , P1_U3470 , P1_R1162_U17 );
nand NAND2_9294 ( P1_R1162_U240 , P1_REG1_REG_6_ , P1_R1162_U18 );
nand NAND2_9295 ( P1_R1162_U241 , P1_R1162_U240 , P1_R1162_U239 );
nand NAND2_9296 ( P1_R1162_U242 , P1_R1162_U221 , P1_R1162_U39 );
nand NAND2_9297 ( P1_R1162_U243 , P1_R1162_U241 , P1_R1162_U111 );
nand NAND2_9298 ( P1_R1162_U244 , P1_U3467 , P1_R1162_U33 );
nand NAND2_9299 ( P1_R1162_U245 , P1_REG1_REG_5_ , P1_R1162_U24 );
nand NAND2_9300 ( P1_R1162_U246 , P1_U3464 , P1_R1162_U22 );
nand NAND2_9301 ( P1_R1162_U247 , P1_REG1_REG_4_ , P1_R1162_U23 );
nand NAND2_9302 ( P1_R1162_U248 , P1_R1162_U247 , P1_R1162_U246 );
nand NAND2_9303 ( P1_R1162_U249 , P1_R1162_U222 , P1_R1162_U42 );
nand NAND2_9304 ( P1_R1162_U250 , P1_R1162_U248 , P1_R1162_U137 );
nand NAND2_9305 ( P1_R1162_U251 , P1_U3461 , P1_R1162_U30 );
nand NAND2_9306 ( P1_R1162_U252 , P1_REG1_REG_3_ , P1_R1162_U31 );
nand NAND2_9307 ( P1_R1162_U253 , P1_R1162_U252 , P1_R1162_U251 );
nand NAND2_9308 ( P1_R1162_U254 , P1_R1162_U223 , P1_R1162_U82 );
nand NAND2_9309 ( P1_R1162_U255 , P1_R1162_U146 , P1_R1162_U253 );
nand NAND2_9310 ( P1_R1162_U256 , P1_U3458 , P1_R1162_U25 );
nand NAND2_9311 ( P1_R1162_U257 , P1_REG1_REG_2_ , P1_R1162_U26 );
nand NAND2_9312 ( P1_R1162_U258 , P1_R1162_U98 , P1_R1162_U83 );
nand NAND2_9313 ( P1_R1162_U259 , P1_R1162_U153 , P1_R1162_U29 );
nand NAND2_9314 ( P1_R1162_U260 , P1_U3443 , P1_R1162_U85 );
nand NAND2_9315 ( P1_R1162_U261 , P1_REG1_REG_19_ , P1_R1162_U84 );
nand NAND2_9316 ( P1_R1162_U262 , P1_U3443 , P1_R1162_U85 );
nand NAND2_9317 ( P1_R1162_U263 , P1_REG1_REG_19_ , P1_R1162_U84 );
nand NAND2_9318 ( P1_R1162_U264 , P1_R1162_U263 , P1_R1162_U262 );
nand NAND2_9319 ( P1_R1162_U265 , P1_U3506 , P1_R1162_U63 );
nand NAND2_9320 ( P1_R1162_U266 , P1_REG1_REG_18_ , P1_R1162_U64 );
nand NAND2_9321 ( P1_R1162_U267 , P1_U3506 , P1_R1162_U63 );
nand NAND2_9322 ( P1_R1162_U268 , P1_REG1_REG_18_ , P1_R1162_U64 );
nand NAND2_9323 ( P1_R1162_U269 , P1_R1162_U268 , P1_R1162_U267 );
nand NAND3_9324 ( P1_R1162_U270 , P1_R1162_U266 , P1_R1162_U265 , P1_R1162_U65 );
nand NAND2_9325 ( P1_R1162_U271 , P1_R1162_U269 , P1_R1162_U188 );
nand NAND2_9326 ( P1_R1162_U272 , P1_U3503 , P1_R1162_U48 );
nand NAND2_9327 ( P1_R1162_U273 , P1_REG1_REG_17_ , P1_R1162_U46 );
nand NAND2_9328 ( P1_R1162_U274 , P1_U3500 , P1_R1162_U44 );
nand NAND2_9329 ( P1_R1162_U275 , P1_REG1_REG_16_ , P1_R1162_U45 );
nand NAND2_9330 ( P1_R1162_U276 , P1_R1162_U275 , P1_R1162_U274 );
nand NAND2_9331 ( P1_R1162_U277 , P1_R1162_U224 , P1_R1162_U66 );
nand NAND2_9332 ( P1_R1162_U278 , P1_R1162_U276 , P1_R1162_U180 );
nand NAND2_9333 ( P1_R1162_U279 , P1_U3497 , P1_R1162_U61 );
nand NAND2_9334 ( P1_R1162_U280 , P1_REG1_REG_15_ , P1_R1162_U62 );
nand NAND2_9335 ( P1_R1162_U281 , P1_U3497 , P1_R1162_U61 );
nand NAND2_9336 ( P1_R1162_U282 , P1_REG1_REG_15_ , P1_R1162_U62 );
nand NAND2_9337 ( P1_R1162_U283 , P1_R1162_U282 , P1_R1162_U281 );
nand NAND3_9338 ( P1_R1162_U284 , P1_R1162_U280 , P1_R1162_U279 , P1_R1162_U86 );
nand NAND2_9339 ( P1_R1162_U285 , P1_R1162_U176 , P1_R1162_U283 );
nand NAND2_9340 ( P1_R1162_U286 , P1_U3494 , P1_R1162_U59 );
nand NAND2_9341 ( P1_R1162_U287 , P1_REG1_REG_14_ , P1_R1162_U60 );
nand NAND2_9342 ( P1_R1162_U288 , P1_U3494 , P1_R1162_U59 );
nand NAND2_9343 ( P1_R1162_U289 , P1_REG1_REG_14_ , P1_R1162_U60 );
nand NAND2_9344 ( P1_R1162_U290 , P1_R1162_U289 , P1_R1162_U288 );
nand NAND3_9345 ( P1_R1162_U291 , P1_R1162_U287 , P1_R1162_U286 , P1_R1162_U87 );
nand NAND2_9346 ( P1_R1162_U292 , P1_R1162_U172 , P1_R1162_U290 );
nand NAND2_9347 ( P1_R1162_U293 , P1_U3491 , P1_R1162_U57 );
nand NAND2_9348 ( P1_R1162_U294 , P1_REG1_REG_13_ , P1_R1162_U58 );
nand NAND2_9349 ( P1_R1162_U295 , P1_U3488 , P1_R1162_U52 );
nand NAND2_9350 ( P1_R1162_U296 , P1_REG1_REG_12_ , P1_R1162_U53 );
nand NAND2_9351 ( P1_R1162_U297 , P1_R1162_U296 , P1_R1162_U295 );
nand NAND2_9352 ( P1_R1162_U298 , P1_R1162_U225 , P1_R1162_U67 );
nand NAND2_9353 ( P1_R1162_U299 , P1_R1162_U297 , P1_R1162_U205 );
nand NAND2_9354 ( P1_R1162_U300 , P1_U3485 , P1_R1162_U54 );
nand NAND2_9355 ( P1_R1162_U301 , P1_REG1_REG_11_ , P1_R1162_U55 );
nand NAND2_9356 ( P1_R1162_U302 , P1_R1162_U301 , P1_R1162_U300 );
nand NAND2_9357 ( P1_R1162_U303 , P1_R1162_U226 , P1_R1162_U88 );
nand NAND2_9358 ( P1_R1162_U304 , P1_R1162_U162 , P1_R1162_U302 );
nand NAND2_9359 ( P1_R1162_U305 , P1_U3482 , P1_R1162_U50 );
nand NAND2_9360 ( P1_R1162_U306 , P1_REG1_REG_10_ , P1_R1162_U51 );
nand NAND2_9361 ( P1_R1162_U307 , P1_U3449 , P1_R1162_U27 );
nand NAND2_9362 ( P1_R1162_U308 , P1_REG1_REG_0_ , P1_R1162_U28 );
and AND2_9363 ( P1_R1117_U6 , P1_R1117_U184 , P1_R1117_U201 );
and AND2_9364 ( P1_R1117_U7 , P1_R1117_U203 , P1_R1117_U202 );
and AND2_9365 ( P1_R1117_U8 , P1_R1117_U179 , P1_R1117_U240 );
and AND2_9366 ( P1_R1117_U9 , P1_R1117_U242 , P1_R1117_U241 );
and AND2_9367 ( P1_R1117_U10 , P1_R1117_U259 , P1_R1117_U258 );
and AND2_9368 ( P1_R1117_U11 , P1_R1117_U285 , P1_R1117_U284 );
and AND2_9369 ( P1_R1117_U12 , P1_R1117_U383 , P1_R1117_U382 );
nand NAND2_9370 ( P1_R1117_U13 , P1_R1117_U340 , P1_R1117_U343 );
nand NAND2_9371 ( P1_R1117_U14 , P1_R1117_U329 , P1_R1117_U332 );
nand NAND2_9372 ( P1_R1117_U15 , P1_R1117_U318 , P1_R1117_U321 );
nand NAND2_9373 ( P1_R1117_U16 , P1_R1117_U310 , P1_R1117_U312 );
nand NAND3_9374 ( P1_R1117_U17 , P1_R1117_U156 , P1_R1117_U175 , P1_R1117_U348 );
nand NAND2_9375 ( P1_R1117_U18 , P1_R1117_U236 , P1_R1117_U238 );
nand NAND2_9376 ( P1_R1117_U19 , P1_R1117_U228 , P1_R1117_U231 );
nand NAND2_9377 ( P1_R1117_U20 , P1_R1117_U220 , P1_R1117_U222 );
nand NAND2_9378 ( P1_R1117_U21 , P1_R1117_U25 , P1_R1117_U346 );
not NOT1_9379 ( P1_R1117_U22 , P1_U3474 );
not NOT1_9380 ( P1_R1117_U23 , P1_U3459 );
not NOT1_9381 ( P1_R1117_U24 , P1_U3451 );
nand NAND2_9382 ( P1_R1117_U25 , P1_U3451 , P1_R1117_U93 );
not NOT1_9383 ( P1_R1117_U26 , P1_U3076 );
not NOT1_9384 ( P1_R1117_U27 , P1_U3462 );
not NOT1_9385 ( P1_R1117_U28 , P1_U3066 );
nand NAND2_9386 ( P1_R1117_U29 , P1_U3066 , P1_R1117_U23 );
not NOT1_9387 ( P1_R1117_U30 , P1_U3062 );
not NOT1_9388 ( P1_R1117_U31 , P1_U3471 );
not NOT1_9389 ( P1_R1117_U32 , P1_U3468 );
not NOT1_9390 ( P1_R1117_U33 , P1_U3465 );
not NOT1_9391 ( P1_R1117_U34 , P1_U3069 );
not NOT1_9392 ( P1_R1117_U35 , P1_U3065 );
not NOT1_9393 ( P1_R1117_U36 , P1_U3058 );
nand NAND2_9394 ( P1_R1117_U37 , P1_U3058 , P1_R1117_U33 );
not NOT1_9395 ( P1_R1117_U38 , P1_U3477 );
not NOT1_9396 ( P1_R1117_U39 , P1_U3068 );
nand NAND2_9397 ( P1_R1117_U40 , P1_U3068 , P1_R1117_U22 );
not NOT1_9398 ( P1_R1117_U41 , P1_U3082 );
not NOT1_9399 ( P1_R1117_U42 , P1_U3480 );
not NOT1_9400 ( P1_R1117_U43 , P1_U3081 );
nand NAND2_9401 ( P1_R1117_U44 , P1_R1117_U209 , P1_R1117_U208 );
nand NAND2_9402 ( P1_R1117_U45 , P1_R1117_U37 , P1_R1117_U224 );
nand NAND2_9403 ( P1_R1117_U46 , P1_R1117_U193 , P1_R1117_U192 );
not NOT1_9404 ( P1_R1117_U47 , P1_U4009 );
not NOT1_9405 ( P1_R1117_U48 , P1_U4013 );
not NOT1_9406 ( P1_R1117_U49 , P1_U3498 );
not NOT1_9407 ( P1_R1117_U50 , P1_U3486 );
not NOT1_9408 ( P1_R1117_U51 , P1_U3483 );
not NOT1_9409 ( P1_R1117_U52 , P1_U3061 );
not NOT1_9410 ( P1_R1117_U53 , P1_U3060 );
nand NAND2_9411 ( P1_R1117_U54 , P1_U3081 , P1_R1117_U42 );
not NOT1_9412 ( P1_R1117_U55 , P1_U3489 );
not NOT1_9413 ( P1_R1117_U56 , P1_U3070 );
not NOT1_9414 ( P1_R1117_U57 , P1_U3492 );
not NOT1_9415 ( P1_R1117_U58 , P1_U3078 );
not NOT1_9416 ( P1_R1117_U59 , P1_U3501 );
not NOT1_9417 ( P1_R1117_U60 , P1_U3495 );
not NOT1_9418 ( P1_R1117_U61 , P1_U3071 );
not NOT1_9419 ( P1_R1117_U62 , P1_U3072 );
not NOT1_9420 ( P1_R1117_U63 , P1_U3077 );
nand NAND2_9421 ( P1_R1117_U64 , P1_U3077 , P1_R1117_U60 );
not NOT1_9422 ( P1_R1117_U65 , P1_U3504 );
not NOT1_9423 ( P1_R1117_U66 , P1_U3067 );
nand NAND2_9424 ( P1_R1117_U67 , P1_R1117_U269 , P1_R1117_U268 );
not NOT1_9425 ( P1_R1117_U68 , P1_U3080 );
not NOT1_9426 ( P1_R1117_U69 , P1_U3509 );
not NOT1_9427 ( P1_R1117_U70 , P1_U3079 );
not NOT1_9428 ( P1_R1117_U71 , P1_U4015 );
not NOT1_9429 ( P1_R1117_U72 , P1_U3074 );
not NOT1_9430 ( P1_R1117_U73 , P1_U4012 );
not NOT1_9431 ( P1_R1117_U74 , P1_U4014 );
not NOT1_9432 ( P1_R1117_U75 , P1_U3064 );
not NOT1_9433 ( P1_R1117_U76 , P1_U3059 );
not NOT1_9434 ( P1_R1117_U77 , P1_U3073 );
nand NAND2_9435 ( P1_R1117_U78 , P1_U3073 , P1_R1117_U74 );
not NOT1_9436 ( P1_R1117_U79 , P1_U4011 );
not NOT1_9437 ( P1_R1117_U80 , P1_U3063 );
not NOT1_9438 ( P1_R1117_U81 , P1_U4010 );
not NOT1_9439 ( P1_R1117_U82 , P1_U3056 );
not NOT1_9440 ( P1_R1117_U83 , P1_U4008 );
not NOT1_9441 ( P1_R1117_U84 , P1_U3055 );
nand NAND2_9442 ( P1_R1117_U85 , P1_U3055 , P1_R1117_U47 );
not NOT1_9443 ( P1_R1117_U86 , P1_U3051 );
not NOT1_9444 ( P1_R1117_U87 , P1_U4007 );
not NOT1_9445 ( P1_R1117_U88 , P1_U3052 );
nand NAND2_9446 ( P1_R1117_U89 , P1_R1117_U299 , P1_R1117_U298 );
nand NAND2_9447 ( P1_R1117_U90 , P1_R1117_U78 , P1_R1117_U314 );
nand NAND2_9448 ( P1_R1117_U91 , P1_R1117_U64 , P1_R1117_U325 );
nand NAND2_9449 ( P1_R1117_U92 , P1_R1117_U54 , P1_R1117_U336 );
not NOT1_9450 ( P1_R1117_U93 , P1_U3075 );
nand NAND2_9451 ( P1_R1117_U94 , P1_R1117_U393 , P1_R1117_U392 );
nand NAND2_9452 ( P1_R1117_U95 , P1_R1117_U407 , P1_R1117_U406 );
nand NAND2_9453 ( P1_R1117_U96 , P1_R1117_U412 , P1_R1117_U411 );
nand NAND2_9454 ( P1_R1117_U97 , P1_R1117_U428 , P1_R1117_U427 );
nand NAND2_9455 ( P1_R1117_U98 , P1_R1117_U433 , P1_R1117_U432 );
nand NAND2_9456 ( P1_R1117_U99 , P1_R1117_U438 , P1_R1117_U437 );
nand NAND2_9457 ( P1_R1117_U100 , P1_R1117_U443 , P1_R1117_U442 );
nand NAND2_9458 ( P1_R1117_U101 , P1_R1117_U448 , P1_R1117_U447 );
nand NAND2_9459 ( P1_R1117_U102 , P1_R1117_U464 , P1_R1117_U463 );
nand NAND2_9460 ( P1_R1117_U103 , P1_R1117_U469 , P1_R1117_U468 );
nand NAND2_9461 ( P1_R1117_U104 , P1_R1117_U352 , P1_R1117_U351 );
nand NAND2_9462 ( P1_R1117_U105 , P1_R1117_U361 , P1_R1117_U360 );
nand NAND2_9463 ( P1_R1117_U106 , P1_R1117_U368 , P1_R1117_U367 );
nand NAND2_9464 ( P1_R1117_U107 , P1_R1117_U372 , P1_R1117_U371 );
nand NAND2_9465 ( P1_R1117_U108 , P1_R1117_U381 , P1_R1117_U380 );
nand NAND2_9466 ( P1_R1117_U109 , P1_R1117_U402 , P1_R1117_U401 );
nand NAND2_9467 ( P1_R1117_U110 , P1_R1117_U419 , P1_R1117_U418 );
nand NAND2_9468 ( P1_R1117_U111 , P1_R1117_U423 , P1_R1117_U422 );
nand NAND2_9469 ( P1_R1117_U112 , P1_R1117_U455 , P1_R1117_U454 );
nand NAND2_9470 ( P1_R1117_U113 , P1_R1117_U459 , P1_R1117_U458 );
nand NAND2_9471 ( P1_R1117_U114 , P1_R1117_U476 , P1_R1117_U475 );
and AND2_9472 ( P1_R1117_U115 , P1_R1117_U195 , P1_R1117_U183 );
and AND2_9473 ( P1_R1117_U116 , P1_R1117_U198 , P1_R1117_U199 );
and AND2_9474 ( P1_R1117_U117 , P1_R1117_U211 , P1_R1117_U185 );
and AND2_9475 ( P1_R1117_U118 , P1_R1117_U214 , P1_R1117_U215 );
and AND3_9476 ( P1_R1117_U119 , P1_R1117_U354 , P1_R1117_U353 , P1_R1117_U40 );
and AND2_9477 ( P1_R1117_U120 , P1_R1117_U357 , P1_R1117_U185 );
and AND2_9478 ( P1_R1117_U121 , P1_R1117_U230 , P1_R1117_U7 );
and AND2_9479 ( P1_R1117_U122 , P1_R1117_U364 , P1_R1117_U184 );
and AND3_9480 ( P1_R1117_U123 , P1_R1117_U374 , P1_R1117_U373 , P1_R1117_U29 );
and AND2_9481 ( P1_R1117_U124 , P1_R1117_U377 , P1_R1117_U183 );
and AND2_9482 ( P1_R1117_U125 , P1_R1117_U217 , P1_R1117_U8 );
and AND2_9483 ( P1_R1117_U126 , P1_R1117_U262 , P1_R1117_U180 );
and AND2_9484 ( P1_R1117_U127 , P1_R1117_U288 , P1_R1117_U181 );
and AND2_9485 ( P1_R1117_U128 , P1_R1117_U304 , P1_R1117_U305 );
and AND2_9486 ( P1_R1117_U129 , P1_R1117_U307 , P1_R1117_U386 );
and AND3_9487 ( P1_R1117_U130 , P1_R1117_U305 , P1_R1117_U304 , P1_R1117_U308 );
nand NAND2_9488 ( P1_R1117_U131 , P1_R1117_U390 , P1_R1117_U389 );
and AND3_9489 ( P1_R1117_U132 , P1_R1117_U395 , P1_R1117_U394 , P1_R1117_U85 );
and AND2_9490 ( P1_R1117_U133 , P1_R1117_U398 , P1_R1117_U182 );
nand NAND2_9491 ( P1_R1117_U134 , P1_R1117_U404 , P1_R1117_U403 );
nand NAND2_9492 ( P1_R1117_U135 , P1_R1117_U409 , P1_R1117_U408 );
and AND2_9493 ( P1_R1117_U136 , P1_R1117_U415 , P1_R1117_U181 );
nand NAND2_9494 ( P1_R1117_U137 , P1_R1117_U425 , P1_R1117_U424 );
nand NAND2_9495 ( P1_R1117_U138 , P1_R1117_U430 , P1_R1117_U429 );
nand NAND2_9496 ( P1_R1117_U139 , P1_R1117_U435 , P1_R1117_U434 );
nand NAND2_9497 ( P1_R1117_U140 , P1_R1117_U440 , P1_R1117_U439 );
nand NAND2_9498 ( P1_R1117_U141 , P1_R1117_U445 , P1_R1117_U444 );
and AND2_9499 ( P1_R1117_U142 , P1_R1117_U451 , P1_R1117_U180 );
nand NAND2_9500 ( P1_R1117_U143 , P1_R1117_U461 , P1_R1117_U460 );
nand NAND2_9501 ( P1_R1117_U144 , P1_R1117_U466 , P1_R1117_U465 );
and AND2_9502 ( P1_R1117_U145 , P1_R1117_U342 , P1_R1117_U9 );
and AND2_9503 ( P1_R1117_U146 , P1_R1117_U472 , P1_R1117_U179 );
and AND2_9504 ( P1_R1117_U147 , P1_R1117_U350 , P1_R1117_U349 );
nand NAND2_9505 ( P1_R1117_U148 , P1_R1117_U118 , P1_R1117_U212 );
and AND2_9506 ( P1_R1117_U149 , P1_R1117_U359 , P1_R1117_U358 );
and AND2_9507 ( P1_R1117_U150 , P1_R1117_U366 , P1_R1117_U365 );
and AND2_9508 ( P1_R1117_U151 , P1_R1117_U370 , P1_R1117_U369 );
nand NAND2_9509 ( P1_R1117_U152 , P1_R1117_U116 , P1_R1117_U196 );
and AND2_9510 ( P1_R1117_U153 , P1_R1117_U379 , P1_R1117_U378 );
not NOT1_9511 ( P1_R1117_U154 , P1_U4018 );
not NOT1_9512 ( P1_R1117_U155 , P1_U3053 );
and AND2_9513 ( P1_R1117_U156 , P1_R1117_U388 , P1_R1117_U387 );
nand NAND2_9514 ( P1_R1117_U157 , P1_R1117_U128 , P1_R1117_U302 );
and AND2_9515 ( P1_R1117_U158 , P1_R1117_U400 , P1_R1117_U399 );
nand NAND2_9516 ( P1_R1117_U159 , P1_R1117_U295 , P1_R1117_U294 );
nand NAND2_9517 ( P1_R1117_U160 , P1_R1117_U291 , P1_R1117_U290 );
and AND2_9518 ( P1_R1117_U161 , P1_R1117_U417 , P1_R1117_U416 );
and AND2_9519 ( P1_R1117_U162 , P1_R1117_U421 , P1_R1117_U420 );
nand NAND2_9520 ( P1_R1117_U163 , P1_R1117_U281 , P1_R1117_U280 );
nand NAND2_9521 ( P1_R1117_U164 , P1_R1117_U277 , P1_R1117_U276 );
not NOT1_9522 ( P1_R1117_U165 , P1_U3456 );
nand NAND2_9523 ( P1_R1117_U166 , P1_R1117_U273 , P1_R1117_U272 );
not NOT1_9524 ( P1_R1117_U167 , P1_U3507 );
nand NAND2_9525 ( P1_R1117_U168 , P1_R1117_U265 , P1_R1117_U264 );
and AND2_9526 ( P1_R1117_U169 , P1_R1117_U453 , P1_R1117_U452 );
and AND2_9527 ( P1_R1117_U170 , P1_R1117_U457 , P1_R1117_U456 );
nand NAND2_9528 ( P1_R1117_U171 , P1_R1117_U255 , P1_R1117_U254 );
nand NAND2_9529 ( P1_R1117_U172 , P1_R1117_U251 , P1_R1117_U250 );
nand NAND2_9530 ( P1_R1117_U173 , P1_R1117_U247 , P1_R1117_U246 );
and AND2_9531 ( P1_R1117_U174 , P1_R1117_U474 , P1_R1117_U473 );
nand NAND2_9532 ( P1_R1117_U175 , P1_R1117_U129 , P1_R1117_U157 );
not NOT1_9533 ( P1_R1117_U176 , P1_R1117_U85 );
not NOT1_9534 ( P1_R1117_U177 , P1_R1117_U29 );
not NOT1_9535 ( P1_R1117_U178 , P1_R1117_U40 );
nand NAND2_9536 ( P1_R1117_U179 , P1_U3483 , P1_R1117_U53 );
nand NAND2_9537 ( P1_R1117_U180 , P1_U3498 , P1_R1117_U62 );
nand NAND2_9538 ( P1_R1117_U181 , P1_U4013 , P1_R1117_U76 );
nand NAND2_9539 ( P1_R1117_U182 , P1_U4009 , P1_R1117_U84 );
nand NAND2_9540 ( P1_R1117_U183 , P1_U3459 , P1_R1117_U28 );
nand NAND2_9541 ( P1_R1117_U184 , P1_U3468 , P1_R1117_U35 );
nand NAND2_9542 ( P1_R1117_U185 , P1_U3474 , P1_R1117_U39 );
not NOT1_9543 ( P1_R1117_U186 , P1_R1117_U64 );
not NOT1_9544 ( P1_R1117_U187 , P1_R1117_U78 );
not NOT1_9545 ( P1_R1117_U188 , P1_R1117_U37 );
not NOT1_9546 ( P1_R1117_U189 , P1_R1117_U54 );
not NOT1_9547 ( P1_R1117_U190 , P1_R1117_U25 );
nand NAND2_9548 ( P1_R1117_U191 , P1_R1117_U190 , P1_R1117_U26 );
nand NAND2_9549 ( P1_R1117_U192 , P1_R1117_U191 , P1_R1117_U165 );
nand NAND2_9550 ( P1_R1117_U193 , P1_U3076 , P1_R1117_U25 );
not NOT1_9551 ( P1_R1117_U194 , P1_R1117_U46 );
nand NAND2_9552 ( P1_R1117_U195 , P1_U3462 , P1_R1117_U30 );
nand NAND2_9553 ( P1_R1117_U196 , P1_R1117_U115 , P1_R1117_U46 );
nand NAND2_9554 ( P1_R1117_U197 , P1_R1117_U30 , P1_R1117_U29 );
nand NAND2_9555 ( P1_R1117_U198 , P1_R1117_U197 , P1_R1117_U27 );
nand NAND2_9556 ( P1_R1117_U199 , P1_U3062 , P1_R1117_U177 );
not NOT1_9557 ( P1_R1117_U200 , P1_R1117_U152 );
nand NAND2_9558 ( P1_R1117_U201 , P1_U3471 , P1_R1117_U34 );
nand NAND2_9559 ( P1_R1117_U202 , P1_U3069 , P1_R1117_U31 );
nand NAND2_9560 ( P1_R1117_U203 , P1_U3065 , P1_R1117_U32 );
nand NAND2_9561 ( P1_R1117_U204 , P1_R1117_U188 , P1_R1117_U6 );
nand NAND2_9562 ( P1_R1117_U205 , P1_R1117_U7 , P1_R1117_U204 );
nand NAND2_9563 ( P1_R1117_U206 , P1_U3465 , P1_R1117_U36 );
nand NAND2_9564 ( P1_R1117_U207 , P1_U3471 , P1_R1117_U34 );
nand NAND3_9565 ( P1_R1117_U208 , P1_R1117_U206 , P1_R1117_U152 , P1_R1117_U6 );
nand NAND2_9566 ( P1_R1117_U209 , P1_R1117_U207 , P1_R1117_U205 );
not NOT1_9567 ( P1_R1117_U210 , P1_R1117_U44 );
nand NAND2_9568 ( P1_R1117_U211 , P1_U3477 , P1_R1117_U41 );
nand NAND2_9569 ( P1_R1117_U212 , P1_R1117_U117 , P1_R1117_U44 );
nand NAND2_9570 ( P1_R1117_U213 , P1_R1117_U41 , P1_R1117_U40 );
nand NAND2_9571 ( P1_R1117_U214 , P1_R1117_U213 , P1_R1117_U38 );
nand NAND2_9572 ( P1_R1117_U215 , P1_U3082 , P1_R1117_U178 );
not NOT1_9573 ( P1_R1117_U216 , P1_R1117_U148 );
nand NAND2_9574 ( P1_R1117_U217 , P1_U3480 , P1_R1117_U43 );
nand NAND2_9575 ( P1_R1117_U218 , P1_R1117_U217 , P1_R1117_U54 );
nand NAND2_9576 ( P1_R1117_U219 , P1_R1117_U210 , P1_R1117_U40 );
nand NAND2_9577 ( P1_R1117_U220 , P1_R1117_U120 , P1_R1117_U219 );
nand NAND2_9578 ( P1_R1117_U221 , P1_R1117_U44 , P1_R1117_U185 );
nand NAND2_9579 ( P1_R1117_U222 , P1_R1117_U119 , P1_R1117_U221 );
nand NAND2_9580 ( P1_R1117_U223 , P1_R1117_U40 , P1_R1117_U185 );
nand NAND2_9581 ( P1_R1117_U224 , P1_R1117_U206 , P1_R1117_U152 );
not NOT1_9582 ( P1_R1117_U225 , P1_R1117_U45 );
nand NAND2_9583 ( P1_R1117_U226 , P1_U3065 , P1_R1117_U32 );
nand NAND2_9584 ( P1_R1117_U227 , P1_R1117_U225 , P1_R1117_U226 );
nand NAND2_9585 ( P1_R1117_U228 , P1_R1117_U122 , P1_R1117_U227 );
nand NAND2_9586 ( P1_R1117_U229 , P1_R1117_U45 , P1_R1117_U184 );
nand NAND2_9587 ( P1_R1117_U230 , P1_U3471 , P1_R1117_U34 );
nand NAND2_9588 ( P1_R1117_U231 , P1_R1117_U121 , P1_R1117_U229 );
nand NAND2_9589 ( P1_R1117_U232 , P1_U3065 , P1_R1117_U32 );
nand NAND2_9590 ( P1_R1117_U233 , P1_R1117_U184 , P1_R1117_U232 );
nand NAND2_9591 ( P1_R1117_U234 , P1_R1117_U206 , P1_R1117_U37 );
nand NAND2_9592 ( P1_R1117_U235 , P1_R1117_U194 , P1_R1117_U29 );
nand NAND2_9593 ( P1_R1117_U236 , P1_R1117_U124 , P1_R1117_U235 );
nand NAND2_9594 ( P1_R1117_U237 , P1_R1117_U46 , P1_R1117_U183 );
nand NAND2_9595 ( P1_R1117_U238 , P1_R1117_U123 , P1_R1117_U237 );
nand NAND2_9596 ( P1_R1117_U239 , P1_R1117_U29 , P1_R1117_U183 );
nand NAND2_9597 ( P1_R1117_U240 , P1_U3486 , P1_R1117_U52 );
nand NAND2_9598 ( P1_R1117_U241 , P1_U3061 , P1_R1117_U50 );
nand NAND2_9599 ( P1_R1117_U242 , P1_U3060 , P1_R1117_U51 );
nand NAND2_9600 ( P1_R1117_U243 , P1_R1117_U189 , P1_R1117_U8 );
nand NAND2_9601 ( P1_R1117_U244 , P1_R1117_U9 , P1_R1117_U243 );
nand NAND2_9602 ( P1_R1117_U245 , P1_U3486 , P1_R1117_U52 );
nand NAND2_9603 ( P1_R1117_U246 , P1_R1117_U125 , P1_R1117_U148 );
nand NAND2_9604 ( P1_R1117_U247 , P1_R1117_U245 , P1_R1117_U244 );
not NOT1_9605 ( P1_R1117_U248 , P1_R1117_U173 );
nand NAND2_9606 ( P1_R1117_U249 , P1_U3489 , P1_R1117_U56 );
nand NAND2_9607 ( P1_R1117_U250 , P1_R1117_U249 , P1_R1117_U173 );
nand NAND2_9608 ( P1_R1117_U251 , P1_U3070 , P1_R1117_U55 );
not NOT1_9609 ( P1_R1117_U252 , P1_R1117_U172 );
nand NAND2_9610 ( P1_R1117_U253 , P1_U3492 , P1_R1117_U58 );
nand NAND2_9611 ( P1_R1117_U254 , P1_R1117_U253 , P1_R1117_U172 );
nand NAND2_9612 ( P1_R1117_U255 , P1_U3078 , P1_R1117_U57 );
not NOT1_9613 ( P1_R1117_U256 , P1_R1117_U171 );
nand NAND2_9614 ( P1_R1117_U257 , P1_U3501 , P1_R1117_U61 );
nand NAND2_9615 ( P1_R1117_U258 , P1_U3071 , P1_R1117_U59 );
nand NAND2_9616 ( P1_R1117_U259 , P1_U3072 , P1_R1117_U49 );
nand NAND2_9617 ( P1_R1117_U260 , P1_R1117_U186 , P1_R1117_U180 );
nand NAND2_9618 ( P1_R1117_U261 , P1_R1117_U10 , P1_R1117_U260 );
nand NAND2_9619 ( P1_R1117_U262 , P1_U3495 , P1_R1117_U63 );
nand NAND2_9620 ( P1_R1117_U263 , P1_U3501 , P1_R1117_U61 );
nand NAND3_9621 ( P1_R1117_U264 , P1_R1117_U171 , P1_R1117_U126 , P1_R1117_U257 );
nand NAND2_9622 ( P1_R1117_U265 , P1_R1117_U263 , P1_R1117_U261 );
not NOT1_9623 ( P1_R1117_U266 , P1_R1117_U168 );
nand NAND2_9624 ( P1_R1117_U267 , P1_U3504 , P1_R1117_U66 );
nand NAND2_9625 ( P1_R1117_U268 , P1_R1117_U267 , P1_R1117_U168 );
nand NAND2_9626 ( P1_R1117_U269 , P1_U3067 , P1_R1117_U65 );
not NOT1_9627 ( P1_R1117_U270 , P1_R1117_U67 );
nand NAND2_9628 ( P1_R1117_U271 , P1_R1117_U270 , P1_R1117_U68 );
nand NAND2_9629 ( P1_R1117_U272 , P1_R1117_U271 , P1_R1117_U167 );
nand NAND2_9630 ( P1_R1117_U273 , P1_U3080 , P1_R1117_U67 );
not NOT1_9631 ( P1_R1117_U274 , P1_R1117_U166 );
nand NAND2_9632 ( P1_R1117_U275 , P1_U3509 , P1_R1117_U70 );
nand NAND2_9633 ( P1_R1117_U276 , P1_R1117_U275 , P1_R1117_U166 );
nand NAND2_9634 ( P1_R1117_U277 , P1_U3079 , P1_R1117_U69 );
not NOT1_9635 ( P1_R1117_U278 , P1_R1117_U164 );
nand NAND2_9636 ( P1_R1117_U279 , P1_U4015 , P1_R1117_U72 );
nand NAND2_9637 ( P1_R1117_U280 , P1_R1117_U279 , P1_R1117_U164 );
nand NAND2_9638 ( P1_R1117_U281 , P1_U3074 , P1_R1117_U71 );
not NOT1_9639 ( P1_R1117_U282 , P1_R1117_U163 );
nand NAND2_9640 ( P1_R1117_U283 , P1_U4012 , P1_R1117_U75 );
nand NAND2_9641 ( P1_R1117_U284 , P1_U3064 , P1_R1117_U73 );
nand NAND2_9642 ( P1_R1117_U285 , P1_U3059 , P1_R1117_U48 );
nand NAND2_9643 ( P1_R1117_U286 , P1_R1117_U187 , P1_R1117_U181 );
nand NAND2_9644 ( P1_R1117_U287 , P1_R1117_U11 , P1_R1117_U286 );
nand NAND2_9645 ( P1_R1117_U288 , P1_U4014 , P1_R1117_U77 );
nand NAND2_9646 ( P1_R1117_U289 , P1_U4012 , P1_R1117_U75 );
nand NAND3_9647 ( P1_R1117_U290 , P1_R1117_U163 , P1_R1117_U127 , P1_R1117_U283 );
nand NAND2_9648 ( P1_R1117_U291 , P1_R1117_U289 , P1_R1117_U287 );
not NOT1_9649 ( P1_R1117_U292 , P1_R1117_U160 );
nand NAND2_9650 ( P1_R1117_U293 , P1_U4011 , P1_R1117_U80 );
nand NAND2_9651 ( P1_R1117_U294 , P1_R1117_U293 , P1_R1117_U160 );
nand NAND2_9652 ( P1_R1117_U295 , P1_U3063 , P1_R1117_U79 );
not NOT1_9653 ( P1_R1117_U296 , P1_R1117_U159 );
nand NAND2_9654 ( P1_R1117_U297 , P1_U4010 , P1_R1117_U82 );
nand NAND2_9655 ( P1_R1117_U298 , P1_R1117_U297 , P1_R1117_U159 );
nand NAND2_9656 ( P1_R1117_U299 , P1_U3056 , P1_R1117_U81 );
not NOT1_9657 ( P1_R1117_U300 , P1_R1117_U89 );
nand NAND2_9658 ( P1_R1117_U301 , P1_U4008 , P1_R1117_U86 );
nand NAND3_9659 ( P1_R1117_U302 , P1_R1117_U89 , P1_R1117_U182 , P1_R1117_U301 );
nand NAND2_9660 ( P1_R1117_U303 , P1_R1117_U86 , P1_R1117_U85 );
nand NAND2_9661 ( P1_R1117_U304 , P1_R1117_U303 , P1_R1117_U83 );
nand NAND2_9662 ( P1_R1117_U305 , P1_U3051 , P1_R1117_U176 );
not NOT1_9663 ( P1_R1117_U306 , P1_R1117_U157 );
nand NAND2_9664 ( P1_R1117_U307 , P1_U4007 , P1_R1117_U88 );
nand NAND2_9665 ( P1_R1117_U308 , P1_U3052 , P1_R1117_U87 );
nand NAND2_9666 ( P1_R1117_U309 , P1_R1117_U300 , P1_R1117_U85 );
nand NAND2_9667 ( P1_R1117_U310 , P1_R1117_U133 , P1_R1117_U309 );
nand NAND2_9668 ( P1_R1117_U311 , P1_R1117_U89 , P1_R1117_U182 );
nand NAND2_9669 ( P1_R1117_U312 , P1_R1117_U132 , P1_R1117_U311 );
nand NAND2_9670 ( P1_R1117_U313 , P1_R1117_U85 , P1_R1117_U182 );
nand NAND2_9671 ( P1_R1117_U314 , P1_R1117_U288 , P1_R1117_U163 );
not NOT1_9672 ( P1_R1117_U315 , P1_R1117_U90 );
nand NAND2_9673 ( P1_R1117_U316 , P1_U3059 , P1_R1117_U48 );
nand NAND2_9674 ( P1_R1117_U317 , P1_R1117_U315 , P1_R1117_U316 );
nand NAND2_9675 ( P1_R1117_U318 , P1_R1117_U136 , P1_R1117_U317 );
nand NAND2_9676 ( P1_R1117_U319 , P1_R1117_U90 , P1_R1117_U181 );
nand NAND2_9677 ( P1_R1117_U320 , P1_U4012 , P1_R1117_U75 );
nand NAND3_9678 ( P1_R1117_U321 , P1_R1117_U320 , P1_R1117_U319 , P1_R1117_U11 );
nand NAND2_9679 ( P1_R1117_U322 , P1_U3059 , P1_R1117_U48 );
nand NAND2_9680 ( P1_R1117_U323 , P1_R1117_U181 , P1_R1117_U322 );
nand NAND2_9681 ( P1_R1117_U324 , P1_R1117_U288 , P1_R1117_U78 );
nand NAND2_9682 ( P1_R1117_U325 , P1_R1117_U262 , P1_R1117_U171 );
not NOT1_9683 ( P1_R1117_U326 , P1_R1117_U91 );
nand NAND2_9684 ( P1_R1117_U327 , P1_U3072 , P1_R1117_U49 );
nand NAND2_9685 ( P1_R1117_U328 , P1_R1117_U326 , P1_R1117_U327 );
nand NAND2_9686 ( P1_R1117_U329 , P1_R1117_U142 , P1_R1117_U328 );
nand NAND2_9687 ( P1_R1117_U330 , P1_R1117_U91 , P1_R1117_U180 );
nand NAND2_9688 ( P1_R1117_U331 , P1_U3501 , P1_R1117_U61 );
nand NAND3_9689 ( P1_R1117_U332 , P1_R1117_U331 , P1_R1117_U330 , P1_R1117_U10 );
nand NAND2_9690 ( P1_R1117_U333 , P1_U3072 , P1_R1117_U49 );
nand NAND2_9691 ( P1_R1117_U334 , P1_R1117_U180 , P1_R1117_U333 );
nand NAND2_9692 ( P1_R1117_U335 , P1_R1117_U262 , P1_R1117_U64 );
nand NAND2_9693 ( P1_R1117_U336 , P1_R1117_U217 , P1_R1117_U148 );
not NOT1_9694 ( P1_R1117_U337 , P1_R1117_U92 );
nand NAND2_9695 ( P1_R1117_U338 , P1_U3060 , P1_R1117_U51 );
nand NAND2_9696 ( P1_R1117_U339 , P1_R1117_U337 , P1_R1117_U338 );
nand NAND2_9697 ( P1_R1117_U340 , P1_R1117_U146 , P1_R1117_U339 );
nand NAND2_9698 ( P1_R1117_U341 , P1_R1117_U92 , P1_R1117_U179 );
nand NAND2_9699 ( P1_R1117_U342 , P1_U3486 , P1_R1117_U52 );
nand NAND2_9700 ( P1_R1117_U343 , P1_R1117_U145 , P1_R1117_U341 );
nand NAND2_9701 ( P1_R1117_U344 , P1_U3060 , P1_R1117_U51 );
nand NAND2_9702 ( P1_R1117_U345 , P1_R1117_U179 , P1_R1117_U344 );
nand NAND2_9703 ( P1_R1117_U346 , P1_U3075 , P1_R1117_U24 );
nand NAND3_9704 ( P1_R1117_U347 , P1_R1117_U89 , P1_R1117_U182 , P1_R1117_U301 );
nand NAND3_9705 ( P1_R1117_U348 , P1_R1117_U12 , P1_R1117_U347 , P1_R1117_U130 );
nand NAND2_9706 ( P1_R1117_U349 , P1_U3480 , P1_R1117_U43 );
nand NAND2_9707 ( P1_R1117_U350 , P1_U3081 , P1_R1117_U42 );
nand NAND2_9708 ( P1_R1117_U351 , P1_R1117_U218 , P1_R1117_U148 );
nand NAND2_9709 ( P1_R1117_U352 , P1_R1117_U216 , P1_R1117_U147 );
nand NAND2_9710 ( P1_R1117_U353 , P1_U3477 , P1_R1117_U41 );
nand NAND2_9711 ( P1_R1117_U354 , P1_U3082 , P1_R1117_U38 );
nand NAND2_9712 ( P1_R1117_U355 , P1_U3477 , P1_R1117_U41 );
nand NAND2_9713 ( P1_R1117_U356 , P1_U3082 , P1_R1117_U38 );
nand NAND2_9714 ( P1_R1117_U357 , P1_R1117_U356 , P1_R1117_U355 );
nand NAND2_9715 ( P1_R1117_U358 , P1_U3474 , P1_R1117_U39 );
nand NAND2_9716 ( P1_R1117_U359 , P1_U3068 , P1_R1117_U22 );
nand NAND2_9717 ( P1_R1117_U360 , P1_R1117_U223 , P1_R1117_U44 );
nand NAND2_9718 ( P1_R1117_U361 , P1_R1117_U149 , P1_R1117_U210 );
nand NAND2_9719 ( P1_R1117_U362 , P1_U3471 , P1_R1117_U34 );
nand NAND2_9720 ( P1_R1117_U363 , P1_U3069 , P1_R1117_U31 );
nand NAND2_9721 ( P1_R1117_U364 , P1_R1117_U363 , P1_R1117_U362 );
nand NAND2_9722 ( P1_R1117_U365 , P1_U3468 , P1_R1117_U35 );
nand NAND2_9723 ( P1_R1117_U366 , P1_U3065 , P1_R1117_U32 );
nand NAND2_9724 ( P1_R1117_U367 , P1_R1117_U233 , P1_R1117_U45 );
nand NAND2_9725 ( P1_R1117_U368 , P1_R1117_U150 , P1_R1117_U225 );
nand NAND2_9726 ( P1_R1117_U369 , P1_U3465 , P1_R1117_U36 );
nand NAND2_9727 ( P1_R1117_U370 , P1_U3058 , P1_R1117_U33 );
nand NAND2_9728 ( P1_R1117_U371 , P1_R1117_U234 , P1_R1117_U152 );
nand NAND2_9729 ( P1_R1117_U372 , P1_R1117_U200 , P1_R1117_U151 );
nand NAND2_9730 ( P1_R1117_U373 , P1_U3462 , P1_R1117_U30 );
nand NAND2_9731 ( P1_R1117_U374 , P1_U3062 , P1_R1117_U27 );
nand NAND2_9732 ( P1_R1117_U375 , P1_U3462 , P1_R1117_U30 );
nand NAND2_9733 ( P1_R1117_U376 , P1_U3062 , P1_R1117_U27 );
nand NAND2_9734 ( P1_R1117_U377 , P1_R1117_U376 , P1_R1117_U375 );
nand NAND2_9735 ( P1_R1117_U378 , P1_U3459 , P1_R1117_U28 );
nand NAND2_9736 ( P1_R1117_U379 , P1_U3066 , P1_R1117_U23 );
nand NAND2_9737 ( P1_R1117_U380 , P1_R1117_U239 , P1_R1117_U46 );
nand NAND2_9738 ( P1_R1117_U381 , P1_R1117_U153 , P1_R1117_U194 );
nand NAND2_9739 ( P1_R1117_U382 , P1_U4018 , P1_R1117_U155 );
nand NAND2_9740 ( P1_R1117_U383 , P1_U3053 , P1_R1117_U154 );
nand NAND2_9741 ( P1_R1117_U384 , P1_U4018 , P1_R1117_U155 );
nand NAND2_9742 ( P1_R1117_U385 , P1_U3053 , P1_R1117_U154 );
nand NAND2_9743 ( P1_R1117_U386 , P1_R1117_U385 , P1_R1117_U384 );
nand NAND3_9744 ( P1_R1117_U387 , P1_U3052 , P1_R1117_U386 , P1_R1117_U87 );
nand NAND3_9745 ( P1_R1117_U388 , P1_R1117_U12 , P1_R1117_U88 , P1_U4007 );
nand NAND2_9746 ( P1_R1117_U389 , P1_U4007 , P1_R1117_U88 );
nand NAND2_9747 ( P1_R1117_U390 , P1_U3052 , P1_R1117_U87 );
not NOT1_9748 ( P1_R1117_U391 , P1_R1117_U131 );
nand NAND2_9749 ( P1_R1117_U392 , P1_R1117_U306 , P1_R1117_U391 );
nand NAND2_9750 ( P1_R1117_U393 , P1_R1117_U131 , P1_R1117_U157 );
nand NAND2_9751 ( P1_R1117_U394 , P1_U4008 , P1_R1117_U86 );
nand NAND2_9752 ( P1_R1117_U395 , P1_U3051 , P1_R1117_U83 );
nand NAND2_9753 ( P1_R1117_U396 , P1_U4008 , P1_R1117_U86 );
nand NAND2_9754 ( P1_R1117_U397 , P1_U3051 , P1_R1117_U83 );
nand NAND2_9755 ( P1_R1117_U398 , P1_R1117_U397 , P1_R1117_U396 );
nand NAND2_9756 ( P1_R1117_U399 , P1_U4009 , P1_R1117_U84 );
nand NAND2_9757 ( P1_R1117_U400 , P1_U3055 , P1_R1117_U47 );
nand NAND2_9758 ( P1_R1117_U401 , P1_R1117_U313 , P1_R1117_U89 );
nand NAND2_9759 ( P1_R1117_U402 , P1_R1117_U158 , P1_R1117_U300 );
nand NAND2_9760 ( P1_R1117_U403 , P1_U4010 , P1_R1117_U82 );
nand NAND2_9761 ( P1_R1117_U404 , P1_U3056 , P1_R1117_U81 );
not NOT1_9762 ( P1_R1117_U405 , P1_R1117_U134 );
nand NAND2_9763 ( P1_R1117_U406 , P1_R1117_U296 , P1_R1117_U405 );
nand NAND2_9764 ( P1_R1117_U407 , P1_R1117_U134 , P1_R1117_U159 );
nand NAND2_9765 ( P1_R1117_U408 , P1_U4011 , P1_R1117_U80 );
nand NAND2_9766 ( P1_R1117_U409 , P1_U3063 , P1_R1117_U79 );
not NOT1_9767 ( P1_R1117_U410 , P1_R1117_U135 );
nand NAND2_9768 ( P1_R1117_U411 , P1_R1117_U292 , P1_R1117_U410 );
nand NAND2_9769 ( P1_R1117_U412 , P1_R1117_U135 , P1_R1117_U160 );
nand NAND2_9770 ( P1_R1117_U413 , P1_U4012 , P1_R1117_U75 );
nand NAND2_9771 ( P1_R1117_U414 , P1_U3064 , P1_R1117_U73 );
nand NAND2_9772 ( P1_R1117_U415 , P1_R1117_U414 , P1_R1117_U413 );
nand NAND2_9773 ( P1_R1117_U416 , P1_U4013 , P1_R1117_U76 );
nand NAND2_9774 ( P1_R1117_U417 , P1_U3059 , P1_R1117_U48 );
nand NAND2_9775 ( P1_R1117_U418 , P1_R1117_U323 , P1_R1117_U90 );
nand NAND2_9776 ( P1_R1117_U419 , P1_R1117_U161 , P1_R1117_U315 );
nand NAND2_9777 ( P1_R1117_U420 , P1_U4014 , P1_R1117_U77 );
nand NAND2_9778 ( P1_R1117_U421 , P1_U3073 , P1_R1117_U74 );
nand NAND2_9779 ( P1_R1117_U422 , P1_R1117_U324 , P1_R1117_U163 );
nand NAND2_9780 ( P1_R1117_U423 , P1_R1117_U282 , P1_R1117_U162 );
nand NAND2_9781 ( P1_R1117_U424 , P1_U4015 , P1_R1117_U72 );
nand NAND2_9782 ( P1_R1117_U425 , P1_U3074 , P1_R1117_U71 );
not NOT1_9783 ( P1_R1117_U426 , P1_R1117_U137 );
nand NAND2_9784 ( P1_R1117_U427 , P1_R1117_U278 , P1_R1117_U426 );
nand NAND2_9785 ( P1_R1117_U428 , P1_R1117_U137 , P1_R1117_U164 );
nand NAND2_9786 ( P1_R1117_U429 , P1_U3456 , P1_R1117_U26 );
nand NAND2_9787 ( P1_R1117_U430 , P1_U3076 , P1_R1117_U165 );
not NOT1_9788 ( P1_R1117_U431 , P1_R1117_U138 );
nand NAND2_9789 ( P1_R1117_U432 , P1_R1117_U431 , P1_R1117_U190 );
nand NAND2_9790 ( P1_R1117_U433 , P1_R1117_U138 , P1_R1117_U25 );
nand NAND2_9791 ( P1_R1117_U434 , P1_U3509 , P1_R1117_U70 );
nand NAND2_9792 ( P1_R1117_U435 , P1_U3079 , P1_R1117_U69 );
not NOT1_9793 ( P1_R1117_U436 , P1_R1117_U139 );
nand NAND2_9794 ( P1_R1117_U437 , P1_R1117_U274 , P1_R1117_U436 );
nand NAND2_9795 ( P1_R1117_U438 , P1_R1117_U139 , P1_R1117_U166 );
nand NAND2_9796 ( P1_R1117_U439 , P1_U3507 , P1_R1117_U68 );
nand NAND2_9797 ( P1_R1117_U440 , P1_U3080 , P1_R1117_U167 );
not NOT1_9798 ( P1_R1117_U441 , P1_R1117_U140 );
nand NAND2_9799 ( P1_R1117_U442 , P1_R1117_U441 , P1_R1117_U270 );
nand NAND2_9800 ( P1_R1117_U443 , P1_R1117_U140 , P1_R1117_U67 );
nand NAND2_9801 ( P1_R1117_U444 , P1_U3504 , P1_R1117_U66 );
nand NAND2_9802 ( P1_R1117_U445 , P1_U3067 , P1_R1117_U65 );
not NOT1_9803 ( P1_R1117_U446 , P1_R1117_U141 );
nand NAND2_9804 ( P1_R1117_U447 , P1_R1117_U266 , P1_R1117_U446 );
nand NAND2_9805 ( P1_R1117_U448 , P1_R1117_U141 , P1_R1117_U168 );
nand NAND2_9806 ( P1_R1117_U449 , P1_U3501 , P1_R1117_U61 );
nand NAND2_9807 ( P1_R1117_U450 , P1_U3071 , P1_R1117_U59 );
nand NAND2_9808 ( P1_R1117_U451 , P1_R1117_U450 , P1_R1117_U449 );
nand NAND2_9809 ( P1_R1117_U452 , P1_U3498 , P1_R1117_U62 );
nand NAND2_9810 ( P1_R1117_U453 , P1_U3072 , P1_R1117_U49 );
nand NAND2_9811 ( P1_R1117_U454 , P1_R1117_U334 , P1_R1117_U91 );
nand NAND2_9812 ( P1_R1117_U455 , P1_R1117_U169 , P1_R1117_U326 );
nand NAND2_9813 ( P1_R1117_U456 , P1_U3495 , P1_R1117_U63 );
nand NAND2_9814 ( P1_R1117_U457 , P1_U3077 , P1_R1117_U60 );
nand NAND2_9815 ( P1_R1117_U458 , P1_R1117_U335 , P1_R1117_U171 );
nand NAND2_9816 ( P1_R1117_U459 , P1_R1117_U256 , P1_R1117_U170 );
nand NAND2_9817 ( P1_R1117_U460 , P1_U3492 , P1_R1117_U58 );
nand NAND2_9818 ( P1_R1117_U461 , P1_U3078 , P1_R1117_U57 );
not NOT1_9819 ( P1_R1117_U462 , P1_R1117_U143 );
nand NAND2_9820 ( P1_R1117_U463 , P1_R1117_U252 , P1_R1117_U462 );
nand NAND2_9821 ( P1_R1117_U464 , P1_R1117_U143 , P1_R1117_U172 );
nand NAND2_9822 ( P1_R1117_U465 , P1_U3489 , P1_R1117_U56 );
nand NAND2_9823 ( P1_R1117_U466 , P1_U3070 , P1_R1117_U55 );
not NOT1_9824 ( P1_R1117_U467 , P1_R1117_U144 );
nand NAND2_9825 ( P1_R1117_U468 , P1_R1117_U248 , P1_R1117_U467 );
nand NAND2_9826 ( P1_R1117_U469 , P1_R1117_U144 , P1_R1117_U173 );
nand NAND2_9827 ( P1_R1117_U470 , P1_U3486 , P1_R1117_U52 );
nand NAND2_9828 ( P1_R1117_U471 , P1_U3061 , P1_R1117_U50 );
nand NAND2_9829 ( P1_R1117_U472 , P1_R1117_U471 , P1_R1117_U470 );
nand NAND2_9830 ( P1_R1117_U473 , P1_U3483 , P1_R1117_U53 );
nand NAND2_9831 ( P1_R1117_U474 , P1_U3060 , P1_R1117_U51 );
nand NAND2_9832 ( P1_R1117_U475 , P1_R1117_U345 , P1_R1117_U92 );
nand NAND2_9833 ( P1_R1117_U476 , P1_R1117_U174 , P1_R1117_U337 );
and AND2_9834 ( P1_R1375_U6 , P1_R1375_U119 , P1_R1375_U120 );
and AND2_9835 ( P1_R1375_U7 , P1_R1375_U137 , P1_R1375_U136 );
and AND4_9836 ( P1_R1375_U8 , P1_R1375_U144 , P1_R1375_U143 , P1_R1375_U142 , P1_R1375_U141 );
and AND2_9837 ( P1_R1375_U9 , P1_R1375_U164 , P1_R1375_U163 );
and AND4_9838 ( P1_R1375_U10 , P1_R1375_U197 , P1_R1375_U196 , P1_R1375_U198 , P1_R1375_U6 );
and AND2_9839 ( P1_R1375_U11 , P1_U4018 , P1_R1375_U20 );
and AND4_9840 ( P1_R1375_U12 , P1_R1375_U207 , P1_R1375_U206 , P1_R1375_U118 , P1_R1375_U117 );
and AND2_9841 ( P1_R1375_U13 , P1_U3451 , P1_R1375_U48 );
and AND3_9842 ( P1_R1375_U14 , P1_R1375_U205 , P1_R1375_U115 , P1_R1375_U204 );
not NOT1_9843 ( P1_R1375_U15 , P1_U4016 );
not NOT1_9844 ( P1_R1375_U16 , P1_U4017 );
not NOT1_9845 ( P1_R1375_U17 , P1_U3054 );
not NOT1_9846 ( P1_R1375_U18 , P1_U4018 );
not NOT1_9847 ( P1_R1375_U19 , P1_U3057 );
not NOT1_9848 ( P1_R1375_U20 , P1_U3053 );
not NOT1_9849 ( P1_R1375_U21 , P1_U3052 );
not NOT1_9850 ( P1_R1375_U22 , P1_U4008 );
not NOT1_9851 ( P1_R1375_U23 , P1_U3055 );
not NOT1_9852 ( P1_R1375_U24 , P1_U4010 );
not NOT1_9853 ( P1_R1375_U25 , P1_U4007 );
not NOT1_9854 ( P1_R1375_U26 , P1_U4009 );
not NOT1_9855 ( P1_R1375_U27 , P1_U4011 );
not NOT1_9856 ( P1_R1375_U28 , P1_U3064 );
not NOT1_9857 ( P1_R1375_U29 , P1_U4012 );
not NOT1_9858 ( P1_R1375_U30 , P1_U3059 );
not NOT1_9859 ( P1_R1375_U31 , P1_U3056 );
not NOT1_9860 ( P1_R1375_U32 , P1_U3063 );
not NOT1_9861 ( P1_R1375_U33 , P1_U3073 );
not NOT1_9862 ( P1_R1375_U34 , P1_U3074 );
not NOT1_9863 ( P1_R1375_U35 , P1_U3504 );
not NOT1_9864 ( P1_R1375_U36 , P1_U3507 );
not NOT1_9865 ( P1_R1375_U37 , P1_U3072 );
not NOT1_9866 ( P1_R1375_U38 , P1_U3077 );
not NOT1_9867 ( P1_R1375_U39 , P1_U3471 );
not NOT1_9868 ( P1_R1375_U40 , P1_U3065 );
not NOT1_9869 ( P1_R1375_U41 , P1_U3081 );
not NOT1_9870 ( P1_R1375_U42 , P1_U3082 );
not NOT1_9871 ( P1_R1375_U43 , P1_U3069 );
not NOT1_9872 ( P1_R1375_U44 , P1_U3068 );
not NOT1_9873 ( P1_R1375_U45 , P1_U3058 );
not NOT1_9874 ( P1_R1375_U46 , P1_U3062 );
not NOT1_9875 ( P1_R1375_U47 , P1_U3451 );
not NOT1_9876 ( P1_R1375_U48 , P1_U3075 );
nand NAND2_9877 ( P1_R1375_U49 , P1_R1375_U147 , P1_R1375_U146 );
not NOT1_9878 ( P1_R1375_U50 , P1_U3456 );
not NOT1_9879 ( P1_R1375_U51 , P1_U3066 );
not NOT1_9880 ( P1_R1375_U52 , P1_U3486 );
not NOT1_9881 ( P1_R1375_U53 , P1_U3489 );
not NOT1_9882 ( P1_R1375_U54 , P1_U3459 );
not NOT1_9883 ( P1_R1375_U55 , P1_U3462 );
not NOT1_9884 ( P1_R1375_U56 , P1_U3468 );
not NOT1_9885 ( P1_R1375_U57 , P1_U3465 );
not NOT1_9886 ( P1_R1375_U58 , P1_U3474 );
not NOT1_9887 ( P1_R1375_U59 , P1_U3477 );
not NOT1_9888 ( P1_R1375_U60 , P1_U3480 );
not NOT1_9889 ( P1_R1375_U61 , P1_U3483 );
not NOT1_9890 ( P1_R1375_U62 , P1_U3060 );
not NOT1_9891 ( P1_R1375_U63 , P1_U3070 );
not NOT1_9892 ( P1_R1375_U64 , P1_U3061 );
not NOT1_9893 ( P1_R1375_U65 , P1_U3078 );
not NOT1_9894 ( P1_R1375_U66 , P1_U3492 );
not NOT1_9895 ( P1_R1375_U67 , P1_U3495 );
not NOT1_9896 ( P1_R1375_U68 , P1_U3498 );
not NOT1_9897 ( P1_R1375_U69 , P1_U3501 );
not NOT1_9898 ( P1_R1375_U70 , P1_U3071 );
not NOT1_9899 ( P1_R1375_U71 , P1_U3067 );
not NOT1_9900 ( P1_R1375_U72 , P1_U3080 );
not NOT1_9901 ( P1_R1375_U73 , P1_U3079 );
not NOT1_9902 ( P1_R1375_U74 , P1_U3509 );
not NOT1_9903 ( P1_R1375_U75 , P1_U4015 );
not NOT1_9904 ( P1_R1375_U76 , P1_U4014 );
not NOT1_9905 ( P1_R1375_U77 , P1_U4013 );
nand NAND2_9906 ( P1_R1375_U78 , P1_R1375_U11 , P1_R1375_U125 );
nand NAND4_9907 ( P1_R1375_U79 , P1_R1375_U124 , P1_R1375_U122 , P1_R1375_U87 , P1_R1375_U12 );
nand NAND2_9908 ( P1_R1375_U80 , P1_R1375_U109 , P1_R1375_U195 );
and AND2_9909 ( P1_R1375_U81 , P1_U4008 , P1_R1375_U113 );
and AND2_9910 ( P1_R1375_U82 , P1_U4010 , P1_R1375_U31 );
and AND2_9911 ( P1_R1375_U83 , P1_U4007 , P1_R1375_U21 );
and AND2_9912 ( P1_R1375_U84 , P1_U4009 , P1_R1375_U23 );
and AND2_9913 ( P1_R1375_U85 , P1_U3064 , P1_R1375_U29 );
and AND2_9914 ( P1_R1375_U86 , P1_U3059 , P1_R1375_U77 );
and AND2_9915 ( P1_R1375_U87 , P1_R1375_U123 , P1_R1375_U121 );
and AND2_9916 ( P1_R1375_U88 , P1_R1375_U129 , P1_R1375_U126 );
and AND3_9917 ( P1_R1375_U89 , P1_R1375_U131 , P1_R1375_U201 , P1_R1375_U128 );
and AND2_9918 ( P1_R1375_U90 , P1_U3065 , P1_R1375_U56 );
and AND2_9919 ( P1_R1375_U91 , P1_R1375_U145 , P1_R1375_U149 );
and AND2_9920 ( P1_R1375_U92 , P1_R1375_U91 , P1_R1375_U140 );
and AND3_9921 ( P1_R1375_U93 , P1_R1375_U153 , P1_R1375_U152 , P1_R1375_U8 );
and AND2_9922 ( P1_R1375_U94 , P1_U3459 , P1_R1375_U51 );
and AND3_9923 ( P1_R1375_U95 , P1_R1375_U161 , P1_R1375_U160 , P1_R1375_U159 );
and AND2_9924 ( P1_R1375_U96 , P1_U3474 , P1_R1375_U44 );
and AND2_9925 ( P1_R1375_U97 , P1_R1375_U171 , P1_R1375_U170 );
and AND2_9926 ( P1_R1375_U98 , P1_R1375_U97 , P1_R1375_U9 );
and AND2_9927 ( P1_R1375_U99 , P1_U3060 , P1_R1375_U61 );
and AND2_9928 ( P1_R1375_U100 , P1_U3061 , P1_R1375_U52 );
and AND3_9929 ( P1_R1375_U101 , P1_R1375_U173 , P1_R1375_U174 , P1_R1375_U102 );
and AND2_9930 ( P1_R1375_U102 , P1_R1375_U177 , P1_R1375_U176 );
and AND2_9931 ( P1_R1375_U103 , P1_R1375_U7 , P1_R1375_U104 );
and AND2_9932 ( P1_R1375_U104 , P1_R1375_U185 , P1_R1375_U186 );
and AND2_9933 ( P1_R1375_U105 , P1_U3071 , P1_R1375_U69 );
and AND2_9934 ( P1_R1375_U106 , P1_U3067 , P1_R1375_U35 );
and AND3_9935 ( P1_R1375_U107 , P1_R1375_U188 , P1_R1375_U190 , P1_R1375_U108 );
and AND2_9936 ( P1_R1375_U108 , P1_R1375_U192 , P1_R1375_U191 );
and AND2_9937 ( P1_R1375_U109 , P1_R1375_U134 , P1_R1375_U133 );
and AND2_9938 ( P1_R1375_U110 , P1_U4015 , P1_R1375_U34 );
and AND2_9939 ( P1_R1375_U111 , P1_R1375_U128 , P1_R1375_U127 );
and AND4_9940 ( P1_R1375_U112 , P1_R1375_U10 , P1_R1375_U131 , P1_R1375_U129 , P1_R1375_U130 );
not NOT1_9941 ( P1_R1375_U113 , P1_U3051 );
nand NAND2_9942 ( P1_R1375_U114 , P1_R1375_U200 , P1_R1375_U199 );
nand NAND2_9943 ( P1_R1375_U115 , P1_U4016 , P1_R1375_U17 );
nand NAND2_9944 ( P1_R1375_U116 , P1_U3053 , P1_R1375_U18 );
nand NAND2_9945 ( P1_R1375_U117 , P1_U3052 , P1_R1375_U25 );
nand NAND2_9946 ( P1_R1375_U118 , P1_U3055 , P1_R1375_U26 );
nand NAND2_9947 ( P1_R1375_U119 , P1_U4011 , P1_R1375_U32 );
nand NAND2_9948 ( P1_R1375_U120 , P1_U4012 , P1_R1375_U28 );
nand NAND2_9949 ( P1_R1375_U121 , P1_R1375_U85 , P1_R1375_U119 );
nand NAND2_9950 ( P1_R1375_U122 , P1_R1375_U86 , P1_R1375_U6 );
nand NAND2_9951 ( P1_R1375_U123 , P1_U3056 , P1_R1375_U24 );
nand NAND2_9952 ( P1_R1375_U124 , P1_U3063 , P1_R1375_U27 );
nand NAND2_9953 ( P1_R1375_U125 , P1_U3057 , P1_R1375_U16 );
nand NAND3_9954 ( P1_R1375_U126 , P1_R1375_U81 , P1_R1375_U117 , P1_R1375_U115 );
nand NAND3_9955 ( P1_R1375_U127 , P1_R1375_U82 , P1_R1375_U12 , P1_R1375_U115 );
nand NAND3_9956 ( P1_R1375_U128 , P1_R1375_U115 , P1_R1375_U19 , P1_U4017 );
nand NAND2_9957 ( P1_R1375_U129 , P1_R1375_U83 , P1_R1375_U115 );
nand NAND3_9958 ( P1_R1375_U130 , P1_R1375_U84 , P1_R1375_U12 , P1_R1375_U115 );
nand NAND2_9959 ( P1_R1375_U131 , P1_U3054 , P1_R1375_U15 );
nand NAND4_9960 ( P1_R1375_U132 , P1_R1375_U79 , P1_R1375_U130 , P1_R1375_U88 , P1_R1375_U127 );
nand NAND2_9961 ( P1_R1375_U133 , P1_U3073 , P1_R1375_U76 );
nand NAND2_9962 ( P1_R1375_U134 , P1_U3074 , P1_R1375_U75 );
nand NAND2_9963 ( P1_R1375_U135 , P1_U3072 , P1_R1375_U68 );
nand NAND2_9964 ( P1_R1375_U136 , P1_U3504 , P1_R1375_U71 );
nand NAND2_9965 ( P1_R1375_U137 , P1_U3507 , P1_R1375_U72 );
nand NAND2_9966 ( P1_R1375_U138 , P1_U3077 , P1_R1375_U67 );
nand NAND2_9967 ( P1_R1375_U139 , P1_U3471 , P1_R1375_U43 );
nand NAND2_9968 ( P1_R1375_U140 , P1_R1375_U90 , P1_R1375_U139 );
nand NAND2_9969 ( P1_R1375_U141 , P1_U3081 , P1_R1375_U60 );
nand NAND2_9970 ( P1_R1375_U142 , P1_U3082 , P1_R1375_U59 );
nand NAND2_9971 ( P1_R1375_U143 , P1_U3069 , P1_R1375_U39 );
nand NAND2_9972 ( P1_R1375_U144 , P1_U3068 , P1_R1375_U58 );
nand NAND2_9973 ( P1_R1375_U145 , P1_U3058 , P1_R1375_U57 );
or OR2_9974 ( P1_R1375_U146 , P1_U3448 , P1_R1375_U13 );
nand NAND2_9975 ( P1_R1375_U147 , P1_U3075 , P1_R1375_U47 );
not NOT1_9976 ( P1_R1375_U148 , P1_R1375_U49 );
nand NAND2_9977 ( P1_R1375_U149 , P1_U3062 , P1_R1375_U55 );
nand NAND2_9978 ( P1_R1375_U150 , P1_U3456 , P1_R1375_U148 );
nand NAND2_9979 ( P1_R1375_U151 , P1_U3076 , P1_R1375_U150 );
nand NAND2_9980 ( P1_R1375_U152 , P1_R1375_U49 , P1_R1375_U50 );
nand NAND2_9981 ( P1_R1375_U153 , P1_U3066 , P1_R1375_U54 );
nand NAND3_9982 ( P1_R1375_U154 , P1_R1375_U92 , P1_R1375_U151 , P1_R1375_U93 );
nand NAND2_9983 ( P1_R1375_U155 , P1_R1375_U94 , P1_R1375_U149 );
nand NAND2_9984 ( P1_R1375_U156 , P1_U3462 , P1_R1375_U46 );
nand NAND2_9985 ( P1_R1375_U157 , P1_R1375_U156 , P1_R1375_U155 );
nand NAND2_9986 ( P1_R1375_U158 , P1_R1375_U157 , P1_R1375_U145 );
nand NAND2_9987 ( P1_R1375_U159 , P1_U3468 , P1_R1375_U40 );
nand NAND2_9988 ( P1_R1375_U160 , P1_U3465 , P1_R1375_U45 );
nand NAND2_9989 ( P1_R1375_U161 , P1_U3471 , P1_R1375_U43 );
nand NAND2_9990 ( P1_R1375_U162 , P1_R1375_U158 , P1_R1375_U95 );
nand NAND2_9991 ( P1_R1375_U163 , P1_U3486 , P1_R1375_U64 );
nand NAND2_9992 ( P1_R1375_U164 , P1_U3489 , P1_R1375_U63 );
nand NAND2_9993 ( P1_R1375_U165 , P1_R1375_U96 , P1_R1375_U142 );
nand NAND2_9994 ( P1_R1375_U166 , P1_U3477 , P1_R1375_U42 );
nand NAND2_9995 ( P1_R1375_U167 , P1_R1375_U166 , P1_R1375_U165 );
nand NAND3_9996 ( P1_R1375_U168 , P1_R1375_U162 , P1_R1375_U140 , P1_R1375_U8 );
nand NAND2_9997 ( P1_R1375_U169 , P1_R1375_U167 , P1_R1375_U141 );
nand NAND2_9998 ( P1_R1375_U170 , P1_U3480 , P1_R1375_U41 );
nand NAND2_9999 ( P1_R1375_U171 , P1_U3483 , P1_R1375_U62 );
nand NAND4_10000 ( P1_R1375_U172 , P1_R1375_U168 , P1_R1375_U169 , P1_R1375_U98 , P1_R1375_U154 );
nand NAND2_10001 ( P1_R1375_U173 , P1_R1375_U99 , P1_R1375_U9 );
nand NAND2_10002 ( P1_R1375_U174 , P1_U3070 , P1_R1375_U53 );
nand NAND2_10003 ( P1_R1375_U175 , P1_U3489 , P1_R1375_U63 );
nand NAND2_10004 ( P1_R1375_U176 , P1_R1375_U100 , P1_R1375_U175 );
nand NAND2_10005 ( P1_R1375_U177 , P1_U3078 , P1_R1375_U66 );
nand NAND2_10006 ( P1_R1375_U178 , P1_R1375_U172 , P1_R1375_U101 );
nand NAND2_10007 ( P1_R1375_U179 , P1_U3492 , P1_R1375_U65 );
nand NAND2_10008 ( P1_R1375_U180 , P1_R1375_U179 , P1_R1375_U178 );
nand NAND2_10009 ( P1_R1375_U181 , P1_R1375_U180 , P1_R1375_U138 );
nand NAND2_10010 ( P1_R1375_U182 , P1_U3495 , P1_R1375_U38 );
nand NAND2_10011 ( P1_R1375_U183 , P1_R1375_U182 , P1_R1375_U181 );
nand NAND2_10012 ( P1_R1375_U184 , P1_R1375_U183 , P1_R1375_U135 );
nand NAND2_10013 ( P1_R1375_U185 , P1_U3498 , P1_R1375_U37 );
nand NAND2_10014 ( P1_R1375_U186 , P1_U3501 , P1_R1375_U70 );
nand NAND2_10015 ( P1_R1375_U187 , P1_R1375_U184 , P1_R1375_U103 );
nand NAND2_10016 ( P1_R1375_U188 , P1_R1375_U105 , P1_R1375_U7 );
nand NAND2_10017 ( P1_R1375_U189 , P1_U3507 , P1_R1375_U72 );
nand NAND2_10018 ( P1_R1375_U190 , P1_R1375_U106 , P1_R1375_U189 );
nand NAND2_10019 ( P1_R1375_U191 , P1_U3080 , P1_R1375_U36 );
nand NAND2_10020 ( P1_R1375_U192 , P1_U3079 , P1_R1375_U74 );
nand NAND2_10021 ( P1_R1375_U193 , P1_R1375_U187 , P1_R1375_U107 );
nand NAND2_10022 ( P1_R1375_U194 , P1_U3509 , P1_R1375_U73 );
nand NAND2_10023 ( P1_R1375_U195 , P1_R1375_U194 , P1_R1375_U193 );
nand NAND2_10024 ( P1_R1375_U196 , P1_R1375_U110 , P1_R1375_U133 );
nand NAND2_10025 ( P1_R1375_U197 , P1_U4014 , P1_R1375_U33 );
nand NAND2_10026 ( P1_R1375_U198 , P1_U4013 , P1_R1375_U30 );
nand NAND2_10027 ( P1_R1375_U199 , P1_U4017 , P1_R1375_U116 );
nand NAND2_10028 ( P1_R1375_U200 , P1_R1375_U19 , P1_R1375_U116 );
nand NAND2_10029 ( P1_R1375_U201 , P1_R1375_U11 , P1_R1375_U202 );
nand NAND2_10030 ( P1_R1375_U202 , P1_U3057 , P1_R1375_U16 );
nand NAND2_10031 ( P1_R1375_U203 , P1_R1375_U132 , P1_R1375_U114 );
nand NAND2_10032 ( P1_R1375_U204 , P1_R1375_U89 , P1_R1375_U203 );
nand NAND5_10033 ( P1_R1375_U205 , P1_R1375_U126 , P1_R1375_U80 , P1_R1375_U78 , P1_R1375_U111 , P1_R1375_U112 );
nand NAND2_10034 ( P1_R1375_U206 , P1_U3051 , P1_R1375_U22 );
nand NAND2_10035 ( P1_R1375_U207 , P1_U4008 , P1_R1375_U113 );
and AND2_10036 ( P1_R1352_U6 , P1_U3057 , P1_R1352_U7 );
not NOT1_10037 ( P1_R1352_U7 , P1_U3054 );
and AND2_10038 ( P1_R1207_U6 , P1_R1207_U184 , P1_R1207_U201 );
and AND2_10039 ( P1_R1207_U7 , P1_R1207_U203 , P1_R1207_U202 );
and AND2_10040 ( P1_R1207_U8 , P1_R1207_U179 , P1_R1207_U240 );
and AND2_10041 ( P1_R1207_U9 , P1_R1207_U242 , P1_R1207_U241 );
and AND2_10042 ( P1_R1207_U10 , P1_R1207_U259 , P1_R1207_U258 );
and AND2_10043 ( P1_R1207_U11 , P1_R1207_U285 , P1_R1207_U284 );
and AND2_10044 ( P1_R1207_U12 , P1_R1207_U383 , P1_R1207_U382 );
nand NAND2_10045 ( P1_R1207_U13 , P1_R1207_U340 , P1_R1207_U343 );
nand NAND2_10046 ( P1_R1207_U14 , P1_R1207_U329 , P1_R1207_U332 );
nand NAND2_10047 ( P1_R1207_U15 , P1_R1207_U318 , P1_R1207_U321 );
nand NAND2_10048 ( P1_R1207_U16 , P1_R1207_U310 , P1_R1207_U312 );
nand NAND3_10049 ( P1_R1207_U17 , P1_R1207_U156 , P1_R1207_U175 , P1_R1207_U348 );
nand NAND2_10050 ( P1_R1207_U18 , P1_R1207_U236 , P1_R1207_U238 );
nand NAND2_10051 ( P1_R1207_U19 , P1_R1207_U228 , P1_R1207_U231 );
nand NAND2_10052 ( P1_R1207_U20 , P1_R1207_U220 , P1_R1207_U222 );
nand NAND2_10053 ( P1_R1207_U21 , P1_R1207_U25 , P1_R1207_U346 );
not NOT1_10054 ( P1_R1207_U22 , P1_U3474 );
not NOT1_10055 ( P1_R1207_U23 , P1_U3459 );
not NOT1_10056 ( P1_R1207_U24 , P1_U3451 );
nand NAND2_10057 ( P1_R1207_U25 , P1_U3451 , P1_R1207_U93 );
not NOT1_10058 ( P1_R1207_U26 , P1_U3076 );
not NOT1_10059 ( P1_R1207_U27 , P1_U3462 );
not NOT1_10060 ( P1_R1207_U28 , P1_U3066 );
nand NAND2_10061 ( P1_R1207_U29 , P1_U3066 , P1_R1207_U23 );
not NOT1_10062 ( P1_R1207_U30 , P1_U3062 );
not NOT1_10063 ( P1_R1207_U31 , P1_U3471 );
not NOT1_10064 ( P1_R1207_U32 , P1_U3468 );
not NOT1_10065 ( P1_R1207_U33 , P1_U3465 );
not NOT1_10066 ( P1_R1207_U34 , P1_U3069 );
not NOT1_10067 ( P1_R1207_U35 , P1_U3065 );
not NOT1_10068 ( P1_R1207_U36 , P1_U3058 );
nand NAND2_10069 ( P1_R1207_U37 , P1_U3058 , P1_R1207_U33 );
not NOT1_10070 ( P1_R1207_U38 , P1_U3477 );
not NOT1_10071 ( P1_R1207_U39 , P1_U3068 );
nand NAND2_10072 ( P1_R1207_U40 , P1_U3068 , P1_R1207_U22 );
not NOT1_10073 ( P1_R1207_U41 , P1_U3082 );
not NOT1_10074 ( P1_R1207_U42 , P1_U3480 );
not NOT1_10075 ( P1_R1207_U43 , P1_U3081 );
nand NAND2_10076 ( P1_R1207_U44 , P1_R1207_U209 , P1_R1207_U208 );
nand NAND2_10077 ( P1_R1207_U45 , P1_R1207_U37 , P1_R1207_U224 );
nand NAND2_10078 ( P1_R1207_U46 , P1_R1207_U193 , P1_R1207_U192 );
not NOT1_10079 ( P1_R1207_U47 , P1_U4009 );
not NOT1_10080 ( P1_R1207_U48 , P1_U4013 );
not NOT1_10081 ( P1_R1207_U49 , P1_U3498 );
not NOT1_10082 ( P1_R1207_U50 , P1_U3486 );
not NOT1_10083 ( P1_R1207_U51 , P1_U3483 );
not NOT1_10084 ( P1_R1207_U52 , P1_U3061 );
not NOT1_10085 ( P1_R1207_U53 , P1_U3060 );
nand NAND2_10086 ( P1_R1207_U54 , P1_U3081 , P1_R1207_U42 );
not NOT1_10087 ( P1_R1207_U55 , P1_U3489 );
not NOT1_10088 ( P1_R1207_U56 , P1_U3070 );
not NOT1_10089 ( P1_R1207_U57 , P1_U3492 );
not NOT1_10090 ( P1_R1207_U58 , P1_U3078 );
not NOT1_10091 ( P1_R1207_U59 , P1_U3501 );
not NOT1_10092 ( P1_R1207_U60 , P1_U3495 );
not NOT1_10093 ( P1_R1207_U61 , P1_U3071 );
not NOT1_10094 ( P1_R1207_U62 , P1_U3072 );
not NOT1_10095 ( P1_R1207_U63 , P1_U3077 );
nand NAND2_10096 ( P1_R1207_U64 , P1_U3077 , P1_R1207_U60 );
not NOT1_10097 ( P1_R1207_U65 , P1_U3504 );
not NOT1_10098 ( P1_R1207_U66 , P1_U3067 );
nand NAND2_10099 ( P1_R1207_U67 , P1_R1207_U269 , P1_R1207_U268 );
not NOT1_10100 ( P1_R1207_U68 , P1_U3080 );
not NOT1_10101 ( P1_R1207_U69 , P1_U3509 );
not NOT1_10102 ( P1_R1207_U70 , P1_U3079 );
not NOT1_10103 ( P1_R1207_U71 , P1_U4015 );
not NOT1_10104 ( P1_R1207_U72 , P1_U3074 );
not NOT1_10105 ( P1_R1207_U73 , P1_U4012 );
not NOT1_10106 ( P1_R1207_U74 , P1_U4014 );
not NOT1_10107 ( P1_R1207_U75 , P1_U3064 );
not NOT1_10108 ( P1_R1207_U76 , P1_U3059 );
not NOT1_10109 ( P1_R1207_U77 , P1_U3073 );
nand NAND2_10110 ( P1_R1207_U78 , P1_U3073 , P1_R1207_U74 );
not NOT1_10111 ( P1_R1207_U79 , P1_U4011 );
not NOT1_10112 ( P1_R1207_U80 , P1_U3063 );
not NOT1_10113 ( P1_R1207_U81 , P1_U4010 );
not NOT1_10114 ( P1_R1207_U82 , P1_U3056 );
not NOT1_10115 ( P1_R1207_U83 , P1_U4008 );
not NOT1_10116 ( P1_R1207_U84 , P1_U3055 );
nand NAND2_10117 ( P1_R1207_U85 , P1_U3055 , P1_R1207_U47 );
not NOT1_10118 ( P1_R1207_U86 , P1_U3051 );
not NOT1_10119 ( P1_R1207_U87 , P1_U4007 );
not NOT1_10120 ( P1_R1207_U88 , P1_U3052 );
nand NAND2_10121 ( P1_R1207_U89 , P1_R1207_U299 , P1_R1207_U298 );
nand NAND2_10122 ( P1_R1207_U90 , P1_R1207_U78 , P1_R1207_U314 );
nand NAND2_10123 ( P1_R1207_U91 , P1_R1207_U64 , P1_R1207_U325 );
nand NAND2_10124 ( P1_R1207_U92 , P1_R1207_U54 , P1_R1207_U336 );
not NOT1_10125 ( P1_R1207_U93 , P1_U3075 );
nand NAND2_10126 ( P1_R1207_U94 , P1_R1207_U393 , P1_R1207_U392 );
nand NAND2_10127 ( P1_R1207_U95 , P1_R1207_U407 , P1_R1207_U406 );
nand NAND2_10128 ( P1_R1207_U96 , P1_R1207_U412 , P1_R1207_U411 );
nand NAND2_10129 ( P1_R1207_U97 , P1_R1207_U428 , P1_R1207_U427 );
nand NAND2_10130 ( P1_R1207_U98 , P1_R1207_U433 , P1_R1207_U432 );
nand NAND2_10131 ( P1_R1207_U99 , P1_R1207_U438 , P1_R1207_U437 );
nand NAND2_10132 ( P1_R1207_U100 , P1_R1207_U443 , P1_R1207_U442 );
nand NAND2_10133 ( P1_R1207_U101 , P1_R1207_U448 , P1_R1207_U447 );
nand NAND2_10134 ( P1_R1207_U102 , P1_R1207_U464 , P1_R1207_U463 );
nand NAND2_10135 ( P1_R1207_U103 , P1_R1207_U469 , P1_R1207_U468 );
nand NAND2_10136 ( P1_R1207_U104 , P1_R1207_U352 , P1_R1207_U351 );
nand NAND2_10137 ( P1_R1207_U105 , P1_R1207_U361 , P1_R1207_U360 );
nand NAND2_10138 ( P1_R1207_U106 , P1_R1207_U368 , P1_R1207_U367 );
nand NAND2_10139 ( P1_R1207_U107 , P1_R1207_U372 , P1_R1207_U371 );
nand NAND2_10140 ( P1_R1207_U108 , P1_R1207_U381 , P1_R1207_U380 );
nand NAND2_10141 ( P1_R1207_U109 , P1_R1207_U402 , P1_R1207_U401 );
nand NAND2_10142 ( P1_R1207_U110 , P1_R1207_U419 , P1_R1207_U418 );
nand NAND2_10143 ( P1_R1207_U111 , P1_R1207_U423 , P1_R1207_U422 );
nand NAND2_10144 ( P1_R1207_U112 , P1_R1207_U455 , P1_R1207_U454 );
nand NAND2_10145 ( P1_R1207_U113 , P1_R1207_U459 , P1_R1207_U458 );
nand NAND2_10146 ( P1_R1207_U114 , P1_R1207_U476 , P1_R1207_U475 );
and AND2_10147 ( P1_R1207_U115 , P1_R1207_U195 , P1_R1207_U183 );
and AND2_10148 ( P1_R1207_U116 , P1_R1207_U198 , P1_R1207_U199 );
and AND2_10149 ( P1_R1207_U117 , P1_R1207_U211 , P1_R1207_U185 );
and AND2_10150 ( P1_R1207_U118 , P1_R1207_U214 , P1_R1207_U215 );
and AND3_10151 ( P1_R1207_U119 , P1_R1207_U354 , P1_R1207_U353 , P1_R1207_U40 );
and AND2_10152 ( P1_R1207_U120 , P1_R1207_U357 , P1_R1207_U185 );
and AND2_10153 ( P1_R1207_U121 , P1_R1207_U230 , P1_R1207_U7 );
and AND2_10154 ( P1_R1207_U122 , P1_R1207_U364 , P1_R1207_U184 );
and AND3_10155 ( P1_R1207_U123 , P1_R1207_U374 , P1_R1207_U373 , P1_R1207_U29 );
and AND2_10156 ( P1_R1207_U124 , P1_R1207_U377 , P1_R1207_U183 );
and AND2_10157 ( P1_R1207_U125 , P1_R1207_U217 , P1_R1207_U8 );
and AND2_10158 ( P1_R1207_U126 , P1_R1207_U262 , P1_R1207_U180 );
and AND2_10159 ( P1_R1207_U127 , P1_R1207_U288 , P1_R1207_U181 );
and AND2_10160 ( P1_R1207_U128 , P1_R1207_U304 , P1_R1207_U305 );
and AND2_10161 ( P1_R1207_U129 , P1_R1207_U307 , P1_R1207_U386 );
and AND3_10162 ( P1_R1207_U130 , P1_R1207_U305 , P1_R1207_U304 , P1_R1207_U308 );
nand NAND2_10163 ( P1_R1207_U131 , P1_R1207_U390 , P1_R1207_U389 );
and AND3_10164 ( P1_R1207_U132 , P1_R1207_U395 , P1_R1207_U394 , P1_R1207_U85 );
and AND2_10165 ( P1_R1207_U133 , P1_R1207_U398 , P1_R1207_U182 );
nand NAND2_10166 ( P1_R1207_U134 , P1_R1207_U404 , P1_R1207_U403 );
nand NAND2_10167 ( P1_R1207_U135 , P1_R1207_U409 , P1_R1207_U408 );
and AND2_10168 ( P1_R1207_U136 , P1_R1207_U415 , P1_R1207_U181 );
nand NAND2_10169 ( P1_R1207_U137 , P1_R1207_U425 , P1_R1207_U424 );
nand NAND2_10170 ( P1_R1207_U138 , P1_R1207_U430 , P1_R1207_U429 );
nand NAND2_10171 ( P1_R1207_U139 , P1_R1207_U435 , P1_R1207_U434 );
nand NAND2_10172 ( P1_R1207_U140 , P1_R1207_U440 , P1_R1207_U439 );
nand NAND2_10173 ( P1_R1207_U141 , P1_R1207_U445 , P1_R1207_U444 );
and AND2_10174 ( P1_R1207_U142 , P1_R1207_U451 , P1_R1207_U180 );
nand NAND2_10175 ( P1_R1207_U143 , P1_R1207_U461 , P1_R1207_U460 );
nand NAND2_10176 ( P1_R1207_U144 , P1_R1207_U466 , P1_R1207_U465 );
and AND2_10177 ( P1_R1207_U145 , P1_R1207_U342 , P1_R1207_U9 );
and AND2_10178 ( P1_R1207_U146 , P1_R1207_U472 , P1_R1207_U179 );
and AND2_10179 ( P1_R1207_U147 , P1_R1207_U350 , P1_R1207_U349 );
nand NAND2_10180 ( P1_R1207_U148 , P1_R1207_U118 , P1_R1207_U212 );
and AND2_10181 ( P1_R1207_U149 , P1_R1207_U359 , P1_R1207_U358 );
and AND2_10182 ( P1_R1207_U150 , P1_R1207_U366 , P1_R1207_U365 );
and AND2_10183 ( P1_R1207_U151 , P1_R1207_U370 , P1_R1207_U369 );
nand NAND2_10184 ( P1_R1207_U152 , P1_R1207_U116 , P1_R1207_U196 );
and AND2_10185 ( P1_R1207_U153 , P1_R1207_U379 , P1_R1207_U378 );
not NOT1_10186 ( P1_R1207_U154 , P1_U4018 );
not NOT1_10187 ( P1_R1207_U155 , P1_U3053 );
and AND2_10188 ( P1_R1207_U156 , P1_R1207_U388 , P1_R1207_U387 );
nand NAND2_10189 ( P1_R1207_U157 , P1_R1207_U128 , P1_R1207_U302 );
and AND2_10190 ( P1_R1207_U158 , P1_R1207_U400 , P1_R1207_U399 );
nand NAND2_10191 ( P1_R1207_U159 , P1_R1207_U295 , P1_R1207_U294 );
nand NAND2_10192 ( P1_R1207_U160 , P1_R1207_U291 , P1_R1207_U290 );
and AND2_10193 ( P1_R1207_U161 , P1_R1207_U417 , P1_R1207_U416 );
and AND2_10194 ( P1_R1207_U162 , P1_R1207_U421 , P1_R1207_U420 );
nand NAND2_10195 ( P1_R1207_U163 , P1_R1207_U281 , P1_R1207_U280 );
nand NAND2_10196 ( P1_R1207_U164 , P1_R1207_U277 , P1_R1207_U276 );
not NOT1_10197 ( P1_R1207_U165 , P1_U3456 );
nand NAND2_10198 ( P1_R1207_U166 , P1_R1207_U273 , P1_R1207_U272 );
not NOT1_10199 ( P1_R1207_U167 , P1_U3507 );
nand NAND2_10200 ( P1_R1207_U168 , P1_R1207_U265 , P1_R1207_U264 );
and AND2_10201 ( P1_R1207_U169 , P1_R1207_U453 , P1_R1207_U452 );
and AND2_10202 ( P1_R1207_U170 , P1_R1207_U457 , P1_R1207_U456 );
nand NAND2_10203 ( P1_R1207_U171 , P1_R1207_U255 , P1_R1207_U254 );
nand NAND2_10204 ( P1_R1207_U172 , P1_R1207_U251 , P1_R1207_U250 );
nand NAND2_10205 ( P1_R1207_U173 , P1_R1207_U247 , P1_R1207_U246 );
and AND2_10206 ( P1_R1207_U174 , P1_R1207_U474 , P1_R1207_U473 );
nand NAND2_10207 ( P1_R1207_U175 , P1_R1207_U129 , P1_R1207_U157 );
not NOT1_10208 ( P1_R1207_U176 , P1_R1207_U85 );
not NOT1_10209 ( P1_R1207_U177 , P1_R1207_U29 );
not NOT1_10210 ( P1_R1207_U178 , P1_R1207_U40 );
nand NAND2_10211 ( P1_R1207_U179 , P1_U3483 , P1_R1207_U53 );
nand NAND2_10212 ( P1_R1207_U180 , P1_U3498 , P1_R1207_U62 );
nand NAND2_10213 ( P1_R1207_U181 , P1_U4013 , P1_R1207_U76 );
nand NAND2_10214 ( P1_R1207_U182 , P1_U4009 , P1_R1207_U84 );
nand NAND2_10215 ( P1_R1207_U183 , P1_U3459 , P1_R1207_U28 );
nand NAND2_10216 ( P1_R1207_U184 , P1_U3468 , P1_R1207_U35 );
nand NAND2_10217 ( P1_R1207_U185 , P1_U3474 , P1_R1207_U39 );
not NOT1_10218 ( P1_R1207_U186 , P1_R1207_U64 );
not NOT1_10219 ( P1_R1207_U187 , P1_R1207_U78 );
not NOT1_10220 ( P1_R1207_U188 , P1_R1207_U37 );
not NOT1_10221 ( P1_R1207_U189 , P1_R1207_U54 );
not NOT1_10222 ( P1_R1207_U190 , P1_R1207_U25 );
nand NAND2_10223 ( P1_R1207_U191 , P1_R1207_U190 , P1_R1207_U26 );
nand NAND2_10224 ( P1_R1207_U192 , P1_R1207_U191 , P1_R1207_U165 );
nand NAND2_10225 ( P1_R1207_U193 , P1_U3076 , P1_R1207_U25 );
not NOT1_10226 ( P1_R1207_U194 , P1_R1207_U46 );
nand NAND2_10227 ( P1_R1207_U195 , P1_U3462 , P1_R1207_U30 );
nand NAND2_10228 ( P1_R1207_U196 , P1_R1207_U115 , P1_R1207_U46 );
nand NAND2_10229 ( P1_R1207_U197 , P1_R1207_U30 , P1_R1207_U29 );
nand NAND2_10230 ( P1_R1207_U198 , P1_R1207_U197 , P1_R1207_U27 );
nand NAND2_10231 ( P1_R1207_U199 , P1_U3062 , P1_R1207_U177 );
not NOT1_10232 ( P1_R1207_U200 , P1_R1207_U152 );
nand NAND2_10233 ( P1_R1207_U201 , P1_U3471 , P1_R1207_U34 );
nand NAND2_10234 ( P1_R1207_U202 , P1_U3069 , P1_R1207_U31 );
nand NAND2_10235 ( P1_R1207_U203 , P1_U3065 , P1_R1207_U32 );
nand NAND2_10236 ( P1_R1207_U204 , P1_R1207_U188 , P1_R1207_U6 );
nand NAND2_10237 ( P1_R1207_U205 , P1_R1207_U7 , P1_R1207_U204 );
nand NAND2_10238 ( P1_R1207_U206 , P1_U3465 , P1_R1207_U36 );
nand NAND2_10239 ( P1_R1207_U207 , P1_U3471 , P1_R1207_U34 );
nand NAND3_10240 ( P1_R1207_U208 , P1_R1207_U206 , P1_R1207_U152 , P1_R1207_U6 );
nand NAND2_10241 ( P1_R1207_U209 , P1_R1207_U207 , P1_R1207_U205 );
not NOT1_10242 ( P1_R1207_U210 , P1_R1207_U44 );
nand NAND2_10243 ( P1_R1207_U211 , P1_U3477 , P1_R1207_U41 );
nand NAND2_10244 ( P1_R1207_U212 , P1_R1207_U117 , P1_R1207_U44 );
nand NAND2_10245 ( P1_R1207_U213 , P1_R1207_U41 , P1_R1207_U40 );
nand NAND2_10246 ( P1_R1207_U214 , P1_R1207_U213 , P1_R1207_U38 );
nand NAND2_10247 ( P1_R1207_U215 , P1_U3082 , P1_R1207_U178 );
not NOT1_10248 ( P1_R1207_U216 , P1_R1207_U148 );
nand NAND2_10249 ( P1_R1207_U217 , P1_U3480 , P1_R1207_U43 );
nand NAND2_10250 ( P1_R1207_U218 , P1_R1207_U217 , P1_R1207_U54 );
nand NAND2_10251 ( P1_R1207_U219 , P1_R1207_U210 , P1_R1207_U40 );
nand NAND2_10252 ( P1_R1207_U220 , P1_R1207_U120 , P1_R1207_U219 );
nand NAND2_10253 ( P1_R1207_U221 , P1_R1207_U44 , P1_R1207_U185 );
nand NAND2_10254 ( P1_R1207_U222 , P1_R1207_U119 , P1_R1207_U221 );
nand NAND2_10255 ( P1_R1207_U223 , P1_R1207_U40 , P1_R1207_U185 );
nand NAND2_10256 ( P1_R1207_U224 , P1_R1207_U206 , P1_R1207_U152 );
not NOT1_10257 ( P1_R1207_U225 , P1_R1207_U45 );
nand NAND2_10258 ( P1_R1207_U226 , P1_U3065 , P1_R1207_U32 );
nand NAND2_10259 ( P1_R1207_U227 , P1_R1207_U225 , P1_R1207_U226 );
nand NAND2_10260 ( P1_R1207_U228 , P1_R1207_U122 , P1_R1207_U227 );
nand NAND2_10261 ( P1_R1207_U229 , P1_R1207_U45 , P1_R1207_U184 );
nand NAND2_10262 ( P1_R1207_U230 , P1_U3471 , P1_R1207_U34 );
nand NAND2_10263 ( P1_R1207_U231 , P1_R1207_U121 , P1_R1207_U229 );
nand NAND2_10264 ( P1_R1207_U232 , P1_U3065 , P1_R1207_U32 );
nand NAND2_10265 ( P1_R1207_U233 , P1_R1207_U184 , P1_R1207_U232 );
nand NAND2_10266 ( P1_R1207_U234 , P1_R1207_U206 , P1_R1207_U37 );
nand NAND2_10267 ( P1_R1207_U235 , P1_R1207_U194 , P1_R1207_U29 );
nand NAND2_10268 ( P1_R1207_U236 , P1_R1207_U124 , P1_R1207_U235 );
nand NAND2_10269 ( P1_R1207_U237 , P1_R1207_U46 , P1_R1207_U183 );
nand NAND2_10270 ( P1_R1207_U238 , P1_R1207_U123 , P1_R1207_U237 );
nand NAND2_10271 ( P1_R1207_U239 , P1_R1207_U29 , P1_R1207_U183 );
nand NAND2_10272 ( P1_R1207_U240 , P1_U3486 , P1_R1207_U52 );
nand NAND2_10273 ( P1_R1207_U241 , P1_U3061 , P1_R1207_U50 );
nand NAND2_10274 ( P1_R1207_U242 , P1_U3060 , P1_R1207_U51 );
nand NAND2_10275 ( P1_R1207_U243 , P1_R1207_U189 , P1_R1207_U8 );
nand NAND2_10276 ( P1_R1207_U244 , P1_R1207_U9 , P1_R1207_U243 );
nand NAND2_10277 ( P1_R1207_U245 , P1_U3486 , P1_R1207_U52 );
nand NAND2_10278 ( P1_R1207_U246 , P1_R1207_U125 , P1_R1207_U148 );
nand NAND2_10279 ( P1_R1207_U247 , P1_R1207_U245 , P1_R1207_U244 );
not NOT1_10280 ( P1_R1207_U248 , P1_R1207_U173 );
nand NAND2_10281 ( P1_R1207_U249 , P1_U3489 , P1_R1207_U56 );
nand NAND2_10282 ( P1_R1207_U250 , P1_R1207_U249 , P1_R1207_U173 );
nand NAND2_10283 ( P1_R1207_U251 , P1_U3070 , P1_R1207_U55 );
not NOT1_10284 ( P1_R1207_U252 , P1_R1207_U172 );
nand NAND2_10285 ( P1_R1207_U253 , P1_U3492 , P1_R1207_U58 );
nand NAND2_10286 ( P1_R1207_U254 , P1_R1207_U253 , P1_R1207_U172 );
nand NAND2_10287 ( P1_R1207_U255 , P1_U3078 , P1_R1207_U57 );
not NOT1_10288 ( P1_R1207_U256 , P1_R1207_U171 );
nand NAND2_10289 ( P1_R1207_U257 , P1_U3501 , P1_R1207_U61 );
nand NAND2_10290 ( P1_R1207_U258 , P1_U3071 , P1_R1207_U59 );
nand NAND2_10291 ( P1_R1207_U259 , P1_U3072 , P1_R1207_U49 );
nand NAND2_10292 ( P1_R1207_U260 , P1_R1207_U186 , P1_R1207_U180 );
nand NAND2_10293 ( P1_R1207_U261 , P1_R1207_U10 , P1_R1207_U260 );
nand NAND2_10294 ( P1_R1207_U262 , P1_U3495 , P1_R1207_U63 );
nand NAND2_10295 ( P1_R1207_U263 , P1_U3501 , P1_R1207_U61 );
nand NAND3_10296 ( P1_R1207_U264 , P1_R1207_U171 , P1_R1207_U126 , P1_R1207_U257 );
nand NAND2_10297 ( P1_R1207_U265 , P1_R1207_U263 , P1_R1207_U261 );
not NOT1_10298 ( P1_R1207_U266 , P1_R1207_U168 );
nand NAND2_10299 ( P1_R1207_U267 , P1_U3504 , P1_R1207_U66 );
nand NAND2_10300 ( P1_R1207_U268 , P1_R1207_U267 , P1_R1207_U168 );
nand NAND2_10301 ( P1_R1207_U269 , P1_U3067 , P1_R1207_U65 );
not NOT1_10302 ( P1_R1207_U270 , P1_R1207_U67 );
nand NAND2_10303 ( P1_R1207_U271 , P1_R1207_U270 , P1_R1207_U68 );
nand NAND2_10304 ( P1_R1207_U272 , P1_R1207_U271 , P1_R1207_U167 );
nand NAND2_10305 ( P1_R1207_U273 , P1_U3080 , P1_R1207_U67 );
not NOT1_10306 ( P1_R1207_U274 , P1_R1207_U166 );
nand NAND2_10307 ( P1_R1207_U275 , P1_U3509 , P1_R1207_U70 );
nand NAND2_10308 ( P1_R1207_U276 , P1_R1207_U275 , P1_R1207_U166 );
nand NAND2_10309 ( P1_R1207_U277 , P1_U3079 , P1_R1207_U69 );
not NOT1_10310 ( P1_R1207_U278 , P1_R1207_U164 );
nand NAND2_10311 ( P1_R1207_U279 , P1_U4015 , P1_R1207_U72 );
nand NAND2_10312 ( P1_R1207_U280 , P1_R1207_U279 , P1_R1207_U164 );
nand NAND2_10313 ( P1_R1207_U281 , P1_U3074 , P1_R1207_U71 );
not NOT1_10314 ( P1_R1207_U282 , P1_R1207_U163 );
nand NAND2_10315 ( P1_R1207_U283 , P1_U4012 , P1_R1207_U75 );
nand NAND2_10316 ( P1_R1207_U284 , P1_U3064 , P1_R1207_U73 );
nand NAND2_10317 ( P1_R1207_U285 , P1_U3059 , P1_R1207_U48 );
nand NAND2_10318 ( P1_R1207_U286 , P1_R1207_U187 , P1_R1207_U181 );
nand NAND2_10319 ( P1_R1207_U287 , P1_R1207_U11 , P1_R1207_U286 );
nand NAND2_10320 ( P1_R1207_U288 , P1_U4014 , P1_R1207_U77 );
nand NAND2_10321 ( P1_R1207_U289 , P1_U4012 , P1_R1207_U75 );
nand NAND3_10322 ( P1_R1207_U290 , P1_R1207_U163 , P1_R1207_U127 , P1_R1207_U283 );
nand NAND2_10323 ( P1_R1207_U291 , P1_R1207_U289 , P1_R1207_U287 );
not NOT1_10324 ( P1_R1207_U292 , P1_R1207_U160 );
nand NAND2_10325 ( P1_R1207_U293 , P1_U4011 , P1_R1207_U80 );
nand NAND2_10326 ( P1_R1207_U294 , P1_R1207_U293 , P1_R1207_U160 );
nand NAND2_10327 ( P1_R1207_U295 , P1_U3063 , P1_R1207_U79 );
not NOT1_10328 ( P1_R1207_U296 , P1_R1207_U159 );
nand NAND2_10329 ( P1_R1207_U297 , P1_U4010 , P1_R1207_U82 );
nand NAND2_10330 ( P1_R1207_U298 , P1_R1207_U297 , P1_R1207_U159 );
nand NAND2_10331 ( P1_R1207_U299 , P1_U3056 , P1_R1207_U81 );
not NOT1_10332 ( P1_R1207_U300 , P1_R1207_U89 );
nand NAND2_10333 ( P1_R1207_U301 , P1_U4008 , P1_R1207_U86 );
nand NAND3_10334 ( P1_R1207_U302 , P1_R1207_U89 , P1_R1207_U182 , P1_R1207_U301 );
nand NAND2_10335 ( P1_R1207_U303 , P1_R1207_U86 , P1_R1207_U85 );
nand NAND2_10336 ( P1_R1207_U304 , P1_R1207_U303 , P1_R1207_U83 );
nand NAND2_10337 ( P1_R1207_U305 , P1_U3051 , P1_R1207_U176 );
not NOT1_10338 ( P1_R1207_U306 , P1_R1207_U157 );
nand NAND2_10339 ( P1_R1207_U307 , P1_U4007 , P1_R1207_U88 );
nand NAND2_10340 ( P1_R1207_U308 , P1_U3052 , P1_R1207_U87 );
nand NAND2_10341 ( P1_R1207_U309 , P1_R1207_U300 , P1_R1207_U85 );
nand NAND2_10342 ( P1_R1207_U310 , P1_R1207_U133 , P1_R1207_U309 );
nand NAND2_10343 ( P1_R1207_U311 , P1_R1207_U89 , P1_R1207_U182 );
nand NAND2_10344 ( P1_R1207_U312 , P1_R1207_U132 , P1_R1207_U311 );
nand NAND2_10345 ( P1_R1207_U313 , P1_R1207_U85 , P1_R1207_U182 );
nand NAND2_10346 ( P1_R1207_U314 , P1_R1207_U288 , P1_R1207_U163 );
not NOT1_10347 ( P1_R1207_U315 , P1_R1207_U90 );
nand NAND2_10348 ( P1_R1207_U316 , P1_U3059 , P1_R1207_U48 );
nand NAND2_10349 ( P1_R1207_U317 , P1_R1207_U315 , P1_R1207_U316 );
nand NAND2_10350 ( P1_R1207_U318 , P1_R1207_U136 , P1_R1207_U317 );
nand NAND2_10351 ( P1_R1207_U319 , P1_R1207_U90 , P1_R1207_U181 );
nand NAND2_10352 ( P1_R1207_U320 , P1_U4012 , P1_R1207_U75 );
nand NAND3_10353 ( P1_R1207_U321 , P1_R1207_U320 , P1_R1207_U319 , P1_R1207_U11 );
nand NAND2_10354 ( P1_R1207_U322 , P1_U3059 , P1_R1207_U48 );
nand NAND2_10355 ( P1_R1207_U323 , P1_R1207_U181 , P1_R1207_U322 );
nand NAND2_10356 ( P1_R1207_U324 , P1_R1207_U288 , P1_R1207_U78 );
nand NAND2_10357 ( P1_R1207_U325 , P1_R1207_U262 , P1_R1207_U171 );
not NOT1_10358 ( P1_R1207_U326 , P1_R1207_U91 );
nand NAND2_10359 ( P1_R1207_U327 , P1_U3072 , P1_R1207_U49 );
nand NAND2_10360 ( P1_R1207_U328 , P1_R1207_U326 , P1_R1207_U327 );
nand NAND2_10361 ( P1_R1207_U329 , P1_R1207_U142 , P1_R1207_U328 );
nand NAND2_10362 ( P1_R1207_U330 , P1_R1207_U91 , P1_R1207_U180 );
nand NAND2_10363 ( P1_R1207_U331 , P1_U3501 , P1_R1207_U61 );
nand NAND3_10364 ( P1_R1207_U332 , P1_R1207_U331 , P1_R1207_U330 , P1_R1207_U10 );
nand NAND2_10365 ( P1_R1207_U333 , P1_U3072 , P1_R1207_U49 );
nand NAND2_10366 ( P1_R1207_U334 , P1_R1207_U180 , P1_R1207_U333 );
nand NAND2_10367 ( P1_R1207_U335 , P1_R1207_U262 , P1_R1207_U64 );
nand NAND2_10368 ( P1_R1207_U336 , P1_R1207_U217 , P1_R1207_U148 );
not NOT1_10369 ( P1_R1207_U337 , P1_R1207_U92 );
nand NAND2_10370 ( P1_R1207_U338 , P1_U3060 , P1_R1207_U51 );
nand NAND2_10371 ( P1_R1207_U339 , P1_R1207_U337 , P1_R1207_U338 );
nand NAND2_10372 ( P1_R1207_U340 , P1_R1207_U146 , P1_R1207_U339 );
nand NAND2_10373 ( P1_R1207_U341 , P1_R1207_U92 , P1_R1207_U179 );
nand NAND2_10374 ( P1_R1207_U342 , P1_U3486 , P1_R1207_U52 );
nand NAND2_10375 ( P1_R1207_U343 , P1_R1207_U145 , P1_R1207_U341 );
nand NAND2_10376 ( P1_R1207_U344 , P1_U3060 , P1_R1207_U51 );
nand NAND2_10377 ( P1_R1207_U345 , P1_R1207_U179 , P1_R1207_U344 );
nand NAND2_10378 ( P1_R1207_U346 , P1_U3075 , P1_R1207_U24 );
nand NAND3_10379 ( P1_R1207_U347 , P1_R1207_U89 , P1_R1207_U182 , P1_R1207_U301 );
nand NAND3_10380 ( P1_R1207_U348 , P1_R1207_U12 , P1_R1207_U347 , P1_R1207_U130 );
nand NAND2_10381 ( P1_R1207_U349 , P1_U3480 , P1_R1207_U43 );
nand NAND2_10382 ( P1_R1207_U350 , P1_U3081 , P1_R1207_U42 );
nand NAND2_10383 ( P1_R1207_U351 , P1_R1207_U218 , P1_R1207_U148 );
nand NAND2_10384 ( P1_R1207_U352 , P1_R1207_U216 , P1_R1207_U147 );
nand NAND2_10385 ( P1_R1207_U353 , P1_U3477 , P1_R1207_U41 );
nand NAND2_10386 ( P1_R1207_U354 , P1_U3082 , P1_R1207_U38 );
nand NAND2_10387 ( P1_R1207_U355 , P1_U3477 , P1_R1207_U41 );
nand NAND2_10388 ( P1_R1207_U356 , P1_U3082 , P1_R1207_U38 );
nand NAND2_10389 ( P1_R1207_U357 , P1_R1207_U356 , P1_R1207_U355 );
nand NAND2_10390 ( P1_R1207_U358 , P1_U3474 , P1_R1207_U39 );
nand NAND2_10391 ( P1_R1207_U359 , P1_U3068 , P1_R1207_U22 );
nand NAND2_10392 ( P1_R1207_U360 , P1_R1207_U223 , P1_R1207_U44 );
nand NAND2_10393 ( P1_R1207_U361 , P1_R1207_U149 , P1_R1207_U210 );
nand NAND2_10394 ( P1_R1207_U362 , P1_U3471 , P1_R1207_U34 );
nand NAND2_10395 ( P1_R1207_U363 , P1_U3069 , P1_R1207_U31 );
nand NAND2_10396 ( P1_R1207_U364 , P1_R1207_U363 , P1_R1207_U362 );
nand NAND2_10397 ( P1_R1207_U365 , P1_U3468 , P1_R1207_U35 );
nand NAND2_10398 ( P1_R1207_U366 , P1_U3065 , P1_R1207_U32 );
nand NAND2_10399 ( P1_R1207_U367 , P1_R1207_U233 , P1_R1207_U45 );
nand NAND2_10400 ( P1_R1207_U368 , P1_R1207_U150 , P1_R1207_U225 );
nand NAND2_10401 ( P1_R1207_U369 , P1_U3465 , P1_R1207_U36 );
nand NAND2_10402 ( P1_R1207_U370 , P1_U3058 , P1_R1207_U33 );
nand NAND2_10403 ( P1_R1207_U371 , P1_R1207_U234 , P1_R1207_U152 );
nand NAND2_10404 ( P1_R1207_U372 , P1_R1207_U200 , P1_R1207_U151 );
nand NAND2_10405 ( P1_R1207_U373 , P1_U3462 , P1_R1207_U30 );
nand NAND2_10406 ( P1_R1207_U374 , P1_U3062 , P1_R1207_U27 );
nand NAND2_10407 ( P1_R1207_U375 , P1_U3462 , P1_R1207_U30 );
nand NAND2_10408 ( P1_R1207_U376 , P1_U3062 , P1_R1207_U27 );
nand NAND2_10409 ( P1_R1207_U377 , P1_R1207_U376 , P1_R1207_U375 );
nand NAND2_10410 ( P1_R1207_U378 , P1_U3459 , P1_R1207_U28 );
nand NAND2_10411 ( P1_R1207_U379 , P1_U3066 , P1_R1207_U23 );
nand NAND2_10412 ( P1_R1207_U380 , P1_R1207_U239 , P1_R1207_U46 );
nand NAND2_10413 ( P1_R1207_U381 , P1_R1207_U153 , P1_R1207_U194 );
nand NAND2_10414 ( P1_R1207_U382 , P1_U4018 , P1_R1207_U155 );
nand NAND2_10415 ( P1_R1207_U383 , P1_U3053 , P1_R1207_U154 );
nand NAND2_10416 ( P1_R1207_U384 , P1_U4018 , P1_R1207_U155 );
nand NAND2_10417 ( P1_R1207_U385 , P1_U3053 , P1_R1207_U154 );
nand NAND2_10418 ( P1_R1207_U386 , P1_R1207_U385 , P1_R1207_U384 );
nand NAND3_10419 ( P1_R1207_U387 , P1_U3052 , P1_R1207_U386 , P1_R1207_U87 );
nand NAND3_10420 ( P1_R1207_U388 , P1_R1207_U12 , P1_R1207_U88 , P1_U4007 );
nand NAND2_10421 ( P1_R1207_U389 , P1_U4007 , P1_R1207_U88 );
nand NAND2_10422 ( P1_R1207_U390 , P1_U3052 , P1_R1207_U87 );
not NOT1_10423 ( P1_R1207_U391 , P1_R1207_U131 );
nand NAND2_10424 ( P1_R1207_U392 , P1_R1207_U306 , P1_R1207_U391 );
nand NAND2_10425 ( P1_R1207_U393 , P1_R1207_U131 , P1_R1207_U157 );
nand NAND2_10426 ( P1_R1207_U394 , P1_U4008 , P1_R1207_U86 );
nand NAND2_10427 ( P1_R1207_U395 , P1_U3051 , P1_R1207_U83 );
nand NAND2_10428 ( P1_R1207_U396 , P1_U4008 , P1_R1207_U86 );
nand NAND2_10429 ( P1_R1207_U397 , P1_U3051 , P1_R1207_U83 );
nand NAND2_10430 ( P1_R1207_U398 , P1_R1207_U397 , P1_R1207_U396 );
nand NAND2_10431 ( P1_R1207_U399 , P1_U4009 , P1_R1207_U84 );
nand NAND2_10432 ( P1_R1207_U400 , P1_U3055 , P1_R1207_U47 );
nand NAND2_10433 ( P1_R1207_U401 , P1_R1207_U313 , P1_R1207_U89 );
nand NAND2_10434 ( P1_R1207_U402 , P1_R1207_U158 , P1_R1207_U300 );
nand NAND2_10435 ( P1_R1207_U403 , P1_U4010 , P1_R1207_U82 );
nand NAND2_10436 ( P1_R1207_U404 , P1_U3056 , P1_R1207_U81 );
not NOT1_10437 ( P1_R1207_U405 , P1_R1207_U134 );
nand NAND2_10438 ( P1_R1207_U406 , P1_R1207_U296 , P1_R1207_U405 );
nand NAND2_10439 ( P1_R1207_U407 , P1_R1207_U134 , P1_R1207_U159 );
nand NAND2_10440 ( P1_R1207_U408 , P1_U4011 , P1_R1207_U80 );
nand NAND2_10441 ( P1_R1207_U409 , P1_U3063 , P1_R1207_U79 );
not NOT1_10442 ( P1_R1207_U410 , P1_R1207_U135 );
nand NAND2_10443 ( P1_R1207_U411 , P1_R1207_U292 , P1_R1207_U410 );
nand NAND2_10444 ( P1_R1207_U412 , P1_R1207_U135 , P1_R1207_U160 );
nand NAND2_10445 ( P1_R1207_U413 , P1_U4012 , P1_R1207_U75 );
nand NAND2_10446 ( P1_R1207_U414 , P1_U3064 , P1_R1207_U73 );
nand NAND2_10447 ( P1_R1207_U415 , P1_R1207_U414 , P1_R1207_U413 );
nand NAND2_10448 ( P1_R1207_U416 , P1_U4013 , P1_R1207_U76 );
nand NAND2_10449 ( P1_R1207_U417 , P1_U3059 , P1_R1207_U48 );
nand NAND2_10450 ( P1_R1207_U418 , P1_R1207_U323 , P1_R1207_U90 );
nand NAND2_10451 ( P1_R1207_U419 , P1_R1207_U161 , P1_R1207_U315 );
nand NAND2_10452 ( P1_R1207_U420 , P1_U4014 , P1_R1207_U77 );
nand NAND2_10453 ( P1_R1207_U421 , P1_U3073 , P1_R1207_U74 );
nand NAND2_10454 ( P1_R1207_U422 , P1_R1207_U324 , P1_R1207_U163 );
nand NAND2_10455 ( P1_R1207_U423 , P1_R1207_U282 , P1_R1207_U162 );
nand NAND2_10456 ( P1_R1207_U424 , P1_U4015 , P1_R1207_U72 );
nand NAND2_10457 ( P1_R1207_U425 , P1_U3074 , P1_R1207_U71 );
not NOT1_10458 ( P1_R1207_U426 , P1_R1207_U137 );
nand NAND2_10459 ( P1_R1207_U427 , P1_R1207_U278 , P1_R1207_U426 );
nand NAND2_10460 ( P1_R1207_U428 , P1_R1207_U137 , P1_R1207_U164 );
nand NAND2_10461 ( P1_R1207_U429 , P1_U3456 , P1_R1207_U26 );
nand NAND2_10462 ( P1_R1207_U430 , P1_U3076 , P1_R1207_U165 );
not NOT1_10463 ( P1_R1207_U431 , P1_R1207_U138 );
nand NAND2_10464 ( P1_R1207_U432 , P1_R1207_U431 , P1_R1207_U190 );
nand NAND2_10465 ( P1_R1207_U433 , P1_R1207_U138 , P1_R1207_U25 );
nand NAND2_10466 ( P1_R1207_U434 , P1_U3509 , P1_R1207_U70 );
nand NAND2_10467 ( P1_R1207_U435 , P1_U3079 , P1_R1207_U69 );
not NOT1_10468 ( P1_R1207_U436 , P1_R1207_U139 );
nand NAND2_10469 ( P1_R1207_U437 , P1_R1207_U274 , P1_R1207_U436 );
nand NAND2_10470 ( P1_R1207_U438 , P1_R1207_U139 , P1_R1207_U166 );
nand NAND2_10471 ( P1_R1207_U439 , P1_U3507 , P1_R1207_U68 );
nand NAND2_10472 ( P1_R1207_U440 , P1_U3080 , P1_R1207_U167 );
not NOT1_10473 ( P1_R1207_U441 , P1_R1207_U140 );
nand NAND2_10474 ( P1_R1207_U442 , P1_R1207_U441 , P1_R1207_U270 );
nand NAND2_10475 ( P1_R1207_U443 , P1_R1207_U140 , P1_R1207_U67 );
nand NAND2_10476 ( P1_R1207_U444 , P1_U3504 , P1_R1207_U66 );
nand NAND2_10477 ( P1_R1207_U445 , P1_U3067 , P1_R1207_U65 );
not NOT1_10478 ( P1_R1207_U446 , P1_R1207_U141 );
nand NAND2_10479 ( P1_R1207_U447 , P1_R1207_U266 , P1_R1207_U446 );
nand NAND2_10480 ( P1_R1207_U448 , P1_R1207_U141 , P1_R1207_U168 );
nand NAND2_10481 ( P1_R1207_U449 , P1_U3501 , P1_R1207_U61 );
nand NAND2_10482 ( P1_R1207_U450 , P1_U3071 , P1_R1207_U59 );
nand NAND2_10483 ( P1_R1207_U451 , P1_R1207_U450 , P1_R1207_U449 );
nand NAND2_10484 ( P1_R1207_U452 , P1_U3498 , P1_R1207_U62 );
nand NAND2_10485 ( P1_R1207_U453 , P1_U3072 , P1_R1207_U49 );
nand NAND2_10486 ( P1_R1207_U454 , P1_R1207_U334 , P1_R1207_U91 );
nand NAND2_10487 ( P1_R1207_U455 , P1_R1207_U169 , P1_R1207_U326 );
nand NAND2_10488 ( P1_R1207_U456 , P1_U3495 , P1_R1207_U63 );
nand NAND2_10489 ( P1_R1207_U457 , P1_U3077 , P1_R1207_U60 );
nand NAND2_10490 ( P1_R1207_U458 , P1_R1207_U335 , P1_R1207_U171 );
nand NAND2_10491 ( P1_R1207_U459 , P1_R1207_U256 , P1_R1207_U170 );
nand NAND2_10492 ( P1_R1207_U460 , P1_U3492 , P1_R1207_U58 );
nand NAND2_10493 ( P1_R1207_U461 , P1_U3078 , P1_R1207_U57 );
not NOT1_10494 ( P1_R1207_U462 , P1_R1207_U143 );
nand NAND2_10495 ( P1_R1207_U463 , P1_R1207_U252 , P1_R1207_U462 );
nand NAND2_10496 ( P1_R1207_U464 , P1_R1207_U143 , P1_R1207_U172 );
nand NAND2_10497 ( P1_R1207_U465 , P1_U3489 , P1_R1207_U56 );
nand NAND2_10498 ( P1_R1207_U466 , P1_U3070 , P1_R1207_U55 );
not NOT1_10499 ( P1_R1207_U467 , P1_R1207_U144 );
nand NAND2_10500 ( P1_R1207_U468 , P1_R1207_U248 , P1_R1207_U467 );
nand NAND2_10501 ( P1_R1207_U469 , P1_R1207_U144 , P1_R1207_U173 );
nand NAND2_10502 ( P1_R1207_U470 , P1_U3486 , P1_R1207_U52 );
nand NAND2_10503 ( P1_R1207_U471 , P1_U3061 , P1_R1207_U50 );
nand NAND2_10504 ( P1_R1207_U472 , P1_R1207_U471 , P1_R1207_U470 );
nand NAND2_10505 ( P1_R1207_U473 , P1_U3483 , P1_R1207_U53 );
nand NAND2_10506 ( P1_R1207_U474 , P1_U3060 , P1_R1207_U51 );
nand NAND2_10507 ( P1_R1207_U475 , P1_R1207_U345 , P1_R1207_U92 );
nand NAND2_10508 ( P1_R1207_U476 , P1_R1207_U174 , P1_R1207_U337 );
and AND2_10509 ( P1_R1165_U4 , P1_R1165_U210 , P1_R1165_U209 );
and AND2_10510 ( P1_R1165_U5 , P1_R1165_U222 , P1_R1165_U221 );
and AND2_10511 ( P1_R1165_U6 , P1_R1165_U253 , P1_R1165_U252 );
and AND2_10512 ( P1_R1165_U7 , P1_R1165_U271 , P1_R1165_U270 );
and AND2_10513 ( P1_R1165_U8 , P1_R1165_U283 , P1_R1165_U282 );
and AND2_10514 ( P1_R1165_U9 , P1_R1165_U507 , P1_R1165_U506 );
and AND2_10515 ( P1_R1165_U10 , P1_R1165_U339 , P1_R1165_U336 );
and AND2_10516 ( P1_R1165_U11 , P1_R1165_U330 , P1_R1165_U327 );
and AND2_10517 ( P1_R1165_U12 , P1_R1165_U323 , P1_R1165_U320 );
and AND3_10518 ( P1_R1165_U13 , P1_R1165_U360 , P1_R1165_U311 , P1_R1165_U314 );
and AND2_10519 ( P1_R1165_U14 , P1_R1165_U245 , P1_R1165_U242 );
and AND2_10520 ( P1_R1165_U15 , P1_R1165_U238 , P1_R1165_U235 );
not NOT1_10521 ( P1_R1165_U16 , P1_U3209 );
not NOT1_10522 ( P1_R1165_U17 , P1_U3173 );
nand NAND2_10523 ( P1_R1165_U18 , P1_U3173 , P1_R1165_U58 );
not NOT1_10524 ( P1_R1165_U19 , P1_U3172 );
not NOT1_10525 ( P1_R1165_U20 , P1_U3175 );
not NOT1_10526 ( P1_R1165_U21 , P1_U3177 );
nand NAND2_10527 ( P1_R1165_U22 , P1_U3177 , P1_R1165_U61 );
not NOT1_10528 ( P1_R1165_U23 , P1_U3176 );
not NOT1_10529 ( P1_R1165_U24 , P1_U3179 );
not NOT1_10530 ( P1_R1165_U25 , P1_U3178 );
not NOT1_10531 ( P1_R1165_U26 , P1_U3174 );
not NOT1_10532 ( P1_R1165_U27 , P1_U3171 );
not NOT1_10533 ( P1_R1165_U28 , P1_U3170 );
nand NAND2_10534 ( P1_R1165_U29 , P1_R1165_U219 , P1_R1165_U218 );
nand NAND2_10535 ( P1_R1165_U30 , P1_R1165_U207 , P1_R1165_U206 );
not NOT1_10536 ( P1_R1165_U31 , P1_U3152 );
not NOT1_10537 ( P1_R1165_U32 , P1_U3153 );
not NOT1_10538 ( P1_R1165_U33 , P1_U3154 );
not NOT1_10539 ( P1_R1165_U34 , P1_U3155 );
not NOT1_10540 ( P1_R1165_U35 , P1_U3163 );
nand NAND2_10541 ( P1_R1165_U36 , P1_U3163 , P1_R1165_U71 );
not NOT1_10542 ( P1_R1165_U37 , P1_U3162 );
not NOT1_10543 ( P1_R1165_U38 , P1_U3169 );
not NOT1_10544 ( P1_R1165_U39 , P1_U3167 );
not NOT1_10545 ( P1_R1165_U40 , P1_U3168 );
nand NAND2_10546 ( P1_R1165_U41 , P1_U3168 , P1_R1165_U74 );
not NOT1_10547 ( P1_R1165_U42 , P1_U3166 );
not NOT1_10548 ( P1_R1165_U43 , P1_U3165 );
not NOT1_10549 ( P1_R1165_U44 , P1_U3164 );
not NOT1_10550 ( P1_R1165_U45 , P1_U3161 );
not NOT1_10551 ( P1_R1165_U46 , P1_U3159 );
not NOT1_10552 ( P1_R1165_U47 , P1_U3160 );
nand NAND2_10553 ( P1_R1165_U48 , P1_U3160 , P1_R1165_U80 );
not NOT1_10554 ( P1_R1165_U49 , P1_U3158 );
not NOT1_10555 ( P1_R1165_U50 , P1_U3157 );
not NOT1_10556 ( P1_R1165_U51 , P1_U3156 );
nand NAND2_10557 ( P1_R1165_U52 , P1_U3153 , P1_R1165_U69 );
nand NAND2_10558 ( P1_R1165_U53 , P1_R1165_U200 , P1_R1165_U309 );
nand NAND2_10559 ( P1_R1165_U54 , P1_R1165_U48 , P1_R1165_U316 );
nand NAND2_10560 ( P1_R1165_U55 , P1_R1165_U268 , P1_R1165_U267 );
nand NAND2_10561 ( P1_R1165_U56 , P1_R1165_U41 , P1_R1165_U332 );
nand NAND2_10562 ( P1_R1165_U57 , P1_R1165_U366 , P1_R1165_U365 );
nand NAND2_10563 ( P1_R1165_U58 , P1_R1165_U395 , P1_R1165_U394 );
nand NAND2_10564 ( P1_R1165_U59 , P1_R1165_U392 , P1_R1165_U391 );
nand NAND2_10565 ( P1_R1165_U60 , P1_R1165_U374 , P1_R1165_U373 );
nand NAND2_10566 ( P1_R1165_U61 , P1_R1165_U386 , P1_R1165_U385 );
nand NAND2_10567 ( P1_R1165_U62 , P1_R1165_U383 , P1_R1165_U382 );
nand NAND2_10568 ( P1_R1165_U63 , P1_R1165_U377 , P1_R1165_U376 );
nand NAND2_10569 ( P1_R1165_U64 , P1_R1165_U380 , P1_R1165_U379 );
nand NAND2_10570 ( P1_R1165_U65 , P1_R1165_U389 , P1_R1165_U388 );
nand NAND2_10571 ( P1_R1165_U66 , P1_R1165_U398 , P1_R1165_U397 );
nand NAND2_10572 ( P1_R1165_U67 , P1_R1165_U438 , P1_R1165_U437 );
nand NAND2_10573 ( P1_R1165_U68 , P1_R1165_U441 , P1_R1165_U440 );
nand NAND2_10574 ( P1_R1165_U69 , P1_R1165_U444 , P1_R1165_U443 );
nand NAND2_10575 ( P1_R1165_U70 , P1_R1165_U447 , P1_R1165_U446 );
nand NAND2_10576 ( P1_R1165_U71 , P1_R1165_U471 , P1_R1165_U470 );
nand NAND2_10577 ( P1_R1165_U72 , P1_R1165_U468 , P1_R1165_U467 );
nand NAND2_10578 ( P1_R1165_U73 , P1_R1165_U450 , P1_R1165_U449 );
nand NAND2_10579 ( P1_R1165_U74 , P1_R1165_U459 , P1_R1165_U458 );
nand NAND2_10580 ( P1_R1165_U75 , P1_R1165_U453 , P1_R1165_U452 );
nand NAND2_10581 ( P1_R1165_U76 , P1_R1165_U456 , P1_R1165_U455 );
nand NAND2_10582 ( P1_R1165_U77 , P1_R1165_U462 , P1_R1165_U461 );
nand NAND2_10583 ( P1_R1165_U78 , P1_R1165_U465 , P1_R1165_U464 );
nand NAND2_10584 ( P1_R1165_U79 , P1_R1165_U474 , P1_R1165_U473 );
nand NAND2_10585 ( P1_R1165_U80 , P1_R1165_U483 , P1_R1165_U482 );
nand NAND2_10586 ( P1_R1165_U81 , P1_R1165_U477 , P1_R1165_U476 );
nand NAND2_10587 ( P1_R1165_U82 , P1_R1165_U480 , P1_R1165_U479 );
nand NAND2_10588 ( P1_R1165_U83 , P1_R1165_U486 , P1_R1165_U485 );
nand NAND2_10589 ( P1_R1165_U84 , P1_R1165_U489 , P1_R1165_U488 );
nand NAND2_10590 ( P1_R1165_U85 , P1_R1165_U495 , P1_R1165_U494 );
nand NAND2_10591 ( P1_R1165_U86 , P1_R1165_U602 , P1_R1165_U601 );
nand NAND2_10592 ( P1_R1165_U87 , P1_R1165_U401 , P1_R1165_U400 );
nand NAND2_10593 ( P1_R1165_U88 , P1_R1165_U408 , P1_R1165_U407 );
nand NAND2_10594 ( P1_R1165_U89 , P1_R1165_U415 , P1_R1165_U414 );
nand NAND2_10595 ( P1_R1165_U90 , P1_R1165_U422 , P1_R1165_U421 );
nand NAND2_10596 ( P1_R1165_U91 , P1_R1165_U429 , P1_R1165_U428 );
nand NAND2_10597 ( P1_R1165_U92 , P1_R1165_U436 , P1_R1165_U435 );
nand NAND2_10598 ( P1_R1165_U93 , P1_R1165_U498 , P1_R1165_U497 );
nand NAND2_10599 ( P1_R1165_U94 , P1_R1165_U505 , P1_R1165_U504 );
nand NAND2_10600 ( P1_R1165_U95 , P1_R1165_U512 , P1_R1165_U511 );
nand NAND2_10601 ( P1_R1165_U96 , P1_R1165_U517 , P1_R1165_U516 );
nand NAND2_10602 ( P1_R1165_U97 , P1_R1165_U524 , P1_R1165_U523 );
nand NAND2_10603 ( P1_R1165_U98 , P1_R1165_U531 , P1_R1165_U530 );
nand NAND2_10604 ( P1_R1165_U99 , P1_R1165_U538 , P1_R1165_U537 );
nand NAND2_10605 ( P1_R1165_U100 , P1_R1165_U545 , P1_R1165_U544 );
nand NAND2_10606 ( P1_R1165_U101 , P1_R1165_U550 , P1_R1165_U549 );
nand NAND2_10607 ( P1_R1165_U102 , P1_R1165_U557 , P1_R1165_U556 );
nand NAND2_10608 ( P1_R1165_U103 , P1_R1165_U564 , P1_R1165_U563 );
nand NAND2_10609 ( P1_R1165_U104 , P1_R1165_U571 , P1_R1165_U570 );
nand NAND2_10610 ( P1_R1165_U105 , P1_R1165_U578 , P1_R1165_U577 );
nand NAND2_10611 ( P1_R1165_U106 , P1_R1165_U585 , P1_R1165_U584 );
nand NAND2_10612 ( P1_R1165_U107 , P1_R1165_U590 , P1_R1165_U589 );
nand NAND2_10613 ( P1_R1165_U108 , P1_R1165_U597 , P1_R1165_U596 );
and AND2_10614 ( P1_R1165_U109 , P1_R1165_U213 , P1_R1165_U212 );
and AND2_10615 ( P1_R1165_U110 , P1_R1165_U226 , P1_R1165_U225 );
and AND3_10616 ( P1_R1165_U111 , P1_R1165_U410 , P1_R1165_U409 , P1_R1165_U18 );
and AND2_10617 ( P1_R1165_U112 , P1_R1165_U237 , P1_R1165_U5 );
and AND3_10618 ( P1_R1165_U113 , P1_R1165_U431 , P1_R1165_U430 , P1_R1165_U22 );
and AND2_10619 ( P1_R1165_U114 , P1_R1165_U244 , P1_R1165_U4 );
and AND2_10620 ( P1_R1165_U115 , P1_R1165_U257 , P1_R1165_U6 );
and AND2_10621 ( P1_R1165_U116 , P1_R1165_U255 , P1_R1165_U195 );
and AND2_10622 ( P1_R1165_U117 , P1_R1165_U275 , P1_R1165_U274 );
and AND2_10623 ( P1_R1165_U118 , P1_R1165_U287 , P1_R1165_U8 );
and AND2_10624 ( P1_R1165_U119 , P1_R1165_U285 , P1_R1165_U196 );
and AND2_10625 ( P1_R1165_U120 , P1_R1165_U359 , P1_R1165_U52 );
and AND2_10626 ( P1_R1165_U121 , P1_R1165_U308 , P1_R1165_U303 );
and AND2_10627 ( P1_R1165_U122 , P1_R1165_U356 , P1_R1165_U307 );
nand NAND2_10628 ( P1_R1165_U123 , P1_R1165_U492 , P1_R1165_U491 );
and AND2_10629 ( P1_R1165_U124 , P1_R1165_U352 , P1_R1165_U52 );
and AND2_10630 ( P1_R1165_U125 , P1_R1165_U442 , P1_R1165_U33 );
and AND2_10631 ( P1_R1165_U126 , P1_R1165_U200 , P1_R1165_U197 );
and AND2_10632 ( P1_R1165_U127 , P1_R1165_U313 , P1_R1165_U193 );
and AND2_10633 ( P1_R1165_U128 , P1_R1165_U9 , P1_R1165_U197 );
and AND3_10634 ( P1_R1165_U129 , P1_R1165_U533 , P1_R1165_U532 , P1_R1165_U196 );
and AND2_10635 ( P1_R1165_U130 , P1_R1165_U322 , P1_R1165_U8 );
and AND3_10636 ( P1_R1165_U131 , P1_R1165_U559 , P1_R1165_U558 , P1_R1165_U36 );
and AND2_10637 ( P1_R1165_U132 , P1_R1165_U329 , P1_R1165_U7 );
and AND3_10638 ( P1_R1165_U133 , P1_R1165_U580 , P1_R1165_U579 , P1_R1165_U195 );
and AND2_10639 ( P1_R1165_U134 , P1_R1165_U338 , P1_R1165_U6 );
nand NAND2_10640 ( P1_R1165_U135 , P1_R1165_U599 , P1_R1165_U598 );
not NOT1_10641 ( P1_R1165_U136 , P1_U3199 );
and AND2_10642 ( P1_R1165_U137 , P1_R1165_U369 , P1_R1165_U368 );
not NOT1_10643 ( P1_R1165_U138 , P1_U3204 );
not NOT1_10644 ( P1_R1165_U139 , P1_U3208 );
not NOT1_10645 ( P1_R1165_U140 , P1_U3207 );
not NOT1_10646 ( P1_R1165_U141 , P1_U3205 );
not NOT1_10647 ( P1_R1165_U142 , P1_U3206 );
not NOT1_10648 ( P1_R1165_U143 , P1_U3203 );
not NOT1_10649 ( P1_R1165_U144 , P1_U3201 );
not NOT1_10650 ( P1_R1165_U145 , P1_U3202 );
not NOT1_10651 ( P1_R1165_U146 , P1_U3200 );
nand NAND2_10652 ( P1_R1165_U147 , P1_R1165_U231 , P1_R1165_U230 );
and AND2_10653 ( P1_R1165_U148 , P1_R1165_U403 , P1_R1165_U402 );
nand NAND2_10654 ( P1_R1165_U149 , P1_R1165_U110 , P1_R1165_U227 );
and AND2_10655 ( P1_R1165_U150 , P1_R1165_U417 , P1_R1165_U416 );
nand NAND2_10656 ( P1_R1165_U151 , P1_R1165_U361 , P1_R1165_U350 );
and AND2_10657 ( P1_R1165_U152 , P1_R1165_U424 , P1_R1165_U423 );
nand NAND2_10658 ( P1_R1165_U153 , P1_R1165_U109 , P1_R1165_U214 );
not NOT1_10659 ( P1_R1165_U154 , P1_U3181 );
not NOT1_10660 ( P1_R1165_U155 , P1_U3183 );
not NOT1_10661 ( P1_R1165_U156 , P1_U3182 );
not NOT1_10662 ( P1_R1165_U157 , P1_U3184 );
not NOT1_10663 ( P1_R1165_U158 , P1_U3198 );
not NOT1_10664 ( P1_R1165_U159 , P1_U3195 );
not NOT1_10665 ( P1_R1165_U160 , P1_U3196 );
not NOT1_10666 ( P1_R1165_U161 , P1_U3197 );
not NOT1_10667 ( P1_R1165_U162 , P1_U3194 );
not NOT1_10668 ( P1_R1165_U163 , P1_U3193 );
not NOT1_10669 ( P1_R1165_U164 , P1_U3191 );
not NOT1_10670 ( P1_R1165_U165 , P1_U3192 );
not NOT1_10671 ( P1_R1165_U166 , P1_U3190 );
not NOT1_10672 ( P1_R1165_U167 , P1_U3187 );
not NOT1_10673 ( P1_R1165_U168 , P1_U3188 );
not NOT1_10674 ( P1_R1165_U169 , P1_U3189 );
not NOT1_10675 ( P1_R1165_U170 , P1_U3186 );
not NOT1_10676 ( P1_R1165_U171 , P1_U3185 );
not NOT1_10677 ( P1_R1165_U172 , P1_U3151 );
not NOT1_10678 ( P1_R1165_U173 , P1_U3180 );
and AND2_10679 ( P1_R1165_U174 , P1_R1165_U500 , P1_R1165_U499 );
nand NAND2_10680 ( P1_R1165_U175 , P1_R1165_U124 , P1_R1165_U304 );
nand NAND2_10681 ( P1_R1165_U176 , P1_R1165_U298 , P1_R1165_U297 );
and AND2_10682 ( P1_R1165_U177 , P1_R1165_U519 , P1_R1165_U518 );
nand NAND2_10683 ( P1_R1165_U178 , P1_R1165_U294 , P1_R1165_U293 );
and AND2_10684 ( P1_R1165_U179 , P1_R1165_U526 , P1_R1165_U525 );
nand NAND2_10685 ( P1_R1165_U180 , P1_R1165_U290 , P1_R1165_U289 );
and AND2_10686 ( P1_R1165_U181 , P1_R1165_U540 , P1_R1165_U539 );
nand NAND2_10687 ( P1_R1165_U182 , P1_R1165_U203 , P1_R1165_U202 );
nand NAND2_10688 ( P1_R1165_U183 , P1_R1165_U280 , P1_R1165_U279 );
and AND2_10689 ( P1_R1165_U184 , P1_R1165_U552 , P1_R1165_U551 );
nand NAND2_10690 ( P1_R1165_U185 , P1_R1165_U117 , P1_R1165_U276 );
and AND2_10691 ( P1_R1165_U186 , P1_R1165_U566 , P1_R1165_U565 );
nand NAND2_10692 ( P1_R1165_U187 , P1_R1165_U264 , P1_R1165_U263 );
and AND2_10693 ( P1_R1165_U188 , P1_R1165_U573 , P1_R1165_U572 );
nand NAND2_10694 ( P1_R1165_U189 , P1_R1165_U260 , P1_R1165_U259 );
nand NAND2_10695 ( P1_R1165_U190 , P1_R1165_U250 , P1_R1165_U249 );
and AND2_10696 ( P1_R1165_U191 , P1_R1165_U592 , P1_R1165_U591 );
nand NAND2_10697 ( P1_R1165_U192 , P1_R1165_U363 , P1_R1165_U353 );
nand NAND2_10698 ( P1_R1165_U193 , P1_R1165_U355 , P1_R1165_U354 );
not NOT1_10699 ( P1_R1165_U194 , P1_R1165_U22 );
nand NAND2_10700 ( P1_R1165_U195 , P1_U3167 , P1_R1165_U76 );
nand NAND2_10701 ( P1_R1165_U196 , P1_U3159 , P1_R1165_U82 );
nand NAND2_10702 ( P1_R1165_U197 , P1_U3154 , P1_R1165_U68 );
not NOT1_10703 ( P1_R1165_U198 , P1_R1165_U41 );
not NOT1_10704 ( P1_R1165_U199 , P1_R1165_U48 );
nand NAND2_10705 ( P1_R1165_U200 , P1_U3155 , P1_R1165_U70 );
or OR2_10706 ( P1_R1165_U201 , P1_U3209 , P1_U3179 );
nand NAND2_10707 ( P1_R1165_U202 , P1_R1165_U63 , P1_R1165_U201 );
nand NAND2_10708 ( P1_R1165_U203 , P1_U3179 , P1_U3209 );
not NOT1_10709 ( P1_R1165_U204 , P1_R1165_U182 );
nand NAND2_10710 ( P1_R1165_U205 , P1_R1165_U381 , P1_R1165_U25 );
nand NAND2_10711 ( P1_R1165_U206 , P1_R1165_U205 , P1_R1165_U182 );
nand NAND2_10712 ( P1_R1165_U207 , P1_U3178 , P1_R1165_U64 );
not NOT1_10713 ( P1_R1165_U208 , P1_R1165_U30 );
nand NAND2_10714 ( P1_R1165_U209 , P1_R1165_U384 , P1_R1165_U23 );
nand NAND2_10715 ( P1_R1165_U210 , P1_R1165_U387 , P1_R1165_U21 );
nand NAND2_10716 ( P1_R1165_U211 , P1_R1165_U23 , P1_R1165_U22 );
nand NAND2_10717 ( P1_R1165_U212 , P1_R1165_U62 , P1_R1165_U211 );
nand NAND2_10718 ( P1_R1165_U213 , P1_U3176 , P1_R1165_U194 );
nand NAND2_10719 ( P1_R1165_U214 , P1_R1165_U4 , P1_R1165_U30 );
not NOT1_10720 ( P1_R1165_U215 , P1_R1165_U153 );
nand NAND2_10721 ( P1_R1165_U216 , P1_R1165_U375 , P1_R1165_U20 );
nand NAND2_10722 ( P1_R1165_U217 , P1_R1165_U390 , P1_R1165_U26 );
nand NAND2_10723 ( P1_R1165_U218 , P1_R1165_U217 , P1_R1165_U151 );
nand NAND2_10724 ( P1_R1165_U219 , P1_U3174 , P1_R1165_U65 );
not NOT1_10725 ( P1_R1165_U220 , P1_R1165_U29 );
nand NAND2_10726 ( P1_R1165_U221 , P1_R1165_U393 , P1_R1165_U19 );
nand NAND2_10727 ( P1_R1165_U222 , P1_R1165_U396 , P1_R1165_U17 );
not NOT1_10728 ( P1_R1165_U223 , P1_R1165_U18 );
nand NAND2_10729 ( P1_R1165_U224 , P1_R1165_U19 , P1_R1165_U18 );
nand NAND2_10730 ( P1_R1165_U225 , P1_R1165_U59 , P1_R1165_U224 );
nand NAND2_10731 ( P1_R1165_U226 , P1_U3172 , P1_R1165_U223 );
nand NAND2_10732 ( P1_R1165_U227 , P1_R1165_U5 , P1_R1165_U29 );
not NOT1_10733 ( P1_R1165_U228 , P1_R1165_U149 );
nand NAND2_10734 ( P1_R1165_U229 , P1_R1165_U399 , P1_R1165_U27 );
nand NAND2_10735 ( P1_R1165_U230 , P1_R1165_U229 , P1_R1165_U149 );
nand NAND2_10736 ( P1_R1165_U231 , P1_U3171 , P1_R1165_U66 );
not NOT1_10737 ( P1_R1165_U232 , P1_R1165_U147 );
nand NAND2_10738 ( P1_R1165_U233 , P1_R1165_U396 , P1_R1165_U17 );
nand NAND2_10739 ( P1_R1165_U234 , P1_R1165_U233 , P1_R1165_U29 );
nand NAND2_10740 ( P1_R1165_U235 , P1_R1165_U111 , P1_R1165_U234 );
nand NAND2_10741 ( P1_R1165_U236 , P1_R1165_U220 , P1_R1165_U18 );
nand NAND2_10742 ( P1_R1165_U237 , P1_U3172 , P1_R1165_U59 );
nand NAND2_10743 ( P1_R1165_U238 , P1_R1165_U112 , P1_R1165_U236 );
nand NAND2_10744 ( P1_R1165_U239 , P1_R1165_U396 , P1_R1165_U17 );
nand NAND2_10745 ( P1_R1165_U240 , P1_R1165_U387 , P1_R1165_U21 );
nand NAND2_10746 ( P1_R1165_U241 , P1_R1165_U240 , P1_R1165_U30 );
nand NAND2_10747 ( P1_R1165_U242 , P1_R1165_U113 , P1_R1165_U241 );
nand NAND2_10748 ( P1_R1165_U243 , P1_R1165_U208 , P1_R1165_U22 );
nand NAND2_10749 ( P1_R1165_U244 , P1_U3176 , P1_R1165_U62 );
nand NAND2_10750 ( P1_R1165_U245 , P1_R1165_U114 , P1_R1165_U243 );
nand NAND2_10751 ( P1_R1165_U246 , P1_R1165_U387 , P1_R1165_U21 );
nand NAND2_10752 ( P1_R1165_U247 , P1_R1165_U367 , P1_R1165_U28 );
nand NAND2_10753 ( P1_R1165_U248 , P1_R1165_U451 , P1_R1165_U38 );
nand NAND2_10754 ( P1_R1165_U249 , P1_R1165_U248 , P1_R1165_U192 );
nand NAND2_10755 ( P1_R1165_U250 , P1_U3169 , P1_R1165_U73 );
not NOT1_10756 ( P1_R1165_U251 , P1_R1165_U190 );
nand NAND2_10757 ( P1_R1165_U252 , P1_R1165_U454 , P1_R1165_U42 );
nand NAND2_10758 ( P1_R1165_U253 , P1_R1165_U457 , P1_R1165_U39 );
nand NAND2_10759 ( P1_R1165_U254 , P1_R1165_U198 , P1_R1165_U6 );
nand NAND2_10760 ( P1_R1165_U255 , P1_U3166 , P1_R1165_U75 );
nand NAND2_10761 ( P1_R1165_U256 , P1_R1165_U116 , P1_R1165_U254 );
nand NAND2_10762 ( P1_R1165_U257 , P1_R1165_U460 , P1_R1165_U40 );
nand NAND2_10763 ( P1_R1165_U258 , P1_R1165_U454 , P1_R1165_U42 );
nand NAND2_10764 ( P1_R1165_U259 , P1_R1165_U115 , P1_R1165_U190 );
nand NAND2_10765 ( P1_R1165_U260 , P1_R1165_U258 , P1_R1165_U256 );
not NOT1_10766 ( P1_R1165_U261 , P1_R1165_U189 );
nand NAND2_10767 ( P1_R1165_U262 , P1_R1165_U463 , P1_R1165_U43 );
nand NAND2_10768 ( P1_R1165_U263 , P1_R1165_U262 , P1_R1165_U189 );
nand NAND2_10769 ( P1_R1165_U264 , P1_U3165 , P1_R1165_U77 );
not NOT1_10770 ( P1_R1165_U265 , P1_R1165_U187 );
nand NAND2_10771 ( P1_R1165_U266 , P1_R1165_U466 , P1_R1165_U44 );
nand NAND2_10772 ( P1_R1165_U267 , P1_R1165_U266 , P1_R1165_U187 );
nand NAND2_10773 ( P1_R1165_U268 , P1_U3164 , P1_R1165_U78 );
not NOT1_10774 ( P1_R1165_U269 , P1_R1165_U55 );
nand NAND2_10775 ( P1_R1165_U270 , P1_R1165_U469 , P1_R1165_U37 );
nand NAND2_10776 ( P1_R1165_U271 , P1_R1165_U472 , P1_R1165_U35 );
not NOT1_10777 ( P1_R1165_U272 , P1_R1165_U36 );
nand NAND2_10778 ( P1_R1165_U273 , P1_R1165_U37 , P1_R1165_U36 );
nand NAND2_10779 ( P1_R1165_U274 , P1_R1165_U72 , P1_R1165_U273 );
nand NAND2_10780 ( P1_R1165_U275 , P1_U3162 , P1_R1165_U272 );
nand NAND2_10781 ( P1_R1165_U276 , P1_R1165_U7 , P1_R1165_U55 );
not NOT1_10782 ( P1_R1165_U277 , P1_R1165_U185 );
nand NAND2_10783 ( P1_R1165_U278 , P1_R1165_U475 , P1_R1165_U45 );
nand NAND2_10784 ( P1_R1165_U279 , P1_R1165_U278 , P1_R1165_U185 );
nand NAND2_10785 ( P1_R1165_U280 , P1_U3161 , P1_R1165_U79 );
not NOT1_10786 ( P1_R1165_U281 , P1_R1165_U183 );
nand NAND2_10787 ( P1_R1165_U282 , P1_R1165_U478 , P1_R1165_U49 );
nand NAND2_10788 ( P1_R1165_U283 , P1_R1165_U481 , P1_R1165_U46 );
nand NAND2_10789 ( P1_R1165_U284 , P1_R1165_U199 , P1_R1165_U8 );
nand NAND2_10790 ( P1_R1165_U285 , P1_U3158 , P1_R1165_U81 );
nand NAND2_10791 ( P1_R1165_U286 , P1_R1165_U119 , P1_R1165_U284 );
nand NAND2_10792 ( P1_R1165_U287 , P1_R1165_U484 , P1_R1165_U47 );
nand NAND2_10793 ( P1_R1165_U288 , P1_R1165_U478 , P1_R1165_U49 );
nand NAND2_10794 ( P1_R1165_U289 , P1_R1165_U118 , P1_R1165_U183 );
nand NAND2_10795 ( P1_R1165_U290 , P1_R1165_U288 , P1_R1165_U286 );
not NOT1_10796 ( P1_R1165_U291 , P1_R1165_U180 );
nand NAND2_10797 ( P1_R1165_U292 , P1_R1165_U487 , P1_R1165_U50 );
nand NAND2_10798 ( P1_R1165_U293 , P1_R1165_U292 , P1_R1165_U180 );
nand NAND2_10799 ( P1_R1165_U294 , P1_U3157 , P1_R1165_U83 );
not NOT1_10800 ( P1_R1165_U295 , P1_R1165_U178 );
nand NAND2_10801 ( P1_R1165_U296 , P1_R1165_U490 , P1_R1165_U51 );
nand NAND2_10802 ( P1_R1165_U297 , P1_R1165_U296 , P1_R1165_U178 );
nand NAND2_10803 ( P1_R1165_U298 , P1_U3156 , P1_R1165_U84 );
not NOT1_10804 ( P1_R1165_U299 , P1_R1165_U176 );
nand NAND2_10805 ( P1_R1165_U300 , P1_R1165_U442 , P1_R1165_U33 );
nand NAND2_10806 ( P1_R1165_U301 , P1_R1165_U200 , P1_R1165_U197 );
not NOT1_10807 ( P1_R1165_U302 , P1_R1165_U52 );
nand NAND2_10808 ( P1_R1165_U303 , P1_R1165_U448 , P1_R1165_U34 );
nand NAND3_10809 ( P1_R1165_U304 , P1_R1165_U176 , P1_R1165_U303 , P1_R1165_U193 );
not NOT1_10810 ( P1_R1165_U305 , P1_R1165_U175 );
nand NAND2_10811 ( P1_R1165_U306 , P1_R1165_U439 , P1_R1165_U31 );
nand NAND2_10812 ( P1_R1165_U307 , P1_U3152 , P1_R1165_U67 );
nand NAND2_10813 ( P1_R1165_U308 , P1_R1165_U439 , P1_R1165_U31 );
nand NAND2_10814 ( P1_R1165_U309 , P1_R1165_U303 , P1_R1165_U176 );
not NOT1_10815 ( P1_R1165_U310 , P1_R1165_U53 );
nand NAND2_10816 ( P1_R1165_U311 , P1_R1165_U125 , P1_R1165_U9 );
nand NAND2_10817 ( P1_R1165_U312 , P1_R1165_U126 , P1_R1165_U309 );
nand NAND2_10818 ( P1_R1165_U313 , P1_U3153 , P1_R1165_U69 );
nand NAND2_10819 ( P1_R1165_U314 , P1_R1165_U127 , P1_R1165_U312 );
nand NAND2_10820 ( P1_R1165_U315 , P1_R1165_U442 , P1_R1165_U33 );
nand NAND2_10821 ( P1_R1165_U316 , P1_R1165_U287 , P1_R1165_U183 );
not NOT1_10822 ( P1_R1165_U317 , P1_R1165_U54 );
nand NAND2_10823 ( P1_R1165_U318 , P1_R1165_U481 , P1_R1165_U46 );
nand NAND2_10824 ( P1_R1165_U319 , P1_R1165_U318 , P1_R1165_U54 );
nand NAND2_10825 ( P1_R1165_U320 , P1_R1165_U129 , P1_R1165_U319 );
nand NAND2_10826 ( P1_R1165_U321 , P1_R1165_U317 , P1_R1165_U196 );
nand NAND2_10827 ( P1_R1165_U322 , P1_U3158 , P1_R1165_U81 );
nand NAND2_10828 ( P1_R1165_U323 , P1_R1165_U130 , P1_R1165_U321 );
nand NAND2_10829 ( P1_R1165_U324 , P1_R1165_U481 , P1_R1165_U46 );
nand NAND2_10830 ( P1_R1165_U325 , P1_R1165_U472 , P1_R1165_U35 );
nand NAND2_10831 ( P1_R1165_U326 , P1_R1165_U325 , P1_R1165_U55 );
nand NAND2_10832 ( P1_R1165_U327 , P1_R1165_U131 , P1_R1165_U326 );
nand NAND2_10833 ( P1_R1165_U328 , P1_R1165_U269 , P1_R1165_U36 );
nand NAND2_10834 ( P1_R1165_U329 , P1_U3162 , P1_R1165_U72 );
nand NAND2_10835 ( P1_R1165_U330 , P1_R1165_U132 , P1_R1165_U328 );
nand NAND2_10836 ( P1_R1165_U331 , P1_R1165_U472 , P1_R1165_U35 );
nand NAND2_10837 ( P1_R1165_U332 , P1_R1165_U257 , P1_R1165_U190 );
not NOT1_10838 ( P1_R1165_U333 , P1_R1165_U56 );
nand NAND2_10839 ( P1_R1165_U334 , P1_R1165_U457 , P1_R1165_U39 );
nand NAND2_10840 ( P1_R1165_U335 , P1_R1165_U334 , P1_R1165_U56 );
nand NAND2_10841 ( P1_R1165_U336 , P1_R1165_U133 , P1_R1165_U335 );
nand NAND2_10842 ( P1_R1165_U337 , P1_R1165_U333 , P1_R1165_U195 );
nand NAND2_10843 ( P1_R1165_U338 , P1_U3166 , P1_R1165_U75 );
nand NAND2_10844 ( P1_R1165_U339 , P1_R1165_U134 , P1_R1165_U337 );
nand NAND2_10845 ( P1_R1165_U340 , P1_R1165_U457 , P1_R1165_U39 );
nand NAND2_10846 ( P1_R1165_U341 , P1_R1165_U239 , P1_R1165_U18 );
nand NAND2_10847 ( P1_R1165_U342 , P1_R1165_U246 , P1_R1165_U22 );
nand NAND2_10848 ( P1_R1165_U343 , P1_R1165_U315 , P1_R1165_U197 );
nand NAND2_10849 ( P1_R1165_U344 , P1_R1165_U303 , P1_R1165_U200 );
nand NAND2_10850 ( P1_R1165_U345 , P1_R1165_U324 , P1_R1165_U196 );
nand NAND2_10851 ( P1_R1165_U346 , P1_R1165_U287 , P1_R1165_U48 );
nand NAND2_10852 ( P1_R1165_U347 , P1_R1165_U331 , P1_R1165_U36 );
nand NAND2_10853 ( P1_R1165_U348 , P1_R1165_U340 , P1_R1165_U195 );
nand NAND2_10854 ( P1_R1165_U349 , P1_R1165_U257 , P1_R1165_U41 );
nand NAND2_10855 ( P1_R1165_U350 , P1_U3175 , P1_R1165_U60 );
nand NAND3_10856 ( P1_R1165_U351 , P1_R1165_U352 , P1_R1165_U304 , P1_R1165_U120 );
nand NAND2_10857 ( P1_R1165_U352 , P1_R1165_U301 , P1_R1165_U193 );
nand NAND2_10858 ( P1_R1165_U353 , P1_U3170 , P1_R1165_U57 );
nand NAND2_10859 ( P1_R1165_U354 , P1_R1165_U69 , P1_R1165_U300 );
nand NAND2_10860 ( P1_R1165_U355 , P1_U3153 , P1_R1165_U300 );
nand NAND3_10861 ( P1_R1165_U356 , P1_R1165_U301 , P1_R1165_U193 , P1_R1165_U308 );
nand NAND3_10862 ( P1_R1165_U357 , P1_R1165_U176 , P1_R1165_U193 , P1_R1165_U121 );
nand NAND2_10863 ( P1_R1165_U358 , P1_R1165_U302 , P1_R1165_U308 );
nand NAND2_10864 ( P1_R1165_U359 , P1_U3152 , P1_R1165_U67 );
nand NAND2_10865 ( P1_R1165_U360 , P1_R1165_U128 , P1_R1165_U310 );
nand NAND2_10866 ( P1_R1165_U361 , P1_R1165_U216 , P1_R1165_U153 );
not NOT1_10867 ( P1_R1165_U362 , P1_R1165_U151 );
nand NAND2_10868 ( P1_R1165_U363 , P1_R1165_U247 , P1_R1165_U147 );
not NOT1_10869 ( P1_R1165_U364 , P1_R1165_U192 );
nand NAND2_10870 ( P1_R1165_U365 , P1_U3209 , P1_R1165_U136 );
nand NAND2_10871 ( P1_R1165_U366 , P1_U3199 , P1_R1165_U16 );
not NOT1_10872 ( P1_R1165_U367 , P1_R1165_U57 );
nand NAND2_10873 ( P1_R1165_U368 , P1_R1165_U367 , P1_U3170 );
nand NAND2_10874 ( P1_R1165_U369 , P1_R1165_U57 , P1_R1165_U28 );
nand NAND2_10875 ( P1_R1165_U370 , P1_R1165_U367 , P1_U3170 );
nand NAND2_10876 ( P1_R1165_U371 , P1_R1165_U57 , P1_R1165_U28 );
nand NAND2_10877 ( P1_R1165_U372 , P1_R1165_U371 , P1_R1165_U370 );
nand NAND2_10878 ( P1_R1165_U373 , P1_U3209 , P1_R1165_U138 );
nand NAND2_10879 ( P1_R1165_U374 , P1_U3204 , P1_R1165_U16 );
not NOT1_10880 ( P1_R1165_U375 , P1_R1165_U60 );
nand NAND2_10881 ( P1_R1165_U376 , P1_U3209 , P1_R1165_U139 );
nand NAND2_10882 ( P1_R1165_U377 , P1_U3208 , P1_R1165_U16 );
not NOT1_10883 ( P1_R1165_U378 , P1_R1165_U63 );
nand NAND2_10884 ( P1_R1165_U379 , P1_U3209 , P1_R1165_U140 );
nand NAND2_10885 ( P1_R1165_U380 , P1_U3207 , P1_R1165_U16 );
not NOT1_10886 ( P1_R1165_U381 , P1_R1165_U64 );
nand NAND2_10887 ( P1_R1165_U382 , P1_U3209 , P1_R1165_U141 );
nand NAND2_10888 ( P1_R1165_U383 , P1_U3205 , P1_R1165_U16 );
not NOT1_10889 ( P1_R1165_U384 , P1_R1165_U62 );
nand NAND2_10890 ( P1_R1165_U385 , P1_U3209 , P1_R1165_U142 );
nand NAND2_10891 ( P1_R1165_U386 , P1_U3206 , P1_R1165_U16 );
not NOT1_10892 ( P1_R1165_U387 , P1_R1165_U61 );
nand NAND2_10893 ( P1_R1165_U388 , P1_U3209 , P1_R1165_U143 );
nand NAND2_10894 ( P1_R1165_U389 , P1_U3203 , P1_R1165_U16 );
not NOT1_10895 ( P1_R1165_U390 , P1_R1165_U65 );
nand NAND2_10896 ( P1_R1165_U391 , P1_U3209 , P1_R1165_U144 );
nand NAND2_10897 ( P1_R1165_U392 , P1_U3201 , P1_R1165_U16 );
not NOT1_10898 ( P1_R1165_U393 , P1_R1165_U59 );
nand NAND2_10899 ( P1_R1165_U394 , P1_U3209 , P1_R1165_U145 );
nand NAND2_10900 ( P1_R1165_U395 , P1_U3202 , P1_R1165_U16 );
not NOT1_10901 ( P1_R1165_U396 , P1_R1165_U58 );
nand NAND2_10902 ( P1_R1165_U397 , P1_U3209 , P1_R1165_U146 );
nand NAND2_10903 ( P1_R1165_U398 , P1_U3200 , P1_R1165_U16 );
not NOT1_10904 ( P1_R1165_U399 , P1_R1165_U66 );
nand NAND2_10905 ( P1_R1165_U400 , P1_R1165_U137 , P1_R1165_U147 );
nand NAND2_10906 ( P1_R1165_U401 , P1_R1165_U232 , P1_R1165_U372 );
nand NAND2_10907 ( P1_R1165_U402 , P1_R1165_U399 , P1_U3171 );
nand NAND2_10908 ( P1_R1165_U403 , P1_R1165_U66 , P1_R1165_U27 );
nand NAND2_10909 ( P1_R1165_U404 , P1_R1165_U399 , P1_U3171 );
nand NAND2_10910 ( P1_R1165_U405 , P1_R1165_U66 , P1_R1165_U27 );
nand NAND2_10911 ( P1_R1165_U406 , P1_R1165_U405 , P1_R1165_U404 );
nand NAND2_10912 ( P1_R1165_U407 , P1_R1165_U148 , P1_R1165_U149 );
nand NAND2_10913 ( P1_R1165_U408 , P1_R1165_U228 , P1_R1165_U406 );
nand NAND2_10914 ( P1_R1165_U409 , P1_R1165_U393 , P1_U3172 );
nand NAND2_10915 ( P1_R1165_U410 , P1_R1165_U59 , P1_R1165_U19 );
nand NAND2_10916 ( P1_R1165_U411 , P1_R1165_U396 , P1_U3173 );
nand NAND2_10917 ( P1_R1165_U412 , P1_R1165_U58 , P1_R1165_U17 );
nand NAND2_10918 ( P1_R1165_U413 , P1_R1165_U412 , P1_R1165_U411 );
nand NAND2_10919 ( P1_R1165_U414 , P1_R1165_U341 , P1_R1165_U29 );
nand NAND2_10920 ( P1_R1165_U415 , P1_R1165_U413 , P1_R1165_U220 );
nand NAND2_10921 ( P1_R1165_U416 , P1_R1165_U390 , P1_U3174 );
nand NAND2_10922 ( P1_R1165_U417 , P1_R1165_U65 , P1_R1165_U26 );
nand NAND2_10923 ( P1_R1165_U418 , P1_R1165_U390 , P1_U3174 );
nand NAND2_10924 ( P1_R1165_U419 , P1_R1165_U65 , P1_R1165_U26 );
nand NAND2_10925 ( P1_R1165_U420 , P1_R1165_U419 , P1_R1165_U418 );
nand NAND2_10926 ( P1_R1165_U421 , P1_R1165_U150 , P1_R1165_U151 );
nand NAND2_10927 ( P1_R1165_U422 , P1_R1165_U362 , P1_R1165_U420 );
nand NAND2_10928 ( P1_R1165_U423 , P1_R1165_U375 , P1_U3175 );
nand NAND2_10929 ( P1_R1165_U424 , P1_R1165_U60 , P1_R1165_U20 );
nand NAND2_10930 ( P1_R1165_U425 , P1_R1165_U375 , P1_U3175 );
nand NAND2_10931 ( P1_R1165_U426 , P1_R1165_U60 , P1_R1165_U20 );
nand NAND2_10932 ( P1_R1165_U427 , P1_R1165_U426 , P1_R1165_U425 );
nand NAND2_10933 ( P1_R1165_U428 , P1_R1165_U152 , P1_R1165_U153 );
nand NAND2_10934 ( P1_R1165_U429 , P1_R1165_U215 , P1_R1165_U427 );
nand NAND2_10935 ( P1_R1165_U430 , P1_R1165_U384 , P1_U3176 );
nand NAND2_10936 ( P1_R1165_U431 , P1_R1165_U62 , P1_R1165_U23 );
nand NAND2_10937 ( P1_R1165_U432 , P1_R1165_U387 , P1_U3177 );
nand NAND2_10938 ( P1_R1165_U433 , P1_R1165_U61 , P1_R1165_U21 );
nand NAND2_10939 ( P1_R1165_U434 , P1_R1165_U433 , P1_R1165_U432 );
nand NAND2_10940 ( P1_R1165_U435 , P1_R1165_U342 , P1_R1165_U30 );
nand NAND2_10941 ( P1_R1165_U436 , P1_R1165_U434 , P1_R1165_U208 );
nand NAND2_10942 ( P1_R1165_U437 , P1_U3209 , P1_R1165_U154 );
nand NAND2_10943 ( P1_R1165_U438 , P1_U3181 , P1_R1165_U16 );
not NOT1_10944 ( P1_R1165_U439 , P1_R1165_U67 );
nand NAND2_10945 ( P1_R1165_U440 , P1_U3209 , P1_R1165_U155 );
nand NAND2_10946 ( P1_R1165_U441 , P1_U3183 , P1_R1165_U16 );
not NOT1_10947 ( P1_R1165_U442 , P1_R1165_U68 );
nand NAND2_10948 ( P1_R1165_U443 , P1_U3209 , P1_R1165_U156 );
nand NAND2_10949 ( P1_R1165_U444 , P1_U3182 , P1_R1165_U16 );
not NOT1_10950 ( P1_R1165_U445 , P1_R1165_U69 );
nand NAND2_10951 ( P1_R1165_U446 , P1_U3209 , P1_R1165_U157 );
nand NAND2_10952 ( P1_R1165_U447 , P1_U3184 , P1_R1165_U16 );
not NOT1_10953 ( P1_R1165_U448 , P1_R1165_U70 );
nand NAND2_10954 ( P1_R1165_U449 , P1_U3209 , P1_R1165_U158 );
nand NAND2_10955 ( P1_R1165_U450 , P1_U3198 , P1_R1165_U16 );
not NOT1_10956 ( P1_R1165_U451 , P1_R1165_U73 );
nand NAND2_10957 ( P1_R1165_U452 , P1_U3209 , P1_R1165_U159 );
nand NAND2_10958 ( P1_R1165_U453 , P1_U3195 , P1_R1165_U16 );
not NOT1_10959 ( P1_R1165_U454 , P1_R1165_U75 );
nand NAND2_10960 ( P1_R1165_U455 , P1_U3209 , P1_R1165_U160 );
nand NAND2_10961 ( P1_R1165_U456 , P1_U3196 , P1_R1165_U16 );
not NOT1_10962 ( P1_R1165_U457 , P1_R1165_U76 );
nand NAND2_10963 ( P1_R1165_U458 , P1_U3209 , P1_R1165_U161 );
nand NAND2_10964 ( P1_R1165_U459 , P1_U3197 , P1_R1165_U16 );
not NOT1_10965 ( P1_R1165_U460 , P1_R1165_U74 );
nand NAND2_10966 ( P1_R1165_U461 , P1_U3209 , P1_R1165_U162 );
nand NAND2_10967 ( P1_R1165_U462 , P1_U3194 , P1_R1165_U16 );
not NOT1_10968 ( P1_R1165_U463 , P1_R1165_U77 );
nand NAND2_10969 ( P1_R1165_U464 , P1_U3209 , P1_R1165_U163 );
nand NAND2_10970 ( P1_R1165_U465 , P1_U3193 , P1_R1165_U16 );
not NOT1_10971 ( P1_R1165_U466 , P1_R1165_U78 );
nand NAND2_10972 ( P1_R1165_U467 , P1_U3209 , P1_R1165_U164 );
nand NAND2_10973 ( P1_R1165_U468 , P1_U3191 , P1_R1165_U16 );
not NOT1_10974 ( P1_R1165_U469 , P1_R1165_U72 );
nand NAND2_10975 ( P1_R1165_U470 , P1_U3209 , P1_R1165_U165 );
nand NAND2_10976 ( P1_R1165_U471 , P1_U3192 , P1_R1165_U16 );
not NOT1_10977 ( P1_R1165_U472 , P1_R1165_U71 );
nand NAND2_10978 ( P1_R1165_U473 , P1_U3209 , P1_R1165_U166 );
nand NAND2_10979 ( P1_R1165_U474 , P1_U3190 , P1_R1165_U16 );
not NOT1_10980 ( P1_R1165_U475 , P1_R1165_U79 );
nand NAND2_10981 ( P1_R1165_U476 , P1_U3209 , P1_R1165_U167 );
nand NAND2_10982 ( P1_R1165_U477 , P1_U3187 , P1_R1165_U16 );
not NOT1_10983 ( P1_R1165_U478 , P1_R1165_U81 );
nand NAND2_10984 ( P1_R1165_U479 , P1_U3209 , P1_R1165_U168 );
nand NAND2_10985 ( P1_R1165_U480 , P1_U3188 , P1_R1165_U16 );
not NOT1_10986 ( P1_R1165_U481 , P1_R1165_U82 );
nand NAND2_10987 ( P1_R1165_U482 , P1_U3209 , P1_R1165_U169 );
nand NAND2_10988 ( P1_R1165_U483 , P1_U3189 , P1_R1165_U16 );
not NOT1_10989 ( P1_R1165_U484 , P1_R1165_U80 );
nand NAND2_10990 ( P1_R1165_U485 , P1_U3209 , P1_R1165_U170 );
nand NAND2_10991 ( P1_R1165_U486 , P1_U3186 , P1_R1165_U16 );
not NOT1_10992 ( P1_R1165_U487 , P1_R1165_U83 );
nand NAND2_10993 ( P1_R1165_U488 , P1_U3209 , P1_R1165_U171 );
nand NAND2_10994 ( P1_R1165_U489 , P1_U3185 , P1_R1165_U16 );
not NOT1_10995 ( P1_R1165_U490 , P1_R1165_U84 );
nand NAND2_10996 ( P1_R1165_U491 , P1_U3209 , P1_R1165_U172 );
nand NAND2_10997 ( P1_R1165_U492 , P1_U3151 , P1_R1165_U16 );
not NOT1_10998 ( P1_R1165_U493 , P1_R1165_U123 );
nand NAND2_10999 ( P1_R1165_U494 , P1_U3180 , P1_R1165_U493 );
nand NAND2_11000 ( P1_R1165_U495 , P1_R1165_U123 , P1_R1165_U173 );
not NOT1_11001 ( P1_R1165_U496 , P1_R1165_U85 );
nand NAND3_11002 ( P1_R1165_U497 , P1_R1165_U351 , P1_R1165_U306 , P1_R1165_U496 );
nand NAND4_11003 ( P1_R1165_U498 , P1_R1165_U358 , P1_R1165_U357 , P1_R1165_U122 , P1_R1165_U85 );
nand NAND2_11004 ( P1_R1165_U499 , P1_R1165_U439 , P1_U3152 );
nand NAND2_11005 ( P1_R1165_U500 , P1_R1165_U67 , P1_R1165_U31 );
nand NAND2_11006 ( P1_R1165_U501 , P1_R1165_U439 , P1_U3152 );
nand NAND2_11007 ( P1_R1165_U502 , P1_R1165_U67 , P1_R1165_U31 );
nand NAND2_11008 ( P1_R1165_U503 , P1_R1165_U502 , P1_R1165_U501 );
nand NAND2_11009 ( P1_R1165_U504 , P1_R1165_U174 , P1_R1165_U175 );
nand NAND2_11010 ( P1_R1165_U505 , P1_R1165_U305 , P1_R1165_U503 );
nand NAND2_11011 ( P1_R1165_U506 , P1_R1165_U445 , P1_U3153 );
nand NAND2_11012 ( P1_R1165_U507 , P1_R1165_U69 , P1_R1165_U32 );
nand NAND2_11013 ( P1_R1165_U508 , P1_R1165_U442 , P1_U3154 );
nand NAND2_11014 ( P1_R1165_U509 , P1_R1165_U68 , P1_R1165_U33 );
nand NAND2_11015 ( P1_R1165_U510 , P1_R1165_U509 , P1_R1165_U508 );
nand NAND2_11016 ( P1_R1165_U511 , P1_R1165_U343 , P1_R1165_U53 );
nand NAND2_11017 ( P1_R1165_U512 , P1_R1165_U510 , P1_R1165_U310 );
nand NAND2_11018 ( P1_R1165_U513 , P1_R1165_U448 , P1_U3155 );
nand NAND2_11019 ( P1_R1165_U514 , P1_R1165_U70 , P1_R1165_U34 );
nand NAND2_11020 ( P1_R1165_U515 , P1_R1165_U514 , P1_R1165_U513 );
nand NAND2_11021 ( P1_R1165_U516 , P1_R1165_U344 , P1_R1165_U176 );
nand NAND2_11022 ( P1_R1165_U517 , P1_R1165_U299 , P1_R1165_U515 );
nand NAND2_11023 ( P1_R1165_U518 , P1_R1165_U490 , P1_U3156 );
nand NAND2_11024 ( P1_R1165_U519 , P1_R1165_U84 , P1_R1165_U51 );
nand NAND2_11025 ( P1_R1165_U520 , P1_R1165_U490 , P1_U3156 );
nand NAND2_11026 ( P1_R1165_U521 , P1_R1165_U84 , P1_R1165_U51 );
nand NAND2_11027 ( P1_R1165_U522 , P1_R1165_U521 , P1_R1165_U520 );
nand NAND2_11028 ( P1_R1165_U523 , P1_R1165_U177 , P1_R1165_U178 );
nand NAND2_11029 ( P1_R1165_U524 , P1_R1165_U295 , P1_R1165_U522 );
nand NAND2_11030 ( P1_R1165_U525 , P1_R1165_U487 , P1_U3157 );
nand NAND2_11031 ( P1_R1165_U526 , P1_R1165_U83 , P1_R1165_U50 );
nand NAND2_11032 ( P1_R1165_U527 , P1_R1165_U487 , P1_U3157 );
nand NAND2_11033 ( P1_R1165_U528 , P1_R1165_U83 , P1_R1165_U50 );
nand NAND2_11034 ( P1_R1165_U529 , P1_R1165_U528 , P1_R1165_U527 );
nand NAND2_11035 ( P1_R1165_U530 , P1_R1165_U179 , P1_R1165_U180 );
nand NAND2_11036 ( P1_R1165_U531 , P1_R1165_U291 , P1_R1165_U529 );
nand NAND2_11037 ( P1_R1165_U532 , P1_R1165_U478 , P1_U3158 );
nand NAND2_11038 ( P1_R1165_U533 , P1_R1165_U81 , P1_R1165_U49 );
nand NAND2_11039 ( P1_R1165_U534 , P1_R1165_U481 , P1_U3159 );
nand NAND2_11040 ( P1_R1165_U535 , P1_R1165_U82 , P1_R1165_U46 );
nand NAND2_11041 ( P1_R1165_U536 , P1_R1165_U535 , P1_R1165_U534 );
nand NAND2_11042 ( P1_R1165_U537 , P1_R1165_U345 , P1_R1165_U54 );
nand NAND2_11043 ( P1_R1165_U538 , P1_R1165_U536 , P1_R1165_U317 );
nand NAND2_11044 ( P1_R1165_U539 , P1_R1165_U381 , P1_U3178 );
nand NAND2_11045 ( P1_R1165_U540 , P1_R1165_U64 , P1_R1165_U25 );
nand NAND2_11046 ( P1_R1165_U541 , P1_R1165_U381 , P1_U3178 );
nand NAND2_11047 ( P1_R1165_U542 , P1_R1165_U64 , P1_R1165_U25 );
nand NAND2_11048 ( P1_R1165_U543 , P1_R1165_U542 , P1_R1165_U541 );
nand NAND2_11049 ( P1_R1165_U544 , P1_R1165_U181 , P1_R1165_U182 );
nand NAND2_11050 ( P1_R1165_U545 , P1_R1165_U204 , P1_R1165_U543 );
nand NAND2_11051 ( P1_R1165_U546 , P1_R1165_U484 , P1_U3160 );
nand NAND2_11052 ( P1_R1165_U547 , P1_R1165_U80 , P1_R1165_U47 );
nand NAND2_11053 ( P1_R1165_U548 , P1_R1165_U547 , P1_R1165_U546 );
nand NAND2_11054 ( P1_R1165_U549 , P1_R1165_U346 , P1_R1165_U183 );
nand NAND2_11055 ( P1_R1165_U550 , P1_R1165_U281 , P1_R1165_U548 );
nand NAND2_11056 ( P1_R1165_U551 , P1_R1165_U475 , P1_U3161 );
nand NAND2_11057 ( P1_R1165_U552 , P1_R1165_U79 , P1_R1165_U45 );
nand NAND2_11058 ( P1_R1165_U553 , P1_R1165_U475 , P1_U3161 );
nand NAND2_11059 ( P1_R1165_U554 , P1_R1165_U79 , P1_R1165_U45 );
nand NAND2_11060 ( P1_R1165_U555 , P1_R1165_U554 , P1_R1165_U553 );
nand NAND2_11061 ( P1_R1165_U556 , P1_R1165_U184 , P1_R1165_U185 );
nand NAND2_11062 ( P1_R1165_U557 , P1_R1165_U277 , P1_R1165_U555 );
nand NAND2_11063 ( P1_R1165_U558 , P1_R1165_U469 , P1_U3162 );
nand NAND2_11064 ( P1_R1165_U559 , P1_R1165_U72 , P1_R1165_U37 );
nand NAND2_11065 ( P1_R1165_U560 , P1_R1165_U472 , P1_U3163 );
nand NAND2_11066 ( P1_R1165_U561 , P1_R1165_U71 , P1_R1165_U35 );
nand NAND2_11067 ( P1_R1165_U562 , P1_R1165_U561 , P1_R1165_U560 );
nand NAND2_11068 ( P1_R1165_U563 , P1_R1165_U347 , P1_R1165_U55 );
nand NAND2_11069 ( P1_R1165_U564 , P1_R1165_U562 , P1_R1165_U269 );
nand NAND2_11070 ( P1_R1165_U565 , P1_R1165_U466 , P1_U3164 );
nand NAND2_11071 ( P1_R1165_U566 , P1_R1165_U78 , P1_R1165_U44 );
nand NAND2_11072 ( P1_R1165_U567 , P1_R1165_U466 , P1_U3164 );
nand NAND2_11073 ( P1_R1165_U568 , P1_R1165_U78 , P1_R1165_U44 );
nand NAND2_11074 ( P1_R1165_U569 , P1_R1165_U568 , P1_R1165_U567 );
nand NAND2_11075 ( P1_R1165_U570 , P1_R1165_U186 , P1_R1165_U187 );
nand NAND2_11076 ( P1_R1165_U571 , P1_R1165_U265 , P1_R1165_U569 );
nand NAND2_11077 ( P1_R1165_U572 , P1_R1165_U463 , P1_U3165 );
nand NAND2_11078 ( P1_R1165_U573 , P1_R1165_U77 , P1_R1165_U43 );
nand NAND2_11079 ( P1_R1165_U574 , P1_R1165_U463 , P1_U3165 );
nand NAND2_11080 ( P1_R1165_U575 , P1_R1165_U77 , P1_R1165_U43 );
nand NAND2_11081 ( P1_R1165_U576 , P1_R1165_U575 , P1_R1165_U574 );
nand NAND2_11082 ( P1_R1165_U577 , P1_R1165_U188 , P1_R1165_U189 );
nand NAND2_11083 ( P1_R1165_U578 , P1_R1165_U261 , P1_R1165_U576 );
nand NAND2_11084 ( P1_R1165_U579 , P1_R1165_U454 , P1_U3166 );
nand NAND2_11085 ( P1_R1165_U580 , P1_R1165_U75 , P1_R1165_U42 );
nand NAND2_11086 ( P1_R1165_U581 , P1_R1165_U457 , P1_U3167 );
nand NAND2_11087 ( P1_R1165_U582 , P1_R1165_U76 , P1_R1165_U39 );
nand NAND2_11088 ( P1_R1165_U583 , P1_R1165_U582 , P1_R1165_U581 );
nand NAND2_11089 ( P1_R1165_U584 , P1_R1165_U348 , P1_R1165_U56 );
nand NAND2_11090 ( P1_R1165_U585 , P1_R1165_U583 , P1_R1165_U333 );
nand NAND2_11091 ( P1_R1165_U586 , P1_R1165_U460 , P1_U3168 );
nand NAND2_11092 ( P1_R1165_U587 , P1_R1165_U74 , P1_R1165_U40 );
nand NAND2_11093 ( P1_R1165_U588 , P1_R1165_U587 , P1_R1165_U586 );
nand NAND2_11094 ( P1_R1165_U589 , P1_R1165_U349 , P1_R1165_U190 );
nand NAND2_11095 ( P1_R1165_U590 , P1_R1165_U251 , P1_R1165_U588 );
nand NAND2_11096 ( P1_R1165_U591 , P1_R1165_U451 , P1_U3169 );
nand NAND2_11097 ( P1_R1165_U592 , P1_R1165_U73 , P1_R1165_U38 );
nand NAND2_11098 ( P1_R1165_U593 , P1_R1165_U451 , P1_U3169 );
nand NAND2_11099 ( P1_R1165_U594 , P1_R1165_U73 , P1_R1165_U38 );
nand NAND2_11100 ( P1_R1165_U595 , P1_R1165_U594 , P1_R1165_U593 );
nand NAND2_11101 ( P1_R1165_U596 , P1_R1165_U191 , P1_R1165_U192 );
nand NAND2_11102 ( P1_R1165_U597 , P1_R1165_U364 , P1_R1165_U595 );
nand NAND2_11103 ( P1_R1165_U598 , P1_U3179 , P1_R1165_U16 );
nand NAND2_11104 ( P1_R1165_U599 , P1_U3209 , P1_R1165_U24 );
not NOT1_11105 ( P1_R1165_U600 , P1_R1165_U135 );
nand NAND2_11106 ( P1_R1165_U601 , P1_R1165_U63 , P1_R1165_U600 );
nand NAND2_11107 ( P1_R1165_U602 , P1_R1165_U135 , P1_R1165_U378 );
and AND2_11108 ( P1_R1150_U6 , P1_R1150_U184 , P1_R1150_U201 );
and AND2_11109 ( P1_R1150_U7 , P1_R1150_U203 , P1_R1150_U202 );
and AND2_11110 ( P1_R1150_U8 , P1_R1150_U179 , P1_R1150_U240 );
and AND2_11111 ( P1_R1150_U9 , P1_R1150_U242 , P1_R1150_U241 );
and AND2_11112 ( P1_R1150_U10 , P1_R1150_U259 , P1_R1150_U258 );
and AND2_11113 ( P1_R1150_U11 , P1_R1150_U285 , P1_R1150_U284 );
and AND2_11114 ( P1_R1150_U12 , P1_R1150_U383 , P1_R1150_U382 );
nand NAND2_11115 ( P1_R1150_U13 , P1_R1150_U340 , P1_R1150_U343 );
nand NAND2_11116 ( P1_R1150_U14 , P1_R1150_U329 , P1_R1150_U332 );
nand NAND2_11117 ( P1_R1150_U15 , P1_R1150_U318 , P1_R1150_U321 );
nand NAND2_11118 ( P1_R1150_U16 , P1_R1150_U310 , P1_R1150_U312 );
nand NAND3_11119 ( P1_R1150_U17 , P1_R1150_U156 , P1_R1150_U175 , P1_R1150_U348 );
nand NAND2_11120 ( P1_R1150_U18 , P1_R1150_U236 , P1_R1150_U238 );
nand NAND2_11121 ( P1_R1150_U19 , P1_R1150_U228 , P1_R1150_U231 );
nand NAND2_11122 ( P1_R1150_U20 , P1_R1150_U220 , P1_R1150_U222 );
nand NAND2_11123 ( P1_R1150_U21 , P1_R1150_U25 , P1_R1150_U346 );
not NOT1_11124 ( P1_R1150_U22 , P1_U3474 );
not NOT1_11125 ( P1_R1150_U23 , P1_U3459 );
not NOT1_11126 ( P1_R1150_U24 , P1_U3451 );
nand NAND2_11127 ( P1_R1150_U25 , P1_U3451 , P1_R1150_U93 );
not NOT1_11128 ( P1_R1150_U26 , P1_U3076 );
not NOT1_11129 ( P1_R1150_U27 , P1_U3462 );
not NOT1_11130 ( P1_R1150_U28 , P1_U3066 );
nand NAND2_11131 ( P1_R1150_U29 , P1_U3066 , P1_R1150_U23 );
not NOT1_11132 ( P1_R1150_U30 , P1_U3062 );
not NOT1_11133 ( P1_R1150_U31 , P1_U3471 );
not NOT1_11134 ( P1_R1150_U32 , P1_U3468 );
not NOT1_11135 ( P1_R1150_U33 , P1_U3465 );
not NOT1_11136 ( P1_R1150_U34 , P1_U3069 );
not NOT1_11137 ( P1_R1150_U35 , P1_U3065 );
not NOT1_11138 ( P1_R1150_U36 , P1_U3058 );
nand NAND2_11139 ( P1_R1150_U37 , P1_U3058 , P1_R1150_U33 );
not NOT1_11140 ( P1_R1150_U38 , P1_U3477 );
not NOT1_11141 ( P1_R1150_U39 , P1_U3068 );
nand NAND2_11142 ( P1_R1150_U40 , P1_U3068 , P1_R1150_U22 );
not NOT1_11143 ( P1_R1150_U41 , P1_U3082 );
not NOT1_11144 ( P1_R1150_U42 , P1_U3480 );
not NOT1_11145 ( P1_R1150_U43 , P1_U3081 );
nand NAND2_11146 ( P1_R1150_U44 , P1_R1150_U209 , P1_R1150_U208 );
nand NAND2_11147 ( P1_R1150_U45 , P1_R1150_U37 , P1_R1150_U224 );
nand NAND2_11148 ( P1_R1150_U46 , P1_R1150_U193 , P1_R1150_U192 );
not NOT1_11149 ( P1_R1150_U47 , P1_U4009 );
not NOT1_11150 ( P1_R1150_U48 , P1_U4013 );
not NOT1_11151 ( P1_R1150_U49 , P1_U3498 );
not NOT1_11152 ( P1_R1150_U50 , P1_U3486 );
not NOT1_11153 ( P1_R1150_U51 , P1_U3483 );
not NOT1_11154 ( P1_R1150_U52 , P1_U3061 );
not NOT1_11155 ( P1_R1150_U53 , P1_U3060 );
nand NAND2_11156 ( P1_R1150_U54 , P1_U3081 , P1_R1150_U42 );
not NOT1_11157 ( P1_R1150_U55 , P1_U3489 );
not NOT1_11158 ( P1_R1150_U56 , P1_U3070 );
not NOT1_11159 ( P1_R1150_U57 , P1_U3492 );
not NOT1_11160 ( P1_R1150_U58 , P1_U3078 );
not NOT1_11161 ( P1_R1150_U59 , P1_U3501 );
not NOT1_11162 ( P1_R1150_U60 , P1_U3495 );
not NOT1_11163 ( P1_R1150_U61 , P1_U3071 );
not NOT1_11164 ( P1_R1150_U62 , P1_U3072 );
not NOT1_11165 ( P1_R1150_U63 , P1_U3077 );
nand NAND2_11166 ( P1_R1150_U64 , P1_U3077 , P1_R1150_U60 );
not NOT1_11167 ( P1_R1150_U65 , P1_U3504 );
not NOT1_11168 ( P1_R1150_U66 , P1_U3067 );
nand NAND2_11169 ( P1_R1150_U67 , P1_R1150_U269 , P1_R1150_U268 );
not NOT1_11170 ( P1_R1150_U68 , P1_U3080 );
not NOT1_11171 ( P1_R1150_U69 , P1_U3509 );
not NOT1_11172 ( P1_R1150_U70 , P1_U3079 );
not NOT1_11173 ( P1_R1150_U71 , P1_U4015 );
not NOT1_11174 ( P1_R1150_U72 , P1_U3074 );
not NOT1_11175 ( P1_R1150_U73 , P1_U4012 );
not NOT1_11176 ( P1_R1150_U74 , P1_U4014 );
not NOT1_11177 ( P1_R1150_U75 , P1_U3064 );
not NOT1_11178 ( P1_R1150_U76 , P1_U3059 );
not NOT1_11179 ( P1_R1150_U77 , P1_U3073 );
nand NAND2_11180 ( P1_R1150_U78 , P1_U3073 , P1_R1150_U74 );
not NOT1_11181 ( P1_R1150_U79 , P1_U4011 );
not NOT1_11182 ( P1_R1150_U80 , P1_U3063 );
not NOT1_11183 ( P1_R1150_U81 , P1_U4010 );
not NOT1_11184 ( P1_R1150_U82 , P1_U3056 );
not NOT1_11185 ( P1_R1150_U83 , P1_U4008 );
not NOT1_11186 ( P1_R1150_U84 , P1_U3055 );
nand NAND2_11187 ( P1_R1150_U85 , P1_U3055 , P1_R1150_U47 );
not NOT1_11188 ( P1_R1150_U86 , P1_U3051 );
not NOT1_11189 ( P1_R1150_U87 , P1_U4007 );
not NOT1_11190 ( P1_R1150_U88 , P1_U3052 );
nand NAND2_11191 ( P1_R1150_U89 , P1_R1150_U299 , P1_R1150_U298 );
nand NAND2_11192 ( P1_R1150_U90 , P1_R1150_U78 , P1_R1150_U314 );
nand NAND2_11193 ( P1_R1150_U91 , P1_R1150_U64 , P1_R1150_U325 );
nand NAND2_11194 ( P1_R1150_U92 , P1_R1150_U54 , P1_R1150_U336 );
not NOT1_11195 ( P1_R1150_U93 , P1_U3075 );
nand NAND2_11196 ( P1_R1150_U94 , P1_R1150_U393 , P1_R1150_U392 );
nand NAND2_11197 ( P1_R1150_U95 , P1_R1150_U407 , P1_R1150_U406 );
nand NAND2_11198 ( P1_R1150_U96 , P1_R1150_U412 , P1_R1150_U411 );
nand NAND2_11199 ( P1_R1150_U97 , P1_R1150_U428 , P1_R1150_U427 );
nand NAND2_11200 ( P1_R1150_U98 , P1_R1150_U433 , P1_R1150_U432 );
nand NAND2_11201 ( P1_R1150_U99 , P1_R1150_U438 , P1_R1150_U437 );
nand NAND2_11202 ( P1_R1150_U100 , P1_R1150_U443 , P1_R1150_U442 );
nand NAND2_11203 ( P1_R1150_U101 , P1_R1150_U448 , P1_R1150_U447 );
nand NAND2_11204 ( P1_R1150_U102 , P1_R1150_U464 , P1_R1150_U463 );
nand NAND2_11205 ( P1_R1150_U103 , P1_R1150_U469 , P1_R1150_U468 );
nand NAND2_11206 ( P1_R1150_U104 , P1_R1150_U352 , P1_R1150_U351 );
nand NAND2_11207 ( P1_R1150_U105 , P1_R1150_U361 , P1_R1150_U360 );
nand NAND2_11208 ( P1_R1150_U106 , P1_R1150_U368 , P1_R1150_U367 );
nand NAND2_11209 ( P1_R1150_U107 , P1_R1150_U372 , P1_R1150_U371 );
nand NAND2_11210 ( P1_R1150_U108 , P1_R1150_U381 , P1_R1150_U380 );
nand NAND2_11211 ( P1_R1150_U109 , P1_R1150_U402 , P1_R1150_U401 );
nand NAND2_11212 ( P1_R1150_U110 , P1_R1150_U419 , P1_R1150_U418 );
nand NAND2_11213 ( P1_R1150_U111 , P1_R1150_U423 , P1_R1150_U422 );
nand NAND2_11214 ( P1_R1150_U112 , P1_R1150_U455 , P1_R1150_U454 );
nand NAND2_11215 ( P1_R1150_U113 , P1_R1150_U459 , P1_R1150_U458 );
nand NAND2_11216 ( P1_R1150_U114 , P1_R1150_U476 , P1_R1150_U475 );
and AND2_11217 ( P1_R1150_U115 , P1_R1150_U195 , P1_R1150_U183 );
and AND2_11218 ( P1_R1150_U116 , P1_R1150_U198 , P1_R1150_U199 );
and AND2_11219 ( P1_R1150_U117 , P1_R1150_U211 , P1_R1150_U185 );
and AND2_11220 ( P1_R1150_U118 , P1_R1150_U214 , P1_R1150_U215 );
and AND3_11221 ( P1_R1150_U119 , P1_R1150_U354 , P1_R1150_U353 , P1_R1150_U40 );
and AND2_11222 ( P1_R1150_U120 , P1_R1150_U357 , P1_R1150_U185 );
and AND2_11223 ( P1_R1150_U121 , P1_R1150_U230 , P1_R1150_U7 );
and AND2_11224 ( P1_R1150_U122 , P1_R1150_U364 , P1_R1150_U184 );
and AND3_11225 ( P1_R1150_U123 , P1_R1150_U374 , P1_R1150_U373 , P1_R1150_U29 );
and AND2_11226 ( P1_R1150_U124 , P1_R1150_U377 , P1_R1150_U183 );
and AND2_11227 ( P1_R1150_U125 , P1_R1150_U217 , P1_R1150_U8 );
and AND2_11228 ( P1_R1150_U126 , P1_R1150_U262 , P1_R1150_U180 );
and AND2_11229 ( P1_R1150_U127 , P1_R1150_U288 , P1_R1150_U181 );
and AND2_11230 ( P1_R1150_U128 , P1_R1150_U304 , P1_R1150_U305 );
and AND2_11231 ( P1_R1150_U129 , P1_R1150_U307 , P1_R1150_U386 );
and AND3_11232 ( P1_R1150_U130 , P1_R1150_U305 , P1_R1150_U304 , P1_R1150_U308 );
nand NAND2_11233 ( P1_R1150_U131 , P1_R1150_U390 , P1_R1150_U389 );
and AND3_11234 ( P1_R1150_U132 , P1_R1150_U395 , P1_R1150_U394 , P1_R1150_U85 );
and AND2_11235 ( P1_R1150_U133 , P1_R1150_U398 , P1_R1150_U182 );
nand NAND2_11236 ( P1_R1150_U134 , P1_R1150_U404 , P1_R1150_U403 );
nand NAND2_11237 ( P1_R1150_U135 , P1_R1150_U409 , P1_R1150_U408 );
and AND2_11238 ( P1_R1150_U136 , P1_R1150_U415 , P1_R1150_U181 );
nand NAND2_11239 ( P1_R1150_U137 , P1_R1150_U425 , P1_R1150_U424 );
nand NAND2_11240 ( P1_R1150_U138 , P1_R1150_U430 , P1_R1150_U429 );
nand NAND2_11241 ( P1_R1150_U139 , P1_R1150_U435 , P1_R1150_U434 );
nand NAND2_11242 ( P1_R1150_U140 , P1_R1150_U440 , P1_R1150_U439 );
nand NAND2_11243 ( P1_R1150_U141 , P1_R1150_U445 , P1_R1150_U444 );
and AND2_11244 ( P1_R1150_U142 , P1_R1150_U451 , P1_R1150_U180 );
nand NAND2_11245 ( P1_R1150_U143 , P1_R1150_U461 , P1_R1150_U460 );
nand NAND2_11246 ( P1_R1150_U144 , P1_R1150_U466 , P1_R1150_U465 );
and AND2_11247 ( P1_R1150_U145 , P1_R1150_U342 , P1_R1150_U9 );
and AND2_11248 ( P1_R1150_U146 , P1_R1150_U472 , P1_R1150_U179 );
and AND2_11249 ( P1_R1150_U147 , P1_R1150_U350 , P1_R1150_U349 );
nand NAND2_11250 ( P1_R1150_U148 , P1_R1150_U118 , P1_R1150_U212 );
and AND2_11251 ( P1_R1150_U149 , P1_R1150_U359 , P1_R1150_U358 );
and AND2_11252 ( P1_R1150_U150 , P1_R1150_U366 , P1_R1150_U365 );
and AND2_11253 ( P1_R1150_U151 , P1_R1150_U370 , P1_R1150_U369 );
nand NAND2_11254 ( P1_R1150_U152 , P1_R1150_U116 , P1_R1150_U196 );
and AND2_11255 ( P1_R1150_U153 , P1_R1150_U379 , P1_R1150_U378 );
not NOT1_11256 ( P1_R1150_U154 , P1_U4018 );
not NOT1_11257 ( P1_R1150_U155 , P1_U3053 );
and AND2_11258 ( P1_R1150_U156 , P1_R1150_U388 , P1_R1150_U387 );
nand NAND2_11259 ( P1_R1150_U157 , P1_R1150_U128 , P1_R1150_U302 );
and AND2_11260 ( P1_R1150_U158 , P1_R1150_U400 , P1_R1150_U399 );
nand NAND2_11261 ( P1_R1150_U159 , P1_R1150_U295 , P1_R1150_U294 );
nand NAND2_11262 ( P1_R1150_U160 , P1_R1150_U291 , P1_R1150_U290 );
and AND2_11263 ( P1_R1150_U161 , P1_R1150_U417 , P1_R1150_U416 );
and AND2_11264 ( P1_R1150_U162 , P1_R1150_U421 , P1_R1150_U420 );
nand NAND2_11265 ( P1_R1150_U163 , P1_R1150_U281 , P1_R1150_U280 );
nand NAND2_11266 ( P1_R1150_U164 , P1_R1150_U277 , P1_R1150_U276 );
not NOT1_11267 ( P1_R1150_U165 , P1_U3456 );
nand NAND2_11268 ( P1_R1150_U166 , P1_R1150_U273 , P1_R1150_U272 );
not NOT1_11269 ( P1_R1150_U167 , P1_U3507 );
nand NAND2_11270 ( P1_R1150_U168 , P1_R1150_U265 , P1_R1150_U264 );
and AND2_11271 ( P1_R1150_U169 , P1_R1150_U453 , P1_R1150_U452 );
and AND2_11272 ( P1_R1150_U170 , P1_R1150_U457 , P1_R1150_U456 );
nand NAND2_11273 ( P1_R1150_U171 , P1_R1150_U255 , P1_R1150_U254 );
nand NAND2_11274 ( P1_R1150_U172 , P1_R1150_U251 , P1_R1150_U250 );
nand NAND2_11275 ( P1_R1150_U173 , P1_R1150_U247 , P1_R1150_U246 );
and AND2_11276 ( P1_R1150_U174 , P1_R1150_U474 , P1_R1150_U473 );
nand NAND2_11277 ( P1_R1150_U175 , P1_R1150_U129 , P1_R1150_U157 );
not NOT1_11278 ( P1_R1150_U176 , P1_R1150_U85 );
not NOT1_11279 ( P1_R1150_U177 , P1_R1150_U29 );
not NOT1_11280 ( P1_R1150_U178 , P1_R1150_U40 );
nand NAND2_11281 ( P1_R1150_U179 , P1_U3483 , P1_R1150_U53 );
nand NAND2_11282 ( P1_R1150_U180 , P1_U3498 , P1_R1150_U62 );
nand NAND2_11283 ( P1_R1150_U181 , P1_U4013 , P1_R1150_U76 );
nand NAND2_11284 ( P1_R1150_U182 , P1_U4009 , P1_R1150_U84 );
nand NAND2_11285 ( P1_R1150_U183 , P1_U3459 , P1_R1150_U28 );
nand NAND2_11286 ( P1_R1150_U184 , P1_U3468 , P1_R1150_U35 );
nand NAND2_11287 ( P1_R1150_U185 , P1_U3474 , P1_R1150_U39 );
not NOT1_11288 ( P1_R1150_U186 , P1_R1150_U64 );
not NOT1_11289 ( P1_R1150_U187 , P1_R1150_U78 );
not NOT1_11290 ( P1_R1150_U188 , P1_R1150_U37 );
not NOT1_11291 ( P1_R1150_U189 , P1_R1150_U54 );
not NOT1_11292 ( P1_R1150_U190 , P1_R1150_U25 );
nand NAND2_11293 ( P1_R1150_U191 , P1_R1150_U190 , P1_R1150_U26 );
nand NAND2_11294 ( P1_R1150_U192 , P1_R1150_U191 , P1_R1150_U165 );
nand NAND2_11295 ( P1_R1150_U193 , P1_U3076 , P1_R1150_U25 );
not NOT1_11296 ( P1_R1150_U194 , P1_R1150_U46 );
nand NAND2_11297 ( P1_R1150_U195 , P1_U3462 , P1_R1150_U30 );
nand NAND2_11298 ( P1_R1150_U196 , P1_R1150_U115 , P1_R1150_U46 );
nand NAND2_11299 ( P1_R1150_U197 , P1_R1150_U30 , P1_R1150_U29 );
nand NAND2_11300 ( P1_R1150_U198 , P1_R1150_U197 , P1_R1150_U27 );
nand NAND2_11301 ( P1_R1150_U199 , P1_U3062 , P1_R1150_U177 );
not NOT1_11302 ( P1_R1150_U200 , P1_R1150_U152 );
nand NAND2_11303 ( P1_R1150_U201 , P1_U3471 , P1_R1150_U34 );
nand NAND2_11304 ( P1_R1150_U202 , P1_U3069 , P1_R1150_U31 );
nand NAND2_11305 ( P1_R1150_U203 , P1_U3065 , P1_R1150_U32 );
nand NAND2_11306 ( P1_R1150_U204 , P1_R1150_U188 , P1_R1150_U6 );
nand NAND2_11307 ( P1_R1150_U205 , P1_R1150_U7 , P1_R1150_U204 );
nand NAND2_11308 ( P1_R1150_U206 , P1_U3465 , P1_R1150_U36 );
nand NAND2_11309 ( P1_R1150_U207 , P1_U3471 , P1_R1150_U34 );
nand NAND3_11310 ( P1_R1150_U208 , P1_R1150_U206 , P1_R1150_U152 , P1_R1150_U6 );
nand NAND2_11311 ( P1_R1150_U209 , P1_R1150_U207 , P1_R1150_U205 );
not NOT1_11312 ( P1_R1150_U210 , P1_R1150_U44 );
nand NAND2_11313 ( P1_R1150_U211 , P1_U3477 , P1_R1150_U41 );
nand NAND2_11314 ( P1_R1150_U212 , P1_R1150_U117 , P1_R1150_U44 );
nand NAND2_11315 ( P1_R1150_U213 , P1_R1150_U41 , P1_R1150_U40 );
nand NAND2_11316 ( P1_R1150_U214 , P1_R1150_U213 , P1_R1150_U38 );
nand NAND2_11317 ( P1_R1150_U215 , P1_U3082 , P1_R1150_U178 );
not NOT1_11318 ( P1_R1150_U216 , P1_R1150_U148 );
nand NAND2_11319 ( P1_R1150_U217 , P1_U3480 , P1_R1150_U43 );
nand NAND2_11320 ( P1_R1150_U218 , P1_R1150_U217 , P1_R1150_U54 );
nand NAND2_11321 ( P1_R1150_U219 , P1_R1150_U210 , P1_R1150_U40 );
nand NAND2_11322 ( P1_R1150_U220 , P1_R1150_U120 , P1_R1150_U219 );
nand NAND2_11323 ( P1_R1150_U221 , P1_R1150_U44 , P1_R1150_U185 );
nand NAND2_11324 ( P1_R1150_U222 , P1_R1150_U119 , P1_R1150_U221 );
nand NAND2_11325 ( P1_R1150_U223 , P1_R1150_U40 , P1_R1150_U185 );
nand NAND2_11326 ( P1_R1150_U224 , P1_R1150_U206 , P1_R1150_U152 );
not NOT1_11327 ( P1_R1150_U225 , P1_R1150_U45 );
nand NAND2_11328 ( P1_R1150_U226 , P1_U3065 , P1_R1150_U32 );
nand NAND2_11329 ( P1_R1150_U227 , P1_R1150_U225 , P1_R1150_U226 );
nand NAND2_11330 ( P1_R1150_U228 , P1_R1150_U122 , P1_R1150_U227 );
nand NAND2_11331 ( P1_R1150_U229 , P1_R1150_U45 , P1_R1150_U184 );
nand NAND2_11332 ( P1_R1150_U230 , P1_U3471 , P1_R1150_U34 );
nand NAND2_11333 ( P1_R1150_U231 , P1_R1150_U121 , P1_R1150_U229 );
nand NAND2_11334 ( P1_R1150_U232 , P1_U3065 , P1_R1150_U32 );
nand NAND2_11335 ( P1_R1150_U233 , P1_R1150_U184 , P1_R1150_U232 );
nand NAND2_11336 ( P1_R1150_U234 , P1_R1150_U206 , P1_R1150_U37 );
nand NAND2_11337 ( P1_R1150_U235 , P1_R1150_U194 , P1_R1150_U29 );
nand NAND2_11338 ( P1_R1150_U236 , P1_R1150_U124 , P1_R1150_U235 );
nand NAND2_11339 ( P1_R1150_U237 , P1_R1150_U46 , P1_R1150_U183 );
nand NAND2_11340 ( P1_R1150_U238 , P1_R1150_U123 , P1_R1150_U237 );
nand NAND2_11341 ( P1_R1150_U239 , P1_R1150_U29 , P1_R1150_U183 );
nand NAND2_11342 ( P1_R1150_U240 , P1_U3486 , P1_R1150_U52 );
nand NAND2_11343 ( P1_R1150_U241 , P1_U3061 , P1_R1150_U50 );
nand NAND2_11344 ( P1_R1150_U242 , P1_U3060 , P1_R1150_U51 );
nand NAND2_11345 ( P1_R1150_U243 , P1_R1150_U189 , P1_R1150_U8 );
nand NAND2_11346 ( P1_R1150_U244 , P1_R1150_U9 , P1_R1150_U243 );
nand NAND2_11347 ( P1_R1150_U245 , P1_U3486 , P1_R1150_U52 );
nand NAND2_11348 ( P1_R1150_U246 , P1_R1150_U125 , P1_R1150_U148 );
nand NAND2_11349 ( P1_R1150_U247 , P1_R1150_U245 , P1_R1150_U244 );
not NOT1_11350 ( P1_R1150_U248 , P1_R1150_U173 );
nand NAND2_11351 ( P1_R1150_U249 , P1_U3489 , P1_R1150_U56 );
nand NAND2_11352 ( P1_R1150_U250 , P1_R1150_U249 , P1_R1150_U173 );
nand NAND2_11353 ( P1_R1150_U251 , P1_U3070 , P1_R1150_U55 );
not NOT1_11354 ( P1_R1150_U252 , P1_R1150_U172 );
nand NAND2_11355 ( P1_R1150_U253 , P1_U3492 , P1_R1150_U58 );
nand NAND2_11356 ( P1_R1150_U254 , P1_R1150_U253 , P1_R1150_U172 );
nand NAND2_11357 ( P1_R1150_U255 , P1_U3078 , P1_R1150_U57 );
not NOT1_11358 ( P1_R1150_U256 , P1_R1150_U171 );
nand NAND2_11359 ( P1_R1150_U257 , P1_U3501 , P1_R1150_U61 );
nand NAND2_11360 ( P1_R1150_U258 , P1_U3071 , P1_R1150_U59 );
nand NAND2_11361 ( P1_R1150_U259 , P1_U3072 , P1_R1150_U49 );
nand NAND2_11362 ( P1_R1150_U260 , P1_R1150_U186 , P1_R1150_U180 );
nand NAND2_11363 ( P1_R1150_U261 , P1_R1150_U10 , P1_R1150_U260 );
nand NAND2_11364 ( P1_R1150_U262 , P1_U3495 , P1_R1150_U63 );
nand NAND2_11365 ( P1_R1150_U263 , P1_U3501 , P1_R1150_U61 );
nand NAND3_11366 ( P1_R1150_U264 , P1_R1150_U171 , P1_R1150_U126 , P1_R1150_U257 );
nand NAND2_11367 ( P1_R1150_U265 , P1_R1150_U263 , P1_R1150_U261 );
not NOT1_11368 ( P1_R1150_U266 , P1_R1150_U168 );
nand NAND2_11369 ( P1_R1150_U267 , P1_U3504 , P1_R1150_U66 );
nand NAND2_11370 ( P1_R1150_U268 , P1_R1150_U267 , P1_R1150_U168 );
nand NAND2_11371 ( P1_R1150_U269 , P1_U3067 , P1_R1150_U65 );
not NOT1_11372 ( P1_R1150_U270 , P1_R1150_U67 );
nand NAND2_11373 ( P1_R1150_U271 , P1_R1150_U270 , P1_R1150_U68 );
nand NAND2_11374 ( P1_R1150_U272 , P1_R1150_U271 , P1_R1150_U167 );
nand NAND2_11375 ( P1_R1150_U273 , P1_U3080 , P1_R1150_U67 );
not NOT1_11376 ( P1_R1150_U274 , P1_R1150_U166 );
nand NAND2_11377 ( P1_R1150_U275 , P1_U3509 , P1_R1150_U70 );
nand NAND2_11378 ( P1_R1150_U276 , P1_R1150_U275 , P1_R1150_U166 );
nand NAND2_11379 ( P1_R1150_U277 , P1_U3079 , P1_R1150_U69 );
not NOT1_11380 ( P1_R1150_U278 , P1_R1150_U164 );
nand NAND2_11381 ( P1_R1150_U279 , P1_U4015 , P1_R1150_U72 );
nand NAND2_11382 ( P1_R1150_U280 , P1_R1150_U279 , P1_R1150_U164 );
nand NAND2_11383 ( P1_R1150_U281 , P1_U3074 , P1_R1150_U71 );
not NOT1_11384 ( P1_R1150_U282 , P1_R1150_U163 );
nand NAND2_11385 ( P1_R1150_U283 , P1_U4012 , P1_R1150_U75 );
nand NAND2_11386 ( P1_R1150_U284 , P1_U3064 , P1_R1150_U73 );
nand NAND2_11387 ( P1_R1150_U285 , P1_U3059 , P1_R1150_U48 );
nand NAND2_11388 ( P1_R1150_U286 , P1_R1150_U187 , P1_R1150_U181 );
nand NAND2_11389 ( P1_R1150_U287 , P1_R1150_U11 , P1_R1150_U286 );
nand NAND2_11390 ( P1_R1150_U288 , P1_U4014 , P1_R1150_U77 );
nand NAND2_11391 ( P1_R1150_U289 , P1_U4012 , P1_R1150_U75 );
nand NAND3_11392 ( P1_R1150_U290 , P1_R1150_U163 , P1_R1150_U127 , P1_R1150_U283 );
nand NAND2_11393 ( P1_R1150_U291 , P1_R1150_U289 , P1_R1150_U287 );
not NOT1_11394 ( P1_R1150_U292 , P1_R1150_U160 );
nand NAND2_11395 ( P1_R1150_U293 , P1_U4011 , P1_R1150_U80 );
nand NAND2_11396 ( P1_R1150_U294 , P1_R1150_U293 , P1_R1150_U160 );
nand NAND2_11397 ( P1_R1150_U295 , P1_U3063 , P1_R1150_U79 );
not NOT1_11398 ( P1_R1150_U296 , P1_R1150_U159 );
nand NAND2_11399 ( P1_R1150_U297 , P1_U4010 , P1_R1150_U82 );
nand NAND2_11400 ( P1_R1150_U298 , P1_R1150_U297 , P1_R1150_U159 );
nand NAND2_11401 ( P1_R1150_U299 , P1_U3056 , P1_R1150_U81 );
not NOT1_11402 ( P1_R1150_U300 , P1_R1150_U89 );
nand NAND2_11403 ( P1_R1150_U301 , P1_U4008 , P1_R1150_U86 );
nand NAND3_11404 ( P1_R1150_U302 , P1_R1150_U89 , P1_R1150_U182 , P1_R1150_U301 );
nand NAND2_11405 ( P1_R1150_U303 , P1_R1150_U86 , P1_R1150_U85 );
nand NAND2_11406 ( P1_R1150_U304 , P1_R1150_U303 , P1_R1150_U83 );
nand NAND2_11407 ( P1_R1150_U305 , P1_U3051 , P1_R1150_U176 );
not NOT1_11408 ( P1_R1150_U306 , P1_R1150_U157 );
nand NAND2_11409 ( P1_R1150_U307 , P1_U4007 , P1_R1150_U88 );
nand NAND2_11410 ( P1_R1150_U308 , P1_U3052 , P1_R1150_U87 );
nand NAND2_11411 ( P1_R1150_U309 , P1_R1150_U300 , P1_R1150_U85 );
nand NAND2_11412 ( P1_R1150_U310 , P1_R1150_U133 , P1_R1150_U309 );
nand NAND2_11413 ( P1_R1150_U311 , P1_R1150_U89 , P1_R1150_U182 );
nand NAND2_11414 ( P1_R1150_U312 , P1_R1150_U132 , P1_R1150_U311 );
nand NAND2_11415 ( P1_R1150_U313 , P1_R1150_U85 , P1_R1150_U182 );
nand NAND2_11416 ( P1_R1150_U314 , P1_R1150_U288 , P1_R1150_U163 );
not NOT1_11417 ( P1_R1150_U315 , P1_R1150_U90 );
nand NAND2_11418 ( P1_R1150_U316 , P1_U3059 , P1_R1150_U48 );
nand NAND2_11419 ( P1_R1150_U317 , P1_R1150_U315 , P1_R1150_U316 );
nand NAND2_11420 ( P1_R1150_U318 , P1_R1150_U136 , P1_R1150_U317 );
nand NAND2_11421 ( P1_R1150_U319 , P1_R1150_U90 , P1_R1150_U181 );
nand NAND2_11422 ( P1_R1150_U320 , P1_U4012 , P1_R1150_U75 );
nand NAND3_11423 ( P1_R1150_U321 , P1_R1150_U320 , P1_R1150_U319 , P1_R1150_U11 );
nand NAND2_11424 ( P1_R1150_U322 , P1_U3059 , P1_R1150_U48 );
nand NAND2_11425 ( P1_R1150_U323 , P1_R1150_U181 , P1_R1150_U322 );
nand NAND2_11426 ( P1_R1150_U324 , P1_R1150_U288 , P1_R1150_U78 );
nand NAND2_11427 ( P1_R1150_U325 , P1_R1150_U262 , P1_R1150_U171 );
not NOT1_11428 ( P1_R1150_U326 , P1_R1150_U91 );
nand NAND2_11429 ( P1_R1150_U327 , P1_U3072 , P1_R1150_U49 );
nand NAND2_11430 ( P1_R1150_U328 , P1_R1150_U326 , P1_R1150_U327 );
nand NAND2_11431 ( P1_R1150_U329 , P1_R1150_U142 , P1_R1150_U328 );
nand NAND2_11432 ( P1_R1150_U330 , P1_R1150_U91 , P1_R1150_U180 );
nand NAND2_11433 ( P1_R1150_U331 , P1_U3501 , P1_R1150_U61 );
nand NAND3_11434 ( P1_R1150_U332 , P1_R1150_U331 , P1_R1150_U330 , P1_R1150_U10 );
nand NAND2_11435 ( P1_R1150_U333 , P1_U3072 , P1_R1150_U49 );
nand NAND2_11436 ( P1_R1150_U334 , P1_R1150_U180 , P1_R1150_U333 );
nand NAND2_11437 ( P1_R1150_U335 , P1_R1150_U262 , P1_R1150_U64 );
nand NAND2_11438 ( P1_R1150_U336 , P1_R1150_U217 , P1_R1150_U148 );
not NOT1_11439 ( P1_R1150_U337 , P1_R1150_U92 );
nand NAND2_11440 ( P1_R1150_U338 , P1_U3060 , P1_R1150_U51 );
nand NAND2_11441 ( P1_R1150_U339 , P1_R1150_U337 , P1_R1150_U338 );
nand NAND2_11442 ( P1_R1150_U340 , P1_R1150_U146 , P1_R1150_U339 );
nand NAND2_11443 ( P1_R1150_U341 , P1_R1150_U92 , P1_R1150_U179 );
nand NAND2_11444 ( P1_R1150_U342 , P1_U3486 , P1_R1150_U52 );
nand NAND2_11445 ( P1_R1150_U343 , P1_R1150_U145 , P1_R1150_U341 );
nand NAND2_11446 ( P1_R1150_U344 , P1_U3060 , P1_R1150_U51 );
nand NAND2_11447 ( P1_R1150_U345 , P1_R1150_U179 , P1_R1150_U344 );
nand NAND2_11448 ( P1_R1150_U346 , P1_U3075 , P1_R1150_U24 );
nand NAND3_11449 ( P1_R1150_U347 , P1_R1150_U89 , P1_R1150_U182 , P1_R1150_U301 );
nand NAND3_11450 ( P1_R1150_U348 , P1_R1150_U12 , P1_R1150_U347 , P1_R1150_U130 );
nand NAND2_11451 ( P1_R1150_U349 , P1_U3480 , P1_R1150_U43 );
nand NAND2_11452 ( P1_R1150_U350 , P1_U3081 , P1_R1150_U42 );
nand NAND2_11453 ( P1_R1150_U351 , P1_R1150_U218 , P1_R1150_U148 );
nand NAND2_11454 ( P1_R1150_U352 , P1_R1150_U216 , P1_R1150_U147 );
nand NAND2_11455 ( P1_R1150_U353 , P1_U3477 , P1_R1150_U41 );
nand NAND2_11456 ( P1_R1150_U354 , P1_U3082 , P1_R1150_U38 );
nand NAND2_11457 ( P1_R1150_U355 , P1_U3477 , P1_R1150_U41 );
nand NAND2_11458 ( P1_R1150_U356 , P1_U3082 , P1_R1150_U38 );
nand NAND2_11459 ( P1_R1150_U357 , P1_R1150_U356 , P1_R1150_U355 );
nand NAND2_11460 ( P1_R1150_U358 , P1_U3474 , P1_R1150_U39 );
nand NAND2_11461 ( P1_R1150_U359 , P1_U3068 , P1_R1150_U22 );
nand NAND2_11462 ( P1_R1150_U360 , P1_R1150_U223 , P1_R1150_U44 );
nand NAND2_11463 ( P1_R1150_U361 , P1_R1150_U149 , P1_R1150_U210 );
nand NAND2_11464 ( P1_R1150_U362 , P1_U3471 , P1_R1150_U34 );
nand NAND2_11465 ( P1_R1150_U363 , P1_U3069 , P1_R1150_U31 );
nand NAND2_11466 ( P1_R1150_U364 , P1_R1150_U363 , P1_R1150_U362 );
nand NAND2_11467 ( P1_R1150_U365 , P1_U3468 , P1_R1150_U35 );
nand NAND2_11468 ( P1_R1150_U366 , P1_U3065 , P1_R1150_U32 );
nand NAND2_11469 ( P1_R1150_U367 , P1_R1150_U233 , P1_R1150_U45 );
nand NAND2_11470 ( P1_R1150_U368 , P1_R1150_U150 , P1_R1150_U225 );
nand NAND2_11471 ( P1_R1150_U369 , P1_U3465 , P1_R1150_U36 );
nand NAND2_11472 ( P1_R1150_U370 , P1_U3058 , P1_R1150_U33 );
nand NAND2_11473 ( P1_R1150_U371 , P1_R1150_U234 , P1_R1150_U152 );
nand NAND2_11474 ( P1_R1150_U372 , P1_R1150_U200 , P1_R1150_U151 );
nand NAND2_11475 ( P1_R1150_U373 , P1_U3462 , P1_R1150_U30 );
nand NAND2_11476 ( P1_R1150_U374 , P1_U3062 , P1_R1150_U27 );
nand NAND2_11477 ( P1_R1150_U375 , P1_U3462 , P1_R1150_U30 );
nand NAND2_11478 ( P1_R1150_U376 , P1_U3062 , P1_R1150_U27 );
nand NAND2_11479 ( P1_R1150_U377 , P1_R1150_U376 , P1_R1150_U375 );
nand NAND2_11480 ( P1_R1150_U378 , P1_U3459 , P1_R1150_U28 );
nand NAND2_11481 ( P1_R1150_U379 , P1_U3066 , P1_R1150_U23 );
nand NAND2_11482 ( P1_R1150_U380 , P1_R1150_U239 , P1_R1150_U46 );
nand NAND2_11483 ( P1_R1150_U381 , P1_R1150_U153 , P1_R1150_U194 );
nand NAND2_11484 ( P1_R1150_U382 , P1_U4018 , P1_R1150_U155 );
nand NAND2_11485 ( P1_R1150_U383 , P1_U3053 , P1_R1150_U154 );
nand NAND2_11486 ( P1_R1150_U384 , P1_U4018 , P1_R1150_U155 );
nand NAND2_11487 ( P1_R1150_U385 , P1_U3053 , P1_R1150_U154 );
nand NAND2_11488 ( P1_R1150_U386 , P1_R1150_U385 , P1_R1150_U384 );
nand NAND3_11489 ( P1_R1150_U387 , P1_U3052 , P1_R1150_U386 , P1_R1150_U87 );
nand NAND3_11490 ( P1_R1150_U388 , P1_R1150_U12 , P1_R1150_U88 , P1_U4007 );
nand NAND2_11491 ( P1_R1150_U389 , P1_U4007 , P1_R1150_U88 );
nand NAND2_11492 ( P1_R1150_U390 , P1_U3052 , P1_R1150_U87 );
not NOT1_11493 ( P1_R1150_U391 , P1_R1150_U131 );
nand NAND2_11494 ( P1_R1150_U392 , P1_R1150_U306 , P1_R1150_U391 );
nand NAND2_11495 ( P1_R1150_U393 , P1_R1150_U131 , P1_R1150_U157 );
nand NAND2_11496 ( P1_R1150_U394 , P1_U4008 , P1_R1150_U86 );
nand NAND2_11497 ( P1_R1150_U395 , P1_U3051 , P1_R1150_U83 );
nand NAND2_11498 ( P1_R1150_U396 , P1_U4008 , P1_R1150_U86 );
nand NAND2_11499 ( P1_R1150_U397 , P1_U3051 , P1_R1150_U83 );
nand NAND2_11500 ( P1_R1150_U398 , P1_R1150_U397 , P1_R1150_U396 );
nand NAND2_11501 ( P1_R1150_U399 , P1_U4009 , P1_R1150_U84 );
nand NAND2_11502 ( P1_R1150_U400 , P1_U3055 , P1_R1150_U47 );
nand NAND2_11503 ( P1_R1150_U401 , P1_R1150_U313 , P1_R1150_U89 );
nand NAND2_11504 ( P1_R1150_U402 , P1_R1150_U158 , P1_R1150_U300 );
nand NAND2_11505 ( P1_R1150_U403 , P1_U4010 , P1_R1150_U82 );
nand NAND2_11506 ( P1_R1150_U404 , P1_U3056 , P1_R1150_U81 );
not NOT1_11507 ( P1_R1150_U405 , P1_R1150_U134 );
nand NAND2_11508 ( P1_R1150_U406 , P1_R1150_U296 , P1_R1150_U405 );
nand NAND2_11509 ( P1_R1150_U407 , P1_R1150_U134 , P1_R1150_U159 );
nand NAND2_11510 ( P1_R1150_U408 , P1_U4011 , P1_R1150_U80 );
nand NAND2_11511 ( P1_R1150_U409 , P1_U3063 , P1_R1150_U79 );
not NOT1_11512 ( P1_R1150_U410 , P1_R1150_U135 );
nand NAND2_11513 ( P1_R1150_U411 , P1_R1150_U292 , P1_R1150_U410 );
nand NAND2_11514 ( P1_R1150_U412 , P1_R1150_U135 , P1_R1150_U160 );
nand NAND2_11515 ( P1_R1150_U413 , P1_U4012 , P1_R1150_U75 );
nand NAND2_11516 ( P1_R1150_U414 , P1_U3064 , P1_R1150_U73 );
nand NAND2_11517 ( P1_R1150_U415 , P1_R1150_U414 , P1_R1150_U413 );
nand NAND2_11518 ( P1_R1150_U416 , P1_U4013 , P1_R1150_U76 );
nand NAND2_11519 ( P1_R1150_U417 , P1_U3059 , P1_R1150_U48 );
nand NAND2_11520 ( P1_R1150_U418 , P1_R1150_U323 , P1_R1150_U90 );
nand NAND2_11521 ( P1_R1150_U419 , P1_R1150_U161 , P1_R1150_U315 );
nand NAND2_11522 ( P1_R1150_U420 , P1_U4014 , P1_R1150_U77 );
nand NAND2_11523 ( P1_R1150_U421 , P1_U3073 , P1_R1150_U74 );
nand NAND2_11524 ( P1_R1150_U422 , P1_R1150_U324 , P1_R1150_U163 );
nand NAND2_11525 ( P1_R1150_U423 , P1_R1150_U282 , P1_R1150_U162 );
nand NAND2_11526 ( P1_R1150_U424 , P1_U4015 , P1_R1150_U72 );
nand NAND2_11527 ( P1_R1150_U425 , P1_U3074 , P1_R1150_U71 );
not NOT1_11528 ( P1_R1150_U426 , P1_R1150_U137 );
nand NAND2_11529 ( P1_R1150_U427 , P1_R1150_U278 , P1_R1150_U426 );
nand NAND2_11530 ( P1_R1150_U428 , P1_R1150_U137 , P1_R1150_U164 );
nand NAND2_11531 ( P1_R1150_U429 , P1_U3456 , P1_R1150_U26 );
nand NAND2_11532 ( P1_R1150_U430 , P1_U3076 , P1_R1150_U165 );
not NOT1_11533 ( P1_R1150_U431 , P1_R1150_U138 );
nand NAND2_11534 ( P1_R1150_U432 , P1_R1150_U431 , P1_R1150_U190 );
nand NAND2_11535 ( P1_R1150_U433 , P1_R1150_U138 , P1_R1150_U25 );
nand NAND2_11536 ( P1_R1150_U434 , P1_U3509 , P1_R1150_U70 );
nand NAND2_11537 ( P1_R1150_U435 , P1_U3079 , P1_R1150_U69 );
not NOT1_11538 ( P1_R1150_U436 , P1_R1150_U139 );
nand NAND2_11539 ( P1_R1150_U437 , P1_R1150_U274 , P1_R1150_U436 );
nand NAND2_11540 ( P1_R1150_U438 , P1_R1150_U139 , P1_R1150_U166 );
nand NAND2_11541 ( P1_R1150_U439 , P1_U3507 , P1_R1150_U68 );
nand NAND2_11542 ( P1_R1150_U440 , P1_U3080 , P1_R1150_U167 );
not NOT1_11543 ( P1_R1150_U441 , P1_R1150_U140 );
nand NAND2_11544 ( P1_R1150_U442 , P1_R1150_U441 , P1_R1150_U270 );
nand NAND2_11545 ( P1_R1150_U443 , P1_R1150_U140 , P1_R1150_U67 );
nand NAND2_11546 ( P1_R1150_U444 , P1_U3504 , P1_R1150_U66 );
nand NAND2_11547 ( P1_R1150_U445 , P1_U3067 , P1_R1150_U65 );
not NOT1_11548 ( P1_R1150_U446 , P1_R1150_U141 );
nand NAND2_11549 ( P1_R1150_U447 , P1_R1150_U266 , P1_R1150_U446 );
nand NAND2_11550 ( P1_R1150_U448 , P1_R1150_U141 , P1_R1150_U168 );
nand NAND2_11551 ( P1_R1150_U449 , P1_U3501 , P1_R1150_U61 );
nand NAND2_11552 ( P1_R1150_U450 , P1_U3071 , P1_R1150_U59 );
nand NAND2_11553 ( P1_R1150_U451 , P1_R1150_U450 , P1_R1150_U449 );
nand NAND2_11554 ( P1_R1150_U452 , P1_U3498 , P1_R1150_U62 );
nand NAND2_11555 ( P1_R1150_U453 , P1_U3072 , P1_R1150_U49 );
nand NAND2_11556 ( P1_R1150_U454 , P1_R1150_U334 , P1_R1150_U91 );
nand NAND2_11557 ( P1_R1150_U455 , P1_R1150_U169 , P1_R1150_U326 );
nand NAND2_11558 ( P1_R1150_U456 , P1_U3495 , P1_R1150_U63 );
nand NAND2_11559 ( P1_R1150_U457 , P1_U3077 , P1_R1150_U60 );
nand NAND2_11560 ( P1_R1150_U458 , P1_R1150_U335 , P1_R1150_U171 );
nand NAND2_11561 ( P1_R1150_U459 , P1_R1150_U256 , P1_R1150_U170 );
nand NAND2_11562 ( P1_R1150_U460 , P1_U3492 , P1_R1150_U58 );
nand NAND2_11563 ( P1_R1150_U461 , P1_U3078 , P1_R1150_U57 );
not NOT1_11564 ( P1_R1150_U462 , P1_R1150_U143 );
nand NAND2_11565 ( P1_R1150_U463 , P1_R1150_U252 , P1_R1150_U462 );
nand NAND2_11566 ( P1_R1150_U464 , P1_R1150_U143 , P1_R1150_U172 );
nand NAND2_11567 ( P1_R1150_U465 , P1_U3489 , P1_R1150_U56 );
nand NAND2_11568 ( P1_R1150_U466 , P1_U3070 , P1_R1150_U55 );
not NOT1_11569 ( P1_R1150_U467 , P1_R1150_U144 );
nand NAND2_11570 ( P1_R1150_U468 , P1_R1150_U248 , P1_R1150_U467 );
nand NAND2_11571 ( P1_R1150_U469 , P1_R1150_U144 , P1_R1150_U173 );
nand NAND2_11572 ( P1_R1150_U470 , P1_U3486 , P1_R1150_U52 );
nand NAND2_11573 ( P1_R1150_U471 , P1_U3061 , P1_R1150_U50 );
nand NAND2_11574 ( P1_R1150_U472 , P1_R1150_U471 , P1_R1150_U470 );
nand NAND2_11575 ( P1_R1150_U473 , P1_U3483 , P1_R1150_U53 );
nand NAND2_11576 ( P1_R1150_U474 , P1_U3060 , P1_R1150_U51 );
nand NAND2_11577 ( P1_R1150_U475 , P1_R1150_U345 , P1_R1150_U92 );
nand NAND2_11578 ( P1_R1150_U476 , P1_R1150_U174 , P1_R1150_U337 );
and AND2_11579 ( P1_R1192_U6 , P1_R1192_U184 , P1_R1192_U201 );
and AND2_11580 ( P1_R1192_U7 , P1_R1192_U203 , P1_R1192_U202 );
and AND2_11581 ( P1_R1192_U8 , P1_R1192_U179 , P1_R1192_U240 );
and AND2_11582 ( P1_R1192_U9 , P1_R1192_U242 , P1_R1192_U241 );
and AND2_11583 ( P1_R1192_U10 , P1_R1192_U259 , P1_R1192_U258 );
and AND2_11584 ( P1_R1192_U11 , P1_R1192_U285 , P1_R1192_U284 );
and AND2_11585 ( P1_R1192_U12 , P1_R1192_U383 , P1_R1192_U382 );
nand NAND2_11586 ( P1_R1192_U13 , P1_R1192_U340 , P1_R1192_U343 );
nand NAND2_11587 ( P1_R1192_U14 , P1_R1192_U329 , P1_R1192_U332 );
nand NAND2_11588 ( P1_R1192_U15 , P1_R1192_U318 , P1_R1192_U321 );
nand NAND2_11589 ( P1_R1192_U16 , P1_R1192_U310 , P1_R1192_U312 );
nand NAND3_11590 ( P1_R1192_U17 , P1_R1192_U156 , P1_R1192_U175 , P1_R1192_U348 );
nand NAND2_11591 ( P1_R1192_U18 , P1_R1192_U236 , P1_R1192_U238 );
nand NAND2_11592 ( P1_R1192_U19 , P1_R1192_U228 , P1_R1192_U231 );
nand NAND2_11593 ( P1_R1192_U20 , P1_R1192_U220 , P1_R1192_U222 );
nand NAND2_11594 ( P1_R1192_U21 , P1_R1192_U25 , P1_R1192_U346 );
not NOT1_11595 ( P1_R1192_U22 , P1_U3474 );
not NOT1_11596 ( P1_R1192_U23 , P1_U3459 );
not NOT1_11597 ( P1_R1192_U24 , P1_U3451 );
nand NAND2_11598 ( P1_R1192_U25 , P1_U3451 , P1_R1192_U93 );
not NOT1_11599 ( P1_R1192_U26 , P1_U3076 );
not NOT1_11600 ( P1_R1192_U27 , P1_U3462 );
not NOT1_11601 ( P1_R1192_U28 , P1_U3066 );
nand NAND2_11602 ( P1_R1192_U29 , P1_U3066 , P1_R1192_U23 );
not NOT1_11603 ( P1_R1192_U30 , P1_U3062 );
not NOT1_11604 ( P1_R1192_U31 , P1_U3471 );
not NOT1_11605 ( P1_R1192_U32 , P1_U3468 );
not NOT1_11606 ( P1_R1192_U33 , P1_U3465 );
not NOT1_11607 ( P1_R1192_U34 , P1_U3069 );
not NOT1_11608 ( P1_R1192_U35 , P1_U3065 );
not NOT1_11609 ( P1_R1192_U36 , P1_U3058 );
nand NAND2_11610 ( P1_R1192_U37 , P1_U3058 , P1_R1192_U33 );
not NOT1_11611 ( P1_R1192_U38 , P1_U3477 );
not NOT1_11612 ( P1_R1192_U39 , P1_U3068 );
nand NAND2_11613 ( P1_R1192_U40 , P1_U3068 , P1_R1192_U22 );
not NOT1_11614 ( P1_R1192_U41 , P1_U3082 );
not NOT1_11615 ( P1_R1192_U42 , P1_U3480 );
not NOT1_11616 ( P1_R1192_U43 , P1_U3081 );
nand NAND2_11617 ( P1_R1192_U44 , P1_R1192_U209 , P1_R1192_U208 );
nand NAND2_11618 ( P1_R1192_U45 , P1_R1192_U37 , P1_R1192_U224 );
nand NAND2_11619 ( P1_R1192_U46 , P1_R1192_U193 , P1_R1192_U192 );
not NOT1_11620 ( P1_R1192_U47 , P1_U4009 );
not NOT1_11621 ( P1_R1192_U48 , P1_U4013 );
not NOT1_11622 ( P1_R1192_U49 , P1_U3498 );
not NOT1_11623 ( P1_R1192_U50 , P1_U3486 );
not NOT1_11624 ( P1_R1192_U51 , P1_U3483 );
not NOT1_11625 ( P1_R1192_U52 , P1_U3061 );
not NOT1_11626 ( P1_R1192_U53 , P1_U3060 );
nand NAND2_11627 ( P1_R1192_U54 , P1_U3081 , P1_R1192_U42 );
not NOT1_11628 ( P1_R1192_U55 , P1_U3489 );
not NOT1_11629 ( P1_R1192_U56 , P1_U3070 );
not NOT1_11630 ( P1_R1192_U57 , P1_U3492 );
not NOT1_11631 ( P1_R1192_U58 , P1_U3078 );
not NOT1_11632 ( P1_R1192_U59 , P1_U3501 );
not NOT1_11633 ( P1_R1192_U60 , P1_U3495 );
not NOT1_11634 ( P1_R1192_U61 , P1_U3071 );
not NOT1_11635 ( P1_R1192_U62 , P1_U3072 );
not NOT1_11636 ( P1_R1192_U63 , P1_U3077 );
nand NAND2_11637 ( P1_R1192_U64 , P1_U3077 , P1_R1192_U60 );
not NOT1_11638 ( P1_R1192_U65 , P1_U3504 );
not NOT1_11639 ( P1_R1192_U66 , P1_U3067 );
nand NAND2_11640 ( P1_R1192_U67 , P1_R1192_U269 , P1_R1192_U268 );
not NOT1_11641 ( P1_R1192_U68 , P1_U3080 );
not NOT1_11642 ( P1_R1192_U69 , P1_U3509 );
not NOT1_11643 ( P1_R1192_U70 , P1_U3079 );
not NOT1_11644 ( P1_R1192_U71 , P1_U4015 );
not NOT1_11645 ( P1_R1192_U72 , P1_U3074 );
not NOT1_11646 ( P1_R1192_U73 , P1_U4012 );
not NOT1_11647 ( P1_R1192_U74 , P1_U4014 );
not NOT1_11648 ( P1_R1192_U75 , P1_U3064 );
not NOT1_11649 ( P1_R1192_U76 , P1_U3059 );
not NOT1_11650 ( P1_R1192_U77 , P1_U3073 );
nand NAND2_11651 ( P1_R1192_U78 , P1_U3073 , P1_R1192_U74 );
not NOT1_11652 ( P1_R1192_U79 , P1_U4011 );
not NOT1_11653 ( P1_R1192_U80 , P1_U3063 );
not NOT1_11654 ( P1_R1192_U81 , P1_U4010 );
not NOT1_11655 ( P1_R1192_U82 , P1_U3056 );
not NOT1_11656 ( P1_R1192_U83 , P1_U4008 );
not NOT1_11657 ( P1_R1192_U84 , P1_U3055 );
nand NAND2_11658 ( P1_R1192_U85 , P1_U3055 , P1_R1192_U47 );
not NOT1_11659 ( P1_R1192_U86 , P1_U3051 );
not NOT1_11660 ( P1_R1192_U87 , P1_U4007 );
not NOT1_11661 ( P1_R1192_U88 , P1_U3052 );
nand NAND2_11662 ( P1_R1192_U89 , P1_R1192_U299 , P1_R1192_U298 );
nand NAND2_11663 ( P1_R1192_U90 , P1_R1192_U78 , P1_R1192_U314 );
nand NAND2_11664 ( P1_R1192_U91 , P1_R1192_U64 , P1_R1192_U325 );
nand NAND2_11665 ( P1_R1192_U92 , P1_R1192_U54 , P1_R1192_U336 );
not NOT1_11666 ( P1_R1192_U93 , P1_U3075 );
nand NAND2_11667 ( P1_R1192_U94 , P1_R1192_U393 , P1_R1192_U392 );
nand NAND2_11668 ( P1_R1192_U95 , P1_R1192_U407 , P1_R1192_U406 );
nand NAND2_11669 ( P1_R1192_U96 , P1_R1192_U412 , P1_R1192_U411 );
nand NAND2_11670 ( P1_R1192_U97 , P1_R1192_U428 , P1_R1192_U427 );
nand NAND2_11671 ( P1_R1192_U98 , P1_R1192_U433 , P1_R1192_U432 );
nand NAND2_11672 ( P1_R1192_U99 , P1_R1192_U438 , P1_R1192_U437 );
nand NAND2_11673 ( P1_R1192_U100 , P1_R1192_U443 , P1_R1192_U442 );
nand NAND2_11674 ( P1_R1192_U101 , P1_R1192_U448 , P1_R1192_U447 );
nand NAND2_11675 ( P1_R1192_U102 , P1_R1192_U464 , P1_R1192_U463 );
nand NAND2_11676 ( P1_R1192_U103 , P1_R1192_U469 , P1_R1192_U468 );
nand NAND2_11677 ( P1_R1192_U104 , P1_R1192_U352 , P1_R1192_U351 );
nand NAND2_11678 ( P1_R1192_U105 , P1_R1192_U361 , P1_R1192_U360 );
nand NAND2_11679 ( P1_R1192_U106 , P1_R1192_U368 , P1_R1192_U367 );
nand NAND2_11680 ( P1_R1192_U107 , P1_R1192_U372 , P1_R1192_U371 );
nand NAND2_11681 ( P1_R1192_U108 , P1_R1192_U381 , P1_R1192_U380 );
nand NAND2_11682 ( P1_R1192_U109 , P1_R1192_U402 , P1_R1192_U401 );
nand NAND2_11683 ( P1_R1192_U110 , P1_R1192_U419 , P1_R1192_U418 );
nand NAND2_11684 ( P1_R1192_U111 , P1_R1192_U423 , P1_R1192_U422 );
nand NAND2_11685 ( P1_R1192_U112 , P1_R1192_U455 , P1_R1192_U454 );
nand NAND2_11686 ( P1_R1192_U113 , P1_R1192_U459 , P1_R1192_U458 );
nand NAND2_11687 ( P1_R1192_U114 , P1_R1192_U476 , P1_R1192_U475 );
and AND2_11688 ( P1_R1192_U115 , P1_R1192_U195 , P1_R1192_U183 );
and AND2_11689 ( P1_R1192_U116 , P1_R1192_U198 , P1_R1192_U199 );
and AND2_11690 ( P1_R1192_U117 , P1_R1192_U211 , P1_R1192_U185 );
and AND2_11691 ( P1_R1192_U118 , P1_R1192_U214 , P1_R1192_U215 );
and AND3_11692 ( P1_R1192_U119 , P1_R1192_U354 , P1_R1192_U353 , P1_R1192_U40 );
and AND2_11693 ( P1_R1192_U120 , P1_R1192_U357 , P1_R1192_U185 );
and AND2_11694 ( P1_R1192_U121 , P1_R1192_U230 , P1_R1192_U7 );
and AND2_11695 ( P1_R1192_U122 , P1_R1192_U364 , P1_R1192_U184 );
and AND3_11696 ( P1_R1192_U123 , P1_R1192_U374 , P1_R1192_U373 , P1_R1192_U29 );
and AND2_11697 ( P1_R1192_U124 , P1_R1192_U377 , P1_R1192_U183 );
and AND2_11698 ( P1_R1192_U125 , P1_R1192_U217 , P1_R1192_U8 );
and AND2_11699 ( P1_R1192_U126 , P1_R1192_U262 , P1_R1192_U180 );
and AND2_11700 ( P1_R1192_U127 , P1_R1192_U288 , P1_R1192_U181 );
and AND2_11701 ( P1_R1192_U128 , P1_R1192_U304 , P1_R1192_U305 );
and AND2_11702 ( P1_R1192_U129 , P1_R1192_U307 , P1_R1192_U386 );
and AND3_11703 ( P1_R1192_U130 , P1_R1192_U305 , P1_R1192_U304 , P1_R1192_U308 );
nand NAND2_11704 ( P1_R1192_U131 , P1_R1192_U390 , P1_R1192_U389 );
and AND3_11705 ( P1_R1192_U132 , P1_R1192_U395 , P1_R1192_U394 , P1_R1192_U85 );
and AND2_11706 ( P1_R1192_U133 , P1_R1192_U398 , P1_R1192_U182 );
nand NAND2_11707 ( P1_R1192_U134 , P1_R1192_U404 , P1_R1192_U403 );
nand NAND2_11708 ( P1_R1192_U135 , P1_R1192_U409 , P1_R1192_U408 );
and AND2_11709 ( P1_R1192_U136 , P1_R1192_U415 , P1_R1192_U181 );
nand NAND2_11710 ( P1_R1192_U137 , P1_R1192_U425 , P1_R1192_U424 );
nand NAND2_11711 ( P1_R1192_U138 , P1_R1192_U430 , P1_R1192_U429 );
nand NAND2_11712 ( P1_R1192_U139 , P1_R1192_U435 , P1_R1192_U434 );
nand NAND2_11713 ( P1_R1192_U140 , P1_R1192_U440 , P1_R1192_U439 );
nand NAND2_11714 ( P1_R1192_U141 , P1_R1192_U445 , P1_R1192_U444 );
and AND2_11715 ( P1_R1192_U142 , P1_R1192_U451 , P1_R1192_U180 );
nand NAND2_11716 ( P1_R1192_U143 , P1_R1192_U461 , P1_R1192_U460 );
nand NAND2_11717 ( P1_R1192_U144 , P1_R1192_U466 , P1_R1192_U465 );
and AND2_11718 ( P1_R1192_U145 , P1_R1192_U342 , P1_R1192_U9 );
and AND2_11719 ( P1_R1192_U146 , P1_R1192_U472 , P1_R1192_U179 );
and AND2_11720 ( P1_R1192_U147 , P1_R1192_U350 , P1_R1192_U349 );
nand NAND2_11721 ( P1_R1192_U148 , P1_R1192_U118 , P1_R1192_U212 );
and AND2_11722 ( P1_R1192_U149 , P1_R1192_U359 , P1_R1192_U358 );
and AND2_11723 ( P1_R1192_U150 , P1_R1192_U366 , P1_R1192_U365 );
and AND2_11724 ( P1_R1192_U151 , P1_R1192_U370 , P1_R1192_U369 );
nand NAND2_11725 ( P1_R1192_U152 , P1_R1192_U116 , P1_R1192_U196 );
and AND2_11726 ( P1_R1192_U153 , P1_R1192_U379 , P1_R1192_U378 );
not NOT1_11727 ( P1_R1192_U154 , P1_U4018 );
not NOT1_11728 ( P1_R1192_U155 , P1_U3053 );
and AND2_11729 ( P1_R1192_U156 , P1_R1192_U388 , P1_R1192_U387 );
nand NAND2_11730 ( P1_R1192_U157 , P1_R1192_U128 , P1_R1192_U302 );
and AND2_11731 ( P1_R1192_U158 , P1_R1192_U400 , P1_R1192_U399 );
nand NAND2_11732 ( P1_R1192_U159 , P1_R1192_U295 , P1_R1192_U294 );
nand NAND2_11733 ( P1_R1192_U160 , P1_R1192_U291 , P1_R1192_U290 );
and AND2_11734 ( P1_R1192_U161 , P1_R1192_U417 , P1_R1192_U416 );
and AND2_11735 ( P1_R1192_U162 , P1_R1192_U421 , P1_R1192_U420 );
nand NAND2_11736 ( P1_R1192_U163 , P1_R1192_U281 , P1_R1192_U280 );
nand NAND2_11737 ( P1_R1192_U164 , P1_R1192_U277 , P1_R1192_U276 );
not NOT1_11738 ( P1_R1192_U165 , P1_U3456 );
nand NAND2_11739 ( P1_R1192_U166 , P1_R1192_U273 , P1_R1192_U272 );
not NOT1_11740 ( P1_R1192_U167 , P1_U3507 );
nand NAND2_11741 ( P1_R1192_U168 , P1_R1192_U265 , P1_R1192_U264 );
and AND2_11742 ( P1_R1192_U169 , P1_R1192_U453 , P1_R1192_U452 );
and AND2_11743 ( P1_R1192_U170 , P1_R1192_U457 , P1_R1192_U456 );
nand NAND2_11744 ( P1_R1192_U171 , P1_R1192_U255 , P1_R1192_U254 );
nand NAND2_11745 ( P1_R1192_U172 , P1_R1192_U251 , P1_R1192_U250 );
nand NAND2_11746 ( P1_R1192_U173 , P1_R1192_U247 , P1_R1192_U246 );
and AND2_11747 ( P1_R1192_U174 , P1_R1192_U474 , P1_R1192_U473 );
nand NAND2_11748 ( P1_R1192_U175 , P1_R1192_U129 , P1_R1192_U157 );
not NOT1_11749 ( P1_R1192_U176 , P1_R1192_U85 );
not NOT1_11750 ( P1_R1192_U177 , P1_R1192_U29 );
not NOT1_11751 ( P1_R1192_U178 , P1_R1192_U40 );
nand NAND2_11752 ( P1_R1192_U179 , P1_U3483 , P1_R1192_U53 );
nand NAND2_11753 ( P1_R1192_U180 , P1_U3498 , P1_R1192_U62 );
nand NAND2_11754 ( P1_R1192_U181 , P1_U4013 , P1_R1192_U76 );
nand NAND2_11755 ( P1_R1192_U182 , P1_U4009 , P1_R1192_U84 );
nand NAND2_11756 ( P1_R1192_U183 , P1_U3459 , P1_R1192_U28 );
nand NAND2_11757 ( P1_R1192_U184 , P1_U3468 , P1_R1192_U35 );
nand NAND2_11758 ( P1_R1192_U185 , P1_U3474 , P1_R1192_U39 );
not NOT1_11759 ( P1_R1192_U186 , P1_R1192_U64 );
not NOT1_11760 ( P1_R1192_U187 , P1_R1192_U78 );
not NOT1_11761 ( P1_R1192_U188 , P1_R1192_U37 );
not NOT1_11762 ( P1_R1192_U189 , P1_R1192_U54 );
not NOT1_11763 ( P1_R1192_U190 , P1_R1192_U25 );
nand NAND2_11764 ( P1_R1192_U191 , P1_R1192_U190 , P1_R1192_U26 );
nand NAND2_11765 ( P1_R1192_U192 , P1_R1192_U191 , P1_R1192_U165 );
nand NAND2_11766 ( P1_R1192_U193 , P1_U3076 , P1_R1192_U25 );
not NOT1_11767 ( P1_R1192_U194 , P1_R1192_U46 );
nand NAND2_11768 ( P1_R1192_U195 , P1_U3462 , P1_R1192_U30 );
nand NAND2_11769 ( P1_R1192_U196 , P1_R1192_U115 , P1_R1192_U46 );
nand NAND2_11770 ( P1_R1192_U197 , P1_R1192_U30 , P1_R1192_U29 );
nand NAND2_11771 ( P1_R1192_U198 , P1_R1192_U197 , P1_R1192_U27 );
nand NAND2_11772 ( P1_R1192_U199 , P1_U3062 , P1_R1192_U177 );
not NOT1_11773 ( P1_R1192_U200 , P1_R1192_U152 );
nand NAND2_11774 ( P1_R1192_U201 , P1_U3471 , P1_R1192_U34 );
nand NAND2_11775 ( P1_R1192_U202 , P1_U3069 , P1_R1192_U31 );
nand NAND2_11776 ( P1_R1192_U203 , P1_U3065 , P1_R1192_U32 );
nand NAND2_11777 ( P1_R1192_U204 , P1_R1192_U188 , P1_R1192_U6 );
nand NAND2_11778 ( P1_R1192_U205 , P1_R1192_U7 , P1_R1192_U204 );
nand NAND2_11779 ( P1_R1192_U206 , P1_U3465 , P1_R1192_U36 );
nand NAND2_11780 ( P1_R1192_U207 , P1_U3471 , P1_R1192_U34 );
nand NAND3_11781 ( P1_R1192_U208 , P1_R1192_U206 , P1_R1192_U152 , P1_R1192_U6 );
nand NAND2_11782 ( P1_R1192_U209 , P1_R1192_U207 , P1_R1192_U205 );
not NOT1_11783 ( P1_R1192_U210 , P1_R1192_U44 );
nand NAND2_11784 ( P1_R1192_U211 , P1_U3477 , P1_R1192_U41 );
nand NAND2_11785 ( P1_R1192_U212 , P1_R1192_U117 , P1_R1192_U44 );
nand NAND2_11786 ( P1_R1192_U213 , P1_R1192_U41 , P1_R1192_U40 );
nand NAND2_11787 ( P1_R1192_U214 , P1_R1192_U213 , P1_R1192_U38 );
nand NAND2_11788 ( P1_R1192_U215 , P1_U3082 , P1_R1192_U178 );
not NOT1_11789 ( P1_R1192_U216 , P1_R1192_U148 );
nand NAND2_11790 ( P1_R1192_U217 , P1_U3480 , P1_R1192_U43 );
nand NAND2_11791 ( P1_R1192_U218 , P1_R1192_U217 , P1_R1192_U54 );
nand NAND2_11792 ( P1_R1192_U219 , P1_R1192_U210 , P1_R1192_U40 );
nand NAND2_11793 ( P1_R1192_U220 , P1_R1192_U120 , P1_R1192_U219 );
nand NAND2_11794 ( P1_R1192_U221 , P1_R1192_U44 , P1_R1192_U185 );
nand NAND2_11795 ( P1_R1192_U222 , P1_R1192_U119 , P1_R1192_U221 );
nand NAND2_11796 ( P1_R1192_U223 , P1_R1192_U40 , P1_R1192_U185 );
nand NAND2_11797 ( P1_R1192_U224 , P1_R1192_U206 , P1_R1192_U152 );
not NOT1_11798 ( P1_R1192_U225 , P1_R1192_U45 );
nand NAND2_11799 ( P1_R1192_U226 , P1_U3065 , P1_R1192_U32 );
nand NAND2_11800 ( P1_R1192_U227 , P1_R1192_U225 , P1_R1192_U226 );
nand NAND2_11801 ( P1_R1192_U228 , P1_R1192_U122 , P1_R1192_U227 );
nand NAND2_11802 ( P1_R1192_U229 , P1_R1192_U45 , P1_R1192_U184 );
nand NAND2_11803 ( P1_R1192_U230 , P1_U3471 , P1_R1192_U34 );
nand NAND2_11804 ( P1_R1192_U231 , P1_R1192_U121 , P1_R1192_U229 );
nand NAND2_11805 ( P1_R1192_U232 , P1_U3065 , P1_R1192_U32 );
nand NAND2_11806 ( P1_R1192_U233 , P1_R1192_U184 , P1_R1192_U232 );
nand NAND2_11807 ( P1_R1192_U234 , P1_R1192_U206 , P1_R1192_U37 );
nand NAND2_11808 ( P1_R1192_U235 , P1_R1192_U194 , P1_R1192_U29 );
nand NAND2_11809 ( P1_R1192_U236 , P1_R1192_U124 , P1_R1192_U235 );
nand NAND2_11810 ( P1_R1192_U237 , P1_R1192_U46 , P1_R1192_U183 );
nand NAND2_11811 ( P1_R1192_U238 , P1_R1192_U123 , P1_R1192_U237 );
nand NAND2_11812 ( P1_R1192_U239 , P1_R1192_U29 , P1_R1192_U183 );
nand NAND2_11813 ( P1_R1192_U240 , P1_U3486 , P1_R1192_U52 );
nand NAND2_11814 ( P1_R1192_U241 , P1_U3061 , P1_R1192_U50 );
nand NAND2_11815 ( P1_R1192_U242 , P1_U3060 , P1_R1192_U51 );
nand NAND2_11816 ( P1_R1192_U243 , P1_R1192_U189 , P1_R1192_U8 );
nand NAND2_11817 ( P1_R1192_U244 , P1_R1192_U9 , P1_R1192_U243 );
nand NAND2_11818 ( P1_R1192_U245 , P1_U3486 , P1_R1192_U52 );
nand NAND2_11819 ( P1_R1192_U246 , P1_R1192_U125 , P1_R1192_U148 );
nand NAND2_11820 ( P1_R1192_U247 , P1_R1192_U245 , P1_R1192_U244 );
not NOT1_11821 ( P1_R1192_U248 , P1_R1192_U173 );
nand NAND2_11822 ( P1_R1192_U249 , P1_U3489 , P1_R1192_U56 );
nand NAND2_11823 ( P1_R1192_U250 , P1_R1192_U249 , P1_R1192_U173 );
nand NAND2_11824 ( P1_R1192_U251 , P1_U3070 , P1_R1192_U55 );
not NOT1_11825 ( P1_R1192_U252 , P1_R1192_U172 );
nand NAND2_11826 ( P1_R1192_U253 , P1_U3492 , P1_R1192_U58 );
nand NAND2_11827 ( P1_R1192_U254 , P1_R1192_U253 , P1_R1192_U172 );
nand NAND2_11828 ( P1_R1192_U255 , P1_U3078 , P1_R1192_U57 );
not NOT1_11829 ( P1_R1192_U256 , P1_R1192_U171 );
nand NAND2_11830 ( P1_R1192_U257 , P1_U3501 , P1_R1192_U61 );
nand NAND2_11831 ( P1_R1192_U258 , P1_U3071 , P1_R1192_U59 );
nand NAND2_11832 ( P1_R1192_U259 , P1_U3072 , P1_R1192_U49 );
nand NAND2_11833 ( P1_R1192_U260 , P1_R1192_U186 , P1_R1192_U180 );
nand NAND2_11834 ( P1_R1192_U261 , P1_R1192_U10 , P1_R1192_U260 );
nand NAND2_11835 ( P1_R1192_U262 , P1_U3495 , P1_R1192_U63 );
nand NAND2_11836 ( P1_R1192_U263 , P1_U3501 , P1_R1192_U61 );
nand NAND3_11837 ( P1_R1192_U264 , P1_R1192_U171 , P1_R1192_U126 , P1_R1192_U257 );
nand NAND2_11838 ( P1_R1192_U265 , P1_R1192_U263 , P1_R1192_U261 );
not NOT1_11839 ( P1_R1192_U266 , P1_R1192_U168 );
nand NAND2_11840 ( P1_R1192_U267 , P1_U3504 , P1_R1192_U66 );
nand NAND2_11841 ( P1_R1192_U268 , P1_R1192_U267 , P1_R1192_U168 );
nand NAND2_11842 ( P1_R1192_U269 , P1_U3067 , P1_R1192_U65 );
not NOT1_11843 ( P1_R1192_U270 , P1_R1192_U67 );
nand NAND2_11844 ( P1_R1192_U271 , P1_R1192_U270 , P1_R1192_U68 );
nand NAND2_11845 ( P1_R1192_U272 , P1_R1192_U271 , P1_R1192_U167 );
nand NAND2_11846 ( P1_R1192_U273 , P1_U3080 , P1_R1192_U67 );
not NOT1_11847 ( P1_R1192_U274 , P1_R1192_U166 );
nand NAND2_11848 ( P1_R1192_U275 , P1_U3509 , P1_R1192_U70 );
nand NAND2_11849 ( P1_R1192_U276 , P1_R1192_U275 , P1_R1192_U166 );
nand NAND2_11850 ( P1_R1192_U277 , P1_U3079 , P1_R1192_U69 );
not NOT1_11851 ( P1_R1192_U278 , P1_R1192_U164 );
nand NAND2_11852 ( P1_R1192_U279 , P1_U4015 , P1_R1192_U72 );
nand NAND2_11853 ( P1_R1192_U280 , P1_R1192_U279 , P1_R1192_U164 );
nand NAND2_11854 ( P1_R1192_U281 , P1_U3074 , P1_R1192_U71 );
not NOT1_11855 ( P1_R1192_U282 , P1_R1192_U163 );
nand NAND2_11856 ( P1_R1192_U283 , P1_U4012 , P1_R1192_U75 );
nand NAND2_11857 ( P1_R1192_U284 , P1_U3064 , P1_R1192_U73 );
nand NAND2_11858 ( P1_R1192_U285 , P1_U3059 , P1_R1192_U48 );
nand NAND2_11859 ( P1_R1192_U286 , P1_R1192_U187 , P1_R1192_U181 );
nand NAND2_11860 ( P1_R1192_U287 , P1_R1192_U11 , P1_R1192_U286 );
nand NAND2_11861 ( P1_R1192_U288 , P1_U4014 , P1_R1192_U77 );
nand NAND2_11862 ( P1_R1192_U289 , P1_U4012 , P1_R1192_U75 );
nand NAND3_11863 ( P1_R1192_U290 , P1_R1192_U163 , P1_R1192_U127 , P1_R1192_U283 );
nand NAND2_11864 ( P1_R1192_U291 , P1_R1192_U289 , P1_R1192_U287 );
not NOT1_11865 ( P1_R1192_U292 , P1_R1192_U160 );
nand NAND2_11866 ( P1_R1192_U293 , P1_U4011 , P1_R1192_U80 );
nand NAND2_11867 ( P1_R1192_U294 , P1_R1192_U293 , P1_R1192_U160 );
nand NAND2_11868 ( P1_R1192_U295 , P1_U3063 , P1_R1192_U79 );
not NOT1_11869 ( P1_R1192_U296 , P1_R1192_U159 );
nand NAND2_11870 ( P1_R1192_U297 , P1_U4010 , P1_R1192_U82 );
nand NAND2_11871 ( P1_R1192_U298 , P1_R1192_U297 , P1_R1192_U159 );
nand NAND2_11872 ( P1_R1192_U299 , P1_U3056 , P1_R1192_U81 );
not NOT1_11873 ( P1_R1192_U300 , P1_R1192_U89 );
nand NAND2_11874 ( P1_R1192_U301 , P1_U4008 , P1_R1192_U86 );
nand NAND3_11875 ( P1_R1192_U302 , P1_R1192_U89 , P1_R1192_U182 , P1_R1192_U301 );
nand NAND2_11876 ( P1_R1192_U303 , P1_R1192_U86 , P1_R1192_U85 );
nand NAND2_11877 ( P1_R1192_U304 , P1_R1192_U303 , P1_R1192_U83 );
nand NAND2_11878 ( P1_R1192_U305 , P1_U3051 , P1_R1192_U176 );
not NOT1_11879 ( P1_R1192_U306 , P1_R1192_U157 );
nand NAND2_11880 ( P1_R1192_U307 , P1_U4007 , P1_R1192_U88 );
nand NAND2_11881 ( P1_R1192_U308 , P1_U3052 , P1_R1192_U87 );
nand NAND2_11882 ( P1_R1192_U309 , P1_R1192_U300 , P1_R1192_U85 );
nand NAND2_11883 ( P1_R1192_U310 , P1_R1192_U133 , P1_R1192_U309 );
nand NAND2_11884 ( P1_R1192_U311 , P1_R1192_U89 , P1_R1192_U182 );
nand NAND2_11885 ( P1_R1192_U312 , P1_R1192_U132 , P1_R1192_U311 );
nand NAND2_11886 ( P1_R1192_U313 , P1_R1192_U85 , P1_R1192_U182 );
nand NAND2_11887 ( P1_R1192_U314 , P1_R1192_U288 , P1_R1192_U163 );
not NOT1_11888 ( P1_R1192_U315 , P1_R1192_U90 );
nand NAND2_11889 ( P1_R1192_U316 , P1_U3059 , P1_R1192_U48 );
nand NAND2_11890 ( P1_R1192_U317 , P1_R1192_U315 , P1_R1192_U316 );
nand NAND2_11891 ( P1_R1192_U318 , P1_R1192_U136 , P1_R1192_U317 );
nand NAND2_11892 ( P1_R1192_U319 , P1_R1192_U90 , P1_R1192_U181 );
nand NAND2_11893 ( P1_R1192_U320 , P1_U4012 , P1_R1192_U75 );
nand NAND3_11894 ( P1_R1192_U321 , P1_R1192_U320 , P1_R1192_U319 , P1_R1192_U11 );
nand NAND2_11895 ( P1_R1192_U322 , P1_U3059 , P1_R1192_U48 );
nand NAND2_11896 ( P1_R1192_U323 , P1_R1192_U181 , P1_R1192_U322 );
nand NAND2_11897 ( P1_R1192_U324 , P1_R1192_U288 , P1_R1192_U78 );
nand NAND2_11898 ( P1_R1192_U325 , P1_R1192_U262 , P1_R1192_U171 );
not NOT1_11899 ( P1_R1192_U326 , P1_R1192_U91 );
nand NAND2_11900 ( P1_R1192_U327 , P1_U3072 , P1_R1192_U49 );
nand NAND2_11901 ( P1_R1192_U328 , P1_R1192_U326 , P1_R1192_U327 );
nand NAND2_11902 ( P1_R1192_U329 , P1_R1192_U142 , P1_R1192_U328 );
nand NAND2_11903 ( P1_R1192_U330 , P1_R1192_U91 , P1_R1192_U180 );
nand NAND2_11904 ( P1_R1192_U331 , P1_U3501 , P1_R1192_U61 );
nand NAND3_11905 ( P1_R1192_U332 , P1_R1192_U331 , P1_R1192_U330 , P1_R1192_U10 );
nand NAND2_11906 ( P1_R1192_U333 , P1_U3072 , P1_R1192_U49 );
nand NAND2_11907 ( P1_R1192_U334 , P1_R1192_U180 , P1_R1192_U333 );
nand NAND2_11908 ( P1_R1192_U335 , P1_R1192_U262 , P1_R1192_U64 );
nand NAND2_11909 ( P1_R1192_U336 , P1_R1192_U217 , P1_R1192_U148 );
not NOT1_11910 ( P1_R1192_U337 , P1_R1192_U92 );
nand NAND2_11911 ( P1_R1192_U338 , P1_U3060 , P1_R1192_U51 );
nand NAND2_11912 ( P1_R1192_U339 , P1_R1192_U337 , P1_R1192_U338 );
nand NAND2_11913 ( P1_R1192_U340 , P1_R1192_U146 , P1_R1192_U339 );
nand NAND2_11914 ( P1_R1192_U341 , P1_R1192_U92 , P1_R1192_U179 );
nand NAND2_11915 ( P1_R1192_U342 , P1_U3486 , P1_R1192_U52 );
nand NAND2_11916 ( P1_R1192_U343 , P1_R1192_U145 , P1_R1192_U341 );
nand NAND2_11917 ( P1_R1192_U344 , P1_U3060 , P1_R1192_U51 );
nand NAND2_11918 ( P1_R1192_U345 , P1_R1192_U179 , P1_R1192_U344 );
nand NAND2_11919 ( P1_R1192_U346 , P1_U3075 , P1_R1192_U24 );
nand NAND3_11920 ( P1_R1192_U347 , P1_R1192_U89 , P1_R1192_U182 , P1_R1192_U301 );
nand NAND3_11921 ( P1_R1192_U348 , P1_R1192_U12 , P1_R1192_U347 , P1_R1192_U130 );
nand NAND2_11922 ( P1_R1192_U349 , P1_U3480 , P1_R1192_U43 );
nand NAND2_11923 ( P1_R1192_U350 , P1_U3081 , P1_R1192_U42 );
nand NAND2_11924 ( P1_R1192_U351 , P1_R1192_U218 , P1_R1192_U148 );
nand NAND2_11925 ( P1_R1192_U352 , P1_R1192_U216 , P1_R1192_U147 );
nand NAND2_11926 ( P1_R1192_U353 , P1_U3477 , P1_R1192_U41 );
nand NAND2_11927 ( P1_R1192_U354 , P1_U3082 , P1_R1192_U38 );
nand NAND2_11928 ( P1_R1192_U355 , P1_U3477 , P1_R1192_U41 );
nand NAND2_11929 ( P1_R1192_U356 , P1_U3082 , P1_R1192_U38 );
nand NAND2_11930 ( P1_R1192_U357 , P1_R1192_U356 , P1_R1192_U355 );
nand NAND2_11931 ( P1_R1192_U358 , P1_U3474 , P1_R1192_U39 );
nand NAND2_11932 ( P1_R1192_U359 , P1_U3068 , P1_R1192_U22 );
nand NAND2_11933 ( P1_R1192_U360 , P1_R1192_U223 , P1_R1192_U44 );
nand NAND2_11934 ( P1_R1192_U361 , P1_R1192_U149 , P1_R1192_U210 );
nand NAND2_11935 ( P1_R1192_U362 , P1_U3471 , P1_R1192_U34 );
nand NAND2_11936 ( P1_R1192_U363 , P1_U3069 , P1_R1192_U31 );
nand NAND2_11937 ( P1_R1192_U364 , P1_R1192_U363 , P1_R1192_U362 );
nand NAND2_11938 ( P1_R1192_U365 , P1_U3468 , P1_R1192_U35 );
nand NAND2_11939 ( P1_R1192_U366 , P1_U3065 , P1_R1192_U32 );
nand NAND2_11940 ( P1_R1192_U367 , P1_R1192_U233 , P1_R1192_U45 );
nand NAND2_11941 ( P1_R1192_U368 , P1_R1192_U150 , P1_R1192_U225 );
nand NAND2_11942 ( P1_R1192_U369 , P1_U3465 , P1_R1192_U36 );
nand NAND2_11943 ( P1_R1192_U370 , P1_U3058 , P1_R1192_U33 );
nand NAND2_11944 ( P1_R1192_U371 , P1_R1192_U234 , P1_R1192_U152 );
nand NAND2_11945 ( P1_R1192_U372 , P1_R1192_U200 , P1_R1192_U151 );
nand NAND2_11946 ( P1_R1192_U373 , P1_U3462 , P1_R1192_U30 );
nand NAND2_11947 ( P1_R1192_U374 , P1_U3062 , P1_R1192_U27 );
nand NAND2_11948 ( P1_R1192_U375 , P1_U3462 , P1_R1192_U30 );
nand NAND2_11949 ( P1_R1192_U376 , P1_U3062 , P1_R1192_U27 );
nand NAND2_11950 ( P1_R1192_U377 , P1_R1192_U376 , P1_R1192_U375 );
nand NAND2_11951 ( P1_R1192_U378 , P1_U3459 , P1_R1192_U28 );
nand NAND2_11952 ( P1_R1192_U379 , P1_U3066 , P1_R1192_U23 );
nand NAND2_11953 ( P1_R1192_U380 , P1_R1192_U239 , P1_R1192_U46 );
nand NAND2_11954 ( P1_R1192_U381 , P1_R1192_U153 , P1_R1192_U194 );
nand NAND2_11955 ( P1_R1192_U382 , P1_U4018 , P1_R1192_U155 );
nand NAND2_11956 ( P1_R1192_U383 , P1_U3053 , P1_R1192_U154 );
nand NAND2_11957 ( P1_R1192_U384 , P1_U4018 , P1_R1192_U155 );
nand NAND2_11958 ( P1_R1192_U385 , P1_U3053 , P1_R1192_U154 );
nand NAND2_11959 ( P1_R1192_U386 , P1_R1192_U385 , P1_R1192_U384 );
nand NAND3_11960 ( P1_R1192_U387 , P1_U3052 , P1_R1192_U386 , P1_R1192_U87 );
nand NAND3_11961 ( P1_R1192_U388 , P1_R1192_U12 , P1_R1192_U88 , P1_U4007 );
nand NAND2_11962 ( P1_R1192_U389 , P1_U4007 , P1_R1192_U88 );
nand NAND2_11963 ( P1_R1192_U390 , P1_U3052 , P1_R1192_U87 );
not NOT1_11964 ( P1_R1192_U391 , P1_R1192_U131 );
nand NAND2_11965 ( P1_R1192_U392 , P1_R1192_U306 , P1_R1192_U391 );
nand NAND2_11966 ( P1_R1192_U393 , P1_R1192_U131 , P1_R1192_U157 );
nand NAND2_11967 ( P1_R1192_U394 , P1_U4008 , P1_R1192_U86 );
nand NAND2_11968 ( P1_R1192_U395 , P1_U3051 , P1_R1192_U83 );
nand NAND2_11969 ( P1_R1192_U396 , P1_U4008 , P1_R1192_U86 );
nand NAND2_11970 ( P1_R1192_U397 , P1_U3051 , P1_R1192_U83 );
nand NAND2_11971 ( P1_R1192_U398 , P1_R1192_U397 , P1_R1192_U396 );
nand NAND2_11972 ( P1_R1192_U399 , P1_U4009 , P1_R1192_U84 );
nand NAND2_11973 ( P1_R1192_U400 , P1_U3055 , P1_R1192_U47 );
nand NAND2_11974 ( P1_R1192_U401 , P1_R1192_U313 , P1_R1192_U89 );
nand NAND2_11975 ( P1_R1192_U402 , P1_R1192_U158 , P1_R1192_U300 );
nand NAND2_11976 ( P1_R1192_U403 , P1_U4010 , P1_R1192_U82 );
nand NAND2_11977 ( P1_R1192_U404 , P1_U3056 , P1_R1192_U81 );
not NOT1_11978 ( P1_R1192_U405 , P1_R1192_U134 );
nand NAND2_11979 ( P1_R1192_U406 , P1_R1192_U296 , P1_R1192_U405 );
nand NAND2_11980 ( P1_R1192_U407 , P1_R1192_U134 , P1_R1192_U159 );
nand NAND2_11981 ( P1_R1192_U408 , P1_U4011 , P1_R1192_U80 );
nand NAND2_11982 ( P1_R1192_U409 , P1_U3063 , P1_R1192_U79 );
not NOT1_11983 ( P1_R1192_U410 , P1_R1192_U135 );
nand NAND2_11984 ( P1_R1192_U411 , P1_R1192_U292 , P1_R1192_U410 );
nand NAND2_11985 ( P1_R1192_U412 , P1_R1192_U135 , P1_R1192_U160 );
nand NAND2_11986 ( P1_R1192_U413 , P1_U4012 , P1_R1192_U75 );
nand NAND2_11987 ( P1_R1192_U414 , P1_U3064 , P1_R1192_U73 );
nand NAND2_11988 ( P1_R1192_U415 , P1_R1192_U414 , P1_R1192_U413 );
nand NAND2_11989 ( P1_R1192_U416 , P1_U4013 , P1_R1192_U76 );
nand NAND2_11990 ( P1_R1192_U417 , P1_U3059 , P1_R1192_U48 );
nand NAND2_11991 ( P1_R1192_U418 , P1_R1192_U323 , P1_R1192_U90 );
nand NAND2_11992 ( P1_R1192_U419 , P1_R1192_U161 , P1_R1192_U315 );
nand NAND2_11993 ( P1_R1192_U420 , P1_U4014 , P1_R1192_U77 );
nand NAND2_11994 ( P1_R1192_U421 , P1_U3073 , P1_R1192_U74 );
nand NAND2_11995 ( P1_R1192_U422 , P1_R1192_U324 , P1_R1192_U163 );
nand NAND2_11996 ( P1_R1192_U423 , P1_R1192_U282 , P1_R1192_U162 );
nand NAND2_11997 ( P1_R1192_U424 , P1_U4015 , P1_R1192_U72 );
nand NAND2_11998 ( P1_R1192_U425 , P1_U3074 , P1_R1192_U71 );
not NOT1_11999 ( P1_R1192_U426 , P1_R1192_U137 );
nand NAND2_12000 ( P1_R1192_U427 , P1_R1192_U278 , P1_R1192_U426 );
nand NAND2_12001 ( P1_R1192_U428 , P1_R1192_U137 , P1_R1192_U164 );
nand NAND2_12002 ( P1_R1192_U429 , P1_U3456 , P1_R1192_U26 );
nand NAND2_12003 ( P1_R1192_U430 , P1_U3076 , P1_R1192_U165 );
not NOT1_12004 ( P1_R1192_U431 , P1_R1192_U138 );
nand NAND2_12005 ( P1_R1192_U432 , P1_R1192_U431 , P1_R1192_U190 );
nand NAND2_12006 ( P1_R1192_U433 , P1_R1192_U138 , P1_R1192_U25 );
nand NAND2_12007 ( P1_R1192_U434 , P1_U3509 , P1_R1192_U70 );
nand NAND2_12008 ( P1_R1192_U435 , P1_U3079 , P1_R1192_U69 );
not NOT1_12009 ( P1_R1192_U436 , P1_R1192_U139 );
nand NAND2_12010 ( P1_R1192_U437 , P1_R1192_U274 , P1_R1192_U436 );
nand NAND2_12011 ( P1_R1192_U438 , P1_R1192_U139 , P1_R1192_U166 );
nand NAND2_12012 ( P1_R1192_U439 , P1_U3507 , P1_R1192_U68 );
nand NAND2_12013 ( P1_R1192_U440 , P1_U3080 , P1_R1192_U167 );
not NOT1_12014 ( P1_R1192_U441 , P1_R1192_U140 );
nand NAND2_12015 ( P1_R1192_U442 , P1_R1192_U441 , P1_R1192_U270 );
nand NAND2_12016 ( P1_R1192_U443 , P1_R1192_U140 , P1_R1192_U67 );
nand NAND2_12017 ( P1_R1192_U444 , P1_U3504 , P1_R1192_U66 );
nand NAND2_12018 ( P1_R1192_U445 , P1_U3067 , P1_R1192_U65 );
not NOT1_12019 ( P1_R1192_U446 , P1_R1192_U141 );
nand NAND2_12020 ( P1_R1192_U447 , P1_R1192_U266 , P1_R1192_U446 );
nand NAND2_12021 ( P1_R1192_U448 , P1_R1192_U141 , P1_R1192_U168 );
nand NAND2_12022 ( P1_R1192_U449 , P1_U3501 , P1_R1192_U61 );
nand NAND2_12023 ( P1_R1192_U450 , P1_U3071 , P1_R1192_U59 );
nand NAND2_12024 ( P1_R1192_U451 , P1_R1192_U450 , P1_R1192_U449 );
nand NAND2_12025 ( P1_R1192_U452 , P1_U3498 , P1_R1192_U62 );
nand NAND2_12026 ( P1_R1192_U453 , P1_U3072 , P1_R1192_U49 );
nand NAND2_12027 ( P1_R1192_U454 , P1_R1192_U334 , P1_R1192_U91 );
nand NAND2_12028 ( P1_R1192_U455 , P1_R1192_U169 , P1_R1192_U326 );
nand NAND2_12029 ( P1_R1192_U456 , P1_U3495 , P1_R1192_U63 );
nand NAND2_12030 ( P1_R1192_U457 , P1_U3077 , P1_R1192_U60 );
nand NAND2_12031 ( P1_R1192_U458 , P1_R1192_U335 , P1_R1192_U171 );
nand NAND2_12032 ( P1_R1192_U459 , P1_R1192_U256 , P1_R1192_U170 );
nand NAND2_12033 ( P1_R1192_U460 , P1_U3492 , P1_R1192_U58 );
nand NAND2_12034 ( P1_R1192_U461 , P1_U3078 , P1_R1192_U57 );
not NOT1_12035 ( P1_R1192_U462 , P1_R1192_U143 );
nand NAND2_12036 ( P1_R1192_U463 , P1_R1192_U252 , P1_R1192_U462 );
nand NAND2_12037 ( P1_R1192_U464 , P1_R1192_U143 , P1_R1192_U172 );
nand NAND2_12038 ( P1_R1192_U465 , P1_U3489 , P1_R1192_U56 );
nand NAND2_12039 ( P1_R1192_U466 , P1_U3070 , P1_R1192_U55 );
not NOT1_12040 ( P1_R1192_U467 , P1_R1192_U144 );
nand NAND2_12041 ( P1_R1192_U468 , P1_R1192_U248 , P1_R1192_U467 );
nand NAND2_12042 ( P1_R1192_U469 , P1_R1192_U144 , P1_R1192_U173 );
nand NAND2_12043 ( P1_R1192_U470 , P1_U3486 , P1_R1192_U52 );
nand NAND2_12044 ( P1_R1192_U471 , P1_U3061 , P1_R1192_U50 );
nand NAND2_12045 ( P1_R1192_U472 , P1_R1192_U471 , P1_R1192_U470 );
nand NAND2_12046 ( P1_R1192_U473 , P1_U3483 , P1_R1192_U53 );
nand NAND2_12047 ( P1_R1192_U474 , P1_U3060 , P1_R1192_U51 );
nand NAND2_12048 ( P1_R1192_U475 , P1_R1192_U345 , P1_R1192_U92 );
nand NAND2_12049 ( P1_R1192_U476 , P1_R1192_U174 , P1_R1192_U337 );
and AND2_12050 ( P1_LT_201_U6 , P1_LT_201_U109 , P1_LT_201_U108 );
and AND2_12051 ( P1_LT_201_U7 , P1_LT_201_U111 , P1_LT_201_U112 );
and AND2_12052 ( P1_LT_201_U8 , P1_LT_201_U113 , P1_LT_201_U114 );
and AND4_12053 ( P1_LT_201_U9 , P1_LT_201_U81 , P1_LT_201_U116 , P1_LT_201_U118 , P1_LT_201_U8 );
and AND2_12054 ( P1_LT_201_U10 , P1_LT_201_U126 , P1_LT_201_U125 );
and AND4_12055 ( P1_LT_201_U11 , P1_LT_201_U127 , P1_LT_201_U124 , P1_LT_201_U84 , P1_LT_201_U85 );
and AND2_12056 ( P1_LT_201_U12 , P1_LT_201_U141 , P1_LT_201_U140 );
and AND2_12057 ( P1_LT_201_U13 , P1_LT_201_U102 , P1_LT_201_U193 );
and AND2_12058 ( P1_LT_201_U14 , P1_LT_201_U189 , P1_LT_201_U104 );
not NOT1_12059 ( P1_LT_201_U15 , P1_U3594 );
not NOT1_12060 ( P1_LT_201_U16 , P1_U3595 );
not NOT1_12061 ( P1_LT_201_U17 , P1_U4017 );
not NOT1_12062 ( P1_LT_201_U18 , P1_U4018 );
not NOT1_12063 ( P1_LT_201_U19 , P1_U3599 );
not NOT1_12064 ( P1_LT_201_U20 , P1_U4011 );
not NOT1_12065 ( P1_LT_201_U21 , P1_U4010 );
not NOT1_12066 ( P1_LT_201_U22 , P1_U3604 );
not NOT1_12067 ( P1_LT_201_U23 , P1_U4014 );
not NOT1_12068 ( P1_LT_201_U24 , P1_U3605 );
not NOT1_12069 ( P1_LT_201_U25 , P1_U4015 );
not NOT1_12070 ( P1_LT_201_U26 , P1_U3509 );
not NOT1_12071 ( P1_LT_201_U27 , P1_U3609 );
not NOT1_12072 ( P1_LT_201_U28 , P1_U3507 );
not NOT1_12073 ( P1_LT_201_U29 , P1_U3610 );
not NOT1_12074 ( P1_LT_201_U30 , P1_U3608 );
not NOT1_12075 ( P1_LT_201_U31 , P1_U3606 );
not NOT1_12076 ( P1_LT_201_U32 , P1_U3504 );
not NOT1_12077 ( P1_LT_201_U33 , P1_U3501 );
not NOT1_12078 ( P1_LT_201_U34 , P1_U3611 );
not NOT1_12079 ( P1_LT_201_U35 , P1_U3612 );
not NOT1_12080 ( P1_LT_201_U36 , P1_U3474 );
not NOT1_12081 ( P1_LT_201_U37 , P1_U3590 );
not NOT1_12082 ( P1_LT_201_U38 , P1_U3471 );
not NOT1_12083 ( P1_LT_201_U39 , P1_U3591 );
not NOT1_12084 ( P1_LT_201_U40 , P1_U3587 );
not NOT1_12085 ( P1_LT_201_U41 , P1_U3617 );
not NOT1_12086 ( P1_LT_201_U42 , P1_U3588 );
not NOT1_12087 ( P1_LT_201_U43 , P1_U3589 );
not NOT1_12088 ( P1_LT_201_U44 , P1_U3592 );
not NOT1_12089 ( P1_LT_201_U45 , P1_U3593 );
nand NAND2_12090 ( P1_LT_201_U46 , P1_U3451 , P1_LT_201_U105 );
not NOT1_12091 ( P1_LT_201_U47 , P1_U3456 );
not NOT1_12092 ( P1_LT_201_U48 , P1_U3596 );
not NOT1_12093 ( P1_LT_201_U49 , P1_U3489 );
not NOT1_12094 ( P1_LT_201_U50 , P1_U3492 );
not NOT1_12095 ( P1_LT_201_U51 , P1_U3459 );
not NOT1_12096 ( P1_LT_201_U52 , P1_U3462 );
not NOT1_12097 ( P1_LT_201_U53 , P1_U3465 );
not NOT1_12098 ( P1_LT_201_U54 , P1_U3468 );
not NOT1_12099 ( P1_LT_201_U55 , P1_U3477 );
not NOT1_12100 ( P1_LT_201_U56 , P1_U3480 );
not NOT1_12101 ( P1_LT_201_U57 , P1_U3483 );
not NOT1_12102 ( P1_LT_201_U58 , P1_U3486 );
not NOT1_12103 ( P1_LT_201_U59 , P1_U3615 );
not NOT1_12104 ( P1_LT_201_U60 , P1_U3616 );
not NOT1_12105 ( P1_LT_201_U61 , P1_U3613 );
not NOT1_12106 ( P1_LT_201_U62 , P1_U3614 );
not NOT1_12107 ( P1_LT_201_U63 , P1_U3495 );
not NOT1_12108 ( P1_LT_201_U64 , P1_U3498 );
not NOT1_12109 ( P1_LT_201_U65 , P1_U4013 );
not NOT1_12110 ( P1_LT_201_U66 , P1_U4012 );
not NOT1_12111 ( P1_LT_201_U67 , P1_U3603 );
not NOT1_12112 ( P1_LT_201_U68 , P1_U3600 );
not NOT1_12113 ( P1_LT_201_U69 , P1_U3602 );
not NOT1_12114 ( P1_LT_201_U70 , P1_U3601 );
not NOT1_12115 ( P1_LT_201_U71 , P1_U4009 );
not NOT1_12116 ( P1_LT_201_U72 , P1_U4008 );
not NOT1_12117 ( P1_LT_201_U73 , P1_U4007 );
not NOT1_12118 ( P1_LT_201_U74 , P1_U3597 );
not NOT1_12119 ( P1_LT_201_U75 , P1_U4016 );
and AND2_12120 ( P1_LT_201_U76 , P1_U4014 , P1_LT_201_U24 );
and AND2_12121 ( P1_LT_201_U77 , P1_U4015 , P1_LT_201_U31 );
and AND2_12122 ( P1_LT_201_U78 , P1_LT_201_U171 , P1_LT_201_U170 );
and AND2_12123 ( P1_LT_201_U79 , P1_U3609 , P1_LT_201_U28 );
and AND2_12124 ( P1_LT_201_U80 , P1_U3610 , P1_LT_201_U32 );
and AND2_12125 ( P1_LT_201_U81 , P1_LT_201_U117 , P1_LT_201_U115 );
and AND2_12126 ( P1_LT_201_U82 , P1_U3590 , P1_LT_201_U38 );
and AND2_12127 ( P1_LT_201_U83 , P1_U3591 , P1_LT_201_U54 );
and AND2_12128 ( P1_LT_201_U84 , P1_LT_201_U129 , P1_LT_201_U128 );
and AND4_12129 ( P1_LT_201_U85 , P1_LT_201_U133 , P1_LT_201_U132 , P1_LT_201_U131 , P1_LT_201_U130 );
and AND2_12130 ( P1_LT_201_U86 , P1_LT_201_U137 , P1_LT_201_U138 );
and AND2_12131 ( P1_LT_201_U87 , P1_LT_201_U86 , P1_LT_201_U136 );
and AND2_12132 ( P1_LT_201_U88 , P1_U3459 , P1_LT_201_U48 );
and AND2_12133 ( P1_LT_201_U89 , P1_U3462 , P1_LT_201_U45 );
and AND3_12134 ( P1_LT_201_U90 , P1_LT_201_U131 , P1_LT_201_U124 , P1_LT_201_U130 );
and AND2_12135 ( P1_LT_201_U91 , P1_LT_201_U154 , P1_LT_201_U139 );
and AND2_12136 ( P1_LT_201_U92 , P1_LT_201_U157 , P1_LT_201_U156 );
and AND2_12137 ( P1_LT_201_U93 , P1_LT_201_U92 , P1_LT_201_U12 );
and AND2_12138 ( P1_LT_201_U94 , P1_U3615 , P1_LT_201_U49 );
and AND2_12139 ( P1_LT_201_U95 , P1_U3616 , P1_LT_201_U58 );
and AND2_12140 ( P1_LT_201_U96 , P1_LT_201_U160 , P1_LT_201_U161 );
and AND2_12141 ( P1_LT_201_U97 , P1_LT_201_U163 , P1_LT_201_U162 );
and AND4_12142 ( P1_LT_201_U98 , P1_LT_201_U174 , P1_LT_201_U173 , P1_LT_201_U120 , P1_LT_201_U121 );
and AND2_12143 ( P1_LT_201_U99 , P1_LT_201_U178 , P1_LT_201_U177 );
and AND2_12144 ( P1_LT_201_U100 , P1_U3603 , P1_LT_201_U66 );
and AND2_12145 ( P1_LT_201_U101 , P1_LT_201_U195 , P1_LT_201_U184 );
and AND2_12146 ( P1_LT_201_U102 , P1_LT_201_U187 , P1_LT_201_U73 );
and AND2_12147 ( P1_LT_201_U103 , P1_U3597 , P1_LT_201_U18 );
and AND3_12148 ( P1_LT_201_U104 , P1_LT_201_U191 , P1_LT_201_U107 , P1_LT_201_U190 );
not NOT1_12149 ( P1_LT_201_U105 , P1_U3618 );
nand NAND2_12150 ( P1_LT_201_U106 , P1_U3594 , P1_LT_201_U75 );
nand NAND3_12151 ( P1_LT_201_U107 , P1_LT_201_U106 , P1_U3595 , P1_LT_201_U17 );
nand NAND2_12152 ( P1_LT_201_U108 , P1_U4017 , P1_LT_201_U16 );
nand NAND2_12153 ( P1_LT_201_U109 , P1_U3594 , P1_LT_201_U75 );
nand NAND2_12154 ( P1_LT_201_U110 , P1_U3599 , P1_LT_201_U72 );
nand NAND2_12155 ( P1_LT_201_U111 , P1_U3509 , P1_LT_201_U30 );
nand NAND2_12156 ( P1_LT_201_U112 , P1_U3507 , P1_LT_201_U27 );
nand NAND2_12157 ( P1_LT_201_U113 , P1_U3604 , P1_LT_201_U65 );
nand NAND2_12158 ( P1_LT_201_U114 , P1_U3605 , P1_LT_201_U23 );
nand NAND2_12159 ( P1_LT_201_U115 , P1_LT_201_U79 , P1_LT_201_U111 );
nand NAND2_12160 ( P1_LT_201_U116 , P1_LT_201_U80 , P1_LT_201_U7 );
nand NAND2_12161 ( P1_LT_201_U117 , P1_U3608 , P1_LT_201_U26 );
nand NAND2_12162 ( P1_LT_201_U118 , P1_U3606 , P1_LT_201_U25 );
nand NAND2_12163 ( P1_LT_201_U119 , P1_U3611 , P1_LT_201_U33 );
nand NAND2_12164 ( P1_LT_201_U120 , P1_U4011 , P1_LT_201_U69 );
nand NAND2_12165 ( P1_LT_201_U121 , P1_U4010 , P1_LT_201_U70 );
nand NAND2_12166 ( P1_LT_201_U122 , P1_U3612 , P1_LT_201_U64 );
nand NAND2_12167 ( P1_LT_201_U123 , P1_U3474 , P1_LT_201_U43 );
nand NAND2_12168 ( P1_LT_201_U124 , P1_LT_201_U82 , P1_LT_201_U123 );
nand NAND2_12169 ( P1_LT_201_U125 , P1_U3471 , P1_LT_201_U37 );
nand NAND2_12170 ( P1_LT_201_U126 , P1_U3474 , P1_LT_201_U43 );
nand NAND2_12171 ( P1_LT_201_U127 , P1_LT_201_U83 , P1_LT_201_U10 );
nand NAND2_12172 ( P1_LT_201_U128 , P1_U3587 , P1_LT_201_U56 );
nand NAND2_12173 ( P1_LT_201_U129 , P1_U3617 , P1_LT_201_U57 );
nand NAND2_12174 ( P1_LT_201_U130 , P1_U3588 , P1_LT_201_U55 );
nand NAND2_12175 ( P1_LT_201_U131 , P1_U3589 , P1_LT_201_U36 );
nand NAND2_12176 ( P1_LT_201_U132 , P1_U3592 , P1_LT_201_U53 );
nand NAND2_12177 ( P1_LT_201_U133 , P1_U3593 , P1_LT_201_U52 );
not NOT1_12178 ( P1_LT_201_U134 , P1_LT_201_U46 );
nand NAND2_12179 ( P1_LT_201_U135 , P1_U3456 , P1_LT_201_U134 );
nand NAND2_12180 ( P1_LT_201_U136 , P1_U3607 , P1_LT_201_U135 );
nand NAND2_12181 ( P1_LT_201_U137 , P1_LT_201_U46 , P1_LT_201_U47 );
nand NAND2_12182 ( P1_LT_201_U138 , P1_U3596 , P1_LT_201_U51 );
nand NAND2_12183 ( P1_LT_201_U139 , P1_LT_201_U87 , P1_LT_201_U11 );
nand NAND2_12184 ( P1_LT_201_U140 , P1_U3489 , P1_LT_201_U59 );
nand NAND2_12185 ( P1_LT_201_U141 , P1_U3492 , P1_LT_201_U62 );
nand NAND2_12186 ( P1_LT_201_U142 , P1_LT_201_U89 , P1_LT_201_U132 );
nand NAND2_12187 ( P1_LT_201_U143 , P1_U3465 , P1_LT_201_U44 );
nand NAND3_12188 ( P1_LT_201_U144 , P1_LT_201_U143 , P1_LT_201_U142 , P1_LT_201_U10 );
nand NAND2_12189 ( P1_LT_201_U145 , P1_LT_201_U144 , P1_LT_201_U127 );
nand NAND2_12190 ( P1_LT_201_U146 , P1_U3468 , P1_LT_201_U39 );
nand NAND2_12191 ( P1_LT_201_U147 , P1_LT_201_U146 , P1_LT_201_U145 );
nand NAND2_12192 ( P1_LT_201_U148 , P1_LT_201_U90 , P1_LT_201_U147 );
nand NAND2_12193 ( P1_LT_201_U149 , P1_U3477 , P1_LT_201_U42 );
nand NAND2_12194 ( P1_LT_201_U150 , P1_LT_201_U149 , P1_LT_201_U148 );
nand NAND2_12195 ( P1_LT_201_U151 , P1_LT_201_U150 , P1_LT_201_U128 );
nand NAND2_12196 ( P1_LT_201_U152 , P1_U3480 , P1_LT_201_U40 );
nand NAND2_12197 ( P1_LT_201_U153 , P1_LT_201_U152 , P1_LT_201_U151 );
nand NAND2_12198 ( P1_LT_201_U154 , P1_LT_201_U88 , P1_LT_201_U11 );
nand NAND2_12199 ( P1_LT_201_U155 , P1_LT_201_U153 , P1_LT_201_U129 );
nand NAND2_12200 ( P1_LT_201_U156 , P1_U3483 , P1_LT_201_U41 );
nand NAND2_12201 ( P1_LT_201_U157 , P1_U3486 , P1_LT_201_U60 );
nand NAND3_12202 ( P1_LT_201_U158 , P1_LT_201_U91 , P1_LT_201_U155 , P1_LT_201_U93 );
nand NAND2_12203 ( P1_LT_201_U159 , P1_U3492 , P1_LT_201_U62 );
nand NAND2_12204 ( P1_LT_201_U160 , P1_LT_201_U94 , P1_LT_201_U159 );
nand NAND2_12205 ( P1_LT_201_U161 , P1_LT_201_U95 , P1_LT_201_U12 );
nand NAND2_12206 ( P1_LT_201_U162 , P1_U3613 , P1_LT_201_U63 );
nand NAND2_12207 ( P1_LT_201_U163 , P1_U3614 , P1_LT_201_U50 );
nand NAND3_12208 ( P1_LT_201_U164 , P1_LT_201_U96 , P1_LT_201_U158 , P1_LT_201_U97 );
nand NAND2_12209 ( P1_LT_201_U165 , P1_U3495 , P1_LT_201_U61 );
nand NAND2_12210 ( P1_LT_201_U166 , P1_LT_201_U165 , P1_LT_201_U164 );
nand NAND2_12211 ( P1_LT_201_U167 , P1_LT_201_U166 , P1_LT_201_U122 );
nand NAND2_12212 ( P1_LT_201_U168 , P1_U3498 , P1_LT_201_U35 );
nand NAND2_12213 ( P1_LT_201_U169 , P1_LT_201_U168 , P1_LT_201_U167 );
nand NAND2_12214 ( P1_LT_201_U170 , P1_U3504 , P1_LT_201_U29 );
nand NAND2_12215 ( P1_LT_201_U171 , P1_U3501 , P1_LT_201_U34 );
nand NAND2_12216 ( P1_LT_201_U172 , P1_LT_201_U78 , P1_LT_201_U7 );
nand NAND2_12217 ( P1_LT_201_U173 , P1_LT_201_U76 , P1_LT_201_U113 );
nand NAND2_12218 ( P1_LT_201_U174 , P1_LT_201_U77 , P1_LT_201_U8 );
nand NAND2_12219 ( P1_LT_201_U175 , P1_LT_201_U9 , P1_LT_201_U172 );
nand NAND3_12220 ( P1_LT_201_U176 , P1_LT_201_U169 , P1_LT_201_U119 , P1_LT_201_U9 );
nand NAND2_12221 ( P1_LT_201_U177 , P1_U4013 , P1_LT_201_U22 );
nand NAND2_12222 ( P1_LT_201_U178 , P1_U4012 , P1_LT_201_U67 );
nand NAND4_12223 ( P1_LT_201_U179 , P1_LT_201_U176 , P1_LT_201_U175 , P1_LT_201_U99 , P1_LT_201_U98 );
nand NAND3_12224 ( P1_LT_201_U180 , P1_LT_201_U120 , P1_LT_201_U100 , P1_LT_201_U121 );
nand NAND2_12225 ( P1_LT_201_U181 , P1_U4010 , P1_LT_201_U70 );
nand NAND2_12226 ( P1_LT_201_U182 , P1_U3602 , P1_LT_201_U20 );
nand NAND2_12227 ( P1_LT_201_U183 , P1_U3601 , P1_LT_201_U21 );
nand NAND2_12228 ( P1_LT_201_U184 , P1_U3600 , P1_LT_201_U71 );
nand NAND3_12229 ( P1_LT_201_U185 , P1_LT_201_U180 , P1_LT_201_U179 , P1_LT_201_U101 );
nand NAND2_12230 ( P1_LT_201_U186 , P1_U4009 , P1_LT_201_U68 );
nand NAND2_12231 ( P1_LT_201_U187 , P1_U4008 , P1_LT_201_U19 );
nand NAND2_12232 ( P1_LT_201_U188 , P1_U4018 , P1_LT_201_U74 );
nand NAND4_12233 ( P1_LT_201_U189 , P1_LT_201_U6 , P1_LT_201_U198 , P1_LT_201_U196 , P1_LT_201_U188 );
nand NAND2_12234 ( P1_LT_201_U190 , P1_LT_201_U103 , P1_LT_201_U6 );
nand NAND2_12235 ( P1_LT_201_U191 , P1_U4016 , P1_LT_201_U15 );
nand NAND2_12236 ( P1_LT_201_U192 , P1_LT_201_U186 , P1_LT_201_U185 );
nand NAND2_12237 ( P1_LT_201_U193 , P1_LT_201_U192 , P1_LT_201_U110 );
nand NAND2_12238 ( P1_LT_201_U194 , P1_LT_201_U183 , P1_LT_201_U182 );
nand NAND2_12239 ( P1_LT_201_U195 , P1_LT_201_U194 , P1_LT_201_U181 );
or OR2_12240 ( P1_LT_201_U196 , P1_U3598 , P1_LT_201_U13 );
nand NAND2_12241 ( P1_LT_201_U197 , P1_LT_201_U187 , P1_LT_201_U193 );
nand NAND2_12242 ( P1_LT_201_U198 , P1_U4007 , P1_LT_201_U197 );
and AND2_12243 ( P1_R1360_U6 , P1_R1360_U111 , P1_R1360_U112 );
and AND2_12244 ( P1_R1360_U7 , P1_R1360_U116 , P1_R1360_U115 );
and AND2_12245 ( P1_R1360_U8 , P1_R1360_U118 , P1_R1360_U119 );
and AND2_12246 ( P1_R1360_U9 , P1_R1360_U123 , P1_R1360_U122 );
and AND5_12247 ( P1_R1360_U10 , P1_R1360_U199 , P1_R1360_U185 , P1_R1360_U186 , P1_R1360_U184 , P1_R1360_U183 );
and AND2_12248 ( P1_R1360_U11 , P1_R1360_U183 , P1_R1360_U104 );
and AND2_12249 ( P1_R1360_U12 , P1_R1360_U203 , P1_R1360_U202 );
and AND2_12250 ( P1_R1360_U13 , P1_R1360_U205 , P1_R1360_U204 );
nand NAND3_12251 ( P1_R1360_U14 , P1_R1360_U108 , P1_R1360_U200 , P1_R1360_U107 );
not NOT1_12252 ( P1_R1360_U15 , P1_U3086 );
not NOT1_12253 ( P1_R1360_U16 , P1_U3085 );
not NOT1_12254 ( P1_R1360_U17 , P1_U3119 );
not NOT1_12255 ( P1_R1360_U18 , P1_U3087 );
not NOT1_12256 ( P1_R1360_U19 , P1_U3088 );
not NOT1_12257 ( P1_R1360_U20 , P1_U3121 );
not NOT1_12258 ( P1_R1360_U21 , P1_U3120 );
not NOT1_12259 ( P1_R1360_U22 , P1_U3118 );
not NOT1_12260 ( P1_R1360_U23 , P1_U3125 );
not NOT1_12261 ( P1_R1360_U24 , P1_U3124 );
not NOT1_12262 ( P1_R1360_U25 , P1_U3095 );
not NOT1_12263 ( P1_R1360_U26 , P1_U3096 );
not NOT1_12264 ( P1_R1360_U27 , P1_U3131 );
not NOT1_12265 ( P1_R1360_U28 , P1_U3130 );
not NOT1_12266 ( P1_R1360_U29 , P1_U3101 );
not NOT1_12267 ( P1_R1360_U30 , P1_U3102 );
not NOT1_12268 ( P1_R1360_U31 , P1_U3137 );
not NOT1_12269 ( P1_R1360_U32 , P1_U3136 );
not NOT1_12270 ( P1_R1360_U33 , P1_U3107 );
not NOT1_12271 ( P1_R1360_U34 , P1_U3140 );
not NOT1_12272 ( P1_R1360_U35 , P1_U3108 );
not NOT1_12273 ( P1_R1360_U36 , P1_U3141 );
not NOT1_12274 ( P1_R1360_U37 , P1_U3110 );
not NOT1_12275 ( P1_R1360_U38 , P1_U3109 );
not NOT1_12276 ( P1_R1360_U39 , P1_U3112 );
not NOT1_12277 ( P1_R1360_U40 , P1_U3111 );
not NOT1_12278 ( P1_R1360_U41 , P1_U3114 );
not NOT1_12279 ( P1_R1360_U42 , P1_U3113 );
not NOT1_12280 ( P1_R1360_U43 , P1_U3115 );
not NOT1_12281 ( P1_R1360_U44 , P1_U3147 );
not NOT1_12282 ( P1_R1360_U45 , P1_U3146 );
not NOT1_12283 ( P1_R1360_U46 , P1_U3145 );
not NOT1_12284 ( P1_R1360_U47 , P1_U3144 );
not NOT1_12285 ( P1_R1360_U48 , P1_U3143 );
not NOT1_12286 ( P1_R1360_U49 , P1_U3142 );
not NOT1_12287 ( P1_R1360_U50 , P1_U3139 );
not NOT1_12288 ( P1_R1360_U51 , P1_U3138 );
not NOT1_12289 ( P1_R1360_U52 , P1_U3106 );
not NOT1_12290 ( P1_R1360_U53 , P1_U3104 );
not NOT1_12291 ( P1_R1360_U54 , P1_U3105 );
not NOT1_12292 ( P1_R1360_U55 , P1_U3103 );
not NOT1_12293 ( P1_R1360_U56 , P1_U3135 );
not NOT1_12294 ( P1_R1360_U57 , P1_U3134 );
not NOT1_12295 ( P1_R1360_U58 , P1_U3133 );
not NOT1_12296 ( P1_R1360_U59 , P1_U3132 );
not NOT1_12297 ( P1_R1360_U60 , P1_U3100 );
not NOT1_12298 ( P1_R1360_U61 , P1_U3099 );
not NOT1_12299 ( P1_R1360_U62 , P1_U3098 );
not NOT1_12300 ( P1_R1360_U63 , P1_U3097 );
not NOT1_12301 ( P1_R1360_U64 , P1_U3129 );
not NOT1_12302 ( P1_R1360_U65 , P1_U3128 );
not NOT1_12303 ( P1_R1360_U66 , P1_U3127 );
not NOT1_12304 ( P1_R1360_U67 , P1_U3126 );
not NOT1_12305 ( P1_R1360_U68 , P1_U3090 );
not NOT1_12306 ( P1_R1360_U69 , P1_U3089 );
not NOT1_12307 ( P1_R1360_U70 , P1_U3093 );
not NOT1_12308 ( P1_R1360_U71 , P1_U3094 );
not NOT1_12309 ( P1_R1360_U72 , P1_U3091 );
not NOT1_12310 ( P1_R1360_U73 , P1_U3092 );
not NOT1_12311 ( P1_R1360_U74 , P1_U3122 );
not NOT1_12312 ( P1_R1360_U75 , P1_U3123 );
not NOT1_12313 ( P1_R1360_U76 , P1_U3150 );
and AND2_12314 ( P1_R1360_U77 , P1_R1360_U18 , P1_U3119 );
and AND2_12315 ( P1_R1360_U78 , P1_R1360_U183 , P1_R1360_U184 );
and AND2_12316 ( P1_R1360_U79 , P1_U3140 , P1_R1360_U35 );
and AND2_12317 ( P1_R1360_U80 , P1_U3141 , P1_R1360_U38 );
and AND4_12318 ( P1_R1360_U81 , P1_R1360_U127 , P1_R1360_U126 , P1_R1360_U125 , P1_R1360_U124 );
and AND3_12319 ( P1_R1360_U82 , P1_R1360_U130 , P1_R1360_U131 , P1_R1360_U129 );
and AND2_12320 ( P1_R1360_U83 , P1_U3147 , P1_R1360_U43 );
and AND2_12321 ( P1_R1360_U84 , P1_R1360_U85 , P1_R1360_U132 );
and AND2_12322 ( P1_R1360_U85 , P1_R1360_U144 , P1_R1360_U143 );
and AND2_12323 ( P1_R1360_U86 , P1_R1360_U121 , P1_R1360_U120 );
and AND2_12324 ( P1_R1360_U87 , P1_R1360_U8 , P1_R1360_U86 );
and AND3_12325 ( P1_R1360_U88 , P1_R1360_U147 , P1_R1360_U146 , P1_R1360_U90 );
and AND2_12326 ( P1_R1360_U89 , P1_R1360_U150 , P1_R1360_U149 );
and AND2_12327 ( P1_R1360_U90 , P1_R1360_U89 , P1_R1360_U9 );
and AND2_12328 ( P1_R1360_U91 , P1_U3106 , P1_R1360_U51 );
and AND2_12329 ( P1_R1360_U92 , P1_U3105 , P1_R1360_U31 );
and AND3_12330 ( P1_R1360_U93 , P1_R1360_U152 , P1_R1360_U153 , P1_R1360_U94 );
and AND2_12331 ( P1_R1360_U94 , P1_R1360_U156 , P1_R1360_U155 );
and AND2_12332 ( P1_R1360_U95 , P1_R1360_U7 , P1_R1360_U96 );
and AND2_12333 ( P1_R1360_U96 , P1_R1360_U164 , P1_R1360_U165 );
and AND2_12334 ( P1_R1360_U97 , P1_U3100 , P1_R1360_U59 );
and AND2_12335 ( P1_R1360_U98 , P1_U3099 , P1_R1360_U27 );
and AND3_12336 ( P1_R1360_U99 , P1_R1360_U167 , P1_R1360_U169 , P1_R1360_U100 );
and AND2_12337 ( P1_R1360_U100 , P1_R1360_U171 , P1_R1360_U170 );
and AND2_12338 ( P1_R1360_U101 , P1_R1360_U179 , P1_R1360_U180 );
and AND2_12339 ( P1_R1360_U102 , P1_U3093 , P1_R1360_U23 );
and AND2_12340 ( P1_R1360_U103 , P1_U3094 , P1_R1360_U67 );
and AND5_12341 ( P1_R1360_U104 , P1_R1360_U181 , P1_R1360_U185 , P1_R1360_U186 , P1_R1360_U106 , P1_R1360_U184 );
and AND2_12342 ( P1_R1360_U105 , P1_R1360_U190 , P1_R1360_U189 );
and AND3_12343 ( P1_R1360_U106 , P1_R1360_U188 , P1_R1360_U187 , P1_R1360_U105 );
and AND3_12344 ( P1_R1360_U107 , P1_R1360_U196 , P1_R1360_U194 , P1_R1360_U195 );
and AND2_12345 ( P1_R1360_U108 , P1_R1360_U201 , P1_R1360_U13 );
not NOT1_12346 ( P1_R1360_U109 , P1_U3117 );
nand NAND2_12347 ( P1_R1360_U110 , P1_U3095 , P1_R1360_U66 );
nand NAND2_12348 ( P1_R1360_U111 , P1_U3124 , P1_R1360_U73 );
nand NAND2_12349 ( P1_R1360_U112 , P1_U3125 , P1_R1360_U70 );
nand NAND2_12350 ( P1_R1360_U113 , P1_U3096 , P1_R1360_U65 );
nand NAND2_12351 ( P1_R1360_U114 , P1_U3101 , P1_R1360_U58 );
nand NAND2_12352 ( P1_R1360_U115 , P1_U3131 , P1_R1360_U61 );
nand NAND2_12353 ( P1_R1360_U116 , P1_U3130 , P1_R1360_U62 );
nand NAND2_12354 ( P1_R1360_U117 , P1_U3102 , P1_R1360_U57 );
nand NAND2_12355 ( P1_R1360_U118 , P1_U3107 , P1_R1360_U50 );
nand NAND2_12356 ( P1_R1360_U119 , P1_U3108 , P1_R1360_U34 );
nand NAND2_12357 ( P1_R1360_U120 , P1_U3110 , P1_R1360_U49 );
nand NAND2_12358 ( P1_R1360_U121 , P1_U3109 , P1_R1360_U36 );
nand NAND2_12359 ( P1_R1360_U122 , P1_U3137 , P1_R1360_U54 );
nand NAND2_12360 ( P1_R1360_U123 , P1_U3136 , P1_R1360_U53 );
nand NAND2_12361 ( P1_R1360_U124 , P1_U3112 , P1_R1360_U47 );
nand NAND2_12362 ( P1_R1360_U125 , P1_U3111 , P1_R1360_U48 );
nand NAND2_12363 ( P1_R1360_U126 , P1_U3114 , P1_R1360_U45 );
nand NAND2_12364 ( P1_R1360_U127 , P1_U3113 , P1_R1360_U46 );
nand NAND2_12365 ( P1_R1360_U128 , P1_U3148 , P1_U3149 );
nand NAND2_12366 ( P1_R1360_U129 , P1_U3116 , P1_R1360_U128 );
or OR2_12367 ( P1_R1360_U130 , P1_U3148 , P1_U3149 );
nand NAND2_12368 ( P1_R1360_U131 , P1_U3115 , P1_R1360_U44 );
nand NAND2_12369 ( P1_R1360_U132 , P1_R1360_U82 , P1_R1360_U81 );
nand NAND2_12370 ( P1_R1360_U133 , P1_R1360_U83 , P1_R1360_U126 );
nand NAND2_12371 ( P1_R1360_U134 , P1_U3146 , P1_R1360_U41 );
nand NAND2_12372 ( P1_R1360_U135 , P1_R1360_U134 , P1_R1360_U133 );
nand NAND2_12373 ( P1_R1360_U136 , P1_R1360_U135 , P1_R1360_U127 );
nand NAND2_12374 ( P1_R1360_U137 , P1_U3145 , P1_R1360_U42 );
nand NAND2_12375 ( P1_R1360_U138 , P1_R1360_U137 , P1_R1360_U136 );
nand NAND2_12376 ( P1_R1360_U139 , P1_R1360_U138 , P1_R1360_U124 );
nand NAND2_12377 ( P1_R1360_U140 , P1_U3144 , P1_R1360_U39 );
nand NAND2_12378 ( P1_R1360_U141 , P1_R1360_U140 , P1_R1360_U139 );
nand NAND2_12379 ( P1_R1360_U142 , P1_R1360_U141 , P1_R1360_U125 );
nand NAND2_12380 ( P1_R1360_U143 , P1_U3143 , P1_R1360_U40 );
nand NAND2_12381 ( P1_R1360_U144 , P1_U3142 , P1_R1360_U37 );
nand NAND2_12382 ( P1_R1360_U145 , P1_R1360_U142 , P1_R1360_U84 );
nand NAND2_12383 ( P1_R1360_U146 , P1_R1360_U79 , P1_R1360_U118 );
nand NAND2_12384 ( P1_R1360_U147 , P1_R1360_U80 , P1_R1360_U8 );
nand NAND2_12385 ( P1_R1360_U148 , P1_R1360_U87 , P1_R1360_U145 );
nand NAND2_12386 ( P1_R1360_U149 , P1_U3139 , P1_R1360_U33 );
nand NAND2_12387 ( P1_R1360_U150 , P1_U3138 , P1_R1360_U52 );
nand NAND2_12388 ( P1_R1360_U151 , P1_R1360_U148 , P1_R1360_U88 );
nand NAND2_12389 ( P1_R1360_U152 , P1_R1360_U91 , P1_R1360_U9 );
nand NAND2_12390 ( P1_R1360_U153 , P1_U3104 , P1_R1360_U32 );
nand NAND2_12391 ( P1_R1360_U154 , P1_U3136 , P1_R1360_U53 );
nand NAND2_12392 ( P1_R1360_U155 , P1_R1360_U92 , P1_R1360_U154 );
nand NAND2_12393 ( P1_R1360_U156 , P1_U3103 , P1_R1360_U56 );
nand NAND2_12394 ( P1_R1360_U157 , P1_R1360_U151 , P1_R1360_U93 );
nand NAND2_12395 ( P1_R1360_U158 , P1_U3135 , P1_R1360_U55 );
nand NAND2_12396 ( P1_R1360_U159 , P1_R1360_U158 , P1_R1360_U157 );
nand NAND2_12397 ( P1_R1360_U160 , P1_R1360_U159 , P1_R1360_U117 );
nand NAND2_12398 ( P1_R1360_U161 , P1_U3134 , P1_R1360_U30 );
nand NAND2_12399 ( P1_R1360_U162 , P1_R1360_U161 , P1_R1360_U160 );
nand NAND2_12400 ( P1_R1360_U163 , P1_R1360_U162 , P1_R1360_U114 );
nand NAND2_12401 ( P1_R1360_U164 , P1_U3133 , P1_R1360_U29 );
nand NAND2_12402 ( P1_R1360_U165 , P1_U3132 , P1_R1360_U60 );
nand NAND2_12403 ( P1_R1360_U166 , P1_R1360_U163 , P1_R1360_U95 );
nand NAND2_12404 ( P1_R1360_U167 , P1_R1360_U97 , P1_R1360_U7 );
nand NAND2_12405 ( P1_R1360_U168 , P1_U3130 , P1_R1360_U62 );
nand NAND2_12406 ( P1_R1360_U169 , P1_R1360_U98 , P1_R1360_U168 );
nand NAND2_12407 ( P1_R1360_U170 , P1_U3098 , P1_R1360_U28 );
nand NAND2_12408 ( P1_R1360_U171 , P1_U3097 , P1_R1360_U64 );
nand NAND2_12409 ( P1_R1360_U172 , P1_R1360_U166 , P1_R1360_U99 );
nand NAND2_12410 ( P1_R1360_U173 , P1_U3129 , P1_R1360_U63 );
nand NAND2_12411 ( P1_R1360_U174 , P1_R1360_U173 , P1_R1360_U172 );
nand NAND2_12412 ( P1_R1360_U175 , P1_R1360_U174 , P1_R1360_U113 );
nand NAND2_12413 ( P1_R1360_U176 , P1_U3128 , P1_R1360_U26 );
nand NAND2_12414 ( P1_R1360_U177 , P1_R1360_U176 , P1_R1360_U175 );
nand NAND2_12415 ( P1_R1360_U178 , P1_R1360_U177 , P1_R1360_U110 );
nand NAND2_12416 ( P1_R1360_U179 , P1_U3127 , P1_R1360_U25 );
nand NAND2_12417 ( P1_R1360_U180 , P1_U3126 , P1_R1360_U71 );
nand NAND3_12418 ( P1_R1360_U181 , P1_R1360_U101 , P1_R1360_U178 , P1_R1360_U6 );
nand NAND2_12419 ( P1_R1360_U182 , P1_U3086 , P1_R1360_U22 );
nand NAND2_12420 ( P1_R1360_U183 , P1_U3087 , P1_R1360_U17 );
nand NAND2_12421 ( P1_R1360_U184 , P1_U3088 , P1_R1360_U21 );
nand NAND2_12422 ( P1_R1360_U185 , P1_U3090 , P1_R1360_U74 );
nand NAND2_12423 ( P1_R1360_U186 , P1_U3089 , P1_R1360_U20 );
nand NAND2_12424 ( P1_R1360_U187 , P1_R1360_U102 , P1_R1360_U111 );
nand NAND2_12425 ( P1_R1360_U188 , P1_R1360_U103 , P1_R1360_U6 );
nand NAND2_12426 ( P1_R1360_U189 , P1_U3091 , P1_R1360_U75 );
nand NAND2_12427 ( P1_R1360_U190 , P1_U3092 , P1_R1360_U24 );
nand NAND2_12428 ( P1_R1360_U191 , P1_U3121 , P1_R1360_U69 );
nand NAND2_12429 ( P1_R1360_U192 , P1_U3120 , P1_R1360_U19 );
nand NAND2_12430 ( P1_R1360_U193 , P1_R1360_U192 , P1_R1360_U191 );
nand NAND3_12431 ( P1_R1360_U194 , P1_R1360_U77 , P1_R1360_U12 , P1_R1360_U182 );
nand NAND4_12432 ( P1_R1360_U195 , P1_R1360_U12 , P1_R1360_U193 , P1_R1360_U78 , P1_R1360_U182 );
nand NAND3_12433 ( P1_R1360_U196 , P1_R1360_U12 , P1_R1360_U15 , P1_U3118 );
nand NAND2_12434 ( P1_R1360_U197 , P1_U3122 , P1_R1360_U68 );
nand NAND2_12435 ( P1_R1360_U198 , P1_U3123 , P1_R1360_U72 );
nand NAND2_12436 ( P1_R1360_U199 , P1_R1360_U198 , P1_R1360_U197 );
nand NAND3_12437 ( P1_R1360_U200 , P1_R1360_U12 , P1_R1360_U11 , P1_R1360_U182 );
nand NAND3_12438 ( P1_R1360_U201 , P1_R1360_U12 , P1_R1360_U10 , P1_R1360_U182 );
nand NAND2_12439 ( P1_R1360_U202 , P1_U3085 , P1_R1360_U109 );
nand NAND2_12440 ( P1_R1360_U203 , P1_U3117 , P1_R1360_U16 );
nand NAND3_12441 ( P1_R1360_U204 , P1_U3150 , P1_U3085 , P1_R1360_U109 );
nand NAND3_12442 ( P1_R1360_U205 , P1_R1360_U76 , P1_R1360_U16 , P1_U3117 );
and AND2_12443 ( P1_R1171_U4 , P1_R1171_U176 , P1_R1171_U175 );
and AND2_12444 ( P1_R1171_U5 , P1_R1171_U177 , P1_R1171_U178 );
and AND2_12445 ( P1_R1171_U6 , P1_R1171_U194 , P1_R1171_U193 );
and AND2_12446 ( P1_R1171_U7 , P1_R1171_U234 , P1_R1171_U233 );
and AND2_12447 ( P1_R1171_U8 , P1_R1171_U243 , P1_R1171_U242 );
and AND2_12448 ( P1_R1171_U9 , P1_R1171_U261 , P1_R1171_U260 );
and AND2_12449 ( P1_R1171_U10 , P1_R1171_U269 , P1_R1171_U268 );
and AND2_12450 ( P1_R1171_U11 , P1_R1171_U348 , P1_R1171_U345 );
and AND2_12451 ( P1_R1171_U12 , P1_R1171_U341 , P1_R1171_U338 );
and AND2_12452 ( P1_R1171_U13 , P1_R1171_U332 , P1_R1171_U329 );
and AND2_12453 ( P1_R1171_U14 , P1_R1171_U323 , P1_R1171_U320 );
and AND2_12454 ( P1_R1171_U15 , P1_R1171_U317 , P1_R1171_U315 );
and AND2_12455 ( P1_R1171_U16 , P1_R1171_U310 , P1_R1171_U307 );
and AND2_12456 ( P1_R1171_U17 , P1_R1171_U232 , P1_R1171_U229 );
and AND2_12457 ( P1_R1171_U18 , P1_R1171_U224 , P1_R1171_U221 );
and AND2_12458 ( P1_R1171_U19 , P1_R1171_U210 , P1_R1171_U207 );
not NOT1_12459 ( P1_R1171_U20 , P1_U3471 );
not NOT1_12460 ( P1_R1171_U21 , P1_U3069 );
not NOT1_12461 ( P1_R1171_U22 , P1_U3068 );
nand NAND2_12462 ( P1_R1171_U23 , P1_U3069 , P1_U3471 );
not NOT1_12463 ( P1_R1171_U24 , P1_U3474 );
not NOT1_12464 ( P1_R1171_U25 , P1_U3465 );
not NOT1_12465 ( P1_R1171_U26 , P1_U3058 );
not NOT1_12466 ( P1_R1171_U27 , P1_U3065 );
not NOT1_12467 ( P1_R1171_U28 , P1_U3459 );
not NOT1_12468 ( P1_R1171_U29 , P1_U3066 );
not NOT1_12469 ( P1_R1171_U30 , P1_U3451 );
not NOT1_12470 ( P1_R1171_U31 , P1_U3075 );
nand NAND2_12471 ( P1_R1171_U32 , P1_U3075 , P1_U3451 );
not NOT1_12472 ( P1_R1171_U33 , P1_U3462 );
not NOT1_12473 ( P1_R1171_U34 , P1_U3062 );
nand NAND2_12474 ( P1_R1171_U35 , P1_U3058 , P1_U3465 );
not NOT1_12475 ( P1_R1171_U36 , P1_U3468 );
not NOT1_12476 ( P1_R1171_U37 , P1_U3477 );
not NOT1_12477 ( P1_R1171_U38 , P1_U3082 );
not NOT1_12478 ( P1_R1171_U39 , P1_U3081 );
not NOT1_12479 ( P1_R1171_U40 , P1_U3480 );
nand NAND2_12480 ( P1_R1171_U41 , P1_R1171_U62 , P1_R1171_U202 );
nand NAND2_12481 ( P1_R1171_U42 , P1_R1171_U118 , P1_R1171_U190 );
nand NAND2_12482 ( P1_R1171_U43 , P1_R1171_U179 , P1_R1171_U180 );
nand NAND2_12483 ( P1_R1171_U44 , P1_U3456 , P1_U3076 );
nand NAND2_12484 ( P1_R1171_U45 , P1_R1171_U122 , P1_R1171_U216 );
nand NAND2_12485 ( P1_R1171_U46 , P1_R1171_U213 , P1_R1171_U212 );
not NOT1_12486 ( P1_R1171_U47 , P1_U4008 );
not NOT1_12487 ( P1_R1171_U48 , P1_U3051 );
not NOT1_12488 ( P1_R1171_U49 , P1_U3055 );
not NOT1_12489 ( P1_R1171_U50 , P1_U4009 );
not NOT1_12490 ( P1_R1171_U51 , P1_U4010 );
not NOT1_12491 ( P1_R1171_U52 , P1_U3056 );
not NOT1_12492 ( P1_R1171_U53 , P1_U4011 );
not NOT1_12493 ( P1_R1171_U54 , P1_U3063 );
not NOT1_12494 ( P1_R1171_U55 , P1_U4014 );
not NOT1_12495 ( P1_R1171_U56 , P1_U3073 );
not NOT1_12496 ( P1_R1171_U57 , P1_U3501 );
not NOT1_12497 ( P1_R1171_U58 , P1_U3071 );
not NOT1_12498 ( P1_R1171_U59 , P1_U3067 );
nand NAND2_12499 ( P1_R1171_U60 , P1_U3071 , P1_U3501 );
not NOT1_12500 ( P1_R1171_U61 , P1_U3504 );
nand NAND2_12501 ( P1_R1171_U62 , P1_U3082 , P1_U3477 );
not NOT1_12502 ( P1_R1171_U63 , P1_U3483 );
not NOT1_12503 ( P1_R1171_U64 , P1_U3060 );
not NOT1_12504 ( P1_R1171_U65 , P1_U3489 );
not NOT1_12505 ( P1_R1171_U66 , P1_U3070 );
not NOT1_12506 ( P1_R1171_U67 , P1_U3486 );
not NOT1_12507 ( P1_R1171_U68 , P1_U3061 );
nand NAND2_12508 ( P1_R1171_U69 , P1_U3061 , P1_U3486 );
not NOT1_12509 ( P1_R1171_U70 , P1_U3492 );
not NOT1_12510 ( P1_R1171_U71 , P1_U3078 );
not NOT1_12511 ( P1_R1171_U72 , P1_U3495 );
not NOT1_12512 ( P1_R1171_U73 , P1_U3077 );
not NOT1_12513 ( P1_R1171_U74 , P1_U3498 );
not NOT1_12514 ( P1_R1171_U75 , P1_U3072 );
not NOT1_12515 ( P1_R1171_U76 , P1_U3507 );
not NOT1_12516 ( P1_R1171_U77 , P1_U3080 );
nand NAND2_12517 ( P1_R1171_U78 , P1_U3080 , P1_U3507 );
not NOT1_12518 ( P1_R1171_U79 , P1_U3509 );
not NOT1_12519 ( P1_R1171_U80 , P1_U3079 );
nand NAND2_12520 ( P1_R1171_U81 , P1_U3079 , P1_U3509 );
not NOT1_12521 ( P1_R1171_U82 , P1_U4015 );
not NOT1_12522 ( P1_R1171_U83 , P1_U4013 );
not NOT1_12523 ( P1_R1171_U84 , P1_U3059 );
not NOT1_12524 ( P1_R1171_U85 , P1_U4012 );
not NOT1_12525 ( P1_R1171_U86 , P1_U3064 );
nand NAND2_12526 ( P1_R1171_U87 , P1_U4009 , P1_U3055 );
not NOT1_12527 ( P1_R1171_U88 , P1_U3052 );
not NOT1_12528 ( P1_R1171_U89 , P1_U4007 );
nand NAND2_12529 ( P1_R1171_U90 , P1_R1171_U303 , P1_R1171_U173 );
not NOT1_12530 ( P1_R1171_U91 , P1_U3074 );
nand NAND2_12531 ( P1_R1171_U92 , P1_R1171_U78 , P1_R1171_U312 );
nand NAND2_12532 ( P1_R1171_U93 , P1_R1171_U258 , P1_R1171_U257 );
nand NAND2_12533 ( P1_R1171_U94 , P1_R1171_U69 , P1_R1171_U334 );
nand NAND2_12534 ( P1_R1171_U95 , P1_R1171_U454 , P1_R1171_U453 );
nand NAND2_12535 ( P1_R1171_U96 , P1_R1171_U501 , P1_R1171_U500 );
nand NAND2_12536 ( P1_R1171_U97 , P1_R1171_U372 , P1_R1171_U371 );
nand NAND2_12537 ( P1_R1171_U98 , P1_R1171_U377 , P1_R1171_U376 );
nand NAND2_12538 ( P1_R1171_U99 , P1_R1171_U384 , P1_R1171_U383 );
nand NAND2_12539 ( P1_R1171_U100 , P1_R1171_U391 , P1_R1171_U390 );
nand NAND2_12540 ( P1_R1171_U101 , P1_R1171_U396 , P1_R1171_U395 );
nand NAND2_12541 ( P1_R1171_U102 , P1_R1171_U405 , P1_R1171_U404 );
nand NAND2_12542 ( P1_R1171_U103 , P1_R1171_U412 , P1_R1171_U411 );
nand NAND2_12543 ( P1_R1171_U104 , P1_R1171_U419 , P1_R1171_U418 );
nand NAND2_12544 ( P1_R1171_U105 , P1_R1171_U426 , P1_R1171_U425 );
nand NAND2_12545 ( P1_R1171_U106 , P1_R1171_U431 , P1_R1171_U430 );
nand NAND2_12546 ( P1_R1171_U107 , P1_R1171_U438 , P1_R1171_U437 );
nand NAND2_12547 ( P1_R1171_U108 , P1_R1171_U445 , P1_R1171_U444 );
nand NAND2_12548 ( P1_R1171_U109 , P1_R1171_U459 , P1_R1171_U458 );
nand NAND2_12549 ( P1_R1171_U110 , P1_R1171_U464 , P1_R1171_U463 );
nand NAND2_12550 ( P1_R1171_U111 , P1_R1171_U471 , P1_R1171_U470 );
nand NAND2_12551 ( P1_R1171_U112 , P1_R1171_U478 , P1_R1171_U477 );
nand NAND2_12552 ( P1_R1171_U113 , P1_R1171_U485 , P1_R1171_U484 );
nand NAND2_12553 ( P1_R1171_U114 , P1_R1171_U492 , P1_R1171_U491 );
nand NAND2_12554 ( P1_R1171_U115 , P1_R1171_U497 , P1_R1171_U496 );
and AND2_12555 ( P1_R1171_U116 , P1_U3459 , P1_U3066 );
and AND2_12556 ( P1_R1171_U117 , P1_R1171_U186 , P1_R1171_U184 );
and AND2_12557 ( P1_R1171_U118 , P1_R1171_U191 , P1_R1171_U189 );
and AND2_12558 ( P1_R1171_U119 , P1_R1171_U198 , P1_R1171_U197 );
and AND3_12559 ( P1_R1171_U120 , P1_R1171_U379 , P1_R1171_U378 , P1_R1171_U23 );
and AND2_12560 ( P1_R1171_U121 , P1_R1171_U209 , P1_R1171_U6 );
and AND2_12561 ( P1_R1171_U122 , P1_R1171_U217 , P1_R1171_U215 );
and AND3_12562 ( P1_R1171_U123 , P1_R1171_U386 , P1_R1171_U385 , P1_R1171_U35 );
and AND2_12563 ( P1_R1171_U124 , P1_R1171_U223 , P1_R1171_U4 );
and AND2_12564 ( P1_R1171_U125 , P1_R1171_U231 , P1_R1171_U178 );
and AND2_12565 ( P1_R1171_U126 , P1_R1171_U201 , P1_R1171_U7 );
and AND2_12566 ( P1_R1171_U127 , P1_R1171_U236 , P1_R1171_U168 );
and AND2_12567 ( P1_R1171_U128 , P1_R1171_U245 , P1_R1171_U169 );
and AND2_12568 ( P1_R1171_U129 , P1_R1171_U265 , P1_R1171_U264 );
and AND2_12569 ( P1_R1171_U130 , P1_R1171_U10 , P1_R1171_U279 );
and AND2_12570 ( P1_R1171_U131 , P1_R1171_U282 , P1_R1171_U277 );
and AND2_12571 ( P1_R1171_U132 , P1_R1171_U298 , P1_R1171_U295 );
and AND2_12572 ( P1_R1171_U133 , P1_R1171_U365 , P1_R1171_U299 );
and AND2_12573 ( P1_R1171_U134 , P1_R1171_U156 , P1_R1171_U275 );
and AND3_12574 ( P1_R1171_U135 , P1_R1171_U466 , P1_R1171_U465 , P1_R1171_U60 );
and AND3_12575 ( P1_R1171_U136 , P1_R1171_U487 , P1_R1171_U486 , P1_R1171_U169 );
and AND2_12576 ( P1_R1171_U137 , P1_R1171_U340 , P1_R1171_U8 );
and AND3_12577 ( P1_R1171_U138 , P1_R1171_U499 , P1_R1171_U498 , P1_R1171_U168 );
and AND2_12578 ( P1_R1171_U139 , P1_R1171_U347 , P1_R1171_U7 );
nand NAND2_12579 ( P1_R1171_U140 , P1_R1171_U119 , P1_R1171_U199 );
nand NAND2_12580 ( P1_R1171_U141 , P1_R1171_U214 , P1_R1171_U226 );
not NOT1_12581 ( P1_R1171_U142 , P1_U3053 );
not NOT1_12582 ( P1_R1171_U143 , P1_U4018 );
and AND2_12583 ( P1_R1171_U144 , P1_R1171_U400 , P1_R1171_U399 );
nand NAND3_12584 ( P1_R1171_U145 , P1_R1171_U301 , P1_R1171_U166 , P1_R1171_U361 );
and AND2_12585 ( P1_R1171_U146 , P1_R1171_U407 , P1_R1171_U406 );
nand NAND3_12586 ( P1_R1171_U147 , P1_R1171_U367 , P1_R1171_U366 , P1_R1171_U133 );
and AND2_12587 ( P1_R1171_U148 , P1_R1171_U414 , P1_R1171_U413 );
nand NAND3_12588 ( P1_R1171_U149 , P1_R1171_U362 , P1_R1171_U296 , P1_R1171_U87 );
and AND2_12589 ( P1_R1171_U150 , P1_R1171_U421 , P1_R1171_U420 );
nand NAND2_12590 ( P1_R1171_U151 , P1_R1171_U290 , P1_R1171_U289 );
and AND2_12591 ( P1_R1171_U152 , P1_R1171_U433 , P1_R1171_U432 );
nand NAND2_12592 ( P1_R1171_U153 , P1_R1171_U286 , P1_R1171_U285 );
and AND2_12593 ( P1_R1171_U154 , P1_R1171_U440 , P1_R1171_U439 );
nand NAND2_12594 ( P1_R1171_U155 , P1_R1171_U131 , P1_R1171_U281 );
and AND2_12595 ( P1_R1171_U156 , P1_R1171_U447 , P1_R1171_U446 );
and AND2_12596 ( P1_R1171_U157 , P1_R1171_U452 , P1_R1171_U451 );
nand NAND2_12597 ( P1_R1171_U158 , P1_R1171_U44 , P1_R1171_U324 );
nand NAND2_12598 ( P1_R1171_U159 , P1_R1171_U129 , P1_R1171_U266 );
and AND2_12599 ( P1_R1171_U160 , P1_R1171_U473 , P1_R1171_U472 );
nand NAND2_12600 ( P1_R1171_U161 , P1_R1171_U254 , P1_R1171_U253 );
and AND2_12601 ( P1_R1171_U162 , P1_R1171_U480 , P1_R1171_U479 );
nand NAND2_12602 ( P1_R1171_U163 , P1_R1171_U250 , P1_R1171_U249 );
nand NAND2_12603 ( P1_R1171_U164 , P1_R1171_U240 , P1_R1171_U239 );
nand NAND2_12604 ( P1_R1171_U165 , P1_R1171_U364 , P1_R1171_U363 );
nand NAND2_12605 ( P1_R1171_U166 , P1_U3052 , P1_R1171_U147 );
not NOT1_12606 ( P1_R1171_U167 , P1_R1171_U35 );
nand NAND2_12607 ( P1_R1171_U168 , P1_U3480 , P1_U3081 );
nand NAND2_12608 ( P1_R1171_U169 , P1_U3070 , P1_U3489 );
nand NAND2_12609 ( P1_R1171_U170 , P1_U3056 , P1_U4010 );
not NOT1_12610 ( P1_R1171_U171 , P1_R1171_U69 );
not NOT1_12611 ( P1_R1171_U172 , P1_R1171_U78 );
nand NAND2_12612 ( P1_R1171_U173 , P1_U3063 , P1_U4011 );
not NOT1_12613 ( P1_R1171_U174 , P1_R1171_U62 );
or OR2_12614 ( P1_R1171_U175 , P1_U3065 , P1_U3468 );
or OR2_12615 ( P1_R1171_U176 , P1_U3058 , P1_U3465 );
or OR2_12616 ( P1_R1171_U177 , P1_U3462 , P1_U3062 );
or OR2_12617 ( P1_R1171_U178 , P1_U3459 , P1_U3066 );
not NOT1_12618 ( P1_R1171_U179 , P1_R1171_U32 );
or OR2_12619 ( P1_R1171_U180 , P1_U3456 , P1_U3076 );
not NOT1_12620 ( P1_R1171_U181 , P1_R1171_U43 );
not NOT1_12621 ( P1_R1171_U182 , P1_R1171_U44 );
nand NAND2_12622 ( P1_R1171_U183 , P1_R1171_U43 , P1_R1171_U44 );
nand NAND2_12623 ( P1_R1171_U184 , P1_R1171_U116 , P1_R1171_U177 );
nand NAND2_12624 ( P1_R1171_U185 , P1_R1171_U5 , P1_R1171_U183 );
nand NAND2_12625 ( P1_R1171_U186 , P1_U3062 , P1_U3462 );
nand NAND2_12626 ( P1_R1171_U187 , P1_R1171_U117 , P1_R1171_U185 );
nand NAND2_12627 ( P1_R1171_U188 , P1_R1171_U36 , P1_R1171_U35 );
nand NAND2_12628 ( P1_R1171_U189 , P1_U3065 , P1_R1171_U188 );
nand NAND2_12629 ( P1_R1171_U190 , P1_R1171_U4 , P1_R1171_U187 );
nand NAND2_12630 ( P1_R1171_U191 , P1_U3468 , P1_R1171_U167 );
not NOT1_12631 ( P1_R1171_U192 , P1_R1171_U42 );
or OR2_12632 ( P1_R1171_U193 , P1_U3068 , P1_U3474 );
or OR2_12633 ( P1_R1171_U194 , P1_U3069 , P1_U3471 );
not NOT1_12634 ( P1_R1171_U195 , P1_R1171_U23 );
nand NAND2_12635 ( P1_R1171_U196 , P1_R1171_U24 , P1_R1171_U23 );
nand NAND2_12636 ( P1_R1171_U197 , P1_U3068 , P1_R1171_U196 );
nand NAND2_12637 ( P1_R1171_U198 , P1_U3474 , P1_R1171_U195 );
nand NAND2_12638 ( P1_R1171_U199 , P1_R1171_U6 , P1_R1171_U42 );
not NOT1_12639 ( P1_R1171_U200 , P1_R1171_U140 );
or OR2_12640 ( P1_R1171_U201 , P1_U3477 , P1_U3082 );
nand NAND2_12641 ( P1_R1171_U202 , P1_R1171_U201 , P1_R1171_U140 );
not NOT1_12642 ( P1_R1171_U203 , P1_R1171_U41 );
or OR2_12643 ( P1_R1171_U204 , P1_U3081 , P1_U3480 );
or OR2_12644 ( P1_R1171_U205 , P1_U3471 , P1_U3069 );
nand NAND2_12645 ( P1_R1171_U206 , P1_R1171_U205 , P1_R1171_U42 );
nand NAND2_12646 ( P1_R1171_U207 , P1_R1171_U120 , P1_R1171_U206 );
nand NAND2_12647 ( P1_R1171_U208 , P1_R1171_U192 , P1_R1171_U23 );
nand NAND2_12648 ( P1_R1171_U209 , P1_U3474 , P1_U3068 );
nand NAND2_12649 ( P1_R1171_U210 , P1_R1171_U121 , P1_R1171_U208 );
or OR2_12650 ( P1_R1171_U211 , P1_U3069 , P1_U3471 );
nand NAND2_12651 ( P1_R1171_U212 , P1_R1171_U182 , P1_R1171_U178 );
nand NAND2_12652 ( P1_R1171_U213 , P1_U3066 , P1_U3459 );
not NOT1_12653 ( P1_R1171_U214 , P1_R1171_U46 );
nand NAND2_12654 ( P1_R1171_U215 , P1_R1171_U181 , P1_R1171_U5 );
nand NAND2_12655 ( P1_R1171_U216 , P1_R1171_U46 , P1_R1171_U177 );
nand NAND2_12656 ( P1_R1171_U217 , P1_U3062 , P1_U3462 );
not NOT1_12657 ( P1_R1171_U218 , P1_R1171_U45 );
or OR2_12658 ( P1_R1171_U219 , P1_U3465 , P1_U3058 );
nand NAND2_12659 ( P1_R1171_U220 , P1_R1171_U219 , P1_R1171_U45 );
nand NAND2_12660 ( P1_R1171_U221 , P1_R1171_U123 , P1_R1171_U220 );
nand NAND2_12661 ( P1_R1171_U222 , P1_R1171_U218 , P1_R1171_U35 );
nand NAND2_12662 ( P1_R1171_U223 , P1_U3468 , P1_U3065 );
nand NAND2_12663 ( P1_R1171_U224 , P1_R1171_U124 , P1_R1171_U222 );
or OR2_12664 ( P1_R1171_U225 , P1_U3058 , P1_U3465 );
nand NAND2_12665 ( P1_R1171_U226 , P1_R1171_U181 , P1_R1171_U178 );
not NOT1_12666 ( P1_R1171_U227 , P1_R1171_U141 );
nand NAND2_12667 ( P1_R1171_U228 , P1_U3062 , P1_U3462 );
nand NAND4_12668 ( P1_R1171_U229 , P1_R1171_U398 , P1_R1171_U397 , P1_R1171_U44 , P1_R1171_U43 );
nand NAND2_12669 ( P1_R1171_U230 , P1_R1171_U44 , P1_R1171_U43 );
nand NAND2_12670 ( P1_R1171_U231 , P1_U3066 , P1_U3459 );
nand NAND2_12671 ( P1_R1171_U232 , P1_R1171_U125 , P1_R1171_U230 );
or OR2_12672 ( P1_R1171_U233 , P1_U3081 , P1_U3480 );
or OR2_12673 ( P1_R1171_U234 , P1_U3060 , P1_U3483 );
nand NAND2_12674 ( P1_R1171_U235 , P1_R1171_U174 , P1_R1171_U7 );
nand NAND2_12675 ( P1_R1171_U236 , P1_U3060 , P1_U3483 );
nand NAND2_12676 ( P1_R1171_U237 , P1_R1171_U127 , P1_R1171_U235 );
or OR2_12677 ( P1_R1171_U238 , P1_U3483 , P1_U3060 );
nand NAND2_12678 ( P1_R1171_U239 , P1_R1171_U126 , P1_R1171_U140 );
nand NAND2_12679 ( P1_R1171_U240 , P1_R1171_U238 , P1_R1171_U237 );
not NOT1_12680 ( P1_R1171_U241 , P1_R1171_U164 );
or OR2_12681 ( P1_R1171_U242 , P1_U3078 , P1_U3492 );
or OR2_12682 ( P1_R1171_U243 , P1_U3070 , P1_U3489 );
nand NAND2_12683 ( P1_R1171_U244 , P1_R1171_U171 , P1_R1171_U8 );
nand NAND2_12684 ( P1_R1171_U245 , P1_U3078 , P1_U3492 );
nand NAND2_12685 ( P1_R1171_U246 , P1_R1171_U128 , P1_R1171_U244 );
or OR2_12686 ( P1_R1171_U247 , P1_U3486 , P1_U3061 );
or OR2_12687 ( P1_R1171_U248 , P1_U3492 , P1_U3078 );
nand NAND3_12688 ( P1_R1171_U249 , P1_R1171_U247 , P1_R1171_U164 , P1_R1171_U8 );
nand NAND2_12689 ( P1_R1171_U250 , P1_R1171_U248 , P1_R1171_U246 );
not NOT1_12690 ( P1_R1171_U251 , P1_R1171_U163 );
or OR2_12691 ( P1_R1171_U252 , P1_U3495 , P1_U3077 );
nand NAND2_12692 ( P1_R1171_U253 , P1_R1171_U252 , P1_R1171_U163 );
nand NAND2_12693 ( P1_R1171_U254 , P1_U3077 , P1_U3495 );
not NOT1_12694 ( P1_R1171_U255 , P1_R1171_U161 );
or OR2_12695 ( P1_R1171_U256 , P1_U3498 , P1_U3072 );
nand NAND2_12696 ( P1_R1171_U257 , P1_R1171_U256 , P1_R1171_U161 );
nand NAND2_12697 ( P1_R1171_U258 , P1_U3072 , P1_U3498 );
not NOT1_12698 ( P1_R1171_U259 , P1_R1171_U93 );
or OR2_12699 ( P1_R1171_U260 , P1_U3067 , P1_U3504 );
or OR2_12700 ( P1_R1171_U261 , P1_U3071 , P1_U3501 );
not NOT1_12701 ( P1_R1171_U262 , P1_R1171_U60 );
nand NAND2_12702 ( P1_R1171_U263 , P1_R1171_U61 , P1_R1171_U60 );
nand NAND2_12703 ( P1_R1171_U264 , P1_U3067 , P1_R1171_U263 );
nand NAND2_12704 ( P1_R1171_U265 , P1_U3504 , P1_R1171_U262 );
nand NAND2_12705 ( P1_R1171_U266 , P1_R1171_U9 , P1_R1171_U93 );
not NOT1_12706 ( P1_R1171_U267 , P1_R1171_U159 );
or OR2_12707 ( P1_R1171_U268 , P1_U3074 , P1_U4015 );
or OR2_12708 ( P1_R1171_U269 , P1_U3079 , P1_U3509 );
or OR2_12709 ( P1_R1171_U270 , P1_U3073 , P1_U4014 );
not NOT1_12710 ( P1_R1171_U271 , P1_R1171_U81 );
nand NAND2_12711 ( P1_R1171_U272 , P1_U4015 , P1_R1171_U271 );
nand NAND2_12712 ( P1_R1171_U273 , P1_R1171_U272 , P1_R1171_U91 );
nand NAND2_12713 ( P1_R1171_U274 , P1_R1171_U81 , P1_R1171_U82 );
nand NAND2_12714 ( P1_R1171_U275 , P1_R1171_U274 , P1_R1171_U273 );
nand NAND2_12715 ( P1_R1171_U276 , P1_R1171_U172 , P1_R1171_U10 );
nand NAND2_12716 ( P1_R1171_U277 , P1_U3073 , P1_U4014 );
nand NAND2_12717 ( P1_R1171_U278 , P1_R1171_U275 , P1_R1171_U276 );
or OR2_12718 ( P1_R1171_U279 , P1_U3507 , P1_U3080 );
or OR2_12719 ( P1_R1171_U280 , P1_U4014 , P1_U3073 );
nand NAND3_12720 ( P1_R1171_U281 , P1_R1171_U270 , P1_R1171_U159 , P1_R1171_U130 );
nand NAND2_12721 ( P1_R1171_U282 , P1_R1171_U280 , P1_R1171_U278 );
not NOT1_12722 ( P1_R1171_U283 , P1_R1171_U155 );
or OR2_12723 ( P1_R1171_U284 , P1_U4013 , P1_U3059 );
nand NAND2_12724 ( P1_R1171_U285 , P1_R1171_U284 , P1_R1171_U155 );
nand NAND2_12725 ( P1_R1171_U286 , P1_U3059 , P1_U4013 );
not NOT1_12726 ( P1_R1171_U287 , P1_R1171_U153 );
or OR2_12727 ( P1_R1171_U288 , P1_U4012 , P1_U3064 );
nand NAND2_12728 ( P1_R1171_U289 , P1_R1171_U288 , P1_R1171_U153 );
nand NAND2_12729 ( P1_R1171_U290 , P1_U3064 , P1_U4012 );
not NOT1_12730 ( P1_R1171_U291 , P1_R1171_U151 );
or OR2_12731 ( P1_R1171_U292 , P1_U3056 , P1_U4010 );
nand NAND2_12732 ( P1_R1171_U293 , P1_R1171_U173 , P1_R1171_U170 );
not NOT1_12733 ( P1_R1171_U294 , P1_R1171_U87 );
or OR2_12734 ( P1_R1171_U295 , P1_U4011 , P1_U3063 );
nand NAND3_12735 ( P1_R1171_U296 , P1_R1171_U151 , P1_R1171_U295 , P1_R1171_U165 );
not NOT1_12736 ( P1_R1171_U297 , P1_R1171_U149 );
or OR2_12737 ( P1_R1171_U298 , P1_U4008 , P1_U3051 );
nand NAND2_12738 ( P1_R1171_U299 , P1_U3051 , P1_U4008 );
not NOT1_12739 ( P1_R1171_U300 , P1_R1171_U147 );
nand NAND2_12740 ( P1_R1171_U301 , P1_U4007 , P1_R1171_U147 );
not NOT1_12741 ( P1_R1171_U302 , P1_R1171_U145 );
nand NAND2_12742 ( P1_R1171_U303 , P1_R1171_U295 , P1_R1171_U151 );
not NOT1_12743 ( P1_R1171_U304 , P1_R1171_U90 );
or OR2_12744 ( P1_R1171_U305 , P1_U4010 , P1_U3056 );
nand NAND2_12745 ( P1_R1171_U306 , P1_R1171_U305 , P1_R1171_U90 );
nand NAND3_12746 ( P1_R1171_U307 , P1_R1171_U306 , P1_R1171_U170 , P1_R1171_U150 );
nand NAND2_12747 ( P1_R1171_U308 , P1_R1171_U304 , P1_R1171_U170 );
nand NAND2_12748 ( P1_R1171_U309 , P1_U4009 , P1_U3055 );
nand NAND3_12749 ( P1_R1171_U310 , P1_R1171_U308 , P1_R1171_U309 , P1_R1171_U165 );
or OR2_12750 ( P1_R1171_U311 , P1_U3056 , P1_U4010 );
nand NAND2_12751 ( P1_R1171_U312 , P1_R1171_U279 , P1_R1171_U159 );
not NOT1_12752 ( P1_R1171_U313 , P1_R1171_U92 );
nand NAND2_12753 ( P1_R1171_U314 , P1_R1171_U10 , P1_R1171_U92 );
nand NAND2_12754 ( P1_R1171_U315 , P1_R1171_U134 , P1_R1171_U314 );
nand NAND2_12755 ( P1_R1171_U316 , P1_R1171_U314 , P1_R1171_U275 );
nand NAND2_12756 ( P1_R1171_U317 , P1_R1171_U450 , P1_R1171_U316 );
or OR2_12757 ( P1_R1171_U318 , P1_U3509 , P1_U3079 );
nand NAND2_12758 ( P1_R1171_U319 , P1_R1171_U318 , P1_R1171_U92 );
nand NAND3_12759 ( P1_R1171_U320 , P1_R1171_U319 , P1_R1171_U81 , P1_R1171_U157 );
nand NAND2_12760 ( P1_R1171_U321 , P1_R1171_U313 , P1_R1171_U81 );
nand NAND2_12761 ( P1_R1171_U322 , P1_U3074 , P1_U4015 );
nand NAND3_12762 ( P1_R1171_U323 , P1_R1171_U322 , P1_R1171_U321 , P1_R1171_U10 );
or OR2_12763 ( P1_R1171_U324 , P1_U3456 , P1_U3076 );
not NOT1_12764 ( P1_R1171_U325 , P1_R1171_U158 );
or OR2_12765 ( P1_R1171_U326 , P1_U3079 , P1_U3509 );
or OR2_12766 ( P1_R1171_U327 , P1_U3501 , P1_U3071 );
nand NAND2_12767 ( P1_R1171_U328 , P1_R1171_U327 , P1_R1171_U93 );
nand NAND2_12768 ( P1_R1171_U329 , P1_R1171_U135 , P1_R1171_U328 );
nand NAND2_12769 ( P1_R1171_U330 , P1_R1171_U259 , P1_R1171_U60 );
nand NAND2_12770 ( P1_R1171_U331 , P1_U3504 , P1_U3067 );
nand NAND3_12771 ( P1_R1171_U332 , P1_R1171_U331 , P1_R1171_U330 , P1_R1171_U9 );
or OR2_12772 ( P1_R1171_U333 , P1_U3071 , P1_U3501 );
nand NAND2_12773 ( P1_R1171_U334 , P1_R1171_U247 , P1_R1171_U164 );
not NOT1_12774 ( P1_R1171_U335 , P1_R1171_U94 );
or OR2_12775 ( P1_R1171_U336 , P1_U3489 , P1_U3070 );
nand NAND2_12776 ( P1_R1171_U337 , P1_R1171_U336 , P1_R1171_U94 );
nand NAND2_12777 ( P1_R1171_U338 , P1_R1171_U136 , P1_R1171_U337 );
nand NAND2_12778 ( P1_R1171_U339 , P1_R1171_U335 , P1_R1171_U169 );
nand NAND2_12779 ( P1_R1171_U340 , P1_U3078 , P1_U3492 );
nand NAND2_12780 ( P1_R1171_U341 , P1_R1171_U137 , P1_R1171_U339 );
or OR2_12781 ( P1_R1171_U342 , P1_U3070 , P1_U3489 );
or OR2_12782 ( P1_R1171_U343 , P1_U3480 , P1_U3081 );
nand NAND2_12783 ( P1_R1171_U344 , P1_R1171_U343 , P1_R1171_U41 );
nand NAND2_12784 ( P1_R1171_U345 , P1_R1171_U138 , P1_R1171_U344 );
nand NAND2_12785 ( P1_R1171_U346 , P1_R1171_U203 , P1_R1171_U168 );
nand NAND2_12786 ( P1_R1171_U347 , P1_U3060 , P1_U3483 );
nand NAND2_12787 ( P1_R1171_U348 , P1_R1171_U139 , P1_R1171_U346 );
nand NAND2_12788 ( P1_R1171_U349 , P1_R1171_U204 , P1_R1171_U168 );
nand NAND2_12789 ( P1_R1171_U350 , P1_R1171_U201 , P1_R1171_U62 );
nand NAND2_12790 ( P1_R1171_U351 , P1_R1171_U211 , P1_R1171_U23 );
nand NAND2_12791 ( P1_R1171_U352 , P1_R1171_U225 , P1_R1171_U35 );
nand NAND2_12792 ( P1_R1171_U353 , P1_R1171_U228 , P1_R1171_U177 );
nand NAND2_12793 ( P1_R1171_U354 , P1_R1171_U311 , P1_R1171_U170 );
nand NAND2_12794 ( P1_R1171_U355 , P1_R1171_U295 , P1_R1171_U173 );
nand NAND2_12795 ( P1_R1171_U356 , P1_R1171_U326 , P1_R1171_U81 );
nand NAND2_12796 ( P1_R1171_U357 , P1_R1171_U279 , P1_R1171_U78 );
nand NAND2_12797 ( P1_R1171_U358 , P1_R1171_U333 , P1_R1171_U60 );
nand NAND2_12798 ( P1_R1171_U359 , P1_R1171_U342 , P1_R1171_U169 );
nand NAND2_12799 ( P1_R1171_U360 , P1_R1171_U247 , P1_R1171_U69 );
nand NAND2_12800 ( P1_R1171_U361 , P1_U4007 , P1_U3052 );
nand NAND2_12801 ( P1_R1171_U362 , P1_R1171_U293 , P1_R1171_U165 );
nand NAND2_12802 ( P1_R1171_U363 , P1_U3055 , P1_R1171_U292 );
nand NAND2_12803 ( P1_R1171_U364 , P1_U4009 , P1_R1171_U292 );
nand NAND3_12804 ( P1_R1171_U365 , P1_R1171_U293 , P1_R1171_U165 , P1_R1171_U298 );
nand NAND3_12805 ( P1_R1171_U366 , P1_R1171_U151 , P1_R1171_U165 , P1_R1171_U132 );
nand NAND2_12806 ( P1_R1171_U367 , P1_R1171_U294 , P1_R1171_U298 );
nand NAND2_12807 ( P1_R1171_U368 , P1_U3081 , P1_R1171_U40 );
nand NAND2_12808 ( P1_R1171_U369 , P1_U3480 , P1_R1171_U39 );
nand NAND2_12809 ( P1_R1171_U370 , P1_R1171_U369 , P1_R1171_U368 );
nand NAND2_12810 ( P1_R1171_U371 , P1_R1171_U349 , P1_R1171_U41 );
nand NAND2_12811 ( P1_R1171_U372 , P1_R1171_U370 , P1_R1171_U203 );
nand NAND2_12812 ( P1_R1171_U373 , P1_U3082 , P1_R1171_U37 );
nand NAND2_12813 ( P1_R1171_U374 , P1_U3477 , P1_R1171_U38 );
nand NAND2_12814 ( P1_R1171_U375 , P1_R1171_U374 , P1_R1171_U373 );
nand NAND2_12815 ( P1_R1171_U376 , P1_R1171_U350 , P1_R1171_U140 );
nand NAND2_12816 ( P1_R1171_U377 , P1_R1171_U200 , P1_R1171_U375 );
nand NAND2_12817 ( P1_R1171_U378 , P1_U3068 , P1_R1171_U24 );
nand NAND2_12818 ( P1_R1171_U379 , P1_U3474 , P1_R1171_U22 );
nand NAND2_12819 ( P1_R1171_U380 , P1_U3069 , P1_R1171_U20 );
nand NAND2_12820 ( P1_R1171_U381 , P1_U3471 , P1_R1171_U21 );
nand NAND2_12821 ( P1_R1171_U382 , P1_R1171_U381 , P1_R1171_U380 );
nand NAND2_12822 ( P1_R1171_U383 , P1_R1171_U351 , P1_R1171_U42 );
nand NAND2_12823 ( P1_R1171_U384 , P1_R1171_U382 , P1_R1171_U192 );
nand NAND2_12824 ( P1_R1171_U385 , P1_U3065 , P1_R1171_U36 );
nand NAND2_12825 ( P1_R1171_U386 , P1_U3468 , P1_R1171_U27 );
nand NAND2_12826 ( P1_R1171_U387 , P1_U3058 , P1_R1171_U25 );
nand NAND2_12827 ( P1_R1171_U388 , P1_U3465 , P1_R1171_U26 );
nand NAND2_12828 ( P1_R1171_U389 , P1_R1171_U388 , P1_R1171_U387 );
nand NAND2_12829 ( P1_R1171_U390 , P1_R1171_U352 , P1_R1171_U45 );
nand NAND2_12830 ( P1_R1171_U391 , P1_R1171_U389 , P1_R1171_U218 );
nand NAND2_12831 ( P1_R1171_U392 , P1_U3062 , P1_R1171_U33 );
nand NAND2_12832 ( P1_R1171_U393 , P1_U3462 , P1_R1171_U34 );
nand NAND2_12833 ( P1_R1171_U394 , P1_R1171_U393 , P1_R1171_U392 );
nand NAND2_12834 ( P1_R1171_U395 , P1_R1171_U353 , P1_R1171_U141 );
nand NAND2_12835 ( P1_R1171_U396 , P1_R1171_U227 , P1_R1171_U394 );
nand NAND2_12836 ( P1_R1171_U397 , P1_U3066 , P1_R1171_U28 );
nand NAND2_12837 ( P1_R1171_U398 , P1_U3459 , P1_R1171_U29 );
nand NAND2_12838 ( P1_R1171_U399 , P1_U3053 , P1_R1171_U143 );
nand NAND2_12839 ( P1_R1171_U400 , P1_U4018 , P1_R1171_U142 );
nand NAND2_12840 ( P1_R1171_U401 , P1_U3053 , P1_R1171_U143 );
nand NAND2_12841 ( P1_R1171_U402 , P1_U4018 , P1_R1171_U142 );
nand NAND2_12842 ( P1_R1171_U403 , P1_R1171_U402 , P1_R1171_U401 );
nand NAND2_12843 ( P1_R1171_U404 , P1_R1171_U144 , P1_R1171_U145 );
nand NAND2_12844 ( P1_R1171_U405 , P1_R1171_U302 , P1_R1171_U403 );
nand NAND2_12845 ( P1_R1171_U406 , P1_U3052 , P1_R1171_U89 );
nand NAND2_12846 ( P1_R1171_U407 , P1_U4007 , P1_R1171_U88 );
nand NAND2_12847 ( P1_R1171_U408 , P1_U3052 , P1_R1171_U89 );
nand NAND2_12848 ( P1_R1171_U409 , P1_U4007 , P1_R1171_U88 );
nand NAND2_12849 ( P1_R1171_U410 , P1_R1171_U409 , P1_R1171_U408 );
nand NAND2_12850 ( P1_R1171_U411 , P1_R1171_U146 , P1_R1171_U147 );
nand NAND2_12851 ( P1_R1171_U412 , P1_R1171_U300 , P1_R1171_U410 );
nand NAND2_12852 ( P1_R1171_U413 , P1_U3051 , P1_R1171_U47 );
nand NAND2_12853 ( P1_R1171_U414 , P1_U4008 , P1_R1171_U48 );
nand NAND2_12854 ( P1_R1171_U415 , P1_U3051 , P1_R1171_U47 );
nand NAND2_12855 ( P1_R1171_U416 , P1_U4008 , P1_R1171_U48 );
nand NAND2_12856 ( P1_R1171_U417 , P1_R1171_U416 , P1_R1171_U415 );
nand NAND2_12857 ( P1_R1171_U418 , P1_R1171_U148 , P1_R1171_U149 );
nand NAND2_12858 ( P1_R1171_U419 , P1_R1171_U297 , P1_R1171_U417 );
nand NAND2_12859 ( P1_R1171_U420 , P1_U3055 , P1_R1171_U50 );
nand NAND2_12860 ( P1_R1171_U421 , P1_U4009 , P1_R1171_U49 );
nand NAND2_12861 ( P1_R1171_U422 , P1_U3056 , P1_R1171_U51 );
nand NAND2_12862 ( P1_R1171_U423 , P1_U4010 , P1_R1171_U52 );
nand NAND2_12863 ( P1_R1171_U424 , P1_R1171_U423 , P1_R1171_U422 );
nand NAND2_12864 ( P1_R1171_U425 , P1_R1171_U354 , P1_R1171_U90 );
nand NAND2_12865 ( P1_R1171_U426 , P1_R1171_U424 , P1_R1171_U304 );
nand NAND2_12866 ( P1_R1171_U427 , P1_U3063 , P1_R1171_U53 );
nand NAND2_12867 ( P1_R1171_U428 , P1_U4011 , P1_R1171_U54 );
nand NAND2_12868 ( P1_R1171_U429 , P1_R1171_U428 , P1_R1171_U427 );
nand NAND2_12869 ( P1_R1171_U430 , P1_R1171_U355 , P1_R1171_U151 );
nand NAND2_12870 ( P1_R1171_U431 , P1_R1171_U291 , P1_R1171_U429 );
nand NAND2_12871 ( P1_R1171_U432 , P1_U3064 , P1_R1171_U85 );
nand NAND2_12872 ( P1_R1171_U433 , P1_U4012 , P1_R1171_U86 );
nand NAND2_12873 ( P1_R1171_U434 , P1_U3064 , P1_R1171_U85 );
nand NAND2_12874 ( P1_R1171_U435 , P1_U4012 , P1_R1171_U86 );
nand NAND2_12875 ( P1_R1171_U436 , P1_R1171_U435 , P1_R1171_U434 );
nand NAND2_12876 ( P1_R1171_U437 , P1_R1171_U152 , P1_R1171_U153 );
nand NAND2_12877 ( P1_R1171_U438 , P1_R1171_U287 , P1_R1171_U436 );
nand NAND2_12878 ( P1_R1171_U439 , P1_U3059 , P1_R1171_U83 );
nand NAND2_12879 ( P1_R1171_U440 , P1_U4013 , P1_R1171_U84 );
nand NAND2_12880 ( P1_R1171_U441 , P1_U3059 , P1_R1171_U83 );
nand NAND2_12881 ( P1_R1171_U442 , P1_U4013 , P1_R1171_U84 );
nand NAND2_12882 ( P1_R1171_U443 , P1_R1171_U442 , P1_R1171_U441 );
nand NAND2_12883 ( P1_R1171_U444 , P1_R1171_U154 , P1_R1171_U155 );
nand NAND2_12884 ( P1_R1171_U445 , P1_R1171_U283 , P1_R1171_U443 );
nand NAND2_12885 ( P1_R1171_U446 , P1_U3073 , P1_R1171_U55 );
nand NAND2_12886 ( P1_R1171_U447 , P1_U4014 , P1_R1171_U56 );
nand NAND2_12887 ( P1_R1171_U448 , P1_U3073 , P1_R1171_U55 );
nand NAND2_12888 ( P1_R1171_U449 , P1_U4014 , P1_R1171_U56 );
nand NAND2_12889 ( P1_R1171_U450 , P1_R1171_U449 , P1_R1171_U448 );
nand NAND2_12890 ( P1_R1171_U451 , P1_U3074 , P1_R1171_U82 );
nand NAND2_12891 ( P1_R1171_U452 , P1_U4015 , P1_R1171_U91 );
nand NAND2_12892 ( P1_R1171_U453 , P1_R1171_U179 , P1_R1171_U158 );
nand NAND2_12893 ( P1_R1171_U454 , P1_R1171_U325 , P1_R1171_U32 );
nand NAND2_12894 ( P1_R1171_U455 , P1_U3079 , P1_R1171_U79 );
nand NAND2_12895 ( P1_R1171_U456 , P1_U3509 , P1_R1171_U80 );
nand NAND2_12896 ( P1_R1171_U457 , P1_R1171_U456 , P1_R1171_U455 );
nand NAND2_12897 ( P1_R1171_U458 , P1_R1171_U356 , P1_R1171_U92 );
nand NAND2_12898 ( P1_R1171_U459 , P1_R1171_U457 , P1_R1171_U313 );
nand NAND2_12899 ( P1_R1171_U460 , P1_U3080 , P1_R1171_U76 );
nand NAND2_12900 ( P1_R1171_U461 , P1_U3507 , P1_R1171_U77 );
nand NAND2_12901 ( P1_R1171_U462 , P1_R1171_U461 , P1_R1171_U460 );
nand NAND2_12902 ( P1_R1171_U463 , P1_R1171_U357 , P1_R1171_U159 );
nand NAND2_12903 ( P1_R1171_U464 , P1_R1171_U267 , P1_R1171_U462 );
nand NAND2_12904 ( P1_R1171_U465 , P1_U3067 , P1_R1171_U61 );
nand NAND2_12905 ( P1_R1171_U466 , P1_U3504 , P1_R1171_U59 );
nand NAND2_12906 ( P1_R1171_U467 , P1_U3071 , P1_R1171_U57 );
nand NAND2_12907 ( P1_R1171_U468 , P1_U3501 , P1_R1171_U58 );
nand NAND2_12908 ( P1_R1171_U469 , P1_R1171_U468 , P1_R1171_U467 );
nand NAND2_12909 ( P1_R1171_U470 , P1_R1171_U358 , P1_R1171_U93 );
nand NAND2_12910 ( P1_R1171_U471 , P1_R1171_U469 , P1_R1171_U259 );
nand NAND2_12911 ( P1_R1171_U472 , P1_U3072 , P1_R1171_U74 );
nand NAND2_12912 ( P1_R1171_U473 , P1_U3498 , P1_R1171_U75 );
nand NAND2_12913 ( P1_R1171_U474 , P1_U3072 , P1_R1171_U74 );
nand NAND2_12914 ( P1_R1171_U475 , P1_U3498 , P1_R1171_U75 );
nand NAND2_12915 ( P1_R1171_U476 , P1_R1171_U475 , P1_R1171_U474 );
nand NAND2_12916 ( P1_R1171_U477 , P1_R1171_U160 , P1_R1171_U161 );
nand NAND2_12917 ( P1_R1171_U478 , P1_R1171_U255 , P1_R1171_U476 );
nand NAND2_12918 ( P1_R1171_U479 , P1_U3077 , P1_R1171_U72 );
nand NAND2_12919 ( P1_R1171_U480 , P1_U3495 , P1_R1171_U73 );
nand NAND2_12920 ( P1_R1171_U481 , P1_U3077 , P1_R1171_U72 );
nand NAND2_12921 ( P1_R1171_U482 , P1_U3495 , P1_R1171_U73 );
nand NAND2_12922 ( P1_R1171_U483 , P1_R1171_U482 , P1_R1171_U481 );
nand NAND2_12923 ( P1_R1171_U484 , P1_R1171_U162 , P1_R1171_U163 );
nand NAND2_12924 ( P1_R1171_U485 , P1_R1171_U251 , P1_R1171_U483 );
nand NAND2_12925 ( P1_R1171_U486 , P1_U3078 , P1_R1171_U70 );
nand NAND2_12926 ( P1_R1171_U487 , P1_U3492 , P1_R1171_U71 );
nand NAND2_12927 ( P1_R1171_U488 , P1_U3070 , P1_R1171_U65 );
nand NAND2_12928 ( P1_R1171_U489 , P1_U3489 , P1_R1171_U66 );
nand NAND2_12929 ( P1_R1171_U490 , P1_R1171_U489 , P1_R1171_U488 );
nand NAND2_12930 ( P1_R1171_U491 , P1_R1171_U359 , P1_R1171_U94 );
nand NAND2_12931 ( P1_R1171_U492 , P1_R1171_U490 , P1_R1171_U335 );
nand NAND2_12932 ( P1_R1171_U493 , P1_U3061 , P1_R1171_U67 );
nand NAND2_12933 ( P1_R1171_U494 , P1_U3486 , P1_R1171_U68 );
nand NAND2_12934 ( P1_R1171_U495 , P1_R1171_U494 , P1_R1171_U493 );
nand NAND2_12935 ( P1_R1171_U496 , P1_R1171_U360 , P1_R1171_U164 );
nand NAND2_12936 ( P1_R1171_U497 , P1_R1171_U241 , P1_R1171_U495 );
nand NAND2_12937 ( P1_R1171_U498 , P1_U3060 , P1_R1171_U63 );
nand NAND2_12938 ( P1_R1171_U499 , P1_U3483 , P1_R1171_U64 );
nand NAND2_12939 ( P1_R1171_U500 , P1_U3075 , P1_R1171_U30 );
nand NAND2_12940 ( P1_R1171_U501 , P1_U3451 , P1_R1171_U31 );
and AND2_12941 ( P1_R1138_U4 , P1_R1138_U176 , P1_R1138_U175 );
and AND2_12942 ( P1_R1138_U5 , P1_R1138_U177 , P1_R1138_U178 );
and AND2_12943 ( P1_R1138_U6 , P1_R1138_U194 , P1_R1138_U193 );
and AND2_12944 ( P1_R1138_U7 , P1_R1138_U234 , P1_R1138_U233 );
and AND2_12945 ( P1_R1138_U8 , P1_R1138_U243 , P1_R1138_U242 );
and AND2_12946 ( P1_R1138_U9 , P1_R1138_U261 , P1_R1138_U260 );
and AND2_12947 ( P1_R1138_U10 , P1_R1138_U269 , P1_R1138_U268 );
and AND2_12948 ( P1_R1138_U11 , P1_R1138_U348 , P1_R1138_U345 );
and AND2_12949 ( P1_R1138_U12 , P1_R1138_U341 , P1_R1138_U338 );
and AND2_12950 ( P1_R1138_U13 , P1_R1138_U332 , P1_R1138_U329 );
and AND2_12951 ( P1_R1138_U14 , P1_R1138_U323 , P1_R1138_U320 );
and AND2_12952 ( P1_R1138_U15 , P1_R1138_U317 , P1_R1138_U315 );
and AND2_12953 ( P1_R1138_U16 , P1_R1138_U310 , P1_R1138_U307 );
and AND2_12954 ( P1_R1138_U17 , P1_R1138_U232 , P1_R1138_U229 );
and AND2_12955 ( P1_R1138_U18 , P1_R1138_U224 , P1_R1138_U221 );
and AND2_12956 ( P1_R1138_U19 , P1_R1138_U210 , P1_R1138_U207 );
not NOT1_12957 ( P1_R1138_U20 , P1_U3471 );
not NOT1_12958 ( P1_R1138_U21 , P1_U3069 );
not NOT1_12959 ( P1_R1138_U22 , P1_U3068 );
nand NAND2_12960 ( P1_R1138_U23 , P1_U3069 , P1_U3471 );
not NOT1_12961 ( P1_R1138_U24 , P1_U3474 );
not NOT1_12962 ( P1_R1138_U25 , P1_U3465 );
not NOT1_12963 ( P1_R1138_U26 , P1_U3058 );
not NOT1_12964 ( P1_R1138_U27 , P1_U3065 );
not NOT1_12965 ( P1_R1138_U28 , P1_U3459 );
not NOT1_12966 ( P1_R1138_U29 , P1_U3066 );
not NOT1_12967 ( P1_R1138_U30 , P1_U3451 );
not NOT1_12968 ( P1_R1138_U31 , P1_U3075 );
nand NAND2_12969 ( P1_R1138_U32 , P1_U3075 , P1_U3451 );
not NOT1_12970 ( P1_R1138_U33 , P1_U3462 );
not NOT1_12971 ( P1_R1138_U34 , P1_U3062 );
nand NAND2_12972 ( P1_R1138_U35 , P1_U3058 , P1_U3465 );
not NOT1_12973 ( P1_R1138_U36 , P1_U3468 );
not NOT1_12974 ( P1_R1138_U37 , P1_U3477 );
not NOT1_12975 ( P1_R1138_U38 , P1_U3082 );
not NOT1_12976 ( P1_R1138_U39 , P1_U3081 );
not NOT1_12977 ( P1_R1138_U40 , P1_U3480 );
nand NAND2_12978 ( P1_R1138_U41 , P1_R1138_U62 , P1_R1138_U202 );
nand NAND2_12979 ( P1_R1138_U42 , P1_R1138_U118 , P1_R1138_U190 );
nand NAND2_12980 ( P1_R1138_U43 , P1_R1138_U179 , P1_R1138_U180 );
nand NAND2_12981 ( P1_R1138_U44 , P1_U3456 , P1_U3076 );
nand NAND2_12982 ( P1_R1138_U45 , P1_R1138_U122 , P1_R1138_U216 );
nand NAND2_12983 ( P1_R1138_U46 , P1_R1138_U213 , P1_R1138_U212 );
not NOT1_12984 ( P1_R1138_U47 , P1_U4008 );
not NOT1_12985 ( P1_R1138_U48 , P1_U3051 );
not NOT1_12986 ( P1_R1138_U49 , P1_U3055 );
not NOT1_12987 ( P1_R1138_U50 , P1_U4009 );
not NOT1_12988 ( P1_R1138_U51 , P1_U4010 );
not NOT1_12989 ( P1_R1138_U52 , P1_U3056 );
not NOT1_12990 ( P1_R1138_U53 , P1_U4011 );
not NOT1_12991 ( P1_R1138_U54 , P1_U3063 );
not NOT1_12992 ( P1_R1138_U55 , P1_U4014 );
not NOT1_12993 ( P1_R1138_U56 , P1_U3073 );
not NOT1_12994 ( P1_R1138_U57 , P1_U3501 );
not NOT1_12995 ( P1_R1138_U58 , P1_U3071 );
not NOT1_12996 ( P1_R1138_U59 , P1_U3067 );
nand NAND2_12997 ( P1_R1138_U60 , P1_U3071 , P1_U3501 );
not NOT1_12998 ( P1_R1138_U61 , P1_U3504 );
nand NAND2_12999 ( P1_R1138_U62 , P1_U3082 , P1_U3477 );
not NOT1_13000 ( P1_R1138_U63 , P1_U3483 );
not NOT1_13001 ( P1_R1138_U64 , P1_U3060 );
not NOT1_13002 ( P1_R1138_U65 , P1_U3489 );
not NOT1_13003 ( P1_R1138_U66 , P1_U3070 );
not NOT1_13004 ( P1_R1138_U67 , P1_U3486 );
not NOT1_13005 ( P1_R1138_U68 , P1_U3061 );
nand NAND2_13006 ( P1_R1138_U69 , P1_U3061 , P1_U3486 );
not NOT1_13007 ( P1_R1138_U70 , P1_U3492 );
not NOT1_13008 ( P1_R1138_U71 , P1_U3078 );
not NOT1_13009 ( P1_R1138_U72 , P1_U3495 );
not NOT1_13010 ( P1_R1138_U73 , P1_U3077 );
not NOT1_13011 ( P1_R1138_U74 , P1_U3498 );
not NOT1_13012 ( P1_R1138_U75 , P1_U3072 );
not NOT1_13013 ( P1_R1138_U76 , P1_U3507 );
not NOT1_13014 ( P1_R1138_U77 , P1_U3080 );
nand NAND2_13015 ( P1_R1138_U78 , P1_U3080 , P1_U3507 );
not NOT1_13016 ( P1_R1138_U79 , P1_U3509 );
not NOT1_13017 ( P1_R1138_U80 , P1_U3079 );
nand NAND2_13018 ( P1_R1138_U81 , P1_U3079 , P1_U3509 );
not NOT1_13019 ( P1_R1138_U82 , P1_U4015 );
not NOT1_13020 ( P1_R1138_U83 , P1_U4013 );
not NOT1_13021 ( P1_R1138_U84 , P1_U3059 );
not NOT1_13022 ( P1_R1138_U85 , P1_U4012 );
not NOT1_13023 ( P1_R1138_U86 , P1_U3064 );
nand NAND2_13024 ( P1_R1138_U87 , P1_U4009 , P1_U3055 );
not NOT1_13025 ( P1_R1138_U88 , P1_U3052 );
not NOT1_13026 ( P1_R1138_U89 , P1_U4007 );
nand NAND2_13027 ( P1_R1138_U90 , P1_R1138_U303 , P1_R1138_U173 );
not NOT1_13028 ( P1_R1138_U91 , P1_U3074 );
nand NAND2_13029 ( P1_R1138_U92 , P1_R1138_U78 , P1_R1138_U312 );
nand NAND2_13030 ( P1_R1138_U93 , P1_R1138_U258 , P1_R1138_U257 );
nand NAND2_13031 ( P1_R1138_U94 , P1_R1138_U69 , P1_R1138_U334 );
nand NAND2_13032 ( P1_R1138_U95 , P1_R1138_U454 , P1_R1138_U453 );
nand NAND2_13033 ( P1_R1138_U96 , P1_R1138_U501 , P1_R1138_U500 );
nand NAND2_13034 ( P1_R1138_U97 , P1_R1138_U372 , P1_R1138_U371 );
nand NAND2_13035 ( P1_R1138_U98 , P1_R1138_U377 , P1_R1138_U376 );
nand NAND2_13036 ( P1_R1138_U99 , P1_R1138_U384 , P1_R1138_U383 );
nand NAND2_13037 ( P1_R1138_U100 , P1_R1138_U391 , P1_R1138_U390 );
nand NAND2_13038 ( P1_R1138_U101 , P1_R1138_U396 , P1_R1138_U395 );
nand NAND2_13039 ( P1_R1138_U102 , P1_R1138_U405 , P1_R1138_U404 );
nand NAND2_13040 ( P1_R1138_U103 , P1_R1138_U412 , P1_R1138_U411 );
nand NAND2_13041 ( P1_R1138_U104 , P1_R1138_U419 , P1_R1138_U418 );
nand NAND2_13042 ( P1_R1138_U105 , P1_R1138_U426 , P1_R1138_U425 );
nand NAND2_13043 ( P1_R1138_U106 , P1_R1138_U431 , P1_R1138_U430 );
nand NAND2_13044 ( P1_R1138_U107 , P1_R1138_U438 , P1_R1138_U437 );
nand NAND2_13045 ( P1_R1138_U108 , P1_R1138_U445 , P1_R1138_U444 );
nand NAND2_13046 ( P1_R1138_U109 , P1_R1138_U459 , P1_R1138_U458 );
nand NAND2_13047 ( P1_R1138_U110 , P1_R1138_U464 , P1_R1138_U463 );
nand NAND2_13048 ( P1_R1138_U111 , P1_R1138_U471 , P1_R1138_U470 );
nand NAND2_13049 ( P1_R1138_U112 , P1_R1138_U478 , P1_R1138_U477 );
nand NAND2_13050 ( P1_R1138_U113 , P1_R1138_U485 , P1_R1138_U484 );
nand NAND2_13051 ( P1_R1138_U114 , P1_R1138_U492 , P1_R1138_U491 );
nand NAND2_13052 ( P1_R1138_U115 , P1_R1138_U497 , P1_R1138_U496 );
and AND2_13053 ( P1_R1138_U116 , P1_U3459 , P1_U3066 );
and AND2_13054 ( P1_R1138_U117 , P1_R1138_U186 , P1_R1138_U184 );
and AND2_13055 ( P1_R1138_U118 , P1_R1138_U191 , P1_R1138_U189 );
and AND2_13056 ( P1_R1138_U119 , P1_R1138_U198 , P1_R1138_U197 );
and AND3_13057 ( P1_R1138_U120 , P1_R1138_U379 , P1_R1138_U378 , P1_R1138_U23 );
and AND2_13058 ( P1_R1138_U121 , P1_R1138_U209 , P1_R1138_U6 );
and AND2_13059 ( P1_R1138_U122 , P1_R1138_U217 , P1_R1138_U215 );
and AND3_13060 ( P1_R1138_U123 , P1_R1138_U386 , P1_R1138_U385 , P1_R1138_U35 );
and AND2_13061 ( P1_R1138_U124 , P1_R1138_U223 , P1_R1138_U4 );
and AND2_13062 ( P1_R1138_U125 , P1_R1138_U231 , P1_R1138_U178 );
and AND2_13063 ( P1_R1138_U126 , P1_R1138_U201 , P1_R1138_U7 );
and AND2_13064 ( P1_R1138_U127 , P1_R1138_U236 , P1_R1138_U168 );
and AND2_13065 ( P1_R1138_U128 , P1_R1138_U245 , P1_R1138_U169 );
and AND2_13066 ( P1_R1138_U129 , P1_R1138_U265 , P1_R1138_U264 );
and AND2_13067 ( P1_R1138_U130 , P1_R1138_U10 , P1_R1138_U279 );
and AND2_13068 ( P1_R1138_U131 , P1_R1138_U282 , P1_R1138_U277 );
and AND2_13069 ( P1_R1138_U132 , P1_R1138_U298 , P1_R1138_U295 );
and AND2_13070 ( P1_R1138_U133 , P1_R1138_U365 , P1_R1138_U299 );
and AND2_13071 ( P1_R1138_U134 , P1_R1138_U156 , P1_R1138_U275 );
and AND3_13072 ( P1_R1138_U135 , P1_R1138_U466 , P1_R1138_U465 , P1_R1138_U60 );
and AND3_13073 ( P1_R1138_U136 , P1_R1138_U487 , P1_R1138_U486 , P1_R1138_U169 );
and AND2_13074 ( P1_R1138_U137 , P1_R1138_U340 , P1_R1138_U8 );
and AND3_13075 ( P1_R1138_U138 , P1_R1138_U499 , P1_R1138_U498 , P1_R1138_U168 );
and AND2_13076 ( P1_R1138_U139 , P1_R1138_U347 , P1_R1138_U7 );
nand NAND2_13077 ( P1_R1138_U140 , P1_R1138_U119 , P1_R1138_U199 );
nand NAND2_13078 ( P1_R1138_U141 , P1_R1138_U214 , P1_R1138_U226 );
not NOT1_13079 ( P1_R1138_U142 , P1_U3053 );
not NOT1_13080 ( P1_R1138_U143 , P1_U4018 );
and AND2_13081 ( P1_R1138_U144 , P1_R1138_U400 , P1_R1138_U399 );
nand NAND3_13082 ( P1_R1138_U145 , P1_R1138_U301 , P1_R1138_U166 , P1_R1138_U361 );
and AND2_13083 ( P1_R1138_U146 , P1_R1138_U407 , P1_R1138_U406 );
nand NAND3_13084 ( P1_R1138_U147 , P1_R1138_U367 , P1_R1138_U366 , P1_R1138_U133 );
and AND2_13085 ( P1_R1138_U148 , P1_R1138_U414 , P1_R1138_U413 );
nand NAND3_13086 ( P1_R1138_U149 , P1_R1138_U362 , P1_R1138_U296 , P1_R1138_U87 );
and AND2_13087 ( P1_R1138_U150 , P1_R1138_U421 , P1_R1138_U420 );
nand NAND2_13088 ( P1_R1138_U151 , P1_R1138_U290 , P1_R1138_U289 );
and AND2_13089 ( P1_R1138_U152 , P1_R1138_U433 , P1_R1138_U432 );
nand NAND2_13090 ( P1_R1138_U153 , P1_R1138_U286 , P1_R1138_U285 );
and AND2_13091 ( P1_R1138_U154 , P1_R1138_U440 , P1_R1138_U439 );
nand NAND2_13092 ( P1_R1138_U155 , P1_R1138_U131 , P1_R1138_U281 );
and AND2_13093 ( P1_R1138_U156 , P1_R1138_U447 , P1_R1138_U446 );
and AND2_13094 ( P1_R1138_U157 , P1_R1138_U452 , P1_R1138_U451 );
nand NAND2_13095 ( P1_R1138_U158 , P1_R1138_U44 , P1_R1138_U324 );
nand NAND2_13096 ( P1_R1138_U159 , P1_R1138_U129 , P1_R1138_U266 );
and AND2_13097 ( P1_R1138_U160 , P1_R1138_U473 , P1_R1138_U472 );
nand NAND2_13098 ( P1_R1138_U161 , P1_R1138_U254 , P1_R1138_U253 );
and AND2_13099 ( P1_R1138_U162 , P1_R1138_U480 , P1_R1138_U479 );
nand NAND2_13100 ( P1_R1138_U163 , P1_R1138_U250 , P1_R1138_U249 );
nand NAND2_13101 ( P1_R1138_U164 , P1_R1138_U240 , P1_R1138_U239 );
nand NAND2_13102 ( P1_R1138_U165 , P1_R1138_U364 , P1_R1138_U363 );
nand NAND2_13103 ( P1_R1138_U166 , P1_U3052 , P1_R1138_U147 );
not NOT1_13104 ( P1_R1138_U167 , P1_R1138_U35 );
nand NAND2_13105 ( P1_R1138_U168 , P1_U3480 , P1_U3081 );
nand NAND2_13106 ( P1_R1138_U169 , P1_U3070 , P1_U3489 );
nand NAND2_13107 ( P1_R1138_U170 , P1_U3056 , P1_U4010 );
not NOT1_13108 ( P1_R1138_U171 , P1_R1138_U69 );
not NOT1_13109 ( P1_R1138_U172 , P1_R1138_U78 );
nand NAND2_13110 ( P1_R1138_U173 , P1_U3063 , P1_U4011 );
not NOT1_13111 ( P1_R1138_U174 , P1_R1138_U62 );
or OR2_13112 ( P1_R1138_U175 , P1_U3065 , P1_U3468 );
or OR2_13113 ( P1_R1138_U176 , P1_U3058 , P1_U3465 );
or OR2_13114 ( P1_R1138_U177 , P1_U3462 , P1_U3062 );
or OR2_13115 ( P1_R1138_U178 , P1_U3459 , P1_U3066 );
not NOT1_13116 ( P1_R1138_U179 , P1_R1138_U32 );
or OR2_13117 ( P1_R1138_U180 , P1_U3456 , P1_U3076 );
not NOT1_13118 ( P1_R1138_U181 , P1_R1138_U43 );
not NOT1_13119 ( P1_R1138_U182 , P1_R1138_U44 );
nand NAND2_13120 ( P1_R1138_U183 , P1_R1138_U43 , P1_R1138_U44 );
nand NAND2_13121 ( P1_R1138_U184 , P1_R1138_U116 , P1_R1138_U177 );
nand NAND2_13122 ( P1_R1138_U185 , P1_R1138_U5 , P1_R1138_U183 );
nand NAND2_13123 ( P1_R1138_U186 , P1_U3062 , P1_U3462 );
nand NAND2_13124 ( P1_R1138_U187 , P1_R1138_U117 , P1_R1138_U185 );
nand NAND2_13125 ( P1_R1138_U188 , P1_R1138_U36 , P1_R1138_U35 );
nand NAND2_13126 ( P1_R1138_U189 , P1_U3065 , P1_R1138_U188 );
nand NAND2_13127 ( P1_R1138_U190 , P1_R1138_U4 , P1_R1138_U187 );
nand NAND2_13128 ( P1_R1138_U191 , P1_U3468 , P1_R1138_U167 );
not NOT1_13129 ( P1_R1138_U192 , P1_R1138_U42 );
or OR2_13130 ( P1_R1138_U193 , P1_U3068 , P1_U3474 );
or OR2_13131 ( P1_R1138_U194 , P1_U3069 , P1_U3471 );
not NOT1_13132 ( P1_R1138_U195 , P1_R1138_U23 );
nand NAND2_13133 ( P1_R1138_U196 , P1_R1138_U24 , P1_R1138_U23 );
nand NAND2_13134 ( P1_R1138_U197 , P1_U3068 , P1_R1138_U196 );
nand NAND2_13135 ( P1_R1138_U198 , P1_U3474 , P1_R1138_U195 );
nand NAND2_13136 ( P1_R1138_U199 , P1_R1138_U6 , P1_R1138_U42 );
not NOT1_13137 ( P1_R1138_U200 , P1_R1138_U140 );
or OR2_13138 ( P1_R1138_U201 , P1_U3477 , P1_U3082 );
nand NAND2_13139 ( P1_R1138_U202 , P1_R1138_U201 , P1_R1138_U140 );
not NOT1_13140 ( P1_R1138_U203 , P1_R1138_U41 );
or OR2_13141 ( P1_R1138_U204 , P1_U3081 , P1_U3480 );
or OR2_13142 ( P1_R1138_U205 , P1_U3471 , P1_U3069 );
nand NAND2_13143 ( P1_R1138_U206 , P1_R1138_U205 , P1_R1138_U42 );
nand NAND2_13144 ( P1_R1138_U207 , P1_R1138_U120 , P1_R1138_U206 );
nand NAND2_13145 ( P1_R1138_U208 , P1_R1138_U192 , P1_R1138_U23 );
nand NAND2_13146 ( P1_R1138_U209 , P1_U3474 , P1_U3068 );
nand NAND2_13147 ( P1_R1138_U210 , P1_R1138_U121 , P1_R1138_U208 );
or OR2_13148 ( P1_R1138_U211 , P1_U3069 , P1_U3471 );
nand NAND2_13149 ( P1_R1138_U212 , P1_R1138_U182 , P1_R1138_U178 );
nand NAND2_13150 ( P1_R1138_U213 , P1_U3066 , P1_U3459 );
not NOT1_13151 ( P1_R1138_U214 , P1_R1138_U46 );
nand NAND2_13152 ( P1_R1138_U215 , P1_R1138_U181 , P1_R1138_U5 );
nand NAND2_13153 ( P1_R1138_U216 , P1_R1138_U46 , P1_R1138_U177 );
nand NAND2_13154 ( P1_R1138_U217 , P1_U3062 , P1_U3462 );
not NOT1_13155 ( P1_R1138_U218 , P1_R1138_U45 );
or OR2_13156 ( P1_R1138_U219 , P1_U3465 , P1_U3058 );
nand NAND2_13157 ( P1_R1138_U220 , P1_R1138_U219 , P1_R1138_U45 );
nand NAND2_13158 ( P1_R1138_U221 , P1_R1138_U123 , P1_R1138_U220 );
nand NAND2_13159 ( P1_R1138_U222 , P1_R1138_U218 , P1_R1138_U35 );
nand NAND2_13160 ( P1_R1138_U223 , P1_U3468 , P1_U3065 );
nand NAND2_13161 ( P1_R1138_U224 , P1_R1138_U124 , P1_R1138_U222 );
or OR2_13162 ( P1_R1138_U225 , P1_U3058 , P1_U3465 );
nand NAND2_13163 ( P1_R1138_U226 , P1_R1138_U181 , P1_R1138_U178 );
not NOT1_13164 ( P1_R1138_U227 , P1_R1138_U141 );
nand NAND2_13165 ( P1_R1138_U228 , P1_U3062 , P1_U3462 );
nand NAND4_13166 ( P1_R1138_U229 , P1_R1138_U398 , P1_R1138_U397 , P1_R1138_U44 , P1_R1138_U43 );
nand NAND2_13167 ( P1_R1138_U230 , P1_R1138_U44 , P1_R1138_U43 );
nand NAND2_13168 ( P1_R1138_U231 , P1_U3066 , P1_U3459 );
nand NAND2_13169 ( P1_R1138_U232 , P1_R1138_U125 , P1_R1138_U230 );
or OR2_13170 ( P1_R1138_U233 , P1_U3081 , P1_U3480 );
or OR2_13171 ( P1_R1138_U234 , P1_U3060 , P1_U3483 );
nand NAND2_13172 ( P1_R1138_U235 , P1_R1138_U174 , P1_R1138_U7 );
nand NAND2_13173 ( P1_R1138_U236 , P1_U3060 , P1_U3483 );
nand NAND2_13174 ( P1_R1138_U237 , P1_R1138_U127 , P1_R1138_U235 );
or OR2_13175 ( P1_R1138_U238 , P1_U3483 , P1_U3060 );
nand NAND2_13176 ( P1_R1138_U239 , P1_R1138_U126 , P1_R1138_U140 );
nand NAND2_13177 ( P1_R1138_U240 , P1_R1138_U238 , P1_R1138_U237 );
not NOT1_13178 ( P1_R1138_U241 , P1_R1138_U164 );
or OR2_13179 ( P1_R1138_U242 , P1_U3078 , P1_U3492 );
or OR2_13180 ( P1_R1138_U243 , P1_U3070 , P1_U3489 );
nand NAND2_13181 ( P1_R1138_U244 , P1_R1138_U171 , P1_R1138_U8 );
nand NAND2_13182 ( P1_R1138_U245 , P1_U3078 , P1_U3492 );
nand NAND2_13183 ( P1_R1138_U246 , P1_R1138_U128 , P1_R1138_U244 );
or OR2_13184 ( P1_R1138_U247 , P1_U3486 , P1_U3061 );
or OR2_13185 ( P1_R1138_U248 , P1_U3492 , P1_U3078 );
nand NAND3_13186 ( P1_R1138_U249 , P1_R1138_U247 , P1_R1138_U164 , P1_R1138_U8 );
nand NAND2_13187 ( P1_R1138_U250 , P1_R1138_U248 , P1_R1138_U246 );
not NOT1_13188 ( P1_R1138_U251 , P1_R1138_U163 );
or OR2_13189 ( P1_R1138_U252 , P1_U3495 , P1_U3077 );
nand NAND2_13190 ( P1_R1138_U253 , P1_R1138_U252 , P1_R1138_U163 );
nand NAND2_13191 ( P1_R1138_U254 , P1_U3077 , P1_U3495 );
not NOT1_13192 ( P1_R1138_U255 , P1_R1138_U161 );
or OR2_13193 ( P1_R1138_U256 , P1_U3498 , P1_U3072 );
nand NAND2_13194 ( P1_R1138_U257 , P1_R1138_U256 , P1_R1138_U161 );
nand NAND2_13195 ( P1_R1138_U258 , P1_U3072 , P1_U3498 );
not NOT1_13196 ( P1_R1138_U259 , P1_R1138_U93 );
or OR2_13197 ( P1_R1138_U260 , P1_U3067 , P1_U3504 );
or OR2_13198 ( P1_R1138_U261 , P1_U3071 , P1_U3501 );
not NOT1_13199 ( P1_R1138_U262 , P1_R1138_U60 );
nand NAND2_13200 ( P1_R1138_U263 , P1_R1138_U61 , P1_R1138_U60 );
nand NAND2_13201 ( P1_R1138_U264 , P1_U3067 , P1_R1138_U263 );
nand NAND2_13202 ( P1_R1138_U265 , P1_U3504 , P1_R1138_U262 );
nand NAND2_13203 ( P1_R1138_U266 , P1_R1138_U9 , P1_R1138_U93 );
not NOT1_13204 ( P1_R1138_U267 , P1_R1138_U159 );
or OR2_13205 ( P1_R1138_U268 , P1_U3074 , P1_U4015 );
or OR2_13206 ( P1_R1138_U269 , P1_U3079 , P1_U3509 );
or OR2_13207 ( P1_R1138_U270 , P1_U3073 , P1_U4014 );
not NOT1_13208 ( P1_R1138_U271 , P1_R1138_U81 );
nand NAND2_13209 ( P1_R1138_U272 , P1_U4015 , P1_R1138_U271 );
nand NAND2_13210 ( P1_R1138_U273 , P1_R1138_U272 , P1_R1138_U91 );
nand NAND2_13211 ( P1_R1138_U274 , P1_R1138_U81 , P1_R1138_U82 );
nand NAND2_13212 ( P1_R1138_U275 , P1_R1138_U274 , P1_R1138_U273 );
nand NAND2_13213 ( P1_R1138_U276 , P1_R1138_U172 , P1_R1138_U10 );
nand NAND2_13214 ( P1_R1138_U277 , P1_U3073 , P1_U4014 );
nand NAND2_13215 ( P1_R1138_U278 , P1_R1138_U275 , P1_R1138_U276 );
or OR2_13216 ( P1_R1138_U279 , P1_U3507 , P1_U3080 );
or OR2_13217 ( P1_R1138_U280 , P1_U4014 , P1_U3073 );
nand NAND3_13218 ( P1_R1138_U281 , P1_R1138_U270 , P1_R1138_U159 , P1_R1138_U130 );
nand NAND2_13219 ( P1_R1138_U282 , P1_R1138_U280 , P1_R1138_U278 );
not NOT1_13220 ( P1_R1138_U283 , P1_R1138_U155 );
or OR2_13221 ( P1_R1138_U284 , P1_U4013 , P1_U3059 );
nand NAND2_13222 ( P1_R1138_U285 , P1_R1138_U284 , P1_R1138_U155 );
nand NAND2_13223 ( P1_R1138_U286 , P1_U3059 , P1_U4013 );
not NOT1_13224 ( P1_R1138_U287 , P1_R1138_U153 );
or OR2_13225 ( P1_R1138_U288 , P1_U4012 , P1_U3064 );
nand NAND2_13226 ( P1_R1138_U289 , P1_R1138_U288 , P1_R1138_U153 );
nand NAND2_13227 ( P1_R1138_U290 , P1_U3064 , P1_U4012 );
not NOT1_13228 ( P1_R1138_U291 , P1_R1138_U151 );
or OR2_13229 ( P1_R1138_U292 , P1_U3056 , P1_U4010 );
nand NAND2_13230 ( P1_R1138_U293 , P1_R1138_U173 , P1_R1138_U170 );
not NOT1_13231 ( P1_R1138_U294 , P1_R1138_U87 );
or OR2_13232 ( P1_R1138_U295 , P1_U4011 , P1_U3063 );
nand NAND3_13233 ( P1_R1138_U296 , P1_R1138_U151 , P1_R1138_U295 , P1_R1138_U165 );
not NOT1_13234 ( P1_R1138_U297 , P1_R1138_U149 );
or OR2_13235 ( P1_R1138_U298 , P1_U4008 , P1_U3051 );
nand NAND2_13236 ( P1_R1138_U299 , P1_U3051 , P1_U4008 );
not NOT1_13237 ( P1_R1138_U300 , P1_R1138_U147 );
nand NAND2_13238 ( P1_R1138_U301 , P1_U4007 , P1_R1138_U147 );
not NOT1_13239 ( P1_R1138_U302 , P1_R1138_U145 );
nand NAND2_13240 ( P1_R1138_U303 , P1_R1138_U295 , P1_R1138_U151 );
not NOT1_13241 ( P1_R1138_U304 , P1_R1138_U90 );
or OR2_13242 ( P1_R1138_U305 , P1_U4010 , P1_U3056 );
nand NAND2_13243 ( P1_R1138_U306 , P1_R1138_U305 , P1_R1138_U90 );
nand NAND3_13244 ( P1_R1138_U307 , P1_R1138_U306 , P1_R1138_U170 , P1_R1138_U150 );
nand NAND2_13245 ( P1_R1138_U308 , P1_R1138_U304 , P1_R1138_U170 );
nand NAND2_13246 ( P1_R1138_U309 , P1_U4009 , P1_U3055 );
nand NAND3_13247 ( P1_R1138_U310 , P1_R1138_U308 , P1_R1138_U309 , P1_R1138_U165 );
or OR2_13248 ( P1_R1138_U311 , P1_U3056 , P1_U4010 );
nand NAND2_13249 ( P1_R1138_U312 , P1_R1138_U279 , P1_R1138_U159 );
not NOT1_13250 ( P1_R1138_U313 , P1_R1138_U92 );
nand NAND2_13251 ( P1_R1138_U314 , P1_R1138_U10 , P1_R1138_U92 );
nand NAND2_13252 ( P1_R1138_U315 , P1_R1138_U134 , P1_R1138_U314 );
nand NAND2_13253 ( P1_R1138_U316 , P1_R1138_U314 , P1_R1138_U275 );
nand NAND2_13254 ( P1_R1138_U317 , P1_R1138_U450 , P1_R1138_U316 );
or OR2_13255 ( P1_R1138_U318 , P1_U3509 , P1_U3079 );
nand NAND2_13256 ( P1_R1138_U319 , P1_R1138_U318 , P1_R1138_U92 );
nand NAND3_13257 ( P1_R1138_U320 , P1_R1138_U319 , P1_R1138_U81 , P1_R1138_U157 );
nand NAND2_13258 ( P1_R1138_U321 , P1_R1138_U313 , P1_R1138_U81 );
nand NAND2_13259 ( P1_R1138_U322 , P1_U3074 , P1_U4015 );
nand NAND3_13260 ( P1_R1138_U323 , P1_R1138_U322 , P1_R1138_U321 , P1_R1138_U10 );
or OR2_13261 ( P1_R1138_U324 , P1_U3456 , P1_U3076 );
not NOT1_13262 ( P1_R1138_U325 , P1_R1138_U158 );
or OR2_13263 ( P1_R1138_U326 , P1_U3079 , P1_U3509 );
or OR2_13264 ( P1_R1138_U327 , P1_U3501 , P1_U3071 );
nand NAND2_13265 ( P1_R1138_U328 , P1_R1138_U327 , P1_R1138_U93 );
nand NAND2_13266 ( P1_R1138_U329 , P1_R1138_U135 , P1_R1138_U328 );
nand NAND2_13267 ( P1_R1138_U330 , P1_R1138_U259 , P1_R1138_U60 );
nand NAND2_13268 ( P1_R1138_U331 , P1_U3504 , P1_U3067 );
nand NAND3_13269 ( P1_R1138_U332 , P1_R1138_U331 , P1_R1138_U330 , P1_R1138_U9 );
or OR2_13270 ( P1_R1138_U333 , P1_U3071 , P1_U3501 );
nand NAND2_13271 ( P1_R1138_U334 , P1_R1138_U247 , P1_R1138_U164 );
not NOT1_13272 ( P1_R1138_U335 , P1_R1138_U94 );
or OR2_13273 ( P1_R1138_U336 , P1_U3489 , P1_U3070 );
nand NAND2_13274 ( P1_R1138_U337 , P1_R1138_U336 , P1_R1138_U94 );
nand NAND2_13275 ( P1_R1138_U338 , P1_R1138_U136 , P1_R1138_U337 );
nand NAND2_13276 ( P1_R1138_U339 , P1_R1138_U335 , P1_R1138_U169 );
nand NAND2_13277 ( P1_R1138_U340 , P1_U3078 , P1_U3492 );
nand NAND2_13278 ( P1_R1138_U341 , P1_R1138_U137 , P1_R1138_U339 );
or OR2_13279 ( P1_R1138_U342 , P1_U3070 , P1_U3489 );
or OR2_13280 ( P1_R1138_U343 , P1_U3480 , P1_U3081 );
nand NAND2_13281 ( P1_R1138_U344 , P1_R1138_U343 , P1_R1138_U41 );
nand NAND2_13282 ( P1_R1138_U345 , P1_R1138_U138 , P1_R1138_U344 );
nand NAND2_13283 ( P1_R1138_U346 , P1_R1138_U203 , P1_R1138_U168 );
nand NAND2_13284 ( P1_R1138_U347 , P1_U3060 , P1_U3483 );
nand NAND2_13285 ( P1_R1138_U348 , P1_R1138_U139 , P1_R1138_U346 );
nand NAND2_13286 ( P1_R1138_U349 , P1_R1138_U204 , P1_R1138_U168 );
nand NAND2_13287 ( P1_R1138_U350 , P1_R1138_U201 , P1_R1138_U62 );
nand NAND2_13288 ( P1_R1138_U351 , P1_R1138_U211 , P1_R1138_U23 );
nand NAND2_13289 ( P1_R1138_U352 , P1_R1138_U225 , P1_R1138_U35 );
nand NAND2_13290 ( P1_R1138_U353 , P1_R1138_U228 , P1_R1138_U177 );
nand NAND2_13291 ( P1_R1138_U354 , P1_R1138_U311 , P1_R1138_U170 );
nand NAND2_13292 ( P1_R1138_U355 , P1_R1138_U295 , P1_R1138_U173 );
nand NAND2_13293 ( P1_R1138_U356 , P1_R1138_U326 , P1_R1138_U81 );
nand NAND2_13294 ( P1_R1138_U357 , P1_R1138_U279 , P1_R1138_U78 );
nand NAND2_13295 ( P1_R1138_U358 , P1_R1138_U333 , P1_R1138_U60 );
nand NAND2_13296 ( P1_R1138_U359 , P1_R1138_U342 , P1_R1138_U169 );
nand NAND2_13297 ( P1_R1138_U360 , P1_R1138_U247 , P1_R1138_U69 );
nand NAND2_13298 ( P1_R1138_U361 , P1_U4007 , P1_U3052 );
nand NAND2_13299 ( P1_R1138_U362 , P1_R1138_U293 , P1_R1138_U165 );
nand NAND2_13300 ( P1_R1138_U363 , P1_U3055 , P1_R1138_U292 );
nand NAND2_13301 ( P1_R1138_U364 , P1_U4009 , P1_R1138_U292 );
nand NAND3_13302 ( P1_R1138_U365 , P1_R1138_U293 , P1_R1138_U165 , P1_R1138_U298 );
nand NAND3_13303 ( P1_R1138_U366 , P1_R1138_U151 , P1_R1138_U165 , P1_R1138_U132 );
nand NAND2_13304 ( P1_R1138_U367 , P1_R1138_U294 , P1_R1138_U298 );
nand NAND2_13305 ( P1_R1138_U368 , P1_U3081 , P1_R1138_U40 );
nand NAND2_13306 ( P1_R1138_U369 , P1_U3480 , P1_R1138_U39 );
nand NAND2_13307 ( P1_R1138_U370 , P1_R1138_U369 , P1_R1138_U368 );
nand NAND2_13308 ( P1_R1138_U371 , P1_R1138_U349 , P1_R1138_U41 );
nand NAND2_13309 ( P1_R1138_U372 , P1_R1138_U370 , P1_R1138_U203 );
nand NAND2_13310 ( P1_R1138_U373 , P1_U3082 , P1_R1138_U37 );
nand NAND2_13311 ( P1_R1138_U374 , P1_U3477 , P1_R1138_U38 );
nand NAND2_13312 ( P1_R1138_U375 , P1_R1138_U374 , P1_R1138_U373 );
nand NAND2_13313 ( P1_R1138_U376 , P1_R1138_U350 , P1_R1138_U140 );
nand NAND2_13314 ( P1_R1138_U377 , P1_R1138_U200 , P1_R1138_U375 );
nand NAND2_13315 ( P1_R1138_U378 , P1_U3068 , P1_R1138_U24 );
nand NAND2_13316 ( P1_R1138_U379 , P1_U3474 , P1_R1138_U22 );
nand NAND2_13317 ( P1_R1138_U380 , P1_U3069 , P1_R1138_U20 );
nand NAND2_13318 ( P1_R1138_U381 , P1_U3471 , P1_R1138_U21 );
nand NAND2_13319 ( P1_R1138_U382 , P1_R1138_U381 , P1_R1138_U380 );
nand NAND2_13320 ( P1_R1138_U383 , P1_R1138_U351 , P1_R1138_U42 );
nand NAND2_13321 ( P1_R1138_U384 , P1_R1138_U382 , P1_R1138_U192 );
nand NAND2_13322 ( P1_R1138_U385 , P1_U3065 , P1_R1138_U36 );
nand NAND2_13323 ( P1_R1138_U386 , P1_U3468 , P1_R1138_U27 );
nand NAND2_13324 ( P1_R1138_U387 , P1_U3058 , P1_R1138_U25 );
nand NAND2_13325 ( P1_R1138_U388 , P1_U3465 , P1_R1138_U26 );
nand NAND2_13326 ( P1_R1138_U389 , P1_R1138_U388 , P1_R1138_U387 );
nand NAND2_13327 ( P1_R1138_U390 , P1_R1138_U352 , P1_R1138_U45 );
nand NAND2_13328 ( P1_R1138_U391 , P1_R1138_U389 , P1_R1138_U218 );
nand NAND2_13329 ( P1_R1138_U392 , P1_U3062 , P1_R1138_U33 );
nand NAND2_13330 ( P1_R1138_U393 , P1_U3462 , P1_R1138_U34 );
nand NAND2_13331 ( P1_R1138_U394 , P1_R1138_U393 , P1_R1138_U392 );
nand NAND2_13332 ( P1_R1138_U395 , P1_R1138_U353 , P1_R1138_U141 );
nand NAND2_13333 ( P1_R1138_U396 , P1_R1138_U227 , P1_R1138_U394 );
nand NAND2_13334 ( P1_R1138_U397 , P1_U3066 , P1_R1138_U28 );
nand NAND2_13335 ( P1_R1138_U398 , P1_U3459 , P1_R1138_U29 );
nand NAND2_13336 ( P1_R1138_U399 , P1_U3053 , P1_R1138_U143 );
nand NAND2_13337 ( P1_R1138_U400 , P1_U4018 , P1_R1138_U142 );
nand NAND2_13338 ( P1_R1138_U401 , P1_U3053 , P1_R1138_U143 );
nand NAND2_13339 ( P1_R1138_U402 , P1_U4018 , P1_R1138_U142 );
nand NAND2_13340 ( P1_R1138_U403 , P1_R1138_U402 , P1_R1138_U401 );
nand NAND2_13341 ( P1_R1138_U404 , P1_R1138_U144 , P1_R1138_U145 );
nand NAND2_13342 ( P1_R1138_U405 , P1_R1138_U302 , P1_R1138_U403 );
nand NAND2_13343 ( P1_R1138_U406 , P1_U3052 , P1_R1138_U89 );
nand NAND2_13344 ( P1_R1138_U407 , P1_U4007 , P1_R1138_U88 );
nand NAND2_13345 ( P1_R1138_U408 , P1_U3052 , P1_R1138_U89 );
nand NAND2_13346 ( P1_R1138_U409 , P1_U4007 , P1_R1138_U88 );
nand NAND2_13347 ( P1_R1138_U410 , P1_R1138_U409 , P1_R1138_U408 );
nand NAND2_13348 ( P1_R1138_U411 , P1_R1138_U146 , P1_R1138_U147 );
nand NAND2_13349 ( P1_R1138_U412 , P1_R1138_U300 , P1_R1138_U410 );
nand NAND2_13350 ( P1_R1138_U413 , P1_U3051 , P1_R1138_U47 );
nand NAND2_13351 ( P1_R1138_U414 , P1_U4008 , P1_R1138_U48 );
nand NAND2_13352 ( P1_R1138_U415 , P1_U3051 , P1_R1138_U47 );
nand NAND2_13353 ( P1_R1138_U416 , P1_U4008 , P1_R1138_U48 );
nand NAND2_13354 ( P1_R1138_U417 , P1_R1138_U416 , P1_R1138_U415 );
nand NAND2_13355 ( P1_R1138_U418 , P1_R1138_U148 , P1_R1138_U149 );
nand NAND2_13356 ( P1_R1138_U419 , P1_R1138_U297 , P1_R1138_U417 );
nand NAND2_13357 ( P1_R1138_U420 , P1_U3055 , P1_R1138_U50 );
nand NAND2_13358 ( P1_R1138_U421 , P1_U4009 , P1_R1138_U49 );
nand NAND2_13359 ( P1_R1138_U422 , P1_U3056 , P1_R1138_U51 );
nand NAND2_13360 ( P1_R1138_U423 , P1_U4010 , P1_R1138_U52 );
nand NAND2_13361 ( P1_R1138_U424 , P1_R1138_U423 , P1_R1138_U422 );
nand NAND2_13362 ( P1_R1138_U425 , P1_R1138_U354 , P1_R1138_U90 );
nand NAND2_13363 ( P1_R1138_U426 , P1_R1138_U424 , P1_R1138_U304 );
nand NAND2_13364 ( P1_R1138_U427 , P1_U3063 , P1_R1138_U53 );
nand NAND2_13365 ( P1_R1138_U428 , P1_U4011 , P1_R1138_U54 );
nand NAND2_13366 ( P1_R1138_U429 , P1_R1138_U428 , P1_R1138_U427 );
nand NAND2_13367 ( P1_R1138_U430 , P1_R1138_U355 , P1_R1138_U151 );
nand NAND2_13368 ( P1_R1138_U431 , P1_R1138_U291 , P1_R1138_U429 );
nand NAND2_13369 ( P1_R1138_U432 , P1_U3064 , P1_R1138_U85 );
nand NAND2_13370 ( P1_R1138_U433 , P1_U4012 , P1_R1138_U86 );
nand NAND2_13371 ( P1_R1138_U434 , P1_U3064 , P1_R1138_U85 );
nand NAND2_13372 ( P1_R1138_U435 , P1_U4012 , P1_R1138_U86 );
nand NAND2_13373 ( P1_R1138_U436 , P1_R1138_U435 , P1_R1138_U434 );
nand NAND2_13374 ( P1_R1138_U437 , P1_R1138_U152 , P1_R1138_U153 );
nand NAND2_13375 ( P1_R1138_U438 , P1_R1138_U287 , P1_R1138_U436 );
nand NAND2_13376 ( P1_R1138_U439 , P1_U3059 , P1_R1138_U83 );
nand NAND2_13377 ( P1_R1138_U440 , P1_U4013 , P1_R1138_U84 );
nand NAND2_13378 ( P1_R1138_U441 , P1_U3059 , P1_R1138_U83 );
nand NAND2_13379 ( P1_R1138_U442 , P1_U4013 , P1_R1138_U84 );
nand NAND2_13380 ( P1_R1138_U443 , P1_R1138_U442 , P1_R1138_U441 );
nand NAND2_13381 ( P1_R1138_U444 , P1_R1138_U154 , P1_R1138_U155 );
nand NAND2_13382 ( P1_R1138_U445 , P1_R1138_U283 , P1_R1138_U443 );
nand NAND2_13383 ( P1_R1138_U446 , P1_U3073 , P1_R1138_U55 );
nand NAND2_13384 ( P1_R1138_U447 , P1_U4014 , P1_R1138_U56 );
nand NAND2_13385 ( P1_R1138_U448 , P1_U3073 , P1_R1138_U55 );
nand NAND2_13386 ( P1_R1138_U449 , P1_U4014 , P1_R1138_U56 );
nand NAND2_13387 ( P1_R1138_U450 , P1_R1138_U449 , P1_R1138_U448 );
nand NAND2_13388 ( P1_R1138_U451 , P1_U3074 , P1_R1138_U82 );
nand NAND2_13389 ( P1_R1138_U452 , P1_U4015 , P1_R1138_U91 );
nand NAND2_13390 ( P1_R1138_U453 , P1_R1138_U179 , P1_R1138_U158 );
nand NAND2_13391 ( P1_R1138_U454 , P1_R1138_U325 , P1_R1138_U32 );
nand NAND2_13392 ( P1_R1138_U455 , P1_U3079 , P1_R1138_U79 );
nand NAND2_13393 ( P1_R1138_U456 , P1_U3509 , P1_R1138_U80 );
nand NAND2_13394 ( P1_R1138_U457 , P1_R1138_U456 , P1_R1138_U455 );
nand NAND2_13395 ( P1_R1138_U458 , P1_R1138_U356 , P1_R1138_U92 );
nand NAND2_13396 ( P1_R1138_U459 , P1_R1138_U457 , P1_R1138_U313 );
nand NAND2_13397 ( P1_R1138_U460 , P1_U3080 , P1_R1138_U76 );
nand NAND2_13398 ( P1_R1138_U461 , P1_U3507 , P1_R1138_U77 );
nand NAND2_13399 ( P1_R1138_U462 , P1_R1138_U461 , P1_R1138_U460 );
nand NAND2_13400 ( P1_R1138_U463 , P1_R1138_U357 , P1_R1138_U159 );
nand NAND2_13401 ( P1_R1138_U464 , P1_R1138_U267 , P1_R1138_U462 );
nand NAND2_13402 ( P1_R1138_U465 , P1_U3067 , P1_R1138_U61 );
nand NAND2_13403 ( P1_R1138_U466 , P1_U3504 , P1_R1138_U59 );
nand NAND2_13404 ( P1_R1138_U467 , P1_U3071 , P1_R1138_U57 );
nand NAND2_13405 ( P1_R1138_U468 , P1_U3501 , P1_R1138_U58 );
nand NAND2_13406 ( P1_R1138_U469 , P1_R1138_U468 , P1_R1138_U467 );
nand NAND2_13407 ( P1_R1138_U470 , P1_R1138_U358 , P1_R1138_U93 );
nand NAND2_13408 ( P1_R1138_U471 , P1_R1138_U469 , P1_R1138_U259 );
nand NAND2_13409 ( P1_R1138_U472 , P1_U3072 , P1_R1138_U74 );
nand NAND2_13410 ( P1_R1138_U473 , P1_U3498 , P1_R1138_U75 );
nand NAND2_13411 ( P1_R1138_U474 , P1_U3072 , P1_R1138_U74 );
nand NAND2_13412 ( P1_R1138_U475 , P1_U3498 , P1_R1138_U75 );
nand NAND2_13413 ( P1_R1138_U476 , P1_R1138_U475 , P1_R1138_U474 );
nand NAND2_13414 ( P1_R1138_U477 , P1_R1138_U160 , P1_R1138_U161 );
nand NAND2_13415 ( P1_R1138_U478 , P1_R1138_U255 , P1_R1138_U476 );
nand NAND2_13416 ( P1_R1138_U479 , P1_U3077 , P1_R1138_U72 );
nand NAND2_13417 ( P1_R1138_U480 , P1_U3495 , P1_R1138_U73 );
nand NAND2_13418 ( P1_R1138_U481 , P1_U3077 , P1_R1138_U72 );
nand NAND2_13419 ( P1_R1138_U482 , P1_U3495 , P1_R1138_U73 );
nand NAND2_13420 ( P1_R1138_U483 , P1_R1138_U482 , P1_R1138_U481 );
nand NAND2_13421 ( P1_R1138_U484 , P1_R1138_U162 , P1_R1138_U163 );
nand NAND2_13422 ( P1_R1138_U485 , P1_R1138_U251 , P1_R1138_U483 );
nand NAND2_13423 ( P1_R1138_U486 , P1_U3078 , P1_R1138_U70 );
nand NAND2_13424 ( P1_R1138_U487 , P1_U3492 , P1_R1138_U71 );
nand NAND2_13425 ( P1_R1138_U488 , P1_U3070 , P1_R1138_U65 );
nand NAND2_13426 ( P1_R1138_U489 , P1_U3489 , P1_R1138_U66 );
nand NAND2_13427 ( P1_R1138_U490 , P1_R1138_U489 , P1_R1138_U488 );
nand NAND2_13428 ( P1_R1138_U491 , P1_R1138_U359 , P1_R1138_U94 );
nand NAND2_13429 ( P1_R1138_U492 , P1_R1138_U490 , P1_R1138_U335 );
nand NAND2_13430 ( P1_R1138_U493 , P1_U3061 , P1_R1138_U67 );
nand NAND2_13431 ( P1_R1138_U494 , P1_U3486 , P1_R1138_U68 );
nand NAND2_13432 ( P1_R1138_U495 , P1_R1138_U494 , P1_R1138_U493 );
nand NAND2_13433 ( P1_R1138_U496 , P1_R1138_U360 , P1_R1138_U164 );
nand NAND2_13434 ( P1_R1138_U497 , P1_R1138_U241 , P1_R1138_U495 );
nand NAND2_13435 ( P1_R1138_U498 , P1_U3060 , P1_R1138_U63 );
nand NAND2_13436 ( P1_R1138_U499 , P1_U3483 , P1_R1138_U64 );
nand NAND2_13437 ( P1_R1138_U500 , P1_U3075 , P1_R1138_U30 );
nand NAND2_13438 ( P1_R1138_U501 , P1_U3451 , P1_R1138_U31 );
and AND2_13439 ( P1_R1222_U4 , P1_R1222_U176 , P1_R1222_U175 );
and AND2_13440 ( P1_R1222_U5 , P1_R1222_U177 , P1_R1222_U178 );
and AND2_13441 ( P1_R1222_U6 , P1_R1222_U194 , P1_R1222_U193 );
and AND2_13442 ( P1_R1222_U7 , P1_R1222_U234 , P1_R1222_U233 );
and AND2_13443 ( P1_R1222_U8 , P1_R1222_U243 , P1_R1222_U242 );
and AND2_13444 ( P1_R1222_U9 , P1_R1222_U261 , P1_R1222_U260 );
and AND2_13445 ( P1_R1222_U10 , P1_R1222_U269 , P1_R1222_U268 );
and AND2_13446 ( P1_R1222_U11 , P1_R1222_U348 , P1_R1222_U345 );
and AND2_13447 ( P1_R1222_U12 , P1_R1222_U341 , P1_R1222_U338 );
and AND2_13448 ( P1_R1222_U13 , P1_R1222_U332 , P1_R1222_U329 );
and AND2_13449 ( P1_R1222_U14 , P1_R1222_U323 , P1_R1222_U320 );
and AND2_13450 ( P1_R1222_U15 , P1_R1222_U317 , P1_R1222_U315 );
and AND2_13451 ( P1_R1222_U16 , P1_R1222_U310 , P1_R1222_U307 );
and AND2_13452 ( P1_R1222_U17 , P1_R1222_U232 , P1_R1222_U229 );
and AND2_13453 ( P1_R1222_U18 , P1_R1222_U224 , P1_R1222_U221 );
and AND2_13454 ( P1_R1222_U19 , P1_R1222_U210 , P1_R1222_U207 );
not NOT1_13455 ( P1_R1222_U20 , P1_U3471 );
not NOT1_13456 ( P1_R1222_U21 , P1_U3069 );
not NOT1_13457 ( P1_R1222_U22 , P1_U3068 );
nand NAND2_13458 ( P1_R1222_U23 , P1_U3069 , P1_U3471 );
not NOT1_13459 ( P1_R1222_U24 , P1_U3474 );
not NOT1_13460 ( P1_R1222_U25 , P1_U3465 );
not NOT1_13461 ( P1_R1222_U26 , P1_U3058 );
not NOT1_13462 ( P1_R1222_U27 , P1_U3065 );
not NOT1_13463 ( P1_R1222_U28 , P1_U3459 );
not NOT1_13464 ( P1_R1222_U29 , P1_U3066 );
not NOT1_13465 ( P1_R1222_U30 , P1_U3451 );
not NOT1_13466 ( P1_R1222_U31 , P1_U3075 );
nand NAND2_13467 ( P1_R1222_U32 , P1_U3075 , P1_U3451 );
not NOT1_13468 ( P1_R1222_U33 , P1_U3462 );
not NOT1_13469 ( P1_R1222_U34 , P1_U3062 );
nand NAND2_13470 ( P1_R1222_U35 , P1_U3058 , P1_U3465 );
not NOT1_13471 ( P1_R1222_U36 , P1_U3468 );
not NOT1_13472 ( P1_R1222_U37 , P1_U3477 );
not NOT1_13473 ( P1_R1222_U38 , P1_U3082 );
not NOT1_13474 ( P1_R1222_U39 , P1_U3081 );
not NOT1_13475 ( P1_R1222_U40 , P1_U3480 );
nand NAND2_13476 ( P1_R1222_U41 , P1_R1222_U62 , P1_R1222_U202 );
nand NAND2_13477 ( P1_R1222_U42 , P1_R1222_U118 , P1_R1222_U190 );
nand NAND2_13478 ( P1_R1222_U43 , P1_R1222_U179 , P1_R1222_U180 );
nand NAND2_13479 ( P1_R1222_U44 , P1_U3456 , P1_U3076 );
nand NAND2_13480 ( P1_R1222_U45 , P1_R1222_U122 , P1_R1222_U216 );
nand NAND2_13481 ( P1_R1222_U46 , P1_R1222_U213 , P1_R1222_U212 );
not NOT1_13482 ( P1_R1222_U47 , P1_U4008 );
not NOT1_13483 ( P1_R1222_U48 , P1_U3051 );
not NOT1_13484 ( P1_R1222_U49 , P1_U3055 );
not NOT1_13485 ( P1_R1222_U50 , P1_U4009 );
not NOT1_13486 ( P1_R1222_U51 , P1_U4010 );
not NOT1_13487 ( P1_R1222_U52 , P1_U3056 );
not NOT1_13488 ( P1_R1222_U53 , P1_U4011 );
not NOT1_13489 ( P1_R1222_U54 , P1_U3063 );
not NOT1_13490 ( P1_R1222_U55 , P1_U4014 );
not NOT1_13491 ( P1_R1222_U56 , P1_U3073 );
not NOT1_13492 ( P1_R1222_U57 , P1_U3501 );
not NOT1_13493 ( P1_R1222_U58 , P1_U3071 );
not NOT1_13494 ( P1_R1222_U59 , P1_U3067 );
nand NAND2_13495 ( P1_R1222_U60 , P1_U3071 , P1_U3501 );
not NOT1_13496 ( P1_R1222_U61 , P1_U3504 );
nand NAND2_13497 ( P1_R1222_U62 , P1_U3082 , P1_U3477 );
not NOT1_13498 ( P1_R1222_U63 , P1_U3483 );
not NOT1_13499 ( P1_R1222_U64 , P1_U3060 );
not NOT1_13500 ( P1_R1222_U65 , P1_U3489 );
not NOT1_13501 ( P1_R1222_U66 , P1_U3070 );
not NOT1_13502 ( P1_R1222_U67 , P1_U3486 );
not NOT1_13503 ( P1_R1222_U68 , P1_U3061 );
nand NAND2_13504 ( P1_R1222_U69 , P1_U3061 , P1_U3486 );
not NOT1_13505 ( P1_R1222_U70 , P1_U3492 );
not NOT1_13506 ( P1_R1222_U71 , P1_U3078 );
not NOT1_13507 ( P1_R1222_U72 , P1_U3495 );
not NOT1_13508 ( P1_R1222_U73 , P1_U3077 );
not NOT1_13509 ( P1_R1222_U74 , P1_U3498 );
not NOT1_13510 ( P1_R1222_U75 , P1_U3072 );
not NOT1_13511 ( P1_R1222_U76 , P1_U3507 );
not NOT1_13512 ( P1_R1222_U77 , P1_U3080 );
nand NAND2_13513 ( P1_R1222_U78 , P1_U3080 , P1_U3507 );
not NOT1_13514 ( P1_R1222_U79 , P1_U3509 );
not NOT1_13515 ( P1_R1222_U80 , P1_U3079 );
nand NAND2_13516 ( P1_R1222_U81 , P1_U3079 , P1_U3509 );
not NOT1_13517 ( P1_R1222_U82 , P1_U4015 );
not NOT1_13518 ( P1_R1222_U83 , P1_U4013 );
not NOT1_13519 ( P1_R1222_U84 , P1_U3059 );
not NOT1_13520 ( P1_R1222_U85 , P1_U4012 );
not NOT1_13521 ( P1_R1222_U86 , P1_U3064 );
nand NAND2_13522 ( P1_R1222_U87 , P1_U4009 , P1_U3055 );
not NOT1_13523 ( P1_R1222_U88 , P1_U3052 );
not NOT1_13524 ( P1_R1222_U89 , P1_U4007 );
nand NAND2_13525 ( P1_R1222_U90 , P1_R1222_U303 , P1_R1222_U173 );
not NOT1_13526 ( P1_R1222_U91 , P1_U3074 );
nand NAND2_13527 ( P1_R1222_U92 , P1_R1222_U78 , P1_R1222_U312 );
nand NAND2_13528 ( P1_R1222_U93 , P1_R1222_U258 , P1_R1222_U257 );
nand NAND2_13529 ( P1_R1222_U94 , P1_R1222_U69 , P1_R1222_U334 );
nand NAND2_13530 ( P1_R1222_U95 , P1_R1222_U454 , P1_R1222_U453 );
nand NAND2_13531 ( P1_R1222_U96 , P1_R1222_U501 , P1_R1222_U500 );
nand NAND2_13532 ( P1_R1222_U97 , P1_R1222_U372 , P1_R1222_U371 );
nand NAND2_13533 ( P1_R1222_U98 , P1_R1222_U377 , P1_R1222_U376 );
nand NAND2_13534 ( P1_R1222_U99 , P1_R1222_U384 , P1_R1222_U383 );
nand NAND2_13535 ( P1_R1222_U100 , P1_R1222_U391 , P1_R1222_U390 );
nand NAND2_13536 ( P1_R1222_U101 , P1_R1222_U396 , P1_R1222_U395 );
nand NAND2_13537 ( P1_R1222_U102 , P1_R1222_U405 , P1_R1222_U404 );
nand NAND2_13538 ( P1_R1222_U103 , P1_R1222_U412 , P1_R1222_U411 );
nand NAND2_13539 ( P1_R1222_U104 , P1_R1222_U419 , P1_R1222_U418 );
nand NAND2_13540 ( P1_R1222_U105 , P1_R1222_U426 , P1_R1222_U425 );
nand NAND2_13541 ( P1_R1222_U106 , P1_R1222_U431 , P1_R1222_U430 );
nand NAND2_13542 ( P1_R1222_U107 , P1_R1222_U438 , P1_R1222_U437 );
nand NAND2_13543 ( P1_R1222_U108 , P1_R1222_U445 , P1_R1222_U444 );
nand NAND2_13544 ( P1_R1222_U109 , P1_R1222_U459 , P1_R1222_U458 );
nand NAND2_13545 ( P1_R1222_U110 , P1_R1222_U464 , P1_R1222_U463 );
nand NAND2_13546 ( P1_R1222_U111 , P1_R1222_U471 , P1_R1222_U470 );
nand NAND2_13547 ( P1_R1222_U112 , P1_R1222_U478 , P1_R1222_U477 );
nand NAND2_13548 ( P1_R1222_U113 , P1_R1222_U485 , P1_R1222_U484 );
nand NAND2_13549 ( P1_R1222_U114 , P1_R1222_U492 , P1_R1222_U491 );
nand NAND2_13550 ( P1_R1222_U115 , P1_R1222_U497 , P1_R1222_U496 );
and AND2_13551 ( P1_R1222_U116 , P1_U3459 , P1_U3066 );
and AND2_13552 ( P1_R1222_U117 , P1_R1222_U186 , P1_R1222_U184 );
and AND2_13553 ( P1_R1222_U118 , P1_R1222_U191 , P1_R1222_U189 );
and AND2_13554 ( P1_R1222_U119 , P1_R1222_U198 , P1_R1222_U197 );
and AND3_13555 ( P1_R1222_U120 , P1_R1222_U379 , P1_R1222_U378 , P1_R1222_U23 );
and AND2_13556 ( P1_R1222_U121 , P1_R1222_U209 , P1_R1222_U6 );
and AND2_13557 ( P1_R1222_U122 , P1_R1222_U217 , P1_R1222_U215 );
and AND3_13558 ( P1_R1222_U123 , P1_R1222_U386 , P1_R1222_U385 , P1_R1222_U35 );
and AND2_13559 ( P1_R1222_U124 , P1_R1222_U223 , P1_R1222_U4 );
and AND2_13560 ( P1_R1222_U125 , P1_R1222_U231 , P1_R1222_U178 );
and AND2_13561 ( P1_R1222_U126 , P1_R1222_U201 , P1_R1222_U7 );
and AND2_13562 ( P1_R1222_U127 , P1_R1222_U236 , P1_R1222_U168 );
and AND2_13563 ( P1_R1222_U128 , P1_R1222_U245 , P1_R1222_U169 );
and AND2_13564 ( P1_R1222_U129 , P1_R1222_U265 , P1_R1222_U264 );
and AND2_13565 ( P1_R1222_U130 , P1_R1222_U10 , P1_R1222_U279 );
and AND2_13566 ( P1_R1222_U131 , P1_R1222_U282 , P1_R1222_U277 );
and AND2_13567 ( P1_R1222_U132 , P1_R1222_U298 , P1_R1222_U295 );
and AND2_13568 ( P1_R1222_U133 , P1_R1222_U365 , P1_R1222_U299 );
and AND2_13569 ( P1_R1222_U134 , P1_R1222_U156 , P1_R1222_U275 );
and AND3_13570 ( P1_R1222_U135 , P1_R1222_U466 , P1_R1222_U465 , P1_R1222_U60 );
and AND3_13571 ( P1_R1222_U136 , P1_R1222_U487 , P1_R1222_U486 , P1_R1222_U169 );
and AND2_13572 ( P1_R1222_U137 , P1_R1222_U340 , P1_R1222_U8 );
and AND3_13573 ( P1_R1222_U138 , P1_R1222_U499 , P1_R1222_U498 , P1_R1222_U168 );
and AND2_13574 ( P1_R1222_U139 , P1_R1222_U347 , P1_R1222_U7 );
nand NAND2_13575 ( P1_R1222_U140 , P1_R1222_U119 , P1_R1222_U199 );
nand NAND2_13576 ( P1_R1222_U141 , P1_R1222_U214 , P1_R1222_U226 );
not NOT1_13577 ( P1_R1222_U142 , P1_U3053 );
not NOT1_13578 ( P1_R1222_U143 , P1_U4018 );
and AND2_13579 ( P1_R1222_U144 , P1_R1222_U400 , P1_R1222_U399 );
nand NAND3_13580 ( P1_R1222_U145 , P1_R1222_U301 , P1_R1222_U166 , P1_R1222_U361 );
and AND2_13581 ( P1_R1222_U146 , P1_R1222_U407 , P1_R1222_U406 );
nand NAND3_13582 ( P1_R1222_U147 , P1_R1222_U367 , P1_R1222_U366 , P1_R1222_U133 );
and AND2_13583 ( P1_R1222_U148 , P1_R1222_U414 , P1_R1222_U413 );
nand NAND3_13584 ( P1_R1222_U149 , P1_R1222_U362 , P1_R1222_U296 , P1_R1222_U87 );
and AND2_13585 ( P1_R1222_U150 , P1_R1222_U421 , P1_R1222_U420 );
nand NAND2_13586 ( P1_R1222_U151 , P1_R1222_U290 , P1_R1222_U289 );
and AND2_13587 ( P1_R1222_U152 , P1_R1222_U433 , P1_R1222_U432 );
nand NAND2_13588 ( P1_R1222_U153 , P1_R1222_U286 , P1_R1222_U285 );
and AND2_13589 ( P1_R1222_U154 , P1_R1222_U440 , P1_R1222_U439 );
nand NAND2_13590 ( P1_R1222_U155 , P1_R1222_U131 , P1_R1222_U281 );
and AND2_13591 ( P1_R1222_U156 , P1_R1222_U447 , P1_R1222_U446 );
and AND2_13592 ( P1_R1222_U157 , P1_R1222_U452 , P1_R1222_U451 );
nand NAND2_13593 ( P1_R1222_U158 , P1_R1222_U44 , P1_R1222_U324 );
nand NAND2_13594 ( P1_R1222_U159 , P1_R1222_U129 , P1_R1222_U266 );
and AND2_13595 ( P1_R1222_U160 , P1_R1222_U473 , P1_R1222_U472 );
nand NAND2_13596 ( P1_R1222_U161 , P1_R1222_U254 , P1_R1222_U253 );
and AND2_13597 ( P1_R1222_U162 , P1_R1222_U480 , P1_R1222_U479 );
nand NAND2_13598 ( P1_R1222_U163 , P1_R1222_U250 , P1_R1222_U249 );
nand NAND2_13599 ( P1_R1222_U164 , P1_R1222_U240 , P1_R1222_U239 );
nand NAND2_13600 ( P1_R1222_U165 , P1_R1222_U364 , P1_R1222_U363 );
nand NAND2_13601 ( P1_R1222_U166 , P1_U3052 , P1_R1222_U147 );
not NOT1_13602 ( P1_R1222_U167 , P1_R1222_U35 );
nand NAND2_13603 ( P1_R1222_U168 , P1_U3480 , P1_U3081 );
nand NAND2_13604 ( P1_R1222_U169 , P1_U3070 , P1_U3489 );
nand NAND2_13605 ( P1_R1222_U170 , P1_U3056 , P1_U4010 );
not NOT1_13606 ( P1_R1222_U171 , P1_R1222_U69 );
not NOT1_13607 ( P1_R1222_U172 , P1_R1222_U78 );
nand NAND2_13608 ( P1_R1222_U173 , P1_U3063 , P1_U4011 );
not NOT1_13609 ( P1_R1222_U174 , P1_R1222_U62 );
or OR2_13610 ( P1_R1222_U175 , P1_U3065 , P1_U3468 );
or OR2_13611 ( P1_R1222_U176 , P1_U3058 , P1_U3465 );
or OR2_13612 ( P1_R1222_U177 , P1_U3462 , P1_U3062 );
or OR2_13613 ( P1_R1222_U178 , P1_U3459 , P1_U3066 );
not NOT1_13614 ( P1_R1222_U179 , P1_R1222_U32 );
or OR2_13615 ( P1_R1222_U180 , P1_U3456 , P1_U3076 );
not NOT1_13616 ( P1_R1222_U181 , P1_R1222_U43 );
not NOT1_13617 ( P1_R1222_U182 , P1_R1222_U44 );
nand NAND2_13618 ( P1_R1222_U183 , P1_R1222_U43 , P1_R1222_U44 );
nand NAND2_13619 ( P1_R1222_U184 , P1_R1222_U116 , P1_R1222_U177 );
nand NAND2_13620 ( P1_R1222_U185 , P1_R1222_U5 , P1_R1222_U183 );
nand NAND2_13621 ( P1_R1222_U186 , P1_U3062 , P1_U3462 );
nand NAND2_13622 ( P1_R1222_U187 , P1_R1222_U117 , P1_R1222_U185 );
nand NAND2_13623 ( P1_R1222_U188 , P1_R1222_U36 , P1_R1222_U35 );
nand NAND2_13624 ( P1_R1222_U189 , P1_U3065 , P1_R1222_U188 );
nand NAND2_13625 ( P1_R1222_U190 , P1_R1222_U4 , P1_R1222_U187 );
nand NAND2_13626 ( P1_R1222_U191 , P1_U3468 , P1_R1222_U167 );
not NOT1_13627 ( P1_R1222_U192 , P1_R1222_U42 );
or OR2_13628 ( P1_R1222_U193 , P1_U3068 , P1_U3474 );
or OR2_13629 ( P1_R1222_U194 , P1_U3069 , P1_U3471 );
not NOT1_13630 ( P1_R1222_U195 , P1_R1222_U23 );
nand NAND2_13631 ( P1_R1222_U196 , P1_R1222_U24 , P1_R1222_U23 );
nand NAND2_13632 ( P1_R1222_U197 , P1_U3068 , P1_R1222_U196 );
nand NAND2_13633 ( P1_R1222_U198 , P1_U3474 , P1_R1222_U195 );
nand NAND2_13634 ( P1_R1222_U199 , P1_R1222_U6 , P1_R1222_U42 );
not NOT1_13635 ( P1_R1222_U200 , P1_R1222_U140 );
or OR2_13636 ( P1_R1222_U201 , P1_U3477 , P1_U3082 );
nand NAND2_13637 ( P1_R1222_U202 , P1_R1222_U201 , P1_R1222_U140 );
not NOT1_13638 ( P1_R1222_U203 , P1_R1222_U41 );
or OR2_13639 ( P1_R1222_U204 , P1_U3081 , P1_U3480 );
or OR2_13640 ( P1_R1222_U205 , P1_U3471 , P1_U3069 );
nand NAND2_13641 ( P1_R1222_U206 , P1_R1222_U205 , P1_R1222_U42 );
nand NAND2_13642 ( P1_R1222_U207 , P1_R1222_U120 , P1_R1222_U206 );
nand NAND2_13643 ( P1_R1222_U208 , P1_R1222_U192 , P1_R1222_U23 );
nand NAND2_13644 ( P1_R1222_U209 , P1_U3474 , P1_U3068 );
nand NAND2_13645 ( P1_R1222_U210 , P1_R1222_U121 , P1_R1222_U208 );
or OR2_13646 ( P1_R1222_U211 , P1_U3069 , P1_U3471 );
nand NAND2_13647 ( P1_R1222_U212 , P1_R1222_U182 , P1_R1222_U178 );
nand NAND2_13648 ( P1_R1222_U213 , P1_U3066 , P1_U3459 );
not NOT1_13649 ( P1_R1222_U214 , P1_R1222_U46 );
nand NAND2_13650 ( P1_R1222_U215 , P1_R1222_U181 , P1_R1222_U5 );
nand NAND2_13651 ( P1_R1222_U216 , P1_R1222_U46 , P1_R1222_U177 );
nand NAND2_13652 ( P1_R1222_U217 , P1_U3062 , P1_U3462 );
not NOT1_13653 ( P1_R1222_U218 , P1_R1222_U45 );
or OR2_13654 ( P1_R1222_U219 , P1_U3465 , P1_U3058 );
nand NAND2_13655 ( P1_R1222_U220 , P1_R1222_U219 , P1_R1222_U45 );
nand NAND2_13656 ( P1_R1222_U221 , P1_R1222_U123 , P1_R1222_U220 );
nand NAND2_13657 ( P1_R1222_U222 , P1_R1222_U218 , P1_R1222_U35 );
nand NAND2_13658 ( P1_R1222_U223 , P1_U3468 , P1_U3065 );
nand NAND2_13659 ( P1_R1222_U224 , P1_R1222_U124 , P1_R1222_U222 );
or OR2_13660 ( P1_R1222_U225 , P1_U3058 , P1_U3465 );
nand NAND2_13661 ( P1_R1222_U226 , P1_R1222_U181 , P1_R1222_U178 );
not NOT1_13662 ( P1_R1222_U227 , P1_R1222_U141 );
nand NAND2_13663 ( P1_R1222_U228 , P1_U3062 , P1_U3462 );
nand NAND4_13664 ( P1_R1222_U229 , P1_R1222_U398 , P1_R1222_U397 , P1_R1222_U44 , P1_R1222_U43 );
nand NAND2_13665 ( P1_R1222_U230 , P1_R1222_U44 , P1_R1222_U43 );
nand NAND2_13666 ( P1_R1222_U231 , P1_U3066 , P1_U3459 );
nand NAND2_13667 ( P1_R1222_U232 , P1_R1222_U125 , P1_R1222_U230 );
or OR2_13668 ( P1_R1222_U233 , P1_U3081 , P1_U3480 );
or OR2_13669 ( P1_R1222_U234 , P1_U3060 , P1_U3483 );
nand NAND2_13670 ( P1_R1222_U235 , P1_R1222_U174 , P1_R1222_U7 );
nand NAND2_13671 ( P1_R1222_U236 , P1_U3060 , P1_U3483 );
nand NAND2_13672 ( P1_R1222_U237 , P1_R1222_U127 , P1_R1222_U235 );
or OR2_13673 ( P1_R1222_U238 , P1_U3483 , P1_U3060 );
nand NAND2_13674 ( P1_R1222_U239 , P1_R1222_U126 , P1_R1222_U140 );
nand NAND2_13675 ( P1_R1222_U240 , P1_R1222_U238 , P1_R1222_U237 );
not NOT1_13676 ( P1_R1222_U241 , P1_R1222_U164 );
or OR2_13677 ( P1_R1222_U242 , P1_U3078 , P1_U3492 );
or OR2_13678 ( P1_R1222_U243 , P1_U3070 , P1_U3489 );
nand NAND2_13679 ( P1_R1222_U244 , P1_R1222_U171 , P1_R1222_U8 );
nand NAND2_13680 ( P1_R1222_U245 , P1_U3078 , P1_U3492 );
nand NAND2_13681 ( P1_R1222_U246 , P1_R1222_U128 , P1_R1222_U244 );
or OR2_13682 ( P1_R1222_U247 , P1_U3486 , P1_U3061 );
or OR2_13683 ( P1_R1222_U248 , P1_U3492 , P1_U3078 );
nand NAND3_13684 ( P1_R1222_U249 , P1_R1222_U247 , P1_R1222_U164 , P1_R1222_U8 );
nand NAND2_13685 ( P1_R1222_U250 , P1_R1222_U248 , P1_R1222_U246 );
not NOT1_13686 ( P1_R1222_U251 , P1_R1222_U163 );
or OR2_13687 ( P1_R1222_U252 , P1_U3495 , P1_U3077 );
nand NAND2_13688 ( P1_R1222_U253 , P1_R1222_U252 , P1_R1222_U163 );
nand NAND2_13689 ( P1_R1222_U254 , P1_U3077 , P1_U3495 );
not NOT1_13690 ( P1_R1222_U255 , P1_R1222_U161 );
or OR2_13691 ( P1_R1222_U256 , P1_U3498 , P1_U3072 );
nand NAND2_13692 ( P1_R1222_U257 , P1_R1222_U256 , P1_R1222_U161 );
nand NAND2_13693 ( P1_R1222_U258 , P1_U3072 , P1_U3498 );
not NOT1_13694 ( P1_R1222_U259 , P1_R1222_U93 );
or OR2_13695 ( P1_R1222_U260 , P1_U3067 , P1_U3504 );
or OR2_13696 ( P1_R1222_U261 , P1_U3071 , P1_U3501 );
not NOT1_13697 ( P1_R1222_U262 , P1_R1222_U60 );
nand NAND2_13698 ( P1_R1222_U263 , P1_R1222_U61 , P1_R1222_U60 );
nand NAND2_13699 ( P1_R1222_U264 , P1_U3067 , P1_R1222_U263 );
nand NAND2_13700 ( P1_R1222_U265 , P1_U3504 , P1_R1222_U262 );
nand NAND2_13701 ( P1_R1222_U266 , P1_R1222_U9 , P1_R1222_U93 );
not NOT1_13702 ( P1_R1222_U267 , P1_R1222_U159 );
or OR2_13703 ( P1_R1222_U268 , P1_U3074 , P1_U4015 );
or OR2_13704 ( P1_R1222_U269 , P1_U3079 , P1_U3509 );
or OR2_13705 ( P1_R1222_U270 , P1_U3073 , P1_U4014 );
not NOT1_13706 ( P1_R1222_U271 , P1_R1222_U81 );
nand NAND2_13707 ( P1_R1222_U272 , P1_U4015 , P1_R1222_U271 );
nand NAND2_13708 ( P1_R1222_U273 , P1_R1222_U272 , P1_R1222_U91 );
nand NAND2_13709 ( P1_R1222_U274 , P1_R1222_U81 , P1_R1222_U82 );
nand NAND2_13710 ( P1_R1222_U275 , P1_R1222_U274 , P1_R1222_U273 );
nand NAND2_13711 ( P1_R1222_U276 , P1_R1222_U172 , P1_R1222_U10 );
nand NAND2_13712 ( P1_R1222_U277 , P1_U3073 , P1_U4014 );
nand NAND2_13713 ( P1_R1222_U278 , P1_R1222_U275 , P1_R1222_U276 );
or OR2_13714 ( P1_R1222_U279 , P1_U3507 , P1_U3080 );
or OR2_13715 ( P1_R1222_U280 , P1_U4014 , P1_U3073 );
nand NAND3_13716 ( P1_R1222_U281 , P1_R1222_U270 , P1_R1222_U159 , P1_R1222_U130 );
nand NAND2_13717 ( P1_R1222_U282 , P1_R1222_U280 , P1_R1222_U278 );
not NOT1_13718 ( P1_R1222_U283 , P1_R1222_U155 );
or OR2_13719 ( P1_R1222_U284 , P1_U4013 , P1_U3059 );
nand NAND2_13720 ( P1_R1222_U285 , P1_R1222_U284 , P1_R1222_U155 );
nand NAND2_13721 ( P1_R1222_U286 , P1_U3059 , P1_U4013 );
not NOT1_13722 ( P1_R1222_U287 , P1_R1222_U153 );
or OR2_13723 ( P1_R1222_U288 , P1_U4012 , P1_U3064 );
nand NAND2_13724 ( P1_R1222_U289 , P1_R1222_U288 , P1_R1222_U153 );
nand NAND2_13725 ( P1_R1222_U290 , P1_U3064 , P1_U4012 );
not NOT1_13726 ( P1_R1222_U291 , P1_R1222_U151 );
or OR2_13727 ( P1_R1222_U292 , P1_U3056 , P1_U4010 );
nand NAND2_13728 ( P1_R1222_U293 , P1_R1222_U173 , P1_R1222_U170 );
not NOT1_13729 ( P1_R1222_U294 , P1_R1222_U87 );
or OR2_13730 ( P1_R1222_U295 , P1_U4011 , P1_U3063 );
nand NAND3_13731 ( P1_R1222_U296 , P1_R1222_U151 , P1_R1222_U295 , P1_R1222_U165 );
not NOT1_13732 ( P1_R1222_U297 , P1_R1222_U149 );
or OR2_13733 ( P1_R1222_U298 , P1_U4008 , P1_U3051 );
nand NAND2_13734 ( P1_R1222_U299 , P1_U3051 , P1_U4008 );
not NOT1_13735 ( P1_R1222_U300 , P1_R1222_U147 );
nand NAND2_13736 ( P1_R1222_U301 , P1_U4007 , P1_R1222_U147 );
not NOT1_13737 ( P1_R1222_U302 , P1_R1222_U145 );
nand NAND2_13738 ( P1_R1222_U303 , P1_R1222_U295 , P1_R1222_U151 );
not NOT1_13739 ( P1_R1222_U304 , P1_R1222_U90 );
or OR2_13740 ( P1_R1222_U305 , P1_U4010 , P1_U3056 );
nand NAND2_13741 ( P1_R1222_U306 , P1_R1222_U305 , P1_R1222_U90 );
nand NAND3_13742 ( P1_R1222_U307 , P1_R1222_U306 , P1_R1222_U170 , P1_R1222_U150 );
nand NAND2_13743 ( P1_R1222_U308 , P1_R1222_U304 , P1_R1222_U170 );
nand NAND2_13744 ( P1_R1222_U309 , P1_U4009 , P1_U3055 );
nand NAND3_13745 ( P1_R1222_U310 , P1_R1222_U308 , P1_R1222_U309 , P1_R1222_U165 );
or OR2_13746 ( P1_R1222_U311 , P1_U3056 , P1_U4010 );
nand NAND2_13747 ( P1_R1222_U312 , P1_R1222_U279 , P1_R1222_U159 );
not NOT1_13748 ( P1_R1222_U313 , P1_R1222_U92 );
nand NAND2_13749 ( P1_R1222_U314 , P1_R1222_U10 , P1_R1222_U92 );
nand NAND2_13750 ( P1_R1222_U315 , P1_R1222_U134 , P1_R1222_U314 );
nand NAND2_13751 ( P1_R1222_U316 , P1_R1222_U314 , P1_R1222_U275 );
nand NAND2_13752 ( P1_R1222_U317 , P1_R1222_U450 , P1_R1222_U316 );
or OR2_13753 ( P1_R1222_U318 , P1_U3509 , P1_U3079 );
nand NAND2_13754 ( P1_R1222_U319 , P1_R1222_U318 , P1_R1222_U92 );
nand NAND3_13755 ( P1_R1222_U320 , P1_R1222_U319 , P1_R1222_U81 , P1_R1222_U157 );
nand NAND2_13756 ( P1_R1222_U321 , P1_R1222_U313 , P1_R1222_U81 );
nand NAND2_13757 ( P1_R1222_U322 , P1_U3074 , P1_U4015 );
nand NAND3_13758 ( P1_R1222_U323 , P1_R1222_U322 , P1_R1222_U321 , P1_R1222_U10 );
or OR2_13759 ( P1_R1222_U324 , P1_U3456 , P1_U3076 );
not NOT1_13760 ( P1_R1222_U325 , P1_R1222_U158 );
or OR2_13761 ( P1_R1222_U326 , P1_U3079 , P1_U3509 );
or OR2_13762 ( P1_R1222_U327 , P1_U3501 , P1_U3071 );
nand NAND2_13763 ( P1_R1222_U328 , P1_R1222_U327 , P1_R1222_U93 );
nand NAND2_13764 ( P1_R1222_U329 , P1_R1222_U135 , P1_R1222_U328 );
nand NAND2_13765 ( P1_R1222_U330 , P1_R1222_U259 , P1_R1222_U60 );
nand NAND2_13766 ( P1_R1222_U331 , P1_U3504 , P1_U3067 );
nand NAND3_13767 ( P1_R1222_U332 , P1_R1222_U331 , P1_R1222_U330 , P1_R1222_U9 );
or OR2_13768 ( P1_R1222_U333 , P1_U3071 , P1_U3501 );
nand NAND2_13769 ( P1_R1222_U334 , P1_R1222_U247 , P1_R1222_U164 );
not NOT1_13770 ( P1_R1222_U335 , P1_R1222_U94 );
or OR2_13771 ( P1_R1222_U336 , P1_U3489 , P1_U3070 );
nand NAND2_13772 ( P1_R1222_U337 , P1_R1222_U336 , P1_R1222_U94 );
nand NAND2_13773 ( P1_R1222_U338 , P1_R1222_U136 , P1_R1222_U337 );
nand NAND2_13774 ( P1_R1222_U339 , P1_R1222_U335 , P1_R1222_U169 );
nand NAND2_13775 ( P1_R1222_U340 , P1_U3078 , P1_U3492 );
nand NAND2_13776 ( P1_R1222_U341 , P1_R1222_U137 , P1_R1222_U339 );
or OR2_13777 ( P1_R1222_U342 , P1_U3070 , P1_U3489 );
or OR2_13778 ( P1_R1222_U343 , P1_U3480 , P1_U3081 );
nand NAND2_13779 ( P1_R1222_U344 , P1_R1222_U343 , P1_R1222_U41 );
nand NAND2_13780 ( P1_R1222_U345 , P1_R1222_U138 , P1_R1222_U344 );
nand NAND2_13781 ( P1_R1222_U346 , P1_R1222_U203 , P1_R1222_U168 );
nand NAND2_13782 ( P1_R1222_U347 , P1_U3060 , P1_U3483 );
nand NAND2_13783 ( P1_R1222_U348 , P1_R1222_U139 , P1_R1222_U346 );
nand NAND2_13784 ( P1_R1222_U349 , P1_R1222_U204 , P1_R1222_U168 );
nand NAND2_13785 ( P1_R1222_U350 , P1_R1222_U201 , P1_R1222_U62 );
nand NAND2_13786 ( P1_R1222_U351 , P1_R1222_U211 , P1_R1222_U23 );
nand NAND2_13787 ( P1_R1222_U352 , P1_R1222_U225 , P1_R1222_U35 );
nand NAND2_13788 ( P1_R1222_U353 , P1_R1222_U228 , P1_R1222_U177 );
nand NAND2_13789 ( P1_R1222_U354 , P1_R1222_U311 , P1_R1222_U170 );
nand NAND2_13790 ( P1_R1222_U355 , P1_R1222_U295 , P1_R1222_U173 );
nand NAND2_13791 ( P1_R1222_U356 , P1_R1222_U326 , P1_R1222_U81 );
nand NAND2_13792 ( P1_R1222_U357 , P1_R1222_U279 , P1_R1222_U78 );
nand NAND2_13793 ( P1_R1222_U358 , P1_R1222_U333 , P1_R1222_U60 );
nand NAND2_13794 ( P1_R1222_U359 , P1_R1222_U342 , P1_R1222_U169 );
nand NAND2_13795 ( P1_R1222_U360 , P1_R1222_U247 , P1_R1222_U69 );
nand NAND2_13796 ( P1_R1222_U361 , P1_U4007 , P1_U3052 );
nand NAND2_13797 ( P1_R1222_U362 , P1_R1222_U293 , P1_R1222_U165 );
nand NAND2_13798 ( P1_R1222_U363 , P1_U3055 , P1_R1222_U292 );
nand NAND2_13799 ( P1_R1222_U364 , P1_U4009 , P1_R1222_U292 );
nand NAND3_13800 ( P1_R1222_U365 , P1_R1222_U293 , P1_R1222_U165 , P1_R1222_U298 );
nand NAND3_13801 ( P1_R1222_U366 , P1_R1222_U151 , P1_R1222_U165 , P1_R1222_U132 );
nand NAND2_13802 ( P1_R1222_U367 , P1_R1222_U294 , P1_R1222_U298 );
nand NAND2_13803 ( P1_R1222_U368 , P1_U3081 , P1_R1222_U40 );
nand NAND2_13804 ( P1_R1222_U369 , P1_U3480 , P1_R1222_U39 );
nand NAND2_13805 ( P1_R1222_U370 , P1_R1222_U369 , P1_R1222_U368 );
nand NAND2_13806 ( P1_R1222_U371 , P1_R1222_U349 , P1_R1222_U41 );
nand NAND2_13807 ( P1_R1222_U372 , P1_R1222_U370 , P1_R1222_U203 );
nand NAND2_13808 ( P1_R1222_U373 , P1_U3082 , P1_R1222_U37 );
nand NAND2_13809 ( P1_R1222_U374 , P1_U3477 , P1_R1222_U38 );
nand NAND2_13810 ( P1_R1222_U375 , P1_R1222_U374 , P1_R1222_U373 );
nand NAND2_13811 ( P1_R1222_U376 , P1_R1222_U350 , P1_R1222_U140 );
nand NAND2_13812 ( P1_R1222_U377 , P1_R1222_U200 , P1_R1222_U375 );
nand NAND2_13813 ( P1_R1222_U378 , P1_U3068 , P1_R1222_U24 );
nand NAND2_13814 ( P1_R1222_U379 , P1_U3474 , P1_R1222_U22 );
nand NAND2_13815 ( P1_R1222_U380 , P1_U3069 , P1_R1222_U20 );
nand NAND2_13816 ( P1_R1222_U381 , P1_U3471 , P1_R1222_U21 );
nand NAND2_13817 ( P1_R1222_U382 , P1_R1222_U381 , P1_R1222_U380 );
nand NAND2_13818 ( P1_R1222_U383 , P1_R1222_U351 , P1_R1222_U42 );
nand NAND2_13819 ( P1_R1222_U384 , P1_R1222_U382 , P1_R1222_U192 );
nand NAND2_13820 ( P1_R1222_U385 , P1_U3065 , P1_R1222_U36 );
nand NAND2_13821 ( P1_R1222_U386 , P1_U3468 , P1_R1222_U27 );
nand NAND2_13822 ( P1_R1222_U387 , P1_U3058 , P1_R1222_U25 );
nand NAND2_13823 ( P1_R1222_U388 , P1_U3465 , P1_R1222_U26 );
nand NAND2_13824 ( P1_R1222_U389 , P1_R1222_U388 , P1_R1222_U387 );
nand NAND2_13825 ( P1_R1222_U390 , P1_R1222_U352 , P1_R1222_U45 );
nand NAND2_13826 ( P1_R1222_U391 , P1_R1222_U389 , P1_R1222_U218 );
nand NAND2_13827 ( P1_R1222_U392 , P1_U3062 , P1_R1222_U33 );
nand NAND2_13828 ( P1_R1222_U393 , P1_U3462 , P1_R1222_U34 );
nand NAND2_13829 ( P1_R1222_U394 , P1_R1222_U393 , P1_R1222_U392 );
nand NAND2_13830 ( P1_R1222_U395 , P1_R1222_U353 , P1_R1222_U141 );
nand NAND2_13831 ( P1_R1222_U396 , P1_R1222_U227 , P1_R1222_U394 );
nand NAND2_13832 ( P1_R1222_U397 , P1_U3066 , P1_R1222_U28 );
nand NAND2_13833 ( P1_R1222_U398 , P1_U3459 , P1_R1222_U29 );
nand NAND2_13834 ( P1_R1222_U399 , P1_U3053 , P1_R1222_U143 );
nand NAND2_13835 ( P1_R1222_U400 , P1_U4018 , P1_R1222_U142 );
nand NAND2_13836 ( P1_R1222_U401 , P1_U3053 , P1_R1222_U143 );
nand NAND2_13837 ( P1_R1222_U402 , P1_U4018 , P1_R1222_U142 );
nand NAND2_13838 ( P1_R1222_U403 , P1_R1222_U402 , P1_R1222_U401 );
nand NAND2_13839 ( P1_R1222_U404 , P1_R1222_U144 , P1_R1222_U145 );
nand NAND2_13840 ( P1_R1222_U405 , P1_R1222_U302 , P1_R1222_U403 );
nand NAND2_13841 ( P1_R1222_U406 , P1_U3052 , P1_R1222_U89 );
nand NAND2_13842 ( P1_R1222_U407 , P1_U4007 , P1_R1222_U88 );
nand NAND2_13843 ( P1_R1222_U408 , P1_U3052 , P1_R1222_U89 );
nand NAND2_13844 ( P1_R1222_U409 , P1_U4007 , P1_R1222_U88 );
nand NAND2_13845 ( P1_R1222_U410 , P1_R1222_U409 , P1_R1222_U408 );
nand NAND2_13846 ( P1_R1222_U411 , P1_R1222_U146 , P1_R1222_U147 );
nand NAND2_13847 ( P1_R1222_U412 , P1_R1222_U300 , P1_R1222_U410 );
nand NAND2_13848 ( P1_R1222_U413 , P1_U3051 , P1_R1222_U47 );
nand NAND2_13849 ( P1_R1222_U414 , P1_U4008 , P1_R1222_U48 );
nand NAND2_13850 ( P1_R1222_U415 , P1_U3051 , P1_R1222_U47 );
nand NAND2_13851 ( P1_R1222_U416 , P1_U4008 , P1_R1222_U48 );
nand NAND2_13852 ( P1_R1222_U417 , P1_R1222_U416 , P1_R1222_U415 );
nand NAND2_13853 ( P1_R1222_U418 , P1_R1222_U148 , P1_R1222_U149 );
nand NAND2_13854 ( P1_R1222_U419 , P1_R1222_U297 , P1_R1222_U417 );
nand NAND2_13855 ( P1_R1222_U420 , P1_U3055 , P1_R1222_U50 );
nand NAND2_13856 ( P1_R1222_U421 , P1_U4009 , P1_R1222_U49 );
nand NAND2_13857 ( P1_R1222_U422 , P1_U3056 , P1_R1222_U51 );
nand NAND2_13858 ( P1_R1222_U423 , P1_U4010 , P1_R1222_U52 );
nand NAND2_13859 ( P1_R1222_U424 , P1_R1222_U423 , P1_R1222_U422 );
nand NAND2_13860 ( P1_R1222_U425 , P1_R1222_U354 , P1_R1222_U90 );
nand NAND2_13861 ( P1_R1222_U426 , P1_R1222_U424 , P1_R1222_U304 );
nand NAND2_13862 ( P1_R1222_U427 , P1_U3063 , P1_R1222_U53 );
nand NAND2_13863 ( P1_R1222_U428 , P1_U4011 , P1_R1222_U54 );
nand NAND2_13864 ( P1_R1222_U429 , P1_R1222_U428 , P1_R1222_U427 );
nand NAND2_13865 ( P1_R1222_U430 , P1_R1222_U355 , P1_R1222_U151 );
nand NAND2_13866 ( P1_R1222_U431 , P1_R1222_U291 , P1_R1222_U429 );
nand NAND2_13867 ( P1_R1222_U432 , P1_U3064 , P1_R1222_U85 );
nand NAND2_13868 ( P1_R1222_U433 , P1_U4012 , P1_R1222_U86 );
nand NAND2_13869 ( P1_R1222_U434 , P1_U3064 , P1_R1222_U85 );
nand NAND2_13870 ( P1_R1222_U435 , P1_U4012 , P1_R1222_U86 );
nand NAND2_13871 ( P1_R1222_U436 , P1_R1222_U435 , P1_R1222_U434 );
nand NAND2_13872 ( P1_R1222_U437 , P1_R1222_U152 , P1_R1222_U153 );
nand NAND2_13873 ( P1_R1222_U438 , P1_R1222_U287 , P1_R1222_U436 );
nand NAND2_13874 ( P1_R1222_U439 , P1_U3059 , P1_R1222_U83 );
nand NAND2_13875 ( P1_R1222_U440 , P1_U4013 , P1_R1222_U84 );
nand NAND2_13876 ( P1_R1222_U441 , P1_U3059 , P1_R1222_U83 );
nand NAND2_13877 ( P1_R1222_U442 , P1_U4013 , P1_R1222_U84 );
nand NAND2_13878 ( P1_R1222_U443 , P1_R1222_U442 , P1_R1222_U441 );
nand NAND2_13879 ( P1_R1222_U444 , P1_R1222_U154 , P1_R1222_U155 );
nand NAND2_13880 ( P1_R1222_U445 , P1_R1222_U283 , P1_R1222_U443 );
nand NAND2_13881 ( P1_R1222_U446 , P1_U3073 , P1_R1222_U55 );
nand NAND2_13882 ( P1_R1222_U447 , P1_U4014 , P1_R1222_U56 );
nand NAND2_13883 ( P1_R1222_U448 , P1_U3073 , P1_R1222_U55 );
nand NAND2_13884 ( P1_R1222_U449 , P1_U4014 , P1_R1222_U56 );
nand NAND2_13885 ( P1_R1222_U450 , P1_R1222_U449 , P1_R1222_U448 );
nand NAND2_13886 ( P1_R1222_U451 , P1_U3074 , P1_R1222_U82 );
nand NAND2_13887 ( P1_R1222_U452 , P1_U4015 , P1_R1222_U91 );
nand NAND2_13888 ( P1_R1222_U453 , P1_R1222_U179 , P1_R1222_U158 );
nand NAND2_13889 ( P1_R1222_U454 , P1_R1222_U325 , P1_R1222_U32 );
nand NAND2_13890 ( P1_R1222_U455 , P1_U3079 , P1_R1222_U79 );
nand NAND2_13891 ( P1_R1222_U456 , P1_U3509 , P1_R1222_U80 );
nand NAND2_13892 ( P1_R1222_U457 , P1_R1222_U456 , P1_R1222_U455 );
nand NAND2_13893 ( P1_R1222_U458 , P1_R1222_U356 , P1_R1222_U92 );
nand NAND2_13894 ( P1_R1222_U459 , P1_R1222_U457 , P1_R1222_U313 );
nand NAND2_13895 ( P1_R1222_U460 , P1_U3080 , P1_R1222_U76 );
nand NAND2_13896 ( P1_R1222_U461 , P1_U3507 , P1_R1222_U77 );
nand NAND2_13897 ( P1_R1222_U462 , P1_R1222_U461 , P1_R1222_U460 );
nand NAND2_13898 ( P1_R1222_U463 , P1_R1222_U357 , P1_R1222_U159 );
nand NAND2_13899 ( P1_R1222_U464 , P1_R1222_U267 , P1_R1222_U462 );
nand NAND2_13900 ( P1_R1222_U465 , P1_U3067 , P1_R1222_U61 );
nand NAND2_13901 ( P1_R1222_U466 , P1_U3504 , P1_R1222_U59 );
nand NAND2_13902 ( P1_R1222_U467 , P1_U3071 , P1_R1222_U57 );
nand NAND2_13903 ( P1_R1222_U468 , P1_U3501 , P1_R1222_U58 );
nand NAND2_13904 ( P1_R1222_U469 , P1_R1222_U468 , P1_R1222_U467 );
nand NAND2_13905 ( P1_R1222_U470 , P1_R1222_U358 , P1_R1222_U93 );
nand NAND2_13906 ( P1_R1222_U471 , P1_R1222_U469 , P1_R1222_U259 );
nand NAND2_13907 ( P1_R1222_U472 , P1_U3072 , P1_R1222_U74 );
nand NAND2_13908 ( P1_R1222_U473 , P1_U3498 , P1_R1222_U75 );
nand NAND2_13909 ( P1_R1222_U474 , P1_U3072 , P1_R1222_U74 );
nand NAND2_13910 ( P1_R1222_U475 , P1_U3498 , P1_R1222_U75 );
nand NAND2_13911 ( P1_R1222_U476 , P1_R1222_U475 , P1_R1222_U474 );
nand NAND2_13912 ( P1_R1222_U477 , P1_R1222_U160 , P1_R1222_U161 );
nand NAND2_13913 ( P1_R1222_U478 , P1_R1222_U255 , P1_R1222_U476 );
nand NAND2_13914 ( P1_R1222_U479 , P1_U3077 , P1_R1222_U72 );
nand NAND2_13915 ( P1_R1222_U480 , P1_U3495 , P1_R1222_U73 );
nand NAND2_13916 ( P1_R1222_U481 , P1_U3077 , P1_R1222_U72 );
nand NAND2_13917 ( P1_R1222_U482 , P1_U3495 , P1_R1222_U73 );
nand NAND2_13918 ( P1_R1222_U483 , P1_R1222_U482 , P1_R1222_U481 );
nand NAND2_13919 ( P1_R1222_U484 , P1_R1222_U162 , P1_R1222_U163 );
nand NAND2_13920 ( P1_R1222_U485 , P1_R1222_U251 , P1_R1222_U483 );
nand NAND2_13921 ( P1_R1222_U486 , P1_U3078 , P1_R1222_U70 );
nand NAND2_13922 ( P1_R1222_U487 , P1_U3492 , P1_R1222_U71 );
nand NAND2_13923 ( P1_R1222_U488 , P1_U3070 , P1_R1222_U65 );
nand NAND2_13924 ( P1_R1222_U489 , P1_U3489 , P1_R1222_U66 );
nand NAND2_13925 ( P1_R1222_U490 , P1_R1222_U489 , P1_R1222_U488 );
nand NAND2_13926 ( P1_R1222_U491 , P1_R1222_U359 , P1_R1222_U94 );
nand NAND2_13927 ( P1_R1222_U492 , P1_R1222_U490 , P1_R1222_U335 );
nand NAND2_13928 ( P1_R1222_U493 , P1_U3061 , P1_R1222_U67 );
nand NAND2_13929 ( P1_R1222_U494 , P1_U3486 , P1_R1222_U68 );
nand NAND2_13930 ( P1_R1222_U495 , P1_R1222_U494 , P1_R1222_U493 );
nand NAND2_13931 ( P1_R1222_U496 , P1_R1222_U360 , P1_R1222_U164 );
nand NAND2_13932 ( P1_R1222_U497 , P1_R1222_U241 , P1_R1222_U495 );
nand NAND2_13933 ( P1_R1222_U498 , P1_U3060 , P1_R1222_U63 );
nand NAND2_13934 ( P1_R1222_U499 , P1_U3483 , P1_R1222_U64 );
nand NAND2_13935 ( P1_R1222_U500 , P1_U3075 , P1_R1222_U30 );
nand NAND2_13936 ( P1_R1222_U501 , P1_U3451 , P1_R1222_U31 );
not NOT1_13937 ( P2_ADD_609_U4 , P2_REG3_REG_3_ );
and AND2_13938 ( P2_ADD_609_U5 , P2_ADD_609_U76 , P2_ADD_609_U104 );
not NOT1_13939 ( P2_ADD_609_U6 , P2_REG3_REG_7_ );
not NOT1_13940 ( P2_ADD_609_U7 , P2_REG3_REG_6_ );
not NOT1_13941 ( P2_ADD_609_U8 , P2_REG3_REG_5_ );
not NOT1_13942 ( P2_ADD_609_U9 , P2_REG3_REG_4_ );
nand NAND5_13943 ( P2_ADD_609_U10 , P2_REG3_REG_7_ , P2_REG3_REG_3_ , P2_REG3_REG_6_ , P2_REG3_REG_4_ , P2_REG3_REG_5_ );
not NOT1_13944 ( P2_ADD_609_U11 , P2_REG3_REG_8_ );
not NOT1_13945 ( P2_ADD_609_U12 , P2_REG3_REG_9_ );
nand NAND2_13946 ( P2_ADD_609_U13 , P2_ADD_609_U74 , P2_ADD_609_U85 );
not NOT1_13947 ( P2_ADD_609_U14 , P2_REG3_REG_11_ );
not NOT1_13948 ( P2_ADD_609_U15 , P2_REG3_REG_10_ );
nand NAND2_13949 ( P2_ADD_609_U16 , P2_ADD_609_U75 , P2_ADD_609_U87 );
not NOT1_13950 ( P2_ADD_609_U17 , P2_REG3_REG_12_ );
nand NAND2_13951 ( P2_ADD_609_U18 , P2_REG3_REG_12_ , P2_ADD_609_U89 );
not NOT1_13952 ( P2_ADD_609_U19 , P2_REG3_REG_13_ );
nand NAND2_13953 ( P2_ADD_609_U20 , P2_REG3_REG_13_ , P2_ADD_609_U90 );
not NOT1_13954 ( P2_ADD_609_U21 , P2_REG3_REG_14_ );
nand NAND2_13955 ( P2_ADD_609_U22 , P2_REG3_REG_14_ , P2_ADD_609_U91 );
not NOT1_13956 ( P2_ADD_609_U23 , P2_REG3_REG_15_ );
nand NAND2_13957 ( P2_ADD_609_U24 , P2_REG3_REG_15_ , P2_ADD_609_U92 );
not NOT1_13958 ( P2_ADD_609_U25 , P2_REG3_REG_16_ );
nand NAND2_13959 ( P2_ADD_609_U26 , P2_REG3_REG_16_ , P2_ADD_609_U93 );
not NOT1_13960 ( P2_ADD_609_U27 , P2_REG3_REG_17_ );
nand NAND2_13961 ( P2_ADD_609_U28 , P2_REG3_REG_17_ , P2_ADD_609_U94 );
not NOT1_13962 ( P2_ADD_609_U29 , P2_REG3_REG_18_ );
nand NAND2_13963 ( P2_ADD_609_U30 , P2_REG3_REG_18_ , P2_ADD_609_U95 );
not NOT1_13964 ( P2_ADD_609_U31 , P2_REG3_REG_19_ );
nand NAND2_13965 ( P2_ADD_609_U32 , P2_REG3_REG_19_ , P2_ADD_609_U96 );
not NOT1_13966 ( P2_ADD_609_U33 , P2_REG3_REG_20_ );
nand NAND2_13967 ( P2_ADD_609_U34 , P2_REG3_REG_20_ , P2_ADD_609_U97 );
not NOT1_13968 ( P2_ADD_609_U35 , P2_REG3_REG_21_ );
nand NAND2_13969 ( P2_ADD_609_U36 , P2_REG3_REG_21_ , P2_ADD_609_U98 );
not NOT1_13970 ( P2_ADD_609_U37 , P2_REG3_REG_22_ );
nand NAND2_13971 ( P2_ADD_609_U38 , P2_REG3_REG_22_ , P2_ADD_609_U99 );
not NOT1_13972 ( P2_ADD_609_U39 , P2_REG3_REG_23_ );
nand NAND2_13973 ( P2_ADD_609_U40 , P2_REG3_REG_23_ , P2_ADD_609_U100 );
not NOT1_13974 ( P2_ADD_609_U41 , P2_REG3_REG_24_ );
nand NAND2_13975 ( P2_ADD_609_U42 , P2_REG3_REG_24_ , P2_ADD_609_U101 );
not NOT1_13976 ( P2_ADD_609_U43 , P2_REG3_REG_25_ );
nand NAND2_13977 ( P2_ADD_609_U44 , P2_REG3_REG_25_ , P2_ADD_609_U102 );
not NOT1_13978 ( P2_ADD_609_U45 , P2_REG3_REG_26_ );
nand NAND2_13979 ( P2_ADD_609_U46 , P2_REG3_REG_26_ , P2_ADD_609_U103 );
not NOT1_13980 ( P2_ADD_609_U47 , P2_REG3_REG_28_ );
not NOT1_13981 ( P2_ADD_609_U48 , P2_REG3_REG_27_ );
nand NAND2_13982 ( P2_ADD_609_U49 , P2_ADD_609_U108 , P2_ADD_609_U107 );
nand NAND2_13983 ( P2_ADD_609_U50 , P2_ADD_609_U110 , P2_ADD_609_U109 );
nand NAND2_13984 ( P2_ADD_609_U51 , P2_ADD_609_U112 , P2_ADD_609_U111 );
nand NAND2_13985 ( P2_ADD_609_U52 , P2_ADD_609_U114 , P2_ADD_609_U113 );
nand NAND2_13986 ( P2_ADD_609_U53 , P2_ADD_609_U116 , P2_ADD_609_U115 );
nand NAND2_13987 ( P2_ADD_609_U54 , P2_ADD_609_U118 , P2_ADD_609_U117 );
nand NAND2_13988 ( P2_ADD_609_U55 , P2_ADD_609_U120 , P2_ADD_609_U119 );
nand NAND2_13989 ( P2_ADD_609_U56 , P2_ADD_609_U122 , P2_ADD_609_U121 );
nand NAND2_13990 ( P2_ADD_609_U57 , P2_ADD_609_U124 , P2_ADD_609_U123 );
nand NAND2_13991 ( P2_ADD_609_U58 , P2_ADD_609_U126 , P2_ADD_609_U125 );
nand NAND2_13992 ( P2_ADD_609_U59 , P2_ADD_609_U128 , P2_ADD_609_U127 );
nand NAND2_13993 ( P2_ADD_609_U60 , P2_ADD_609_U130 , P2_ADD_609_U129 );
nand NAND2_13994 ( P2_ADD_609_U61 , P2_ADD_609_U132 , P2_ADD_609_U131 );
nand NAND2_13995 ( P2_ADD_609_U62 , P2_ADD_609_U134 , P2_ADD_609_U133 );
nand NAND2_13996 ( P2_ADD_609_U63 , P2_ADD_609_U136 , P2_ADD_609_U135 );
nand NAND2_13997 ( P2_ADD_609_U64 , P2_ADD_609_U138 , P2_ADD_609_U137 );
nand NAND2_13998 ( P2_ADD_609_U65 , P2_ADD_609_U140 , P2_ADD_609_U139 );
nand NAND2_13999 ( P2_ADD_609_U66 , P2_ADD_609_U142 , P2_ADD_609_U141 );
nand NAND2_14000 ( P2_ADD_609_U67 , P2_ADD_609_U144 , P2_ADD_609_U143 );
nand NAND2_14001 ( P2_ADD_609_U68 , P2_ADD_609_U146 , P2_ADD_609_U145 );
nand NAND2_14002 ( P2_ADD_609_U69 , P2_ADD_609_U148 , P2_ADD_609_U147 );
nand NAND2_14003 ( P2_ADD_609_U70 , P2_ADD_609_U150 , P2_ADD_609_U149 );
nand NAND2_14004 ( P2_ADD_609_U71 , P2_ADD_609_U152 , P2_ADD_609_U151 );
nand NAND2_14005 ( P2_ADD_609_U72 , P2_ADD_609_U154 , P2_ADD_609_U153 );
nand NAND2_14006 ( P2_ADD_609_U73 , P2_ADD_609_U156 , P2_ADD_609_U155 );
and AND2_14007 ( P2_ADD_609_U74 , P2_REG3_REG_8_ , P2_REG3_REG_9_ );
and AND2_14008 ( P2_ADD_609_U75 , P2_REG3_REG_11_ , P2_REG3_REG_10_ );
and AND2_14009 ( P2_ADD_609_U76 , P2_REG3_REG_28_ , P2_REG3_REG_27_ );
nand NAND2_14010 ( P2_ADD_609_U77 , P2_REG3_REG_8_ , P2_ADD_609_U85 );
nand NAND4_14011 ( P2_ADD_609_U78 , P2_REG3_REG_4_ , P2_REG3_REG_5_ , P2_REG3_REG_6_ , P2_REG3_REG_3_ );
nand NAND3_14012 ( P2_ADD_609_U79 , P2_REG3_REG_5_ , P2_REG3_REG_3_ , P2_REG3_REG_4_ );
nand NAND2_14013 ( P2_ADD_609_U80 , P2_REG3_REG_4_ , P2_REG3_REG_3_ );
nand NAND2_14014 ( P2_ADD_609_U81 , P2_REG3_REG_27_ , P2_ADD_609_U104 );
nand NAND2_14015 ( P2_ADD_609_U82 , P2_REG3_REG_10_ , P2_ADD_609_U87 );
not NOT1_14016 ( P2_ADD_609_U83 , P2_ADD_609_U80 );
not NOT1_14017 ( P2_ADD_609_U84 , P2_ADD_609_U78 );
not NOT1_14018 ( P2_ADD_609_U85 , P2_ADD_609_U10 );
not NOT1_14019 ( P2_ADD_609_U86 , P2_ADD_609_U77 );
not NOT1_14020 ( P2_ADD_609_U87 , P2_ADD_609_U13 );
not NOT1_14021 ( P2_ADD_609_U88 , P2_ADD_609_U82 );
not NOT1_14022 ( P2_ADD_609_U89 , P2_ADD_609_U16 );
not NOT1_14023 ( P2_ADD_609_U90 , P2_ADD_609_U18 );
not NOT1_14024 ( P2_ADD_609_U91 , P2_ADD_609_U20 );
not NOT1_14025 ( P2_ADD_609_U92 , P2_ADD_609_U22 );
not NOT1_14026 ( P2_ADD_609_U93 , P2_ADD_609_U24 );
not NOT1_14027 ( P2_ADD_609_U94 , P2_ADD_609_U26 );
not NOT1_14028 ( P2_ADD_609_U95 , P2_ADD_609_U28 );
not NOT1_14029 ( P2_ADD_609_U96 , P2_ADD_609_U30 );
not NOT1_14030 ( P2_ADD_609_U97 , P2_ADD_609_U32 );
not NOT1_14031 ( P2_ADD_609_U98 , P2_ADD_609_U34 );
not NOT1_14032 ( P2_ADD_609_U99 , P2_ADD_609_U36 );
not NOT1_14033 ( P2_ADD_609_U100 , P2_ADD_609_U38 );
not NOT1_14034 ( P2_ADD_609_U101 , P2_ADD_609_U40 );
not NOT1_14035 ( P2_ADD_609_U102 , P2_ADD_609_U42 );
not NOT1_14036 ( P2_ADD_609_U103 , P2_ADD_609_U44 );
not NOT1_14037 ( P2_ADD_609_U104 , P2_ADD_609_U46 );
not NOT1_14038 ( P2_ADD_609_U105 , P2_ADD_609_U81 );
not NOT1_14039 ( P2_ADD_609_U106 , P2_ADD_609_U79 );
nand NAND2_14040 ( P2_ADD_609_U107 , P2_REG3_REG_9_ , P2_ADD_609_U77 );
nand NAND2_14041 ( P2_ADD_609_U108 , P2_ADD_609_U86 , P2_ADD_609_U12 );
nand NAND2_14042 ( P2_ADD_609_U109 , P2_REG3_REG_8_ , P2_ADD_609_U10 );
nand NAND2_14043 ( P2_ADD_609_U110 , P2_ADD_609_U85 , P2_ADD_609_U11 );
nand NAND2_14044 ( P2_ADD_609_U111 , P2_REG3_REG_7_ , P2_ADD_609_U78 );
nand NAND2_14045 ( P2_ADD_609_U112 , P2_ADD_609_U84 , P2_ADD_609_U6 );
nand NAND2_14046 ( P2_ADD_609_U113 , P2_REG3_REG_6_ , P2_ADD_609_U79 );
nand NAND2_14047 ( P2_ADD_609_U114 , P2_ADD_609_U106 , P2_ADD_609_U7 );
nand NAND2_14048 ( P2_ADD_609_U115 , P2_REG3_REG_5_ , P2_ADD_609_U80 );
nand NAND2_14049 ( P2_ADD_609_U116 , P2_ADD_609_U83 , P2_ADD_609_U8 );
nand NAND2_14050 ( P2_ADD_609_U117 , P2_REG3_REG_4_ , P2_ADD_609_U4 );
nand NAND2_14051 ( P2_ADD_609_U118 , P2_REG3_REG_3_ , P2_ADD_609_U9 );
nand NAND2_14052 ( P2_ADD_609_U119 , P2_REG3_REG_28_ , P2_ADD_609_U81 );
nand NAND2_14053 ( P2_ADD_609_U120 , P2_ADD_609_U105 , P2_ADD_609_U47 );
nand NAND2_14054 ( P2_ADD_609_U121 , P2_REG3_REG_27_ , P2_ADD_609_U46 );
nand NAND2_14055 ( P2_ADD_609_U122 , P2_ADD_609_U104 , P2_ADD_609_U48 );
nand NAND2_14056 ( P2_ADD_609_U123 , P2_REG3_REG_26_ , P2_ADD_609_U44 );
nand NAND2_14057 ( P2_ADD_609_U124 , P2_ADD_609_U103 , P2_ADD_609_U45 );
nand NAND2_14058 ( P2_ADD_609_U125 , P2_REG3_REG_25_ , P2_ADD_609_U42 );
nand NAND2_14059 ( P2_ADD_609_U126 , P2_ADD_609_U102 , P2_ADD_609_U43 );
nand NAND2_14060 ( P2_ADD_609_U127 , P2_REG3_REG_24_ , P2_ADD_609_U40 );
nand NAND2_14061 ( P2_ADD_609_U128 , P2_ADD_609_U101 , P2_ADD_609_U41 );
nand NAND2_14062 ( P2_ADD_609_U129 , P2_REG3_REG_23_ , P2_ADD_609_U38 );
nand NAND2_14063 ( P2_ADD_609_U130 , P2_ADD_609_U100 , P2_ADD_609_U39 );
nand NAND2_14064 ( P2_ADD_609_U131 , P2_REG3_REG_22_ , P2_ADD_609_U36 );
nand NAND2_14065 ( P2_ADD_609_U132 , P2_ADD_609_U99 , P2_ADD_609_U37 );
nand NAND2_14066 ( P2_ADD_609_U133 , P2_REG3_REG_21_ , P2_ADD_609_U34 );
nand NAND2_14067 ( P2_ADD_609_U134 , P2_ADD_609_U98 , P2_ADD_609_U35 );
nand NAND2_14068 ( P2_ADD_609_U135 , P2_REG3_REG_20_ , P2_ADD_609_U32 );
nand NAND2_14069 ( P2_ADD_609_U136 , P2_ADD_609_U97 , P2_ADD_609_U33 );
nand NAND2_14070 ( P2_ADD_609_U137 , P2_REG3_REG_19_ , P2_ADD_609_U30 );
nand NAND2_14071 ( P2_ADD_609_U138 , P2_ADD_609_U96 , P2_ADD_609_U31 );
nand NAND2_14072 ( P2_ADD_609_U139 , P2_REG3_REG_18_ , P2_ADD_609_U28 );
nand NAND2_14073 ( P2_ADD_609_U140 , P2_ADD_609_U95 , P2_ADD_609_U29 );
nand NAND2_14074 ( P2_ADD_609_U141 , P2_REG3_REG_17_ , P2_ADD_609_U26 );
nand NAND2_14075 ( P2_ADD_609_U142 , P2_ADD_609_U94 , P2_ADD_609_U27 );
nand NAND2_14076 ( P2_ADD_609_U143 , P2_REG3_REG_16_ , P2_ADD_609_U24 );
nand NAND2_14077 ( P2_ADD_609_U144 , P2_ADD_609_U93 , P2_ADD_609_U25 );
nand NAND2_14078 ( P2_ADD_609_U145 , P2_REG3_REG_15_ , P2_ADD_609_U22 );
nand NAND2_14079 ( P2_ADD_609_U146 , P2_ADD_609_U92 , P2_ADD_609_U23 );
nand NAND2_14080 ( P2_ADD_609_U147 , P2_REG3_REG_14_ , P2_ADD_609_U20 );
nand NAND2_14081 ( P2_ADD_609_U148 , P2_ADD_609_U91 , P2_ADD_609_U21 );
nand NAND2_14082 ( P2_ADD_609_U149 , P2_REG3_REG_13_ , P2_ADD_609_U18 );
nand NAND2_14083 ( P2_ADD_609_U150 , P2_ADD_609_U90 , P2_ADD_609_U19 );
nand NAND2_14084 ( P2_ADD_609_U151 , P2_REG3_REG_12_ , P2_ADD_609_U16 );
nand NAND2_14085 ( P2_ADD_609_U152 , P2_ADD_609_U89 , P2_ADD_609_U17 );
nand NAND2_14086 ( P2_ADD_609_U153 , P2_REG3_REG_11_ , P2_ADD_609_U82 );
nand NAND2_14087 ( P2_ADD_609_U154 , P2_ADD_609_U88 , P2_ADD_609_U14 );
nand NAND2_14088 ( P2_ADD_609_U155 , P2_REG3_REG_10_ , P2_ADD_609_U13 );
nand NAND2_14089 ( P2_ADD_609_U156 , P2_ADD_609_U87 , P2_ADD_609_U15 );
and AND4_14090 ( P2_R1340_U6 , P2_R1340_U179 , P2_R1340_U176 , P2_R1340_U175 , P2_R1340_U173 );
not NOT1_14091 ( P2_R1340_U7 , P2_U3456 );
not NOT1_14092 ( P2_R1340_U8 , P2_U3459 );
not NOT1_14093 ( P2_R1340_U9 , P2_U3462 );
not NOT1_14094 ( P2_R1340_U10 , P2_U3182 );
not NOT1_14095 ( P2_R1340_U11 , P2_U3181 );
not NOT1_14096 ( P2_R1340_U12 , P2_U3180 );
not NOT1_14097 ( P2_R1340_U13 , P2_U3179 );
not NOT1_14098 ( P2_R1340_U14 , P2_U3178 );
not NOT1_14099 ( P2_R1340_U15 , P2_U3177 );
not NOT1_14100 ( P2_R1340_U16 , P2_U3465 );
not NOT1_14101 ( P2_R1340_U17 , P2_U3468 );
not NOT1_14102 ( P2_R1340_U18 , P2_U3471 );
not NOT1_14103 ( P2_R1340_U19 , P2_U3474 );
not NOT1_14104 ( P2_R1340_U20 , P2_U3477 );
not NOT1_14105 ( P2_R1340_U21 , P2_U3480 );
not NOT1_14106 ( P2_R1340_U22 , P2_U3176 );
not NOT1_14107 ( P2_R1340_U23 , P2_U3175 );
not NOT1_14108 ( P2_R1340_U24 , P2_U3174 );
not NOT1_14109 ( P2_R1340_U25 , P2_U3173 );
not NOT1_14110 ( P2_R1340_U26 , P2_U3172 );
not NOT1_14111 ( P2_R1340_U27 , P2_U3171 );
not NOT1_14112 ( P2_R1340_U28 , P2_U3483 );
not NOT1_14113 ( P2_R1340_U29 , P2_U3486 );
not NOT1_14114 ( P2_R1340_U30 , P2_U3489 );
not NOT1_14115 ( P2_R1340_U31 , P2_U3492 );
not NOT1_14116 ( P2_R1340_U32 , P2_U3495 );
not NOT1_14117 ( P2_R1340_U33 , P2_U3498 );
not NOT1_14118 ( P2_R1340_U34 , P2_U3170 );
not NOT1_14119 ( P2_R1340_U35 , P2_U3169 );
not NOT1_14120 ( P2_R1340_U36 , P2_U3168 );
not NOT1_14121 ( P2_R1340_U37 , P2_U3167 );
not NOT1_14122 ( P2_R1340_U38 , P2_U3501 );
not NOT1_14123 ( P2_R1340_U39 , P2_U3504 );
not NOT1_14124 ( P2_R1340_U40 , P2_U3166 );
not NOT1_14125 ( P2_R1340_U41 , P2_U3165 );
not NOT1_14126 ( P2_R1340_U42 , P2_U3506 );
not NOT1_14127 ( P2_R1340_U43 , P2_U3976 );
not NOT1_14128 ( P2_R1340_U44 , P2_U3164 );
not NOT1_14129 ( P2_R1340_U45 , P2_U3163 );
not NOT1_14130 ( P2_R1340_U46 , P2_U3975 );
not NOT1_14131 ( P2_R1340_U47 , P2_U3974 );
not NOT1_14132 ( P2_R1340_U48 , P2_U3162 );
not NOT1_14133 ( P2_R1340_U49 , P2_U3161 );
not NOT1_14134 ( P2_R1340_U50 , P2_U3973 );
not NOT1_14135 ( P2_R1340_U51 , P2_U3972 );
not NOT1_14136 ( P2_R1340_U52 , P2_U3160 );
not NOT1_14137 ( P2_R1340_U53 , P2_U3159 );
not NOT1_14138 ( P2_R1340_U54 , P2_U3971 );
not NOT1_14139 ( P2_R1340_U55 , P2_U3970 );
not NOT1_14140 ( P2_R1340_U56 , P2_U3158 );
not NOT1_14141 ( P2_R1340_U57 , P2_U3157 );
not NOT1_14142 ( P2_R1340_U58 , P2_U3969 );
not NOT1_14143 ( P2_R1340_U59 , P2_U3968 );
not NOT1_14144 ( P2_R1340_U60 , P2_U3156 );
not NOT1_14145 ( P2_R1340_U61 , P2_U3155 );
not NOT1_14146 ( P2_R1340_U62 , P2_U3979 );
not NOT1_14147 ( P2_R1340_U63 , P2_U3153 );
not NOT1_14148 ( P2_R1340_U64 , P2_U3977 );
and AND3_14149 ( P2_R1340_U65 , P2_R1340_U99 , P2_R1340_U100 , P2_R1340_U98 );
and AND3_14150 ( P2_R1340_U66 , P2_R1340_U105 , P2_R1340_U104 , P2_R1340_U178 );
and AND2_14151 ( P2_R1340_U67 , P2_U3181 , P2_R1340_U8 );
and AND4_14152 ( P2_R1340_U68 , P2_R1340_U106 , P2_R1340_U103 , P2_R1340_U102 , P2_R1340_U69 );
and AND3_14153 ( P2_R1340_U69 , P2_R1340_U111 , P2_R1340_U107 , P2_R1340_U112 );
and AND2_14154 ( P2_R1340_U70 , P2_U3468 , P2_R1340_U14 );
and AND4_14155 ( P2_R1340_U71 , P2_R1340_U113 , P2_R1340_U110 , P2_R1340_U109 , P2_R1340_U72 );
and AND3_14156 ( P2_R1340_U72 , P2_R1340_U118 , P2_R1340_U114 , P2_R1340_U119 );
and AND2_14157 ( P2_R1340_U73 , P2_U3175 , P2_R1340_U20 );
and AND4_14158 ( P2_R1340_U74 , P2_R1340_U120 , P2_R1340_U117 , P2_R1340_U116 , P2_R1340_U75 );
and AND3_14159 ( P2_R1340_U75 , P2_R1340_U125 , P2_R1340_U121 , P2_R1340_U126 );
and AND2_14160 ( P2_R1340_U76 , P2_U3486 , P2_R1340_U26 );
and AND4_14161 ( P2_R1340_U77 , P2_R1340_U127 , P2_R1340_U124 , P2_R1340_U123 , P2_R1340_U78 );
and AND3_14162 ( P2_R1340_U78 , P2_R1340_U132 , P2_R1340_U128 , P2_R1340_U133 );
and AND2_14163 ( P2_R1340_U79 , P2_U3169 , P2_R1340_U32 );
and AND3_14164 ( P2_R1340_U80 , P2_R1340_U81 , P2_R1340_U131 , P2_R1340_U130 );
and AND2_14165 ( P2_R1340_U81 , P2_R1340_U135 , P2_R1340_U134 );
and AND2_14166 ( P2_R1340_U82 , P2_R1340_U137 , P2_R1340_U138 );
and AND2_14167 ( P2_R1340_U83 , P2_R1340_U140 , P2_R1340_U141 );
and AND2_14168 ( P2_R1340_U84 , P2_R1340_U143 , P2_R1340_U144 );
and AND2_14169 ( P2_R1340_U85 , P2_R1340_U146 , P2_R1340_U147 );
and AND2_14170 ( P2_R1340_U86 , P2_R1340_U149 , P2_R1340_U150 );
and AND2_14171 ( P2_R1340_U87 , P2_R1340_U152 , P2_R1340_U153 );
and AND2_14172 ( P2_R1340_U88 , P2_R1340_U155 , P2_R1340_U156 );
and AND2_14173 ( P2_R1340_U89 , P2_R1340_U158 , P2_R1340_U159 );
and AND2_14174 ( P2_R1340_U90 , P2_R1340_U161 , P2_R1340_U162 );
and AND2_14175 ( P2_R1340_U91 , P2_R1340_U164 , P2_R1340_U165 );
and AND2_14176 ( P2_R1340_U92 , P2_R1340_U170 , P2_R1340_U171 );
and AND2_14177 ( P2_R1340_U93 , P2_R1340_U177 , P2_R1340_U174 );
and AND2_14178 ( P2_R1340_U94 , P2_U3154 , P2_R1340_U177 );
not NOT1_14179 ( P2_R1340_U95 , P2_U3978 );
not NOT1_14180 ( P2_R1340_U96 , P2_U3183 );
not NOT1_14181 ( P2_R1340_U97 , P2_U3184 );
nand NAND3_14182 ( P2_R1340_U98 , P2_R1340_U97 , P2_R1340_U96 , P2_U3448 );
nand NAND2_14183 ( P2_R1340_U99 , P2_U3453 , P2_R1340_U96 );
nand NAND2_14184 ( P2_R1340_U100 , P2_U3456 , P2_R1340_U10 );
nand NAND2_14185 ( P2_R1340_U101 , P2_R1340_U66 , P2_R1340_U65 );
nand NAND4_14186 ( P2_R1340_U102 , P2_U3182 , P2_R1340_U105 , P2_R1340_U104 , P2_R1340_U7 );
nand NAND2_14187 ( P2_R1340_U103 , P2_R1340_U67 , P2_R1340_U105 );
nand NAND2_14188 ( P2_R1340_U104 , P2_U3459 , P2_R1340_U11 );
nand NAND2_14189 ( P2_R1340_U105 , P2_U3462 , P2_R1340_U12 );
nand NAND2_14190 ( P2_R1340_U106 , P2_U3180 , P2_R1340_U9 );
nand NAND2_14191 ( P2_R1340_U107 , P2_U3179 , P2_R1340_U16 );
nand NAND2_14192 ( P2_R1340_U108 , P2_R1340_U101 , P2_R1340_U68 );
nand NAND4_14193 ( P2_R1340_U109 , P2_U3465 , P2_R1340_U112 , P2_R1340_U111 , P2_R1340_U13 );
nand NAND2_14194 ( P2_R1340_U110 , P2_R1340_U70 , P2_R1340_U112 );
nand NAND2_14195 ( P2_R1340_U111 , P2_U3178 , P2_R1340_U17 );
nand NAND2_14196 ( P2_R1340_U112 , P2_U3177 , P2_R1340_U18 );
nand NAND2_14197 ( P2_R1340_U113 , P2_U3471 , P2_R1340_U15 );
nand NAND2_14198 ( P2_R1340_U114 , P2_U3474 , P2_R1340_U22 );
nand NAND2_14199 ( P2_R1340_U115 , P2_R1340_U108 , P2_R1340_U71 );
nand NAND4_14200 ( P2_R1340_U116 , P2_U3176 , P2_R1340_U119 , P2_R1340_U118 , P2_R1340_U19 );
nand NAND2_14201 ( P2_R1340_U117 , P2_R1340_U73 , P2_R1340_U119 );
nand NAND2_14202 ( P2_R1340_U118 , P2_U3477 , P2_R1340_U23 );
nand NAND2_14203 ( P2_R1340_U119 , P2_U3480 , P2_R1340_U24 );
nand NAND2_14204 ( P2_R1340_U120 , P2_U3174 , P2_R1340_U21 );
nand NAND2_14205 ( P2_R1340_U121 , P2_U3173 , P2_R1340_U28 );
nand NAND2_14206 ( P2_R1340_U122 , P2_R1340_U115 , P2_R1340_U74 );
nand NAND4_14207 ( P2_R1340_U123 , P2_U3483 , P2_R1340_U126 , P2_R1340_U125 , P2_R1340_U25 );
nand NAND2_14208 ( P2_R1340_U124 , P2_R1340_U76 , P2_R1340_U126 );
nand NAND2_14209 ( P2_R1340_U125 , P2_U3172 , P2_R1340_U29 );
nand NAND2_14210 ( P2_R1340_U126 , P2_U3171 , P2_R1340_U30 );
nand NAND2_14211 ( P2_R1340_U127 , P2_U3489 , P2_R1340_U27 );
nand NAND2_14212 ( P2_R1340_U128 , P2_U3492 , P2_R1340_U34 );
nand NAND2_14213 ( P2_R1340_U129 , P2_R1340_U122 , P2_R1340_U77 );
nand NAND4_14214 ( P2_R1340_U130 , P2_U3170 , P2_R1340_U133 , P2_R1340_U132 , P2_R1340_U31 );
nand NAND2_14215 ( P2_R1340_U131 , P2_R1340_U79 , P2_R1340_U133 );
nand NAND2_14216 ( P2_R1340_U132 , P2_U3495 , P2_R1340_U35 );
nand NAND2_14217 ( P2_R1340_U133 , P2_U3498 , P2_R1340_U36 );
nand NAND2_14218 ( P2_R1340_U134 , P2_U3168 , P2_R1340_U33 );
nand NAND2_14219 ( P2_R1340_U135 , P2_U3167 , P2_R1340_U38 );
nand NAND2_14220 ( P2_R1340_U136 , P2_R1340_U129 , P2_R1340_U80 );
nand NAND2_14221 ( P2_R1340_U137 , P2_U3501 , P2_R1340_U37 );
nand NAND2_14222 ( P2_R1340_U138 , P2_U3504 , P2_R1340_U40 );
nand NAND2_14223 ( P2_R1340_U139 , P2_R1340_U82 , P2_R1340_U136 );
nand NAND2_14224 ( P2_R1340_U140 , P2_U3166 , P2_R1340_U39 );
nand NAND2_14225 ( P2_R1340_U141 , P2_U3165 , P2_R1340_U42 );
nand NAND2_14226 ( P2_R1340_U142 , P2_R1340_U83 , P2_R1340_U139 );
nand NAND2_14227 ( P2_R1340_U143 , P2_U3506 , P2_R1340_U41 );
nand NAND2_14228 ( P2_R1340_U144 , P2_U3976 , P2_R1340_U44 );
nand NAND2_14229 ( P2_R1340_U145 , P2_R1340_U84 , P2_R1340_U142 );
nand NAND2_14230 ( P2_R1340_U146 , P2_U3164 , P2_R1340_U43 );
nand NAND2_14231 ( P2_R1340_U147 , P2_U3163 , P2_R1340_U46 );
nand NAND2_14232 ( P2_R1340_U148 , P2_R1340_U85 , P2_R1340_U145 );
nand NAND2_14233 ( P2_R1340_U149 , P2_U3975 , P2_R1340_U45 );
nand NAND2_14234 ( P2_R1340_U150 , P2_U3974 , P2_R1340_U48 );
nand NAND2_14235 ( P2_R1340_U151 , P2_R1340_U86 , P2_R1340_U148 );
nand NAND2_14236 ( P2_R1340_U152 , P2_U3162 , P2_R1340_U47 );
nand NAND2_14237 ( P2_R1340_U153 , P2_U3161 , P2_R1340_U50 );
nand NAND2_14238 ( P2_R1340_U154 , P2_R1340_U87 , P2_R1340_U151 );
nand NAND2_14239 ( P2_R1340_U155 , P2_U3973 , P2_R1340_U49 );
nand NAND2_14240 ( P2_R1340_U156 , P2_U3972 , P2_R1340_U52 );
nand NAND2_14241 ( P2_R1340_U157 , P2_R1340_U88 , P2_R1340_U154 );
nand NAND2_14242 ( P2_R1340_U158 , P2_U3160 , P2_R1340_U51 );
nand NAND2_14243 ( P2_R1340_U159 , P2_U3159 , P2_R1340_U54 );
nand NAND2_14244 ( P2_R1340_U160 , P2_R1340_U89 , P2_R1340_U157 );
nand NAND2_14245 ( P2_R1340_U161 , P2_U3971 , P2_R1340_U53 );
nand NAND2_14246 ( P2_R1340_U162 , P2_U3970 , P2_R1340_U56 );
nand NAND2_14247 ( P2_R1340_U163 , P2_R1340_U90 , P2_R1340_U160 );
nand NAND2_14248 ( P2_R1340_U164 , P2_U3158 , P2_R1340_U55 );
nand NAND2_14249 ( P2_R1340_U165 , P2_U3157 , P2_R1340_U58 );
nand NAND2_14250 ( P2_R1340_U166 , P2_R1340_U91 , P2_R1340_U163 );
nand NAND2_14251 ( P2_R1340_U167 , P2_U3969 , P2_R1340_U57 );
nand NAND2_14252 ( P2_R1340_U168 , P2_U3968 , P2_R1340_U60 );
nand NAND3_14253 ( P2_R1340_U169 , P2_R1340_U167 , P2_R1340_U166 , P2_R1340_U168 );
nand NAND2_14254 ( P2_R1340_U170 , P2_U3156 , P2_R1340_U59 );
nand NAND2_14255 ( P2_R1340_U171 , P2_U3155 , P2_R1340_U62 );
nand NAND2_14256 ( P2_R1340_U172 , P2_R1340_U92 , P2_R1340_U169 );
nand NAND3_14257 ( P2_R1340_U173 , P2_R1340_U172 , P2_R1340_U95 , P2_R1340_U93 );
nand NAND2_14258 ( P2_R1340_U174 , P2_U3979 , P2_R1340_U61 );
nand NAND2_14259 ( P2_R1340_U175 , P2_U3977 , P2_R1340_U63 );
nand NAND3_14260 ( P2_R1340_U176 , P2_R1340_U177 , P2_U3154 , P2_R1340_U95 );
nand NAND2_14261 ( P2_R1340_U177 , P2_U3153 , P2_R1340_U64 );
nand NAND3_14262 ( P2_R1340_U178 , P2_U3448 , P2_U3453 , P2_R1340_U97 );
nand NAND3_14263 ( P2_R1340_U179 , P2_R1340_U174 , P2_R1340_U172 , P2_R1340_U94 );
and AND2_14264 ( P2_SUB_598_U6 , P2_SUB_598_U57 , P2_SUB_598_U56 );
nor nor_14265 ( P2_SUB_598_U7 , P2_IR_REG_25_ , P2_IR_REG_26_ , P2_IR_REG_27_ );
nor nor_14266 ( P2_SUB_598_U8 , P2_IR_REG_25_ , P2_IR_REG_26_ );
and AND4_14267 ( P2_SUB_598_U9 , P2_SUB_598_U55 , P2_SUB_598_U54 , P2_SUB_598_U53 , P2_SUB_598_U52 );
nor nor_14268 ( P2_SUB_598_U10 , P2_IR_REG_12_ , P2_IR_REG_9_ , P2_IR_REG_10_ , P2_IR_REG_11_ );
and AND2_14269 ( P2_SUB_598_U11 , P2_SUB_598_U142 , P2_SUB_598_U47 );
and AND2_14270 ( P2_SUB_598_U12 , P2_SUB_598_U140 , P2_SUB_598_U111 );
and AND2_14271 ( P2_SUB_598_U13 , P2_SUB_598_U139 , P2_SUB_598_U43 );
and AND2_14272 ( P2_SUB_598_U14 , P2_SUB_598_U138 , P2_SUB_598_U44 );
and AND2_14273 ( P2_SUB_598_U15 , P2_SUB_598_U136 , P2_SUB_598_U114 );
and AND2_14274 ( P2_SUB_598_U16 , P2_SUB_598_U135 , P2_SUB_598_U96 );
and AND2_14275 ( P2_SUB_598_U17 , P2_SUB_598_U134 , P2_SUB_598_U125 );
and AND2_14276 ( P2_SUB_598_U18 , P2_SUB_598_U132 , P2_SUB_598_U126 );
and AND2_14277 ( P2_SUB_598_U19 , P2_SUB_598_U131 , P2_SUB_598_U91 );
and AND2_14278 ( P2_SUB_598_U20 , P2_SUB_598_U64 , P2_SUB_598_U144 );
and AND2_14279 ( P2_SUB_598_U21 , P2_SUB_598_U130 , P2_SUB_598_U89 );
and AND2_14280 ( P2_SUB_598_U22 , P2_SUB_598_U124 , P2_SUB_598_U116 );
and AND2_14281 ( P2_SUB_598_U23 , P2_SUB_598_U123 , P2_SUB_598_U117 );
and AND2_14282 ( P2_SUB_598_U24 , P2_SUB_598_U122 , P2_SUB_598_U34 );
and AND2_14283 ( P2_SUB_598_U25 , P2_SUB_598_U109 , P2_SUB_598_U101 );
and AND2_14284 ( P2_SUB_598_U26 , P2_SUB_598_U108 , P2_SUB_598_U30 );
and AND2_14285 ( P2_SUB_598_U27 , P2_SUB_598_U107 , P2_SUB_598_U32 );
and AND2_14286 ( P2_SUB_598_U28 , P2_SUB_598_U105 , P2_SUB_598_U103 );
and AND2_14287 ( P2_SUB_598_U29 , P2_SUB_598_U104 , P2_SUB_598_U31 );
or OR5_14288 ( P2_SUB_598_U30 , P2_IR_REG_1_ , P2_IR_REG_0_ , P2_IR_REG_2_ , P2_IR_REG_3_ , P2_IR_REG_4_ );
nand NAND2_14289 ( P2_SUB_598_U31 , P2_SUB_598_U50 , P2_SUB_598_U148 );
nand NAND2_14290 ( P2_SUB_598_U32 , P2_SUB_598_U51 , P2_SUB_598_U148 );
not NOT1_14291 ( P2_SUB_598_U33 , P2_IR_REG_7_ );
or OR3_14292 ( P2_SUB_598_U34 , P2_IR_REG_1_ , P2_IR_REG_0_ , P2_IR_REG_2_ );
not NOT1_14293 ( P2_SUB_598_U35 , P2_IR_REG_3_ );
nand NAND2_14294 ( P2_SUB_598_U36 , P2_SUB_598_U6 , P2_SUB_598_U9 );
nand NAND2_14295 ( P2_SUB_598_U37 , P2_SUB_598_U58 , P2_SUB_598_U147 );
nand NAND2_14296 ( P2_SUB_598_U38 , P2_SUB_598_U118 , P2_SUB_598_U80 );
not NOT1_14297 ( P2_SUB_598_U39 , P2_IR_REG_25_ );
nand NAND2_14298 ( P2_SUB_598_U40 , P2_SUB_598_U62 , P2_SUB_598_U9 );
not NOT1_14299 ( P2_SUB_598_U41 , P2_IR_REG_23_ );
not NOT1_14300 ( P2_SUB_598_U42 , P2_IR_REG_21_ );
nand NAND2_14301 ( P2_SUB_598_U43 , P2_SUB_598_U10 , P2_SUB_598_U149 );
nand NAND2_14302 ( P2_SUB_598_U44 , P2_SUB_598_U69 , P2_SUB_598_U112 );
not NOT1_14303 ( P2_SUB_598_U45 , P2_IR_REG_16_ );
not NOT1_14304 ( P2_SUB_598_U46 , P2_IR_REG_15_ );
nand NAND2_14305 ( P2_SUB_598_U47 , P2_SUB_598_U70 , P2_SUB_598_U149 );
not NOT1_14306 ( P2_SUB_598_U48 , P2_IR_REG_11_ );
nand NAND2_14307 ( P2_SUB_598_U49 , P2_SUB_598_U169 , P2_SUB_598_U168 );
nor nor_14308 ( P2_SUB_598_U50 , P2_IR_REG_5_ , P2_IR_REG_6_ , P2_IR_REG_7_ , P2_IR_REG_8_ );
nor nor_14309 ( P2_SUB_598_U51 , P2_IR_REG_5_ , P2_IR_REG_6_ );
nor nor_14310 ( P2_SUB_598_U52 , P2_IR_REG_13_ , P2_IR_REG_14_ , P2_IR_REG_12_ , P2_IR_REG_10_ , P2_IR_REG_11_ );
nor nor_14311 ( P2_SUB_598_U53 , P2_IR_REG_15_ , P2_IR_REG_16_ , P2_IR_REG_1_ , P2_IR_REG_0_ );
nor nor_14312 ( P2_SUB_598_U54 , P2_IR_REG_2_ , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ );
nor nor_14313 ( P2_SUB_598_U55 , P2_IR_REG_6_ , P2_IR_REG_7_ , P2_IR_REG_8_ , P2_IR_REG_9_ );
nor nor_14314 ( P2_SUB_598_U56 , P2_IR_REG_17_ , P2_IR_REG_18_ , P2_IR_REG_19_ , P2_IR_REG_20_ );
nor nor_14315 ( P2_SUB_598_U57 , P2_IR_REG_21_ , P2_IR_REG_22_ , P2_IR_REG_23_ , P2_IR_REG_24_ );
and AND2_14316 ( P2_SUB_598_U58 , P2_SUB_598_U7 , P2_SUB_598_U82 );
nor nor_14317 ( P2_SUB_598_U59 , P2_IR_REG_17_ , P2_IR_REG_18_ );
nor nor_14318 ( P2_SUB_598_U60 , P2_IR_REG_19_ , P2_IR_REG_20_ );
nor nor_14319 ( P2_SUB_598_U61 , P2_IR_REG_21_ , P2_IR_REG_22_ );
and AND3_14320 ( P2_SUB_598_U62 , P2_SUB_598_U60 , P2_SUB_598_U59 , P2_SUB_598_U61 );
nor nor_14321 ( P2_SUB_598_U63 , P2_IR_REG_17_ , P2_IR_REG_18_ , P2_IR_REG_19_ , P2_IR_REG_20_ );
and AND2_14322 ( P2_SUB_598_U64 , P2_SUB_598_U143 , P2_SUB_598_U40 );
nor nor_14323 ( P2_SUB_598_U65 , P2_IR_REG_19_ , P2_IR_REG_17_ , P2_IR_REG_18_ );
nor nor_14324 ( P2_SUB_598_U66 , P2_IR_REG_17_ , P2_IR_REG_18_ );
nor nor_14325 ( P2_SUB_598_U67 , P2_IR_REG_15_ , P2_IR_REG_13_ , P2_IR_REG_14_ );
and AND3_14326 ( P2_SUB_598_U68 , P2_SUB_598_U10 , P2_SUB_598_U45 , P2_SUB_598_U67 );
nor nor_14327 ( P2_SUB_598_U69 , P2_IR_REG_13_ , P2_IR_REG_14_ );
nor nor_14328 ( P2_SUB_598_U70 , P2_IR_REG_10_ , P2_IR_REG_9_ );
not NOT1_14329 ( P2_SUB_598_U71 , P2_IR_REG_9_ );
and AND2_14330 ( P2_SUB_598_U72 , P2_SUB_598_U151 , P2_SUB_598_U150 );
not NOT1_14331 ( P2_SUB_598_U73 , P2_IR_REG_5_ );
and AND2_14332 ( P2_SUB_598_U74 , P2_SUB_598_U153 , P2_SUB_598_U152 );
not NOT1_14333 ( P2_SUB_598_U75 , P2_IR_REG_31_ );
nand NAND2_14334 ( P2_SUB_598_U76 , P2_SUB_598_U119 , P2_SUB_598_U78 );
and AND2_14335 ( P2_SUB_598_U77 , P2_SUB_598_U155 , P2_SUB_598_U154 );
not NOT1_14336 ( P2_SUB_598_U78 , P2_IR_REG_30_ );
and AND2_14337 ( P2_SUB_598_U79 , P2_SUB_598_U157 , P2_SUB_598_U156 );
not NOT1_14338 ( P2_SUB_598_U80 , P2_IR_REG_29_ );
and AND2_14339 ( P2_SUB_598_U81 , P2_SUB_598_U159 , P2_SUB_598_U158 );
not NOT1_14340 ( P2_SUB_598_U82 , P2_IR_REG_28_ );
nand NAND3_14341 ( P2_SUB_598_U83 , P2_SUB_598_U6 , P2_SUB_598_U7 , P2_SUB_598_U9 );
and AND2_14342 ( P2_SUB_598_U84 , P2_SUB_598_U161 , P2_SUB_598_U160 );
not NOT1_14343 ( P2_SUB_598_U85 , P2_IR_REG_27_ );
nand NAND3_14344 ( P2_SUB_598_U86 , P2_SUB_598_U6 , P2_SUB_598_U8 , P2_SUB_598_U9 );
and AND2_14345 ( P2_SUB_598_U87 , P2_SUB_598_U163 , P2_SUB_598_U162 );
not NOT1_14346 ( P2_SUB_598_U88 , P2_IR_REG_24_ );
nand NAND2_14347 ( P2_SUB_598_U89 , P2_SUB_598_U128 , P2_SUB_598_U41 );
and AND2_14348 ( P2_SUB_598_U90 , P2_SUB_598_U165 , P2_SUB_598_U164 );
nand NAND2_14349 ( P2_SUB_598_U91 , P2_SUB_598_U63 , P2_SUB_598_U9 );
and AND2_14350 ( P2_SUB_598_U92 , P2_SUB_598_U167 , P2_SUB_598_U166 );
not NOT1_14351 ( P2_SUB_598_U93 , P2_IR_REG_1_ );
not NOT1_14352 ( P2_SUB_598_U94 , P2_IR_REG_0_ );
not NOT1_14353 ( P2_SUB_598_U95 , P2_IR_REG_17_ );
nand NAND2_14354 ( P2_SUB_598_U96 , P2_SUB_598_U68 , P2_SUB_598_U149 );
and AND2_14355 ( P2_SUB_598_U97 , P2_SUB_598_U171 , P2_SUB_598_U170 );
not NOT1_14356 ( P2_SUB_598_U98 , P2_IR_REG_13_ );
and AND2_14357 ( P2_SUB_598_U99 , P2_SUB_598_U173 , P2_SUB_598_U172 );
not NOT1_14358 ( P2_SUB_598_U100 , P2_SUB_598_U34 );
nand NAND2_14359 ( P2_SUB_598_U101 , P2_SUB_598_U100 , P2_SUB_598_U35 );
not NOT1_14360 ( P2_SUB_598_U102 , P2_SUB_598_U32 );
nand NAND2_14361 ( P2_SUB_598_U103 , P2_SUB_598_U102 , P2_SUB_598_U33 );
nand NAND2_14362 ( P2_SUB_598_U104 , P2_IR_REG_8_ , P2_SUB_598_U103 );
nand NAND2_14363 ( P2_SUB_598_U105 , P2_IR_REG_7_ , P2_SUB_598_U32 );
nand NAND2_14364 ( P2_SUB_598_U106 , P2_SUB_598_U148 , P2_SUB_598_U73 );
nand NAND2_14365 ( P2_SUB_598_U107 , P2_IR_REG_6_ , P2_SUB_598_U106 );
nand NAND2_14366 ( P2_SUB_598_U108 , P2_IR_REG_4_ , P2_SUB_598_U101 );
nand NAND2_14367 ( P2_SUB_598_U109 , P2_IR_REG_3_ , P2_SUB_598_U34 );
not NOT1_14368 ( P2_SUB_598_U110 , P2_SUB_598_U47 );
nand NAND2_14369 ( P2_SUB_598_U111 , P2_SUB_598_U110 , P2_SUB_598_U48 );
not NOT1_14370 ( P2_SUB_598_U112 , P2_SUB_598_U43 );
not NOT1_14371 ( P2_SUB_598_U113 , P2_SUB_598_U44 );
nand NAND2_14372 ( P2_SUB_598_U114 , P2_SUB_598_U113 , P2_SUB_598_U46 );
not NOT1_14373 ( P2_SUB_598_U115 , P2_SUB_598_U96 );
nand NAND2_14374 ( P2_SUB_598_U116 , P2_SUB_598_U147 , P2_SUB_598_U39 );
nand NAND2_14375 ( P2_SUB_598_U117 , P2_SUB_598_U8 , P2_SUB_598_U147 );
not NOT1_14376 ( P2_SUB_598_U118 , P2_SUB_598_U37 );
not NOT1_14377 ( P2_SUB_598_U119 , P2_SUB_598_U38 );
not NOT1_14378 ( P2_SUB_598_U120 , P2_SUB_598_U76 );
or OR2_14379 ( P2_SUB_598_U121 , P2_IR_REG_1_ , P2_IR_REG_0_ );
nand NAND2_14380 ( P2_SUB_598_U122 , P2_IR_REG_2_ , P2_SUB_598_U121 );
nand NAND2_14381 ( P2_SUB_598_U123 , P2_IR_REG_26_ , P2_SUB_598_U116 );
nand NAND2_14382 ( P2_SUB_598_U124 , P2_IR_REG_25_ , P2_SUB_598_U36 );
nand NAND2_14383 ( P2_SUB_598_U125 , P2_SUB_598_U66 , P2_SUB_598_U9 );
nand NAND2_14384 ( P2_SUB_598_U126 , P2_SUB_598_U65 , P2_SUB_598_U9 );
not NOT1_14385 ( P2_SUB_598_U127 , P2_SUB_598_U91 );
not NOT1_14386 ( P2_SUB_598_U128 , P2_SUB_598_U40 );
not NOT1_14387 ( P2_SUB_598_U129 , P2_SUB_598_U89 );
nand NAND2_14388 ( P2_SUB_598_U130 , P2_IR_REG_23_ , P2_SUB_598_U40 );
nand NAND2_14389 ( P2_SUB_598_U131 , P2_IR_REG_20_ , P2_SUB_598_U126 );
nand NAND2_14390 ( P2_SUB_598_U132 , P2_IR_REG_19_ , P2_SUB_598_U125 );
nand NAND2_14391 ( P2_SUB_598_U133 , P2_SUB_598_U9 , P2_SUB_598_U95 );
nand NAND2_14392 ( P2_SUB_598_U134 , P2_IR_REG_18_ , P2_SUB_598_U133 );
nand NAND2_14393 ( P2_SUB_598_U135 , P2_IR_REG_16_ , P2_SUB_598_U114 );
nand NAND2_14394 ( P2_SUB_598_U136 , P2_IR_REG_15_ , P2_SUB_598_U44 );
nand NAND2_14395 ( P2_SUB_598_U137 , P2_SUB_598_U112 , P2_SUB_598_U98 );
nand NAND2_14396 ( P2_SUB_598_U138 , P2_IR_REG_14_ , P2_SUB_598_U137 );
nand NAND2_14397 ( P2_SUB_598_U139 , P2_IR_REG_12_ , P2_SUB_598_U111 );
nand NAND2_14398 ( P2_SUB_598_U140 , P2_IR_REG_11_ , P2_SUB_598_U47 );
nand NAND2_14399 ( P2_SUB_598_U141 , P2_SUB_598_U149 , P2_SUB_598_U71 );
nand NAND2_14400 ( P2_SUB_598_U142 , P2_IR_REG_10_ , P2_SUB_598_U141 );
nand NAND2_14401 ( P2_SUB_598_U143 , P2_IR_REG_21_ , P2_IR_REG_22_ );
nand NAND2_14402 ( P2_SUB_598_U144 , P2_IR_REG_22_ , P2_SUB_598_U91 );
not NOT1_14403 ( P2_SUB_598_U145 , P2_SUB_598_U86 );
not NOT1_14404 ( P2_SUB_598_U146 , P2_SUB_598_U83 );
not NOT1_14405 ( P2_SUB_598_U147 , P2_SUB_598_U36 );
not NOT1_14406 ( P2_SUB_598_U148 , P2_SUB_598_U30 );
not NOT1_14407 ( P2_SUB_598_U149 , P2_SUB_598_U31 );
nand NAND2_14408 ( P2_SUB_598_U150 , P2_IR_REG_9_ , P2_SUB_598_U31 );
nand NAND2_14409 ( P2_SUB_598_U151 , P2_SUB_598_U149 , P2_SUB_598_U71 );
nand NAND2_14410 ( P2_SUB_598_U152 , P2_IR_REG_5_ , P2_SUB_598_U30 );
nand NAND2_14411 ( P2_SUB_598_U153 , P2_SUB_598_U148 , P2_SUB_598_U73 );
nand NAND2_14412 ( P2_SUB_598_U154 , P2_IR_REG_31_ , P2_SUB_598_U76 );
nand NAND2_14413 ( P2_SUB_598_U155 , P2_SUB_598_U120 , P2_SUB_598_U75 );
nand NAND2_14414 ( P2_SUB_598_U156 , P2_IR_REG_30_ , P2_SUB_598_U38 );
nand NAND2_14415 ( P2_SUB_598_U157 , P2_SUB_598_U119 , P2_SUB_598_U78 );
nand NAND2_14416 ( P2_SUB_598_U158 , P2_IR_REG_29_ , P2_SUB_598_U37 );
nand NAND2_14417 ( P2_SUB_598_U159 , P2_SUB_598_U118 , P2_SUB_598_U80 );
nand NAND2_14418 ( P2_SUB_598_U160 , P2_IR_REG_28_ , P2_SUB_598_U83 );
nand NAND2_14419 ( P2_SUB_598_U161 , P2_SUB_598_U146 , P2_SUB_598_U82 );
nand NAND2_14420 ( P2_SUB_598_U162 , P2_IR_REG_27_ , P2_SUB_598_U86 );
nand NAND2_14421 ( P2_SUB_598_U163 , P2_SUB_598_U145 , P2_SUB_598_U85 );
nand NAND2_14422 ( P2_SUB_598_U164 , P2_IR_REG_24_ , P2_SUB_598_U89 );
nand NAND2_14423 ( P2_SUB_598_U165 , P2_SUB_598_U129 , P2_SUB_598_U88 );
nand NAND2_14424 ( P2_SUB_598_U166 , P2_IR_REG_21_ , P2_SUB_598_U91 );
nand NAND2_14425 ( P2_SUB_598_U167 , P2_SUB_598_U127 , P2_SUB_598_U42 );
nand NAND2_14426 ( P2_SUB_598_U168 , P2_IR_REG_1_ , P2_SUB_598_U94 );
nand NAND2_14427 ( P2_SUB_598_U169 , P2_IR_REG_0_ , P2_SUB_598_U93 );
nand NAND2_14428 ( P2_SUB_598_U170 , P2_IR_REG_17_ , P2_SUB_598_U96 );
nand NAND2_14429 ( P2_SUB_598_U171 , P2_SUB_598_U115 , P2_SUB_598_U95 );
nand NAND2_14430 ( P2_SUB_598_U172 , P2_IR_REG_13_ , P2_SUB_598_U43 );
nand NAND2_14431 ( P2_SUB_598_U173 , P2_SUB_598_U112 , P2_SUB_598_U98 );
and AND2_14432 ( P2_R1299_U6 , P2_U3059 , P2_R1299_U7 );
not NOT1_14433 ( P2_R1299_U7 , P2_U3056 );
and AND2_14434 ( P2_R1312_U6 , P2_R1312_U129 , P2_R1312_U130 );
and AND2_14435 ( P2_R1312_U7 , P2_R1312_U131 , P2_R1312_U132 );
and AND4_14436 ( P2_R1312_U8 , P2_R1312_U96 , P2_R1312_U134 , P2_R1312_U136 , P2_R1312_U7 );
and AND2_14437 ( P2_R1312_U9 , P2_R1312_U143 , P2_R1312_U144 );
and AND2_14438 ( P2_R1312_U10 , P2_R1312_U146 , P2_R1312_U145 );
and AND3_14439 ( P2_R1312_U11 , P2_R1312_U99 , P2_R1312_U147 , P2_R1312_U100 );
and AND2_14440 ( P2_R1312_U12 , P2_R1312_U101 , P2_R1312_U11 );
and AND2_14441 ( P2_R1312_U13 , P2_R1312_U162 , P2_R1312_U161 );
and AND2_14442 ( P2_R1312_U14 , P2_R1312_U128 , P2_R1312_U127 );
and AND2_14443 ( P2_R1312_U15 , P2_R1312_U85 , P2_R1312_U20 );
and AND2_14444 ( P2_R1312_U16 , P2_R1312_U87 , P2_R1312_U20 );
and AND2_14445 ( P2_R1312_U17 , P2_R1312_U89 , P2_R1312_U20 );
and AND2_14446 ( P2_R1312_U18 , P2_R1312_U90 , P2_R1312_U20 );
and AND2_14447 ( P2_R1312_U19 , P2_R1312_U119 , P2_R1312_U20 );
and AND2_14448 ( P2_R1312_U20 , P2_R1312_U207 , P2_R1312_U206 );
nand NAND4_14449 ( P2_R1312_U21 , P2_R1312_U204 , P2_R1312_U203 , P2_R1312_U14 , P2_R1312_U120 );
not NOT1_14450 ( P2_R1312_U22 , P2_U3117 );
not NOT1_14451 ( P2_R1312_U23 , P2_U3085 );
not NOT1_14452 ( P2_R1312_U24 , P2_U3118 );
not NOT1_14453 ( P2_R1312_U25 , P2_U3086 );
not NOT1_14454 ( P2_R1312_U26 , P2_U3119 );
not NOT1_14455 ( P2_R1312_U27 , P2_U3087 );
not NOT1_14456 ( P2_R1312_U28 , P2_U3088 );
not NOT1_14457 ( P2_R1312_U29 , P2_U3090 );
not NOT1_14458 ( P2_R1312_U30 , P2_U3089 );
not NOT1_14459 ( P2_R1312_U31 , P2_U3123 );
not NOT1_14460 ( P2_R1312_U32 , P2_U3122 );
not NOT1_14461 ( P2_R1312_U33 , P2_U3121 );
not NOT1_14462 ( P2_R1312_U34 , P2_U3120 );
not NOT1_14463 ( P2_R1312_U35 , P2_U3125 );
not NOT1_14464 ( P2_R1312_U36 , P2_U3124 );
not NOT1_14465 ( P2_R1312_U37 , P2_U3095 );
not NOT1_14466 ( P2_R1312_U38 , P2_U3128 );
not NOT1_14467 ( P2_R1312_U39 , P2_U3096 );
not NOT1_14468 ( P2_R1312_U40 , P2_U3129 );
not NOT1_14469 ( P2_R1312_U41 , P2_U3130 );
not NOT1_14470 ( P2_R1312_U42 , P2_U3099 );
not NOT1_14471 ( P2_R1312_U43 , P2_U3131 );
not NOT1_14472 ( P2_R1312_U44 , P2_U3100 );
not NOT1_14473 ( P2_R1312_U45 , P2_U3098 );
not NOT1_14474 ( P2_R1312_U46 , P2_U3097 );
not NOT1_14475 ( P2_R1312_U47 , P2_U3132 );
not NOT1_14476 ( P2_R1312_U48 , P2_U3133 );
not NOT1_14477 ( P2_R1312_U49 , P2_U3101 );
not NOT1_14478 ( P2_R1312_U50 , P2_U3102 );
not NOT1_14479 ( P2_R1312_U51 , P2_U3142 );
not NOT1_14480 ( P2_R1312_U52 , P2_U3111 );
not NOT1_14481 ( P2_R1312_U53 , P2_U3108 );
not NOT1_14482 ( P2_R1312_U54 , P2_U3107 );
not NOT1_14483 ( P2_R1312_U55 , P2_U3143 );
not NOT1_14484 ( P2_R1312_U56 , P2_U3112 );
not NOT1_14485 ( P2_R1312_U57 , P2_U3110 );
not NOT1_14486 ( P2_R1312_U58 , P2_U3109 );
not NOT1_14487 ( P2_R1312_U59 , P2_U3113 );
not NOT1_14488 ( P2_R1312_U60 , P2_U3114 );
not NOT1_14489 ( P2_R1312_U61 , P2_U3115 );
not NOT1_14490 ( P2_R1312_U62 , P2_U3137 );
not NOT1_14491 ( P2_R1312_U63 , P2_U3136 );
not NOT1_14492 ( P2_R1312_U64 , P2_U3140 );
not NOT1_14493 ( P2_R1312_U65 , P2_U3141 );
not NOT1_14494 ( P2_R1312_U66 , P2_U3147 );
not NOT1_14495 ( P2_R1312_U67 , P2_U3146 );
not NOT1_14496 ( P2_R1312_U68 , P2_U3144 );
not NOT1_14497 ( P2_R1312_U69 , P2_U3145 );
not NOT1_14498 ( P2_R1312_U70 , P2_U3139 );
not NOT1_14499 ( P2_R1312_U71 , P2_U3138 );
not NOT1_14500 ( P2_R1312_U72 , P2_U3105 );
not NOT1_14501 ( P2_R1312_U73 , P2_U3106 );
not NOT1_14502 ( P2_R1312_U74 , P2_U3103 );
not NOT1_14503 ( P2_R1312_U75 , P2_U3104 );
not NOT1_14504 ( P2_R1312_U76 , P2_U3135 );
not NOT1_14505 ( P2_R1312_U77 , P2_U3134 );
not NOT1_14506 ( P2_R1312_U78 , P2_U3127 );
not NOT1_14507 ( P2_R1312_U79 , P2_U3126 );
not NOT1_14508 ( P2_R1312_U80 , P2_U3094 );
not NOT1_14509 ( P2_R1312_U81 , P2_U3093 );
not NOT1_14510 ( P2_R1312_U82 , P2_U3091 );
not NOT1_14511 ( P2_R1312_U83 , P2_U3092 );
and AND2_14512 ( P2_R1312_U84 , P2_R1312_U27 , P2_U3119 );
and AND5_14513 ( P2_R1312_U85 , P2_R1312_U124 , P2_R1312_U82 , P2_U3123 , P2_R1312_U125 , P2_R1312_U123 );
and AND2_14514 ( P2_R1312_U86 , P2_U3122 , P2_R1312_U29 );
and AND3_14515 ( P2_R1312_U87 , P2_R1312_U86 , P2_R1312_U125 , P2_R1312_U123 );
and AND2_14516 ( P2_R1312_U88 , P2_U3121 , P2_R1312_U30 );
and AND2_14517 ( P2_R1312_U89 , P2_R1312_U88 , P2_R1312_U123 );
and AND2_14518 ( P2_R1312_U90 , P2_U3120 , P2_R1312_U28 );
and AND2_14519 ( P2_R1312_U91 , P2_U3128 , P2_R1312_U39 );
and AND2_14520 ( P2_R1312_U92 , P2_U3129 , P2_R1312_U46 );
and AND2_14521 ( P2_R1312_U93 , P2_R1312_U182 , P2_R1312_U181 );
and AND2_14522 ( P2_R1312_U94 , P2_U3099 , P2_R1312_U43 );
and AND2_14523 ( P2_R1312_U95 , P2_U3100 , P2_R1312_U47 );
and AND2_14524 ( P2_R1312_U96 , P2_R1312_U135 , P2_R1312_U133 );
and AND2_14525 ( P2_R1312_U97 , P2_U3111 , P2_R1312_U55 );
and AND2_14526 ( P2_R1312_U98 , P2_U3112 , P2_R1312_U68 );
and AND2_14527 ( P2_R1312_U99 , P2_R1312_U148 , P2_R1312_U142 );
and AND2_14528 ( P2_R1312_U100 , P2_R1312_U9 , P2_R1312_U149 );
and AND2_14529 ( P2_R1312_U101 , P2_R1312_U151 , P2_R1312_U150 );
and AND3_14530 ( P2_R1312_U102 , P2_R1312_U154 , P2_R1312_U155 , P2_R1312_U153 );
and AND2_14531 ( P2_R1312_U103 , P2_U3140 , P2_R1312_U53 );
and AND2_14532 ( P2_R1312_U104 , P2_U3141 , P2_R1312_U58 );
and AND2_14533 ( P2_R1312_U105 , P2_U3147 , P2_R1312_U61 );
and AND2_14534 ( P2_R1312_U106 , P2_U3146 , P2_R1312_U60 );
and AND2_14535 ( P2_R1312_U107 , P2_R1312_U13 , P2_R1312_U108 );
and AND2_14536 ( P2_R1312_U108 , P2_R1312_U167 , P2_R1312_U168 );
and AND2_14537 ( P2_R1312_U109 , P2_R1312_U166 , P2_R1312_U107 );
and AND2_14538 ( P2_R1312_U110 , P2_U3105 , P2_R1312_U62 );
and AND2_14539 ( P2_R1312_U111 , P2_U3106 , P2_R1312_U71 );
and AND2_14540 ( P2_R1312_U112 , P2_R1312_U171 , P2_R1312_U114 );
and AND2_14541 ( P2_R1312_U113 , P2_R1312_U112 , P2_R1312_U172 );
and AND2_14542 ( P2_R1312_U114 , P2_R1312_U174 , P2_R1312_U173 );
and AND3_14543 ( P2_R1312_U115 , P2_R1312_U185 , P2_R1312_U184 , P2_R1312_U138 );
and AND2_14544 ( P2_R1312_U116 , P2_R1312_U117 , P2_R1312_U186 );
and AND2_14545 ( P2_R1312_U117 , P2_R1312_U189 , P2_R1312_U188 );
and AND3_14546 ( P2_R1312_U118 , P2_R1312_U196 , P2_R1312_U194 , P2_R1312_U195 );
and AND5_14547 ( P2_R1312_U119 , P2_R1312_U190 , P2_R1312_U124 , P2_R1312_U118 , P2_R1312_U125 , P2_R1312_U123 );
and AND4_14548 ( P2_R1312_U120 , P2_R1312_U202 , P2_R1312_U201 , P2_R1312_U200 , P2_R1312_U199 );
nand NAND2_14549 ( P2_R1312_U121 , P2_R1312_U198 , P2_R1312_U197 );
nand NAND2_14550 ( P2_R1312_U122 , P2_U3087 , P2_R1312_U26 );
nand NAND2_14551 ( P2_R1312_U123 , P2_U3088 , P2_R1312_U34 );
nand NAND2_14552 ( P2_R1312_U124 , P2_U3090 , P2_R1312_U32 );
nand NAND2_14553 ( P2_R1312_U125 , P2_U3089 , P2_R1312_U33 );
nand NAND2_14554 ( P2_R1312_U126 , P2_U3086 , P2_R1312_U24 );
nand NAND3_14555 ( P2_R1312_U127 , P2_R1312_U209 , P2_R1312_U208 , P2_R1312_U205 );
nand NAND3_14556 ( P2_R1312_U128 , P2_R1312_U20 , P2_U3118 , P2_R1312_U25 );
nand NAND2_14557 ( P2_R1312_U129 , P2_U3130 , P2_R1312_U45 );
nand NAND2_14558 ( P2_R1312_U130 , P2_U3131 , P2_R1312_U42 );
nand NAND2_14559 ( P2_R1312_U131 , P2_U3095 , P2_R1312_U78 );
nand NAND2_14560 ( P2_R1312_U132 , P2_U3096 , P2_R1312_U38 );
nand NAND2_14561 ( P2_R1312_U133 , P2_R1312_U94 , P2_R1312_U129 );
nand NAND2_14562 ( P2_R1312_U134 , P2_R1312_U95 , P2_R1312_U6 );
nand NAND2_14563 ( P2_R1312_U135 , P2_U3098 , P2_R1312_U41 );
nand NAND2_14564 ( P2_R1312_U136 , P2_U3097 , P2_R1312_U40 );
nand NAND2_14565 ( P2_R1312_U137 , P2_U3101 , P2_R1312_U48 );
nand NAND2_14566 ( P2_R1312_U138 , P2_U3125 , P2_R1312_U81 );
nand NAND2_14567 ( P2_R1312_U139 , P2_U3124 , P2_R1312_U83 );
nand NAND2_14568 ( P2_R1312_U140 , P2_U3102 , P2_R1312_U77 );
nand NAND2_14569 ( P2_R1312_U141 , P2_U3142 , P2_R1312_U57 );
nand NAND2_14570 ( P2_R1312_U142 , P2_R1312_U97 , P2_R1312_U141 );
nand NAND2_14571 ( P2_R1312_U143 , P2_U3107 , P2_R1312_U70 );
nand NAND2_14572 ( P2_R1312_U144 , P2_U3108 , P2_R1312_U64 );
nand NAND2_14573 ( P2_R1312_U145 , P2_U3143 , P2_R1312_U52 );
nand NAND2_14574 ( P2_R1312_U146 , P2_U3142 , P2_R1312_U57 );
nand NAND2_14575 ( P2_R1312_U147 , P2_R1312_U98 , P2_R1312_U10 );
nand NAND2_14576 ( P2_R1312_U148 , P2_U3110 , P2_R1312_U51 );
nand NAND2_14577 ( P2_R1312_U149 , P2_U3109 , P2_R1312_U65 );
nand NAND2_14578 ( P2_R1312_U150 , P2_U3113 , P2_R1312_U69 );
nand NAND2_14579 ( P2_R1312_U151 , P2_U3114 , P2_R1312_U67 );
nand NAND2_14580 ( P2_R1312_U152 , P2_U3148 , P2_U3149 );
nand NAND2_14581 ( P2_R1312_U153 , P2_U3116 , P2_R1312_U152 );
or OR2_14582 ( P2_R1312_U154 , P2_U3148 , P2_U3149 );
nand NAND2_14583 ( P2_R1312_U155 , P2_U3115 , P2_R1312_U66 );
nand NAND2_14584 ( P2_R1312_U156 , P2_R1312_U102 , P2_R1312_U12 );
nand NAND2_14585 ( P2_R1312_U157 , P2_R1312_U106 , P2_R1312_U150 );
nand NAND2_14586 ( P2_R1312_U158 , P2_U3144 , P2_R1312_U56 );
nand NAND2_14587 ( P2_R1312_U159 , P2_U3145 , P2_R1312_U59 );
nand NAND4_14588 ( P2_R1312_U160 , P2_R1312_U10 , P2_R1312_U159 , P2_R1312_U158 , P2_R1312_U157 );
nand NAND2_14589 ( P2_R1312_U161 , P2_U3137 , P2_R1312_U72 );
nand NAND2_14590 ( P2_R1312_U162 , P2_U3136 , P2_R1312_U75 );
nand NAND2_14591 ( P2_R1312_U163 , P2_R1312_U103 , P2_R1312_U143 );
nand NAND2_14592 ( P2_R1312_U164 , P2_R1312_U104 , P2_R1312_U9 );
nand NAND2_14593 ( P2_R1312_U165 , P2_R1312_U105 , P2_R1312_U12 );
nand NAND2_14594 ( P2_R1312_U166 , P2_R1312_U11 , P2_R1312_U160 );
nand NAND2_14595 ( P2_R1312_U167 , P2_U3139 , P2_R1312_U54 );
nand NAND2_14596 ( P2_R1312_U168 , P2_U3138 , P2_R1312_U73 );
nand NAND5_14597 ( P2_R1312_U169 , P2_R1312_U165 , P2_R1312_U164 , P2_R1312_U163 , P2_R1312_U156 , P2_R1312_U109 );
nand NAND2_14598 ( P2_R1312_U170 , P2_U3136 , P2_R1312_U75 );
nand NAND2_14599 ( P2_R1312_U171 , P2_R1312_U110 , P2_R1312_U170 );
nand NAND2_14600 ( P2_R1312_U172 , P2_R1312_U111 , P2_R1312_U13 );
nand NAND2_14601 ( P2_R1312_U173 , P2_U3103 , P2_R1312_U76 );
nand NAND2_14602 ( P2_R1312_U174 , P2_U3104 , P2_R1312_U63 );
nand NAND2_14603 ( P2_R1312_U175 , P2_R1312_U169 , P2_R1312_U113 );
nand NAND2_14604 ( P2_R1312_U176 , P2_U3135 , P2_R1312_U74 );
nand NAND2_14605 ( P2_R1312_U177 , P2_R1312_U176 , P2_R1312_U175 );
nand NAND2_14606 ( P2_R1312_U178 , P2_R1312_U177 , P2_R1312_U140 );
nand NAND2_14607 ( P2_R1312_U179 , P2_U3134 , P2_R1312_U50 );
nand NAND2_14608 ( P2_R1312_U180 , P2_R1312_U179 , P2_R1312_U178 );
nand NAND2_14609 ( P2_R1312_U181 , P2_U3132 , P2_R1312_U44 );
nand NAND2_14610 ( P2_R1312_U182 , P2_U3133 , P2_R1312_U49 );
nand NAND2_14611 ( P2_R1312_U183 , P2_R1312_U93 , P2_R1312_U6 );
nand NAND2_14612 ( P2_R1312_U184 , P2_R1312_U91 , P2_R1312_U131 );
nand NAND2_14613 ( P2_R1312_U185 , P2_R1312_U92 , P2_R1312_U7 );
nand NAND2_14614 ( P2_R1312_U186 , P2_R1312_U8 , P2_R1312_U183 );
nand NAND3_14615 ( P2_R1312_U187 , P2_R1312_U180 , P2_R1312_U137 , P2_R1312_U8 );
nand NAND2_14616 ( P2_R1312_U188 , P2_U3127 , P2_R1312_U37 );
nand NAND2_14617 ( P2_R1312_U189 , P2_U3126 , P2_R1312_U80 );
nand NAND4_14618 ( P2_R1312_U190 , P2_R1312_U187 , P2_R1312_U116 , P2_R1312_U115 , P2_R1312_U139 );
nand NAND2_14619 ( P2_R1312_U191 , P2_U3094 , P2_R1312_U79 );
nand NAND2_14620 ( P2_R1312_U192 , P2_U3093 , P2_R1312_U35 );
nand NAND2_14621 ( P2_R1312_U193 , P2_R1312_U192 , P2_R1312_U191 );
nand NAND3_14622 ( P2_R1312_U194 , P2_R1312_U193 , P2_R1312_U138 , P2_R1312_U139 );
nand NAND2_14623 ( P2_R1312_U195 , P2_U3091 , P2_R1312_U31 );
nand NAND2_14624 ( P2_R1312_U196 , P2_U3092 , P2_R1312_U36 );
nand NAND2_14625 ( P2_R1312_U197 , P2_U3118 , P2_R1312_U122 );
nand NAND2_14626 ( P2_R1312_U198 , P2_R1312_U122 , P2_R1312_U25 );
nand NAND3_14627 ( P2_R1312_U199 , P2_R1312_U84 , P2_R1312_U20 , P2_R1312_U126 );
nand NAND2_14628 ( P2_R1312_U200 , P2_R1312_U15 , P2_R1312_U121 );
nand NAND2_14629 ( P2_R1312_U201 , P2_R1312_U16 , P2_R1312_U121 );
nand NAND2_14630 ( P2_R1312_U202 , P2_R1312_U17 , P2_R1312_U121 );
nand NAND2_14631 ( P2_R1312_U203 , P2_R1312_U18 , P2_R1312_U121 );
nand NAND2_14632 ( P2_R1312_U204 , P2_R1312_U19 , P2_R1312_U121 );
nand NAND2_14633 ( P2_R1312_U205 , P2_U3085 , P2_U3117 );
nand NAND2_14634 ( P2_R1312_U206 , P2_U3085 , P2_R1312_U22 );
nand NAND2_14635 ( P2_R1312_U207 , P2_U3117 , P2_R1312_U23 );
or OR2_14636 ( P2_R1312_U208 , P2_U3150 , P2_U3117 );
nand NAND2_14637 ( P2_R1312_U209 , P2_U3150 , P2_R1312_U23 );
not NOT1_14638 ( P2_R1335_U6 , P2_U3059 );
not NOT1_14639 ( P2_R1335_U7 , P2_U3056 );
and AND2_14640 ( P2_R1335_U8 , P2_R1335_U10 , P2_R1335_U9 );
nand NAND2_14641 ( P2_R1335_U9 , P2_U3056 , P2_R1335_U6 );
nand NAND2_14642 ( P2_R1335_U10 , P2_U3059 , P2_R1335_U7 );
and AND2_14643 ( P2_R1209_U4 , P2_R1209_U95 , P2_R1209_U94 );
and AND2_14644 ( P2_R1209_U5 , P2_R1209_U96 , P2_R1209_U97 );
and AND2_14645 ( P2_R1209_U6 , P2_R1209_U113 , P2_R1209_U112 );
and AND2_14646 ( P2_R1209_U7 , P2_R1209_U155 , P2_R1209_U154 );
and AND2_14647 ( P2_R1209_U8 , P2_R1209_U164 , P2_R1209_U163 );
and AND2_14648 ( P2_R1209_U9 , P2_R1209_U182 , P2_R1209_U181 );
and AND2_14649 ( P2_R1209_U10 , P2_R1209_U218 , P2_R1209_U215 );
and AND2_14650 ( P2_R1209_U11 , P2_R1209_U211 , P2_R1209_U208 );
and AND2_14651 ( P2_R1209_U12 , P2_R1209_U202 , P2_R1209_U199 );
and AND2_14652 ( P2_R1209_U13 , P2_R1209_U196 , P2_R1209_U192 );
and AND2_14653 ( P2_R1209_U14 , P2_R1209_U151 , P2_R1209_U148 );
and AND2_14654 ( P2_R1209_U15 , P2_R1209_U143 , P2_R1209_U140 );
and AND2_14655 ( P2_R1209_U16 , P2_R1209_U129 , P2_R1209_U126 );
not NOT1_14656 ( P2_R1209_U17 , P2_REG1_REG_6_ );
not NOT1_14657 ( P2_R1209_U18 , P2_U3467 );
not NOT1_14658 ( P2_R1209_U19 , P2_U3470 );
nand NAND2_14659 ( P2_R1209_U20 , P2_U3467 , P2_REG1_REG_6_ );
not NOT1_14660 ( P2_R1209_U21 , P2_REG1_REG_7_ );
not NOT1_14661 ( P2_R1209_U22 , P2_REG1_REG_4_ );
not NOT1_14662 ( P2_R1209_U23 , P2_U3461 );
not NOT1_14663 ( P2_R1209_U24 , P2_U3464 );
not NOT1_14664 ( P2_R1209_U25 , P2_REG1_REG_2_ );
not NOT1_14665 ( P2_R1209_U26 , P2_U3455 );
not NOT1_14666 ( P2_R1209_U27 , P2_REG1_REG_0_ );
not NOT1_14667 ( P2_R1209_U28 , P2_U3446 );
nand NAND2_14668 ( P2_R1209_U29 , P2_U3446 , P2_REG1_REG_0_ );
not NOT1_14669 ( P2_R1209_U30 , P2_REG1_REG_3_ );
not NOT1_14670 ( P2_R1209_U31 , P2_U3458 );
nand NAND2_14671 ( P2_R1209_U32 , P2_U3461 , P2_REG1_REG_4_ );
not NOT1_14672 ( P2_R1209_U33 , P2_REG1_REG_5_ );
not NOT1_14673 ( P2_R1209_U34 , P2_REG1_REG_8_ );
not NOT1_14674 ( P2_R1209_U35 , P2_U3473 );
not NOT1_14675 ( P2_R1209_U36 , P2_U3476 );
not NOT1_14676 ( P2_R1209_U37 , P2_REG1_REG_9_ );
nand NAND2_14677 ( P2_R1209_U38 , P2_R1209_U49 , P2_R1209_U121 );
nand NAND3_14678 ( P2_R1209_U39 , P2_R1209_U110 , P2_R1209_U108 , P2_R1209_U109 );
nand NAND2_14679 ( P2_R1209_U40 , P2_R1209_U98 , P2_R1209_U99 );
nand NAND2_14680 ( P2_R1209_U41 , P2_REG1_REG_1_ , P2_U3452 );
nand NAND3_14681 ( P2_R1209_U42 , P2_R1209_U136 , P2_R1209_U134 , P2_R1209_U135 );
nand NAND2_14682 ( P2_R1209_U43 , P2_R1209_U132 , P2_R1209_U131 );
not NOT1_14683 ( P2_R1209_U44 , P2_REG1_REG_16_ );
not NOT1_14684 ( P2_R1209_U45 , P2_U3497 );
not NOT1_14685 ( P2_R1209_U46 , P2_U3500 );
nand NAND2_14686 ( P2_R1209_U47 , P2_U3497 , P2_REG1_REG_16_ );
not NOT1_14687 ( P2_R1209_U48 , P2_REG1_REG_17_ );
nand NAND2_14688 ( P2_R1209_U49 , P2_U3473 , P2_REG1_REG_8_ );
not NOT1_14689 ( P2_R1209_U50 , P2_REG1_REG_10_ );
not NOT1_14690 ( P2_R1209_U51 , P2_U3479 );
not NOT1_14691 ( P2_R1209_U52 , P2_REG1_REG_12_ );
not NOT1_14692 ( P2_R1209_U53 , P2_U3485 );
not NOT1_14693 ( P2_R1209_U54 , P2_REG1_REG_11_ );
not NOT1_14694 ( P2_R1209_U55 , P2_U3482 );
nand NAND2_14695 ( P2_R1209_U56 , P2_U3482 , P2_REG1_REG_11_ );
not NOT1_14696 ( P2_R1209_U57 , P2_REG1_REG_13_ );
not NOT1_14697 ( P2_R1209_U58 , P2_U3488 );
not NOT1_14698 ( P2_R1209_U59 , P2_REG1_REG_14_ );
not NOT1_14699 ( P2_R1209_U60 , P2_U3491 );
not NOT1_14700 ( P2_R1209_U61 , P2_REG1_REG_15_ );
not NOT1_14701 ( P2_R1209_U62 , P2_U3494 );
not NOT1_14702 ( P2_R1209_U63 , P2_REG1_REG_18_ );
not NOT1_14703 ( P2_R1209_U64 , P2_U3503 );
nand NAND3_14704 ( P2_R1209_U65 , P2_R1209_U186 , P2_R1209_U185 , P2_R1209_U187 );
nand NAND2_14705 ( P2_R1209_U66 , P2_R1209_U179 , P2_R1209_U178 );
nand NAND2_14706 ( P2_R1209_U67 , P2_R1209_U56 , P2_R1209_U204 );
nand NAND2_14707 ( P2_R1209_U68 , P2_R1209_U259 , P2_R1209_U258 );
nand NAND2_14708 ( P2_R1209_U69 , P2_R1209_U308 , P2_R1209_U307 );
nand NAND2_14709 ( P2_R1209_U70 , P2_R1209_U231 , P2_R1209_U230 );
nand NAND2_14710 ( P2_R1209_U71 , P2_R1209_U236 , P2_R1209_U235 );
nand NAND2_14711 ( P2_R1209_U72 , P2_R1209_U243 , P2_R1209_U242 );
nand NAND2_14712 ( P2_R1209_U73 , P2_R1209_U250 , P2_R1209_U249 );
nand NAND2_14713 ( P2_R1209_U74 , P2_R1209_U255 , P2_R1209_U254 );
nand NAND2_14714 ( P2_R1209_U75 , P2_R1209_U271 , P2_R1209_U270 );
nand NAND2_14715 ( P2_R1209_U76 , P2_R1209_U278 , P2_R1209_U277 );
nand NAND2_14716 ( P2_R1209_U77 , P2_R1209_U285 , P2_R1209_U284 );
nand NAND2_14717 ( P2_R1209_U78 , P2_R1209_U292 , P2_R1209_U291 );
nand NAND2_14718 ( P2_R1209_U79 , P2_R1209_U299 , P2_R1209_U298 );
nand NAND2_14719 ( P2_R1209_U80 , P2_R1209_U304 , P2_R1209_U303 );
nand NAND3_14720 ( P2_R1209_U81 , P2_R1209_U117 , P2_R1209_U116 , P2_R1209_U118 );
nand NAND2_14721 ( P2_R1209_U82 , P2_R1209_U133 , P2_R1209_U145 );
nand NAND2_14722 ( P2_R1209_U83 , P2_R1209_U41 , P2_R1209_U152 );
not NOT1_14723 ( P2_R1209_U84 , P2_U3445 );
not NOT1_14724 ( P2_R1209_U85 , P2_REG1_REG_19_ );
nand NAND2_14725 ( P2_R1209_U86 , P2_R1209_U175 , P2_R1209_U174 );
nand NAND2_14726 ( P2_R1209_U87 , P2_R1209_U171 , P2_R1209_U170 );
nand NAND2_14727 ( P2_R1209_U88 , P2_R1209_U161 , P2_R1209_U160 );
not NOT1_14728 ( P2_R1209_U89 , P2_R1209_U32 );
nand NAND2_14729 ( P2_R1209_U90 , P2_REG1_REG_9_ , P2_U3476 );
nand NAND2_14730 ( P2_R1209_U91 , P2_U3485 , P2_REG1_REG_12_ );
not NOT1_14731 ( P2_R1209_U92 , P2_R1209_U56 );
not NOT1_14732 ( P2_R1209_U93 , P2_R1209_U49 );
or OR2_14733 ( P2_R1209_U94 , P2_U3464 , P2_REG1_REG_5_ );
or OR2_14734 ( P2_R1209_U95 , P2_U3461 , P2_REG1_REG_4_ );
or OR2_14735 ( P2_R1209_U96 , P2_REG1_REG_3_ , P2_U3458 );
or OR2_14736 ( P2_R1209_U97 , P2_REG1_REG_2_ , P2_U3455 );
not NOT1_14737 ( P2_R1209_U98 , P2_R1209_U29 );
or OR2_14738 ( P2_R1209_U99 , P2_REG1_REG_1_ , P2_U3452 );
not NOT1_14739 ( P2_R1209_U100 , P2_R1209_U40 );
not NOT1_14740 ( P2_R1209_U101 , P2_R1209_U41 );
nand NAND2_14741 ( P2_R1209_U102 , P2_R1209_U40 , P2_R1209_U41 );
nand NAND3_14742 ( P2_R1209_U103 , P2_REG1_REG_2_ , P2_U3455 , P2_R1209_U96 );
nand NAND2_14743 ( P2_R1209_U104 , P2_R1209_U5 , P2_R1209_U102 );
nand NAND2_14744 ( P2_R1209_U105 , P2_U3458 , P2_REG1_REG_3_ );
nand NAND3_14745 ( P2_R1209_U106 , P2_R1209_U105 , P2_R1209_U103 , P2_R1209_U104 );
nand NAND2_14746 ( P2_R1209_U107 , P2_R1209_U33 , P2_R1209_U32 );
nand NAND2_14747 ( P2_R1209_U108 , P2_U3464 , P2_R1209_U107 );
nand NAND2_14748 ( P2_R1209_U109 , P2_R1209_U4 , P2_R1209_U106 );
nand NAND2_14749 ( P2_R1209_U110 , P2_REG1_REG_5_ , P2_R1209_U89 );
not NOT1_14750 ( P2_R1209_U111 , P2_R1209_U39 );
or OR2_14751 ( P2_R1209_U112 , P2_U3470 , P2_REG1_REG_7_ );
or OR2_14752 ( P2_R1209_U113 , P2_U3467 , P2_REG1_REG_6_ );
not NOT1_14753 ( P2_R1209_U114 , P2_R1209_U20 );
nand NAND2_14754 ( P2_R1209_U115 , P2_R1209_U21 , P2_R1209_U20 );
nand NAND2_14755 ( P2_R1209_U116 , P2_U3470 , P2_R1209_U115 );
nand NAND2_14756 ( P2_R1209_U117 , P2_REG1_REG_7_ , P2_R1209_U114 );
nand NAND2_14757 ( P2_R1209_U118 , P2_R1209_U6 , P2_R1209_U39 );
not NOT1_14758 ( P2_R1209_U119 , P2_R1209_U81 );
or OR2_14759 ( P2_R1209_U120 , P2_REG1_REG_8_ , P2_U3473 );
nand NAND2_14760 ( P2_R1209_U121 , P2_R1209_U120 , P2_R1209_U81 );
not NOT1_14761 ( P2_R1209_U122 , P2_R1209_U38 );
or OR2_14762 ( P2_R1209_U123 , P2_U3476 , P2_REG1_REG_9_ );
or OR2_14763 ( P2_R1209_U124 , P2_REG1_REG_6_ , P2_U3467 );
nand NAND2_14764 ( P2_R1209_U125 , P2_R1209_U124 , P2_R1209_U39 );
nand NAND4_14765 ( P2_R1209_U126 , P2_R1209_U238 , P2_R1209_U237 , P2_R1209_U20 , P2_R1209_U125 );
nand NAND2_14766 ( P2_R1209_U127 , P2_R1209_U111 , P2_R1209_U20 );
nand NAND2_14767 ( P2_R1209_U128 , P2_REG1_REG_7_ , P2_U3470 );
nand NAND3_14768 ( P2_R1209_U129 , P2_R1209_U128 , P2_R1209_U6 , P2_R1209_U127 );
or OR2_14769 ( P2_R1209_U130 , P2_U3467 , P2_REG1_REG_6_ );
nand NAND2_14770 ( P2_R1209_U131 , P2_R1209_U101 , P2_R1209_U97 );
nand NAND2_14771 ( P2_R1209_U132 , P2_U3455 , P2_REG1_REG_2_ );
not NOT1_14772 ( P2_R1209_U133 , P2_R1209_U43 );
nand NAND2_14773 ( P2_R1209_U134 , P2_R1209_U100 , P2_R1209_U5 );
nand NAND2_14774 ( P2_R1209_U135 , P2_R1209_U43 , P2_R1209_U96 );
nand NAND2_14775 ( P2_R1209_U136 , P2_U3458 , P2_REG1_REG_3_ );
not NOT1_14776 ( P2_R1209_U137 , P2_R1209_U42 );
or OR2_14777 ( P2_R1209_U138 , P2_REG1_REG_4_ , P2_U3461 );
nand NAND2_14778 ( P2_R1209_U139 , P2_R1209_U138 , P2_R1209_U42 );
nand NAND4_14779 ( P2_R1209_U140 , P2_R1209_U245 , P2_R1209_U244 , P2_R1209_U32 , P2_R1209_U139 );
nand NAND2_14780 ( P2_R1209_U141 , P2_R1209_U137 , P2_R1209_U32 );
nand NAND2_14781 ( P2_R1209_U142 , P2_REG1_REG_5_ , P2_U3464 );
nand NAND3_14782 ( P2_R1209_U143 , P2_R1209_U142 , P2_R1209_U4 , P2_R1209_U141 );
or OR2_14783 ( P2_R1209_U144 , P2_U3461 , P2_REG1_REG_4_ );
nand NAND2_14784 ( P2_R1209_U145 , P2_R1209_U100 , P2_R1209_U97 );
not NOT1_14785 ( P2_R1209_U146 , P2_R1209_U82 );
nand NAND2_14786 ( P2_R1209_U147 , P2_U3458 , P2_REG1_REG_3_ );
nand NAND4_14787 ( P2_R1209_U148 , P2_R1209_U257 , P2_R1209_U256 , P2_R1209_U41 , P2_R1209_U40 );
nand NAND2_14788 ( P2_R1209_U149 , P2_R1209_U41 , P2_R1209_U40 );
nand NAND2_14789 ( P2_R1209_U150 , P2_U3455 , P2_REG1_REG_2_ );
nand NAND3_14790 ( P2_R1209_U151 , P2_R1209_U150 , P2_R1209_U97 , P2_R1209_U149 );
or OR2_14791 ( P2_R1209_U152 , P2_REG1_REG_1_ , P2_U3452 );
not NOT1_14792 ( P2_R1209_U153 , P2_R1209_U83 );
or OR2_14793 ( P2_R1209_U154 , P2_U3476 , P2_REG1_REG_9_ );
or OR2_14794 ( P2_R1209_U155 , P2_U3479 , P2_REG1_REG_10_ );
nand NAND2_14795 ( P2_R1209_U156 , P2_R1209_U93 , P2_R1209_U7 );
nand NAND2_14796 ( P2_R1209_U157 , P2_U3479 , P2_REG1_REG_10_ );
nand NAND3_14797 ( P2_R1209_U158 , P2_R1209_U157 , P2_R1209_U90 , P2_R1209_U156 );
or OR2_14798 ( P2_R1209_U159 , P2_REG1_REG_10_ , P2_U3479 );
nand NAND3_14799 ( P2_R1209_U160 , P2_R1209_U120 , P2_R1209_U7 , P2_R1209_U81 );
nand NAND2_14800 ( P2_R1209_U161 , P2_R1209_U159 , P2_R1209_U158 );
not NOT1_14801 ( P2_R1209_U162 , P2_R1209_U88 );
or OR2_14802 ( P2_R1209_U163 , P2_U3488 , P2_REG1_REG_13_ );
or OR2_14803 ( P2_R1209_U164 , P2_U3485 , P2_REG1_REG_12_ );
nand NAND2_14804 ( P2_R1209_U165 , P2_R1209_U92 , P2_R1209_U8 );
nand NAND2_14805 ( P2_R1209_U166 , P2_U3488 , P2_REG1_REG_13_ );
nand NAND3_14806 ( P2_R1209_U167 , P2_R1209_U166 , P2_R1209_U91 , P2_R1209_U165 );
or OR2_14807 ( P2_R1209_U168 , P2_REG1_REG_11_ , P2_U3482 );
or OR2_14808 ( P2_R1209_U169 , P2_REG1_REG_13_ , P2_U3488 );
nand NAND3_14809 ( P2_R1209_U170 , P2_R1209_U168 , P2_R1209_U8 , P2_R1209_U88 );
nand NAND2_14810 ( P2_R1209_U171 , P2_R1209_U169 , P2_R1209_U167 );
not NOT1_14811 ( P2_R1209_U172 , P2_R1209_U87 );
or OR2_14812 ( P2_R1209_U173 , P2_REG1_REG_14_ , P2_U3491 );
nand NAND2_14813 ( P2_R1209_U174 , P2_R1209_U173 , P2_R1209_U87 );
nand NAND2_14814 ( P2_R1209_U175 , P2_U3491 , P2_REG1_REG_14_ );
not NOT1_14815 ( P2_R1209_U176 , P2_R1209_U86 );
or OR2_14816 ( P2_R1209_U177 , P2_REG1_REG_15_ , P2_U3494 );
nand NAND2_14817 ( P2_R1209_U178 , P2_R1209_U177 , P2_R1209_U86 );
nand NAND2_14818 ( P2_R1209_U179 , P2_U3494 , P2_REG1_REG_15_ );
not NOT1_14819 ( P2_R1209_U180 , P2_R1209_U66 );
or OR2_14820 ( P2_R1209_U181 , P2_U3500 , P2_REG1_REG_17_ );
or OR2_14821 ( P2_R1209_U182 , P2_U3497 , P2_REG1_REG_16_ );
not NOT1_14822 ( P2_R1209_U183 , P2_R1209_U47 );
nand NAND2_14823 ( P2_R1209_U184 , P2_R1209_U48 , P2_R1209_U47 );
nand NAND2_14824 ( P2_R1209_U185 , P2_U3500 , P2_R1209_U184 );
nand NAND2_14825 ( P2_R1209_U186 , P2_REG1_REG_17_ , P2_R1209_U183 );
nand NAND2_14826 ( P2_R1209_U187 , P2_R1209_U9 , P2_R1209_U66 );
not NOT1_14827 ( P2_R1209_U188 , P2_R1209_U65 );
or OR2_14828 ( P2_R1209_U189 , P2_REG1_REG_18_ , P2_U3503 );
nand NAND2_14829 ( P2_R1209_U190 , P2_R1209_U189 , P2_R1209_U65 );
nand NAND2_14830 ( P2_R1209_U191 , P2_U3503 , P2_REG1_REG_18_ );
nand NAND4_14831 ( P2_R1209_U192 , P2_R1209_U261 , P2_R1209_U260 , P2_R1209_U191 , P2_R1209_U190 );
nand NAND2_14832 ( P2_R1209_U193 , P2_U3503 , P2_REG1_REG_18_ );
nand NAND2_14833 ( P2_R1209_U194 , P2_R1209_U188 , P2_R1209_U193 );
or OR2_14834 ( P2_R1209_U195 , P2_U3503 , P2_REG1_REG_18_ );
nand NAND3_14835 ( P2_R1209_U196 , P2_R1209_U195 , P2_R1209_U264 , P2_R1209_U194 );
or OR2_14836 ( P2_R1209_U197 , P2_REG1_REG_16_ , P2_U3497 );
nand NAND2_14837 ( P2_R1209_U198 , P2_R1209_U197 , P2_R1209_U66 );
nand NAND4_14838 ( P2_R1209_U199 , P2_R1209_U273 , P2_R1209_U272 , P2_R1209_U47 , P2_R1209_U198 );
nand NAND2_14839 ( P2_R1209_U200 , P2_R1209_U180 , P2_R1209_U47 );
nand NAND2_14840 ( P2_R1209_U201 , P2_REG1_REG_17_ , P2_U3500 );
nand NAND3_14841 ( P2_R1209_U202 , P2_R1209_U201 , P2_R1209_U9 , P2_R1209_U200 );
or OR2_14842 ( P2_R1209_U203 , P2_U3497 , P2_REG1_REG_16_ );
nand NAND2_14843 ( P2_R1209_U204 , P2_R1209_U168 , P2_R1209_U88 );
not NOT1_14844 ( P2_R1209_U205 , P2_R1209_U67 );
or OR2_14845 ( P2_R1209_U206 , P2_REG1_REG_12_ , P2_U3485 );
nand NAND2_14846 ( P2_R1209_U207 , P2_R1209_U206 , P2_R1209_U67 );
nand NAND4_14847 ( P2_R1209_U208 , P2_R1209_U294 , P2_R1209_U293 , P2_R1209_U91 , P2_R1209_U207 );
nand NAND2_14848 ( P2_R1209_U209 , P2_R1209_U205 , P2_R1209_U91 );
nand NAND2_14849 ( P2_R1209_U210 , P2_U3488 , P2_REG1_REG_13_ );
nand NAND3_14850 ( P2_R1209_U211 , P2_R1209_U210 , P2_R1209_U8 , P2_R1209_U209 );
or OR2_14851 ( P2_R1209_U212 , P2_U3485 , P2_REG1_REG_12_ );
or OR2_14852 ( P2_R1209_U213 , P2_REG1_REG_9_ , P2_U3476 );
nand NAND2_14853 ( P2_R1209_U214 , P2_R1209_U213 , P2_R1209_U38 );
nand NAND4_14854 ( P2_R1209_U215 , P2_R1209_U306 , P2_R1209_U305 , P2_R1209_U90 , P2_R1209_U214 );
nand NAND2_14855 ( P2_R1209_U216 , P2_R1209_U122 , P2_R1209_U90 );
nand NAND2_14856 ( P2_R1209_U217 , P2_U3479 , P2_REG1_REG_10_ );
nand NAND3_14857 ( P2_R1209_U218 , P2_R1209_U217 , P2_R1209_U7 , P2_R1209_U216 );
nand NAND2_14858 ( P2_R1209_U219 , P2_R1209_U123 , P2_R1209_U90 );
nand NAND2_14859 ( P2_R1209_U220 , P2_R1209_U120 , P2_R1209_U49 );
nand NAND2_14860 ( P2_R1209_U221 , P2_R1209_U130 , P2_R1209_U20 );
nand NAND2_14861 ( P2_R1209_U222 , P2_R1209_U144 , P2_R1209_U32 );
nand NAND2_14862 ( P2_R1209_U223 , P2_R1209_U147 , P2_R1209_U96 );
nand NAND2_14863 ( P2_R1209_U224 , P2_R1209_U203 , P2_R1209_U47 );
nand NAND2_14864 ( P2_R1209_U225 , P2_R1209_U212 , P2_R1209_U91 );
nand NAND2_14865 ( P2_R1209_U226 , P2_R1209_U168 , P2_R1209_U56 );
nand NAND2_14866 ( P2_R1209_U227 , P2_U3476 , P2_R1209_U37 );
nand NAND2_14867 ( P2_R1209_U228 , P2_REG1_REG_9_ , P2_R1209_U36 );
nand NAND2_14868 ( P2_R1209_U229 , P2_R1209_U228 , P2_R1209_U227 );
nand NAND2_14869 ( P2_R1209_U230 , P2_R1209_U219 , P2_R1209_U38 );
nand NAND2_14870 ( P2_R1209_U231 , P2_R1209_U229 , P2_R1209_U122 );
nand NAND2_14871 ( P2_R1209_U232 , P2_U3473 , P2_R1209_U34 );
nand NAND2_14872 ( P2_R1209_U233 , P2_REG1_REG_8_ , P2_R1209_U35 );
nand NAND2_14873 ( P2_R1209_U234 , P2_R1209_U233 , P2_R1209_U232 );
nand NAND2_14874 ( P2_R1209_U235 , P2_R1209_U220 , P2_R1209_U81 );
nand NAND2_14875 ( P2_R1209_U236 , P2_R1209_U119 , P2_R1209_U234 );
nand NAND2_14876 ( P2_R1209_U237 , P2_U3470 , P2_R1209_U21 );
nand NAND2_14877 ( P2_R1209_U238 , P2_REG1_REG_7_ , P2_R1209_U19 );
nand NAND2_14878 ( P2_R1209_U239 , P2_U3467 , P2_R1209_U17 );
nand NAND2_14879 ( P2_R1209_U240 , P2_REG1_REG_6_ , P2_R1209_U18 );
nand NAND2_14880 ( P2_R1209_U241 , P2_R1209_U240 , P2_R1209_U239 );
nand NAND2_14881 ( P2_R1209_U242 , P2_R1209_U221 , P2_R1209_U39 );
nand NAND2_14882 ( P2_R1209_U243 , P2_R1209_U241 , P2_R1209_U111 );
nand NAND2_14883 ( P2_R1209_U244 , P2_U3464 , P2_R1209_U33 );
nand NAND2_14884 ( P2_R1209_U245 , P2_REG1_REG_5_ , P2_R1209_U24 );
nand NAND2_14885 ( P2_R1209_U246 , P2_U3461 , P2_R1209_U22 );
nand NAND2_14886 ( P2_R1209_U247 , P2_REG1_REG_4_ , P2_R1209_U23 );
nand NAND2_14887 ( P2_R1209_U248 , P2_R1209_U247 , P2_R1209_U246 );
nand NAND2_14888 ( P2_R1209_U249 , P2_R1209_U222 , P2_R1209_U42 );
nand NAND2_14889 ( P2_R1209_U250 , P2_R1209_U248 , P2_R1209_U137 );
nand NAND2_14890 ( P2_R1209_U251 , P2_U3458 , P2_R1209_U30 );
nand NAND2_14891 ( P2_R1209_U252 , P2_REG1_REG_3_ , P2_R1209_U31 );
nand NAND2_14892 ( P2_R1209_U253 , P2_R1209_U252 , P2_R1209_U251 );
nand NAND2_14893 ( P2_R1209_U254 , P2_R1209_U223 , P2_R1209_U82 );
nand NAND2_14894 ( P2_R1209_U255 , P2_R1209_U146 , P2_R1209_U253 );
nand NAND2_14895 ( P2_R1209_U256 , P2_U3455 , P2_R1209_U25 );
nand NAND2_14896 ( P2_R1209_U257 , P2_REG1_REG_2_ , P2_R1209_U26 );
nand NAND2_14897 ( P2_R1209_U258 , P2_R1209_U98 , P2_R1209_U83 );
nand NAND2_14898 ( P2_R1209_U259 , P2_R1209_U153 , P2_R1209_U29 );
nand NAND2_14899 ( P2_R1209_U260 , P2_U3445 , P2_R1209_U85 );
nand NAND2_14900 ( P2_R1209_U261 , P2_REG1_REG_19_ , P2_R1209_U84 );
nand NAND2_14901 ( P2_R1209_U262 , P2_U3445 , P2_R1209_U85 );
nand NAND2_14902 ( P2_R1209_U263 , P2_REG1_REG_19_ , P2_R1209_U84 );
nand NAND2_14903 ( P2_R1209_U264 , P2_R1209_U263 , P2_R1209_U262 );
nand NAND2_14904 ( P2_R1209_U265 , P2_U3503 , P2_R1209_U63 );
nand NAND2_14905 ( P2_R1209_U266 , P2_REG1_REG_18_ , P2_R1209_U64 );
nand NAND2_14906 ( P2_R1209_U267 , P2_U3503 , P2_R1209_U63 );
nand NAND2_14907 ( P2_R1209_U268 , P2_REG1_REG_18_ , P2_R1209_U64 );
nand NAND2_14908 ( P2_R1209_U269 , P2_R1209_U268 , P2_R1209_U267 );
nand NAND3_14909 ( P2_R1209_U270 , P2_R1209_U266 , P2_R1209_U265 , P2_R1209_U65 );
nand NAND2_14910 ( P2_R1209_U271 , P2_R1209_U269 , P2_R1209_U188 );
nand NAND2_14911 ( P2_R1209_U272 , P2_U3500 , P2_R1209_U48 );
nand NAND2_14912 ( P2_R1209_U273 , P2_REG1_REG_17_ , P2_R1209_U46 );
nand NAND2_14913 ( P2_R1209_U274 , P2_U3497 , P2_R1209_U44 );
nand NAND2_14914 ( P2_R1209_U275 , P2_REG1_REG_16_ , P2_R1209_U45 );
nand NAND2_14915 ( P2_R1209_U276 , P2_R1209_U275 , P2_R1209_U274 );
nand NAND2_14916 ( P2_R1209_U277 , P2_R1209_U224 , P2_R1209_U66 );
nand NAND2_14917 ( P2_R1209_U278 , P2_R1209_U276 , P2_R1209_U180 );
nand NAND2_14918 ( P2_R1209_U279 , P2_U3494 , P2_R1209_U61 );
nand NAND2_14919 ( P2_R1209_U280 , P2_REG1_REG_15_ , P2_R1209_U62 );
nand NAND2_14920 ( P2_R1209_U281 , P2_U3494 , P2_R1209_U61 );
nand NAND2_14921 ( P2_R1209_U282 , P2_REG1_REG_15_ , P2_R1209_U62 );
nand NAND2_14922 ( P2_R1209_U283 , P2_R1209_U282 , P2_R1209_U281 );
nand NAND3_14923 ( P2_R1209_U284 , P2_R1209_U280 , P2_R1209_U279 , P2_R1209_U86 );
nand NAND2_14924 ( P2_R1209_U285 , P2_R1209_U176 , P2_R1209_U283 );
nand NAND2_14925 ( P2_R1209_U286 , P2_U3491 , P2_R1209_U59 );
nand NAND2_14926 ( P2_R1209_U287 , P2_REG1_REG_14_ , P2_R1209_U60 );
nand NAND2_14927 ( P2_R1209_U288 , P2_U3491 , P2_R1209_U59 );
nand NAND2_14928 ( P2_R1209_U289 , P2_REG1_REG_14_ , P2_R1209_U60 );
nand NAND2_14929 ( P2_R1209_U290 , P2_R1209_U289 , P2_R1209_U288 );
nand NAND3_14930 ( P2_R1209_U291 , P2_R1209_U287 , P2_R1209_U286 , P2_R1209_U87 );
nand NAND2_14931 ( P2_R1209_U292 , P2_R1209_U172 , P2_R1209_U290 );
nand NAND2_14932 ( P2_R1209_U293 , P2_U3488 , P2_R1209_U57 );
nand NAND2_14933 ( P2_R1209_U294 , P2_REG1_REG_13_ , P2_R1209_U58 );
nand NAND2_14934 ( P2_R1209_U295 , P2_U3485 , P2_R1209_U52 );
nand NAND2_14935 ( P2_R1209_U296 , P2_REG1_REG_12_ , P2_R1209_U53 );
nand NAND2_14936 ( P2_R1209_U297 , P2_R1209_U296 , P2_R1209_U295 );
nand NAND2_14937 ( P2_R1209_U298 , P2_R1209_U225 , P2_R1209_U67 );
nand NAND2_14938 ( P2_R1209_U299 , P2_R1209_U297 , P2_R1209_U205 );
nand NAND2_14939 ( P2_R1209_U300 , P2_U3482 , P2_R1209_U54 );
nand NAND2_14940 ( P2_R1209_U301 , P2_REG1_REG_11_ , P2_R1209_U55 );
nand NAND2_14941 ( P2_R1209_U302 , P2_R1209_U301 , P2_R1209_U300 );
nand NAND2_14942 ( P2_R1209_U303 , P2_R1209_U226 , P2_R1209_U88 );
nand NAND2_14943 ( P2_R1209_U304 , P2_R1209_U162 , P2_R1209_U302 );
nand NAND2_14944 ( P2_R1209_U305 , P2_U3479 , P2_R1209_U50 );
nand NAND2_14945 ( P2_R1209_U306 , P2_REG1_REG_10_ , P2_R1209_U51 );
nand NAND2_14946 ( P2_R1209_U307 , P2_U3446 , P2_R1209_U27 );
nand NAND2_14947 ( P2_R1209_U308 , P2_REG1_REG_0_ , P2_R1209_U28 );
and AND2_14948 ( P2_R1170_U4 , P2_R1170_U95 , P2_R1170_U94 );
and AND2_14949 ( P2_R1170_U5 , P2_R1170_U96 , P2_R1170_U97 );
and AND2_14950 ( P2_R1170_U6 , P2_R1170_U113 , P2_R1170_U112 );
and AND2_14951 ( P2_R1170_U7 , P2_R1170_U155 , P2_R1170_U154 );
and AND2_14952 ( P2_R1170_U8 , P2_R1170_U164 , P2_R1170_U163 );
and AND2_14953 ( P2_R1170_U9 , P2_R1170_U182 , P2_R1170_U181 );
and AND2_14954 ( P2_R1170_U10 , P2_R1170_U218 , P2_R1170_U215 );
and AND2_14955 ( P2_R1170_U11 , P2_R1170_U211 , P2_R1170_U208 );
and AND2_14956 ( P2_R1170_U12 , P2_R1170_U202 , P2_R1170_U199 );
and AND2_14957 ( P2_R1170_U13 , P2_R1170_U196 , P2_R1170_U192 );
and AND2_14958 ( P2_R1170_U14 , P2_R1170_U151 , P2_R1170_U148 );
and AND2_14959 ( P2_R1170_U15 , P2_R1170_U143 , P2_R1170_U140 );
and AND2_14960 ( P2_R1170_U16 , P2_R1170_U129 , P2_R1170_U126 );
not NOT1_14961 ( P2_R1170_U17 , P2_REG2_REG_6_ );
not NOT1_14962 ( P2_R1170_U18 , P2_U3467 );
not NOT1_14963 ( P2_R1170_U19 , P2_U3470 );
nand NAND2_14964 ( P2_R1170_U20 , P2_U3467 , P2_REG2_REG_6_ );
not NOT1_14965 ( P2_R1170_U21 , P2_REG2_REG_7_ );
not NOT1_14966 ( P2_R1170_U22 , P2_REG2_REG_4_ );
not NOT1_14967 ( P2_R1170_U23 , P2_U3461 );
not NOT1_14968 ( P2_R1170_U24 , P2_U3464 );
not NOT1_14969 ( P2_R1170_U25 , P2_REG2_REG_2_ );
not NOT1_14970 ( P2_R1170_U26 , P2_U3455 );
not NOT1_14971 ( P2_R1170_U27 , P2_REG2_REG_0_ );
not NOT1_14972 ( P2_R1170_U28 , P2_U3446 );
nand NAND2_14973 ( P2_R1170_U29 , P2_U3446 , P2_REG2_REG_0_ );
not NOT1_14974 ( P2_R1170_U30 , P2_REG2_REG_3_ );
not NOT1_14975 ( P2_R1170_U31 , P2_U3458 );
nand NAND2_14976 ( P2_R1170_U32 , P2_U3461 , P2_REG2_REG_4_ );
not NOT1_14977 ( P2_R1170_U33 , P2_REG2_REG_5_ );
not NOT1_14978 ( P2_R1170_U34 , P2_REG2_REG_8_ );
not NOT1_14979 ( P2_R1170_U35 , P2_U3473 );
not NOT1_14980 ( P2_R1170_U36 , P2_U3476 );
not NOT1_14981 ( P2_R1170_U37 , P2_REG2_REG_9_ );
nand NAND2_14982 ( P2_R1170_U38 , P2_R1170_U49 , P2_R1170_U121 );
nand NAND3_14983 ( P2_R1170_U39 , P2_R1170_U110 , P2_R1170_U108 , P2_R1170_U109 );
nand NAND2_14984 ( P2_R1170_U40 , P2_R1170_U98 , P2_R1170_U99 );
nand NAND2_14985 ( P2_R1170_U41 , P2_REG2_REG_1_ , P2_U3452 );
nand NAND3_14986 ( P2_R1170_U42 , P2_R1170_U136 , P2_R1170_U134 , P2_R1170_U135 );
nand NAND2_14987 ( P2_R1170_U43 , P2_R1170_U132 , P2_R1170_U131 );
not NOT1_14988 ( P2_R1170_U44 , P2_REG2_REG_16_ );
not NOT1_14989 ( P2_R1170_U45 , P2_U3497 );
not NOT1_14990 ( P2_R1170_U46 , P2_U3500 );
nand NAND2_14991 ( P2_R1170_U47 , P2_U3497 , P2_REG2_REG_16_ );
not NOT1_14992 ( P2_R1170_U48 , P2_REG2_REG_17_ );
nand NAND2_14993 ( P2_R1170_U49 , P2_U3473 , P2_REG2_REG_8_ );
not NOT1_14994 ( P2_R1170_U50 , P2_REG2_REG_10_ );
not NOT1_14995 ( P2_R1170_U51 , P2_U3479 );
not NOT1_14996 ( P2_R1170_U52 , P2_REG2_REG_12_ );
not NOT1_14997 ( P2_R1170_U53 , P2_U3485 );
not NOT1_14998 ( P2_R1170_U54 , P2_REG2_REG_11_ );
not NOT1_14999 ( P2_R1170_U55 , P2_U3482 );
nand NAND2_15000 ( P2_R1170_U56 , P2_U3482 , P2_REG2_REG_11_ );
not NOT1_15001 ( P2_R1170_U57 , P2_REG2_REG_13_ );
not NOT1_15002 ( P2_R1170_U58 , P2_U3488 );
not NOT1_15003 ( P2_R1170_U59 , P2_REG2_REG_14_ );
not NOT1_15004 ( P2_R1170_U60 , P2_U3491 );
not NOT1_15005 ( P2_R1170_U61 , P2_REG2_REG_15_ );
not NOT1_15006 ( P2_R1170_U62 , P2_U3494 );
not NOT1_15007 ( P2_R1170_U63 , P2_REG2_REG_18_ );
not NOT1_15008 ( P2_R1170_U64 , P2_U3503 );
nand NAND3_15009 ( P2_R1170_U65 , P2_R1170_U186 , P2_R1170_U185 , P2_R1170_U187 );
nand NAND2_15010 ( P2_R1170_U66 , P2_R1170_U179 , P2_R1170_U178 );
nand NAND2_15011 ( P2_R1170_U67 , P2_R1170_U56 , P2_R1170_U204 );
nand NAND2_15012 ( P2_R1170_U68 , P2_R1170_U259 , P2_R1170_U258 );
nand NAND2_15013 ( P2_R1170_U69 , P2_R1170_U308 , P2_R1170_U307 );
nand NAND2_15014 ( P2_R1170_U70 , P2_R1170_U231 , P2_R1170_U230 );
nand NAND2_15015 ( P2_R1170_U71 , P2_R1170_U236 , P2_R1170_U235 );
nand NAND2_15016 ( P2_R1170_U72 , P2_R1170_U243 , P2_R1170_U242 );
nand NAND2_15017 ( P2_R1170_U73 , P2_R1170_U250 , P2_R1170_U249 );
nand NAND2_15018 ( P2_R1170_U74 , P2_R1170_U255 , P2_R1170_U254 );
nand NAND2_15019 ( P2_R1170_U75 , P2_R1170_U271 , P2_R1170_U270 );
nand NAND2_15020 ( P2_R1170_U76 , P2_R1170_U278 , P2_R1170_U277 );
nand NAND2_15021 ( P2_R1170_U77 , P2_R1170_U285 , P2_R1170_U284 );
nand NAND2_15022 ( P2_R1170_U78 , P2_R1170_U292 , P2_R1170_U291 );
nand NAND2_15023 ( P2_R1170_U79 , P2_R1170_U299 , P2_R1170_U298 );
nand NAND2_15024 ( P2_R1170_U80 , P2_R1170_U304 , P2_R1170_U303 );
nand NAND3_15025 ( P2_R1170_U81 , P2_R1170_U117 , P2_R1170_U116 , P2_R1170_U118 );
nand NAND2_15026 ( P2_R1170_U82 , P2_R1170_U133 , P2_R1170_U145 );
nand NAND2_15027 ( P2_R1170_U83 , P2_R1170_U41 , P2_R1170_U152 );
not NOT1_15028 ( P2_R1170_U84 , P2_U3445 );
not NOT1_15029 ( P2_R1170_U85 , P2_REG2_REG_19_ );
nand NAND2_15030 ( P2_R1170_U86 , P2_R1170_U175 , P2_R1170_U174 );
nand NAND2_15031 ( P2_R1170_U87 , P2_R1170_U171 , P2_R1170_U170 );
nand NAND2_15032 ( P2_R1170_U88 , P2_R1170_U161 , P2_R1170_U160 );
not NOT1_15033 ( P2_R1170_U89 , P2_R1170_U32 );
nand NAND2_15034 ( P2_R1170_U90 , P2_REG2_REG_9_ , P2_U3476 );
nand NAND2_15035 ( P2_R1170_U91 , P2_U3485 , P2_REG2_REG_12_ );
not NOT1_15036 ( P2_R1170_U92 , P2_R1170_U56 );
not NOT1_15037 ( P2_R1170_U93 , P2_R1170_U49 );
or OR2_15038 ( P2_R1170_U94 , P2_U3464 , P2_REG2_REG_5_ );
or OR2_15039 ( P2_R1170_U95 , P2_U3461 , P2_REG2_REG_4_ );
or OR2_15040 ( P2_R1170_U96 , P2_REG2_REG_3_ , P2_U3458 );
or OR2_15041 ( P2_R1170_U97 , P2_REG2_REG_2_ , P2_U3455 );
not NOT1_15042 ( P2_R1170_U98 , P2_R1170_U29 );
or OR2_15043 ( P2_R1170_U99 , P2_REG2_REG_1_ , P2_U3452 );
not NOT1_15044 ( P2_R1170_U100 , P2_R1170_U40 );
not NOT1_15045 ( P2_R1170_U101 , P2_R1170_U41 );
nand NAND2_15046 ( P2_R1170_U102 , P2_R1170_U40 , P2_R1170_U41 );
nand NAND3_15047 ( P2_R1170_U103 , P2_REG2_REG_2_ , P2_U3455 , P2_R1170_U96 );
nand NAND2_15048 ( P2_R1170_U104 , P2_R1170_U5 , P2_R1170_U102 );
nand NAND2_15049 ( P2_R1170_U105 , P2_U3458 , P2_REG2_REG_3_ );
nand NAND3_15050 ( P2_R1170_U106 , P2_R1170_U105 , P2_R1170_U103 , P2_R1170_U104 );
nand NAND2_15051 ( P2_R1170_U107 , P2_R1170_U33 , P2_R1170_U32 );
nand NAND2_15052 ( P2_R1170_U108 , P2_U3464 , P2_R1170_U107 );
nand NAND2_15053 ( P2_R1170_U109 , P2_R1170_U4 , P2_R1170_U106 );
nand NAND2_15054 ( P2_R1170_U110 , P2_REG2_REG_5_ , P2_R1170_U89 );
not NOT1_15055 ( P2_R1170_U111 , P2_R1170_U39 );
or OR2_15056 ( P2_R1170_U112 , P2_U3470 , P2_REG2_REG_7_ );
or OR2_15057 ( P2_R1170_U113 , P2_U3467 , P2_REG2_REG_6_ );
not NOT1_15058 ( P2_R1170_U114 , P2_R1170_U20 );
nand NAND2_15059 ( P2_R1170_U115 , P2_R1170_U21 , P2_R1170_U20 );
nand NAND2_15060 ( P2_R1170_U116 , P2_U3470 , P2_R1170_U115 );
nand NAND2_15061 ( P2_R1170_U117 , P2_REG2_REG_7_ , P2_R1170_U114 );
nand NAND2_15062 ( P2_R1170_U118 , P2_R1170_U6 , P2_R1170_U39 );
not NOT1_15063 ( P2_R1170_U119 , P2_R1170_U81 );
or OR2_15064 ( P2_R1170_U120 , P2_REG2_REG_8_ , P2_U3473 );
nand NAND2_15065 ( P2_R1170_U121 , P2_R1170_U120 , P2_R1170_U81 );
not NOT1_15066 ( P2_R1170_U122 , P2_R1170_U38 );
or OR2_15067 ( P2_R1170_U123 , P2_U3476 , P2_REG2_REG_9_ );
or OR2_15068 ( P2_R1170_U124 , P2_REG2_REG_6_ , P2_U3467 );
nand NAND2_15069 ( P2_R1170_U125 , P2_R1170_U124 , P2_R1170_U39 );
nand NAND4_15070 ( P2_R1170_U126 , P2_R1170_U238 , P2_R1170_U237 , P2_R1170_U20 , P2_R1170_U125 );
nand NAND2_15071 ( P2_R1170_U127 , P2_R1170_U111 , P2_R1170_U20 );
nand NAND2_15072 ( P2_R1170_U128 , P2_REG2_REG_7_ , P2_U3470 );
nand NAND3_15073 ( P2_R1170_U129 , P2_R1170_U128 , P2_R1170_U6 , P2_R1170_U127 );
or OR2_15074 ( P2_R1170_U130 , P2_U3467 , P2_REG2_REG_6_ );
nand NAND2_15075 ( P2_R1170_U131 , P2_R1170_U101 , P2_R1170_U97 );
nand NAND2_15076 ( P2_R1170_U132 , P2_U3455 , P2_REG2_REG_2_ );
not NOT1_15077 ( P2_R1170_U133 , P2_R1170_U43 );
nand NAND2_15078 ( P2_R1170_U134 , P2_R1170_U100 , P2_R1170_U5 );
nand NAND2_15079 ( P2_R1170_U135 , P2_R1170_U43 , P2_R1170_U96 );
nand NAND2_15080 ( P2_R1170_U136 , P2_U3458 , P2_REG2_REG_3_ );
not NOT1_15081 ( P2_R1170_U137 , P2_R1170_U42 );
or OR2_15082 ( P2_R1170_U138 , P2_REG2_REG_4_ , P2_U3461 );
nand NAND2_15083 ( P2_R1170_U139 , P2_R1170_U138 , P2_R1170_U42 );
nand NAND4_15084 ( P2_R1170_U140 , P2_R1170_U245 , P2_R1170_U244 , P2_R1170_U32 , P2_R1170_U139 );
nand NAND2_15085 ( P2_R1170_U141 , P2_R1170_U137 , P2_R1170_U32 );
nand NAND2_15086 ( P2_R1170_U142 , P2_REG2_REG_5_ , P2_U3464 );
nand NAND3_15087 ( P2_R1170_U143 , P2_R1170_U142 , P2_R1170_U4 , P2_R1170_U141 );
or OR2_15088 ( P2_R1170_U144 , P2_U3461 , P2_REG2_REG_4_ );
nand NAND2_15089 ( P2_R1170_U145 , P2_R1170_U100 , P2_R1170_U97 );
not NOT1_15090 ( P2_R1170_U146 , P2_R1170_U82 );
nand NAND2_15091 ( P2_R1170_U147 , P2_U3458 , P2_REG2_REG_3_ );
nand NAND4_15092 ( P2_R1170_U148 , P2_R1170_U257 , P2_R1170_U256 , P2_R1170_U41 , P2_R1170_U40 );
nand NAND2_15093 ( P2_R1170_U149 , P2_R1170_U41 , P2_R1170_U40 );
nand NAND2_15094 ( P2_R1170_U150 , P2_U3455 , P2_REG2_REG_2_ );
nand NAND3_15095 ( P2_R1170_U151 , P2_R1170_U150 , P2_R1170_U97 , P2_R1170_U149 );
or OR2_15096 ( P2_R1170_U152 , P2_REG2_REG_1_ , P2_U3452 );
not NOT1_15097 ( P2_R1170_U153 , P2_R1170_U83 );
or OR2_15098 ( P2_R1170_U154 , P2_U3476 , P2_REG2_REG_9_ );
or OR2_15099 ( P2_R1170_U155 , P2_U3479 , P2_REG2_REG_10_ );
nand NAND2_15100 ( P2_R1170_U156 , P2_R1170_U93 , P2_R1170_U7 );
nand NAND2_15101 ( P2_R1170_U157 , P2_U3479 , P2_REG2_REG_10_ );
nand NAND3_15102 ( P2_R1170_U158 , P2_R1170_U157 , P2_R1170_U90 , P2_R1170_U156 );
or OR2_15103 ( P2_R1170_U159 , P2_REG2_REG_10_ , P2_U3479 );
nand NAND3_15104 ( P2_R1170_U160 , P2_R1170_U120 , P2_R1170_U7 , P2_R1170_U81 );
nand NAND2_15105 ( P2_R1170_U161 , P2_R1170_U159 , P2_R1170_U158 );
not NOT1_15106 ( P2_R1170_U162 , P2_R1170_U88 );
or OR2_15107 ( P2_R1170_U163 , P2_U3488 , P2_REG2_REG_13_ );
or OR2_15108 ( P2_R1170_U164 , P2_U3485 , P2_REG2_REG_12_ );
nand NAND2_15109 ( P2_R1170_U165 , P2_R1170_U92 , P2_R1170_U8 );
nand NAND2_15110 ( P2_R1170_U166 , P2_U3488 , P2_REG2_REG_13_ );
nand NAND3_15111 ( P2_R1170_U167 , P2_R1170_U166 , P2_R1170_U91 , P2_R1170_U165 );
or OR2_15112 ( P2_R1170_U168 , P2_REG2_REG_11_ , P2_U3482 );
or OR2_15113 ( P2_R1170_U169 , P2_REG2_REG_13_ , P2_U3488 );
nand NAND3_15114 ( P2_R1170_U170 , P2_R1170_U168 , P2_R1170_U8 , P2_R1170_U88 );
nand NAND2_15115 ( P2_R1170_U171 , P2_R1170_U169 , P2_R1170_U167 );
not NOT1_15116 ( P2_R1170_U172 , P2_R1170_U87 );
or OR2_15117 ( P2_R1170_U173 , P2_REG2_REG_14_ , P2_U3491 );
nand NAND2_15118 ( P2_R1170_U174 , P2_R1170_U173 , P2_R1170_U87 );
nand NAND2_15119 ( P2_R1170_U175 , P2_U3491 , P2_REG2_REG_14_ );
not NOT1_15120 ( P2_R1170_U176 , P2_R1170_U86 );
or OR2_15121 ( P2_R1170_U177 , P2_REG2_REG_15_ , P2_U3494 );
nand NAND2_15122 ( P2_R1170_U178 , P2_R1170_U177 , P2_R1170_U86 );
nand NAND2_15123 ( P2_R1170_U179 , P2_U3494 , P2_REG2_REG_15_ );
not NOT1_15124 ( P2_R1170_U180 , P2_R1170_U66 );
or OR2_15125 ( P2_R1170_U181 , P2_U3500 , P2_REG2_REG_17_ );
or OR2_15126 ( P2_R1170_U182 , P2_U3497 , P2_REG2_REG_16_ );
not NOT1_15127 ( P2_R1170_U183 , P2_R1170_U47 );
nand NAND2_15128 ( P2_R1170_U184 , P2_R1170_U48 , P2_R1170_U47 );
nand NAND2_15129 ( P2_R1170_U185 , P2_U3500 , P2_R1170_U184 );
nand NAND2_15130 ( P2_R1170_U186 , P2_REG2_REG_17_ , P2_R1170_U183 );
nand NAND2_15131 ( P2_R1170_U187 , P2_R1170_U9 , P2_R1170_U66 );
not NOT1_15132 ( P2_R1170_U188 , P2_R1170_U65 );
or OR2_15133 ( P2_R1170_U189 , P2_REG2_REG_18_ , P2_U3503 );
nand NAND2_15134 ( P2_R1170_U190 , P2_R1170_U189 , P2_R1170_U65 );
nand NAND2_15135 ( P2_R1170_U191 , P2_U3503 , P2_REG2_REG_18_ );
nand NAND4_15136 ( P2_R1170_U192 , P2_R1170_U261 , P2_R1170_U260 , P2_R1170_U191 , P2_R1170_U190 );
nand NAND2_15137 ( P2_R1170_U193 , P2_U3503 , P2_REG2_REG_18_ );
nand NAND2_15138 ( P2_R1170_U194 , P2_R1170_U188 , P2_R1170_U193 );
or OR2_15139 ( P2_R1170_U195 , P2_U3503 , P2_REG2_REG_18_ );
nand NAND3_15140 ( P2_R1170_U196 , P2_R1170_U195 , P2_R1170_U264 , P2_R1170_U194 );
or OR2_15141 ( P2_R1170_U197 , P2_REG2_REG_16_ , P2_U3497 );
nand NAND2_15142 ( P2_R1170_U198 , P2_R1170_U197 , P2_R1170_U66 );
nand NAND4_15143 ( P2_R1170_U199 , P2_R1170_U273 , P2_R1170_U272 , P2_R1170_U47 , P2_R1170_U198 );
nand NAND2_15144 ( P2_R1170_U200 , P2_R1170_U180 , P2_R1170_U47 );
nand NAND2_15145 ( P2_R1170_U201 , P2_REG2_REG_17_ , P2_U3500 );
nand NAND3_15146 ( P2_R1170_U202 , P2_R1170_U201 , P2_R1170_U9 , P2_R1170_U200 );
or OR2_15147 ( P2_R1170_U203 , P2_U3497 , P2_REG2_REG_16_ );
nand NAND2_15148 ( P2_R1170_U204 , P2_R1170_U168 , P2_R1170_U88 );
not NOT1_15149 ( P2_R1170_U205 , P2_R1170_U67 );
or OR2_15150 ( P2_R1170_U206 , P2_REG2_REG_12_ , P2_U3485 );
nand NAND2_15151 ( P2_R1170_U207 , P2_R1170_U206 , P2_R1170_U67 );
nand NAND4_15152 ( P2_R1170_U208 , P2_R1170_U294 , P2_R1170_U293 , P2_R1170_U91 , P2_R1170_U207 );
nand NAND2_15153 ( P2_R1170_U209 , P2_R1170_U205 , P2_R1170_U91 );
nand NAND2_15154 ( P2_R1170_U210 , P2_U3488 , P2_REG2_REG_13_ );
nand NAND3_15155 ( P2_R1170_U211 , P2_R1170_U210 , P2_R1170_U8 , P2_R1170_U209 );
or OR2_15156 ( P2_R1170_U212 , P2_U3485 , P2_REG2_REG_12_ );
or OR2_15157 ( P2_R1170_U213 , P2_REG2_REG_9_ , P2_U3476 );
nand NAND2_15158 ( P2_R1170_U214 , P2_R1170_U213 , P2_R1170_U38 );
nand NAND4_15159 ( P2_R1170_U215 , P2_R1170_U306 , P2_R1170_U305 , P2_R1170_U90 , P2_R1170_U214 );
nand NAND2_15160 ( P2_R1170_U216 , P2_R1170_U122 , P2_R1170_U90 );
nand NAND2_15161 ( P2_R1170_U217 , P2_U3479 , P2_REG2_REG_10_ );
nand NAND3_15162 ( P2_R1170_U218 , P2_R1170_U217 , P2_R1170_U7 , P2_R1170_U216 );
nand NAND2_15163 ( P2_R1170_U219 , P2_R1170_U123 , P2_R1170_U90 );
nand NAND2_15164 ( P2_R1170_U220 , P2_R1170_U120 , P2_R1170_U49 );
nand NAND2_15165 ( P2_R1170_U221 , P2_R1170_U130 , P2_R1170_U20 );
nand NAND2_15166 ( P2_R1170_U222 , P2_R1170_U144 , P2_R1170_U32 );
nand NAND2_15167 ( P2_R1170_U223 , P2_R1170_U147 , P2_R1170_U96 );
nand NAND2_15168 ( P2_R1170_U224 , P2_R1170_U203 , P2_R1170_U47 );
nand NAND2_15169 ( P2_R1170_U225 , P2_R1170_U212 , P2_R1170_U91 );
nand NAND2_15170 ( P2_R1170_U226 , P2_R1170_U168 , P2_R1170_U56 );
nand NAND2_15171 ( P2_R1170_U227 , P2_U3476 , P2_R1170_U37 );
nand NAND2_15172 ( P2_R1170_U228 , P2_REG2_REG_9_ , P2_R1170_U36 );
nand NAND2_15173 ( P2_R1170_U229 , P2_R1170_U228 , P2_R1170_U227 );
nand NAND2_15174 ( P2_R1170_U230 , P2_R1170_U219 , P2_R1170_U38 );
nand NAND2_15175 ( P2_R1170_U231 , P2_R1170_U229 , P2_R1170_U122 );
nand NAND2_15176 ( P2_R1170_U232 , P2_U3473 , P2_R1170_U34 );
nand NAND2_15177 ( P2_R1170_U233 , P2_REG2_REG_8_ , P2_R1170_U35 );
nand NAND2_15178 ( P2_R1170_U234 , P2_R1170_U233 , P2_R1170_U232 );
nand NAND2_15179 ( P2_R1170_U235 , P2_R1170_U220 , P2_R1170_U81 );
nand NAND2_15180 ( P2_R1170_U236 , P2_R1170_U119 , P2_R1170_U234 );
nand NAND2_15181 ( P2_R1170_U237 , P2_U3470 , P2_R1170_U21 );
nand NAND2_15182 ( P2_R1170_U238 , P2_REG2_REG_7_ , P2_R1170_U19 );
nand NAND2_15183 ( P2_R1170_U239 , P2_U3467 , P2_R1170_U17 );
nand NAND2_15184 ( P2_R1170_U240 , P2_REG2_REG_6_ , P2_R1170_U18 );
nand NAND2_15185 ( P2_R1170_U241 , P2_R1170_U240 , P2_R1170_U239 );
nand NAND2_15186 ( P2_R1170_U242 , P2_R1170_U221 , P2_R1170_U39 );
nand NAND2_15187 ( P2_R1170_U243 , P2_R1170_U241 , P2_R1170_U111 );
nand NAND2_15188 ( P2_R1170_U244 , P2_U3464 , P2_R1170_U33 );
nand NAND2_15189 ( P2_R1170_U245 , P2_REG2_REG_5_ , P2_R1170_U24 );
nand NAND2_15190 ( P2_R1170_U246 , P2_U3461 , P2_R1170_U22 );
nand NAND2_15191 ( P2_R1170_U247 , P2_REG2_REG_4_ , P2_R1170_U23 );
nand NAND2_15192 ( P2_R1170_U248 , P2_R1170_U247 , P2_R1170_U246 );
nand NAND2_15193 ( P2_R1170_U249 , P2_R1170_U222 , P2_R1170_U42 );
nand NAND2_15194 ( P2_R1170_U250 , P2_R1170_U248 , P2_R1170_U137 );
nand NAND2_15195 ( P2_R1170_U251 , P2_U3458 , P2_R1170_U30 );
nand NAND2_15196 ( P2_R1170_U252 , P2_REG2_REG_3_ , P2_R1170_U31 );
nand NAND2_15197 ( P2_R1170_U253 , P2_R1170_U252 , P2_R1170_U251 );
nand NAND2_15198 ( P2_R1170_U254 , P2_R1170_U223 , P2_R1170_U82 );
nand NAND2_15199 ( P2_R1170_U255 , P2_R1170_U146 , P2_R1170_U253 );
nand NAND2_15200 ( P2_R1170_U256 , P2_U3455 , P2_R1170_U25 );
nand NAND2_15201 ( P2_R1170_U257 , P2_REG2_REG_2_ , P2_R1170_U26 );
nand NAND2_15202 ( P2_R1170_U258 , P2_R1170_U98 , P2_R1170_U83 );
nand NAND2_15203 ( P2_R1170_U259 , P2_R1170_U153 , P2_R1170_U29 );
nand NAND2_15204 ( P2_R1170_U260 , P2_U3445 , P2_R1170_U85 );
nand NAND2_15205 ( P2_R1170_U261 , P2_REG2_REG_19_ , P2_R1170_U84 );
nand NAND2_15206 ( P2_R1170_U262 , P2_U3445 , P2_R1170_U85 );
nand NAND2_15207 ( P2_R1170_U263 , P2_REG2_REG_19_ , P2_R1170_U84 );
nand NAND2_15208 ( P2_R1170_U264 , P2_R1170_U263 , P2_R1170_U262 );
nand NAND2_15209 ( P2_R1170_U265 , P2_U3503 , P2_R1170_U63 );
nand NAND2_15210 ( P2_R1170_U266 , P2_REG2_REG_18_ , P2_R1170_U64 );
nand NAND2_15211 ( P2_R1170_U267 , P2_U3503 , P2_R1170_U63 );
nand NAND2_15212 ( P2_R1170_U268 , P2_REG2_REG_18_ , P2_R1170_U64 );
nand NAND2_15213 ( P2_R1170_U269 , P2_R1170_U268 , P2_R1170_U267 );
nand NAND3_15214 ( P2_R1170_U270 , P2_R1170_U266 , P2_R1170_U265 , P2_R1170_U65 );
nand NAND2_15215 ( P2_R1170_U271 , P2_R1170_U269 , P2_R1170_U188 );
nand NAND2_15216 ( P2_R1170_U272 , P2_U3500 , P2_R1170_U48 );
nand NAND2_15217 ( P2_R1170_U273 , P2_REG2_REG_17_ , P2_R1170_U46 );
nand NAND2_15218 ( P2_R1170_U274 , P2_U3497 , P2_R1170_U44 );
nand NAND2_15219 ( P2_R1170_U275 , P2_REG2_REG_16_ , P2_R1170_U45 );
nand NAND2_15220 ( P2_R1170_U276 , P2_R1170_U275 , P2_R1170_U274 );
nand NAND2_15221 ( P2_R1170_U277 , P2_R1170_U224 , P2_R1170_U66 );
nand NAND2_15222 ( P2_R1170_U278 , P2_R1170_U276 , P2_R1170_U180 );
nand NAND2_15223 ( P2_R1170_U279 , P2_U3494 , P2_R1170_U61 );
nand NAND2_15224 ( P2_R1170_U280 , P2_REG2_REG_15_ , P2_R1170_U62 );
nand NAND2_15225 ( P2_R1170_U281 , P2_U3494 , P2_R1170_U61 );
nand NAND2_15226 ( P2_R1170_U282 , P2_REG2_REG_15_ , P2_R1170_U62 );
nand NAND2_15227 ( P2_R1170_U283 , P2_R1170_U282 , P2_R1170_U281 );
nand NAND3_15228 ( P2_R1170_U284 , P2_R1170_U280 , P2_R1170_U279 , P2_R1170_U86 );
nand NAND2_15229 ( P2_R1170_U285 , P2_R1170_U176 , P2_R1170_U283 );
nand NAND2_15230 ( P2_R1170_U286 , P2_U3491 , P2_R1170_U59 );
nand NAND2_15231 ( P2_R1170_U287 , P2_REG2_REG_14_ , P2_R1170_U60 );
nand NAND2_15232 ( P2_R1170_U288 , P2_U3491 , P2_R1170_U59 );
nand NAND2_15233 ( P2_R1170_U289 , P2_REG2_REG_14_ , P2_R1170_U60 );
nand NAND2_15234 ( P2_R1170_U290 , P2_R1170_U289 , P2_R1170_U288 );
nand NAND3_15235 ( P2_R1170_U291 , P2_R1170_U287 , P2_R1170_U286 , P2_R1170_U87 );
nand NAND2_15236 ( P2_R1170_U292 , P2_R1170_U172 , P2_R1170_U290 );
nand NAND2_15237 ( P2_R1170_U293 , P2_U3488 , P2_R1170_U57 );
nand NAND2_15238 ( P2_R1170_U294 , P2_REG2_REG_13_ , P2_R1170_U58 );
nand NAND2_15239 ( P2_R1170_U295 , P2_U3485 , P2_R1170_U52 );
nand NAND2_15240 ( P2_R1170_U296 , P2_REG2_REG_12_ , P2_R1170_U53 );
nand NAND2_15241 ( P2_R1170_U297 , P2_R1170_U296 , P2_R1170_U295 );
nand NAND2_15242 ( P2_R1170_U298 , P2_R1170_U225 , P2_R1170_U67 );
nand NAND2_15243 ( P2_R1170_U299 , P2_R1170_U297 , P2_R1170_U205 );
nand NAND2_15244 ( P2_R1170_U300 , P2_U3482 , P2_R1170_U54 );
nand NAND2_15245 ( P2_R1170_U301 , P2_REG2_REG_11_ , P2_R1170_U55 );
nand NAND2_15246 ( P2_R1170_U302 , P2_R1170_U301 , P2_R1170_U300 );
nand NAND2_15247 ( P2_R1170_U303 , P2_R1170_U226 , P2_R1170_U88 );
nand NAND2_15248 ( P2_R1170_U304 , P2_R1170_U162 , P2_R1170_U302 );
nand NAND2_15249 ( P2_R1170_U305 , P2_U3479 , P2_R1170_U50 );
nand NAND2_15250 ( P2_R1170_U306 , P2_REG2_REG_10_ , P2_R1170_U51 );
nand NAND2_15251 ( P2_R1170_U307 , P2_U3446 , P2_R1170_U27 );
nand NAND2_15252 ( P2_R1170_U308 , P2_REG2_REG_0_ , P2_R1170_U28 );
and AND2_15253 ( P2_R1275_U6 , P2_R1275_U135 , P2_R1275_U35 );
and AND2_15254 ( P2_R1275_U7 , P2_R1275_U133 , P2_R1275_U36 );
and AND2_15255 ( P2_R1275_U8 , P2_R1275_U132 , P2_R1275_U37 );
and AND2_15256 ( P2_R1275_U9 , P2_R1275_U131 , P2_R1275_U38 );
and AND2_15257 ( P2_R1275_U10 , P2_R1275_U129 , P2_R1275_U39 );
and AND2_15258 ( P2_R1275_U11 , P2_R1275_U128 , P2_R1275_U40 );
and AND2_15259 ( P2_R1275_U12 , P2_R1275_U127 , P2_R1275_U41 );
and AND2_15260 ( P2_R1275_U13 , P2_R1275_U125 , P2_R1275_U42 );
and AND2_15261 ( P2_R1275_U14 , P2_R1275_U123 , P2_R1275_U43 );
and AND2_15262 ( P2_R1275_U15 , P2_R1275_U121 , P2_R1275_U44 );
and AND2_15263 ( P2_R1275_U16 , P2_R1275_U119 , P2_R1275_U45 );
and AND2_15264 ( P2_R1275_U17 , P2_R1275_U117 , P2_R1275_U46 );
and AND2_15265 ( P2_R1275_U18 , P2_R1275_U115 , P2_R1275_U25 );
and AND2_15266 ( P2_R1275_U19 , P2_R1275_U113 , P2_R1275_U67 );
and AND2_15267 ( P2_R1275_U20 , P2_R1275_U98 , P2_R1275_U26 );
and AND2_15268 ( P2_R1275_U21 , P2_R1275_U97 , P2_R1275_U27 );
and AND2_15269 ( P2_R1275_U22 , P2_R1275_U96 , P2_R1275_U28 );
and AND2_15270 ( P2_R1275_U23 , P2_R1275_U94 , P2_R1275_U29 );
and AND2_15271 ( P2_R1275_U24 , P2_R1275_U93 , P2_R1275_U30 );
or OR3_15272 ( P2_R1275_U25 , P2_U3453 , P2_U3448 , P2_U3456 );
nand NAND2_15273 ( P2_R1275_U26 , P2_R1275_U87 , P2_R1275_U34 );
nand NAND2_15274 ( P2_R1275_U27 , P2_R1275_U88 , P2_R1275_U33 );
nand NAND2_15275 ( P2_R1275_U28 , P2_R1275_U56 , P2_R1275_U89 );
nand NAND2_15276 ( P2_R1275_U29 , P2_R1275_U90 , P2_R1275_U32 );
nand NAND2_15277 ( P2_R1275_U30 , P2_R1275_U91 , P2_R1275_U31 );
not NOT1_15278 ( P2_R1275_U31 , P2_U3474 );
not NOT1_15279 ( P2_R1275_U32 , P2_U3471 );
not NOT1_15280 ( P2_R1275_U33 , P2_U3462 );
not NOT1_15281 ( P2_R1275_U34 , P2_U3459 );
nand NAND2_15282 ( P2_R1275_U35 , P2_R1275_U57 , P2_R1275_U92 );
nand NAND2_15283 ( P2_R1275_U36 , P2_R1275_U99 , P2_R1275_U54 );
nand NAND2_15284 ( P2_R1275_U37 , P2_R1275_U100 , P2_R1275_U53 );
nand NAND2_15285 ( P2_R1275_U38 , P2_R1275_U58 , P2_R1275_U101 );
nand NAND2_15286 ( P2_R1275_U39 , P2_R1275_U102 , P2_R1275_U52 );
nand NAND2_15287 ( P2_R1275_U40 , P2_R1275_U103 , P2_R1275_U51 );
nand NAND2_15288 ( P2_R1275_U41 , P2_R1275_U59 , P2_R1275_U104 );
nand NAND2_15289 ( P2_R1275_U42 , P2_R1275_U60 , P2_R1275_U105 );
nand NAND2_15290 ( P2_R1275_U43 , P2_R1275_U61 , P2_R1275_U106 );
nand NAND3_15291 ( P2_R1275_U44 , P2_R1275_U107 , P2_R1275_U75 , P2_R1275_U50 );
nand NAND3_15292 ( P2_R1275_U45 , P2_R1275_U108 , P2_R1275_U73 , P2_R1275_U49 );
nand NAND3_15293 ( P2_R1275_U46 , P2_R1275_U109 , P2_R1275_U71 , P2_R1275_U48 );
not NOT1_15294 ( P2_R1275_U47 , P2_U3978 );
not NOT1_15295 ( P2_R1275_U48 , P2_U3968 );
not NOT1_15296 ( P2_R1275_U49 , P2_U3970 );
not NOT1_15297 ( P2_R1275_U50 , P2_U3972 );
not NOT1_15298 ( P2_R1275_U51 , P2_U3498 );
not NOT1_15299 ( P2_R1275_U52 , P2_U3495 );
not NOT1_15300 ( P2_R1275_U53 , P2_U3486 );
not NOT1_15301 ( P2_R1275_U54 , P2_U3483 );
nand NAND2_15302 ( P2_R1275_U55 , P2_R1275_U153 , P2_R1275_U152 );
nor nor_15303 ( P2_R1275_U56 , P2_U3465 , P2_U3468 );
nor nor_15304 ( P2_R1275_U57 , P2_U3480 , P2_U3477 );
nor nor_15305 ( P2_R1275_U58 , P2_U3489 , P2_U3492 );
nor nor_15306 ( P2_R1275_U59 , P2_U3501 , P2_U3504 );
nor nor_15307 ( P2_R1275_U60 , P2_U3506 , P2_U3976 );
nor nor_15308 ( P2_R1275_U61 , P2_U3975 , P2_U3974 );
not NOT1_15309 ( P2_R1275_U62 , P2_U3477 );
and AND2_15310 ( P2_R1275_U63 , P2_R1275_U137 , P2_R1275_U136 );
not NOT1_15311 ( P2_R1275_U64 , P2_U3465 );
and AND2_15312 ( P2_R1275_U65 , P2_R1275_U139 , P2_R1275_U138 );
not NOT1_15313 ( P2_R1275_U66 , P2_U3977 );
nand NAND3_15314 ( P2_R1275_U67 , P2_R1275_U110 , P2_R1275_U69 , P2_R1275_U47 );
and AND2_15315 ( P2_R1275_U68 , P2_R1275_U141 , P2_R1275_U140 );
not NOT1_15316 ( P2_R1275_U69 , P2_U3979 );
and AND2_15317 ( P2_R1275_U70 , P2_R1275_U143 , P2_R1275_U142 );
not NOT1_15318 ( P2_R1275_U71 , P2_U3969 );
and AND2_15319 ( P2_R1275_U72 , P2_R1275_U145 , P2_R1275_U144 );
not NOT1_15320 ( P2_R1275_U73 , P2_U3971 );
and AND2_15321 ( P2_R1275_U74 , P2_R1275_U147 , P2_R1275_U146 );
not NOT1_15322 ( P2_R1275_U75 , P2_U3973 );
and AND2_15323 ( P2_R1275_U76 , P2_R1275_U149 , P2_R1275_U148 );
not NOT1_15324 ( P2_R1275_U77 , P2_U3975 );
and AND2_15325 ( P2_R1275_U78 , P2_R1275_U151 , P2_R1275_U150 );
not NOT1_15326 ( P2_R1275_U79 , P2_U3453 );
not NOT1_15327 ( P2_R1275_U80 , P2_U3448 );
not NOT1_15328 ( P2_R1275_U81 , P2_U3506 );
and AND2_15329 ( P2_R1275_U82 , P2_R1275_U155 , P2_R1275_U154 );
not NOT1_15330 ( P2_R1275_U83 , P2_U3501 );
and AND2_15331 ( P2_R1275_U84 , P2_R1275_U157 , P2_R1275_U156 );
not NOT1_15332 ( P2_R1275_U85 , P2_U3489 );
and AND2_15333 ( P2_R1275_U86 , P2_R1275_U159 , P2_R1275_U158 );
not NOT1_15334 ( P2_R1275_U87 , P2_R1275_U25 );
not NOT1_15335 ( P2_R1275_U88 , P2_R1275_U26 );
not NOT1_15336 ( P2_R1275_U89 , P2_R1275_U27 );
not NOT1_15337 ( P2_R1275_U90 , P2_R1275_U28 );
not NOT1_15338 ( P2_R1275_U91 , P2_R1275_U29 );
not NOT1_15339 ( P2_R1275_U92 , P2_R1275_U30 );
nand NAND2_15340 ( P2_R1275_U93 , P2_U3474 , P2_R1275_U29 );
nand NAND2_15341 ( P2_R1275_U94 , P2_U3471 , P2_R1275_U28 );
nand NAND2_15342 ( P2_R1275_U95 , P2_R1275_U89 , P2_R1275_U64 );
nand NAND2_15343 ( P2_R1275_U96 , P2_U3468 , P2_R1275_U95 );
nand NAND2_15344 ( P2_R1275_U97 , P2_U3462 , P2_R1275_U26 );
nand NAND2_15345 ( P2_R1275_U98 , P2_U3459 , P2_R1275_U25 );
not NOT1_15346 ( P2_R1275_U99 , P2_R1275_U35 );
not NOT1_15347 ( P2_R1275_U100 , P2_R1275_U36 );
not NOT1_15348 ( P2_R1275_U101 , P2_R1275_U37 );
not NOT1_15349 ( P2_R1275_U102 , P2_R1275_U38 );
not NOT1_15350 ( P2_R1275_U103 , P2_R1275_U39 );
not NOT1_15351 ( P2_R1275_U104 , P2_R1275_U40 );
not NOT1_15352 ( P2_R1275_U105 , P2_R1275_U41 );
not NOT1_15353 ( P2_R1275_U106 , P2_R1275_U42 );
not NOT1_15354 ( P2_R1275_U107 , P2_R1275_U43 );
not NOT1_15355 ( P2_R1275_U108 , P2_R1275_U44 );
not NOT1_15356 ( P2_R1275_U109 , P2_R1275_U45 );
not NOT1_15357 ( P2_R1275_U110 , P2_R1275_U46 );
not NOT1_15358 ( P2_R1275_U111 , P2_R1275_U67 );
nand NAND2_15359 ( P2_R1275_U112 , P2_R1275_U110 , P2_R1275_U69 );
nand NAND2_15360 ( P2_R1275_U113 , P2_U3978 , P2_R1275_U112 );
or OR2_15361 ( P2_R1275_U114 , P2_U3453 , P2_U3448 );
nand NAND2_15362 ( P2_R1275_U115 , P2_U3456 , P2_R1275_U114 );
nand NAND2_15363 ( P2_R1275_U116 , P2_R1275_U109 , P2_R1275_U71 );
nand NAND2_15364 ( P2_R1275_U117 , P2_U3968 , P2_R1275_U116 );
nand NAND2_15365 ( P2_R1275_U118 , P2_R1275_U108 , P2_R1275_U73 );
nand NAND2_15366 ( P2_R1275_U119 , P2_U3970 , P2_R1275_U118 );
nand NAND2_15367 ( P2_R1275_U120 , P2_R1275_U107 , P2_R1275_U75 );
nand NAND2_15368 ( P2_R1275_U121 , P2_U3972 , P2_R1275_U120 );
nand NAND2_15369 ( P2_R1275_U122 , P2_R1275_U106 , P2_R1275_U77 );
nand NAND2_15370 ( P2_R1275_U123 , P2_U3974 , P2_R1275_U122 );
nand NAND2_15371 ( P2_R1275_U124 , P2_R1275_U105 , P2_R1275_U81 );
nand NAND2_15372 ( P2_R1275_U125 , P2_U3976 , P2_R1275_U124 );
nand NAND2_15373 ( P2_R1275_U126 , P2_R1275_U104 , P2_R1275_U83 );
nand NAND2_15374 ( P2_R1275_U127 , P2_U3504 , P2_R1275_U126 );
nand NAND2_15375 ( P2_R1275_U128 , P2_U3498 , P2_R1275_U39 );
nand NAND2_15376 ( P2_R1275_U129 , P2_U3495 , P2_R1275_U38 );
nand NAND2_15377 ( P2_R1275_U130 , P2_R1275_U101 , P2_R1275_U85 );
nand NAND2_15378 ( P2_R1275_U131 , P2_U3492 , P2_R1275_U130 );
nand NAND2_15379 ( P2_R1275_U132 , P2_U3486 , P2_R1275_U36 );
nand NAND2_15380 ( P2_R1275_U133 , P2_U3483 , P2_R1275_U35 );
nand NAND2_15381 ( P2_R1275_U134 , P2_R1275_U92 , P2_R1275_U62 );
nand NAND2_15382 ( P2_R1275_U135 , P2_U3480 , P2_R1275_U134 );
nand NAND2_15383 ( P2_R1275_U136 , P2_U3477 , P2_R1275_U30 );
nand NAND2_15384 ( P2_R1275_U137 , P2_R1275_U92 , P2_R1275_U62 );
nand NAND2_15385 ( P2_R1275_U138 , P2_U3465 , P2_R1275_U27 );
nand NAND2_15386 ( P2_R1275_U139 , P2_R1275_U89 , P2_R1275_U64 );
nand NAND2_15387 ( P2_R1275_U140 , P2_U3977 , P2_R1275_U67 );
nand NAND2_15388 ( P2_R1275_U141 , P2_R1275_U111 , P2_R1275_U66 );
nand NAND2_15389 ( P2_R1275_U142 , P2_U3979 , P2_R1275_U46 );
nand NAND2_15390 ( P2_R1275_U143 , P2_R1275_U110 , P2_R1275_U69 );
nand NAND2_15391 ( P2_R1275_U144 , P2_U3969 , P2_R1275_U45 );
nand NAND2_15392 ( P2_R1275_U145 , P2_R1275_U109 , P2_R1275_U71 );
nand NAND2_15393 ( P2_R1275_U146 , P2_U3971 , P2_R1275_U44 );
nand NAND2_15394 ( P2_R1275_U147 , P2_R1275_U108 , P2_R1275_U73 );
nand NAND2_15395 ( P2_R1275_U148 , P2_U3973 , P2_R1275_U43 );
nand NAND2_15396 ( P2_R1275_U149 , P2_R1275_U107 , P2_R1275_U75 );
nand NAND2_15397 ( P2_R1275_U150 , P2_U3975 , P2_R1275_U42 );
nand NAND2_15398 ( P2_R1275_U151 , P2_R1275_U106 , P2_R1275_U77 );
nand NAND2_15399 ( P2_R1275_U152 , P2_U3453 , P2_R1275_U80 );
nand NAND2_15400 ( P2_R1275_U153 , P2_U3448 , P2_R1275_U79 );
nand NAND2_15401 ( P2_R1275_U154 , P2_U3506 , P2_R1275_U41 );
nand NAND2_15402 ( P2_R1275_U155 , P2_R1275_U105 , P2_R1275_U81 );
nand NAND2_15403 ( P2_R1275_U156 , P2_U3501 , P2_R1275_U40 );
nand NAND2_15404 ( P2_R1275_U157 , P2_R1275_U104 , P2_R1275_U83 );
nand NAND2_15405 ( P2_R1275_U158 , P2_U3489 , P2_R1275_U37 );
nand NAND2_15406 ( P2_R1275_U159 , P2_R1275_U101 , P2_R1275_U85 );
and AND2_15407 ( P2_LT_719_U6 , P2_LT_719_U115 , P2_LT_719_U116 );
and AND4_15408 ( P2_LT_719_U7 , P2_LT_719_U122 , P2_LT_719_U121 , P2_LT_719_U120 , P2_LT_719_U118 );
and AND2_15409 ( P2_LT_719_U8 , P2_LT_719_U75 , P2_LT_719_U7 );
and AND2_15410 ( P2_LT_719_U9 , P2_LT_719_U8 , P2_LT_719_U126 );
and AND3_15411 ( P2_LT_719_U10 , P2_LT_719_U111 , P2_LT_719_U112 , P2_LT_719_U109 );
and AND4_15412 ( P2_LT_719_U11 , P2_LT_719_U186 , P2_LT_719_U185 , P2_LT_719_U105 , P2_LT_719_U106 );
not NOT1_15413 ( P2_LT_719_U12 , P2_U3979 );
not NOT1_15414 ( P2_LT_719_U13 , P2_U3592 );
not NOT1_15415 ( P2_LT_719_U14 , P2_U3599 );
not NOT1_15416 ( P2_LT_719_U15 , P2_U3600 );
not NOT1_15417 ( P2_LT_719_U16 , P2_U3974 );
not NOT1_15418 ( P2_LT_719_U17 , P2_U3606 );
not NOT1_15419 ( P2_LT_719_U18 , P2_U3605 );
not NOT1_15420 ( P2_LT_719_U19 , P2_U3498 );
not NOT1_15421 ( P2_LT_719_U20 , P2_U3495 );
not NOT1_15422 ( P2_LT_719_U21 , P2_U3492 );
not NOT1_15423 ( P2_LT_719_U22 , P2_U3611 );
not NOT1_15424 ( P2_LT_719_U23 , P2_U3480 );
not NOT1_15425 ( P2_LT_719_U24 , P2_U3477 );
not NOT1_15426 ( P2_LT_719_U25 , P2_U3471 );
not NOT1_15427 ( P2_LT_719_U26 , P2_U3474 );
not NOT1_15428 ( P2_LT_719_U27 , P2_U3468 );
not NOT1_15429 ( P2_LT_719_U28 , P2_U3465 );
not NOT1_15430 ( P2_LT_719_U29 , P2_U3462 );
not NOT1_15431 ( P2_LT_719_U30 , P2_U3459 );
not NOT1_15432 ( P2_LT_719_U31 , P2_U3604 );
not NOT1_15433 ( P2_LT_719_U32 , P2_U3456 );
not NOT1_15434 ( P2_LT_719_U33 , P2_U3453 );
not NOT1_15435 ( P2_LT_719_U34 , P2_U3612 );
not NOT1_15436 ( P2_LT_719_U35 , P2_U3593 );
not NOT1_15437 ( P2_LT_719_U36 , P2_U3590 );
not NOT1_15438 ( P2_LT_719_U37 , P2_U3589 );
not NOT1_15439 ( P2_LT_719_U38 , P2_U3588 );
not NOT1_15440 ( P2_LT_719_U39 , P2_U3587 );
not NOT1_15441 ( P2_LT_719_U40 , P2_U3586 );
not NOT1_15442 ( P2_LT_719_U41 , P2_U3585 );
not NOT1_15443 ( P2_LT_719_U42 , P2_U3584 );
not NOT1_15444 ( P2_LT_719_U43 , P2_U3614 );
not NOT1_15445 ( P2_LT_719_U44 , P2_U3613 );
not NOT1_15446 ( P2_LT_719_U45 , P2_U3486 );
not NOT1_15447 ( P2_LT_719_U46 , P2_U3483 );
not NOT1_15448 ( P2_LT_719_U47 , P2_U3489 );
not NOT1_15449 ( P2_LT_719_U48 , P2_U3610 );
not NOT1_15450 ( P2_LT_719_U49 , P2_U3609 );
not NOT1_15451 ( P2_LT_719_U50 , P2_U3608 );
not NOT1_15452 ( P2_LT_719_U51 , P2_U3607 );
not NOT1_15453 ( P2_LT_719_U52 , P2_U3975 );
not NOT1_15454 ( P2_LT_719_U53 , P2_U3504 );
not NOT1_15455 ( P2_LT_719_U54 , P2_U3501 );
not NOT1_15456 ( P2_LT_719_U55 , P2_U3506 );
not NOT1_15457 ( P2_LT_719_U56 , P2_U3976 );
not NOT1_15458 ( P2_LT_719_U57 , P2_U3603 );
not NOT1_15459 ( P2_LT_719_U58 , P2_U3602 );
not NOT1_15460 ( P2_LT_719_U59 , P2_U3601 );
not NOT1_15461 ( P2_LT_719_U60 , P2_U3973 );
not NOT1_15462 ( P2_LT_719_U61 , P2_U3972 );
nand NAND2_15463 ( P2_LT_719_U62 , P2_LT_719_U179 , P2_LT_719_U178 );
not NOT1_15464 ( P2_LT_719_U63 , P2_U3598 );
not NOT1_15465 ( P2_LT_719_U64 , P2_U3970 );
not NOT1_15466 ( P2_LT_719_U65 , P2_U3591 );
not NOT1_15467 ( P2_LT_719_U66 , P2_U3969 );
not NOT1_15468 ( P2_LT_719_U67 , P2_U3968 );
not NOT1_15469 ( P2_LT_719_U68 , P2_U3978 );
not NOT1_15470 ( P2_LT_719_U69 , P2_U3594 );
not NOT1_15471 ( P2_LT_719_U70 , P2_U3596 );
not NOT1_15472 ( P2_LT_719_U71 , P2_U3597 );
not NOT1_15473 ( P2_LT_719_U72 , P2_U3977 );
not NOT1_15474 ( P2_LT_719_U73 , P2_U3595 );
and AND2_15475 ( P2_LT_719_U74 , P2_U3448 , P2_LT_719_U107 );
and AND3_15476 ( P2_LT_719_U75 , P2_LT_719_U124 , P2_LT_719_U123 , P2_LT_719_U125 );
and AND2_15477 ( P2_LT_719_U76 , P2_LT_719_U128 , P2_LT_719_U129 );
and AND2_15478 ( P2_LT_719_U77 , P2_LT_719_U76 , P2_LT_719_U127 );
and AND2_15479 ( P2_LT_719_U78 , P2_U3593 , P2_LT_719_U32 );
and AND2_15480 ( P2_LT_719_U79 , P2_U3590 , P2_LT_719_U30 );
and AND2_15481 ( P2_LT_719_U80 , P2_LT_719_U124 , P2_LT_719_U123 );
and AND2_15482 ( P2_LT_719_U81 , P2_LT_719_U140 , P2_LT_719_U141 );
and AND2_15483 ( P2_LT_719_U82 , P2_LT_719_U120 , P2_LT_719_U118 );
and AND2_15484 ( P2_LT_719_U83 , P2_LT_719_U146 , P2_LT_719_U84 );
and AND2_15485 ( P2_LT_719_U84 , P2_LT_719_U148 , P2_LT_719_U147 );
and AND2_15486 ( P2_LT_719_U85 , P2_LT_719_U145 , P2_LT_719_U83 );
and AND2_15487 ( P2_LT_719_U86 , P2_U3483 , P2_LT_719_U44 );
and AND2_15488 ( P2_LT_719_U87 , P2_LT_719_U151 , P2_LT_719_U88 );
and AND2_15489 ( P2_LT_719_U88 , P2_LT_719_U152 , P2_LT_719_U150 );
and AND2_15490 ( P2_LT_719_U89 , P2_LT_719_U155 , P2_LT_719_U132 );
and AND2_15491 ( P2_LT_719_U90 , P2_LT_719_U153 , P2_LT_719_U117 );
and AND2_15492 ( P2_LT_719_U91 , P2_LT_719_U6 , P2_LT_719_U92 );
and AND2_15493 ( P2_LT_719_U92 , P2_LT_719_U161 , P2_LT_719_U162 );
and AND2_15494 ( P2_LT_719_U93 , P2_U3504 , P2_LT_719_U17 );
and AND2_15495 ( P2_LT_719_U94 , P2_U3501 , P2_LT_719_U51 );
and AND2_15496 ( P2_LT_719_U95 , P2_LT_719_U164 , P2_LT_719_U166 );
and AND4_15497 ( P2_LT_719_U96 , P2_LT_719_U168 , P2_LT_719_U167 , P2_LT_719_U169 , P2_LT_719_U95 );
and AND2_15498 ( P2_LT_719_U97 , P2_U3603 , P2_LT_719_U56 );
and AND3_15499 ( P2_LT_719_U98 , P2_LT_719_U171 , P2_LT_719_U172 , P2_LT_719_U173 );
and AND2_15500 ( P2_LT_719_U99 , P2_LT_719_U176 , P2_LT_719_U165 );
and AND2_15501 ( P2_LT_719_U100 , P2_LT_719_U174 , P2_LT_719_U113 );
and AND2_15502 ( P2_LT_719_U101 , P2_LT_719_U10 , P2_LT_719_U184 );
and AND2_15503 ( P2_LT_719_U102 , P2_U3594 , P2_LT_719_U12 );
and AND2_15504 ( P2_LT_719_U103 , P2_LT_719_U104 , P2_LT_719_U109 );
and AND2_15505 ( P2_LT_719_U104 , P2_U3595 , P2_LT_719_U67 );
and AND2_15506 ( P2_LT_719_U105 , P2_LT_719_U189 , P2_LT_719_U188 );
and AND3_15507 ( P2_LT_719_U106 , P2_LT_719_U191 , P2_LT_719_U192 , P2_LT_719_U190 );
not NOT1_15508 ( P2_LT_719_U107 , P2_U3615 );
nand NAND2_15509 ( P2_LT_719_U108 , P2_LT_719_U194 , P2_LT_719_U193 );
nand NAND2_15510 ( P2_LT_719_U109 , P2_U3591 , P2_LT_719_U72 );
nand NAND2_15511 ( P2_LT_719_U110 , P2_U3979 , P2_LT_719_U69 );
nand NAND2_15512 ( P2_LT_719_U111 , P2_U3969 , P2_LT_719_U70 );
nand NAND2_15513 ( P2_LT_719_U112 , P2_U3968 , P2_LT_719_U73 );
nand NAND2_15514 ( P2_LT_719_U113 , P2_U3599 , P2_LT_719_U61 );
nand NAND2_15515 ( P2_LT_719_U114 , P2_U3498 , P2_LT_719_U50 );
nand NAND2_15516 ( P2_LT_719_U115 , P2_U3605 , P2_LT_719_U55 );
nand NAND2_15517 ( P2_LT_719_U116 , P2_U3606 , P2_LT_719_U53 );
nand NAND2_15518 ( P2_LT_719_U117 , P2_U3495 , P2_LT_719_U49 );
nand NAND2_15519 ( P2_LT_719_U118 , P2_U3480 , P2_LT_719_U43 );
nand NAND2_15520 ( P2_LT_719_U119 , P2_U3604 , P2_LT_719_U33 );
nand NAND2_15521 ( P2_LT_719_U120 , P2_U3477 , P2_LT_719_U42 );
nand NAND2_15522 ( P2_LT_719_U121 , P2_U3471 , P2_LT_719_U40 );
nand NAND2_15523 ( P2_LT_719_U122 , P2_U3474 , P2_LT_719_U41 );
nand NAND2_15524 ( P2_LT_719_U123 , P2_U3468 , P2_LT_719_U39 );
nand NAND2_15525 ( P2_LT_719_U124 , P2_U3465 , P2_LT_719_U38 );
nand NAND2_15526 ( P2_LT_719_U125 , P2_U3462 , P2_LT_719_U37 );
nand NAND2_15527 ( P2_LT_719_U126 , P2_U3459 , P2_LT_719_U36 );
nand NAND2_15528 ( P2_LT_719_U127 , P2_LT_719_U74 , P2_LT_719_U119 );
nand NAND2_15529 ( P2_LT_719_U128 , P2_U3456 , P2_LT_719_U35 );
nand NAND2_15530 ( P2_LT_719_U129 , P2_U3453 , P2_LT_719_U31 );
nand NAND2_15531 ( P2_LT_719_U130 , P2_LT_719_U77 , P2_LT_719_U9 );
nand NAND2_15532 ( P2_LT_719_U131 , P2_U3612 , P2_LT_719_U45 );
nand NAND2_15533 ( P2_LT_719_U132 , P2_U3611 , P2_LT_719_U47 );
nand NAND2_15534 ( P2_LT_719_U133 , P2_U3585 , P2_LT_719_U26 );
nand NAND2_15535 ( P2_LT_719_U134 , P2_U3584 , P2_LT_719_U24 );
nand NAND2_15536 ( P2_LT_719_U135 , P2_LT_719_U134 , P2_LT_719_U133 );
nand NAND2_15537 ( P2_LT_719_U136 , P2_U3589 , P2_LT_719_U29 );
nand NAND2_15538 ( P2_LT_719_U137 , P2_U3588 , P2_LT_719_U28 );
nand NAND2_15539 ( P2_LT_719_U138 , P2_LT_719_U137 , P2_LT_719_U136 );
nand NAND2_15540 ( P2_LT_719_U139 , P2_LT_719_U80 , P2_LT_719_U138 );
nand NAND2_15541 ( P2_LT_719_U140 , P2_U3587 , P2_LT_719_U27 );
nand NAND2_15542 ( P2_LT_719_U141 , P2_U3586 , P2_LT_719_U25 );
nand NAND2_15543 ( P2_LT_719_U142 , P2_LT_719_U81 , P2_LT_719_U139 );
nand NAND2_15544 ( P2_LT_719_U143 , P2_LT_719_U78 , P2_LT_719_U9 );
nand NAND2_15545 ( P2_LT_719_U144 , P2_LT_719_U79 , P2_LT_719_U8 );
nand NAND2_15546 ( P2_LT_719_U145 , P2_LT_719_U7 , P2_LT_719_U142 );
nand NAND2_15547 ( P2_LT_719_U146 , P2_LT_719_U82 , P2_LT_719_U135 );
nand NAND2_15548 ( P2_LT_719_U147 , P2_U3614 , P2_LT_719_U23 );
nand NAND2_15549 ( P2_LT_719_U148 , P2_U3613 , P2_LT_719_U46 );
nand NAND5_15550 ( P2_LT_719_U149 , P2_LT_719_U144 , P2_LT_719_U143 , P2_LT_719_U131 , P2_LT_719_U130 , P2_LT_719_U85 );
nand NAND2_15551 ( P2_LT_719_U150 , P2_U3486 , P2_LT_719_U34 );
nand NAND2_15552 ( P2_LT_719_U151 , P2_LT_719_U86 , P2_LT_719_U131 );
nand NAND2_15553 ( P2_LT_719_U152 , P2_U3489 , P2_LT_719_U22 );
nand NAND2_15554 ( P2_LT_719_U153 , P2_U3492 , P2_LT_719_U48 );
nand NAND2_15555 ( P2_LT_719_U154 , P2_LT_719_U149 , P2_LT_719_U87 );
nand NAND2_15556 ( P2_LT_719_U155 , P2_U3610 , P2_LT_719_U21 );
nand NAND2_15557 ( P2_LT_719_U156 , P2_LT_719_U89 , P2_LT_719_U154 );
nand NAND2_15558 ( P2_LT_719_U157 , P2_LT_719_U90 , P2_LT_719_U156 );
nand NAND2_15559 ( P2_LT_719_U158 , P2_U3609 , P2_LT_719_U20 );
nand NAND2_15560 ( P2_LT_719_U159 , P2_LT_719_U158 , P2_LT_719_U157 );
nand NAND2_15561 ( P2_LT_719_U160 , P2_LT_719_U159 , P2_LT_719_U114 );
nand NAND2_15562 ( P2_LT_719_U161 , P2_U3608 , P2_LT_719_U19 );
nand NAND2_15563 ( P2_LT_719_U162 , P2_U3607 , P2_LT_719_U54 );
nand NAND2_15564 ( P2_LT_719_U163 , P2_LT_719_U160 , P2_LT_719_U91 );
nand NAND2_15565 ( P2_LT_719_U164 , P2_U3975 , P2_LT_719_U58 );
nand NAND2_15566 ( P2_LT_719_U165 , P2_U3974 , P2_LT_719_U59 );
nand NAND2_15567 ( P2_LT_719_U166 , P2_LT_719_U93 , P2_LT_719_U115 );
nand NAND2_15568 ( P2_LT_719_U167 , P2_LT_719_U94 , P2_LT_719_U6 );
nand NAND2_15569 ( P2_LT_719_U168 , P2_U3506 , P2_LT_719_U18 );
nand NAND2_15570 ( P2_LT_719_U169 , P2_U3976 , P2_LT_719_U57 );
nand NAND2_15571 ( P2_LT_719_U170 , P2_LT_719_U163 , P2_LT_719_U96 );
nand NAND2_15572 ( P2_LT_719_U171 , P2_LT_719_U97 , P2_LT_719_U164 );
nand NAND2_15573 ( P2_LT_719_U172 , P2_U3602 , P2_LT_719_U52 );
nand NAND2_15574 ( P2_LT_719_U173 , P2_U3601 , P2_LT_719_U16 );
nand NAND2_15575 ( P2_LT_719_U174 , P2_U3600 , P2_LT_719_U60 );
nand NAND2_15576 ( P2_LT_719_U175 , P2_LT_719_U170 , P2_LT_719_U98 );
nand NAND2_15577 ( P2_LT_719_U176 , P2_U3973 , P2_LT_719_U15 );
nand NAND2_15578 ( P2_LT_719_U177 , P2_LT_719_U99 , P2_LT_719_U175 );
nand NAND2_15579 ( P2_LT_719_U178 , P2_LT_719_U100 , P2_LT_719_U177 );
nand NAND2_15580 ( P2_LT_719_U179 , P2_U3972 , P2_LT_719_U14 );
not NOT1_15581 ( P2_LT_719_U180 , P2_LT_719_U62 );
nand NAND2_15582 ( P2_LT_719_U181 , P2_U3598 , P2_LT_719_U180 );
nand NAND2_15583 ( P2_LT_719_U182 , P2_U3971 , P2_LT_719_U181 );
nand NAND2_15584 ( P2_LT_719_U183 , P2_LT_719_U62 , P2_LT_719_U63 );
nand NAND2_15585 ( P2_LT_719_U184 , P2_U3970 , P2_LT_719_U71 );
nand NAND4_15586 ( P2_LT_719_U185 , P2_LT_719_U182 , P2_LT_719_U183 , P2_LT_719_U108 , P2_LT_719_U101 );
nand NAND3_15587 ( P2_LT_719_U186 , P2_LT_719_U109 , P2_U3592 , P2_LT_719_U68 );
nand NAND2_15588 ( P2_LT_719_U187 , P2_U3978 , P2_LT_719_U13 );
nand NAND3_15589 ( P2_LT_719_U188 , P2_LT_719_U109 , P2_LT_719_U102 , P2_LT_719_U187 );
nand NAND4_15590 ( P2_LT_719_U189 , P2_U3596 , P2_LT_719_U10 , P2_LT_719_U108 , P2_LT_719_U66 );
nand NAND4_15591 ( P2_LT_719_U190 , P2_U3597 , P2_LT_719_U10 , P2_LT_719_U108 , P2_LT_719_U64 );
nand NAND2_15592 ( P2_LT_719_U191 , P2_U3977 , P2_LT_719_U65 );
nand NAND2_15593 ( P2_LT_719_U192 , P2_LT_719_U108 , P2_LT_719_U103 );
nand NAND2_15594 ( P2_LT_719_U193 , P2_U3592 , P2_LT_719_U110 );
nand NAND2_15595 ( P2_LT_719_U194 , P2_LT_719_U110 , P2_LT_719_U68 );
and AND2_15596 ( P2_R1179_U6 , P2_R1179_U205 , P2_R1179_U204 );
and AND2_15597 ( P2_R1179_U7 , P2_R1179_U244 , P2_R1179_U243 );
and AND2_15598 ( P2_R1179_U8 , P2_R1179_U261 , P2_R1179_U260 );
and AND2_15599 ( P2_R1179_U9 , P2_R1179_U285 , P2_R1179_U284 );
and AND2_15600 ( P2_R1179_U10 , P2_R1179_U384 , P2_R1179_U383 );
nand NAND2_15601 ( P2_R1179_U11 , P2_R1179_U340 , P2_R1179_U343 );
nand NAND2_15602 ( P2_R1179_U12 , P2_R1179_U329 , P2_R1179_U332 );
nand NAND2_15603 ( P2_R1179_U13 , P2_R1179_U318 , P2_R1179_U321 );
nand NAND2_15604 ( P2_R1179_U14 , P2_R1179_U310 , P2_R1179_U312 );
nand NAND3_15605 ( P2_R1179_U15 , P2_R1179_U349 , P2_R1179_U177 , P2_R1179_U156 );
nand NAND2_15606 ( P2_R1179_U16 , P2_R1179_U238 , P2_R1179_U240 );
nand NAND2_15607 ( P2_R1179_U17 , P2_R1179_U230 , P2_R1179_U233 );
nand NAND2_15608 ( P2_R1179_U18 , P2_R1179_U222 , P2_R1179_U224 );
nand NAND2_15609 ( P2_R1179_U19 , P2_R1179_U166 , P2_R1179_U346 );
not NOT1_15610 ( P2_R1179_U20 , P2_U3471 );
not NOT1_15611 ( P2_R1179_U21 , P2_U3465 );
not NOT1_15612 ( P2_R1179_U22 , P2_U3456 );
not NOT1_15613 ( P2_R1179_U23 , P2_U3448 );
not NOT1_15614 ( P2_R1179_U24 , P2_U3078 );
not NOT1_15615 ( P2_R1179_U25 , P2_U3459 );
not NOT1_15616 ( P2_R1179_U26 , P2_U3068 );
nand NAND2_15617 ( P2_R1179_U27 , P2_U3068 , P2_R1179_U22 );
not NOT1_15618 ( P2_R1179_U28 , P2_U3064 );
not NOT1_15619 ( P2_R1179_U29 , P2_U3468 );
not NOT1_15620 ( P2_R1179_U30 , P2_U3462 );
not NOT1_15621 ( P2_R1179_U31 , P2_U3071 );
not NOT1_15622 ( P2_R1179_U32 , P2_U3067 );
not NOT1_15623 ( P2_R1179_U33 , P2_U3060 );
nand NAND2_15624 ( P2_R1179_U34 , P2_U3060 , P2_R1179_U30 );
not NOT1_15625 ( P2_R1179_U35 , P2_U3474 );
not NOT1_15626 ( P2_R1179_U36 , P2_U3070 );
nand NAND2_15627 ( P2_R1179_U37 , P2_U3070 , P2_R1179_U20 );
not NOT1_15628 ( P2_R1179_U38 , P2_U3084 );
not NOT1_15629 ( P2_R1179_U39 , P2_U3477 );
not NOT1_15630 ( P2_R1179_U40 , P2_U3083 );
nand NAND2_15631 ( P2_R1179_U41 , P2_R1179_U211 , P2_R1179_U210 );
nand NAND2_15632 ( P2_R1179_U42 , P2_R1179_U34 , P2_R1179_U226 );
nand NAND3_15633 ( P2_R1179_U43 , P2_R1179_U195 , P2_R1179_U179 , P2_R1179_U347 );
not NOT1_15634 ( P2_R1179_U44 , P2_U3970 );
not NOT1_15635 ( P2_R1179_U45 , P2_U3974 );
not NOT1_15636 ( P2_R1179_U46 , P2_U3495 );
not NOT1_15637 ( P2_R1179_U47 , P2_U3480 );
not NOT1_15638 ( P2_R1179_U48 , P2_U3483 );
not NOT1_15639 ( P2_R1179_U49 , P2_U3063 );
not NOT1_15640 ( P2_R1179_U50 , P2_U3062 );
nand NAND2_15641 ( P2_R1179_U51 , P2_U3083 , P2_R1179_U39 );
not NOT1_15642 ( P2_R1179_U52 , P2_U3486 );
not NOT1_15643 ( P2_R1179_U53 , P2_U3072 );
not NOT1_15644 ( P2_R1179_U54 , P2_U3489 );
not NOT1_15645 ( P2_R1179_U55 , P2_U3080 );
not NOT1_15646 ( P2_R1179_U56 , P2_U3498 );
not NOT1_15647 ( P2_R1179_U57 , P2_U3492 );
not NOT1_15648 ( P2_R1179_U58 , P2_U3073 );
not NOT1_15649 ( P2_R1179_U59 , P2_U3074 );
not NOT1_15650 ( P2_R1179_U60 , P2_U3079 );
nand NAND2_15651 ( P2_R1179_U61 , P2_U3079 , P2_R1179_U57 );
not NOT1_15652 ( P2_R1179_U62 , P2_U3501 );
not NOT1_15653 ( P2_R1179_U63 , P2_U3069 );
not NOT1_15654 ( P2_R1179_U64 , P2_U3082 );
not NOT1_15655 ( P2_R1179_U65 , P2_U3506 );
not NOT1_15656 ( P2_R1179_U66 , P2_U3081 );
not NOT1_15657 ( P2_R1179_U67 , P2_U3976 );
not NOT1_15658 ( P2_R1179_U68 , P2_U3076 );
not NOT1_15659 ( P2_R1179_U69 , P2_U3973 );
not NOT1_15660 ( P2_R1179_U70 , P2_U3975 );
not NOT1_15661 ( P2_R1179_U71 , P2_U3066 );
not NOT1_15662 ( P2_R1179_U72 , P2_U3061 );
not NOT1_15663 ( P2_R1179_U73 , P2_U3075 );
nand NAND2_15664 ( P2_R1179_U74 , P2_U3075 , P2_R1179_U70 );
not NOT1_15665 ( P2_R1179_U75 , P2_U3972 );
not NOT1_15666 ( P2_R1179_U76 , P2_U3065 );
not NOT1_15667 ( P2_R1179_U77 , P2_U3971 );
not NOT1_15668 ( P2_R1179_U78 , P2_U3058 );
not NOT1_15669 ( P2_R1179_U79 , P2_U3969 );
not NOT1_15670 ( P2_R1179_U80 , P2_U3057 );
nand NAND2_15671 ( P2_R1179_U81 , P2_U3057 , P2_R1179_U44 );
not NOT1_15672 ( P2_R1179_U82 , P2_U3053 );
not NOT1_15673 ( P2_R1179_U83 , P2_U3968 );
not NOT1_15674 ( P2_R1179_U84 , P2_U3054 );
nand NAND2_15675 ( P2_R1179_U85 , P2_R1179_U299 , P2_R1179_U298 );
nand NAND2_15676 ( P2_R1179_U86 , P2_R1179_U74 , P2_R1179_U314 );
nand NAND2_15677 ( P2_R1179_U87 , P2_R1179_U61 , P2_R1179_U325 );
nand NAND2_15678 ( P2_R1179_U88 , P2_R1179_U51 , P2_R1179_U336 );
not NOT1_15679 ( P2_R1179_U89 , P2_U3077 );
nand NAND2_15680 ( P2_R1179_U90 , P2_R1179_U394 , P2_R1179_U393 );
nand NAND2_15681 ( P2_R1179_U91 , P2_R1179_U408 , P2_R1179_U407 );
nand NAND2_15682 ( P2_R1179_U92 , P2_R1179_U413 , P2_R1179_U412 );
nand NAND2_15683 ( P2_R1179_U93 , P2_R1179_U429 , P2_R1179_U428 );
nand NAND2_15684 ( P2_R1179_U94 , P2_R1179_U434 , P2_R1179_U433 );
nand NAND2_15685 ( P2_R1179_U95 , P2_R1179_U439 , P2_R1179_U438 );
nand NAND2_15686 ( P2_R1179_U96 , P2_R1179_U444 , P2_R1179_U443 );
nand NAND2_15687 ( P2_R1179_U97 , P2_R1179_U449 , P2_R1179_U448 );
nand NAND2_15688 ( P2_R1179_U98 , P2_R1179_U465 , P2_R1179_U464 );
nand NAND2_15689 ( P2_R1179_U99 , P2_R1179_U470 , P2_R1179_U469 );
nand NAND2_15690 ( P2_R1179_U100 , P2_R1179_U353 , P2_R1179_U352 );
nand NAND2_15691 ( P2_R1179_U101 , P2_R1179_U362 , P2_R1179_U361 );
nand NAND2_15692 ( P2_R1179_U102 , P2_R1179_U369 , P2_R1179_U368 );
nand NAND2_15693 ( P2_R1179_U103 , P2_R1179_U373 , P2_R1179_U372 );
nand NAND2_15694 ( P2_R1179_U104 , P2_R1179_U382 , P2_R1179_U381 );
nand NAND2_15695 ( P2_R1179_U105 , P2_R1179_U403 , P2_R1179_U402 );
nand NAND2_15696 ( P2_R1179_U106 , P2_R1179_U420 , P2_R1179_U419 );
nand NAND2_15697 ( P2_R1179_U107 , P2_R1179_U424 , P2_R1179_U423 );
nand NAND2_15698 ( P2_R1179_U108 , P2_R1179_U456 , P2_R1179_U455 );
nand NAND2_15699 ( P2_R1179_U109 , P2_R1179_U460 , P2_R1179_U459 );
nand NAND2_15700 ( P2_R1179_U110 , P2_R1179_U477 , P2_R1179_U476 );
and AND2_15701 ( P2_R1179_U111 , P2_R1179_U197 , P2_R1179_U187 );
and AND2_15702 ( P2_R1179_U112 , P2_R1179_U200 , P2_R1179_U201 );
and AND3_15703 ( P2_R1179_U113 , P2_R1179_U208 , P2_R1179_U203 , P2_R1179_U188 );
and AND2_15704 ( P2_R1179_U114 , P2_R1179_U213 , P2_R1179_U189 );
and AND2_15705 ( P2_R1179_U115 , P2_R1179_U216 , P2_R1179_U217 );
and AND3_15706 ( P2_R1179_U116 , P2_R1179_U355 , P2_R1179_U354 , P2_R1179_U37 );
and AND2_15707 ( P2_R1179_U117 , P2_R1179_U358 , P2_R1179_U189 );
and AND2_15708 ( P2_R1179_U118 , P2_R1179_U232 , P2_R1179_U6 );
and AND2_15709 ( P2_R1179_U119 , P2_R1179_U365 , P2_R1179_U188 );
and AND3_15710 ( P2_R1179_U120 , P2_R1179_U375 , P2_R1179_U374 , P2_R1179_U27 );
and AND2_15711 ( P2_R1179_U121 , P2_R1179_U378 , P2_R1179_U187 );
and AND3_15712 ( P2_R1179_U122 , P2_R1179_U242 , P2_R1179_U219 , P2_R1179_U183 );
and AND3_15713 ( P2_R1179_U123 , P2_R1179_U264 , P2_R1179_U184 , P2_R1179_U259 );
and AND3_15714 ( P2_R1179_U124 , P2_R1179_U288 , P2_R1179_U185 , P2_R1179_U283 );
and AND2_15715 ( P2_R1179_U125 , P2_R1179_U301 , P2_R1179_U186 );
and AND2_15716 ( P2_R1179_U126 , P2_R1179_U304 , P2_R1179_U305 );
and AND2_15717 ( P2_R1179_U127 , P2_R1179_U304 , P2_R1179_U305 );
and AND2_15718 ( P2_R1179_U128 , P2_R1179_U10 , P2_R1179_U308 );
nand NAND2_15719 ( P2_R1179_U129 , P2_R1179_U391 , P2_R1179_U390 );
and AND3_15720 ( P2_R1179_U130 , P2_R1179_U396 , P2_R1179_U395 , P2_R1179_U81 );
and AND2_15721 ( P2_R1179_U131 , P2_R1179_U399 , P2_R1179_U186 );
nand NAND2_15722 ( P2_R1179_U132 , P2_R1179_U405 , P2_R1179_U404 );
nand NAND2_15723 ( P2_R1179_U133 , P2_R1179_U410 , P2_R1179_U409 );
and AND2_15724 ( P2_R1179_U134 , P2_R1179_U320 , P2_R1179_U9 );
and AND2_15725 ( P2_R1179_U135 , P2_R1179_U416 , P2_R1179_U185 );
nand NAND2_15726 ( P2_R1179_U136 , P2_R1179_U426 , P2_R1179_U425 );
nand NAND2_15727 ( P2_R1179_U137 , P2_R1179_U431 , P2_R1179_U430 );
nand NAND2_15728 ( P2_R1179_U138 , P2_R1179_U436 , P2_R1179_U435 );
nand NAND2_15729 ( P2_R1179_U139 , P2_R1179_U441 , P2_R1179_U440 );
nand NAND2_15730 ( P2_R1179_U140 , P2_R1179_U446 , P2_R1179_U445 );
and AND2_15731 ( P2_R1179_U141 , P2_R1179_U331 , P2_R1179_U8 );
and AND2_15732 ( P2_R1179_U142 , P2_R1179_U452 , P2_R1179_U184 );
nand NAND2_15733 ( P2_R1179_U143 , P2_R1179_U462 , P2_R1179_U461 );
nand NAND2_15734 ( P2_R1179_U144 , P2_R1179_U467 , P2_R1179_U466 );
and AND2_15735 ( P2_R1179_U145 , P2_R1179_U342 , P2_R1179_U7 );
and AND2_15736 ( P2_R1179_U146 , P2_R1179_U473 , P2_R1179_U183 );
and AND2_15737 ( P2_R1179_U147 , P2_R1179_U351 , P2_R1179_U350 );
nand NAND2_15738 ( P2_R1179_U148 , P2_R1179_U115 , P2_R1179_U214 );
and AND2_15739 ( P2_R1179_U149 , P2_R1179_U360 , P2_R1179_U359 );
and AND2_15740 ( P2_R1179_U150 , P2_R1179_U367 , P2_R1179_U366 );
and AND2_15741 ( P2_R1179_U151 , P2_R1179_U371 , P2_R1179_U370 );
nand NAND2_15742 ( P2_R1179_U152 , P2_R1179_U112 , P2_R1179_U198 );
and AND2_15743 ( P2_R1179_U153 , P2_R1179_U380 , P2_R1179_U379 );
not NOT1_15744 ( P2_R1179_U154 , P2_U3979 );
not NOT1_15745 ( P2_R1179_U155 , P2_U3055 );
and AND2_15746 ( P2_R1179_U156 , P2_R1179_U389 , P2_R1179_U388 );
nand NAND2_15747 ( P2_R1179_U157 , P2_R1179_U126 , P2_R1179_U302 );
and AND2_15748 ( P2_R1179_U158 , P2_R1179_U401 , P2_R1179_U400 );
nand NAND2_15749 ( P2_R1179_U159 , P2_R1179_U295 , P2_R1179_U294 );
nand NAND2_15750 ( P2_R1179_U160 , P2_R1179_U291 , P2_R1179_U290 );
and AND2_15751 ( P2_R1179_U161 , P2_R1179_U418 , P2_R1179_U417 );
and AND2_15752 ( P2_R1179_U162 , P2_R1179_U422 , P2_R1179_U421 );
nand NAND2_15753 ( P2_R1179_U163 , P2_R1179_U281 , P2_R1179_U280 );
nand NAND2_15754 ( P2_R1179_U164 , P2_R1179_U277 , P2_R1179_U276 );
not NOT1_15755 ( P2_R1179_U165 , P2_U3453 );
nand NAND2_15756 ( P2_R1179_U166 , P2_U3448 , P2_R1179_U89 );
nand NAND3_15757 ( P2_R1179_U167 , P2_R1179_U273 , P2_R1179_U178 , P2_R1179_U348 );
not NOT1_15758 ( P2_R1179_U168 , P2_U3504 );
nand NAND2_15759 ( P2_R1179_U169 , P2_R1179_U271 , P2_R1179_U270 );
nand NAND2_15760 ( P2_R1179_U170 , P2_R1179_U267 , P2_R1179_U266 );
and AND2_15761 ( P2_R1179_U171 , P2_R1179_U454 , P2_R1179_U453 );
and AND2_15762 ( P2_R1179_U172 , P2_R1179_U458 , P2_R1179_U457 );
nand NAND2_15763 ( P2_R1179_U173 , P2_R1179_U257 , P2_R1179_U256 );
nand NAND2_15764 ( P2_R1179_U174 , P2_R1179_U253 , P2_R1179_U252 );
nand NAND2_15765 ( P2_R1179_U175 , P2_R1179_U249 , P2_R1179_U248 );
and AND2_15766 ( P2_R1179_U176 , P2_R1179_U475 , P2_R1179_U474 );
nand NAND3_15767 ( P2_R1179_U177 , P2_R1179_U307 , P2_R1179_U157 , P2_R1179_U387 );
nand NAND2_15768 ( P2_R1179_U178 , P2_R1179_U169 , P2_R1179_U168 );
nand NAND2_15769 ( P2_R1179_U179 , P2_R1179_U166 , P2_R1179_U165 );
not NOT1_15770 ( P2_R1179_U180 , P2_R1179_U81 );
not NOT1_15771 ( P2_R1179_U181 , P2_R1179_U27 );
not NOT1_15772 ( P2_R1179_U182 , P2_R1179_U37 );
nand NAND2_15773 ( P2_R1179_U183 , P2_U3480 , P2_R1179_U50 );
nand NAND2_15774 ( P2_R1179_U184 , P2_U3495 , P2_R1179_U59 );
nand NAND2_15775 ( P2_R1179_U185 , P2_U3974 , P2_R1179_U72 );
nand NAND2_15776 ( P2_R1179_U186 , P2_U3970 , P2_R1179_U80 );
nand NAND2_15777 ( P2_R1179_U187 , P2_U3456 , P2_R1179_U26 );
nand NAND2_15778 ( P2_R1179_U188 , P2_U3465 , P2_R1179_U32 );
nand NAND2_15779 ( P2_R1179_U189 , P2_U3471 , P2_R1179_U36 );
not NOT1_15780 ( P2_R1179_U190 , P2_R1179_U61 );
not NOT1_15781 ( P2_R1179_U191 , P2_R1179_U74 );
not NOT1_15782 ( P2_R1179_U192 , P2_R1179_U34 );
not NOT1_15783 ( P2_R1179_U193 , P2_R1179_U51 );
not NOT1_15784 ( P2_R1179_U194 , P2_R1179_U166 );
nand NAND2_15785 ( P2_R1179_U195 , P2_U3078 , P2_R1179_U166 );
not NOT1_15786 ( P2_R1179_U196 , P2_R1179_U43 );
nand NAND2_15787 ( P2_R1179_U197 , P2_U3459 , P2_R1179_U28 );
nand NAND2_15788 ( P2_R1179_U198 , P2_R1179_U111 , P2_R1179_U43 );
nand NAND2_15789 ( P2_R1179_U199 , P2_R1179_U28 , P2_R1179_U27 );
nand NAND2_15790 ( P2_R1179_U200 , P2_R1179_U199 , P2_R1179_U25 );
nand NAND2_15791 ( P2_R1179_U201 , P2_U3064 , P2_R1179_U181 );
not NOT1_15792 ( P2_R1179_U202 , P2_R1179_U152 );
nand NAND2_15793 ( P2_R1179_U203 , P2_U3468 , P2_R1179_U31 );
nand NAND2_15794 ( P2_R1179_U204 , P2_U3071 , P2_R1179_U29 );
nand NAND2_15795 ( P2_R1179_U205 , P2_U3067 , P2_R1179_U21 );
nand NAND2_15796 ( P2_R1179_U206 , P2_R1179_U192 , P2_R1179_U188 );
nand NAND2_15797 ( P2_R1179_U207 , P2_R1179_U6 , P2_R1179_U206 );
nand NAND2_15798 ( P2_R1179_U208 , P2_U3462 , P2_R1179_U33 );
nand NAND2_15799 ( P2_R1179_U209 , P2_U3468 , P2_R1179_U31 );
nand NAND2_15800 ( P2_R1179_U210 , P2_R1179_U152 , P2_R1179_U113 );
nand NAND2_15801 ( P2_R1179_U211 , P2_R1179_U209 , P2_R1179_U207 );
not NOT1_15802 ( P2_R1179_U212 , P2_R1179_U41 );
nand NAND2_15803 ( P2_R1179_U213 , P2_U3474 , P2_R1179_U38 );
nand NAND2_15804 ( P2_R1179_U214 , P2_R1179_U114 , P2_R1179_U41 );
nand NAND2_15805 ( P2_R1179_U215 , P2_R1179_U38 , P2_R1179_U37 );
nand NAND2_15806 ( P2_R1179_U216 , P2_R1179_U215 , P2_R1179_U35 );
nand NAND2_15807 ( P2_R1179_U217 , P2_U3084 , P2_R1179_U182 );
not NOT1_15808 ( P2_R1179_U218 , P2_R1179_U148 );
nand NAND2_15809 ( P2_R1179_U219 , P2_U3477 , P2_R1179_U40 );
nand NAND2_15810 ( P2_R1179_U220 , P2_R1179_U219 , P2_R1179_U51 );
nand NAND2_15811 ( P2_R1179_U221 , P2_R1179_U212 , P2_R1179_U37 );
nand NAND2_15812 ( P2_R1179_U222 , P2_R1179_U117 , P2_R1179_U221 );
nand NAND2_15813 ( P2_R1179_U223 , P2_R1179_U41 , P2_R1179_U189 );
nand NAND2_15814 ( P2_R1179_U224 , P2_R1179_U116 , P2_R1179_U223 );
nand NAND2_15815 ( P2_R1179_U225 , P2_R1179_U37 , P2_R1179_U189 );
nand NAND2_15816 ( P2_R1179_U226 , P2_R1179_U208 , P2_R1179_U152 );
not NOT1_15817 ( P2_R1179_U227 , P2_R1179_U42 );
nand NAND2_15818 ( P2_R1179_U228 , P2_U3067 , P2_R1179_U21 );
nand NAND2_15819 ( P2_R1179_U229 , P2_R1179_U227 , P2_R1179_U228 );
nand NAND2_15820 ( P2_R1179_U230 , P2_R1179_U119 , P2_R1179_U229 );
nand NAND2_15821 ( P2_R1179_U231 , P2_R1179_U42 , P2_R1179_U188 );
nand NAND2_15822 ( P2_R1179_U232 , P2_U3468 , P2_R1179_U31 );
nand NAND2_15823 ( P2_R1179_U233 , P2_R1179_U118 , P2_R1179_U231 );
nand NAND2_15824 ( P2_R1179_U234 , P2_U3067 , P2_R1179_U21 );
nand NAND2_15825 ( P2_R1179_U235 , P2_R1179_U188 , P2_R1179_U234 );
nand NAND2_15826 ( P2_R1179_U236 , P2_R1179_U208 , P2_R1179_U34 );
nand NAND2_15827 ( P2_R1179_U237 , P2_R1179_U196 , P2_R1179_U27 );
nand NAND2_15828 ( P2_R1179_U238 , P2_R1179_U121 , P2_R1179_U237 );
nand NAND2_15829 ( P2_R1179_U239 , P2_R1179_U43 , P2_R1179_U187 );
nand NAND2_15830 ( P2_R1179_U240 , P2_R1179_U120 , P2_R1179_U239 );
nand NAND2_15831 ( P2_R1179_U241 , P2_R1179_U27 , P2_R1179_U187 );
nand NAND2_15832 ( P2_R1179_U242 , P2_U3483 , P2_R1179_U49 );
nand NAND2_15833 ( P2_R1179_U243 , P2_U3063 , P2_R1179_U48 );
nand NAND2_15834 ( P2_R1179_U244 , P2_U3062 , P2_R1179_U47 );
nand NAND2_15835 ( P2_R1179_U245 , P2_R1179_U193 , P2_R1179_U183 );
nand NAND2_15836 ( P2_R1179_U246 , P2_R1179_U7 , P2_R1179_U245 );
nand NAND2_15837 ( P2_R1179_U247 , P2_U3483 , P2_R1179_U49 );
nand NAND2_15838 ( P2_R1179_U248 , P2_R1179_U148 , P2_R1179_U122 );
nand NAND2_15839 ( P2_R1179_U249 , P2_R1179_U247 , P2_R1179_U246 );
not NOT1_15840 ( P2_R1179_U250 , P2_R1179_U175 );
nand NAND2_15841 ( P2_R1179_U251 , P2_U3486 , P2_R1179_U53 );
nand NAND2_15842 ( P2_R1179_U252 , P2_R1179_U251 , P2_R1179_U175 );
nand NAND2_15843 ( P2_R1179_U253 , P2_U3072 , P2_R1179_U52 );
not NOT1_15844 ( P2_R1179_U254 , P2_R1179_U174 );
nand NAND2_15845 ( P2_R1179_U255 , P2_U3489 , P2_R1179_U55 );
nand NAND2_15846 ( P2_R1179_U256 , P2_R1179_U255 , P2_R1179_U174 );
nand NAND2_15847 ( P2_R1179_U257 , P2_U3080 , P2_R1179_U54 );
not NOT1_15848 ( P2_R1179_U258 , P2_R1179_U173 );
nand NAND2_15849 ( P2_R1179_U259 , P2_U3498 , P2_R1179_U58 );
nand NAND2_15850 ( P2_R1179_U260 , P2_U3073 , P2_R1179_U56 );
nand NAND2_15851 ( P2_R1179_U261 , P2_U3074 , P2_R1179_U46 );
nand NAND2_15852 ( P2_R1179_U262 , P2_R1179_U190 , P2_R1179_U184 );
nand NAND2_15853 ( P2_R1179_U263 , P2_R1179_U8 , P2_R1179_U262 );
nand NAND2_15854 ( P2_R1179_U264 , P2_U3492 , P2_R1179_U60 );
nand NAND2_15855 ( P2_R1179_U265 , P2_U3498 , P2_R1179_U58 );
nand NAND2_15856 ( P2_R1179_U266 , P2_R1179_U173 , P2_R1179_U123 );
nand NAND2_15857 ( P2_R1179_U267 , P2_R1179_U265 , P2_R1179_U263 );
not NOT1_15858 ( P2_R1179_U268 , P2_R1179_U170 );
nand NAND2_15859 ( P2_R1179_U269 , P2_U3501 , P2_R1179_U63 );
nand NAND2_15860 ( P2_R1179_U270 , P2_R1179_U269 , P2_R1179_U170 );
nand NAND2_15861 ( P2_R1179_U271 , P2_U3069 , P2_R1179_U62 );
not NOT1_15862 ( P2_R1179_U272 , P2_R1179_U169 );
nand NAND2_15863 ( P2_R1179_U273 , P2_U3082 , P2_R1179_U169 );
not NOT1_15864 ( P2_R1179_U274 , P2_R1179_U167 );
nand NAND2_15865 ( P2_R1179_U275 , P2_U3506 , P2_R1179_U66 );
nand NAND2_15866 ( P2_R1179_U276 , P2_R1179_U275 , P2_R1179_U167 );
nand NAND2_15867 ( P2_R1179_U277 , P2_U3081 , P2_R1179_U65 );
not NOT1_15868 ( P2_R1179_U278 , P2_R1179_U164 );
nand NAND2_15869 ( P2_R1179_U279 , P2_U3976 , P2_R1179_U68 );
nand NAND2_15870 ( P2_R1179_U280 , P2_R1179_U279 , P2_R1179_U164 );
nand NAND2_15871 ( P2_R1179_U281 , P2_U3076 , P2_R1179_U67 );
not NOT1_15872 ( P2_R1179_U282 , P2_R1179_U163 );
nand NAND2_15873 ( P2_R1179_U283 , P2_U3973 , P2_R1179_U71 );
nand NAND2_15874 ( P2_R1179_U284 , P2_U3066 , P2_R1179_U69 );
nand NAND2_15875 ( P2_R1179_U285 , P2_U3061 , P2_R1179_U45 );
nand NAND2_15876 ( P2_R1179_U286 , P2_R1179_U191 , P2_R1179_U185 );
nand NAND2_15877 ( P2_R1179_U287 , P2_R1179_U9 , P2_R1179_U286 );
nand NAND2_15878 ( P2_R1179_U288 , P2_U3975 , P2_R1179_U73 );
nand NAND2_15879 ( P2_R1179_U289 , P2_U3973 , P2_R1179_U71 );
nand NAND2_15880 ( P2_R1179_U290 , P2_R1179_U163 , P2_R1179_U124 );
nand NAND2_15881 ( P2_R1179_U291 , P2_R1179_U289 , P2_R1179_U287 );
not NOT1_15882 ( P2_R1179_U292 , P2_R1179_U160 );
nand NAND2_15883 ( P2_R1179_U293 , P2_U3972 , P2_R1179_U76 );
nand NAND2_15884 ( P2_R1179_U294 , P2_R1179_U293 , P2_R1179_U160 );
nand NAND2_15885 ( P2_R1179_U295 , P2_U3065 , P2_R1179_U75 );
not NOT1_15886 ( P2_R1179_U296 , P2_R1179_U159 );
nand NAND2_15887 ( P2_R1179_U297 , P2_U3971 , P2_R1179_U78 );
nand NAND2_15888 ( P2_R1179_U298 , P2_R1179_U297 , P2_R1179_U159 );
nand NAND2_15889 ( P2_R1179_U299 , P2_U3058 , P2_R1179_U77 );
not NOT1_15890 ( P2_R1179_U300 , P2_R1179_U85 );
nand NAND2_15891 ( P2_R1179_U301 , P2_U3969 , P2_R1179_U82 );
nand NAND2_15892 ( P2_R1179_U302 , P2_R1179_U125 , P2_R1179_U85 );
nand NAND2_15893 ( P2_R1179_U303 , P2_R1179_U82 , P2_R1179_U81 );
nand NAND2_15894 ( P2_R1179_U304 , P2_R1179_U303 , P2_R1179_U79 );
nand NAND2_15895 ( P2_R1179_U305 , P2_U3053 , P2_R1179_U180 );
not NOT1_15896 ( P2_R1179_U306 , P2_R1179_U157 );
nand NAND2_15897 ( P2_R1179_U307 , P2_U3968 , P2_R1179_U84 );
nand NAND2_15898 ( P2_R1179_U308 , P2_U3054 , P2_R1179_U83 );
nand NAND2_15899 ( P2_R1179_U309 , P2_R1179_U300 , P2_R1179_U81 );
nand NAND2_15900 ( P2_R1179_U310 , P2_R1179_U131 , P2_R1179_U309 );
nand NAND2_15901 ( P2_R1179_U311 , P2_R1179_U85 , P2_R1179_U186 );
nand NAND2_15902 ( P2_R1179_U312 , P2_R1179_U130 , P2_R1179_U311 );
nand NAND2_15903 ( P2_R1179_U313 , P2_R1179_U81 , P2_R1179_U186 );
nand NAND2_15904 ( P2_R1179_U314 , P2_R1179_U288 , P2_R1179_U163 );
not NOT1_15905 ( P2_R1179_U315 , P2_R1179_U86 );
nand NAND2_15906 ( P2_R1179_U316 , P2_U3061 , P2_R1179_U45 );
nand NAND2_15907 ( P2_R1179_U317 , P2_R1179_U315 , P2_R1179_U316 );
nand NAND2_15908 ( P2_R1179_U318 , P2_R1179_U135 , P2_R1179_U317 );
nand NAND2_15909 ( P2_R1179_U319 , P2_R1179_U86 , P2_R1179_U185 );
nand NAND2_15910 ( P2_R1179_U320 , P2_U3973 , P2_R1179_U71 );
nand NAND2_15911 ( P2_R1179_U321 , P2_R1179_U134 , P2_R1179_U319 );
nand NAND2_15912 ( P2_R1179_U322 , P2_U3061 , P2_R1179_U45 );
nand NAND2_15913 ( P2_R1179_U323 , P2_R1179_U185 , P2_R1179_U322 );
nand NAND2_15914 ( P2_R1179_U324 , P2_R1179_U288 , P2_R1179_U74 );
nand NAND2_15915 ( P2_R1179_U325 , P2_R1179_U264 , P2_R1179_U173 );
not NOT1_15916 ( P2_R1179_U326 , P2_R1179_U87 );
nand NAND2_15917 ( P2_R1179_U327 , P2_U3074 , P2_R1179_U46 );
nand NAND2_15918 ( P2_R1179_U328 , P2_R1179_U326 , P2_R1179_U327 );
nand NAND2_15919 ( P2_R1179_U329 , P2_R1179_U142 , P2_R1179_U328 );
nand NAND2_15920 ( P2_R1179_U330 , P2_R1179_U87 , P2_R1179_U184 );
nand NAND2_15921 ( P2_R1179_U331 , P2_U3498 , P2_R1179_U58 );
nand NAND2_15922 ( P2_R1179_U332 , P2_R1179_U141 , P2_R1179_U330 );
nand NAND2_15923 ( P2_R1179_U333 , P2_U3074 , P2_R1179_U46 );
nand NAND2_15924 ( P2_R1179_U334 , P2_R1179_U184 , P2_R1179_U333 );
nand NAND2_15925 ( P2_R1179_U335 , P2_R1179_U264 , P2_R1179_U61 );
nand NAND2_15926 ( P2_R1179_U336 , P2_R1179_U219 , P2_R1179_U148 );
not NOT1_15927 ( P2_R1179_U337 , P2_R1179_U88 );
nand NAND2_15928 ( P2_R1179_U338 , P2_U3062 , P2_R1179_U47 );
nand NAND2_15929 ( P2_R1179_U339 , P2_R1179_U337 , P2_R1179_U338 );
nand NAND2_15930 ( P2_R1179_U340 , P2_R1179_U146 , P2_R1179_U339 );
nand NAND2_15931 ( P2_R1179_U341 , P2_R1179_U88 , P2_R1179_U183 );
nand NAND2_15932 ( P2_R1179_U342 , P2_U3483 , P2_R1179_U49 );
nand NAND2_15933 ( P2_R1179_U343 , P2_R1179_U145 , P2_R1179_U341 );
nand NAND2_15934 ( P2_R1179_U344 , P2_U3062 , P2_R1179_U47 );
nand NAND2_15935 ( P2_R1179_U345 , P2_R1179_U183 , P2_R1179_U344 );
nand NAND2_15936 ( P2_R1179_U346 , P2_U3077 , P2_R1179_U23 );
nand NAND2_15937 ( P2_R1179_U347 , P2_U3078 , P2_R1179_U165 );
nand NAND2_15938 ( P2_R1179_U348 , P2_U3082 , P2_R1179_U168 );
nand NAND3_15939 ( P2_R1179_U349 , P2_R1179_U127 , P2_R1179_U302 , P2_R1179_U128 );
nand NAND2_15940 ( P2_R1179_U350 , P2_U3477 , P2_R1179_U40 );
nand NAND2_15941 ( P2_R1179_U351 , P2_U3083 , P2_R1179_U39 );
nand NAND2_15942 ( P2_R1179_U352 , P2_R1179_U220 , P2_R1179_U148 );
nand NAND2_15943 ( P2_R1179_U353 , P2_R1179_U218 , P2_R1179_U147 );
nand NAND2_15944 ( P2_R1179_U354 , P2_U3474 , P2_R1179_U38 );
nand NAND2_15945 ( P2_R1179_U355 , P2_U3084 , P2_R1179_U35 );
nand NAND2_15946 ( P2_R1179_U356 , P2_U3474 , P2_R1179_U38 );
nand NAND2_15947 ( P2_R1179_U357 , P2_U3084 , P2_R1179_U35 );
nand NAND2_15948 ( P2_R1179_U358 , P2_R1179_U357 , P2_R1179_U356 );
nand NAND2_15949 ( P2_R1179_U359 , P2_U3471 , P2_R1179_U36 );
nand NAND2_15950 ( P2_R1179_U360 , P2_U3070 , P2_R1179_U20 );
nand NAND2_15951 ( P2_R1179_U361 , P2_R1179_U225 , P2_R1179_U41 );
nand NAND2_15952 ( P2_R1179_U362 , P2_R1179_U149 , P2_R1179_U212 );
nand NAND2_15953 ( P2_R1179_U363 , P2_U3468 , P2_R1179_U31 );
nand NAND2_15954 ( P2_R1179_U364 , P2_U3071 , P2_R1179_U29 );
nand NAND2_15955 ( P2_R1179_U365 , P2_R1179_U364 , P2_R1179_U363 );
nand NAND2_15956 ( P2_R1179_U366 , P2_U3465 , P2_R1179_U32 );
nand NAND2_15957 ( P2_R1179_U367 , P2_U3067 , P2_R1179_U21 );
nand NAND2_15958 ( P2_R1179_U368 , P2_R1179_U235 , P2_R1179_U42 );
nand NAND2_15959 ( P2_R1179_U369 , P2_R1179_U150 , P2_R1179_U227 );
nand NAND2_15960 ( P2_R1179_U370 , P2_U3462 , P2_R1179_U33 );
nand NAND2_15961 ( P2_R1179_U371 , P2_U3060 , P2_R1179_U30 );
nand NAND2_15962 ( P2_R1179_U372 , P2_R1179_U236 , P2_R1179_U152 );
nand NAND2_15963 ( P2_R1179_U373 , P2_R1179_U202 , P2_R1179_U151 );
nand NAND2_15964 ( P2_R1179_U374 , P2_U3459 , P2_R1179_U28 );
nand NAND2_15965 ( P2_R1179_U375 , P2_U3064 , P2_R1179_U25 );
nand NAND2_15966 ( P2_R1179_U376 , P2_U3459 , P2_R1179_U28 );
nand NAND2_15967 ( P2_R1179_U377 , P2_U3064 , P2_R1179_U25 );
nand NAND2_15968 ( P2_R1179_U378 , P2_R1179_U377 , P2_R1179_U376 );
nand NAND2_15969 ( P2_R1179_U379 , P2_U3456 , P2_R1179_U26 );
nand NAND2_15970 ( P2_R1179_U380 , P2_U3068 , P2_R1179_U22 );
nand NAND2_15971 ( P2_R1179_U381 , P2_R1179_U241 , P2_R1179_U43 );
nand NAND2_15972 ( P2_R1179_U382 , P2_R1179_U153 , P2_R1179_U196 );
nand NAND2_15973 ( P2_R1179_U383 , P2_U3979 , P2_R1179_U155 );
nand NAND2_15974 ( P2_R1179_U384 , P2_U3055 , P2_R1179_U154 );
nand NAND2_15975 ( P2_R1179_U385 , P2_U3979 , P2_R1179_U155 );
nand NAND2_15976 ( P2_R1179_U386 , P2_U3055 , P2_R1179_U154 );
nand NAND2_15977 ( P2_R1179_U387 , P2_R1179_U386 , P2_R1179_U385 );
nand NAND3_15978 ( P2_R1179_U388 , P2_U3968 , P2_R1179_U10 , P2_R1179_U84 );
nand NAND3_15979 ( P2_R1179_U389 , P2_R1179_U387 , P2_R1179_U83 , P2_U3054 );
nand NAND2_15980 ( P2_R1179_U390 , P2_U3968 , P2_R1179_U84 );
nand NAND2_15981 ( P2_R1179_U391 , P2_U3054 , P2_R1179_U83 );
not NOT1_15982 ( P2_R1179_U392 , P2_R1179_U129 );
nand NAND2_15983 ( P2_R1179_U393 , P2_R1179_U306 , P2_R1179_U392 );
nand NAND2_15984 ( P2_R1179_U394 , P2_R1179_U129 , P2_R1179_U157 );
nand NAND2_15985 ( P2_R1179_U395 , P2_U3969 , P2_R1179_U82 );
nand NAND2_15986 ( P2_R1179_U396 , P2_U3053 , P2_R1179_U79 );
nand NAND2_15987 ( P2_R1179_U397 , P2_U3969 , P2_R1179_U82 );
nand NAND2_15988 ( P2_R1179_U398 , P2_U3053 , P2_R1179_U79 );
nand NAND2_15989 ( P2_R1179_U399 , P2_R1179_U398 , P2_R1179_U397 );
nand NAND2_15990 ( P2_R1179_U400 , P2_U3970 , P2_R1179_U80 );
nand NAND2_15991 ( P2_R1179_U401 , P2_U3057 , P2_R1179_U44 );
nand NAND2_15992 ( P2_R1179_U402 , P2_R1179_U313 , P2_R1179_U85 );
nand NAND2_15993 ( P2_R1179_U403 , P2_R1179_U158 , P2_R1179_U300 );
nand NAND2_15994 ( P2_R1179_U404 , P2_U3971 , P2_R1179_U78 );
nand NAND2_15995 ( P2_R1179_U405 , P2_U3058 , P2_R1179_U77 );
not NOT1_15996 ( P2_R1179_U406 , P2_R1179_U132 );
nand NAND2_15997 ( P2_R1179_U407 , P2_R1179_U296 , P2_R1179_U406 );
nand NAND2_15998 ( P2_R1179_U408 , P2_R1179_U132 , P2_R1179_U159 );
nand NAND2_15999 ( P2_R1179_U409 , P2_U3972 , P2_R1179_U76 );
nand NAND2_16000 ( P2_R1179_U410 , P2_U3065 , P2_R1179_U75 );
not NOT1_16001 ( P2_R1179_U411 , P2_R1179_U133 );
nand NAND2_16002 ( P2_R1179_U412 , P2_R1179_U292 , P2_R1179_U411 );
nand NAND2_16003 ( P2_R1179_U413 , P2_R1179_U133 , P2_R1179_U160 );
nand NAND2_16004 ( P2_R1179_U414 , P2_U3973 , P2_R1179_U71 );
nand NAND2_16005 ( P2_R1179_U415 , P2_U3066 , P2_R1179_U69 );
nand NAND2_16006 ( P2_R1179_U416 , P2_R1179_U415 , P2_R1179_U414 );
nand NAND2_16007 ( P2_R1179_U417 , P2_U3974 , P2_R1179_U72 );
nand NAND2_16008 ( P2_R1179_U418 , P2_U3061 , P2_R1179_U45 );
nand NAND2_16009 ( P2_R1179_U419 , P2_R1179_U323 , P2_R1179_U86 );
nand NAND2_16010 ( P2_R1179_U420 , P2_R1179_U161 , P2_R1179_U315 );
nand NAND2_16011 ( P2_R1179_U421 , P2_U3975 , P2_R1179_U73 );
nand NAND2_16012 ( P2_R1179_U422 , P2_U3075 , P2_R1179_U70 );
nand NAND2_16013 ( P2_R1179_U423 , P2_R1179_U324 , P2_R1179_U163 );
nand NAND2_16014 ( P2_R1179_U424 , P2_R1179_U282 , P2_R1179_U162 );
nand NAND2_16015 ( P2_R1179_U425 , P2_U3976 , P2_R1179_U68 );
nand NAND2_16016 ( P2_R1179_U426 , P2_U3076 , P2_R1179_U67 );
not NOT1_16017 ( P2_R1179_U427 , P2_R1179_U136 );
nand NAND2_16018 ( P2_R1179_U428 , P2_R1179_U278 , P2_R1179_U427 );
nand NAND2_16019 ( P2_R1179_U429 , P2_R1179_U136 , P2_R1179_U164 );
nand NAND2_16020 ( P2_R1179_U430 , P2_U3453 , P2_R1179_U24 );
nand NAND2_16021 ( P2_R1179_U431 , P2_U3078 , P2_R1179_U165 );
not NOT1_16022 ( P2_R1179_U432 , P2_R1179_U137 );
nand NAND2_16023 ( P2_R1179_U433 , P2_R1179_U194 , P2_R1179_U432 );
nand NAND2_16024 ( P2_R1179_U434 , P2_R1179_U137 , P2_R1179_U166 );
nand NAND2_16025 ( P2_R1179_U435 , P2_U3506 , P2_R1179_U66 );
nand NAND2_16026 ( P2_R1179_U436 , P2_U3081 , P2_R1179_U65 );
not NOT1_16027 ( P2_R1179_U437 , P2_R1179_U138 );
nand NAND2_16028 ( P2_R1179_U438 , P2_R1179_U274 , P2_R1179_U437 );
nand NAND2_16029 ( P2_R1179_U439 , P2_R1179_U138 , P2_R1179_U167 );
nand NAND2_16030 ( P2_R1179_U440 , P2_U3504 , P2_R1179_U64 );
nand NAND2_16031 ( P2_R1179_U441 , P2_U3082 , P2_R1179_U168 );
not NOT1_16032 ( P2_R1179_U442 , P2_R1179_U139 );
nand NAND2_16033 ( P2_R1179_U443 , P2_R1179_U272 , P2_R1179_U442 );
nand NAND2_16034 ( P2_R1179_U444 , P2_R1179_U139 , P2_R1179_U169 );
nand NAND2_16035 ( P2_R1179_U445 , P2_U3501 , P2_R1179_U63 );
nand NAND2_16036 ( P2_R1179_U446 , P2_U3069 , P2_R1179_U62 );
not NOT1_16037 ( P2_R1179_U447 , P2_R1179_U140 );
nand NAND2_16038 ( P2_R1179_U448 , P2_R1179_U268 , P2_R1179_U447 );
nand NAND2_16039 ( P2_R1179_U449 , P2_R1179_U140 , P2_R1179_U170 );
nand NAND2_16040 ( P2_R1179_U450 , P2_U3498 , P2_R1179_U58 );
nand NAND2_16041 ( P2_R1179_U451 , P2_U3073 , P2_R1179_U56 );
nand NAND2_16042 ( P2_R1179_U452 , P2_R1179_U451 , P2_R1179_U450 );
nand NAND2_16043 ( P2_R1179_U453 , P2_U3495 , P2_R1179_U59 );
nand NAND2_16044 ( P2_R1179_U454 , P2_U3074 , P2_R1179_U46 );
nand NAND2_16045 ( P2_R1179_U455 , P2_R1179_U334 , P2_R1179_U87 );
nand NAND2_16046 ( P2_R1179_U456 , P2_R1179_U171 , P2_R1179_U326 );
nand NAND2_16047 ( P2_R1179_U457 , P2_U3492 , P2_R1179_U60 );
nand NAND2_16048 ( P2_R1179_U458 , P2_U3079 , P2_R1179_U57 );
nand NAND2_16049 ( P2_R1179_U459 , P2_R1179_U335 , P2_R1179_U173 );
nand NAND2_16050 ( P2_R1179_U460 , P2_R1179_U258 , P2_R1179_U172 );
nand NAND2_16051 ( P2_R1179_U461 , P2_U3489 , P2_R1179_U55 );
nand NAND2_16052 ( P2_R1179_U462 , P2_U3080 , P2_R1179_U54 );
not NOT1_16053 ( P2_R1179_U463 , P2_R1179_U143 );
nand NAND2_16054 ( P2_R1179_U464 , P2_R1179_U254 , P2_R1179_U463 );
nand NAND2_16055 ( P2_R1179_U465 , P2_R1179_U143 , P2_R1179_U174 );
nand NAND2_16056 ( P2_R1179_U466 , P2_U3486 , P2_R1179_U53 );
nand NAND2_16057 ( P2_R1179_U467 , P2_U3072 , P2_R1179_U52 );
not NOT1_16058 ( P2_R1179_U468 , P2_R1179_U144 );
nand NAND2_16059 ( P2_R1179_U469 , P2_R1179_U250 , P2_R1179_U468 );
nand NAND2_16060 ( P2_R1179_U470 , P2_R1179_U144 , P2_R1179_U175 );
nand NAND2_16061 ( P2_R1179_U471 , P2_U3483 , P2_R1179_U49 );
nand NAND2_16062 ( P2_R1179_U472 , P2_U3063 , P2_R1179_U48 );
nand NAND2_16063 ( P2_R1179_U473 , P2_R1179_U472 , P2_R1179_U471 );
nand NAND2_16064 ( P2_R1179_U474 , P2_U3480 , P2_R1179_U50 );
nand NAND2_16065 ( P2_R1179_U475 , P2_U3062 , P2_R1179_U47 );
nand NAND2_16066 ( P2_R1179_U476 , P2_R1179_U345 , P2_R1179_U88 );
nand NAND2_16067 ( P2_R1179_U477 , P2_R1179_U176 , P2_R1179_U337 );
and AND2_16068 ( P2_R1215_U4 , P2_R1215_U179 , P2_R1215_U178 );
and AND2_16069 ( P2_R1215_U5 , P2_R1215_U197 , P2_R1215_U196 );
and AND2_16070 ( P2_R1215_U6 , P2_R1215_U237 , P2_R1215_U236 );
and AND2_16071 ( P2_R1215_U7 , P2_R1215_U246 , P2_R1215_U245 );
and AND2_16072 ( P2_R1215_U8 , P2_R1215_U264 , P2_R1215_U263 );
and AND2_16073 ( P2_R1215_U9 , P2_R1215_U272 , P2_R1215_U271 );
and AND2_16074 ( P2_R1215_U10 , P2_R1215_U351 , P2_R1215_U348 );
and AND2_16075 ( P2_R1215_U11 , P2_R1215_U344 , P2_R1215_U341 );
and AND2_16076 ( P2_R1215_U12 , P2_R1215_U335 , P2_R1215_U332 );
and AND2_16077 ( P2_R1215_U13 , P2_R1215_U326 , P2_R1215_U323 );
and AND2_16078 ( P2_R1215_U14 , P2_R1215_U320 , P2_R1215_U318 );
and AND2_16079 ( P2_R1215_U15 , P2_R1215_U313 , P2_R1215_U310 );
and AND2_16080 ( P2_R1215_U16 , P2_R1215_U235 , P2_R1215_U232 );
and AND2_16081 ( P2_R1215_U17 , P2_R1215_U227 , P2_R1215_U224 );
and AND2_16082 ( P2_R1215_U18 , P2_R1215_U213 , P2_R1215_U210 );
not NOT1_16083 ( P2_R1215_U19 , P2_U3468 );
not NOT1_16084 ( P2_R1215_U20 , P2_U3071 );
not NOT1_16085 ( P2_R1215_U21 , P2_U3070 );
nand NAND2_16086 ( P2_R1215_U22 , P2_U3071 , P2_U3468 );
not NOT1_16087 ( P2_R1215_U23 , P2_U3471 );
not NOT1_16088 ( P2_R1215_U24 , P2_U3462 );
not NOT1_16089 ( P2_R1215_U25 , P2_U3060 );
not NOT1_16090 ( P2_R1215_U26 , P2_U3067 );
not NOT1_16091 ( P2_R1215_U27 , P2_U3456 );
not NOT1_16092 ( P2_R1215_U28 , P2_U3068 );
not NOT1_16093 ( P2_R1215_U29 , P2_U3448 );
not NOT1_16094 ( P2_R1215_U30 , P2_U3077 );
nand NAND2_16095 ( P2_R1215_U31 , P2_U3077 , P2_U3448 );
not NOT1_16096 ( P2_R1215_U32 , P2_U3459 );
not NOT1_16097 ( P2_R1215_U33 , P2_U3064 );
nand NAND2_16098 ( P2_R1215_U34 , P2_U3060 , P2_U3462 );
not NOT1_16099 ( P2_R1215_U35 , P2_U3465 );
not NOT1_16100 ( P2_R1215_U36 , P2_U3474 );
not NOT1_16101 ( P2_R1215_U37 , P2_U3084 );
not NOT1_16102 ( P2_R1215_U38 , P2_U3083 );
not NOT1_16103 ( P2_R1215_U39 , P2_U3477 );
nand NAND2_16104 ( P2_R1215_U40 , P2_R1215_U61 , P2_R1215_U205 );
nand NAND2_16105 ( P2_R1215_U41 , P2_R1215_U117 , P2_R1215_U193 );
nand NAND2_16106 ( P2_R1215_U42 , P2_R1215_U182 , P2_R1215_U183 );
nand NAND2_16107 ( P2_R1215_U43 , P2_U3453 , P2_U3078 );
nand NAND2_16108 ( P2_R1215_U44 , P2_R1215_U122 , P2_R1215_U219 );
nand NAND2_16109 ( P2_R1215_U45 , P2_R1215_U216 , P2_R1215_U215 );
not NOT1_16110 ( P2_R1215_U46 , P2_U3969 );
not NOT1_16111 ( P2_R1215_U47 , P2_U3053 );
not NOT1_16112 ( P2_R1215_U48 , P2_U3057 );
not NOT1_16113 ( P2_R1215_U49 , P2_U3970 );
not NOT1_16114 ( P2_R1215_U50 , P2_U3971 );
not NOT1_16115 ( P2_R1215_U51 , P2_U3058 );
not NOT1_16116 ( P2_R1215_U52 , P2_U3972 );
not NOT1_16117 ( P2_R1215_U53 , P2_U3065 );
not NOT1_16118 ( P2_R1215_U54 , P2_U3975 );
not NOT1_16119 ( P2_R1215_U55 , P2_U3075 );
not NOT1_16120 ( P2_R1215_U56 , P2_U3498 );
not NOT1_16121 ( P2_R1215_U57 , P2_U3073 );
not NOT1_16122 ( P2_R1215_U58 , P2_U3069 );
nand NAND2_16123 ( P2_R1215_U59 , P2_U3073 , P2_U3498 );
not NOT1_16124 ( P2_R1215_U60 , P2_U3501 );
nand NAND2_16125 ( P2_R1215_U61 , P2_U3084 , P2_U3474 );
not NOT1_16126 ( P2_R1215_U62 , P2_U3480 );
not NOT1_16127 ( P2_R1215_U63 , P2_U3062 );
not NOT1_16128 ( P2_R1215_U64 , P2_U3486 );
not NOT1_16129 ( P2_R1215_U65 , P2_U3072 );
not NOT1_16130 ( P2_R1215_U66 , P2_U3483 );
not NOT1_16131 ( P2_R1215_U67 , P2_U3063 );
nand NAND2_16132 ( P2_R1215_U68 , P2_U3063 , P2_U3483 );
not NOT1_16133 ( P2_R1215_U69 , P2_U3489 );
not NOT1_16134 ( P2_R1215_U70 , P2_U3080 );
not NOT1_16135 ( P2_R1215_U71 , P2_U3492 );
not NOT1_16136 ( P2_R1215_U72 , P2_U3079 );
not NOT1_16137 ( P2_R1215_U73 , P2_U3495 );
not NOT1_16138 ( P2_R1215_U74 , P2_U3074 );
not NOT1_16139 ( P2_R1215_U75 , P2_U3504 );
not NOT1_16140 ( P2_R1215_U76 , P2_U3082 );
nand NAND2_16141 ( P2_R1215_U77 , P2_U3082 , P2_U3504 );
not NOT1_16142 ( P2_R1215_U78 , P2_U3506 );
not NOT1_16143 ( P2_R1215_U79 , P2_U3081 );
nand NAND2_16144 ( P2_R1215_U80 , P2_U3081 , P2_U3506 );
not NOT1_16145 ( P2_R1215_U81 , P2_U3976 );
not NOT1_16146 ( P2_R1215_U82 , P2_U3974 );
not NOT1_16147 ( P2_R1215_U83 , P2_U3061 );
not NOT1_16148 ( P2_R1215_U84 , P2_U3973 );
not NOT1_16149 ( P2_R1215_U85 , P2_U3066 );
nand NAND2_16150 ( P2_R1215_U86 , P2_U3970 , P2_U3057 );
not NOT1_16151 ( P2_R1215_U87 , P2_U3054 );
not NOT1_16152 ( P2_R1215_U88 , P2_U3968 );
nand NAND2_16153 ( P2_R1215_U89 , P2_R1215_U306 , P2_R1215_U176 );
not NOT1_16154 ( P2_R1215_U90 , P2_U3076 );
nand NAND2_16155 ( P2_R1215_U91 , P2_R1215_U77 , P2_R1215_U315 );
nand NAND2_16156 ( P2_R1215_U92 , P2_R1215_U261 , P2_R1215_U260 );
nand NAND2_16157 ( P2_R1215_U93 , P2_R1215_U68 , P2_R1215_U337 );
nand NAND2_16158 ( P2_R1215_U94 , P2_R1215_U457 , P2_R1215_U456 );
nand NAND2_16159 ( P2_R1215_U95 , P2_R1215_U504 , P2_R1215_U503 );
nand NAND2_16160 ( P2_R1215_U96 , P2_R1215_U375 , P2_R1215_U374 );
nand NAND2_16161 ( P2_R1215_U97 , P2_R1215_U380 , P2_R1215_U379 );
nand NAND2_16162 ( P2_R1215_U98 , P2_R1215_U387 , P2_R1215_U386 );
nand NAND2_16163 ( P2_R1215_U99 , P2_R1215_U394 , P2_R1215_U393 );
nand NAND2_16164 ( P2_R1215_U100 , P2_R1215_U399 , P2_R1215_U398 );
nand NAND2_16165 ( P2_R1215_U101 , P2_R1215_U408 , P2_R1215_U407 );
nand NAND2_16166 ( P2_R1215_U102 , P2_R1215_U415 , P2_R1215_U414 );
nand NAND2_16167 ( P2_R1215_U103 , P2_R1215_U422 , P2_R1215_U421 );
nand NAND2_16168 ( P2_R1215_U104 , P2_R1215_U429 , P2_R1215_U428 );
nand NAND2_16169 ( P2_R1215_U105 , P2_R1215_U434 , P2_R1215_U433 );
nand NAND2_16170 ( P2_R1215_U106 , P2_R1215_U441 , P2_R1215_U440 );
nand NAND2_16171 ( P2_R1215_U107 , P2_R1215_U448 , P2_R1215_U447 );
nand NAND2_16172 ( P2_R1215_U108 , P2_R1215_U462 , P2_R1215_U461 );
nand NAND2_16173 ( P2_R1215_U109 , P2_R1215_U467 , P2_R1215_U466 );
nand NAND2_16174 ( P2_R1215_U110 , P2_R1215_U474 , P2_R1215_U473 );
nand NAND2_16175 ( P2_R1215_U111 , P2_R1215_U481 , P2_R1215_U480 );
nand NAND2_16176 ( P2_R1215_U112 , P2_R1215_U488 , P2_R1215_U487 );
nand NAND2_16177 ( P2_R1215_U113 , P2_R1215_U495 , P2_R1215_U494 );
nand NAND2_16178 ( P2_R1215_U114 , P2_R1215_U500 , P2_R1215_U499 );
and AND2_16179 ( P2_R1215_U115 , P2_R1215_U189 , P2_R1215_U187 );
and AND2_16180 ( P2_R1215_U116 , P2_R1215_U4 , P2_R1215_U180 );
and AND2_16181 ( P2_R1215_U117 , P2_R1215_U194 , P2_R1215_U192 );
and AND2_16182 ( P2_R1215_U118 , P2_R1215_U201 , P2_R1215_U200 );
and AND3_16183 ( P2_R1215_U119 , P2_R1215_U382 , P2_R1215_U381 , P2_R1215_U22 );
and AND2_16184 ( P2_R1215_U120 , P2_R1215_U212 , P2_R1215_U5 );
and AND2_16185 ( P2_R1215_U121 , P2_R1215_U181 , P2_R1215_U180 );
and AND2_16186 ( P2_R1215_U122 , P2_R1215_U220 , P2_R1215_U218 );
and AND3_16187 ( P2_R1215_U123 , P2_R1215_U389 , P2_R1215_U388 , P2_R1215_U34 );
and AND2_16188 ( P2_R1215_U124 , P2_R1215_U226 , P2_R1215_U4 );
and AND2_16189 ( P2_R1215_U125 , P2_R1215_U234 , P2_R1215_U181 );
and AND2_16190 ( P2_R1215_U126 , P2_R1215_U204 , P2_R1215_U6 );
and AND2_16191 ( P2_R1215_U127 , P2_R1215_U239 , P2_R1215_U171 );
and AND2_16192 ( P2_R1215_U128 , P2_R1215_U250 , P2_R1215_U7 );
and AND2_16193 ( P2_R1215_U129 , P2_R1215_U248 , P2_R1215_U172 );
and AND2_16194 ( P2_R1215_U130 , P2_R1215_U268 , P2_R1215_U267 );
and AND3_16195 ( P2_R1215_U131 , P2_R1215_U9 , P2_R1215_U282 , P2_R1215_U273 );
and AND2_16196 ( P2_R1215_U132 , P2_R1215_U285 , P2_R1215_U280 );
and AND2_16197 ( P2_R1215_U133 , P2_R1215_U301 , P2_R1215_U298 );
and AND2_16198 ( P2_R1215_U134 , P2_R1215_U368 , P2_R1215_U302 );
and AND3_16199 ( P2_R1215_U135 , P2_R1215_U424 , P2_R1215_U423 , P2_R1215_U173 );
and AND2_16200 ( P2_R1215_U136 , P2_R1215_U160 , P2_R1215_U278 );
and AND3_16201 ( P2_R1215_U137 , P2_R1215_U455 , P2_R1215_U454 , P2_R1215_U80 );
and AND2_16202 ( P2_R1215_U138 , P2_R1215_U325 , P2_R1215_U9 );
and AND3_16203 ( P2_R1215_U139 , P2_R1215_U469 , P2_R1215_U468 , P2_R1215_U59 );
and AND2_16204 ( P2_R1215_U140 , P2_R1215_U334 , P2_R1215_U8 );
and AND3_16205 ( P2_R1215_U141 , P2_R1215_U490 , P2_R1215_U489 , P2_R1215_U172 );
and AND2_16206 ( P2_R1215_U142 , P2_R1215_U343 , P2_R1215_U7 );
and AND3_16207 ( P2_R1215_U143 , P2_R1215_U502 , P2_R1215_U501 , P2_R1215_U171 );
and AND2_16208 ( P2_R1215_U144 , P2_R1215_U350 , P2_R1215_U6 );
nand NAND2_16209 ( P2_R1215_U145 , P2_R1215_U118 , P2_R1215_U202 );
nand NAND2_16210 ( P2_R1215_U146 , P2_R1215_U217 , P2_R1215_U229 );
not NOT1_16211 ( P2_R1215_U147 , P2_U3055 );
not NOT1_16212 ( P2_R1215_U148 , P2_U3979 );
and AND2_16213 ( P2_R1215_U149 , P2_R1215_U403 , P2_R1215_U402 );
nand NAND3_16214 ( P2_R1215_U150 , P2_R1215_U304 , P2_R1215_U169 , P2_R1215_U364 );
and AND2_16215 ( P2_R1215_U151 , P2_R1215_U410 , P2_R1215_U409 );
nand NAND3_16216 ( P2_R1215_U152 , P2_R1215_U370 , P2_R1215_U369 , P2_R1215_U134 );
and AND2_16217 ( P2_R1215_U153 , P2_R1215_U417 , P2_R1215_U416 );
nand NAND3_16218 ( P2_R1215_U154 , P2_R1215_U365 , P2_R1215_U299 , P2_R1215_U86 );
nand NAND2_16219 ( P2_R1215_U155 , P2_R1215_U293 , P2_R1215_U292 );
and AND2_16220 ( P2_R1215_U156 , P2_R1215_U436 , P2_R1215_U435 );
nand NAND2_16221 ( P2_R1215_U157 , P2_R1215_U289 , P2_R1215_U288 );
and AND2_16222 ( P2_R1215_U158 , P2_R1215_U443 , P2_R1215_U442 );
nand NAND2_16223 ( P2_R1215_U159 , P2_R1215_U132 , P2_R1215_U284 );
and AND2_16224 ( P2_R1215_U160 , P2_R1215_U450 , P2_R1215_U449 );
nand NAND2_16225 ( P2_R1215_U161 , P2_R1215_U43 , P2_R1215_U327 );
nand NAND2_16226 ( P2_R1215_U162 , P2_R1215_U130 , P2_R1215_U269 );
and AND2_16227 ( P2_R1215_U163 , P2_R1215_U476 , P2_R1215_U475 );
nand NAND2_16228 ( P2_R1215_U164 , P2_R1215_U257 , P2_R1215_U256 );
and AND2_16229 ( P2_R1215_U165 , P2_R1215_U483 , P2_R1215_U482 );
nand NAND2_16230 ( P2_R1215_U166 , P2_R1215_U253 , P2_R1215_U252 );
nand NAND2_16231 ( P2_R1215_U167 , P2_R1215_U243 , P2_R1215_U242 );
nand NAND2_16232 ( P2_R1215_U168 , P2_R1215_U367 , P2_R1215_U366 );
nand NAND2_16233 ( P2_R1215_U169 , P2_U3054 , P2_R1215_U152 );
not NOT1_16234 ( P2_R1215_U170 , P2_R1215_U34 );
nand NAND2_16235 ( P2_R1215_U171 , P2_U3477 , P2_U3083 );
nand NAND2_16236 ( P2_R1215_U172 , P2_U3072 , P2_U3486 );
nand NAND2_16237 ( P2_R1215_U173 , P2_U3058 , P2_U3971 );
not NOT1_16238 ( P2_R1215_U174 , P2_R1215_U68 );
not NOT1_16239 ( P2_R1215_U175 , P2_R1215_U77 );
nand NAND2_16240 ( P2_R1215_U176 , P2_U3065 , P2_U3972 );
not NOT1_16241 ( P2_R1215_U177 , P2_R1215_U61 );
or OR2_16242 ( P2_R1215_U178 , P2_U3067 , P2_U3465 );
or OR2_16243 ( P2_R1215_U179 , P2_U3060 , P2_U3462 );
or OR2_16244 ( P2_R1215_U180 , P2_U3459 , P2_U3064 );
or OR2_16245 ( P2_R1215_U181 , P2_U3456 , P2_U3068 );
not NOT1_16246 ( P2_R1215_U182 , P2_R1215_U31 );
or OR2_16247 ( P2_R1215_U183 , P2_U3453 , P2_U3078 );
not NOT1_16248 ( P2_R1215_U184 , P2_R1215_U42 );
not NOT1_16249 ( P2_R1215_U185 , P2_R1215_U43 );
nand NAND2_16250 ( P2_R1215_U186 , P2_R1215_U42 , P2_R1215_U43 );
nand NAND2_16251 ( P2_R1215_U187 , P2_U3068 , P2_U3456 );
nand NAND2_16252 ( P2_R1215_U188 , P2_R1215_U186 , P2_R1215_U181 );
nand NAND2_16253 ( P2_R1215_U189 , P2_U3064 , P2_U3459 );
nand NAND2_16254 ( P2_R1215_U190 , P2_R1215_U115 , P2_R1215_U188 );
nand NAND2_16255 ( P2_R1215_U191 , P2_R1215_U35 , P2_R1215_U34 );
nand NAND2_16256 ( P2_R1215_U192 , P2_U3067 , P2_R1215_U191 );
nand NAND2_16257 ( P2_R1215_U193 , P2_R1215_U116 , P2_R1215_U190 );
nand NAND2_16258 ( P2_R1215_U194 , P2_U3465 , P2_R1215_U170 );
not NOT1_16259 ( P2_R1215_U195 , P2_R1215_U41 );
or OR2_16260 ( P2_R1215_U196 , P2_U3070 , P2_U3471 );
or OR2_16261 ( P2_R1215_U197 , P2_U3071 , P2_U3468 );
not NOT1_16262 ( P2_R1215_U198 , P2_R1215_U22 );
nand NAND2_16263 ( P2_R1215_U199 , P2_R1215_U23 , P2_R1215_U22 );
nand NAND2_16264 ( P2_R1215_U200 , P2_U3070 , P2_R1215_U199 );
nand NAND2_16265 ( P2_R1215_U201 , P2_U3471 , P2_R1215_U198 );
nand NAND2_16266 ( P2_R1215_U202 , P2_R1215_U5 , P2_R1215_U41 );
not NOT1_16267 ( P2_R1215_U203 , P2_R1215_U145 );
or OR2_16268 ( P2_R1215_U204 , P2_U3474 , P2_U3084 );
nand NAND2_16269 ( P2_R1215_U205 , P2_R1215_U204 , P2_R1215_U145 );
not NOT1_16270 ( P2_R1215_U206 , P2_R1215_U40 );
or OR2_16271 ( P2_R1215_U207 , P2_U3083 , P2_U3477 );
or OR2_16272 ( P2_R1215_U208 , P2_U3468 , P2_U3071 );
nand NAND2_16273 ( P2_R1215_U209 , P2_R1215_U208 , P2_R1215_U41 );
nand NAND2_16274 ( P2_R1215_U210 , P2_R1215_U119 , P2_R1215_U209 );
nand NAND2_16275 ( P2_R1215_U211 , P2_R1215_U195 , P2_R1215_U22 );
nand NAND2_16276 ( P2_R1215_U212 , P2_U3471 , P2_U3070 );
nand NAND2_16277 ( P2_R1215_U213 , P2_R1215_U120 , P2_R1215_U211 );
or OR2_16278 ( P2_R1215_U214 , P2_U3071 , P2_U3468 );
nand NAND2_16279 ( P2_R1215_U215 , P2_R1215_U185 , P2_R1215_U181 );
nand NAND2_16280 ( P2_R1215_U216 , P2_U3068 , P2_U3456 );
not NOT1_16281 ( P2_R1215_U217 , P2_R1215_U45 );
nand NAND2_16282 ( P2_R1215_U218 , P2_R1215_U121 , P2_R1215_U184 );
nand NAND2_16283 ( P2_R1215_U219 , P2_R1215_U45 , P2_R1215_U180 );
nand NAND2_16284 ( P2_R1215_U220 , P2_U3064 , P2_U3459 );
not NOT1_16285 ( P2_R1215_U221 , P2_R1215_U44 );
or OR2_16286 ( P2_R1215_U222 , P2_U3462 , P2_U3060 );
nand NAND2_16287 ( P2_R1215_U223 , P2_R1215_U222 , P2_R1215_U44 );
nand NAND2_16288 ( P2_R1215_U224 , P2_R1215_U123 , P2_R1215_U223 );
nand NAND2_16289 ( P2_R1215_U225 , P2_R1215_U221 , P2_R1215_U34 );
nand NAND2_16290 ( P2_R1215_U226 , P2_U3465 , P2_U3067 );
nand NAND2_16291 ( P2_R1215_U227 , P2_R1215_U124 , P2_R1215_U225 );
or OR2_16292 ( P2_R1215_U228 , P2_U3060 , P2_U3462 );
nand NAND2_16293 ( P2_R1215_U229 , P2_R1215_U184 , P2_R1215_U181 );
not NOT1_16294 ( P2_R1215_U230 , P2_R1215_U146 );
nand NAND2_16295 ( P2_R1215_U231 , P2_U3064 , P2_U3459 );
nand NAND4_16296 ( P2_R1215_U232 , P2_R1215_U401 , P2_R1215_U400 , P2_R1215_U43 , P2_R1215_U42 );
nand NAND2_16297 ( P2_R1215_U233 , P2_R1215_U43 , P2_R1215_U42 );
nand NAND2_16298 ( P2_R1215_U234 , P2_U3068 , P2_U3456 );
nand NAND2_16299 ( P2_R1215_U235 , P2_R1215_U125 , P2_R1215_U233 );
or OR2_16300 ( P2_R1215_U236 , P2_U3083 , P2_U3477 );
or OR2_16301 ( P2_R1215_U237 , P2_U3062 , P2_U3480 );
nand NAND2_16302 ( P2_R1215_U238 , P2_R1215_U177 , P2_R1215_U6 );
nand NAND2_16303 ( P2_R1215_U239 , P2_U3062 , P2_U3480 );
nand NAND2_16304 ( P2_R1215_U240 , P2_R1215_U127 , P2_R1215_U238 );
or OR2_16305 ( P2_R1215_U241 , P2_U3480 , P2_U3062 );
nand NAND2_16306 ( P2_R1215_U242 , P2_R1215_U126 , P2_R1215_U145 );
nand NAND2_16307 ( P2_R1215_U243 , P2_R1215_U241 , P2_R1215_U240 );
not NOT1_16308 ( P2_R1215_U244 , P2_R1215_U167 );
or OR2_16309 ( P2_R1215_U245 , P2_U3080 , P2_U3489 );
or OR2_16310 ( P2_R1215_U246 , P2_U3072 , P2_U3486 );
nand NAND2_16311 ( P2_R1215_U247 , P2_R1215_U174 , P2_R1215_U7 );
nand NAND2_16312 ( P2_R1215_U248 , P2_U3080 , P2_U3489 );
nand NAND2_16313 ( P2_R1215_U249 , P2_R1215_U129 , P2_R1215_U247 );
or OR2_16314 ( P2_R1215_U250 , P2_U3483 , P2_U3063 );
or OR2_16315 ( P2_R1215_U251 , P2_U3489 , P2_U3080 );
nand NAND2_16316 ( P2_R1215_U252 , P2_R1215_U128 , P2_R1215_U167 );
nand NAND2_16317 ( P2_R1215_U253 , P2_R1215_U251 , P2_R1215_U249 );
not NOT1_16318 ( P2_R1215_U254 , P2_R1215_U166 );
or OR2_16319 ( P2_R1215_U255 , P2_U3492 , P2_U3079 );
nand NAND2_16320 ( P2_R1215_U256 , P2_R1215_U255 , P2_R1215_U166 );
nand NAND2_16321 ( P2_R1215_U257 , P2_U3079 , P2_U3492 );
not NOT1_16322 ( P2_R1215_U258 , P2_R1215_U164 );
or OR2_16323 ( P2_R1215_U259 , P2_U3495 , P2_U3074 );
nand NAND2_16324 ( P2_R1215_U260 , P2_R1215_U259 , P2_R1215_U164 );
nand NAND2_16325 ( P2_R1215_U261 , P2_U3074 , P2_U3495 );
not NOT1_16326 ( P2_R1215_U262 , P2_R1215_U92 );
or OR2_16327 ( P2_R1215_U263 , P2_U3069 , P2_U3501 );
or OR2_16328 ( P2_R1215_U264 , P2_U3073 , P2_U3498 );
not NOT1_16329 ( P2_R1215_U265 , P2_R1215_U59 );
nand NAND2_16330 ( P2_R1215_U266 , P2_R1215_U60 , P2_R1215_U59 );
nand NAND2_16331 ( P2_R1215_U267 , P2_U3069 , P2_R1215_U266 );
nand NAND2_16332 ( P2_R1215_U268 , P2_U3501 , P2_R1215_U265 );
nand NAND2_16333 ( P2_R1215_U269 , P2_R1215_U8 , P2_R1215_U92 );
not NOT1_16334 ( P2_R1215_U270 , P2_R1215_U162 );
or OR2_16335 ( P2_R1215_U271 , P2_U3076 , P2_U3976 );
or OR2_16336 ( P2_R1215_U272 , P2_U3081 , P2_U3506 );
or OR2_16337 ( P2_R1215_U273 , P2_U3075 , P2_U3975 );
not NOT1_16338 ( P2_R1215_U274 , P2_R1215_U80 );
nand NAND2_16339 ( P2_R1215_U275 , P2_U3976 , P2_R1215_U274 );
nand NAND2_16340 ( P2_R1215_U276 , P2_R1215_U275 , P2_R1215_U90 );
nand NAND2_16341 ( P2_R1215_U277 , P2_R1215_U80 , P2_R1215_U81 );
nand NAND2_16342 ( P2_R1215_U278 , P2_R1215_U277 , P2_R1215_U276 );
nand NAND2_16343 ( P2_R1215_U279 , P2_R1215_U175 , P2_R1215_U9 );
nand NAND2_16344 ( P2_R1215_U280 , P2_U3075 , P2_U3975 );
nand NAND2_16345 ( P2_R1215_U281 , P2_R1215_U278 , P2_R1215_U279 );
or OR2_16346 ( P2_R1215_U282 , P2_U3504 , P2_U3082 );
or OR2_16347 ( P2_R1215_U283 , P2_U3975 , P2_U3075 );
nand NAND2_16348 ( P2_R1215_U284 , P2_R1215_U162 , P2_R1215_U131 );
nand NAND2_16349 ( P2_R1215_U285 , P2_R1215_U283 , P2_R1215_U281 );
not NOT1_16350 ( P2_R1215_U286 , P2_R1215_U159 );
or OR2_16351 ( P2_R1215_U287 , P2_U3974 , P2_U3061 );
nand NAND2_16352 ( P2_R1215_U288 , P2_R1215_U287 , P2_R1215_U159 );
nand NAND2_16353 ( P2_R1215_U289 , P2_U3061 , P2_U3974 );
not NOT1_16354 ( P2_R1215_U290 , P2_R1215_U157 );
or OR2_16355 ( P2_R1215_U291 , P2_U3973 , P2_U3066 );
nand NAND2_16356 ( P2_R1215_U292 , P2_R1215_U291 , P2_R1215_U157 );
nand NAND2_16357 ( P2_R1215_U293 , P2_U3066 , P2_U3973 );
not NOT1_16358 ( P2_R1215_U294 , P2_R1215_U155 );
or OR2_16359 ( P2_R1215_U295 , P2_U3058 , P2_U3971 );
nand NAND2_16360 ( P2_R1215_U296 , P2_R1215_U176 , P2_R1215_U173 );
not NOT1_16361 ( P2_R1215_U297 , P2_R1215_U86 );
or OR2_16362 ( P2_R1215_U298 , P2_U3972 , P2_U3065 );
nand NAND3_16363 ( P2_R1215_U299 , P2_R1215_U155 , P2_R1215_U298 , P2_R1215_U168 );
not NOT1_16364 ( P2_R1215_U300 , P2_R1215_U154 );
or OR2_16365 ( P2_R1215_U301 , P2_U3969 , P2_U3053 );
nand NAND2_16366 ( P2_R1215_U302 , P2_U3053 , P2_U3969 );
not NOT1_16367 ( P2_R1215_U303 , P2_R1215_U152 );
nand NAND2_16368 ( P2_R1215_U304 , P2_U3968 , P2_R1215_U152 );
not NOT1_16369 ( P2_R1215_U305 , P2_R1215_U150 );
nand NAND2_16370 ( P2_R1215_U306 , P2_R1215_U298 , P2_R1215_U155 );
not NOT1_16371 ( P2_R1215_U307 , P2_R1215_U89 );
or OR2_16372 ( P2_R1215_U308 , P2_U3971 , P2_U3058 );
nand NAND2_16373 ( P2_R1215_U309 , P2_R1215_U308 , P2_R1215_U89 );
nand NAND2_16374 ( P2_R1215_U310 , P2_R1215_U135 , P2_R1215_U309 );
nand NAND2_16375 ( P2_R1215_U311 , P2_R1215_U307 , P2_R1215_U173 );
nand NAND2_16376 ( P2_R1215_U312 , P2_U3970 , P2_U3057 );
nand NAND3_16377 ( P2_R1215_U313 , P2_R1215_U311 , P2_R1215_U312 , P2_R1215_U168 );
or OR2_16378 ( P2_R1215_U314 , P2_U3058 , P2_U3971 );
nand NAND2_16379 ( P2_R1215_U315 , P2_R1215_U282 , P2_R1215_U162 );
not NOT1_16380 ( P2_R1215_U316 , P2_R1215_U91 );
nand NAND2_16381 ( P2_R1215_U317 , P2_R1215_U9 , P2_R1215_U91 );
nand NAND2_16382 ( P2_R1215_U318 , P2_R1215_U136 , P2_R1215_U317 );
nand NAND2_16383 ( P2_R1215_U319 , P2_R1215_U317 , P2_R1215_U278 );
nand NAND2_16384 ( P2_R1215_U320 , P2_R1215_U453 , P2_R1215_U319 );
or OR2_16385 ( P2_R1215_U321 , P2_U3506 , P2_U3081 );
nand NAND2_16386 ( P2_R1215_U322 , P2_R1215_U321 , P2_R1215_U91 );
nand NAND2_16387 ( P2_R1215_U323 , P2_R1215_U137 , P2_R1215_U322 );
nand NAND2_16388 ( P2_R1215_U324 , P2_R1215_U316 , P2_R1215_U80 );
nand NAND2_16389 ( P2_R1215_U325 , P2_U3076 , P2_U3976 );
nand NAND2_16390 ( P2_R1215_U326 , P2_R1215_U138 , P2_R1215_U324 );
or OR2_16391 ( P2_R1215_U327 , P2_U3453 , P2_U3078 );
not NOT1_16392 ( P2_R1215_U328 , P2_R1215_U161 );
or OR2_16393 ( P2_R1215_U329 , P2_U3081 , P2_U3506 );
or OR2_16394 ( P2_R1215_U330 , P2_U3498 , P2_U3073 );
nand NAND2_16395 ( P2_R1215_U331 , P2_R1215_U330 , P2_R1215_U92 );
nand NAND2_16396 ( P2_R1215_U332 , P2_R1215_U139 , P2_R1215_U331 );
nand NAND2_16397 ( P2_R1215_U333 , P2_R1215_U262 , P2_R1215_U59 );
nand NAND2_16398 ( P2_R1215_U334 , P2_U3501 , P2_U3069 );
nand NAND2_16399 ( P2_R1215_U335 , P2_R1215_U140 , P2_R1215_U333 );
or OR2_16400 ( P2_R1215_U336 , P2_U3073 , P2_U3498 );
nand NAND2_16401 ( P2_R1215_U337 , P2_R1215_U250 , P2_R1215_U167 );
not NOT1_16402 ( P2_R1215_U338 , P2_R1215_U93 );
or OR2_16403 ( P2_R1215_U339 , P2_U3486 , P2_U3072 );
nand NAND2_16404 ( P2_R1215_U340 , P2_R1215_U339 , P2_R1215_U93 );
nand NAND2_16405 ( P2_R1215_U341 , P2_R1215_U141 , P2_R1215_U340 );
nand NAND2_16406 ( P2_R1215_U342 , P2_R1215_U338 , P2_R1215_U172 );
nand NAND2_16407 ( P2_R1215_U343 , P2_U3080 , P2_U3489 );
nand NAND2_16408 ( P2_R1215_U344 , P2_R1215_U142 , P2_R1215_U342 );
or OR2_16409 ( P2_R1215_U345 , P2_U3072 , P2_U3486 );
or OR2_16410 ( P2_R1215_U346 , P2_U3477 , P2_U3083 );
nand NAND2_16411 ( P2_R1215_U347 , P2_R1215_U346 , P2_R1215_U40 );
nand NAND2_16412 ( P2_R1215_U348 , P2_R1215_U143 , P2_R1215_U347 );
nand NAND2_16413 ( P2_R1215_U349 , P2_R1215_U206 , P2_R1215_U171 );
nand NAND2_16414 ( P2_R1215_U350 , P2_U3062 , P2_U3480 );
nand NAND2_16415 ( P2_R1215_U351 , P2_R1215_U144 , P2_R1215_U349 );
nand NAND2_16416 ( P2_R1215_U352 , P2_R1215_U207 , P2_R1215_U171 );
nand NAND2_16417 ( P2_R1215_U353 , P2_R1215_U204 , P2_R1215_U61 );
nand NAND2_16418 ( P2_R1215_U354 , P2_R1215_U214 , P2_R1215_U22 );
nand NAND2_16419 ( P2_R1215_U355 , P2_R1215_U228 , P2_R1215_U34 );
nand NAND2_16420 ( P2_R1215_U356 , P2_R1215_U231 , P2_R1215_U180 );
nand NAND2_16421 ( P2_R1215_U357 , P2_R1215_U314 , P2_R1215_U173 );
nand NAND2_16422 ( P2_R1215_U358 , P2_R1215_U298 , P2_R1215_U176 );
nand NAND2_16423 ( P2_R1215_U359 , P2_R1215_U329 , P2_R1215_U80 );
nand NAND2_16424 ( P2_R1215_U360 , P2_R1215_U282 , P2_R1215_U77 );
nand NAND2_16425 ( P2_R1215_U361 , P2_R1215_U336 , P2_R1215_U59 );
nand NAND2_16426 ( P2_R1215_U362 , P2_R1215_U345 , P2_R1215_U172 );
nand NAND2_16427 ( P2_R1215_U363 , P2_R1215_U250 , P2_R1215_U68 );
nand NAND2_16428 ( P2_R1215_U364 , P2_U3968 , P2_U3054 );
nand NAND2_16429 ( P2_R1215_U365 , P2_R1215_U296 , P2_R1215_U168 );
nand NAND2_16430 ( P2_R1215_U366 , P2_U3057 , P2_R1215_U295 );
nand NAND2_16431 ( P2_R1215_U367 , P2_U3970 , P2_R1215_U295 );
nand NAND3_16432 ( P2_R1215_U368 , P2_R1215_U296 , P2_R1215_U168 , P2_R1215_U301 );
nand NAND3_16433 ( P2_R1215_U369 , P2_R1215_U155 , P2_R1215_U168 , P2_R1215_U133 );
nand NAND2_16434 ( P2_R1215_U370 , P2_R1215_U297 , P2_R1215_U301 );
nand NAND2_16435 ( P2_R1215_U371 , P2_U3083 , P2_R1215_U39 );
nand NAND2_16436 ( P2_R1215_U372 , P2_U3477 , P2_R1215_U38 );
nand NAND2_16437 ( P2_R1215_U373 , P2_R1215_U372 , P2_R1215_U371 );
nand NAND2_16438 ( P2_R1215_U374 , P2_R1215_U352 , P2_R1215_U40 );
nand NAND2_16439 ( P2_R1215_U375 , P2_R1215_U373 , P2_R1215_U206 );
nand NAND2_16440 ( P2_R1215_U376 , P2_U3084 , P2_R1215_U36 );
nand NAND2_16441 ( P2_R1215_U377 , P2_U3474 , P2_R1215_U37 );
nand NAND2_16442 ( P2_R1215_U378 , P2_R1215_U377 , P2_R1215_U376 );
nand NAND2_16443 ( P2_R1215_U379 , P2_R1215_U353 , P2_R1215_U145 );
nand NAND2_16444 ( P2_R1215_U380 , P2_R1215_U203 , P2_R1215_U378 );
nand NAND2_16445 ( P2_R1215_U381 , P2_U3070 , P2_R1215_U23 );
nand NAND2_16446 ( P2_R1215_U382 , P2_U3471 , P2_R1215_U21 );
nand NAND2_16447 ( P2_R1215_U383 , P2_U3071 , P2_R1215_U19 );
nand NAND2_16448 ( P2_R1215_U384 , P2_U3468 , P2_R1215_U20 );
nand NAND2_16449 ( P2_R1215_U385 , P2_R1215_U384 , P2_R1215_U383 );
nand NAND2_16450 ( P2_R1215_U386 , P2_R1215_U354 , P2_R1215_U41 );
nand NAND2_16451 ( P2_R1215_U387 , P2_R1215_U385 , P2_R1215_U195 );
nand NAND2_16452 ( P2_R1215_U388 , P2_U3067 , P2_R1215_U35 );
nand NAND2_16453 ( P2_R1215_U389 , P2_U3465 , P2_R1215_U26 );
nand NAND2_16454 ( P2_R1215_U390 , P2_U3060 , P2_R1215_U24 );
nand NAND2_16455 ( P2_R1215_U391 , P2_U3462 , P2_R1215_U25 );
nand NAND2_16456 ( P2_R1215_U392 , P2_R1215_U391 , P2_R1215_U390 );
nand NAND2_16457 ( P2_R1215_U393 , P2_R1215_U355 , P2_R1215_U44 );
nand NAND2_16458 ( P2_R1215_U394 , P2_R1215_U392 , P2_R1215_U221 );
nand NAND2_16459 ( P2_R1215_U395 , P2_U3064 , P2_R1215_U32 );
nand NAND2_16460 ( P2_R1215_U396 , P2_U3459 , P2_R1215_U33 );
nand NAND2_16461 ( P2_R1215_U397 , P2_R1215_U396 , P2_R1215_U395 );
nand NAND2_16462 ( P2_R1215_U398 , P2_R1215_U356 , P2_R1215_U146 );
nand NAND2_16463 ( P2_R1215_U399 , P2_R1215_U230 , P2_R1215_U397 );
nand NAND2_16464 ( P2_R1215_U400 , P2_U3068 , P2_R1215_U27 );
nand NAND2_16465 ( P2_R1215_U401 , P2_U3456 , P2_R1215_U28 );
nand NAND2_16466 ( P2_R1215_U402 , P2_U3055 , P2_R1215_U148 );
nand NAND2_16467 ( P2_R1215_U403 , P2_U3979 , P2_R1215_U147 );
nand NAND2_16468 ( P2_R1215_U404 , P2_U3055 , P2_R1215_U148 );
nand NAND2_16469 ( P2_R1215_U405 , P2_U3979 , P2_R1215_U147 );
nand NAND2_16470 ( P2_R1215_U406 , P2_R1215_U405 , P2_R1215_U404 );
nand NAND2_16471 ( P2_R1215_U407 , P2_R1215_U149 , P2_R1215_U150 );
nand NAND2_16472 ( P2_R1215_U408 , P2_R1215_U305 , P2_R1215_U406 );
nand NAND2_16473 ( P2_R1215_U409 , P2_U3054 , P2_R1215_U88 );
nand NAND2_16474 ( P2_R1215_U410 , P2_U3968 , P2_R1215_U87 );
nand NAND2_16475 ( P2_R1215_U411 , P2_U3054 , P2_R1215_U88 );
nand NAND2_16476 ( P2_R1215_U412 , P2_U3968 , P2_R1215_U87 );
nand NAND2_16477 ( P2_R1215_U413 , P2_R1215_U412 , P2_R1215_U411 );
nand NAND2_16478 ( P2_R1215_U414 , P2_R1215_U151 , P2_R1215_U152 );
nand NAND2_16479 ( P2_R1215_U415 , P2_R1215_U303 , P2_R1215_U413 );
nand NAND2_16480 ( P2_R1215_U416 , P2_U3053 , P2_R1215_U46 );
nand NAND2_16481 ( P2_R1215_U417 , P2_U3969 , P2_R1215_U47 );
nand NAND2_16482 ( P2_R1215_U418 , P2_U3053 , P2_R1215_U46 );
nand NAND2_16483 ( P2_R1215_U419 , P2_U3969 , P2_R1215_U47 );
nand NAND2_16484 ( P2_R1215_U420 , P2_R1215_U419 , P2_R1215_U418 );
nand NAND2_16485 ( P2_R1215_U421 , P2_R1215_U153 , P2_R1215_U154 );
nand NAND2_16486 ( P2_R1215_U422 , P2_R1215_U300 , P2_R1215_U420 );
nand NAND2_16487 ( P2_R1215_U423 , P2_U3057 , P2_R1215_U49 );
nand NAND2_16488 ( P2_R1215_U424 , P2_U3970 , P2_R1215_U48 );
nand NAND2_16489 ( P2_R1215_U425 , P2_U3058 , P2_R1215_U50 );
nand NAND2_16490 ( P2_R1215_U426 , P2_U3971 , P2_R1215_U51 );
nand NAND2_16491 ( P2_R1215_U427 , P2_R1215_U426 , P2_R1215_U425 );
nand NAND2_16492 ( P2_R1215_U428 , P2_R1215_U357 , P2_R1215_U89 );
nand NAND2_16493 ( P2_R1215_U429 , P2_R1215_U427 , P2_R1215_U307 );
nand NAND2_16494 ( P2_R1215_U430 , P2_U3065 , P2_R1215_U52 );
nand NAND2_16495 ( P2_R1215_U431 , P2_U3972 , P2_R1215_U53 );
nand NAND2_16496 ( P2_R1215_U432 , P2_R1215_U431 , P2_R1215_U430 );
nand NAND2_16497 ( P2_R1215_U433 , P2_R1215_U358 , P2_R1215_U155 );
nand NAND2_16498 ( P2_R1215_U434 , P2_R1215_U294 , P2_R1215_U432 );
nand NAND2_16499 ( P2_R1215_U435 , P2_U3066 , P2_R1215_U84 );
nand NAND2_16500 ( P2_R1215_U436 , P2_U3973 , P2_R1215_U85 );
nand NAND2_16501 ( P2_R1215_U437 , P2_U3066 , P2_R1215_U84 );
nand NAND2_16502 ( P2_R1215_U438 , P2_U3973 , P2_R1215_U85 );
nand NAND2_16503 ( P2_R1215_U439 , P2_R1215_U438 , P2_R1215_U437 );
nand NAND2_16504 ( P2_R1215_U440 , P2_R1215_U156 , P2_R1215_U157 );
nand NAND2_16505 ( P2_R1215_U441 , P2_R1215_U290 , P2_R1215_U439 );
nand NAND2_16506 ( P2_R1215_U442 , P2_U3061 , P2_R1215_U82 );
nand NAND2_16507 ( P2_R1215_U443 , P2_U3974 , P2_R1215_U83 );
nand NAND2_16508 ( P2_R1215_U444 , P2_U3061 , P2_R1215_U82 );
nand NAND2_16509 ( P2_R1215_U445 , P2_U3974 , P2_R1215_U83 );
nand NAND2_16510 ( P2_R1215_U446 , P2_R1215_U445 , P2_R1215_U444 );
nand NAND2_16511 ( P2_R1215_U447 , P2_R1215_U158 , P2_R1215_U159 );
nand NAND2_16512 ( P2_R1215_U448 , P2_R1215_U286 , P2_R1215_U446 );
nand NAND2_16513 ( P2_R1215_U449 , P2_U3075 , P2_R1215_U54 );
nand NAND2_16514 ( P2_R1215_U450 , P2_U3975 , P2_R1215_U55 );
nand NAND2_16515 ( P2_R1215_U451 , P2_U3075 , P2_R1215_U54 );
nand NAND2_16516 ( P2_R1215_U452 , P2_U3975 , P2_R1215_U55 );
nand NAND2_16517 ( P2_R1215_U453 , P2_R1215_U452 , P2_R1215_U451 );
nand NAND2_16518 ( P2_R1215_U454 , P2_U3076 , P2_R1215_U81 );
nand NAND2_16519 ( P2_R1215_U455 , P2_U3976 , P2_R1215_U90 );
nand NAND2_16520 ( P2_R1215_U456 , P2_R1215_U182 , P2_R1215_U161 );
nand NAND2_16521 ( P2_R1215_U457 , P2_R1215_U328 , P2_R1215_U31 );
nand NAND2_16522 ( P2_R1215_U458 , P2_U3081 , P2_R1215_U78 );
nand NAND2_16523 ( P2_R1215_U459 , P2_U3506 , P2_R1215_U79 );
nand NAND2_16524 ( P2_R1215_U460 , P2_R1215_U459 , P2_R1215_U458 );
nand NAND2_16525 ( P2_R1215_U461 , P2_R1215_U359 , P2_R1215_U91 );
nand NAND2_16526 ( P2_R1215_U462 , P2_R1215_U460 , P2_R1215_U316 );
nand NAND2_16527 ( P2_R1215_U463 , P2_U3082 , P2_R1215_U75 );
nand NAND2_16528 ( P2_R1215_U464 , P2_U3504 , P2_R1215_U76 );
nand NAND2_16529 ( P2_R1215_U465 , P2_R1215_U464 , P2_R1215_U463 );
nand NAND2_16530 ( P2_R1215_U466 , P2_R1215_U360 , P2_R1215_U162 );
nand NAND2_16531 ( P2_R1215_U467 , P2_R1215_U270 , P2_R1215_U465 );
nand NAND2_16532 ( P2_R1215_U468 , P2_U3069 , P2_R1215_U60 );
nand NAND2_16533 ( P2_R1215_U469 , P2_U3501 , P2_R1215_U58 );
nand NAND2_16534 ( P2_R1215_U470 , P2_U3073 , P2_R1215_U56 );
nand NAND2_16535 ( P2_R1215_U471 , P2_U3498 , P2_R1215_U57 );
nand NAND2_16536 ( P2_R1215_U472 , P2_R1215_U471 , P2_R1215_U470 );
nand NAND2_16537 ( P2_R1215_U473 , P2_R1215_U361 , P2_R1215_U92 );
nand NAND2_16538 ( P2_R1215_U474 , P2_R1215_U472 , P2_R1215_U262 );
nand NAND2_16539 ( P2_R1215_U475 , P2_U3074 , P2_R1215_U73 );
nand NAND2_16540 ( P2_R1215_U476 , P2_U3495 , P2_R1215_U74 );
nand NAND2_16541 ( P2_R1215_U477 , P2_U3074 , P2_R1215_U73 );
nand NAND2_16542 ( P2_R1215_U478 , P2_U3495 , P2_R1215_U74 );
nand NAND2_16543 ( P2_R1215_U479 , P2_R1215_U478 , P2_R1215_U477 );
nand NAND2_16544 ( P2_R1215_U480 , P2_R1215_U163 , P2_R1215_U164 );
nand NAND2_16545 ( P2_R1215_U481 , P2_R1215_U258 , P2_R1215_U479 );
nand NAND2_16546 ( P2_R1215_U482 , P2_U3079 , P2_R1215_U71 );
nand NAND2_16547 ( P2_R1215_U483 , P2_U3492 , P2_R1215_U72 );
nand NAND2_16548 ( P2_R1215_U484 , P2_U3079 , P2_R1215_U71 );
nand NAND2_16549 ( P2_R1215_U485 , P2_U3492 , P2_R1215_U72 );
nand NAND2_16550 ( P2_R1215_U486 , P2_R1215_U485 , P2_R1215_U484 );
nand NAND2_16551 ( P2_R1215_U487 , P2_R1215_U165 , P2_R1215_U166 );
nand NAND2_16552 ( P2_R1215_U488 , P2_R1215_U254 , P2_R1215_U486 );
nand NAND2_16553 ( P2_R1215_U489 , P2_U3080 , P2_R1215_U69 );
nand NAND2_16554 ( P2_R1215_U490 , P2_U3489 , P2_R1215_U70 );
nand NAND2_16555 ( P2_R1215_U491 , P2_U3072 , P2_R1215_U64 );
nand NAND2_16556 ( P2_R1215_U492 , P2_U3486 , P2_R1215_U65 );
nand NAND2_16557 ( P2_R1215_U493 , P2_R1215_U492 , P2_R1215_U491 );
nand NAND2_16558 ( P2_R1215_U494 , P2_R1215_U362 , P2_R1215_U93 );
nand NAND2_16559 ( P2_R1215_U495 , P2_R1215_U493 , P2_R1215_U338 );
nand NAND2_16560 ( P2_R1215_U496 , P2_U3063 , P2_R1215_U66 );
nand NAND2_16561 ( P2_R1215_U497 , P2_U3483 , P2_R1215_U67 );
nand NAND2_16562 ( P2_R1215_U498 , P2_R1215_U497 , P2_R1215_U496 );
nand NAND2_16563 ( P2_R1215_U499 , P2_R1215_U363 , P2_R1215_U167 );
nand NAND2_16564 ( P2_R1215_U500 , P2_R1215_U244 , P2_R1215_U498 );
nand NAND2_16565 ( P2_R1215_U501 , P2_U3062 , P2_R1215_U62 );
nand NAND2_16566 ( P2_R1215_U502 , P2_U3480 , P2_R1215_U63 );
nand NAND2_16567 ( P2_R1215_U503 , P2_U3077 , P2_R1215_U29 );
nand NAND2_16568 ( P2_R1215_U504 , P2_U3448 , P2_R1215_U30 );
and AND2_16569 ( P2_R1164_U4 , P2_R1164_U179 , P2_R1164_U178 );
and AND2_16570 ( P2_R1164_U5 , P2_R1164_U197 , P2_R1164_U196 );
and AND2_16571 ( P2_R1164_U6 , P2_R1164_U237 , P2_R1164_U236 );
and AND2_16572 ( P2_R1164_U7 , P2_R1164_U246 , P2_R1164_U245 );
and AND2_16573 ( P2_R1164_U8 , P2_R1164_U264 , P2_R1164_U263 );
and AND2_16574 ( P2_R1164_U9 , P2_R1164_U272 , P2_R1164_U271 );
and AND2_16575 ( P2_R1164_U10 , P2_R1164_U351 , P2_R1164_U348 );
and AND2_16576 ( P2_R1164_U11 , P2_R1164_U344 , P2_R1164_U341 );
and AND2_16577 ( P2_R1164_U12 , P2_R1164_U335 , P2_R1164_U332 );
and AND2_16578 ( P2_R1164_U13 , P2_R1164_U326 , P2_R1164_U323 );
and AND2_16579 ( P2_R1164_U14 , P2_R1164_U320 , P2_R1164_U318 );
and AND2_16580 ( P2_R1164_U15 , P2_R1164_U313 , P2_R1164_U310 );
and AND2_16581 ( P2_R1164_U16 , P2_R1164_U235 , P2_R1164_U232 );
and AND2_16582 ( P2_R1164_U17 , P2_R1164_U227 , P2_R1164_U224 );
and AND2_16583 ( P2_R1164_U18 , P2_R1164_U213 , P2_R1164_U210 );
not NOT1_16584 ( P2_R1164_U19 , P2_U3468 );
not NOT1_16585 ( P2_R1164_U20 , P2_U3071 );
not NOT1_16586 ( P2_R1164_U21 , P2_U3070 );
nand NAND2_16587 ( P2_R1164_U22 , P2_U3071 , P2_U3468 );
not NOT1_16588 ( P2_R1164_U23 , P2_U3471 );
not NOT1_16589 ( P2_R1164_U24 , P2_U3462 );
not NOT1_16590 ( P2_R1164_U25 , P2_U3060 );
not NOT1_16591 ( P2_R1164_U26 , P2_U3067 );
not NOT1_16592 ( P2_R1164_U27 , P2_U3456 );
not NOT1_16593 ( P2_R1164_U28 , P2_U3068 );
not NOT1_16594 ( P2_R1164_U29 , P2_U3448 );
not NOT1_16595 ( P2_R1164_U30 , P2_U3077 );
nand NAND2_16596 ( P2_R1164_U31 , P2_U3077 , P2_U3448 );
not NOT1_16597 ( P2_R1164_U32 , P2_U3459 );
not NOT1_16598 ( P2_R1164_U33 , P2_U3064 );
nand NAND2_16599 ( P2_R1164_U34 , P2_U3060 , P2_U3462 );
not NOT1_16600 ( P2_R1164_U35 , P2_U3465 );
not NOT1_16601 ( P2_R1164_U36 , P2_U3474 );
not NOT1_16602 ( P2_R1164_U37 , P2_U3084 );
not NOT1_16603 ( P2_R1164_U38 , P2_U3083 );
not NOT1_16604 ( P2_R1164_U39 , P2_U3477 );
nand NAND2_16605 ( P2_R1164_U40 , P2_R1164_U63 , P2_R1164_U205 );
nand NAND2_16606 ( P2_R1164_U41 , P2_R1164_U117 , P2_R1164_U193 );
nand NAND2_16607 ( P2_R1164_U42 , P2_R1164_U182 , P2_R1164_U183 );
nand NAND2_16608 ( P2_R1164_U43 , P2_U3453 , P2_U3078 );
nand NAND2_16609 ( P2_R1164_U44 , P2_R1164_U122 , P2_R1164_U219 );
nand NAND2_16610 ( P2_R1164_U45 , P2_R1164_U216 , P2_R1164_U215 );
not NOT1_16611 ( P2_R1164_U46 , P2_U3969 );
not NOT1_16612 ( P2_R1164_U47 , P2_U3053 );
not NOT1_16613 ( P2_R1164_U48 , P2_U3057 );
not NOT1_16614 ( P2_R1164_U49 , P2_U3970 );
not NOT1_16615 ( P2_R1164_U50 , P2_U3971 );
not NOT1_16616 ( P2_R1164_U51 , P2_U3058 );
not NOT1_16617 ( P2_R1164_U52 , P2_U3972 );
not NOT1_16618 ( P2_R1164_U53 , P2_U3065 );
not NOT1_16619 ( P2_R1164_U54 , P2_U3975 );
not NOT1_16620 ( P2_R1164_U55 , P2_U3075 );
not NOT1_16621 ( P2_R1164_U56 , P2_U3498 );
not NOT1_16622 ( P2_R1164_U57 , P2_U3073 );
not NOT1_16623 ( P2_R1164_U58 , P2_U3069 );
nand NAND2_16624 ( P2_R1164_U59 , P2_U3073 , P2_U3498 );
not NOT1_16625 ( P2_R1164_U60 , P2_U3501 );
not NOT1_16626 ( P2_R1164_U61 , P2_U3480 );
not NOT1_16627 ( P2_R1164_U62 , P2_U3062 );
nand NAND2_16628 ( P2_R1164_U63 , P2_U3084 , P2_U3474 );
not NOT1_16629 ( P2_R1164_U64 , P2_U3486 );
not NOT1_16630 ( P2_R1164_U65 , P2_U3072 );
not NOT1_16631 ( P2_R1164_U66 , P2_U3483 );
not NOT1_16632 ( P2_R1164_U67 , P2_U3063 );
nand NAND2_16633 ( P2_R1164_U68 , P2_U3063 , P2_U3483 );
not NOT1_16634 ( P2_R1164_U69 , P2_U3489 );
not NOT1_16635 ( P2_R1164_U70 , P2_U3080 );
not NOT1_16636 ( P2_R1164_U71 , P2_U3492 );
not NOT1_16637 ( P2_R1164_U72 , P2_U3079 );
not NOT1_16638 ( P2_R1164_U73 , P2_U3495 );
not NOT1_16639 ( P2_R1164_U74 , P2_U3074 );
not NOT1_16640 ( P2_R1164_U75 , P2_U3504 );
not NOT1_16641 ( P2_R1164_U76 , P2_U3082 );
nand NAND2_16642 ( P2_R1164_U77 , P2_U3082 , P2_U3504 );
not NOT1_16643 ( P2_R1164_U78 , P2_U3506 );
not NOT1_16644 ( P2_R1164_U79 , P2_U3081 );
nand NAND2_16645 ( P2_R1164_U80 , P2_U3081 , P2_U3506 );
not NOT1_16646 ( P2_R1164_U81 , P2_U3976 );
not NOT1_16647 ( P2_R1164_U82 , P2_U3974 );
not NOT1_16648 ( P2_R1164_U83 , P2_U3061 );
not NOT1_16649 ( P2_R1164_U84 , P2_U3973 );
not NOT1_16650 ( P2_R1164_U85 , P2_U3066 );
nand NAND2_16651 ( P2_R1164_U86 , P2_U3970 , P2_U3057 );
not NOT1_16652 ( P2_R1164_U87 , P2_U3054 );
not NOT1_16653 ( P2_R1164_U88 , P2_U3968 );
nand NAND2_16654 ( P2_R1164_U89 , P2_R1164_U306 , P2_R1164_U176 );
not NOT1_16655 ( P2_R1164_U90 , P2_U3076 );
nand NAND2_16656 ( P2_R1164_U91 , P2_R1164_U77 , P2_R1164_U315 );
nand NAND2_16657 ( P2_R1164_U92 , P2_R1164_U261 , P2_R1164_U260 );
nand NAND2_16658 ( P2_R1164_U93 , P2_R1164_U68 , P2_R1164_U337 );
nand NAND2_16659 ( P2_R1164_U94 , P2_R1164_U457 , P2_R1164_U456 );
nand NAND2_16660 ( P2_R1164_U95 , P2_R1164_U504 , P2_R1164_U503 );
nand NAND2_16661 ( P2_R1164_U96 , P2_R1164_U375 , P2_R1164_U374 );
nand NAND2_16662 ( P2_R1164_U97 , P2_R1164_U380 , P2_R1164_U379 );
nand NAND2_16663 ( P2_R1164_U98 , P2_R1164_U387 , P2_R1164_U386 );
nand NAND2_16664 ( P2_R1164_U99 , P2_R1164_U394 , P2_R1164_U393 );
nand NAND2_16665 ( P2_R1164_U100 , P2_R1164_U399 , P2_R1164_U398 );
nand NAND2_16666 ( P2_R1164_U101 , P2_R1164_U408 , P2_R1164_U407 );
nand NAND2_16667 ( P2_R1164_U102 , P2_R1164_U415 , P2_R1164_U414 );
nand NAND2_16668 ( P2_R1164_U103 , P2_R1164_U422 , P2_R1164_U421 );
nand NAND2_16669 ( P2_R1164_U104 , P2_R1164_U429 , P2_R1164_U428 );
nand NAND2_16670 ( P2_R1164_U105 , P2_R1164_U434 , P2_R1164_U433 );
nand NAND2_16671 ( P2_R1164_U106 , P2_R1164_U441 , P2_R1164_U440 );
nand NAND2_16672 ( P2_R1164_U107 , P2_R1164_U448 , P2_R1164_U447 );
nand NAND2_16673 ( P2_R1164_U108 , P2_R1164_U462 , P2_R1164_U461 );
nand NAND2_16674 ( P2_R1164_U109 , P2_R1164_U467 , P2_R1164_U466 );
nand NAND2_16675 ( P2_R1164_U110 , P2_R1164_U474 , P2_R1164_U473 );
nand NAND2_16676 ( P2_R1164_U111 , P2_R1164_U481 , P2_R1164_U480 );
nand NAND2_16677 ( P2_R1164_U112 , P2_R1164_U488 , P2_R1164_U487 );
nand NAND2_16678 ( P2_R1164_U113 , P2_R1164_U495 , P2_R1164_U494 );
nand NAND2_16679 ( P2_R1164_U114 , P2_R1164_U500 , P2_R1164_U499 );
and AND2_16680 ( P2_R1164_U115 , P2_R1164_U189 , P2_R1164_U187 );
and AND2_16681 ( P2_R1164_U116 , P2_R1164_U4 , P2_R1164_U180 );
and AND2_16682 ( P2_R1164_U117 , P2_R1164_U194 , P2_R1164_U192 );
and AND2_16683 ( P2_R1164_U118 , P2_R1164_U201 , P2_R1164_U200 );
and AND3_16684 ( P2_R1164_U119 , P2_R1164_U382 , P2_R1164_U381 , P2_R1164_U22 );
and AND2_16685 ( P2_R1164_U120 , P2_R1164_U212 , P2_R1164_U5 );
and AND2_16686 ( P2_R1164_U121 , P2_R1164_U181 , P2_R1164_U180 );
and AND2_16687 ( P2_R1164_U122 , P2_R1164_U220 , P2_R1164_U218 );
and AND3_16688 ( P2_R1164_U123 , P2_R1164_U389 , P2_R1164_U388 , P2_R1164_U34 );
and AND2_16689 ( P2_R1164_U124 , P2_R1164_U226 , P2_R1164_U4 );
and AND2_16690 ( P2_R1164_U125 , P2_R1164_U234 , P2_R1164_U181 );
and AND2_16691 ( P2_R1164_U126 , P2_R1164_U204 , P2_R1164_U6 );
and AND2_16692 ( P2_R1164_U127 , P2_R1164_U243 , P2_R1164_U239 );
and AND2_16693 ( P2_R1164_U128 , P2_R1164_U250 , P2_R1164_U7 );
and AND2_16694 ( P2_R1164_U129 , P2_R1164_U248 , P2_R1164_U172 );
and AND2_16695 ( P2_R1164_U130 , P2_R1164_U268 , P2_R1164_U267 );
and AND3_16696 ( P2_R1164_U131 , P2_R1164_U9 , P2_R1164_U282 , P2_R1164_U273 );
and AND2_16697 ( P2_R1164_U132 , P2_R1164_U285 , P2_R1164_U280 );
and AND2_16698 ( P2_R1164_U133 , P2_R1164_U301 , P2_R1164_U298 );
and AND2_16699 ( P2_R1164_U134 , P2_R1164_U368 , P2_R1164_U302 );
and AND3_16700 ( P2_R1164_U135 , P2_R1164_U424 , P2_R1164_U423 , P2_R1164_U173 );
and AND2_16701 ( P2_R1164_U136 , P2_R1164_U160 , P2_R1164_U278 );
and AND3_16702 ( P2_R1164_U137 , P2_R1164_U455 , P2_R1164_U454 , P2_R1164_U80 );
and AND2_16703 ( P2_R1164_U138 , P2_R1164_U325 , P2_R1164_U9 );
and AND3_16704 ( P2_R1164_U139 , P2_R1164_U469 , P2_R1164_U468 , P2_R1164_U59 );
and AND2_16705 ( P2_R1164_U140 , P2_R1164_U334 , P2_R1164_U8 );
and AND3_16706 ( P2_R1164_U141 , P2_R1164_U490 , P2_R1164_U489 , P2_R1164_U172 );
and AND2_16707 ( P2_R1164_U142 , P2_R1164_U343 , P2_R1164_U7 );
and AND3_16708 ( P2_R1164_U143 , P2_R1164_U502 , P2_R1164_U501 , P2_R1164_U171 );
and AND2_16709 ( P2_R1164_U144 , P2_R1164_U350 , P2_R1164_U6 );
nand NAND2_16710 ( P2_R1164_U145 , P2_R1164_U118 , P2_R1164_U202 );
nand NAND2_16711 ( P2_R1164_U146 , P2_R1164_U217 , P2_R1164_U229 );
not NOT1_16712 ( P2_R1164_U147 , P2_U3055 );
not NOT1_16713 ( P2_R1164_U148 , P2_U3979 );
and AND2_16714 ( P2_R1164_U149 , P2_R1164_U403 , P2_R1164_U402 );
nand NAND3_16715 ( P2_R1164_U150 , P2_R1164_U304 , P2_R1164_U169 , P2_R1164_U364 );
and AND2_16716 ( P2_R1164_U151 , P2_R1164_U410 , P2_R1164_U409 );
nand NAND3_16717 ( P2_R1164_U152 , P2_R1164_U370 , P2_R1164_U369 , P2_R1164_U134 );
and AND2_16718 ( P2_R1164_U153 , P2_R1164_U417 , P2_R1164_U416 );
nand NAND3_16719 ( P2_R1164_U154 , P2_R1164_U365 , P2_R1164_U299 , P2_R1164_U86 );
nand NAND2_16720 ( P2_R1164_U155 , P2_R1164_U293 , P2_R1164_U292 );
and AND2_16721 ( P2_R1164_U156 , P2_R1164_U436 , P2_R1164_U435 );
nand NAND2_16722 ( P2_R1164_U157 , P2_R1164_U289 , P2_R1164_U288 );
and AND2_16723 ( P2_R1164_U158 , P2_R1164_U443 , P2_R1164_U442 );
nand NAND2_16724 ( P2_R1164_U159 , P2_R1164_U132 , P2_R1164_U284 );
and AND2_16725 ( P2_R1164_U160 , P2_R1164_U450 , P2_R1164_U449 );
nand NAND2_16726 ( P2_R1164_U161 , P2_R1164_U43 , P2_R1164_U327 );
nand NAND2_16727 ( P2_R1164_U162 , P2_R1164_U130 , P2_R1164_U269 );
and AND2_16728 ( P2_R1164_U163 , P2_R1164_U476 , P2_R1164_U475 );
nand NAND2_16729 ( P2_R1164_U164 , P2_R1164_U257 , P2_R1164_U256 );
and AND2_16730 ( P2_R1164_U165 , P2_R1164_U483 , P2_R1164_U482 );
nand NAND2_16731 ( P2_R1164_U166 , P2_R1164_U253 , P2_R1164_U252 );
nand NAND2_16732 ( P2_R1164_U167 , P2_R1164_U127 , P2_R1164_U242 );
nand NAND2_16733 ( P2_R1164_U168 , P2_R1164_U367 , P2_R1164_U366 );
nand NAND2_16734 ( P2_R1164_U169 , P2_U3054 , P2_R1164_U152 );
not NOT1_16735 ( P2_R1164_U170 , P2_R1164_U34 );
nand NAND2_16736 ( P2_R1164_U171 , P2_U3477 , P2_U3083 );
nand NAND2_16737 ( P2_R1164_U172 , P2_U3072 , P2_U3486 );
nand NAND2_16738 ( P2_R1164_U173 , P2_U3058 , P2_U3971 );
not NOT1_16739 ( P2_R1164_U174 , P2_R1164_U68 );
not NOT1_16740 ( P2_R1164_U175 , P2_R1164_U77 );
nand NAND2_16741 ( P2_R1164_U176 , P2_U3065 , P2_U3972 );
not NOT1_16742 ( P2_R1164_U177 , P2_R1164_U63 );
or OR2_16743 ( P2_R1164_U178 , P2_U3067 , P2_U3465 );
or OR2_16744 ( P2_R1164_U179 , P2_U3060 , P2_U3462 );
or OR2_16745 ( P2_R1164_U180 , P2_U3459 , P2_U3064 );
or OR2_16746 ( P2_R1164_U181 , P2_U3456 , P2_U3068 );
not NOT1_16747 ( P2_R1164_U182 , P2_R1164_U31 );
or OR2_16748 ( P2_R1164_U183 , P2_U3453 , P2_U3078 );
not NOT1_16749 ( P2_R1164_U184 , P2_R1164_U42 );
not NOT1_16750 ( P2_R1164_U185 , P2_R1164_U43 );
nand NAND2_16751 ( P2_R1164_U186 , P2_R1164_U42 , P2_R1164_U43 );
nand NAND2_16752 ( P2_R1164_U187 , P2_U3068 , P2_U3456 );
nand NAND2_16753 ( P2_R1164_U188 , P2_R1164_U186 , P2_R1164_U181 );
nand NAND2_16754 ( P2_R1164_U189 , P2_U3064 , P2_U3459 );
nand NAND2_16755 ( P2_R1164_U190 , P2_R1164_U115 , P2_R1164_U188 );
nand NAND2_16756 ( P2_R1164_U191 , P2_R1164_U35 , P2_R1164_U34 );
nand NAND2_16757 ( P2_R1164_U192 , P2_U3067 , P2_R1164_U191 );
nand NAND2_16758 ( P2_R1164_U193 , P2_R1164_U116 , P2_R1164_U190 );
nand NAND2_16759 ( P2_R1164_U194 , P2_U3465 , P2_R1164_U170 );
not NOT1_16760 ( P2_R1164_U195 , P2_R1164_U41 );
or OR2_16761 ( P2_R1164_U196 , P2_U3070 , P2_U3471 );
or OR2_16762 ( P2_R1164_U197 , P2_U3071 , P2_U3468 );
not NOT1_16763 ( P2_R1164_U198 , P2_R1164_U22 );
nand NAND2_16764 ( P2_R1164_U199 , P2_R1164_U23 , P2_R1164_U22 );
nand NAND2_16765 ( P2_R1164_U200 , P2_U3070 , P2_R1164_U199 );
nand NAND2_16766 ( P2_R1164_U201 , P2_U3471 , P2_R1164_U198 );
nand NAND2_16767 ( P2_R1164_U202 , P2_R1164_U5 , P2_R1164_U41 );
not NOT1_16768 ( P2_R1164_U203 , P2_R1164_U145 );
or OR2_16769 ( P2_R1164_U204 , P2_U3474 , P2_U3084 );
nand NAND2_16770 ( P2_R1164_U205 , P2_R1164_U204 , P2_R1164_U145 );
not NOT1_16771 ( P2_R1164_U206 , P2_R1164_U40 );
or OR2_16772 ( P2_R1164_U207 , P2_U3083 , P2_U3477 );
or OR2_16773 ( P2_R1164_U208 , P2_U3468 , P2_U3071 );
nand NAND2_16774 ( P2_R1164_U209 , P2_R1164_U208 , P2_R1164_U41 );
nand NAND2_16775 ( P2_R1164_U210 , P2_R1164_U119 , P2_R1164_U209 );
nand NAND2_16776 ( P2_R1164_U211 , P2_R1164_U195 , P2_R1164_U22 );
nand NAND2_16777 ( P2_R1164_U212 , P2_U3471 , P2_U3070 );
nand NAND2_16778 ( P2_R1164_U213 , P2_R1164_U120 , P2_R1164_U211 );
or OR2_16779 ( P2_R1164_U214 , P2_U3071 , P2_U3468 );
nand NAND2_16780 ( P2_R1164_U215 , P2_R1164_U185 , P2_R1164_U181 );
nand NAND2_16781 ( P2_R1164_U216 , P2_U3068 , P2_U3456 );
not NOT1_16782 ( P2_R1164_U217 , P2_R1164_U45 );
nand NAND2_16783 ( P2_R1164_U218 , P2_R1164_U121 , P2_R1164_U184 );
nand NAND2_16784 ( P2_R1164_U219 , P2_R1164_U45 , P2_R1164_U180 );
nand NAND2_16785 ( P2_R1164_U220 , P2_U3064 , P2_U3459 );
not NOT1_16786 ( P2_R1164_U221 , P2_R1164_U44 );
or OR2_16787 ( P2_R1164_U222 , P2_U3462 , P2_U3060 );
nand NAND2_16788 ( P2_R1164_U223 , P2_R1164_U222 , P2_R1164_U44 );
nand NAND2_16789 ( P2_R1164_U224 , P2_R1164_U123 , P2_R1164_U223 );
nand NAND2_16790 ( P2_R1164_U225 , P2_R1164_U221 , P2_R1164_U34 );
nand NAND2_16791 ( P2_R1164_U226 , P2_U3465 , P2_U3067 );
nand NAND2_16792 ( P2_R1164_U227 , P2_R1164_U124 , P2_R1164_U225 );
or OR2_16793 ( P2_R1164_U228 , P2_U3060 , P2_U3462 );
nand NAND2_16794 ( P2_R1164_U229 , P2_R1164_U184 , P2_R1164_U181 );
not NOT1_16795 ( P2_R1164_U230 , P2_R1164_U146 );
nand NAND2_16796 ( P2_R1164_U231 , P2_U3064 , P2_U3459 );
nand NAND4_16797 ( P2_R1164_U232 , P2_R1164_U401 , P2_R1164_U400 , P2_R1164_U43 , P2_R1164_U42 );
nand NAND2_16798 ( P2_R1164_U233 , P2_R1164_U43 , P2_R1164_U42 );
nand NAND2_16799 ( P2_R1164_U234 , P2_U3068 , P2_U3456 );
nand NAND2_16800 ( P2_R1164_U235 , P2_R1164_U125 , P2_R1164_U233 );
or OR2_16801 ( P2_R1164_U236 , P2_U3083 , P2_U3477 );
or OR2_16802 ( P2_R1164_U237 , P2_U3062 , P2_U3480 );
nand NAND2_16803 ( P2_R1164_U238 , P2_R1164_U177 , P2_R1164_U6 );
nand NAND2_16804 ( P2_R1164_U239 , P2_U3062 , P2_U3480 );
nand NAND2_16805 ( P2_R1164_U240 , P2_R1164_U171 , P2_R1164_U238 );
or OR2_16806 ( P2_R1164_U241 , P2_U3480 , P2_U3062 );
nand NAND2_16807 ( P2_R1164_U242 , P2_R1164_U126 , P2_R1164_U145 );
nand NAND2_16808 ( P2_R1164_U243 , P2_R1164_U241 , P2_R1164_U240 );
not NOT1_16809 ( P2_R1164_U244 , P2_R1164_U167 );
or OR2_16810 ( P2_R1164_U245 , P2_U3080 , P2_U3489 );
or OR2_16811 ( P2_R1164_U246 , P2_U3072 , P2_U3486 );
nand NAND2_16812 ( P2_R1164_U247 , P2_R1164_U174 , P2_R1164_U7 );
nand NAND2_16813 ( P2_R1164_U248 , P2_U3080 , P2_U3489 );
nand NAND2_16814 ( P2_R1164_U249 , P2_R1164_U129 , P2_R1164_U247 );
or OR2_16815 ( P2_R1164_U250 , P2_U3483 , P2_U3063 );
or OR2_16816 ( P2_R1164_U251 , P2_U3489 , P2_U3080 );
nand NAND2_16817 ( P2_R1164_U252 , P2_R1164_U128 , P2_R1164_U167 );
nand NAND2_16818 ( P2_R1164_U253 , P2_R1164_U251 , P2_R1164_U249 );
not NOT1_16819 ( P2_R1164_U254 , P2_R1164_U166 );
or OR2_16820 ( P2_R1164_U255 , P2_U3492 , P2_U3079 );
nand NAND2_16821 ( P2_R1164_U256 , P2_R1164_U255 , P2_R1164_U166 );
nand NAND2_16822 ( P2_R1164_U257 , P2_U3079 , P2_U3492 );
not NOT1_16823 ( P2_R1164_U258 , P2_R1164_U164 );
or OR2_16824 ( P2_R1164_U259 , P2_U3495 , P2_U3074 );
nand NAND2_16825 ( P2_R1164_U260 , P2_R1164_U259 , P2_R1164_U164 );
nand NAND2_16826 ( P2_R1164_U261 , P2_U3074 , P2_U3495 );
not NOT1_16827 ( P2_R1164_U262 , P2_R1164_U92 );
or OR2_16828 ( P2_R1164_U263 , P2_U3069 , P2_U3501 );
or OR2_16829 ( P2_R1164_U264 , P2_U3073 , P2_U3498 );
not NOT1_16830 ( P2_R1164_U265 , P2_R1164_U59 );
nand NAND2_16831 ( P2_R1164_U266 , P2_R1164_U60 , P2_R1164_U59 );
nand NAND2_16832 ( P2_R1164_U267 , P2_U3069 , P2_R1164_U266 );
nand NAND2_16833 ( P2_R1164_U268 , P2_U3501 , P2_R1164_U265 );
nand NAND2_16834 ( P2_R1164_U269 , P2_R1164_U8 , P2_R1164_U92 );
not NOT1_16835 ( P2_R1164_U270 , P2_R1164_U162 );
or OR2_16836 ( P2_R1164_U271 , P2_U3076 , P2_U3976 );
or OR2_16837 ( P2_R1164_U272 , P2_U3081 , P2_U3506 );
or OR2_16838 ( P2_R1164_U273 , P2_U3075 , P2_U3975 );
not NOT1_16839 ( P2_R1164_U274 , P2_R1164_U80 );
nand NAND2_16840 ( P2_R1164_U275 , P2_U3976 , P2_R1164_U274 );
nand NAND2_16841 ( P2_R1164_U276 , P2_R1164_U275 , P2_R1164_U90 );
nand NAND2_16842 ( P2_R1164_U277 , P2_R1164_U80 , P2_R1164_U81 );
nand NAND2_16843 ( P2_R1164_U278 , P2_R1164_U277 , P2_R1164_U276 );
nand NAND2_16844 ( P2_R1164_U279 , P2_R1164_U175 , P2_R1164_U9 );
nand NAND2_16845 ( P2_R1164_U280 , P2_U3075 , P2_U3975 );
nand NAND2_16846 ( P2_R1164_U281 , P2_R1164_U278 , P2_R1164_U279 );
or OR2_16847 ( P2_R1164_U282 , P2_U3504 , P2_U3082 );
or OR2_16848 ( P2_R1164_U283 , P2_U3975 , P2_U3075 );
nand NAND2_16849 ( P2_R1164_U284 , P2_R1164_U162 , P2_R1164_U131 );
nand NAND2_16850 ( P2_R1164_U285 , P2_R1164_U283 , P2_R1164_U281 );
not NOT1_16851 ( P2_R1164_U286 , P2_R1164_U159 );
or OR2_16852 ( P2_R1164_U287 , P2_U3974 , P2_U3061 );
nand NAND2_16853 ( P2_R1164_U288 , P2_R1164_U287 , P2_R1164_U159 );
nand NAND2_16854 ( P2_R1164_U289 , P2_U3061 , P2_U3974 );
not NOT1_16855 ( P2_R1164_U290 , P2_R1164_U157 );
or OR2_16856 ( P2_R1164_U291 , P2_U3973 , P2_U3066 );
nand NAND2_16857 ( P2_R1164_U292 , P2_R1164_U291 , P2_R1164_U157 );
nand NAND2_16858 ( P2_R1164_U293 , P2_U3066 , P2_U3973 );
not NOT1_16859 ( P2_R1164_U294 , P2_R1164_U155 );
or OR2_16860 ( P2_R1164_U295 , P2_U3058 , P2_U3971 );
nand NAND2_16861 ( P2_R1164_U296 , P2_R1164_U176 , P2_R1164_U173 );
not NOT1_16862 ( P2_R1164_U297 , P2_R1164_U86 );
or OR2_16863 ( P2_R1164_U298 , P2_U3972 , P2_U3065 );
nand NAND3_16864 ( P2_R1164_U299 , P2_R1164_U155 , P2_R1164_U298 , P2_R1164_U168 );
not NOT1_16865 ( P2_R1164_U300 , P2_R1164_U154 );
or OR2_16866 ( P2_R1164_U301 , P2_U3969 , P2_U3053 );
nand NAND2_16867 ( P2_R1164_U302 , P2_U3053 , P2_U3969 );
not NOT1_16868 ( P2_R1164_U303 , P2_R1164_U152 );
nand NAND2_16869 ( P2_R1164_U304 , P2_U3968 , P2_R1164_U152 );
not NOT1_16870 ( P2_R1164_U305 , P2_R1164_U150 );
nand NAND2_16871 ( P2_R1164_U306 , P2_R1164_U298 , P2_R1164_U155 );
not NOT1_16872 ( P2_R1164_U307 , P2_R1164_U89 );
or OR2_16873 ( P2_R1164_U308 , P2_U3971 , P2_U3058 );
nand NAND2_16874 ( P2_R1164_U309 , P2_R1164_U308 , P2_R1164_U89 );
nand NAND2_16875 ( P2_R1164_U310 , P2_R1164_U135 , P2_R1164_U309 );
nand NAND2_16876 ( P2_R1164_U311 , P2_R1164_U307 , P2_R1164_U173 );
nand NAND2_16877 ( P2_R1164_U312 , P2_U3970 , P2_U3057 );
nand NAND3_16878 ( P2_R1164_U313 , P2_R1164_U311 , P2_R1164_U312 , P2_R1164_U168 );
or OR2_16879 ( P2_R1164_U314 , P2_U3058 , P2_U3971 );
nand NAND2_16880 ( P2_R1164_U315 , P2_R1164_U282 , P2_R1164_U162 );
not NOT1_16881 ( P2_R1164_U316 , P2_R1164_U91 );
nand NAND2_16882 ( P2_R1164_U317 , P2_R1164_U9 , P2_R1164_U91 );
nand NAND2_16883 ( P2_R1164_U318 , P2_R1164_U136 , P2_R1164_U317 );
nand NAND2_16884 ( P2_R1164_U319 , P2_R1164_U317 , P2_R1164_U278 );
nand NAND2_16885 ( P2_R1164_U320 , P2_R1164_U453 , P2_R1164_U319 );
or OR2_16886 ( P2_R1164_U321 , P2_U3506 , P2_U3081 );
nand NAND2_16887 ( P2_R1164_U322 , P2_R1164_U321 , P2_R1164_U91 );
nand NAND2_16888 ( P2_R1164_U323 , P2_R1164_U137 , P2_R1164_U322 );
nand NAND2_16889 ( P2_R1164_U324 , P2_R1164_U316 , P2_R1164_U80 );
nand NAND2_16890 ( P2_R1164_U325 , P2_U3076 , P2_U3976 );
nand NAND2_16891 ( P2_R1164_U326 , P2_R1164_U138 , P2_R1164_U324 );
or OR2_16892 ( P2_R1164_U327 , P2_U3453 , P2_U3078 );
not NOT1_16893 ( P2_R1164_U328 , P2_R1164_U161 );
or OR2_16894 ( P2_R1164_U329 , P2_U3081 , P2_U3506 );
or OR2_16895 ( P2_R1164_U330 , P2_U3498 , P2_U3073 );
nand NAND2_16896 ( P2_R1164_U331 , P2_R1164_U330 , P2_R1164_U92 );
nand NAND2_16897 ( P2_R1164_U332 , P2_R1164_U139 , P2_R1164_U331 );
nand NAND2_16898 ( P2_R1164_U333 , P2_R1164_U262 , P2_R1164_U59 );
nand NAND2_16899 ( P2_R1164_U334 , P2_U3501 , P2_U3069 );
nand NAND2_16900 ( P2_R1164_U335 , P2_R1164_U140 , P2_R1164_U333 );
or OR2_16901 ( P2_R1164_U336 , P2_U3073 , P2_U3498 );
nand NAND2_16902 ( P2_R1164_U337 , P2_R1164_U250 , P2_R1164_U167 );
not NOT1_16903 ( P2_R1164_U338 , P2_R1164_U93 );
or OR2_16904 ( P2_R1164_U339 , P2_U3486 , P2_U3072 );
nand NAND2_16905 ( P2_R1164_U340 , P2_R1164_U339 , P2_R1164_U93 );
nand NAND2_16906 ( P2_R1164_U341 , P2_R1164_U141 , P2_R1164_U340 );
nand NAND2_16907 ( P2_R1164_U342 , P2_R1164_U338 , P2_R1164_U172 );
nand NAND2_16908 ( P2_R1164_U343 , P2_U3080 , P2_U3489 );
nand NAND2_16909 ( P2_R1164_U344 , P2_R1164_U142 , P2_R1164_U342 );
or OR2_16910 ( P2_R1164_U345 , P2_U3072 , P2_U3486 );
or OR2_16911 ( P2_R1164_U346 , P2_U3477 , P2_U3083 );
nand NAND2_16912 ( P2_R1164_U347 , P2_R1164_U346 , P2_R1164_U40 );
nand NAND2_16913 ( P2_R1164_U348 , P2_R1164_U143 , P2_R1164_U347 );
nand NAND2_16914 ( P2_R1164_U349 , P2_R1164_U206 , P2_R1164_U171 );
nand NAND2_16915 ( P2_R1164_U350 , P2_U3062 , P2_U3480 );
nand NAND2_16916 ( P2_R1164_U351 , P2_R1164_U144 , P2_R1164_U349 );
nand NAND2_16917 ( P2_R1164_U352 , P2_R1164_U207 , P2_R1164_U171 );
nand NAND2_16918 ( P2_R1164_U353 , P2_R1164_U204 , P2_R1164_U63 );
nand NAND2_16919 ( P2_R1164_U354 , P2_R1164_U214 , P2_R1164_U22 );
nand NAND2_16920 ( P2_R1164_U355 , P2_R1164_U228 , P2_R1164_U34 );
nand NAND2_16921 ( P2_R1164_U356 , P2_R1164_U231 , P2_R1164_U180 );
nand NAND2_16922 ( P2_R1164_U357 , P2_R1164_U314 , P2_R1164_U173 );
nand NAND2_16923 ( P2_R1164_U358 , P2_R1164_U298 , P2_R1164_U176 );
nand NAND2_16924 ( P2_R1164_U359 , P2_R1164_U329 , P2_R1164_U80 );
nand NAND2_16925 ( P2_R1164_U360 , P2_R1164_U282 , P2_R1164_U77 );
nand NAND2_16926 ( P2_R1164_U361 , P2_R1164_U336 , P2_R1164_U59 );
nand NAND2_16927 ( P2_R1164_U362 , P2_R1164_U345 , P2_R1164_U172 );
nand NAND2_16928 ( P2_R1164_U363 , P2_R1164_U250 , P2_R1164_U68 );
nand NAND2_16929 ( P2_R1164_U364 , P2_U3968 , P2_U3054 );
nand NAND2_16930 ( P2_R1164_U365 , P2_R1164_U296 , P2_R1164_U168 );
nand NAND2_16931 ( P2_R1164_U366 , P2_U3057 , P2_R1164_U295 );
nand NAND2_16932 ( P2_R1164_U367 , P2_U3970 , P2_R1164_U295 );
nand NAND3_16933 ( P2_R1164_U368 , P2_R1164_U296 , P2_R1164_U168 , P2_R1164_U301 );
nand NAND3_16934 ( P2_R1164_U369 , P2_R1164_U155 , P2_R1164_U168 , P2_R1164_U133 );
nand NAND2_16935 ( P2_R1164_U370 , P2_R1164_U297 , P2_R1164_U301 );
nand NAND2_16936 ( P2_R1164_U371 , P2_U3083 , P2_R1164_U39 );
nand NAND2_16937 ( P2_R1164_U372 , P2_U3477 , P2_R1164_U38 );
nand NAND2_16938 ( P2_R1164_U373 , P2_R1164_U372 , P2_R1164_U371 );
nand NAND2_16939 ( P2_R1164_U374 , P2_R1164_U352 , P2_R1164_U40 );
nand NAND2_16940 ( P2_R1164_U375 , P2_R1164_U373 , P2_R1164_U206 );
nand NAND2_16941 ( P2_R1164_U376 , P2_U3084 , P2_R1164_U36 );
nand NAND2_16942 ( P2_R1164_U377 , P2_U3474 , P2_R1164_U37 );
nand NAND2_16943 ( P2_R1164_U378 , P2_R1164_U377 , P2_R1164_U376 );
nand NAND2_16944 ( P2_R1164_U379 , P2_R1164_U353 , P2_R1164_U145 );
nand NAND2_16945 ( P2_R1164_U380 , P2_R1164_U203 , P2_R1164_U378 );
nand NAND2_16946 ( P2_R1164_U381 , P2_U3070 , P2_R1164_U23 );
nand NAND2_16947 ( P2_R1164_U382 , P2_U3471 , P2_R1164_U21 );
nand NAND2_16948 ( P2_R1164_U383 , P2_U3071 , P2_R1164_U19 );
nand NAND2_16949 ( P2_R1164_U384 , P2_U3468 , P2_R1164_U20 );
nand NAND2_16950 ( P2_R1164_U385 , P2_R1164_U384 , P2_R1164_U383 );
nand NAND2_16951 ( P2_R1164_U386 , P2_R1164_U354 , P2_R1164_U41 );
nand NAND2_16952 ( P2_R1164_U387 , P2_R1164_U385 , P2_R1164_U195 );
nand NAND2_16953 ( P2_R1164_U388 , P2_U3067 , P2_R1164_U35 );
nand NAND2_16954 ( P2_R1164_U389 , P2_U3465 , P2_R1164_U26 );
nand NAND2_16955 ( P2_R1164_U390 , P2_U3060 , P2_R1164_U24 );
nand NAND2_16956 ( P2_R1164_U391 , P2_U3462 , P2_R1164_U25 );
nand NAND2_16957 ( P2_R1164_U392 , P2_R1164_U391 , P2_R1164_U390 );
nand NAND2_16958 ( P2_R1164_U393 , P2_R1164_U355 , P2_R1164_U44 );
nand NAND2_16959 ( P2_R1164_U394 , P2_R1164_U392 , P2_R1164_U221 );
nand NAND2_16960 ( P2_R1164_U395 , P2_U3064 , P2_R1164_U32 );
nand NAND2_16961 ( P2_R1164_U396 , P2_U3459 , P2_R1164_U33 );
nand NAND2_16962 ( P2_R1164_U397 , P2_R1164_U396 , P2_R1164_U395 );
nand NAND2_16963 ( P2_R1164_U398 , P2_R1164_U356 , P2_R1164_U146 );
nand NAND2_16964 ( P2_R1164_U399 , P2_R1164_U230 , P2_R1164_U397 );
nand NAND2_16965 ( P2_R1164_U400 , P2_U3068 , P2_R1164_U27 );
nand NAND2_16966 ( P2_R1164_U401 , P2_U3456 , P2_R1164_U28 );
nand NAND2_16967 ( P2_R1164_U402 , P2_U3055 , P2_R1164_U148 );
nand NAND2_16968 ( P2_R1164_U403 , P2_U3979 , P2_R1164_U147 );
nand NAND2_16969 ( P2_R1164_U404 , P2_U3055 , P2_R1164_U148 );
nand NAND2_16970 ( P2_R1164_U405 , P2_U3979 , P2_R1164_U147 );
nand NAND2_16971 ( P2_R1164_U406 , P2_R1164_U405 , P2_R1164_U404 );
nand NAND2_16972 ( P2_R1164_U407 , P2_R1164_U149 , P2_R1164_U150 );
nand NAND2_16973 ( P2_R1164_U408 , P2_R1164_U305 , P2_R1164_U406 );
nand NAND2_16974 ( P2_R1164_U409 , P2_U3054 , P2_R1164_U88 );
nand NAND2_16975 ( P2_R1164_U410 , P2_U3968 , P2_R1164_U87 );
nand NAND2_16976 ( P2_R1164_U411 , P2_U3054 , P2_R1164_U88 );
nand NAND2_16977 ( P2_R1164_U412 , P2_U3968 , P2_R1164_U87 );
nand NAND2_16978 ( P2_R1164_U413 , P2_R1164_U412 , P2_R1164_U411 );
nand NAND2_16979 ( P2_R1164_U414 , P2_R1164_U151 , P2_R1164_U152 );
nand NAND2_16980 ( P2_R1164_U415 , P2_R1164_U303 , P2_R1164_U413 );
nand NAND2_16981 ( P2_R1164_U416 , P2_U3053 , P2_R1164_U46 );
nand NAND2_16982 ( P2_R1164_U417 , P2_U3969 , P2_R1164_U47 );
nand NAND2_16983 ( P2_R1164_U418 , P2_U3053 , P2_R1164_U46 );
nand NAND2_16984 ( P2_R1164_U419 , P2_U3969 , P2_R1164_U47 );
nand NAND2_16985 ( P2_R1164_U420 , P2_R1164_U419 , P2_R1164_U418 );
nand NAND2_16986 ( P2_R1164_U421 , P2_R1164_U153 , P2_R1164_U154 );
nand NAND2_16987 ( P2_R1164_U422 , P2_R1164_U300 , P2_R1164_U420 );
nand NAND2_16988 ( P2_R1164_U423 , P2_U3057 , P2_R1164_U49 );
nand NAND2_16989 ( P2_R1164_U424 , P2_U3970 , P2_R1164_U48 );
nand NAND2_16990 ( P2_R1164_U425 , P2_U3058 , P2_R1164_U50 );
nand NAND2_16991 ( P2_R1164_U426 , P2_U3971 , P2_R1164_U51 );
nand NAND2_16992 ( P2_R1164_U427 , P2_R1164_U426 , P2_R1164_U425 );
nand NAND2_16993 ( P2_R1164_U428 , P2_R1164_U357 , P2_R1164_U89 );
nand NAND2_16994 ( P2_R1164_U429 , P2_R1164_U427 , P2_R1164_U307 );
nand NAND2_16995 ( P2_R1164_U430 , P2_U3065 , P2_R1164_U52 );
nand NAND2_16996 ( P2_R1164_U431 , P2_U3972 , P2_R1164_U53 );
nand NAND2_16997 ( P2_R1164_U432 , P2_R1164_U431 , P2_R1164_U430 );
nand NAND2_16998 ( P2_R1164_U433 , P2_R1164_U358 , P2_R1164_U155 );
nand NAND2_16999 ( P2_R1164_U434 , P2_R1164_U294 , P2_R1164_U432 );
nand NAND2_17000 ( P2_R1164_U435 , P2_U3066 , P2_R1164_U84 );
nand NAND2_17001 ( P2_R1164_U436 , P2_U3973 , P2_R1164_U85 );
nand NAND2_17002 ( P2_R1164_U437 , P2_U3066 , P2_R1164_U84 );
nand NAND2_17003 ( P2_R1164_U438 , P2_U3973 , P2_R1164_U85 );
nand NAND2_17004 ( P2_R1164_U439 , P2_R1164_U438 , P2_R1164_U437 );
nand NAND2_17005 ( P2_R1164_U440 , P2_R1164_U156 , P2_R1164_U157 );
nand NAND2_17006 ( P2_R1164_U441 , P2_R1164_U290 , P2_R1164_U439 );
nand NAND2_17007 ( P2_R1164_U442 , P2_U3061 , P2_R1164_U82 );
nand NAND2_17008 ( P2_R1164_U443 , P2_U3974 , P2_R1164_U83 );
nand NAND2_17009 ( P2_R1164_U444 , P2_U3061 , P2_R1164_U82 );
nand NAND2_17010 ( P2_R1164_U445 , P2_U3974 , P2_R1164_U83 );
nand NAND2_17011 ( P2_R1164_U446 , P2_R1164_U445 , P2_R1164_U444 );
nand NAND2_17012 ( P2_R1164_U447 , P2_R1164_U158 , P2_R1164_U159 );
nand NAND2_17013 ( P2_R1164_U448 , P2_R1164_U286 , P2_R1164_U446 );
nand NAND2_17014 ( P2_R1164_U449 , P2_U3075 , P2_R1164_U54 );
nand NAND2_17015 ( P2_R1164_U450 , P2_U3975 , P2_R1164_U55 );
nand NAND2_17016 ( P2_R1164_U451 , P2_U3075 , P2_R1164_U54 );
nand NAND2_17017 ( P2_R1164_U452 , P2_U3975 , P2_R1164_U55 );
nand NAND2_17018 ( P2_R1164_U453 , P2_R1164_U452 , P2_R1164_U451 );
nand NAND2_17019 ( P2_R1164_U454 , P2_U3076 , P2_R1164_U81 );
nand NAND2_17020 ( P2_R1164_U455 , P2_U3976 , P2_R1164_U90 );
nand NAND2_17021 ( P2_R1164_U456 , P2_R1164_U182 , P2_R1164_U161 );
nand NAND2_17022 ( P2_R1164_U457 , P2_R1164_U328 , P2_R1164_U31 );
nand NAND2_17023 ( P2_R1164_U458 , P2_U3081 , P2_R1164_U78 );
nand NAND2_17024 ( P2_R1164_U459 , P2_U3506 , P2_R1164_U79 );
nand NAND2_17025 ( P2_R1164_U460 , P2_R1164_U459 , P2_R1164_U458 );
nand NAND2_17026 ( P2_R1164_U461 , P2_R1164_U359 , P2_R1164_U91 );
nand NAND2_17027 ( P2_R1164_U462 , P2_R1164_U460 , P2_R1164_U316 );
nand NAND2_17028 ( P2_R1164_U463 , P2_U3082 , P2_R1164_U75 );
nand NAND2_17029 ( P2_R1164_U464 , P2_U3504 , P2_R1164_U76 );
nand NAND2_17030 ( P2_R1164_U465 , P2_R1164_U464 , P2_R1164_U463 );
nand NAND2_17031 ( P2_R1164_U466 , P2_R1164_U360 , P2_R1164_U162 );
nand NAND2_17032 ( P2_R1164_U467 , P2_R1164_U270 , P2_R1164_U465 );
nand NAND2_17033 ( P2_R1164_U468 , P2_U3069 , P2_R1164_U60 );
nand NAND2_17034 ( P2_R1164_U469 , P2_U3501 , P2_R1164_U58 );
nand NAND2_17035 ( P2_R1164_U470 , P2_U3073 , P2_R1164_U56 );
nand NAND2_17036 ( P2_R1164_U471 , P2_U3498 , P2_R1164_U57 );
nand NAND2_17037 ( P2_R1164_U472 , P2_R1164_U471 , P2_R1164_U470 );
nand NAND2_17038 ( P2_R1164_U473 , P2_R1164_U361 , P2_R1164_U92 );
nand NAND2_17039 ( P2_R1164_U474 , P2_R1164_U472 , P2_R1164_U262 );
nand NAND2_17040 ( P2_R1164_U475 , P2_U3074 , P2_R1164_U73 );
nand NAND2_17041 ( P2_R1164_U476 , P2_U3495 , P2_R1164_U74 );
nand NAND2_17042 ( P2_R1164_U477 , P2_U3074 , P2_R1164_U73 );
nand NAND2_17043 ( P2_R1164_U478 , P2_U3495 , P2_R1164_U74 );
nand NAND2_17044 ( P2_R1164_U479 , P2_R1164_U478 , P2_R1164_U477 );
nand NAND2_17045 ( P2_R1164_U480 , P2_R1164_U163 , P2_R1164_U164 );
nand NAND2_17046 ( P2_R1164_U481 , P2_R1164_U258 , P2_R1164_U479 );
nand NAND2_17047 ( P2_R1164_U482 , P2_U3079 , P2_R1164_U71 );
nand NAND2_17048 ( P2_R1164_U483 , P2_U3492 , P2_R1164_U72 );
nand NAND2_17049 ( P2_R1164_U484 , P2_U3079 , P2_R1164_U71 );
nand NAND2_17050 ( P2_R1164_U485 , P2_U3492 , P2_R1164_U72 );
nand NAND2_17051 ( P2_R1164_U486 , P2_R1164_U485 , P2_R1164_U484 );
nand NAND2_17052 ( P2_R1164_U487 , P2_R1164_U165 , P2_R1164_U166 );
nand NAND2_17053 ( P2_R1164_U488 , P2_R1164_U254 , P2_R1164_U486 );
nand NAND2_17054 ( P2_R1164_U489 , P2_U3080 , P2_R1164_U69 );
nand NAND2_17055 ( P2_R1164_U490 , P2_U3489 , P2_R1164_U70 );
nand NAND2_17056 ( P2_R1164_U491 , P2_U3072 , P2_R1164_U64 );
nand NAND2_17057 ( P2_R1164_U492 , P2_U3486 , P2_R1164_U65 );
nand NAND2_17058 ( P2_R1164_U493 , P2_R1164_U492 , P2_R1164_U491 );
nand NAND2_17059 ( P2_R1164_U494 , P2_R1164_U362 , P2_R1164_U93 );
nand NAND2_17060 ( P2_R1164_U495 , P2_R1164_U493 , P2_R1164_U338 );
nand NAND2_17061 ( P2_R1164_U496 , P2_U3063 , P2_R1164_U66 );
nand NAND2_17062 ( P2_R1164_U497 , P2_U3483 , P2_R1164_U67 );
nand NAND2_17063 ( P2_R1164_U498 , P2_R1164_U497 , P2_R1164_U496 );
nand NAND2_17064 ( P2_R1164_U499 , P2_R1164_U363 , P2_R1164_U167 );
nand NAND2_17065 ( P2_R1164_U500 , P2_R1164_U244 , P2_R1164_U498 );
nand NAND2_17066 ( P2_R1164_U501 , P2_U3062 , P2_R1164_U61 );
nand NAND2_17067 ( P2_R1164_U502 , P2_U3480 , P2_R1164_U62 );
nand NAND2_17068 ( P2_R1164_U503 , P2_U3077 , P2_R1164_U29 );
nand NAND2_17069 ( P2_R1164_U504 , P2_U3448 , P2_R1164_U30 );
and AND2_17070 ( P2_R1233_U4 , P2_R1233_U179 , P2_R1233_U178 );
and AND2_17071 ( P2_R1233_U5 , P2_R1233_U197 , P2_R1233_U196 );
and AND2_17072 ( P2_R1233_U6 , P2_R1233_U237 , P2_R1233_U236 );
and AND2_17073 ( P2_R1233_U7 , P2_R1233_U246 , P2_R1233_U245 );
and AND2_17074 ( P2_R1233_U8 , P2_R1233_U264 , P2_R1233_U263 );
and AND2_17075 ( P2_R1233_U9 , P2_R1233_U272 , P2_R1233_U271 );
and AND2_17076 ( P2_R1233_U10 , P2_R1233_U351 , P2_R1233_U348 );
and AND2_17077 ( P2_R1233_U11 , P2_R1233_U344 , P2_R1233_U341 );
and AND2_17078 ( P2_R1233_U12 , P2_R1233_U335 , P2_R1233_U332 );
and AND2_17079 ( P2_R1233_U13 , P2_R1233_U326 , P2_R1233_U323 );
and AND2_17080 ( P2_R1233_U14 , P2_R1233_U320 , P2_R1233_U318 );
and AND2_17081 ( P2_R1233_U15 , P2_R1233_U313 , P2_R1233_U310 );
and AND2_17082 ( P2_R1233_U16 , P2_R1233_U235 , P2_R1233_U232 );
and AND2_17083 ( P2_R1233_U17 , P2_R1233_U227 , P2_R1233_U224 );
and AND2_17084 ( P2_R1233_U18 , P2_R1233_U213 , P2_R1233_U210 );
not NOT1_17085 ( P2_R1233_U19 , P2_U3468 );
not NOT1_17086 ( P2_R1233_U20 , P2_U3071 );
not NOT1_17087 ( P2_R1233_U21 , P2_U3070 );
nand NAND2_17088 ( P2_R1233_U22 , P2_U3071 , P2_U3468 );
not NOT1_17089 ( P2_R1233_U23 , P2_U3471 );
not NOT1_17090 ( P2_R1233_U24 , P2_U3462 );
not NOT1_17091 ( P2_R1233_U25 , P2_U3060 );
not NOT1_17092 ( P2_R1233_U26 , P2_U3067 );
not NOT1_17093 ( P2_R1233_U27 , P2_U3456 );
not NOT1_17094 ( P2_R1233_U28 , P2_U3068 );
not NOT1_17095 ( P2_R1233_U29 , P2_U3448 );
not NOT1_17096 ( P2_R1233_U30 , P2_U3077 );
nand NAND2_17097 ( P2_R1233_U31 , P2_U3077 , P2_U3448 );
not NOT1_17098 ( P2_R1233_U32 , P2_U3459 );
not NOT1_17099 ( P2_R1233_U33 , P2_U3064 );
nand NAND2_17100 ( P2_R1233_U34 , P2_U3060 , P2_U3462 );
not NOT1_17101 ( P2_R1233_U35 , P2_U3465 );
not NOT1_17102 ( P2_R1233_U36 , P2_U3474 );
not NOT1_17103 ( P2_R1233_U37 , P2_U3084 );
not NOT1_17104 ( P2_R1233_U38 , P2_U3083 );
not NOT1_17105 ( P2_R1233_U39 , P2_U3477 );
nand NAND2_17106 ( P2_R1233_U40 , P2_R1233_U63 , P2_R1233_U205 );
nand NAND2_17107 ( P2_R1233_U41 , P2_R1233_U117 , P2_R1233_U193 );
nand NAND2_17108 ( P2_R1233_U42 , P2_R1233_U182 , P2_R1233_U183 );
nand NAND2_17109 ( P2_R1233_U43 , P2_U3453 , P2_U3078 );
nand NAND2_17110 ( P2_R1233_U44 , P2_R1233_U122 , P2_R1233_U219 );
nand NAND2_17111 ( P2_R1233_U45 , P2_R1233_U216 , P2_R1233_U215 );
not NOT1_17112 ( P2_R1233_U46 , P2_U3969 );
not NOT1_17113 ( P2_R1233_U47 , P2_U3053 );
not NOT1_17114 ( P2_R1233_U48 , P2_U3057 );
not NOT1_17115 ( P2_R1233_U49 , P2_U3970 );
not NOT1_17116 ( P2_R1233_U50 , P2_U3971 );
not NOT1_17117 ( P2_R1233_U51 , P2_U3058 );
not NOT1_17118 ( P2_R1233_U52 , P2_U3972 );
not NOT1_17119 ( P2_R1233_U53 , P2_U3065 );
not NOT1_17120 ( P2_R1233_U54 , P2_U3975 );
not NOT1_17121 ( P2_R1233_U55 , P2_U3075 );
not NOT1_17122 ( P2_R1233_U56 , P2_U3498 );
not NOT1_17123 ( P2_R1233_U57 , P2_U3073 );
not NOT1_17124 ( P2_R1233_U58 , P2_U3069 );
nand NAND2_17125 ( P2_R1233_U59 , P2_U3073 , P2_U3498 );
not NOT1_17126 ( P2_R1233_U60 , P2_U3501 );
not NOT1_17127 ( P2_R1233_U61 , P2_U3480 );
not NOT1_17128 ( P2_R1233_U62 , P2_U3062 );
nand NAND2_17129 ( P2_R1233_U63 , P2_U3084 , P2_U3474 );
not NOT1_17130 ( P2_R1233_U64 , P2_U3486 );
not NOT1_17131 ( P2_R1233_U65 , P2_U3072 );
not NOT1_17132 ( P2_R1233_U66 , P2_U3483 );
not NOT1_17133 ( P2_R1233_U67 , P2_U3063 );
nand NAND2_17134 ( P2_R1233_U68 , P2_U3063 , P2_U3483 );
not NOT1_17135 ( P2_R1233_U69 , P2_U3489 );
not NOT1_17136 ( P2_R1233_U70 , P2_U3080 );
not NOT1_17137 ( P2_R1233_U71 , P2_U3492 );
not NOT1_17138 ( P2_R1233_U72 , P2_U3079 );
not NOT1_17139 ( P2_R1233_U73 , P2_U3495 );
not NOT1_17140 ( P2_R1233_U74 , P2_U3074 );
not NOT1_17141 ( P2_R1233_U75 , P2_U3504 );
not NOT1_17142 ( P2_R1233_U76 , P2_U3082 );
nand NAND2_17143 ( P2_R1233_U77 , P2_U3082 , P2_U3504 );
not NOT1_17144 ( P2_R1233_U78 , P2_U3506 );
not NOT1_17145 ( P2_R1233_U79 , P2_U3081 );
nand NAND2_17146 ( P2_R1233_U80 , P2_U3081 , P2_U3506 );
not NOT1_17147 ( P2_R1233_U81 , P2_U3976 );
not NOT1_17148 ( P2_R1233_U82 , P2_U3974 );
not NOT1_17149 ( P2_R1233_U83 , P2_U3061 );
not NOT1_17150 ( P2_R1233_U84 , P2_U3973 );
not NOT1_17151 ( P2_R1233_U85 , P2_U3066 );
nand NAND2_17152 ( P2_R1233_U86 , P2_U3970 , P2_U3057 );
not NOT1_17153 ( P2_R1233_U87 , P2_U3054 );
not NOT1_17154 ( P2_R1233_U88 , P2_U3968 );
nand NAND2_17155 ( P2_R1233_U89 , P2_R1233_U306 , P2_R1233_U176 );
not NOT1_17156 ( P2_R1233_U90 , P2_U3076 );
nand NAND2_17157 ( P2_R1233_U91 , P2_R1233_U77 , P2_R1233_U315 );
nand NAND2_17158 ( P2_R1233_U92 , P2_R1233_U261 , P2_R1233_U260 );
nand NAND2_17159 ( P2_R1233_U93 , P2_R1233_U68 , P2_R1233_U337 );
nand NAND2_17160 ( P2_R1233_U94 , P2_R1233_U457 , P2_R1233_U456 );
nand NAND2_17161 ( P2_R1233_U95 , P2_R1233_U504 , P2_R1233_U503 );
nand NAND2_17162 ( P2_R1233_U96 , P2_R1233_U375 , P2_R1233_U374 );
nand NAND2_17163 ( P2_R1233_U97 , P2_R1233_U380 , P2_R1233_U379 );
nand NAND2_17164 ( P2_R1233_U98 , P2_R1233_U387 , P2_R1233_U386 );
nand NAND2_17165 ( P2_R1233_U99 , P2_R1233_U394 , P2_R1233_U393 );
nand NAND2_17166 ( P2_R1233_U100 , P2_R1233_U399 , P2_R1233_U398 );
nand NAND2_17167 ( P2_R1233_U101 , P2_R1233_U408 , P2_R1233_U407 );
nand NAND2_17168 ( P2_R1233_U102 , P2_R1233_U415 , P2_R1233_U414 );
nand NAND2_17169 ( P2_R1233_U103 , P2_R1233_U422 , P2_R1233_U421 );
nand NAND2_17170 ( P2_R1233_U104 , P2_R1233_U429 , P2_R1233_U428 );
nand NAND2_17171 ( P2_R1233_U105 , P2_R1233_U434 , P2_R1233_U433 );
nand NAND2_17172 ( P2_R1233_U106 , P2_R1233_U441 , P2_R1233_U440 );
nand NAND2_17173 ( P2_R1233_U107 , P2_R1233_U448 , P2_R1233_U447 );
nand NAND2_17174 ( P2_R1233_U108 , P2_R1233_U462 , P2_R1233_U461 );
nand NAND2_17175 ( P2_R1233_U109 , P2_R1233_U467 , P2_R1233_U466 );
nand NAND2_17176 ( P2_R1233_U110 , P2_R1233_U474 , P2_R1233_U473 );
nand NAND2_17177 ( P2_R1233_U111 , P2_R1233_U481 , P2_R1233_U480 );
nand NAND2_17178 ( P2_R1233_U112 , P2_R1233_U488 , P2_R1233_U487 );
nand NAND2_17179 ( P2_R1233_U113 , P2_R1233_U495 , P2_R1233_U494 );
nand NAND2_17180 ( P2_R1233_U114 , P2_R1233_U500 , P2_R1233_U499 );
and AND2_17181 ( P2_R1233_U115 , P2_R1233_U189 , P2_R1233_U187 );
and AND2_17182 ( P2_R1233_U116 , P2_R1233_U4 , P2_R1233_U180 );
and AND2_17183 ( P2_R1233_U117 , P2_R1233_U194 , P2_R1233_U192 );
and AND2_17184 ( P2_R1233_U118 , P2_R1233_U201 , P2_R1233_U200 );
and AND3_17185 ( P2_R1233_U119 , P2_R1233_U382 , P2_R1233_U381 , P2_R1233_U22 );
and AND2_17186 ( P2_R1233_U120 , P2_R1233_U212 , P2_R1233_U5 );
and AND2_17187 ( P2_R1233_U121 , P2_R1233_U181 , P2_R1233_U180 );
and AND2_17188 ( P2_R1233_U122 , P2_R1233_U220 , P2_R1233_U218 );
and AND3_17189 ( P2_R1233_U123 , P2_R1233_U389 , P2_R1233_U388 , P2_R1233_U34 );
and AND2_17190 ( P2_R1233_U124 , P2_R1233_U226 , P2_R1233_U4 );
and AND2_17191 ( P2_R1233_U125 , P2_R1233_U234 , P2_R1233_U181 );
and AND2_17192 ( P2_R1233_U126 , P2_R1233_U204 , P2_R1233_U6 );
and AND2_17193 ( P2_R1233_U127 , P2_R1233_U243 , P2_R1233_U239 );
and AND2_17194 ( P2_R1233_U128 , P2_R1233_U250 , P2_R1233_U7 );
and AND2_17195 ( P2_R1233_U129 , P2_R1233_U248 , P2_R1233_U172 );
and AND2_17196 ( P2_R1233_U130 , P2_R1233_U268 , P2_R1233_U267 );
and AND3_17197 ( P2_R1233_U131 , P2_R1233_U9 , P2_R1233_U282 , P2_R1233_U273 );
and AND2_17198 ( P2_R1233_U132 , P2_R1233_U285 , P2_R1233_U280 );
and AND2_17199 ( P2_R1233_U133 , P2_R1233_U301 , P2_R1233_U298 );
and AND2_17200 ( P2_R1233_U134 , P2_R1233_U368 , P2_R1233_U302 );
and AND3_17201 ( P2_R1233_U135 , P2_R1233_U424 , P2_R1233_U423 , P2_R1233_U173 );
and AND2_17202 ( P2_R1233_U136 , P2_R1233_U160 , P2_R1233_U278 );
and AND3_17203 ( P2_R1233_U137 , P2_R1233_U455 , P2_R1233_U454 , P2_R1233_U80 );
and AND2_17204 ( P2_R1233_U138 , P2_R1233_U325 , P2_R1233_U9 );
and AND3_17205 ( P2_R1233_U139 , P2_R1233_U469 , P2_R1233_U468 , P2_R1233_U59 );
and AND2_17206 ( P2_R1233_U140 , P2_R1233_U334 , P2_R1233_U8 );
and AND3_17207 ( P2_R1233_U141 , P2_R1233_U490 , P2_R1233_U489 , P2_R1233_U172 );
and AND2_17208 ( P2_R1233_U142 , P2_R1233_U343 , P2_R1233_U7 );
and AND3_17209 ( P2_R1233_U143 , P2_R1233_U502 , P2_R1233_U501 , P2_R1233_U171 );
and AND2_17210 ( P2_R1233_U144 , P2_R1233_U350 , P2_R1233_U6 );
nand NAND2_17211 ( P2_R1233_U145 , P2_R1233_U118 , P2_R1233_U202 );
nand NAND2_17212 ( P2_R1233_U146 , P2_R1233_U217 , P2_R1233_U229 );
not NOT1_17213 ( P2_R1233_U147 , P2_U3055 );
not NOT1_17214 ( P2_R1233_U148 , P2_U3979 );
and AND2_17215 ( P2_R1233_U149 , P2_R1233_U403 , P2_R1233_U402 );
nand NAND3_17216 ( P2_R1233_U150 , P2_R1233_U304 , P2_R1233_U169 , P2_R1233_U364 );
and AND2_17217 ( P2_R1233_U151 , P2_R1233_U410 , P2_R1233_U409 );
nand NAND3_17218 ( P2_R1233_U152 , P2_R1233_U370 , P2_R1233_U369 , P2_R1233_U134 );
and AND2_17219 ( P2_R1233_U153 , P2_R1233_U417 , P2_R1233_U416 );
nand NAND3_17220 ( P2_R1233_U154 , P2_R1233_U365 , P2_R1233_U299 , P2_R1233_U86 );
nand NAND2_17221 ( P2_R1233_U155 , P2_R1233_U293 , P2_R1233_U292 );
and AND2_17222 ( P2_R1233_U156 , P2_R1233_U436 , P2_R1233_U435 );
nand NAND2_17223 ( P2_R1233_U157 , P2_R1233_U289 , P2_R1233_U288 );
and AND2_17224 ( P2_R1233_U158 , P2_R1233_U443 , P2_R1233_U442 );
nand NAND2_17225 ( P2_R1233_U159 , P2_R1233_U132 , P2_R1233_U284 );
and AND2_17226 ( P2_R1233_U160 , P2_R1233_U450 , P2_R1233_U449 );
nand NAND2_17227 ( P2_R1233_U161 , P2_R1233_U43 , P2_R1233_U327 );
nand NAND2_17228 ( P2_R1233_U162 , P2_R1233_U130 , P2_R1233_U269 );
and AND2_17229 ( P2_R1233_U163 , P2_R1233_U476 , P2_R1233_U475 );
nand NAND2_17230 ( P2_R1233_U164 , P2_R1233_U257 , P2_R1233_U256 );
and AND2_17231 ( P2_R1233_U165 , P2_R1233_U483 , P2_R1233_U482 );
nand NAND2_17232 ( P2_R1233_U166 , P2_R1233_U253 , P2_R1233_U252 );
nand NAND2_17233 ( P2_R1233_U167 , P2_R1233_U127 , P2_R1233_U242 );
nand NAND2_17234 ( P2_R1233_U168 , P2_R1233_U367 , P2_R1233_U366 );
nand NAND2_17235 ( P2_R1233_U169 , P2_U3054 , P2_R1233_U152 );
not NOT1_17236 ( P2_R1233_U170 , P2_R1233_U34 );
nand NAND2_17237 ( P2_R1233_U171 , P2_U3477 , P2_U3083 );
nand NAND2_17238 ( P2_R1233_U172 , P2_U3072 , P2_U3486 );
nand NAND2_17239 ( P2_R1233_U173 , P2_U3058 , P2_U3971 );
not NOT1_17240 ( P2_R1233_U174 , P2_R1233_U68 );
not NOT1_17241 ( P2_R1233_U175 , P2_R1233_U77 );
nand NAND2_17242 ( P2_R1233_U176 , P2_U3065 , P2_U3972 );
not NOT1_17243 ( P2_R1233_U177 , P2_R1233_U63 );
or OR2_17244 ( P2_R1233_U178 , P2_U3067 , P2_U3465 );
or OR2_17245 ( P2_R1233_U179 , P2_U3060 , P2_U3462 );
or OR2_17246 ( P2_R1233_U180 , P2_U3459 , P2_U3064 );
or OR2_17247 ( P2_R1233_U181 , P2_U3456 , P2_U3068 );
not NOT1_17248 ( P2_R1233_U182 , P2_R1233_U31 );
or OR2_17249 ( P2_R1233_U183 , P2_U3453 , P2_U3078 );
not NOT1_17250 ( P2_R1233_U184 , P2_R1233_U42 );
not NOT1_17251 ( P2_R1233_U185 , P2_R1233_U43 );
nand NAND2_17252 ( P2_R1233_U186 , P2_R1233_U42 , P2_R1233_U43 );
nand NAND2_17253 ( P2_R1233_U187 , P2_U3068 , P2_U3456 );
nand NAND2_17254 ( P2_R1233_U188 , P2_R1233_U186 , P2_R1233_U181 );
nand NAND2_17255 ( P2_R1233_U189 , P2_U3064 , P2_U3459 );
nand NAND2_17256 ( P2_R1233_U190 , P2_R1233_U115 , P2_R1233_U188 );
nand NAND2_17257 ( P2_R1233_U191 , P2_R1233_U35 , P2_R1233_U34 );
nand NAND2_17258 ( P2_R1233_U192 , P2_U3067 , P2_R1233_U191 );
nand NAND2_17259 ( P2_R1233_U193 , P2_R1233_U116 , P2_R1233_U190 );
nand NAND2_17260 ( P2_R1233_U194 , P2_U3465 , P2_R1233_U170 );
not NOT1_17261 ( P2_R1233_U195 , P2_R1233_U41 );
or OR2_17262 ( P2_R1233_U196 , P2_U3070 , P2_U3471 );
or OR2_17263 ( P2_R1233_U197 , P2_U3071 , P2_U3468 );
not NOT1_17264 ( P2_R1233_U198 , P2_R1233_U22 );
nand NAND2_17265 ( P2_R1233_U199 , P2_R1233_U23 , P2_R1233_U22 );
nand NAND2_17266 ( P2_R1233_U200 , P2_U3070 , P2_R1233_U199 );
nand NAND2_17267 ( P2_R1233_U201 , P2_U3471 , P2_R1233_U198 );
nand NAND2_17268 ( P2_R1233_U202 , P2_R1233_U5 , P2_R1233_U41 );
not NOT1_17269 ( P2_R1233_U203 , P2_R1233_U145 );
or OR2_17270 ( P2_R1233_U204 , P2_U3474 , P2_U3084 );
nand NAND2_17271 ( P2_R1233_U205 , P2_R1233_U204 , P2_R1233_U145 );
not NOT1_17272 ( P2_R1233_U206 , P2_R1233_U40 );
or OR2_17273 ( P2_R1233_U207 , P2_U3083 , P2_U3477 );
or OR2_17274 ( P2_R1233_U208 , P2_U3468 , P2_U3071 );
nand NAND2_17275 ( P2_R1233_U209 , P2_R1233_U208 , P2_R1233_U41 );
nand NAND2_17276 ( P2_R1233_U210 , P2_R1233_U119 , P2_R1233_U209 );
nand NAND2_17277 ( P2_R1233_U211 , P2_R1233_U195 , P2_R1233_U22 );
nand NAND2_17278 ( P2_R1233_U212 , P2_U3471 , P2_U3070 );
nand NAND2_17279 ( P2_R1233_U213 , P2_R1233_U120 , P2_R1233_U211 );
or OR2_17280 ( P2_R1233_U214 , P2_U3071 , P2_U3468 );
nand NAND2_17281 ( P2_R1233_U215 , P2_R1233_U185 , P2_R1233_U181 );
nand NAND2_17282 ( P2_R1233_U216 , P2_U3068 , P2_U3456 );
not NOT1_17283 ( P2_R1233_U217 , P2_R1233_U45 );
nand NAND2_17284 ( P2_R1233_U218 , P2_R1233_U121 , P2_R1233_U184 );
nand NAND2_17285 ( P2_R1233_U219 , P2_R1233_U45 , P2_R1233_U180 );
nand NAND2_17286 ( P2_R1233_U220 , P2_U3064 , P2_U3459 );
not NOT1_17287 ( P2_R1233_U221 , P2_R1233_U44 );
or OR2_17288 ( P2_R1233_U222 , P2_U3462 , P2_U3060 );
nand NAND2_17289 ( P2_R1233_U223 , P2_R1233_U222 , P2_R1233_U44 );
nand NAND2_17290 ( P2_R1233_U224 , P2_R1233_U123 , P2_R1233_U223 );
nand NAND2_17291 ( P2_R1233_U225 , P2_R1233_U221 , P2_R1233_U34 );
nand NAND2_17292 ( P2_R1233_U226 , P2_U3465 , P2_U3067 );
nand NAND2_17293 ( P2_R1233_U227 , P2_R1233_U124 , P2_R1233_U225 );
or OR2_17294 ( P2_R1233_U228 , P2_U3060 , P2_U3462 );
nand NAND2_17295 ( P2_R1233_U229 , P2_R1233_U184 , P2_R1233_U181 );
not NOT1_17296 ( P2_R1233_U230 , P2_R1233_U146 );
nand NAND2_17297 ( P2_R1233_U231 , P2_U3064 , P2_U3459 );
nand NAND4_17298 ( P2_R1233_U232 , P2_R1233_U401 , P2_R1233_U400 , P2_R1233_U43 , P2_R1233_U42 );
nand NAND2_17299 ( P2_R1233_U233 , P2_R1233_U43 , P2_R1233_U42 );
nand NAND2_17300 ( P2_R1233_U234 , P2_U3068 , P2_U3456 );
nand NAND2_17301 ( P2_R1233_U235 , P2_R1233_U125 , P2_R1233_U233 );
or OR2_17302 ( P2_R1233_U236 , P2_U3083 , P2_U3477 );
or OR2_17303 ( P2_R1233_U237 , P2_U3062 , P2_U3480 );
nand NAND2_17304 ( P2_R1233_U238 , P2_R1233_U177 , P2_R1233_U6 );
nand NAND2_17305 ( P2_R1233_U239 , P2_U3062 , P2_U3480 );
nand NAND2_17306 ( P2_R1233_U240 , P2_R1233_U171 , P2_R1233_U238 );
or OR2_17307 ( P2_R1233_U241 , P2_U3480 , P2_U3062 );
nand NAND2_17308 ( P2_R1233_U242 , P2_R1233_U126 , P2_R1233_U145 );
nand NAND2_17309 ( P2_R1233_U243 , P2_R1233_U241 , P2_R1233_U240 );
not NOT1_17310 ( P2_R1233_U244 , P2_R1233_U167 );
or OR2_17311 ( P2_R1233_U245 , P2_U3080 , P2_U3489 );
or OR2_17312 ( P2_R1233_U246 , P2_U3072 , P2_U3486 );
nand NAND2_17313 ( P2_R1233_U247 , P2_R1233_U174 , P2_R1233_U7 );
nand NAND2_17314 ( P2_R1233_U248 , P2_U3080 , P2_U3489 );
nand NAND2_17315 ( P2_R1233_U249 , P2_R1233_U129 , P2_R1233_U247 );
or OR2_17316 ( P2_R1233_U250 , P2_U3483 , P2_U3063 );
or OR2_17317 ( P2_R1233_U251 , P2_U3489 , P2_U3080 );
nand NAND2_17318 ( P2_R1233_U252 , P2_R1233_U128 , P2_R1233_U167 );
nand NAND2_17319 ( P2_R1233_U253 , P2_R1233_U251 , P2_R1233_U249 );
not NOT1_17320 ( P2_R1233_U254 , P2_R1233_U166 );
or OR2_17321 ( P2_R1233_U255 , P2_U3492 , P2_U3079 );
nand NAND2_17322 ( P2_R1233_U256 , P2_R1233_U255 , P2_R1233_U166 );
nand NAND2_17323 ( P2_R1233_U257 , P2_U3079 , P2_U3492 );
not NOT1_17324 ( P2_R1233_U258 , P2_R1233_U164 );
or OR2_17325 ( P2_R1233_U259 , P2_U3495 , P2_U3074 );
nand NAND2_17326 ( P2_R1233_U260 , P2_R1233_U259 , P2_R1233_U164 );
nand NAND2_17327 ( P2_R1233_U261 , P2_U3074 , P2_U3495 );
not NOT1_17328 ( P2_R1233_U262 , P2_R1233_U92 );
or OR2_17329 ( P2_R1233_U263 , P2_U3069 , P2_U3501 );
or OR2_17330 ( P2_R1233_U264 , P2_U3073 , P2_U3498 );
not NOT1_17331 ( P2_R1233_U265 , P2_R1233_U59 );
nand NAND2_17332 ( P2_R1233_U266 , P2_R1233_U60 , P2_R1233_U59 );
nand NAND2_17333 ( P2_R1233_U267 , P2_U3069 , P2_R1233_U266 );
nand NAND2_17334 ( P2_R1233_U268 , P2_U3501 , P2_R1233_U265 );
nand NAND2_17335 ( P2_R1233_U269 , P2_R1233_U8 , P2_R1233_U92 );
not NOT1_17336 ( P2_R1233_U270 , P2_R1233_U162 );
or OR2_17337 ( P2_R1233_U271 , P2_U3076 , P2_U3976 );
or OR2_17338 ( P2_R1233_U272 , P2_U3081 , P2_U3506 );
or OR2_17339 ( P2_R1233_U273 , P2_U3075 , P2_U3975 );
not NOT1_17340 ( P2_R1233_U274 , P2_R1233_U80 );
nand NAND2_17341 ( P2_R1233_U275 , P2_U3976 , P2_R1233_U274 );
nand NAND2_17342 ( P2_R1233_U276 , P2_R1233_U275 , P2_R1233_U90 );
nand NAND2_17343 ( P2_R1233_U277 , P2_R1233_U80 , P2_R1233_U81 );
nand NAND2_17344 ( P2_R1233_U278 , P2_R1233_U277 , P2_R1233_U276 );
nand NAND2_17345 ( P2_R1233_U279 , P2_R1233_U175 , P2_R1233_U9 );
nand NAND2_17346 ( P2_R1233_U280 , P2_U3075 , P2_U3975 );
nand NAND2_17347 ( P2_R1233_U281 , P2_R1233_U278 , P2_R1233_U279 );
or OR2_17348 ( P2_R1233_U282 , P2_U3504 , P2_U3082 );
or OR2_17349 ( P2_R1233_U283 , P2_U3975 , P2_U3075 );
nand NAND2_17350 ( P2_R1233_U284 , P2_R1233_U162 , P2_R1233_U131 );
nand NAND2_17351 ( P2_R1233_U285 , P2_R1233_U283 , P2_R1233_U281 );
not NOT1_17352 ( P2_R1233_U286 , P2_R1233_U159 );
or OR2_17353 ( P2_R1233_U287 , P2_U3974 , P2_U3061 );
nand NAND2_17354 ( P2_R1233_U288 , P2_R1233_U287 , P2_R1233_U159 );
nand NAND2_17355 ( P2_R1233_U289 , P2_U3061 , P2_U3974 );
not NOT1_17356 ( P2_R1233_U290 , P2_R1233_U157 );
or OR2_17357 ( P2_R1233_U291 , P2_U3973 , P2_U3066 );
nand NAND2_17358 ( P2_R1233_U292 , P2_R1233_U291 , P2_R1233_U157 );
nand NAND2_17359 ( P2_R1233_U293 , P2_U3066 , P2_U3973 );
not NOT1_17360 ( P2_R1233_U294 , P2_R1233_U155 );
or OR2_17361 ( P2_R1233_U295 , P2_U3058 , P2_U3971 );
nand NAND2_17362 ( P2_R1233_U296 , P2_R1233_U176 , P2_R1233_U173 );
not NOT1_17363 ( P2_R1233_U297 , P2_R1233_U86 );
or OR2_17364 ( P2_R1233_U298 , P2_U3972 , P2_U3065 );
nand NAND3_17365 ( P2_R1233_U299 , P2_R1233_U155 , P2_R1233_U298 , P2_R1233_U168 );
not NOT1_17366 ( P2_R1233_U300 , P2_R1233_U154 );
or OR2_17367 ( P2_R1233_U301 , P2_U3969 , P2_U3053 );
nand NAND2_17368 ( P2_R1233_U302 , P2_U3053 , P2_U3969 );
not NOT1_17369 ( P2_R1233_U303 , P2_R1233_U152 );
nand NAND2_17370 ( P2_R1233_U304 , P2_U3968 , P2_R1233_U152 );
not NOT1_17371 ( P2_R1233_U305 , P2_R1233_U150 );
nand NAND2_17372 ( P2_R1233_U306 , P2_R1233_U298 , P2_R1233_U155 );
not NOT1_17373 ( P2_R1233_U307 , P2_R1233_U89 );
or OR2_17374 ( P2_R1233_U308 , P2_U3971 , P2_U3058 );
nand NAND2_17375 ( P2_R1233_U309 , P2_R1233_U308 , P2_R1233_U89 );
nand NAND2_17376 ( P2_R1233_U310 , P2_R1233_U135 , P2_R1233_U309 );
nand NAND2_17377 ( P2_R1233_U311 , P2_R1233_U307 , P2_R1233_U173 );
nand NAND2_17378 ( P2_R1233_U312 , P2_U3970 , P2_U3057 );
nand NAND3_17379 ( P2_R1233_U313 , P2_R1233_U311 , P2_R1233_U312 , P2_R1233_U168 );
or OR2_17380 ( P2_R1233_U314 , P2_U3058 , P2_U3971 );
nand NAND2_17381 ( P2_R1233_U315 , P2_R1233_U282 , P2_R1233_U162 );
not NOT1_17382 ( P2_R1233_U316 , P2_R1233_U91 );
nand NAND2_17383 ( P2_R1233_U317 , P2_R1233_U9 , P2_R1233_U91 );
nand NAND2_17384 ( P2_R1233_U318 , P2_R1233_U136 , P2_R1233_U317 );
nand NAND2_17385 ( P2_R1233_U319 , P2_R1233_U317 , P2_R1233_U278 );
nand NAND2_17386 ( P2_R1233_U320 , P2_R1233_U453 , P2_R1233_U319 );
or OR2_17387 ( P2_R1233_U321 , P2_U3506 , P2_U3081 );
nand NAND2_17388 ( P2_R1233_U322 , P2_R1233_U321 , P2_R1233_U91 );
nand NAND2_17389 ( P2_R1233_U323 , P2_R1233_U137 , P2_R1233_U322 );
nand NAND2_17390 ( P2_R1233_U324 , P2_R1233_U316 , P2_R1233_U80 );
nand NAND2_17391 ( P2_R1233_U325 , P2_U3076 , P2_U3976 );
nand NAND2_17392 ( P2_R1233_U326 , P2_R1233_U138 , P2_R1233_U324 );
or OR2_17393 ( P2_R1233_U327 , P2_U3453 , P2_U3078 );
not NOT1_17394 ( P2_R1233_U328 , P2_R1233_U161 );
or OR2_17395 ( P2_R1233_U329 , P2_U3081 , P2_U3506 );
or OR2_17396 ( P2_R1233_U330 , P2_U3498 , P2_U3073 );
nand NAND2_17397 ( P2_R1233_U331 , P2_R1233_U330 , P2_R1233_U92 );
nand NAND2_17398 ( P2_R1233_U332 , P2_R1233_U139 , P2_R1233_U331 );
nand NAND2_17399 ( P2_R1233_U333 , P2_R1233_U262 , P2_R1233_U59 );
nand NAND2_17400 ( P2_R1233_U334 , P2_U3501 , P2_U3069 );
nand NAND2_17401 ( P2_R1233_U335 , P2_R1233_U140 , P2_R1233_U333 );
or OR2_17402 ( P2_R1233_U336 , P2_U3073 , P2_U3498 );
nand NAND2_17403 ( P2_R1233_U337 , P2_R1233_U250 , P2_R1233_U167 );
not NOT1_17404 ( P2_R1233_U338 , P2_R1233_U93 );
or OR2_17405 ( P2_R1233_U339 , P2_U3486 , P2_U3072 );
nand NAND2_17406 ( P2_R1233_U340 , P2_R1233_U339 , P2_R1233_U93 );
nand NAND2_17407 ( P2_R1233_U341 , P2_R1233_U141 , P2_R1233_U340 );
nand NAND2_17408 ( P2_R1233_U342 , P2_R1233_U338 , P2_R1233_U172 );
nand NAND2_17409 ( P2_R1233_U343 , P2_U3080 , P2_U3489 );
nand NAND2_17410 ( P2_R1233_U344 , P2_R1233_U142 , P2_R1233_U342 );
or OR2_17411 ( P2_R1233_U345 , P2_U3072 , P2_U3486 );
or OR2_17412 ( P2_R1233_U346 , P2_U3477 , P2_U3083 );
nand NAND2_17413 ( P2_R1233_U347 , P2_R1233_U346 , P2_R1233_U40 );
nand NAND2_17414 ( P2_R1233_U348 , P2_R1233_U143 , P2_R1233_U347 );
nand NAND2_17415 ( P2_R1233_U349 , P2_R1233_U206 , P2_R1233_U171 );
nand NAND2_17416 ( P2_R1233_U350 , P2_U3062 , P2_U3480 );
nand NAND2_17417 ( P2_R1233_U351 , P2_R1233_U144 , P2_R1233_U349 );
nand NAND2_17418 ( P2_R1233_U352 , P2_R1233_U207 , P2_R1233_U171 );
nand NAND2_17419 ( P2_R1233_U353 , P2_R1233_U204 , P2_R1233_U63 );
nand NAND2_17420 ( P2_R1233_U354 , P2_R1233_U214 , P2_R1233_U22 );
nand NAND2_17421 ( P2_R1233_U355 , P2_R1233_U228 , P2_R1233_U34 );
nand NAND2_17422 ( P2_R1233_U356 , P2_R1233_U231 , P2_R1233_U180 );
nand NAND2_17423 ( P2_R1233_U357 , P2_R1233_U314 , P2_R1233_U173 );
nand NAND2_17424 ( P2_R1233_U358 , P2_R1233_U298 , P2_R1233_U176 );
nand NAND2_17425 ( P2_R1233_U359 , P2_R1233_U329 , P2_R1233_U80 );
nand NAND2_17426 ( P2_R1233_U360 , P2_R1233_U282 , P2_R1233_U77 );
nand NAND2_17427 ( P2_R1233_U361 , P2_R1233_U336 , P2_R1233_U59 );
nand NAND2_17428 ( P2_R1233_U362 , P2_R1233_U345 , P2_R1233_U172 );
nand NAND2_17429 ( P2_R1233_U363 , P2_R1233_U250 , P2_R1233_U68 );
nand NAND2_17430 ( P2_R1233_U364 , P2_U3968 , P2_U3054 );
nand NAND2_17431 ( P2_R1233_U365 , P2_R1233_U296 , P2_R1233_U168 );
nand NAND2_17432 ( P2_R1233_U366 , P2_U3057 , P2_R1233_U295 );
nand NAND2_17433 ( P2_R1233_U367 , P2_U3970 , P2_R1233_U295 );
nand NAND3_17434 ( P2_R1233_U368 , P2_R1233_U296 , P2_R1233_U168 , P2_R1233_U301 );
nand NAND3_17435 ( P2_R1233_U369 , P2_R1233_U155 , P2_R1233_U168 , P2_R1233_U133 );
nand NAND2_17436 ( P2_R1233_U370 , P2_R1233_U297 , P2_R1233_U301 );
nand NAND2_17437 ( P2_R1233_U371 , P2_U3083 , P2_R1233_U39 );
nand NAND2_17438 ( P2_R1233_U372 , P2_U3477 , P2_R1233_U38 );
nand NAND2_17439 ( P2_R1233_U373 , P2_R1233_U372 , P2_R1233_U371 );
nand NAND2_17440 ( P2_R1233_U374 , P2_R1233_U352 , P2_R1233_U40 );
nand NAND2_17441 ( P2_R1233_U375 , P2_R1233_U373 , P2_R1233_U206 );
nand NAND2_17442 ( P2_R1233_U376 , P2_U3084 , P2_R1233_U36 );
nand NAND2_17443 ( P2_R1233_U377 , P2_U3474 , P2_R1233_U37 );
nand NAND2_17444 ( P2_R1233_U378 , P2_R1233_U377 , P2_R1233_U376 );
nand NAND2_17445 ( P2_R1233_U379 , P2_R1233_U353 , P2_R1233_U145 );
nand NAND2_17446 ( P2_R1233_U380 , P2_R1233_U203 , P2_R1233_U378 );
nand NAND2_17447 ( P2_R1233_U381 , P2_U3070 , P2_R1233_U23 );
nand NAND2_17448 ( P2_R1233_U382 , P2_U3471 , P2_R1233_U21 );
nand NAND2_17449 ( P2_R1233_U383 , P2_U3071 , P2_R1233_U19 );
nand NAND2_17450 ( P2_R1233_U384 , P2_U3468 , P2_R1233_U20 );
nand NAND2_17451 ( P2_R1233_U385 , P2_R1233_U384 , P2_R1233_U383 );
nand NAND2_17452 ( P2_R1233_U386 , P2_R1233_U354 , P2_R1233_U41 );
nand NAND2_17453 ( P2_R1233_U387 , P2_R1233_U385 , P2_R1233_U195 );
nand NAND2_17454 ( P2_R1233_U388 , P2_U3067 , P2_R1233_U35 );
nand NAND2_17455 ( P2_R1233_U389 , P2_U3465 , P2_R1233_U26 );
nand NAND2_17456 ( P2_R1233_U390 , P2_U3060 , P2_R1233_U24 );
nand NAND2_17457 ( P2_R1233_U391 , P2_U3462 , P2_R1233_U25 );
nand NAND2_17458 ( P2_R1233_U392 , P2_R1233_U391 , P2_R1233_U390 );
nand NAND2_17459 ( P2_R1233_U393 , P2_R1233_U355 , P2_R1233_U44 );
nand NAND2_17460 ( P2_R1233_U394 , P2_R1233_U392 , P2_R1233_U221 );
nand NAND2_17461 ( P2_R1233_U395 , P2_U3064 , P2_R1233_U32 );
nand NAND2_17462 ( P2_R1233_U396 , P2_U3459 , P2_R1233_U33 );
nand NAND2_17463 ( P2_R1233_U397 , P2_R1233_U396 , P2_R1233_U395 );
nand NAND2_17464 ( P2_R1233_U398 , P2_R1233_U356 , P2_R1233_U146 );
nand NAND2_17465 ( P2_R1233_U399 , P2_R1233_U230 , P2_R1233_U397 );
nand NAND2_17466 ( P2_R1233_U400 , P2_U3068 , P2_R1233_U27 );
nand NAND2_17467 ( P2_R1233_U401 , P2_U3456 , P2_R1233_U28 );
nand NAND2_17468 ( P2_R1233_U402 , P2_U3055 , P2_R1233_U148 );
nand NAND2_17469 ( P2_R1233_U403 , P2_U3979 , P2_R1233_U147 );
nand NAND2_17470 ( P2_R1233_U404 , P2_U3055 , P2_R1233_U148 );
nand NAND2_17471 ( P2_R1233_U405 , P2_U3979 , P2_R1233_U147 );
nand NAND2_17472 ( P2_R1233_U406 , P2_R1233_U405 , P2_R1233_U404 );
nand NAND2_17473 ( P2_R1233_U407 , P2_R1233_U149 , P2_R1233_U150 );
nand NAND2_17474 ( P2_R1233_U408 , P2_R1233_U305 , P2_R1233_U406 );
nand NAND2_17475 ( P2_R1233_U409 , P2_U3054 , P2_R1233_U88 );
nand NAND2_17476 ( P2_R1233_U410 , P2_U3968 , P2_R1233_U87 );
nand NAND2_17477 ( P2_R1233_U411 , P2_U3054 , P2_R1233_U88 );
nand NAND2_17478 ( P2_R1233_U412 , P2_U3968 , P2_R1233_U87 );
nand NAND2_17479 ( P2_R1233_U413 , P2_R1233_U412 , P2_R1233_U411 );
nand NAND2_17480 ( P2_R1233_U414 , P2_R1233_U151 , P2_R1233_U152 );
nand NAND2_17481 ( P2_R1233_U415 , P2_R1233_U303 , P2_R1233_U413 );
nand NAND2_17482 ( P2_R1233_U416 , P2_U3053 , P2_R1233_U46 );
nand NAND2_17483 ( P2_R1233_U417 , P2_U3969 , P2_R1233_U47 );
nand NAND2_17484 ( P2_R1233_U418 , P2_U3053 , P2_R1233_U46 );
nand NAND2_17485 ( P2_R1233_U419 , P2_U3969 , P2_R1233_U47 );
nand NAND2_17486 ( P2_R1233_U420 , P2_R1233_U419 , P2_R1233_U418 );
nand NAND2_17487 ( P2_R1233_U421 , P2_R1233_U153 , P2_R1233_U154 );
nand NAND2_17488 ( P2_R1233_U422 , P2_R1233_U300 , P2_R1233_U420 );
nand NAND2_17489 ( P2_R1233_U423 , P2_U3057 , P2_R1233_U49 );
nand NAND2_17490 ( P2_R1233_U424 , P2_U3970 , P2_R1233_U48 );
nand NAND2_17491 ( P2_R1233_U425 , P2_U3058 , P2_R1233_U50 );
nand NAND2_17492 ( P2_R1233_U426 , P2_U3971 , P2_R1233_U51 );
nand NAND2_17493 ( P2_R1233_U427 , P2_R1233_U426 , P2_R1233_U425 );
nand NAND2_17494 ( P2_R1233_U428 , P2_R1233_U357 , P2_R1233_U89 );
nand NAND2_17495 ( P2_R1233_U429 , P2_R1233_U427 , P2_R1233_U307 );
nand NAND2_17496 ( P2_R1233_U430 , P2_U3065 , P2_R1233_U52 );
nand NAND2_17497 ( P2_R1233_U431 , P2_U3972 , P2_R1233_U53 );
nand NAND2_17498 ( P2_R1233_U432 , P2_R1233_U431 , P2_R1233_U430 );
nand NAND2_17499 ( P2_R1233_U433 , P2_R1233_U358 , P2_R1233_U155 );
nand NAND2_17500 ( P2_R1233_U434 , P2_R1233_U294 , P2_R1233_U432 );
nand NAND2_17501 ( P2_R1233_U435 , P2_U3066 , P2_R1233_U84 );
nand NAND2_17502 ( P2_R1233_U436 , P2_U3973 , P2_R1233_U85 );
nand NAND2_17503 ( P2_R1233_U437 , P2_U3066 , P2_R1233_U84 );
nand NAND2_17504 ( P2_R1233_U438 , P2_U3973 , P2_R1233_U85 );
nand NAND2_17505 ( P2_R1233_U439 , P2_R1233_U438 , P2_R1233_U437 );
nand NAND2_17506 ( P2_R1233_U440 , P2_R1233_U156 , P2_R1233_U157 );
nand NAND2_17507 ( P2_R1233_U441 , P2_R1233_U290 , P2_R1233_U439 );
nand NAND2_17508 ( P2_R1233_U442 , P2_U3061 , P2_R1233_U82 );
nand NAND2_17509 ( P2_R1233_U443 , P2_U3974 , P2_R1233_U83 );
nand NAND2_17510 ( P2_R1233_U444 , P2_U3061 , P2_R1233_U82 );
nand NAND2_17511 ( P2_R1233_U445 , P2_U3974 , P2_R1233_U83 );
nand NAND2_17512 ( P2_R1233_U446 , P2_R1233_U445 , P2_R1233_U444 );
nand NAND2_17513 ( P2_R1233_U447 , P2_R1233_U158 , P2_R1233_U159 );
nand NAND2_17514 ( P2_R1233_U448 , P2_R1233_U286 , P2_R1233_U446 );
nand NAND2_17515 ( P2_R1233_U449 , P2_U3075 , P2_R1233_U54 );
nand NAND2_17516 ( P2_R1233_U450 , P2_U3975 , P2_R1233_U55 );
nand NAND2_17517 ( P2_R1233_U451 , P2_U3075 , P2_R1233_U54 );
nand NAND2_17518 ( P2_R1233_U452 , P2_U3975 , P2_R1233_U55 );
nand NAND2_17519 ( P2_R1233_U453 , P2_R1233_U452 , P2_R1233_U451 );
nand NAND2_17520 ( P2_R1233_U454 , P2_U3076 , P2_R1233_U81 );
nand NAND2_17521 ( P2_R1233_U455 , P2_U3976 , P2_R1233_U90 );
nand NAND2_17522 ( P2_R1233_U456 , P2_R1233_U182 , P2_R1233_U161 );
nand NAND2_17523 ( P2_R1233_U457 , P2_R1233_U328 , P2_R1233_U31 );
nand NAND2_17524 ( P2_R1233_U458 , P2_U3081 , P2_R1233_U78 );
nand NAND2_17525 ( P2_R1233_U459 , P2_U3506 , P2_R1233_U79 );
nand NAND2_17526 ( P2_R1233_U460 , P2_R1233_U459 , P2_R1233_U458 );
nand NAND2_17527 ( P2_R1233_U461 , P2_R1233_U359 , P2_R1233_U91 );
nand NAND2_17528 ( P2_R1233_U462 , P2_R1233_U460 , P2_R1233_U316 );
nand NAND2_17529 ( P2_R1233_U463 , P2_U3082 , P2_R1233_U75 );
nand NAND2_17530 ( P2_R1233_U464 , P2_U3504 , P2_R1233_U76 );
nand NAND2_17531 ( P2_R1233_U465 , P2_R1233_U464 , P2_R1233_U463 );
nand NAND2_17532 ( P2_R1233_U466 , P2_R1233_U360 , P2_R1233_U162 );
nand NAND2_17533 ( P2_R1233_U467 , P2_R1233_U270 , P2_R1233_U465 );
nand NAND2_17534 ( P2_R1233_U468 , P2_U3069 , P2_R1233_U60 );
nand NAND2_17535 ( P2_R1233_U469 , P2_U3501 , P2_R1233_U58 );
nand NAND2_17536 ( P2_R1233_U470 , P2_U3073 , P2_R1233_U56 );
nand NAND2_17537 ( P2_R1233_U471 , P2_U3498 , P2_R1233_U57 );
nand NAND2_17538 ( P2_R1233_U472 , P2_R1233_U471 , P2_R1233_U470 );
nand NAND2_17539 ( P2_R1233_U473 , P2_R1233_U361 , P2_R1233_U92 );
nand NAND2_17540 ( P2_R1233_U474 , P2_R1233_U472 , P2_R1233_U262 );
nand NAND2_17541 ( P2_R1233_U475 , P2_U3074 , P2_R1233_U73 );
nand NAND2_17542 ( P2_R1233_U476 , P2_U3495 , P2_R1233_U74 );
nand NAND2_17543 ( P2_R1233_U477 , P2_U3074 , P2_R1233_U73 );
nand NAND2_17544 ( P2_R1233_U478 , P2_U3495 , P2_R1233_U74 );
nand NAND2_17545 ( P2_R1233_U479 , P2_R1233_U478 , P2_R1233_U477 );
nand NAND2_17546 ( P2_R1233_U480 , P2_R1233_U163 , P2_R1233_U164 );
nand NAND2_17547 ( P2_R1233_U481 , P2_R1233_U258 , P2_R1233_U479 );
nand NAND2_17548 ( P2_R1233_U482 , P2_U3079 , P2_R1233_U71 );
nand NAND2_17549 ( P2_R1233_U483 , P2_U3492 , P2_R1233_U72 );
nand NAND2_17550 ( P2_R1233_U484 , P2_U3079 , P2_R1233_U71 );
nand NAND2_17551 ( P2_R1233_U485 , P2_U3492 , P2_R1233_U72 );
nand NAND2_17552 ( P2_R1233_U486 , P2_R1233_U485 , P2_R1233_U484 );
nand NAND2_17553 ( P2_R1233_U487 , P2_R1233_U165 , P2_R1233_U166 );
nand NAND2_17554 ( P2_R1233_U488 , P2_R1233_U254 , P2_R1233_U486 );
nand NAND2_17555 ( P2_R1233_U489 , P2_U3080 , P2_R1233_U69 );
nand NAND2_17556 ( P2_R1233_U490 , P2_U3489 , P2_R1233_U70 );
nand NAND2_17557 ( P2_R1233_U491 , P2_U3072 , P2_R1233_U64 );
nand NAND2_17558 ( P2_R1233_U492 , P2_U3486 , P2_R1233_U65 );
nand NAND2_17559 ( P2_R1233_U493 , P2_R1233_U492 , P2_R1233_U491 );
nand NAND2_17560 ( P2_R1233_U494 , P2_R1233_U362 , P2_R1233_U93 );
nand NAND2_17561 ( P2_R1233_U495 , P2_R1233_U493 , P2_R1233_U338 );
nand NAND2_17562 ( P2_R1233_U496 , P2_U3063 , P2_R1233_U66 );
nand NAND2_17563 ( P2_R1233_U497 , P2_U3483 , P2_R1233_U67 );
nand NAND2_17564 ( P2_R1233_U498 , P2_R1233_U497 , P2_R1233_U496 );
nand NAND2_17565 ( P2_R1233_U499 , P2_R1233_U363 , P2_R1233_U167 );
nand NAND2_17566 ( P2_R1233_U500 , P2_R1233_U244 , P2_R1233_U498 );
nand NAND2_17567 ( P2_R1233_U501 , P2_U3062 , P2_R1233_U61 );
nand NAND2_17568 ( P2_R1233_U502 , P2_U3480 , P2_R1233_U62 );
nand NAND2_17569 ( P2_R1233_U503 , P2_U3077 , P2_R1233_U29 );
nand NAND2_17570 ( P2_R1233_U504 , P2_U3448 , P2_R1233_U30 );
and AND2_17571 ( P2_R1176_U4 , P2_R1176_U211 , P2_R1176_U210 );
and AND2_17572 ( P2_R1176_U5 , P2_R1176_U224 , P2_R1176_U223 );
and AND2_17573 ( P2_R1176_U6 , P2_R1176_U256 , P2_R1176_U255 );
and AND2_17574 ( P2_R1176_U7 , P2_R1176_U274 , P2_R1176_U273 );
and AND2_17575 ( P2_R1176_U8 , P2_R1176_U286 , P2_R1176_U285 );
and AND2_17576 ( P2_R1176_U9 , P2_R1176_U344 , P2_R1176_U341 );
and AND2_17577 ( P2_R1176_U10 , P2_R1176_U335 , P2_R1176_U332 );
and AND2_17578 ( P2_R1176_U11 , P2_R1176_U328 , P2_R1176_U325 );
and AND2_17579 ( P2_R1176_U12 , P2_R1176_U319 , P2_R1176_U316 );
and AND2_17580 ( P2_R1176_U13 , P2_R1176_U247 , P2_R1176_U244 );
and AND2_17581 ( P2_R1176_U14 , P2_R1176_U240 , P2_R1176_U237 );
not NOT1_17582 ( P2_R1176_U15 , P2_U3214 );
not NOT1_17583 ( P2_R1176_U16 , P2_U3207 );
nand NAND2_17584 ( P2_R1176_U17 , P2_U3207 , P2_R1176_U56 );
not NOT1_17585 ( P2_R1176_U18 , P2_U3206 );
not NOT1_17586 ( P2_R1176_U19 , P2_U3211 );
nand NAND2_17587 ( P2_R1176_U20 , P2_U3211 , P2_R1176_U58 );
not NOT1_17588 ( P2_R1176_U21 , P2_U3210 );
not NOT1_17589 ( P2_R1176_U22 , P2_U3213 );
not NOT1_17590 ( P2_R1176_U23 , P2_U3212 );
not NOT1_17591 ( P2_R1176_U24 , P2_U3209 );
not NOT1_17592 ( P2_R1176_U25 , P2_U3208 );
not NOT1_17593 ( P2_R1176_U26 , P2_U3205 );
not NOT1_17594 ( P2_R1176_U27 , P2_U3204 );
nand NAND2_17595 ( P2_R1176_U28 , P2_R1176_U221 , P2_R1176_U220 );
nand NAND2_17596 ( P2_R1176_U29 , P2_R1176_U208 , P2_R1176_U207 );
not NOT1_17597 ( P2_R1176_U30 , P2_U3186 );
not NOT1_17598 ( P2_R1176_U31 , P2_U3187 );
not NOT1_17599 ( P2_R1176_U32 , P2_U3188 );
not NOT1_17600 ( P2_R1176_U33 , P2_U3189 );
not NOT1_17601 ( P2_R1176_U34 , P2_U3197 );
nand NAND2_17602 ( P2_R1176_U35 , P2_U3197 , P2_R1176_U69 );
not NOT1_17603 ( P2_R1176_U36 , P2_U3196 );
not NOT1_17604 ( P2_R1176_U37 , P2_U3203 );
not NOT1_17605 ( P2_R1176_U38 , P2_U3201 );
not NOT1_17606 ( P2_R1176_U39 , P2_U3202 );
nand NAND2_17607 ( P2_R1176_U40 , P2_U3202 , P2_R1176_U72 );
not NOT1_17608 ( P2_R1176_U41 , P2_U3200 );
not NOT1_17609 ( P2_R1176_U42 , P2_U3199 );
not NOT1_17610 ( P2_R1176_U43 , P2_U3198 );
not NOT1_17611 ( P2_R1176_U44 , P2_U3195 );
not NOT1_17612 ( P2_R1176_U45 , P2_U3193 );
not NOT1_17613 ( P2_R1176_U46 , P2_U3194 );
nand NAND2_17614 ( P2_R1176_U47 , P2_U3194 , P2_R1176_U78 );
not NOT1_17615 ( P2_R1176_U48 , P2_U3192 );
not NOT1_17616 ( P2_R1176_U49 , P2_U3191 );
not NOT1_17617 ( P2_R1176_U50 , P2_U3190 );
nand NAND2_17618 ( P2_R1176_U51 , P2_U3187 , P2_R1176_U67 );
nand NAND2_17619 ( P2_R1176_U52 , P2_R1176_U47 , P2_R1176_U321 );
nand NAND2_17620 ( P2_R1176_U53 , P2_R1176_U271 , P2_R1176_U270 );
nand NAND2_17621 ( P2_R1176_U54 , P2_R1176_U40 , P2_R1176_U337 );
nand NAND2_17622 ( P2_R1176_U55 , P2_R1176_U366 , P2_R1176_U365 );
nand NAND2_17623 ( P2_R1176_U56 , P2_R1176_U395 , P2_R1176_U394 );
nand NAND2_17624 ( P2_R1176_U57 , P2_R1176_U392 , P2_R1176_U391 );
nand NAND2_17625 ( P2_R1176_U58 , P2_R1176_U386 , P2_R1176_U385 );
nand NAND2_17626 ( P2_R1176_U59 , P2_R1176_U383 , P2_R1176_U382 );
nand NAND2_17627 ( P2_R1176_U60 , P2_R1176_U377 , P2_R1176_U376 );
nand NAND2_17628 ( P2_R1176_U61 , P2_R1176_U380 , P2_R1176_U379 );
nand NAND2_17629 ( P2_R1176_U62 , P2_R1176_U374 , P2_R1176_U373 );
nand NAND2_17630 ( P2_R1176_U63 , P2_R1176_U389 , P2_R1176_U388 );
nand NAND2_17631 ( P2_R1176_U64 , P2_R1176_U398 , P2_R1176_U397 );
nand NAND2_17632 ( P2_R1176_U65 , P2_R1176_U438 , P2_R1176_U437 );
nand NAND2_17633 ( P2_R1176_U66 , P2_R1176_U483 , P2_R1176_U482 );
nand NAND2_17634 ( P2_R1176_U67 , P2_R1176_U486 , P2_R1176_U485 );
nand NAND2_17635 ( P2_R1176_U68 , P2_R1176_U489 , P2_R1176_U488 );
nand NAND2_17636 ( P2_R1176_U69 , P2_R1176_U462 , P2_R1176_U461 );
nand NAND2_17637 ( P2_R1176_U70 , P2_R1176_U459 , P2_R1176_U458 );
nand NAND2_17638 ( P2_R1176_U71 , P2_R1176_U441 , P2_R1176_U440 );
nand NAND2_17639 ( P2_R1176_U72 , P2_R1176_U450 , P2_R1176_U449 );
nand NAND2_17640 ( P2_R1176_U73 , P2_R1176_U444 , P2_R1176_U443 );
nand NAND2_17641 ( P2_R1176_U74 , P2_R1176_U447 , P2_R1176_U446 );
nand NAND2_17642 ( P2_R1176_U75 , P2_R1176_U453 , P2_R1176_U452 );
nand NAND2_17643 ( P2_R1176_U76 , P2_R1176_U456 , P2_R1176_U455 );
nand NAND2_17644 ( P2_R1176_U77 , P2_R1176_U465 , P2_R1176_U464 );
nand NAND2_17645 ( P2_R1176_U78 , P2_R1176_U474 , P2_R1176_U473 );
nand NAND2_17646 ( P2_R1176_U79 , P2_R1176_U468 , P2_R1176_U467 );
nand NAND2_17647 ( P2_R1176_U80 , P2_R1176_U471 , P2_R1176_U470 );
nand NAND2_17648 ( P2_R1176_U81 , P2_R1176_U477 , P2_R1176_U476 );
nand NAND2_17649 ( P2_R1176_U82 , P2_R1176_U480 , P2_R1176_U479 );
nand NAND2_17650 ( P2_R1176_U83 , P2_R1176_U495 , P2_R1176_U494 );
nand NAND2_17651 ( P2_R1176_U84 , P2_R1176_U602 , P2_R1176_U601 );
nand NAND2_17652 ( P2_R1176_U85 , P2_R1176_U401 , P2_R1176_U400 );
nand NAND2_17653 ( P2_R1176_U86 , P2_R1176_U408 , P2_R1176_U407 );
nand NAND2_17654 ( P2_R1176_U87 , P2_R1176_U415 , P2_R1176_U414 );
nand NAND2_17655 ( P2_R1176_U88 , P2_R1176_U422 , P2_R1176_U421 );
nand NAND2_17656 ( P2_R1176_U89 , P2_R1176_U429 , P2_R1176_U428 );
nand NAND2_17657 ( P2_R1176_U90 , P2_R1176_U436 , P2_R1176_U435 );
nand NAND2_17658 ( P2_R1176_U91 , P2_R1176_U498 , P2_R1176_U497 );
nand NAND2_17659 ( P2_R1176_U92 , P2_R1176_U505 , P2_R1176_U504 );
nand NAND2_17660 ( P2_R1176_U93 , P2_R1176_U512 , P2_R1176_U511 );
nand NAND2_17661 ( P2_R1176_U94 , P2_R1176_U517 , P2_R1176_U516 );
nand NAND2_17662 ( P2_R1176_U95 , P2_R1176_U524 , P2_R1176_U523 );
nand NAND2_17663 ( P2_R1176_U96 , P2_R1176_U531 , P2_R1176_U530 );
nand NAND2_17664 ( P2_R1176_U97 , P2_R1176_U538 , P2_R1176_U537 );
nand NAND2_17665 ( P2_R1176_U98 , P2_R1176_U545 , P2_R1176_U544 );
nand NAND2_17666 ( P2_R1176_U99 , P2_R1176_U550 , P2_R1176_U549 );
nand NAND2_17667 ( P2_R1176_U100 , P2_R1176_U557 , P2_R1176_U556 );
nand NAND2_17668 ( P2_R1176_U101 , P2_R1176_U564 , P2_R1176_U563 );
nand NAND2_17669 ( P2_R1176_U102 , P2_R1176_U571 , P2_R1176_U570 );
nand NAND2_17670 ( P2_R1176_U103 , P2_R1176_U578 , P2_R1176_U577 );
nand NAND2_17671 ( P2_R1176_U104 , P2_R1176_U585 , P2_R1176_U584 );
nand NAND2_17672 ( P2_R1176_U105 , P2_R1176_U590 , P2_R1176_U589 );
nand NAND2_17673 ( P2_R1176_U106 , P2_R1176_U597 , P2_R1176_U596 );
and AND2_17674 ( P2_R1176_U107 , P2_R1176_U214 , P2_R1176_U213 );
and AND2_17675 ( P2_R1176_U108 , P2_R1176_U228 , P2_R1176_U227 );
and AND3_17676 ( P2_R1176_U109 , P2_R1176_U410 , P2_R1176_U409 , P2_R1176_U17 );
and AND2_17677 ( P2_R1176_U110 , P2_R1176_U239 , P2_R1176_U5 );
and AND3_17678 ( P2_R1176_U111 , P2_R1176_U431 , P2_R1176_U430 , P2_R1176_U20 );
and AND2_17679 ( P2_R1176_U112 , P2_R1176_U246 , P2_R1176_U4 );
and AND2_17680 ( P2_R1176_U113 , P2_R1176_U260 , P2_R1176_U6 );
and AND2_17681 ( P2_R1176_U114 , P2_R1176_U258 , P2_R1176_U196 );
and AND2_17682 ( P2_R1176_U115 , P2_R1176_U278 , P2_R1176_U277 );
and AND2_17683 ( P2_R1176_U116 , P2_R1176_U290 , P2_R1176_U8 );
and AND2_17684 ( P2_R1176_U117 , P2_R1176_U288 , P2_R1176_U197 );
and AND2_17685 ( P2_R1176_U118 , P2_R1176_U306 , P2_R1176_U192 );
and AND2_17686 ( P2_R1176_U119 , P2_R1176_U364 , P2_R1176_U51 );
and AND2_17687 ( P2_R1176_U120 , P2_R1176_U311 , P2_R1176_U306 );
and AND2_17688 ( P2_R1176_U121 , P2_R1176_U361 , P2_R1176_U310 );
nand NAND2_17689 ( P2_R1176_U122 , P2_R1176_U492 , P2_R1176_U491 );
and AND2_17690 ( P2_R1176_U123 , P2_R1176_U357 , P2_R1176_U51 );
and AND3_17691 ( P2_R1176_U124 , P2_R1176_U507 , P2_R1176_U506 , P2_R1176_U198 );
and AND2_17692 ( P2_R1176_U125 , P2_R1176_U201 , P2_R1176_U198 );
and AND2_17693 ( P2_R1176_U126 , P2_R1176_U318 , P2_R1176_U192 );
and AND3_17694 ( P2_R1176_U127 , P2_R1176_U533 , P2_R1176_U532 , P2_R1176_U197 );
and AND2_17695 ( P2_R1176_U128 , P2_R1176_U327 , P2_R1176_U8 );
and AND3_17696 ( P2_R1176_U129 , P2_R1176_U559 , P2_R1176_U558 , P2_R1176_U35 );
and AND2_17697 ( P2_R1176_U130 , P2_R1176_U334 , P2_R1176_U7 );
and AND3_17698 ( P2_R1176_U131 , P2_R1176_U580 , P2_R1176_U579 , P2_R1176_U196 );
and AND2_17699 ( P2_R1176_U132 , P2_R1176_U343 , P2_R1176_U6 );
nand NAND2_17700 ( P2_R1176_U133 , P2_R1176_U599 , P2_R1176_U598 );
not NOT1_17701 ( P2_R1176_U134 , P2_U3477 );
and AND2_17702 ( P2_R1176_U135 , P2_R1176_U369 , P2_R1176_U368 );
not NOT1_17703 ( P2_R1176_U136 , P2_U3462 );
not NOT1_17704 ( P2_R1176_U137 , P2_U3448 );
not NOT1_17705 ( P2_R1176_U138 , P2_U3453 );
not NOT1_17706 ( P2_R1176_U139 , P2_U3459 );
not NOT1_17707 ( P2_R1176_U140 , P2_U3456 );
not NOT1_17708 ( P2_R1176_U141 , P2_U3465 );
not NOT1_17709 ( P2_R1176_U142 , P2_U3471 );
not NOT1_17710 ( P2_R1176_U143 , P2_U3468 );
not NOT1_17711 ( P2_R1176_U144 , P2_U3474 );
nand NAND2_17712 ( P2_R1176_U145 , P2_R1176_U233 , P2_R1176_U232 );
and AND2_17713 ( P2_R1176_U146 , P2_R1176_U403 , P2_R1176_U402 );
nand NAND2_17714 ( P2_R1176_U147 , P2_R1176_U108 , P2_R1176_U229 );
and AND2_17715 ( P2_R1176_U148 , P2_R1176_U417 , P2_R1176_U416 );
nand NAND3_17716 ( P2_R1176_U149 , P2_R1176_U217 , P2_R1176_U194 , P2_R1176_U355 );
and AND2_17717 ( P2_R1176_U150 , P2_R1176_U424 , P2_R1176_U423 );
nand NAND2_17718 ( P2_R1176_U151 , P2_R1176_U107 , P2_R1176_U215 );
not NOT1_17719 ( P2_R1176_U152 , P2_U3969 );
not NOT1_17720 ( P2_R1176_U153 , P2_U3480 );
not NOT1_17721 ( P2_R1176_U154 , P2_U3489 );
not NOT1_17722 ( P2_R1176_U155 , P2_U3486 );
not NOT1_17723 ( P2_R1176_U156 , P2_U3483 );
not NOT1_17724 ( P2_R1176_U157 , P2_U3492 );
not NOT1_17725 ( P2_R1176_U158 , P2_U3495 );
not NOT1_17726 ( P2_R1176_U159 , P2_U3501 );
not NOT1_17727 ( P2_R1176_U160 , P2_U3498 );
not NOT1_17728 ( P2_R1176_U161 , P2_U3504 );
not NOT1_17729 ( P2_R1176_U162 , P2_U3975 );
not NOT1_17730 ( P2_R1176_U163 , P2_U3976 );
not NOT1_17731 ( P2_R1176_U164 , P2_U3506 );
not NOT1_17732 ( P2_R1176_U165 , P2_U3974 );
not NOT1_17733 ( P2_R1176_U166 , P2_U3973 );
not NOT1_17734 ( P2_R1176_U167 , P2_U3971 );
not NOT1_17735 ( P2_R1176_U168 , P2_U3970 );
not NOT1_17736 ( P2_R1176_U169 , P2_U3972 );
not NOT1_17737 ( P2_R1176_U170 , P2_U3185 );
not NOT1_17738 ( P2_R1176_U171 , P2_U3968 );
and AND2_17739 ( P2_R1176_U172 , P2_R1176_U500 , P2_R1176_U499 );
nand NAND2_17740 ( P2_R1176_U173 , P2_R1176_U123 , P2_R1176_U307 );
nand NAND2_17741 ( P2_R1176_U174 , P2_R1176_U201 , P2_R1176_U312 );
nand NAND2_17742 ( P2_R1176_U175 , P2_R1176_U301 , P2_R1176_U300 );
and AND2_17743 ( P2_R1176_U176 , P2_R1176_U519 , P2_R1176_U518 );
nand NAND2_17744 ( P2_R1176_U177 , P2_R1176_U297 , P2_R1176_U296 );
and AND2_17745 ( P2_R1176_U178 , P2_R1176_U526 , P2_R1176_U525 );
nand NAND2_17746 ( P2_R1176_U179 , P2_R1176_U293 , P2_R1176_U292 );
and AND2_17747 ( P2_R1176_U180 , P2_R1176_U540 , P2_R1176_U539 );
nand NAND2_17748 ( P2_R1176_U181 , P2_R1176_U204 , P2_R1176_U203 );
nand NAND2_17749 ( P2_R1176_U182 , P2_R1176_U283 , P2_R1176_U282 );
and AND2_17750 ( P2_R1176_U183 , P2_R1176_U552 , P2_R1176_U551 );
nand NAND2_17751 ( P2_R1176_U184 , P2_R1176_U115 , P2_R1176_U279 );
and AND2_17752 ( P2_R1176_U185 , P2_R1176_U566 , P2_R1176_U565 );
nand NAND2_17753 ( P2_R1176_U186 , P2_R1176_U267 , P2_R1176_U266 );
and AND2_17754 ( P2_R1176_U187 , P2_R1176_U573 , P2_R1176_U572 );
nand NAND2_17755 ( P2_R1176_U188 , P2_R1176_U263 , P2_R1176_U262 );
nand NAND2_17756 ( P2_R1176_U189 , P2_R1176_U253 , P2_R1176_U252 );
and AND2_17757 ( P2_R1176_U190 , P2_R1176_U592 , P2_R1176_U591 );
nand NAND3_17758 ( P2_R1176_U191 , P2_R1176_U249 , P2_R1176_U193 , P2_R1176_U360 );
nand NAND2_17759 ( P2_R1176_U192 , P2_R1176_U359 , P2_R1176_U358 );
nand NAND2_17760 ( P2_R1176_U193 , P2_R1176_U55 , P2_R1176_U145 );
nand NAND2_17761 ( P2_R1176_U194 , P2_R1176_U62 , P2_R1176_U151 );
not NOT1_17762 ( P2_R1176_U195 , P2_R1176_U20 );
nand NAND2_17763 ( P2_R1176_U196 , P2_U3201 , P2_R1176_U74 );
nand NAND2_17764 ( P2_R1176_U197 , P2_U3193 , P2_R1176_U80 );
nand NAND2_17765 ( P2_R1176_U198 , P2_U3188 , P2_R1176_U66 );
not NOT1_17766 ( P2_R1176_U199 , P2_R1176_U40 );
not NOT1_17767 ( P2_R1176_U200 , P2_R1176_U47 );
nand NAND2_17768 ( P2_R1176_U201 , P2_U3189 , P2_R1176_U68 );
nand NAND2_17769 ( P2_R1176_U202 , P2_R1176_U378 , P2_R1176_U15 );
nand NAND2_17770 ( P2_R1176_U203 , P2_U3213 , P2_R1176_U202 );
nand NAND2_17771 ( P2_R1176_U204 , P2_U3214 , P2_R1176_U60 );
not NOT1_17772 ( P2_R1176_U205 , P2_R1176_U181 );
nand NAND2_17773 ( P2_R1176_U206 , P2_R1176_U381 , P2_R1176_U23 );
nand NAND2_17774 ( P2_R1176_U207 , P2_R1176_U206 , P2_R1176_U181 );
nand NAND2_17775 ( P2_R1176_U208 , P2_U3212 , P2_R1176_U61 );
not NOT1_17776 ( P2_R1176_U209 , P2_R1176_U29 );
nand NAND2_17777 ( P2_R1176_U210 , P2_R1176_U384 , P2_R1176_U21 );
nand NAND2_17778 ( P2_R1176_U211 , P2_R1176_U387 , P2_R1176_U19 );
nand NAND2_17779 ( P2_R1176_U212 , P2_R1176_U21 , P2_R1176_U20 );
nand NAND2_17780 ( P2_R1176_U213 , P2_R1176_U59 , P2_R1176_U212 );
nand NAND2_17781 ( P2_R1176_U214 , P2_U3210 , P2_R1176_U195 );
nand NAND2_17782 ( P2_R1176_U215 , P2_R1176_U4 , P2_R1176_U29 );
not NOT1_17783 ( P2_R1176_U216 , P2_R1176_U151 );
nand NAND2_17784 ( P2_R1176_U217 , P2_U3209 , P2_R1176_U151 );
not NOT1_17785 ( P2_R1176_U218 , P2_R1176_U149 );
nand NAND2_17786 ( P2_R1176_U219 , P2_R1176_U390 , P2_R1176_U25 );
nand NAND2_17787 ( P2_R1176_U220 , P2_R1176_U219 , P2_R1176_U149 );
nand NAND2_17788 ( P2_R1176_U221 , P2_U3208 , P2_R1176_U63 );
not NOT1_17789 ( P2_R1176_U222 , P2_R1176_U28 );
nand NAND2_17790 ( P2_R1176_U223 , P2_R1176_U393 , P2_R1176_U18 );
nand NAND2_17791 ( P2_R1176_U224 , P2_R1176_U396 , P2_R1176_U16 );
not NOT1_17792 ( P2_R1176_U225 , P2_R1176_U17 );
nand NAND2_17793 ( P2_R1176_U226 , P2_R1176_U18 , P2_R1176_U17 );
nand NAND2_17794 ( P2_R1176_U227 , P2_R1176_U57 , P2_R1176_U226 );
nand NAND2_17795 ( P2_R1176_U228 , P2_U3206 , P2_R1176_U225 );
nand NAND2_17796 ( P2_R1176_U229 , P2_R1176_U5 , P2_R1176_U28 );
not NOT1_17797 ( P2_R1176_U230 , P2_R1176_U147 );
nand NAND2_17798 ( P2_R1176_U231 , P2_R1176_U399 , P2_R1176_U26 );
nand NAND2_17799 ( P2_R1176_U232 , P2_R1176_U231 , P2_R1176_U147 );
nand NAND2_17800 ( P2_R1176_U233 , P2_U3205 , P2_R1176_U64 );
not NOT1_17801 ( P2_R1176_U234 , P2_R1176_U145 );
nand NAND2_17802 ( P2_R1176_U235 , P2_R1176_U396 , P2_R1176_U16 );
nand NAND2_17803 ( P2_R1176_U236 , P2_R1176_U235 , P2_R1176_U28 );
nand NAND2_17804 ( P2_R1176_U237 , P2_R1176_U109 , P2_R1176_U236 );
nand NAND2_17805 ( P2_R1176_U238 , P2_R1176_U222 , P2_R1176_U17 );
nand NAND2_17806 ( P2_R1176_U239 , P2_U3206 , P2_R1176_U57 );
nand NAND2_17807 ( P2_R1176_U240 , P2_R1176_U110 , P2_R1176_U238 );
nand NAND2_17808 ( P2_R1176_U241 , P2_R1176_U396 , P2_R1176_U16 );
nand NAND2_17809 ( P2_R1176_U242 , P2_R1176_U387 , P2_R1176_U19 );
nand NAND2_17810 ( P2_R1176_U243 , P2_R1176_U242 , P2_R1176_U29 );
nand NAND2_17811 ( P2_R1176_U244 , P2_R1176_U111 , P2_R1176_U243 );
nand NAND2_17812 ( P2_R1176_U245 , P2_R1176_U209 , P2_R1176_U20 );
nand NAND2_17813 ( P2_R1176_U246 , P2_U3210 , P2_R1176_U59 );
nand NAND2_17814 ( P2_R1176_U247 , P2_R1176_U112 , P2_R1176_U245 );
nand NAND2_17815 ( P2_R1176_U248 , P2_R1176_U387 , P2_R1176_U19 );
nand NAND2_17816 ( P2_R1176_U249 , P2_U3204 , P2_R1176_U145 );
not NOT1_17817 ( P2_R1176_U250 , P2_R1176_U191 );
nand NAND2_17818 ( P2_R1176_U251 , P2_R1176_U442 , P2_R1176_U37 );
nand NAND2_17819 ( P2_R1176_U252 , P2_R1176_U251 , P2_R1176_U191 );
nand NAND2_17820 ( P2_R1176_U253 , P2_U3203 , P2_R1176_U71 );
not NOT1_17821 ( P2_R1176_U254 , P2_R1176_U189 );
nand NAND2_17822 ( P2_R1176_U255 , P2_R1176_U445 , P2_R1176_U41 );
nand NAND2_17823 ( P2_R1176_U256 , P2_R1176_U448 , P2_R1176_U38 );
nand NAND2_17824 ( P2_R1176_U257 , P2_R1176_U199 , P2_R1176_U6 );
nand NAND2_17825 ( P2_R1176_U258 , P2_U3200 , P2_R1176_U73 );
nand NAND2_17826 ( P2_R1176_U259 , P2_R1176_U114 , P2_R1176_U257 );
nand NAND2_17827 ( P2_R1176_U260 , P2_R1176_U451 , P2_R1176_U39 );
nand NAND2_17828 ( P2_R1176_U261 , P2_R1176_U445 , P2_R1176_U41 );
nand NAND2_17829 ( P2_R1176_U262 , P2_R1176_U113 , P2_R1176_U189 );
nand NAND2_17830 ( P2_R1176_U263 , P2_R1176_U261 , P2_R1176_U259 );
not NOT1_17831 ( P2_R1176_U264 , P2_R1176_U188 );
nand NAND2_17832 ( P2_R1176_U265 , P2_R1176_U454 , P2_R1176_U42 );
nand NAND2_17833 ( P2_R1176_U266 , P2_R1176_U265 , P2_R1176_U188 );
nand NAND2_17834 ( P2_R1176_U267 , P2_U3199 , P2_R1176_U75 );
not NOT1_17835 ( P2_R1176_U268 , P2_R1176_U186 );
nand NAND2_17836 ( P2_R1176_U269 , P2_R1176_U457 , P2_R1176_U43 );
nand NAND2_17837 ( P2_R1176_U270 , P2_R1176_U269 , P2_R1176_U186 );
nand NAND2_17838 ( P2_R1176_U271 , P2_U3198 , P2_R1176_U76 );
not NOT1_17839 ( P2_R1176_U272 , P2_R1176_U53 );
nand NAND2_17840 ( P2_R1176_U273 , P2_R1176_U460 , P2_R1176_U36 );
nand NAND2_17841 ( P2_R1176_U274 , P2_R1176_U463 , P2_R1176_U34 );
not NOT1_17842 ( P2_R1176_U275 , P2_R1176_U35 );
nand NAND2_17843 ( P2_R1176_U276 , P2_R1176_U36 , P2_R1176_U35 );
nand NAND2_17844 ( P2_R1176_U277 , P2_R1176_U70 , P2_R1176_U276 );
nand NAND2_17845 ( P2_R1176_U278 , P2_U3196 , P2_R1176_U275 );
nand NAND2_17846 ( P2_R1176_U279 , P2_R1176_U7 , P2_R1176_U53 );
not NOT1_17847 ( P2_R1176_U280 , P2_R1176_U184 );
nand NAND2_17848 ( P2_R1176_U281 , P2_R1176_U466 , P2_R1176_U44 );
nand NAND2_17849 ( P2_R1176_U282 , P2_R1176_U281 , P2_R1176_U184 );
nand NAND2_17850 ( P2_R1176_U283 , P2_U3195 , P2_R1176_U77 );
not NOT1_17851 ( P2_R1176_U284 , P2_R1176_U182 );
nand NAND2_17852 ( P2_R1176_U285 , P2_R1176_U469 , P2_R1176_U48 );
nand NAND2_17853 ( P2_R1176_U286 , P2_R1176_U472 , P2_R1176_U45 );
nand NAND2_17854 ( P2_R1176_U287 , P2_R1176_U200 , P2_R1176_U8 );
nand NAND2_17855 ( P2_R1176_U288 , P2_U3192 , P2_R1176_U79 );
nand NAND2_17856 ( P2_R1176_U289 , P2_R1176_U117 , P2_R1176_U287 );
nand NAND2_17857 ( P2_R1176_U290 , P2_R1176_U475 , P2_R1176_U46 );
nand NAND2_17858 ( P2_R1176_U291 , P2_R1176_U469 , P2_R1176_U48 );
nand NAND2_17859 ( P2_R1176_U292 , P2_R1176_U116 , P2_R1176_U182 );
nand NAND2_17860 ( P2_R1176_U293 , P2_R1176_U291 , P2_R1176_U289 );
not NOT1_17861 ( P2_R1176_U294 , P2_R1176_U179 );
nand NAND2_17862 ( P2_R1176_U295 , P2_R1176_U478 , P2_R1176_U49 );
nand NAND2_17863 ( P2_R1176_U296 , P2_R1176_U295 , P2_R1176_U179 );
nand NAND2_17864 ( P2_R1176_U297 , P2_U3191 , P2_R1176_U81 );
not NOT1_17865 ( P2_R1176_U298 , P2_R1176_U177 );
nand NAND2_17866 ( P2_R1176_U299 , P2_R1176_U481 , P2_R1176_U50 );
nand NAND2_17867 ( P2_R1176_U300 , P2_R1176_U299 , P2_R1176_U177 );
nand NAND2_17868 ( P2_R1176_U301 , P2_U3190 , P2_R1176_U82 );
not NOT1_17869 ( P2_R1176_U302 , P2_R1176_U175 );
nand NAND2_17870 ( P2_R1176_U303 , P2_R1176_U484 , P2_R1176_U32 );
nand NAND2_17871 ( P2_R1176_U304 , P2_R1176_U201 , P2_R1176_U198 );
not NOT1_17872 ( P2_R1176_U305 , P2_R1176_U51 );
nand NAND2_17873 ( P2_R1176_U306 , P2_R1176_U490 , P2_R1176_U33 );
nand NAND2_17874 ( P2_R1176_U307 , P2_R1176_U118 , P2_R1176_U175 );
not NOT1_17875 ( P2_R1176_U308 , P2_R1176_U173 );
nand NAND2_17876 ( P2_R1176_U309 , P2_R1176_U439 , P2_R1176_U30 );
nand NAND2_17877 ( P2_R1176_U310 , P2_U3186 , P2_R1176_U65 );
nand NAND2_17878 ( P2_R1176_U311 , P2_R1176_U439 , P2_R1176_U30 );
nand NAND2_17879 ( P2_R1176_U312 , P2_R1176_U306 , P2_R1176_U175 );
not NOT1_17880 ( P2_R1176_U313 , P2_R1176_U174 );
nand NAND2_17881 ( P2_R1176_U314 , P2_R1176_U484 , P2_R1176_U32 );
nand NAND2_17882 ( P2_R1176_U315 , P2_R1176_U314 , P2_R1176_U174 );
nand NAND2_17883 ( P2_R1176_U316 , P2_R1176_U124 , P2_R1176_U315 );
nand NAND2_17884 ( P2_R1176_U317 , P2_R1176_U125 , P2_R1176_U312 );
nand NAND2_17885 ( P2_R1176_U318 , P2_U3187 , P2_R1176_U67 );
nand NAND2_17886 ( P2_R1176_U319 , P2_R1176_U126 , P2_R1176_U317 );
nand NAND2_17887 ( P2_R1176_U320 , P2_R1176_U484 , P2_R1176_U32 );
nand NAND2_17888 ( P2_R1176_U321 , P2_R1176_U290 , P2_R1176_U182 );
not NOT1_17889 ( P2_R1176_U322 , P2_R1176_U52 );
nand NAND2_17890 ( P2_R1176_U323 , P2_R1176_U472 , P2_R1176_U45 );
nand NAND2_17891 ( P2_R1176_U324 , P2_R1176_U323 , P2_R1176_U52 );
nand NAND2_17892 ( P2_R1176_U325 , P2_R1176_U127 , P2_R1176_U324 );
nand NAND2_17893 ( P2_R1176_U326 , P2_R1176_U322 , P2_R1176_U197 );
nand NAND2_17894 ( P2_R1176_U327 , P2_U3192 , P2_R1176_U79 );
nand NAND2_17895 ( P2_R1176_U328 , P2_R1176_U128 , P2_R1176_U326 );
nand NAND2_17896 ( P2_R1176_U329 , P2_R1176_U472 , P2_R1176_U45 );
nand NAND2_17897 ( P2_R1176_U330 , P2_R1176_U463 , P2_R1176_U34 );
nand NAND2_17898 ( P2_R1176_U331 , P2_R1176_U330 , P2_R1176_U53 );
nand NAND2_17899 ( P2_R1176_U332 , P2_R1176_U129 , P2_R1176_U331 );
nand NAND2_17900 ( P2_R1176_U333 , P2_R1176_U272 , P2_R1176_U35 );
nand NAND2_17901 ( P2_R1176_U334 , P2_U3196 , P2_R1176_U70 );
nand NAND2_17902 ( P2_R1176_U335 , P2_R1176_U130 , P2_R1176_U333 );
nand NAND2_17903 ( P2_R1176_U336 , P2_R1176_U463 , P2_R1176_U34 );
nand NAND2_17904 ( P2_R1176_U337 , P2_R1176_U260 , P2_R1176_U189 );
not NOT1_17905 ( P2_R1176_U338 , P2_R1176_U54 );
nand NAND2_17906 ( P2_R1176_U339 , P2_R1176_U448 , P2_R1176_U38 );
nand NAND2_17907 ( P2_R1176_U340 , P2_R1176_U339 , P2_R1176_U54 );
nand NAND2_17908 ( P2_R1176_U341 , P2_R1176_U131 , P2_R1176_U340 );
nand NAND2_17909 ( P2_R1176_U342 , P2_R1176_U338 , P2_R1176_U196 );
nand NAND2_17910 ( P2_R1176_U343 , P2_U3200 , P2_R1176_U73 );
nand NAND2_17911 ( P2_R1176_U344 , P2_R1176_U132 , P2_R1176_U342 );
nand NAND2_17912 ( P2_R1176_U345 , P2_R1176_U448 , P2_R1176_U38 );
nand NAND2_17913 ( P2_R1176_U346 , P2_R1176_U241 , P2_R1176_U17 );
nand NAND2_17914 ( P2_R1176_U347 , P2_R1176_U248 , P2_R1176_U20 );
nand NAND2_17915 ( P2_R1176_U348 , P2_R1176_U320 , P2_R1176_U198 );
nand NAND2_17916 ( P2_R1176_U349 , P2_R1176_U306 , P2_R1176_U201 );
nand NAND2_17917 ( P2_R1176_U350 , P2_R1176_U329 , P2_R1176_U197 );
nand NAND2_17918 ( P2_R1176_U351 , P2_R1176_U290 , P2_R1176_U47 );
nand NAND2_17919 ( P2_R1176_U352 , P2_R1176_U336 , P2_R1176_U35 );
nand NAND2_17920 ( P2_R1176_U353 , P2_R1176_U345 , P2_R1176_U196 );
nand NAND2_17921 ( P2_R1176_U354 , P2_R1176_U260 , P2_R1176_U40 );
nand NAND2_17922 ( P2_R1176_U355 , P2_U3209 , P2_R1176_U62 );
nand NAND3_17923 ( P2_R1176_U356 , P2_R1176_U357 , P2_R1176_U307 , P2_R1176_U119 );
nand NAND2_17924 ( P2_R1176_U357 , P2_R1176_U304 , P2_R1176_U192 );
nand NAND2_17925 ( P2_R1176_U358 , P2_R1176_U67 , P2_R1176_U303 );
nand NAND2_17926 ( P2_R1176_U359 , P2_U3187 , P2_R1176_U303 );
nand NAND2_17927 ( P2_R1176_U360 , P2_U3204 , P2_R1176_U55 );
nand NAND3_17928 ( P2_R1176_U361 , P2_R1176_U304 , P2_R1176_U192 , P2_R1176_U311 );
nand NAND3_17929 ( P2_R1176_U362 , P2_R1176_U175 , P2_R1176_U192 , P2_R1176_U120 );
nand NAND2_17930 ( P2_R1176_U363 , P2_R1176_U305 , P2_R1176_U311 );
nand NAND2_17931 ( P2_R1176_U364 , P2_U3186 , P2_R1176_U65 );
nand NAND2_17932 ( P2_R1176_U365 , P2_U3214 , P2_R1176_U134 );
nand NAND2_17933 ( P2_R1176_U366 , P2_U3477 , P2_R1176_U15 );
not NOT1_17934 ( P2_R1176_U367 , P2_R1176_U55 );
nand NAND2_17935 ( P2_R1176_U368 , P2_R1176_U367 , P2_U3204 );
nand NAND2_17936 ( P2_R1176_U369 , P2_R1176_U55 , P2_R1176_U27 );
nand NAND2_17937 ( P2_R1176_U370 , P2_R1176_U367 , P2_U3204 );
nand NAND2_17938 ( P2_R1176_U371 , P2_R1176_U55 , P2_R1176_U27 );
nand NAND2_17939 ( P2_R1176_U372 , P2_R1176_U371 , P2_R1176_U370 );
nand NAND2_17940 ( P2_R1176_U373 , P2_U3214 , P2_R1176_U136 );
nand NAND2_17941 ( P2_R1176_U374 , P2_U3462 , P2_R1176_U15 );
not NOT1_17942 ( P2_R1176_U375 , P2_R1176_U62 );
nand NAND2_17943 ( P2_R1176_U376 , P2_U3214 , P2_R1176_U137 );
nand NAND2_17944 ( P2_R1176_U377 , P2_U3448 , P2_R1176_U15 );
not NOT1_17945 ( P2_R1176_U378 , P2_R1176_U60 );
nand NAND2_17946 ( P2_R1176_U379 , P2_U3214 , P2_R1176_U138 );
nand NAND2_17947 ( P2_R1176_U380 , P2_U3453 , P2_R1176_U15 );
not NOT1_17948 ( P2_R1176_U381 , P2_R1176_U61 );
nand NAND2_17949 ( P2_R1176_U382 , P2_U3214 , P2_R1176_U139 );
nand NAND2_17950 ( P2_R1176_U383 , P2_U3459 , P2_R1176_U15 );
not NOT1_17951 ( P2_R1176_U384 , P2_R1176_U59 );
nand NAND2_17952 ( P2_R1176_U385 , P2_U3214 , P2_R1176_U140 );
nand NAND2_17953 ( P2_R1176_U386 , P2_U3456 , P2_R1176_U15 );
not NOT1_17954 ( P2_R1176_U387 , P2_R1176_U58 );
nand NAND2_17955 ( P2_R1176_U388 , P2_U3214 , P2_R1176_U141 );
nand NAND2_17956 ( P2_R1176_U389 , P2_U3465 , P2_R1176_U15 );
not NOT1_17957 ( P2_R1176_U390 , P2_R1176_U63 );
nand NAND2_17958 ( P2_R1176_U391 , P2_U3214 , P2_R1176_U142 );
nand NAND2_17959 ( P2_R1176_U392 , P2_U3471 , P2_R1176_U15 );
not NOT1_17960 ( P2_R1176_U393 , P2_R1176_U57 );
nand NAND2_17961 ( P2_R1176_U394 , P2_U3214 , P2_R1176_U143 );
nand NAND2_17962 ( P2_R1176_U395 , P2_U3468 , P2_R1176_U15 );
not NOT1_17963 ( P2_R1176_U396 , P2_R1176_U56 );
nand NAND2_17964 ( P2_R1176_U397 , P2_U3214 , P2_R1176_U144 );
nand NAND2_17965 ( P2_R1176_U398 , P2_U3474 , P2_R1176_U15 );
not NOT1_17966 ( P2_R1176_U399 , P2_R1176_U64 );
nand NAND2_17967 ( P2_R1176_U400 , P2_R1176_U135 , P2_R1176_U145 );
nand NAND2_17968 ( P2_R1176_U401 , P2_R1176_U234 , P2_R1176_U372 );
nand NAND2_17969 ( P2_R1176_U402 , P2_R1176_U399 , P2_U3205 );
nand NAND2_17970 ( P2_R1176_U403 , P2_R1176_U64 , P2_R1176_U26 );
nand NAND2_17971 ( P2_R1176_U404 , P2_R1176_U399 , P2_U3205 );
nand NAND2_17972 ( P2_R1176_U405 , P2_R1176_U64 , P2_R1176_U26 );
nand NAND2_17973 ( P2_R1176_U406 , P2_R1176_U405 , P2_R1176_U404 );
nand NAND2_17974 ( P2_R1176_U407 , P2_R1176_U146 , P2_R1176_U147 );
nand NAND2_17975 ( P2_R1176_U408 , P2_R1176_U230 , P2_R1176_U406 );
nand NAND2_17976 ( P2_R1176_U409 , P2_R1176_U393 , P2_U3206 );
nand NAND2_17977 ( P2_R1176_U410 , P2_R1176_U57 , P2_R1176_U18 );
nand NAND2_17978 ( P2_R1176_U411 , P2_R1176_U396 , P2_U3207 );
nand NAND2_17979 ( P2_R1176_U412 , P2_R1176_U56 , P2_R1176_U16 );
nand NAND2_17980 ( P2_R1176_U413 , P2_R1176_U412 , P2_R1176_U411 );
nand NAND2_17981 ( P2_R1176_U414 , P2_R1176_U346 , P2_R1176_U28 );
nand NAND2_17982 ( P2_R1176_U415 , P2_R1176_U413 , P2_R1176_U222 );
nand NAND2_17983 ( P2_R1176_U416 , P2_R1176_U390 , P2_U3208 );
nand NAND2_17984 ( P2_R1176_U417 , P2_R1176_U63 , P2_R1176_U25 );
nand NAND2_17985 ( P2_R1176_U418 , P2_R1176_U390 , P2_U3208 );
nand NAND2_17986 ( P2_R1176_U419 , P2_R1176_U63 , P2_R1176_U25 );
nand NAND2_17987 ( P2_R1176_U420 , P2_R1176_U419 , P2_R1176_U418 );
nand NAND2_17988 ( P2_R1176_U421 , P2_R1176_U148 , P2_R1176_U149 );
nand NAND2_17989 ( P2_R1176_U422 , P2_R1176_U218 , P2_R1176_U420 );
nand NAND2_17990 ( P2_R1176_U423 , P2_R1176_U375 , P2_U3209 );
nand NAND2_17991 ( P2_R1176_U424 , P2_R1176_U62 , P2_R1176_U24 );
nand NAND2_17992 ( P2_R1176_U425 , P2_R1176_U375 , P2_U3209 );
nand NAND2_17993 ( P2_R1176_U426 , P2_R1176_U62 , P2_R1176_U24 );
nand NAND2_17994 ( P2_R1176_U427 , P2_R1176_U426 , P2_R1176_U425 );
nand NAND2_17995 ( P2_R1176_U428 , P2_R1176_U150 , P2_R1176_U151 );
nand NAND2_17996 ( P2_R1176_U429 , P2_R1176_U216 , P2_R1176_U427 );
nand NAND2_17997 ( P2_R1176_U430 , P2_R1176_U384 , P2_U3210 );
nand NAND2_17998 ( P2_R1176_U431 , P2_R1176_U59 , P2_R1176_U21 );
nand NAND2_17999 ( P2_R1176_U432 , P2_R1176_U387 , P2_U3211 );
nand NAND2_18000 ( P2_R1176_U433 , P2_R1176_U58 , P2_R1176_U19 );
nand NAND2_18001 ( P2_R1176_U434 , P2_R1176_U433 , P2_R1176_U432 );
nand NAND2_18002 ( P2_R1176_U435 , P2_R1176_U347 , P2_R1176_U29 );
nand NAND2_18003 ( P2_R1176_U436 , P2_R1176_U434 , P2_R1176_U209 );
nand NAND2_18004 ( P2_R1176_U437 , P2_U3214 , P2_R1176_U152 );
nand NAND2_18005 ( P2_R1176_U438 , P2_U3969 , P2_R1176_U15 );
not NOT1_18006 ( P2_R1176_U439 , P2_R1176_U65 );
nand NAND2_18007 ( P2_R1176_U440 , P2_U3214 , P2_R1176_U153 );
nand NAND2_18008 ( P2_R1176_U441 , P2_U3480 , P2_R1176_U15 );
not NOT1_18009 ( P2_R1176_U442 , P2_R1176_U71 );
nand NAND2_18010 ( P2_R1176_U443 , P2_U3214 , P2_R1176_U154 );
nand NAND2_18011 ( P2_R1176_U444 , P2_U3489 , P2_R1176_U15 );
not NOT1_18012 ( P2_R1176_U445 , P2_R1176_U73 );
nand NAND2_18013 ( P2_R1176_U446 , P2_U3214 , P2_R1176_U155 );
nand NAND2_18014 ( P2_R1176_U447 , P2_U3486 , P2_R1176_U15 );
not NOT1_18015 ( P2_R1176_U448 , P2_R1176_U74 );
nand NAND2_18016 ( P2_R1176_U449 , P2_U3214 , P2_R1176_U156 );
nand NAND2_18017 ( P2_R1176_U450 , P2_U3483 , P2_R1176_U15 );
not NOT1_18018 ( P2_R1176_U451 , P2_R1176_U72 );
nand NAND2_18019 ( P2_R1176_U452 , P2_U3214 , P2_R1176_U157 );
nand NAND2_18020 ( P2_R1176_U453 , P2_U3492 , P2_R1176_U15 );
not NOT1_18021 ( P2_R1176_U454 , P2_R1176_U75 );
nand NAND2_18022 ( P2_R1176_U455 , P2_U3214 , P2_R1176_U158 );
nand NAND2_18023 ( P2_R1176_U456 , P2_U3495 , P2_R1176_U15 );
not NOT1_18024 ( P2_R1176_U457 , P2_R1176_U76 );
nand NAND2_18025 ( P2_R1176_U458 , P2_U3214 , P2_R1176_U159 );
nand NAND2_18026 ( P2_R1176_U459 , P2_U3501 , P2_R1176_U15 );
not NOT1_18027 ( P2_R1176_U460 , P2_R1176_U70 );
nand NAND2_18028 ( P2_R1176_U461 , P2_U3214 , P2_R1176_U160 );
nand NAND2_18029 ( P2_R1176_U462 , P2_U3498 , P2_R1176_U15 );
not NOT1_18030 ( P2_R1176_U463 , P2_R1176_U69 );
nand NAND2_18031 ( P2_R1176_U464 , P2_U3214 , P2_R1176_U161 );
nand NAND2_18032 ( P2_R1176_U465 , P2_U3504 , P2_R1176_U15 );
not NOT1_18033 ( P2_R1176_U466 , P2_R1176_U77 );
nand NAND2_18034 ( P2_R1176_U467 , P2_U3214 , P2_R1176_U162 );
nand NAND2_18035 ( P2_R1176_U468 , P2_U3975 , P2_R1176_U15 );
not NOT1_18036 ( P2_R1176_U469 , P2_R1176_U79 );
nand NAND2_18037 ( P2_R1176_U470 , P2_U3214 , P2_R1176_U163 );
nand NAND2_18038 ( P2_R1176_U471 , P2_U3976 , P2_R1176_U15 );
not NOT1_18039 ( P2_R1176_U472 , P2_R1176_U80 );
nand NAND2_18040 ( P2_R1176_U473 , P2_U3214 , P2_R1176_U164 );
nand NAND2_18041 ( P2_R1176_U474 , P2_U3506 , P2_R1176_U15 );
not NOT1_18042 ( P2_R1176_U475 , P2_R1176_U78 );
nand NAND2_18043 ( P2_R1176_U476 , P2_U3214 , P2_R1176_U165 );
nand NAND2_18044 ( P2_R1176_U477 , P2_U3974 , P2_R1176_U15 );
not NOT1_18045 ( P2_R1176_U478 , P2_R1176_U81 );
nand NAND2_18046 ( P2_R1176_U479 , P2_U3214 , P2_R1176_U166 );
nand NAND2_18047 ( P2_R1176_U480 , P2_U3973 , P2_R1176_U15 );
not NOT1_18048 ( P2_R1176_U481 , P2_R1176_U82 );
nand NAND2_18049 ( P2_R1176_U482 , P2_U3214 , P2_R1176_U167 );
nand NAND2_18050 ( P2_R1176_U483 , P2_U3971 , P2_R1176_U15 );
not NOT1_18051 ( P2_R1176_U484 , P2_R1176_U66 );
nand NAND2_18052 ( P2_R1176_U485 , P2_U3214 , P2_R1176_U168 );
nand NAND2_18053 ( P2_R1176_U486 , P2_U3970 , P2_R1176_U15 );
not NOT1_18054 ( P2_R1176_U487 , P2_R1176_U67 );
nand NAND2_18055 ( P2_R1176_U488 , P2_U3214 , P2_R1176_U169 );
nand NAND2_18056 ( P2_R1176_U489 , P2_U3972 , P2_R1176_U15 );
not NOT1_18057 ( P2_R1176_U490 , P2_R1176_U68 );
nand NAND2_18058 ( P2_R1176_U491 , P2_U3214 , P2_R1176_U170 );
nand NAND2_18059 ( P2_R1176_U492 , P2_U3185 , P2_R1176_U15 );
not NOT1_18060 ( P2_R1176_U493 , P2_R1176_U122 );
nand NAND2_18061 ( P2_R1176_U494 , P2_U3968 , P2_R1176_U493 );
nand NAND2_18062 ( P2_R1176_U495 , P2_R1176_U122 , P2_R1176_U171 );
not NOT1_18063 ( P2_R1176_U496 , P2_R1176_U83 );
nand NAND3_18064 ( P2_R1176_U497 , P2_R1176_U356 , P2_R1176_U309 , P2_R1176_U496 );
nand NAND4_18065 ( P2_R1176_U498 , P2_R1176_U363 , P2_R1176_U362 , P2_R1176_U121 , P2_R1176_U83 );
nand NAND2_18066 ( P2_R1176_U499 , P2_R1176_U439 , P2_U3186 );
nand NAND2_18067 ( P2_R1176_U500 , P2_R1176_U65 , P2_R1176_U30 );
nand NAND2_18068 ( P2_R1176_U501 , P2_R1176_U439 , P2_U3186 );
nand NAND2_18069 ( P2_R1176_U502 , P2_R1176_U65 , P2_R1176_U30 );
nand NAND2_18070 ( P2_R1176_U503 , P2_R1176_U502 , P2_R1176_U501 );
nand NAND2_18071 ( P2_R1176_U504 , P2_R1176_U172 , P2_R1176_U173 );
nand NAND2_18072 ( P2_R1176_U505 , P2_R1176_U308 , P2_R1176_U503 );
nand NAND2_18073 ( P2_R1176_U506 , P2_R1176_U487 , P2_U3187 );
nand NAND2_18074 ( P2_R1176_U507 , P2_R1176_U67 , P2_R1176_U31 );
nand NAND2_18075 ( P2_R1176_U508 , P2_R1176_U484 , P2_U3188 );
nand NAND2_18076 ( P2_R1176_U509 , P2_R1176_U66 , P2_R1176_U32 );
nand NAND2_18077 ( P2_R1176_U510 , P2_R1176_U509 , P2_R1176_U508 );
nand NAND2_18078 ( P2_R1176_U511 , P2_R1176_U348 , P2_R1176_U174 );
nand NAND2_18079 ( P2_R1176_U512 , P2_R1176_U313 , P2_R1176_U510 );
nand NAND2_18080 ( P2_R1176_U513 , P2_R1176_U490 , P2_U3189 );
nand NAND2_18081 ( P2_R1176_U514 , P2_R1176_U68 , P2_R1176_U33 );
nand NAND2_18082 ( P2_R1176_U515 , P2_R1176_U514 , P2_R1176_U513 );
nand NAND2_18083 ( P2_R1176_U516 , P2_R1176_U349 , P2_R1176_U175 );
nand NAND2_18084 ( P2_R1176_U517 , P2_R1176_U302 , P2_R1176_U515 );
nand NAND2_18085 ( P2_R1176_U518 , P2_R1176_U481 , P2_U3190 );
nand NAND2_18086 ( P2_R1176_U519 , P2_R1176_U82 , P2_R1176_U50 );
nand NAND2_18087 ( P2_R1176_U520 , P2_R1176_U481 , P2_U3190 );
nand NAND2_18088 ( P2_R1176_U521 , P2_R1176_U82 , P2_R1176_U50 );
nand NAND2_18089 ( P2_R1176_U522 , P2_R1176_U521 , P2_R1176_U520 );
nand NAND2_18090 ( P2_R1176_U523 , P2_R1176_U176 , P2_R1176_U177 );
nand NAND2_18091 ( P2_R1176_U524 , P2_R1176_U298 , P2_R1176_U522 );
nand NAND2_18092 ( P2_R1176_U525 , P2_R1176_U478 , P2_U3191 );
nand NAND2_18093 ( P2_R1176_U526 , P2_R1176_U81 , P2_R1176_U49 );
nand NAND2_18094 ( P2_R1176_U527 , P2_R1176_U478 , P2_U3191 );
nand NAND2_18095 ( P2_R1176_U528 , P2_R1176_U81 , P2_R1176_U49 );
nand NAND2_18096 ( P2_R1176_U529 , P2_R1176_U528 , P2_R1176_U527 );
nand NAND2_18097 ( P2_R1176_U530 , P2_R1176_U178 , P2_R1176_U179 );
nand NAND2_18098 ( P2_R1176_U531 , P2_R1176_U294 , P2_R1176_U529 );
nand NAND2_18099 ( P2_R1176_U532 , P2_R1176_U469 , P2_U3192 );
nand NAND2_18100 ( P2_R1176_U533 , P2_R1176_U79 , P2_R1176_U48 );
nand NAND2_18101 ( P2_R1176_U534 , P2_R1176_U472 , P2_U3193 );
nand NAND2_18102 ( P2_R1176_U535 , P2_R1176_U80 , P2_R1176_U45 );
nand NAND2_18103 ( P2_R1176_U536 , P2_R1176_U535 , P2_R1176_U534 );
nand NAND2_18104 ( P2_R1176_U537 , P2_R1176_U350 , P2_R1176_U52 );
nand NAND2_18105 ( P2_R1176_U538 , P2_R1176_U536 , P2_R1176_U322 );
nand NAND2_18106 ( P2_R1176_U539 , P2_R1176_U381 , P2_U3212 );
nand NAND2_18107 ( P2_R1176_U540 , P2_R1176_U61 , P2_R1176_U23 );
nand NAND2_18108 ( P2_R1176_U541 , P2_R1176_U381 , P2_U3212 );
nand NAND2_18109 ( P2_R1176_U542 , P2_R1176_U61 , P2_R1176_U23 );
nand NAND2_18110 ( P2_R1176_U543 , P2_R1176_U542 , P2_R1176_U541 );
nand NAND2_18111 ( P2_R1176_U544 , P2_R1176_U180 , P2_R1176_U181 );
nand NAND2_18112 ( P2_R1176_U545 , P2_R1176_U205 , P2_R1176_U543 );
nand NAND2_18113 ( P2_R1176_U546 , P2_R1176_U475 , P2_U3194 );
nand NAND2_18114 ( P2_R1176_U547 , P2_R1176_U78 , P2_R1176_U46 );
nand NAND2_18115 ( P2_R1176_U548 , P2_R1176_U547 , P2_R1176_U546 );
nand NAND2_18116 ( P2_R1176_U549 , P2_R1176_U351 , P2_R1176_U182 );
nand NAND2_18117 ( P2_R1176_U550 , P2_R1176_U284 , P2_R1176_U548 );
nand NAND2_18118 ( P2_R1176_U551 , P2_R1176_U466 , P2_U3195 );
nand NAND2_18119 ( P2_R1176_U552 , P2_R1176_U77 , P2_R1176_U44 );
nand NAND2_18120 ( P2_R1176_U553 , P2_R1176_U466 , P2_U3195 );
nand NAND2_18121 ( P2_R1176_U554 , P2_R1176_U77 , P2_R1176_U44 );
nand NAND2_18122 ( P2_R1176_U555 , P2_R1176_U554 , P2_R1176_U553 );
nand NAND2_18123 ( P2_R1176_U556 , P2_R1176_U183 , P2_R1176_U184 );
nand NAND2_18124 ( P2_R1176_U557 , P2_R1176_U280 , P2_R1176_U555 );
nand NAND2_18125 ( P2_R1176_U558 , P2_R1176_U460 , P2_U3196 );
nand NAND2_18126 ( P2_R1176_U559 , P2_R1176_U70 , P2_R1176_U36 );
nand NAND2_18127 ( P2_R1176_U560 , P2_R1176_U463 , P2_U3197 );
nand NAND2_18128 ( P2_R1176_U561 , P2_R1176_U69 , P2_R1176_U34 );
nand NAND2_18129 ( P2_R1176_U562 , P2_R1176_U561 , P2_R1176_U560 );
nand NAND2_18130 ( P2_R1176_U563 , P2_R1176_U352 , P2_R1176_U53 );
nand NAND2_18131 ( P2_R1176_U564 , P2_R1176_U562 , P2_R1176_U272 );
nand NAND2_18132 ( P2_R1176_U565 , P2_R1176_U457 , P2_U3198 );
nand NAND2_18133 ( P2_R1176_U566 , P2_R1176_U76 , P2_R1176_U43 );
nand NAND2_18134 ( P2_R1176_U567 , P2_R1176_U457 , P2_U3198 );
nand NAND2_18135 ( P2_R1176_U568 , P2_R1176_U76 , P2_R1176_U43 );
nand NAND2_18136 ( P2_R1176_U569 , P2_R1176_U568 , P2_R1176_U567 );
nand NAND2_18137 ( P2_R1176_U570 , P2_R1176_U185 , P2_R1176_U186 );
nand NAND2_18138 ( P2_R1176_U571 , P2_R1176_U268 , P2_R1176_U569 );
nand NAND2_18139 ( P2_R1176_U572 , P2_R1176_U454 , P2_U3199 );
nand NAND2_18140 ( P2_R1176_U573 , P2_R1176_U75 , P2_R1176_U42 );
nand NAND2_18141 ( P2_R1176_U574 , P2_R1176_U454 , P2_U3199 );
nand NAND2_18142 ( P2_R1176_U575 , P2_R1176_U75 , P2_R1176_U42 );
nand NAND2_18143 ( P2_R1176_U576 , P2_R1176_U575 , P2_R1176_U574 );
nand NAND2_18144 ( P2_R1176_U577 , P2_R1176_U187 , P2_R1176_U188 );
nand NAND2_18145 ( P2_R1176_U578 , P2_R1176_U264 , P2_R1176_U576 );
nand NAND2_18146 ( P2_R1176_U579 , P2_R1176_U445 , P2_U3200 );
nand NAND2_18147 ( P2_R1176_U580 , P2_R1176_U73 , P2_R1176_U41 );
nand NAND2_18148 ( P2_R1176_U581 , P2_R1176_U448 , P2_U3201 );
nand NAND2_18149 ( P2_R1176_U582 , P2_R1176_U74 , P2_R1176_U38 );
nand NAND2_18150 ( P2_R1176_U583 , P2_R1176_U582 , P2_R1176_U581 );
nand NAND2_18151 ( P2_R1176_U584 , P2_R1176_U353 , P2_R1176_U54 );
nand NAND2_18152 ( P2_R1176_U585 , P2_R1176_U583 , P2_R1176_U338 );
nand NAND2_18153 ( P2_R1176_U586 , P2_R1176_U451 , P2_U3202 );
nand NAND2_18154 ( P2_R1176_U587 , P2_R1176_U72 , P2_R1176_U39 );
nand NAND2_18155 ( P2_R1176_U588 , P2_R1176_U587 , P2_R1176_U586 );
nand NAND2_18156 ( P2_R1176_U589 , P2_R1176_U354 , P2_R1176_U189 );
nand NAND2_18157 ( P2_R1176_U590 , P2_R1176_U254 , P2_R1176_U588 );
nand NAND2_18158 ( P2_R1176_U591 , P2_R1176_U442 , P2_U3203 );
nand NAND2_18159 ( P2_R1176_U592 , P2_R1176_U71 , P2_R1176_U37 );
nand NAND2_18160 ( P2_R1176_U593 , P2_R1176_U442 , P2_U3203 );
nand NAND2_18161 ( P2_R1176_U594 , P2_R1176_U71 , P2_R1176_U37 );
nand NAND2_18162 ( P2_R1176_U595 , P2_R1176_U594 , P2_R1176_U593 );
nand NAND2_18163 ( P2_R1176_U596 , P2_R1176_U190 , P2_R1176_U191 );
nand NAND2_18164 ( P2_R1176_U597 , P2_R1176_U250 , P2_R1176_U595 );
nand NAND2_18165 ( P2_R1176_U598 , P2_U3213 , P2_R1176_U15 );
nand NAND2_18166 ( P2_R1176_U599 , P2_U3214 , P2_R1176_U22 );
not NOT1_18167 ( P2_R1176_U600 , P2_R1176_U133 );
nand NAND2_18168 ( P2_R1176_U601 , P2_R1176_U60 , P2_R1176_U600 );
nand NAND2_18169 ( P2_R1176_U602 , P2_R1176_U133 , P2_R1176_U378 );
and AND2_18170 ( P2_R1131_U4 , P2_R1131_U179 , P2_R1131_U178 );
and AND2_18171 ( P2_R1131_U5 , P2_R1131_U197 , P2_R1131_U196 );
and AND2_18172 ( P2_R1131_U6 , P2_R1131_U237 , P2_R1131_U236 );
and AND2_18173 ( P2_R1131_U7 , P2_R1131_U246 , P2_R1131_U245 );
and AND2_18174 ( P2_R1131_U8 , P2_R1131_U264 , P2_R1131_U263 );
and AND2_18175 ( P2_R1131_U9 , P2_R1131_U272 , P2_R1131_U271 );
and AND2_18176 ( P2_R1131_U10 , P2_R1131_U351 , P2_R1131_U348 );
and AND2_18177 ( P2_R1131_U11 , P2_R1131_U344 , P2_R1131_U341 );
and AND2_18178 ( P2_R1131_U12 , P2_R1131_U335 , P2_R1131_U332 );
and AND2_18179 ( P2_R1131_U13 , P2_R1131_U326 , P2_R1131_U323 );
and AND2_18180 ( P2_R1131_U14 , P2_R1131_U320 , P2_R1131_U318 );
and AND2_18181 ( P2_R1131_U15 , P2_R1131_U313 , P2_R1131_U310 );
and AND2_18182 ( P2_R1131_U16 , P2_R1131_U235 , P2_R1131_U232 );
and AND2_18183 ( P2_R1131_U17 , P2_R1131_U227 , P2_R1131_U224 );
and AND2_18184 ( P2_R1131_U18 , P2_R1131_U213 , P2_R1131_U210 );
not NOT1_18185 ( P2_R1131_U19 , P2_U3468 );
not NOT1_18186 ( P2_R1131_U20 , P2_U3071 );
not NOT1_18187 ( P2_R1131_U21 , P2_U3070 );
nand NAND2_18188 ( P2_R1131_U22 , P2_U3071 , P2_U3468 );
not NOT1_18189 ( P2_R1131_U23 , P2_U3471 );
not NOT1_18190 ( P2_R1131_U24 , P2_U3462 );
not NOT1_18191 ( P2_R1131_U25 , P2_U3060 );
not NOT1_18192 ( P2_R1131_U26 , P2_U3067 );
not NOT1_18193 ( P2_R1131_U27 , P2_U3456 );
not NOT1_18194 ( P2_R1131_U28 , P2_U3068 );
not NOT1_18195 ( P2_R1131_U29 , P2_U3448 );
not NOT1_18196 ( P2_R1131_U30 , P2_U3077 );
nand NAND2_18197 ( P2_R1131_U31 , P2_U3077 , P2_U3448 );
not NOT1_18198 ( P2_R1131_U32 , P2_U3459 );
not NOT1_18199 ( P2_R1131_U33 , P2_U3064 );
nand NAND2_18200 ( P2_R1131_U34 , P2_U3060 , P2_U3462 );
not NOT1_18201 ( P2_R1131_U35 , P2_U3465 );
not NOT1_18202 ( P2_R1131_U36 , P2_U3474 );
not NOT1_18203 ( P2_R1131_U37 , P2_U3084 );
not NOT1_18204 ( P2_R1131_U38 , P2_U3083 );
not NOT1_18205 ( P2_R1131_U39 , P2_U3477 );
nand NAND2_18206 ( P2_R1131_U40 , P2_R1131_U61 , P2_R1131_U205 );
nand NAND2_18207 ( P2_R1131_U41 , P2_R1131_U117 , P2_R1131_U193 );
nand NAND2_18208 ( P2_R1131_U42 , P2_R1131_U182 , P2_R1131_U183 );
nand NAND2_18209 ( P2_R1131_U43 , P2_U3453 , P2_U3078 );
nand NAND2_18210 ( P2_R1131_U44 , P2_R1131_U122 , P2_R1131_U219 );
nand NAND2_18211 ( P2_R1131_U45 , P2_R1131_U216 , P2_R1131_U215 );
not NOT1_18212 ( P2_R1131_U46 , P2_U3969 );
not NOT1_18213 ( P2_R1131_U47 , P2_U3053 );
not NOT1_18214 ( P2_R1131_U48 , P2_U3057 );
not NOT1_18215 ( P2_R1131_U49 , P2_U3970 );
not NOT1_18216 ( P2_R1131_U50 , P2_U3971 );
not NOT1_18217 ( P2_R1131_U51 , P2_U3058 );
not NOT1_18218 ( P2_R1131_U52 , P2_U3972 );
not NOT1_18219 ( P2_R1131_U53 , P2_U3065 );
not NOT1_18220 ( P2_R1131_U54 , P2_U3975 );
not NOT1_18221 ( P2_R1131_U55 , P2_U3075 );
not NOT1_18222 ( P2_R1131_U56 , P2_U3498 );
not NOT1_18223 ( P2_R1131_U57 , P2_U3073 );
not NOT1_18224 ( P2_R1131_U58 , P2_U3069 );
nand NAND2_18225 ( P2_R1131_U59 , P2_U3073 , P2_U3498 );
not NOT1_18226 ( P2_R1131_U60 , P2_U3501 );
nand NAND2_18227 ( P2_R1131_U61 , P2_U3084 , P2_U3474 );
not NOT1_18228 ( P2_R1131_U62 , P2_U3480 );
not NOT1_18229 ( P2_R1131_U63 , P2_U3062 );
not NOT1_18230 ( P2_R1131_U64 , P2_U3486 );
not NOT1_18231 ( P2_R1131_U65 , P2_U3072 );
not NOT1_18232 ( P2_R1131_U66 , P2_U3483 );
not NOT1_18233 ( P2_R1131_U67 , P2_U3063 );
nand NAND2_18234 ( P2_R1131_U68 , P2_U3063 , P2_U3483 );
not NOT1_18235 ( P2_R1131_U69 , P2_U3489 );
not NOT1_18236 ( P2_R1131_U70 , P2_U3080 );
not NOT1_18237 ( P2_R1131_U71 , P2_U3492 );
not NOT1_18238 ( P2_R1131_U72 , P2_U3079 );
not NOT1_18239 ( P2_R1131_U73 , P2_U3495 );
not NOT1_18240 ( P2_R1131_U74 , P2_U3074 );
not NOT1_18241 ( P2_R1131_U75 , P2_U3504 );
not NOT1_18242 ( P2_R1131_U76 , P2_U3082 );
nand NAND2_18243 ( P2_R1131_U77 , P2_U3082 , P2_U3504 );
not NOT1_18244 ( P2_R1131_U78 , P2_U3506 );
not NOT1_18245 ( P2_R1131_U79 , P2_U3081 );
nand NAND2_18246 ( P2_R1131_U80 , P2_U3081 , P2_U3506 );
not NOT1_18247 ( P2_R1131_U81 , P2_U3976 );
not NOT1_18248 ( P2_R1131_U82 , P2_U3974 );
not NOT1_18249 ( P2_R1131_U83 , P2_U3061 );
not NOT1_18250 ( P2_R1131_U84 , P2_U3973 );
not NOT1_18251 ( P2_R1131_U85 , P2_U3066 );
nand NAND2_18252 ( P2_R1131_U86 , P2_U3970 , P2_U3057 );
not NOT1_18253 ( P2_R1131_U87 , P2_U3054 );
not NOT1_18254 ( P2_R1131_U88 , P2_U3968 );
nand NAND2_18255 ( P2_R1131_U89 , P2_R1131_U306 , P2_R1131_U176 );
not NOT1_18256 ( P2_R1131_U90 , P2_U3076 );
nand NAND2_18257 ( P2_R1131_U91 , P2_R1131_U77 , P2_R1131_U315 );
nand NAND2_18258 ( P2_R1131_U92 , P2_R1131_U261 , P2_R1131_U260 );
nand NAND2_18259 ( P2_R1131_U93 , P2_R1131_U68 , P2_R1131_U337 );
nand NAND2_18260 ( P2_R1131_U94 , P2_R1131_U457 , P2_R1131_U456 );
nand NAND2_18261 ( P2_R1131_U95 , P2_R1131_U504 , P2_R1131_U503 );
nand NAND2_18262 ( P2_R1131_U96 , P2_R1131_U375 , P2_R1131_U374 );
nand NAND2_18263 ( P2_R1131_U97 , P2_R1131_U380 , P2_R1131_U379 );
nand NAND2_18264 ( P2_R1131_U98 , P2_R1131_U387 , P2_R1131_U386 );
nand NAND2_18265 ( P2_R1131_U99 , P2_R1131_U394 , P2_R1131_U393 );
nand NAND2_18266 ( P2_R1131_U100 , P2_R1131_U399 , P2_R1131_U398 );
nand NAND2_18267 ( P2_R1131_U101 , P2_R1131_U408 , P2_R1131_U407 );
nand NAND2_18268 ( P2_R1131_U102 , P2_R1131_U415 , P2_R1131_U414 );
nand NAND2_18269 ( P2_R1131_U103 , P2_R1131_U422 , P2_R1131_U421 );
nand NAND2_18270 ( P2_R1131_U104 , P2_R1131_U429 , P2_R1131_U428 );
nand NAND2_18271 ( P2_R1131_U105 , P2_R1131_U434 , P2_R1131_U433 );
nand NAND2_18272 ( P2_R1131_U106 , P2_R1131_U441 , P2_R1131_U440 );
nand NAND2_18273 ( P2_R1131_U107 , P2_R1131_U448 , P2_R1131_U447 );
nand NAND2_18274 ( P2_R1131_U108 , P2_R1131_U462 , P2_R1131_U461 );
nand NAND2_18275 ( P2_R1131_U109 , P2_R1131_U467 , P2_R1131_U466 );
nand NAND2_18276 ( P2_R1131_U110 , P2_R1131_U474 , P2_R1131_U473 );
nand NAND2_18277 ( P2_R1131_U111 , P2_R1131_U481 , P2_R1131_U480 );
nand NAND2_18278 ( P2_R1131_U112 , P2_R1131_U488 , P2_R1131_U487 );
nand NAND2_18279 ( P2_R1131_U113 , P2_R1131_U495 , P2_R1131_U494 );
nand NAND2_18280 ( P2_R1131_U114 , P2_R1131_U500 , P2_R1131_U499 );
and AND2_18281 ( P2_R1131_U115 , P2_R1131_U189 , P2_R1131_U187 );
and AND2_18282 ( P2_R1131_U116 , P2_R1131_U4 , P2_R1131_U180 );
and AND2_18283 ( P2_R1131_U117 , P2_R1131_U194 , P2_R1131_U192 );
and AND2_18284 ( P2_R1131_U118 , P2_R1131_U201 , P2_R1131_U200 );
and AND3_18285 ( P2_R1131_U119 , P2_R1131_U382 , P2_R1131_U381 , P2_R1131_U22 );
and AND2_18286 ( P2_R1131_U120 , P2_R1131_U212 , P2_R1131_U5 );
and AND2_18287 ( P2_R1131_U121 , P2_R1131_U181 , P2_R1131_U180 );
and AND2_18288 ( P2_R1131_U122 , P2_R1131_U220 , P2_R1131_U218 );
and AND3_18289 ( P2_R1131_U123 , P2_R1131_U389 , P2_R1131_U388 , P2_R1131_U34 );
and AND2_18290 ( P2_R1131_U124 , P2_R1131_U226 , P2_R1131_U4 );
and AND2_18291 ( P2_R1131_U125 , P2_R1131_U234 , P2_R1131_U181 );
and AND2_18292 ( P2_R1131_U126 , P2_R1131_U204 , P2_R1131_U6 );
and AND2_18293 ( P2_R1131_U127 , P2_R1131_U239 , P2_R1131_U171 );
and AND2_18294 ( P2_R1131_U128 , P2_R1131_U250 , P2_R1131_U7 );
and AND2_18295 ( P2_R1131_U129 , P2_R1131_U248 , P2_R1131_U172 );
and AND2_18296 ( P2_R1131_U130 , P2_R1131_U268 , P2_R1131_U267 );
and AND3_18297 ( P2_R1131_U131 , P2_R1131_U9 , P2_R1131_U282 , P2_R1131_U273 );
and AND2_18298 ( P2_R1131_U132 , P2_R1131_U285 , P2_R1131_U280 );
and AND2_18299 ( P2_R1131_U133 , P2_R1131_U301 , P2_R1131_U298 );
and AND2_18300 ( P2_R1131_U134 , P2_R1131_U368 , P2_R1131_U302 );
and AND3_18301 ( P2_R1131_U135 , P2_R1131_U424 , P2_R1131_U423 , P2_R1131_U173 );
and AND2_18302 ( P2_R1131_U136 , P2_R1131_U160 , P2_R1131_U278 );
and AND3_18303 ( P2_R1131_U137 , P2_R1131_U455 , P2_R1131_U454 , P2_R1131_U80 );
and AND2_18304 ( P2_R1131_U138 , P2_R1131_U325 , P2_R1131_U9 );
and AND3_18305 ( P2_R1131_U139 , P2_R1131_U469 , P2_R1131_U468 , P2_R1131_U59 );
and AND2_18306 ( P2_R1131_U140 , P2_R1131_U334 , P2_R1131_U8 );
and AND3_18307 ( P2_R1131_U141 , P2_R1131_U490 , P2_R1131_U489 , P2_R1131_U172 );
and AND2_18308 ( P2_R1131_U142 , P2_R1131_U343 , P2_R1131_U7 );
and AND3_18309 ( P2_R1131_U143 , P2_R1131_U502 , P2_R1131_U501 , P2_R1131_U171 );
and AND2_18310 ( P2_R1131_U144 , P2_R1131_U350 , P2_R1131_U6 );
nand NAND2_18311 ( P2_R1131_U145 , P2_R1131_U118 , P2_R1131_U202 );
nand NAND2_18312 ( P2_R1131_U146 , P2_R1131_U217 , P2_R1131_U229 );
not NOT1_18313 ( P2_R1131_U147 , P2_U3055 );
not NOT1_18314 ( P2_R1131_U148 , P2_U3979 );
and AND2_18315 ( P2_R1131_U149 , P2_R1131_U403 , P2_R1131_U402 );
nand NAND3_18316 ( P2_R1131_U150 , P2_R1131_U304 , P2_R1131_U169 , P2_R1131_U364 );
and AND2_18317 ( P2_R1131_U151 , P2_R1131_U410 , P2_R1131_U409 );
nand NAND3_18318 ( P2_R1131_U152 , P2_R1131_U370 , P2_R1131_U369 , P2_R1131_U134 );
and AND2_18319 ( P2_R1131_U153 , P2_R1131_U417 , P2_R1131_U416 );
nand NAND3_18320 ( P2_R1131_U154 , P2_R1131_U365 , P2_R1131_U299 , P2_R1131_U86 );
nand NAND2_18321 ( P2_R1131_U155 , P2_R1131_U293 , P2_R1131_U292 );
and AND2_18322 ( P2_R1131_U156 , P2_R1131_U436 , P2_R1131_U435 );
nand NAND2_18323 ( P2_R1131_U157 , P2_R1131_U289 , P2_R1131_U288 );
and AND2_18324 ( P2_R1131_U158 , P2_R1131_U443 , P2_R1131_U442 );
nand NAND2_18325 ( P2_R1131_U159 , P2_R1131_U132 , P2_R1131_U284 );
and AND2_18326 ( P2_R1131_U160 , P2_R1131_U450 , P2_R1131_U449 );
nand NAND2_18327 ( P2_R1131_U161 , P2_R1131_U43 , P2_R1131_U327 );
nand NAND2_18328 ( P2_R1131_U162 , P2_R1131_U130 , P2_R1131_U269 );
and AND2_18329 ( P2_R1131_U163 , P2_R1131_U476 , P2_R1131_U475 );
nand NAND2_18330 ( P2_R1131_U164 , P2_R1131_U257 , P2_R1131_U256 );
and AND2_18331 ( P2_R1131_U165 , P2_R1131_U483 , P2_R1131_U482 );
nand NAND2_18332 ( P2_R1131_U166 , P2_R1131_U253 , P2_R1131_U252 );
nand NAND2_18333 ( P2_R1131_U167 , P2_R1131_U243 , P2_R1131_U242 );
nand NAND2_18334 ( P2_R1131_U168 , P2_R1131_U367 , P2_R1131_U366 );
nand NAND2_18335 ( P2_R1131_U169 , P2_U3054 , P2_R1131_U152 );
not NOT1_18336 ( P2_R1131_U170 , P2_R1131_U34 );
nand NAND2_18337 ( P2_R1131_U171 , P2_U3477 , P2_U3083 );
nand NAND2_18338 ( P2_R1131_U172 , P2_U3072 , P2_U3486 );
nand NAND2_18339 ( P2_R1131_U173 , P2_U3058 , P2_U3971 );
not NOT1_18340 ( P2_R1131_U174 , P2_R1131_U68 );
not NOT1_18341 ( P2_R1131_U175 , P2_R1131_U77 );
nand NAND2_18342 ( P2_R1131_U176 , P2_U3065 , P2_U3972 );
not NOT1_18343 ( P2_R1131_U177 , P2_R1131_U61 );
or OR2_18344 ( P2_R1131_U178 , P2_U3067 , P2_U3465 );
or OR2_18345 ( P2_R1131_U179 , P2_U3060 , P2_U3462 );
or OR2_18346 ( P2_R1131_U180 , P2_U3459 , P2_U3064 );
or OR2_18347 ( P2_R1131_U181 , P2_U3456 , P2_U3068 );
not NOT1_18348 ( P2_R1131_U182 , P2_R1131_U31 );
or OR2_18349 ( P2_R1131_U183 , P2_U3453 , P2_U3078 );
not NOT1_18350 ( P2_R1131_U184 , P2_R1131_U42 );
not NOT1_18351 ( P2_R1131_U185 , P2_R1131_U43 );
nand NAND2_18352 ( P2_R1131_U186 , P2_R1131_U42 , P2_R1131_U43 );
nand NAND2_18353 ( P2_R1131_U187 , P2_U3068 , P2_U3456 );
nand NAND2_18354 ( P2_R1131_U188 , P2_R1131_U186 , P2_R1131_U181 );
nand NAND2_18355 ( P2_R1131_U189 , P2_U3064 , P2_U3459 );
nand NAND2_18356 ( P2_R1131_U190 , P2_R1131_U115 , P2_R1131_U188 );
nand NAND2_18357 ( P2_R1131_U191 , P2_R1131_U35 , P2_R1131_U34 );
nand NAND2_18358 ( P2_R1131_U192 , P2_U3067 , P2_R1131_U191 );
nand NAND2_18359 ( P2_R1131_U193 , P2_R1131_U116 , P2_R1131_U190 );
nand NAND2_18360 ( P2_R1131_U194 , P2_U3465 , P2_R1131_U170 );
not NOT1_18361 ( P2_R1131_U195 , P2_R1131_U41 );
or OR2_18362 ( P2_R1131_U196 , P2_U3070 , P2_U3471 );
or OR2_18363 ( P2_R1131_U197 , P2_U3071 , P2_U3468 );
not NOT1_18364 ( P2_R1131_U198 , P2_R1131_U22 );
nand NAND2_18365 ( P2_R1131_U199 , P2_R1131_U23 , P2_R1131_U22 );
nand NAND2_18366 ( P2_R1131_U200 , P2_U3070 , P2_R1131_U199 );
nand NAND2_18367 ( P2_R1131_U201 , P2_U3471 , P2_R1131_U198 );
nand NAND2_18368 ( P2_R1131_U202 , P2_R1131_U5 , P2_R1131_U41 );
not NOT1_18369 ( P2_R1131_U203 , P2_R1131_U145 );
or OR2_18370 ( P2_R1131_U204 , P2_U3474 , P2_U3084 );
nand NAND2_18371 ( P2_R1131_U205 , P2_R1131_U204 , P2_R1131_U145 );
not NOT1_18372 ( P2_R1131_U206 , P2_R1131_U40 );
or OR2_18373 ( P2_R1131_U207 , P2_U3083 , P2_U3477 );
or OR2_18374 ( P2_R1131_U208 , P2_U3468 , P2_U3071 );
nand NAND2_18375 ( P2_R1131_U209 , P2_R1131_U208 , P2_R1131_U41 );
nand NAND2_18376 ( P2_R1131_U210 , P2_R1131_U119 , P2_R1131_U209 );
nand NAND2_18377 ( P2_R1131_U211 , P2_R1131_U195 , P2_R1131_U22 );
nand NAND2_18378 ( P2_R1131_U212 , P2_U3471 , P2_U3070 );
nand NAND2_18379 ( P2_R1131_U213 , P2_R1131_U120 , P2_R1131_U211 );
or OR2_18380 ( P2_R1131_U214 , P2_U3071 , P2_U3468 );
nand NAND2_18381 ( P2_R1131_U215 , P2_R1131_U185 , P2_R1131_U181 );
nand NAND2_18382 ( P2_R1131_U216 , P2_U3068 , P2_U3456 );
not NOT1_18383 ( P2_R1131_U217 , P2_R1131_U45 );
nand NAND2_18384 ( P2_R1131_U218 , P2_R1131_U121 , P2_R1131_U184 );
nand NAND2_18385 ( P2_R1131_U219 , P2_R1131_U45 , P2_R1131_U180 );
nand NAND2_18386 ( P2_R1131_U220 , P2_U3064 , P2_U3459 );
not NOT1_18387 ( P2_R1131_U221 , P2_R1131_U44 );
or OR2_18388 ( P2_R1131_U222 , P2_U3462 , P2_U3060 );
nand NAND2_18389 ( P2_R1131_U223 , P2_R1131_U222 , P2_R1131_U44 );
nand NAND2_18390 ( P2_R1131_U224 , P2_R1131_U123 , P2_R1131_U223 );
nand NAND2_18391 ( P2_R1131_U225 , P2_R1131_U221 , P2_R1131_U34 );
nand NAND2_18392 ( P2_R1131_U226 , P2_U3465 , P2_U3067 );
nand NAND2_18393 ( P2_R1131_U227 , P2_R1131_U124 , P2_R1131_U225 );
or OR2_18394 ( P2_R1131_U228 , P2_U3060 , P2_U3462 );
nand NAND2_18395 ( P2_R1131_U229 , P2_R1131_U184 , P2_R1131_U181 );
not NOT1_18396 ( P2_R1131_U230 , P2_R1131_U146 );
nand NAND2_18397 ( P2_R1131_U231 , P2_U3064 , P2_U3459 );
nand NAND4_18398 ( P2_R1131_U232 , P2_R1131_U401 , P2_R1131_U400 , P2_R1131_U43 , P2_R1131_U42 );
nand NAND2_18399 ( P2_R1131_U233 , P2_R1131_U43 , P2_R1131_U42 );
nand NAND2_18400 ( P2_R1131_U234 , P2_U3068 , P2_U3456 );
nand NAND2_18401 ( P2_R1131_U235 , P2_R1131_U125 , P2_R1131_U233 );
or OR2_18402 ( P2_R1131_U236 , P2_U3083 , P2_U3477 );
or OR2_18403 ( P2_R1131_U237 , P2_U3062 , P2_U3480 );
nand NAND2_18404 ( P2_R1131_U238 , P2_R1131_U177 , P2_R1131_U6 );
nand NAND2_18405 ( P2_R1131_U239 , P2_U3062 , P2_U3480 );
nand NAND2_18406 ( P2_R1131_U240 , P2_R1131_U127 , P2_R1131_U238 );
or OR2_18407 ( P2_R1131_U241 , P2_U3480 , P2_U3062 );
nand NAND2_18408 ( P2_R1131_U242 , P2_R1131_U126 , P2_R1131_U145 );
nand NAND2_18409 ( P2_R1131_U243 , P2_R1131_U241 , P2_R1131_U240 );
not NOT1_18410 ( P2_R1131_U244 , P2_R1131_U167 );
or OR2_18411 ( P2_R1131_U245 , P2_U3080 , P2_U3489 );
or OR2_18412 ( P2_R1131_U246 , P2_U3072 , P2_U3486 );
nand NAND2_18413 ( P2_R1131_U247 , P2_R1131_U174 , P2_R1131_U7 );
nand NAND2_18414 ( P2_R1131_U248 , P2_U3080 , P2_U3489 );
nand NAND2_18415 ( P2_R1131_U249 , P2_R1131_U129 , P2_R1131_U247 );
or OR2_18416 ( P2_R1131_U250 , P2_U3483 , P2_U3063 );
or OR2_18417 ( P2_R1131_U251 , P2_U3489 , P2_U3080 );
nand NAND2_18418 ( P2_R1131_U252 , P2_R1131_U128 , P2_R1131_U167 );
nand NAND2_18419 ( P2_R1131_U253 , P2_R1131_U251 , P2_R1131_U249 );
not NOT1_18420 ( P2_R1131_U254 , P2_R1131_U166 );
or OR2_18421 ( P2_R1131_U255 , P2_U3492 , P2_U3079 );
nand NAND2_18422 ( P2_R1131_U256 , P2_R1131_U255 , P2_R1131_U166 );
nand NAND2_18423 ( P2_R1131_U257 , P2_U3079 , P2_U3492 );
not NOT1_18424 ( P2_R1131_U258 , P2_R1131_U164 );
or OR2_18425 ( P2_R1131_U259 , P2_U3495 , P2_U3074 );
nand NAND2_18426 ( P2_R1131_U260 , P2_R1131_U259 , P2_R1131_U164 );
nand NAND2_18427 ( P2_R1131_U261 , P2_U3074 , P2_U3495 );
not NOT1_18428 ( P2_R1131_U262 , P2_R1131_U92 );
or OR2_18429 ( P2_R1131_U263 , P2_U3069 , P2_U3501 );
or OR2_18430 ( P2_R1131_U264 , P2_U3073 , P2_U3498 );
not NOT1_18431 ( P2_R1131_U265 , P2_R1131_U59 );
nand NAND2_18432 ( P2_R1131_U266 , P2_R1131_U60 , P2_R1131_U59 );
nand NAND2_18433 ( P2_R1131_U267 , P2_U3069 , P2_R1131_U266 );
nand NAND2_18434 ( P2_R1131_U268 , P2_U3501 , P2_R1131_U265 );
nand NAND2_18435 ( P2_R1131_U269 , P2_R1131_U8 , P2_R1131_U92 );
not NOT1_18436 ( P2_R1131_U270 , P2_R1131_U162 );
or OR2_18437 ( P2_R1131_U271 , P2_U3076 , P2_U3976 );
or OR2_18438 ( P2_R1131_U272 , P2_U3081 , P2_U3506 );
or OR2_18439 ( P2_R1131_U273 , P2_U3075 , P2_U3975 );
not NOT1_18440 ( P2_R1131_U274 , P2_R1131_U80 );
nand NAND2_18441 ( P2_R1131_U275 , P2_U3976 , P2_R1131_U274 );
nand NAND2_18442 ( P2_R1131_U276 , P2_R1131_U275 , P2_R1131_U90 );
nand NAND2_18443 ( P2_R1131_U277 , P2_R1131_U80 , P2_R1131_U81 );
nand NAND2_18444 ( P2_R1131_U278 , P2_R1131_U277 , P2_R1131_U276 );
nand NAND2_18445 ( P2_R1131_U279 , P2_R1131_U175 , P2_R1131_U9 );
nand NAND2_18446 ( P2_R1131_U280 , P2_U3075 , P2_U3975 );
nand NAND2_18447 ( P2_R1131_U281 , P2_R1131_U278 , P2_R1131_U279 );
or OR2_18448 ( P2_R1131_U282 , P2_U3504 , P2_U3082 );
or OR2_18449 ( P2_R1131_U283 , P2_U3975 , P2_U3075 );
nand NAND2_18450 ( P2_R1131_U284 , P2_R1131_U162 , P2_R1131_U131 );
nand NAND2_18451 ( P2_R1131_U285 , P2_R1131_U283 , P2_R1131_U281 );
not NOT1_18452 ( P2_R1131_U286 , P2_R1131_U159 );
or OR2_18453 ( P2_R1131_U287 , P2_U3974 , P2_U3061 );
nand NAND2_18454 ( P2_R1131_U288 , P2_R1131_U287 , P2_R1131_U159 );
nand NAND2_18455 ( P2_R1131_U289 , P2_U3061 , P2_U3974 );
not NOT1_18456 ( P2_R1131_U290 , P2_R1131_U157 );
or OR2_18457 ( P2_R1131_U291 , P2_U3973 , P2_U3066 );
nand NAND2_18458 ( P2_R1131_U292 , P2_R1131_U291 , P2_R1131_U157 );
nand NAND2_18459 ( P2_R1131_U293 , P2_U3066 , P2_U3973 );
not NOT1_18460 ( P2_R1131_U294 , P2_R1131_U155 );
or OR2_18461 ( P2_R1131_U295 , P2_U3058 , P2_U3971 );
nand NAND2_18462 ( P2_R1131_U296 , P2_R1131_U176 , P2_R1131_U173 );
not NOT1_18463 ( P2_R1131_U297 , P2_R1131_U86 );
or OR2_18464 ( P2_R1131_U298 , P2_U3972 , P2_U3065 );
nand NAND3_18465 ( P2_R1131_U299 , P2_R1131_U155 , P2_R1131_U298 , P2_R1131_U168 );
not NOT1_18466 ( P2_R1131_U300 , P2_R1131_U154 );
or OR2_18467 ( P2_R1131_U301 , P2_U3969 , P2_U3053 );
nand NAND2_18468 ( P2_R1131_U302 , P2_U3053 , P2_U3969 );
not NOT1_18469 ( P2_R1131_U303 , P2_R1131_U152 );
nand NAND2_18470 ( P2_R1131_U304 , P2_U3968 , P2_R1131_U152 );
not NOT1_18471 ( P2_R1131_U305 , P2_R1131_U150 );
nand NAND2_18472 ( P2_R1131_U306 , P2_R1131_U298 , P2_R1131_U155 );
not NOT1_18473 ( P2_R1131_U307 , P2_R1131_U89 );
or OR2_18474 ( P2_R1131_U308 , P2_U3971 , P2_U3058 );
nand NAND2_18475 ( P2_R1131_U309 , P2_R1131_U308 , P2_R1131_U89 );
nand NAND2_18476 ( P2_R1131_U310 , P2_R1131_U135 , P2_R1131_U309 );
nand NAND2_18477 ( P2_R1131_U311 , P2_R1131_U307 , P2_R1131_U173 );
nand NAND2_18478 ( P2_R1131_U312 , P2_U3970 , P2_U3057 );
nand NAND3_18479 ( P2_R1131_U313 , P2_R1131_U311 , P2_R1131_U312 , P2_R1131_U168 );
or OR2_18480 ( P2_R1131_U314 , P2_U3058 , P2_U3971 );
nand NAND2_18481 ( P2_R1131_U315 , P2_R1131_U282 , P2_R1131_U162 );
not NOT1_18482 ( P2_R1131_U316 , P2_R1131_U91 );
nand NAND2_18483 ( P2_R1131_U317 , P2_R1131_U9 , P2_R1131_U91 );
nand NAND2_18484 ( P2_R1131_U318 , P2_R1131_U136 , P2_R1131_U317 );
nand NAND2_18485 ( P2_R1131_U319 , P2_R1131_U317 , P2_R1131_U278 );
nand NAND2_18486 ( P2_R1131_U320 , P2_R1131_U453 , P2_R1131_U319 );
or OR2_18487 ( P2_R1131_U321 , P2_U3506 , P2_U3081 );
nand NAND2_18488 ( P2_R1131_U322 , P2_R1131_U321 , P2_R1131_U91 );
nand NAND2_18489 ( P2_R1131_U323 , P2_R1131_U137 , P2_R1131_U322 );
nand NAND2_18490 ( P2_R1131_U324 , P2_R1131_U316 , P2_R1131_U80 );
nand NAND2_18491 ( P2_R1131_U325 , P2_U3076 , P2_U3976 );
nand NAND2_18492 ( P2_R1131_U326 , P2_R1131_U138 , P2_R1131_U324 );
or OR2_18493 ( P2_R1131_U327 , P2_U3453 , P2_U3078 );
not NOT1_18494 ( P2_R1131_U328 , P2_R1131_U161 );
or OR2_18495 ( P2_R1131_U329 , P2_U3081 , P2_U3506 );
or OR2_18496 ( P2_R1131_U330 , P2_U3498 , P2_U3073 );
nand NAND2_18497 ( P2_R1131_U331 , P2_R1131_U330 , P2_R1131_U92 );
nand NAND2_18498 ( P2_R1131_U332 , P2_R1131_U139 , P2_R1131_U331 );
nand NAND2_18499 ( P2_R1131_U333 , P2_R1131_U262 , P2_R1131_U59 );
nand NAND2_18500 ( P2_R1131_U334 , P2_U3501 , P2_U3069 );
nand NAND2_18501 ( P2_R1131_U335 , P2_R1131_U140 , P2_R1131_U333 );
or OR2_18502 ( P2_R1131_U336 , P2_U3073 , P2_U3498 );
nand NAND2_18503 ( P2_R1131_U337 , P2_R1131_U250 , P2_R1131_U167 );
not NOT1_18504 ( P2_R1131_U338 , P2_R1131_U93 );
or OR2_18505 ( P2_R1131_U339 , P2_U3486 , P2_U3072 );
nand NAND2_18506 ( P2_R1131_U340 , P2_R1131_U339 , P2_R1131_U93 );
nand NAND2_18507 ( P2_R1131_U341 , P2_R1131_U141 , P2_R1131_U340 );
nand NAND2_18508 ( P2_R1131_U342 , P2_R1131_U338 , P2_R1131_U172 );
nand NAND2_18509 ( P2_R1131_U343 , P2_U3080 , P2_U3489 );
nand NAND2_18510 ( P2_R1131_U344 , P2_R1131_U142 , P2_R1131_U342 );
or OR2_18511 ( P2_R1131_U345 , P2_U3072 , P2_U3486 );
or OR2_18512 ( P2_R1131_U346 , P2_U3477 , P2_U3083 );
nand NAND2_18513 ( P2_R1131_U347 , P2_R1131_U346 , P2_R1131_U40 );
nand NAND2_18514 ( P2_R1131_U348 , P2_R1131_U143 , P2_R1131_U347 );
nand NAND2_18515 ( P2_R1131_U349 , P2_R1131_U206 , P2_R1131_U171 );
nand NAND2_18516 ( P2_R1131_U350 , P2_U3062 , P2_U3480 );
nand NAND2_18517 ( P2_R1131_U351 , P2_R1131_U144 , P2_R1131_U349 );
nand NAND2_18518 ( P2_R1131_U352 , P2_R1131_U207 , P2_R1131_U171 );
nand NAND2_18519 ( P2_R1131_U353 , P2_R1131_U204 , P2_R1131_U61 );
nand NAND2_18520 ( P2_R1131_U354 , P2_R1131_U214 , P2_R1131_U22 );
nand NAND2_18521 ( P2_R1131_U355 , P2_R1131_U228 , P2_R1131_U34 );
nand NAND2_18522 ( P2_R1131_U356 , P2_R1131_U231 , P2_R1131_U180 );
nand NAND2_18523 ( P2_R1131_U357 , P2_R1131_U314 , P2_R1131_U173 );
nand NAND2_18524 ( P2_R1131_U358 , P2_R1131_U298 , P2_R1131_U176 );
nand NAND2_18525 ( P2_R1131_U359 , P2_R1131_U329 , P2_R1131_U80 );
nand NAND2_18526 ( P2_R1131_U360 , P2_R1131_U282 , P2_R1131_U77 );
nand NAND2_18527 ( P2_R1131_U361 , P2_R1131_U336 , P2_R1131_U59 );
nand NAND2_18528 ( P2_R1131_U362 , P2_R1131_U345 , P2_R1131_U172 );
nand NAND2_18529 ( P2_R1131_U363 , P2_R1131_U250 , P2_R1131_U68 );
nand NAND2_18530 ( P2_R1131_U364 , P2_U3968 , P2_U3054 );
nand NAND2_18531 ( P2_R1131_U365 , P2_R1131_U296 , P2_R1131_U168 );
nand NAND2_18532 ( P2_R1131_U366 , P2_U3057 , P2_R1131_U295 );
nand NAND2_18533 ( P2_R1131_U367 , P2_U3970 , P2_R1131_U295 );
nand NAND3_18534 ( P2_R1131_U368 , P2_R1131_U296 , P2_R1131_U168 , P2_R1131_U301 );
nand NAND3_18535 ( P2_R1131_U369 , P2_R1131_U155 , P2_R1131_U168 , P2_R1131_U133 );
nand NAND2_18536 ( P2_R1131_U370 , P2_R1131_U297 , P2_R1131_U301 );
nand NAND2_18537 ( P2_R1131_U371 , P2_U3083 , P2_R1131_U39 );
nand NAND2_18538 ( P2_R1131_U372 , P2_U3477 , P2_R1131_U38 );
nand NAND2_18539 ( P2_R1131_U373 , P2_R1131_U372 , P2_R1131_U371 );
nand NAND2_18540 ( P2_R1131_U374 , P2_R1131_U352 , P2_R1131_U40 );
nand NAND2_18541 ( P2_R1131_U375 , P2_R1131_U373 , P2_R1131_U206 );
nand NAND2_18542 ( P2_R1131_U376 , P2_U3084 , P2_R1131_U36 );
nand NAND2_18543 ( P2_R1131_U377 , P2_U3474 , P2_R1131_U37 );
nand NAND2_18544 ( P2_R1131_U378 , P2_R1131_U377 , P2_R1131_U376 );
nand NAND2_18545 ( P2_R1131_U379 , P2_R1131_U353 , P2_R1131_U145 );
nand NAND2_18546 ( P2_R1131_U380 , P2_R1131_U203 , P2_R1131_U378 );
nand NAND2_18547 ( P2_R1131_U381 , P2_U3070 , P2_R1131_U23 );
nand NAND2_18548 ( P2_R1131_U382 , P2_U3471 , P2_R1131_U21 );
nand NAND2_18549 ( P2_R1131_U383 , P2_U3071 , P2_R1131_U19 );
nand NAND2_18550 ( P2_R1131_U384 , P2_U3468 , P2_R1131_U20 );
nand NAND2_18551 ( P2_R1131_U385 , P2_R1131_U384 , P2_R1131_U383 );
nand NAND2_18552 ( P2_R1131_U386 , P2_R1131_U354 , P2_R1131_U41 );
nand NAND2_18553 ( P2_R1131_U387 , P2_R1131_U385 , P2_R1131_U195 );
nand NAND2_18554 ( P2_R1131_U388 , P2_U3067 , P2_R1131_U35 );
nand NAND2_18555 ( P2_R1131_U389 , P2_U3465 , P2_R1131_U26 );
nand NAND2_18556 ( P2_R1131_U390 , P2_U3060 , P2_R1131_U24 );
nand NAND2_18557 ( P2_R1131_U391 , P2_U3462 , P2_R1131_U25 );
nand NAND2_18558 ( P2_R1131_U392 , P2_R1131_U391 , P2_R1131_U390 );
nand NAND2_18559 ( P2_R1131_U393 , P2_R1131_U355 , P2_R1131_U44 );
nand NAND2_18560 ( P2_R1131_U394 , P2_R1131_U392 , P2_R1131_U221 );
nand NAND2_18561 ( P2_R1131_U395 , P2_U3064 , P2_R1131_U32 );
nand NAND2_18562 ( P2_R1131_U396 , P2_U3459 , P2_R1131_U33 );
nand NAND2_18563 ( P2_R1131_U397 , P2_R1131_U396 , P2_R1131_U395 );
nand NAND2_18564 ( P2_R1131_U398 , P2_R1131_U356 , P2_R1131_U146 );
nand NAND2_18565 ( P2_R1131_U399 , P2_R1131_U230 , P2_R1131_U397 );
nand NAND2_18566 ( P2_R1131_U400 , P2_U3068 , P2_R1131_U27 );
nand NAND2_18567 ( P2_R1131_U401 , P2_U3456 , P2_R1131_U28 );
nand NAND2_18568 ( P2_R1131_U402 , P2_U3055 , P2_R1131_U148 );
nand NAND2_18569 ( P2_R1131_U403 , P2_U3979 , P2_R1131_U147 );
nand NAND2_18570 ( P2_R1131_U404 , P2_U3055 , P2_R1131_U148 );
nand NAND2_18571 ( P2_R1131_U405 , P2_U3979 , P2_R1131_U147 );
nand NAND2_18572 ( P2_R1131_U406 , P2_R1131_U405 , P2_R1131_U404 );
nand NAND2_18573 ( P2_R1131_U407 , P2_R1131_U149 , P2_R1131_U150 );
nand NAND2_18574 ( P2_R1131_U408 , P2_R1131_U305 , P2_R1131_U406 );
nand NAND2_18575 ( P2_R1131_U409 , P2_U3054 , P2_R1131_U88 );
nand NAND2_18576 ( P2_R1131_U410 , P2_U3968 , P2_R1131_U87 );
nand NAND2_18577 ( P2_R1131_U411 , P2_U3054 , P2_R1131_U88 );
nand NAND2_18578 ( P2_R1131_U412 , P2_U3968 , P2_R1131_U87 );
nand NAND2_18579 ( P2_R1131_U413 , P2_R1131_U412 , P2_R1131_U411 );
nand NAND2_18580 ( P2_R1131_U414 , P2_R1131_U151 , P2_R1131_U152 );
nand NAND2_18581 ( P2_R1131_U415 , P2_R1131_U303 , P2_R1131_U413 );
nand NAND2_18582 ( P2_R1131_U416 , P2_U3053 , P2_R1131_U46 );
nand NAND2_18583 ( P2_R1131_U417 , P2_U3969 , P2_R1131_U47 );
nand NAND2_18584 ( P2_R1131_U418 , P2_U3053 , P2_R1131_U46 );
nand NAND2_18585 ( P2_R1131_U419 , P2_U3969 , P2_R1131_U47 );
nand NAND2_18586 ( P2_R1131_U420 , P2_R1131_U419 , P2_R1131_U418 );
nand NAND2_18587 ( P2_R1131_U421 , P2_R1131_U153 , P2_R1131_U154 );
nand NAND2_18588 ( P2_R1131_U422 , P2_R1131_U300 , P2_R1131_U420 );
nand NAND2_18589 ( P2_R1131_U423 , P2_U3057 , P2_R1131_U49 );
nand NAND2_18590 ( P2_R1131_U424 , P2_U3970 , P2_R1131_U48 );
nand NAND2_18591 ( P2_R1131_U425 , P2_U3058 , P2_R1131_U50 );
nand NAND2_18592 ( P2_R1131_U426 , P2_U3971 , P2_R1131_U51 );
nand NAND2_18593 ( P2_R1131_U427 , P2_R1131_U426 , P2_R1131_U425 );
nand NAND2_18594 ( P2_R1131_U428 , P2_R1131_U357 , P2_R1131_U89 );
nand NAND2_18595 ( P2_R1131_U429 , P2_R1131_U427 , P2_R1131_U307 );
nand NAND2_18596 ( P2_R1131_U430 , P2_U3065 , P2_R1131_U52 );
nand NAND2_18597 ( P2_R1131_U431 , P2_U3972 , P2_R1131_U53 );
nand NAND2_18598 ( P2_R1131_U432 , P2_R1131_U431 , P2_R1131_U430 );
nand NAND2_18599 ( P2_R1131_U433 , P2_R1131_U358 , P2_R1131_U155 );
nand NAND2_18600 ( P2_R1131_U434 , P2_R1131_U294 , P2_R1131_U432 );
nand NAND2_18601 ( P2_R1131_U435 , P2_U3066 , P2_R1131_U84 );
nand NAND2_18602 ( P2_R1131_U436 , P2_U3973 , P2_R1131_U85 );
nand NAND2_18603 ( P2_R1131_U437 , P2_U3066 , P2_R1131_U84 );
nand NAND2_18604 ( P2_R1131_U438 , P2_U3973 , P2_R1131_U85 );
nand NAND2_18605 ( P2_R1131_U439 , P2_R1131_U438 , P2_R1131_U437 );
nand NAND2_18606 ( P2_R1131_U440 , P2_R1131_U156 , P2_R1131_U157 );
nand NAND2_18607 ( P2_R1131_U441 , P2_R1131_U290 , P2_R1131_U439 );
nand NAND2_18608 ( P2_R1131_U442 , P2_U3061 , P2_R1131_U82 );
nand NAND2_18609 ( P2_R1131_U443 , P2_U3974 , P2_R1131_U83 );
nand NAND2_18610 ( P2_R1131_U444 , P2_U3061 , P2_R1131_U82 );
nand NAND2_18611 ( P2_R1131_U445 , P2_U3974 , P2_R1131_U83 );
nand NAND2_18612 ( P2_R1131_U446 , P2_R1131_U445 , P2_R1131_U444 );
nand NAND2_18613 ( P2_R1131_U447 , P2_R1131_U158 , P2_R1131_U159 );
nand NAND2_18614 ( P2_R1131_U448 , P2_R1131_U286 , P2_R1131_U446 );
nand NAND2_18615 ( P2_R1131_U449 , P2_U3075 , P2_R1131_U54 );
nand NAND2_18616 ( P2_R1131_U450 , P2_U3975 , P2_R1131_U55 );
nand NAND2_18617 ( P2_R1131_U451 , P2_U3075 , P2_R1131_U54 );
nand NAND2_18618 ( P2_R1131_U452 , P2_U3975 , P2_R1131_U55 );
nand NAND2_18619 ( P2_R1131_U453 , P2_R1131_U452 , P2_R1131_U451 );
nand NAND2_18620 ( P2_R1131_U454 , P2_U3076 , P2_R1131_U81 );
nand NAND2_18621 ( P2_R1131_U455 , P2_U3976 , P2_R1131_U90 );
nand NAND2_18622 ( P2_R1131_U456 , P2_R1131_U182 , P2_R1131_U161 );
nand NAND2_18623 ( P2_R1131_U457 , P2_R1131_U328 , P2_R1131_U31 );
nand NAND2_18624 ( P2_R1131_U458 , P2_U3081 , P2_R1131_U78 );
nand NAND2_18625 ( P2_R1131_U459 , P2_U3506 , P2_R1131_U79 );
nand NAND2_18626 ( P2_R1131_U460 , P2_R1131_U459 , P2_R1131_U458 );
nand NAND2_18627 ( P2_R1131_U461 , P2_R1131_U359 , P2_R1131_U91 );
nand NAND2_18628 ( P2_R1131_U462 , P2_R1131_U460 , P2_R1131_U316 );
nand NAND2_18629 ( P2_R1131_U463 , P2_U3082 , P2_R1131_U75 );
nand NAND2_18630 ( P2_R1131_U464 , P2_U3504 , P2_R1131_U76 );
nand NAND2_18631 ( P2_R1131_U465 , P2_R1131_U464 , P2_R1131_U463 );
nand NAND2_18632 ( P2_R1131_U466 , P2_R1131_U360 , P2_R1131_U162 );
nand NAND2_18633 ( P2_R1131_U467 , P2_R1131_U270 , P2_R1131_U465 );
nand NAND2_18634 ( P2_R1131_U468 , P2_U3069 , P2_R1131_U60 );
nand NAND2_18635 ( P2_R1131_U469 , P2_U3501 , P2_R1131_U58 );
nand NAND2_18636 ( P2_R1131_U470 , P2_U3073 , P2_R1131_U56 );
nand NAND2_18637 ( P2_R1131_U471 , P2_U3498 , P2_R1131_U57 );
nand NAND2_18638 ( P2_R1131_U472 , P2_R1131_U471 , P2_R1131_U470 );
nand NAND2_18639 ( P2_R1131_U473 , P2_R1131_U361 , P2_R1131_U92 );
nand NAND2_18640 ( P2_R1131_U474 , P2_R1131_U472 , P2_R1131_U262 );
nand NAND2_18641 ( P2_R1131_U475 , P2_U3074 , P2_R1131_U73 );
nand NAND2_18642 ( P2_R1131_U476 , P2_U3495 , P2_R1131_U74 );
nand NAND2_18643 ( P2_R1131_U477 , P2_U3074 , P2_R1131_U73 );
nand NAND2_18644 ( P2_R1131_U478 , P2_U3495 , P2_R1131_U74 );
nand NAND2_18645 ( P2_R1131_U479 , P2_R1131_U478 , P2_R1131_U477 );
nand NAND2_18646 ( P2_R1131_U480 , P2_R1131_U163 , P2_R1131_U164 );
nand NAND2_18647 ( P2_R1131_U481 , P2_R1131_U258 , P2_R1131_U479 );
nand NAND2_18648 ( P2_R1131_U482 , P2_U3079 , P2_R1131_U71 );
nand NAND2_18649 ( P2_R1131_U483 , P2_U3492 , P2_R1131_U72 );
nand NAND2_18650 ( P2_R1131_U484 , P2_U3079 , P2_R1131_U71 );
nand NAND2_18651 ( P2_R1131_U485 , P2_U3492 , P2_R1131_U72 );
nand NAND2_18652 ( P2_R1131_U486 , P2_R1131_U485 , P2_R1131_U484 );
nand NAND2_18653 ( P2_R1131_U487 , P2_R1131_U165 , P2_R1131_U166 );
nand NAND2_18654 ( P2_R1131_U488 , P2_R1131_U254 , P2_R1131_U486 );
nand NAND2_18655 ( P2_R1131_U489 , P2_U3080 , P2_R1131_U69 );
nand NAND2_18656 ( P2_R1131_U490 , P2_U3489 , P2_R1131_U70 );
nand NAND2_18657 ( P2_R1131_U491 , P2_U3072 , P2_R1131_U64 );
nand NAND2_18658 ( P2_R1131_U492 , P2_U3486 , P2_R1131_U65 );
nand NAND2_18659 ( P2_R1131_U493 , P2_R1131_U492 , P2_R1131_U491 );
nand NAND2_18660 ( P2_R1131_U494 , P2_R1131_U362 , P2_R1131_U93 );
nand NAND2_18661 ( P2_R1131_U495 , P2_R1131_U493 , P2_R1131_U338 );
nand NAND2_18662 ( P2_R1131_U496 , P2_U3063 , P2_R1131_U66 );
nand NAND2_18663 ( P2_R1131_U497 , P2_U3483 , P2_R1131_U67 );
nand NAND2_18664 ( P2_R1131_U498 , P2_R1131_U497 , P2_R1131_U496 );
nand NAND2_18665 ( P2_R1131_U499 , P2_R1131_U363 , P2_R1131_U167 );
nand NAND2_18666 ( P2_R1131_U500 , P2_R1131_U244 , P2_R1131_U498 );
nand NAND2_18667 ( P2_R1131_U501 , P2_U3062 , P2_R1131_U62 );
nand NAND2_18668 ( P2_R1131_U502 , P2_U3480 , P2_R1131_U63 );
nand NAND2_18669 ( P2_R1131_U503 , P2_U3077 , P2_R1131_U29 );
nand NAND2_18670 ( P2_R1131_U504 , P2_U3448 , P2_R1131_U30 );
and AND2_18671 ( P2_R1146_U6 , P2_R1146_U205 , P2_R1146_U204 );
and AND2_18672 ( P2_R1146_U7 , P2_R1146_U244 , P2_R1146_U243 );
and AND2_18673 ( P2_R1146_U8 , P2_R1146_U261 , P2_R1146_U260 );
and AND2_18674 ( P2_R1146_U9 , P2_R1146_U285 , P2_R1146_U284 );
and AND2_18675 ( P2_R1146_U10 , P2_R1146_U384 , P2_R1146_U383 );
nand NAND2_18676 ( P2_R1146_U11 , P2_R1146_U340 , P2_R1146_U343 );
nand NAND2_18677 ( P2_R1146_U12 , P2_R1146_U329 , P2_R1146_U332 );
nand NAND2_18678 ( P2_R1146_U13 , P2_R1146_U318 , P2_R1146_U321 );
nand NAND2_18679 ( P2_R1146_U14 , P2_R1146_U310 , P2_R1146_U312 );
nand NAND3_18680 ( P2_R1146_U15 , P2_R1146_U349 , P2_R1146_U177 , P2_R1146_U156 );
nand NAND2_18681 ( P2_R1146_U16 , P2_R1146_U238 , P2_R1146_U240 );
nand NAND2_18682 ( P2_R1146_U17 , P2_R1146_U230 , P2_R1146_U233 );
nand NAND2_18683 ( P2_R1146_U18 , P2_R1146_U222 , P2_R1146_U224 );
nand NAND2_18684 ( P2_R1146_U19 , P2_R1146_U166 , P2_R1146_U346 );
not NOT1_18685 ( P2_R1146_U20 , P2_U3471 );
not NOT1_18686 ( P2_R1146_U21 , P2_U3465 );
not NOT1_18687 ( P2_R1146_U22 , P2_U3456 );
not NOT1_18688 ( P2_R1146_U23 , P2_U3448 );
not NOT1_18689 ( P2_R1146_U24 , P2_U3078 );
not NOT1_18690 ( P2_R1146_U25 , P2_U3459 );
not NOT1_18691 ( P2_R1146_U26 , P2_U3068 );
nand NAND2_18692 ( P2_R1146_U27 , P2_U3068 , P2_R1146_U22 );
not NOT1_18693 ( P2_R1146_U28 , P2_U3064 );
not NOT1_18694 ( P2_R1146_U29 , P2_U3468 );
not NOT1_18695 ( P2_R1146_U30 , P2_U3462 );
not NOT1_18696 ( P2_R1146_U31 , P2_U3071 );
not NOT1_18697 ( P2_R1146_U32 , P2_U3067 );
not NOT1_18698 ( P2_R1146_U33 , P2_U3060 );
nand NAND2_18699 ( P2_R1146_U34 , P2_U3060 , P2_R1146_U30 );
not NOT1_18700 ( P2_R1146_U35 , P2_U3474 );
not NOT1_18701 ( P2_R1146_U36 , P2_U3070 );
nand NAND2_18702 ( P2_R1146_U37 , P2_U3070 , P2_R1146_U20 );
not NOT1_18703 ( P2_R1146_U38 , P2_U3084 );
not NOT1_18704 ( P2_R1146_U39 , P2_U3477 );
not NOT1_18705 ( P2_R1146_U40 , P2_U3083 );
nand NAND2_18706 ( P2_R1146_U41 , P2_R1146_U211 , P2_R1146_U210 );
nand NAND2_18707 ( P2_R1146_U42 , P2_R1146_U34 , P2_R1146_U226 );
nand NAND3_18708 ( P2_R1146_U43 , P2_R1146_U195 , P2_R1146_U179 , P2_R1146_U347 );
not NOT1_18709 ( P2_R1146_U44 , P2_U3970 );
not NOT1_18710 ( P2_R1146_U45 , P2_U3974 );
not NOT1_18711 ( P2_R1146_U46 , P2_U3495 );
not NOT1_18712 ( P2_R1146_U47 , P2_U3480 );
not NOT1_18713 ( P2_R1146_U48 , P2_U3483 );
not NOT1_18714 ( P2_R1146_U49 , P2_U3063 );
not NOT1_18715 ( P2_R1146_U50 , P2_U3062 );
nand NAND2_18716 ( P2_R1146_U51 , P2_U3083 , P2_R1146_U39 );
not NOT1_18717 ( P2_R1146_U52 , P2_U3486 );
not NOT1_18718 ( P2_R1146_U53 , P2_U3072 );
not NOT1_18719 ( P2_R1146_U54 , P2_U3489 );
not NOT1_18720 ( P2_R1146_U55 , P2_U3080 );
not NOT1_18721 ( P2_R1146_U56 , P2_U3498 );
not NOT1_18722 ( P2_R1146_U57 , P2_U3492 );
not NOT1_18723 ( P2_R1146_U58 , P2_U3073 );
not NOT1_18724 ( P2_R1146_U59 , P2_U3074 );
not NOT1_18725 ( P2_R1146_U60 , P2_U3079 );
nand NAND2_18726 ( P2_R1146_U61 , P2_U3079 , P2_R1146_U57 );
not NOT1_18727 ( P2_R1146_U62 , P2_U3501 );
not NOT1_18728 ( P2_R1146_U63 , P2_U3069 );
not NOT1_18729 ( P2_R1146_U64 , P2_U3082 );
not NOT1_18730 ( P2_R1146_U65 , P2_U3506 );
not NOT1_18731 ( P2_R1146_U66 , P2_U3081 );
not NOT1_18732 ( P2_R1146_U67 , P2_U3976 );
not NOT1_18733 ( P2_R1146_U68 , P2_U3076 );
not NOT1_18734 ( P2_R1146_U69 , P2_U3973 );
not NOT1_18735 ( P2_R1146_U70 , P2_U3975 );
not NOT1_18736 ( P2_R1146_U71 , P2_U3066 );
not NOT1_18737 ( P2_R1146_U72 , P2_U3061 );
not NOT1_18738 ( P2_R1146_U73 , P2_U3075 );
nand NAND2_18739 ( P2_R1146_U74 , P2_U3075 , P2_R1146_U70 );
not NOT1_18740 ( P2_R1146_U75 , P2_U3972 );
not NOT1_18741 ( P2_R1146_U76 , P2_U3065 );
not NOT1_18742 ( P2_R1146_U77 , P2_U3971 );
not NOT1_18743 ( P2_R1146_U78 , P2_U3058 );
not NOT1_18744 ( P2_R1146_U79 , P2_U3969 );
not NOT1_18745 ( P2_R1146_U80 , P2_U3057 );
nand NAND2_18746 ( P2_R1146_U81 , P2_U3057 , P2_R1146_U44 );
not NOT1_18747 ( P2_R1146_U82 , P2_U3053 );
not NOT1_18748 ( P2_R1146_U83 , P2_U3968 );
not NOT1_18749 ( P2_R1146_U84 , P2_U3054 );
nand NAND2_18750 ( P2_R1146_U85 , P2_R1146_U299 , P2_R1146_U298 );
nand NAND2_18751 ( P2_R1146_U86 , P2_R1146_U74 , P2_R1146_U314 );
nand NAND2_18752 ( P2_R1146_U87 , P2_R1146_U61 , P2_R1146_U325 );
nand NAND2_18753 ( P2_R1146_U88 , P2_R1146_U51 , P2_R1146_U336 );
not NOT1_18754 ( P2_R1146_U89 , P2_U3077 );
nand NAND2_18755 ( P2_R1146_U90 , P2_R1146_U394 , P2_R1146_U393 );
nand NAND2_18756 ( P2_R1146_U91 , P2_R1146_U408 , P2_R1146_U407 );
nand NAND2_18757 ( P2_R1146_U92 , P2_R1146_U413 , P2_R1146_U412 );
nand NAND2_18758 ( P2_R1146_U93 , P2_R1146_U429 , P2_R1146_U428 );
nand NAND2_18759 ( P2_R1146_U94 , P2_R1146_U434 , P2_R1146_U433 );
nand NAND2_18760 ( P2_R1146_U95 , P2_R1146_U439 , P2_R1146_U438 );
nand NAND2_18761 ( P2_R1146_U96 , P2_R1146_U444 , P2_R1146_U443 );
nand NAND2_18762 ( P2_R1146_U97 , P2_R1146_U449 , P2_R1146_U448 );
nand NAND2_18763 ( P2_R1146_U98 , P2_R1146_U465 , P2_R1146_U464 );
nand NAND2_18764 ( P2_R1146_U99 , P2_R1146_U470 , P2_R1146_U469 );
nand NAND2_18765 ( P2_R1146_U100 , P2_R1146_U353 , P2_R1146_U352 );
nand NAND2_18766 ( P2_R1146_U101 , P2_R1146_U362 , P2_R1146_U361 );
nand NAND2_18767 ( P2_R1146_U102 , P2_R1146_U369 , P2_R1146_U368 );
nand NAND2_18768 ( P2_R1146_U103 , P2_R1146_U373 , P2_R1146_U372 );
nand NAND2_18769 ( P2_R1146_U104 , P2_R1146_U382 , P2_R1146_U381 );
nand NAND2_18770 ( P2_R1146_U105 , P2_R1146_U403 , P2_R1146_U402 );
nand NAND2_18771 ( P2_R1146_U106 , P2_R1146_U420 , P2_R1146_U419 );
nand NAND2_18772 ( P2_R1146_U107 , P2_R1146_U424 , P2_R1146_U423 );
nand NAND2_18773 ( P2_R1146_U108 , P2_R1146_U456 , P2_R1146_U455 );
nand NAND2_18774 ( P2_R1146_U109 , P2_R1146_U460 , P2_R1146_U459 );
nand NAND2_18775 ( P2_R1146_U110 , P2_R1146_U477 , P2_R1146_U476 );
and AND2_18776 ( P2_R1146_U111 , P2_R1146_U197 , P2_R1146_U187 );
and AND2_18777 ( P2_R1146_U112 , P2_R1146_U200 , P2_R1146_U201 );
and AND3_18778 ( P2_R1146_U113 , P2_R1146_U208 , P2_R1146_U203 , P2_R1146_U188 );
and AND2_18779 ( P2_R1146_U114 , P2_R1146_U213 , P2_R1146_U189 );
and AND2_18780 ( P2_R1146_U115 , P2_R1146_U216 , P2_R1146_U217 );
and AND3_18781 ( P2_R1146_U116 , P2_R1146_U355 , P2_R1146_U354 , P2_R1146_U37 );
and AND2_18782 ( P2_R1146_U117 , P2_R1146_U358 , P2_R1146_U189 );
and AND2_18783 ( P2_R1146_U118 , P2_R1146_U232 , P2_R1146_U6 );
and AND2_18784 ( P2_R1146_U119 , P2_R1146_U365 , P2_R1146_U188 );
and AND3_18785 ( P2_R1146_U120 , P2_R1146_U375 , P2_R1146_U374 , P2_R1146_U27 );
and AND2_18786 ( P2_R1146_U121 , P2_R1146_U378 , P2_R1146_U187 );
and AND3_18787 ( P2_R1146_U122 , P2_R1146_U242 , P2_R1146_U219 , P2_R1146_U183 );
and AND3_18788 ( P2_R1146_U123 , P2_R1146_U264 , P2_R1146_U184 , P2_R1146_U259 );
and AND3_18789 ( P2_R1146_U124 , P2_R1146_U288 , P2_R1146_U185 , P2_R1146_U283 );
and AND2_18790 ( P2_R1146_U125 , P2_R1146_U301 , P2_R1146_U186 );
and AND2_18791 ( P2_R1146_U126 , P2_R1146_U304 , P2_R1146_U305 );
and AND2_18792 ( P2_R1146_U127 , P2_R1146_U304 , P2_R1146_U305 );
and AND2_18793 ( P2_R1146_U128 , P2_R1146_U10 , P2_R1146_U308 );
nand NAND2_18794 ( P2_R1146_U129 , P2_R1146_U391 , P2_R1146_U390 );
and AND3_18795 ( P2_R1146_U130 , P2_R1146_U396 , P2_R1146_U395 , P2_R1146_U81 );
and AND2_18796 ( P2_R1146_U131 , P2_R1146_U399 , P2_R1146_U186 );
nand NAND2_18797 ( P2_R1146_U132 , P2_R1146_U405 , P2_R1146_U404 );
nand NAND2_18798 ( P2_R1146_U133 , P2_R1146_U410 , P2_R1146_U409 );
and AND2_18799 ( P2_R1146_U134 , P2_R1146_U320 , P2_R1146_U9 );
and AND2_18800 ( P2_R1146_U135 , P2_R1146_U416 , P2_R1146_U185 );
nand NAND2_18801 ( P2_R1146_U136 , P2_R1146_U426 , P2_R1146_U425 );
nand NAND2_18802 ( P2_R1146_U137 , P2_R1146_U431 , P2_R1146_U430 );
nand NAND2_18803 ( P2_R1146_U138 , P2_R1146_U436 , P2_R1146_U435 );
nand NAND2_18804 ( P2_R1146_U139 , P2_R1146_U441 , P2_R1146_U440 );
nand NAND2_18805 ( P2_R1146_U140 , P2_R1146_U446 , P2_R1146_U445 );
and AND2_18806 ( P2_R1146_U141 , P2_R1146_U331 , P2_R1146_U8 );
and AND2_18807 ( P2_R1146_U142 , P2_R1146_U452 , P2_R1146_U184 );
nand NAND2_18808 ( P2_R1146_U143 , P2_R1146_U462 , P2_R1146_U461 );
nand NAND2_18809 ( P2_R1146_U144 , P2_R1146_U467 , P2_R1146_U466 );
and AND2_18810 ( P2_R1146_U145 , P2_R1146_U342 , P2_R1146_U7 );
and AND2_18811 ( P2_R1146_U146 , P2_R1146_U473 , P2_R1146_U183 );
and AND2_18812 ( P2_R1146_U147 , P2_R1146_U351 , P2_R1146_U350 );
nand NAND2_18813 ( P2_R1146_U148 , P2_R1146_U115 , P2_R1146_U214 );
and AND2_18814 ( P2_R1146_U149 , P2_R1146_U360 , P2_R1146_U359 );
and AND2_18815 ( P2_R1146_U150 , P2_R1146_U367 , P2_R1146_U366 );
and AND2_18816 ( P2_R1146_U151 , P2_R1146_U371 , P2_R1146_U370 );
nand NAND2_18817 ( P2_R1146_U152 , P2_R1146_U112 , P2_R1146_U198 );
and AND2_18818 ( P2_R1146_U153 , P2_R1146_U380 , P2_R1146_U379 );
not NOT1_18819 ( P2_R1146_U154 , P2_U3979 );
not NOT1_18820 ( P2_R1146_U155 , P2_U3055 );
and AND2_18821 ( P2_R1146_U156 , P2_R1146_U389 , P2_R1146_U388 );
nand NAND2_18822 ( P2_R1146_U157 , P2_R1146_U126 , P2_R1146_U302 );
and AND2_18823 ( P2_R1146_U158 , P2_R1146_U401 , P2_R1146_U400 );
nand NAND2_18824 ( P2_R1146_U159 , P2_R1146_U295 , P2_R1146_U294 );
nand NAND2_18825 ( P2_R1146_U160 , P2_R1146_U291 , P2_R1146_U290 );
and AND2_18826 ( P2_R1146_U161 , P2_R1146_U418 , P2_R1146_U417 );
and AND2_18827 ( P2_R1146_U162 , P2_R1146_U422 , P2_R1146_U421 );
nand NAND2_18828 ( P2_R1146_U163 , P2_R1146_U281 , P2_R1146_U280 );
nand NAND2_18829 ( P2_R1146_U164 , P2_R1146_U277 , P2_R1146_U276 );
not NOT1_18830 ( P2_R1146_U165 , P2_U3453 );
nand NAND2_18831 ( P2_R1146_U166 , P2_U3448 , P2_R1146_U89 );
nand NAND3_18832 ( P2_R1146_U167 , P2_R1146_U273 , P2_R1146_U178 , P2_R1146_U348 );
not NOT1_18833 ( P2_R1146_U168 , P2_U3504 );
nand NAND2_18834 ( P2_R1146_U169 , P2_R1146_U271 , P2_R1146_U270 );
nand NAND2_18835 ( P2_R1146_U170 , P2_R1146_U267 , P2_R1146_U266 );
and AND2_18836 ( P2_R1146_U171 , P2_R1146_U454 , P2_R1146_U453 );
and AND2_18837 ( P2_R1146_U172 , P2_R1146_U458 , P2_R1146_U457 );
nand NAND2_18838 ( P2_R1146_U173 , P2_R1146_U257 , P2_R1146_U256 );
nand NAND2_18839 ( P2_R1146_U174 , P2_R1146_U253 , P2_R1146_U252 );
nand NAND2_18840 ( P2_R1146_U175 , P2_R1146_U249 , P2_R1146_U248 );
and AND2_18841 ( P2_R1146_U176 , P2_R1146_U475 , P2_R1146_U474 );
nand NAND3_18842 ( P2_R1146_U177 , P2_R1146_U307 , P2_R1146_U157 , P2_R1146_U387 );
nand NAND2_18843 ( P2_R1146_U178 , P2_R1146_U169 , P2_R1146_U168 );
nand NAND2_18844 ( P2_R1146_U179 , P2_R1146_U166 , P2_R1146_U165 );
not NOT1_18845 ( P2_R1146_U180 , P2_R1146_U81 );
not NOT1_18846 ( P2_R1146_U181 , P2_R1146_U27 );
not NOT1_18847 ( P2_R1146_U182 , P2_R1146_U37 );
nand NAND2_18848 ( P2_R1146_U183 , P2_U3480 , P2_R1146_U50 );
nand NAND2_18849 ( P2_R1146_U184 , P2_U3495 , P2_R1146_U59 );
nand NAND2_18850 ( P2_R1146_U185 , P2_U3974 , P2_R1146_U72 );
nand NAND2_18851 ( P2_R1146_U186 , P2_U3970 , P2_R1146_U80 );
nand NAND2_18852 ( P2_R1146_U187 , P2_U3456 , P2_R1146_U26 );
nand NAND2_18853 ( P2_R1146_U188 , P2_U3465 , P2_R1146_U32 );
nand NAND2_18854 ( P2_R1146_U189 , P2_U3471 , P2_R1146_U36 );
not NOT1_18855 ( P2_R1146_U190 , P2_R1146_U61 );
not NOT1_18856 ( P2_R1146_U191 , P2_R1146_U74 );
not NOT1_18857 ( P2_R1146_U192 , P2_R1146_U34 );
not NOT1_18858 ( P2_R1146_U193 , P2_R1146_U51 );
not NOT1_18859 ( P2_R1146_U194 , P2_R1146_U166 );
nand NAND2_18860 ( P2_R1146_U195 , P2_U3078 , P2_R1146_U166 );
not NOT1_18861 ( P2_R1146_U196 , P2_R1146_U43 );
nand NAND2_18862 ( P2_R1146_U197 , P2_U3459 , P2_R1146_U28 );
nand NAND2_18863 ( P2_R1146_U198 , P2_R1146_U111 , P2_R1146_U43 );
nand NAND2_18864 ( P2_R1146_U199 , P2_R1146_U28 , P2_R1146_U27 );
nand NAND2_18865 ( P2_R1146_U200 , P2_R1146_U199 , P2_R1146_U25 );
nand NAND2_18866 ( P2_R1146_U201 , P2_U3064 , P2_R1146_U181 );
not NOT1_18867 ( P2_R1146_U202 , P2_R1146_U152 );
nand NAND2_18868 ( P2_R1146_U203 , P2_U3468 , P2_R1146_U31 );
nand NAND2_18869 ( P2_R1146_U204 , P2_U3071 , P2_R1146_U29 );
nand NAND2_18870 ( P2_R1146_U205 , P2_U3067 , P2_R1146_U21 );
nand NAND2_18871 ( P2_R1146_U206 , P2_R1146_U192 , P2_R1146_U188 );
nand NAND2_18872 ( P2_R1146_U207 , P2_R1146_U6 , P2_R1146_U206 );
nand NAND2_18873 ( P2_R1146_U208 , P2_U3462 , P2_R1146_U33 );
nand NAND2_18874 ( P2_R1146_U209 , P2_U3468 , P2_R1146_U31 );
nand NAND2_18875 ( P2_R1146_U210 , P2_R1146_U152 , P2_R1146_U113 );
nand NAND2_18876 ( P2_R1146_U211 , P2_R1146_U209 , P2_R1146_U207 );
not NOT1_18877 ( P2_R1146_U212 , P2_R1146_U41 );
nand NAND2_18878 ( P2_R1146_U213 , P2_U3474 , P2_R1146_U38 );
nand NAND2_18879 ( P2_R1146_U214 , P2_R1146_U114 , P2_R1146_U41 );
nand NAND2_18880 ( P2_R1146_U215 , P2_R1146_U38 , P2_R1146_U37 );
nand NAND2_18881 ( P2_R1146_U216 , P2_R1146_U215 , P2_R1146_U35 );
nand NAND2_18882 ( P2_R1146_U217 , P2_U3084 , P2_R1146_U182 );
not NOT1_18883 ( P2_R1146_U218 , P2_R1146_U148 );
nand NAND2_18884 ( P2_R1146_U219 , P2_U3477 , P2_R1146_U40 );
nand NAND2_18885 ( P2_R1146_U220 , P2_R1146_U219 , P2_R1146_U51 );
nand NAND2_18886 ( P2_R1146_U221 , P2_R1146_U212 , P2_R1146_U37 );
nand NAND2_18887 ( P2_R1146_U222 , P2_R1146_U117 , P2_R1146_U221 );
nand NAND2_18888 ( P2_R1146_U223 , P2_R1146_U41 , P2_R1146_U189 );
nand NAND2_18889 ( P2_R1146_U224 , P2_R1146_U116 , P2_R1146_U223 );
nand NAND2_18890 ( P2_R1146_U225 , P2_R1146_U37 , P2_R1146_U189 );
nand NAND2_18891 ( P2_R1146_U226 , P2_R1146_U208 , P2_R1146_U152 );
not NOT1_18892 ( P2_R1146_U227 , P2_R1146_U42 );
nand NAND2_18893 ( P2_R1146_U228 , P2_U3067 , P2_R1146_U21 );
nand NAND2_18894 ( P2_R1146_U229 , P2_R1146_U227 , P2_R1146_U228 );
nand NAND2_18895 ( P2_R1146_U230 , P2_R1146_U119 , P2_R1146_U229 );
nand NAND2_18896 ( P2_R1146_U231 , P2_R1146_U42 , P2_R1146_U188 );
nand NAND2_18897 ( P2_R1146_U232 , P2_U3468 , P2_R1146_U31 );
nand NAND2_18898 ( P2_R1146_U233 , P2_R1146_U118 , P2_R1146_U231 );
nand NAND2_18899 ( P2_R1146_U234 , P2_U3067 , P2_R1146_U21 );
nand NAND2_18900 ( P2_R1146_U235 , P2_R1146_U188 , P2_R1146_U234 );
nand NAND2_18901 ( P2_R1146_U236 , P2_R1146_U208 , P2_R1146_U34 );
nand NAND2_18902 ( P2_R1146_U237 , P2_R1146_U196 , P2_R1146_U27 );
nand NAND2_18903 ( P2_R1146_U238 , P2_R1146_U121 , P2_R1146_U237 );
nand NAND2_18904 ( P2_R1146_U239 , P2_R1146_U43 , P2_R1146_U187 );
nand NAND2_18905 ( P2_R1146_U240 , P2_R1146_U120 , P2_R1146_U239 );
nand NAND2_18906 ( P2_R1146_U241 , P2_R1146_U27 , P2_R1146_U187 );
nand NAND2_18907 ( P2_R1146_U242 , P2_U3483 , P2_R1146_U49 );
nand NAND2_18908 ( P2_R1146_U243 , P2_U3063 , P2_R1146_U48 );
nand NAND2_18909 ( P2_R1146_U244 , P2_U3062 , P2_R1146_U47 );
nand NAND2_18910 ( P2_R1146_U245 , P2_R1146_U193 , P2_R1146_U183 );
nand NAND2_18911 ( P2_R1146_U246 , P2_R1146_U7 , P2_R1146_U245 );
nand NAND2_18912 ( P2_R1146_U247 , P2_U3483 , P2_R1146_U49 );
nand NAND2_18913 ( P2_R1146_U248 , P2_R1146_U148 , P2_R1146_U122 );
nand NAND2_18914 ( P2_R1146_U249 , P2_R1146_U247 , P2_R1146_U246 );
not NOT1_18915 ( P2_R1146_U250 , P2_R1146_U175 );
nand NAND2_18916 ( P2_R1146_U251 , P2_U3486 , P2_R1146_U53 );
nand NAND2_18917 ( P2_R1146_U252 , P2_R1146_U251 , P2_R1146_U175 );
nand NAND2_18918 ( P2_R1146_U253 , P2_U3072 , P2_R1146_U52 );
not NOT1_18919 ( P2_R1146_U254 , P2_R1146_U174 );
nand NAND2_18920 ( P2_R1146_U255 , P2_U3489 , P2_R1146_U55 );
nand NAND2_18921 ( P2_R1146_U256 , P2_R1146_U255 , P2_R1146_U174 );
nand NAND2_18922 ( P2_R1146_U257 , P2_U3080 , P2_R1146_U54 );
not NOT1_18923 ( P2_R1146_U258 , P2_R1146_U173 );
nand NAND2_18924 ( P2_R1146_U259 , P2_U3498 , P2_R1146_U58 );
nand NAND2_18925 ( P2_R1146_U260 , P2_U3073 , P2_R1146_U56 );
nand NAND2_18926 ( P2_R1146_U261 , P2_U3074 , P2_R1146_U46 );
nand NAND2_18927 ( P2_R1146_U262 , P2_R1146_U190 , P2_R1146_U184 );
nand NAND2_18928 ( P2_R1146_U263 , P2_R1146_U8 , P2_R1146_U262 );
nand NAND2_18929 ( P2_R1146_U264 , P2_U3492 , P2_R1146_U60 );
nand NAND2_18930 ( P2_R1146_U265 , P2_U3498 , P2_R1146_U58 );
nand NAND2_18931 ( P2_R1146_U266 , P2_R1146_U173 , P2_R1146_U123 );
nand NAND2_18932 ( P2_R1146_U267 , P2_R1146_U265 , P2_R1146_U263 );
not NOT1_18933 ( P2_R1146_U268 , P2_R1146_U170 );
nand NAND2_18934 ( P2_R1146_U269 , P2_U3501 , P2_R1146_U63 );
nand NAND2_18935 ( P2_R1146_U270 , P2_R1146_U269 , P2_R1146_U170 );
nand NAND2_18936 ( P2_R1146_U271 , P2_U3069 , P2_R1146_U62 );
not NOT1_18937 ( P2_R1146_U272 , P2_R1146_U169 );
nand NAND2_18938 ( P2_R1146_U273 , P2_U3082 , P2_R1146_U169 );
not NOT1_18939 ( P2_R1146_U274 , P2_R1146_U167 );
nand NAND2_18940 ( P2_R1146_U275 , P2_U3506 , P2_R1146_U66 );
nand NAND2_18941 ( P2_R1146_U276 , P2_R1146_U275 , P2_R1146_U167 );
nand NAND2_18942 ( P2_R1146_U277 , P2_U3081 , P2_R1146_U65 );
not NOT1_18943 ( P2_R1146_U278 , P2_R1146_U164 );
nand NAND2_18944 ( P2_R1146_U279 , P2_U3976 , P2_R1146_U68 );
nand NAND2_18945 ( P2_R1146_U280 , P2_R1146_U279 , P2_R1146_U164 );
nand NAND2_18946 ( P2_R1146_U281 , P2_U3076 , P2_R1146_U67 );
not NOT1_18947 ( P2_R1146_U282 , P2_R1146_U163 );
nand NAND2_18948 ( P2_R1146_U283 , P2_U3973 , P2_R1146_U71 );
nand NAND2_18949 ( P2_R1146_U284 , P2_U3066 , P2_R1146_U69 );
nand NAND2_18950 ( P2_R1146_U285 , P2_U3061 , P2_R1146_U45 );
nand NAND2_18951 ( P2_R1146_U286 , P2_R1146_U191 , P2_R1146_U185 );
nand NAND2_18952 ( P2_R1146_U287 , P2_R1146_U9 , P2_R1146_U286 );
nand NAND2_18953 ( P2_R1146_U288 , P2_U3975 , P2_R1146_U73 );
nand NAND2_18954 ( P2_R1146_U289 , P2_U3973 , P2_R1146_U71 );
nand NAND2_18955 ( P2_R1146_U290 , P2_R1146_U163 , P2_R1146_U124 );
nand NAND2_18956 ( P2_R1146_U291 , P2_R1146_U289 , P2_R1146_U287 );
not NOT1_18957 ( P2_R1146_U292 , P2_R1146_U160 );
nand NAND2_18958 ( P2_R1146_U293 , P2_U3972 , P2_R1146_U76 );
nand NAND2_18959 ( P2_R1146_U294 , P2_R1146_U293 , P2_R1146_U160 );
nand NAND2_18960 ( P2_R1146_U295 , P2_U3065 , P2_R1146_U75 );
not NOT1_18961 ( P2_R1146_U296 , P2_R1146_U159 );
nand NAND2_18962 ( P2_R1146_U297 , P2_U3971 , P2_R1146_U78 );
nand NAND2_18963 ( P2_R1146_U298 , P2_R1146_U297 , P2_R1146_U159 );
nand NAND2_18964 ( P2_R1146_U299 , P2_U3058 , P2_R1146_U77 );
not NOT1_18965 ( P2_R1146_U300 , P2_R1146_U85 );
nand NAND2_18966 ( P2_R1146_U301 , P2_U3969 , P2_R1146_U82 );
nand NAND2_18967 ( P2_R1146_U302 , P2_R1146_U125 , P2_R1146_U85 );
nand NAND2_18968 ( P2_R1146_U303 , P2_R1146_U82 , P2_R1146_U81 );
nand NAND2_18969 ( P2_R1146_U304 , P2_R1146_U303 , P2_R1146_U79 );
nand NAND2_18970 ( P2_R1146_U305 , P2_U3053 , P2_R1146_U180 );
not NOT1_18971 ( P2_R1146_U306 , P2_R1146_U157 );
nand NAND2_18972 ( P2_R1146_U307 , P2_U3968 , P2_R1146_U84 );
nand NAND2_18973 ( P2_R1146_U308 , P2_U3054 , P2_R1146_U83 );
nand NAND2_18974 ( P2_R1146_U309 , P2_R1146_U300 , P2_R1146_U81 );
nand NAND2_18975 ( P2_R1146_U310 , P2_R1146_U131 , P2_R1146_U309 );
nand NAND2_18976 ( P2_R1146_U311 , P2_R1146_U85 , P2_R1146_U186 );
nand NAND2_18977 ( P2_R1146_U312 , P2_R1146_U130 , P2_R1146_U311 );
nand NAND2_18978 ( P2_R1146_U313 , P2_R1146_U81 , P2_R1146_U186 );
nand NAND2_18979 ( P2_R1146_U314 , P2_R1146_U288 , P2_R1146_U163 );
not NOT1_18980 ( P2_R1146_U315 , P2_R1146_U86 );
nand NAND2_18981 ( P2_R1146_U316 , P2_U3061 , P2_R1146_U45 );
nand NAND2_18982 ( P2_R1146_U317 , P2_R1146_U315 , P2_R1146_U316 );
nand NAND2_18983 ( P2_R1146_U318 , P2_R1146_U135 , P2_R1146_U317 );
nand NAND2_18984 ( P2_R1146_U319 , P2_R1146_U86 , P2_R1146_U185 );
nand NAND2_18985 ( P2_R1146_U320 , P2_U3973 , P2_R1146_U71 );
nand NAND2_18986 ( P2_R1146_U321 , P2_R1146_U134 , P2_R1146_U319 );
nand NAND2_18987 ( P2_R1146_U322 , P2_U3061 , P2_R1146_U45 );
nand NAND2_18988 ( P2_R1146_U323 , P2_R1146_U185 , P2_R1146_U322 );
nand NAND2_18989 ( P2_R1146_U324 , P2_R1146_U288 , P2_R1146_U74 );
nand NAND2_18990 ( P2_R1146_U325 , P2_R1146_U264 , P2_R1146_U173 );
not NOT1_18991 ( P2_R1146_U326 , P2_R1146_U87 );
nand NAND2_18992 ( P2_R1146_U327 , P2_U3074 , P2_R1146_U46 );
nand NAND2_18993 ( P2_R1146_U328 , P2_R1146_U326 , P2_R1146_U327 );
nand NAND2_18994 ( P2_R1146_U329 , P2_R1146_U142 , P2_R1146_U328 );
nand NAND2_18995 ( P2_R1146_U330 , P2_R1146_U87 , P2_R1146_U184 );
nand NAND2_18996 ( P2_R1146_U331 , P2_U3498 , P2_R1146_U58 );
nand NAND2_18997 ( P2_R1146_U332 , P2_R1146_U141 , P2_R1146_U330 );
nand NAND2_18998 ( P2_R1146_U333 , P2_U3074 , P2_R1146_U46 );
nand NAND2_18999 ( P2_R1146_U334 , P2_R1146_U184 , P2_R1146_U333 );
nand NAND2_19000 ( P2_R1146_U335 , P2_R1146_U264 , P2_R1146_U61 );
nand NAND2_19001 ( P2_R1146_U336 , P2_R1146_U219 , P2_R1146_U148 );
not NOT1_19002 ( P2_R1146_U337 , P2_R1146_U88 );
nand NAND2_19003 ( P2_R1146_U338 , P2_U3062 , P2_R1146_U47 );
nand NAND2_19004 ( P2_R1146_U339 , P2_R1146_U337 , P2_R1146_U338 );
nand NAND2_19005 ( P2_R1146_U340 , P2_R1146_U146 , P2_R1146_U339 );
nand NAND2_19006 ( P2_R1146_U341 , P2_R1146_U88 , P2_R1146_U183 );
nand NAND2_19007 ( P2_R1146_U342 , P2_U3483 , P2_R1146_U49 );
nand NAND2_19008 ( P2_R1146_U343 , P2_R1146_U145 , P2_R1146_U341 );
nand NAND2_19009 ( P2_R1146_U344 , P2_U3062 , P2_R1146_U47 );
nand NAND2_19010 ( P2_R1146_U345 , P2_R1146_U183 , P2_R1146_U344 );
nand NAND2_19011 ( P2_R1146_U346 , P2_U3077 , P2_R1146_U23 );
nand NAND2_19012 ( P2_R1146_U347 , P2_U3078 , P2_R1146_U165 );
nand NAND2_19013 ( P2_R1146_U348 , P2_U3082 , P2_R1146_U168 );
nand NAND3_19014 ( P2_R1146_U349 , P2_R1146_U127 , P2_R1146_U302 , P2_R1146_U128 );
nand NAND2_19015 ( P2_R1146_U350 , P2_U3477 , P2_R1146_U40 );
nand NAND2_19016 ( P2_R1146_U351 , P2_U3083 , P2_R1146_U39 );
nand NAND2_19017 ( P2_R1146_U352 , P2_R1146_U220 , P2_R1146_U148 );
nand NAND2_19018 ( P2_R1146_U353 , P2_R1146_U218 , P2_R1146_U147 );
nand NAND2_19019 ( P2_R1146_U354 , P2_U3474 , P2_R1146_U38 );
nand NAND2_19020 ( P2_R1146_U355 , P2_U3084 , P2_R1146_U35 );
nand NAND2_19021 ( P2_R1146_U356 , P2_U3474 , P2_R1146_U38 );
nand NAND2_19022 ( P2_R1146_U357 , P2_U3084 , P2_R1146_U35 );
nand NAND2_19023 ( P2_R1146_U358 , P2_R1146_U357 , P2_R1146_U356 );
nand NAND2_19024 ( P2_R1146_U359 , P2_U3471 , P2_R1146_U36 );
nand NAND2_19025 ( P2_R1146_U360 , P2_U3070 , P2_R1146_U20 );
nand NAND2_19026 ( P2_R1146_U361 , P2_R1146_U225 , P2_R1146_U41 );
nand NAND2_19027 ( P2_R1146_U362 , P2_R1146_U149 , P2_R1146_U212 );
nand NAND2_19028 ( P2_R1146_U363 , P2_U3468 , P2_R1146_U31 );
nand NAND2_19029 ( P2_R1146_U364 , P2_U3071 , P2_R1146_U29 );
nand NAND2_19030 ( P2_R1146_U365 , P2_R1146_U364 , P2_R1146_U363 );
nand NAND2_19031 ( P2_R1146_U366 , P2_U3465 , P2_R1146_U32 );
nand NAND2_19032 ( P2_R1146_U367 , P2_U3067 , P2_R1146_U21 );
nand NAND2_19033 ( P2_R1146_U368 , P2_R1146_U235 , P2_R1146_U42 );
nand NAND2_19034 ( P2_R1146_U369 , P2_R1146_U150 , P2_R1146_U227 );
nand NAND2_19035 ( P2_R1146_U370 , P2_U3462 , P2_R1146_U33 );
nand NAND2_19036 ( P2_R1146_U371 , P2_U3060 , P2_R1146_U30 );
nand NAND2_19037 ( P2_R1146_U372 , P2_R1146_U236 , P2_R1146_U152 );
nand NAND2_19038 ( P2_R1146_U373 , P2_R1146_U202 , P2_R1146_U151 );
nand NAND2_19039 ( P2_R1146_U374 , P2_U3459 , P2_R1146_U28 );
nand NAND2_19040 ( P2_R1146_U375 , P2_U3064 , P2_R1146_U25 );
nand NAND2_19041 ( P2_R1146_U376 , P2_U3459 , P2_R1146_U28 );
nand NAND2_19042 ( P2_R1146_U377 , P2_U3064 , P2_R1146_U25 );
nand NAND2_19043 ( P2_R1146_U378 , P2_R1146_U377 , P2_R1146_U376 );
nand NAND2_19044 ( P2_R1146_U379 , P2_U3456 , P2_R1146_U26 );
nand NAND2_19045 ( P2_R1146_U380 , P2_U3068 , P2_R1146_U22 );
nand NAND2_19046 ( P2_R1146_U381 , P2_R1146_U241 , P2_R1146_U43 );
nand NAND2_19047 ( P2_R1146_U382 , P2_R1146_U153 , P2_R1146_U196 );
nand NAND2_19048 ( P2_R1146_U383 , P2_U3979 , P2_R1146_U155 );
nand NAND2_19049 ( P2_R1146_U384 , P2_U3055 , P2_R1146_U154 );
nand NAND2_19050 ( P2_R1146_U385 , P2_U3979 , P2_R1146_U155 );
nand NAND2_19051 ( P2_R1146_U386 , P2_U3055 , P2_R1146_U154 );
nand NAND2_19052 ( P2_R1146_U387 , P2_R1146_U386 , P2_R1146_U385 );
nand NAND3_19053 ( P2_R1146_U388 , P2_U3968 , P2_R1146_U10 , P2_R1146_U84 );
nand NAND3_19054 ( P2_R1146_U389 , P2_R1146_U387 , P2_R1146_U83 , P2_U3054 );
nand NAND2_19055 ( P2_R1146_U390 , P2_U3968 , P2_R1146_U84 );
nand NAND2_19056 ( P2_R1146_U391 , P2_U3054 , P2_R1146_U83 );
not NOT1_19057 ( P2_R1146_U392 , P2_R1146_U129 );
nand NAND2_19058 ( P2_R1146_U393 , P2_R1146_U306 , P2_R1146_U392 );
nand NAND2_19059 ( P2_R1146_U394 , P2_R1146_U129 , P2_R1146_U157 );
nand NAND2_19060 ( P2_R1146_U395 , P2_U3969 , P2_R1146_U82 );
nand NAND2_19061 ( P2_R1146_U396 , P2_U3053 , P2_R1146_U79 );
nand NAND2_19062 ( P2_R1146_U397 , P2_U3969 , P2_R1146_U82 );
nand NAND2_19063 ( P2_R1146_U398 , P2_U3053 , P2_R1146_U79 );
nand NAND2_19064 ( P2_R1146_U399 , P2_R1146_U398 , P2_R1146_U397 );
nand NAND2_19065 ( P2_R1146_U400 , P2_U3970 , P2_R1146_U80 );
nand NAND2_19066 ( P2_R1146_U401 , P2_U3057 , P2_R1146_U44 );
nand NAND2_19067 ( P2_R1146_U402 , P2_R1146_U313 , P2_R1146_U85 );
nand NAND2_19068 ( P2_R1146_U403 , P2_R1146_U158 , P2_R1146_U300 );
nand NAND2_19069 ( P2_R1146_U404 , P2_U3971 , P2_R1146_U78 );
nand NAND2_19070 ( P2_R1146_U405 , P2_U3058 , P2_R1146_U77 );
not NOT1_19071 ( P2_R1146_U406 , P2_R1146_U132 );
nand NAND2_19072 ( P2_R1146_U407 , P2_R1146_U296 , P2_R1146_U406 );
nand NAND2_19073 ( P2_R1146_U408 , P2_R1146_U132 , P2_R1146_U159 );
nand NAND2_19074 ( P2_R1146_U409 , P2_U3972 , P2_R1146_U76 );
nand NAND2_19075 ( P2_R1146_U410 , P2_U3065 , P2_R1146_U75 );
not NOT1_19076 ( P2_R1146_U411 , P2_R1146_U133 );
nand NAND2_19077 ( P2_R1146_U412 , P2_R1146_U292 , P2_R1146_U411 );
nand NAND2_19078 ( P2_R1146_U413 , P2_R1146_U133 , P2_R1146_U160 );
nand NAND2_19079 ( P2_R1146_U414 , P2_U3973 , P2_R1146_U71 );
nand NAND2_19080 ( P2_R1146_U415 , P2_U3066 , P2_R1146_U69 );
nand NAND2_19081 ( P2_R1146_U416 , P2_R1146_U415 , P2_R1146_U414 );
nand NAND2_19082 ( P2_R1146_U417 , P2_U3974 , P2_R1146_U72 );
nand NAND2_19083 ( P2_R1146_U418 , P2_U3061 , P2_R1146_U45 );
nand NAND2_19084 ( P2_R1146_U419 , P2_R1146_U323 , P2_R1146_U86 );
nand NAND2_19085 ( P2_R1146_U420 , P2_R1146_U161 , P2_R1146_U315 );
nand NAND2_19086 ( P2_R1146_U421 , P2_U3975 , P2_R1146_U73 );
nand NAND2_19087 ( P2_R1146_U422 , P2_U3075 , P2_R1146_U70 );
nand NAND2_19088 ( P2_R1146_U423 , P2_R1146_U324 , P2_R1146_U163 );
nand NAND2_19089 ( P2_R1146_U424 , P2_R1146_U282 , P2_R1146_U162 );
nand NAND2_19090 ( P2_R1146_U425 , P2_U3976 , P2_R1146_U68 );
nand NAND2_19091 ( P2_R1146_U426 , P2_U3076 , P2_R1146_U67 );
not NOT1_19092 ( P2_R1146_U427 , P2_R1146_U136 );
nand NAND2_19093 ( P2_R1146_U428 , P2_R1146_U278 , P2_R1146_U427 );
nand NAND2_19094 ( P2_R1146_U429 , P2_R1146_U136 , P2_R1146_U164 );
nand NAND2_19095 ( P2_R1146_U430 , P2_U3453 , P2_R1146_U24 );
nand NAND2_19096 ( P2_R1146_U431 , P2_U3078 , P2_R1146_U165 );
not NOT1_19097 ( P2_R1146_U432 , P2_R1146_U137 );
nand NAND2_19098 ( P2_R1146_U433 , P2_R1146_U194 , P2_R1146_U432 );
nand NAND2_19099 ( P2_R1146_U434 , P2_R1146_U137 , P2_R1146_U166 );
nand NAND2_19100 ( P2_R1146_U435 , P2_U3506 , P2_R1146_U66 );
nand NAND2_19101 ( P2_R1146_U436 , P2_U3081 , P2_R1146_U65 );
not NOT1_19102 ( P2_R1146_U437 , P2_R1146_U138 );
nand NAND2_19103 ( P2_R1146_U438 , P2_R1146_U274 , P2_R1146_U437 );
nand NAND2_19104 ( P2_R1146_U439 , P2_R1146_U138 , P2_R1146_U167 );
nand NAND2_19105 ( P2_R1146_U440 , P2_U3504 , P2_R1146_U64 );
nand NAND2_19106 ( P2_R1146_U441 , P2_U3082 , P2_R1146_U168 );
not NOT1_19107 ( P2_R1146_U442 , P2_R1146_U139 );
nand NAND2_19108 ( P2_R1146_U443 , P2_R1146_U272 , P2_R1146_U442 );
nand NAND2_19109 ( P2_R1146_U444 , P2_R1146_U139 , P2_R1146_U169 );
nand NAND2_19110 ( P2_R1146_U445 , P2_U3501 , P2_R1146_U63 );
nand NAND2_19111 ( P2_R1146_U446 , P2_U3069 , P2_R1146_U62 );
not NOT1_19112 ( P2_R1146_U447 , P2_R1146_U140 );
nand NAND2_19113 ( P2_R1146_U448 , P2_R1146_U268 , P2_R1146_U447 );
nand NAND2_19114 ( P2_R1146_U449 , P2_R1146_U140 , P2_R1146_U170 );
nand NAND2_19115 ( P2_R1146_U450 , P2_U3498 , P2_R1146_U58 );
nand NAND2_19116 ( P2_R1146_U451 , P2_U3073 , P2_R1146_U56 );
nand NAND2_19117 ( P2_R1146_U452 , P2_R1146_U451 , P2_R1146_U450 );
nand NAND2_19118 ( P2_R1146_U453 , P2_U3495 , P2_R1146_U59 );
nand NAND2_19119 ( P2_R1146_U454 , P2_U3074 , P2_R1146_U46 );
nand NAND2_19120 ( P2_R1146_U455 , P2_R1146_U334 , P2_R1146_U87 );
nand NAND2_19121 ( P2_R1146_U456 , P2_R1146_U171 , P2_R1146_U326 );
nand NAND2_19122 ( P2_R1146_U457 , P2_U3492 , P2_R1146_U60 );
nand NAND2_19123 ( P2_R1146_U458 , P2_U3079 , P2_R1146_U57 );
nand NAND2_19124 ( P2_R1146_U459 , P2_R1146_U335 , P2_R1146_U173 );
nand NAND2_19125 ( P2_R1146_U460 , P2_R1146_U258 , P2_R1146_U172 );
nand NAND2_19126 ( P2_R1146_U461 , P2_U3489 , P2_R1146_U55 );
nand NAND2_19127 ( P2_R1146_U462 , P2_U3080 , P2_R1146_U54 );
not NOT1_19128 ( P2_R1146_U463 , P2_R1146_U143 );
nand NAND2_19129 ( P2_R1146_U464 , P2_R1146_U254 , P2_R1146_U463 );
nand NAND2_19130 ( P2_R1146_U465 , P2_R1146_U143 , P2_R1146_U174 );
nand NAND2_19131 ( P2_R1146_U466 , P2_U3486 , P2_R1146_U53 );
nand NAND2_19132 ( P2_R1146_U467 , P2_U3072 , P2_R1146_U52 );
not NOT1_19133 ( P2_R1146_U468 , P2_R1146_U144 );
nand NAND2_19134 ( P2_R1146_U469 , P2_R1146_U250 , P2_R1146_U468 );
nand NAND2_19135 ( P2_R1146_U470 , P2_R1146_U144 , P2_R1146_U175 );
nand NAND2_19136 ( P2_R1146_U471 , P2_U3483 , P2_R1146_U49 );
nand NAND2_19137 ( P2_R1146_U472 , P2_U3063 , P2_R1146_U48 );
nand NAND2_19138 ( P2_R1146_U473 , P2_R1146_U472 , P2_R1146_U471 );
nand NAND2_19139 ( P2_R1146_U474 , P2_U3480 , P2_R1146_U50 );
nand NAND2_19140 ( P2_R1146_U475 , P2_U3062 , P2_R1146_U47 );
nand NAND2_19141 ( P2_R1146_U476 , P2_R1146_U345 , P2_R1146_U88 );
nand NAND2_19142 ( P2_R1146_U477 , P2_R1146_U176 , P2_R1146_U337 );
and AND2_19143 ( P2_R1203_U6 , P2_R1203_U205 , P2_R1203_U204 );
and AND2_19144 ( P2_R1203_U7 , P2_R1203_U244 , P2_R1203_U243 );
and AND2_19145 ( P2_R1203_U8 , P2_R1203_U261 , P2_R1203_U260 );
and AND2_19146 ( P2_R1203_U9 , P2_R1203_U285 , P2_R1203_U284 );
and AND2_19147 ( P2_R1203_U10 , P2_R1203_U384 , P2_R1203_U383 );
nand NAND2_19148 ( P2_R1203_U11 , P2_R1203_U340 , P2_R1203_U343 );
nand NAND2_19149 ( P2_R1203_U12 , P2_R1203_U329 , P2_R1203_U332 );
nand NAND2_19150 ( P2_R1203_U13 , P2_R1203_U318 , P2_R1203_U321 );
nand NAND2_19151 ( P2_R1203_U14 , P2_R1203_U310 , P2_R1203_U312 );
nand NAND3_19152 ( P2_R1203_U15 , P2_R1203_U349 , P2_R1203_U177 , P2_R1203_U156 );
nand NAND2_19153 ( P2_R1203_U16 , P2_R1203_U238 , P2_R1203_U240 );
nand NAND2_19154 ( P2_R1203_U17 , P2_R1203_U230 , P2_R1203_U233 );
nand NAND2_19155 ( P2_R1203_U18 , P2_R1203_U222 , P2_R1203_U224 );
nand NAND2_19156 ( P2_R1203_U19 , P2_R1203_U166 , P2_R1203_U346 );
not NOT1_19157 ( P2_R1203_U20 , P2_U3471 );
not NOT1_19158 ( P2_R1203_U21 , P2_U3465 );
not NOT1_19159 ( P2_R1203_U22 , P2_U3456 );
not NOT1_19160 ( P2_R1203_U23 , P2_U3448 );
not NOT1_19161 ( P2_R1203_U24 , P2_U3078 );
not NOT1_19162 ( P2_R1203_U25 , P2_U3459 );
not NOT1_19163 ( P2_R1203_U26 , P2_U3068 );
nand NAND2_19164 ( P2_R1203_U27 , P2_U3068 , P2_R1203_U22 );
not NOT1_19165 ( P2_R1203_U28 , P2_U3064 );
not NOT1_19166 ( P2_R1203_U29 , P2_U3468 );
not NOT1_19167 ( P2_R1203_U30 , P2_U3462 );
not NOT1_19168 ( P2_R1203_U31 , P2_U3071 );
not NOT1_19169 ( P2_R1203_U32 , P2_U3067 );
not NOT1_19170 ( P2_R1203_U33 , P2_U3060 );
nand NAND2_19171 ( P2_R1203_U34 , P2_U3060 , P2_R1203_U30 );
not NOT1_19172 ( P2_R1203_U35 , P2_U3474 );
not NOT1_19173 ( P2_R1203_U36 , P2_U3070 );
nand NAND2_19174 ( P2_R1203_U37 , P2_U3070 , P2_R1203_U20 );
not NOT1_19175 ( P2_R1203_U38 , P2_U3084 );
not NOT1_19176 ( P2_R1203_U39 , P2_U3477 );
not NOT1_19177 ( P2_R1203_U40 , P2_U3083 );
nand NAND2_19178 ( P2_R1203_U41 , P2_R1203_U211 , P2_R1203_U210 );
nand NAND2_19179 ( P2_R1203_U42 , P2_R1203_U34 , P2_R1203_U226 );
nand NAND3_19180 ( P2_R1203_U43 , P2_R1203_U195 , P2_R1203_U179 , P2_R1203_U347 );
not NOT1_19181 ( P2_R1203_U44 , P2_U3970 );
not NOT1_19182 ( P2_R1203_U45 , P2_U3974 );
not NOT1_19183 ( P2_R1203_U46 , P2_U3495 );
not NOT1_19184 ( P2_R1203_U47 , P2_U3480 );
not NOT1_19185 ( P2_R1203_U48 , P2_U3483 );
not NOT1_19186 ( P2_R1203_U49 , P2_U3063 );
not NOT1_19187 ( P2_R1203_U50 , P2_U3062 );
nand NAND2_19188 ( P2_R1203_U51 , P2_U3083 , P2_R1203_U39 );
not NOT1_19189 ( P2_R1203_U52 , P2_U3486 );
not NOT1_19190 ( P2_R1203_U53 , P2_U3072 );
not NOT1_19191 ( P2_R1203_U54 , P2_U3489 );
not NOT1_19192 ( P2_R1203_U55 , P2_U3080 );
not NOT1_19193 ( P2_R1203_U56 , P2_U3498 );
not NOT1_19194 ( P2_R1203_U57 , P2_U3492 );
not NOT1_19195 ( P2_R1203_U58 , P2_U3073 );
not NOT1_19196 ( P2_R1203_U59 , P2_U3074 );
not NOT1_19197 ( P2_R1203_U60 , P2_U3079 );
nand NAND2_19198 ( P2_R1203_U61 , P2_U3079 , P2_R1203_U57 );
not NOT1_19199 ( P2_R1203_U62 , P2_U3501 );
not NOT1_19200 ( P2_R1203_U63 , P2_U3069 );
not NOT1_19201 ( P2_R1203_U64 , P2_U3082 );
not NOT1_19202 ( P2_R1203_U65 , P2_U3506 );
not NOT1_19203 ( P2_R1203_U66 , P2_U3081 );
not NOT1_19204 ( P2_R1203_U67 , P2_U3976 );
not NOT1_19205 ( P2_R1203_U68 , P2_U3076 );
not NOT1_19206 ( P2_R1203_U69 , P2_U3973 );
not NOT1_19207 ( P2_R1203_U70 , P2_U3975 );
not NOT1_19208 ( P2_R1203_U71 , P2_U3066 );
not NOT1_19209 ( P2_R1203_U72 , P2_U3061 );
not NOT1_19210 ( P2_R1203_U73 , P2_U3075 );
nand NAND2_19211 ( P2_R1203_U74 , P2_U3075 , P2_R1203_U70 );
not NOT1_19212 ( P2_R1203_U75 , P2_U3972 );
not NOT1_19213 ( P2_R1203_U76 , P2_U3065 );
not NOT1_19214 ( P2_R1203_U77 , P2_U3971 );
not NOT1_19215 ( P2_R1203_U78 , P2_U3058 );
not NOT1_19216 ( P2_R1203_U79 , P2_U3969 );
not NOT1_19217 ( P2_R1203_U80 , P2_U3057 );
nand NAND2_19218 ( P2_R1203_U81 , P2_U3057 , P2_R1203_U44 );
not NOT1_19219 ( P2_R1203_U82 , P2_U3053 );
not NOT1_19220 ( P2_R1203_U83 , P2_U3968 );
not NOT1_19221 ( P2_R1203_U84 , P2_U3054 );
nand NAND2_19222 ( P2_R1203_U85 , P2_R1203_U299 , P2_R1203_U298 );
nand NAND2_19223 ( P2_R1203_U86 , P2_R1203_U74 , P2_R1203_U314 );
nand NAND2_19224 ( P2_R1203_U87 , P2_R1203_U61 , P2_R1203_U325 );
nand NAND2_19225 ( P2_R1203_U88 , P2_R1203_U51 , P2_R1203_U336 );
not NOT1_19226 ( P2_R1203_U89 , P2_U3077 );
nand NAND2_19227 ( P2_R1203_U90 , P2_R1203_U394 , P2_R1203_U393 );
nand NAND2_19228 ( P2_R1203_U91 , P2_R1203_U408 , P2_R1203_U407 );
nand NAND2_19229 ( P2_R1203_U92 , P2_R1203_U413 , P2_R1203_U412 );
nand NAND2_19230 ( P2_R1203_U93 , P2_R1203_U429 , P2_R1203_U428 );
nand NAND2_19231 ( P2_R1203_U94 , P2_R1203_U434 , P2_R1203_U433 );
nand NAND2_19232 ( P2_R1203_U95 , P2_R1203_U439 , P2_R1203_U438 );
nand NAND2_19233 ( P2_R1203_U96 , P2_R1203_U444 , P2_R1203_U443 );
nand NAND2_19234 ( P2_R1203_U97 , P2_R1203_U449 , P2_R1203_U448 );
nand NAND2_19235 ( P2_R1203_U98 , P2_R1203_U465 , P2_R1203_U464 );
nand NAND2_19236 ( P2_R1203_U99 , P2_R1203_U470 , P2_R1203_U469 );
nand NAND2_19237 ( P2_R1203_U100 , P2_R1203_U353 , P2_R1203_U352 );
nand NAND2_19238 ( P2_R1203_U101 , P2_R1203_U362 , P2_R1203_U361 );
nand NAND2_19239 ( P2_R1203_U102 , P2_R1203_U369 , P2_R1203_U368 );
nand NAND2_19240 ( P2_R1203_U103 , P2_R1203_U373 , P2_R1203_U372 );
nand NAND2_19241 ( P2_R1203_U104 , P2_R1203_U382 , P2_R1203_U381 );
nand NAND2_19242 ( P2_R1203_U105 , P2_R1203_U403 , P2_R1203_U402 );
nand NAND2_19243 ( P2_R1203_U106 , P2_R1203_U420 , P2_R1203_U419 );
nand NAND2_19244 ( P2_R1203_U107 , P2_R1203_U424 , P2_R1203_U423 );
nand NAND2_19245 ( P2_R1203_U108 , P2_R1203_U456 , P2_R1203_U455 );
nand NAND2_19246 ( P2_R1203_U109 , P2_R1203_U460 , P2_R1203_U459 );
nand NAND2_19247 ( P2_R1203_U110 , P2_R1203_U477 , P2_R1203_U476 );
and AND2_19248 ( P2_R1203_U111 , P2_R1203_U197 , P2_R1203_U187 );
and AND2_19249 ( P2_R1203_U112 , P2_R1203_U200 , P2_R1203_U201 );
and AND3_19250 ( P2_R1203_U113 , P2_R1203_U208 , P2_R1203_U203 , P2_R1203_U188 );
and AND2_19251 ( P2_R1203_U114 , P2_R1203_U213 , P2_R1203_U189 );
and AND2_19252 ( P2_R1203_U115 , P2_R1203_U216 , P2_R1203_U217 );
and AND3_19253 ( P2_R1203_U116 , P2_R1203_U355 , P2_R1203_U354 , P2_R1203_U37 );
and AND2_19254 ( P2_R1203_U117 , P2_R1203_U358 , P2_R1203_U189 );
and AND2_19255 ( P2_R1203_U118 , P2_R1203_U232 , P2_R1203_U6 );
and AND2_19256 ( P2_R1203_U119 , P2_R1203_U365 , P2_R1203_U188 );
and AND3_19257 ( P2_R1203_U120 , P2_R1203_U375 , P2_R1203_U374 , P2_R1203_U27 );
and AND2_19258 ( P2_R1203_U121 , P2_R1203_U378 , P2_R1203_U187 );
and AND3_19259 ( P2_R1203_U122 , P2_R1203_U242 , P2_R1203_U219 , P2_R1203_U183 );
and AND3_19260 ( P2_R1203_U123 , P2_R1203_U264 , P2_R1203_U184 , P2_R1203_U259 );
and AND3_19261 ( P2_R1203_U124 , P2_R1203_U288 , P2_R1203_U185 , P2_R1203_U283 );
and AND2_19262 ( P2_R1203_U125 , P2_R1203_U301 , P2_R1203_U186 );
and AND2_19263 ( P2_R1203_U126 , P2_R1203_U304 , P2_R1203_U305 );
and AND2_19264 ( P2_R1203_U127 , P2_R1203_U304 , P2_R1203_U305 );
and AND2_19265 ( P2_R1203_U128 , P2_R1203_U10 , P2_R1203_U308 );
nand NAND2_19266 ( P2_R1203_U129 , P2_R1203_U391 , P2_R1203_U390 );
and AND3_19267 ( P2_R1203_U130 , P2_R1203_U396 , P2_R1203_U395 , P2_R1203_U81 );
and AND2_19268 ( P2_R1203_U131 , P2_R1203_U399 , P2_R1203_U186 );
nand NAND2_19269 ( P2_R1203_U132 , P2_R1203_U405 , P2_R1203_U404 );
nand NAND2_19270 ( P2_R1203_U133 , P2_R1203_U410 , P2_R1203_U409 );
and AND2_19271 ( P2_R1203_U134 , P2_R1203_U320 , P2_R1203_U9 );
and AND2_19272 ( P2_R1203_U135 , P2_R1203_U416 , P2_R1203_U185 );
nand NAND2_19273 ( P2_R1203_U136 , P2_R1203_U426 , P2_R1203_U425 );
nand NAND2_19274 ( P2_R1203_U137 , P2_R1203_U431 , P2_R1203_U430 );
nand NAND2_19275 ( P2_R1203_U138 , P2_R1203_U436 , P2_R1203_U435 );
nand NAND2_19276 ( P2_R1203_U139 , P2_R1203_U441 , P2_R1203_U440 );
nand NAND2_19277 ( P2_R1203_U140 , P2_R1203_U446 , P2_R1203_U445 );
and AND2_19278 ( P2_R1203_U141 , P2_R1203_U331 , P2_R1203_U8 );
and AND2_19279 ( P2_R1203_U142 , P2_R1203_U452 , P2_R1203_U184 );
nand NAND2_19280 ( P2_R1203_U143 , P2_R1203_U462 , P2_R1203_U461 );
nand NAND2_19281 ( P2_R1203_U144 , P2_R1203_U467 , P2_R1203_U466 );
and AND2_19282 ( P2_R1203_U145 , P2_R1203_U342 , P2_R1203_U7 );
and AND2_19283 ( P2_R1203_U146 , P2_R1203_U473 , P2_R1203_U183 );
and AND2_19284 ( P2_R1203_U147 , P2_R1203_U351 , P2_R1203_U350 );
nand NAND2_19285 ( P2_R1203_U148 , P2_R1203_U115 , P2_R1203_U214 );
and AND2_19286 ( P2_R1203_U149 , P2_R1203_U360 , P2_R1203_U359 );
and AND2_19287 ( P2_R1203_U150 , P2_R1203_U367 , P2_R1203_U366 );
and AND2_19288 ( P2_R1203_U151 , P2_R1203_U371 , P2_R1203_U370 );
nand NAND2_19289 ( P2_R1203_U152 , P2_R1203_U112 , P2_R1203_U198 );
and AND2_19290 ( P2_R1203_U153 , P2_R1203_U380 , P2_R1203_U379 );
not NOT1_19291 ( P2_R1203_U154 , P2_U3979 );
not NOT1_19292 ( P2_R1203_U155 , P2_U3055 );
and AND2_19293 ( P2_R1203_U156 , P2_R1203_U389 , P2_R1203_U388 );
nand NAND2_19294 ( P2_R1203_U157 , P2_R1203_U126 , P2_R1203_U302 );
and AND2_19295 ( P2_R1203_U158 , P2_R1203_U401 , P2_R1203_U400 );
nand NAND2_19296 ( P2_R1203_U159 , P2_R1203_U295 , P2_R1203_U294 );
nand NAND2_19297 ( P2_R1203_U160 , P2_R1203_U291 , P2_R1203_U290 );
and AND2_19298 ( P2_R1203_U161 , P2_R1203_U418 , P2_R1203_U417 );
and AND2_19299 ( P2_R1203_U162 , P2_R1203_U422 , P2_R1203_U421 );
nand NAND2_19300 ( P2_R1203_U163 , P2_R1203_U281 , P2_R1203_U280 );
nand NAND2_19301 ( P2_R1203_U164 , P2_R1203_U277 , P2_R1203_U276 );
not NOT1_19302 ( P2_R1203_U165 , P2_U3453 );
nand NAND2_19303 ( P2_R1203_U166 , P2_U3448 , P2_R1203_U89 );
nand NAND3_19304 ( P2_R1203_U167 , P2_R1203_U273 , P2_R1203_U178 , P2_R1203_U348 );
not NOT1_19305 ( P2_R1203_U168 , P2_U3504 );
nand NAND2_19306 ( P2_R1203_U169 , P2_R1203_U271 , P2_R1203_U270 );
nand NAND2_19307 ( P2_R1203_U170 , P2_R1203_U267 , P2_R1203_U266 );
and AND2_19308 ( P2_R1203_U171 , P2_R1203_U454 , P2_R1203_U453 );
and AND2_19309 ( P2_R1203_U172 , P2_R1203_U458 , P2_R1203_U457 );
nand NAND2_19310 ( P2_R1203_U173 , P2_R1203_U257 , P2_R1203_U256 );
nand NAND2_19311 ( P2_R1203_U174 , P2_R1203_U253 , P2_R1203_U252 );
nand NAND2_19312 ( P2_R1203_U175 , P2_R1203_U249 , P2_R1203_U248 );
and AND2_19313 ( P2_R1203_U176 , P2_R1203_U475 , P2_R1203_U474 );
nand NAND3_19314 ( P2_R1203_U177 , P2_R1203_U307 , P2_R1203_U157 , P2_R1203_U387 );
nand NAND2_19315 ( P2_R1203_U178 , P2_R1203_U169 , P2_R1203_U168 );
nand NAND2_19316 ( P2_R1203_U179 , P2_R1203_U166 , P2_R1203_U165 );
not NOT1_19317 ( P2_R1203_U180 , P2_R1203_U81 );
not NOT1_19318 ( P2_R1203_U181 , P2_R1203_U27 );
not NOT1_19319 ( P2_R1203_U182 , P2_R1203_U37 );
nand NAND2_19320 ( P2_R1203_U183 , P2_U3480 , P2_R1203_U50 );
nand NAND2_19321 ( P2_R1203_U184 , P2_U3495 , P2_R1203_U59 );
nand NAND2_19322 ( P2_R1203_U185 , P2_U3974 , P2_R1203_U72 );
nand NAND2_19323 ( P2_R1203_U186 , P2_U3970 , P2_R1203_U80 );
nand NAND2_19324 ( P2_R1203_U187 , P2_U3456 , P2_R1203_U26 );
nand NAND2_19325 ( P2_R1203_U188 , P2_U3465 , P2_R1203_U32 );
nand NAND2_19326 ( P2_R1203_U189 , P2_U3471 , P2_R1203_U36 );
not NOT1_19327 ( P2_R1203_U190 , P2_R1203_U61 );
not NOT1_19328 ( P2_R1203_U191 , P2_R1203_U74 );
not NOT1_19329 ( P2_R1203_U192 , P2_R1203_U34 );
not NOT1_19330 ( P2_R1203_U193 , P2_R1203_U51 );
not NOT1_19331 ( P2_R1203_U194 , P2_R1203_U166 );
nand NAND2_19332 ( P2_R1203_U195 , P2_U3078 , P2_R1203_U166 );
not NOT1_19333 ( P2_R1203_U196 , P2_R1203_U43 );
nand NAND2_19334 ( P2_R1203_U197 , P2_U3459 , P2_R1203_U28 );
nand NAND2_19335 ( P2_R1203_U198 , P2_R1203_U111 , P2_R1203_U43 );
nand NAND2_19336 ( P2_R1203_U199 , P2_R1203_U28 , P2_R1203_U27 );
nand NAND2_19337 ( P2_R1203_U200 , P2_R1203_U199 , P2_R1203_U25 );
nand NAND2_19338 ( P2_R1203_U201 , P2_U3064 , P2_R1203_U181 );
not NOT1_19339 ( P2_R1203_U202 , P2_R1203_U152 );
nand NAND2_19340 ( P2_R1203_U203 , P2_U3468 , P2_R1203_U31 );
nand NAND2_19341 ( P2_R1203_U204 , P2_U3071 , P2_R1203_U29 );
nand NAND2_19342 ( P2_R1203_U205 , P2_U3067 , P2_R1203_U21 );
nand NAND2_19343 ( P2_R1203_U206 , P2_R1203_U192 , P2_R1203_U188 );
nand NAND2_19344 ( P2_R1203_U207 , P2_R1203_U6 , P2_R1203_U206 );
nand NAND2_19345 ( P2_R1203_U208 , P2_U3462 , P2_R1203_U33 );
nand NAND2_19346 ( P2_R1203_U209 , P2_U3468 , P2_R1203_U31 );
nand NAND2_19347 ( P2_R1203_U210 , P2_R1203_U152 , P2_R1203_U113 );
nand NAND2_19348 ( P2_R1203_U211 , P2_R1203_U209 , P2_R1203_U207 );
not NOT1_19349 ( P2_R1203_U212 , P2_R1203_U41 );
nand NAND2_19350 ( P2_R1203_U213 , P2_U3474 , P2_R1203_U38 );
nand NAND2_19351 ( P2_R1203_U214 , P2_R1203_U114 , P2_R1203_U41 );
nand NAND2_19352 ( P2_R1203_U215 , P2_R1203_U38 , P2_R1203_U37 );
nand NAND2_19353 ( P2_R1203_U216 , P2_R1203_U215 , P2_R1203_U35 );
nand NAND2_19354 ( P2_R1203_U217 , P2_U3084 , P2_R1203_U182 );
not NOT1_19355 ( P2_R1203_U218 , P2_R1203_U148 );
nand NAND2_19356 ( P2_R1203_U219 , P2_U3477 , P2_R1203_U40 );
nand NAND2_19357 ( P2_R1203_U220 , P2_R1203_U219 , P2_R1203_U51 );
nand NAND2_19358 ( P2_R1203_U221 , P2_R1203_U212 , P2_R1203_U37 );
nand NAND2_19359 ( P2_R1203_U222 , P2_R1203_U117 , P2_R1203_U221 );
nand NAND2_19360 ( P2_R1203_U223 , P2_R1203_U41 , P2_R1203_U189 );
nand NAND2_19361 ( P2_R1203_U224 , P2_R1203_U116 , P2_R1203_U223 );
nand NAND2_19362 ( P2_R1203_U225 , P2_R1203_U37 , P2_R1203_U189 );
nand NAND2_19363 ( P2_R1203_U226 , P2_R1203_U208 , P2_R1203_U152 );
not NOT1_19364 ( P2_R1203_U227 , P2_R1203_U42 );
nand NAND2_19365 ( P2_R1203_U228 , P2_U3067 , P2_R1203_U21 );
nand NAND2_19366 ( P2_R1203_U229 , P2_R1203_U227 , P2_R1203_U228 );
nand NAND2_19367 ( P2_R1203_U230 , P2_R1203_U119 , P2_R1203_U229 );
nand NAND2_19368 ( P2_R1203_U231 , P2_R1203_U42 , P2_R1203_U188 );
nand NAND2_19369 ( P2_R1203_U232 , P2_U3468 , P2_R1203_U31 );
nand NAND2_19370 ( P2_R1203_U233 , P2_R1203_U118 , P2_R1203_U231 );
nand NAND2_19371 ( P2_R1203_U234 , P2_U3067 , P2_R1203_U21 );
nand NAND2_19372 ( P2_R1203_U235 , P2_R1203_U188 , P2_R1203_U234 );
nand NAND2_19373 ( P2_R1203_U236 , P2_R1203_U208 , P2_R1203_U34 );
nand NAND2_19374 ( P2_R1203_U237 , P2_R1203_U196 , P2_R1203_U27 );
nand NAND2_19375 ( P2_R1203_U238 , P2_R1203_U121 , P2_R1203_U237 );
nand NAND2_19376 ( P2_R1203_U239 , P2_R1203_U43 , P2_R1203_U187 );
nand NAND2_19377 ( P2_R1203_U240 , P2_R1203_U120 , P2_R1203_U239 );
nand NAND2_19378 ( P2_R1203_U241 , P2_R1203_U27 , P2_R1203_U187 );
nand NAND2_19379 ( P2_R1203_U242 , P2_U3483 , P2_R1203_U49 );
nand NAND2_19380 ( P2_R1203_U243 , P2_U3063 , P2_R1203_U48 );
nand NAND2_19381 ( P2_R1203_U244 , P2_U3062 , P2_R1203_U47 );
nand NAND2_19382 ( P2_R1203_U245 , P2_R1203_U193 , P2_R1203_U183 );
nand NAND2_19383 ( P2_R1203_U246 , P2_R1203_U7 , P2_R1203_U245 );
nand NAND2_19384 ( P2_R1203_U247 , P2_U3483 , P2_R1203_U49 );
nand NAND2_19385 ( P2_R1203_U248 , P2_R1203_U148 , P2_R1203_U122 );
nand NAND2_19386 ( P2_R1203_U249 , P2_R1203_U247 , P2_R1203_U246 );
not NOT1_19387 ( P2_R1203_U250 , P2_R1203_U175 );
nand NAND2_19388 ( P2_R1203_U251 , P2_U3486 , P2_R1203_U53 );
nand NAND2_19389 ( P2_R1203_U252 , P2_R1203_U251 , P2_R1203_U175 );
nand NAND2_19390 ( P2_R1203_U253 , P2_U3072 , P2_R1203_U52 );
not NOT1_19391 ( P2_R1203_U254 , P2_R1203_U174 );
nand NAND2_19392 ( P2_R1203_U255 , P2_U3489 , P2_R1203_U55 );
nand NAND2_19393 ( P2_R1203_U256 , P2_R1203_U255 , P2_R1203_U174 );
nand NAND2_19394 ( P2_R1203_U257 , P2_U3080 , P2_R1203_U54 );
not NOT1_19395 ( P2_R1203_U258 , P2_R1203_U173 );
nand NAND2_19396 ( P2_R1203_U259 , P2_U3498 , P2_R1203_U58 );
nand NAND2_19397 ( P2_R1203_U260 , P2_U3073 , P2_R1203_U56 );
nand NAND2_19398 ( P2_R1203_U261 , P2_U3074 , P2_R1203_U46 );
nand NAND2_19399 ( P2_R1203_U262 , P2_R1203_U190 , P2_R1203_U184 );
nand NAND2_19400 ( P2_R1203_U263 , P2_R1203_U8 , P2_R1203_U262 );
nand NAND2_19401 ( P2_R1203_U264 , P2_U3492 , P2_R1203_U60 );
nand NAND2_19402 ( P2_R1203_U265 , P2_U3498 , P2_R1203_U58 );
nand NAND2_19403 ( P2_R1203_U266 , P2_R1203_U173 , P2_R1203_U123 );
nand NAND2_19404 ( P2_R1203_U267 , P2_R1203_U265 , P2_R1203_U263 );
not NOT1_19405 ( P2_R1203_U268 , P2_R1203_U170 );
nand NAND2_19406 ( P2_R1203_U269 , P2_U3501 , P2_R1203_U63 );
nand NAND2_19407 ( P2_R1203_U270 , P2_R1203_U269 , P2_R1203_U170 );
nand NAND2_19408 ( P2_R1203_U271 , P2_U3069 , P2_R1203_U62 );
not NOT1_19409 ( P2_R1203_U272 , P2_R1203_U169 );
nand NAND2_19410 ( P2_R1203_U273 , P2_U3082 , P2_R1203_U169 );
not NOT1_19411 ( P2_R1203_U274 , P2_R1203_U167 );
nand NAND2_19412 ( P2_R1203_U275 , P2_U3506 , P2_R1203_U66 );
nand NAND2_19413 ( P2_R1203_U276 , P2_R1203_U275 , P2_R1203_U167 );
nand NAND2_19414 ( P2_R1203_U277 , P2_U3081 , P2_R1203_U65 );
not NOT1_19415 ( P2_R1203_U278 , P2_R1203_U164 );
nand NAND2_19416 ( P2_R1203_U279 , P2_U3976 , P2_R1203_U68 );
nand NAND2_19417 ( P2_R1203_U280 , P2_R1203_U279 , P2_R1203_U164 );
nand NAND2_19418 ( P2_R1203_U281 , P2_U3076 , P2_R1203_U67 );
not NOT1_19419 ( P2_R1203_U282 , P2_R1203_U163 );
nand NAND2_19420 ( P2_R1203_U283 , P2_U3973 , P2_R1203_U71 );
nand NAND2_19421 ( P2_R1203_U284 , P2_U3066 , P2_R1203_U69 );
nand NAND2_19422 ( P2_R1203_U285 , P2_U3061 , P2_R1203_U45 );
nand NAND2_19423 ( P2_R1203_U286 , P2_R1203_U191 , P2_R1203_U185 );
nand NAND2_19424 ( P2_R1203_U287 , P2_R1203_U9 , P2_R1203_U286 );
nand NAND2_19425 ( P2_R1203_U288 , P2_U3975 , P2_R1203_U73 );
nand NAND2_19426 ( P2_R1203_U289 , P2_U3973 , P2_R1203_U71 );
nand NAND2_19427 ( P2_R1203_U290 , P2_R1203_U163 , P2_R1203_U124 );
nand NAND2_19428 ( P2_R1203_U291 , P2_R1203_U289 , P2_R1203_U287 );
not NOT1_19429 ( P2_R1203_U292 , P2_R1203_U160 );
nand NAND2_19430 ( P2_R1203_U293 , P2_U3972 , P2_R1203_U76 );
nand NAND2_19431 ( P2_R1203_U294 , P2_R1203_U293 , P2_R1203_U160 );
nand NAND2_19432 ( P2_R1203_U295 , P2_U3065 , P2_R1203_U75 );
not NOT1_19433 ( P2_R1203_U296 , P2_R1203_U159 );
nand NAND2_19434 ( P2_R1203_U297 , P2_U3971 , P2_R1203_U78 );
nand NAND2_19435 ( P2_R1203_U298 , P2_R1203_U297 , P2_R1203_U159 );
nand NAND2_19436 ( P2_R1203_U299 , P2_U3058 , P2_R1203_U77 );
not NOT1_19437 ( P2_R1203_U300 , P2_R1203_U85 );
nand NAND2_19438 ( P2_R1203_U301 , P2_U3969 , P2_R1203_U82 );
nand NAND2_19439 ( P2_R1203_U302 , P2_R1203_U125 , P2_R1203_U85 );
nand NAND2_19440 ( P2_R1203_U303 , P2_R1203_U82 , P2_R1203_U81 );
nand NAND2_19441 ( P2_R1203_U304 , P2_R1203_U303 , P2_R1203_U79 );
nand NAND2_19442 ( P2_R1203_U305 , P2_U3053 , P2_R1203_U180 );
not NOT1_19443 ( P2_R1203_U306 , P2_R1203_U157 );
nand NAND2_19444 ( P2_R1203_U307 , P2_U3968 , P2_R1203_U84 );
nand NAND2_19445 ( P2_R1203_U308 , P2_U3054 , P2_R1203_U83 );
nand NAND2_19446 ( P2_R1203_U309 , P2_R1203_U300 , P2_R1203_U81 );
nand NAND2_19447 ( P2_R1203_U310 , P2_R1203_U131 , P2_R1203_U309 );
nand NAND2_19448 ( P2_R1203_U311 , P2_R1203_U85 , P2_R1203_U186 );
nand NAND2_19449 ( P2_R1203_U312 , P2_R1203_U130 , P2_R1203_U311 );
nand NAND2_19450 ( P2_R1203_U313 , P2_R1203_U81 , P2_R1203_U186 );
nand NAND2_19451 ( P2_R1203_U314 , P2_R1203_U288 , P2_R1203_U163 );
not NOT1_19452 ( P2_R1203_U315 , P2_R1203_U86 );
nand NAND2_19453 ( P2_R1203_U316 , P2_U3061 , P2_R1203_U45 );
nand NAND2_19454 ( P2_R1203_U317 , P2_R1203_U315 , P2_R1203_U316 );
nand NAND2_19455 ( P2_R1203_U318 , P2_R1203_U135 , P2_R1203_U317 );
nand NAND2_19456 ( P2_R1203_U319 , P2_R1203_U86 , P2_R1203_U185 );
nand NAND2_19457 ( P2_R1203_U320 , P2_U3973 , P2_R1203_U71 );
nand NAND2_19458 ( P2_R1203_U321 , P2_R1203_U134 , P2_R1203_U319 );
nand NAND2_19459 ( P2_R1203_U322 , P2_U3061 , P2_R1203_U45 );
nand NAND2_19460 ( P2_R1203_U323 , P2_R1203_U185 , P2_R1203_U322 );
nand NAND2_19461 ( P2_R1203_U324 , P2_R1203_U288 , P2_R1203_U74 );
nand NAND2_19462 ( P2_R1203_U325 , P2_R1203_U264 , P2_R1203_U173 );
not NOT1_19463 ( P2_R1203_U326 , P2_R1203_U87 );
nand NAND2_19464 ( P2_R1203_U327 , P2_U3074 , P2_R1203_U46 );
nand NAND2_19465 ( P2_R1203_U328 , P2_R1203_U326 , P2_R1203_U327 );
nand NAND2_19466 ( P2_R1203_U329 , P2_R1203_U142 , P2_R1203_U328 );
nand NAND2_19467 ( P2_R1203_U330 , P2_R1203_U87 , P2_R1203_U184 );
nand NAND2_19468 ( P2_R1203_U331 , P2_U3498 , P2_R1203_U58 );
nand NAND2_19469 ( P2_R1203_U332 , P2_R1203_U141 , P2_R1203_U330 );
nand NAND2_19470 ( P2_R1203_U333 , P2_U3074 , P2_R1203_U46 );
nand NAND2_19471 ( P2_R1203_U334 , P2_R1203_U184 , P2_R1203_U333 );
nand NAND2_19472 ( P2_R1203_U335 , P2_R1203_U264 , P2_R1203_U61 );
nand NAND2_19473 ( P2_R1203_U336 , P2_R1203_U219 , P2_R1203_U148 );
not NOT1_19474 ( P2_R1203_U337 , P2_R1203_U88 );
nand NAND2_19475 ( P2_R1203_U338 , P2_U3062 , P2_R1203_U47 );
nand NAND2_19476 ( P2_R1203_U339 , P2_R1203_U337 , P2_R1203_U338 );
nand NAND2_19477 ( P2_R1203_U340 , P2_R1203_U146 , P2_R1203_U339 );
nand NAND2_19478 ( P2_R1203_U341 , P2_R1203_U88 , P2_R1203_U183 );
nand NAND2_19479 ( P2_R1203_U342 , P2_U3483 , P2_R1203_U49 );
nand NAND2_19480 ( P2_R1203_U343 , P2_R1203_U145 , P2_R1203_U341 );
nand NAND2_19481 ( P2_R1203_U344 , P2_U3062 , P2_R1203_U47 );
nand NAND2_19482 ( P2_R1203_U345 , P2_R1203_U183 , P2_R1203_U344 );
nand NAND2_19483 ( P2_R1203_U346 , P2_U3077 , P2_R1203_U23 );
nand NAND2_19484 ( P2_R1203_U347 , P2_U3078 , P2_R1203_U165 );
nand NAND2_19485 ( P2_R1203_U348 , P2_U3082 , P2_R1203_U168 );
nand NAND3_19486 ( P2_R1203_U349 , P2_R1203_U127 , P2_R1203_U302 , P2_R1203_U128 );
nand NAND2_19487 ( P2_R1203_U350 , P2_U3477 , P2_R1203_U40 );
nand NAND2_19488 ( P2_R1203_U351 , P2_U3083 , P2_R1203_U39 );
nand NAND2_19489 ( P2_R1203_U352 , P2_R1203_U220 , P2_R1203_U148 );
nand NAND2_19490 ( P2_R1203_U353 , P2_R1203_U218 , P2_R1203_U147 );
nand NAND2_19491 ( P2_R1203_U354 , P2_U3474 , P2_R1203_U38 );
nand NAND2_19492 ( P2_R1203_U355 , P2_U3084 , P2_R1203_U35 );
nand NAND2_19493 ( P2_R1203_U356 , P2_U3474 , P2_R1203_U38 );
nand NAND2_19494 ( P2_R1203_U357 , P2_U3084 , P2_R1203_U35 );
nand NAND2_19495 ( P2_R1203_U358 , P2_R1203_U357 , P2_R1203_U356 );
nand NAND2_19496 ( P2_R1203_U359 , P2_U3471 , P2_R1203_U36 );
nand NAND2_19497 ( P2_R1203_U360 , P2_U3070 , P2_R1203_U20 );
nand NAND2_19498 ( P2_R1203_U361 , P2_R1203_U225 , P2_R1203_U41 );
nand NAND2_19499 ( P2_R1203_U362 , P2_R1203_U149 , P2_R1203_U212 );
nand NAND2_19500 ( P2_R1203_U363 , P2_U3468 , P2_R1203_U31 );
nand NAND2_19501 ( P2_R1203_U364 , P2_U3071 , P2_R1203_U29 );
nand NAND2_19502 ( P2_R1203_U365 , P2_R1203_U364 , P2_R1203_U363 );
nand NAND2_19503 ( P2_R1203_U366 , P2_U3465 , P2_R1203_U32 );
nand NAND2_19504 ( P2_R1203_U367 , P2_U3067 , P2_R1203_U21 );
nand NAND2_19505 ( P2_R1203_U368 , P2_R1203_U235 , P2_R1203_U42 );
nand NAND2_19506 ( P2_R1203_U369 , P2_R1203_U150 , P2_R1203_U227 );
nand NAND2_19507 ( P2_R1203_U370 , P2_U3462 , P2_R1203_U33 );
nand NAND2_19508 ( P2_R1203_U371 , P2_U3060 , P2_R1203_U30 );
nand NAND2_19509 ( P2_R1203_U372 , P2_R1203_U236 , P2_R1203_U152 );
nand NAND2_19510 ( P2_R1203_U373 , P2_R1203_U202 , P2_R1203_U151 );
nand NAND2_19511 ( P2_R1203_U374 , P2_U3459 , P2_R1203_U28 );
nand NAND2_19512 ( P2_R1203_U375 , P2_U3064 , P2_R1203_U25 );
nand NAND2_19513 ( P2_R1203_U376 , P2_U3459 , P2_R1203_U28 );
nand NAND2_19514 ( P2_R1203_U377 , P2_U3064 , P2_R1203_U25 );
nand NAND2_19515 ( P2_R1203_U378 , P2_R1203_U377 , P2_R1203_U376 );
nand NAND2_19516 ( P2_R1203_U379 , P2_U3456 , P2_R1203_U26 );
nand NAND2_19517 ( P2_R1203_U380 , P2_U3068 , P2_R1203_U22 );
nand NAND2_19518 ( P2_R1203_U381 , P2_R1203_U241 , P2_R1203_U43 );
nand NAND2_19519 ( P2_R1203_U382 , P2_R1203_U153 , P2_R1203_U196 );
nand NAND2_19520 ( P2_R1203_U383 , P2_U3979 , P2_R1203_U155 );
nand NAND2_19521 ( P2_R1203_U384 , P2_U3055 , P2_R1203_U154 );
nand NAND2_19522 ( P2_R1203_U385 , P2_U3979 , P2_R1203_U155 );
nand NAND2_19523 ( P2_R1203_U386 , P2_U3055 , P2_R1203_U154 );
nand NAND2_19524 ( P2_R1203_U387 , P2_R1203_U386 , P2_R1203_U385 );
nand NAND3_19525 ( P2_R1203_U388 , P2_U3968 , P2_R1203_U10 , P2_R1203_U84 );
nand NAND3_19526 ( P2_R1203_U389 , P2_R1203_U387 , P2_R1203_U83 , P2_U3054 );
nand NAND2_19527 ( P2_R1203_U390 , P2_U3968 , P2_R1203_U84 );
nand NAND2_19528 ( P2_R1203_U391 , P2_U3054 , P2_R1203_U83 );
not NOT1_19529 ( P2_R1203_U392 , P2_R1203_U129 );
nand NAND2_19530 ( P2_R1203_U393 , P2_R1203_U306 , P2_R1203_U392 );
nand NAND2_19531 ( P2_R1203_U394 , P2_R1203_U129 , P2_R1203_U157 );
nand NAND2_19532 ( P2_R1203_U395 , P2_U3969 , P2_R1203_U82 );
nand NAND2_19533 ( P2_R1203_U396 , P2_U3053 , P2_R1203_U79 );
nand NAND2_19534 ( P2_R1203_U397 , P2_U3969 , P2_R1203_U82 );
nand NAND2_19535 ( P2_R1203_U398 , P2_U3053 , P2_R1203_U79 );
nand NAND2_19536 ( P2_R1203_U399 , P2_R1203_U398 , P2_R1203_U397 );
nand NAND2_19537 ( P2_R1203_U400 , P2_U3970 , P2_R1203_U80 );
nand NAND2_19538 ( P2_R1203_U401 , P2_U3057 , P2_R1203_U44 );
nand NAND2_19539 ( P2_R1203_U402 , P2_R1203_U313 , P2_R1203_U85 );
nand NAND2_19540 ( P2_R1203_U403 , P2_R1203_U158 , P2_R1203_U300 );
nand NAND2_19541 ( P2_R1203_U404 , P2_U3971 , P2_R1203_U78 );
nand NAND2_19542 ( P2_R1203_U405 , P2_U3058 , P2_R1203_U77 );
not NOT1_19543 ( P2_R1203_U406 , P2_R1203_U132 );
nand NAND2_19544 ( P2_R1203_U407 , P2_R1203_U296 , P2_R1203_U406 );
nand NAND2_19545 ( P2_R1203_U408 , P2_R1203_U132 , P2_R1203_U159 );
nand NAND2_19546 ( P2_R1203_U409 , P2_U3972 , P2_R1203_U76 );
nand NAND2_19547 ( P2_R1203_U410 , P2_U3065 , P2_R1203_U75 );
not NOT1_19548 ( P2_R1203_U411 , P2_R1203_U133 );
nand NAND2_19549 ( P2_R1203_U412 , P2_R1203_U292 , P2_R1203_U411 );
nand NAND2_19550 ( P2_R1203_U413 , P2_R1203_U133 , P2_R1203_U160 );
nand NAND2_19551 ( P2_R1203_U414 , P2_U3973 , P2_R1203_U71 );
nand NAND2_19552 ( P2_R1203_U415 , P2_U3066 , P2_R1203_U69 );
nand NAND2_19553 ( P2_R1203_U416 , P2_R1203_U415 , P2_R1203_U414 );
nand NAND2_19554 ( P2_R1203_U417 , P2_U3974 , P2_R1203_U72 );
nand NAND2_19555 ( P2_R1203_U418 , P2_U3061 , P2_R1203_U45 );
nand NAND2_19556 ( P2_R1203_U419 , P2_R1203_U323 , P2_R1203_U86 );
nand NAND2_19557 ( P2_R1203_U420 , P2_R1203_U161 , P2_R1203_U315 );
nand NAND2_19558 ( P2_R1203_U421 , P2_U3975 , P2_R1203_U73 );
nand NAND2_19559 ( P2_R1203_U422 , P2_U3075 , P2_R1203_U70 );
nand NAND2_19560 ( P2_R1203_U423 , P2_R1203_U324 , P2_R1203_U163 );
nand NAND2_19561 ( P2_R1203_U424 , P2_R1203_U282 , P2_R1203_U162 );
nand NAND2_19562 ( P2_R1203_U425 , P2_U3976 , P2_R1203_U68 );
nand NAND2_19563 ( P2_R1203_U426 , P2_U3076 , P2_R1203_U67 );
not NOT1_19564 ( P2_R1203_U427 , P2_R1203_U136 );
nand NAND2_19565 ( P2_R1203_U428 , P2_R1203_U278 , P2_R1203_U427 );
nand NAND2_19566 ( P2_R1203_U429 , P2_R1203_U136 , P2_R1203_U164 );
nand NAND2_19567 ( P2_R1203_U430 , P2_U3453 , P2_R1203_U24 );
nand NAND2_19568 ( P2_R1203_U431 , P2_U3078 , P2_R1203_U165 );
not NOT1_19569 ( P2_R1203_U432 , P2_R1203_U137 );
nand NAND2_19570 ( P2_R1203_U433 , P2_R1203_U194 , P2_R1203_U432 );
nand NAND2_19571 ( P2_R1203_U434 , P2_R1203_U137 , P2_R1203_U166 );
nand NAND2_19572 ( P2_R1203_U435 , P2_U3506 , P2_R1203_U66 );
nand NAND2_19573 ( P2_R1203_U436 , P2_U3081 , P2_R1203_U65 );
not NOT1_19574 ( P2_R1203_U437 , P2_R1203_U138 );
nand NAND2_19575 ( P2_R1203_U438 , P2_R1203_U274 , P2_R1203_U437 );
nand NAND2_19576 ( P2_R1203_U439 , P2_R1203_U138 , P2_R1203_U167 );
nand NAND2_19577 ( P2_R1203_U440 , P2_U3504 , P2_R1203_U64 );
nand NAND2_19578 ( P2_R1203_U441 , P2_U3082 , P2_R1203_U168 );
not NOT1_19579 ( P2_R1203_U442 , P2_R1203_U139 );
nand NAND2_19580 ( P2_R1203_U443 , P2_R1203_U272 , P2_R1203_U442 );
nand NAND2_19581 ( P2_R1203_U444 , P2_R1203_U139 , P2_R1203_U169 );
nand NAND2_19582 ( P2_R1203_U445 , P2_U3501 , P2_R1203_U63 );
nand NAND2_19583 ( P2_R1203_U446 , P2_U3069 , P2_R1203_U62 );
not NOT1_19584 ( P2_R1203_U447 , P2_R1203_U140 );
nand NAND2_19585 ( P2_R1203_U448 , P2_R1203_U268 , P2_R1203_U447 );
nand NAND2_19586 ( P2_R1203_U449 , P2_R1203_U140 , P2_R1203_U170 );
nand NAND2_19587 ( P2_R1203_U450 , P2_U3498 , P2_R1203_U58 );
nand NAND2_19588 ( P2_R1203_U451 , P2_U3073 , P2_R1203_U56 );
nand NAND2_19589 ( P2_R1203_U452 , P2_R1203_U451 , P2_R1203_U450 );
nand NAND2_19590 ( P2_R1203_U453 , P2_U3495 , P2_R1203_U59 );
nand NAND2_19591 ( P2_R1203_U454 , P2_U3074 , P2_R1203_U46 );
nand NAND2_19592 ( P2_R1203_U455 , P2_R1203_U334 , P2_R1203_U87 );
nand NAND2_19593 ( P2_R1203_U456 , P2_R1203_U171 , P2_R1203_U326 );
nand NAND2_19594 ( P2_R1203_U457 , P2_U3492 , P2_R1203_U60 );
nand NAND2_19595 ( P2_R1203_U458 , P2_U3079 , P2_R1203_U57 );
nand NAND2_19596 ( P2_R1203_U459 , P2_R1203_U335 , P2_R1203_U173 );
nand NAND2_19597 ( P2_R1203_U460 , P2_R1203_U258 , P2_R1203_U172 );
nand NAND2_19598 ( P2_R1203_U461 , P2_U3489 , P2_R1203_U55 );
nand NAND2_19599 ( P2_R1203_U462 , P2_U3080 , P2_R1203_U54 );
not NOT1_19600 ( P2_R1203_U463 , P2_R1203_U143 );
nand NAND2_19601 ( P2_R1203_U464 , P2_R1203_U254 , P2_R1203_U463 );
nand NAND2_19602 ( P2_R1203_U465 , P2_R1203_U143 , P2_R1203_U174 );
nand NAND2_19603 ( P2_R1203_U466 , P2_U3486 , P2_R1203_U53 );
nand NAND2_19604 ( P2_R1203_U467 , P2_U3072 , P2_R1203_U52 );
not NOT1_19605 ( P2_R1203_U468 , P2_R1203_U144 );
nand NAND2_19606 ( P2_R1203_U469 , P2_R1203_U250 , P2_R1203_U468 );
nand NAND2_19607 ( P2_R1203_U470 , P2_R1203_U144 , P2_R1203_U175 );
nand NAND2_19608 ( P2_R1203_U471 , P2_U3483 , P2_R1203_U49 );
nand NAND2_19609 ( P2_R1203_U472 , P2_U3063 , P2_R1203_U48 );
nand NAND2_19610 ( P2_R1203_U473 , P2_R1203_U472 , P2_R1203_U471 );
nand NAND2_19611 ( P2_R1203_U474 , P2_U3480 , P2_R1203_U50 );
nand NAND2_19612 ( P2_R1203_U475 , P2_U3062 , P2_R1203_U47 );
nand NAND2_19613 ( P2_R1203_U476 , P2_R1203_U345 , P2_R1203_U88 );
nand NAND2_19614 ( P2_R1203_U477 , P2_R1203_U176 , P2_R1203_U337 );
and AND2_19615 ( P2_R1113_U6 , P2_R1113_U205 , P2_R1113_U204 );
and AND2_19616 ( P2_R1113_U7 , P2_R1113_U244 , P2_R1113_U243 );
and AND2_19617 ( P2_R1113_U8 , P2_R1113_U261 , P2_R1113_U260 );
and AND2_19618 ( P2_R1113_U9 , P2_R1113_U285 , P2_R1113_U284 );
and AND2_19619 ( P2_R1113_U10 , P2_R1113_U384 , P2_R1113_U383 );
nand NAND2_19620 ( P2_R1113_U11 , P2_R1113_U340 , P2_R1113_U343 );
nand NAND2_19621 ( P2_R1113_U12 , P2_R1113_U329 , P2_R1113_U332 );
nand NAND2_19622 ( P2_R1113_U13 , P2_R1113_U318 , P2_R1113_U321 );
nand NAND2_19623 ( P2_R1113_U14 , P2_R1113_U310 , P2_R1113_U312 );
nand NAND3_19624 ( P2_R1113_U15 , P2_R1113_U349 , P2_R1113_U177 , P2_R1113_U156 );
nand NAND2_19625 ( P2_R1113_U16 , P2_R1113_U238 , P2_R1113_U240 );
nand NAND2_19626 ( P2_R1113_U17 , P2_R1113_U230 , P2_R1113_U233 );
nand NAND2_19627 ( P2_R1113_U18 , P2_R1113_U222 , P2_R1113_U224 );
nand NAND2_19628 ( P2_R1113_U19 , P2_R1113_U166 , P2_R1113_U346 );
not NOT1_19629 ( P2_R1113_U20 , P2_U3471 );
not NOT1_19630 ( P2_R1113_U21 , P2_U3465 );
not NOT1_19631 ( P2_R1113_U22 , P2_U3456 );
not NOT1_19632 ( P2_R1113_U23 , P2_U3448 );
not NOT1_19633 ( P2_R1113_U24 , P2_U3078 );
not NOT1_19634 ( P2_R1113_U25 , P2_U3459 );
not NOT1_19635 ( P2_R1113_U26 , P2_U3068 );
nand NAND2_19636 ( P2_R1113_U27 , P2_U3068 , P2_R1113_U22 );
not NOT1_19637 ( P2_R1113_U28 , P2_U3064 );
not NOT1_19638 ( P2_R1113_U29 , P2_U3468 );
not NOT1_19639 ( P2_R1113_U30 , P2_U3462 );
not NOT1_19640 ( P2_R1113_U31 , P2_U3071 );
not NOT1_19641 ( P2_R1113_U32 , P2_U3067 );
not NOT1_19642 ( P2_R1113_U33 , P2_U3060 );
nand NAND2_19643 ( P2_R1113_U34 , P2_U3060 , P2_R1113_U30 );
not NOT1_19644 ( P2_R1113_U35 , P2_U3474 );
not NOT1_19645 ( P2_R1113_U36 , P2_U3070 );
nand NAND2_19646 ( P2_R1113_U37 , P2_U3070 , P2_R1113_U20 );
not NOT1_19647 ( P2_R1113_U38 , P2_U3084 );
not NOT1_19648 ( P2_R1113_U39 , P2_U3477 );
not NOT1_19649 ( P2_R1113_U40 , P2_U3083 );
nand NAND2_19650 ( P2_R1113_U41 , P2_R1113_U211 , P2_R1113_U210 );
nand NAND2_19651 ( P2_R1113_U42 , P2_R1113_U34 , P2_R1113_U226 );
nand NAND3_19652 ( P2_R1113_U43 , P2_R1113_U195 , P2_R1113_U179 , P2_R1113_U347 );
not NOT1_19653 ( P2_R1113_U44 , P2_U3970 );
not NOT1_19654 ( P2_R1113_U45 , P2_U3974 );
not NOT1_19655 ( P2_R1113_U46 , P2_U3495 );
not NOT1_19656 ( P2_R1113_U47 , P2_U3480 );
not NOT1_19657 ( P2_R1113_U48 , P2_U3483 );
not NOT1_19658 ( P2_R1113_U49 , P2_U3063 );
not NOT1_19659 ( P2_R1113_U50 , P2_U3062 );
nand NAND2_19660 ( P2_R1113_U51 , P2_U3083 , P2_R1113_U39 );
not NOT1_19661 ( P2_R1113_U52 , P2_U3486 );
not NOT1_19662 ( P2_R1113_U53 , P2_U3072 );
not NOT1_19663 ( P2_R1113_U54 , P2_U3489 );
not NOT1_19664 ( P2_R1113_U55 , P2_U3080 );
not NOT1_19665 ( P2_R1113_U56 , P2_U3498 );
not NOT1_19666 ( P2_R1113_U57 , P2_U3492 );
not NOT1_19667 ( P2_R1113_U58 , P2_U3073 );
not NOT1_19668 ( P2_R1113_U59 , P2_U3074 );
not NOT1_19669 ( P2_R1113_U60 , P2_U3079 );
nand NAND2_19670 ( P2_R1113_U61 , P2_U3079 , P2_R1113_U57 );
not NOT1_19671 ( P2_R1113_U62 , P2_U3501 );
not NOT1_19672 ( P2_R1113_U63 , P2_U3069 );
not NOT1_19673 ( P2_R1113_U64 , P2_U3082 );
not NOT1_19674 ( P2_R1113_U65 , P2_U3506 );
not NOT1_19675 ( P2_R1113_U66 , P2_U3081 );
not NOT1_19676 ( P2_R1113_U67 , P2_U3976 );
not NOT1_19677 ( P2_R1113_U68 , P2_U3076 );
not NOT1_19678 ( P2_R1113_U69 , P2_U3973 );
not NOT1_19679 ( P2_R1113_U70 , P2_U3975 );
not NOT1_19680 ( P2_R1113_U71 , P2_U3066 );
not NOT1_19681 ( P2_R1113_U72 , P2_U3061 );
not NOT1_19682 ( P2_R1113_U73 , P2_U3075 );
nand NAND2_19683 ( P2_R1113_U74 , P2_U3075 , P2_R1113_U70 );
not NOT1_19684 ( P2_R1113_U75 , P2_U3972 );
not NOT1_19685 ( P2_R1113_U76 , P2_U3065 );
not NOT1_19686 ( P2_R1113_U77 , P2_U3971 );
not NOT1_19687 ( P2_R1113_U78 , P2_U3058 );
not NOT1_19688 ( P2_R1113_U79 , P2_U3969 );
not NOT1_19689 ( P2_R1113_U80 , P2_U3057 );
nand NAND2_19690 ( P2_R1113_U81 , P2_U3057 , P2_R1113_U44 );
not NOT1_19691 ( P2_R1113_U82 , P2_U3053 );
not NOT1_19692 ( P2_R1113_U83 , P2_U3968 );
not NOT1_19693 ( P2_R1113_U84 , P2_U3054 );
nand NAND2_19694 ( P2_R1113_U85 , P2_R1113_U299 , P2_R1113_U298 );
nand NAND2_19695 ( P2_R1113_U86 , P2_R1113_U74 , P2_R1113_U314 );
nand NAND2_19696 ( P2_R1113_U87 , P2_R1113_U61 , P2_R1113_U325 );
nand NAND2_19697 ( P2_R1113_U88 , P2_R1113_U51 , P2_R1113_U336 );
not NOT1_19698 ( P2_R1113_U89 , P2_U3077 );
nand NAND2_19699 ( P2_R1113_U90 , P2_R1113_U394 , P2_R1113_U393 );
nand NAND2_19700 ( P2_R1113_U91 , P2_R1113_U408 , P2_R1113_U407 );
nand NAND2_19701 ( P2_R1113_U92 , P2_R1113_U413 , P2_R1113_U412 );
nand NAND2_19702 ( P2_R1113_U93 , P2_R1113_U429 , P2_R1113_U428 );
nand NAND2_19703 ( P2_R1113_U94 , P2_R1113_U434 , P2_R1113_U433 );
nand NAND2_19704 ( P2_R1113_U95 , P2_R1113_U439 , P2_R1113_U438 );
nand NAND2_19705 ( P2_R1113_U96 , P2_R1113_U444 , P2_R1113_U443 );
nand NAND2_19706 ( P2_R1113_U97 , P2_R1113_U449 , P2_R1113_U448 );
nand NAND2_19707 ( P2_R1113_U98 , P2_R1113_U465 , P2_R1113_U464 );
nand NAND2_19708 ( P2_R1113_U99 , P2_R1113_U470 , P2_R1113_U469 );
nand NAND2_19709 ( P2_R1113_U100 , P2_R1113_U353 , P2_R1113_U352 );
nand NAND2_19710 ( P2_R1113_U101 , P2_R1113_U362 , P2_R1113_U361 );
nand NAND2_19711 ( P2_R1113_U102 , P2_R1113_U369 , P2_R1113_U368 );
nand NAND2_19712 ( P2_R1113_U103 , P2_R1113_U373 , P2_R1113_U372 );
nand NAND2_19713 ( P2_R1113_U104 , P2_R1113_U382 , P2_R1113_U381 );
nand NAND2_19714 ( P2_R1113_U105 , P2_R1113_U403 , P2_R1113_U402 );
nand NAND2_19715 ( P2_R1113_U106 , P2_R1113_U420 , P2_R1113_U419 );
nand NAND2_19716 ( P2_R1113_U107 , P2_R1113_U424 , P2_R1113_U423 );
nand NAND2_19717 ( P2_R1113_U108 , P2_R1113_U456 , P2_R1113_U455 );
nand NAND2_19718 ( P2_R1113_U109 , P2_R1113_U460 , P2_R1113_U459 );
nand NAND2_19719 ( P2_R1113_U110 , P2_R1113_U477 , P2_R1113_U476 );
and AND2_19720 ( P2_R1113_U111 , P2_R1113_U197 , P2_R1113_U187 );
and AND2_19721 ( P2_R1113_U112 , P2_R1113_U200 , P2_R1113_U201 );
and AND3_19722 ( P2_R1113_U113 , P2_R1113_U208 , P2_R1113_U203 , P2_R1113_U188 );
and AND2_19723 ( P2_R1113_U114 , P2_R1113_U213 , P2_R1113_U189 );
and AND2_19724 ( P2_R1113_U115 , P2_R1113_U216 , P2_R1113_U217 );
and AND3_19725 ( P2_R1113_U116 , P2_R1113_U355 , P2_R1113_U354 , P2_R1113_U37 );
and AND2_19726 ( P2_R1113_U117 , P2_R1113_U358 , P2_R1113_U189 );
and AND2_19727 ( P2_R1113_U118 , P2_R1113_U232 , P2_R1113_U6 );
and AND2_19728 ( P2_R1113_U119 , P2_R1113_U365 , P2_R1113_U188 );
and AND3_19729 ( P2_R1113_U120 , P2_R1113_U375 , P2_R1113_U374 , P2_R1113_U27 );
and AND2_19730 ( P2_R1113_U121 , P2_R1113_U378 , P2_R1113_U187 );
and AND3_19731 ( P2_R1113_U122 , P2_R1113_U242 , P2_R1113_U219 , P2_R1113_U183 );
and AND3_19732 ( P2_R1113_U123 , P2_R1113_U264 , P2_R1113_U184 , P2_R1113_U259 );
and AND3_19733 ( P2_R1113_U124 , P2_R1113_U288 , P2_R1113_U185 , P2_R1113_U283 );
and AND2_19734 ( P2_R1113_U125 , P2_R1113_U301 , P2_R1113_U186 );
and AND2_19735 ( P2_R1113_U126 , P2_R1113_U304 , P2_R1113_U305 );
and AND2_19736 ( P2_R1113_U127 , P2_R1113_U304 , P2_R1113_U305 );
and AND2_19737 ( P2_R1113_U128 , P2_R1113_U10 , P2_R1113_U308 );
nand NAND2_19738 ( P2_R1113_U129 , P2_R1113_U391 , P2_R1113_U390 );
and AND3_19739 ( P2_R1113_U130 , P2_R1113_U396 , P2_R1113_U395 , P2_R1113_U81 );
and AND2_19740 ( P2_R1113_U131 , P2_R1113_U399 , P2_R1113_U186 );
nand NAND2_19741 ( P2_R1113_U132 , P2_R1113_U405 , P2_R1113_U404 );
nand NAND2_19742 ( P2_R1113_U133 , P2_R1113_U410 , P2_R1113_U409 );
and AND2_19743 ( P2_R1113_U134 , P2_R1113_U320 , P2_R1113_U9 );
and AND2_19744 ( P2_R1113_U135 , P2_R1113_U416 , P2_R1113_U185 );
nand NAND2_19745 ( P2_R1113_U136 , P2_R1113_U426 , P2_R1113_U425 );
nand NAND2_19746 ( P2_R1113_U137 , P2_R1113_U431 , P2_R1113_U430 );
nand NAND2_19747 ( P2_R1113_U138 , P2_R1113_U436 , P2_R1113_U435 );
nand NAND2_19748 ( P2_R1113_U139 , P2_R1113_U441 , P2_R1113_U440 );
nand NAND2_19749 ( P2_R1113_U140 , P2_R1113_U446 , P2_R1113_U445 );
and AND2_19750 ( P2_R1113_U141 , P2_R1113_U331 , P2_R1113_U8 );
and AND2_19751 ( P2_R1113_U142 , P2_R1113_U452 , P2_R1113_U184 );
nand NAND2_19752 ( P2_R1113_U143 , P2_R1113_U462 , P2_R1113_U461 );
nand NAND2_19753 ( P2_R1113_U144 , P2_R1113_U467 , P2_R1113_U466 );
and AND2_19754 ( P2_R1113_U145 , P2_R1113_U342 , P2_R1113_U7 );
and AND2_19755 ( P2_R1113_U146 , P2_R1113_U473 , P2_R1113_U183 );
and AND2_19756 ( P2_R1113_U147 , P2_R1113_U351 , P2_R1113_U350 );
nand NAND2_19757 ( P2_R1113_U148 , P2_R1113_U115 , P2_R1113_U214 );
and AND2_19758 ( P2_R1113_U149 , P2_R1113_U360 , P2_R1113_U359 );
and AND2_19759 ( P2_R1113_U150 , P2_R1113_U367 , P2_R1113_U366 );
and AND2_19760 ( P2_R1113_U151 , P2_R1113_U371 , P2_R1113_U370 );
nand NAND2_19761 ( P2_R1113_U152 , P2_R1113_U112 , P2_R1113_U198 );
and AND2_19762 ( P2_R1113_U153 , P2_R1113_U380 , P2_R1113_U379 );
not NOT1_19763 ( P2_R1113_U154 , P2_U3979 );
not NOT1_19764 ( P2_R1113_U155 , P2_U3055 );
and AND2_19765 ( P2_R1113_U156 , P2_R1113_U389 , P2_R1113_U388 );
nand NAND2_19766 ( P2_R1113_U157 , P2_R1113_U126 , P2_R1113_U302 );
and AND2_19767 ( P2_R1113_U158 , P2_R1113_U401 , P2_R1113_U400 );
nand NAND2_19768 ( P2_R1113_U159 , P2_R1113_U295 , P2_R1113_U294 );
nand NAND2_19769 ( P2_R1113_U160 , P2_R1113_U291 , P2_R1113_U290 );
and AND2_19770 ( P2_R1113_U161 , P2_R1113_U418 , P2_R1113_U417 );
and AND2_19771 ( P2_R1113_U162 , P2_R1113_U422 , P2_R1113_U421 );
nand NAND2_19772 ( P2_R1113_U163 , P2_R1113_U281 , P2_R1113_U280 );
nand NAND2_19773 ( P2_R1113_U164 , P2_R1113_U277 , P2_R1113_U276 );
not NOT1_19774 ( P2_R1113_U165 , P2_U3453 );
nand NAND2_19775 ( P2_R1113_U166 , P2_U3448 , P2_R1113_U89 );
nand NAND3_19776 ( P2_R1113_U167 , P2_R1113_U273 , P2_R1113_U178 , P2_R1113_U348 );
not NOT1_19777 ( P2_R1113_U168 , P2_U3504 );
nand NAND2_19778 ( P2_R1113_U169 , P2_R1113_U271 , P2_R1113_U270 );
nand NAND2_19779 ( P2_R1113_U170 , P2_R1113_U267 , P2_R1113_U266 );
and AND2_19780 ( P2_R1113_U171 , P2_R1113_U454 , P2_R1113_U453 );
and AND2_19781 ( P2_R1113_U172 , P2_R1113_U458 , P2_R1113_U457 );
nand NAND2_19782 ( P2_R1113_U173 , P2_R1113_U257 , P2_R1113_U256 );
nand NAND2_19783 ( P2_R1113_U174 , P2_R1113_U253 , P2_R1113_U252 );
nand NAND2_19784 ( P2_R1113_U175 , P2_R1113_U249 , P2_R1113_U248 );
and AND2_19785 ( P2_R1113_U176 , P2_R1113_U475 , P2_R1113_U474 );
nand NAND3_19786 ( P2_R1113_U177 , P2_R1113_U307 , P2_R1113_U157 , P2_R1113_U387 );
nand NAND2_19787 ( P2_R1113_U178 , P2_R1113_U169 , P2_R1113_U168 );
nand NAND2_19788 ( P2_R1113_U179 , P2_R1113_U166 , P2_R1113_U165 );
not NOT1_19789 ( P2_R1113_U180 , P2_R1113_U81 );
not NOT1_19790 ( P2_R1113_U181 , P2_R1113_U27 );
not NOT1_19791 ( P2_R1113_U182 , P2_R1113_U37 );
nand NAND2_19792 ( P2_R1113_U183 , P2_U3480 , P2_R1113_U50 );
nand NAND2_19793 ( P2_R1113_U184 , P2_U3495 , P2_R1113_U59 );
nand NAND2_19794 ( P2_R1113_U185 , P2_U3974 , P2_R1113_U72 );
nand NAND2_19795 ( P2_R1113_U186 , P2_U3970 , P2_R1113_U80 );
nand NAND2_19796 ( P2_R1113_U187 , P2_U3456 , P2_R1113_U26 );
nand NAND2_19797 ( P2_R1113_U188 , P2_U3465 , P2_R1113_U32 );
nand NAND2_19798 ( P2_R1113_U189 , P2_U3471 , P2_R1113_U36 );
not NOT1_19799 ( P2_R1113_U190 , P2_R1113_U61 );
not NOT1_19800 ( P2_R1113_U191 , P2_R1113_U74 );
not NOT1_19801 ( P2_R1113_U192 , P2_R1113_U34 );
not NOT1_19802 ( P2_R1113_U193 , P2_R1113_U51 );
not NOT1_19803 ( P2_R1113_U194 , P2_R1113_U166 );
nand NAND2_19804 ( P2_R1113_U195 , P2_U3078 , P2_R1113_U166 );
not NOT1_19805 ( P2_R1113_U196 , P2_R1113_U43 );
nand NAND2_19806 ( P2_R1113_U197 , P2_U3459 , P2_R1113_U28 );
nand NAND2_19807 ( P2_R1113_U198 , P2_R1113_U111 , P2_R1113_U43 );
nand NAND2_19808 ( P2_R1113_U199 , P2_R1113_U28 , P2_R1113_U27 );
nand NAND2_19809 ( P2_R1113_U200 , P2_R1113_U199 , P2_R1113_U25 );
nand NAND2_19810 ( P2_R1113_U201 , P2_U3064 , P2_R1113_U181 );
not NOT1_19811 ( P2_R1113_U202 , P2_R1113_U152 );
nand NAND2_19812 ( P2_R1113_U203 , P2_U3468 , P2_R1113_U31 );
nand NAND2_19813 ( P2_R1113_U204 , P2_U3071 , P2_R1113_U29 );
nand NAND2_19814 ( P2_R1113_U205 , P2_U3067 , P2_R1113_U21 );
nand NAND2_19815 ( P2_R1113_U206 , P2_R1113_U192 , P2_R1113_U188 );
nand NAND2_19816 ( P2_R1113_U207 , P2_R1113_U6 , P2_R1113_U206 );
nand NAND2_19817 ( P2_R1113_U208 , P2_U3462 , P2_R1113_U33 );
nand NAND2_19818 ( P2_R1113_U209 , P2_U3468 , P2_R1113_U31 );
nand NAND2_19819 ( P2_R1113_U210 , P2_R1113_U152 , P2_R1113_U113 );
nand NAND2_19820 ( P2_R1113_U211 , P2_R1113_U209 , P2_R1113_U207 );
not NOT1_19821 ( P2_R1113_U212 , P2_R1113_U41 );
nand NAND2_19822 ( P2_R1113_U213 , P2_U3474 , P2_R1113_U38 );
nand NAND2_19823 ( P2_R1113_U214 , P2_R1113_U114 , P2_R1113_U41 );
nand NAND2_19824 ( P2_R1113_U215 , P2_R1113_U38 , P2_R1113_U37 );
nand NAND2_19825 ( P2_R1113_U216 , P2_R1113_U215 , P2_R1113_U35 );
nand NAND2_19826 ( P2_R1113_U217 , P2_U3084 , P2_R1113_U182 );
not NOT1_19827 ( P2_R1113_U218 , P2_R1113_U148 );
nand NAND2_19828 ( P2_R1113_U219 , P2_U3477 , P2_R1113_U40 );
nand NAND2_19829 ( P2_R1113_U220 , P2_R1113_U219 , P2_R1113_U51 );
nand NAND2_19830 ( P2_R1113_U221 , P2_R1113_U212 , P2_R1113_U37 );
nand NAND2_19831 ( P2_R1113_U222 , P2_R1113_U117 , P2_R1113_U221 );
nand NAND2_19832 ( P2_R1113_U223 , P2_R1113_U41 , P2_R1113_U189 );
nand NAND2_19833 ( P2_R1113_U224 , P2_R1113_U116 , P2_R1113_U223 );
nand NAND2_19834 ( P2_R1113_U225 , P2_R1113_U37 , P2_R1113_U189 );
nand NAND2_19835 ( P2_R1113_U226 , P2_R1113_U208 , P2_R1113_U152 );
not NOT1_19836 ( P2_R1113_U227 , P2_R1113_U42 );
nand NAND2_19837 ( P2_R1113_U228 , P2_U3067 , P2_R1113_U21 );
nand NAND2_19838 ( P2_R1113_U229 , P2_R1113_U227 , P2_R1113_U228 );
nand NAND2_19839 ( P2_R1113_U230 , P2_R1113_U119 , P2_R1113_U229 );
nand NAND2_19840 ( P2_R1113_U231 , P2_R1113_U42 , P2_R1113_U188 );
nand NAND2_19841 ( P2_R1113_U232 , P2_U3468 , P2_R1113_U31 );
nand NAND2_19842 ( P2_R1113_U233 , P2_R1113_U118 , P2_R1113_U231 );
nand NAND2_19843 ( P2_R1113_U234 , P2_U3067 , P2_R1113_U21 );
nand NAND2_19844 ( P2_R1113_U235 , P2_R1113_U188 , P2_R1113_U234 );
nand NAND2_19845 ( P2_R1113_U236 , P2_R1113_U208 , P2_R1113_U34 );
nand NAND2_19846 ( P2_R1113_U237 , P2_R1113_U196 , P2_R1113_U27 );
nand NAND2_19847 ( P2_R1113_U238 , P2_R1113_U121 , P2_R1113_U237 );
nand NAND2_19848 ( P2_R1113_U239 , P2_R1113_U43 , P2_R1113_U187 );
nand NAND2_19849 ( P2_R1113_U240 , P2_R1113_U120 , P2_R1113_U239 );
nand NAND2_19850 ( P2_R1113_U241 , P2_R1113_U27 , P2_R1113_U187 );
nand NAND2_19851 ( P2_R1113_U242 , P2_U3483 , P2_R1113_U49 );
nand NAND2_19852 ( P2_R1113_U243 , P2_U3063 , P2_R1113_U48 );
nand NAND2_19853 ( P2_R1113_U244 , P2_U3062 , P2_R1113_U47 );
nand NAND2_19854 ( P2_R1113_U245 , P2_R1113_U193 , P2_R1113_U183 );
nand NAND2_19855 ( P2_R1113_U246 , P2_R1113_U7 , P2_R1113_U245 );
nand NAND2_19856 ( P2_R1113_U247 , P2_U3483 , P2_R1113_U49 );
nand NAND2_19857 ( P2_R1113_U248 , P2_R1113_U148 , P2_R1113_U122 );
nand NAND2_19858 ( P2_R1113_U249 , P2_R1113_U247 , P2_R1113_U246 );
not NOT1_19859 ( P2_R1113_U250 , P2_R1113_U175 );
nand NAND2_19860 ( P2_R1113_U251 , P2_U3486 , P2_R1113_U53 );
nand NAND2_19861 ( P2_R1113_U252 , P2_R1113_U251 , P2_R1113_U175 );
nand NAND2_19862 ( P2_R1113_U253 , P2_U3072 , P2_R1113_U52 );
not NOT1_19863 ( P2_R1113_U254 , P2_R1113_U174 );
nand NAND2_19864 ( P2_R1113_U255 , P2_U3489 , P2_R1113_U55 );
nand NAND2_19865 ( P2_R1113_U256 , P2_R1113_U255 , P2_R1113_U174 );
nand NAND2_19866 ( P2_R1113_U257 , P2_U3080 , P2_R1113_U54 );
not NOT1_19867 ( P2_R1113_U258 , P2_R1113_U173 );
nand NAND2_19868 ( P2_R1113_U259 , P2_U3498 , P2_R1113_U58 );
nand NAND2_19869 ( P2_R1113_U260 , P2_U3073 , P2_R1113_U56 );
nand NAND2_19870 ( P2_R1113_U261 , P2_U3074 , P2_R1113_U46 );
nand NAND2_19871 ( P2_R1113_U262 , P2_R1113_U190 , P2_R1113_U184 );
nand NAND2_19872 ( P2_R1113_U263 , P2_R1113_U8 , P2_R1113_U262 );
nand NAND2_19873 ( P2_R1113_U264 , P2_U3492 , P2_R1113_U60 );
nand NAND2_19874 ( P2_R1113_U265 , P2_U3498 , P2_R1113_U58 );
nand NAND2_19875 ( P2_R1113_U266 , P2_R1113_U173 , P2_R1113_U123 );
nand NAND2_19876 ( P2_R1113_U267 , P2_R1113_U265 , P2_R1113_U263 );
not NOT1_19877 ( P2_R1113_U268 , P2_R1113_U170 );
nand NAND2_19878 ( P2_R1113_U269 , P2_U3501 , P2_R1113_U63 );
nand NAND2_19879 ( P2_R1113_U270 , P2_R1113_U269 , P2_R1113_U170 );
nand NAND2_19880 ( P2_R1113_U271 , P2_U3069 , P2_R1113_U62 );
not NOT1_19881 ( P2_R1113_U272 , P2_R1113_U169 );
nand NAND2_19882 ( P2_R1113_U273 , P2_U3082 , P2_R1113_U169 );
not NOT1_19883 ( P2_R1113_U274 , P2_R1113_U167 );
nand NAND2_19884 ( P2_R1113_U275 , P2_U3506 , P2_R1113_U66 );
nand NAND2_19885 ( P2_R1113_U276 , P2_R1113_U275 , P2_R1113_U167 );
nand NAND2_19886 ( P2_R1113_U277 , P2_U3081 , P2_R1113_U65 );
not NOT1_19887 ( P2_R1113_U278 , P2_R1113_U164 );
nand NAND2_19888 ( P2_R1113_U279 , P2_U3976 , P2_R1113_U68 );
nand NAND2_19889 ( P2_R1113_U280 , P2_R1113_U279 , P2_R1113_U164 );
nand NAND2_19890 ( P2_R1113_U281 , P2_U3076 , P2_R1113_U67 );
not NOT1_19891 ( P2_R1113_U282 , P2_R1113_U163 );
nand NAND2_19892 ( P2_R1113_U283 , P2_U3973 , P2_R1113_U71 );
nand NAND2_19893 ( P2_R1113_U284 , P2_U3066 , P2_R1113_U69 );
nand NAND2_19894 ( P2_R1113_U285 , P2_U3061 , P2_R1113_U45 );
nand NAND2_19895 ( P2_R1113_U286 , P2_R1113_U191 , P2_R1113_U185 );
nand NAND2_19896 ( P2_R1113_U287 , P2_R1113_U9 , P2_R1113_U286 );
nand NAND2_19897 ( P2_R1113_U288 , P2_U3975 , P2_R1113_U73 );
nand NAND2_19898 ( P2_R1113_U289 , P2_U3973 , P2_R1113_U71 );
nand NAND2_19899 ( P2_R1113_U290 , P2_R1113_U163 , P2_R1113_U124 );
nand NAND2_19900 ( P2_R1113_U291 , P2_R1113_U289 , P2_R1113_U287 );
not NOT1_19901 ( P2_R1113_U292 , P2_R1113_U160 );
nand NAND2_19902 ( P2_R1113_U293 , P2_U3972 , P2_R1113_U76 );
nand NAND2_19903 ( P2_R1113_U294 , P2_R1113_U293 , P2_R1113_U160 );
nand NAND2_19904 ( P2_R1113_U295 , P2_U3065 , P2_R1113_U75 );
not NOT1_19905 ( P2_R1113_U296 , P2_R1113_U159 );
nand NAND2_19906 ( P2_R1113_U297 , P2_U3971 , P2_R1113_U78 );
nand NAND2_19907 ( P2_R1113_U298 , P2_R1113_U297 , P2_R1113_U159 );
nand NAND2_19908 ( P2_R1113_U299 , P2_U3058 , P2_R1113_U77 );
not NOT1_19909 ( P2_R1113_U300 , P2_R1113_U85 );
nand NAND2_19910 ( P2_R1113_U301 , P2_U3969 , P2_R1113_U82 );
nand NAND2_19911 ( P2_R1113_U302 , P2_R1113_U125 , P2_R1113_U85 );
nand NAND2_19912 ( P2_R1113_U303 , P2_R1113_U82 , P2_R1113_U81 );
nand NAND2_19913 ( P2_R1113_U304 , P2_R1113_U303 , P2_R1113_U79 );
nand NAND2_19914 ( P2_R1113_U305 , P2_U3053 , P2_R1113_U180 );
not NOT1_19915 ( P2_R1113_U306 , P2_R1113_U157 );
nand NAND2_19916 ( P2_R1113_U307 , P2_U3968 , P2_R1113_U84 );
nand NAND2_19917 ( P2_R1113_U308 , P2_U3054 , P2_R1113_U83 );
nand NAND2_19918 ( P2_R1113_U309 , P2_R1113_U300 , P2_R1113_U81 );
nand NAND2_19919 ( P2_R1113_U310 , P2_R1113_U131 , P2_R1113_U309 );
nand NAND2_19920 ( P2_R1113_U311 , P2_R1113_U85 , P2_R1113_U186 );
nand NAND2_19921 ( P2_R1113_U312 , P2_R1113_U130 , P2_R1113_U311 );
nand NAND2_19922 ( P2_R1113_U313 , P2_R1113_U81 , P2_R1113_U186 );
nand NAND2_19923 ( P2_R1113_U314 , P2_R1113_U288 , P2_R1113_U163 );
not NOT1_19924 ( P2_R1113_U315 , P2_R1113_U86 );
nand NAND2_19925 ( P2_R1113_U316 , P2_U3061 , P2_R1113_U45 );
nand NAND2_19926 ( P2_R1113_U317 , P2_R1113_U315 , P2_R1113_U316 );
nand NAND2_19927 ( P2_R1113_U318 , P2_R1113_U135 , P2_R1113_U317 );
nand NAND2_19928 ( P2_R1113_U319 , P2_R1113_U86 , P2_R1113_U185 );
nand NAND2_19929 ( P2_R1113_U320 , P2_U3973 , P2_R1113_U71 );
nand NAND2_19930 ( P2_R1113_U321 , P2_R1113_U134 , P2_R1113_U319 );
nand NAND2_19931 ( P2_R1113_U322 , P2_U3061 , P2_R1113_U45 );
nand NAND2_19932 ( P2_R1113_U323 , P2_R1113_U185 , P2_R1113_U322 );
nand NAND2_19933 ( P2_R1113_U324 , P2_R1113_U288 , P2_R1113_U74 );
nand NAND2_19934 ( P2_R1113_U325 , P2_R1113_U264 , P2_R1113_U173 );
not NOT1_19935 ( P2_R1113_U326 , P2_R1113_U87 );
nand NAND2_19936 ( P2_R1113_U327 , P2_U3074 , P2_R1113_U46 );
nand NAND2_19937 ( P2_R1113_U328 , P2_R1113_U326 , P2_R1113_U327 );
nand NAND2_19938 ( P2_R1113_U329 , P2_R1113_U142 , P2_R1113_U328 );
nand NAND2_19939 ( P2_R1113_U330 , P2_R1113_U87 , P2_R1113_U184 );
nand NAND2_19940 ( P2_R1113_U331 , P2_U3498 , P2_R1113_U58 );
nand NAND2_19941 ( P2_R1113_U332 , P2_R1113_U141 , P2_R1113_U330 );
nand NAND2_19942 ( P2_R1113_U333 , P2_U3074 , P2_R1113_U46 );
nand NAND2_19943 ( P2_R1113_U334 , P2_R1113_U184 , P2_R1113_U333 );
nand NAND2_19944 ( P2_R1113_U335 , P2_R1113_U264 , P2_R1113_U61 );
nand NAND2_19945 ( P2_R1113_U336 , P2_R1113_U219 , P2_R1113_U148 );
not NOT1_19946 ( P2_R1113_U337 , P2_R1113_U88 );
nand NAND2_19947 ( P2_R1113_U338 , P2_U3062 , P2_R1113_U47 );
nand NAND2_19948 ( P2_R1113_U339 , P2_R1113_U337 , P2_R1113_U338 );
nand NAND2_19949 ( P2_R1113_U340 , P2_R1113_U146 , P2_R1113_U339 );
nand NAND2_19950 ( P2_R1113_U341 , P2_R1113_U88 , P2_R1113_U183 );
nand NAND2_19951 ( P2_R1113_U342 , P2_U3483 , P2_R1113_U49 );
nand NAND2_19952 ( P2_R1113_U343 , P2_R1113_U145 , P2_R1113_U341 );
nand NAND2_19953 ( P2_R1113_U344 , P2_U3062 , P2_R1113_U47 );
nand NAND2_19954 ( P2_R1113_U345 , P2_R1113_U183 , P2_R1113_U344 );
nand NAND2_19955 ( P2_R1113_U346 , P2_U3077 , P2_R1113_U23 );
nand NAND2_19956 ( P2_R1113_U347 , P2_U3078 , P2_R1113_U165 );
nand NAND2_19957 ( P2_R1113_U348 , P2_U3082 , P2_R1113_U168 );
nand NAND3_19958 ( P2_R1113_U349 , P2_R1113_U127 , P2_R1113_U302 , P2_R1113_U128 );
nand NAND2_19959 ( P2_R1113_U350 , P2_U3477 , P2_R1113_U40 );
nand NAND2_19960 ( P2_R1113_U351 , P2_U3083 , P2_R1113_U39 );
nand NAND2_19961 ( P2_R1113_U352 , P2_R1113_U220 , P2_R1113_U148 );
nand NAND2_19962 ( P2_R1113_U353 , P2_R1113_U218 , P2_R1113_U147 );
nand NAND2_19963 ( P2_R1113_U354 , P2_U3474 , P2_R1113_U38 );
nand NAND2_19964 ( P2_R1113_U355 , P2_U3084 , P2_R1113_U35 );
nand NAND2_19965 ( P2_R1113_U356 , P2_U3474 , P2_R1113_U38 );
nand NAND2_19966 ( P2_R1113_U357 , P2_U3084 , P2_R1113_U35 );
nand NAND2_19967 ( P2_R1113_U358 , P2_R1113_U357 , P2_R1113_U356 );
nand NAND2_19968 ( P2_R1113_U359 , P2_U3471 , P2_R1113_U36 );
nand NAND2_19969 ( P2_R1113_U360 , P2_U3070 , P2_R1113_U20 );
nand NAND2_19970 ( P2_R1113_U361 , P2_R1113_U225 , P2_R1113_U41 );
nand NAND2_19971 ( P2_R1113_U362 , P2_R1113_U149 , P2_R1113_U212 );
nand NAND2_19972 ( P2_R1113_U363 , P2_U3468 , P2_R1113_U31 );
nand NAND2_19973 ( P2_R1113_U364 , P2_U3071 , P2_R1113_U29 );
nand NAND2_19974 ( P2_R1113_U365 , P2_R1113_U364 , P2_R1113_U363 );
nand NAND2_19975 ( P2_R1113_U366 , P2_U3465 , P2_R1113_U32 );
nand NAND2_19976 ( P2_R1113_U367 , P2_U3067 , P2_R1113_U21 );
nand NAND2_19977 ( P2_R1113_U368 , P2_R1113_U235 , P2_R1113_U42 );
nand NAND2_19978 ( P2_R1113_U369 , P2_R1113_U150 , P2_R1113_U227 );
nand NAND2_19979 ( P2_R1113_U370 , P2_U3462 , P2_R1113_U33 );
nand NAND2_19980 ( P2_R1113_U371 , P2_U3060 , P2_R1113_U30 );
nand NAND2_19981 ( P2_R1113_U372 , P2_R1113_U236 , P2_R1113_U152 );
nand NAND2_19982 ( P2_R1113_U373 , P2_R1113_U202 , P2_R1113_U151 );
nand NAND2_19983 ( P2_R1113_U374 , P2_U3459 , P2_R1113_U28 );
nand NAND2_19984 ( P2_R1113_U375 , P2_U3064 , P2_R1113_U25 );
nand NAND2_19985 ( P2_R1113_U376 , P2_U3459 , P2_R1113_U28 );
nand NAND2_19986 ( P2_R1113_U377 , P2_U3064 , P2_R1113_U25 );
nand NAND2_19987 ( P2_R1113_U378 , P2_R1113_U377 , P2_R1113_U376 );
nand NAND2_19988 ( P2_R1113_U379 , P2_U3456 , P2_R1113_U26 );
nand NAND2_19989 ( P2_R1113_U380 , P2_U3068 , P2_R1113_U22 );
nand NAND2_19990 ( P2_R1113_U381 , P2_R1113_U241 , P2_R1113_U43 );
nand NAND2_19991 ( P2_R1113_U382 , P2_R1113_U153 , P2_R1113_U196 );
nand NAND2_19992 ( P2_R1113_U383 , P2_U3979 , P2_R1113_U155 );
nand NAND2_19993 ( P2_R1113_U384 , P2_U3055 , P2_R1113_U154 );
nand NAND2_19994 ( P2_R1113_U385 , P2_U3979 , P2_R1113_U155 );
nand NAND2_19995 ( P2_R1113_U386 , P2_U3055 , P2_R1113_U154 );
nand NAND2_19996 ( P2_R1113_U387 , P2_R1113_U386 , P2_R1113_U385 );
nand NAND3_19997 ( P2_R1113_U388 , P2_U3968 , P2_R1113_U10 , P2_R1113_U84 );
nand NAND3_19998 ( P2_R1113_U389 , P2_R1113_U387 , P2_R1113_U83 , P2_U3054 );
nand NAND2_19999 ( P2_R1113_U390 , P2_U3968 , P2_R1113_U84 );
nand NAND2_20000 ( P2_R1113_U391 , P2_U3054 , P2_R1113_U83 );
not NOT1_20001 ( P2_R1113_U392 , P2_R1113_U129 );
nand NAND2_20002 ( P2_R1113_U393 , P2_R1113_U306 , P2_R1113_U392 );
nand NAND2_20003 ( P2_R1113_U394 , P2_R1113_U129 , P2_R1113_U157 );
nand NAND2_20004 ( P2_R1113_U395 , P2_U3969 , P2_R1113_U82 );
nand NAND2_20005 ( P2_R1113_U396 , P2_U3053 , P2_R1113_U79 );
nand NAND2_20006 ( P2_R1113_U397 , P2_U3969 , P2_R1113_U82 );
nand NAND2_20007 ( P2_R1113_U398 , P2_U3053 , P2_R1113_U79 );
nand NAND2_20008 ( P2_R1113_U399 , P2_R1113_U398 , P2_R1113_U397 );
nand NAND2_20009 ( P2_R1113_U400 , P2_U3970 , P2_R1113_U80 );
nand NAND2_20010 ( P2_R1113_U401 , P2_U3057 , P2_R1113_U44 );
nand NAND2_20011 ( P2_R1113_U402 , P2_R1113_U313 , P2_R1113_U85 );
nand NAND2_20012 ( P2_R1113_U403 , P2_R1113_U158 , P2_R1113_U300 );
nand NAND2_20013 ( P2_R1113_U404 , P2_U3971 , P2_R1113_U78 );
nand NAND2_20014 ( P2_R1113_U405 , P2_U3058 , P2_R1113_U77 );
not NOT1_20015 ( P2_R1113_U406 , P2_R1113_U132 );
nand NAND2_20016 ( P2_R1113_U407 , P2_R1113_U296 , P2_R1113_U406 );
nand NAND2_20017 ( P2_R1113_U408 , P2_R1113_U132 , P2_R1113_U159 );
nand NAND2_20018 ( P2_R1113_U409 , P2_U3972 , P2_R1113_U76 );
nand NAND2_20019 ( P2_R1113_U410 , P2_U3065 , P2_R1113_U75 );
not NOT1_20020 ( P2_R1113_U411 , P2_R1113_U133 );
nand NAND2_20021 ( P2_R1113_U412 , P2_R1113_U292 , P2_R1113_U411 );
nand NAND2_20022 ( P2_R1113_U413 , P2_R1113_U133 , P2_R1113_U160 );
nand NAND2_20023 ( P2_R1113_U414 , P2_U3973 , P2_R1113_U71 );
nand NAND2_20024 ( P2_R1113_U415 , P2_U3066 , P2_R1113_U69 );
nand NAND2_20025 ( P2_R1113_U416 , P2_R1113_U415 , P2_R1113_U414 );
nand NAND2_20026 ( P2_R1113_U417 , P2_U3974 , P2_R1113_U72 );
nand NAND2_20027 ( P2_R1113_U418 , P2_U3061 , P2_R1113_U45 );

endmodule
