// b14
// 277 inputs  (32 PIs + 245 PPIs)
// 299 outputs (54 POs + 245 PPOs)
// 9821 gates (8236 gates + 1531 inverters + 54 buffers )
// ( 1281 AND + 216 OR + 6721 NAND + 18 NOR + 54 BUFF )
// Time: Wed Mar 25 17:47:49 2009
// All copyrigh from NCKU EE TestLAB, Taiwan. [2008.12. WCL]

module b14_ras ( U3352 , U3351 , U3350 , U3349 , U3348 , U3347 ,
             U3346 , U3345 , U3344 , U3343 , U3342 , U3341 ,
             U3340 , U3339 , U3338 , U3337 , U3336 , U3335 ,
             U3334 , U3333 , U3332 , U3331 , U3330 , U3329 ,
             U3328 , U3327 , U3326 , U3325 , U3324 , U3323 ,
             U3322 , U3321 , U3458 , U3459 , U3320 , U3319 ,
             U3318 , U3317 , U3316 , U3315 , U3314 , U3313 ,
             U3312 , U3311 , U3310 , U3309 , U3308 , U3307 ,
             U3306 , U3305 , U3304 , U3303 , U3302 , U3301 ,
             U3300 , U3299 , U3298 , U3297 , U3296 , U3295 ,
             U3294 , U3293 , U3292 , U3291 , U3467 , U3469 ,
             U3471 , U3473 , U3475 , U3477 , U3479 , U3481 ,
             U3483 , U3485 , U3487 , U3489 , U3491 , U3493 ,
             U3495 , U3497 , U3499 , U3501 , U3503 , U3505 ,
             U3506 , U3507 , U3508 , U3509 , U3510 , U3511 ,
             U3512 , U3513 , U3514 , U3515 , U3516 , U3517 ,
             U3518 , U3519 , U3520 , U3521 , U3522 , U3523 ,
             U3524 , U3525 , U3526 , U3527 , U3528 , U3529 ,
             U3530 , U3531 , U3532 , U3533 , U3534 , U3535 ,
             U3536 , U3537 , U3538 , U3539 , U3540 , U3541 ,
             U3542 , U3543 , U3544 , U3545 , U3546 , U3547 ,
             U3548 , U3549 , U3290 , U3289 , U3288 , U3287 ,
             U3286 , U3285 , U3284 , U3283 , U3282 , U3281 ,
             U3280 , U3279 , U3278 , U3277 , U3276 , U3275 ,
             U3274 , U3273 , U3272 , U3271 , U3270 , U3269 ,
             U3268 , U3267 , U3266 , U3265 , U3264 , U3263 ,
             U3262 , U3354 , U3261 , U3260 , U3259 , U3258 ,
             U3257 , U3256 , U3255 , U3254 , U3253 , U3252 ,
             U3251 , U3250 , U3249 , U3248 , U3247 , U3246 ,
             U3245 , U3244 , U3243 , U3242 , U3241 , U3240 ,
             U3550 , U3551 , U3552 , U3553 , U3554 , U3555 ,
             U3556 , U3557 , U3558 , U3559 , U3560 , U3561 ,
             U3562 , U3563 , U3564 , U3565 , U3566 , U3567 ,
             U3568 , U3569 , U3570 , U3571 , U3572 , U3573 ,
             U3574 , U3575 , U3576 , U3577 , U3578 , U3579 ,
             U3580 , U3581 , U3239 , U3238 , U3237 , U3236 ,
             U3235 , U3234 , U3233 , U3232 , U3231 , U3230 ,
             U3229 , U3228 , U3227 , U3226 , U3225 , U3224 ,
             U3223 , U3222 , U3221 , U3220 , U3219 , U3218 ,
             U3217 , U3216 , U3215 , U3214 , U3213 , U3212 ,
             U3211 , U3210 , U3149 , U3148 , U4043 , ADDR_REG_19_ ,
             ADDR_REG_18_ , ADDR_REG_17_ , ADDR_REG_16_ , ADDR_REG_15_ , ADDR_REG_14_ , ADDR_REG_13_ ,
             ADDR_REG_12_ , ADDR_REG_11_ , ADDR_REG_10_ , ADDR_REG_9_ , ADDR_REG_8_ , ADDR_REG_7_ ,
             ADDR_REG_6_ , ADDR_REG_5_ , ADDR_REG_4_ , ADDR_REG_3_ , ADDR_REG_2_ , ADDR_REG_1_ ,
             ADDR_REG_0_ , DATAO_REG_31_ , DATAO_REG_30_ , DATAO_REG_29_ , DATAO_REG_28_ , DATAO_REG_27_ ,
             DATAO_REG_26_ , DATAO_REG_25_ , DATAO_REG_24_ , DATAO_REG_23_ , DATAO_REG_22_ , DATAO_REG_21_ ,
             DATAO_REG_20_ , DATAO_REG_19_ , DATAO_REG_18_ , DATAO_REG_17_ , DATAO_REG_16_ , DATAO_REG_15_ ,
             DATAO_REG_14_ , DATAO_REG_13_ , DATAO_REG_12_ , DATAO_REG_11_ , DATAO_REG_10_ , DATAO_REG_9_ ,
             DATAO_REG_8_ , DATAO_REG_7_ , DATAO_REG_6_ , DATAO_REG_5_ , DATAO_REG_4_ , DATAO_REG_3_ ,
             DATAO_REG_2_ , DATAO_REG_1_ , DATAO_REG_0_ , RD_REG , WR_REG ,
             IR_REG_0_ , IR_REG_1_ , IR_REG_2_ , IR_REG_3_ , IR_REG_4_ , IR_REG_5_ ,
             IR_REG_6_ , IR_REG_7_ , IR_REG_8_ , IR_REG_9_ , IR_REG_10_ , IR_REG_11_ ,
             IR_REG_12_ , IR_REG_13_ , IR_REG_14_ , IR_REG_15_ , IR_REG_16_ , IR_REG_17_ ,
             IR_REG_18_ , IR_REG_19_ , IR_REG_20_ , IR_REG_21_ , IR_REG_22_ , IR_REG_23_ ,
             IR_REG_24_ , IR_REG_25_ , IR_REG_26_ , IR_REG_27_ , IR_REG_28_ , IR_REG_29_ ,
             IR_REG_30_ , IR_REG_31_ , D_REG_0_ , D_REG_1_ , D_REG_2_ , D_REG_3_ ,
             D_REG_4_ , D_REG_5_ , D_REG_6_ , D_REG_7_ , D_REG_8_ , D_REG_9_ ,
             D_REG_10_ , D_REG_11_ , D_REG_12_ , D_REG_13_ , D_REG_14_ , D_REG_15_ ,
             D_REG_16_ , D_REG_17_ , D_REG_18_ , D_REG_19_ , D_REG_20_ , D_REG_21_ ,
             D_REG_22_ , D_REG_23_ , D_REG_24_ , D_REG_25_ , D_REG_26_ , D_REG_27_ ,
             D_REG_28_ , D_REG_29_ , D_REG_30_ , D_REG_31_ , REG0_REG_0_ , REG0_REG_1_ ,
             REG0_REG_2_ , REG0_REG_3_ , REG0_REG_4_ , REG0_REG_5_ , REG0_REG_6_ , REG0_REG_7_ ,
             REG0_REG_8_ , REG0_REG_9_ , REG0_REG_10_ , REG0_REG_11_ , REG0_REG_12_ , REG0_REG_13_ ,
             REG0_REG_14_ , REG0_REG_15_ , REG0_REG_16_ , REG0_REG_17_ , REG0_REG_18_ , REG0_REG_19_ ,
             REG0_REG_20_ , REG0_REG_21_ , REG0_REG_22_ , REG0_REG_23_ , REG0_REG_24_ , REG0_REG_25_ ,
             REG0_REG_26_ , REG0_REG_27_ , REG0_REG_28_ , REG0_REG_29_ , REG0_REG_30_ , REG0_REG_31_ ,
             REG1_REG_0_ , REG1_REG_1_ , REG1_REG_2_ , REG1_REG_3_ , REG1_REG_4_ , REG1_REG_5_ ,
             REG1_REG_6_ , REG1_REG_7_ , REG1_REG_8_ , REG1_REG_9_ , REG1_REG_10_ , REG1_REG_11_ ,
             REG1_REG_12_ , REG1_REG_13_ , REG1_REG_14_ , REG1_REG_15_ , REG1_REG_16_ , REG1_REG_17_ ,
             REG1_REG_18_ , REG1_REG_19_ , REG1_REG_20_ , REG1_REG_21_ , REG1_REG_22_ , REG1_REG_23_ ,
             REG1_REG_24_ , REG1_REG_25_ , REG1_REG_26_ , REG1_REG_27_ , REG1_REG_28_ , REG1_REG_29_ ,
             REG1_REG_30_ , REG1_REG_31_ , REG2_REG_0_ , REG2_REG_1_ , REG2_REG_2_ , REG2_REG_3_ ,
             REG2_REG_4_ , REG2_REG_5_ , REG2_REG_6_ , REG2_REG_7_ , REG2_REG_8_ , REG2_REG_9_ ,
             REG2_REG_10_ , REG2_REG_11_ , REG2_REG_12_ , REG2_REG_13_ , REG2_REG_14_ , REG2_REG_15_ ,
             REG2_REG_16_ , REG2_REG_17_ , REG2_REG_18_ , REG2_REG_19_ , REG2_REG_20_ , REG2_REG_21_ ,
             REG2_REG_22_ , REG2_REG_23_ , REG2_REG_24_ , REG2_REG_25_ , REG2_REG_26_ , REG2_REG_27_ ,
             REG2_REG_28_ , REG2_REG_29_ , REG2_REG_30_ , REG2_REG_31_ , ADDR_REG_19__EXTRA , ADDR_REG_18__EXTRA ,
             ADDR_REG_17__EXTRA , ADDR_REG_16__EXTRA , ADDR_REG_15__EXTRA , ADDR_REG_14__EXTRA , ADDR_REG_13__EXTRA , ADDR_REG_12__EXTRA ,
             ADDR_REG_11__EXTRA , ADDR_REG_10__EXTRA , ADDR_REG_9__EXTRA , ADDR_REG_8__EXTRA , ADDR_REG_7__EXTRA , ADDR_REG_6__EXTRA ,
             ADDR_REG_5__EXTRA , ADDR_REG_4__EXTRA , ADDR_REG_3__EXTRA , ADDR_REG_2__EXTRA , ADDR_REG_1__EXTRA , ADDR_REG_0__EXTRA ,
             DATAO_REG_0__EXTRA , DATAO_REG_1__EXTRA , DATAO_REG_2__EXTRA , DATAO_REG_3__EXTRA , DATAO_REG_4__EXTRA , DATAO_REG_5__EXTRA ,
             DATAO_REG_6__EXTRA , DATAO_REG_7__EXTRA , DATAO_REG_8__EXTRA , DATAO_REG_9__EXTRA , DATAO_REG_10__EXTRA , DATAO_REG_11__EXTRA ,
             DATAO_REG_12__EXTRA , DATAO_REG_13__EXTRA , DATAO_REG_14__EXTRA , DATAO_REG_15__EXTRA , DATAO_REG_16__EXTRA , DATAO_REG_17__EXTRA ,
             DATAO_REG_18__EXTRA , DATAO_REG_19__EXTRA , DATAO_REG_20__EXTRA , DATAO_REG_21__EXTRA , DATAO_REG_22__EXTRA , DATAO_REG_23__EXTRA ,
             DATAO_REG_24__EXTRA , DATAO_REG_25__EXTRA , DATAO_REG_26__EXTRA , DATAO_REG_27__EXTRA , DATAO_REG_28__EXTRA , DATAO_REG_29__EXTRA ,
             DATAO_REG_30__EXTRA , DATAO_REG_31__EXTRA , B_REG , REG3_REG_15_ , REG3_REG_26_ , REG3_REG_6_ ,
             REG3_REG_18_ , REG3_REG_2_ , REG3_REG_11_ , REG3_REG_22_ , REG3_REG_13_ , REG3_REG_20_ ,
             REG3_REG_0_ , REG3_REG_9_ , REG3_REG_4_ , REG3_REG_24_ , REG3_REG_17_ , REG3_REG_5_ ,
             REG3_REG_16_ , REG3_REG_25_ , REG3_REG_12_ , REG3_REG_21_ , REG3_REG_1_ , REG3_REG_8_ ,
             REG3_REG_28_ , REG3_REG_19_ , REG3_REG_3_ , REG3_REG_10_ , REG3_REG_23_ , REG3_REG_14_ ,
             REG3_REG_27_ , REG3_REG_7_ , STATE_REG , RD_REG_EXTRA , WR_REG_EXTRA , DATAI_31_ ,
             DATAI_30_ , DATAI_29_ , DATAI_28_ , DATAI_27_ , DATAI_26_ , DATAI_25_ ,
             DATAI_24_ , DATAI_23_ , DATAI_22_ , DATAI_21_ , DATAI_20_ , DATAI_19_ ,
             DATAI_18_ , DATAI_17_ , DATAI_16_ , DATAI_15_ , DATAI_14_ , DATAI_13_ ,
             DATAI_12_ , DATAI_11_ , DATAI_10_ , DATAI_9_ , DATAI_8_ , DATAI_7_ ,
             DATAI_6_ , DATAI_5_ , DATAI_4_ , DATAI_3_ , DATAI_2_ , DATAI_1_ ,
             DATAI_0_ );


output U3352 , U3351 , U3350 , U3349 , U3348 , U3347 , U3346;
output U3345 , U3344 , U3343 , U3342 , U3341 , U3340 , U3339;
output U3338 , U3337 , U3336 , U3335 , U3334 , U3333 , U3332;
output U3331 , U3330 , U3329 , U3328 , U3327 , U3326 , U3325;
output U3324 , U3323 , U3322 , U3321 , U3458 , U3459 , U3320;
output U3319 , U3318 , U3317 , U3316 , U3315 , U3314 , U3313;
output U3312 , U3311 , U3310 , U3309 , U3308 , U3307 , U3306;
output U3305 , U3304 , U3303 , U3302 , U3301 , U3300 , U3299;
output U3298 , U3297 , U3296 , U3295 , U3294 , U3293 , U3292;
output U3291 , U3467 , U3469 , U3471 , U3473 , U3475 , U3477;
output U3479 , U3481 , U3483 , U3485 , U3487 , U3489 , U3491;
output U3493 , U3495 , U3497 , U3499 , U3501 , U3503 , U3505;
output U3506 , U3507 , U3508 , U3509 , U3510 , U3511 , U3512;
output U3513 , U3514 , U3515 , U3516 , U3517 , U3518 , U3519;
output U3520 , U3521 , U3522 , U3523 , U3524 , U3525 , U3526;
output U3527 , U3528 , U3529 , U3530 , U3531 , U3532 , U3533;
output U3534 , U3535 , U3536 , U3537 , U3538 , U3539 , U3540;
output U3541 , U3542 , U3543 , U3544 , U3545 , U3546 , U3547;
output U3548 , U3549 , U3290 , U3289 , U3288 , U3287 , U3286;
output U3285 , U3284 , U3283 , U3282 , U3281 , U3280 , U3279;
output U3278 , U3277 , U3276 , U3275 , U3274 , U3273 , U3272;
output U3271 , U3270 , U3269 , U3268 , U3267 , U3266 , U3265;
output U3264 , U3263 , U3262 , U3354 , U3261 , U3260 , U3259;
output U3258 , U3257 , U3256 , U3255 , U3254 , U3253 , U3252;
output U3251 , U3250 , U3249 , U3248 , U3247 , U3246 , U3245;
output U3244 , U3243 , U3242 , U3241 , U3240 , U3550 , U3551;
output U3552 , U3553 , U3554 , U3555 , U3556 , U3557 , U3558;
output U3559 , U3560 , U3561 , U3562 , U3563 , U3564 , U3565;
output U3566 , U3567 , U3568 , U3569 , U3570 , U3571 , U3572;
output U3573 , U3574 , U3575 , U3576 , U3577 , U3578 , U3579;
output U3580 , U3581 , U3239 , U3238 , U3237 , U3236 , U3235;
output U3234 , U3233 , U3232 , U3231 , U3230 , U3229 , U3228;
output U3227 , U3226 , U3225 , U3224 , U3223 , U3222 , U3221;
output U3220 , U3219 , U3218 , U3217 , U3216 , U3215 , U3214;
output U3213 , U3212 , U3211 , U3210 , U3149 , U3148 , U4043;
output ADDR_REG_19_ , ADDR_REG_18_ , ADDR_REG_17_ , ADDR_REG_16_ , ADDR_REG_15_ , ADDR_REG_14_;
output ADDR_REG_13_ , ADDR_REG_12_ , ADDR_REG_11_ , ADDR_REG_10_ , ADDR_REG_9_ , ADDR_REG_8_;
output ADDR_REG_7_ , ADDR_REG_6_ , ADDR_REG_5_ , ADDR_REG_4_ , ADDR_REG_3_ , ADDR_REG_2_;
output ADDR_REG_1_ , ADDR_REG_0_ , DATAO_REG_31_ , DATAO_REG_30_ , DATAO_REG_29_ , DATAO_REG_28_;
output DATAO_REG_27_ , DATAO_REG_26_ , DATAO_REG_25_ , DATAO_REG_24_ , DATAO_REG_23_ , DATAO_REG_22_;
output DATAO_REG_21_ , DATAO_REG_20_ , DATAO_REG_19_ , DATAO_REG_18_ , DATAO_REG_17_ , DATAO_REG_16_;
output DATAO_REG_15_ , DATAO_REG_14_ , DATAO_REG_13_ , DATAO_REG_12_ , DATAO_REG_11_ , DATAO_REG_10_;
output DATAO_REG_9_ , DATAO_REG_8_ , DATAO_REG_7_ , DATAO_REG_6_ , DATAO_REG_5_ , DATAO_REG_4_;
output DATAO_REG_3_ , DATAO_REG_2_ , DATAO_REG_1_ , DATAO_REG_0_ , RD_REG , WR_REG;



input IR_REG_0_ , IR_REG_1_ , IR_REG_2_ , IR_REG_3_ , IR_REG_4_ , IR_REG_5_;
input IR_REG_6_ , IR_REG_7_ , IR_REG_8_ , IR_REG_9_ , IR_REG_10_ , IR_REG_11_;
input IR_REG_12_ , IR_REG_13_ , IR_REG_14_ , IR_REG_15_ , IR_REG_16_ , IR_REG_17_;
input IR_REG_18_ , IR_REG_19_ , IR_REG_20_ , IR_REG_21_ , IR_REG_22_ , IR_REG_23_;
input IR_REG_24_ , IR_REG_25_ , IR_REG_26_ , IR_REG_27_ , IR_REG_28_ , IR_REG_29_;
input IR_REG_30_ , IR_REG_31_ , D_REG_0_ , D_REG_1_ , D_REG_2_ , D_REG_3_;
input D_REG_4_ , D_REG_5_ , D_REG_6_ , D_REG_7_ , D_REG_8_ , D_REG_9_;
input D_REG_10_ , D_REG_11_ , D_REG_12_ , D_REG_13_ , D_REG_14_ , D_REG_15_;
input D_REG_16_ , D_REG_17_ , D_REG_18_ , D_REG_19_ , D_REG_20_ , D_REG_21_;
input D_REG_22_ , D_REG_23_ , D_REG_24_ , D_REG_25_ , D_REG_26_ , D_REG_27_;
input D_REG_28_ , D_REG_29_ , D_REG_30_ , D_REG_31_ , REG0_REG_0_ , REG0_REG_1_;
input REG0_REG_2_ , REG0_REG_3_ , REG0_REG_4_ , REG0_REG_5_ , REG0_REG_6_ , REG0_REG_7_;
input REG0_REG_8_ , REG0_REG_9_ , REG0_REG_10_ , REG0_REG_11_ , REG0_REG_12_ , REG0_REG_13_;
input REG0_REG_14_ , REG0_REG_15_ , REG0_REG_16_ , REG0_REG_17_ , REG0_REG_18_ , REG0_REG_19_;
input REG0_REG_20_ , REG0_REG_21_ , REG0_REG_22_ , REG0_REG_23_ , REG0_REG_24_ , REG0_REG_25_;
input REG0_REG_26_ , REG0_REG_27_ , REG0_REG_28_ , REG0_REG_29_ , REG0_REG_30_ , REG0_REG_31_;
input REG1_REG_0_ , REG1_REG_1_ , REG1_REG_2_ , REG1_REG_3_ , REG1_REG_4_ , REG1_REG_5_;
input REG1_REG_6_ , REG1_REG_7_ , REG1_REG_8_ , REG1_REG_9_ , REG1_REG_10_ , REG1_REG_11_;
input REG1_REG_12_ , REG1_REG_13_ , REG1_REG_14_ , REG1_REG_15_ , REG1_REG_16_ , REG1_REG_17_;
input REG1_REG_18_ , REG1_REG_19_ , REG1_REG_20_ , REG1_REG_21_ , REG1_REG_22_ , REG1_REG_23_;
input REG1_REG_24_ , REG1_REG_25_ , REG1_REG_26_ , REG1_REG_27_ , REG1_REG_28_ , REG1_REG_29_;
input REG1_REG_30_ , REG1_REG_31_ , REG2_REG_0_ , REG2_REG_1_ , REG2_REG_2_ , REG2_REG_3_;
input REG2_REG_4_ , REG2_REG_5_ , REG2_REG_6_ , REG2_REG_7_ , REG2_REG_8_ , REG2_REG_9_;
input REG2_REG_10_ , REG2_REG_11_ , REG2_REG_12_ , REG2_REG_13_ , REG2_REG_14_ , REG2_REG_15_;
input REG2_REG_16_ , REG2_REG_17_ , REG2_REG_18_ , REG2_REG_19_ , REG2_REG_20_ , REG2_REG_21_;
input REG2_REG_22_ , REG2_REG_23_ , REG2_REG_24_ , REG2_REG_25_ , REG2_REG_26_ , REG2_REG_27_;
input REG2_REG_28_ , REG2_REG_29_ , REG2_REG_30_ , REG2_REG_31_ , ADDR_REG_19__EXTRA , ADDR_REG_18__EXTRA;
input ADDR_REG_17__EXTRA , ADDR_REG_16__EXTRA , ADDR_REG_15__EXTRA , ADDR_REG_14__EXTRA , ADDR_REG_13__EXTRA , ADDR_REG_12__EXTRA;
input ADDR_REG_11__EXTRA , ADDR_REG_10__EXTRA , ADDR_REG_9__EXTRA , ADDR_REG_8__EXTRA , ADDR_REG_7__EXTRA , ADDR_REG_6__EXTRA;
input ADDR_REG_5__EXTRA , ADDR_REG_4__EXTRA , ADDR_REG_3__EXTRA , ADDR_REG_2__EXTRA , ADDR_REG_1__EXTRA , ADDR_REG_0__EXTRA;
input DATAO_REG_0__EXTRA , DATAO_REG_1__EXTRA , DATAO_REG_2__EXTRA , DATAO_REG_3__EXTRA , DATAO_REG_4__EXTRA , DATAO_REG_5__EXTRA;
input DATAO_REG_6__EXTRA , DATAO_REG_7__EXTRA , DATAO_REG_8__EXTRA , DATAO_REG_9__EXTRA , DATAO_REG_10__EXTRA , DATAO_REG_11__EXTRA;
input DATAO_REG_12__EXTRA , DATAO_REG_13__EXTRA , DATAO_REG_14__EXTRA , DATAO_REG_15__EXTRA , DATAO_REG_16__EXTRA , DATAO_REG_17__EXTRA;
input DATAO_REG_18__EXTRA , DATAO_REG_19__EXTRA , DATAO_REG_20__EXTRA , DATAO_REG_21__EXTRA , DATAO_REG_22__EXTRA , DATAO_REG_23__EXTRA;
input DATAO_REG_24__EXTRA , DATAO_REG_25__EXTRA , DATAO_REG_26__EXTRA , DATAO_REG_27__EXTRA , DATAO_REG_28__EXTRA , DATAO_REG_29__EXTRA;
input DATAO_REG_30__EXTRA , DATAO_REG_31__EXTRA , B_REG , REG3_REG_15_ , REG3_REG_26_ , REG3_REG_6_;
input REG3_REG_18_ , REG3_REG_2_ , REG3_REG_11_ , REG3_REG_22_ , REG3_REG_13_ , REG3_REG_20_;
input REG3_REG_0_ , REG3_REG_9_ , REG3_REG_4_ , REG3_REG_24_ , REG3_REG_17_ , REG3_REG_5_;
input REG3_REG_16_ , REG3_REG_25_ , REG3_REG_12_ , REG3_REG_21_ , REG3_REG_1_ , REG3_REG_8_;
input REG3_REG_28_ , REG3_REG_19_ , REG3_REG_3_ , REG3_REG_10_ , REG3_REG_23_ , REG3_REG_14_;
input REG3_REG_27_ , REG3_REG_7_ , STATE_REG , RD_REG_EXTRA , WR_REG_EXTRA;
input DATAI_31_ , DATAI_30_ , DATAI_29_ , DATAI_28_ , DATAI_27_ , DATAI_26_;
input DATAI_25_ , DATAI_24_ , DATAI_23_ , DATAI_22_ , DATAI_21_ , DATAI_20_;
input DATAI_19_ , DATAI_18_ , DATAI_17_ , DATAI_16_ , DATAI_15_ , DATAI_14_;
input DATAI_13_ , DATAI_12_ , DATAI_11_ , DATAI_10_ , DATAI_9_ , DATAI_8_;
input DATAI_7_ , DATAI_6_ , DATAI_5_ , DATAI_4_ , DATAI_3_ , DATAI_2_;
input DATAI_1_ , DATAI_0_;

wire R1222_U519 , R1222_U518 , R1222_U517 , U3014 , U3015 , U3016 , U3017 , U3018 , U3019 , U3020;
wire U3021 , U3022 , U3023 , U3024 , U3025 , U3026 , U3027 , U3028 , U3029 , U3030;
wire U3031 , U3032 , U3033 , U3034 , U3035 , U3036 , U3037 , U3038 , U3039 , U3040;
wire U3041 , U3042 , U3043 , U3044 , U3045 , U3046 , U3047 , U3048 , U3049 , U3050;
wire U3051 , U3052 , U3053 , U3054 , U3055 , U3056 , U3057 , U3058 , U3059 , U3060;
wire U3061 , U3062 , U3063 , U3064 , U3065 , U3066 , U3067 , U3068 , U3069 , U3070;
wire U3071 , U3072 , U3073 , U3074 , U3075 , U3076 , U3077 , U3078 , U3079 , U3080;
wire U3081 , U3082 , U3083 , U3084 , U3085 , U3086 , U3087 , U3088 , U3089 , U3090;
wire U3091 , U3092 , U3093 , U3094 , U3095 , U3096 , U3097 , U3098 , U3099 , U3100;
wire U3101 , U3102 , U3103 , U3104 , U3105 , U3106 , U3107 , U3108 , U3109 , U3110;
wire U3111 , U3112 , U3113 , U3114 , U3115 , U3116 , U3117 , U3118 , U3119 , U3120;
wire U3121 , U3122 , U3123 , U3124 , U3125 , U3126 , U3127 , U3128 , U3129 , U3130;
wire U3131 , U3132 , U3133 , U3134 , U3135 , U3136 , U3137 , U3138 , U3139 , U3140;
wire U3141 , U3142 , U3143 , U3144 , U3145 , U3146 , U3147 , U3150 , U3151 , U3152;
wire U3153 , U3154 , U3155 , U3156 , U3157 , U3158 , U3159 , U3160 , U3161 , U3162;
wire U3163 , U3164 , U3165 , U3166 , U3167 , U3168 , U3169 , U3170 , U3171 , U3172;
wire U3173 , U3174 , U3175 , U3176 , U3177 , U3178 , U3179 , U3180 , U3181 , U3182;
wire U3183 , U3184 , U3185 , U3186 , U3187 , U3188 , U3189 , U3190 , U3191 , U3192;
wire U3193 , U3194 , U3195 , U3196 , U3197 , U3198 , U3199 , U3200 , U3201 , U3202;
wire U3203 , U3204 , U3205 , U3206 , U3207 , U3208 , U3209 , U3353 , U3355 , U3356;
wire U3357 , U3358 , U3359 , U3360 , U3361 , U3362 , U3363 , U3364 , U3365 , U3366;
wire U3367 , U3368 , U3369 , U3370 , U3371 , U3372 , U3373 , U3374 , U3375 , U3376;
wire U3377 , U3378 , U3379 , U3380 , U3381 , U3382 , U3383 , U3384 , U3385 , U3386;
wire U3387 , U3388 , U3389 , U3390 , U3391 , U3392 , U3393 , U3394 , U3395 , U3396;
wire U3397 , U3398 , U3399 , U3400 , U3401 , U3402 , U3403 , U3404 , U3405 , U3406;
wire U3407 , U3408 , U3409 , U3410 , U3411 , U3412 , U3413 , U3414 , U3415 , U3416;
wire U3417 , U3418 , U3419 , U3420 , U3421 , U3422 , U3423 , U3424 , U3425 , U3426;
wire U3427 , U3428 , U3429 , U3430 , U3431 , U3432 , U3433 , U3434 , U3435 , U3436;
wire U3437 , U3438 , U3439 , U3440 , U3441 , U3442 , U3443 , U3444 , U3445 , U3446;
wire U3447 , U3448 , U3449 , U3450 , U3451 , U3452 , U3453 , U3454 , U3455 , U3456;
wire U3457 , U3460 , U3461 , U3462 , U3463 , U3464 , U3465 , U3466 , U3468 , U3470;
wire U3472 , U3474 , U3476 , U3478 , U3480 , U3482 , U3484 , U3486 , U3488 , U3490;
wire U3492 , U3494 , U3496 , U3498 , U3500 , U3502 , U3504 , U3582 , U3583 , U3584;
wire U3585 , U3586 , U3587 , U3588 , U3589 , U3590 , U3591 , U3592 , U3593 , U3594;
wire U3595 , U3596 , U3597 , U3598 , U3599 , U3600 , U3601 , U3602 , U3603 , U3604;
wire U3605 , U3606 , U3607 , U3608 , U3609 , U3610 , U3611 , U3612 , U3613 , U3614;
wire U3615 , U3616 , U3617 , U3618 , U3619 , U3620 , U3621 , U3622 , U3623 , U3624;
wire U3625 , U3626 , U3627 , U3628 , U3629 , U3630 , U3631 , U3632 , U3633 , U3634;
wire U3635 , U3636 , U3637 , U3638 , U3639 , U3640 , U3641 , U3642 , U3643 , U3644;
wire U3645 , U3646 , U3647 , U3648 , U3649 , U3650 , U3651 , U3652 , U3653 , U3654;
wire U3655 , U3656 , U3657 , U3658 , U3659 , U3660 , U3661 , U3662 , U3663 , U3664;
wire U3665 , U3666 , U3667 , U3668 , U3669 , U3670 , U3671 , U3672 , U3673 , U3674;
wire U3675 , U3676 , U3677 , U3678 , U3679 , U3680 , U3681 , U3682 , U3683 , U3684;
wire U3685 , U3686 , U3687 , U3688 , U3689 , U3690 , U3691 , U3692 , U3693 , U3694;
wire U3695 , U3696 , U3697 , U3698 , U3699 , U3700 , U3701 , U3702 , U3703 , U3704;
wire U3705 , U3706 , U3707 , U3708 , U3709 , U3710 , U3711 , U3712 , U3713 , U3714;
wire U3715 , U3716 , U3717 , U3718 , U3719 , U3720 , U3721 , U3722 , U3723 , U3724;
wire U3725 , U3726 , U3727 , U3728 , U3729 , U3730 , U3731 , U3732 , U3733 , U3734;
wire U3735 , U3736 , U3737 , U3738 , U3739 , U3740 , U3741 , U3742 , U3743 , U3744;
wire U3745 , U3746 , U3747 , U3748 , U3749 , U3750 , U3751 , U3752 , U3753 , U3754;
wire U3755 , U3756 , U3757 , U3758 , U3759 , U3760 , U3761 , U3762 , U3763 , U3764;
wire U3765 , U3766 , U3767 , U3768 , U3769 , U3770 , U3771 , U3772 , U3773 , U3774;
wire U3775 , U3776 , U3777 , U3778 , U3779 , U3780 , U3781 , U3782 , U3783 , U3784;
wire U3785 , U3786 , U3787 , U3788 , U3789 , U3790 , U3791 , U3792 , U3793 , U3794;
wire U3795 , U3796 , U3797 , U3798 , U3799 , U3800 , U3801 , U3802 , U3803 , U3804;
wire U3805 , U3806 , U3807 , U3808 , U3809 , U3810 , U3811 , U3812 , U3813 , U3814;
wire U3815 , U3816 , U3817 , U3818 , U3819 , U3820 , U3821 , U3822 , U3823 , U3824;
wire U3825 , U3826 , U3827 , U3828 , U3829 , U3830 , U3831 , U3832 , U3833 , U3834;
wire U3835 , U3836 , U3837 , U3838 , U3839 , U3840 , U3841 , U3842 , U3843 , U3844;
wire U3845 , U3846 , U3847 , U3848 , U3849 , U3850 , U3851 , U3852 , U3853 , U3854;
wire U3855 , U3856 , U3857 , U3858 , U3859 , U3860 , U3861 , U3862 , U3863 , U3864;
wire U3865 , U3866 , U3867 , U3868 , U3869 , U3870 , U3871 , U3872 , U3873 , U3874;
wire U3875 , U3876 , U3877 , U3878 , U3879 , U3880 , U3881 , U3882 , U3883 , U3884;
wire U3885 , U3886 , U3887 , U3888 , U3889 , U3890 , U3891 , U3892 , U3893 , U3894;
wire U3895 , U3896 , U3897 , U3898 , U3899 , U3900 , U3901 , U3902 , U3903 , U3904;
wire U3905 , U3906 , U3907 , U3908 , U3909 , U3910 , U3911 , U3912 , U3913 , U3914;
wire U3915 , U3916 , U3917 , U3918 , U3919 , U3920 , U3921 , U3922 , U3923 , U3924;
wire U3925 , U3926 , U3927 , U3928 , U3929 , U3930 , U3931 , U3932 , U3933 , U3934;
wire U3935 , U3936 , U3937 , U3938 , U3939 , U3940 , U3941 , U3942 , U3943 , U3944;
wire U3945 , U3946 , U3947 , U3948 , U3949 , U3950 , U3951 , U3952 , U3953 , U3954;
wire U3955 , U3956 , U3957 , U3958 , U3959 , U3960 , U3961 , U3962 , U3963 , U3964;
wire U3965 , U3966 , U3967 , U3968 , U3969 , U3970 , U3971 , U3972 , U3973 , U3974;
wire U3975 , U3976 , U3977 , U3978 , U3979 , U3980 , U3981 , U3982 , U3983 , U3984;
wire U3985 , U3986 , U3987 , U3988 , U3989 , U3990 , U3991 , U3992 , U3993 , U3994;
wire U3995 , U3996 , U3997 , U3998 , U3999 , U4000 , U4001 , U4002 , U4003 , U4004;
wire U4005 , U4006 , U4007 , U4008 , U4009 , U4010 , U4011 , U4012 , U4013 , U4014;
wire U4015 , U4016 , U4017 , U4018 , U4019 , U4020 , U4021 , U4022 , U4023 , U4024;
wire U4025 , U4026 , U4027 , U4028 , U4029 , U4030 , U4031 , U4032 , U4033 , U4034;
wire U4035 , U4036 , U4037 , U4038 , U4039 , U4040 , U4041 , U4042 , U4044 , U4045;
wire U4046 , U4047 , U4048 , U4049 , U4050 , U4051 , U4052 , U4053 , U4054 , U4055;
wire U4056 , U4057 , U4058 , U4059 , U4060 , U4061 , U4062 , U4063 , U4064 , U4065;
wire U4066 , U4067 , U4068 , U4069 , U4070 , U4071 , U4072 , U4073 , U4074 , U4075;
wire U4076 , U4077 , U4078 , U4079 , U4080 , U4081 , U4082 , U4083 , U4084 , U4085;
wire U4086 , U4087 , U4088 , U4089 , U4090 , U4091 , U4092 , U4093 , U4094 , U4095;
wire U4096 , U4097 , U4098 , U4099 , U4100 , U4101 , U4102 , U4103 , U4104 , U4105;
wire U4106 , U4107 , U4108 , U4109 , U4110 , U4111 , U4112 , U4113 , U4114 , U4115;
wire U4116 , U4117 , U4118 , U4119 , U4120 , U4121 , U4122 , U4123 , U4124 , U4125;
wire U4126 , U4127 , U4128 , U4129 , U4130 , U4131 , U4132 , U4133 , U4134 , U4135;
wire U4136 , U4137 , U4138 , U4139 , U4140 , U4141 , U4142 , U4143 , U4144 , U4145;
wire U4146 , U4147 , U4148 , U4149 , U4150 , U4151 , U4152 , U4153 , U4154 , U4155;
wire U4156 , U4157 , U4158 , U4159 , U4160 , U4161 , U4162 , U4163 , U4164 , U4165;
wire U4166 , U4167 , U4168 , U4169 , U4170 , U4171 , U4172 , U4173 , U4174 , U4175;
wire U4176 , U4177 , U4178 , U4179 , U4180 , U4181 , U4182 , U4183 , U4184 , U4185;
wire U4186 , U4187 , U4188 , U4189 , U4190 , U4191 , U4192 , U4193 , U4194 , U4195;
wire U4196 , U4197 , U4198 , U4199 , U4200 , U4201 , U4202 , U4203 , U4204 , U4205;
wire U4206 , U4207 , U4208 , U4209 , U4210 , U4211 , U4212 , U4213 , U4214 , U4215;
wire U4216 , U4217 , U4218 , U4219 , U4220 , U4221 , U4222 , U4223 , U4224 , U4225;
wire U4226 , U4227 , U4228 , U4229 , U4230 , U4231 , U4232 , U4233 , U4234 , U4235;
wire U4236 , U4237 , U4238 , U4239 , U4240 , U4241 , U4242 , U4243 , U4244 , U4245;
wire U4246 , U4247 , U4248 , U4249 , U4250 , U4251 , U4252 , U4253 , U4254 , U4255;
wire U4256 , U4257 , U4258 , U4259 , U4260 , U4261 , U4262 , U4263 , U4264 , U4265;
wire U4266 , U4267 , U4268 , U4269 , U4270 , U4271 , U4272 , U4273 , U4274 , U4275;
wire U4276 , U4277 , U4278 , U4279 , U4280 , U4281 , U4282 , U4283 , U4284 , U4285;
wire U4286 , U4287 , U4288 , U4289 , U4290 , U4291 , U4292 , U4293 , U4294 , U4295;
wire U4296 , U4297 , U4298 , U4299 , U4300 , U4301 , U4302 , U4303 , U4304 , U4305;
wire U4306 , U4307 , U4308 , U4309 , U4310 , U4311 , U4312 , U4313 , U4314 , U4315;
wire U4316 , U4317 , U4318 , U4319 , U4320 , U4321 , U4322 , U4323 , U4324 , U4325;
wire U4326 , U4327 , U4328 , U4329 , U4330 , U4331 , U4332 , U4333 , U4334 , U4335;
wire U4336 , U4337 , U4338 , U4339 , U4340 , U4341 , U4342 , U4343 , U4344 , U4345;
wire U4346 , U4347 , U4348 , U4349 , U4350 , U4351 , U4352 , U4353 , U4354 , U4355;
wire U4356 , U4357 , U4358 , U4359 , U4360 , U4361 , U4362 , U4363 , U4364 , U4365;
wire U4366 , U4367 , U4368 , U4369 , U4370 , U4371 , U4372 , U4373 , U4374 , U4375;
wire U4376 , U4377 , U4378 , U4379 , U4380 , U4381 , U4382 , U4383 , U4384 , U4385;
wire U4386 , U4387 , U4388 , U4389 , U4390 , U4391 , U4392 , U4393 , U4394 , U4395;
wire U4396 , U4397 , U4398 , U4399 , U4400 , U4401 , U4402 , U4403 , U4404 , U4405;
wire U4406 , U4407 , U4408 , U4409 , U4410 , U4411 , U4412 , U4413 , U4414 , U4415;
wire U4416 , U4417 , U4418 , U4419 , U4420 , U4421 , U4422 , U4423 , U4424 , U4425;
wire U4426 , U4427 , U4428 , U4429 , U4430 , U4431 , U4432 , U4433 , U4434 , U4435;
wire U4436 , U4437 , U4438 , U4439 , U4440 , U4441 , U4442 , U4443 , U4444 , U4445;
wire U4446 , U4447 , U4448 , U4449 , U4450 , U4451 , U4452 , U4453 , U4454 , U4455;
wire U4456 , U4457 , U4458 , U4459 , U4460 , U4461 , U4462 , U4463 , U4464 , U4465;
wire U4466 , U4467 , U4468 , U4469 , U4470 , U4471 , U4472 , U4473 , U4474 , U4475;
wire U4476 , U4477 , U4478 , U4479 , U4480 , U4481 , U4482 , U4483 , U4484 , U4485;
wire U4486 , U4487 , U4488 , U4489 , U4490 , U4491 , U4492 , U4493 , U4494 , U4495;
wire U4496 , U4497 , U4498 , U4499 , U4500 , U4501 , U4502 , U4503 , U4504 , U4505;
wire U4506 , U4507 , U4508 , U4509 , U4510 , U4511 , U4512 , U4513 , U4514 , U4515;
wire U4516 , U4517 , U4518 , U4519 , U4520 , U4521 , U4522 , U4523 , U4524 , U4525;
wire U4526 , U4527 , U4528 , U4529 , U4530 , U4531 , U4532 , U4533 , U4534 , U4535;
wire U4536 , U4537 , U4538 , U4539 , U4540 , U4541 , U4542 , U4543 , U4544 , U4545;
wire U4546 , U4547 , U4548 , U4549 , U4550 , U4551 , U4552 , U4553 , U4554 , U4555;
wire U4556 , U4557 , U4558 , U4559 , U4560 , U4561 , U4562 , U4563 , U4564 , U4565;
wire U4566 , U4567 , U4568 , U4569 , U4570 , U4571 , U4572 , U4573 , U4574 , U4575;
wire U4576 , U4577 , U4578 , U4579 , U4580 , U4581 , U4582 , U4583 , U4584 , U4585;
wire U4586 , U4587 , U4588 , U4589 , U4590 , U4591 , U4592 , U4593 , U4594 , U4595;
wire U4596 , U4597 , U4598 , U4599 , U4600 , U4601 , U4602 , U4603 , U4604 , U4605;
wire U4606 , U4607 , U4608 , U4609 , U4610 , U4611 , U4612 , U4613 , U4614 , U4615;
wire U4616 , U4617 , U4618 , U4619 , U4620 , U4621 , U4622 , U4623 , U4624 , U4625;
wire U4626 , U4627 , U4628 , U4629 , U4630 , U4631 , U4632 , U4633 , U4634 , U4635;
wire U4636 , U4637 , U4638 , U4639 , U4640 , U4641 , U4642 , U4643 , U4644 , U4645;
wire U4646 , U4647 , U4648 , U4649 , U4650 , U4651 , U4652 , U4653 , U4654 , U4655;
wire U4656 , U4657 , U4658 , U4659 , U4660 , U4661 , U4662 , U4663 , U4664 , U4665;
wire U4666 , U4667 , U4668 , U4669 , U4670 , U4671 , U4672 , U4673 , U4674 , U4675;
wire U4676 , U4677 , U4678 , U4679 , U4680 , U4681 , U4682 , U4683 , U4684 , U4685;
wire U4686 , U4687 , U4688 , U4689 , U4690 , U4691 , U4692 , U4693 , U4694 , U4695;
wire U4696 , U4697 , U4698 , U4699 , U4700 , U4701 , U4702 , U4703 , U4704 , U4705;
wire U4706 , U4707 , U4708 , U4709 , U4710 , U4711 , U4712 , U4713 , U4714 , U4715;
wire U4716 , U4717 , U4718 , U4719 , U4720 , U4721 , U4722 , U4723 , U4724 , U4725;
wire U4726 , U4727 , U4728 , U4729 , U4730 , U4731 , U4732 , U4733 , U4734 , U4735;
wire U4736 , U4737 , U4738 , U4739 , U4740 , U4741 , U4742 , U4743 , U4744 , U4745;
wire U4746 , U4747 , U4748 , U4749 , U4750 , U4751 , U4752 , U4753 , U4754 , U4755;
wire U4756 , U4757 , U4758 , U4759 , U4760 , U4761 , U4762 , U4763 , U4764 , U4765;
wire U4766 , U4767 , U4768 , U4769 , U4770 , U4771 , U4772 , U4773 , U4774 , U4775;
wire U4776 , U4777 , U4778 , U4779 , U4780 , U4781 , U4782 , U4783 , U4784 , U4785;
wire U4786 , U4787 , U4788 , U4789 , U4790 , U4791 , U4792 , U4793 , U4794 , U4795;
wire U4796 , U4797 , U4798 , U4799 , U4800 , U4801 , U4802 , U4803 , U4804 , U4805;
wire U4806 , U4807 , U4808 , U4809 , U4810 , U4811 , U4812 , U4813 , U4814 , U4815;
wire U4816 , U4817 , U4818 , U4819 , U4820 , U4821 , U4822 , U4823 , U4824 , U4825;
wire U4826 , U4827 , U4828 , U4829 , U4830 , U4831 , U4832 , U4833 , U4834 , U4835;
wire U4836 , U4837 , U4838 , U4839 , U4840 , U4841 , U4842 , U4843 , U4844 , U4845;
wire U4846 , U4847 , U4848 , U4849 , U4850 , U4851 , U4852 , U4853 , U4854 , U4855;
wire U4856 , U4857 , U4858 , U4859 , U4860 , U4861 , U4862 , U4863 , U4864 , U4865;
wire U4866 , U4867 , U4868 , U4869 , U4870 , U4871 , U4872 , U4873 , U4874 , U4875;
wire U4876 , U4877 , U4878 , U4879 , U4880 , U4881 , U4882 , U4883 , U4884 , U4885;
wire U4886 , U4887 , U4888 , U4889 , U4890 , U4891 , U4892 , U4893 , U4894 , U4895;
wire U4896 , U4897 , U4898 , U4899 , U4900 , U4901 , U4902 , U4903 , U4904 , U4905;
wire U4906 , U4907 , U4908 , U4909 , U4910 , U4911 , U4912 , U4913 , U4914 , U4915;
wire U4916 , U4917 , U4918 , U4919 , U4920 , U4921 , U4922 , U4923 , U4924 , U4925;
wire U4926 , U4927 , U4928 , U4929 , U4930 , U4931 , U4932 , U4933 , U4934 , U4935;
wire U4936 , U4937 , U4938 , U4939 , U4940 , U4941 , U4942 , U4943 , U4944 , U4945;
wire U4946 , U4947 , U4948 , U4949 , U4950 , U4951 , U4952 , U4953 , U4954 , U4955;
wire U4956 , U4957 , U4958 , U4959 , U4960 , U4961 , U4962 , U4963 , U4964 , U4965;
wire U4966 , U4967 , U4968 , U4969 , U4970 , U4971 , U4972 , U4973 , U4974 , U4975;
wire U4976 , U4977 , U4978 , U4979 , U4980 , U4981 , U4982 , U4983 , U4984 , U4985;
wire U4986 , U4987 , U4988 , U4989 , U4990 , U4991 , U4992 , U4993 , U4994 , U4995;
wire U4996 , U4997 , U4998 , U4999 , U5000 , U5001 , U5002 , U5003 , U5004 , U5005;
wire U5006 , U5007 , U5008 , U5009 , U5010 , U5011 , U5012 , U5013 , U5014 , U5015;
wire U5016 , U5017 , U5018 , U5019 , U5020 , U5021 , U5022 , U5023 , U5024 , U5025;
wire U5026 , U5027 , U5028 , U5029 , U5030 , U5031 , U5032 , U5033 , U5034 , U5035;
wire U5036 , U5037 , U5038 , U5039 , U5040 , U5041 , U5042 , U5043 , U5044 , U5045;
wire U5046 , U5047 , U5048 , U5049 , U5050 , U5051 , U5052 , U5053 , U5054 , U5055;
wire U5056 , U5057 , U5058 , U5059 , U5060 , U5061 , U5062 , U5063 , U5064 , U5065;
wire U5066 , U5067 , U5068 , U5069 , U5070 , U5071 , U5072 , U5073 , U5074 , U5075;
wire U5076 , U5077 , U5078 , U5079 , U5080 , U5081 , U5082 , U5083 , U5084 , U5085;
wire U5086 , U5087 , U5088 , U5089 , U5090 , U5091 , U5092 , U5093 , U5094 , U5095;
wire U5096 , U5097 , U5098 , U5099 , U5100 , U5101 , U5102 , U5103 , U5104 , U5105;
wire U5106 , U5107 , U5108 , U5109 , U5110 , U5111 , U5112 , U5113 , U5114 , U5115;
wire U5116 , U5117 , U5118 , U5119 , U5120 , U5121 , U5122 , U5123 , U5124 , U5125;
wire U5126 , U5127 , U5128 , U5129 , U5130 , U5131 , U5132 , U5133 , U5134 , U5135;
wire U5136 , U5137 , U5138 , U5139 , U5140 , U5141 , U5142 , U5143 , U5144 , U5145;
wire U5146 , U5147 , U5148 , U5149 , U5150 , U5151 , U5152 , U5153 , U5154 , U5155;
wire U5156 , U5157 , U5158 , U5159 , U5160 , U5161 , U5162 , U5163 , U5164 , U5165;
wire U5166 , U5167 , U5168 , U5169 , U5170 , U5171 , U5172 , U5173 , U5174 , U5175;
wire U5176 , U5177 , U5178 , U5179 , U5180 , U5181 , U5182 , U5183 , U5184 , U5185;
wire U5186 , U5187 , U5188 , U5189 , U5190 , U5191 , U5192 , U5193 , U5194 , U5195;
wire U5196 , U5197 , U5198 , U5199 , U5200 , U5201 , U5202 , U5203 , U5204 , U5205;
wire U5206 , U5207 , U5208 , U5209 , U5210 , U5211 , U5212 , U5213 , U5214 , U5215;
wire U5216 , U5217 , U5218 , U5219 , U5220 , U5221 , U5222 , U5223 , U5224 , U5225;
wire U5226 , U5227 , U5228 , U5229 , U5230 , U5231 , U5232 , U5233 , U5234 , U5235;
wire U5236 , U5237 , U5238 , U5239 , U5240 , U5241 , U5242 , U5243 , U5244 , U5245;
wire U5246 , U5247 , U5248 , U5249 , U5250 , U5251 , U5252 , U5253 , U5254 , U5255;
wire U5256 , U5257 , U5258 , U5259 , U5260 , U5261 , U5262 , U5263 , U5264 , U5265;
wire U5266 , U5267 , U5268 , U5269 , U5270 , U5271 , U5272 , U5273 , U5274 , U5275;
wire U5276 , U5277 , U5278 , U5279 , U5280 , U5281 , U5282 , U5283 , U5284 , U5285;
wire U5286 , U5287 , U5288 , U5289 , U5290 , U5291 , U5292 , U5293 , U5294 , U5295;
wire U5296 , U5297 , U5298 , U5299 , U5300 , U5301 , U5302 , U5303 , U5304 , U5305;
wire U5306 , U5307 , U5308 , U5309 , U5310 , U5311 , U5312 , U5313 , U5314 , U5315;
wire U5316 , U5317 , U5318 , U5319 , U5320 , U5321 , U5322 , U5323 , U5324 , U5325;
wire U5326 , U5327 , U5328 , U5329 , U5330 , U5331 , U5332 , U5333 , U5334 , U5335;
wire U5336 , U5337 , U5338 , U5339 , U5340 , U5341 , U5342 , U5343 , U5344 , U5345;
wire U5346 , U5347 , U5348 , U5349 , U5350 , U5351 , U5352 , U5353 , U5354 , U5355;
wire U5356 , U5357 , U5358 , U5359 , U5360 , U5361 , U5362 , U5363 , U5364 , U5365;
wire U5366 , U5367 , U5368 , U5369 , U5370 , U5371 , U5372 , U5373 , U5374 , U5375;
wire U5376 , U5377 , U5378 , U5379 , U5380 , U5381 , U5382 , U5383 , U5384 , U5385;
wire U5386 , U5387 , U5388 , U5389 , U5390 , U5391 , U5392 , U5393 , U5394 , U5395;
wire U5396 , U5397 , U5398 , U5399 , U5400 , U5401 , U5402 , U5403 , U5404 , U5405;
wire U5406 , U5407 , U5408 , U5409 , U5410 , U5411 , U5412 , U5413 , U5414 , U5415;
wire U5416 , U5417 , U5418 , U5419 , U5420 , U5421 , U5422 , U5423 , U5424 , U5425;
wire U5426 , U5427 , U5428 , U5429 , U5430 , U5431 , U5432 , U5433 , U5434 , U5435;
wire U5436 , U5437 , U5438 , U5439 , U5440 , U5441 , U5442 , U5443 , U5444 , U5445;
wire U5446 , U5447 , U5448 , U5449 , U5450 , U5451 , U5452 , U5453 , U5454 , U5455;
wire U5456 , U5457 , U5458 , U5459 , U5460 , U5461 , U5462 , U5463 , U5464 , U5465;
wire U5466 , U5467 , U5468 , U5469 , U5470 , U5471 , U5472 , U5473 , U5474 , U5475;
wire U5476 , U5477 , U5478 , U5479 , U5480 , U5481 , U5482 , U5483 , U5484 , U5485;
wire U5486 , U5487 , U5488 , U5489 , U5490 , U5491 , U5492 , U5493 , U5494 , U5495;
wire U5496 , U5497 , U5498 , U5499 , U5500 , U5501 , U5502 , U5503 , U5504 , U5505;
wire U5506 , U5507 , U5508 , U5509 , U5510 , U5511 , U5512 , U5513 , U5514 , U5515;
wire U5516 , U5517 , U5518 , U5519 , U5520 , U5521 , U5522 , U5523 , U5524 , U5525;
wire U5526 , U5527 , U5528 , U5529 , U5530 , U5531 , U5532 , U5533 , U5534 , U5535;
wire U5536 , U5537 , U5538 , U5539 , U5540 , U5541 , U5542 , U5543 , U5544 , U5545;
wire U5546 , U5547 , U5548 , U5549 , U5550 , U5551 , U5552 , U5553 , U5554 , U5555;
wire U5556 , U5557 , U5558 , U5559 , U5560 , U5561 , U5562 , U5563 , U5564 , U5565;
wire U5566 , U5567 , U5568 , U5569 , U5570 , U5571 , U5572 , U5573 , U5574 , U5575;
wire U5576 , U5577 , U5578 , U5579 , U5580 , U5581 , U5582 , U5583 , U5584 , U5585;
wire U5586 , U5587 , U5588 , U5589 , U5590 , U5591 , U5592 , U5593 , U5594 , U5595;
wire U5596 , U5597 , U5598 , U5599 , U5600 , U5601 , U5602 , U5603 , U5604 , U5605;
wire U5606 , U5607 , U5608 , U5609 , U5610 , U5611 , U5612 , U5613 , U5614 , U5615;
wire U5616 , U5617 , U5618 , U5619 , U5620 , U5621 , U5622 , U5623 , U5624 , U5625;
wire U5626 , U5627 , U5628 , U5629 , U5630 , U5631 , U5632 , U5633 , U5634 , U5635;
wire U5636 , U5637 , U5638 , U5639 , U5640 , U5641 , U5642 , U5643 , U5644 , U5645;
wire U5646 , U5647 , U5648 , U5649 , U5650 , U5651 , U5652 , U5653 , U5654 , U5655;
wire U5656 , U5657 , U5658 , U5659 , U5660 , U5661 , U5662 , U5663 , U5664 , U5665;
wire U5666 , U5667 , U5668 , U5669 , U5670 , U5671 , U5672 , U5673 , U5674 , U5675;
wire U5676 , U5677 , U5678 , U5679 , U5680 , U5681 , U5682 , U5683 , U5684 , U5685;
wire U5686 , U5687 , U5688 , U5689 , U5690 , U5691 , U5692 , U5693 , U5694 , U5695;
wire U5696 , U5697 , U5698 , U5699 , U5700 , U5701 , U5702 , U5703 , U5704 , U5705;
wire U5706 , U5707 , U5708 , U5709 , U5710 , U5711 , U5712 , U5713 , U5714 , U5715;
wire U5716 , U5717 , U5718 , U5719 , U5720 , U5721 , U5722 , U5723 , U5724 , U5725;
wire U5726 , U5727 , U5728 , U5729 , U5730 , U5731 , U5732 , U5733 , U5734 , U5735;
wire U5736 , U5737 , U5738 , U5739 , U5740 , U5741 , U5742 , U5743 , U5744 , U5745;
wire U5746 , U5747 , U5748 , U5749 , U5750 , U5751 , U5752 , U5753 , U5754 , U5755;
wire U5756 , U5757 , U5758 , U5759 , U5760 , U5761 , U5762 , U5763 , U5764 , U5765;
wire U5766 , U5767 , U5768 , U5769 , U5770 , U5771 , U5772 , U5773 , U5774 , U5775;
wire U5776 , U5777 , U5778 , U5779 , U5780 , U5781 , U5782 , U5783 , U5784 , U5785;
wire U5786 , U5787 , U5788 , U5789 , U5790 , U5791 , U5792 , U5793 , U5794 , U5795;
wire U5796 , U5797 , U5798 , U5799 , U5800 , U5801 , U5802 , U5803 , U5804 , U5805;
wire U5806 , U5807 , U5808 , U5809 , U5810 , U5811 , U5812 , U5813 , U5814 , U5815;
wire U5816 , U5817 , U5818 , U5819 , U5820 , U5821 , U5822 , U5823 , U5824 , U5825;
wire U5826 , U5827 , U5828 , U5829 , U5830 , U5831 , U5832 , U5833 , U5834 , U5835;
wire U5836 , U5837 , U5838 , U5839 , U5840 , U5841 , U5842 , U5843 , U5844 , U5845;
wire U5846 , U5847 , U5848 , U5849 , U5850 , U5851 , U5852 , U5853 , U5854 , U5855;
wire U5856 , U5857 , U5858 , U5859 , U5860 , U5861 , U5862 , U5863 , U5864 , U5865;
wire U5866 , U5867 , U5868 , U5869 , U5870 , U5871 , U5872 , U5873 , U5874 , U5875;
wire U5876 , U5877 , U5878 , U5879 , U5880 , U5881 , U5882 , U5883 , U5884 , U5885;
wire U5886 , U5887 , U5888 , U5889 , U5890 , U5891 , U5892 , U5893 , U5894 , U5895;
wire U5896 , U5897 , U5898 , U5899 , U5900 , U5901 , U5902 , U5903 , U5904 , U5905;
wire U5906 , U5907 , U5908 , U5909 , U5910 , U5911 , U5912 , U5913 , U5914 , U5915;
wire U5916 , U5917 , U5918 , U5919 , U5920 , U5921 , U5922 , U5923 , U5924 , U5925;
wire U5926 , U5927 , U5928 , U5929 , U5930 , U5931 , U5932 , U5933 , U5934 , U5935;
wire U5936 , U5937 , U5938 , U5939 , U5940 , U5941 , U5942 , U5943 , U5944 , U5945;
wire U5946 , U5947 , U5948 , U5949 , U5950 , U5951 , U5952 , U5953 , U5954 , U5955;
wire U5956 , U5957 , U5958 , U5959 , U5960 , U5961 , U5962 , U5963 , U5964 , U5965;
wire U5966 , U5967 , U5968 , U5969 , U5970 , U5971 , U5972 , U5973 , U5974 , U5975;
wire U5976 , U5977 , U5978 , U5979 , U5980 , U5981 , U5982 , U5983 , U5984 , U5985;
wire U5986 , U5987 , U5988 , U5989 , U5990 , U5991 , U5992 , U5993 , U5994 , U5995;
wire U5996 , U5997 , U5998 , U5999 , U6000 , U6001 , U6002 , U6003 , U6004 , U6005;
wire U6006 , U6007 , U6008 , U6009 , U6010 , U6011 , U6012 , U6013 , U6014 , U6015;
wire U6016 , U6017 , U6018 , U6019 , U6020 , U6021 , U6022 , U6023 , U6024 , U6025;
wire U6026 , U6027 , U6028 , U6029 , U6030 , U6031 , U6032 , U6033 , U6034 , U6035;
wire U6036 , U6037 , U6038 , U6039 , U6040 , U6041 , U6042 , U6043 , U6044 , U6045;
wire U6046 , U6047 , U6048 , U6049 , U6050 , U6051 , U6052 , U6053 , U6054 , U6055;
wire U6056 , U6057 , U6058 , U6059 , U6060 , U6061 , U6062 , U6063 , U6064 , U6065;
wire U6066 , U6067 , U6068 , U6069 , U6070 , U6071 , U6072 , U6073 , U6074 , U6075;
wire U6076 , U6077 , U6078 , U6079 , U6080 , U6081 , U6082 , U6083 , U6084 , U6085;
wire U6086 , U6087 , U6088 , U6089 , U6090 , U6091 , U6092 , U6093 , U6094 , U6095;
wire U6096 , U6097 , U6098 , U6099 , U6100 , U6101 , U6102 , U6103 , U6104 , U6105;
wire U6106 , U6107 , U6108 , U6109 , U6110 , U6111 , U6112 , U6113 , U6114 , U6115;
wire U6116 , U6117 , U6118 , U6119 , U6120 , U6121 , U6122 , U6123 , U6124 , U6125;
wire U6126 , U6127 , U6128 , U6129 , U6130 , U6131 , U6132 , U6133 , U6134 , U6135;
wire U6136 , U6137 , U6138 , U6139 , U6140 , U6141 , U6142 , U6143 , U6144 , U6145;
wire U6146 , U6147 , U6148 , U6149 , U6150 , U6151 , U6152 , U6153 , U6154 , U6155;
wire U6156 , U6157 , U6158 , U6159 , U6160 , U6161 , U6162 , U6163 , U6164 , U6165;
wire U6166 , U6167 , U6168 , U6169 , U6170 , U6171 , U6172 , U6173 , U6174 , U6175;
wire U6176 , U6177 , U6178 , U6179 , U6180 , U6181 , U6182 , U6183 , U6184 , U6185;
wire U6186 , U6187 , U6188 , U6189 , U6190 , U6191 , U6192 , U6193 , U6194 , U6195;
wire U6196 , U6197 , U6198 , U6199 , U6200 , U6201 , U6202 , U6203 , U6204 , U6205;
wire U6206 , U6207 , U6208 , U6209 , U6210 , U6211 , U6212 , U6213 , U6214 , U6215;
wire U6216 , U6217 , U6218 , U6219 , U6220 , U6221 , U6222 , U6223 , U6224 , U6225;
wire U6226 , U6227 , U6228 , U6229 , U6230 , U6231 , U6232 , U6233 , U6234 , U6235;
wire U6236 , U6237 , U6238 , U6239 , U6240 , U6241 , U6242 , U6243 , U6244 , U6245;
wire U6246 , U6247 , U6248 , U6249 , U6250 , U6251 , U6252 , U6253 , U6254 , U6255;
wire U6256 , U6257 , U6258 , U6259 , U6260 , U6261 , U6262 , U6263 , U6264 , U6265;
wire U6266 , U6267 , U6268 , U6269 , U6270 , U6271 , U6272 , U6273 , U6274 , U6275;
wire U6276 , U6277 , U6278 , U6279 , U6280 , U6281 , U6282 , U6283 , U6284 , U6285;
wire U6286 , U6287 , U6288 , U6289 , U6290 , U6291 , U6292 , U6293 , U6294 , U6295;
wire U6296 , U6297 , U6298 , U6299 , U6300 , U6301 , U6302 , U6303 , U6304 , U6305;
wire U6306 , U6307 , U6308 , U6309 , U6310 , U6311 , U6312 , U6313 , U6314 , U6315;
wire U6316 , U6317 , U6318 , U6319 , U6320 , U6321 , U6322 , U6323 , R1222_U516 , R1222_U515;
wire R1222_U514 , R1222_U513 , R1222_U512 , R1222_U511 , R1222_U510 , R1222_U509 , R1222_U508 , R1222_U507 , R1222_U506 , R1222_U505;
wire R1222_U504 , R1222_U503 , R1222_U502 , R1222_U501 , R1222_U500 , R1222_U499 , R1222_U498 , R1222_U497 , R1222_U496 , R1222_U495;
wire SUB_84_U4 , SUB_84_U5 , SUB_84_U6 , SUB_84_U7 , SUB_84_U8 , SUB_84_U9 , SUB_84_U10 , SUB_84_U11 , SUB_84_U12 , SUB_84_U13;
wire SUB_84_U14 , SUB_84_U15 , SUB_84_U16 , SUB_84_U17 , SUB_84_U18 , SUB_84_U19 , SUB_84_U20 , SUB_84_U21 , SUB_84_U22 , SUB_84_U23;
wire SUB_84_U24 , SUB_84_U25 , SUB_84_U26 , SUB_84_U27 , SUB_84_U28 , SUB_84_U29 , SUB_84_U30 , SUB_84_U31 , SUB_84_U32 , SUB_84_U33;
wire SUB_84_U34 , SUB_84_U35 , SUB_84_U36 , SUB_84_U37 , SUB_84_U38 , SUB_84_U39 , SUB_84_U40 , SUB_84_U41 , SUB_84_U42 , SUB_84_U43;
wire SUB_84_U44 , SUB_84_U45 , SUB_84_U46 , SUB_84_U47 , SUB_84_U48 , SUB_84_U49 , SUB_84_U50 , SUB_84_U51 , SUB_84_U52 , SUB_84_U53;
wire SUB_84_U54 , SUB_84_U55 , SUB_84_U56 , SUB_84_U57 , SUB_84_U58 , SUB_84_U59 , SUB_84_U60 , SUB_84_U61 , SUB_84_U62 , SUB_84_U63;
wire SUB_84_U64 , SUB_84_U65 , SUB_84_U66 , SUB_84_U67 , SUB_84_U68 , SUB_84_U69 , SUB_84_U70 , SUB_84_U71 , SUB_84_U72 , SUB_84_U73;
wire SUB_84_U74 , SUB_84_U75 , SUB_84_U76 , SUB_84_U77 , SUB_84_U78 , SUB_84_U79 , SUB_84_U80 , SUB_84_U81 , SUB_84_U82 , SUB_84_U83;
wire SUB_84_U84 , SUB_84_U85 , SUB_84_U86 , SUB_84_U87 , SUB_84_U88 , SUB_84_U89 , SUB_84_U90 , SUB_84_U91 , SUB_84_U92 , SUB_84_U93;
wire SUB_84_U94 , SUB_84_U95 , SUB_84_U96 , SUB_84_U97 , SUB_84_U98 , SUB_84_U99 , SUB_84_U100 , SUB_84_U101 , SUB_84_U102 , SUB_84_U103;
wire SUB_84_U104 , SUB_84_U105 , SUB_84_U106 , SUB_84_U107 , SUB_84_U108 , SUB_84_U109 , SUB_84_U110 , SUB_84_U111 , SUB_84_U112 , SUB_84_U113;
wire SUB_84_U114 , SUB_84_U115 , SUB_84_U116 , SUB_84_U117 , SUB_84_U118 , SUB_84_U119 , SUB_84_U120 , SUB_84_U121 , SUB_84_U122 , SUB_84_U123;
wire SUB_84_U124 , SUB_84_U125 , SUB_84_U126 , SUB_84_U127 , SUB_84_U128 , SUB_84_U129 , SUB_84_U130 , SUB_84_U131 , SUB_84_U132 , SUB_84_U133;
wire SUB_84_U134 , SUB_84_U135 , SUB_84_U136 , SUB_84_U137 , SUB_84_U138 , SUB_84_U139 , SUB_84_U140 , SUB_84_U141 , SUB_84_U142 , SUB_84_U143;
wire SUB_84_U144 , SUB_84_U145 , SUB_84_U146 , SUB_84_U147 , SUB_84_U148 , SUB_84_U149 , SUB_84_U150 , SUB_84_U151 , SUB_84_U152 , SUB_84_U153;
wire SUB_84_U154 , SUB_84_U155 , SUB_84_U156 , SUB_84_U157 , SUB_84_U158 , SUB_84_U159 , SUB_84_U160 , SUB_84_U161 , ADD_95_U4 , ADD_95_U5;
wire ADD_95_U6 , ADD_95_U7 , ADD_95_U8 , ADD_95_U9 , ADD_95_U10 , ADD_95_U11 , ADD_95_U12 , ADD_95_U13 , ADD_95_U14 , ADD_95_U15;
wire ADD_95_U16 , ADD_95_U17 , ADD_95_U18 , ADD_95_U19 , ADD_95_U20 , ADD_95_U21 , ADD_95_U22 , ADD_95_U23 , ADD_95_U24 , ADD_95_U25;
wire ADD_95_U26 , ADD_95_U27 , ADD_95_U28 , ADD_95_U29 , ADD_95_U30 , ADD_95_U31 , ADD_95_U32 , ADD_95_U33 , ADD_95_U34 , ADD_95_U35;
wire ADD_95_U36 , ADD_95_U37 , ADD_95_U38 , ADD_95_U39 , ADD_95_U40 , ADD_95_U41 , ADD_95_U42 , ADD_95_U43 , ADD_95_U44 , ADD_95_U45;
wire ADD_95_U46 , ADD_95_U47 , ADD_95_U48 , ADD_95_U49 , ADD_95_U50 , ADD_95_U51 , ADD_95_U52 , ADD_95_U53 , ADD_95_U54 , ADD_95_U55;
wire ADD_95_U56 , ADD_95_U57 , ADD_95_U58 , ADD_95_U59 , ADD_95_U60 , ADD_95_U61 , ADD_95_U62 , ADD_95_U63 , ADD_95_U64 , ADD_95_U65;
wire ADD_95_U66 , ADD_95_U67 , ADD_95_U68 , ADD_95_U69 , ADD_95_U70 , ADD_95_U71 , ADD_95_U72 , ADD_95_U73 , ADD_95_U74 , ADD_95_U75;
wire ADD_95_U76 , ADD_95_U77 , ADD_95_U78 , ADD_95_U79 , ADD_95_U80 , ADD_95_U81 , ADD_95_U82 , ADD_95_U83 , ADD_95_U84 , ADD_95_U85;
wire ADD_95_U86 , ADD_95_U87 , ADD_95_U88 , ADD_95_U89 , ADD_95_U90 , ADD_95_U91 , ADD_95_U92 , ADD_95_U93 , ADD_95_U94 , ADD_95_U95;
wire ADD_95_U96 , ADD_95_U97 , ADD_95_U98 , ADD_95_U99 , ADD_95_U100 , ADD_95_U101 , ADD_95_U102 , ADD_95_U103 , ADD_95_U104 , ADD_95_U105;
wire ADD_95_U106 , ADD_95_U107 , ADD_95_U108 , ADD_95_U109 , ADD_95_U110 , ADD_95_U111 , ADD_95_U112 , ADD_95_U113 , ADD_95_U114 , ADD_95_U115;
wire ADD_95_U116 , ADD_95_U117 , ADD_95_U118 , ADD_95_U119 , ADD_95_U120 , ADD_95_U121 , ADD_95_U122 , ADD_95_U123 , ADD_95_U124 , ADD_95_U125;
wire ADD_95_U126 , ADD_95_U127 , ADD_95_U128 , ADD_95_U129 , ADD_95_U130 , ADD_95_U131 , ADD_95_U132 , ADD_95_U133 , ADD_95_U134 , ADD_95_U135;
wire ADD_95_U136 , ADD_95_U137 , ADD_95_U138 , ADD_95_U139 , ADD_95_U140 , ADD_95_U141 , ADD_95_U142 , ADD_95_U143 , ADD_95_U144 , ADD_95_U145;
wire ADD_95_U146 , ADD_95_U147 , ADD_95_U148 , ADD_95_U149 , ADD_95_U150 , ADD_95_U151 , ADD_95_U152 , ADD_95_U153 , ADD_95_U154 , ADD_95_U155;
wire ADD_95_U156 , ADD_95_U157 , ADD_95_U158 , ADD_95_U159 , R395_U6 , R395_U7 , R395_U8 , R395_U9 , R395_U10 , R395_U11;
wire R395_U12 , R395_U13 , R395_U14 , R395_U15 , R395_U16 , R395_U17 , R395_U18 , R395_U19 , R395_U20 , R395_U21;
wire R395_U22 , R395_U23 , R395_U24 , R395_U25 , R395_U26 , R395_U27 , R395_U28 , R395_U29 , R395_U30 , R395_U31;
wire R395_U32 , R395_U33 , R395_U34 , R395_U35 , R395_U36 , R395_U37 , R395_U38 , R395_U39 , R395_U40 , R395_U41;
wire R395_U42 , R395_U43 , R395_U44 , R395_U45 , R395_U46 , R395_U47 , R395_U48 , R395_U49 , R395_U50 , R395_U51;
wire R395_U52 , R395_U53 , R395_U54 , R395_U55 , R395_U56 , R395_U57 , R395_U58 , R395_U59 , R395_U60 , R395_U61;
wire R395_U62 , R395_U63 , R395_U64 , R395_U65 , R395_U66 , R395_U67 , R395_U68 , R395_U69 , R395_U70 , R395_U71;
wire R395_U72 , R395_U73 , R395_U74 , R395_U75 , R395_U76 , R395_U77 , R395_U78 , R395_U79 , R395_U80 , R395_U81;
wire R395_U82 , R395_U83 , R395_U84 , R395_U85 , R395_U86 , R395_U87 , R395_U88 , R395_U89 , R395_U90 , R395_U91;
wire R395_U92 , R395_U93 , R395_U94 , R395_U95 , R395_U96 , R395_U97 , R395_U98 , R395_U99 , R395_U100 , R395_U101;
wire R395_U102 , R395_U103 , R395_U104 , R395_U105 , R395_U106 , R395_U107 , R395_U108 , R395_U109 , R395_U110 , R395_U111;
wire R395_U112 , R395_U113 , R395_U114 , R395_U115 , R395_U116 , R395_U117 , R395_U118 , R395_U119 , R395_U120 , R395_U121;
wire R395_U122 , R395_U123 , R395_U124 , R395_U125 , R395_U126 , R395_U127 , R395_U128 , R395_U129 , R395_U130 , R395_U131;
wire R395_U132 , R395_U133 , R395_U134 , R395_U135 , R395_U136 , R395_U137 , R395_U138 , R395_U139 , R395_U140 , R395_U141;
wire R395_U142 , R395_U143 , R395_U144 , R395_U145 , R395_U146 , R395_U147 , R395_U148 , R395_U149 , R395_U150 , R395_U151;
wire R395_U152 , R395_U153 , R395_U154 , R395_U155 , R395_U156 , R395_U157 , R395_U158 , R395_U159 , R395_U160 , R395_U161;
wire R395_U162 , R395_U163 , R395_U164 , R395_U165 , R395_U166 , R395_U167 , R395_U168 , R395_U169 , R395_U170 , R395_U171;
wire R395_U172 , R395_U173 , R395_U174 , R395_U175 , R395_U176 , R395_U177 , R395_U178 , R395_U179 , R395_U180 , R395_U181;
wire R395_U182 , R395_U183 , R395_U184 , R395_U185 , R395_U186 , R395_U187 , R395_U188 , R1105_U4 , R1105_U5 , R1105_U6;
wire R1105_U7 , R1105_U8 , R1105_U9 , R1105_U10 , R1105_U11 , R1105_U12 , R1105_U13 , R1105_U14 , R1105_U15 , R1105_U16;
wire R1105_U17 , R1105_U18 , R1105_U19 , R1105_U20 , R1105_U21 , R1105_U22 , R1105_U23 , R1105_U24 , R1105_U25 , R1105_U26;
wire R1105_U27 , R1105_U28 , R1105_U29 , R1105_U30 , R1105_U31 , R1105_U32 , R1105_U33 , R1105_U34 , R1105_U35 , R1105_U36;
wire R1105_U37 , R1105_U38 , R1105_U39 , R1105_U40 , R1105_U41 , R1105_U42 , R1105_U43 , R1105_U44 , R1105_U45 , R1105_U46;
wire R1105_U47 , R1105_U48 , R1105_U49 , R1105_U50 , R1105_U51 , R1105_U52 , R1105_U53 , R1105_U54 , R1105_U55 , R1105_U56;
wire R1105_U57 , R1105_U58 , R1105_U59 , R1105_U60 , R1105_U61 , R1105_U62 , R1105_U63 , R1105_U64 , R1105_U65 , R1105_U66;
wire R1105_U67 , R1105_U68 , R1105_U69 , R1105_U70 , R1105_U71 , R1105_U72 , R1105_U73 , R1105_U74 , R1105_U75 , R1105_U76;
wire R1105_U77 , R1105_U78 , R1105_U79 , R1105_U80 , R1105_U81 , R1105_U82 , R1105_U83 , R1105_U84 , R1105_U85 , R1105_U86;
wire R1105_U87 , R1105_U88 , R1105_U89 , R1105_U90 , R1105_U91 , R1105_U92 , R1105_U93 , R1105_U94 , R1105_U95 , R1105_U96;
wire R1105_U97 , R1105_U98 , R1105_U99 , R1105_U100 , R1105_U101 , R1105_U102 , R1105_U103 , R1105_U104 , R1105_U105 , R1105_U106;
wire R1105_U107 , R1105_U108 , R1105_U109 , R1105_U110 , R1105_U111 , R1105_U112 , R1105_U113 , R1105_U114 , R1105_U115 , R1105_U116;
wire R1105_U117 , R1105_U118 , R1105_U119 , R1105_U120 , R1105_U121 , R1105_U122 , R1105_U123 , R1105_U124 , R1105_U125 , R1105_U126;
wire R1105_U127 , R1105_U128 , R1105_U129 , R1105_U130 , R1105_U131 , R1105_U132 , R1105_U133 , R1105_U134 , R1105_U135 , R1105_U136;
wire R1105_U137 , R1105_U138 , R1105_U139 , R1105_U140 , R1105_U141 , R1105_U142 , R1105_U143 , R1105_U144 , R1105_U145 , R1105_U146;
wire R1105_U147 , R1105_U148 , R1105_U149 , R1105_U150 , R1105_U151 , R1105_U152 , R1105_U153 , R1105_U154 , R1105_U155 , R1105_U156;
wire R1105_U157 , R1105_U158 , R1105_U159 , R1105_U160 , R1105_U161 , R1105_U162 , R1105_U163 , R1105_U164 , R1105_U165 , R1105_U166;
wire R1105_U167 , R1105_U168 , R1105_U169 , R1105_U170 , R1105_U171 , R1105_U172 , R1105_U173 , R1105_U174 , R1105_U175 , R1105_U176;
wire R1105_U177 , R1105_U178 , R1105_U179 , R1105_U180 , R1105_U181 , R1105_U182 , R1105_U183 , R1105_U184 , R1105_U185 , R1105_U186;
wire R1105_U187 , R1105_U188 , R1105_U189 , R1105_U190 , R1105_U191 , R1105_U192 , R1105_U193 , R1105_U194 , R1105_U195 , R1105_U196;
wire R1105_U197 , R1105_U198 , R1105_U199 , R1105_U200 , R1105_U201 , R1105_U202 , R1105_U203 , R1105_U204 , R1105_U205 , R1105_U206;
wire R1105_U207 , R1105_U208 , R1105_U209 , R1105_U210 , R1105_U211 , R1105_U212 , R1105_U213 , R1105_U214 , R1105_U215 , R1105_U216;
wire R1105_U217 , R1105_U218 , R1105_U219 , R1105_U220 , R1105_U221 , R1105_U222 , R1105_U223 , R1105_U224 , R1105_U225 , R1105_U226;
wire R1105_U227 , R1105_U228 , R1105_U229 , R1105_U230 , R1105_U231 , R1105_U232 , R1105_U233 , R1105_U234 , R1105_U235 , R1105_U236;
wire R1105_U237 , R1105_U238 , R1105_U239 , R1105_U240 , R1105_U241 , R1105_U242 , R1105_U243 , R1105_U244 , R1105_U245 , R1105_U246;
wire R1105_U247 , R1105_U248 , R1105_U249 , R1105_U250 , R1105_U251 , R1105_U252 , R1105_U253 , R1105_U254 , R1105_U255 , R1105_U256;
wire R1105_U257 , R1105_U258 , R1105_U259 , R1105_U260 , R1105_U261 , R1105_U262 , R1105_U263 , R1105_U264 , R1105_U265 , R1105_U266;
wire R1105_U267 , R1105_U268 , R1105_U269 , R1105_U270 , R1105_U271 , R1105_U272 , R1105_U273 , R1105_U274 , R1105_U275 , R1105_U276;
wire R1105_U277 , R1105_U278 , R1105_U279 , R1105_U280 , R1105_U281 , R1105_U282 , R1105_U283 , R1105_U284 , R1105_U285 , R1105_U286;
wire R1105_U287 , R1105_U288 , R1105_U289 , R1105_U290 , R1105_U291 , R1105_U292 , R1105_U293 , R1105_U294 , R1105_U295 , R1105_U296;
wire R1105_U297 , R1105_U298 , R1105_U299 , R1105_U300 , R1105_U301 , R1105_U302 , R1105_U303 , R1105_U304 , R1105_U305 , R1105_U306;
wire R1105_U307 , R1105_U308 , R1105_U309 , R1105_U310 , R1105_U311 , R1309_U6 , R1309_U7 , R1309_U8 , R1309_U9 , R1309_U10;
wire R1282_U6 , R1282_U7 , R1282_U8 , R1282_U9 , R1282_U10 , R1282_U11 , R1282_U12 , R1282_U13 , R1282_U14 , R1282_U15;
wire R1282_U16 , R1282_U17 , R1282_U18 , R1282_U19 , R1282_U20 , R1282_U21 , R1282_U22 , R1282_U23 , R1282_U24 , R1282_U25;
wire R1282_U26 , R1282_U27 , R1282_U28 , R1282_U29 , R1282_U30 , R1282_U31 , R1282_U32 , R1282_U33 , R1282_U34 , R1282_U35;
wire R1282_U36 , R1282_U37 , R1282_U38 , R1282_U39 , R1282_U40 , R1282_U41 , R1282_U42 , R1282_U43 , R1282_U44 , R1282_U45;
wire R1282_U46 , R1282_U47 , R1282_U48 , R1282_U49 , R1282_U50 , R1282_U51 , R1282_U52 , R1282_U53 , R1282_U54 , R1282_U55;
wire R1282_U56 , R1282_U57 , R1282_U58 , R1282_U59 , R1282_U60 , R1282_U61 , R1282_U62 , R1282_U63 , R1282_U64 , R1282_U65;
wire R1282_U66 , R1282_U67 , R1282_U68 , R1282_U69 , R1282_U70 , R1282_U71 , R1282_U72 , R1282_U73 , R1282_U74 , R1282_U75;
wire R1282_U76 , R1282_U77 , R1282_U78 , R1282_U79 , R1282_U80 , R1282_U81 , R1282_U82 , R1282_U83 , R1282_U84 , R1282_U85;
wire R1282_U86 , R1282_U87 , R1282_U88 , R1282_U89 , R1282_U90 , R1282_U91 , R1282_U92 , R1282_U93 , R1282_U94 , R1282_U95;
wire R1282_U96 , R1282_U97 , R1282_U98 , R1282_U99 , R1282_U100 , R1282_U101 , R1282_U102 , R1282_U103 , R1282_U104 , R1282_U105;
wire R1282_U106 , R1282_U107 , R1282_U108 , R1282_U109 , R1282_U110 , R1282_U111 , R1282_U112 , R1282_U113 , R1282_U114 , R1282_U115;
wire R1282_U116 , R1282_U117 , R1282_U118 , R1282_U119 , R1282_U120 , R1282_U121 , R1282_U122 , R1282_U123 , R1282_U124 , R1282_U125;
wire R1282_U126 , R1282_U127 , R1282_U128 , R1282_U129 , R1282_U130 , R1282_U131 , R1282_U132 , R1282_U133 , R1282_U134 , R1282_U135;
wire R1282_U136 , R1282_U137 , R1282_U138 , R1282_U139 , R1282_U140 , R1282_U141 , R1282_U142 , R1282_U143 , R1282_U144 , R1282_U145;
wire R1282_U146 , R1282_U147 , R1282_U148 , R1282_U149 , R1282_U150 , R1282_U151 , R1282_U152 , R1282_U153 , R1282_U154 , R1282_U155;
wire R1282_U156 , R1282_U157 , R1282_U158 , R1282_U159 , R1282_U160 , R1282_U161 , R1282_U162 , R1282_U163 , R1282_U164 , R1282_U165;
wire R1282_U166 , R1282_U167 , R1282_U168 , R1282_U169 , R1282_U170 , R1282_U171 , R1282_U172 , R1282_U173 , R1282_U174 , R1282_U175;
wire R1282_U176 , R1282_U177 , R1282_U178 , R1282_U179 , R1282_U180 , R1240_U4 , R1240_U5 , R1240_U6 , R1240_U7 , R1240_U8;
wire R1240_U9 , R1240_U10 , R1240_U11 , R1240_U12 , R1240_U13 , R1240_U14 , R1240_U15 , R1240_U16 , R1240_U17 , R1240_U18;
wire R1240_U19 , R1240_U20 , R1240_U21 , R1240_U22 , R1240_U23 , R1240_U24 , R1240_U25 , R1240_U26 , R1240_U27 , R1240_U28;
wire R1240_U29 , R1240_U30 , R1240_U31 , R1240_U32 , R1240_U33 , R1240_U34 , R1240_U35 , R1240_U36 , R1240_U37 , R1240_U38;
wire R1240_U39 , R1240_U40 , R1240_U41 , R1240_U42 , R1240_U43 , R1240_U44 , R1240_U45 , R1240_U46 , R1240_U47 , R1240_U48;
wire R1240_U49 , R1240_U50 , R1240_U51 , R1240_U52 , R1240_U53 , R1240_U54 , R1240_U55 , R1240_U56 , R1240_U57 , R1240_U58;
wire R1240_U59 , R1240_U60 , R1240_U61 , R1240_U62 , R1240_U63 , R1240_U64 , R1240_U65 , R1240_U66 , R1240_U67 , R1240_U68;
wire R1240_U69 , R1240_U70 , R1240_U71 , R1240_U72 , R1240_U73 , R1240_U74 , R1240_U75 , R1240_U76 , R1240_U77 , R1240_U78;
wire R1240_U79 , R1240_U80 , R1240_U81 , R1240_U82 , R1240_U83 , R1240_U84 , R1240_U85 , R1240_U86 , R1240_U87 , R1240_U88;
wire R1240_U89 , R1240_U90 , R1240_U91 , R1240_U92 , R1240_U93 , R1240_U94 , R1240_U95 , R1240_U96 , R1240_U97 , R1240_U98;
wire R1240_U99 , R1240_U100 , R1240_U101 , R1240_U102 , R1240_U103 , R1240_U104 , R1240_U105 , R1240_U106 , R1240_U107 , R1240_U108;
wire R1240_U109 , R1240_U110 , R1240_U111 , R1240_U112 , R1240_U113 , R1240_U114 , R1240_U115 , R1240_U116 , R1240_U117 , R1240_U118;
wire R1240_U119 , R1240_U120 , R1240_U121 , R1240_U122 , R1240_U123 , R1240_U124 , R1240_U125 , R1240_U126 , R1240_U127 , R1240_U128;
wire R1240_U129 , R1240_U130 , R1240_U131 , R1240_U132 , R1240_U133 , R1240_U134 , R1240_U135 , R1240_U136 , R1240_U137 , R1240_U138;
wire R1240_U139 , R1240_U140 , R1240_U141 , R1240_U142 , R1240_U143 , R1240_U144 , R1240_U145 , R1240_U146 , R1240_U147 , R1240_U148;
wire R1240_U149 , R1240_U150 , R1240_U151 , R1240_U152 , R1240_U153 , R1240_U154 , R1240_U155 , R1240_U156 , R1240_U157 , R1240_U158;
wire R1240_U159 , R1240_U160 , R1240_U161 , R1240_U162 , R1240_U163 , R1240_U164 , R1240_U165 , R1240_U166 , R1240_U167 , R1240_U168;
wire R1240_U169 , R1240_U170 , R1240_U171 , R1240_U172 , R1240_U173 , R1240_U174 , R1240_U175 , R1240_U176 , R1240_U177 , R1240_U178;
wire R1240_U179 , R1240_U180 , R1240_U181 , R1240_U182 , R1240_U183 , R1240_U184 , R1240_U185 , R1240_U186 , R1240_U187 , R1240_U188;
wire R1240_U189 , R1240_U190 , R1240_U191 , R1240_U192 , R1240_U193 , R1240_U194 , R1240_U195 , R1240_U196 , R1240_U197 , R1240_U198;
wire R1240_U199 , R1240_U200 , R1240_U201 , R1240_U202 , R1240_U203 , R1240_U204 , R1240_U205 , R1240_U206 , R1240_U207 , R1240_U208;
wire R1240_U209 , R1240_U210 , R1240_U211 , R1240_U212 , R1240_U213 , R1240_U214 , R1240_U215 , R1240_U216 , R1240_U217 , R1240_U218;
wire R1240_U219 , R1240_U220 , R1240_U221 , R1240_U222 , R1240_U223 , R1240_U224 , R1240_U225 , R1240_U226 , R1240_U227 , R1240_U228;
wire R1240_U229 , R1240_U230 , R1240_U231 , R1240_U232 , R1240_U233 , R1240_U234 , R1240_U235 , R1240_U236 , R1240_U237 , R1240_U238;
wire R1240_U239 , R1240_U240 , R1240_U241 , R1240_U242 , R1240_U243 , R1240_U244 , R1240_U245 , R1240_U246 , R1240_U247 , R1240_U248;
wire R1240_U249 , R1240_U250 , R1240_U251 , R1240_U252 , R1240_U253 , R1240_U254 , R1240_U255 , R1240_U256 , R1240_U257 , R1240_U258;
wire R1240_U259 , R1240_U260 , R1240_U261 , R1240_U262 , R1240_U263 , R1240_U264 , R1240_U265 , R1240_U266 , R1240_U267 , R1240_U268;
wire R1240_U269 , R1240_U270 , R1240_U271 , R1240_U272 , R1240_U273 , R1240_U274 , R1240_U275 , R1240_U276 , R1240_U277 , R1240_U278;
wire R1240_U279 , R1240_U280 , R1240_U281 , R1240_U282 , R1240_U283 , R1240_U284 , R1240_U285 , R1240_U286 , R1240_U287 , R1240_U288;
wire R1240_U289 , R1240_U290 , R1240_U291 , R1240_U292 , R1240_U293 , R1240_U294 , R1240_U295 , R1240_U296 , R1240_U297 , R1240_U298;
wire R1240_U299 , R1240_U300 , R1240_U301 , R1240_U302 , R1240_U303 , R1240_U304 , R1240_U305 , R1240_U306 , R1240_U307 , R1240_U308;
wire R1240_U309 , R1240_U310 , R1240_U311 , R1240_U312 , R1240_U313 , R1240_U314 , R1240_U315 , R1240_U316 , R1240_U317 , R1240_U318;
wire R1240_U319 , R1240_U320 , R1240_U321 , R1240_U322 , R1240_U323 , R1240_U324 , R1240_U325 , R1240_U326 , R1240_U327 , R1240_U328;
wire R1240_U329 , R1240_U330 , R1240_U331 , R1240_U332 , R1240_U333 , R1240_U334 , R1240_U335 , R1240_U336 , R1240_U337 , R1240_U338;
wire R1240_U339 , R1240_U340 , R1240_U341 , R1240_U342 , R1240_U343 , R1240_U344 , R1240_U345 , R1240_U346 , R1240_U347 , R1240_U348;
wire R1240_U349 , R1240_U350 , R1240_U351 , R1240_U352 , R1240_U353 , R1240_U354 , R1240_U355 , R1240_U356 , R1240_U357 , R1240_U358;
wire R1240_U359 , R1240_U360 , R1240_U361 , R1240_U362 , R1240_U363 , R1240_U364 , R1240_U365 , R1240_U366 , R1240_U367 , R1240_U368;
wire R1240_U369 , R1240_U370 , R1240_U371 , R1240_U372 , R1240_U373 , R1240_U374 , R1240_U375 , R1240_U376 , R1240_U377 , R1240_U378;
wire R1240_U379 , R1240_U380 , R1240_U381 , R1240_U382 , R1240_U383 , R1240_U384 , R1240_U385 , R1240_U386 , R1240_U387 , R1240_U388;
wire R1240_U389 , R1240_U390 , R1240_U391 , R1240_U392 , R1240_U393 , R1240_U394 , R1240_U395 , R1240_U396 , R1240_U397 , R1240_U398;
wire R1240_U399 , R1240_U400 , R1240_U401 , R1240_U402 , R1240_U403 , R1240_U404 , R1240_U405 , R1240_U406 , R1240_U407 , R1240_U408;
wire R1240_U409 , R1240_U410 , R1240_U411 , R1240_U412 , R1240_U413 , R1240_U414 , R1240_U415 , R1240_U416 , R1240_U417 , R1240_U418;
wire R1240_U419 , R1240_U420 , R1240_U421 , R1240_U422 , R1240_U423 , R1240_U424 , R1240_U425 , R1240_U426 , R1240_U427 , R1240_U428;
wire R1240_U429 , R1240_U430 , R1240_U431 , R1240_U432 , R1240_U433 , R1240_U434 , R1240_U435 , R1240_U436 , R1240_U437 , R1240_U438;
wire R1240_U439 , R1240_U440 , R1240_U441 , R1240_U442 , R1240_U443 , R1240_U444 , R1240_U445 , R1240_U446 , R1240_U447 , R1240_U448;
wire R1240_U449 , R1240_U450 , R1240_U451 , R1240_U452 , R1240_U453 , R1240_U454 , R1240_U455 , R1240_U456 , R1240_U457 , R1240_U458;
wire R1240_U459 , R1240_U460 , R1240_U461 , R1240_U462 , R1240_U463 , R1240_U464 , R1240_U465 , R1240_U466 , R1240_U467 , R1240_U468;
wire R1240_U469 , R1240_U470 , R1240_U471 , R1240_U472 , R1240_U473 , R1240_U474 , R1240_U475 , R1240_U476 , R1240_U477 , R1240_U478;
wire R1240_U479 , R1240_U480 , R1240_U481 , R1240_U482 , R1240_U483 , R1240_U484 , R1240_U485 , R1240_U486 , R1240_U487 , R1240_U488;
wire R1240_U489 , R1240_U490 , R1240_U491 , R1240_U492 , R1240_U493 , R1240_U494 , R1240_U495 , R1240_U496 , R1240_U497 , R1240_U498;
wire R1240_U499 , R1240_U500 , R1240_U501 , R1240_U502 , R1240_U503 , R1240_U504 , R1240_U505 , R1240_U506 , R1240_U507 , R1240_U508;
wire R1240_U509 , R1240_U510 , R1240_U511 , R1240_U512 , R1240_U513 , R1240_U514 , R1240_U515 , R1240_U516 , R1240_U517 , R1240_U518;
wire R1240_U519 , R1240_U520 , R1240_U521 , R1240_U522 , R1240_U523 , R1240_U524 , R1240_U525 , R1240_U526 , R1240_U527 , R1240_U528;
wire R1240_U529 , R1240_U530 , R1240_U531 , R1162_U4 , R1162_U5 , R1162_U6 , R1162_U7 , R1162_U8 , R1162_U9 , R1162_U10;
wire R1162_U11 , R1162_U12 , R1162_U13 , R1162_U14 , R1162_U15 , R1162_U16 , R1162_U17 , R1162_U18 , R1162_U19 , R1162_U20;
wire R1162_U21 , R1162_U22 , R1162_U23 , R1162_U24 , R1162_U25 , R1162_U26 , R1162_U27 , R1162_U28 , R1162_U29 , R1162_U30;
wire R1162_U31 , R1162_U32 , R1162_U33 , R1162_U34 , R1162_U35 , R1162_U36 , R1162_U37 , R1162_U38 , R1162_U39 , R1162_U40;
wire R1162_U41 , R1162_U42 , R1162_U43 , R1162_U44 , R1162_U45 , R1162_U46 , R1162_U47 , R1162_U48 , R1162_U49 , R1162_U50;
wire R1162_U51 , R1162_U52 , R1162_U53 , R1162_U54 , R1162_U55 , R1162_U56 , R1162_U57 , R1162_U58 , R1162_U59 , R1162_U60;
wire R1162_U61 , R1162_U62 , R1162_U63 , R1162_U64 , R1162_U65 , R1162_U66 , R1162_U67 , R1162_U68 , R1162_U69 , R1162_U70;
wire R1162_U71 , R1162_U72 , R1162_U73 , R1162_U74 , R1162_U75 , R1162_U76 , R1162_U77 , R1162_U78 , R1162_U79 , R1162_U80;
wire R1162_U81 , R1162_U82 , R1162_U83 , R1162_U84 , R1162_U85 , R1162_U86 , R1162_U87 , R1162_U88 , R1162_U89 , R1162_U90;
wire R1162_U91 , R1162_U92 , R1162_U93 , R1162_U94 , R1162_U95 , R1162_U96 , R1162_U97 , R1162_U98 , R1162_U99 , R1162_U100;
wire R1162_U101 , R1162_U102 , R1162_U103 , R1162_U104 , R1162_U105 , R1162_U106 , R1162_U107 , R1162_U108 , R1162_U109 , R1162_U110;
wire R1162_U111 , R1162_U112 , R1162_U113 , R1162_U114 , R1162_U115 , R1162_U116 , R1162_U117 , R1162_U118 , R1162_U119 , R1162_U120;
wire R1162_U121 , R1162_U122 , R1162_U123 , R1162_U124 , R1162_U125 , R1162_U126 , R1162_U127 , R1162_U128 , R1162_U129 , R1162_U130;
wire R1162_U131 , R1162_U132 , R1162_U133 , R1162_U134 , R1162_U135 , R1162_U136 , R1162_U137 , R1162_U138 , R1162_U139 , R1162_U140;
wire R1162_U141 , R1162_U142 , R1162_U143 , R1162_U144 , R1162_U145 , R1162_U146 , R1162_U147 , R1162_U148 , R1162_U149 , R1162_U150;
wire R1162_U151 , R1162_U152 , R1162_U153 , R1162_U154 , R1162_U155 , R1162_U156 , R1162_U157 , R1162_U158 , R1162_U159 , R1162_U160;
wire R1162_U161 , R1162_U162 , R1162_U163 , R1162_U164 , R1162_U165 , R1162_U166 , R1162_U167 , R1162_U168 , R1162_U169 , R1162_U170;
wire R1162_U171 , R1162_U172 , R1162_U173 , R1162_U174 , R1162_U175 , R1162_U176 , R1162_U177 , R1162_U178 , R1162_U179 , R1162_U180;
wire R1162_U181 , R1162_U182 , R1162_U183 , R1162_U184 , R1162_U185 , R1162_U186 , R1162_U187 , R1162_U188 , R1162_U189 , R1162_U190;
wire R1162_U191 , R1162_U192 , R1162_U193 , R1162_U194 , R1162_U195 , R1162_U196 , R1162_U197 , R1162_U198 , R1162_U199 , R1162_U200;
wire R1162_U201 , R1162_U202 , R1162_U203 , R1162_U204 , R1162_U205 , R1162_U206 , R1162_U207 , R1162_U208 , R1162_U209 , R1162_U210;
wire R1162_U211 , R1162_U212 , R1162_U213 , R1162_U214 , R1162_U215 , R1162_U216 , R1162_U217 , R1162_U218 , R1162_U219 , R1162_U220;
wire R1162_U221 , R1162_U222 , R1162_U223 , R1162_U224 , R1162_U225 , R1162_U226 , R1162_U227 , R1162_U228 , R1162_U229 , R1162_U230;
wire R1162_U231 , R1162_U232 , R1162_U233 , R1162_U234 , R1162_U235 , R1162_U236 , R1162_U237 , R1162_U238 , R1162_U239 , R1162_U240;
wire R1162_U241 , R1162_U242 , R1162_U243 , R1162_U244 , R1162_U245 , R1162_U246 , R1162_U247 , R1162_U248 , R1162_U249 , R1162_U250;
wire R1162_U251 , R1162_U252 , R1162_U253 , R1162_U254 , R1162_U255 , R1162_U256 , R1162_U257 , R1162_U258 , R1162_U259 , R1162_U260;
wire R1162_U261 , R1162_U262 , R1162_U263 , R1162_U264 , R1162_U265 , R1162_U266 , R1162_U267 , R1162_U268 , R1162_U269 , R1162_U270;
wire R1162_U271 , R1162_U272 , R1162_U273 , R1162_U274 , R1162_U275 , R1162_U276 , R1162_U277 , R1162_U278 , R1162_U279 , R1162_U280;
wire R1162_U281 , R1162_U282 , R1162_U283 , R1162_U284 , R1162_U285 , R1162_U286 , R1162_U287 , R1162_U288 , R1162_U289 , R1162_U290;
wire R1117_U6 , R1117_U7 , R1117_U8 , R1117_U9 , R1117_U10 , R1117_U11 , R1117_U12 , R1117_U13 , R1117_U14 , R1117_U15;
wire R1117_U16 , R1117_U17 , R1117_U18 , R1117_U19 , R1117_U20 , R1117_U21 , R1117_U22 , R1117_U23 , R1117_U24 , R1117_U25;
wire R1117_U26 , R1117_U27 , R1117_U28 , R1117_U29 , R1117_U30 , R1117_U31 , R1117_U32 , R1117_U33 , R1117_U34 , R1117_U35;
wire R1117_U36 , R1117_U37 , R1117_U38 , R1117_U39 , R1117_U40 , R1117_U41 , R1117_U42 , R1117_U43 , R1117_U44 , R1117_U45;
wire R1117_U46 , R1117_U47 , R1117_U48 , R1117_U49 , R1117_U50 , R1117_U51 , R1117_U52 , R1117_U53 , R1117_U54 , R1117_U55;
wire R1117_U56 , R1117_U57 , R1117_U58 , R1117_U59 , R1117_U60 , R1117_U61 , R1117_U62 , R1117_U63 , R1117_U64 , R1117_U65;
wire R1117_U66 , R1117_U67 , R1117_U68 , R1117_U69 , R1117_U70 , R1117_U71 , R1117_U72 , R1117_U73 , R1117_U74 , R1117_U75;
wire R1117_U76 , R1117_U77 , R1117_U78 , R1117_U79 , R1117_U80 , R1117_U81 , R1117_U82 , R1117_U83 , R1117_U84 , R1117_U85;
wire R1117_U86 , R1117_U87 , R1117_U88 , R1117_U89 , R1117_U90 , R1117_U91 , R1117_U92 , R1117_U93 , R1117_U94 , R1117_U95;
wire R1117_U96 , R1117_U97 , R1117_U98 , R1117_U99 , R1117_U100 , R1117_U101 , R1117_U102 , R1117_U103 , R1117_U104 , R1117_U105;
wire R1117_U106 , R1117_U107 , R1117_U108 , R1117_U109 , R1117_U110 , R1117_U111 , R1117_U112 , R1117_U113 , R1117_U114 , R1117_U115;
wire R1117_U116 , R1117_U117 , R1117_U118 , R1117_U119 , R1117_U120 , R1117_U121 , R1117_U122 , R1117_U123 , R1117_U124 , R1117_U125;
wire R1117_U126 , R1117_U127 , R1117_U128 , R1117_U129 , R1117_U130 , R1117_U131 , R1117_U132 , R1117_U133 , R1117_U134 , R1117_U135;
wire R1117_U136 , R1117_U137 , R1117_U138 , R1117_U139 , R1117_U140 , R1117_U141 , R1117_U142 , R1117_U143 , R1117_U144 , R1117_U145;
wire R1117_U146 , R1117_U147 , R1117_U148 , R1117_U149 , R1117_U150 , R1117_U151 , R1117_U152 , R1117_U153 , R1117_U154 , R1117_U155;
wire R1117_U156 , R1117_U157 , R1117_U158 , R1117_U159 , R1117_U160 , R1117_U161 , R1117_U162 , R1117_U163 , R1117_U164 , R1117_U165;
wire R1117_U166 , R1117_U167 , R1117_U168 , R1117_U169 , R1117_U170 , R1117_U171 , R1117_U172 , R1117_U173 , R1117_U174 , R1117_U175;
wire R1117_U176 , R1117_U177 , R1117_U178 , R1117_U179 , R1117_U180 , R1117_U181 , R1117_U182 , R1117_U183 , R1117_U184 , R1117_U185;
wire R1117_U186 , R1117_U187 , R1117_U188 , R1117_U189 , R1117_U190 , R1117_U191 , R1117_U192 , R1117_U193 , R1117_U194 , R1117_U195;
wire R1117_U196 , R1117_U197 , R1117_U198 , R1117_U199 , R1117_U200 , R1117_U201 , R1117_U202 , R1117_U203 , R1117_U204 , R1117_U205;
wire R1117_U206 , R1117_U207 , R1117_U208 , R1117_U209 , R1117_U210 , R1117_U211 , R1117_U212 , R1117_U213 , R1117_U214 , R1117_U215;
wire R1117_U216 , R1117_U217 , R1117_U218 , R1117_U219 , R1117_U220 , R1117_U221 , R1117_U222 , R1117_U223 , R1117_U224 , R1117_U225;
wire R1117_U226 , R1117_U227 , R1117_U228 , R1117_U229 , R1117_U230 , R1117_U231 , R1117_U232 , R1117_U233 , R1117_U234 , R1117_U235;
wire R1117_U236 , R1117_U237 , R1117_U238 , R1117_U239 , R1117_U240 , R1117_U241 , R1117_U242 , R1117_U243 , R1117_U244 , R1117_U245;
wire R1117_U246 , R1117_U247 , R1117_U248 , R1117_U249 , R1117_U250 , R1117_U251 , R1117_U252 , R1117_U253 , R1117_U254 , R1117_U255;
wire R1117_U256 , R1117_U257 , R1117_U258 , R1117_U259 , R1117_U260 , R1117_U261 , R1117_U262 , R1117_U263 , R1117_U264 , R1117_U265;
wire R1117_U266 , R1117_U267 , R1117_U268 , R1117_U269 , R1117_U270 , R1117_U271 , R1117_U272 , R1117_U273 , R1117_U274 , R1117_U275;
wire R1117_U276 , R1117_U277 , R1117_U278 , R1117_U279 , R1117_U280 , R1117_U281 , R1117_U282 , R1117_U283 , R1117_U284 , R1117_U285;
wire R1117_U286 , R1117_U287 , R1117_U288 , R1117_U289 , R1117_U290 , R1117_U291 , R1117_U292 , R1117_U293 , R1117_U294 , R1117_U295;
wire R1117_U296 , R1117_U297 , R1117_U298 , R1117_U299 , R1117_U300 , R1117_U301 , R1117_U302 , R1117_U303 , R1117_U304 , R1117_U305;
wire R1117_U306 , R1117_U307 , R1117_U308 , R1117_U309 , R1117_U310 , R1117_U311 , R1117_U312 , R1117_U313 , R1117_U314 , R1117_U315;
wire R1117_U316 , R1117_U317 , R1117_U318 , R1117_U319 , R1117_U320 , R1117_U321 , R1117_U322 , R1117_U323 , R1117_U324 , R1117_U325;
wire R1117_U326 , R1117_U327 , R1117_U328 , R1117_U329 , R1117_U330 , R1117_U331 , R1117_U332 , R1117_U333 , R1117_U334 , R1117_U335;
wire R1117_U336 , R1117_U337 , R1117_U338 , R1117_U339 , R1117_U340 , R1117_U341 , R1117_U342 , R1117_U343 , R1117_U344 , R1117_U345;
wire R1117_U346 , R1117_U347 , R1117_U348 , R1117_U349 , R1117_U350 , R1117_U351 , R1117_U352 , R1117_U353 , R1117_U354 , R1117_U355;
wire R1117_U356 , R1117_U357 , R1117_U358 , R1117_U359 , R1117_U360 , R1117_U361 , R1117_U362 , R1117_U363 , R1117_U364 , R1117_U365;
wire R1117_U366 , R1117_U367 , R1117_U368 , R1117_U369 , R1117_U370 , R1117_U371 , R1117_U372 , R1117_U373 , R1117_U374 , R1117_U375;
wire R1117_U376 , R1117_U377 , R1117_U378 , R1117_U379 , R1117_U380 , R1117_U381 , R1117_U382 , R1117_U383 , R1117_U384 , R1117_U385;
wire R1117_U386 , R1117_U387 , R1117_U388 , R1117_U389 , R1117_U390 , R1117_U391 , R1117_U392 , R1117_U393 , R1117_U394 , R1117_U395;
wire R1117_U396 , R1117_U397 , R1117_U398 , R1117_U399 , R1117_U400 , R1117_U401 , R1117_U402 , R1117_U403 , R1117_U404 , R1117_U405;
wire R1117_U406 , R1117_U407 , R1117_U408 , R1117_U409 , R1117_U410 , R1117_U411 , R1117_U412 , R1117_U413 , R1117_U414 , R1117_U415;
wire R1117_U416 , R1117_U417 , R1117_U418 , R1117_U419 , R1117_U420 , R1117_U421 , R1117_U422 , R1117_U423 , R1117_U424 , R1117_U425;
wire R1117_U426 , R1117_U427 , R1117_U428 , R1117_U429 , R1117_U430 , R1117_U431 , R1117_U432 , R1117_U433 , R1117_U434 , R1117_U435;
wire R1117_U436 , R1117_U437 , R1117_U438 , R1117_U439 , R1117_U440 , R1117_U441 , R1117_U442 , R1117_U443 , R1117_U444 , R1117_U445;
wire R1117_U446 , R1117_U447 , R1117_U448 , R1117_U449 , R1117_U450 , R1117_U451 , R1117_U452 , R1117_U453 , R1117_U454 , R1117_U455;
wire R1117_U456 , R1117_U457 , R1117_U458 , R1117_U459 , R1117_U460 , R1117_U461 , R1117_U462 , R1117_U463 , R1117_U464 , R1117_U465;
wire R1117_U466 , R1117_U467 , R1117_U468 , R1117_U469 , R1117_U470 , R1117_U471 , R1117_U472 , R1117_U473 , R1117_U474 , R1117_U475;
wire R1117_U476 , R1117_U477 , R1117_U478 , R1117_U479 , R1117_U480 , R1117_U481 , R1117_U482 , R1117_U483 , R1117_U484 , R1117_U485;
wire R1117_U486 , R1117_U487 , R1117_U488 , R1117_U489 , R1117_U490 , R1117_U491 , R1117_U492 , R1117_U493 , R1117_U494 , R1117_U495;
wire R1117_U496 , R1117_U497 , R1117_U498 , R1117_U499 , R1117_U500 , R1117_U501 , R1117_U502 , R1117_U503 , R1117_U504 , R1117_U505;
wire R1117_U506 , R1117_U507 , R1117_U508 , R1117_U509 , R1117_U510 , R1117_U511 , R1117_U512 , R1117_U513 , R1117_U514 , R1117_U515;
wire R1375_U6 , R1375_U7 , R1375_U8 , R1375_U9 , R1375_U10 , R1375_U11 , R1375_U12 , R1375_U13 , R1375_U14 , R1375_U15;
wire R1375_U16 , R1375_U17 , R1375_U18 , R1375_U19 , R1375_U20 , R1375_U21 , R1375_U22 , R1375_U23 , R1375_U24 , R1375_U25;
wire R1375_U26 , R1375_U27 , R1375_U28 , R1375_U29 , R1375_U30 , R1375_U31 , R1375_U32 , R1375_U33 , R1375_U34 , R1375_U35;
wire R1375_U36 , R1375_U37 , R1375_U38 , R1375_U39 , R1375_U40 , R1375_U41 , R1375_U42 , R1375_U43 , R1375_U44 , R1375_U45;
wire R1375_U46 , R1375_U47 , R1375_U48 , R1375_U49 , R1375_U50 , R1375_U51 , R1375_U52 , R1375_U53 , R1375_U54 , R1375_U55;
wire R1375_U56 , R1375_U57 , R1375_U58 , R1375_U59 , R1375_U60 , R1375_U61 , R1375_U62 , R1375_U63 , R1375_U64 , R1375_U65;
wire R1375_U66 , R1375_U67 , R1375_U68 , R1375_U69 , R1375_U70 , R1375_U71 , R1375_U72 , R1375_U73 , R1375_U74 , R1375_U75;
wire R1375_U76 , R1375_U77 , R1375_U78 , R1375_U79 , R1375_U80 , R1375_U81 , R1375_U82 , R1375_U83 , R1375_U84 , R1375_U85;
wire R1375_U86 , R1375_U87 , R1375_U88 , R1375_U89 , R1375_U90 , R1375_U91 , R1375_U92 , R1375_U93 , R1375_U94 , R1375_U95;
wire R1375_U96 , R1375_U97 , R1375_U98 , R1375_U99 , R1375_U100 , R1375_U101 , R1375_U102 , R1375_U103 , R1375_U104 , R1375_U105;
wire R1375_U106 , R1375_U107 , R1375_U108 , R1375_U109 , R1375_U110 , R1375_U111 , R1375_U112 , R1375_U113 , R1375_U114 , R1375_U115;
wire R1375_U116 , R1375_U117 , R1375_U118 , R1375_U119 , R1375_U120 , R1375_U121 , R1375_U122 , R1375_U123 , R1375_U124 , R1375_U125;
wire R1375_U126 , R1375_U127 , R1375_U128 , R1375_U129 , R1375_U130 , R1375_U131 , R1375_U132 , R1375_U133 , R1375_U134 , R1375_U135;
wire R1375_U136 , R1375_U137 , R1375_U138 , R1375_U139 , R1375_U140 , R1375_U141 , R1375_U142 , R1375_U143 , R1375_U144 , R1375_U145;
wire R1375_U146 , R1375_U147 , R1375_U148 , R1375_U149 , R1375_U150 , R1375_U151 , R1375_U152 , R1375_U153 , R1375_U154 , R1375_U155;
wire R1375_U156 , R1375_U157 , R1375_U158 , R1375_U159 , R1375_U160 , R1375_U161 , R1375_U162 , R1375_U163 , R1375_U164 , R1375_U165;
wire R1375_U166 , R1375_U167 , R1375_U168 , R1375_U169 , R1375_U170 , R1375_U171 , R1375_U172 , R1375_U173 , R1375_U174 , R1375_U175;
wire R1375_U176 , R1375_U177 , R1375_U178 , R1375_U179 , R1375_U180 , R1375_U181 , R1375_U182 , R1375_U183 , R1375_U184 , R1375_U185;
wire R1375_U186 , R1375_U187 , R1375_U188 , R1375_U189 , R1375_U190 , R1375_U191 , R1375_U192 , R1375_U193 , R1375_U194 , R1375_U195;
wire R1375_U196 , R1375_U197 , R1375_U198 , R1375_U199 , R1375_U200 , R1375_U201 , R1375_U202 , R1375_U203 , R1375_U204 , R1375_U205;
wire R1375_U206 , R1375_U207 , R1375_U208 , R1375_U209 , R1375_U210 , R1375_U211 , R1375_U212 , R1375_U213 , R1375_U214 , R1375_U215;
wire R1375_U216 , R1375_U217 , R1375_U218 , R1375_U219 , R1375_U220 , R1375_U221 , R1375_U222 , R1375_U223 , R1375_U224 , R1375_U225;
wire R1352_U6 , R1352_U7 , R1207_U6 , R1207_U7 , R1207_U8 , R1207_U9 , R1207_U10 , R1207_U11 , R1207_U12 , R1207_U13;
wire R1207_U14 , R1207_U15 , R1207_U16 , R1207_U17 , R1207_U18 , R1207_U19 , R1207_U20 , R1207_U21 , R1207_U22 , R1207_U23;
wire R1207_U24 , R1207_U25 , R1207_U26 , R1207_U27 , R1207_U28 , R1207_U29 , R1207_U30 , R1207_U31 , R1207_U32 , R1207_U33;
wire R1207_U34 , R1207_U35 , R1207_U36 , R1207_U37 , R1207_U38 , R1207_U39 , R1207_U40 , R1207_U41 , R1207_U42 , R1207_U43;
wire R1207_U44 , R1207_U45 , R1207_U46 , R1207_U47 , R1207_U48 , R1207_U49 , R1207_U50 , R1207_U51 , R1207_U52 , R1207_U53;
wire R1207_U54 , R1207_U55 , R1207_U56 , R1207_U57 , R1207_U58 , R1207_U59 , R1207_U60 , R1207_U61 , R1207_U62 , R1207_U63;
wire R1207_U64 , R1207_U65 , R1207_U66 , R1207_U67 , R1207_U68 , R1207_U69 , R1207_U70 , R1207_U71 , R1207_U72 , R1207_U73;
wire R1207_U74 , R1207_U75 , R1207_U76 , R1207_U77 , R1207_U78 , R1207_U79 , R1207_U80 , R1207_U81 , R1207_U82 , R1207_U83;
wire R1207_U84 , R1207_U85 , R1207_U86 , R1207_U87 , R1207_U88 , R1207_U89 , R1207_U90 , R1207_U91 , R1207_U92 , R1207_U93;
wire R1207_U94 , R1207_U95 , R1207_U96 , R1207_U97 , R1207_U98 , R1207_U99 , R1207_U100 , R1207_U101 , R1207_U102 , R1207_U103;
wire R1207_U104 , R1207_U105 , R1207_U106 , R1207_U107 , R1207_U108 , R1207_U109 , R1207_U110 , R1207_U111 , R1207_U112 , R1207_U113;
wire R1207_U114 , R1207_U115 , R1207_U116 , R1207_U117 , R1207_U118 , R1207_U119 , R1207_U120 , R1207_U121 , R1207_U122 , R1207_U123;
wire R1207_U124 , R1207_U125 , R1207_U126 , R1207_U127 , R1207_U128 , R1207_U129 , R1207_U130 , R1207_U131 , R1207_U132 , R1207_U133;
wire R1207_U134 , R1207_U135 , R1207_U136 , R1207_U137 , R1207_U138 , R1207_U139 , R1207_U140 , R1207_U141 , R1207_U142 , R1207_U143;
wire R1207_U144 , R1207_U145 , R1207_U146 , R1207_U147 , R1207_U148 , R1207_U149 , R1207_U150 , R1207_U151 , R1207_U152 , R1207_U153;
wire R1207_U154 , R1207_U155 , R1207_U156 , R1207_U157 , R1207_U158 , R1207_U159 , R1207_U160 , R1207_U161 , R1207_U162 , R1207_U163;
wire R1207_U164 , R1207_U165 , R1207_U166 , R1207_U167 , R1207_U168 , R1207_U169 , R1207_U170 , R1207_U171 , R1207_U172 , R1207_U173;
wire R1207_U174 , R1207_U175 , R1207_U176 , R1207_U177 , R1207_U178 , R1207_U179 , R1207_U180 , R1207_U181 , R1207_U182 , R1207_U183;
wire R1207_U184 , R1207_U185 , R1207_U186 , R1207_U187 , R1207_U188 , R1207_U189 , R1207_U190 , R1207_U191 , R1207_U192 , R1207_U193;
wire R1207_U194 , R1207_U195 , R1207_U196 , R1207_U197 , R1207_U198 , R1207_U199 , R1207_U200 , R1207_U201 , R1207_U202 , R1207_U203;
wire R1207_U204 , R1207_U205 , R1207_U206 , R1207_U207 , R1207_U208 , R1207_U209 , R1207_U210 , R1207_U211 , R1207_U212 , R1207_U213;
wire R1207_U214 , R1207_U215 , R1207_U216 , R1207_U217 , R1207_U218 , R1207_U219 , R1207_U220 , R1207_U221 , R1207_U222 , R1207_U223;
wire R1207_U224 , R1207_U225 , R1207_U226 , R1207_U227 , R1207_U228 , R1207_U229 , R1207_U230 , R1207_U231 , R1207_U232 , R1207_U233;
wire R1207_U234 , R1207_U235 , R1207_U236 , R1207_U237 , R1207_U238 , R1207_U239 , R1207_U240 , R1207_U241 , R1207_U242 , R1207_U243;
wire R1207_U244 , R1207_U245 , R1207_U246 , R1207_U247 , R1207_U248 , R1207_U249 , R1207_U250 , R1207_U251 , R1207_U252 , R1207_U253;
wire R1207_U254 , R1207_U255 , R1207_U256 , R1207_U257 , R1207_U258 , R1207_U259 , R1207_U260 , R1207_U261 , R1207_U262 , R1207_U263;
wire R1207_U264 , R1207_U265 , R1207_U266 , R1207_U267 , R1207_U268 , R1207_U269 , R1207_U270 , R1207_U271 , R1207_U272 , R1207_U273;
wire R1207_U274 , R1207_U275 , R1207_U276 , R1207_U277 , R1207_U278 , R1207_U279 , R1207_U280 , R1207_U281 , R1207_U282 , R1207_U283;
wire R1207_U284 , R1207_U285 , R1207_U286 , R1207_U287 , R1207_U288 , R1207_U289 , R1207_U290 , R1207_U291 , R1207_U292 , R1207_U293;
wire R1207_U294 , R1207_U295 , R1207_U296 , R1207_U297 , R1207_U298 , R1207_U299 , R1207_U300 , R1207_U301 , R1207_U302 , R1207_U303;
wire R1207_U304 , R1207_U305 , R1207_U306 , R1207_U307 , R1207_U308 , R1207_U309 , R1207_U310 , R1207_U311 , R1207_U312 , R1207_U313;
wire R1207_U314 , R1207_U315 , R1207_U316 , R1207_U317 , R1207_U318 , R1207_U319 , R1207_U320 , R1207_U321 , R1207_U322 , R1207_U323;
wire R1207_U324 , R1207_U325 , R1207_U326 , R1207_U327 , R1207_U328 , R1207_U329 , R1207_U330 , R1207_U331 , R1207_U332 , R1207_U333;
wire R1207_U334 , R1207_U335 , R1207_U336 , R1207_U337 , R1207_U338 , R1207_U339 , R1207_U340 , R1207_U341 , R1207_U342 , R1207_U343;
wire R1207_U344 , R1207_U345 , R1207_U346 , R1207_U347 , R1207_U348 , R1207_U349 , R1207_U350 , R1207_U351 , R1207_U352 , R1207_U353;
wire R1207_U354 , R1207_U355 , R1207_U356 , R1207_U357 , R1207_U358 , R1207_U359 , R1207_U360 , R1207_U361 , R1207_U362 , R1207_U363;
wire R1207_U364 , R1207_U365 , R1207_U366 , R1207_U367 , R1207_U368 , R1207_U369 , R1207_U370 , R1207_U371 , R1207_U372 , R1207_U373;
wire R1207_U374 , R1207_U375 , R1207_U376 , R1207_U377 , R1207_U378 , R1207_U379 , R1207_U380 , R1207_U381 , R1207_U382 , R1207_U383;
wire R1207_U384 , R1207_U385 , R1207_U386 , R1207_U387 , R1207_U388 , R1207_U389 , R1207_U390 , R1207_U391 , R1207_U392 , R1207_U393;
wire R1207_U394 , R1207_U395 , R1207_U396 , R1207_U397 , R1207_U398 , R1207_U399 , R1207_U400 , R1207_U401 , R1207_U402 , R1207_U403;
wire R1207_U404 , R1207_U405 , R1207_U406 , R1207_U407 , R1207_U408 , R1207_U409 , R1207_U410 , R1207_U411 , R1207_U412 , R1207_U413;
wire R1207_U414 , R1207_U415 , R1207_U416 , R1207_U417 , R1207_U418 , R1207_U419 , R1207_U420 , R1207_U421 , R1207_U422 , R1207_U423;
wire R1207_U424 , R1207_U425 , R1207_U426 , R1207_U427 , R1207_U428 , R1207_U429 , R1207_U430 , R1207_U431 , R1207_U432 , R1207_U433;
wire R1207_U434 , R1207_U435 , R1207_U436 , R1207_U437 , R1207_U438 , R1207_U439 , R1207_U440 , R1207_U441 , R1207_U442 , R1207_U443;
wire R1207_U444 , R1207_U445 , R1207_U446 , R1207_U447 , R1207_U448 , R1207_U449 , R1207_U450 , R1207_U451 , R1207_U452 , R1207_U453;
wire R1207_U454 , R1207_U455 , R1207_U456 , R1207_U457 , R1207_U458 , R1207_U459 , R1207_U460 , R1207_U461 , R1207_U462 , R1207_U463;
wire R1207_U464 , R1207_U465 , R1207_U466 , R1207_U467 , R1207_U468 , R1207_U469 , R1207_U470 , R1207_U471 , R1207_U472 , R1207_U473;
wire R1207_U474 , R1207_U475 , R1207_U476 , R1207_U477 , R1207_U478 , R1207_U479 , R1207_U480 , R1207_U481 , R1207_U482 , R1207_U483;
wire R1207_U484 , R1207_U485 , R1207_U486 , R1207_U487 , R1207_U488 , R1207_U489 , R1207_U490 , R1207_U491 , R1207_U492 , R1207_U493;
wire R1207_U494 , R1207_U495 , R1207_U496 , R1207_U497 , R1207_U498 , R1207_U499 , R1207_U500 , R1207_U501 , R1207_U502 , R1207_U503;
wire R1207_U504 , R1207_U505 , R1207_U506 , R1207_U507 , R1207_U508 , R1207_U509 , R1207_U510 , R1207_U511 , R1207_U512 , R1207_U513;
wire R1207_U514 , R1207_U515 , R1207_U516 , R1207_U517 , R1207_U518 , R1207_U519 , R1207_U520 , R1165_U4 , R1165_U5 , R1165_U6;
wire R1165_U7 , R1165_U8 , R1165_U9 , R1165_U10 , R1165_U11 , R1165_U12 , R1165_U13 , R1165_U14 , R1165_U15 , R1165_U16;
wire R1165_U17 , R1165_U18 , R1165_U19 , R1165_U20 , R1165_U21 , R1165_U22 , R1165_U23 , R1165_U24 , R1165_U25 , R1165_U26;
wire R1165_U27 , R1165_U28 , R1165_U29 , R1165_U30 , R1165_U31 , R1165_U32 , R1165_U33 , R1165_U34 , R1165_U35 , R1165_U36;
wire R1165_U37 , R1165_U38 , R1165_U39 , R1165_U40 , R1165_U41 , R1165_U42 , R1165_U43 , R1165_U44 , R1165_U45 , R1165_U46;
wire R1165_U47 , R1165_U48 , R1165_U49 , R1165_U50 , R1165_U51 , R1165_U52 , R1165_U53 , R1165_U54 , R1165_U55 , R1165_U56;
wire R1165_U57 , R1165_U58 , R1165_U59 , R1165_U60 , R1165_U61 , R1165_U62 , R1165_U63 , R1165_U64 , R1165_U65 , R1165_U66;
wire R1165_U67 , R1165_U68 , R1165_U69 , R1165_U70 , R1165_U71 , R1165_U72 , R1165_U73 , R1165_U74 , R1165_U75 , R1165_U76;
wire R1165_U77 , R1165_U78 , R1165_U79 , R1165_U80 , R1165_U81 , R1165_U82 , R1165_U83 , R1165_U84 , R1165_U85 , R1165_U86;
wire R1165_U87 , R1165_U88 , R1165_U89 , R1165_U90 , R1165_U91 , R1165_U92 , R1165_U93 , R1165_U94 , R1165_U95 , R1165_U96;
wire R1165_U97 , R1165_U98 , R1165_U99 , R1165_U100 , R1165_U101 , R1165_U102 , R1165_U103 , R1165_U104 , R1165_U105 , R1165_U106;
wire R1165_U107 , R1165_U108 , R1165_U109 , R1165_U110 , R1165_U111 , R1165_U112 , R1165_U113 , R1165_U114 , R1165_U115 , R1165_U116;
wire R1165_U117 , R1165_U118 , R1165_U119 , R1165_U120 , R1165_U121 , R1165_U122 , R1165_U123 , R1165_U124 , R1165_U125 , R1165_U126;
wire R1165_U127 , R1165_U128 , R1165_U129 , R1165_U130 , R1165_U131 , R1165_U132 , R1165_U133 , R1165_U134 , R1165_U135 , R1165_U136;
wire R1165_U137 , R1165_U138 , R1165_U139 , R1165_U140 , R1165_U141 , R1165_U142 , R1165_U143 , R1165_U144 , R1165_U145 , R1165_U146;
wire R1165_U147 , R1165_U148 , R1165_U149 , R1165_U150 , R1165_U151 , R1165_U152 , R1165_U153 , R1165_U154 , R1165_U155 , R1165_U156;
wire R1165_U157 , R1165_U158 , R1165_U159 , R1165_U160 , R1165_U161 , R1165_U162 , R1165_U163 , R1165_U164 , R1165_U165 , R1165_U166;
wire R1165_U167 , R1165_U168 , R1165_U169 , R1165_U170 , R1165_U171 , R1165_U172 , R1165_U173 , R1165_U174 , R1165_U175 , R1165_U176;
wire R1165_U177 , R1165_U178 , R1165_U179 , R1165_U180 , R1165_U181 , R1165_U182 , R1165_U183 , R1165_U184 , R1165_U185 , R1165_U186;
wire R1165_U187 , R1165_U188 , R1165_U189 , R1165_U190 , R1165_U191 , R1165_U192 , R1165_U193 , R1165_U194 , R1165_U195 , R1165_U196;
wire R1165_U197 , R1165_U198 , R1165_U199 , R1165_U200 , R1165_U201 , R1165_U202 , R1165_U203 , R1165_U204 , R1165_U205 , R1165_U206;
wire R1165_U207 , R1165_U208 , R1165_U209 , R1165_U210 , R1165_U211 , R1165_U212 , R1165_U213 , R1165_U214 , R1165_U215 , R1165_U216;
wire R1165_U217 , R1165_U218 , R1165_U219 , R1165_U220 , R1165_U221 , R1165_U222 , R1165_U223 , R1165_U224 , R1165_U225 , R1165_U226;
wire R1165_U227 , R1165_U228 , R1165_U229 , R1165_U230 , R1165_U231 , R1165_U232 , R1165_U233 , R1165_U234 , R1165_U235 , R1165_U236;
wire R1165_U237 , R1165_U238 , R1165_U239 , R1165_U240 , R1165_U241 , R1165_U242 , R1165_U243 , R1165_U244 , R1165_U245 , R1165_U246;
wire R1165_U247 , R1165_U248 , R1165_U249 , R1165_U250 , R1165_U251 , R1165_U252 , R1165_U253 , R1165_U254 , R1165_U255 , R1165_U256;
wire R1165_U257 , R1165_U258 , R1165_U259 , R1165_U260 , R1165_U261 , R1165_U262 , R1165_U263 , R1165_U264 , R1165_U265 , R1165_U266;
wire R1165_U267 , R1165_U268 , R1165_U269 , R1165_U270 , R1165_U271 , R1165_U272 , R1165_U273 , R1165_U274 , R1165_U275 , R1165_U276;
wire R1165_U277 , R1165_U278 , R1165_U279 , R1165_U280 , R1165_U281 , R1165_U282 , R1165_U283 , R1165_U284 , R1165_U285 , R1165_U286;
wire R1165_U287 , R1165_U288 , R1165_U289 , R1165_U290 , R1165_U291 , R1165_U292 , R1165_U293 , R1165_U294 , R1165_U295 , R1165_U296;
wire R1165_U297 , R1165_U298 , R1165_U299 , R1165_U300 , R1165_U301 , R1165_U302 , R1165_U303 , R1165_U304 , R1165_U305 , R1165_U306;
wire R1165_U307 , R1165_U308 , R1165_U309 , R1165_U310 , R1165_U311 , R1165_U312 , R1165_U313 , R1165_U314 , R1165_U315 , R1165_U316;
wire R1165_U317 , R1165_U318 , R1165_U319 , R1165_U320 , R1165_U321 , R1165_U322 , R1165_U323 , R1165_U324 , R1165_U325 , R1165_U326;
wire R1165_U327 , R1165_U328 , R1165_U329 , R1165_U330 , R1165_U331 , R1165_U332 , R1165_U333 , R1165_U334 , R1165_U335 , R1165_U336;
wire R1165_U337 , R1165_U338 , R1165_U339 , R1165_U340 , R1165_U341 , R1165_U342 , R1165_U343 , R1165_U344 , R1165_U345 , R1165_U346;
wire R1165_U347 , R1165_U348 , R1165_U349 , R1165_U350 , R1165_U351 , R1165_U352 , R1165_U353 , R1165_U354 , R1165_U355 , R1165_U356;
wire R1165_U357 , R1165_U358 , R1165_U359 , R1165_U360 , R1165_U361 , R1165_U362 , R1165_U363 , R1165_U364 , R1165_U365 , R1165_U366;
wire R1165_U367 , R1165_U368 , R1165_U369 , R1165_U370 , R1165_U371 , R1165_U372 , R1165_U373 , R1165_U374 , R1165_U375 , R1165_U376;
wire R1165_U377 , R1165_U378 , R1165_U379 , R1165_U380 , R1165_U381 , R1165_U382 , R1165_U383 , R1165_U384 , R1165_U385 , R1165_U386;
wire R1165_U387 , R1165_U388 , R1165_U389 , R1165_U390 , R1165_U391 , R1165_U392 , R1165_U393 , R1165_U394 , R1165_U395 , R1165_U396;
wire R1165_U397 , R1165_U398 , R1165_U399 , R1165_U400 , R1165_U401 , R1165_U402 , R1165_U403 , R1165_U404 , R1165_U405 , R1165_U406;
wire R1165_U407 , R1165_U408 , R1165_U409 , R1165_U410 , R1165_U411 , R1165_U412 , R1165_U413 , R1165_U414 , R1165_U415 , R1165_U416;
wire R1165_U417 , R1165_U418 , R1165_U419 , R1165_U420 , R1165_U421 , R1165_U422 , R1165_U423 , R1165_U424 , R1165_U425 , R1165_U426;
wire R1165_U427 , R1165_U428 , R1165_U429 , R1165_U430 , R1165_U431 , R1165_U432 , R1165_U433 , R1165_U434 , R1165_U435 , R1165_U436;
wire R1165_U437 , R1165_U438 , R1165_U439 , R1165_U440 , R1165_U441 , R1165_U442 , R1165_U443 , R1165_U444 , R1165_U445 , R1165_U446;
wire R1165_U447 , R1165_U448 , R1165_U449 , R1165_U450 , R1165_U451 , R1165_U452 , R1165_U453 , R1165_U454 , R1165_U455 , R1165_U456;
wire R1165_U457 , R1165_U458 , R1165_U459 , R1165_U460 , R1165_U461 , R1165_U462 , R1165_U463 , R1165_U464 , R1165_U465 , R1165_U466;
wire R1165_U467 , R1165_U468 , R1165_U469 , R1165_U470 , R1165_U471 , R1165_U472 , R1165_U473 , R1165_U474 , R1165_U475 , R1165_U476;
wire R1165_U477 , R1165_U478 , R1165_U479 , R1165_U480 , R1165_U481 , R1165_U482 , R1165_U483 , R1165_U484 , R1165_U485 , R1165_U486;
wire R1165_U487 , R1165_U488 , R1165_U489 , R1165_U490 , R1165_U491 , R1165_U492 , R1165_U493 , R1165_U494 , R1165_U495 , R1165_U496;
wire R1165_U497 , R1165_U498 , R1165_U499 , R1165_U500 , R1165_U501 , R1165_U502 , R1165_U503 , R1165_U504 , R1165_U505 , R1165_U506;
wire R1165_U507 , R1165_U508 , R1165_U509 , R1165_U510 , R1165_U511 , R1165_U512 , R1165_U513 , R1165_U514 , R1165_U515 , R1165_U516;
wire R1165_U517 , R1165_U518 , R1165_U519 , R1165_U520 , R1165_U521 , R1165_U522 , R1165_U523 , R1165_U524 , R1165_U525 , R1165_U526;
wire R1165_U527 , R1165_U528 , R1165_U529 , R1165_U530 , R1165_U531 , R1165_U532 , R1165_U533 , R1165_U534 , R1165_U535 , R1165_U536;
wire R1165_U537 , R1165_U538 , R1165_U539 , R1165_U540 , R1165_U541 , R1165_U542 , R1165_U543 , R1165_U544 , R1165_U545 , R1165_U546;
wire R1165_U547 , R1165_U548 , R1165_U549 , R1165_U550 , R1165_U551 , R1165_U552 , R1165_U553 , R1165_U554 , R1165_U555 , R1165_U556;
wire R1165_U557 , R1165_U558 , R1165_U559 , R1165_U560 , R1165_U561 , R1165_U562 , R1165_U563 , R1165_U564 , R1165_U565 , R1165_U566;
wire R1165_U567 , R1165_U568 , R1165_U569 , R1165_U570 , R1165_U571 , R1165_U572 , R1165_U573 , R1165_U574 , R1165_U575 , R1165_U576;
wire R1165_U577 , R1165_U578 , R1165_U579 , R1165_U580 , R1165_U581 , R1165_U582 , R1165_U583 , R1165_U584 , R1165_U585 , R1165_U586;
wire R1165_U587 , R1165_U588 , R1165_U589 , R1165_U590 , R1165_U591 , R1165_U592 , R1165_U593 , R1165_U594 , R1165_U595 , R1165_U596;
wire R1165_U597 , R1165_U598 , R1165_U599 , R1165_U600 , R1165_U601 , R1165_U602 , R1165_U603 , R1165_U604 , R1165_U605 , R1165_U606;
wire R1165_U607 , R1165_U608 , R1165_U609 , R1165_U610 , R1165_U611 , R1165_U612 , R1165_U613 , R1150_U6 , R1150_U7 , R1150_U8;
wire R1150_U9 , R1150_U10 , R1150_U11 , R1150_U12 , R1150_U13 , R1150_U14 , R1150_U15 , R1150_U16 , R1150_U17 , R1150_U18;
wire R1150_U19 , R1150_U20 , R1150_U21 , R1150_U22 , R1150_U23 , R1150_U24 , R1150_U25 , R1150_U26 , R1150_U27 , R1150_U28;
wire R1150_U29 , R1150_U30 , R1150_U31 , R1150_U32 , R1150_U33 , R1150_U34 , R1150_U35 , R1150_U36 , R1150_U37 , R1150_U38;
wire R1150_U39 , R1150_U40 , R1150_U41 , R1150_U42 , R1150_U43 , R1150_U44 , R1150_U45 , R1150_U46 , R1150_U47 , R1150_U48;
wire R1150_U49 , R1150_U50 , R1150_U51 , R1150_U52 , R1150_U53 , R1150_U54 , R1150_U55 , R1150_U56 , R1150_U57 , R1150_U58;
wire R1150_U59 , R1150_U60 , R1150_U61 , R1150_U62 , R1150_U63 , R1150_U64 , R1150_U65 , R1150_U66 , R1150_U67 , R1150_U68;
wire R1150_U69 , R1150_U70 , R1150_U71 , R1150_U72 , R1150_U73 , R1150_U74 , R1150_U75 , R1150_U76 , R1150_U77 , R1150_U78;
wire R1150_U79 , R1150_U80 , R1150_U81 , R1150_U82 , R1150_U83 , R1150_U84 , R1150_U85 , R1150_U86 , R1150_U87 , R1150_U88;
wire R1150_U89 , R1150_U90 , R1150_U91 , R1150_U92 , R1150_U93 , R1150_U94 , R1150_U95 , R1150_U96 , R1150_U97 , R1150_U98;
wire R1150_U99 , R1150_U100 , R1150_U101 , R1150_U102 , R1150_U103 , R1150_U104 , R1150_U105 , R1150_U106 , R1150_U107 , R1150_U108;
wire R1150_U109 , R1150_U110 , R1150_U111 , R1150_U112 , R1150_U113 , R1150_U114 , R1150_U115 , R1150_U116 , R1150_U117 , R1150_U118;
wire R1150_U119 , R1150_U120 , R1150_U121 , R1150_U122 , R1150_U123 , R1150_U124 , R1150_U125 , R1150_U126 , R1150_U127 , R1150_U128;
wire R1150_U129 , R1150_U130 , R1150_U131 , R1150_U132 , R1150_U133 , R1150_U134 , R1150_U135 , R1150_U136 , R1150_U137 , R1150_U138;
wire R1150_U139 , R1150_U140 , R1150_U141 , R1150_U142 , R1150_U143 , R1150_U144 , R1150_U145 , R1150_U146 , R1150_U147 , R1150_U148;
wire R1150_U149 , R1150_U150 , R1150_U151 , R1150_U152 , R1150_U153 , R1150_U154 , R1150_U155 , R1150_U156 , R1150_U157 , R1150_U158;
wire R1150_U159 , R1150_U160 , R1150_U161 , R1150_U162 , R1150_U163 , R1150_U164 , R1150_U165 , R1150_U166 , R1150_U167 , R1150_U168;
wire R1150_U169 , R1150_U170 , R1150_U171 , R1150_U172 , R1150_U173 , R1150_U174 , R1150_U175 , R1150_U176 , R1150_U177 , R1150_U178;
wire R1150_U179 , R1150_U180 , R1150_U181 , R1150_U182 , R1150_U183 , R1150_U184 , R1150_U185 , R1150_U186 , R1150_U187 , R1150_U188;
wire R1150_U189 , R1150_U190 , R1150_U191 , R1150_U192 , R1150_U193 , R1150_U194 , R1150_U195 , R1150_U196 , R1150_U197 , R1150_U198;
wire R1150_U199 , R1150_U200 , R1150_U201 , R1150_U202 , R1150_U203 , R1150_U204 , R1150_U205 , R1150_U206 , R1150_U207 , R1150_U208;
wire R1150_U209 , R1150_U210 , R1150_U211 , R1150_U212 , R1150_U213 , R1150_U214 , R1150_U215 , R1150_U216 , R1150_U217 , R1150_U218;
wire R1150_U219 , R1150_U220 , R1150_U221 , R1150_U222 , R1150_U223 , R1150_U224 , R1150_U225 , R1150_U226 , R1150_U227 , R1150_U228;
wire R1150_U229 , R1150_U230 , R1150_U231 , R1150_U232 , R1150_U233 , R1150_U234 , R1150_U235 , R1150_U236 , R1150_U237 , R1150_U238;
wire R1150_U239 , R1150_U240 , R1150_U241 , R1150_U242 , R1150_U243 , R1150_U244 , R1150_U245 , R1150_U246 , R1150_U247 , R1150_U248;
wire R1150_U249 , R1150_U250 , R1150_U251 , R1150_U252 , R1150_U253 , R1150_U254 , R1150_U255 , R1150_U256 , R1150_U257 , R1150_U258;
wire R1150_U259 , R1150_U260 , R1150_U261 , R1150_U262 , R1150_U263 , R1150_U264 , R1150_U265 , R1150_U266 , R1150_U267 , R1150_U268;
wire R1150_U269 , R1150_U270 , R1150_U271 , R1150_U272 , R1150_U273 , R1150_U274 , R1150_U275 , R1150_U276 , R1150_U277 , R1150_U278;
wire R1150_U279 , R1150_U280 , R1150_U281 , R1150_U282 , R1150_U283 , R1150_U284 , R1150_U285 , R1150_U286 , R1150_U287 , R1150_U288;
wire R1150_U289 , R1150_U290 , R1150_U291 , R1150_U292 , R1150_U293 , R1150_U294 , R1150_U295 , R1150_U296 , R1150_U297 , R1150_U298;
wire R1150_U299 , R1150_U300 , R1150_U301 , R1150_U302 , R1150_U303 , R1150_U304 , R1150_U305 , R1150_U306 , R1150_U307 , R1150_U308;
wire R1150_U309 , R1150_U310 , R1150_U311 , R1150_U312 , R1150_U313 , R1150_U314 , R1150_U315 , R1150_U316 , R1150_U317 , R1150_U318;
wire R1150_U319 , R1150_U320 , R1150_U321 , R1150_U322 , R1150_U323 , R1150_U324 , R1150_U325 , R1150_U326 , R1150_U327 , R1150_U328;
wire R1150_U329 , R1150_U330 , R1150_U331 , R1150_U332 , R1150_U333 , R1150_U334 , R1150_U335 , R1150_U336 , R1150_U337 , R1150_U338;
wire R1150_U339 , R1150_U340 , R1150_U341 , R1150_U342 , R1150_U343 , R1150_U344 , R1150_U345 , R1150_U346 , R1150_U347 , R1150_U348;
wire R1150_U349 , R1150_U350 , R1150_U351 , R1150_U352 , R1150_U353 , R1150_U354 , R1150_U355 , R1150_U356 , R1150_U357 , R1150_U358;
wire R1150_U359 , R1150_U360 , R1150_U361 , R1150_U362 , R1150_U363 , R1150_U364 , R1150_U365 , R1150_U366 , R1150_U367 , R1150_U368;
wire R1150_U369 , R1150_U370 , R1150_U371 , R1150_U372 , R1150_U373 , R1150_U374 , R1150_U375 , R1150_U376 , R1150_U377 , R1150_U378;
wire R1150_U379 , R1150_U380 , R1150_U381 , R1150_U382 , R1150_U383 , R1150_U384 , R1150_U385 , R1150_U386 , R1150_U387 , R1150_U388;
wire R1150_U389 , R1150_U390 , R1150_U391 , R1150_U392 , R1150_U393 , R1150_U394 , R1150_U395 , R1150_U396 , R1150_U397 , R1150_U398;
wire R1150_U399 , R1150_U400 , R1150_U401 , R1150_U402 , R1150_U403 , R1150_U404 , R1150_U405 , R1150_U406 , R1150_U407 , R1150_U408;
wire R1150_U409 , R1150_U410 , R1150_U411 , R1150_U412 , R1150_U413 , R1150_U414 , R1150_U415 , R1150_U416 , R1150_U417 , R1150_U418;
wire R1150_U419 , R1150_U420 , R1150_U421 , R1150_U422 , R1150_U423 , R1150_U424 , R1150_U425 , R1150_U426 , R1150_U427 , R1150_U428;
wire R1150_U429 , R1150_U430 , R1150_U431 , R1150_U432 , R1150_U433 , R1150_U434 , R1150_U435 , R1150_U436 , R1150_U437 , R1150_U438;
wire R1150_U439 , R1150_U440 , R1150_U441 , R1150_U442 , R1150_U443 , R1150_U444 , R1150_U445 , R1150_U446 , R1150_U447 , R1150_U448;
wire R1150_U449 , R1150_U450 , R1150_U451 , R1150_U452 , R1150_U453 , R1150_U454 , R1150_U455 , R1150_U456 , R1150_U457 , R1150_U458;
wire R1150_U459 , R1150_U460 , R1150_U461 , R1150_U462 , R1150_U463 , R1150_U464 , R1150_U465 , R1150_U466 , R1150_U467 , R1150_U468;
wire R1150_U469 , R1150_U470 , R1150_U471 , R1150_U472 , R1150_U473 , R1150_U474 , R1150_U475 , R1150_U476 , R1150_U477 , R1150_U478;
wire R1150_U479 , R1150_U480 , R1150_U481 , R1150_U482 , R1150_U483 , R1150_U484 , R1150_U485 , R1150_U486 , R1150_U487 , R1150_U488;
wire R1150_U489 , R1150_U490 , R1150_U491 , R1150_U492 , R1150_U493 , R1150_U494 , R1150_U495 , R1150_U496 , R1150_U497 , R1150_U498;
wire R1150_U499 , R1150_U500 , R1150_U501 , R1150_U502 , R1150_U503 , R1150_U504 , R1150_U505 , R1150_U506 , R1150_U507 , R1150_U508;
wire R1150_U509 , R1150_U510 , R1150_U511 , R1192_U6 , R1192_U7 , R1192_U8 , R1192_U9 , R1192_U10 , R1192_U11 , R1192_U12;
wire R1192_U13 , R1192_U14 , R1192_U15 , R1192_U16 , R1192_U17 , R1192_U18 , R1192_U19 , R1192_U20 , R1192_U21 , R1192_U22;
wire R1192_U23 , R1192_U24 , R1192_U25 , R1192_U26 , R1192_U27 , R1192_U28 , R1192_U29 , R1192_U30 , R1192_U31 , R1192_U32;
wire R1192_U33 , R1192_U34 , R1192_U35 , R1192_U36 , R1192_U37 , R1192_U38 , R1192_U39 , R1192_U40 , R1192_U41 , R1192_U42;
wire R1192_U43 , R1192_U44 , R1192_U45 , R1192_U46 , R1192_U47 , R1192_U48 , R1192_U49 , R1192_U50 , R1192_U51 , R1192_U52;
wire R1192_U53 , R1192_U54 , R1192_U55 , R1192_U56 , R1192_U57 , R1192_U58 , R1192_U59 , R1192_U60 , R1192_U61 , R1192_U62;
wire R1192_U63 , R1192_U64 , R1192_U65 , R1192_U66 , R1192_U67 , R1192_U68 , R1192_U69 , R1192_U70 , R1192_U71 , R1192_U72;
wire R1192_U73 , R1192_U74 , R1192_U75 , R1192_U76 , R1192_U77 , R1192_U78 , R1192_U79 , R1192_U80 , R1192_U81 , R1192_U82;
wire R1192_U83 , R1192_U84 , R1192_U85 , R1192_U86 , R1192_U87 , R1192_U88 , R1192_U89 , R1192_U90 , R1192_U91 , R1192_U92;
wire R1192_U93 , R1192_U94 , R1192_U95 , R1192_U96 , R1192_U97 , R1192_U98 , R1192_U99 , R1192_U100 , R1192_U101 , R1192_U102;
wire R1192_U103 , R1192_U104 , R1192_U105 , R1192_U106 , R1192_U107 , R1192_U108 , R1192_U109 , R1192_U110 , R1192_U111 , R1192_U112;
wire R1192_U113 , R1192_U114 , R1192_U115 , R1192_U116 , R1192_U117 , R1192_U118 , R1192_U119 , R1192_U120 , R1192_U121 , R1192_U122;
wire R1192_U123 , R1192_U124 , R1192_U125 , R1192_U126 , R1192_U127 , R1192_U128 , R1192_U129 , R1192_U130 , R1192_U131 , R1192_U132;
wire R1192_U133 , R1192_U134 , R1192_U135 , R1192_U136 , R1192_U137 , R1192_U138 , R1192_U139 , R1192_U140 , R1192_U141 , R1192_U142;
wire R1192_U143 , R1192_U144 , R1192_U145 , R1192_U146 , R1192_U147 , R1192_U148 , R1192_U149 , R1192_U150 , R1192_U151 , R1192_U152;
wire R1192_U153 , R1192_U154 , R1192_U155 , R1192_U156 , R1192_U157 , R1192_U158 , R1192_U159 , R1192_U160 , R1192_U161 , R1192_U162;
wire R1192_U163 , R1192_U164 , R1192_U165 , R1192_U166 , R1192_U167 , R1192_U168 , R1192_U169 , R1192_U170 , R1192_U171 , R1192_U172;
wire R1192_U173 , R1192_U174 , R1192_U175 , R1192_U176 , R1192_U177 , R1192_U178 , R1192_U179 , R1192_U180 , R1192_U181 , R1192_U182;
wire R1192_U183 , R1192_U184 , R1192_U185 , R1192_U186 , R1192_U187 , R1192_U188 , R1192_U189 , R1192_U190 , R1192_U191 , R1192_U192;
wire R1192_U193 , R1192_U194 , R1192_U195 , R1192_U196 , R1192_U197 , R1192_U198 , R1192_U199 , R1192_U200 , R1192_U201 , R1192_U202;
wire R1192_U203 , R1192_U204 , R1192_U205 , R1192_U206 , R1192_U207 , R1192_U208 , R1192_U209 , R1192_U210 , R1192_U211 , R1192_U212;
wire R1192_U213 , R1192_U214 , R1192_U215 , R1192_U216 , R1192_U217 , R1192_U218 , R1192_U219 , R1192_U220 , R1192_U221 , R1192_U222;
wire R1192_U223 , R1192_U224 , R1192_U225 , R1192_U226 , R1192_U227 , R1192_U228 , R1192_U229 , R1192_U230 , R1192_U231 , R1192_U232;
wire R1192_U233 , R1192_U234 , R1192_U235 , R1192_U236 , R1192_U237 , R1192_U238 , R1192_U239 , R1192_U240 , R1192_U241 , R1192_U242;
wire R1192_U243 , R1192_U244 , R1192_U245 , R1192_U246 , R1192_U247 , R1192_U248 , R1192_U249 , R1192_U250 , R1192_U251 , R1192_U252;
wire R1192_U253 , R1192_U254 , R1192_U255 , R1192_U256 , R1192_U257 , R1192_U258 , R1192_U259 , R1192_U260 , R1192_U261 , R1192_U262;
wire R1192_U263 , R1192_U264 , R1192_U265 , R1192_U266 , R1192_U267 , R1192_U268 , R1192_U269 , R1192_U270 , R1192_U271 , R1192_U272;
wire R1192_U273 , R1192_U274 , R1192_U275 , R1192_U276 , R1192_U277 , R1192_U278 , R1192_U279 , R1192_U280 , R1192_U281 , R1192_U282;
wire R1192_U283 , R1192_U284 , R1192_U285 , R1192_U286 , R1192_U287 , R1192_U288 , R1192_U289 , R1192_U290 , R1192_U291 , R1192_U292;
wire R1192_U293 , R1192_U294 , R1192_U295 , R1192_U296 , R1192_U297 , R1192_U298 , R1192_U299 , R1192_U300 , R1192_U301 , R1192_U302;
wire R1192_U303 , R1192_U304 , R1192_U305 , R1192_U306 , R1192_U307 , R1192_U308 , R1192_U309 , R1192_U310 , R1192_U311 , R1192_U312;
wire R1192_U313 , R1192_U314 , R1192_U315 , R1192_U316 , R1192_U317 , R1192_U318 , R1192_U319 , R1192_U320 , R1192_U321 , R1192_U322;
wire R1192_U323 , R1192_U324 , R1192_U325 , R1192_U326 , R1192_U327 , R1192_U328 , R1192_U329 , R1192_U330 , R1192_U331 , R1192_U332;
wire R1192_U333 , R1192_U334 , R1192_U335 , R1192_U336 , R1192_U337 , R1192_U338 , R1192_U339 , R1192_U340 , R1192_U341 , R1192_U342;
wire R1192_U343 , R1192_U344 , R1192_U345 , R1192_U346 , R1192_U347 , R1192_U348 , R1192_U349 , R1192_U350 , R1192_U351 , R1192_U352;
wire R1192_U353 , R1192_U354 , R1192_U355 , R1192_U356 , R1192_U357 , R1192_U358 , R1192_U359 , R1192_U360 , R1192_U361 , R1192_U362;
wire R1192_U363 , R1192_U364 , R1192_U365 , R1192_U366 , R1192_U367 , R1192_U368 , R1192_U369 , R1192_U370 , R1192_U371 , R1192_U372;
wire R1192_U373 , R1192_U374 , R1192_U375 , R1192_U376 , R1192_U377 , R1192_U378 , R1192_U379 , R1192_U380 , R1192_U381 , R1192_U382;
wire R1192_U383 , R1192_U384 , R1192_U385 , R1192_U386 , R1192_U387 , R1192_U388 , R1192_U389 , R1192_U390 , R1192_U391 , R1192_U392;
wire R1192_U393 , R1192_U394 , R1192_U395 , R1192_U396 , R1192_U397 , R1192_U398 , R1192_U399 , R1192_U400 , R1192_U401 , R1192_U402;
wire R1192_U403 , R1192_U404 , R1192_U405 , R1192_U406 , R1192_U407 , R1192_U408 , R1192_U409 , R1192_U410 , R1192_U411 , R1192_U412;
wire R1192_U413 , R1192_U414 , R1192_U415 , R1192_U416 , R1192_U417 , R1192_U418 , R1192_U419 , R1192_U420 , R1192_U421 , R1192_U422;
wire R1192_U423 , R1192_U424 , R1192_U425 , R1192_U426 , R1192_U427 , R1192_U428 , R1192_U429 , R1192_U430 , R1192_U431 , R1192_U432;
wire R1192_U433 , R1192_U434 , R1192_U435 , R1192_U436 , R1192_U437 , R1192_U438 , R1192_U439 , R1192_U440 , R1192_U441 , R1192_U442;
wire R1192_U443 , R1192_U444 , R1192_U445 , R1192_U446 , R1192_U447 , R1192_U448 , R1192_U449 , R1192_U450 , R1192_U451 , R1192_U452;
wire R1192_U453 , R1192_U454 , R1192_U455 , R1192_U456 , R1192_U457 , R1192_U458 , R1192_U459 , R1192_U460 , R1192_U461 , R1192_U462;
wire R1192_U463 , R1192_U464 , R1192_U465 , R1192_U466 , R1192_U467 , R1192_U468 , R1192_U469 , R1192_U470 , R1192_U471 , R1192_U472;
wire R1192_U473 , R1192_U474 , R1192_U475 , R1192_U476 , R1192_U477 , R1192_U478 , R1192_U479 , R1192_U480 , R1192_U481 , R1192_U482;
wire R1192_U483 , R1192_U484 , R1192_U485 , R1192_U486 , R1192_U487 , R1192_U488 , R1192_U489 , R1192_U490 , R1192_U491 , R1192_U492;
wire R1192_U493 , R1192_U494 , R1192_U495 , R1192_U496 , R1192_U497 , R1192_U498 , R1192_U499 , R1192_U500 , R1192_U501 , R1192_U502;
wire R1192_U503 , R1192_U504 , R1192_U505 , R1192_U506 , R1192_U507 , R1192_U508 , R1192_U509 , R1192_U510 , R1192_U511 , R1192_U512;
wire R1192_U513 , R1192_U514 , R1192_U515 , R1192_U516 , R1192_U517 , R1192_U518 , R1192_U519 , R1192_U520 , R1347_U6 , R1347_U7;
wire R1347_U8 , R1347_U9 , R1347_U10 , R1347_U11 , R1347_U12 , R1347_U13 , R1347_U14 , R1347_U15 , R1347_U16 , R1347_U17;
wire R1347_U18 , R1347_U19 , R1347_U20 , R1347_U21 , R1347_U22 , R1347_U23 , R1347_U24 , R1347_U25 , R1347_U26 , R1347_U27;
wire R1347_U28 , R1347_U29 , R1347_U30 , R1347_U31 , R1347_U32 , R1347_U33 , R1347_U34 , R1347_U35 , R1347_U36 , R1347_U37;
wire R1347_U38 , R1347_U39 , R1347_U40 , R1347_U41 , R1347_U42 , R1347_U43 , R1347_U44 , R1347_U45 , R1347_U46 , R1347_U47;
wire R1347_U48 , R1347_U49 , R1347_U50 , R1347_U51 , R1347_U52 , R1347_U53 , R1347_U54 , R1347_U55 , R1347_U56 , R1347_U57;
wire R1347_U58 , R1347_U59 , R1347_U60 , R1347_U61 , R1347_U62 , R1347_U63 , R1347_U64 , R1347_U65 , R1347_U66 , R1347_U67;
wire R1347_U68 , R1347_U69 , R1347_U70 , R1347_U71 , R1347_U72 , R1347_U73 , R1347_U74 , R1347_U75 , R1347_U76 , R1347_U77;
wire R1347_U78 , R1347_U79 , R1347_U80 , R1347_U81 , R1347_U82 , R1347_U83 , R1347_U84 , R1347_U85 , R1347_U86 , R1347_U87;
wire R1347_U88 , R1347_U89 , R1347_U90 , R1347_U91 , R1347_U92 , R1347_U93 , R1347_U94 , R1347_U95 , R1347_U96 , R1347_U97;
wire R1347_U98 , R1347_U99 , R1347_U100 , R1347_U101 , R1347_U102 , R1347_U103 , R1347_U104 , R1347_U105 , R1347_U106 , R1347_U107;
wire R1347_U108 , R1347_U109 , R1347_U110 , R1347_U111 , R1347_U112 , R1347_U113 , R1347_U114 , R1347_U115 , R1347_U116 , R1347_U117;
wire R1347_U118 , R1347_U119 , R1347_U120 , R1347_U121 , R1347_U122 , R1347_U123 , R1347_U124 , R1347_U125 , R1347_U126 , R1347_U127;
wire R1347_U128 , R1347_U129 , R1347_U130 , R1347_U131 , R1347_U132 , R1347_U133 , R1347_U134 , R1347_U135 , R1347_U136 , R1347_U137;
wire R1347_U138 , R1347_U139 , R1347_U140 , R1347_U141 , R1347_U142 , R1347_U143 , R1347_U144 , R1347_U145 , R1347_U146 , R1347_U147;
wire R1347_U148 , R1347_U149 , R1347_U150 , R1347_U151 , R1347_U152 , R1347_U153 , R1347_U154 , R1347_U155 , R1347_U156 , R1347_U157;
wire R1347_U158 , R1347_U159 , R1347_U160 , R1347_U161 , R1347_U162 , R1347_U163 , R1347_U164 , R1347_U165 , R1347_U166 , R1347_U167;
wire R1347_U168 , R1347_U169 , R1347_U170 , R1347_U171 , R1347_U172 , R1347_U173 , R1347_U174 , R1347_U175 , R1347_U176 , R1347_U177;
wire R1347_U178 , R1347_U179 , R1347_U180 , R1347_U181 , R1347_U182 , R1347_U183 , R1347_U184 , R1347_U185 , R1347_U186 , R1347_U187;
wire R1347_U188 , R1347_U189 , R1347_U190 , R1347_U191 , R1347_U192 , R1347_U193 , R1347_U194 , R1347_U195 , R1347_U196 , R1347_U197;
wire R1347_U198 , R1347_U199 , R1347_U200 , R1347_U201 , R1347_U202 , R1347_U203 , R1347_U204 , R1347_U205 , R1347_U206 , R1347_U207;
wire R1347_U208 , R1347_U209 , R1347_U210 , R1347_U211 , R1347_U212 , R1171_U4 , R1171_U5 , R1171_U6 , R1171_U7 , R1171_U8;
wire R1171_U9 , R1171_U10 , R1171_U11 , R1171_U12 , R1171_U13 , R1171_U14 , R1171_U15 , R1171_U16 , R1171_U17 , R1171_U18;
wire R1171_U19 , R1171_U20 , R1171_U21 , R1171_U22 , R1171_U23 , R1171_U24 , R1171_U25 , R1171_U26 , R1171_U27 , R1171_U28;
wire R1171_U29 , R1171_U30 , R1171_U31 , R1171_U32 , R1171_U33 , R1171_U34 , R1171_U35 , R1171_U36 , R1171_U37 , R1171_U38;
wire R1171_U39 , R1171_U40 , R1171_U41 , R1171_U42 , R1171_U43 , R1171_U44 , R1171_U45 , R1171_U46 , R1171_U47 , R1171_U48;
wire R1171_U49 , R1171_U50 , R1171_U51 , R1171_U52 , R1171_U53 , R1171_U54 , R1171_U55 , R1171_U56 , R1171_U57 , R1171_U58;
wire R1171_U59 , R1171_U60 , R1171_U61 , R1171_U62 , R1171_U63 , R1171_U64 , R1171_U65 , R1171_U66 , R1171_U67 , R1171_U68;
wire R1171_U69 , R1171_U70 , R1171_U71 , R1171_U72 , R1171_U73 , R1171_U74 , R1171_U75 , R1171_U76 , R1171_U77 , R1171_U78;
wire R1171_U79 , R1171_U80 , R1171_U81 , R1171_U82 , R1171_U83 , R1171_U84 , R1171_U85 , R1171_U86 , R1171_U87 , R1171_U88;
wire R1171_U89 , R1171_U90 , R1171_U91 , R1171_U92 , R1171_U93 , R1171_U94 , R1171_U95 , R1171_U96 , R1171_U97 , R1171_U98;
wire R1171_U99 , R1171_U100 , R1171_U101 , R1171_U102 , R1171_U103 , R1171_U104 , R1171_U105 , R1171_U106 , R1171_U107 , R1171_U108;
wire R1171_U109 , R1171_U110 , R1171_U111 , R1171_U112 , R1171_U113 , R1171_U114 , R1171_U115 , R1171_U116 , R1171_U117 , R1171_U118;
wire R1171_U119 , R1171_U120 , R1171_U121 , R1171_U122 , R1171_U123 , R1171_U124 , R1171_U125 , R1171_U126 , R1171_U127 , R1171_U128;
wire R1171_U129 , R1171_U130 , R1171_U131 , R1171_U132 , R1171_U133 , R1171_U134 , R1171_U135 , R1171_U136 , R1171_U137 , R1171_U138;
wire R1171_U139 , R1171_U140 , R1171_U141 , R1171_U142 , R1171_U143 , R1171_U144 , R1171_U145 , R1171_U146 , R1171_U147 , R1171_U148;
wire R1171_U149 , R1171_U150 , R1171_U151 , R1171_U152 , R1171_U153 , R1171_U154 , R1171_U155 , R1171_U156 , R1171_U157 , R1171_U158;
wire R1171_U159 , R1171_U160 , R1171_U161 , R1171_U162 , R1171_U163 , R1171_U164 , R1171_U165 , R1171_U166 , R1171_U167 , R1171_U168;
wire R1171_U169 , R1171_U170 , R1171_U171 , R1171_U172 , R1171_U173 , R1171_U174 , R1171_U175 , R1171_U176 , R1171_U177 , R1171_U178;
wire R1171_U179 , R1171_U180 , R1171_U181 , R1171_U182 , R1171_U183 , R1171_U184 , R1171_U185 , R1171_U186 , R1171_U187 , R1171_U188;
wire R1171_U189 , R1171_U190 , R1171_U191 , R1171_U192 , R1171_U193 , R1171_U194 , R1171_U195 , R1171_U196 , R1171_U197 , R1171_U198;
wire R1171_U199 , R1171_U200 , R1171_U201 , R1171_U202 , R1171_U203 , R1171_U204 , R1171_U205 , R1171_U206 , R1171_U207 , R1171_U208;
wire R1171_U209 , R1171_U210 , R1171_U211 , R1171_U212 , R1171_U213 , R1171_U214 , R1171_U215 , R1171_U216 , R1171_U217 , R1171_U218;
wire R1171_U219 , R1171_U220 , R1171_U221 , R1171_U222 , R1171_U223 , R1171_U224 , R1171_U225 , R1171_U226 , R1171_U227 , R1171_U228;
wire R1171_U229 , R1171_U230 , R1171_U231 , R1171_U232 , R1171_U233 , R1171_U234 , R1171_U235 , R1171_U236 , R1171_U237 , R1171_U238;
wire R1171_U239 , R1171_U240 , R1171_U241 , R1171_U242 , R1171_U243 , R1171_U244 , R1171_U245 , R1171_U246 , R1171_U247 , R1171_U248;
wire R1171_U249 , R1171_U250 , R1171_U251 , R1171_U252 , R1171_U253 , R1171_U254 , R1171_U255 , R1171_U256 , R1171_U257 , R1171_U258;
wire R1171_U259 , R1171_U260 , R1171_U261 , R1171_U262 , R1171_U263 , R1171_U264 , R1171_U265 , R1171_U266 , R1171_U267 , R1171_U268;
wire R1171_U269 , R1171_U270 , R1171_U271 , R1171_U272 , R1171_U273 , R1171_U274 , R1171_U275 , R1171_U276 , R1171_U277 , R1171_U278;
wire R1171_U279 , R1171_U280 , R1171_U281 , R1171_U282 , R1171_U283 , R1171_U284 , R1171_U285 , R1171_U286 , R1171_U287 , R1171_U288;
wire R1171_U289 , R1171_U290 , R1171_U291 , R1171_U292 , R1171_U293 , R1171_U294 , R1171_U295 , R1171_U296 , R1171_U297 , R1171_U298;
wire R1171_U299 , R1171_U300 , R1171_U301 , R1171_U302 , R1171_U303 , R1171_U304 , R1171_U305 , R1171_U306 , R1171_U307 , R1171_U308;
wire R1171_U309 , R1171_U310 , R1171_U311 , R1171_U312 , R1171_U313 , R1171_U314 , R1171_U315 , R1171_U316 , R1171_U317 , R1171_U318;
wire R1171_U319 , R1171_U320 , R1171_U321 , R1171_U322 , R1171_U323 , R1171_U324 , R1171_U325 , R1171_U326 , R1171_U327 , R1171_U328;
wire R1171_U329 , R1171_U330 , R1171_U331 , R1171_U332 , R1171_U333 , R1171_U334 , R1171_U335 , R1171_U336 , R1171_U337 , R1171_U338;
wire R1171_U339 , R1171_U340 , R1171_U341 , R1171_U342 , R1171_U343 , R1171_U344 , R1171_U345 , R1171_U346 , R1171_U347 , R1171_U348;
wire R1171_U349 , R1171_U350 , R1171_U351 , R1171_U352 , R1171_U353 , R1171_U354 , R1171_U355 , R1171_U356 , R1171_U357 , R1171_U358;
wire R1171_U359 , R1171_U360 , R1171_U361 , R1171_U362 , R1171_U363 , R1171_U364 , R1171_U365 , R1171_U366 , R1171_U367 , R1171_U368;
wire R1171_U369 , R1171_U370 , R1171_U371 , R1171_U372 , R1171_U373 , R1171_U374 , R1171_U375 , R1171_U376 , R1171_U377 , R1171_U378;
wire R1171_U379 , R1171_U380 , R1171_U381 , R1171_U382 , R1171_U383 , R1171_U384 , R1171_U385 , R1171_U386 , R1171_U387 , R1171_U388;
wire R1171_U389 , R1171_U390 , R1171_U391 , R1171_U392 , R1171_U393 , R1171_U394 , R1171_U395 , R1171_U396 , R1171_U397 , R1171_U398;
wire R1171_U399 , R1171_U400 , R1171_U401 , R1171_U402 , R1171_U403 , R1171_U404 , R1171_U405 , R1171_U406 , R1171_U407 , R1171_U408;
wire R1171_U409 , R1171_U410 , R1171_U411 , R1171_U412 , R1171_U413 , R1171_U414 , R1171_U415 , R1171_U416 , R1171_U417 , R1171_U418;
wire R1171_U419 , R1171_U420 , R1171_U421 , R1171_U422 , R1171_U423 , R1171_U424 , R1171_U425 , R1171_U426 , R1171_U427 , R1171_U428;
wire R1171_U429 , R1171_U430 , R1171_U431 , R1171_U432 , R1171_U433 , R1171_U434 , R1171_U435 , R1171_U436 , R1171_U437 , R1171_U438;
wire R1171_U439 , R1171_U440 , R1171_U441 , R1171_U442 , R1171_U443 , R1171_U444 , R1171_U445 , R1171_U446 , R1171_U447 , R1171_U448;
wire R1171_U449 , R1171_U450 , R1171_U451 , R1171_U452 , R1171_U453 , R1171_U454 , R1171_U455 , R1171_U456 , R1171_U457 , R1171_U458;
wire R1171_U459 , R1171_U460 , R1171_U461 , R1171_U462 , R1171_U463 , R1171_U464 , R1171_U465 , R1171_U466 , R1171_U467 , R1171_U468;
wire R1171_U469 , R1171_U470 , R1171_U471 , R1171_U472 , R1171_U473 , R1171_U474 , R1171_U475 , R1171_U476 , R1171_U477 , R1171_U478;
wire R1171_U479 , R1171_U480 , R1171_U481 , R1171_U482 , R1171_U483 , R1171_U484 , R1171_U485 , R1171_U486 , R1171_U487 , R1171_U488;
wire R1171_U489 , R1171_U490 , R1171_U491 , R1171_U492 , R1171_U493 , R1171_U494 , R1171_U495 , R1171_U496 , R1171_U497 , R1171_U498;
wire R1171_U499 , R1171_U500 , R1171_U501 , R1171_U502 , R1171_U503 , R1171_U504 , R1171_U505 , R1171_U506 , R1171_U507 , R1171_U508;
wire R1171_U509 , R1171_U510 , R1171_U511 , R1171_U512 , R1171_U513 , R1171_U514 , R1171_U515 , R1171_U516 , R1171_U517 , R1171_U518;
wire R1171_U519 , R1171_U520 , R1171_U521 , R1171_U522 , R1171_U523 , R1171_U524 , R1171_U525 , R1171_U526 , R1171_U527 , R1171_U528;
wire R1171_U529 , R1171_U530 , R1171_U531 , R1138_U4 , R1138_U5 , R1138_U6 , R1138_U7 , R1138_U8 , R1138_U9 , R1138_U10;
wire R1138_U11 , R1138_U12 , R1138_U13 , R1138_U14 , R1138_U15 , R1138_U16 , R1138_U17 , R1138_U18 , R1138_U19 , R1138_U20;
wire R1138_U21 , R1138_U22 , R1138_U23 , R1138_U24 , R1138_U25 , R1138_U26 , R1138_U27 , R1138_U28 , R1138_U29 , R1138_U30;
wire R1138_U31 , R1138_U32 , R1138_U33 , R1138_U34 , R1138_U35 , R1138_U36 , R1138_U37 , R1138_U38 , R1138_U39 , R1138_U40;
wire R1138_U41 , R1138_U42 , R1138_U43 , R1138_U44 , R1138_U45 , R1138_U46 , R1138_U47 , R1138_U48 , R1138_U49 , R1138_U50;
wire R1138_U51 , R1138_U52 , R1138_U53 , R1138_U54 , R1138_U55 , R1138_U56 , R1138_U57 , R1138_U58 , R1138_U59 , R1138_U60;
wire R1138_U61 , R1138_U62 , R1138_U63 , R1138_U64 , R1138_U65 , R1138_U66 , R1138_U67 , R1138_U68 , R1138_U69 , R1138_U70;
wire R1138_U71 , R1138_U72 , R1138_U73 , R1138_U74 , R1138_U75 , R1138_U76 , R1138_U77 , R1138_U78 , R1138_U79 , R1138_U80;
wire R1138_U81 , R1138_U82 , R1138_U83 , R1138_U84 , R1138_U85 , R1138_U86 , R1138_U87 , R1138_U88 , R1138_U89 , R1138_U90;
wire R1138_U91 , R1138_U92 , R1138_U93 , R1138_U94 , R1138_U95 , R1138_U96 , R1138_U97 , R1138_U98 , R1138_U99 , R1138_U100;
wire R1138_U101 , R1138_U102 , R1138_U103 , R1138_U104 , R1138_U105 , R1138_U106 , R1138_U107 , R1138_U108 , R1138_U109 , R1138_U110;
wire R1138_U111 , R1138_U112 , R1138_U113 , R1138_U114 , R1138_U115 , R1138_U116 , R1138_U117 , R1138_U118 , R1138_U119 , R1138_U120;
wire R1138_U121 , R1138_U122 , R1138_U123 , R1138_U124 , R1138_U125 , R1138_U126 , R1138_U127 , R1138_U128 , R1138_U129 , R1138_U130;
wire R1138_U131 , R1138_U132 , R1138_U133 , R1138_U134 , R1138_U135 , R1138_U136 , R1138_U137 , R1138_U138 , R1138_U139 , R1138_U140;
wire R1138_U141 , R1138_U142 , R1138_U143 , R1138_U144 , R1138_U145 , R1138_U146 , R1138_U147 , R1138_U148 , R1138_U149 , R1138_U150;
wire R1138_U151 , R1138_U152 , R1138_U153 , R1138_U154 , R1138_U155 , R1138_U156 , R1138_U157 , R1138_U158 , R1138_U159 , R1138_U160;
wire R1138_U161 , R1138_U162 , R1138_U163 , R1138_U164 , R1138_U165 , R1138_U166 , R1138_U167 , R1138_U168 , R1138_U169 , R1138_U170;
wire R1138_U171 , R1138_U172 , R1138_U173 , R1138_U174 , R1138_U175 , R1138_U176 , R1138_U177 , R1138_U178 , R1138_U179 , R1138_U180;
wire R1138_U181 , R1138_U182 , R1138_U183 , R1138_U184 , R1138_U185 , R1138_U186 , R1138_U187 , R1138_U188 , R1138_U189 , R1138_U190;
wire R1138_U191 , R1138_U192 , R1138_U193 , R1138_U194 , R1138_U195 , R1138_U196 , R1138_U197 , R1138_U198 , R1138_U199 , R1138_U200;
wire R1138_U201 , R1138_U202 , R1138_U203 , R1138_U204 , R1138_U205 , R1138_U206 , R1138_U207 , R1138_U208 , R1138_U209 , R1138_U210;
wire R1138_U211 , R1138_U212 , R1138_U213 , R1138_U214 , R1138_U215 , R1138_U216 , R1138_U217 , R1138_U218 , R1138_U219 , R1138_U220;
wire R1138_U221 , R1138_U222 , R1138_U223 , R1138_U224 , R1138_U225 , R1138_U226 , R1138_U227 , R1138_U228 , R1138_U229 , R1138_U230;
wire R1138_U231 , R1138_U232 , R1138_U233 , R1138_U234 , R1138_U235 , R1138_U236 , R1138_U237 , R1138_U238 , R1138_U239 , R1138_U240;
wire R1138_U241 , R1138_U242 , R1138_U243 , R1138_U244 , R1138_U245 , R1138_U246 , R1138_U247 , R1138_U248 , R1138_U249 , R1138_U250;
wire R1138_U251 , R1138_U252 , R1138_U253 , R1138_U254 , R1138_U255 , R1138_U256 , R1138_U257 , R1138_U258 , R1138_U259 , R1138_U260;
wire R1138_U261 , R1138_U262 , R1138_U263 , R1138_U264 , R1138_U265 , R1138_U266 , R1138_U267 , R1138_U268 , R1138_U269 , R1138_U270;
wire R1138_U271 , R1138_U272 , R1138_U273 , R1138_U274 , R1138_U275 , R1138_U276 , R1138_U277 , R1138_U278 , R1138_U279 , R1138_U280;
wire R1138_U281 , R1138_U282 , R1138_U283 , R1138_U284 , R1138_U285 , R1138_U286 , R1138_U287 , R1138_U288 , R1138_U289 , R1138_U290;
wire R1138_U291 , R1138_U292 , R1138_U293 , R1138_U294 , R1138_U295 , R1138_U296 , R1138_U297 , R1138_U298 , R1138_U299 , R1138_U300;
wire R1138_U301 , R1138_U302 , R1138_U303 , R1138_U304 , R1138_U305 , R1138_U306 , R1138_U307 , R1138_U308 , R1138_U309 , R1138_U310;
wire R1138_U311 , R1138_U312 , R1138_U313 , R1138_U314 , R1138_U315 , R1138_U316 , R1138_U317 , R1138_U318 , R1138_U319 , R1138_U320;
wire R1138_U321 , R1138_U322 , R1138_U323 , R1138_U324 , R1138_U325 , R1138_U326 , R1138_U327 , R1138_U328 , R1138_U329 , R1138_U330;
wire R1138_U331 , R1138_U332 , R1138_U333 , R1138_U334 , R1138_U335 , R1138_U336 , R1138_U337 , R1138_U338 , R1138_U339 , R1138_U340;
wire R1138_U341 , R1138_U342 , R1138_U343 , R1138_U344 , R1138_U345 , R1138_U346 , R1138_U347 , R1138_U348 , R1138_U349 , R1138_U350;
wire R1138_U351 , R1138_U352 , R1138_U353 , R1138_U354 , R1138_U355 , R1138_U356 , R1138_U357 , R1138_U358 , R1138_U359 , R1138_U360;
wire R1138_U361 , R1138_U362 , R1138_U363 , R1138_U364 , R1138_U365 , R1138_U366 , R1138_U367 , R1138_U368 , R1138_U369 , R1138_U370;
wire R1138_U371 , R1138_U372 , R1138_U373 , R1138_U374 , R1138_U375 , R1138_U376 , R1138_U377 , R1138_U378 , R1138_U379 , R1138_U380;
wire R1138_U381 , R1138_U382 , R1138_U383 , R1138_U384 , R1138_U385 , R1138_U386 , R1138_U387 , R1138_U388 , R1138_U389 , R1138_U390;
wire R1138_U391 , R1138_U392 , R1138_U393 , R1138_U394 , R1138_U395 , R1138_U396 , R1138_U397 , R1138_U398 , R1138_U399 , R1138_U400;
wire R1138_U401 , R1138_U402 , R1138_U403 , R1138_U404 , R1138_U405 , R1138_U406 , R1138_U407 , R1138_U408 , R1138_U409 , R1138_U410;
wire R1138_U411 , R1138_U412 , R1138_U413 , R1138_U414 , R1138_U415 , R1138_U416 , R1138_U417 , R1138_U418 , R1138_U419 , R1138_U420;
wire R1138_U421 , R1138_U422 , R1138_U423 , R1138_U424 , R1138_U425 , R1138_U426 , R1138_U427 , R1138_U428 , R1138_U429 , R1138_U430;
wire R1138_U431 , R1138_U432 , R1138_U433 , R1138_U434 , R1138_U435 , R1138_U436 , R1138_U437 , R1138_U438 , R1138_U439 , R1138_U440;
wire R1138_U441 , R1138_U442 , R1138_U443 , R1138_U444 , R1138_U445 , R1138_U446 , R1138_U447 , R1138_U448 , R1138_U449 , R1138_U450;
wire R1138_U451 , R1138_U452 , R1138_U453 , R1138_U454 , R1138_U455 , R1138_U456 , R1138_U457 , R1138_U458 , R1138_U459 , R1138_U460;
wire R1138_U461 , R1138_U462 , R1138_U463 , R1138_U464 , R1138_U465 , R1138_U466 , R1138_U467 , R1138_U468 , R1138_U469 , R1138_U470;
wire R1138_U471 , R1138_U472 , R1138_U473 , R1138_U474 , R1138_U475 , R1138_U476 , R1138_U477 , R1138_U478 , R1138_U479 , R1138_U480;
wire R1138_U481 , R1138_U482 , R1138_U483 , R1138_U484 , R1138_U485 , R1138_U486 , R1138_U487 , R1138_U488 , R1138_U489 , R1138_U490;
wire R1138_U491 , R1138_U492 , R1138_U493 , R1138_U494 , R1138_U495 , R1138_U496 , R1138_U497 , R1138_U498 , R1138_U499 , R1138_U500;
wire R1138_U501 , R1138_U502 , R1138_U503 , R1138_U504 , R1138_U505 , R1138_U506 , R1138_U507 , R1138_U508 , R1138_U509 , R1138_U510;
wire R1138_U511 , R1138_U512 , R1138_U513 , R1138_U514 , R1138_U515 , R1138_U516 , R1138_U517 , R1138_U518 , R1138_U519 , R1138_U520;
wire R1138_U521 , R1138_U522 , R1138_U523 , R1138_U524 , R1138_U525 , R1138_U526 , R1138_U527 , R1138_U528 , R1138_U529 , R1138_U530;
wire R1138_U531 , R1222_U4 , R1222_U5 , R1222_U6 , R1222_U7 , R1222_U8 , R1222_U9 , R1222_U10 , R1222_U11 , R1222_U12;
wire R1222_U13 , R1222_U14 , R1222_U15 , R1222_U16 , R1222_U17 , R1222_U18 , R1222_U19 , R1222_U20 , R1222_U21 , R1222_U22;
wire R1222_U23 , R1222_U24 , R1222_U25 , R1222_U26 , R1222_U27 , R1222_U28 , R1222_U29 , R1222_U30 , R1222_U31 , R1222_U32;
wire R1222_U33 , R1222_U34 , R1222_U35 , R1222_U36 , R1222_U37 , R1222_U38 , R1222_U39 , R1222_U40 , R1222_U41 , R1222_U42;
wire R1222_U43 , R1222_U44 , R1222_U45 , R1222_U46 , R1222_U47 , R1222_U48 , R1222_U49 , R1222_U50 , R1222_U51 , R1222_U52;
wire R1222_U53 , R1222_U54 , R1222_U55 , R1222_U56 , R1222_U57 , R1222_U58 , R1222_U59 , R1222_U60 , R1222_U61 , R1222_U62;
wire R1222_U63 , R1222_U64 , R1222_U65 , R1222_U66 , R1222_U67 , R1222_U68 , R1222_U69 , R1222_U70 , R1222_U71 , R1222_U72;
wire R1222_U73 , R1222_U74 , R1222_U75 , R1222_U76 , R1222_U77 , R1222_U78 , R1222_U79 , R1222_U80 , R1222_U81 , R1222_U82;
wire R1222_U83 , R1222_U84 , R1222_U85 , R1222_U86 , R1222_U87 , R1222_U88 , R1222_U89 , R1222_U90 , R1222_U91 , R1222_U92;
wire R1222_U93 , R1222_U94 , R1222_U95 , R1222_U96 , R1222_U97 , R1222_U98 , R1222_U99 , R1222_U100 , R1222_U101 , R1222_U102;
wire R1222_U103 , R1222_U104 , R1222_U105 , R1222_U106 , R1222_U107 , R1222_U108 , R1222_U109 , R1222_U110 , R1222_U111 , R1222_U112;
wire R1222_U113 , R1222_U114 , R1222_U115 , R1222_U116 , R1222_U117 , R1222_U118 , R1222_U119 , R1222_U120 , R1222_U121 , R1222_U122;
wire R1222_U123 , R1222_U124 , R1222_U125 , R1222_U126 , R1222_U127 , R1222_U128 , R1222_U129 , R1222_U130 , R1222_U131 , R1222_U132;
wire R1222_U133 , R1222_U134 , R1222_U135 , R1222_U136 , R1222_U137 , R1222_U138 , R1222_U139 , R1222_U140 , R1222_U141 , R1222_U142;
wire R1222_U143 , R1222_U144 , R1222_U145 , R1222_U146 , R1222_U147 , R1222_U148 , R1222_U149 , R1222_U150 , R1222_U151 , R1222_U152;
wire R1222_U153 , R1222_U154 , R1222_U155 , R1222_U156 , R1222_U157 , R1222_U158 , R1222_U159 , R1222_U160 , R1222_U161 , R1222_U162;
wire R1222_U163 , R1222_U164 , R1222_U165 , R1222_U166 , R1222_U167 , R1222_U168 , R1222_U169 , R1222_U170 , R1222_U171 , R1222_U172;
wire R1222_U173 , R1222_U174 , R1222_U175 , R1222_U176 , R1222_U177 , R1222_U178 , R1222_U179 , R1222_U180 , R1222_U181 , R1222_U182;
wire R1222_U183 , R1222_U184 , R1222_U185 , R1222_U186 , R1222_U187 , R1222_U188 , R1222_U189 , R1222_U190 , R1222_U191 , R1222_U192;
wire R1222_U193 , R1222_U194 , R1222_U195 , R1222_U196 , R1222_U197 , R1222_U198 , R1222_U199 , R1222_U200 , R1222_U201 , R1222_U202;
wire R1222_U203 , R1222_U204 , R1222_U205 , R1222_U206 , R1222_U207 , R1222_U208 , R1222_U209 , R1222_U210 , R1222_U211 , R1222_U212;
wire R1222_U213 , R1222_U214 , R1222_U215 , R1222_U216 , R1222_U217 , R1222_U218 , R1222_U219 , R1222_U220 , R1222_U221 , R1222_U222;
wire R1222_U223 , R1222_U224 , R1222_U225 , R1222_U226 , R1222_U227 , R1222_U228 , R1222_U229 , R1222_U230 , R1222_U231 , R1222_U232;
wire R1222_U233 , R1222_U234 , R1222_U235 , R1222_U236 , R1222_U237 , R1222_U238 , R1222_U239 , R1222_U240 , R1222_U241 , R1222_U242;
wire R1222_U243 , R1222_U244 , R1222_U245 , R1222_U246 , R1222_U247 , R1222_U248 , R1222_U249 , R1222_U250 , R1222_U251 , R1222_U252;
wire R1222_U253 , R1222_U254 , R1222_U255 , R1222_U256 , R1222_U257 , R1222_U258 , R1222_U259 , R1222_U260 , R1222_U261 , R1222_U262;
wire R1222_U263 , R1222_U264 , R1222_U265 , R1222_U266 , R1222_U267 , R1222_U268 , R1222_U269 , R1222_U270 , R1222_U271 , R1222_U272;
wire R1222_U273 , R1222_U274 , R1222_U275 , R1222_U276 , R1222_U277 , R1222_U278 , R1222_U279 , R1222_U280 , R1222_U281 , R1222_U282;
wire R1222_U283 , R1222_U284 , R1222_U285 , R1222_U286 , R1222_U287 , R1222_U288 , R1222_U289 , R1222_U290 , R1222_U291 , R1222_U292;
wire R1222_U293 , R1222_U294 , R1222_U295 , R1222_U296 , R1222_U297 , R1222_U298 , R1222_U299 , R1222_U300 , R1222_U301 , R1222_U302;
wire R1222_U303 , R1222_U304 , R1222_U305 , R1222_U306 , R1222_U307 , R1222_U308 , R1222_U309 , R1222_U310 , R1222_U311 , R1222_U312;
wire R1222_U313 , R1222_U314 , R1222_U315 , R1222_U316 , R1222_U317 , R1222_U318 , R1222_U319 , R1222_U320 , R1222_U321 , R1222_U322;
wire R1222_U323 , R1222_U324 , R1222_U325 , R1222_U326 , R1222_U327 , R1222_U328 , R1222_U329 , R1222_U330 , R1222_U331 , R1222_U332;
wire R1222_U333 , R1222_U334 , R1222_U335 , R1222_U336 , R1222_U337 , R1222_U338 , R1222_U339 , R1222_U340 , R1222_U341 , R1222_U342;
wire R1222_U343 , R1222_U344 , R1222_U345 , R1222_U346 , R1222_U347 , R1222_U348 , R1222_U349 , R1222_U350 , R1222_U351 , R1222_U352;
wire R1222_U353 , R1222_U354 , R1222_U355 , R1222_U356 , R1222_U357 , R1222_U358 , R1222_U359 , R1222_U360 , R1222_U361 , R1222_U362;
wire R1222_U363 , R1222_U364 , R1222_U365 , R1222_U366 , R1222_U367 , R1222_U368 , R1222_U369 , R1222_U370 , R1222_U371 , R1222_U372;
wire R1222_U373 , R1222_U374 , R1222_U375 , R1222_U376 , R1222_U377 , R1222_U378 , R1222_U379 , R1222_U380 , R1222_U381 , R1222_U382;
wire R1222_U383 , R1222_U384 , R1222_U385 , R1222_U386 , R1222_U387 , R1222_U388 , R1222_U389 , R1222_U390 , R1222_U391 , R1222_U392;
wire R1222_U393 , R1222_U394 , R1222_U395 , R1222_U396 , R1222_U397 , R1222_U398 , R1222_U399 , R1222_U400 , R1222_U401 , R1222_U402;
wire R1222_U403 , R1222_U404 , R1222_U405 , R1222_U406 , R1222_U407 , R1222_U408 , R1222_U409 , R1222_U410 , R1222_U411 , R1222_U412;
wire R1222_U413 , R1222_U414 , R1222_U415 , R1222_U416 , R1222_U417 , R1222_U418 , R1222_U419 , R1222_U420 , R1222_U421 , R1222_U422;
wire R1222_U423 , R1222_U424 , R1222_U425 , R1222_U426 , R1222_U427 , R1222_U428 , R1222_U429 , R1222_U430 , R1222_U431 , R1222_U432;
wire R1222_U433 , R1222_U434 , R1222_U435 , R1222_U436 , R1222_U437 , R1222_U438 , R1222_U439 , R1222_U440 , R1222_U441 , R1222_U442;
wire R1222_U443 , R1222_U444 , R1222_U445 , R1222_U446 , R1222_U447 , R1222_U448 , R1222_U449 , R1222_U450 , R1222_U451 , R1222_U452;
wire R1222_U453 , R1222_U454 , R1222_U455 , R1222_U456 , R1222_U457 , R1222_U458 , R1222_U459 , R1222_U460 , R1222_U461 , R1222_U462;
wire R1222_U463 , R1222_U464 , R1222_U465 , R1222_U466 , R1222_U467 , R1222_U468 , R1222_U469 , R1222_U470 , R1222_U471 , R1222_U472;
wire R1222_U473 , R1222_U474 , R1222_U475 , R1222_U476 , R1222_U477 , R1222_U478 , R1222_U479 , R1222_U480 , R1222_U481 , R1222_U482;
wire R1222_U483 , R1222_U484 , R1222_U485 , R1222_U486 , R1222_U487 , R1222_U488 , R1222_U489 , R1222_U490 , R1222_U491 , R1222_U492;
wire R1222_U493 , R1222_U494;


nand NAND2_1 ( R1222_U519 , U3464 , R1222_U42 );
nand NAND2_2 ( R1222_U518 , U3074 , R1222_U41 );
nand NAND2_3 ( R1222_U517 , U3486 , R1222_U71 );
and AND2_4 ( U3014 , U4201 , U3431 );
and AND2_5 ( U3015 , U4011 , U3456 );
and AND2_6 ( U3016 , U3454 , U3455 );
and AND2_7 ( U3017 , U3659 , U3654 );
and AND2_8 ( U3018 , U3462 , U3463 );
and AND2_9 ( U3019 , U5826 , U3462 );
and AND2_10 ( U3020 , U5823 , U3463 );
and AND2_11 ( U3021 , U5823 , U5826 );
and AND2_12 ( U3022 , U5613 , U3355 );
and AND2_13 ( U3023 , U3047 , STATE_REG );
and AND3_14 ( U3024 , U5820 , U5805 , U5808 );
and AND2_15 ( U3025 , U3845 , U3421 );
and AND2_16 ( U3026 , U4042 , U5799 );
and AND2_17 ( U3027 , U4010 , U5820 );
and AND2_18 ( U3028 , U3908 , U4028 );
and AND2_19 ( U3029 , U3357 , STATE_REG );
and AND2_20 ( U3030 , U4019 , U4044 );
and AND2_21 ( U3031 , U4044 , U4021 );
and AND2_22 ( U3032 , U4012 , U4044 );
and AND2_23 ( U3033 , U4020 , U4044 );
and AND2_24 ( U3034 , U4042 , U3454 );
and AND2_25 ( U3035 , U4028 , U5799 );
and AND2_26 ( U3036 , U4044 , U3026 );
and AND2_27 ( U3037 , U4028 , U3454 );
and AND2_28 ( U3038 , U5802 , U4938 );
and AND2_29 ( U3039 , U3025 , U5802 );
and AND2_30 ( U3040 , U5799 , U4938 );
and AND2_31 ( U3041 , U3025 , U5799 );
and AND2_32 ( U3042 , U3016 , U4938 );
and AND2_33 ( U3043 , U3025 , U3016 );
and AND2_34 ( U3044 , U3023 , U3421 );
and AND2_35 ( U3045 , U5170 , STATE_REG );
and AND2_36 ( U3046 , U3023 , U5172 );
and AND2_37 ( U3047 , U5748 , U3355 );
and AND2_38 ( U3048 , U3660 , U3017 );
and AND5_39 ( U3049 , U4759 , U4758 , U4762 , U4766 , U4765 );
nand NAND4_40 ( U3050 , U4696 , U4697 , U4695 , U4698 );
nand NAND4_41 ( U3051 , U4715 , U4716 , U4714 , U4717 );
nand NAND4_42 ( U3052 , U4736 , U4735 , U4734 , U4733 );
nand NAND3_43 ( U3053 , U4773 , U4774 , U4772 );
nand NAND4_44 ( U3054 , U4677 , U4678 , U4676 , U4679 );
nand NAND4_45 ( U3055 , U4658 , U4659 , U4657 , U4660 );
nand NAND3_46 ( U3056 , U4753 , U4754 , U4752 );
nand NAND4_47 ( U3057 , U4261 , U4260 , U4259 , U4258 );
nand NAND4_48 ( U3058 , U4601 , U4602 , U4600 , U4603 );
nand NAND4_49 ( U3059 , U4375 , U4374 , U4373 , U4372 );
nand NAND4_50 ( U3060 , U4394 , U4393 , U4392 , U4391 );
nand NAND4_51 ( U3061 , U4242 , U4241 , U4240 , U4239 );
nand NAND4_52 ( U3062 , U4639 , U4640 , U4638 , U4641 );
nand NAND4_53 ( U3063 , U4620 , U4621 , U4619 , U4622 );
nand NAND4_54 ( U3064 , U4280 , U4279 , U4278 , U4277 );
nand NAND4_55 ( U3065 , U4218 , U4217 , U4216 , U4215 );
nand NAND4_56 ( U3066 , U4508 , U4507 , U4506 , U4505 );
nand NAND4_57 ( U3067 , U4318 , U4317 , U4316 , U4315 );
nand NAND4_58 ( U3068 , U4299 , U4298 , U4297 , U4296 );
nand NAND4_59 ( U3069 , U4413 , U4412 , U4411 , U4410 );
nand NAND4_60 ( U3070 , U4489 , U4488 , U4487 , U4486 );
nand NAND4_61 ( U3071 , U4470 , U4469 , U4468 , U4467 );
nand NAND4_62 ( U3072 , U4582 , U4583 , U4581 , U4584 );
nand NAND4_63 ( U3073 , U4565 , U4564 , U4563 , U4562 );
nand NAND4_64 ( U3074 , U4223 , U4222 , U4221 , U4220 );
nand NAND4_65 ( U3075 , U4199 , U4198 , U4197 , U4196 );
nand NAND4_66 ( U3076 , U4451 , U4450 , U4449 , U4448 );
nand NAND4_67 ( U3077 , U4432 , U4431 , U4430 , U4429 );
nand NAND4_68 ( U3078 , U4546 , U4545 , U4544 , U4543 );
nand NAND4_69 ( U3079 , U4527 , U4526 , U4525 , U4524 );
nand NAND4_70 ( U3080 , U4356 , U4355 , U4354 , U4353 );
nand NAND4_71 ( U3081 , U4337 , U4336 , U4335 , U4334 );
nand NAND2_72 ( U3082 , U5538 , U5537 );
nand NAND2_73 ( U3083 , U5540 , U5539 );
nand NAND3_74 ( U3084 , U5545 , U5544 , U5546 );
nand NAND3_75 ( U3085 , U5548 , U5547 , U5549 );
nand NAND3_76 ( U3086 , U5552 , U5550 , U5551 );
nand NAND3_77 ( U3087 , U5554 , U5553 , U5555 );
nand NAND3_78 ( U3088 , U5558 , U5556 , U5557 );
nand NAND3_79 ( U3089 , U5560 , U5559 , U5561 );
nand NAND3_80 ( U3090 , U5564 , U5562 , U5563 );
nand NAND3_81 ( U3091 , U5566 , U5565 , U5567 );
nand NAND3_82 ( U3092 , U5570 , U5568 , U5569 );
nand NAND3_83 ( U3093 , U5572 , U5571 , U5573 );
nand NAND3_84 ( U3094 , U5579 , U5577 , U5578 );
nand NAND3_85 ( U3095 , U5581 , U5580 , U5582 );
nand NAND3_86 ( U3096 , U5584 , U5583 , U5585 );
nand NAND3_87 ( U3097 , U5587 , U5586 , U5588 );
nand NAND3_88 ( U3098 , U5590 , U5589 , U5591 );
nand NAND3_89 ( U3099 , U5593 , U5592 , U5594 );
nand NAND3_90 ( U3100 , U5596 , U5595 , U5597 );
nand NAND3_91 ( U3101 , U5599 , U5598 , U5600 );
nand NAND3_92 ( U3102 , U5602 , U5601 , U5603 );
nand NAND3_93 ( U3103 , U5605 , U5604 , U5606 );
nand NAND3_94 ( U3104 , U5520 , U5519 , U5521 );
nand NAND3_95 ( U3105 , U5523 , U5522 , U5524 );
nand NAND3_96 ( U3106 , U5526 , U5525 , U5527 );
nand NAND3_97 ( U3107 , U5529 , U5528 , U5530 );
nand NAND3_98 ( U3108 , U5532 , U5531 , U5533 );
nand NAND3_99 ( U3109 , U5535 , U5534 , U5536 );
nand NAND3_100 ( U3110 , U5542 , U5541 , U5543 );
nand NAND3_101 ( U3111 , U5575 , U5574 , U5576 );
nand NAND3_102 ( U3112 , U5608 , U5607 , U5609 );
nand NAND2_103 ( U3113 , U5611 , U5610 );
nand NAND2_104 ( U3114 , U3926 , U5441 );
nand NAND2_105 ( U3115 , U3927 , U5444 );
nand NAND2_106 ( U3116 , U5450 , U3929 );
nand NAND2_107 ( U3117 , U5453 , U3931 );
nand NAND2_108 ( U3118 , U5456 , U3933 );
nand NAND2_109 ( U3119 , U5459 , U3935 );
nand NAND2_110 ( U3120 , U5462 , U3937 );
nand NAND2_111 ( U3121 , U5465 , U3939 );
nand NAND2_112 ( U3122 , U5468 , U3941 );
nand NAND2_113 ( U3123 , U5471 , U3943 );
nand NAND2_114 ( U3124 , U5474 , U3945 );
nand NAND2_115 ( U3125 , U5477 , U3947 );
nand NAND2_116 ( U3126 , U5484 , U3950 );
nand NAND2_117 ( U3127 , U5487 , U3951 );
nand NAND2_118 ( U3128 , U5490 , U3952 );
nand NAND2_119 ( U3129 , U5493 , U3953 );
nand NAND2_120 ( U3130 , U5496 , U3954 );
nand NAND2_121 ( U3131 , U5499 , U3955 );
nand NAND2_122 ( U3132 , U5502 , U3956 );
nand NAND2_123 ( U3133 , U5505 , U3957 );
nand NAND2_124 ( U3134 , U5508 , U3958 );
nand NAND2_125 ( U3135 , U5511 , U3959 );
nand NAND2_126 ( U3136 , U5424 , U3920 );
nand NAND2_127 ( U3137 , U5427 , U3921 );
nand NAND2_128 ( U3138 , U5430 , U3922 );
nand NAND2_129 ( U3139 , U5433 , U3923 );
nand NAND2_130 ( U3140 , U5436 , U3924 );
nand NAND2_131 ( U3141 , U5439 , U3925 );
nand NAND2_132 ( U3142 , U5448 , U3928 );
nand NAND2_133 ( U3143 , U5481 , U3949 );
nand NAND2_134 ( U3144 , U5514 , U3960 );
nand NAND2_135 ( U3145 , U5517 , U3961 );
nand NAND2_136 ( U3146 , U4201 , U5748 );
nand NAND2_137 ( U3147 , U5808 , U3372 );
nand NAND2_138 ( U3148 , U4062 , STATE_REG );
not NOT1_139 ( U3149 , STATE_REG );
nand NAND2_140 ( U3150 , U5693 , U5692 );
nand NAND2_141 ( U3151 , U5695 , U5694 );
nand NAND2_142 ( U3152 , U5697 , U5696 );
nand NAND2_143 ( U3153 , U5699 , U5698 );
nand NAND2_144 ( U3154 , U5701 , U5700 );
nand NAND2_145 ( U3155 , U5703 , U5702 );
nand NAND2_146 ( U3156 , U5705 , U5704 );
nand NAND2_147 ( U3157 , U5707 , U5706 );
nand NAND2_148 ( U3158 , U5709 , U5708 );
nand NAND2_149 ( U3159 , U5713 , U5712 );
nand NAND2_150 ( U3160 , U5715 , U5714 );
nand NAND2_151 ( U3161 , U5717 , U5716 );
nand NAND2_152 ( U3162 , U5719 , U5718 );
nand NAND2_153 ( U3163 , U5721 , U5720 );
nand NAND2_154 ( U3164 , U5723 , U5722 );
nand NAND2_155 ( U3165 , U5725 , U5724 );
nand NAND2_156 ( U3166 , U5727 , U5726 );
nand NAND2_157 ( U3167 , U5729 , U5728 );
nand NAND2_158 ( U3168 , U5731 , U5730 );
nand NAND2_159 ( U3169 , U5679 , U5678 );
nand NAND2_160 ( U3170 , U5681 , U5680 );
nand NAND2_161 ( U3171 , U5683 , U5682 );
nand NAND2_162 ( U3172 , U5685 , U5684 );
nand NAND2_163 ( U3173 , U5687 , U5686 );
nand NAND2_164 ( U3174 , U5689 , U5688 );
nand NAND2_165 ( U3175 , U5691 , U5690 );
nand NAND2_166 ( U3176 , U5711 , U5710 );
nand NAND2_167 ( U3177 , U5733 , U5732 );
nand NAND2_168 ( U3178 , U3966 , U5735 );
nand NAND2_169 ( U3179 , U5634 , U5633 );
nand NAND2_170 ( U3180 , U5636 , U5635 );
nand NAND2_171 ( U3181 , U5638 , U5637 );
nand NAND2_172 ( U3182 , U5640 , U5639 );
nand NAND2_173 ( U3183 , U5642 , U5641 );
nand NAND2_174 ( U3184 , U5644 , U5643 );
nand NAND2_175 ( U3185 , U5646 , U5645 );
nand NAND2_176 ( U3186 , U5648 , U5647 );
nand NAND2_177 ( U3187 , U5650 , U5649 );
nand NAND2_178 ( U3188 , U5654 , U5653 );
nand NAND2_179 ( U3189 , U5656 , U5655 );
nand NAND2_180 ( U3190 , U5658 , U5657 );
nand NAND2_181 ( U3191 , U5660 , U5659 );
nand NAND2_182 ( U3192 , U5662 , U5661 );
nand NAND2_183 ( U3193 , U5664 , U5663 );
nand NAND2_184 ( U3194 , U5666 , U5665 );
nand NAND2_185 ( U3195 , U5668 , U5667 );
nand NAND2_186 ( U3196 , U5670 , U5669 );
nand NAND2_187 ( U3197 , U5672 , U5671 );
nand NAND2_188 ( U3198 , U5620 , U5619 );
nand NAND2_189 ( U3199 , U5622 , U5621 );
nand NAND2_190 ( U3200 , U5624 , U5623 );
nand NAND2_191 ( U3201 , U5626 , U5625 );
nand NAND2_192 ( U3202 , U5628 , U5627 );
nand NAND2_193 ( U3203 , U5630 , U5629 );
nand NAND2_194 ( U3204 , U5632 , U5631 );
nand NAND2_195 ( U3205 , U5652 , U5651 );
nand NAND2_196 ( U3206 , U5674 , U5673 );
nand NAND2_197 ( U3207 , U3965 , U5675 );
and AND2_198 ( U3208 , U5612 , U3355 );
nand NAND3_199 ( U3209 , U6259 , U6258 , U5422 );
nand NAND5_200 ( U3210 , U5416 , U5415 , U5419 , U5417 , U5418 );
nand NAND5_201 ( U3211 , U5407 , U5406 , U5410 , U5408 , U5409 );
nand NAND5_202 ( U3212 , U5398 , U5397 , U5401 , U5399 , U5400 );
nand NAND5_203 ( U3213 , U5389 , U5388 , U5392 , U5390 , U5391 );
nand NAND5_204 ( U3214 , U5380 , U5379 , U5383 , U5381 , U5382 );
nand NAND3_205 ( U3215 , U3918 , U5371 , U5372 );
nand NAND5_206 ( U3216 , U5362 , U5361 , U5365 , U5363 , U5364 );
nand NAND5_207 ( U3217 , U5353 , U5352 , U5356 , U5354 , U5355 );
nand NAND5_208 ( U3218 , U5344 , U5343 , U5347 , U5345 , U5346 );
nand NAND3_209 ( U3219 , U3916 , U5335 , U5336 );
nand NAND5_210 ( U3220 , U5326 , U5325 , U5329 , U5327 , U5328 );
nand NAND5_211 ( U3221 , U5317 , U5316 , U5320 , U5318 , U5319 );
nand NAND5_212 ( U3222 , U5308 , U5307 , U5311 , U5309 , U5310 );
nand NAND5_213 ( U3223 , U5299 , U5298 , U5302 , U5300 , U5301 );
nand NAND4_214 ( U3224 , U5290 , U5289 , U5291 , U3915 );
nand NAND5_215 ( U3225 , U5281 , U5280 , U5284 , U5282 , U5283 );
nand NAND5_216 ( U3226 , U5272 , U5271 , U5275 , U5273 , U5274 );
nand NAND4_217 ( U3227 , U5263 , U5262 , U3914 , U5264 );
nand NAND5_218 ( U3228 , U5254 , U5253 , U5257 , U5255 , U5256 );
nand NAND3_219 ( U3229 , U3913 , U5246 , U3912 );
nand NAND5_220 ( U3230 , U5237 , U5236 , U5240 , U5238 , U5239 );
nand NAND5_221 ( U3231 , U5228 , U5227 , U5231 , U5229 , U5230 );
nand NAND5_222 ( U3232 , U5219 , U5218 , U5222 , U5220 , U5221 );
nand NAND5_223 ( U3233 , U5210 , U5209 , U5213 , U5211 , U5212 );
nand NAND3_224 ( U3234 , U3909 , U5201 , U5202 );
nand NAND5_225 ( U3235 , U5192 , U5191 , U5195 , U5193 , U5194 );
nand NAND5_226 ( U3236 , U5183 , U5182 , U5186 , U5184 , U5185 );
nand NAND5_227 ( U3237 , U5174 , U5173 , U5177 , U5175 , U5176 );
nand NAND5_228 ( U3238 , U5161 , U5160 , U5164 , U5162 , U5163 );
nand NAND2_229 ( U3239 , U3904 , U5147 );
nand NAND2_230 ( U3240 , U3890 , U3889 );
nand NAND2_231 ( U3241 , U3888 , U3887 );
nand NAND2_232 ( U3242 , U3886 , U3885 );
nand NAND2_233 ( U3243 , U3883 , U3882 );
nand NAND2_234 ( U3244 , U3881 , U3880 );
nand NAND2_235 ( U3245 , U3878 , U3877 );
nand NAND2_236 ( U3246 , U3876 , U3875 );
nand NAND2_237 ( U3247 , U3874 , U3873 );
nand NAND4_238 ( U3248 , U3872 , U3871 , U5054 , U5050 );
nand NAND4_239 ( U3249 , U3870 , U3869 , U5044 , U5040 );
nand NAND4_240 ( U3250 , U3868 , U3867 , U5034 , U5030 );
nand NAND4_241 ( U3251 , U3866 , U3865 , U5024 , U5020 );
nand NAND4_242 ( U3252 , U3864 , U3863 , U5014 , U5010 );
nand NAND4_243 ( U3253 , U3862 , U3861 , U5004 , U5000 );
nand NAND4_244 ( U3254 , U3860 , U3859 , U4994 , U4990 );
nand NAND4_245 ( U3255 , U3858 , U3857 , U4984 , U4980 );
nand NAND4_246 ( U3256 , U3856 , U3855 , U4974 , U4970 );
nand NAND4_247 ( U3257 , U3854 , U3853 , U4964 , U4960 );
nand NAND2_248 ( U3258 , U3852 , U3850 );
nand NAND2_249 ( U3259 , U3848 , U3846 );
nand NAND3_250 ( U3260 , U4937 , U4936 , U4004 );
nand NAND3_251 ( U3261 , U4935 , U4934 , U4003 );
nand NAND4_252 ( U3262 , U3836 , U3837 , U4927 , U4000 );
nand NAND4_253 ( U3263 , U3834 , U3835 , U4922 , U3999 );
nand NAND4_254 ( U3264 , U3832 , U3833 , U4917 , U3998 );
nand NAND4_255 ( U3265 , U3830 , U3831 , U4912 , U3997 );
nand NAND4_256 ( U3266 , U3828 , U3829 , U4907 , U3996 );
nand NAND4_257 ( U3267 , U3826 , U3827 , U4902 , U3995 );
nand NAND4_258 ( U3268 , U3824 , U3825 , U4897 , U3994 );
nand NAND4_259 ( U3269 , U3822 , U3823 , U4892 , U3993 );
nand NAND4_260 ( U3270 , U3820 , U3821 , U4887 , U3992 );
nand NAND4_261 ( U3271 , U3818 , U3819 , U4882 , U3991 );
nand NAND4_262 ( U3272 , U3816 , U3817 , U4877 , U3990 );
nand NAND4_263 ( U3273 , U3814 , U3815 , U4872 , U3989 );
nand NAND4_264 ( U3274 , U3812 , U3813 , U4867 , U3988 );
nand NAND4_265 ( U3275 , U3810 , U3811 , U4862 , U3987 );
nand NAND3_266 ( U3276 , U3809 , U3808 , U3986 );
nand NAND4_267 ( U3277 , U3806 , U3807 , U4852 , U3985 );
nand NAND3_268 ( U3278 , U3805 , U3804 , U3984 );
nand NAND3_269 ( U3279 , U3803 , U3802 , U3983 );
nand NAND3_270 ( U3280 , U3801 , U3800 , U3982 );
nand NAND3_271 ( U3281 , U3799 , U3798 , U3981 );
nand NAND3_272 ( U3282 , U3797 , U3796 , U3980 );
nand NAND3_273 ( U3283 , U3795 , U3794 , U3979 );
nand NAND3_274 ( U3284 , U3793 , U3792 , U3978 );
nand NAND3_275 ( U3285 , U3791 , U3790 , U3977 );
nand NAND2_276 ( U3286 , U3789 , U3788 );
nand NAND2_277 ( U3287 , U3787 , U3786 );
nand NAND2_278 ( U3288 , U3785 , U3784 );
nand NAND2_279 ( U3289 , U3783 , U3782 );
nand NAND2_280 ( U3290 , U3781 , U3780 );
and AND2_281 ( U3291 , D_REG_31_ , U3968 );
and AND2_282 ( U3292 , D_REG_30_ , U3968 );
and AND2_283 ( U3293 , D_REG_29_ , U3968 );
and AND2_284 ( U3294 , D_REG_28_ , U3968 );
and AND2_285 ( U3295 , D_REG_27_ , U3968 );
and AND2_286 ( U3296 , D_REG_26_ , U3968 );
and AND2_287 ( U3297 , D_REG_25_ , U3968 );
and AND2_288 ( U3298 , D_REG_24_ , U3968 );
and AND2_289 ( U3299 , D_REG_23_ , U3968 );
and AND2_290 ( U3300 , D_REG_22_ , U3968 );
and AND2_291 ( U3301 , D_REG_21_ , U3968 );
and AND2_292 ( U3302 , D_REG_20_ , U3968 );
and AND2_293 ( U3303 , D_REG_19_ , U3968 );
and AND2_294 ( U3304 , D_REG_18_ , U3968 );
and AND2_295 ( U3305 , D_REG_17_ , U3968 );
and AND2_296 ( U3306 , D_REG_16_ , U3968 );
and AND2_297 ( U3307 , D_REG_15_ , U3968 );
and AND2_298 ( U3308 , D_REG_14_ , U3968 );
and AND2_299 ( U3309 , D_REG_13_ , U3968 );
and AND2_300 ( U3310 , D_REG_12_ , U3968 );
and AND2_301 ( U3311 , D_REG_11_ , U3968 );
and AND2_302 ( U3312 , D_REG_10_ , U3968 );
and AND2_303 ( U3313 , D_REG_9_ , U3968 );
and AND2_304 ( U3314 , D_REG_8_ , U3968 );
and AND2_305 ( U3315 , D_REG_7_ , U3968 );
and AND2_306 ( U3316 , D_REG_6_ , U3968 );
and AND2_307 ( U3317 , D_REG_5_ , U3968 );
and AND2_308 ( U3318 , D_REG_4_ , U3968 );
and AND2_309 ( U3319 , D_REG_3_ , U3968 );
and AND2_310 ( U3320 , D_REG_2_ , U3968 );
nand NAND2_311 ( U3321 , U3645 , U4159 );
nand NAND2_312 ( U3322 , U3644 , U4156 );
nand NAND2_313 ( U3323 , U3643 , U4153 );
nand NAND2_314 ( U3324 , U3642 , U4150 );
nand NAND2_315 ( U3325 , U3641 , U4147 );
nand NAND2_316 ( U3326 , U3640 , U4144 );
nand NAND2_317 ( U3327 , U3639 , U4141 );
nand NAND2_318 ( U3328 , U3638 , U4138 );
nand NAND2_319 ( U3329 , U3637 , U4135 );
nand NAND2_320 ( U3330 , U3636 , U4132 );
nand NAND2_321 ( U3331 , U3635 , U4129 );
nand NAND2_322 ( U3332 , U3634 , U4126 );
nand NAND2_323 ( U3333 , U3633 , U4123 );
nand NAND2_324 ( U3334 , U3632 , U4120 );
nand NAND2_325 ( U3335 , U3631 , U4117 );
nand NAND2_326 ( U3336 , U3630 , U4114 );
nand NAND2_327 ( U3337 , U3629 , U4111 );
nand NAND2_328 ( U3338 , U3628 , U4108 );
nand NAND2_329 ( U3339 , U3627 , U4105 );
nand NAND2_330 ( U3340 , U3626 , U4102 );
nand NAND2_331 ( U3341 , U3625 , U4099 );
nand NAND2_332 ( U3342 , U3624 , U4096 );
nand NAND2_333 ( U3343 , U3623 , U4093 );
nand NAND2_334 ( U3344 , U3622 , U4090 );
nand NAND2_335 ( U3345 , U3621 , U4087 );
nand NAND2_336 ( U3346 , U3620 , U4084 );
nand NAND2_337 ( U3347 , U3619 , U4081 );
nand NAND2_338 ( U3348 , U3618 , U4078 );
nand NAND2_339 ( U3349 , U3617 , U4075 );
nand NAND2_340 ( U3350 , U3616 , U4072 );
nand NAND2_341 ( U3351 , U3615 , U4069 );
nand NAND2_342 ( U3352 , U3614 , U4066 );
nand NAND2_343 ( U3353 , U4055 , U5805 );
nand NAND5_344 ( U3354 , U4932 , U4930 , U4933 , U4931 , U4001 );
nand NAND3_345 ( U3355 , U3433 , U3432 , U3434 );
nand NAND2_346 ( U3356 , U4059 , U5748 );
nand NAND2_347 ( U3357 , STATE_REG , U3967 );
nand NAND2_348 ( U3358 , U3432 , U5757 );
not NOT1_349 ( U3359 , B_REG );
nand NAND3_350 ( U3360 , U5810 , U5809 , U3432 );
nand NAND2_351 ( U3361 , U5820 , U3456 );
nand NAND2_352 ( U3362 , U4201 , U3461 );
nand NAND3_353 ( U3363 , U3461 , U3456 , U3460 );
nand NAND3_354 ( U3364 , U5817 , U3456 , U3460 );
nand NAND2_355 ( U3365 , U3460 , U3457 );
nand NAND2_356 ( U3366 , U4056 , U3461 );
nand NAND2_357 ( U3367 , U4056 , U5817 );
nand NAND2_358 ( U3368 , U4201 , U5817 );
nand NAND2_359 ( U3369 , U4015 , U5808 );
nand NAND3_360 ( U3370 , U5817 , U5820 , U3457 );
nand NAND2_361 ( U3371 , U4011 , U5805 );
nand NAND2_362 ( U3372 , U5805 , U3461 );
nand NAND2_363 ( U3373 , U3457 , U3456 );
nand NAND2_364 ( U3374 , U5808 , U3460 );
nand NAND5_365 ( U3375 , U4207 , U4206 , U4208 , U3647 , U3646 );
not NOT1_366 ( U3376 , REG2_REG_0_ );
nand NAND4_367 ( U3377 , U4226 , U4225 , U3662 , U3664 );
nand NAND4_368 ( U3378 , U4245 , U4244 , U3666 , U3668 );
nand NAND4_369 ( U3379 , U4264 , U4263 , U3670 , U3672 );
nand NAND4_370 ( U3380 , U4283 , U4282 , U3674 , U3676 );
nand NAND4_371 ( U3381 , U4302 , U4301 , U3678 , U3680 );
nand NAND4_372 ( U3382 , U4321 , U4320 , U3682 , U3684 );
nand NAND4_373 ( U3383 , U4340 , U4339 , U3686 , U3688 );
nand NAND4_374 ( U3384 , U4359 , U4358 , U3690 , U3692 );
nand NAND4_375 ( U3385 , U4378 , U4377 , U3694 , U3696 );
nand NAND4_376 ( U3386 , U4397 , U4396 , U3698 , U3700 );
nand NAND4_377 ( U3387 , U4416 , U4415 , U3702 , U3704 );
nand NAND4_378 ( U3388 , U4435 , U4434 , U3706 , U3708 );
nand NAND4_379 ( U3389 , U4454 , U4453 , U3710 , U3712 );
nand NAND4_380 ( U3390 , U4473 , U4472 , U3714 , U3716 );
nand NAND4_381 ( U3391 , U4492 , U4491 , U3718 , U3720 );
nand NAND4_382 ( U3392 , U4511 , U4510 , U3722 , U3724 );
nand NAND4_383 ( U3393 , U4530 , U4529 , U3726 , U3728 );
nand NAND4_384 ( U3394 , U4549 , U4548 , U3730 , U3732 );
nand NAND4_385 ( U3395 , U4568 , U4567 , U3734 , U3736 );
nand NAND2_386 ( U3396 , DATAI_20_ , U3969 );
nand NAND4_387 ( U3397 , U4587 , U4586 , U3738 , U3740 );
nand NAND2_388 ( U3398 , DATAI_21_ , U3969 );
nand NAND4_389 ( U3399 , U4606 , U4605 , U3742 , U3744 );
nand NAND2_390 ( U3400 , DATAI_22_ , U3969 );
nand NAND4_391 ( U3401 , U4625 , U4624 , U3746 , U3748 );
nand NAND2_392 ( U3402 , DATAI_23_ , U3969 );
nand NAND4_393 ( U3403 , U4644 , U4643 , U3750 , U3752 );
nand NAND2_394 ( U3404 , DATAI_24_ , U3969 );
nand NAND4_395 ( U3405 , U4663 , U4662 , U3754 , U3756 );
nand NAND2_396 ( U3406 , DATAI_25_ , U3969 );
nand NAND4_397 ( U3407 , U4682 , U4681 , U3758 , U3760 );
nand NAND2_398 ( U3408 , DATAI_26_ , U3969 );
nand NAND4_399 ( U3409 , U4701 , U4700 , U3762 , U3764 );
nand NAND2_400 ( U3410 , DATAI_27_ , U3969 );
nand NAND4_401 ( U3411 , U4720 , U4719 , U3766 , U3768 );
nand NAND2_402 ( U3412 , DATAI_28_ , U3969 );
nand NAND4_403 ( U3413 , U4739 , U4738 , U3770 , U3772 );
nand NAND2_404 ( U3414 , DATAI_29_ , U3969 );
nand NAND2_405 ( U3415 , DATAI_30_ , U3969 );
nand NAND2_406 ( U3416 , DATAI_31_ , U3969 );
nand NAND2_407 ( U3417 , U3023 , U4784 );
nand NAND3_408 ( U3418 , U5820 , U4010 , U5808 );
nand NAND3_409 ( U3419 , U3461 , U5820 , U3457 );
nand NAND2_410 ( U3420 , U3024 , U5817 );
nand NAND2_411 ( U3421 , U3356 , U4063 );
nand NAND2_412 ( U3422 , U4054 , STATE_REG );
nand NAND2_413 ( U3423 , U3015 , U3016 );
not NOT1_414 ( U3424 , R395_U6 );
nand NAND2_415 ( U3425 , U3901 , U3900 );
nand NAND2_416 ( U3426 , U3023 , U4021 );
nand NAND2_417 ( U3427 , U3905 , U3017 );
nand NAND2_418 ( U3428 , U3015 , U3023 );
nand NAND2_419 ( U3429 , U3907 , U5158 );
nand NAND2_420 ( U3430 , U5808 , U3461 );
nand NAND2_421 ( U3431 , U5747 , U5746 );
nand NAND2_422 ( U3432 , U5753 , U5752 );
nand NAND2_423 ( U3433 , U5756 , U5755 );
nand NAND2_424 ( U3434 , U5750 , U5749 );
nand NAND2_425 ( U3435 , U5759 , U5758 );
nand NAND2_426 ( U3436 , U5761 , U5760 );
nand NAND2_427 ( U3437 , U5763 , U5762 );
nand NAND2_428 ( U3438 , U5765 , U5764 );
nand NAND2_429 ( U3439 , U5767 , U5766 );
nand NAND2_430 ( U3440 , U5769 , U5768 );
nand NAND2_431 ( U3441 , U5771 , U5770 );
nand NAND2_432 ( U3442 , U5773 , U5772 );
nand NAND2_433 ( U3443 , U5775 , U5774 );
nand NAND2_434 ( U3444 , U5777 , U5776 );
nand NAND2_435 ( U3445 , U5779 , U5778 );
nand NAND2_436 ( U3446 , U5781 , U5780 );
nand NAND2_437 ( U3447 , U5783 , U5782 );
nand NAND2_438 ( U3448 , U5785 , U5784 );
nand NAND2_439 ( U3449 , U5787 , U5786 );
nand NAND2_440 ( U3450 , U5789 , U5788 );
nand NAND2_441 ( U3451 , U5791 , U5790 );
nand NAND2_442 ( U3452 , U5793 , U5792 );
nand NAND2_443 ( U3453 , U5795 , U5794 );
nand NAND2_444 ( U3454 , U5798 , U5797 );
nand NAND2_445 ( U3455 , U5801 , U5800 );
nand NAND2_446 ( U3456 , U5804 , U5803 );
nand NAND2_447 ( U3457 , U5807 , U5806 );
nand NAND2_448 ( U3458 , U5812 , U5811 );
nand NAND2_449 ( U3459 , U5814 , U5813 );
nand NAND2_450 ( U3460 , U5819 , U5818 );
nand NAND2_451 ( U3461 , U5816 , U5815 );
nand NAND2_452 ( U3462 , U5822 , U5821 );
nand NAND2_453 ( U3463 , U5825 , U5824 );
nand NAND2_454 ( U3464 , U5828 , U5827 );
nand NAND2_455 ( U3465 , U5836 , U5835 );
nand NAND2_456 ( U3466 , U5833 , U5832 );
nand NAND2_457 ( U3467 , U5839 , U5838 );
nand NAND2_458 ( U3468 , U5841 , U5840 );
nand NAND2_459 ( U3469 , U5844 , U5843 );
nand NAND2_460 ( U3470 , U5846 , U5845 );
nand NAND2_461 ( U3471 , U5849 , U5848 );
nand NAND2_462 ( U3472 , U5851 , U5850 );
nand NAND2_463 ( U3473 , U5854 , U5853 );
nand NAND2_464 ( U3474 , U5856 , U5855 );
nand NAND2_465 ( U3475 , U5859 , U5858 );
nand NAND2_466 ( U3476 , U5861 , U5860 );
nand NAND2_467 ( U3477 , U5864 , U5863 );
nand NAND2_468 ( U3478 , U5866 , U5865 );
nand NAND2_469 ( U3479 , U5869 , U5868 );
nand NAND2_470 ( U3480 , U5871 , U5870 );
nand NAND2_471 ( U3481 , U5874 , U5873 );
nand NAND2_472 ( U3482 , U5876 , U5875 );
nand NAND2_473 ( U3483 , U5879 , U5878 );
nand NAND2_474 ( U3484 , U5881 , U5880 );
nand NAND2_475 ( U3485 , U5884 , U5883 );
nand NAND2_476 ( U3486 , U5886 , U5885 );
nand NAND2_477 ( U3487 , U5889 , U5888 );
nand NAND2_478 ( U3488 , U5891 , U5890 );
nand NAND2_479 ( U3489 , U5894 , U5893 );
nand NAND2_480 ( U3490 , U5896 , U5895 );
nand NAND2_481 ( U3491 , U5899 , U5898 );
nand NAND2_482 ( U3492 , U5901 , U5900 );
nand NAND2_483 ( U3493 , U5904 , U5903 );
nand NAND2_484 ( U3494 , U5906 , U5905 );
nand NAND2_485 ( U3495 , U5909 , U5908 );
nand NAND2_486 ( U3496 , U5911 , U5910 );
nand NAND2_487 ( U3497 , U5914 , U5913 );
nand NAND2_488 ( U3498 , U5916 , U5915 );
nand NAND2_489 ( U3499 , U5919 , U5918 );
nand NAND2_490 ( U3500 , U5921 , U5920 );
nand NAND2_491 ( U3501 , U5924 , U5923 );
nand NAND2_492 ( U3502 , U5926 , U5925 );
nand NAND2_493 ( U3503 , U5929 , U5928 );
nand NAND2_494 ( U3504 , U5931 , U5930 );
nand NAND2_495 ( U3505 , U5934 , U5933 );
nand NAND2_496 ( U3506 , U5936 , U5935 );
nand NAND2_497 ( U3507 , U5938 , U5937 );
nand NAND2_498 ( U3508 , U5940 , U5939 );
nand NAND2_499 ( U3509 , U5942 , U5941 );
nand NAND2_500 ( U3510 , U5944 , U5943 );
nand NAND2_501 ( U3511 , U5946 , U5945 );
nand NAND2_502 ( U3512 , U5948 , U5947 );
nand NAND2_503 ( U3513 , U5950 , U5949 );
nand NAND2_504 ( U3514 , U5952 , U5951 );
nand NAND2_505 ( U3515 , U5954 , U5953 );
nand NAND2_506 ( U3516 , U5956 , U5955 );
nand NAND2_507 ( U3517 , U5958 , U5957 );
nand NAND2_508 ( U3518 , U5960 , U5959 );
nand NAND2_509 ( U3519 , U5962 , U5961 );
nand NAND2_510 ( U3520 , U5964 , U5963 );
nand NAND2_511 ( U3521 , U5966 , U5965 );
nand NAND2_512 ( U3522 , U5968 , U5967 );
nand NAND2_513 ( U3523 , U5970 , U5969 );
nand NAND2_514 ( U3524 , U5972 , U5971 );
nand NAND2_515 ( U3525 , U5974 , U5973 );
nand NAND2_516 ( U3526 , U5976 , U5975 );
nand NAND2_517 ( U3527 , U5978 , U5977 );
nand NAND2_518 ( U3528 , U5980 , U5979 );
nand NAND2_519 ( U3529 , U5982 , U5981 );
nand NAND2_520 ( U3530 , U5984 , U5983 );
nand NAND2_521 ( U3531 , U5986 , U5985 );
nand NAND2_522 ( U3532 , U5988 , U5987 );
nand NAND2_523 ( U3533 , U5990 , U5989 );
nand NAND2_524 ( U3534 , U5992 , U5991 );
nand NAND2_525 ( U3535 , U5994 , U5993 );
nand NAND2_526 ( U3536 , U5996 , U5995 );
nand NAND2_527 ( U3537 , U5998 , U5997 );
nand NAND2_528 ( U3538 , U6000 , U5999 );
nand NAND2_529 ( U3539 , U6002 , U6001 );
nand NAND2_530 ( U3540 , U6004 , U6003 );
nand NAND2_531 ( U3541 , U6006 , U6005 );
nand NAND2_532 ( U3542 , U6008 , U6007 );
nand NAND2_533 ( U3543 , U6010 , U6009 );
nand NAND2_534 ( U3544 , U6012 , U6011 );
nand NAND2_535 ( U3545 , U6014 , U6013 );
nand NAND2_536 ( U3546 , U6016 , U6015 );
nand NAND2_537 ( U3547 , U6018 , U6017 );
nand NAND2_538 ( U3548 , U6020 , U6019 );
nand NAND2_539 ( U3549 , U6022 , U6021 );
nand NAND2_540 ( U3550 , U6088 , U6087 );
nand NAND2_541 ( U3551 , U6090 , U6089 );
nand NAND2_542 ( U3552 , U6092 , U6091 );
nand NAND2_543 ( U3553 , U6094 , U6093 );
nand NAND2_544 ( U3554 , U6096 , U6095 );
nand NAND2_545 ( U3555 , U6098 , U6097 );
nand NAND2_546 ( U3556 , U6100 , U6099 );
nand NAND2_547 ( U3557 , U6102 , U6101 );
nand NAND2_548 ( U3558 , U6104 , U6103 );
nand NAND2_549 ( U3559 , U6106 , U6105 );
nand NAND2_550 ( U3560 , U6108 , U6107 );
nand NAND2_551 ( U3561 , U6110 , U6109 );
nand NAND2_552 ( U3562 , U6112 , U6111 );
nand NAND2_553 ( U3563 , U6114 , U6113 );
nand NAND2_554 ( U3564 , U6116 , U6115 );
nand NAND2_555 ( U3565 , U6118 , U6117 );
nand NAND2_556 ( U3566 , U6120 , U6119 );
nand NAND2_557 ( U3567 , U6122 , U6121 );
nand NAND2_558 ( U3568 , U6124 , U6123 );
nand NAND2_559 ( U3569 , U6126 , U6125 );
nand NAND2_560 ( U3570 , U6128 , U6127 );
nand NAND2_561 ( U3571 , U6130 , U6129 );
nand NAND2_562 ( U3572 , U6132 , U6131 );
nand NAND2_563 ( U3573 , U6134 , U6133 );
nand NAND2_564 ( U3574 , U6136 , U6135 );
nand NAND2_565 ( U3575 , U6138 , U6137 );
nand NAND2_566 ( U3576 , U6140 , U6139 );
nand NAND2_567 ( U3577 , U6142 , U6141 );
nand NAND2_568 ( U3578 , U6144 , U6143 );
nand NAND2_569 ( U3579 , U6146 , U6145 );
nand NAND2_570 ( U3580 , U6148 , U6147 );
nand NAND2_571 ( U3581 , U6150 , U6149 );
nand NAND2_572 ( U3582 , U6261 , U6260 );
nand NAND2_573 ( U3583 , U6263 , U6262 );
nand NAND2_574 ( U3584 , U6265 , U6264 );
nand NAND2_575 ( U3585 , U6267 , U6266 );
nand NAND2_576 ( U3586 , U6269 , U6268 );
nand NAND2_577 ( U3587 , U6271 , U6270 );
nand NAND2_578 ( U3588 , U6273 , U6272 );
nand NAND2_579 ( U3589 , U6275 , U6274 );
nand NAND2_580 ( U3590 , U6277 , U6276 );
nand NAND2_581 ( U3591 , U6279 , U6278 );
nand NAND2_582 ( U3592 , U6281 , U6280 );
nand NAND2_583 ( U3593 , U6283 , U6282 );
nand NAND2_584 ( U3594 , U6285 , U6284 );
nand NAND2_585 ( U3595 , U6287 , U6286 );
nand NAND2_586 ( U3596 , U6289 , U6288 );
nand NAND2_587 ( U3597 , U6291 , U6290 );
nand NAND2_588 ( U3598 , U6293 , U6292 );
nand NAND2_589 ( U3599 , U6295 , U6294 );
nand NAND2_590 ( U3600 , U6297 , U6296 );
nand NAND2_591 ( U3601 , U6299 , U6298 );
nand NAND2_592 ( U3602 , U6301 , U6300 );
nand NAND2_593 ( U3603 , U6303 , U6302 );
nand NAND2_594 ( U3604 , U6305 , U6304 );
nand NAND2_595 ( U3605 , U6307 , U6306 );
nand NAND2_596 ( U3606 , U6309 , U6308 );
nand NAND2_597 ( U3607 , U6311 , U6310 );
nand NAND2_598 ( U3608 , U6313 , U6312 );
nand NAND2_599 ( U3609 , U6315 , U6314 );
nand NAND2_600 ( U3610 , U6317 , U6316 );
nand NAND2_601 ( U3611 , U6319 , U6318 );
nand NAND2_602 ( U3612 , U6321 , U6320 );
nand NAND2_603 ( U3613 , U6323 , U6322 );
and AND2_604 ( U3614 , U4067 , U4065 );
and AND2_605 ( U3615 , U4070 , U4068 );
and AND2_606 ( U3616 , U4073 , U4071 );
and AND2_607 ( U3617 , U4076 , U4074 );
and AND2_608 ( U3618 , U4079 , U4077 );
and AND2_609 ( U3619 , U4082 , U4080 );
and AND2_610 ( U3620 , U4085 , U4083 );
and AND2_611 ( U3621 , U4088 , U4086 );
and AND2_612 ( U3622 , U4091 , U4089 );
and AND2_613 ( U3623 , U4094 , U4092 );
and AND2_614 ( U3624 , U4097 , U4095 );
and AND2_615 ( U3625 , U4100 , U4098 );
and AND2_616 ( U3626 , U4103 , U4101 );
and AND2_617 ( U3627 , U4106 , U4104 );
and AND2_618 ( U3628 , U4109 , U4107 );
and AND2_619 ( U3629 , U4112 , U4110 );
and AND2_620 ( U3630 , U4115 , U4113 );
and AND2_621 ( U3631 , U4118 , U4116 );
and AND2_622 ( U3632 , U4121 , U4119 );
and AND2_623 ( U3633 , U4124 , U4122 );
and AND2_624 ( U3634 , U4127 , U4125 );
and AND2_625 ( U3635 , U4130 , U4128 );
and AND2_626 ( U3636 , U4133 , U4131 );
and AND2_627 ( U3637 , U4136 , U4134 );
and AND2_628 ( U3638 , U4139 , U4137 );
and AND2_629 ( U3639 , U4142 , U4140 );
and AND2_630 ( U3640 , U4145 , U4143 );
and AND2_631 ( U3641 , U4148 , U4146 );
and AND2_632 ( U3642 , U4151 , U4149 );
and AND2_633 ( U3643 , U4154 , U4152 );
and AND2_634 ( U3644 , U4157 , U4155 );
and AND2_635 ( U3645 , U4160 , U4158 );
and AND2_636 ( U3646 , U4203 , U4202 );
and AND2_637 ( U3647 , U4205 , U4204 );
and AND2_638 ( U3648 , U4212 , U4210 );
and AND3_639 ( U3649 , U4213 , U4211 , U3648 );
and AND4_640 ( U3650 , U4167 , U4166 , U4165 , U4164 );
and AND4_641 ( U3651 , U4171 , U4170 , U4169 , U4168 );
and AND4_642 ( U3652 , U4175 , U4174 , U4173 , U4172 );
and AND3_643 ( U3653 , U4177 , U4176 , U4178 );
and AND4_644 ( U3654 , U3653 , U3652 , U3651 , U3650 );
and AND4_645 ( U3655 , U4182 , U4181 , U4180 , U4179 );
and AND4_646 ( U3656 , U4186 , U4185 , U4184 , U4183 );
and AND4_647 ( U3657 , U4190 , U4189 , U4188 , U4187 );
and AND3_648 ( U3658 , U4192 , U4191 , U4193 );
and AND4_649 ( U3659 , U3658 , U3657 , U3656 , U3655 );
and AND2_650 ( U3660 , U5834 , U4195 );
and AND2_651 ( U3661 , U5837 , U3023 );
and AND2_652 ( U3662 , U4228 , U4227 );
and AND2_653 ( U3663 , U4230 , U4229 );
and AND3_654 ( U3664 , U4232 , U4231 , U3663 );
and AND4_655 ( U3665 , U4235 , U4236 , U4237 , U4234 );
and AND2_656 ( U3666 , U4247 , U4246 );
and AND2_657 ( U3667 , U4249 , U4248 );
and AND3_658 ( U3668 , U4251 , U4250 , U3667 );
and AND4_659 ( U3669 , U4254 , U4255 , U4256 , U4253 );
and AND2_660 ( U3670 , U4266 , U4265 );
and AND2_661 ( U3671 , U4268 , U4267 );
and AND3_662 ( U3672 , U4270 , U4269 , U3671 );
and AND4_663 ( U3673 , U4273 , U4274 , U4275 , U4272 );
and AND2_664 ( U3674 , U4285 , U4284 );
and AND2_665 ( U3675 , U4287 , U4286 );
and AND3_666 ( U3676 , U4289 , U4288 , U3675 );
and AND4_667 ( U3677 , U4292 , U4293 , U4294 , U4291 );
and AND2_668 ( U3678 , U4304 , U4303 );
and AND2_669 ( U3679 , U4306 , U4305 );
and AND3_670 ( U3680 , U4308 , U4307 , U3679 );
and AND4_671 ( U3681 , U4311 , U4312 , U4313 , U4310 );
and AND2_672 ( U3682 , U4323 , U4322 );
and AND2_673 ( U3683 , U4325 , U4324 );
and AND3_674 ( U3684 , U4327 , U4326 , U3683 );
and AND4_675 ( U3685 , U4330 , U4331 , U4332 , U4329 );
and AND2_676 ( U3686 , U4342 , U4341 );
and AND2_677 ( U3687 , U4344 , U4343 );
and AND3_678 ( U3688 , U4346 , U4345 , U3687 );
and AND4_679 ( U3689 , U4349 , U4350 , U4351 , U4348 );
and AND2_680 ( U3690 , U4361 , U4360 );
and AND2_681 ( U3691 , U4363 , U4362 );
and AND3_682 ( U3692 , U4365 , U4364 , U3691 );
and AND4_683 ( U3693 , U4368 , U4369 , U4370 , U4367 );
and AND2_684 ( U3694 , U4380 , U4379 );
and AND2_685 ( U3695 , U4382 , U4381 );
and AND3_686 ( U3696 , U4384 , U4383 , U3695 );
and AND4_687 ( U3697 , U4387 , U4388 , U4389 , U4386 );
and AND2_688 ( U3698 , U4399 , U4398 );
and AND2_689 ( U3699 , U4401 , U4400 );
and AND3_690 ( U3700 , U4403 , U4402 , U3699 );
and AND4_691 ( U3701 , U4406 , U4407 , U4408 , U4405 );
and AND2_692 ( U3702 , U4418 , U4417 );
and AND2_693 ( U3703 , U4420 , U4419 );
and AND3_694 ( U3704 , U4422 , U4421 , U3703 );
and AND4_695 ( U3705 , U4425 , U4426 , U4427 , U4424 );
and AND2_696 ( U3706 , U4437 , U4436 );
and AND2_697 ( U3707 , U4439 , U4438 );
and AND3_698 ( U3708 , U4441 , U4440 , U3707 );
and AND4_699 ( U3709 , U4444 , U4445 , U4446 , U4443 );
and AND2_700 ( U3710 , U4456 , U4455 );
and AND2_701 ( U3711 , U4458 , U4457 );
and AND3_702 ( U3712 , U4460 , U4459 , U3711 );
and AND4_703 ( U3713 , U4463 , U4464 , U4465 , U4462 );
and AND2_704 ( U3714 , U4475 , U4474 );
and AND2_705 ( U3715 , U4477 , U4476 );
and AND3_706 ( U3716 , U4479 , U4478 , U3715 );
and AND4_707 ( U3717 , U4482 , U4483 , U4484 , U4481 );
and AND2_708 ( U3718 , U4494 , U4493 );
and AND2_709 ( U3719 , U4496 , U4495 );
and AND3_710 ( U3720 , U4498 , U4497 , U3719 );
and AND4_711 ( U3721 , U4501 , U4502 , U4503 , U4500 );
and AND2_712 ( U3722 , U4513 , U4512 );
and AND2_713 ( U3723 , U4515 , U4514 );
and AND3_714 ( U3724 , U4517 , U4516 , U3723 );
and AND4_715 ( U3725 , U4520 , U4521 , U4522 , U4519 );
and AND2_716 ( U3726 , U4532 , U4531 );
and AND2_717 ( U3727 , U4534 , U4533 );
and AND3_718 ( U3728 , U4536 , U4535 , U3727 );
and AND4_719 ( U3729 , U4539 , U4540 , U4541 , U4538 );
and AND2_720 ( U3730 , U4551 , U4550 );
and AND2_721 ( U3731 , U4553 , U4552 );
and AND3_722 ( U3732 , U4555 , U4554 , U3731 );
and AND4_723 ( U3733 , U4558 , U4559 , U4560 , U4557 );
and AND2_724 ( U3734 , U4570 , U4569 );
and AND2_725 ( U3735 , U4572 , U4571 );
and AND3_726 ( U3736 , U4574 , U4573 , U3735 );
and AND4_727 ( U3737 , U4577 , U4578 , U4579 , U4576 );
and AND2_728 ( U3738 , U4589 , U4588 );
and AND2_729 ( U3739 , U4591 , U4590 );
and AND3_730 ( U3740 , U4593 , U4592 , U3739 );
and AND4_731 ( U3741 , U4596 , U4597 , U4598 , U4595 );
and AND2_732 ( U3742 , U4608 , U4607 );
and AND2_733 ( U3743 , U4610 , U4609 );
and AND3_734 ( U3744 , U4612 , U4611 , U3743 );
and AND4_735 ( U3745 , U4615 , U4616 , U4617 , U4614 );
and AND2_736 ( U3746 , U4627 , U4626 );
and AND2_737 ( U3747 , U4629 , U4628 );
and AND3_738 ( U3748 , U4631 , U4630 , U3747 );
and AND4_739 ( U3749 , U4634 , U4635 , U4636 , U4633 );
and AND2_740 ( U3750 , U4646 , U4645 );
and AND2_741 ( U3751 , U4648 , U4647 );
and AND3_742 ( U3752 , U4650 , U4649 , U3751 );
and AND4_743 ( U3753 , U4653 , U4654 , U4655 , U4652 );
and AND2_744 ( U3754 , U4665 , U4664 );
and AND2_745 ( U3755 , U4667 , U4666 );
and AND3_746 ( U3756 , U4669 , U4668 , U3755 );
and AND4_747 ( U3757 , U4672 , U4673 , U4674 , U4671 );
and AND2_748 ( U3758 , U4684 , U4683 );
and AND2_749 ( U3759 , U4686 , U4685 );
and AND3_750 ( U3760 , U4688 , U4687 , U3759 );
and AND4_751 ( U3761 , U4691 , U4692 , U4693 , U4690 );
and AND2_752 ( U3762 , U4703 , U4702 );
and AND2_753 ( U3763 , U4705 , U4704 );
and AND3_754 ( U3764 , U4707 , U4706 , U3763 );
and AND4_755 ( U3765 , U4710 , U4711 , U4712 , U4709 );
and AND2_756 ( U3766 , U4722 , U4721 );
and AND2_757 ( U3767 , U4724 , U4723 );
and AND3_758 ( U3768 , U4726 , U4725 , U3767 );
and AND4_759 ( U3769 , U4729 , U4730 , U4731 , U4728 );
and AND2_760 ( U3770 , U4741 , U4740 );
and AND2_761 ( U3771 , U4743 , U4742 );
and AND3_762 ( U3772 , U4745 , U4744 , U3771 );
and AND4_763 ( U3773 , U4748 , U4749 , U4750 , U4747 );
and AND2_764 ( U3774 , U4757 , U4042 );
and AND4_765 ( U3775 , U4764 , U4763 , U4761 , U4760 );
and AND3_766 ( U3776 , U4769 , U4770 , U4768 );
and AND2_767 ( U3777 , U4042 , U4757 );
and AND2_768 ( U3778 , U3023 , U3465 );
and AND3_769 ( U3779 , U5837 , U4025 , U3466 );
and AND3_770 ( U3780 , U4786 , U4785 , U4787 );
and AND3_771 ( U3781 , U4789 , U4788 , U3972 );
and AND3_772 ( U3782 , U4791 , U4790 , U4792 );
and AND3_773 ( U3783 , U4794 , U4793 , U3973 );
and AND3_774 ( U3784 , U4796 , U4795 , U4797 );
and AND3_775 ( U3785 , U4799 , U4798 , U3974 );
and AND3_776 ( U3786 , U4801 , U4800 , U4802 );
and AND3_777 ( U3787 , U4804 , U4803 , U3975 );
and AND3_778 ( U3788 , U4806 , U4805 , U4807 );
and AND3_779 ( U3789 , U4809 , U4808 , U3976 );
and AND3_780 ( U3790 , U4811 , U4810 , U4812 );
and AND2_781 ( U3791 , U4814 , U4813 );
and AND3_782 ( U3792 , U4816 , U4815 , U4817 );
and AND2_783 ( U3793 , U4819 , U4818 );
and AND3_784 ( U3794 , U4821 , U4820 , U4822 );
and AND2_785 ( U3795 , U4824 , U4823 );
and AND3_786 ( U3796 , U4826 , U4825 , U4827 );
and AND2_787 ( U3797 , U4829 , U4828 );
and AND3_788 ( U3798 , U4831 , U4830 , U4832 );
and AND2_789 ( U3799 , U4834 , U4833 );
and AND3_790 ( U3800 , U4836 , U4835 , U4837 );
and AND2_791 ( U3801 , U4839 , U4838 );
and AND3_792 ( U3802 , U4841 , U4840 , U4842 );
and AND2_793 ( U3803 , U4844 , U4843 );
and AND3_794 ( U3804 , U4846 , U4845 , U4847 );
and AND2_795 ( U3805 , U4849 , U4848 );
and AND2_796 ( U3806 , U4851 , U4850 );
and AND2_797 ( U3807 , U4854 , U4853 );
and AND3_798 ( U3808 , U4856 , U4855 , U4857 );
and AND2_799 ( U3809 , U4859 , U4858 );
and AND2_800 ( U3810 , U4861 , U4860 );
and AND2_801 ( U3811 , U4864 , U4863 );
and AND2_802 ( U3812 , U4866 , U4865 );
and AND2_803 ( U3813 , U4869 , U4868 );
and AND2_804 ( U3814 , U4871 , U4870 );
and AND2_805 ( U3815 , U4874 , U4873 );
and AND2_806 ( U3816 , U4876 , U4875 );
and AND2_807 ( U3817 , U4879 , U4878 );
and AND2_808 ( U3818 , U4881 , U4880 );
and AND2_809 ( U3819 , U4884 , U4883 );
and AND2_810 ( U3820 , U4886 , U4885 );
and AND2_811 ( U3821 , U4889 , U4888 );
and AND2_812 ( U3822 , U4891 , U4890 );
and AND2_813 ( U3823 , U4894 , U4893 );
and AND2_814 ( U3824 , U4896 , U4895 );
and AND2_815 ( U3825 , U4899 , U4898 );
and AND2_816 ( U3826 , U4901 , U4900 );
and AND2_817 ( U3827 , U4904 , U4903 );
and AND2_818 ( U3828 , U4906 , U4905 );
and AND2_819 ( U3829 , U4909 , U4908 );
and AND2_820 ( U3830 , U4911 , U4910 );
and AND2_821 ( U3831 , U4914 , U4913 );
and AND2_822 ( U3832 , U4916 , U4915 );
and AND2_823 ( U3833 , U4919 , U4918 );
and AND2_824 ( U3834 , U4921 , U4920 );
and AND2_825 ( U3835 , U4924 , U4923 );
and AND2_826 ( U3836 , U4926 , U4925 );
and AND2_827 ( U3837 , U4929 , U4928 );
and AND3_828 ( U3838 , U5738 , U5737 , U5739 );
and AND3_829 ( U3839 , U3419 , U3370 , U3367 );
and AND3_830 ( U3840 , U3368 , U3362 , U3366 );
and AND2_831 ( U3841 , U3363 , U3364 );
and AND2_832 ( U3842 , U3841 , U3420 );
and AND2_833 ( U3843 , U3353 , U3418 );
and AND2_834 ( U3844 , U3040 , U3461 );
and AND2_835 ( U3845 , U3431 , STATE_REG );
and AND4_836 ( U3846 , U4940 , U4939 , U4943 , U4941 );
and AND2_837 ( U3847 , U4947 , U4944 );
and AND3_838 ( U3848 , U4945 , U3847 , U4946 );
and AND2_839 ( U3849 , U3040 , U3444 );
and AND4_840 ( U3850 , U4949 , U4948 , U4951 , U4950 );
and AND2_841 ( U3851 , U4955 , U4952 );
and AND3_842 ( U3852 , U4953 , U3851 , U4954 );
and AND2_843 ( U3853 , U4961 , U4962 );
and AND2_844 ( U3854 , U4965 , U4963 );
and AND2_845 ( U3855 , U4971 , U4972 );
and AND2_846 ( U3856 , U4975 , U4973 );
and AND2_847 ( U3857 , U4981 , U4982 );
and AND2_848 ( U3858 , U4985 , U4983 );
and AND2_849 ( U3859 , U4991 , U4992 );
and AND2_850 ( U3860 , U4995 , U4993 );
and AND2_851 ( U3861 , U5001 , U5002 );
and AND2_852 ( U3862 , U5005 , U5003 );
and AND2_853 ( U3863 , U5011 , U5012 );
and AND2_854 ( U3864 , U5015 , U5013 );
and AND2_855 ( U3865 , U5021 , U5022 );
and AND2_856 ( U3866 , U5025 , U5023 );
and AND2_857 ( U3867 , U5031 , U5032 );
and AND2_858 ( U3868 , U5035 , U5033 );
and AND2_859 ( U3869 , U5041 , U5042 );
and AND2_860 ( U3870 , U5045 , U5043 );
and AND2_861 ( U3871 , U5051 , U5052 );
and AND2_862 ( U3872 , U5055 , U5053 );
and AND3_863 ( U3873 , U5061 , U5062 , U5060 );
and AND3_864 ( U3874 , U5064 , U5063 , U5065 );
and AND3_865 ( U3875 , U5071 , U5072 , U5070 );
and AND3_866 ( U3876 , U5074 , U5073 , U5075 );
and AND3_867 ( U3877 , U5081 , U5082 , U5080 );
and AND3_868 ( U3878 , U5084 , U5083 , U5085 );
and AND2_869 ( U3879 , U5090 , U4053 );
and AND3_870 ( U3880 , U5092 , U5091 , U3879 );
and AND3_871 ( U3881 , U5094 , U5093 , U5095 );
and AND3_872 ( U3882 , U5101 , U5102 , U5100 );
and AND3_873 ( U3883 , U5104 , U5103 , U5105 );
and AND2_874 ( U3884 , U5110 , U4053 );
and AND3_875 ( U3885 , U5112 , U5111 , U3884 );
and AND3_876 ( U3886 , U5114 , U5113 , U5115 );
and AND3_877 ( U3887 , U5121 , U5122 , U5120 );
and AND3_878 ( U3888 , U5124 , U5123 , U5125 );
and AND3_879 ( U3889 , U5131 , U5132 , U5130 );
and AND3_880 ( U3890 , U5134 , U5133 , U5135 );
and AND4_881 ( U3891 , U6210 , U6207 , U6204 , U6201 );
and AND4_882 ( U3892 , U6222 , U6219 , U6216 , U6213 );
and AND4_883 ( U3893 , U6234 , U6231 , U6228 , U6225 );
and AND4_884 ( U3894 , U6246 , U6243 , U6240 , U6237 );
and AND4_885 ( U3895 , U6174 , U6171 , U6168 , U6165 );
and AND3_886 ( U3896 , U6159 , U6156 , U6162 );
and AND4_887 ( U3897 , U6192 , U6189 , U6186 , U6183 );
and AND2_888 ( U3898 , U6180 , U6177 );
and AND2_889 ( U3899 , U6198 , U6195 );
and AND5_890 ( U3900 , U3895 , U3896 , U6153 , U3897 , U3898 );
and AND5_891 ( U3901 , U3894 , U3893 , U3892 , U3891 , U3899 );
and AND4_892 ( U3902 , U6255 , U6254 , U5141 , U5140 );
and AND2_893 ( U3903 , U3356 , STATE_REG );
and AND2_894 ( U3904 , U5148 , U5146 );
and AND2_895 ( U3905 , U3465 , U3466 );
and AND3_896 ( U3906 , U3371 , U3420 , U4008 );
and AND3_897 ( U3907 , U3356 , U4025 , U5748 );
and AND2_898 ( U3908 , U3023 , U5157 );
and AND2_899 ( U3909 , U3910 , U5200 );
and AND2_900 ( U3910 , U5204 , U5203 );
and AND2_901 ( U3911 , U4049 , U3075 );
and AND2_902 ( U3912 , U5245 , U5244 );
and AND2_903 ( U3913 , U5248 , U5247 );
and AND2_904 ( U3914 , U5266 , U5265 );
and AND2_905 ( U3915 , U5293 , U5292 );
and AND2_906 ( U3916 , U3917 , U5334 );
and AND2_907 ( U3917 , U5338 , U5337 );
and AND2_908 ( U3918 , U3919 , U5370 );
and AND2_909 ( U3919 , U5374 , U5373 );
and AND3_910 ( U3920 , U3431 , U5423 , U5425 );
and AND3_911 ( U3921 , U3431 , U5426 , U5428 );
and AND3_912 ( U3922 , U3431 , U5429 , U5431 );
and AND3_913 ( U3923 , U3431 , U5432 , U5434 );
and AND3_914 ( U3924 , U3431 , U5435 , U5437 );
and AND3_915 ( U3925 , U3431 , U5438 , U5440 );
and AND2_916 ( U3926 , U5442 , U5443 );
and AND2_917 ( U3927 , U5445 , U5446 );
and AND3_918 ( U3928 , U3431 , U5447 , U5449 );
and AND2_919 ( U3929 , U5452 , U3930 );
and AND2_920 ( U3930 , U3431 , U5451 );
and AND2_921 ( U3931 , U5455 , U3932 );
and AND2_922 ( U3932 , U3431 , U5454 );
and AND2_923 ( U3933 , U5458 , U3934 );
and AND2_924 ( U3934 , U3431 , U5457 );
and AND2_925 ( U3935 , U5461 , U3936 );
and AND2_926 ( U3936 , U3431 , U5460 );
and AND2_927 ( U3937 , U5464 , U3938 );
and AND2_928 ( U3938 , U3431 , U5463 );
and AND2_929 ( U3939 , U5467 , U3940 );
and AND2_930 ( U3940 , U3431 , U5466 );
and AND2_931 ( U3941 , U5470 , U3942 );
and AND2_932 ( U3942 , U3431 , U5469 );
and AND2_933 ( U3943 , U5473 , U3944 );
and AND2_934 ( U3944 , U3431 , U5472 );
and AND2_935 ( U3945 , U5476 , U3946 );
and AND2_936 ( U3946 , U3431 , U5475 );
and AND2_937 ( U3947 , U5479 , U3948 );
and AND2_938 ( U3948 , U3431 , U5478 );
and AND3_939 ( U3949 , U3431 , U5480 , U5482 );
and AND3_940 ( U3950 , U3431 , U5483 , U5485 );
and AND3_941 ( U3951 , U3431 , U5486 , U5488 );
and AND3_942 ( U3952 , U3431 , U5489 , U5491 );
and AND3_943 ( U3953 , U3431 , U5492 , U5494 );
and AND3_944 ( U3954 , U3431 , U5495 , U5497 );
and AND3_945 ( U3955 , U3431 , U5498 , U5500 );
and AND3_946 ( U3956 , U3431 , U5501 , U5503 );
and AND3_947 ( U3957 , U3431 , U5504 , U5506 );
and AND3_948 ( U3958 , U3431 , U5507 , U5509 );
and AND3_949 ( U3959 , U3431 , U5510 , U5512 );
and AND3_950 ( U3960 , U3431 , U5513 , U5515 );
and AND3_951 ( U3961 , U3431 , U5516 , U5518 );
and AND2_952 ( U3962 , U5808 , U5805 );
and AND2_953 ( U3963 , U3365 , U3430 );
and AND2_954 ( U3964 , U5616 , U4026 );
and AND2_955 ( U3965 , U5676 , U5677 );
and AND2_956 ( U3966 , U5736 , U5734 );
not NOT1_957 ( U3967 , IR_REG_31_ );
nand NAND2_958 ( U3968 , U3023 , U3360 );
nand NAND2_959 ( U3969 , U5802 , U5799 );
nand NAND2_960 ( U3970 , U3661 , U3048 );
nand NAND2_961 ( U3971 , U3778 , U3048 );
and AND2_962 ( U3972 , U6024 , U6023 );
and AND2_963 ( U3973 , U6026 , U6025 );
and AND2_964 ( U3974 , U6028 , U6027 );
and AND2_965 ( U3975 , U6030 , U6029 );
and AND2_966 ( U3976 , U6032 , U6031 );
and AND2_967 ( U3977 , U6034 , U6033 );
and AND2_968 ( U3978 , U6036 , U6035 );
and AND2_969 ( U3979 , U6038 , U6037 );
and AND2_970 ( U3980 , U6040 , U6039 );
and AND2_971 ( U3981 , U6042 , U6041 );
and AND2_972 ( U3982 , U6044 , U6043 );
and AND2_973 ( U3983 , U6046 , U6045 );
and AND2_974 ( U3984 , U6048 , U6047 );
and AND2_975 ( U3985 , U6050 , U6049 );
and AND2_976 ( U3986 , U6052 , U6051 );
and AND2_977 ( U3987 , U6054 , U6053 );
and AND2_978 ( U3988 , U6056 , U6055 );
and AND2_979 ( U3989 , U6058 , U6057 );
and AND2_980 ( U3990 , U6060 , U6059 );
and AND2_981 ( U3991 , U6062 , U6061 );
and AND2_982 ( U3992 , U6064 , U6063 );
and AND2_983 ( U3993 , U6066 , U6065 );
and AND2_984 ( U3994 , U6068 , U6067 );
and AND2_985 ( U3995 , U6070 , U6069 );
and AND2_986 ( U3996 , U6072 , U6071 );
and AND2_987 ( U3997 , U6074 , U6073 );
and AND2_988 ( U3998 , U6076 , U6075 );
and AND2_989 ( U3999 , U6078 , U6077 );
and AND2_990 ( U4000 , U6080 , U6079 );
and AND2_991 ( U4001 , U6082 , U6081 );
nand NAND2_992 ( U4002 , U3777 , U3053 );
and AND2_993 ( U4003 , U6084 , U6083 );
and AND2_994 ( U4004 , U6086 , U6085 );
not NOT1_995 ( U4005 , R1375_U26 );
and AND2_996 ( U4006 , U6251 , U6250 );
not NOT1_997 ( U4007 , R1347_U13 );
nand NAND2_998 ( U4008 , U4013 , U5805 );
not NOT1_999 ( U4009 , R1352_U6 );
not NOT1_1000 ( U4010 , U3372 );
not NOT1_1001 ( U4011 , U3370 );
not NOT1_1002 ( U4012 , U3419 );
not NOT1_1003 ( U4013 , U3367 );
not NOT1_1004 ( U4014 , U3366 );
not NOT1_1005 ( U4015 , U3368 );
not NOT1_1006 ( U4016 , U3362 );
not NOT1_1007 ( U4017 , U3364 );
not NOT1_1008 ( U4018 , U3363 );
not NOT1_1009 ( U4019 , U3420 );
not NOT1_1010 ( U4020 , U3418 );
not NOT1_1011 ( U4021 , U3353 );
not NOT1_1012 ( U4022 , U3371 );
not NOT1_1013 ( U4023 , U4008 );
not NOT1_1014 ( U4024 , U3369 );
nand NAND2_1015 ( U4025 , U4042 , U4782 );
nand NAND2_1016 ( U4026 , U3962 , U3355 );
not NOT1_1017 ( U4027 , U3969 );
not NOT1_1018 ( U4028 , U3427 );
not NOT1_1019 ( U4029 , U3412 );
not NOT1_1020 ( U4030 , U3410 );
not NOT1_1021 ( U4031 , U3408 );
not NOT1_1022 ( U4032 , U3406 );
not NOT1_1023 ( U4033 , U3404 );
not NOT1_1024 ( U4034 , U3402 );
not NOT1_1025 ( U4035 , U3400 );
not NOT1_1026 ( U4036 , U3398 );
not NOT1_1027 ( U4037 , U3396 );
not NOT1_1028 ( U4038 , U3416 );
not NOT1_1029 ( U4039 , U3415 );
not NOT1_1030 ( U4040 , U3414 );
not NOT1_1031 ( U4041 , U3423 );
not NOT1_1032 ( U4042 , U3373 );
not NOT1_1033 ( U4043 , U3422 );
not NOT1_1034 ( U4044 , U3417 );
not NOT1_1035 ( U4045 , U3971 );
not NOT1_1036 ( U4046 , U3970 );
not NOT1_1037 ( U4047 , U3968 );
not NOT1_1038 ( U4048 , U4002 );
not NOT1_1039 ( U4049 , U3428 );
nand NAND2_1040 ( U4050 , U3429 , STATE_REG );
nand NAND2_1041 ( U4051 , U4020 , U3023 );
not NOT1_1042 ( U4052 , U3426 );
nand NAND2_1043 ( U4053 , U4043 , U3209 );
not NOT1_1044 ( U4054 , U3356 );
not NOT1_1045 ( U4055 , U3374 );
not NOT1_1046 ( U4056 , U3365 );
not NOT1_1047 ( U4057 , U3430 );
not NOT1_1048 ( U4058 , U3358 );
not NOT1_1049 ( U4059 , U3355 );
nand NAND2_1050 ( U4060 , U3047 , U3373 );
nand NAND2_1051 ( U4061 , U5748 , U4060 );
nand NAND2_1052 ( U4062 , U4061 , U3969 );
not NOT1_1053 ( U4063 , U3148 );
not NOT1_1054 ( U4064 , U3357 );
nand NAND2_1055 ( U4065 , DATAI_0_ , U3149 );
nand NAND2_1056 ( U4066 , U3029 , IR_REG_0_ );
nand NAND2_1057 ( U4067 , U4064 , IR_REG_0_ );
nand NAND2_1058 ( U4068 , DATAI_1_ , U3149 );
nand NAND2_1059 ( U4069 , U3029 , SUB_84_U48 );
nand NAND2_1060 ( U4070 , U4064 , IR_REG_1_ );
nand NAND2_1061 ( U4071 , DATAI_2_ , U3149 );
nand NAND2_1062 ( U4072 , U3029 , SUB_84_U20 );
nand NAND2_1063 ( U4073 , U4064 , IR_REG_2_ );
nand NAND2_1064 ( U4074 , DATAI_3_ , U3149 );
nand NAND2_1065 ( U4075 , U3029 , SUB_84_U21 );
nand NAND2_1066 ( U4076 , U4064 , IR_REG_3_ );
nand NAND2_1067 ( U4077 , DATAI_4_ , U3149 );
nand NAND2_1068 ( U4078 , U3029 , SUB_84_U70 );
nand NAND2_1069 ( U4079 , U4064 , IR_REG_4_ );
nand NAND2_1070 ( U4080 , DATAI_5_ , U3149 );
nand NAND2_1071 ( U4081 , U3029 , SUB_84_U22 );
nand NAND2_1072 ( U4082 , U4064 , IR_REG_5_ );
nand NAND2_1073 ( U4083 , DATAI_6_ , U3149 );
nand NAND2_1074 ( U4084 , U3029 , SUB_84_U23 );
nand NAND2_1075 ( U4085 , U4064 , IR_REG_6_ );
nand NAND2_1076 ( U4086 , DATAI_7_ , U3149 );
nand NAND2_1077 ( U4087 , U3029 , SUB_84_U24 );
nand NAND2_1078 ( U4088 , U4064 , IR_REG_7_ );
nand NAND2_1079 ( U4089 , DATAI_8_ , U3149 );
nand NAND2_1080 ( U4090 , U3029 , SUB_84_U68 );
nand NAND2_1081 ( U4091 , U4064 , IR_REG_8_ );
nand NAND2_1082 ( U4092 , DATAI_9_ , U3149 );
nand NAND2_1083 ( U4093 , U3029 , SUB_84_U25 );
nand NAND2_1084 ( U4094 , U4064 , IR_REG_9_ );
nand NAND2_1085 ( U4095 , DATAI_10_ , U3149 );
nand NAND2_1086 ( U4096 , U3029 , SUB_84_U6 );
nand NAND2_1087 ( U4097 , U4064 , IR_REG_10_ );
nand NAND2_1088 ( U4098 , DATAI_11_ , U3149 );
nand NAND2_1089 ( U4099 , U3029 , SUB_84_U7 );
nand NAND2_1090 ( U4100 , U4064 , IR_REG_11_ );
nand NAND2_1091 ( U4101 , DATAI_12_ , U3149 );
nand NAND2_1092 ( U4102 , U3029 , SUB_84_U89 );
nand NAND2_1093 ( U4103 , U4064 , IR_REG_12_ );
nand NAND2_1094 ( U4104 , DATAI_13_ , U3149 );
nand NAND2_1095 ( U4105 , U3029 , SUB_84_U8 );
nand NAND2_1096 ( U4106 , U4064 , IR_REG_13_ );
nand NAND2_1097 ( U4107 , DATAI_14_ , U3149 );
nand NAND2_1098 ( U4108 , U3029 , SUB_84_U9 );
nand NAND2_1099 ( U4109 , U4064 , IR_REG_14_ );
nand NAND2_1100 ( U4110 , DATAI_15_ , U3149 );
nand NAND2_1101 ( U4111 , U3029 , SUB_84_U10 );
nand NAND2_1102 ( U4112 , U4064 , IR_REG_15_ );
nand NAND2_1103 ( U4113 , DATAI_16_ , U3149 );
nand NAND2_1104 ( U4114 , U3029 , SUB_84_U87 );
nand NAND2_1105 ( U4115 , U4064 , IR_REG_16_ );
nand NAND2_1106 ( U4116 , DATAI_17_ , U3149 );
nand NAND2_1107 ( U4117 , U3029 , SUB_84_U11 );
nand NAND2_1108 ( U4118 , U4064 , IR_REG_17_ );
nand NAND2_1109 ( U4119 , DATAI_18_ , U3149 );
nand NAND2_1110 ( U4120 , U3029 , SUB_84_U12 );
nand NAND2_1111 ( U4121 , U4064 , IR_REG_18_ );
nand NAND2_1112 ( U4122 , DATAI_19_ , U3149 );
nand NAND2_1113 ( U4123 , SUB_84_U13 , U3029 );
nand NAND2_1114 ( U4124 , IR_REG_19_ , U4064 );
nand NAND2_1115 ( U4125 , DATAI_20_ , U3149 );
nand NAND2_1116 ( U4126 , SUB_84_U83 , U3029 );
nand NAND2_1117 ( U4127 , IR_REG_20_ , U4064 );
nand NAND2_1118 ( U4128 , DATAI_21_ , U3149 );
nand NAND2_1119 ( U4129 , U3029 , SUB_84_U14 );
nand NAND2_1120 ( U4130 , U4064 , IR_REG_21_ );
nand NAND2_1121 ( U4131 , DATAI_22_ , U3149 );
nand NAND2_1122 ( U4132 , U3029 , SUB_84_U15 );
nand NAND2_1123 ( U4133 , U4064 , IR_REG_22_ );
nand NAND2_1124 ( U4134 , DATAI_23_ , U3149 );
nand NAND2_1125 ( U4135 , U3029 , SUB_84_U81 );
nand NAND2_1126 ( U4136 , U4064 , IR_REG_23_ );
nand NAND2_1127 ( U4137 , DATAI_24_ , U3149 );
nand NAND2_1128 ( U4138 , U3029 , SUB_84_U78 );
nand NAND2_1129 ( U4139 , U4064 , IR_REG_24_ );
nand NAND2_1130 ( U4140 , DATAI_25_ , U3149 );
nand NAND2_1131 ( U4141 , U3029 , SUB_84_U16 );
nand NAND2_1132 ( U4142 , U4064 , IR_REG_25_ );
nand NAND2_1133 ( U4143 , DATAI_26_ , U3149 );
nand NAND2_1134 ( U4144 , U3029 , SUB_84_U17 );
nand NAND2_1135 ( U4145 , U4064 , IR_REG_26_ );
nand NAND2_1136 ( U4146 , DATAI_27_ , U3149 );
nand NAND2_1137 ( U4147 , U3029 , SUB_84_U76 );
nand NAND2_1138 ( U4148 , U4064 , IR_REG_27_ );
nand NAND2_1139 ( U4149 , DATAI_28_ , U3149 );
nand NAND2_1140 ( U4150 , U3029 , SUB_84_U18 );
nand NAND2_1141 ( U4151 , U4064 , IR_REG_28_ );
nand NAND2_1142 ( U4152 , DATAI_29_ , U3149 );
nand NAND2_1143 ( U4153 , SUB_84_U19 , U3029 );
nand NAND2_1144 ( U4154 , IR_REG_29_ , U4064 );
nand NAND2_1145 ( U4155 , DATAI_30_ , U3149 );
nand NAND2_1146 ( U4156 , SUB_84_U73 , U3029 );
nand NAND2_1147 ( U4157 , IR_REG_30_ , U4064 );
nand NAND2_1148 ( U4158 , DATAI_31_ , U3149 );
nand NAND2_1149 ( U4159 , SUB_84_U49 , U3029 );
nand NAND2_1150 ( U4160 , IR_REG_31_ , U4064 );
not NOT1_1151 ( U4161 , U3360 );
nand NAND2_1152 ( U4162 , U3358 , U5751 );
nand NAND2_1153 ( U4163 , U3358 , U5757 );
nand NAND2_1154 ( U4164 , U4161 , D_REG_10_ );
nand NAND2_1155 ( U4165 , U4161 , D_REG_11_ );
nand NAND2_1156 ( U4166 , U4161 , D_REG_12_ );
nand NAND2_1157 ( U4167 , U4161 , D_REG_13_ );
nand NAND2_1158 ( U4168 , U4161 , D_REG_14_ );
nand NAND2_1159 ( U4169 , U4161 , D_REG_15_ );
nand NAND2_1160 ( U4170 , U4161 , D_REG_16_ );
nand NAND2_1161 ( U4171 , U4161 , D_REG_17_ );
nand NAND2_1162 ( U4172 , U4161 , D_REG_18_ );
nand NAND2_1163 ( U4173 , U4161 , D_REG_19_ );
nand NAND2_1164 ( U4174 , U4161 , D_REG_20_ );
nand NAND2_1165 ( U4175 , U4161 , D_REG_21_ );
nand NAND2_1166 ( U4176 , U4161 , D_REG_22_ );
nand NAND2_1167 ( U4177 , U4161 , D_REG_23_ );
nand NAND2_1168 ( U4178 , U4161 , D_REG_24_ );
nand NAND2_1169 ( U4179 , U4161 , D_REG_25_ );
nand NAND2_1170 ( U4180 , U4161 , D_REG_26_ );
nand NAND2_1171 ( U4181 , U4161 , D_REG_27_ );
nand NAND2_1172 ( U4182 , U4161 , D_REG_28_ );
nand NAND2_1173 ( U4183 , U4161 , D_REG_29_ );
nand NAND2_1174 ( U4184 , U4161 , D_REG_2_ );
nand NAND2_1175 ( U4185 , U4161 , D_REG_30_ );
nand NAND2_1176 ( U4186 , U4161 , D_REG_31_ );
nand NAND2_1177 ( U4187 , U4161 , D_REG_3_ );
nand NAND2_1178 ( U4188 , U4161 , D_REG_4_ );
nand NAND2_1179 ( U4189 , U4161 , D_REG_5_ );
nand NAND2_1180 ( U4190 , U4161 , D_REG_6_ );
nand NAND2_1181 ( U4191 , U4161 , D_REG_7_ );
nand NAND2_1182 ( U4192 , U4161 , D_REG_8_ );
nand NAND2_1183 ( U4193 , U4161 , D_REG_9_ );
nand NAND2_1184 ( U4194 , U5820 , U5817 );
nand NAND4_1185 ( U4195 , U4194 , U3374 , U5831 , U5830 );
nand NAND2_1186 ( U4196 , U3019 , REG2_REG_1_ );
nand NAND2_1187 ( U4197 , U3020 , REG1_REG_1_ );
nand NAND2_1188 ( U4198 , U3021 , REG0_REG_1_ );
nand NAND2_1189 ( U4199 , REG3_REG_1_ , U3018 );
not NOT1_1190 ( U4200 , U3075 );
not NOT1_1191 ( U4201 , U3361 );
nand NAND2_1192 ( U4202 , U4016 , R1150_U31 );
nand NAND2_1193 ( U4203 , U4018 , R1117_U30 );
nand NAND2_1194 ( U4204 , U4017 , R1138_U108 );
nand NAND2_1195 ( U4205 , U4014 , R1192_U32 );
nand NAND2_1196 ( U4206 , U4013 , R1207_U32 );
nand NAND2_1197 ( U4207 , U4024 , R1171_U108 );
nand NAND2_1198 ( U4208 , U4022 , R1240_U108 );
not NOT1_1199 ( U4209 , U3375 );
nand NAND2_1200 ( U4210 , R1222_U104 , U3027 );
nand NAND2_1201 ( U4211 , U3026 , U3075 );
nand NAND2_1202 ( U4212 , U3464 , U3024 );
nand NAND2_1203 ( U4213 , U3464 , U4021 );
nand NAND2_1204 ( U4214 , U3649 , U4209 );
nand NAND2_1205 ( U4215 , REG2_REG_2_ , U3019 );
nand NAND2_1206 ( U4216 , REG1_REG_2_ , U3020 );
nand NAND2_1207 ( U4217 , REG0_REG_2_ , U3021 );
nand NAND2_1208 ( U4218 , REG3_REG_2_ , U3018 );
not NOT1_1209 ( U4219 , U3065 );
nand NAND2_1210 ( U4220 , REG0_REG_0_ , U3021 );
nand NAND2_1211 ( U4221 , REG1_REG_0_ , U3020 );
nand NAND2_1212 ( U4222 , REG2_REG_0_ , U3019 );
nand NAND2_1213 ( U4223 , REG3_REG_0_ , U3018 );
not NOT1_1214 ( U4224 , U3074 );
nand NAND2_1215 ( U4225 , U3034 , U3074 );
nand NAND2_1216 ( U4226 , R1150_U114 , U4016 );
nand NAND2_1217 ( U4227 , R1117_U113 , U4018 );
nand NAND2_1218 ( U4228 , R1138_U107 , U4017 );
nand NAND2_1219 ( U4229 , R1192_U114 , U4014 );
nand NAND2_1220 ( U4230 , R1207_U114 , U4013 );
nand NAND2_1221 ( U4231 , R1171_U107 , U4024 );
nand NAND2_1222 ( U4232 , R1240_U107 , U4022 );
not NOT1_1223 ( U4233 , U3377 );
nand NAND2_1224 ( U4234 , R1222_U103 , U3027 );
nand NAND2_1225 ( U4235 , U3026 , U3065 );
nand NAND2_1226 ( U4236 , R1282_U31 , U3024 );
nand NAND2_1227 ( U4237 , U3468 , U4021 );
nand NAND2_1228 ( U4238 , U3665 , U4233 );
nand NAND2_1229 ( U4239 , REG2_REG_3_ , U3019 );
nand NAND2_1230 ( U4240 , REG1_REG_3_ , U3020 );
nand NAND2_1231 ( U4241 , REG0_REG_3_ , U3021 );
nand NAND2_1232 ( U4242 , ADD_95_U4 , U3018 );
not NOT1_1233 ( U4243 , U3061 );
nand NAND2_1234 ( U4244 , U3034 , U3075 );
nand NAND2_1235 ( U4245 , R1150_U124 , U4016 );
nand NAND2_1236 ( U4246 , R1117_U123 , U4018 );
nand NAND2_1237 ( U4247 , R1138_U24 , U4017 );
nand NAND2_1238 ( U4248 , R1192_U124 , U4014 );
nand NAND2_1239 ( U4249 , R1207_U124 , U4013 );
nand NAND2_1240 ( U4250 , R1171_U24 , U4024 );
nand NAND2_1241 ( U4251 , R1240_U24 , U4022 );
not NOT1_1242 ( U4252 , U3378 );
nand NAND2_1243 ( U4253 , R1222_U23 , U3027 );
nand NAND2_1244 ( U4254 , U3026 , U3061 );
nand NAND2_1245 ( U4255 , R1282_U6 , U3024 );
nand NAND2_1246 ( U4256 , U3470 , U4021 );
nand NAND2_1247 ( U4257 , U3669 , U4252 );
nand NAND2_1248 ( U4258 , REG2_REG_4_ , U3019 );
nand NAND2_1249 ( U4259 , REG1_REG_4_ , U3020 );
nand NAND2_1250 ( U4260 , REG0_REG_4_ , U3021 );
nand NAND2_1251 ( U4261 , ADD_95_U51 , U3018 );
not NOT1_1252 ( U4262 , U3057 );
nand NAND2_1253 ( U4263 , U3034 , U3065 );
nand NAND2_1254 ( U4264 , R1150_U28 , U4016 );
nand NAND2_1255 ( U4265 , R1117_U27 , U4018 );
nand NAND2_1256 ( U4266 , R1138_U113 , U4017 );
nand NAND2_1257 ( U4267 , R1192_U29 , U4014 );
nand NAND2_1258 ( U4268 , R1207_U29 , U4013 );
nand NAND2_1259 ( U4269 , R1171_U113 , U4024 );
nand NAND2_1260 ( U4270 , R1240_U113 , U4022 );
not NOT1_1261 ( U4271 , U3379 );
nand NAND2_1262 ( U4272 , R1222_U109 , U3027 );
nand NAND2_1263 ( U4273 , U3026 , U3057 );
nand NAND2_1264 ( U4274 , R1282_U7 , U3024 );
nand NAND2_1265 ( U4275 , U3472 , U4021 );
nand NAND2_1266 ( U4276 , U3673 , U4271 );
nand NAND2_1267 ( U4277 , REG2_REG_5_ , U3019 );
nand NAND2_1268 ( U4278 , REG1_REG_5_ , U3020 );
nand NAND2_1269 ( U4279 , REG0_REG_5_ , U3021 );
nand NAND2_1270 ( U4280 , ADD_95_U50 , U3018 );
not NOT1_1271 ( U4281 , U3064 );
nand NAND2_1272 ( U4282 , U3034 , U3061 );
nand NAND2_1273 ( U4283 , R1150_U123 , U4016 );
nand NAND2_1274 ( U4284 , R1117_U122 , U4018 );
nand NAND2_1275 ( U4285 , R1138_U112 , U4017 );
nand NAND2_1276 ( U4286 , R1192_U123 , U4014 );
nand NAND2_1277 ( U4287 , R1207_U123 , U4013 );
nand NAND2_1278 ( U4288 , R1171_U112 , U4024 );
nand NAND2_1279 ( U4289 , R1240_U112 , U4022 );
not NOT1_1280 ( U4290 , U3380 );
nand NAND2_1281 ( U4291 , R1222_U108 , U3027 );
nand NAND2_1282 ( U4292 , U3026 , U3064 );
nand NAND2_1283 ( U4293 , R1282_U8 , U3024 );
nand NAND2_1284 ( U4294 , U3474 , U4021 );
nand NAND2_1285 ( U4295 , U3677 , U4290 );
nand NAND2_1286 ( U4296 , REG2_REG_6_ , U3019 );
nand NAND2_1287 ( U4297 , REG1_REG_6_ , U3020 );
nand NAND2_1288 ( U4298 , REG0_REG_6_ , U3021 );
nand NAND2_1289 ( U4299 , ADD_95_U49 , U3018 );
not NOT1_1290 ( U4300 , U3068 );
nand NAND2_1291 ( U4301 , U3034 , U3057 );
nand NAND2_1292 ( U4302 , R1150_U122 , U4016 );
nand NAND2_1293 ( U4303 , R1117_U121 , U4018 );
nand NAND2_1294 ( U4304 , R1138_U25 , U4017 );
nand NAND2_1295 ( U4305 , R1192_U122 , U4014 );
nand NAND2_1296 ( U4306 , R1207_U122 , U4013 );
nand NAND2_1297 ( U4307 , R1171_U25 , U4024 );
nand NAND2_1298 ( U4308 , R1240_U25 , U4022 );
not NOT1_1299 ( U4309 , U3381 );
nand NAND2_1300 ( U4310 , R1222_U24 , U3027 );
nand NAND2_1301 ( U4311 , U3026 , U3068 );
nand NAND2_1302 ( U4312 , R1282_U9 , U3024 );
nand NAND2_1303 ( U4313 , U3476 , U4021 );
nand NAND2_1304 ( U4314 , U3681 , U4309 );
nand NAND2_1305 ( U4315 , REG2_REG_7_ , U3019 );
nand NAND2_1306 ( U4316 , REG1_REG_7_ , U3020 );
nand NAND2_1307 ( U4317 , REG0_REG_7_ , U3021 );
nand NAND2_1308 ( U4318 , ADD_95_U48 , U3018 );
not NOT1_1309 ( U4319 , U3067 );
nand NAND2_1310 ( U4320 , U3034 , U3064 );
nand NAND2_1311 ( U4321 , R1150_U29 , U4016 );
nand NAND2_1312 ( U4322 , R1117_U28 , U4018 );
nand NAND2_1313 ( U4323 , R1138_U111 , U4017 );
nand NAND2_1314 ( U4324 , R1192_U30 , U4014 );
nand NAND2_1315 ( U4325 , R1207_U30 , U4013 );
nand NAND2_1316 ( U4326 , R1171_U111 , U4024 );
nand NAND2_1317 ( U4327 , R1240_U111 , U4022 );
not NOT1_1318 ( U4328 , U3382 );
nand NAND2_1319 ( U4329 , R1222_U107 , U3027 );
nand NAND2_1320 ( U4330 , U3026 , U3067 );
nand NAND2_1321 ( U4331 , R1282_U10 , U3024 );
nand NAND2_1322 ( U4332 , U3478 , U4021 );
nand NAND2_1323 ( U4333 , U3685 , U4328 );
nand NAND2_1324 ( U4334 , REG2_REG_8_ , U3019 );
nand NAND2_1325 ( U4335 , REG1_REG_8_ , U3020 );
nand NAND2_1326 ( U4336 , REG0_REG_8_ , U3021 );
nand NAND2_1327 ( U4337 , ADD_95_U47 , U3018 );
not NOT1_1328 ( U4338 , U3081 );
nand NAND2_1329 ( U4339 , U3034 , U3068 );
nand NAND2_1330 ( U4340 , R1150_U121 , U4016 );
nand NAND2_1331 ( U4341 , R1117_U120 , U4018 );
nand NAND2_1332 ( U4342 , R1138_U26 , U4017 );
nand NAND2_1333 ( U4343 , R1192_U121 , U4014 );
nand NAND2_1334 ( U4344 , R1207_U121 , U4013 );
nand NAND2_1335 ( U4345 , R1171_U26 , U4024 );
nand NAND2_1336 ( U4346 , R1240_U26 , U4022 );
not NOT1_1337 ( U4347 , U3383 );
nand NAND2_1338 ( U4348 , R1222_U25 , U3027 );
nand NAND2_1339 ( U4349 , U3026 , U3081 );
nand NAND2_1340 ( U4350 , R1282_U11 , U3024 );
nand NAND2_1341 ( U4351 , U3480 , U4021 );
nand NAND2_1342 ( U4352 , U3689 , U4347 );
nand NAND2_1343 ( U4353 , REG2_REG_9_ , U3019 );
nand NAND2_1344 ( U4354 , REG1_REG_9_ , U3020 );
nand NAND2_1345 ( U4355 , REG0_REG_9_ , U3021 );
nand NAND2_1346 ( U4356 , ADD_95_U46 , U3018 );
not NOT1_1347 ( U4357 , U3080 );
nand NAND2_1348 ( U4358 , U3034 , U3067 );
nand NAND2_1349 ( U4359 , R1150_U30 , U4016 );
nand NAND2_1350 ( U4360 , R1117_U29 , U4018 );
nand NAND2_1351 ( U4361 , R1138_U110 , U4017 );
nand NAND2_1352 ( U4362 , R1192_U31 , U4014 );
nand NAND2_1353 ( U4363 , R1207_U31 , U4013 );
nand NAND2_1354 ( U4364 , R1171_U110 , U4024 );
nand NAND2_1355 ( U4365 , R1240_U110 , U4022 );
not NOT1_1356 ( U4366 , U3384 );
nand NAND2_1357 ( U4367 , R1222_U106 , U3027 );
nand NAND2_1358 ( U4368 , U3026 , U3080 );
nand NAND2_1359 ( U4369 , R1282_U36 , U3024 );
nand NAND2_1360 ( U4370 , U3482 , U4021 );
nand NAND2_1361 ( U4371 , U3693 , U4366 );
nand NAND2_1362 ( U4372 , REG2_REG_10_ , U3019 );
nand NAND2_1363 ( U4373 , REG1_REG_10_ , U3020 );
nand NAND2_1364 ( U4374 , REG0_REG_10_ , U3021 );
nand NAND2_1365 ( U4375 , ADD_95_U70 , U3018 );
not NOT1_1366 ( U4376 , U3059 );
nand NAND2_1367 ( U4377 , U3034 , U3081 );
nand NAND2_1368 ( U4378 , R1150_U120 , U4016 );
nand NAND2_1369 ( U4379 , R1117_U119 , U4018 );
nand NAND2_1370 ( U4380 , R1138_U109 , U4017 );
nand NAND2_1371 ( U4381 , R1192_U120 , U4014 );
nand NAND2_1372 ( U4382 , R1207_U120 , U4013 );
nand NAND2_1373 ( U4383 , R1171_U109 , U4024 );
nand NAND2_1374 ( U4384 , R1240_U109 , U4022 );
not NOT1_1375 ( U4385 , U3385 );
nand NAND2_1376 ( U4386 , R1222_U105 , U3027 );
nand NAND2_1377 ( U4387 , U3026 , U3059 );
nand NAND2_1378 ( U4388 , R1282_U33 , U3024 );
nand NAND2_1379 ( U4389 , U3484 , U4021 );
nand NAND2_1380 ( U4390 , U3697 , U4385 );
nand NAND2_1381 ( U4391 , REG2_REG_11_ , U3019 );
nand NAND2_1382 ( U4392 , REG1_REG_11_ , U3020 );
nand NAND2_1383 ( U4393 , REG0_REG_11_ , U3021 );
nand NAND2_1384 ( U4394 , ADD_95_U69 , U3018 );
not NOT1_1385 ( U4395 , U3060 );
nand NAND2_1386 ( U4396 , U3034 , U3080 );
nand NAND2_1387 ( U4397 , R1150_U130 , U4016 );
nand NAND2_1388 ( U4398 , R1117_U129 , U4018 );
nand NAND2_1389 ( U4399 , R1138_U18 , U4017 );
nand NAND2_1390 ( U4400 , R1192_U130 , U4014 );
nand NAND2_1391 ( U4401 , R1207_U130 , U4013 );
nand NAND2_1392 ( U4402 , R1171_U18 , U4024 );
nand NAND2_1393 ( U4403 , R1240_U18 , U4022 );
not NOT1_1394 ( U4404 , U3386 );
nand NAND2_1395 ( U4405 , R1222_U17 , U3027 );
nand NAND2_1396 ( U4406 , U3026 , U3060 );
nand NAND2_1397 ( U4407 , R1282_U94 , U3024 );
nand NAND2_1398 ( U4408 , U3486 , U4021 );
nand NAND2_1399 ( U4409 , U3701 , U4404 );
nand NAND2_1400 ( U4410 , REG2_REG_12_ , U3019 );
nand NAND2_1401 ( U4411 , REG1_REG_12_ , U3020 );
nand NAND2_1402 ( U4412 , REG0_REG_12_ , U3021 );
nand NAND2_1403 ( U4413 , ADD_95_U68 , U3018 );
not NOT1_1404 ( U4414 , U3069 );
nand NAND2_1405 ( U4415 , U3034 , U3059 );
nand NAND2_1406 ( U4416 , R1150_U23 , U4016 );
nand NAND2_1407 ( U4417 , R1117_U23 , U4018 );
nand NAND2_1408 ( U4418 , R1138_U127 , U4017 );
nand NAND2_1409 ( U4419 , R1192_U24 , U4014 );
nand NAND2_1410 ( U4420 , R1207_U24 , U4013 );
nand NAND2_1411 ( U4421 , R1171_U127 , U4024 );
nand NAND2_1412 ( U4422 , R1240_U127 , U4022 );
not NOT1_1413 ( U4423 , U3387 );
nand NAND2_1414 ( U4424 , R1222_U123 , U3027 );
nand NAND2_1415 ( U4425 , U3026 , U3069 );
nand NAND2_1416 ( U4426 , R1282_U91 , U3024 );
nand NAND2_1417 ( U4427 , U3488 , U4021 );
nand NAND2_1418 ( U4428 , U3705 , U4423 );
nand NAND2_1419 ( U4429 , REG2_REG_13_ , U3019 );
nand NAND2_1420 ( U4430 , REG1_REG_13_ , U3020 );
nand NAND2_1421 ( U4431 , REG0_REG_13_ , U3021 );
nand NAND2_1422 ( U4432 , ADD_95_U67 , U3018 );
not NOT1_1423 ( U4433 , U3077 );
nand NAND2_1424 ( U4434 , U3034 , U3060 );
nand NAND2_1425 ( U4435 , R1150_U119 , U4016 );
nand NAND2_1426 ( U4436 , R1117_U118 , U4018 );
nand NAND2_1427 ( U4437 , R1138_U126 , U4017 );
nand NAND2_1428 ( U4438 , R1192_U119 , U4014 );
nand NAND2_1429 ( U4439 , R1207_U119 , U4013 );
nand NAND2_1430 ( U4440 , R1171_U126 , U4024 );
nand NAND2_1431 ( U4441 , R1240_U126 , U4022 );
not NOT1_1432 ( U4442 , U3388 );
nand NAND2_1433 ( U4443 , R1222_U122 , U3027 );
nand NAND2_1434 ( U4444 , U3026 , U3077 );
nand NAND2_1435 ( U4445 , R1282_U89 , U3024 );
nand NAND2_1436 ( U4446 , U3490 , U4021 );
nand NAND2_1437 ( U4447 , U3709 , U4442 );
nand NAND2_1438 ( U4448 , REG2_REG_14_ , U3019 );
nand NAND2_1439 ( U4449 , REG1_REG_14_ , U3020 );
nand NAND2_1440 ( U4450 , REG0_REG_14_ , U3021 );
nand NAND2_1441 ( U4451 , ADD_95_U66 , U3018 );
not NOT1_1442 ( U4452 , U3076 );
nand NAND2_1443 ( U4453 , U3034 , U3069 );
nand NAND2_1444 ( U4454 , R1150_U118 , U4016 );
nand NAND2_1445 ( U4455 , R1117_U117 , U4018 );
nand NAND2_1446 ( U4456 , R1138_U19 , U4017 );
nand NAND2_1447 ( U4457 , R1192_U118 , U4014 );
nand NAND2_1448 ( U4458 , R1207_U118 , U4013 );
nand NAND2_1449 ( U4459 , R1171_U19 , U4024 );
nand NAND2_1450 ( U4460 , R1240_U19 , U4022 );
not NOT1_1451 ( U4461 , U3389 );
nand NAND2_1452 ( U4462 , R1222_U18 , U3027 );
nand NAND2_1453 ( U4463 , U3026 , U3076 );
nand NAND2_1454 ( U4464 , R1282_U86 , U3024 );
nand NAND2_1455 ( U4465 , U3492 , U4021 );
nand NAND2_1456 ( U4466 , U3713 , U4461 );
nand NAND2_1457 ( U4467 , REG2_REG_15_ , U3019 );
nand NAND2_1458 ( U4468 , REG1_REG_15_ , U3020 );
nand NAND2_1459 ( U4469 , REG0_REG_15_ , U3021 );
nand NAND2_1460 ( U4470 , ADD_95_U65 , U3018 );
not NOT1_1461 ( U4471 , U3071 );
nand NAND2_1462 ( U4472 , U3034 , U3077 );
nand NAND2_1463 ( U4473 , R1150_U129 , U4016 );
nand NAND2_1464 ( U4474 , R1117_U128 , U4018 );
nand NAND2_1465 ( U4475 , R1138_U125 , U4017 );
nand NAND2_1466 ( U4476 , R1192_U129 , U4014 );
nand NAND2_1467 ( U4477 , R1207_U129 , U4013 );
nand NAND2_1468 ( U4478 , R1171_U125 , U4024 );
nand NAND2_1469 ( U4479 , R1240_U125 , U4022 );
not NOT1_1470 ( U4480 , U3390 );
nand NAND2_1471 ( U4481 , R1222_U121 , U3027 );
nand NAND2_1472 ( U4482 , U3026 , U3071 );
nand NAND2_1473 ( U4483 , R1282_U84 , U3024 );
nand NAND2_1474 ( U4484 , U3494 , U4021 );
nand NAND2_1475 ( U4485 , U3717 , U4480 );
nand NAND2_1476 ( U4486 , REG2_REG_16_ , U3019 );
nand NAND2_1477 ( U4487 , REG1_REG_16_ , U3020 );
nand NAND2_1478 ( U4488 , REG0_REG_16_ , U3021 );
nand NAND2_1479 ( U4489 , ADD_95_U64 , U3018 );
not NOT1_1480 ( U4490 , U3070 );
nand NAND2_1481 ( U4491 , U3034 , U3076 );
nand NAND2_1482 ( U4492 , R1150_U128 , U4016 );
nand NAND2_1483 ( U4493 , R1117_U127 , U4018 );
nand NAND2_1484 ( U4494 , R1138_U124 , U4017 );
nand NAND2_1485 ( U4495 , R1192_U128 , U4014 );
nand NAND2_1486 ( U4496 , R1207_U128 , U4013 );
nand NAND2_1487 ( U4497 , R1171_U124 , U4024 );
nand NAND2_1488 ( U4498 , R1240_U124 , U4022 );
not NOT1_1489 ( U4499 , U3391 );
nand NAND2_1490 ( U4500 , R1222_U120 , U3027 );
nand NAND2_1491 ( U4501 , U3026 , U3070 );
nand NAND2_1492 ( U4502 , R1282_U81 , U3024 );
nand NAND2_1493 ( U4503 , U3496 , U4021 );
nand NAND2_1494 ( U4504 , U3721 , U4499 );
nand NAND2_1495 ( U4505 , REG2_REG_17_ , U3019 );
nand NAND2_1496 ( U4506 , REG1_REG_17_ , U3020 );
nand NAND2_1497 ( U4507 , REG0_REG_17_ , U3021 );
nand NAND2_1498 ( U4508 , ADD_95_U63 , U3018 );
not NOT1_1499 ( U4509 , U3066 );
nand NAND2_1500 ( U4510 , U3034 , U3071 );
nand NAND2_1501 ( U4511 , R1150_U24 , U4016 );
nand NAND2_1502 ( U4512 , R1117_U24 , U4018 );
nand NAND2_1503 ( U4513 , R1138_U123 , U4017 );
nand NAND2_1504 ( U4514 , R1192_U25 , U4014 );
nand NAND2_1505 ( U4515 , R1207_U25 , U4013 );
nand NAND2_1506 ( U4516 , R1171_U123 , U4024 );
nand NAND2_1507 ( U4517 , R1240_U123 , U4022 );
not NOT1_1508 ( U4518 , U3392 );
nand NAND2_1509 ( U4519 , R1222_U119 , U3027 );
nand NAND2_1510 ( U4520 , U3026 , U3066 );
nand NAND2_1511 ( U4521 , R1282_U79 , U3024 );
nand NAND2_1512 ( U4522 , U3498 , U4021 );
nand NAND2_1513 ( U4523 , U3725 , U4518 );
nand NAND2_1514 ( U4524 , REG2_REG_18_ , U3019 );
nand NAND2_1515 ( U4525 , REG1_REG_18_ , U3020 );
nand NAND2_1516 ( U4526 , REG0_REG_18_ , U3021 );
nand NAND2_1517 ( U4527 , ADD_95_U62 , U3018 );
not NOT1_1518 ( U4528 , U3079 );
nand NAND2_1519 ( U4529 , U3034 , U3070 );
nand NAND2_1520 ( U4530 , R1150_U117 , U4016 );
nand NAND2_1521 ( U4531 , R1117_U116 , U4018 );
nand NAND2_1522 ( U4532 , R1138_U20 , U4017 );
nand NAND2_1523 ( U4533 , R1192_U117 , U4014 );
nand NAND2_1524 ( U4534 , R1207_U117 , U4013 );
nand NAND2_1525 ( U4535 , R1171_U20 , U4024 );
nand NAND2_1526 ( U4536 , R1240_U20 , U4022 );
not NOT1_1527 ( U4537 , U3393 );
nand NAND2_1528 ( U4538 , R1222_U19 , U3027 );
nand NAND2_1529 ( U4539 , U3026 , U3079 );
nand NAND2_1530 ( U4540 , R1282_U76 , U3024 );
nand NAND2_1531 ( U4541 , U3500 , U4021 );
nand NAND2_1532 ( U4542 , U3729 , U4537 );
nand NAND2_1533 ( U4543 , REG2_REG_19_ , U3019 );
nand NAND2_1534 ( U4544 , REG1_REG_19_ , U3020 );
nand NAND2_1535 ( U4545 , REG0_REG_19_ , U3021 );
nand NAND2_1536 ( U4546 , ADD_95_U61 , U3018 );
not NOT1_1537 ( U4547 , U3078 );
nand NAND2_1538 ( U4548 , U3034 , U3066 );
nand NAND2_1539 ( U4549 , R1150_U116 , U4016 );
nand NAND2_1540 ( U4550 , R1117_U115 , U4018 );
nand NAND2_1541 ( U4551 , R1138_U122 , U4017 );
nand NAND2_1542 ( U4552 , R1192_U116 , U4014 );
nand NAND2_1543 ( U4553 , R1207_U116 , U4013 );
nand NAND2_1544 ( U4554 , R1171_U122 , U4024 );
nand NAND2_1545 ( U4555 , R1240_U122 , U4022 );
not NOT1_1546 ( U4556 , U3394 );
nand NAND2_1547 ( U4557 , R1222_U118 , U3027 );
nand NAND2_1548 ( U4558 , U3026 , U3078 );
nand NAND2_1549 ( U4559 , R1282_U74 , U3024 );
nand NAND2_1550 ( U4560 , U3502 , U4021 );
nand NAND2_1551 ( U4561 , U3733 , U4556 );
nand NAND2_1552 ( U4562 , REG2_REG_20_ , U3019 );
nand NAND2_1553 ( U4563 , REG1_REG_20_ , U3020 );
nand NAND2_1554 ( U4564 , REG0_REG_20_ , U3021 );
nand NAND2_1555 ( U4565 , ADD_95_U60 , U3018 );
not NOT1_1556 ( U4566 , U3073 );
nand NAND2_1557 ( U4567 , U3034 , U3079 );
nand NAND2_1558 ( U4568 , R1150_U115 , U4016 );
nand NAND2_1559 ( U4569 , R1117_U114 , U4018 );
nand NAND2_1560 ( U4570 , R1138_U121 , U4017 );
nand NAND2_1561 ( U4571 , R1192_U115 , U4014 );
nand NAND2_1562 ( U4572 , R1207_U115 , U4013 );
nand NAND2_1563 ( U4573 , R1171_U121 , U4024 );
nand NAND2_1564 ( U4574 , R1240_U121 , U4022 );
not NOT1_1565 ( U4575 , U3395 );
nand NAND2_1566 ( U4576 , R1222_U117 , U3027 );
nand NAND2_1567 ( U4577 , U3026 , U3073 );
nand NAND2_1568 ( U4578 , R1282_U71 , U3024 );
nand NAND2_1569 ( U4579 , U3504 , U4021 );
nand NAND2_1570 ( U4580 , U3737 , U4575 );
nand NAND2_1571 ( U4581 , REG2_REG_21_ , U3019 );
nand NAND2_1572 ( U4582 , REG1_REG_21_ , U3020 );
nand NAND2_1573 ( U4583 , REG0_REG_21_ , U3021 );
nand NAND2_1574 ( U4584 , ADD_95_U59 , U3018 );
not NOT1_1575 ( U4585 , U3072 );
nand NAND2_1576 ( U4586 , U3034 , U3078 );
nand NAND2_1577 ( U4587 , R1150_U113 , U4016 );
nand NAND2_1578 ( U4588 , R1117_U112 , U4018 );
nand NAND2_1579 ( U4589 , R1138_U21 , U4017 );
nand NAND2_1580 ( U4590 , R1192_U113 , U4014 );
nand NAND2_1581 ( U4591 , R1207_U113 , U4013 );
nand NAND2_1582 ( U4592 , R1171_U21 , U4024 );
nand NAND2_1583 ( U4593 , R1240_U21 , U4022 );
not NOT1_1584 ( U4594 , U3397 );
nand NAND2_1585 ( U4595 , R1222_U20 , U3027 );
nand NAND2_1586 ( U4596 , U3026 , U3072 );
nand NAND2_1587 ( U4597 , R1282_U67 , U3024 );
nand NAND2_1588 ( U4598 , U4037 , U4021 );
nand NAND2_1589 ( U4599 , U3741 , U4594 );
nand NAND2_1590 ( U4600 , REG2_REG_22_ , U3019 );
nand NAND2_1591 ( U4601 , REG1_REG_22_ , U3020 );
nand NAND2_1592 ( U4602 , REG0_REG_22_ , U3021 );
nand NAND2_1593 ( U4603 , ADD_95_U58 , U3018 );
not NOT1_1594 ( U4604 , U3058 );
nand NAND2_1595 ( U4605 , U3034 , U3073 );
nand NAND2_1596 ( U4606 , R1150_U127 , U4016 );
nand NAND2_1597 ( U4607 , R1117_U126 , U4018 );
nand NAND2_1598 ( U4608 , R1138_U22 , U4017 );
nand NAND2_1599 ( U4609 , R1192_U127 , U4014 );
nand NAND2_1600 ( U4610 , R1207_U127 , U4013 );
nand NAND2_1601 ( U4611 , R1171_U22 , U4024 );
nand NAND2_1602 ( U4612 , R1240_U22 , U4022 );
not NOT1_1603 ( U4613 , U3399 );
nand NAND2_1604 ( U4614 , R1222_U21 , U3027 );
nand NAND2_1605 ( U4615 , U3026 , U3058 );
nand NAND2_1606 ( U4616 , R1282_U64 , U3024 );
nand NAND2_1607 ( U4617 , U4036 , U4021 );
nand NAND2_1608 ( U4618 , U3745 , U4613 );
nand NAND2_1609 ( U4619 , REG2_REG_23_ , U3019 );
nand NAND2_1610 ( U4620 , REG1_REG_23_ , U3020 );
nand NAND2_1611 ( U4621 , REG0_REG_23_ , U3021 );
nand NAND2_1612 ( U4622 , ADD_95_U57 , U3018 );
not NOT1_1613 ( U4623 , U3063 );
nand NAND2_1614 ( U4624 , U3034 , U3072 );
nand NAND2_1615 ( U4625 , R1150_U126 , U4016 );
nand NAND2_1616 ( U4626 , R1117_U125 , U4018 );
nand NAND2_1617 ( U4627 , R1138_U120 , U4017 );
nand NAND2_1618 ( U4628 , R1192_U126 , U4014 );
nand NAND2_1619 ( U4629 , R1207_U126 , U4013 );
nand NAND2_1620 ( U4630 , R1171_U120 , U4024 );
nand NAND2_1621 ( U4631 , R1240_U120 , U4022 );
not NOT1_1622 ( U4632 , U3401 );
nand NAND2_1623 ( U4633 , R1222_U116 , U3027 );
nand NAND2_1624 ( U4634 , U3026 , U3063 );
nand NAND2_1625 ( U4635 , R1282_U62 , U3024 );
nand NAND2_1626 ( U4636 , U4035 , U4021 );
nand NAND2_1627 ( U4637 , U3749 , U4632 );
nand NAND2_1628 ( U4638 , REG2_REG_24_ , U3019 );
nand NAND2_1629 ( U4639 , REG1_REG_24_ , U3020 );
nand NAND2_1630 ( U4640 , REG0_REG_24_ , U3021 );
nand NAND2_1631 ( U4641 , ADD_95_U56 , U3018 );
not NOT1_1632 ( U4642 , U3062 );
nand NAND2_1633 ( U4643 , U3034 , U3058 );
nand NAND2_1634 ( U4644 , R1150_U25 , U4016 );
nand NAND2_1635 ( U4645 , R1117_U25 , U4018 );
nand NAND2_1636 ( U4646 , R1138_U119 , U4017 );
nand NAND2_1637 ( U4647 , R1192_U26 , U4014 );
nand NAND2_1638 ( U4648 , R1207_U26 , U4013 );
nand NAND2_1639 ( U4649 , R1171_U119 , U4024 );
nand NAND2_1640 ( U4650 , R1240_U119 , U4022 );
not NOT1_1641 ( U4651 , U3403 );
nand NAND2_1642 ( U4652 , R1222_U115 , U3027 );
nand NAND2_1643 ( U4653 , U3026 , U3062 );
nand NAND2_1644 ( U4654 , R1282_U59 , U3024 );
nand NAND2_1645 ( U4655 , U4034 , U4021 );
nand NAND2_1646 ( U4656 , U3753 , U4651 );
nand NAND2_1647 ( U4657 , REG2_REG_25_ , U3019 );
nand NAND2_1648 ( U4658 , REG1_REG_25_ , U3020 );
nand NAND2_1649 ( U4659 , REG0_REG_25_ , U3021 );
nand NAND2_1650 ( U4660 , ADD_95_U55 , U3018 );
not NOT1_1651 ( U4661 , U3055 );
nand NAND2_1652 ( U4662 , U3034 , U3063 );
nand NAND2_1653 ( U4663 , R1150_U112 , U4016 );
nand NAND2_1654 ( U4664 , R1117_U111 , U4018 );
nand NAND2_1655 ( U4665 , R1138_U118 , U4017 );
nand NAND2_1656 ( U4666 , R1192_U112 , U4014 );
nand NAND2_1657 ( U4667 , R1207_U112 , U4013 );
nand NAND2_1658 ( U4668 , R1171_U118 , U4024 );
nand NAND2_1659 ( U4669 , R1240_U118 , U4022 );
not NOT1_1660 ( U4670 , U3405 );
nand NAND2_1661 ( U4671 , R1222_U114 , U3027 );
nand NAND2_1662 ( U4672 , U3026 , U3055 );
nand NAND2_1663 ( U4673 , R1282_U57 , U3024 );
nand NAND2_1664 ( U4674 , U4033 , U4021 );
nand NAND2_1665 ( U4675 , U3757 , U4670 );
nand NAND2_1666 ( U4676 , REG2_REG_26_ , U3019 );
nand NAND2_1667 ( U4677 , REG1_REG_26_ , U3020 );
nand NAND2_1668 ( U4678 , REG0_REG_26_ , U3021 );
nand NAND2_1669 ( U4679 , ADD_95_U54 , U3018 );
not NOT1_1670 ( U4680 , U3054 );
nand NAND2_1671 ( U4681 , U3034 , U3062 );
nand NAND2_1672 ( U4682 , R1150_U111 , U4016 );
nand NAND2_1673 ( U4683 , R1117_U110 , U4018 );
nand NAND2_1674 ( U4684 , R1138_U117 , U4017 );
nand NAND2_1675 ( U4685 , R1192_U111 , U4014 );
nand NAND2_1676 ( U4686 , R1207_U111 , U4013 );
nand NAND2_1677 ( U4687 , R1171_U117 , U4024 );
nand NAND2_1678 ( U4688 , R1240_U117 , U4022 );
not NOT1_1679 ( U4689 , U3407 );
nand NAND2_1680 ( U4690 , R1222_U113 , U3027 );
nand NAND2_1681 ( U4691 , U3026 , U3054 );
nand NAND2_1682 ( U4692 , R1282_U54 , U3024 );
nand NAND2_1683 ( U4693 , U4032 , U4021 );
nand NAND2_1684 ( U4694 , U3761 , U4689 );
nand NAND2_1685 ( U4695 , REG2_REG_27_ , U3019 );
nand NAND2_1686 ( U4696 , REG1_REG_27_ , U3020 );
nand NAND2_1687 ( U4697 , REG0_REG_27_ , U3021 );
nand NAND2_1688 ( U4698 , ADD_95_U53 , U3018 );
not NOT1_1689 ( U4699 , U3050 );
nand NAND2_1690 ( U4700 , U3034 , U3055 );
nand NAND2_1691 ( U4701 , R1150_U125 , U4016 );
nand NAND2_1692 ( U4702 , R1117_U124 , U4018 );
nand NAND2_1693 ( U4703 , R1138_U23 , U4017 );
nand NAND2_1694 ( U4704 , R1192_U125 , U4014 );
nand NAND2_1695 ( U4705 , R1207_U125 , U4013 );
nand NAND2_1696 ( U4706 , R1171_U23 , U4024 );
nand NAND2_1697 ( U4707 , R1240_U23 , U4022 );
not NOT1_1698 ( U4708 , U3409 );
nand NAND2_1699 ( U4709 , R1222_U22 , U3027 );
nand NAND2_1700 ( U4710 , U3026 , U3050 );
nand NAND2_1701 ( U4711 , R1282_U52 , U3024 );
nand NAND2_1702 ( U4712 , U4031 , U4021 );
nand NAND2_1703 ( U4713 , U3765 , U4708 );
nand NAND2_1704 ( U4714 , REG2_REG_28_ , U3019 );
nand NAND2_1705 ( U4715 , REG1_REG_28_ , U3020 );
nand NAND2_1706 ( U4716 , REG0_REG_28_ , U3021 );
nand NAND2_1707 ( U4717 , ADD_95_U52 , U3018 );
not NOT1_1708 ( U4718 , U3051 );
nand NAND2_1709 ( U4719 , U3034 , U3054 );
nand NAND2_1710 ( U4720 , R1150_U26 , U4016 );
nand NAND2_1711 ( U4721 , R1117_U31 , U4018 );
nand NAND2_1712 ( U4722 , R1138_U116 , U4017 );
nand NAND2_1713 ( U4723 , R1192_U27 , U4014 );
nand NAND2_1714 ( U4724 , R1207_U27 , U4013 );
nand NAND2_1715 ( U4725 , R1171_U116 , U4024 );
nand NAND2_1716 ( U4726 , R1240_U116 , U4022 );
not NOT1_1717 ( U4727 , U3411 );
nand NAND2_1718 ( U4728 , R1222_U112 , U3027 );
nand NAND2_1719 ( U4729 , U3026 , U3051 );
nand NAND2_1720 ( U4730 , R1282_U49 , U3024 );
nand NAND2_1721 ( U4731 , U4030 , U4021 );
nand NAND2_1722 ( U4732 , U3769 , U4727 );
nand NAND2_1723 ( U4733 , ADD_95_U5 , U3018 );
nand NAND2_1724 ( U4734 , REG2_REG_29_ , U3019 );
nand NAND2_1725 ( U4735 , REG1_REG_29_ , U3020 );
nand NAND2_1726 ( U4736 , REG0_REG_29_ , U3021 );
not NOT1_1727 ( U4737 , U3052 );
nand NAND2_1728 ( U4738 , U3034 , U3050 );
nand NAND2_1729 ( U4739 , R1150_U110 , U4016 );
nand NAND2_1730 ( U4740 , R1117_U109 , U4018 );
nand NAND2_1731 ( U4741 , R1138_U115 , U4017 );
nand NAND2_1732 ( U4742 , R1192_U110 , U4014 );
nand NAND2_1733 ( U4743 , R1207_U110 , U4013 );
nand NAND2_1734 ( U4744 , R1171_U115 , U4024 );
nand NAND2_1735 ( U4745 , R1240_U115 , U4022 );
not NOT1_1736 ( U4746 , U3413 );
nand NAND2_1737 ( U4747 , R1222_U111 , U3027 );
nand NAND2_1738 ( U4748 , U3026 , U3052 );
nand NAND2_1739 ( U4749 , R1282_U47 , U3024 );
nand NAND2_1740 ( U4750 , U4029 , U4021 );
nand NAND2_1741 ( U4751 , U3773 , U4746 );
nand NAND2_1742 ( U4752 , REG2_REG_30_ , U3019 );
nand NAND2_1743 ( U4753 , REG1_REG_30_ , U3020 );
nand NAND2_1744 ( U4754 , REG0_REG_30_ , U3021 );
not NOT1_1745 ( U4755 , U3056 );
nand NAND2_1746 ( U4756 , U5799 , U3359 );
nand NAND2_1747 ( U4757 , U3969 , U4756 );
nand NAND2_1748 ( U4758 , U3774 , U3056 );
nand NAND2_1749 ( U4759 , U3034 , U3051 );
nand NAND2_1750 ( U4760 , R1150_U27 , U4016 );
nand NAND2_1751 ( U4761 , R1117_U26 , U4018 );
nand NAND2_1752 ( U4762 , R1138_U114 , U4017 );
nand NAND2_1753 ( U4763 , R1192_U28 , U4014 );
nand NAND2_1754 ( U4764 , R1207_U28 , U4013 );
nand NAND2_1755 ( U4765 , R1171_U114 , U4024 );
nand NAND2_1756 ( U4766 , R1240_U114 , U4022 );
nand NAND3_1757 ( U4767 , U3049 , U5740 , U3838 );
nand NAND2_1758 ( U4768 , R1222_U110 , U3027 );
nand NAND2_1759 ( U4769 , R1282_U44 , U3024 );
nand NAND2_1760 ( U4770 , U4040 , U4021 );
nand NAND3_1761 ( U4771 , U3776 , U3049 , U3775 );
nand NAND2_1762 ( U4772 , REG2_REG_31_ , U3019 );
nand NAND2_1763 ( U4773 , REG1_REG_31_ , U3020 );
nand NAND2_1764 ( U4774 , REG0_REG_31_ , U3021 );
not NOT1_1765 ( U4775 , U3053 );
nand NAND2_1766 ( U4776 , R1282_U42 , U3024 );
nand NAND2_1767 ( U4777 , U4039 , U4021 );
nand NAND3_1768 ( U4778 , U4777 , U4002 , U4776 );
nand NAND2_1769 ( U4779 , R1282_U39 , U3024 );
nand NAND2_1770 ( U4780 , U4038 , U4021 );
nand NAND3_1771 ( U4781 , U4780 , U4002 , U4779 );
nand NAND2_1772 ( U4782 , U5820 , U5817 );
nand NAND2_1773 ( U4783 , U3779 , U3017 );
nand NAND2_1774 ( U4784 , U3418 , U4783 );
nand NAND2_1775 ( U4785 , U3036 , U3075 );
nand NAND2_1776 ( U4786 , U3033 , REG3_REG_0_ );
nand NAND2_1777 ( U4787 , U3032 , R1222_U104 );
nand NAND2_1778 ( U4788 , U3031 , U3464 );
nand NAND2_1779 ( U4789 , U3030 , U3464 );
nand NAND2_1780 ( U4790 , U3036 , U3065 );
nand NAND2_1781 ( U4791 , U3033 , REG3_REG_1_ );
nand NAND2_1782 ( U4792 , U3032 , R1222_U103 );
nand NAND2_1783 ( U4793 , U3031 , U3468 );
nand NAND2_1784 ( U4794 , U3030 , R1282_U31 );
nand NAND2_1785 ( U4795 , U3036 , U3061 );
nand NAND2_1786 ( U4796 , U3033 , REG3_REG_2_ );
nand NAND2_1787 ( U4797 , U3032 , R1222_U23 );
nand NAND2_1788 ( U4798 , U3031 , U3470 );
nand NAND2_1789 ( U4799 , U3030 , R1282_U6 );
nand NAND2_1790 ( U4800 , U3036 , U3057 );
nand NAND2_1791 ( U4801 , U3033 , ADD_95_U4 );
nand NAND2_1792 ( U4802 , U3032 , R1222_U109 );
nand NAND2_1793 ( U4803 , U3031 , U3472 );
nand NAND2_1794 ( U4804 , U3030 , R1282_U7 );
nand NAND2_1795 ( U4805 , U3036 , U3064 );
nand NAND2_1796 ( U4806 , U3033 , ADD_95_U51 );
nand NAND2_1797 ( U4807 , U3032 , R1222_U108 );
nand NAND2_1798 ( U4808 , U3031 , U3474 );
nand NAND2_1799 ( U4809 , U3030 , R1282_U8 );
nand NAND2_1800 ( U4810 , U3036 , U3068 );
nand NAND2_1801 ( U4811 , U3033 , ADD_95_U50 );
nand NAND2_1802 ( U4812 , U3032 , R1222_U24 );
nand NAND2_1803 ( U4813 , U3031 , U3476 );
nand NAND2_1804 ( U4814 , U3030 , R1282_U9 );
nand NAND2_1805 ( U4815 , U3036 , U3067 );
nand NAND2_1806 ( U4816 , U3033 , ADD_95_U49 );
nand NAND2_1807 ( U4817 , U3032 , R1222_U107 );
nand NAND2_1808 ( U4818 , U3031 , U3478 );
nand NAND2_1809 ( U4819 , U3030 , R1282_U10 );
nand NAND2_1810 ( U4820 , U3036 , U3081 );
nand NAND2_1811 ( U4821 , U3033 , ADD_95_U48 );
nand NAND2_1812 ( U4822 , U3032 , R1222_U25 );
nand NAND2_1813 ( U4823 , U3031 , U3480 );
nand NAND2_1814 ( U4824 , U3030 , R1282_U11 );
nand NAND2_1815 ( U4825 , U3036 , U3080 );
nand NAND2_1816 ( U4826 , U3033 , ADD_95_U47 );
nand NAND2_1817 ( U4827 , U3032 , R1222_U106 );
nand NAND2_1818 ( U4828 , U3031 , U3482 );
nand NAND2_1819 ( U4829 , U3030 , R1282_U36 );
nand NAND2_1820 ( U4830 , U3036 , U3059 );
nand NAND2_1821 ( U4831 , U3033 , ADD_95_U46 );
nand NAND2_1822 ( U4832 , U3032 , R1222_U105 );
nand NAND2_1823 ( U4833 , U3031 , U3484 );
nand NAND2_1824 ( U4834 , U3030 , R1282_U33 );
nand NAND2_1825 ( U4835 , U3036 , U3060 );
nand NAND2_1826 ( U4836 , U3033 , ADD_95_U70 );
nand NAND2_1827 ( U4837 , U3032 , R1222_U17 );
nand NAND2_1828 ( U4838 , U3031 , U3486 );
nand NAND2_1829 ( U4839 , U3030 , R1282_U94 );
nand NAND2_1830 ( U4840 , U3036 , U3069 );
nand NAND2_1831 ( U4841 , U3033 , ADD_95_U69 );
nand NAND2_1832 ( U4842 , U3032 , R1222_U123 );
nand NAND2_1833 ( U4843 , U3031 , U3488 );
nand NAND2_1834 ( U4844 , U3030 , R1282_U91 );
nand NAND2_1835 ( U4845 , U3036 , U3077 );
nand NAND2_1836 ( U4846 , U3033 , ADD_95_U68 );
nand NAND2_1837 ( U4847 , U3032 , R1222_U122 );
nand NAND2_1838 ( U4848 , U3031 , U3490 );
nand NAND2_1839 ( U4849 , U3030 , R1282_U89 );
nand NAND2_1840 ( U4850 , U3036 , U3076 );
nand NAND2_1841 ( U4851 , U3033 , ADD_95_U67 );
nand NAND2_1842 ( U4852 , U3032 , R1222_U18 );
nand NAND2_1843 ( U4853 , U3031 , U3492 );
nand NAND2_1844 ( U4854 , U3030 , R1282_U86 );
nand NAND2_1845 ( U4855 , U3036 , U3071 );
nand NAND2_1846 ( U4856 , U3033 , ADD_95_U66 );
nand NAND2_1847 ( U4857 , U3032 , R1222_U121 );
nand NAND2_1848 ( U4858 , U3031 , U3494 );
nand NAND2_1849 ( U4859 , U3030 , R1282_U84 );
nand NAND2_1850 ( U4860 , U3036 , U3070 );
nand NAND2_1851 ( U4861 , U3033 , ADD_95_U65 );
nand NAND2_1852 ( U4862 , U3032 , R1222_U120 );
nand NAND2_1853 ( U4863 , U3031 , U3496 );
nand NAND2_1854 ( U4864 , U3030 , R1282_U81 );
nand NAND2_1855 ( U4865 , U3036 , U3066 );
nand NAND2_1856 ( U4866 , U3033 , ADD_95_U64 );
nand NAND2_1857 ( U4867 , U3032 , R1222_U119 );
nand NAND2_1858 ( U4868 , U3031 , U3498 );
nand NAND2_1859 ( U4869 , U3030 , R1282_U79 );
nand NAND2_1860 ( U4870 , U3036 , U3079 );
nand NAND2_1861 ( U4871 , U3033 , ADD_95_U63 );
nand NAND2_1862 ( U4872 , U3032 , R1222_U19 );
nand NAND2_1863 ( U4873 , U3031 , U3500 );
nand NAND2_1864 ( U4874 , U3030 , R1282_U76 );
nand NAND2_1865 ( U4875 , U3036 , U3078 );
nand NAND2_1866 ( U4876 , U3033 , ADD_95_U62 );
nand NAND2_1867 ( U4877 , U3032 , R1222_U118 );
nand NAND2_1868 ( U4878 , U3031 , U3502 );
nand NAND2_1869 ( U4879 , U3030 , R1282_U74 );
nand NAND2_1870 ( U4880 , U3036 , U3073 );
nand NAND2_1871 ( U4881 , U3033 , ADD_95_U61 );
nand NAND2_1872 ( U4882 , U3032 , R1222_U117 );
nand NAND2_1873 ( U4883 , U3031 , U3504 );
nand NAND2_1874 ( U4884 , U3030 , R1282_U71 );
nand NAND2_1875 ( U4885 , U3036 , U3072 );
nand NAND2_1876 ( U4886 , U3033 , ADD_95_U60 );
nand NAND2_1877 ( U4887 , U3032 , R1222_U20 );
nand NAND2_1878 ( U4888 , U3031 , U4037 );
nand NAND2_1879 ( U4889 , U3030 , R1282_U67 );
nand NAND2_1880 ( U4890 , U3036 , U3058 );
nand NAND2_1881 ( U4891 , U3033 , ADD_95_U59 );
nand NAND2_1882 ( U4892 , U3032 , R1222_U21 );
nand NAND2_1883 ( U4893 , U3031 , U4036 );
nand NAND2_1884 ( U4894 , U3030 , R1282_U64 );
nand NAND2_1885 ( U4895 , U3036 , U3063 );
nand NAND2_1886 ( U4896 , U3033 , ADD_95_U58 );
nand NAND2_1887 ( U4897 , U3032 , R1222_U116 );
nand NAND2_1888 ( U4898 , U3031 , U4035 );
nand NAND2_1889 ( U4899 , U3030 , R1282_U62 );
nand NAND2_1890 ( U4900 , U3036 , U3062 );
nand NAND2_1891 ( U4901 , U3033 , ADD_95_U57 );
nand NAND2_1892 ( U4902 , U3032 , R1222_U115 );
nand NAND2_1893 ( U4903 , U3031 , U4034 );
nand NAND2_1894 ( U4904 , U3030 , R1282_U59 );
nand NAND2_1895 ( U4905 , U3036 , U3055 );
nand NAND2_1896 ( U4906 , U3033 , ADD_95_U56 );
nand NAND2_1897 ( U4907 , U3032 , R1222_U114 );
nand NAND2_1898 ( U4908 , U3031 , U4033 );
nand NAND2_1899 ( U4909 , U3030 , R1282_U57 );
nand NAND2_1900 ( U4910 , U3036 , U3054 );
nand NAND2_1901 ( U4911 , U3033 , ADD_95_U55 );
nand NAND2_1902 ( U4912 , U3032 , R1222_U113 );
nand NAND2_1903 ( U4913 , U3031 , U4032 );
nand NAND2_1904 ( U4914 , U3030 , R1282_U54 );
nand NAND2_1905 ( U4915 , U3036 , U3050 );
nand NAND2_1906 ( U4916 , U3033 , ADD_95_U54 );
nand NAND2_1907 ( U4917 , U3032 , R1222_U22 );
nand NAND2_1908 ( U4918 , U3031 , U4031 );
nand NAND2_1909 ( U4919 , U3030 , R1282_U52 );
nand NAND2_1910 ( U4920 , U3036 , U3051 );
nand NAND2_1911 ( U4921 , U3033 , ADD_95_U53 );
nand NAND2_1912 ( U4922 , U3032 , R1222_U112 );
nand NAND2_1913 ( U4923 , U3031 , U4030 );
nand NAND2_1914 ( U4924 , U3030 , R1282_U49 );
nand NAND2_1915 ( U4925 , U3036 , U3052 );
nand NAND2_1916 ( U4926 , U3033 , ADD_95_U52 );
nand NAND2_1917 ( U4927 , U3032 , R1222_U111 );
nand NAND2_1918 ( U4928 , U3031 , U4029 );
nand NAND2_1919 ( U4929 , U3030 , R1282_U47 );
nand NAND2_1920 ( U4930 , U3033 , ADD_95_U5 );
nand NAND2_1921 ( U4931 , U3032 , R1222_U110 );
nand NAND2_1922 ( U4932 , U3031 , U4040 );
nand NAND2_1923 ( U4933 , U3030 , R1282_U44 );
nand NAND2_1924 ( U4934 , U3031 , U4039 );
nand NAND2_1925 ( U4935 , U3030 , R1282_U42 );
nand NAND2_1926 ( U4936 , U3031 , U4038 );
nand NAND2_1927 ( U4937 , U3030 , R1282_U39 );
nand NAND4_1928 ( U4938 , U3843 , U3842 , U3840 , U3839 );
nand NAND3_1929 ( U4939 , U3042 , U3044 , R1105_U4 );
nand NAND2_1930 ( U4940 , U3844 , U3044 );
nand NAND3_1931 ( U4941 , U3038 , U3044 , R1162_U4 );
not NOT1_1932 ( U4942 , U3421 );
nand NAND2_1933 ( U4943 , U3043 , R1105_U4 );
nand NAND2_1934 ( U4944 , REG3_REG_19_ , U3149 );
nand NAND2_1935 ( U4945 , U3041 , U3461 );
nand NAND2_1936 ( U4946 , U3039 , R1162_U4 );
nand NAND2_1937 ( U4947 , ADDR_REG_19_ , U4942 );
nand NAND3_1938 ( U4948 , U3042 , U3044 , R1105_U55 );
nand NAND2_1939 ( U4949 , U3849 , U3044 );
nand NAND3_1940 ( U4950 , U3038 , U3044 , R1162_U62 );
nand NAND2_1941 ( U4951 , R1105_U55 , U3043 );
nand NAND2_1942 ( U4952 , REG3_REG_18_ , U3149 );
nand NAND2_1943 ( U4953 , U3041 , U3444 );
nand NAND2_1944 ( U4954 , R1162_U62 , U3039 );
nand NAND2_1945 ( U4955 , ADDR_REG_18_ , U4942 );
nand NAND2_1946 ( U4956 , R1105_U56 , U3042 );
nand NAND2_1947 ( U4957 , U3040 , U3445 );
nand NAND2_1948 ( U4958 , R1162_U63 , U3038 );
nand NAND3_1949 ( U4959 , U4957 , U4956 , U4958 );
nand NAND2_1950 ( U4960 , U3044 , U4959 );
nand NAND2_1951 ( U4961 , R1105_U56 , U3043 );
nand NAND2_1952 ( U4962 , REG3_REG_17_ , U3149 );
nand NAND2_1953 ( U4963 , U3041 , U3445 );
nand NAND2_1954 ( U4964 , R1162_U63 , U3039 );
nand NAND2_1955 ( U4965 , ADDR_REG_17_ , U4942 );
nand NAND2_1956 ( U4966 , R1105_U57 , U3042 );
nand NAND2_1957 ( U4967 , U3040 , U3446 );
nand NAND2_1958 ( U4968 , R1162_U64 , U3038 );
nand NAND3_1959 ( U4969 , U4967 , U4966 , U4968 );
nand NAND2_1960 ( U4970 , U3044 , U4969 );
nand NAND2_1961 ( U4971 , R1105_U57 , U3043 );
nand NAND2_1962 ( U4972 , REG3_REG_16_ , U3149 );
nand NAND2_1963 ( U4973 , U3041 , U3446 );
nand NAND2_1964 ( U4974 , R1162_U64 , U3039 );
nand NAND2_1965 ( U4975 , ADDR_REG_16_ , U4942 );
nand NAND2_1966 ( U4976 , R1105_U58 , U3042 );
nand NAND2_1967 ( U4977 , U3040 , U3447 );
nand NAND2_1968 ( U4978 , R1162_U65 , U3038 );
nand NAND3_1969 ( U4979 , U4977 , U4976 , U4978 );
nand NAND2_1970 ( U4980 , U3044 , U4979 );
nand NAND2_1971 ( U4981 , R1105_U58 , U3043 );
nand NAND2_1972 ( U4982 , REG3_REG_15_ , U3149 );
nand NAND2_1973 ( U4983 , U3041 , U3447 );
nand NAND2_1974 ( U4984 , R1162_U65 , U3039 );
nand NAND2_1975 ( U4985 , ADDR_REG_15_ , U4942 );
nand NAND2_1976 ( U4986 , R1105_U59 , U3042 );
nand NAND2_1977 ( U4987 , U3040 , U3448 );
nand NAND2_1978 ( U4988 , R1162_U66 , U3038 );
nand NAND3_1979 ( U4989 , U4987 , U4986 , U4988 );
nand NAND2_1980 ( U4990 , U3044 , U4989 );
nand NAND2_1981 ( U4991 , R1105_U59 , U3043 );
nand NAND2_1982 ( U4992 , REG3_REG_14_ , U3149 );
nand NAND2_1983 ( U4993 , U3041 , U3448 );
nand NAND2_1984 ( U4994 , R1162_U66 , U3039 );
nand NAND2_1985 ( U4995 , ADDR_REG_14_ , U4942 );
nand NAND2_1986 ( U4996 , R1105_U60 , U3042 );
nand NAND2_1987 ( U4997 , U3040 , U3449 );
nand NAND2_1988 ( U4998 , R1162_U67 , U3038 );
nand NAND3_1989 ( U4999 , U4997 , U4996 , U4998 );
nand NAND2_1990 ( U5000 , U3044 , U4999 );
nand NAND2_1991 ( U5001 , R1105_U60 , U3043 );
nand NAND2_1992 ( U5002 , REG3_REG_13_ , U3149 );
nand NAND2_1993 ( U5003 , U3041 , U3449 );
nand NAND2_1994 ( U5004 , R1162_U67 , U3039 );
nand NAND2_1995 ( U5005 , ADDR_REG_13_ , U4942 );
nand NAND2_1996 ( U5006 , R1105_U61 , U3042 );
nand NAND2_1997 ( U5007 , U3040 , U3450 );
nand NAND2_1998 ( U5008 , R1162_U68 , U3038 );
nand NAND3_1999 ( U5009 , U5007 , U5006 , U5008 );
nand NAND2_2000 ( U5010 , U3044 , U5009 );
nand NAND2_2001 ( U5011 , R1105_U61 , U3043 );
nand NAND2_2002 ( U5012 , REG3_REG_12_ , U3149 );
nand NAND2_2003 ( U5013 , U3041 , U3450 );
nand NAND2_2004 ( U5014 , R1162_U68 , U3039 );
nand NAND2_2005 ( U5015 , ADDR_REG_12_ , U4942 );
nand NAND2_2006 ( U5016 , R1105_U62 , U3042 );
nand NAND2_2007 ( U5017 , U3040 , U3451 );
nand NAND2_2008 ( U5018 , R1162_U69 , U3038 );
nand NAND3_2009 ( U5019 , U5017 , U5016 , U5018 );
nand NAND2_2010 ( U5020 , U3044 , U5019 );
nand NAND2_2011 ( U5021 , R1105_U62 , U3043 );
nand NAND2_2012 ( U5022 , REG3_REG_11_ , U3149 );
nand NAND2_2013 ( U5023 , U3041 , U3451 );
nand NAND2_2014 ( U5024 , R1162_U69 , U3039 );
nand NAND2_2015 ( U5025 , ADDR_REG_11_ , U4942 );
nand NAND2_2016 ( U5026 , R1105_U63 , U3042 );
nand NAND2_2017 ( U5027 , U3040 , U3452 );
nand NAND2_2018 ( U5028 , R1162_U70 , U3038 );
nand NAND3_2019 ( U5029 , U5027 , U5026 , U5028 );
nand NAND2_2020 ( U5030 , U3044 , U5029 );
nand NAND2_2021 ( U5031 , R1105_U63 , U3043 );
nand NAND2_2022 ( U5032 , REG3_REG_10_ , U3149 );
nand NAND2_2023 ( U5033 , U3041 , U3452 );
nand NAND2_2024 ( U5034 , R1162_U70 , U3039 );
nand NAND2_2025 ( U5035 , ADDR_REG_10_ , U4942 );
nand NAND2_2026 ( U5036 , R1105_U47 , U3042 );
nand NAND2_2027 ( U5037 , U3040 , U3435 );
nand NAND2_2028 ( U5038 , R1162_U54 , U3038 );
nand NAND3_2029 ( U5039 , U5037 , U5036 , U5038 );
nand NAND2_2030 ( U5040 , U3044 , U5039 );
nand NAND2_2031 ( U5041 , R1105_U47 , U3043 );
nand NAND2_2032 ( U5042 , REG3_REG_9_ , U3149 );
nand NAND2_2033 ( U5043 , U3041 , U3435 );
nand NAND2_2034 ( U5044 , R1162_U54 , U3039 );
nand NAND2_2035 ( U5045 , ADDR_REG_9_ , U4942 );
nand NAND2_2036 ( U5046 , R1105_U48 , U3042 );
nand NAND2_2037 ( U5047 , U3040 , U3436 );
nand NAND2_2038 ( U5048 , R1162_U55 , U3038 );
nand NAND3_2039 ( U5049 , U5047 , U5046 , U5048 );
nand NAND2_2040 ( U5050 , U3044 , U5049 );
nand NAND2_2041 ( U5051 , R1105_U48 , U3043 );
nand NAND2_2042 ( U5052 , REG3_REG_8_ , U3149 );
nand NAND2_2043 ( U5053 , U3041 , U3436 );
nand NAND2_2044 ( U5054 , R1162_U55 , U3039 );
nand NAND2_2045 ( U5055 , ADDR_REG_8_ , U4942 );
nand NAND2_2046 ( U5056 , R1105_U49 , U3042 );
nand NAND2_2047 ( U5057 , U3040 , U3437 );
nand NAND2_2048 ( U5058 , R1162_U56 , U3038 );
nand NAND3_2049 ( U5059 , U5057 , U5056 , U5058 );
nand NAND2_2050 ( U5060 , U3044 , U5059 );
nand NAND2_2051 ( U5061 , R1105_U49 , U3043 );
nand NAND2_2052 ( U5062 , REG3_REG_7_ , U3149 );
nand NAND2_2053 ( U5063 , U3041 , U3437 );
nand NAND2_2054 ( U5064 , R1162_U56 , U3039 );
nand NAND2_2055 ( U5065 , ADDR_REG_7_ , U4942 );
nand NAND2_2056 ( U5066 , R1105_U50 , U3042 );
nand NAND2_2057 ( U5067 , U3040 , U3438 );
nand NAND2_2058 ( U5068 , R1162_U57 , U3038 );
nand NAND3_2059 ( U5069 , U5067 , U5066 , U5068 );
nand NAND2_2060 ( U5070 , U3044 , U5069 );
nand NAND2_2061 ( U5071 , R1105_U50 , U3043 );
nand NAND2_2062 ( U5072 , REG3_REG_6_ , U3149 );
nand NAND2_2063 ( U5073 , U3041 , U3438 );
nand NAND2_2064 ( U5074 , R1162_U57 , U3039 );
nand NAND2_2065 ( U5075 , ADDR_REG_6_ , U4942 );
nand NAND2_2066 ( U5076 , R1105_U51 , U3042 );
nand NAND2_2067 ( U5077 , U3040 , U3439 );
nand NAND2_2068 ( U5078 , R1162_U58 , U3038 );
nand NAND3_2069 ( U5079 , U5077 , U5076 , U5078 );
nand NAND2_2070 ( U5080 , U3044 , U5079 );
nand NAND2_2071 ( U5081 , R1105_U51 , U3043 );
nand NAND2_2072 ( U5082 , REG3_REG_5_ , U3149 );
nand NAND2_2073 ( U5083 , U3041 , U3439 );
nand NAND2_2074 ( U5084 , R1162_U58 , U3039 );
nand NAND2_2075 ( U5085 , ADDR_REG_5_ , U4942 );
nand NAND2_2076 ( U5086 , R1105_U52 , U3042 );
nand NAND2_2077 ( U5087 , U3040 , U3440 );
nand NAND2_2078 ( U5088 , R1162_U59 , U3038 );
nand NAND3_2079 ( U5089 , U5087 , U5086 , U5088 );
nand NAND2_2080 ( U5090 , U3044 , U5089 );
nand NAND2_2081 ( U5091 , R1105_U52 , U3043 );
nand NAND2_2082 ( U5092 , REG3_REG_4_ , U3149 );
nand NAND2_2083 ( U5093 , U3041 , U3440 );
nand NAND2_2084 ( U5094 , R1162_U59 , U3039 );
nand NAND2_2085 ( U5095 , ADDR_REG_4_ , U4942 );
nand NAND2_2086 ( U5096 , R1105_U53 , U3042 );
nand NAND2_2087 ( U5097 , U3040 , U3441 );
nand NAND2_2088 ( U5098 , R1162_U60 , U3038 );
nand NAND3_2089 ( U5099 , U5097 , U5096 , U5098 );
nand NAND2_2090 ( U5100 , U3044 , U5099 );
nand NAND2_2091 ( U5101 , R1105_U53 , U3043 );
nand NAND2_2092 ( U5102 , REG3_REG_3_ , U3149 );
nand NAND2_2093 ( U5103 , U3041 , U3441 );
nand NAND2_2094 ( U5104 , R1162_U60 , U3039 );
nand NAND2_2095 ( U5105 , ADDR_REG_3_ , U4942 );
nand NAND2_2096 ( U5106 , R1105_U54 , U3042 );
nand NAND2_2097 ( U5107 , U3040 , U3442 );
nand NAND2_2098 ( U5108 , R1162_U61 , U3038 );
nand NAND3_2099 ( U5109 , U5107 , U5106 , U5108 );
nand NAND2_2100 ( U5110 , U3044 , U5109 );
nand NAND2_2101 ( U5111 , R1105_U54 , U3043 );
nand NAND2_2102 ( U5112 , REG3_REG_2_ , U3149 );
nand NAND2_2103 ( U5113 , U3041 , U3442 );
nand NAND2_2104 ( U5114 , R1162_U61 , U3039 );
nand NAND2_2105 ( U5115 , ADDR_REG_2_ , U4942 );
nand NAND2_2106 ( U5116 , R1105_U5 , U3042 );
nand NAND2_2107 ( U5117 , U3040 , U3443 );
nand NAND2_2108 ( U5118 , R1162_U5 , U3038 );
nand NAND3_2109 ( U5119 , U5117 , U5116 , U5118 );
nand NAND2_2110 ( U5120 , U3044 , U5119 );
nand NAND2_2111 ( U5121 , R1105_U5 , U3043 );
nand NAND2_2112 ( U5122 , REG3_REG_1_ , U3149 );
nand NAND2_2113 ( U5123 , U3041 , U3443 );
nand NAND2_2114 ( U5124 , R1162_U5 , U3039 );
nand NAND2_2115 ( U5125 , ADDR_REG_1_ , U4942 );
nand NAND2_2116 ( U5126 , R1105_U46 , U3042 );
nand NAND2_2117 ( U5127 , U3040 , U3453 );
nand NAND2_2118 ( U5128 , R1162_U53 , U3038 );
nand NAND3_2119 ( U5129 , U5127 , U5126 , U5128 );
nand NAND2_2120 ( U5130 , U3044 , U5129 );
nand NAND2_2121 ( U5131 , R1105_U46 , U3043 );
nand NAND2_2122 ( U5132 , REG3_REG_0_ , U3149 );
nand NAND2_2123 ( U5133 , U3041 , U3453 );
nand NAND2_2124 ( U5134 , R1162_U53 , U3039 );
nand NAND2_2125 ( U5135 , ADDR_REG_0_ , U4942 );
nand NAND3_2126 ( U5136 , U6257 , U6256 , U3903 );
not NOT1_2127 ( U5137 , U3425 );
nand NAND2_2128 ( U5138 , U5137 , U4055 );
nand NAND2_2129 ( U5139 , U4006 , U5138 );
nand NAND2_2130 ( U5140 , U4020 , U3424 );
nand NAND2_2131 ( U5141 , U4012 , U4005 );
nand NAND3_2132 ( U5142 , U6253 , U6252 , U3902 );
nand NAND3_2133 ( U5143 , U3461 , U3014 , U4005 );
nand NAND2_2134 ( U5144 , U3431 , U5142 );
nand NAND2_2135 ( U5145 , U5144 , U5143 );
nand NAND3_2136 ( U5146 , U4041 , U3023 , R395_U6 );
nand NAND2_2137 ( U5147 , U5145 , STATE_REG );
nand NAND2_2138 ( U5148 , B_REG , U5136 );
nand NAND2_2139 ( U5149 , U3037 , U3076 );
nand NAND2_2140 ( U5150 , U3035 , U3070 );
nand NAND2_2141 ( U5151 , ADD_95_U65 , U3427 );
nand NAND3_2142 ( U5152 , U5150 , U5149 , U5151 );
nand NAND3_2143 ( U5153 , U3364 , U3363 , U3362 );
nand NAND2_2144 ( U5154 , U3419 , U3366 );
nand NAND2_2145 ( U5155 , U5805 , U5154 );
nand NAND2_2146 ( U5156 , U5808 , U5153 );
nand NAND4_2147 ( U5157 , U5156 , U3369 , U5155 , U3906 );
nand NAND2_2148 ( U5158 , U5157 , U3427 );
not NOT1_2149 ( U5159 , U3429 );
nand NAND2_2150 ( U5160 , U3496 , U5744 );
nand NAND2_2151 ( U5161 , ADD_95_U65 , U5743 );
nand NAND2_2152 ( U5162 , U4049 , U5152 );
nand NAND2_2153 ( U5163 , R1165_U109 , U3028 );
nand NAND2_2154 ( U5164 , REG3_REG_15_ , U3149 );
nand NAND2_2155 ( U5165 , U3037 , U3055 );
nand NAND2_2156 ( U5166 , U3035 , U3050 );
nand NAND2_2157 ( U5167 , ADD_95_U54 , U3427 );
nand NAND3_2158 ( U5168 , U5166 , U5165 , U5167 );
nand NAND2_2159 ( U5169 , U4021 , U3427 );
nand NAND2_2160 ( U5170 , U5159 , U5169 );
nand NAND2_2161 ( U5171 , U4028 , U4021 );
nand NAND2_2162 ( U5172 , U3418 , U5171 );
nand NAND2_2163 ( U5173 , U3046 , U4031 );
nand NAND2_2164 ( U5174 , U3045 , ADD_95_U54 );
nand NAND2_2165 ( U5175 , U4049 , U5168 );
nand NAND2_2166 ( U5176 , R1165_U15 , U3028 );
nand NAND2_2167 ( U5177 , REG3_REG_26_ , U3149 );
nand NAND2_2168 ( U5178 , U3037 , U3064 );
nand NAND2_2169 ( U5179 , U3035 , U3067 );
nand NAND2_2170 ( U5180 , ADD_95_U49 , U3427 );
nand NAND3_2171 ( U5181 , U5179 , U5178 , U5180 );
nand NAND2_2172 ( U5182 , U3478 , U5744 );
nand NAND2_2173 ( U5183 , ADD_95_U49 , U5743 );
nand NAND2_2174 ( U5184 , U4049 , U5181 );
nand NAND2_2175 ( U5185 , R1165_U94 , U3028 );
nand NAND2_2176 ( U5186 , REG3_REG_6_ , U3149 );
nand NAND2_2177 ( U5187 , U3037 , U3066 );
nand NAND2_2178 ( U5188 , U3035 , U3078 );
nand NAND2_2179 ( U5189 , ADD_95_U62 , U3427 );
nand NAND3_2180 ( U5190 , U5188 , U5187 , U5189 );
nand NAND2_2181 ( U5191 , U3502 , U5744 );
nand NAND2_2182 ( U5192 , ADD_95_U62 , U5743 );
nand NAND2_2183 ( U5193 , U4049 , U5190 );
nand NAND2_2184 ( U5194 , R1165_U107 , U3028 );
nand NAND2_2185 ( U5195 , REG3_REG_18_ , U3149 );
nand NAND2_2186 ( U5196 , U3037 , U3075 );
nand NAND2_2187 ( U5197 , U3035 , U3061 );
nand NAND2_2188 ( U5198 , REG3_REG_2_ , U3427 );
nand NAND3_2189 ( U5199 , U5197 , U5196 , U5198 );
nand NAND2_2190 ( U5200 , U3470 , U5744 );
nand NAND2_2191 ( U5201 , REG3_REG_2_ , U5743 );
nand NAND2_2192 ( U5202 , U4049 , U5199 );
nand NAND2_2193 ( U5203 , R1165_U97 , U3028 );
nand NAND2_2194 ( U5204 , REG3_REG_2_ , U3149 );
nand NAND2_2195 ( U5205 , U3037 , U3059 );
nand NAND2_2196 ( U5206 , U3035 , U3069 );
nand NAND2_2197 ( U5207 , ADD_95_U69 , U3427 );
nand NAND3_2198 ( U5208 , U5206 , U5205 , U5207 );
nand NAND2_2199 ( U5209 , U3488 , U5744 );
nand NAND2_2200 ( U5210 , ADD_95_U69 , U5743 );
nand NAND2_2201 ( U5211 , U4049 , U5208 );
nand NAND2_2202 ( U5212 , R1165_U112 , U3028 );
nand NAND2_2203 ( U5213 , REG3_REG_11_ , U3149 );
nand NAND2_2204 ( U5214 , U3037 , U3072 );
nand NAND2_2205 ( U5215 , U3035 , U3063 );
nand NAND2_2206 ( U5216 , ADD_95_U58 , U3427 );
nand NAND3_2207 ( U5217 , U5215 , U5214 , U5216 );
nand NAND2_2208 ( U5218 , U3046 , U4035 );
nand NAND2_2209 ( U5219 , U3045 , ADD_95_U58 );
nand NAND2_2210 ( U5220 , U4049 , U5217 );
nand NAND2_2211 ( U5221 , R1165_U103 , U3028 );
nand NAND2_2212 ( U5222 , REG3_REG_22_ , U3149 );
nand NAND2_2213 ( U5223 , U3037 , U3069 );
nand NAND2_2214 ( U5224 , U3035 , U3076 );
nand NAND2_2215 ( U5225 , ADD_95_U67 , U3427 );
nand NAND3_2216 ( U5226 , U5224 , U5223 , U5225 );
nand NAND2_2217 ( U5227 , U3492 , U5744 );
nand NAND2_2218 ( U5228 , ADD_95_U67 , U5743 );
nand NAND2_2219 ( U5229 , U4049 , U5226 );
nand NAND2_2220 ( U5230 , R1165_U12 , U3028 );
nand NAND2_2221 ( U5231 , REG3_REG_13_ , U3149 );
nand NAND2_2222 ( U5232 , U3037 , U3078 );
nand NAND2_2223 ( U5233 , U3035 , U3072 );
nand NAND2_2224 ( U5234 , ADD_95_U60 , U3427 );
nand NAND3_2225 ( U5235 , U5233 , U5232 , U5234 );
nand NAND2_2226 ( U5236 , U3046 , U4037 );
nand NAND2_2227 ( U5237 , U3045 , ADD_95_U60 );
nand NAND2_2228 ( U5238 , U4049 , U5235 );
nand NAND2_2229 ( U5239 , R1165_U104 , U3028 );
nand NAND2_2230 ( U5240 , REG3_REG_20_ , U3149 );
nand NAND2_2231 ( U5241 , U3428 , U3426 );
nand NAND2_2232 ( U5242 , U5241 , U3427 );
nand NAND2_2233 ( U5243 , U4050 , U5242 );
nand NAND2_2234 ( U5244 , U3911 , U3035 );
nand NAND2_2235 ( U5245 , U3464 , U5744 );
nand NAND2_2236 ( U5246 , REG3_REG_0_ , U5243 );
nand NAND2_2237 ( U5247 , R1165_U91 , U3028 );
nand NAND2_2238 ( U5248 , REG3_REG_0_ , U3149 );
nand NAND2_2239 ( U5249 , U3037 , U3081 );
nand NAND2_2240 ( U5250 , U3035 , U3059 );
nand NAND2_2241 ( U5251 , ADD_95_U46 , U3427 );
nand NAND3_2242 ( U5252 , U5250 , U5249 , U5251 );
nand NAND2_2243 ( U5253 , U3484 , U5744 );
nand NAND2_2244 ( U5254 , ADD_95_U46 , U5743 );
nand NAND2_2245 ( U5255 , U4049 , U5252 );
nand NAND2_2246 ( U5256 , R1165_U92 , U3028 );
nand NAND2_2247 ( U5257 , REG3_REG_9_ , U3149 );
nand NAND2_2248 ( U5258 , U3037 , U3061 );
nand NAND2_2249 ( U5259 , U3035 , U3064 );
nand NAND2_2250 ( U5260 , ADD_95_U51 , U3427 );
nand NAND3_2251 ( U5261 , U5259 , U5258 , U5260 );
nand NAND2_2252 ( U5262 , U3474 , U5744 );
nand NAND2_2253 ( U5263 , ADD_95_U51 , U5743 );
nand NAND2_2254 ( U5264 , U4049 , U5261 );
nand NAND2_2255 ( U5265 , R1165_U96 , U3028 );
nand NAND2_2256 ( U5266 , REG3_REG_4_ , U3149 );
nand NAND2_2257 ( U5267 , U3037 , U3063 );
nand NAND2_2258 ( U5268 , U3035 , U3055 );
nand NAND2_2259 ( U5269 , ADD_95_U56 , U3427 );
nand NAND3_2260 ( U5270 , U5268 , U5267 , U5269 );
nand NAND2_2261 ( U5271 , U3046 , U4033 );
nand NAND2_2262 ( U5272 , U3045 , ADD_95_U56 );
nand NAND2_2263 ( U5273 , U4049 , U5270 );
nand NAND2_2264 ( U5274 , R1165_U101 , U3028 );
nand NAND2_2265 ( U5275 , REG3_REG_24_ , U3149 );
nand NAND2_2266 ( U5276 , U3037 , U3070 );
nand NAND2_2267 ( U5277 , U3035 , U3079 );
nand NAND2_2268 ( U5278 , ADD_95_U63 , U3427 );
nand NAND3_2269 ( U5279 , U5277 , U5276 , U5278 );
nand NAND2_2270 ( U5280 , U3500 , U5744 );
nand NAND2_2271 ( U5281 , ADD_95_U63 , U5743 );
nand NAND2_2272 ( U5282 , U4049 , U5279 );
nand NAND2_2273 ( U5283 , R1165_U13 , U3028 );
nand NAND2_2274 ( U5284 , REG3_REG_17_ , U3149 );
nand NAND2_2275 ( U5285 , U3037 , U3057 );
nand NAND2_2276 ( U5286 , U3035 , U3068 );
nand NAND2_2277 ( U5287 , ADD_95_U50 , U3427 );
nand NAND3_2278 ( U5288 , U5286 , U5285 , U5287 );
nand NAND2_2279 ( U5289 , U3476 , U5744 );
nand NAND2_2280 ( U5290 , ADD_95_U50 , U5743 );
nand NAND2_2281 ( U5291 , U4049 , U5288 );
nand NAND2_2282 ( U5292 , R1165_U95 , U3028 );
nand NAND2_2283 ( U5293 , REG3_REG_5_ , U3149 );
nand NAND2_2284 ( U5294 , U3037 , U3071 );
nand NAND2_2285 ( U5295 , U3035 , U3066 );
nand NAND2_2286 ( U5296 , ADD_95_U64 , U3427 );
nand NAND3_2287 ( U5297 , U5295 , U5294 , U5296 );
nand NAND2_2288 ( U5298 , U3498 , U5744 );
nand NAND2_2289 ( U5299 , ADD_95_U64 , U5743 );
nand NAND2_2290 ( U5300 , U4049 , U5297 );
nand NAND2_2291 ( U5301 , R1165_U108 , U3028 );
nand NAND2_2292 ( U5302 , REG3_REG_16_ , U3149 );
nand NAND2_2293 ( U5303 , U3037 , U3062 );
nand NAND2_2294 ( U5304 , U3035 , U3054 );
nand NAND2_2295 ( U5305 , ADD_95_U55 , U3427 );
nand NAND3_2296 ( U5306 , U5304 , U5303 , U5305 );
nand NAND2_2297 ( U5307 , U3046 , U4032 );
nand NAND2_2298 ( U5308 , U3045 , ADD_95_U55 );
nand NAND2_2299 ( U5309 , U4049 , U5306 );
nand NAND2_2300 ( U5310 , R1165_U100 , U3028 );
nand NAND2_2301 ( U5311 , REG3_REG_25_ , U3149 );
nand NAND2_2302 ( U5312 , U3037 , U3060 );
nand NAND2_2303 ( U5313 , U3035 , U3077 );
nand NAND2_2304 ( U5314 , ADD_95_U68 , U3427 );
nand NAND3_2305 ( U5315 , U5313 , U5312 , U5314 );
nand NAND2_2306 ( U5316 , U3490 , U5744 );
nand NAND2_2307 ( U5317 , ADD_95_U68 , U5743 );
nand NAND2_2308 ( U5318 , U4049 , U5315 );
nand NAND2_2309 ( U5319 , R1165_U111 , U3028 );
nand NAND2_2310 ( U5320 , REG3_REG_12_ , U3149 );
nand NAND2_2311 ( U5321 , U3037 , U3073 );
nand NAND2_2312 ( U5322 , U3035 , U3058 );
nand NAND2_2313 ( U5323 , ADD_95_U59 , U3427 );
nand NAND3_2314 ( U5324 , U5322 , U5321 , U5323 );
nand NAND2_2315 ( U5325 , U3046 , U4036 );
nand NAND2_2316 ( U5326 , U3045 , ADD_95_U59 );
nand NAND2_2317 ( U5327 , U4049 , U5324 );
nand NAND2_2318 ( U5328 , R1165_U14 , U3028 );
nand NAND2_2319 ( U5329 , REG3_REG_21_ , U3149 );
nand NAND2_2320 ( U5330 , U3037 , U3074 );
nand NAND2_2321 ( U5331 , U3035 , U3065 );
nand NAND2_2322 ( U5332 , REG3_REG_1_ , U3427 );
nand NAND3_2323 ( U5333 , U5331 , U5330 , U5332 );
nand NAND2_2324 ( U5334 , U3468 , U5744 );
nand NAND2_2325 ( U5335 , REG3_REG_1_ , U5743 );
nand NAND2_2326 ( U5336 , U4049 , U5333 );
nand NAND2_2327 ( U5337 , R1165_U105 , U3028 );
nand NAND2_2328 ( U5338 , REG3_REG_1_ , U3149 );
nand NAND2_2329 ( U5339 , U3037 , U3067 );
nand NAND2_2330 ( U5340 , U3035 , U3080 );
nand NAND2_2331 ( U5341 , ADD_95_U47 , U3427 );
nand NAND3_2332 ( U5342 , U5340 , U5339 , U5341 );
nand NAND2_2333 ( U5343 , U3482 , U5744 );
nand NAND2_2334 ( U5344 , ADD_95_U47 , U5743 );
nand NAND2_2335 ( U5345 , U4049 , U5342 );
nand NAND2_2336 ( U5346 , R1165_U93 , U3028 );
nand NAND2_2337 ( U5347 , REG3_REG_8_ , U3149 );
nand NAND2_2338 ( U5348 , U3037 , U3050 );
nand NAND2_2339 ( U5349 , U3035 , U3052 );
nand NAND2_2340 ( U5350 , ADD_95_U52 , U3427 );
nand NAND3_2341 ( U5351 , U5349 , U5348 , U5350 );
nand NAND2_2342 ( U5352 , U3046 , U4029 );
nand NAND2_2343 ( U5353 , U3045 , ADD_95_U52 );
nand NAND2_2344 ( U5354 , U4049 , U5351 );
nand NAND2_2345 ( U5355 , R1165_U98 , U3028 );
nand NAND2_2346 ( U5356 , REG3_REG_28_ , U3149 );
nand NAND2_2347 ( U5357 , U3037 , U3079 );
nand NAND2_2348 ( U5358 , U3035 , U3073 );
nand NAND2_2349 ( U5359 , ADD_95_U61 , U3427 );
nand NAND3_2350 ( U5360 , U5358 , U5357 , U5359 );
nand NAND2_2351 ( U5361 , U3504 , U5744 );
nand NAND2_2352 ( U5362 , ADD_95_U61 , U5743 );
nand NAND2_2353 ( U5363 , U4049 , U5360 );
nand NAND2_2354 ( U5364 , R1165_U106 , U3028 );
nand NAND2_2355 ( U5365 , REG3_REG_19_ , U3149 );
nand NAND2_2356 ( U5366 , U3037 , U3065 );
nand NAND2_2357 ( U5367 , U3035 , U3057 );
nand NAND2_2358 ( U5368 , ADD_95_U4 , U3427 );
nand NAND3_2359 ( U5369 , U5367 , U5366 , U5368 );
nand NAND2_2360 ( U5370 , U3472 , U5744 );
nand NAND2_2361 ( U5371 , ADD_95_U4 , U5743 );
nand NAND2_2362 ( U5372 , U4049 , U5369 );
nand NAND2_2363 ( U5373 , R1165_U16 , U3028 );
nand NAND2_2364 ( U5374 , REG3_REG_3_ , U3149 );
nand NAND2_2365 ( U5375 , U3037 , U3080 );
nand NAND2_2366 ( U5376 , U3035 , U3060 );
nand NAND2_2367 ( U5377 , ADD_95_U70 , U3427 );
nand NAND3_2368 ( U5378 , U5376 , U5375 , U5377 );
nand NAND2_2369 ( U5379 , U3486 , U5744 );
nand NAND2_2370 ( U5380 , ADD_95_U70 , U5743 );
nand NAND2_2371 ( U5381 , U4049 , U5378 );
nand NAND2_2372 ( U5382 , R1165_U113 , U3028 );
nand NAND2_2373 ( U5383 , REG3_REG_10_ , U3149 );
nand NAND2_2374 ( U5384 , U3037 , U3058 );
nand NAND2_2375 ( U5385 , U3035 , U3062 );
nand NAND2_2376 ( U5386 , ADD_95_U57 , U3427 );
nand NAND3_2377 ( U5387 , U5385 , U5384 , U5386 );
nand NAND2_2378 ( U5388 , U3046 , U4034 );
nand NAND2_2379 ( U5389 , U3045 , ADD_95_U57 );
nand NAND2_2380 ( U5390 , U4049 , U5387 );
nand NAND2_2381 ( U5391 , R1165_U102 , U3028 );
nand NAND2_2382 ( U5392 , REG3_REG_23_ , U3149 );
nand NAND2_2383 ( U5393 , U3037 , U3077 );
nand NAND2_2384 ( U5394 , U3035 , U3071 );
nand NAND2_2385 ( U5395 , ADD_95_U66 , U3427 );
nand NAND3_2386 ( U5396 , U5394 , U5393 , U5395 );
nand NAND2_2387 ( U5397 , U3494 , U5744 );
nand NAND2_2388 ( U5398 , ADD_95_U66 , U5743 );
nand NAND2_2389 ( U5399 , U4049 , U5396 );
nand NAND2_2390 ( U5400 , R1165_U110 , U3028 );
nand NAND2_2391 ( U5401 , REG3_REG_14_ , U3149 );
nand NAND2_2392 ( U5402 , U3037 , U3054 );
nand NAND2_2393 ( U5403 , U3035 , U3051 );
nand NAND2_2394 ( U5404 , ADD_95_U53 , U3427 );
nand NAND3_2395 ( U5405 , U5403 , U5402 , U5404 );
nand NAND2_2396 ( U5406 , U3046 , U4030 );
nand NAND2_2397 ( U5407 , U3045 , ADD_95_U53 );
nand NAND2_2398 ( U5408 , U4049 , U5405 );
nand NAND2_2399 ( U5409 , R1165_U99 , U3028 );
nand NAND2_2400 ( U5410 , REG3_REG_27_ , U3149 );
nand NAND2_2401 ( U5411 , U3037 , U3068 );
nand NAND2_2402 ( U5412 , U3035 , U3081 );
nand NAND2_2403 ( U5413 , ADD_95_U48 , U3427 );
nand NAND3_2404 ( U5414 , U5412 , U5411 , U5413 );
nand NAND2_2405 ( U5415 , U3480 , U5744 );
nand NAND2_2406 ( U5416 , ADD_95_U48 , U5743 );
nand NAND2_2407 ( U5417 , U4049 , U5414 );
nand NAND2_2408 ( U5418 , R1165_U17 , U3028 );
nand NAND2_2409 ( U5419 , REG3_REG_7_ , U3149 );
nand NAND2_2410 ( U5420 , U3455 , U3376 );
nand NAND2_2411 ( U5421 , U3454 , U5420 );
nand NAND3_2412 ( U5422 , U5802 , U3454 , R1165_U91 );
nand NAND2_2413 ( U5423 , U3014 , U3484 );
nand NAND2_2414 ( U5424 , U3582 , U3460 );
nand NAND2_2415 ( U5425 , U5805 , U3080 );
nand NAND2_2416 ( U5426 , U3014 , U3482 );
nand NAND2_2417 ( U5427 , U3583 , U3460 );
nand NAND2_2418 ( U5428 , U5805 , U3081 );
nand NAND2_2419 ( U5429 , U3014 , U3480 );
nand NAND2_2420 ( U5430 , U3584 , U3460 );
nand NAND2_2421 ( U5431 , U5805 , U3067 );
nand NAND2_2422 ( U5432 , U3014 , U3478 );
nand NAND2_2423 ( U5433 , U3585 , U3460 );
nand NAND2_2424 ( U5434 , U5805 , U3068 );
nand NAND2_2425 ( U5435 , U3014 , U3476 );
nand NAND2_2426 ( U5436 , U3586 , U3460 );
nand NAND2_2427 ( U5437 , U5805 , U3064 );
nand NAND2_2428 ( U5438 , U3014 , U3474 );
nand NAND2_2429 ( U5439 , U3587 , U3460 );
nand NAND2_2430 ( U5440 , U5805 , U3057 );
nand NAND2_2431 ( U5441 , U3588 , U3460 );
nand NAND2_2432 ( U5442 , U3014 , U4038 );
nand NAND2_2433 ( U5443 , U5805 , U3053 );
nand NAND2_2434 ( U5444 , U3589 , U3460 );
nand NAND2_2435 ( U5445 , U3014 , U4039 );
nand NAND2_2436 ( U5446 , U5805 , U3056 );
nand NAND2_2437 ( U5447 , U3014 , U3472 );
nand NAND2_2438 ( U5448 , U3590 , U3460 );
nand NAND2_2439 ( U5449 , U5805 , U3061 );
nand NAND2_2440 ( U5450 , U3591 , U3460 );
nand NAND2_2441 ( U5451 , U3014 , U4040 );
nand NAND2_2442 ( U5452 , U5805 , U3052 );
nand NAND2_2443 ( U5453 , U3592 , U3460 );
nand NAND2_2444 ( U5454 , U3014 , U4029 );
nand NAND2_2445 ( U5455 , U5805 , U3051 );
nand NAND2_2446 ( U5456 , U3593 , U3460 );
nand NAND2_2447 ( U5457 , U3014 , U4030 );
nand NAND2_2448 ( U5458 , U5805 , U3050 );
nand NAND2_2449 ( U5459 , U3594 , U3460 );
nand NAND2_2450 ( U5460 , U3014 , U4031 );
nand NAND2_2451 ( U5461 , U5805 , U3054 );
nand NAND2_2452 ( U5462 , U3595 , U3460 );
nand NAND2_2453 ( U5463 , U3014 , U4032 );
nand NAND2_2454 ( U5464 , U5805 , U3055 );
nand NAND2_2455 ( U5465 , U3596 , U3460 );
nand NAND2_2456 ( U5466 , U3014 , U4033 );
nand NAND2_2457 ( U5467 , U5805 , U3062 );
nand NAND2_2458 ( U5468 , U3597 , U3460 );
nand NAND2_2459 ( U5469 , U3014 , U4034 );
nand NAND2_2460 ( U5470 , U5805 , U3063 );
nand NAND2_2461 ( U5471 , U3598 , U3460 );
nand NAND2_2462 ( U5472 , U3014 , U4035 );
nand NAND2_2463 ( U5473 , U5805 , U3058 );
nand NAND2_2464 ( U5474 , U3599 , U3460 );
nand NAND2_2465 ( U5475 , U3014 , U4036 );
nand NAND2_2466 ( U5476 , U5805 , U3072 );
nand NAND2_2467 ( U5477 , U3600 , U3460 );
nand NAND2_2468 ( U5478 , U3014 , U4037 );
nand NAND2_2469 ( U5479 , U5805 , U3073 );
nand NAND2_2470 ( U5480 , U3014 , U3470 );
nand NAND2_2471 ( U5481 , U3601 , U3460 );
nand NAND2_2472 ( U5482 , U5805 , U3065 );
nand NAND2_2473 ( U5483 , U3014 , U3504 );
nand NAND2_2474 ( U5484 , U3602 , U3460 );
nand NAND2_2475 ( U5485 , U5805 , U3078 );
nand NAND2_2476 ( U5486 , U3014 , U3502 );
nand NAND2_2477 ( U5487 , U3603 , U3460 );
nand NAND2_2478 ( U5488 , U5805 , U3079 );
nand NAND2_2479 ( U5489 , U3014 , U3500 );
nand NAND2_2480 ( U5490 , U3604 , U3460 );
nand NAND2_2481 ( U5491 , U5805 , U3066 );
nand NAND2_2482 ( U5492 , U3014 , U3498 );
nand NAND2_2483 ( U5493 , U3605 , U3460 );
nand NAND2_2484 ( U5494 , U5805 , U3070 );
nand NAND2_2485 ( U5495 , U3014 , U3496 );
nand NAND2_2486 ( U5496 , U3606 , U3460 );
nand NAND2_2487 ( U5497 , U5805 , U3071 );
nand NAND2_2488 ( U5498 , U3014 , U3494 );
nand NAND2_2489 ( U5499 , U3607 , U3460 );
nand NAND2_2490 ( U5500 , U5805 , U3076 );
nand NAND2_2491 ( U5501 , U3014 , U3492 );
nand NAND2_2492 ( U5502 , U3608 , U3460 );
nand NAND2_2493 ( U5503 , U5805 , U3077 );
nand NAND2_2494 ( U5504 , U3014 , U3490 );
nand NAND2_2495 ( U5505 , U3609 , U3460 );
nand NAND2_2496 ( U5506 , U5805 , U3069 );
nand NAND2_2497 ( U5507 , U3014 , U3488 );
nand NAND2_2498 ( U5508 , U3610 , U3460 );
nand NAND2_2499 ( U5509 , U5805 , U3060 );
nand NAND2_2500 ( U5510 , U3014 , U3486 );
nand NAND2_2501 ( U5511 , U3611 , U3460 );
nand NAND2_2502 ( U5512 , U5805 , U3059 );
nand NAND2_2503 ( U5513 , U3014 , U3468 );
nand NAND2_2504 ( U5514 , U3612 , U3460 );
nand NAND2_2505 ( U5515 , U5805 , U3075 );
nand NAND2_2506 ( U5516 , U3014 , U3464 );
nand NAND2_2507 ( U5517 , U3613 , U3460 );
nand NAND2_2508 ( U5518 , U5805 , U3074 );
nand NAND2_2509 ( U5519 , U3484 , U3361 );
nand NAND2_2510 ( U5520 , U3014 , U3080 );
nand NAND2_2511 ( U5521 , U5748 , U3081 );
nand NAND2_2512 ( U5522 , U3482 , U3361 );
nand NAND2_2513 ( U5523 , U3014 , U3081 );
nand NAND2_2514 ( U5524 , U5748 , U3067 );
nand NAND2_2515 ( U5525 , U3480 , U3361 );
nand NAND2_2516 ( U5526 , U3014 , U3067 );
nand NAND2_2517 ( U5527 , U5748 , U3068 );
nand NAND2_2518 ( U5528 , U3478 , U3361 );
nand NAND2_2519 ( U5529 , U3014 , U3068 );
nand NAND2_2520 ( U5530 , U5748 , U3064 );
nand NAND2_2521 ( U5531 , U3476 , U3361 );
nand NAND2_2522 ( U5532 , U3014 , U3064 );
nand NAND2_2523 ( U5533 , U5748 , U3057 );
nand NAND2_2524 ( U5534 , U3474 , U3361 );
nand NAND2_2525 ( U5535 , U3014 , U3057 );
nand NAND2_2526 ( U5536 , U5748 , U3061 );
nand NAND2_2527 ( U5537 , U4038 , U3361 );
nand NAND2_2528 ( U5538 , U3014 , U3053 );
nand NAND2_2529 ( U5539 , U4039 , U3361 );
nand NAND2_2530 ( U5540 , U3014 , U3056 );
nand NAND2_2531 ( U5541 , U3472 , U3361 );
nand NAND2_2532 ( U5542 , U3014 , U3061 );
nand NAND2_2533 ( U5543 , U5748 , U3065 );
nand NAND2_2534 ( U5544 , U4040 , U3361 );
nand NAND2_2535 ( U5545 , U3014 , U3052 );
nand NAND2_2536 ( U5546 , U5748 , U3051 );
nand NAND2_2537 ( U5547 , U4029 , U3361 );
nand NAND2_2538 ( U5548 , U3014 , U3051 );
nand NAND2_2539 ( U5549 , U5748 , U3050 );
nand NAND2_2540 ( U5550 , U4030 , U3361 );
nand NAND2_2541 ( U5551 , U3014 , U3050 );
nand NAND2_2542 ( U5552 , U5748 , U3054 );
nand NAND2_2543 ( U5553 , U4031 , U3361 );
nand NAND2_2544 ( U5554 , U3014 , U3054 );
nand NAND2_2545 ( U5555 , U5748 , U3055 );
nand NAND2_2546 ( U5556 , U4032 , U3361 );
nand NAND2_2547 ( U5557 , U3014 , U3055 );
nand NAND2_2548 ( U5558 , U5748 , U3062 );
nand NAND2_2549 ( U5559 , U4033 , U3361 );
nand NAND2_2550 ( U5560 , U3014 , U3062 );
nand NAND2_2551 ( U5561 , U5748 , U3063 );
nand NAND2_2552 ( U5562 , U4034 , U3361 );
nand NAND2_2553 ( U5563 , U3014 , U3063 );
nand NAND2_2554 ( U5564 , U5748 , U3058 );
nand NAND2_2555 ( U5565 , U4035 , U3361 );
nand NAND2_2556 ( U5566 , U3014 , U3058 );
nand NAND2_2557 ( U5567 , U5748 , U3072 );
nand NAND2_2558 ( U5568 , U4036 , U3361 );
nand NAND2_2559 ( U5569 , U3014 , U3072 );
nand NAND2_2560 ( U5570 , U5748 , U3073 );
nand NAND2_2561 ( U5571 , U4037 , U3361 );
nand NAND2_2562 ( U5572 , U3014 , U3073 );
nand NAND2_2563 ( U5573 , U5748 , U3078 );
nand NAND2_2564 ( U5574 , U3470 , U3361 );
nand NAND2_2565 ( U5575 , U3014 , U3065 );
nand NAND2_2566 ( U5576 , U5748 , U3075 );
nand NAND2_2567 ( U5577 , U3504 , U3361 );
nand NAND2_2568 ( U5578 , U3014 , U3078 );
nand NAND2_2569 ( U5579 , U5748 , U3079 );
nand NAND2_2570 ( U5580 , U3502 , U3361 );
nand NAND2_2571 ( U5581 , U3014 , U3079 );
nand NAND2_2572 ( U5582 , U5748 , U3066 );
nand NAND2_2573 ( U5583 , U3500 , U3361 );
nand NAND2_2574 ( U5584 , U3014 , U3066 );
nand NAND2_2575 ( U5585 , U5748 , U3070 );
nand NAND2_2576 ( U5586 , U3498 , U3361 );
nand NAND2_2577 ( U5587 , U3014 , U3070 );
nand NAND2_2578 ( U5588 , U5748 , U3071 );
nand NAND2_2579 ( U5589 , U3496 , U3361 );
nand NAND2_2580 ( U5590 , U3014 , U3071 );
nand NAND2_2581 ( U5591 , U5748 , U3076 );
nand NAND2_2582 ( U5592 , U3494 , U3361 );
nand NAND2_2583 ( U5593 , U3014 , U3076 );
nand NAND2_2584 ( U5594 , U5748 , U3077 );
nand NAND2_2585 ( U5595 , U3492 , U3361 );
nand NAND2_2586 ( U5596 , U3014 , U3077 );
nand NAND2_2587 ( U5597 , U5748 , U3069 );
nand NAND2_2588 ( U5598 , U3490 , U3361 );
nand NAND2_2589 ( U5599 , U3014 , U3069 );
nand NAND2_2590 ( U5600 , U5748 , U3060 );
nand NAND2_2591 ( U5601 , U3488 , U3361 );
nand NAND2_2592 ( U5602 , U3014 , U3060 );
nand NAND2_2593 ( U5603 , U5748 , U3059 );
nand NAND2_2594 ( U5604 , U3486 , U3361 );
nand NAND2_2595 ( U5605 , U3014 , U3059 );
nand NAND2_2596 ( U5606 , U5748 , U3080 );
nand NAND2_2597 ( U5607 , U3468 , U3361 );
nand NAND2_2598 ( U5608 , U3014 , U3075 );
nand NAND2_2599 ( U5609 , U5748 , U3074 );
nand NAND2_2600 ( U5610 , U3464 , U3361 );
nand NAND2_2601 ( U5611 , U3014 , U3074 );
nand NAND2_2602 ( U5612 , U3963 , U4026 );
nand NAND2_2603 ( U5613 , U3370 , U3419 );
nand NAND4_2604 ( U5614 , U3374 , U3368 , U3366 , U3367 );
nand NAND2_2605 ( U5615 , U5614 , U3355 );
nand NAND2_2606 ( U5616 , U4057 , U3355 );
nand NAND2_2607 ( U5617 , U5616 , U5615 );
nand NAND2_2608 ( U5618 , U3964 , U5615 );
nand NAND2_2609 ( U5619 , U3484 , U5618 );
nand NAND2_2610 ( U5620 , U3022 , U3080 );
nand NAND2_2611 ( U5621 , U3482 , U5618 );
nand NAND2_2612 ( U5622 , U3022 , U3081 );
nand NAND2_2613 ( U5623 , U3480 , U5618 );
nand NAND2_2614 ( U5624 , U3022 , U3067 );
nand NAND2_2615 ( U5625 , U3478 , U5618 );
nand NAND2_2616 ( U5626 , U3022 , U3068 );
nand NAND2_2617 ( U5627 , U3476 , U5618 );
nand NAND2_2618 ( U5628 , U3022 , U3064 );
nand NAND2_2619 ( U5629 , U3474 , U5618 );
nand NAND2_2620 ( U5630 , U3022 , U3057 );
nand NAND2_2621 ( U5631 , U3472 , U5618 );
nand NAND2_2622 ( U5632 , U3022 , U3061 );
nand NAND2_2623 ( U5633 , U4029 , U5618 );
nand NAND2_2624 ( U5634 , U3022 , U3051 );
nand NAND2_2625 ( U5635 , U4030 , U5618 );
nand NAND2_2626 ( U5636 , U3022 , U3050 );
nand NAND2_2627 ( U5637 , U4031 , U5618 );
nand NAND2_2628 ( U5638 , U3022 , U3054 );
nand NAND2_2629 ( U5639 , U4032 , U5618 );
nand NAND2_2630 ( U5640 , U3022 , U3055 );
nand NAND2_2631 ( U5641 , U4033 , U5618 );
nand NAND2_2632 ( U5642 , U3022 , U3062 );
nand NAND2_2633 ( U5643 , U4034 , U5618 );
nand NAND2_2634 ( U5644 , U3022 , U3063 );
nand NAND2_2635 ( U5645 , U4035 , U5618 );
nand NAND2_2636 ( U5646 , U3022 , U3058 );
nand NAND2_2637 ( U5647 , U4036 , U5618 );
nand NAND2_2638 ( U5648 , U3022 , U3072 );
nand NAND2_2639 ( U5649 , U4037 , U5618 );
nand NAND2_2640 ( U5650 , U3022 , U3073 );
nand NAND2_2641 ( U5651 , U3470 , U5618 );
nand NAND2_2642 ( U5652 , U3022 , U3065 );
nand NAND2_2643 ( U5653 , U3504 , U5618 );
nand NAND2_2644 ( U5654 , U3022 , U3078 );
nand NAND2_2645 ( U5655 , U3502 , U5618 );
nand NAND2_2646 ( U5656 , U3022 , U3079 );
nand NAND2_2647 ( U5657 , U3500 , U5618 );
nand NAND2_2648 ( U5658 , U3022 , U3066 );
nand NAND2_2649 ( U5659 , U3498 , U5618 );
nand NAND2_2650 ( U5660 , U3022 , U3070 );
nand NAND2_2651 ( U5661 , U3496 , U5618 );
nand NAND2_2652 ( U5662 , U3022 , U3071 );
nand NAND2_2653 ( U5663 , U3494 , U5618 );
nand NAND2_2654 ( U5664 , U3022 , U3076 );
nand NAND2_2655 ( U5665 , U3492 , U5618 );
nand NAND2_2656 ( U5666 , U3022 , U3077 );
nand NAND2_2657 ( U5667 , U3490 , U5618 );
nand NAND2_2658 ( U5668 , U3022 , U3069 );
nand NAND2_2659 ( U5669 , U3488 , U5618 );
nand NAND2_2660 ( U5670 , U3022 , U3060 );
nand NAND2_2661 ( U5671 , U3486 , U5618 );
nand NAND2_2662 ( U5672 , U3022 , U3059 );
nand NAND2_2663 ( U5673 , U3468 , U5618 );
nand NAND2_2664 ( U5674 , U3022 , U3075 );
nand NAND2_2665 ( U5675 , U3464 , U5618 );
nand NAND2_2666 ( U5676 , U3022 , U3074 );
nand NAND2_2667 ( U5677 , REG1_REG_0_ , U4059 );
nand NAND2_2668 ( U5678 , U3022 , U3484 );
nand NAND2_2669 ( U5679 , U5617 , U3080 );
nand NAND2_2670 ( U5680 , U3022 , U3482 );
nand NAND2_2671 ( U5681 , U5617 , U3081 );
nand NAND2_2672 ( U5682 , U3022 , U3480 );
nand NAND2_2673 ( U5683 , U5617 , U3067 );
nand NAND2_2674 ( U5684 , U3022 , U3478 );
nand NAND2_2675 ( U5685 , U5617 , U3068 );
nand NAND2_2676 ( U5686 , U3022 , U3476 );
nand NAND2_2677 ( U5687 , U5617 , U3064 );
nand NAND2_2678 ( U5688 , U3022 , U3474 );
nand NAND2_2679 ( U5689 , U5617 , U3057 );
nand NAND2_2680 ( U5690 , U3022 , U3472 );
nand NAND2_2681 ( U5691 , U5617 , U3061 );
nand NAND2_2682 ( U5692 , U3022 , U4029 );
nand NAND2_2683 ( U5693 , U5617 , U3051 );
nand NAND2_2684 ( U5694 , U3022 , U4030 );
nand NAND2_2685 ( U5695 , U5617 , U3050 );
nand NAND2_2686 ( U5696 , U3022 , U4031 );
nand NAND2_2687 ( U5697 , U5617 , U3054 );
nand NAND2_2688 ( U5698 , U3022 , U4032 );
nand NAND2_2689 ( U5699 , U5617 , U3055 );
nand NAND2_2690 ( U5700 , U3022 , U4033 );
nand NAND2_2691 ( U5701 , U5617 , U3062 );
nand NAND2_2692 ( U5702 , U3022 , U4034 );
nand NAND2_2693 ( U5703 , U5617 , U3063 );
nand NAND2_2694 ( U5704 , U3022 , U4035 );
nand NAND2_2695 ( U5705 , U5617 , U3058 );
nand NAND2_2696 ( U5706 , U3022 , U4036 );
nand NAND2_2697 ( U5707 , U5617 , U3072 );
nand NAND2_2698 ( U5708 , U3022 , U4037 );
nand NAND2_2699 ( U5709 , U5617 , U3073 );
nand NAND2_2700 ( U5710 , U3022 , U3470 );
nand NAND2_2701 ( U5711 , U5617 , U3065 );
nand NAND2_2702 ( U5712 , U3022 , U3504 );
nand NAND2_2703 ( U5713 , U5617 , U3078 );
nand NAND2_2704 ( U5714 , U3022 , U3502 );
nand NAND2_2705 ( U5715 , U5617 , U3079 );
nand NAND2_2706 ( U5716 , U3022 , U3500 );
nand NAND2_2707 ( U5717 , U5617 , U3066 );
nand NAND2_2708 ( U5718 , U3022 , U3498 );
nand NAND2_2709 ( U5719 , U5617 , U3070 );
nand NAND2_2710 ( U5720 , U3022 , U3496 );
nand NAND2_2711 ( U5721 , U5617 , U3071 );
nand NAND2_2712 ( U5722 , U3022 , U3494 );
nand NAND2_2713 ( U5723 , U5617 , U3076 );
nand NAND2_2714 ( U5724 , U3022 , U3492 );
nand NAND2_2715 ( U5725 , U5617 , U3077 );
nand NAND2_2716 ( U5726 , U3022 , U3490 );
nand NAND2_2717 ( U5727 , U5617 , U3069 );
nand NAND2_2718 ( U5728 , U3022 , U3488 );
nand NAND2_2719 ( U5729 , U5617 , U3060 );
nand NAND2_2720 ( U5730 , U3022 , U3486 );
nand NAND2_2721 ( U5731 , U5617 , U3059 );
nand NAND2_2722 ( U5732 , U3022 , U3468 );
nand NAND2_2723 ( U5733 , U5617 , U3075 );
nand NAND2_2724 ( U5734 , U3022 , U3464 );
nand NAND2_2725 ( U5735 , U5617 , U3074 );
nand NAND2_2726 ( U5736 , U4059 , U3453 );
nand NAND2_2727 ( U5737 , R1207_U28 , U4013 );
nand NAND2_2728 ( U5738 , R1192_U28 , U4014 );
nand NAND2_2729 ( U5739 , R1150_U27 , U4016 );
nand NAND2_2730 ( U5740 , R1117_U26 , U4018 );
nand NAND2_2731 ( U5741 , U4052 , U3427 );
nand NAND2_2732 ( U5742 , U4028 , U4052 );
nand NAND2_2733 ( U5743 , U5741 , U4050 );
nand NAND2_2734 ( U5744 , U5742 , U4051 );
nand NAND2_2735 ( U5745 , U5754 , U5751 );
nand NAND2_2736 ( U5746 , IR_REG_23_ , U3967 );
nand NAND2_2737 ( U5747 , IR_REG_31_ , SUB_84_U81 );
not NOT1_2738 ( U5748 , U3431 );
nand NAND2_2739 ( U5749 , IR_REG_24_ , U3967 );
nand NAND2_2740 ( U5750 , IR_REG_31_ , SUB_84_U78 );
not NOT1_2741 ( U5751 , U3434 );
nand NAND2_2742 ( U5752 , IR_REG_26_ , U3967 );
nand NAND2_2743 ( U5753 , IR_REG_31_ , SUB_84_U17 );
not NOT1_2744 ( U5754 , U3432 );
nand NAND2_2745 ( U5755 , IR_REG_25_ , U3967 );
nand NAND2_2746 ( U5756 , IR_REG_31_ , SUB_84_U16 );
not NOT1_2747 ( U5757 , U3433 );
nand NAND2_2748 ( U5758 , IR_REG_9_ , U3967 );
nand NAND2_2749 ( U5759 , IR_REG_31_ , SUB_84_U25 );
nand NAND2_2750 ( U5760 , IR_REG_8_ , U3967 );
nand NAND2_2751 ( U5761 , IR_REG_31_ , SUB_84_U68 );
nand NAND2_2752 ( U5762 , IR_REG_7_ , U3967 );
nand NAND2_2753 ( U5763 , IR_REG_31_ , SUB_84_U24 );
nand NAND2_2754 ( U5764 , IR_REG_6_ , U3967 );
nand NAND2_2755 ( U5765 , IR_REG_31_ , SUB_84_U23 );
nand NAND2_2756 ( U5766 , IR_REG_5_ , U3967 );
nand NAND2_2757 ( U5767 , IR_REG_31_ , SUB_84_U22 );
nand NAND2_2758 ( U5768 , IR_REG_4_ , U3967 );
nand NAND2_2759 ( U5769 , IR_REG_31_ , SUB_84_U70 );
nand NAND2_2760 ( U5770 , IR_REG_3_ , U3967 );
nand NAND2_2761 ( U5771 , IR_REG_31_ , SUB_84_U21 );
nand NAND2_2762 ( U5772 , IR_REG_2_ , U3967 );
nand NAND2_2763 ( U5773 , IR_REG_31_ , SUB_84_U20 );
nand NAND2_2764 ( U5774 , IR_REG_1_ , U3967 );
nand NAND2_2765 ( U5775 , IR_REG_31_ , SUB_84_U48 );
nand NAND2_2766 ( U5776 , IR_REG_18_ , U3967 );
nand NAND2_2767 ( U5777 , IR_REG_31_ , SUB_84_U12 );
nand NAND2_2768 ( U5778 , IR_REG_17_ , U3967 );
nand NAND2_2769 ( U5779 , IR_REG_31_ , SUB_84_U11 );
nand NAND2_2770 ( U5780 , IR_REG_16_ , U3967 );
nand NAND2_2771 ( U5781 , IR_REG_31_ , SUB_84_U87 );
nand NAND2_2772 ( U5782 , IR_REG_15_ , U3967 );
nand NAND2_2773 ( U5783 , IR_REG_31_ , SUB_84_U10 );
nand NAND2_2774 ( U5784 , IR_REG_14_ , U3967 );
nand NAND2_2775 ( U5785 , IR_REG_31_ , SUB_84_U9 );
nand NAND2_2776 ( U5786 , IR_REG_13_ , U3967 );
nand NAND2_2777 ( U5787 , IR_REG_31_ , SUB_84_U8 );
nand NAND2_2778 ( U5788 , IR_REG_12_ , U3967 );
nand NAND2_2779 ( U5789 , IR_REG_31_ , SUB_84_U89 );
nand NAND2_2780 ( U5790 , IR_REG_11_ , U3967 );
nand NAND2_2781 ( U5791 , IR_REG_31_ , SUB_84_U7 );
nand NAND2_2782 ( U5792 , IR_REG_10_ , U3967 );
nand NAND2_2783 ( U5793 , IR_REG_31_ , SUB_84_U6 );
nand NAND2_2784 ( U5794 , IR_REG_0_ , U3967 );
nand NAND2_2785 ( U5795 , IR_REG_31_ , IR_REG_0_ );
not NOT1_2786 ( U5796 , U3453 );
nand NAND2_2787 ( U5797 , IR_REG_28_ , U3967 );
nand NAND2_2788 ( U5798 , IR_REG_31_ , SUB_84_U18 );
not NOT1_2789 ( U5799 , U3454 );
nand NAND2_2790 ( U5800 , IR_REG_27_ , U3967 );
nand NAND2_2791 ( U5801 , IR_REG_31_ , SUB_84_U76 );
not NOT1_2792 ( U5802 , U3455 );
nand NAND2_2793 ( U5803 , IR_REG_22_ , U3967 );
nand NAND2_2794 ( U5804 , IR_REG_31_ , SUB_84_U15 );
not NOT1_2795 ( U5805 , U3456 );
nand NAND2_2796 ( U5806 , IR_REG_21_ , U3967 );
nand NAND2_2797 ( U5807 , IR_REG_31_ , SUB_84_U14 );
not NOT1_2798 ( U5808 , U3457 );
nand NAND2_2799 ( U5809 , U3434 , U3359 );
nand NAND3_2800 ( U5810 , U4058 , U5751 , B_REG );
nand NAND2_2801 ( U5811 , D_REG_0_ , U3968 );
nand NAND2_2802 ( U5812 , U4047 , U4162 );
nand NAND2_2803 ( U5813 , D_REG_1_ , U3968 );
nand NAND2_2804 ( U5814 , U4047 , U4163 );
nand NAND2_2805 ( U5815 , IR_REG_19_ , U3967 );
nand NAND2_2806 ( U5816 , IR_REG_31_ , SUB_84_U13 );
not NOT1_2807 ( U5817 , U3461 );
nand NAND2_2808 ( U5818 , IR_REG_20_ , U3967 );
nand NAND2_2809 ( U5819 , IR_REG_31_ , SUB_84_U83 );
not NOT1_2810 ( U5820 , U3460 );
nand NAND2_2811 ( U5821 , IR_REG_30_ , U3967 );
nand NAND2_2812 ( U5822 , IR_REG_31_ , SUB_84_U73 );
not NOT1_2813 ( U5823 , U3462 );
nand NAND2_2814 ( U5824 , IR_REG_29_ , U3967 );
nand NAND2_2815 ( U5825 , IR_REG_31_ , SUB_84_U19 );
not NOT1_2816 ( U5826 , U3463 );
nand NAND2_2817 ( U5827 , DATAI_0_ , U3969 );
nand NAND2_2818 ( U5828 , U4027 , U3453 );
not NOT1_2819 ( U5829 , U3464 );
nand NAND2_2820 ( U5830 , U3456 , U5808 );
nand NAND2_2821 ( U5831 , U3457 , U5805 );
nand NAND2_2822 ( U5832 , D_REG_1_ , U4161 );
nand NAND2_2823 ( U5833 , U4163 , U3360 );
not NOT1_2824 ( U5834 , U3466 );
nand NAND2_2825 ( U5835 , U5745 , U3360 );
nand NAND2_2826 ( U5836 , D_REG_0_ , U4161 );
not NOT1_2827 ( U5837 , U3465 );
nand NAND2_2828 ( U5838 , REG0_REG_0_ , U3970 );
nand NAND2_2829 ( U5839 , U4046 , U4214 );
nand NAND2_2830 ( U5840 , DATAI_1_ , U3969 );
nand NAND2_2831 ( U5841 , U4027 , U3443 );
not NOT1_2832 ( U5842 , U3468 );
nand NAND2_2833 ( U5843 , REG0_REG_1_ , U3970 );
nand NAND2_2834 ( U5844 , U4046 , U4238 );
nand NAND2_2835 ( U5845 , DATAI_2_ , U3969 );
nand NAND2_2836 ( U5846 , U4027 , U3442 );
not NOT1_2837 ( U5847 , U3470 );
nand NAND2_2838 ( U5848 , REG0_REG_2_ , U3970 );
nand NAND2_2839 ( U5849 , U4046 , U4257 );
nand NAND2_2840 ( U5850 , DATAI_3_ , U3969 );
nand NAND2_2841 ( U5851 , U4027 , U3441 );
not NOT1_2842 ( U5852 , U3472 );
nand NAND2_2843 ( U5853 , REG0_REG_3_ , U3970 );
nand NAND2_2844 ( U5854 , U4046 , U4276 );
nand NAND2_2845 ( U5855 , DATAI_4_ , U3969 );
nand NAND2_2846 ( U5856 , U4027 , U3440 );
not NOT1_2847 ( U5857 , U3474 );
nand NAND2_2848 ( U5858 , REG0_REG_4_ , U3970 );
nand NAND2_2849 ( U5859 , U4046 , U4295 );
nand NAND2_2850 ( U5860 , DATAI_5_ , U3969 );
nand NAND2_2851 ( U5861 , U4027 , U3439 );
not NOT1_2852 ( U5862 , U3476 );
nand NAND2_2853 ( U5863 , REG0_REG_5_ , U3970 );
nand NAND2_2854 ( U5864 , U4046 , U4314 );
nand NAND2_2855 ( U5865 , DATAI_6_ , U3969 );
nand NAND2_2856 ( U5866 , U4027 , U3438 );
not NOT1_2857 ( U5867 , U3478 );
nand NAND2_2858 ( U5868 , REG0_REG_6_ , U3970 );
nand NAND2_2859 ( U5869 , U4046 , U4333 );
nand NAND2_2860 ( U5870 , DATAI_7_ , U3969 );
nand NAND2_2861 ( U5871 , U4027 , U3437 );
not NOT1_2862 ( U5872 , U3480 );
nand NAND2_2863 ( U5873 , REG0_REG_7_ , U3970 );
nand NAND2_2864 ( U5874 , U4046 , U4352 );
nand NAND2_2865 ( U5875 , DATAI_8_ , U3969 );
nand NAND2_2866 ( U5876 , U4027 , U3436 );
not NOT1_2867 ( U5877 , U3482 );
nand NAND2_2868 ( U5878 , REG0_REG_8_ , U3970 );
nand NAND2_2869 ( U5879 , U4046 , U4371 );
nand NAND2_2870 ( U5880 , DATAI_9_ , U3969 );
nand NAND2_2871 ( U5881 , U4027 , U3435 );
not NOT1_2872 ( U5882 , U3484 );
nand NAND2_2873 ( U5883 , REG0_REG_9_ , U3970 );
nand NAND2_2874 ( U5884 , U4046 , U4390 );
nand NAND2_2875 ( U5885 , DATAI_10_ , U3969 );
nand NAND2_2876 ( U5886 , U4027 , U3452 );
not NOT1_2877 ( U5887 , U3486 );
nand NAND2_2878 ( U5888 , REG0_REG_10_ , U3970 );
nand NAND2_2879 ( U5889 , U4046 , U4409 );
nand NAND2_2880 ( U5890 , DATAI_11_ , U3969 );
nand NAND2_2881 ( U5891 , U4027 , U3451 );
not NOT1_2882 ( U5892 , U3488 );
nand NAND2_2883 ( U5893 , REG0_REG_11_ , U3970 );
nand NAND2_2884 ( U5894 , U4046 , U4428 );
nand NAND2_2885 ( U5895 , DATAI_12_ , U3969 );
nand NAND2_2886 ( U5896 , U4027 , U3450 );
not NOT1_2887 ( U5897 , U3490 );
nand NAND2_2888 ( U5898 , REG0_REG_12_ , U3970 );
nand NAND2_2889 ( U5899 , U4046 , U4447 );
nand NAND2_2890 ( U5900 , DATAI_13_ , U3969 );
nand NAND2_2891 ( U5901 , U4027 , U3449 );
not NOT1_2892 ( U5902 , U3492 );
nand NAND2_2893 ( U5903 , REG0_REG_13_ , U3970 );
nand NAND2_2894 ( U5904 , U4046 , U4466 );
nand NAND2_2895 ( U5905 , DATAI_14_ , U3969 );
nand NAND2_2896 ( U5906 , U4027 , U3448 );
not NOT1_2897 ( U5907 , U3494 );
nand NAND2_2898 ( U5908 , REG0_REG_14_ , U3970 );
nand NAND2_2899 ( U5909 , U4046 , U4485 );
nand NAND2_2900 ( U5910 , DATAI_15_ , U3969 );
nand NAND2_2901 ( U5911 , U4027 , U3447 );
not NOT1_2902 ( U5912 , U3496 );
nand NAND2_2903 ( U5913 , REG0_REG_15_ , U3970 );
nand NAND2_2904 ( U5914 , U4046 , U4504 );
nand NAND2_2905 ( U5915 , DATAI_16_ , U3969 );
nand NAND2_2906 ( U5916 , U4027 , U3446 );
not NOT1_2907 ( U5917 , U3498 );
nand NAND2_2908 ( U5918 , REG0_REG_16_ , U3970 );
nand NAND2_2909 ( U5919 , U4046 , U4523 );
nand NAND2_2910 ( U5920 , DATAI_17_ , U3969 );
nand NAND2_2911 ( U5921 , U4027 , U3445 );
not NOT1_2912 ( U5922 , U3500 );
nand NAND2_2913 ( U5923 , REG0_REG_17_ , U3970 );
nand NAND2_2914 ( U5924 , U4046 , U4542 );
nand NAND2_2915 ( U5925 , DATAI_18_ , U3969 );
nand NAND2_2916 ( U5926 , U4027 , U3444 );
not NOT1_2917 ( U5927 , U3502 );
nand NAND2_2918 ( U5928 , REG0_REG_18_ , U3970 );
nand NAND2_2919 ( U5929 , U4046 , U4561 );
nand NAND2_2920 ( U5930 , DATAI_19_ , U3969 );
nand NAND2_2921 ( U5931 , U4027 , U3461 );
not NOT1_2922 ( U5932 , U3504 );
nand NAND2_2923 ( U5933 , REG0_REG_19_ , U3970 );
nand NAND2_2924 ( U5934 , U4046 , U4580 );
nand NAND2_2925 ( U5935 , REG0_REG_20_ , U3970 );
nand NAND2_2926 ( U5936 , U4046 , U4599 );
nand NAND2_2927 ( U5937 , REG0_REG_21_ , U3970 );
nand NAND2_2928 ( U5938 , U4046 , U4618 );
nand NAND2_2929 ( U5939 , REG0_REG_22_ , U3970 );
nand NAND2_2930 ( U5940 , U4046 , U4637 );
nand NAND2_2931 ( U5941 , REG0_REG_23_ , U3970 );
nand NAND2_2932 ( U5942 , U4046 , U4656 );
nand NAND2_2933 ( U5943 , REG0_REG_24_ , U3970 );
nand NAND2_2934 ( U5944 , U4046 , U4675 );
nand NAND2_2935 ( U5945 , REG0_REG_25_ , U3970 );
nand NAND2_2936 ( U5946 , U4046 , U4694 );
nand NAND2_2937 ( U5947 , REG0_REG_26_ , U3970 );
nand NAND2_2938 ( U5948 , U4046 , U4713 );
nand NAND2_2939 ( U5949 , REG0_REG_27_ , U3970 );
nand NAND2_2940 ( U5950 , U4046 , U4732 );
nand NAND2_2941 ( U5951 , REG0_REG_28_ , U3970 );
nand NAND2_2942 ( U5952 , U4046 , U4751 );
nand NAND2_2943 ( U5953 , REG0_REG_29_ , U3970 );
nand NAND2_2944 ( U5954 , U4046 , U4771 );
nand NAND2_2945 ( U5955 , REG0_REG_30_ , U3970 );
nand NAND2_2946 ( U5956 , U4046 , U4778 );
nand NAND2_2947 ( U5957 , REG0_REG_31_ , U3970 );
nand NAND2_2948 ( U5958 , U4046 , U4781 );
nand NAND2_2949 ( U5959 , REG1_REG_0_ , U3971 );
nand NAND2_2950 ( U5960 , U4045 , U4214 );
nand NAND2_2951 ( U5961 , REG1_REG_1_ , U3971 );
nand NAND2_2952 ( U5962 , U4045 , U4238 );
nand NAND2_2953 ( U5963 , REG1_REG_2_ , U3971 );
nand NAND2_2954 ( U5964 , U4045 , U4257 );
nand NAND2_2955 ( U5965 , REG1_REG_3_ , U3971 );
nand NAND2_2956 ( U5966 , U4045 , U4276 );
nand NAND2_2957 ( U5967 , REG1_REG_4_ , U3971 );
nand NAND2_2958 ( U5968 , U4045 , U4295 );
nand NAND2_2959 ( U5969 , REG1_REG_5_ , U3971 );
nand NAND2_2960 ( U5970 , U4045 , U4314 );
nand NAND2_2961 ( U5971 , REG1_REG_6_ , U3971 );
nand NAND2_2962 ( U5972 , U4045 , U4333 );
nand NAND2_2963 ( U5973 , REG1_REG_7_ , U3971 );
nand NAND2_2964 ( U5974 , U4045 , U4352 );
nand NAND2_2965 ( U5975 , REG1_REG_8_ , U3971 );
nand NAND2_2966 ( U5976 , U4045 , U4371 );
nand NAND2_2967 ( U5977 , REG1_REG_9_ , U3971 );
nand NAND2_2968 ( U5978 , U4045 , U4390 );
nand NAND2_2969 ( U5979 , REG1_REG_10_ , U3971 );
nand NAND2_2970 ( U5980 , U4045 , U4409 );
nand NAND2_2971 ( U5981 , REG1_REG_11_ , U3971 );
nand NAND2_2972 ( U5982 , U4045 , U4428 );
nand NAND2_2973 ( U5983 , REG1_REG_12_ , U3971 );
nand NAND2_2974 ( U5984 , U4045 , U4447 );
nand NAND2_2975 ( U5985 , REG1_REG_13_ , U3971 );
nand NAND2_2976 ( U5986 , U4045 , U4466 );
nand NAND2_2977 ( U5987 , REG1_REG_14_ , U3971 );
nand NAND2_2978 ( U5988 , U4045 , U4485 );
nand NAND2_2979 ( U5989 , REG1_REG_15_ , U3971 );
nand NAND2_2980 ( U5990 , U4045 , U4504 );
nand NAND2_2981 ( U5991 , REG1_REG_16_ , U3971 );
nand NAND2_2982 ( U5992 , U4045 , U4523 );
nand NAND2_2983 ( U5993 , REG1_REG_17_ , U3971 );
nand NAND2_2984 ( U5994 , U4045 , U4542 );
nand NAND2_2985 ( U5995 , REG1_REG_18_ , U3971 );
nand NAND2_2986 ( U5996 , U4045 , U4561 );
nand NAND2_2987 ( U5997 , REG1_REG_19_ , U3971 );
nand NAND2_2988 ( U5998 , U4045 , U4580 );
nand NAND2_2989 ( U5999 , REG1_REG_20_ , U3971 );
nand NAND2_2990 ( U6000 , U4045 , U4599 );
nand NAND2_2991 ( U6001 , REG1_REG_21_ , U3971 );
nand NAND2_2992 ( U6002 , U4045 , U4618 );
nand NAND2_2993 ( U6003 , REG1_REG_22_ , U3971 );
nand NAND2_2994 ( U6004 , U4045 , U4637 );
nand NAND2_2995 ( U6005 , REG1_REG_23_ , U3971 );
nand NAND2_2996 ( U6006 , U4045 , U4656 );
nand NAND2_2997 ( U6007 , REG1_REG_24_ , U3971 );
nand NAND2_2998 ( U6008 , U4045 , U4675 );
nand NAND2_2999 ( U6009 , REG1_REG_25_ , U3971 );
nand NAND2_3000 ( U6010 , U4045 , U4694 );
nand NAND2_3001 ( U6011 , REG1_REG_26_ , U3971 );
nand NAND2_3002 ( U6012 , U4045 , U4713 );
nand NAND2_3003 ( U6013 , REG1_REG_27_ , U3971 );
nand NAND2_3004 ( U6014 , U4045 , U4732 );
nand NAND2_3005 ( U6015 , REG1_REG_28_ , U3971 );
nand NAND2_3006 ( U6016 , U4045 , U4751 );
nand NAND2_3007 ( U6017 , REG1_REG_29_ , U3971 );
nand NAND2_3008 ( U6018 , U4045 , U4771 );
nand NAND2_3009 ( U6019 , REG1_REG_30_ , U3971 );
nand NAND2_3010 ( U6020 , U4045 , U4778 );
nand NAND2_3011 ( U6021 , REG1_REG_31_ , U3971 );
nand NAND2_3012 ( U6022 , U4045 , U4781 );
nand NAND2_3013 ( U6023 , REG2_REG_0_ , U3417 );
nand NAND2_3014 ( U6024 , U4044 , U3375 );
nand NAND2_3015 ( U6025 , REG2_REG_1_ , U3417 );
nand NAND2_3016 ( U6026 , U4044 , U3377 );
nand NAND2_3017 ( U6027 , REG2_REG_2_ , U3417 );
nand NAND2_3018 ( U6028 , U4044 , U3378 );
nand NAND2_3019 ( U6029 , REG2_REG_3_ , U3417 );
nand NAND2_3020 ( U6030 , U4044 , U3379 );
nand NAND2_3021 ( U6031 , REG2_REG_4_ , U3417 );
nand NAND2_3022 ( U6032 , U4044 , U3380 );
nand NAND2_3023 ( U6033 , REG2_REG_5_ , U3417 );
nand NAND2_3024 ( U6034 , U4044 , U3381 );
nand NAND2_3025 ( U6035 , REG2_REG_6_ , U3417 );
nand NAND2_3026 ( U6036 , U4044 , U3382 );
nand NAND2_3027 ( U6037 , REG2_REG_7_ , U3417 );
nand NAND2_3028 ( U6038 , U4044 , U3383 );
nand NAND2_3029 ( U6039 , REG2_REG_8_ , U3417 );
nand NAND2_3030 ( U6040 , U4044 , U3384 );
nand NAND2_3031 ( U6041 , REG2_REG_9_ , U3417 );
nand NAND2_3032 ( U6042 , U4044 , U3385 );
nand NAND2_3033 ( U6043 , REG2_REG_10_ , U3417 );
nand NAND2_3034 ( U6044 , U4044 , U3386 );
nand NAND2_3035 ( U6045 , REG2_REG_11_ , U3417 );
nand NAND2_3036 ( U6046 , U4044 , U3387 );
nand NAND2_3037 ( U6047 , REG2_REG_12_ , U3417 );
nand NAND2_3038 ( U6048 , U4044 , U3388 );
nand NAND2_3039 ( U6049 , REG2_REG_13_ , U3417 );
nand NAND2_3040 ( U6050 , U4044 , U3389 );
nand NAND2_3041 ( U6051 , REG2_REG_14_ , U3417 );
nand NAND2_3042 ( U6052 , U4044 , U3390 );
nand NAND2_3043 ( U6053 , REG2_REG_15_ , U3417 );
nand NAND2_3044 ( U6054 , U4044 , U3391 );
nand NAND2_3045 ( U6055 , REG2_REG_16_ , U3417 );
nand NAND2_3046 ( U6056 , U4044 , U3392 );
nand NAND2_3047 ( U6057 , REG2_REG_17_ , U3417 );
nand NAND2_3048 ( U6058 , U4044 , U3393 );
nand NAND2_3049 ( U6059 , REG2_REG_18_ , U3417 );
nand NAND2_3050 ( U6060 , U4044 , U3394 );
nand NAND2_3051 ( U6061 , REG2_REG_19_ , U3417 );
nand NAND2_3052 ( U6062 , U4044 , U3395 );
nand NAND2_3053 ( U6063 , REG2_REG_20_ , U3417 );
nand NAND2_3054 ( U6064 , U4044 , U3397 );
nand NAND2_3055 ( U6065 , REG2_REG_21_ , U3417 );
nand NAND2_3056 ( U6066 , U4044 , U3399 );
nand NAND2_3057 ( U6067 , REG2_REG_22_ , U3417 );
nand NAND2_3058 ( U6068 , U4044 , U3401 );
nand NAND2_3059 ( U6069 , REG2_REG_23_ , U3417 );
nand NAND2_3060 ( U6070 , U4044 , U3403 );
nand NAND2_3061 ( U6071 , REG2_REG_24_ , U3417 );
nand NAND2_3062 ( U6072 , U4044 , U3405 );
nand NAND2_3063 ( U6073 , REG2_REG_25_ , U3417 );
nand NAND2_3064 ( U6074 , U4044 , U3407 );
nand NAND2_3065 ( U6075 , REG2_REG_26_ , U3417 );
nand NAND2_3066 ( U6076 , U4044 , U3409 );
nand NAND2_3067 ( U6077 , REG2_REG_27_ , U3417 );
nand NAND2_3068 ( U6078 , U4044 , U3411 );
nand NAND2_3069 ( U6079 , REG2_REG_28_ , U3417 );
nand NAND2_3070 ( U6080 , U4044 , U3413 );
nand NAND2_3071 ( U6081 , REG2_REG_29_ , U3417 );
nand NAND2_3072 ( U6082 , U4044 , U4767 );
nand NAND2_3073 ( U6083 , REG2_REG_30_ , U3417 );
nand NAND2_3074 ( U6084 , U4048 , U4044 );
nand NAND2_3075 ( U6085 , REG2_REG_31_ , U3417 );
nand NAND2_3076 ( U6086 , U4048 , U4044 );
nand NAND2_3077 ( U6087 , DATAO_REG_0_ , U3422 );
nand NAND2_3078 ( U6088 , U4043 , U3074 );
nand NAND2_3079 ( U6089 , DATAO_REG_1_ , U3422 );
nand NAND2_3080 ( U6090 , U4043 , U3075 );
nand NAND2_3081 ( U6091 , DATAO_REG_2_ , U3422 );
nand NAND2_3082 ( U6092 , U4043 , U3065 );
nand NAND2_3083 ( U6093 , DATAO_REG_3_ , U3422 );
nand NAND2_3084 ( U6094 , U4043 , U3061 );
nand NAND2_3085 ( U6095 , DATAO_REG_4_ , U3422 );
nand NAND2_3086 ( U6096 , U4043 , U3057 );
nand NAND2_3087 ( U6097 , DATAO_REG_5_ , U3422 );
nand NAND2_3088 ( U6098 , U4043 , U3064 );
nand NAND2_3089 ( U6099 , DATAO_REG_6_ , U3422 );
nand NAND2_3090 ( U6100 , U4043 , U3068 );
nand NAND2_3091 ( U6101 , DATAO_REG_7_ , U3422 );
nand NAND2_3092 ( U6102 , U4043 , U3067 );
nand NAND2_3093 ( U6103 , DATAO_REG_8_ , U3422 );
nand NAND2_3094 ( U6104 , U4043 , U3081 );
nand NAND2_3095 ( U6105 , DATAO_REG_9_ , U3422 );
nand NAND2_3096 ( U6106 , U4043 , U3080 );
nand NAND2_3097 ( U6107 , DATAO_REG_10_ , U3422 );
nand NAND2_3098 ( U6108 , U4043 , U3059 );
nand NAND2_3099 ( U6109 , DATAO_REG_11_ , U3422 );
nand NAND2_3100 ( U6110 , U4043 , U3060 );
nand NAND2_3101 ( U6111 , DATAO_REG_12_ , U3422 );
nand NAND2_3102 ( U6112 , U4043 , U3069 );
nand NAND2_3103 ( U6113 , DATAO_REG_13_ , U3422 );
nand NAND2_3104 ( U6114 , U4043 , U3077 );
nand NAND2_3105 ( U6115 , DATAO_REG_14_ , U3422 );
nand NAND2_3106 ( U6116 , U4043 , U3076 );
nand NAND2_3107 ( U6117 , DATAO_REG_15_ , U3422 );
nand NAND2_3108 ( U6118 , U4043 , U3071 );
nand NAND2_3109 ( U6119 , DATAO_REG_16_ , U3422 );
nand NAND2_3110 ( U6120 , U4043 , U3070 );
nand NAND2_3111 ( U6121 , DATAO_REG_17_ , U3422 );
nand NAND2_3112 ( U6122 , U4043 , U3066 );
nand NAND2_3113 ( U6123 , DATAO_REG_18_ , U3422 );
nand NAND2_3114 ( U6124 , U4043 , U3079 );
nand NAND2_3115 ( U6125 , DATAO_REG_19_ , U3422 );
nand NAND2_3116 ( U6126 , U4043 , U3078 );
nand NAND2_3117 ( U6127 , DATAO_REG_20_ , U3422 );
nand NAND2_3118 ( U6128 , U4043 , U3073 );
nand NAND2_3119 ( U6129 , DATAO_REG_21_ , U3422 );
nand NAND2_3120 ( U6130 , U4043 , U3072 );
nand NAND2_3121 ( U6131 , DATAO_REG_22_ , U3422 );
nand NAND2_3122 ( U6132 , U4043 , U3058 );
nand NAND2_3123 ( U6133 , DATAO_REG_23_ , U3422 );
nand NAND2_3124 ( U6134 , U4043 , U3063 );
nand NAND2_3125 ( U6135 , DATAO_REG_24_ , U3422 );
nand NAND2_3126 ( U6136 , U4043 , U3062 );
nand NAND2_3127 ( U6137 , DATAO_REG_25_ , U3422 );
nand NAND2_3128 ( U6138 , U4043 , U3055 );
nand NAND2_3129 ( U6139 , DATAO_REG_26_ , U3422 );
nand NAND2_3130 ( U6140 , U4043 , U3054 );
nand NAND2_3131 ( U6141 , DATAO_REG_27_ , U3422 );
nand NAND2_3132 ( U6142 , U4043 , U3050 );
nand NAND2_3133 ( U6143 , DATAO_REG_28_ , U3422 );
nand NAND2_3134 ( U6144 , U4043 , U3051 );
nand NAND2_3135 ( U6145 , DATAO_REG_29_ , U3422 );
nand NAND2_3136 ( U6146 , U4043 , U3052 );
nand NAND2_3137 ( U6147 , DATAO_REG_30_ , U3422 );
nand NAND2_3138 ( U6148 , U4043 , U3056 );
nand NAND2_3139 ( U6149 , DATAO_REG_31_ , U3422 );
nand NAND2_3140 ( U6150 , U4043 , U3053 );
nand NAND2_3141 ( U6151 , U4040 , U3052 );
nand NAND2_3142 ( U6152 , U3414 , U4737 );
nand NAND2_3143 ( U6153 , U6152 , U6151 );
nand NAND2_3144 ( U6154 , U4038 , U3053 );
nand NAND2_3145 ( U6155 , U3416 , U4775 );
nand NAND2_3146 ( U6156 , U6155 , U6154 );
nand NAND2_3147 ( U6157 , U4039 , U3056 );
nand NAND2_3148 ( U6158 , U3415 , U4755 );
nand NAND2_3149 ( U6159 , U6158 , U6157 );
nand NAND2_3150 ( U6160 , U4037 , U3073 );
nand NAND2_3151 ( U6161 , U3396 , U4566 );
nand NAND2_3152 ( U6162 , U6161 , U6160 );
nand NAND2_3153 ( U6163 , U5892 , U4395 );
nand NAND2_3154 ( U6164 , U3488 , U3060 );
nand NAND2_3155 ( U6165 , U6164 , U6163 );
nand NAND2_3156 ( U6166 , U5887 , U4376 );
nand NAND2_3157 ( U6167 , U3486 , U3059 );
nand NAND2_3158 ( U6168 , U6167 , U6166 );
nand NAND2_3159 ( U6169 , U5857 , U4262 );
nand NAND2_3160 ( U6170 , U3474 , U3057 );
nand NAND2_3161 ( U6171 , U6170 , U6169 );
nand NAND2_3162 ( U6172 , U5932 , U4547 );
nand NAND2_3163 ( U6173 , U3504 , U3078 );
nand NAND2_3164 ( U6174 , U6173 , U6172 );
nand NAND2_3165 ( U6175 , U4032 , U3055 );
nand NAND2_3166 ( U6176 , U3406 , U4661 );
nand NAND2_3167 ( U6177 , U6176 , U6175 );
nand NAND2_3168 ( U6178 , U4031 , U3054 );
nand NAND2_3169 ( U6179 , U3408 , U4680 );
nand NAND2_3170 ( U6180 , U6179 , U6178 );
nand NAND2_3171 ( U6181 , U4036 , U3072 );
nand NAND2_3172 ( U6182 , U3398 , U4585 );
nand NAND2_3173 ( U6183 , U6182 , U6181 );
nand NAND2_3174 ( U6184 , U4035 , U3058 );
nand NAND2_3175 ( U6185 , U3400 , U4604 );
nand NAND2_3176 ( U6186 , U6185 , U6184 );
nand NAND2_3177 ( U6187 , U4034 , U3063 );
nand NAND2_3178 ( U6188 , U3402 , U4623 );
nand NAND2_3179 ( U6189 , U6188 , U6187 );
nand NAND2_3180 ( U6190 , U4033 , U3062 );
nand NAND2_3181 ( U6191 , U3404 , U4642 );
nand NAND2_3182 ( U6192 , U6191 , U6190 );
nand NAND2_3183 ( U6193 , U4030 , U3050 );
nand NAND2_3184 ( U6194 , U3410 , U4699 );
nand NAND2_3185 ( U6195 , U6194 , U6193 );
nand NAND2_3186 ( U6196 , U4029 , U3051 );
nand NAND2_3187 ( U6197 , U3412 , U4718 );
nand NAND2_3188 ( U6198 , U6197 , U6196 );
nand NAND2_3189 ( U6199 , U5877 , U4338 );
nand NAND2_3190 ( U6200 , U3482 , U3081 );
nand NAND2_3191 ( U6201 , U6200 , U6199 );
nand NAND2_3192 ( U6202 , U5882 , U4357 );
nand NAND2_3193 ( U6203 , U3484 , U3080 );
nand NAND2_3194 ( U6204 , U6203 , U6202 );
nand NAND2_3195 ( U6205 , U5927 , U4528 );
nand NAND2_3196 ( U6206 , U3502 , U3079 );
nand NAND2_3197 ( U6207 , U6206 , U6205 );
nand NAND2_3198 ( U6208 , U5902 , U4433 );
nand NAND2_3199 ( U6209 , U3492 , U3077 );
nand NAND2_3200 ( U6210 , U6209 , U6208 );
nand NAND2_3201 ( U6211 , U5907 , U4452 );
nand NAND2_3202 ( U6212 , U3494 , U3076 );
nand NAND2_3203 ( U6213 , U6212 , U6211 );
nand NAND2_3204 ( U6214 , U5842 , U4200 );
nand NAND2_3205 ( U6215 , U3468 , U3075 );
nand NAND2_3206 ( U6216 , U6215 , U6214 );
nand NAND2_3207 ( U6217 , U5829 , U4224 );
nand NAND2_3208 ( U6218 , U3464 , U3074 );
nand NAND2_3209 ( U6219 , U6218 , U6217 );
nand NAND2_3210 ( U6220 , U5912 , U4471 );
nand NAND2_3211 ( U6221 , U3496 , U3071 );
nand NAND2_3212 ( U6222 , U6221 , U6220 );
nand NAND2_3213 ( U6223 , U5917 , U4490 );
nand NAND2_3214 ( U6224 , U3498 , U3070 );
nand NAND2_3215 ( U6225 , U6224 , U6223 );
nand NAND2_3216 ( U6226 , U5897 , U4414 );
nand NAND2_3217 ( U6227 , U3490 , U3069 );
nand NAND2_3218 ( U6228 , U6227 , U6226 );
nand NAND2_3219 ( U6229 , U5867 , U4300 );
nand NAND2_3220 ( U6230 , U3478 , U3068 );
nand NAND2_3221 ( U6231 , U6230 , U6229 );
nand NAND2_3222 ( U6232 , U5872 , U4319 );
nand NAND2_3223 ( U6233 , U3480 , U3067 );
nand NAND2_3224 ( U6234 , U6233 , U6232 );
nand NAND2_3225 ( U6235 , U5922 , U4509 );
nand NAND2_3226 ( U6236 , U3500 , U3066 );
nand NAND2_3227 ( U6237 , U6236 , U6235 );
nand NAND2_3228 ( U6238 , U5847 , U4219 );
nand NAND2_3229 ( U6239 , U3470 , U3065 );
nand NAND2_3230 ( U6240 , U6239 , U6238 );
nand NAND2_3231 ( U6241 , U5862 , U4281 );
nand NAND2_3232 ( U6242 , U3476 , U3064 );
nand NAND2_3233 ( U6243 , U6242 , U6241 );
nand NAND2_3234 ( U6244 , U5852 , U4243 );
nand NAND2_3235 ( U6245 , U3472 , U3061 );
nand NAND2_3236 ( U6246 , U6245 , U6244 );
nand NAND2_3237 ( U6247 , U4042 , U3424 );
nand NAND2_3238 ( U6248 , R1375_U26 , U3373 );
nand NAND2_3239 ( U6249 , U6248 , U6247 );
nand NAND2_3240 ( U6250 , U6249 , U5820 );
nand NAND3_3241 ( U6251 , R395_U6 , U4042 , U3460 );
nand NAND2_3242 ( U6252 , U5817 , U5139 );
nand NAND3_3243 ( U6253 , U4055 , U3425 , U3461 );
nand NAND2_3244 ( U6254 , U4014 , U4007 );
nand NAND2_3245 ( U6255 , U4023 , R1347_U13 );
nand NAND2_3246 ( U6256 , U5748 , U3423 );
nand NAND2_3247 ( U6257 , U3456 , U3431 );
nand NAND2_3248 ( U6258 , U3453 , U5421 );
nand NAND3_3249 ( U6259 , U3016 , REG2_REG_0_ , U5796 );
nand NAND2_3250 ( U6260 , U3080 , R1352_U6 );
nand NAND2_3251 ( U6261 , U3080 , U4009 );
nand NAND2_3252 ( U6262 , U3081 , R1352_U6 );
nand NAND2_3253 ( U6263 , U3081 , U4009 );
nand NAND2_3254 ( U6264 , U3067 , R1352_U6 );
nand NAND2_3255 ( U6265 , U3067 , U4009 );
nand NAND2_3256 ( U6266 , U3068 , R1352_U6 );
nand NAND2_3257 ( U6267 , U3068 , U4009 );
nand NAND2_3258 ( U6268 , U3064 , R1352_U6 );
nand NAND2_3259 ( U6269 , U3064 , U4009 );
nand NAND2_3260 ( U6270 , U3057 , R1352_U6 );
nand NAND2_3261 ( U6271 , U3057 , U4009 );
nand NAND2_3262 ( U6272 , R1309_U8 , R1352_U6 );
nand NAND2_3263 ( U6273 , U3053 , U4009 );
nand NAND2_3264 ( U6274 , R1309_U6 , R1352_U6 );
nand NAND2_3265 ( U6275 , U3056 , U4009 );
nand NAND2_3266 ( U6276 , U3061 , R1352_U6 );
nand NAND2_3267 ( U6277 , U3061 , U4009 );
nand NAND2_3268 ( U6278 , U3052 , R1352_U6 );
nand NAND2_3269 ( U6279 , U3052 , U4009 );
nand NAND2_3270 ( U6280 , U3051 , R1352_U6 );
nand NAND2_3271 ( U6281 , U3051 , U4009 );
nand NAND2_3272 ( U6282 , U3050 , R1352_U6 );
nand NAND2_3273 ( U6283 , U3050 , U4009 );
nand NAND2_3274 ( U6284 , U3054 , R1352_U6 );
nand NAND2_3275 ( U6285 , U3054 , U4009 );
nand NAND2_3276 ( U6286 , U3055 , R1352_U6 );
nand NAND2_3277 ( U6287 , U3055 , U4009 );
nand NAND2_3278 ( U6288 , U3062 , R1352_U6 );
nand NAND2_3279 ( U6289 , U3062 , U4009 );
nand NAND2_3280 ( U6290 , U3063 , R1352_U6 );
nand NAND2_3281 ( U6291 , U3063 , U4009 );
nand NAND2_3282 ( U6292 , U3058 , R1352_U6 );
nand NAND2_3283 ( U6293 , U3058 , U4009 );
nand NAND2_3284 ( U6294 , U3072 , R1352_U6 );
nand NAND2_3285 ( U6295 , U3072 , U4009 );
nand NAND2_3286 ( U6296 , U3073 , R1352_U6 );
nand NAND2_3287 ( U6297 , U3073 , U4009 );
nand NAND2_3288 ( U6298 , U3065 , R1352_U6 );
nand NAND2_3289 ( U6299 , U3065 , U4009 );
nand NAND2_3290 ( U6300 , U3078 , R1352_U6 );
nand NAND2_3291 ( U6301 , U3078 , U4009 );
nand NAND2_3292 ( U6302 , U3079 , R1352_U6 );
nand NAND2_3293 ( U6303 , U3079 , U4009 );
nand NAND2_3294 ( U6304 , U3066 , R1352_U6 );
nand NAND2_3295 ( U6305 , U3066 , U4009 );
nand NAND2_3296 ( U6306 , U3070 , R1352_U6 );
nand NAND2_3297 ( U6307 , U3070 , U4009 );
nand NAND2_3298 ( U6308 , U3071 , R1352_U6 );
nand NAND2_3299 ( U6309 , U3071 , U4009 );
nand NAND2_3300 ( U6310 , U3076 , R1352_U6 );
nand NAND2_3301 ( U6311 , U3076 , U4009 );
nand NAND2_3302 ( U6312 , U3077 , R1352_U6 );
nand NAND2_3303 ( U6313 , U3077 , U4009 );
nand NAND2_3304 ( U6314 , U3069 , R1352_U6 );
nand NAND2_3305 ( U6315 , U3069 , U4009 );
nand NAND2_3306 ( U6316 , U3060 , R1352_U6 );
nand NAND2_3307 ( U6317 , U3060 , U4009 );
nand NAND2_3308 ( U6318 , U3059 , R1352_U6 );
nand NAND2_3309 ( U6319 , U3059 , U4009 );
nand NAND2_3310 ( U6320 , U3075 , R1352_U6 );
nand NAND2_3311 ( U6321 , U3075 , U4009 );
nand NAND2_3312 ( U6322 , U3074 , R1352_U6 );
nand NAND2_3313 ( U6323 , U3074 , U4009 );
nand NAND2_3314 ( R1222_U516 , U3059 , R1222_U70 );
nand NAND2_3315 ( R1222_U515 , R1222_U378 , R1222_U513 );
nand NAND2_3316 ( R1222_U514 , R1222_U179 , R1222_U359 );
nand NAND2_3317 ( R1222_U513 , R1222_U512 , R1222_U511 );
nand NAND2_3318 ( R1222_U512 , U3488 , R1222_U75 );
nand NAND2_3319 ( R1222_U511 , U3060 , R1222_U74 );
nand NAND2_3320 ( R1222_U510 , R1222_U508 , R1222_U334 );
nand NAND2_3321 ( R1222_U509 , R1222_U358 , R1222_U102 );
nand NAND2_3322 ( R1222_U508 , R1222_U507 , R1222_U506 );
nand NAND2_3323 ( R1222_U507 , U3490 , R1222_U73 );
nand NAND2_3324 ( R1222_U506 , U3069 , R1222_U72 );
nand NAND2_3325 ( R1222_U505 , U3492 , R1222_U78 );
nand NAND2_3326 ( R1222_U504 , U3077 , R1222_U77 );
nand NAND2_3327 ( R1222_U503 , R1222_U254 , R1222_U501 );
nand NAND2_3328 ( R1222_U502 , R1222_U177 , R1222_U178 );
nand NAND2_3329 ( R1222_U501 , R1222_U500 , R1222_U499 );
nand NAND2_3330 ( R1222_U500 , U3494 , R1222_U80 );
nand NAND2_3331 ( R1222_U499 , U3076 , R1222_U79 );
nand NAND2_3332 ( R1222_U498 , U3494 , R1222_U80 );
nand NAND2_3333 ( R1222_U497 , U3076 , R1222_U79 );
nand NAND2_3334 ( R1222_U496 , R1222_U257 , R1222_U494 );
nand NAND2_3335 ( R1222_U495 , R1222_U175 , R1222_U176 );
nor nor_3336 ( SUB_84_U4 , IR_REG_26_ , IR_REG_27_ , IR_REG_24_ , IR_REG_25_ );
and AND2_3337 ( SUB_84_U5 , SUB_84_U55 , SUB_84_U54 );
and AND2_3338 ( SUB_84_U6 , SUB_84_U138 , SUB_84_U103 );
and AND2_3339 ( SUB_84_U7 , SUB_84_U137 , SUB_84_U46 );
and AND2_3340 ( SUB_84_U8 , SUB_84_U136 , SUB_84_U32 );
and AND2_3341 ( SUB_84_U9 , SUB_84_U134 , SUB_84_U106 );
and AND2_3342 ( SUB_84_U10 , SUB_84_U133 , SUB_84_U43 );
and AND2_3343 ( SUB_84_U11 , SUB_84_U132 , SUB_84_U38 );
and AND2_3344 ( SUB_84_U12 , SUB_84_U130 , SUB_84_U122 );
and AND2_3345 ( SUB_84_U13 , SUB_84_U129 , SUB_84_U39 );
and AND2_3346 ( SUB_84_U14 , SUB_84_U128 , SUB_84_U40 );
and AND2_3347 ( SUB_84_U15 , SUB_84_U126 , SUB_84_U80 );
and AND2_3348 ( SUB_84_U16 , SUB_84_U120 , SUB_84_U36 );
and AND2_3349 ( SUB_84_U17 , SUB_84_U118 , SUB_84_U75 );
and AND2_3350 ( SUB_84_U18 , SUB_84_U115 , SUB_84_U109 );
and AND2_3351 ( SUB_84_U19 , SUB_84_U113 , SUB_84_U33 );
and AND2_3352 ( SUB_84_U20 , SUB_84_U112 , SUB_84_U29 );
and AND2_3353 ( SUB_84_U21 , SUB_84_U102 , SUB_84_U30 );
and AND2_3354 ( SUB_84_U22 , SUB_84_U101 , SUB_84_U26 );
and AND2_3355 ( SUB_84_U23 , SUB_84_U99 , SUB_84_U93 );
and AND2_3356 ( SUB_84_U24 , SUB_84_U98 , SUB_84_U27 );
and AND2_3357 ( SUB_84_U25 , SUB_84_U97 , SUB_84_U45 );
nand NAND2_3358 ( SUB_84_U26 , SUB_84_U51 , SUB_84_U50 );
nand NAND2_3359 ( SUB_84_U27 , SUB_84_U53 , SUB_84_U92 );
not NOT1_3360 ( SUB_84_U28 , IR_REG_6_ );
or OR3_3361 ( SUB_84_U29 , IR_REG_1_ , IR_REG_0_ , IR_REG_2_ );
nand NAND2_3362 ( SUB_84_U30 , SUB_84_U90 , SUB_84_U31 );
not NOT1_3363 ( SUB_84_U31 , IR_REG_3_ );
nand NAND4_3364 ( SUB_84_U32 , SUB_84_U59 , SUB_84_U58 , SUB_84_U57 , SUB_84_U56 );
nand NAND4_3365 ( SUB_84_U33 , SUB_84_U105 , SUB_84_U4 , SUB_84_U60 , SUB_84_U5 );
nand NAND2_3366 ( SUB_84_U34 , SUB_84_U105 , SUB_84_U5 );
not NOT1_3367 ( SUB_84_U35 , IR_REG_28_ );
nand NAND2_3368 ( SUB_84_U36 , SUB_84_U61 , SUB_84_U108 );
not NOT1_3369 ( SUB_84_U37 , IR_REG_26_ );
nand NAND2_3370 ( SUB_84_U38 , SUB_84_U62 , SUB_84_U105 );
nand NAND2_3371 ( SUB_84_U39 , SUB_84_U63 , SUB_84_U121 );
nand NAND2_3372 ( SUB_84_U40 , SUB_84_U64 , SUB_84_U123 );
not NOT1_3373 ( SUB_84_U41 , IR_REG_22_ );
not NOT1_3374 ( SUB_84_U42 , IR_REG_18_ );
nand NAND2_3375 ( SUB_84_U43 , SUB_84_U65 , SUB_84_U105 );
not NOT1_3376 ( SUB_84_U44 , IR_REG_14_ );
nand NAND2_3377 ( SUB_84_U45 , SUB_84_U52 , SUB_84_U92 );
nand NAND2_3378 ( SUB_84_U46 , SUB_84_U66 , SUB_84_U95 );
not NOT1_3379 ( SUB_84_U47 , IR_REG_10_ );
nand NAND2_3380 ( SUB_84_U48 , SUB_84_U157 , SUB_84_U156 );
nand NAND2_3381 ( SUB_84_U49 , SUB_84_U145 , SUB_84_U144 );
nor nor_3382 ( SUB_84_U50 , IR_REG_2_ , IR_REG_1_ , IR_REG_0_ );
nor nor_3383 ( SUB_84_U51 , IR_REG_5_ , IR_REG_3_ , IR_REG_4_ );
nor nor_3384 ( SUB_84_U52 , IR_REG_6_ , IR_REG_7_ , IR_REG_8_ , IR_REG_9_ );
nor nor_3385 ( SUB_84_U53 , IR_REG_6_ , IR_REG_7_ );
nor nor_3386 ( SUB_84_U54 , IR_REG_17_ , IR_REG_18_ , IR_REG_16_ , IR_REG_14_ , IR_REG_15_ );
nor nor_3387 ( SUB_84_U55 , IR_REG_22_ , IR_REG_23_ , IR_REG_21_ , IR_REG_19_ , IR_REG_20_ );
nor nor_3388 ( SUB_84_U56 , IR_REG_10_ , IR_REG_11_ , IR_REG_12_ , IR_REG_13_ );
nor nor_3389 ( SUB_84_U57 , IR_REG_2_ , IR_REG_1_ , IR_REG_0_ );
nor nor_3390 ( SUB_84_U58 , IR_REG_3_ , IR_REG_4_ , IR_REG_5_ , IR_REG_6_ );
nor nor_3391 ( SUB_84_U59 , IR_REG_9_ , IR_REG_7_ , IR_REG_8_ );
nor nor_3392 ( SUB_84_U60 , IR_REG_28_ , IR_REG_29_ );
nor nor_3393 ( SUB_84_U61 , IR_REG_24_ , IR_REG_25_ );
nor nor_3394 ( SUB_84_U62 , IR_REG_14_ , IR_REG_15_ , IR_REG_16_ , IR_REG_17_ );
nor nor_3395 ( SUB_84_U63 , IR_REG_18_ , IR_REG_19_ );
nor nor_3396 ( SUB_84_U64 , IR_REG_20_ , IR_REG_21_ );
nor nor_3397 ( SUB_84_U65 , IR_REG_14_ , IR_REG_15_ );
nor nor_3398 ( SUB_84_U66 , IR_REG_10_ , IR_REG_11_ );
not NOT1_3399 ( SUB_84_U67 , IR_REG_8_ );
and AND2_3400 ( SUB_84_U68 , SUB_84_U141 , SUB_84_U140 );
not NOT1_3401 ( SUB_84_U69 , IR_REG_4_ );
and AND2_3402 ( SUB_84_U70 , SUB_84_U143 , SUB_84_U142 );
not NOT1_3403 ( SUB_84_U71 , IR_REG_31_ );
not NOT1_3404 ( SUB_84_U72 , IR_REG_30_ );
and AND2_3405 ( SUB_84_U73 , SUB_84_U147 , SUB_84_U146 );
not NOT1_3406 ( SUB_84_U74 , IR_REG_27_ );
nand NAND2_3407 ( SUB_84_U75 , SUB_84_U116 , SUB_84_U37 );
and AND2_3408 ( SUB_84_U76 , SUB_84_U149 , SUB_84_U148 );
not NOT1_3409 ( SUB_84_U77 , IR_REG_24_ );
and AND2_3410 ( SUB_84_U78 , SUB_84_U151 , SUB_84_U150 );
not NOT1_3411 ( SUB_84_U79 , IR_REG_23_ );
nand NAND2_3412 ( SUB_84_U80 , SUB_84_U124 , SUB_84_U41 );
and AND2_3413 ( SUB_84_U81 , SUB_84_U153 , SUB_84_U152 );
not NOT1_3414 ( SUB_84_U82 , IR_REG_20_ );
and AND2_3415 ( SUB_84_U83 , SUB_84_U155 , SUB_84_U154 );
not NOT1_3416 ( SUB_84_U84 , IR_REG_1_ );
not NOT1_3417 ( SUB_84_U85 , IR_REG_0_ );
not NOT1_3418 ( SUB_84_U86 , IR_REG_16_ );
and AND2_3419 ( SUB_84_U87 , SUB_84_U159 , SUB_84_U158 );
not NOT1_3420 ( SUB_84_U88 , IR_REG_12_ );
and AND2_3421 ( SUB_84_U89 , SUB_84_U161 , SUB_84_U160 );
not NOT1_3422 ( SUB_84_U90 , SUB_84_U29 );
not NOT1_3423 ( SUB_84_U91 , SUB_84_U30 );
not NOT1_3424 ( SUB_84_U92 , SUB_84_U26 );
nand NAND2_3425 ( SUB_84_U93 , SUB_84_U92 , SUB_84_U28 );
not NOT1_3426 ( SUB_84_U94 , SUB_84_U27 );
not NOT1_3427 ( SUB_84_U95 , SUB_84_U45 );
nand NAND2_3428 ( SUB_84_U96 , SUB_84_U94 , SUB_84_U67 );
nand NAND2_3429 ( SUB_84_U97 , IR_REG_9_ , SUB_84_U96 );
nand NAND2_3430 ( SUB_84_U98 , IR_REG_7_ , SUB_84_U93 );
nand NAND2_3431 ( SUB_84_U99 , IR_REG_6_ , SUB_84_U26 );
nand NAND2_3432 ( SUB_84_U100 , SUB_84_U91 , SUB_84_U69 );
nand NAND2_3433 ( SUB_84_U101 , IR_REG_5_ , SUB_84_U100 );
nand NAND2_3434 ( SUB_84_U102 , IR_REG_3_ , SUB_84_U29 );
nand NAND2_3435 ( SUB_84_U103 , SUB_84_U95 , SUB_84_U47 );
not NOT1_3436 ( SUB_84_U104 , SUB_84_U46 );
not NOT1_3437 ( SUB_84_U105 , SUB_84_U32 );
nand NAND2_3438 ( SUB_84_U106 , SUB_84_U105 , SUB_84_U44 );
not NOT1_3439 ( SUB_84_U107 , SUB_84_U43 );
not NOT1_3440 ( SUB_84_U108 , SUB_84_U34 );
nand NAND4_3441 ( SUB_84_U109 , SUB_84_U105 , SUB_84_U4 , SUB_84_U5 , SUB_84_U35 );
not NOT1_3442 ( SUB_84_U110 , SUB_84_U33 );
or OR2_3443 ( SUB_84_U111 , IR_REG_1_ , IR_REG_0_ );
nand NAND2_3444 ( SUB_84_U112 , IR_REG_2_ , SUB_84_U111 );
nand NAND2_3445 ( SUB_84_U113 , IR_REG_29_ , SUB_84_U109 );
nand NAND2_3446 ( SUB_84_U114 , SUB_84_U108 , SUB_84_U4 );
nand NAND2_3447 ( SUB_84_U115 , IR_REG_28_ , SUB_84_U114 );
not NOT1_3448 ( SUB_84_U116 , SUB_84_U36 );
not NOT1_3449 ( SUB_84_U117 , SUB_84_U75 );
nand NAND2_3450 ( SUB_84_U118 , IR_REG_26_ , SUB_84_U36 );
nand NAND2_3451 ( SUB_84_U119 , SUB_84_U108 , SUB_84_U77 );
nand NAND2_3452 ( SUB_84_U120 , IR_REG_25_ , SUB_84_U119 );
not NOT1_3453 ( SUB_84_U121 , SUB_84_U38 );
nand NAND2_3454 ( SUB_84_U122 , SUB_84_U121 , SUB_84_U42 );
not NOT1_3455 ( SUB_84_U123 , SUB_84_U39 );
not NOT1_3456 ( SUB_84_U124 , SUB_84_U40 );
not NOT1_3457 ( SUB_84_U125 , SUB_84_U80 );
nand NAND2_3458 ( SUB_84_U126 , IR_REG_22_ , SUB_84_U40 );
nand NAND2_3459 ( SUB_84_U127 , SUB_84_U123 , SUB_84_U82 );
nand NAND2_3460 ( SUB_84_U128 , IR_REG_21_ , SUB_84_U127 );
nand NAND2_3461 ( SUB_84_U129 , IR_REG_19_ , SUB_84_U122 );
nand NAND2_3462 ( SUB_84_U130 , IR_REG_18_ , SUB_84_U38 );
nand NAND2_3463 ( SUB_84_U131 , SUB_84_U107 , SUB_84_U86 );
nand NAND2_3464 ( SUB_84_U132 , IR_REG_17_ , SUB_84_U131 );
nand NAND2_3465 ( SUB_84_U133 , IR_REG_15_ , SUB_84_U106 );
nand NAND2_3466 ( SUB_84_U134 , IR_REG_14_ , SUB_84_U32 );
nand NAND2_3467 ( SUB_84_U135 , SUB_84_U104 , SUB_84_U88 );
nand NAND2_3468 ( SUB_84_U136 , IR_REG_13_ , SUB_84_U135 );
nand NAND2_3469 ( SUB_84_U137 , IR_REG_11_ , SUB_84_U103 );
nand NAND2_3470 ( SUB_84_U138 , IR_REG_10_ , SUB_84_U45 );
nand NAND2_3471 ( SUB_84_U139 , SUB_84_U110 , SUB_84_U72 );
nand NAND2_3472 ( SUB_84_U140 , IR_REG_8_ , SUB_84_U27 );
nand NAND2_3473 ( SUB_84_U141 , SUB_84_U94 , SUB_84_U67 );
nand NAND2_3474 ( SUB_84_U142 , IR_REG_4_ , SUB_84_U30 );
nand NAND2_3475 ( SUB_84_U143 , SUB_84_U91 , SUB_84_U69 );
nand NAND2_3476 ( SUB_84_U144 , SUB_84_U139 , SUB_84_U71 );
nand NAND3_3477 ( SUB_84_U145 , SUB_84_U110 , SUB_84_U72 , IR_REG_31_ );
nand NAND2_3478 ( SUB_84_U146 , IR_REG_30_ , SUB_84_U33 );
nand NAND2_3479 ( SUB_84_U147 , SUB_84_U110 , SUB_84_U72 );
nand NAND2_3480 ( SUB_84_U148 , IR_REG_27_ , SUB_84_U75 );
nand NAND2_3481 ( SUB_84_U149 , SUB_84_U117 , SUB_84_U74 );
nand NAND2_3482 ( SUB_84_U150 , IR_REG_24_ , SUB_84_U34 );
nand NAND2_3483 ( SUB_84_U151 , SUB_84_U108 , SUB_84_U77 );
nand NAND2_3484 ( SUB_84_U152 , IR_REG_23_ , SUB_84_U80 );
nand NAND2_3485 ( SUB_84_U153 , SUB_84_U125 , SUB_84_U79 );
nand NAND2_3486 ( SUB_84_U154 , IR_REG_20_ , SUB_84_U39 );
nand NAND2_3487 ( SUB_84_U155 , SUB_84_U123 , SUB_84_U82 );
nand NAND2_3488 ( SUB_84_U156 , IR_REG_1_ , SUB_84_U85 );
nand NAND2_3489 ( SUB_84_U157 , IR_REG_0_ , SUB_84_U84 );
nand NAND2_3490 ( SUB_84_U158 , IR_REG_16_ , SUB_84_U43 );
nand NAND2_3491 ( SUB_84_U159 , SUB_84_U107 , SUB_84_U86 );
nand NAND2_3492 ( SUB_84_U160 , IR_REG_12_ , SUB_84_U46 );
nand NAND2_3493 ( SUB_84_U161 , SUB_84_U104 , SUB_84_U88 );
not NOT1_3494 ( ADD_95_U4 , REG3_REG_3_ );
and AND2_3495 ( ADD_95_U5 , ADD_95_U76 , ADD_95_U107 );
not NOT1_3496 ( ADD_95_U6 , REG3_REG_7_ );
not NOT1_3497 ( ADD_95_U7 , REG3_REG_6_ );
not NOT1_3498 ( ADD_95_U8 , REG3_REG_5_ );
not NOT1_3499 ( ADD_95_U9 , REG3_REG_4_ );
nand NAND5_3500 ( ADD_95_U10 , REG3_REG_7_ , REG3_REG_3_ , REG3_REG_6_ , REG3_REG_4_ , REG3_REG_5_ );
not NOT1_3501 ( ADD_95_U11 , REG3_REG_8_ );
not NOT1_3502 ( ADD_95_U12 , REG3_REG_9_ );
nand NAND2_3503 ( ADD_95_U13 , ADD_95_U71 , ADD_95_U88 );
not NOT1_3504 ( ADD_95_U14 , REG3_REG_11_ );
not NOT1_3505 ( ADD_95_U15 , REG3_REG_10_ );
nand NAND2_3506 ( ADD_95_U16 , ADD_95_U72 , ADD_95_U90 );
not NOT1_3507 ( ADD_95_U17 , REG3_REG_13_ );
not NOT1_3508 ( ADD_95_U18 , REG3_REG_12_ );
nand NAND2_3509 ( ADD_95_U19 , ADD_95_U73 , ADD_95_U92 );
not NOT1_3510 ( ADD_95_U20 , REG3_REG_15_ );
not NOT1_3511 ( ADD_95_U21 , REG3_REG_14_ );
nand NAND2_3512 ( ADD_95_U22 , ADD_95_U74 , ADD_95_U94 );
not NOT1_3513 ( ADD_95_U23 , REG3_REG_17_ );
not NOT1_3514 ( ADD_95_U24 , REG3_REG_16_ );
nand NAND2_3515 ( ADD_95_U25 , ADD_95_U75 , ADD_95_U96 );
not NOT1_3516 ( ADD_95_U26 , REG3_REG_18_ );
nand NAND2_3517 ( ADD_95_U27 , REG3_REG_18_ , ADD_95_U98 );
not NOT1_3518 ( ADD_95_U28 , REG3_REG_19_ );
nand NAND2_3519 ( ADD_95_U29 , REG3_REG_19_ , ADD_95_U99 );
not NOT1_3520 ( ADD_95_U30 , REG3_REG_20_ );
nand NAND2_3521 ( ADD_95_U31 , REG3_REG_20_ , ADD_95_U100 );
not NOT1_3522 ( ADD_95_U32 , REG3_REG_21_ );
nand NAND2_3523 ( ADD_95_U33 , REG3_REG_21_ , ADD_95_U101 );
not NOT1_3524 ( ADD_95_U34 , REG3_REG_22_ );
nand NAND2_3525 ( ADD_95_U35 , REG3_REG_22_ , ADD_95_U102 );
not NOT1_3526 ( ADD_95_U36 , REG3_REG_23_ );
nand NAND2_3527 ( ADD_95_U37 , REG3_REG_23_ , ADD_95_U103 );
not NOT1_3528 ( ADD_95_U38 , REG3_REG_24_ );
nand NAND2_3529 ( ADD_95_U39 , REG3_REG_24_ , ADD_95_U104 );
not NOT1_3530 ( ADD_95_U40 , REG3_REG_25_ );
nand NAND2_3531 ( ADD_95_U41 , REG3_REG_25_ , ADD_95_U105 );
not NOT1_3532 ( ADD_95_U42 , REG3_REG_26_ );
nand NAND2_3533 ( ADD_95_U43 , REG3_REG_26_ , ADD_95_U106 );
not NOT1_3534 ( ADD_95_U44 , REG3_REG_28_ );
not NOT1_3535 ( ADD_95_U45 , REG3_REG_27_ );
nand NAND2_3536 ( ADD_95_U46 , ADD_95_U111 , ADD_95_U110 );
nand NAND2_3537 ( ADD_95_U47 , ADD_95_U113 , ADD_95_U112 );
nand NAND2_3538 ( ADD_95_U48 , ADD_95_U115 , ADD_95_U114 );
nand NAND2_3539 ( ADD_95_U49 , ADD_95_U117 , ADD_95_U116 );
nand NAND2_3540 ( ADD_95_U50 , ADD_95_U119 , ADD_95_U118 );
nand NAND2_3541 ( ADD_95_U51 , ADD_95_U121 , ADD_95_U120 );
nand NAND2_3542 ( ADD_95_U52 , ADD_95_U123 , ADD_95_U122 );
nand NAND2_3543 ( ADD_95_U53 , ADD_95_U125 , ADD_95_U124 );
nand NAND2_3544 ( ADD_95_U54 , ADD_95_U127 , ADD_95_U126 );
nand NAND2_3545 ( ADD_95_U55 , ADD_95_U129 , ADD_95_U128 );
nand NAND2_3546 ( ADD_95_U56 , ADD_95_U131 , ADD_95_U130 );
nand NAND2_3547 ( ADD_95_U57 , ADD_95_U133 , ADD_95_U132 );
nand NAND2_3548 ( ADD_95_U58 , ADD_95_U135 , ADD_95_U134 );
nand NAND2_3549 ( ADD_95_U59 , ADD_95_U137 , ADD_95_U136 );
nand NAND2_3550 ( ADD_95_U60 , ADD_95_U139 , ADD_95_U138 );
nand NAND2_3551 ( ADD_95_U61 , ADD_95_U141 , ADD_95_U140 );
nand NAND2_3552 ( ADD_95_U62 , ADD_95_U143 , ADD_95_U142 );
nand NAND2_3553 ( ADD_95_U63 , ADD_95_U145 , ADD_95_U144 );
nand NAND2_3554 ( ADD_95_U64 , ADD_95_U147 , ADD_95_U146 );
nand NAND2_3555 ( ADD_95_U65 , ADD_95_U149 , ADD_95_U148 );
nand NAND2_3556 ( ADD_95_U66 , ADD_95_U151 , ADD_95_U150 );
nand NAND2_3557 ( ADD_95_U67 , ADD_95_U153 , ADD_95_U152 );
nand NAND2_3558 ( ADD_95_U68 , ADD_95_U155 , ADD_95_U154 );
nand NAND2_3559 ( ADD_95_U69 , ADD_95_U157 , ADD_95_U156 );
nand NAND2_3560 ( ADD_95_U70 , ADD_95_U159 , ADD_95_U158 );
and AND2_3561 ( ADD_95_U71 , REG3_REG_8_ , REG3_REG_9_ );
and AND2_3562 ( ADD_95_U72 , REG3_REG_11_ , REG3_REG_10_ );
and AND2_3563 ( ADD_95_U73 , REG3_REG_13_ , REG3_REG_12_ );
and AND2_3564 ( ADD_95_U74 , REG3_REG_15_ , REG3_REG_14_ );
and AND2_3565 ( ADD_95_U75 , REG3_REG_17_ , REG3_REG_16_ );
and AND2_3566 ( ADD_95_U76 , REG3_REG_28_ , REG3_REG_27_ );
nand NAND2_3567 ( ADD_95_U77 , REG3_REG_8_ , ADD_95_U88 );
nand NAND4_3568 ( ADD_95_U78 , REG3_REG_4_ , REG3_REG_5_ , REG3_REG_6_ , REG3_REG_3_ );
nand NAND3_3569 ( ADD_95_U79 , REG3_REG_5_ , REG3_REG_3_ , REG3_REG_4_ );
nand NAND2_3570 ( ADD_95_U80 , REG3_REG_4_ , REG3_REG_3_ );
nand NAND2_3571 ( ADD_95_U81 , REG3_REG_27_ , ADD_95_U107 );
nand NAND2_3572 ( ADD_95_U82 , REG3_REG_16_ , ADD_95_U96 );
nand NAND2_3573 ( ADD_95_U83 , REG3_REG_14_ , ADD_95_U94 );
nand NAND2_3574 ( ADD_95_U84 , REG3_REG_12_ , ADD_95_U92 );
nand NAND2_3575 ( ADD_95_U85 , REG3_REG_10_ , ADD_95_U90 );
not NOT1_3576 ( ADD_95_U86 , ADD_95_U80 );
not NOT1_3577 ( ADD_95_U87 , ADD_95_U78 );
not NOT1_3578 ( ADD_95_U88 , ADD_95_U10 );
not NOT1_3579 ( ADD_95_U89 , ADD_95_U77 );
not NOT1_3580 ( ADD_95_U90 , ADD_95_U13 );
not NOT1_3581 ( ADD_95_U91 , ADD_95_U85 );
not NOT1_3582 ( ADD_95_U92 , ADD_95_U16 );
not NOT1_3583 ( ADD_95_U93 , ADD_95_U84 );
not NOT1_3584 ( ADD_95_U94 , ADD_95_U19 );
not NOT1_3585 ( ADD_95_U95 , ADD_95_U83 );
not NOT1_3586 ( ADD_95_U96 , ADD_95_U22 );
not NOT1_3587 ( ADD_95_U97 , ADD_95_U82 );
not NOT1_3588 ( ADD_95_U98 , ADD_95_U25 );
not NOT1_3589 ( ADD_95_U99 , ADD_95_U27 );
not NOT1_3590 ( ADD_95_U100 , ADD_95_U29 );
not NOT1_3591 ( ADD_95_U101 , ADD_95_U31 );
not NOT1_3592 ( ADD_95_U102 , ADD_95_U33 );
not NOT1_3593 ( ADD_95_U103 , ADD_95_U35 );
not NOT1_3594 ( ADD_95_U104 , ADD_95_U37 );
not NOT1_3595 ( ADD_95_U105 , ADD_95_U39 );
not NOT1_3596 ( ADD_95_U106 , ADD_95_U41 );
not NOT1_3597 ( ADD_95_U107 , ADD_95_U43 );
not NOT1_3598 ( ADD_95_U108 , ADD_95_U81 );
not NOT1_3599 ( ADD_95_U109 , ADD_95_U79 );
nand NAND2_3600 ( ADD_95_U110 , REG3_REG_9_ , ADD_95_U77 );
nand NAND2_3601 ( ADD_95_U111 , ADD_95_U89 , ADD_95_U12 );
nand NAND2_3602 ( ADD_95_U112 , REG3_REG_8_ , ADD_95_U10 );
nand NAND2_3603 ( ADD_95_U113 , ADD_95_U88 , ADD_95_U11 );
nand NAND2_3604 ( ADD_95_U114 , REG3_REG_7_ , ADD_95_U78 );
nand NAND2_3605 ( ADD_95_U115 , ADD_95_U87 , ADD_95_U6 );
nand NAND2_3606 ( ADD_95_U116 , REG3_REG_6_ , ADD_95_U79 );
nand NAND2_3607 ( ADD_95_U117 , ADD_95_U109 , ADD_95_U7 );
nand NAND2_3608 ( ADD_95_U118 , REG3_REG_5_ , ADD_95_U80 );
nand NAND2_3609 ( ADD_95_U119 , ADD_95_U86 , ADD_95_U8 );
nand NAND2_3610 ( ADD_95_U120 , REG3_REG_4_ , ADD_95_U4 );
nand NAND2_3611 ( ADD_95_U121 , REG3_REG_3_ , ADD_95_U9 );
nand NAND2_3612 ( ADD_95_U122 , REG3_REG_28_ , ADD_95_U81 );
nand NAND2_3613 ( ADD_95_U123 , ADD_95_U108 , ADD_95_U44 );
nand NAND2_3614 ( ADD_95_U124 , REG3_REG_27_ , ADD_95_U43 );
nand NAND2_3615 ( ADD_95_U125 , ADD_95_U107 , ADD_95_U45 );
nand NAND2_3616 ( ADD_95_U126 , REG3_REG_26_ , ADD_95_U41 );
nand NAND2_3617 ( ADD_95_U127 , ADD_95_U106 , ADD_95_U42 );
nand NAND2_3618 ( ADD_95_U128 , REG3_REG_25_ , ADD_95_U39 );
nand NAND2_3619 ( ADD_95_U129 , ADD_95_U105 , ADD_95_U40 );
nand NAND2_3620 ( ADD_95_U130 , REG3_REG_24_ , ADD_95_U37 );
nand NAND2_3621 ( ADD_95_U131 , ADD_95_U104 , ADD_95_U38 );
nand NAND2_3622 ( ADD_95_U132 , REG3_REG_23_ , ADD_95_U35 );
nand NAND2_3623 ( ADD_95_U133 , ADD_95_U103 , ADD_95_U36 );
nand NAND2_3624 ( ADD_95_U134 , REG3_REG_22_ , ADD_95_U33 );
nand NAND2_3625 ( ADD_95_U135 , ADD_95_U102 , ADD_95_U34 );
nand NAND2_3626 ( ADD_95_U136 , REG3_REG_21_ , ADD_95_U31 );
nand NAND2_3627 ( ADD_95_U137 , ADD_95_U101 , ADD_95_U32 );
nand NAND2_3628 ( ADD_95_U138 , REG3_REG_20_ , ADD_95_U29 );
nand NAND2_3629 ( ADD_95_U139 , ADD_95_U100 , ADD_95_U30 );
nand NAND2_3630 ( ADD_95_U140 , REG3_REG_19_ , ADD_95_U27 );
nand NAND2_3631 ( ADD_95_U141 , ADD_95_U99 , ADD_95_U28 );
nand NAND2_3632 ( ADD_95_U142 , REG3_REG_18_ , ADD_95_U25 );
nand NAND2_3633 ( ADD_95_U143 , ADD_95_U98 , ADD_95_U26 );
nand NAND2_3634 ( ADD_95_U144 , REG3_REG_17_ , ADD_95_U82 );
nand NAND2_3635 ( ADD_95_U145 , ADD_95_U97 , ADD_95_U23 );
nand NAND2_3636 ( ADD_95_U146 , REG3_REG_16_ , ADD_95_U22 );
nand NAND2_3637 ( ADD_95_U147 , ADD_95_U96 , ADD_95_U24 );
nand NAND2_3638 ( ADD_95_U148 , REG3_REG_15_ , ADD_95_U83 );
nand NAND2_3639 ( ADD_95_U149 , ADD_95_U95 , ADD_95_U20 );
nand NAND2_3640 ( ADD_95_U150 , REG3_REG_14_ , ADD_95_U19 );
nand NAND2_3641 ( ADD_95_U151 , ADD_95_U94 , ADD_95_U21 );
nand NAND2_3642 ( ADD_95_U152 , REG3_REG_13_ , ADD_95_U84 );
nand NAND2_3643 ( ADD_95_U153 , ADD_95_U93 , ADD_95_U17 );
nand NAND2_3644 ( ADD_95_U154 , REG3_REG_12_ , ADD_95_U16 );
nand NAND2_3645 ( ADD_95_U155 , ADD_95_U92 , ADD_95_U18 );
nand NAND2_3646 ( ADD_95_U156 , REG3_REG_11_ , ADD_95_U85 );
nand NAND2_3647 ( ADD_95_U157 , ADD_95_U91 , ADD_95_U14 );
nand NAND2_3648 ( ADD_95_U158 , REG3_REG_10_ , ADD_95_U13 );
nand NAND2_3649 ( ADD_95_U159 , ADD_95_U90 , ADD_95_U15 );
nand NAND2_3650 ( R395_U6 , R395_U99 , R395_U183 );
not NOT1_3651 ( R395_U7 , U3111 );
not NOT1_3652 ( R395_U8 , U3110 );
not NOT1_3653 ( R395_U9 , U3109 );
not NOT1_3654 ( R395_U10 , U3143 );
not NOT1_3655 ( R395_U11 , U3142 );
not NOT1_3656 ( R395_U12 , U3141 );
not NOT1_3657 ( R395_U13 , U3140 );
not NOT1_3658 ( R395_U14 , U3139 );
not NOT1_3659 ( R395_U15 , U3138 );
not NOT1_3660 ( R395_U16 , U3108 );
not NOT1_3661 ( R395_U17 , U3107 );
not NOT1_3662 ( R395_U18 , U3106 );
not NOT1_3663 ( R395_U19 , U3105 );
not NOT1_3664 ( R395_U20 , U3104 );
not NOT1_3665 ( R395_U21 , U3103 );
not NOT1_3666 ( R395_U22 , U3137 );
not NOT1_3667 ( R395_U23 , U3136 );
not NOT1_3668 ( R395_U24 , U3135 );
not NOT1_3669 ( R395_U25 , U3134 );
not NOT1_3670 ( R395_U26 , U3133 );
not NOT1_3671 ( R395_U27 , U3132 );
not NOT1_3672 ( R395_U28 , U3102 );
not NOT1_3673 ( R395_U29 , U3101 );
not NOT1_3674 ( R395_U30 , U3100 );
not NOT1_3675 ( R395_U31 , U3099 );
not NOT1_3676 ( R395_U32 , U3131 );
not NOT1_3677 ( R395_U33 , U3130 );
not NOT1_3678 ( R395_U34 , U3098 );
not NOT1_3679 ( R395_U35 , U3097 );
not NOT1_3680 ( R395_U36 , U3129 );
not NOT1_3681 ( R395_U37 , U3128 );
not NOT1_3682 ( R395_U38 , U3096 );
not NOT1_3683 ( R395_U39 , U3095 );
not NOT1_3684 ( R395_U40 , U3127 );
not NOT1_3685 ( R395_U41 , U3126 );
not NOT1_3686 ( R395_U42 , U3094 );
not NOT1_3687 ( R395_U43 , U3093 );
not NOT1_3688 ( R395_U44 , U3125 );
not NOT1_3689 ( R395_U45 , U3124 );
not NOT1_3690 ( R395_U46 , U3092 );
not NOT1_3691 ( R395_U47 , U3091 );
not NOT1_3692 ( R395_U48 , U3123 );
not NOT1_3693 ( R395_U49 , U3122 );
not NOT1_3694 ( R395_U50 , U3090 );
not NOT1_3695 ( R395_U51 , U3089 );
not NOT1_3696 ( R395_U52 , U3121 );
not NOT1_3697 ( R395_U53 , U3120 );
not NOT1_3698 ( R395_U54 , U3088 );
not NOT1_3699 ( R395_U55 , U3087 );
not NOT1_3700 ( R395_U56 , U3119 );
not NOT1_3701 ( R395_U57 , U3118 );
not NOT1_3702 ( R395_U58 , U3086 );
not NOT1_3703 ( R395_U59 , U3085 );
not NOT1_3704 ( R395_U60 , U3117 );
not NOT1_3705 ( R395_U61 , U3116 );
not NOT1_3706 ( R395_U62 , U3084 );
not NOT1_3707 ( R395_U63 , U3083 );
not NOT1_3708 ( R395_U64 , U3115 );
not NOT1_3709 ( R395_U65 , U3114 );
not NOT1_3710 ( R395_U66 , U3146 );
and AND3_3711 ( R395_U67 , R395_U103 , R395_U104 , R395_U102 );
and AND3_3712 ( R395_U68 , R395_U109 , R395_U108 , R395_U184 );
and AND2_3713 ( R395_U69 , U3142 , R395_U8 );
and AND3_3714 ( R395_U70 , R395_U110 , R395_U107 , R395_U106 );
and AND3_3715 ( R395_U71 , R395_U115 , R395_U111 , R395_U116 );
and AND2_3716 ( R395_U72 , U3107 , R395_U14 );
and AND4_3717 ( R395_U73 , R395_U117 , R395_U114 , R395_U113 , R395_U74 );
and AND3_3718 ( R395_U74 , R395_U122 , R395_U118 , R395_U123 );
and AND2_3719 ( R395_U75 , U3136 , R395_U20 );
and AND4_3720 ( R395_U76 , R395_U124 , R395_U121 , R395_U120 , R395_U77 );
and AND3_3721 ( R395_U77 , R395_U129 , R395_U125 , R395_U130 );
and AND2_3722 ( R395_U78 , U3101 , R395_U26 );
and AND3_3723 ( R395_U79 , R395_U80 , R395_U128 , R395_U127 );
and AND2_3724 ( R395_U80 , R395_U132 , R395_U131 );
and AND2_3725 ( R395_U81 , R395_U134 , R395_U135 );
and AND2_3726 ( R395_U82 , R395_U137 , R395_U138 );
and AND2_3727 ( R395_U83 , R395_U140 , R395_U141 );
and AND2_3728 ( R395_U84 , R395_U143 , R395_U144 );
and AND2_3729 ( R395_U85 , R395_U146 , R395_U147 );
and AND2_3730 ( R395_U86 , R395_U149 , R395_U150 );
and AND2_3731 ( R395_U87 , R395_U152 , R395_U153 );
and AND2_3732 ( R395_U88 , R395_U155 , R395_U156 );
and AND2_3733 ( R395_U89 , R395_U158 , R395_U159 );
and AND2_3734 ( R395_U90 , R395_U161 , R395_U162 );
and AND2_3735 ( R395_U91 , R395_U164 , R395_U165 );
and AND2_3736 ( R395_U92 , R395_U167 , R395_U168 );
and AND2_3737 ( R395_U93 , R395_U170 , R395_U171 );
and AND2_3738 ( R395_U94 , R395_U173 , R395_U174 );
and AND2_3739 ( R395_U95 , R395_U176 , R395_U177 );
and AND2_3740 ( R395_U96 , R395_U179 , R395_U180 );
and AND3_3741 ( R395_U97 , R395_U186 , R395_U185 , R395_U182 );
not NOT1_3742 ( R395_U98 , U3082 );
and AND2_3743 ( R395_U99 , R395_U188 , R395_U187 );
not NOT1_3744 ( R395_U100 , U3144 );
not NOT1_3745 ( R395_U101 , U3145 );
nand NAND3_3746 ( R395_U102 , R395_U101 , R395_U100 , U3113 );
nand NAND2_3747 ( R395_U103 , U3112 , R395_U100 );
nand NAND2_3748 ( R395_U104 , U3111 , R395_U10 );
nand NAND2_3749 ( R395_U105 , R395_U68 , R395_U67 );
nand NAND4_3750 ( R395_U106 , U3143 , R395_U109 , R395_U108 , R395_U7 );
nand NAND2_3751 ( R395_U107 , R395_U69 , R395_U109 );
nand NAND2_3752 ( R395_U108 , U3110 , R395_U11 );
nand NAND2_3753 ( R395_U109 , U3109 , R395_U12 );
nand NAND2_3754 ( R395_U110 , U3141 , R395_U9 );
nand NAND2_3755 ( R395_U111 , U3140 , R395_U16 );
nand NAND3_3756 ( R395_U112 , R395_U105 , R395_U71 , R395_U70 );
nand NAND4_3757 ( R395_U113 , U3108 , R395_U116 , R395_U115 , R395_U13 );
nand NAND2_3758 ( R395_U114 , R395_U72 , R395_U116 );
nand NAND2_3759 ( R395_U115 , U3139 , R395_U17 );
nand NAND2_3760 ( R395_U116 , U3138 , R395_U18 );
nand NAND2_3761 ( R395_U117 , U3106 , R395_U15 );
nand NAND2_3762 ( R395_U118 , U3105 , R395_U22 );
nand NAND2_3763 ( R395_U119 , R395_U112 , R395_U73 );
nand NAND4_3764 ( R395_U120 , U3137 , R395_U123 , R395_U122 , R395_U19 );
nand NAND2_3765 ( R395_U121 , R395_U75 , R395_U123 );
nand NAND2_3766 ( R395_U122 , U3104 , R395_U23 );
nand NAND2_3767 ( R395_U123 , U3103 , R395_U24 );
nand NAND2_3768 ( R395_U124 , U3135 , R395_U21 );
nand NAND2_3769 ( R395_U125 , U3134 , R395_U28 );
nand NAND2_3770 ( R395_U126 , R395_U119 , R395_U76 );
nand NAND4_3771 ( R395_U127 , U3102 , R395_U130 , R395_U129 , R395_U25 );
nand NAND2_3772 ( R395_U128 , R395_U78 , R395_U130 );
nand NAND2_3773 ( R395_U129 , U3133 , R395_U29 );
nand NAND2_3774 ( R395_U130 , U3132 , R395_U30 );
nand NAND2_3775 ( R395_U131 , U3100 , R395_U27 );
nand NAND2_3776 ( R395_U132 , U3099 , R395_U32 );
nand NAND2_3777 ( R395_U133 , R395_U126 , R395_U79 );
nand NAND2_3778 ( R395_U134 , U3131 , R395_U31 );
nand NAND2_3779 ( R395_U135 , U3130 , R395_U34 );
nand NAND2_3780 ( R395_U136 , R395_U81 , R395_U133 );
nand NAND2_3781 ( R395_U137 , U3098 , R395_U33 );
nand NAND2_3782 ( R395_U138 , U3097 , R395_U36 );
nand NAND2_3783 ( R395_U139 , R395_U82 , R395_U136 );
nand NAND2_3784 ( R395_U140 , U3129 , R395_U35 );
nand NAND2_3785 ( R395_U141 , U3128 , R395_U38 );
nand NAND2_3786 ( R395_U142 , R395_U83 , R395_U139 );
nand NAND2_3787 ( R395_U143 , U3096 , R395_U37 );
nand NAND2_3788 ( R395_U144 , U3095 , R395_U40 );
nand NAND2_3789 ( R395_U145 , R395_U84 , R395_U142 );
nand NAND2_3790 ( R395_U146 , U3127 , R395_U39 );
nand NAND2_3791 ( R395_U147 , U3126 , R395_U42 );
nand NAND2_3792 ( R395_U148 , R395_U85 , R395_U145 );
nand NAND2_3793 ( R395_U149 , U3094 , R395_U41 );
nand NAND2_3794 ( R395_U150 , U3093 , R395_U44 );
nand NAND2_3795 ( R395_U151 , R395_U86 , R395_U148 );
nand NAND2_3796 ( R395_U152 , U3125 , R395_U43 );
nand NAND2_3797 ( R395_U153 , U3124 , R395_U46 );
nand NAND2_3798 ( R395_U154 , R395_U87 , R395_U151 );
nand NAND2_3799 ( R395_U155 , U3092 , R395_U45 );
nand NAND2_3800 ( R395_U156 , U3091 , R395_U48 );
nand NAND2_3801 ( R395_U157 , R395_U88 , R395_U154 );
nand NAND2_3802 ( R395_U158 , U3123 , R395_U47 );
nand NAND2_3803 ( R395_U159 , U3122 , R395_U50 );
nand NAND2_3804 ( R395_U160 , R395_U89 , R395_U157 );
nand NAND2_3805 ( R395_U161 , U3090 , R395_U49 );
nand NAND2_3806 ( R395_U162 , U3089 , R395_U52 );
nand NAND2_3807 ( R395_U163 , R395_U90 , R395_U160 );
nand NAND2_3808 ( R395_U164 , U3121 , R395_U51 );
nand NAND2_3809 ( R395_U165 , U3120 , R395_U54 );
nand NAND2_3810 ( R395_U166 , R395_U91 , R395_U163 );
nand NAND2_3811 ( R395_U167 , U3088 , R395_U53 );
nand NAND2_3812 ( R395_U168 , U3087 , R395_U56 );
nand NAND2_3813 ( R395_U169 , R395_U92 , R395_U166 );
nand NAND2_3814 ( R395_U170 , U3119 , R395_U55 );
nand NAND2_3815 ( R395_U171 , U3118 , R395_U58 );
nand NAND2_3816 ( R395_U172 , R395_U93 , R395_U169 );
nand NAND2_3817 ( R395_U173 , U3086 , R395_U57 );
nand NAND2_3818 ( R395_U174 , U3085 , R395_U60 );
nand NAND2_3819 ( R395_U175 , R395_U94 , R395_U172 );
nand NAND2_3820 ( R395_U176 , U3117 , R395_U59 );
nand NAND2_3821 ( R395_U177 , U3116 , R395_U62 );
nand NAND2_3822 ( R395_U178 , R395_U95 , R395_U175 );
nand NAND2_3823 ( R395_U179 , U3084 , R395_U61 );
nand NAND2_3824 ( R395_U180 , U3083 , R395_U64 );
nand NAND2_3825 ( R395_U181 , R395_U96 , R395_U178 );
nand NAND2_3826 ( R395_U182 , U3115 , R395_U63 );
nand NAND2_3827 ( R395_U183 , R395_U97 , R395_U181 );
nand NAND3_3828 ( R395_U184 , U3113 , U3112 , R395_U101 );
nand NAND2_3829 ( R395_U185 , U3114 , R395_U98 );
nand NAND2_3830 ( R395_U186 , U3082 , R395_U65 );
nand NAND3_3831 ( R395_U187 , U3146 , U3114 , R395_U98 );
nand NAND3_3832 ( R395_U188 , R395_U66 , R395_U65 , U3082 );
and AND2_3833 ( R1105_U4 , R1105_U179 , R1105_U175 );
nand NAND2_3834 ( R1105_U5 , R1105_U83 , R1105_U180 );
not NOT1_3835 ( R1105_U6 , REG2_REG_0_ );
not NOT1_3836 ( R1105_U7 , U3453 );
not NOT1_3837 ( R1105_U8 , REG2_REG_1_ );
nand NAND2_3838 ( R1105_U9 , U3453 , REG2_REG_0_ );
not NOT1_3839 ( R1105_U10 , U3443 );
not NOT1_3840 ( R1105_U11 , REG2_REG_2_ );
not NOT1_3841 ( R1105_U12 , U3442 );
not NOT1_3842 ( R1105_U13 , REG2_REG_3_ );
not NOT1_3843 ( R1105_U14 , U3441 );
not NOT1_3844 ( R1105_U15 , REG2_REG_4_ );
not NOT1_3845 ( R1105_U16 , U3440 );
not NOT1_3846 ( R1105_U17 , REG2_REG_5_ );
not NOT1_3847 ( R1105_U18 , U3439 );
not NOT1_3848 ( R1105_U19 , REG2_REG_6_ );
not NOT1_3849 ( R1105_U20 , U3438 );
not NOT1_3850 ( R1105_U21 , REG2_REG_7_ );
not NOT1_3851 ( R1105_U22 , U3437 );
not NOT1_3852 ( R1105_U23 , REG2_REG_8_ );
not NOT1_3853 ( R1105_U24 , U3436 );
not NOT1_3854 ( R1105_U25 , U3435 );
not NOT1_3855 ( R1105_U26 , REG2_REG_9_ );
not NOT1_3856 ( R1105_U27 , REG2_REG_10_ );
not NOT1_3857 ( R1105_U28 , U3452 );
not NOT1_3858 ( R1105_U29 , REG2_REG_11_ );
not NOT1_3859 ( R1105_U30 , U3451 );
not NOT1_3860 ( R1105_U31 , REG2_REG_12_ );
not NOT1_3861 ( R1105_U32 , U3450 );
not NOT1_3862 ( R1105_U33 , REG2_REG_13_ );
not NOT1_3863 ( R1105_U34 , U3449 );
not NOT1_3864 ( R1105_U35 , REG2_REG_14_ );
not NOT1_3865 ( R1105_U36 , U3448 );
not NOT1_3866 ( R1105_U37 , REG2_REG_15_ );
not NOT1_3867 ( R1105_U38 , U3447 );
not NOT1_3868 ( R1105_U39 , REG2_REG_16_ );
not NOT1_3869 ( R1105_U40 , U3446 );
not NOT1_3870 ( R1105_U41 , REG2_REG_17_ );
not NOT1_3871 ( R1105_U42 , U3445 );
not NOT1_3872 ( R1105_U43 , REG2_REG_18_ );
not NOT1_3873 ( R1105_U44 , U3444 );
nand NAND2_3874 ( R1105_U45 , R1105_U170 , R1105_U169 );
nand NAND2_3875 ( R1105_U46 , R1105_U311 , R1105_U310 );
nand NAND2_3876 ( R1105_U47 , R1105_U187 , R1105_U186 );
nand NAND2_3877 ( R1105_U48 , R1105_U194 , R1105_U193 );
nand NAND2_3878 ( R1105_U49 , R1105_U201 , R1105_U200 );
nand NAND2_3879 ( R1105_U50 , R1105_U208 , R1105_U207 );
nand NAND2_3880 ( R1105_U51 , R1105_U215 , R1105_U214 );
nand NAND2_3881 ( R1105_U52 , R1105_U222 , R1105_U221 );
nand NAND2_3882 ( R1105_U53 , R1105_U229 , R1105_U228 );
nand NAND2_3883 ( R1105_U54 , R1105_U236 , R1105_U235 );
nand NAND2_3884 ( R1105_U55 , R1105_U253 , R1105_U252 );
nand NAND2_3885 ( R1105_U56 , R1105_U260 , R1105_U259 );
nand NAND2_3886 ( R1105_U57 , R1105_U267 , R1105_U266 );
nand NAND2_3887 ( R1105_U58 , R1105_U274 , R1105_U273 );
nand NAND2_3888 ( R1105_U59 , R1105_U281 , R1105_U280 );
nand NAND2_3889 ( R1105_U60 , R1105_U288 , R1105_U287 );
nand NAND2_3890 ( R1105_U61 , R1105_U295 , R1105_U294 );
nand NAND2_3891 ( R1105_U62 , R1105_U302 , R1105_U301 );
nand NAND2_3892 ( R1105_U63 , R1105_U309 , R1105_U308 );
and AND3_3893 ( R1105_U64 , R1105_U243 , R1105_U242 , R1105_U174 );
and AND2_3894 ( R1105_U65 , R1105_U178 , R1105_U246 );
and AND2_3895 ( R1105_U66 , R1105_U182 , R1105_U181 );
nand NAND2_3896 ( R1105_U67 , R1105_U134 , R1105_U133 );
and AND2_3897 ( R1105_U68 , R1105_U189 , R1105_U188 );
nand NAND2_3898 ( R1105_U69 , R1105_U130 , R1105_U129 );
and AND2_3899 ( R1105_U70 , R1105_U196 , R1105_U195 );
nand NAND2_3900 ( R1105_U71 , R1105_U126 , R1105_U125 );
and AND2_3901 ( R1105_U72 , R1105_U203 , R1105_U202 );
nand NAND2_3902 ( R1105_U73 , R1105_U122 , R1105_U121 );
and AND2_3903 ( R1105_U74 , R1105_U210 , R1105_U209 );
nand NAND2_3904 ( R1105_U75 , R1105_U118 , R1105_U117 );
and AND2_3905 ( R1105_U76 , R1105_U217 , R1105_U216 );
nand NAND2_3906 ( R1105_U77 , R1105_U114 , R1105_U113 );
and AND2_3907 ( R1105_U78 , R1105_U224 , R1105_U223 );
nand NAND2_3908 ( R1105_U79 , R1105_U110 , R1105_U109 );
and AND2_3909 ( R1105_U80 , R1105_U231 , R1105_U230 );
nand NAND2_3910 ( R1105_U81 , R1105_U82 , R1105_U106 );
nand NAND2_3911 ( R1105_U82 , U3443 , R1105_U104 );
and AND2_3912 ( R1105_U83 , R1105_U241 , R1105_U240 );
not NOT1_3913 ( R1105_U84 , U3461 );
not NOT1_3914 ( R1105_U85 , REG2_REG_19_ );
and AND2_3915 ( R1105_U86 , R1105_U248 , R1105_U247 );
and AND2_3916 ( R1105_U87 , R1105_U255 , R1105_U254 );
nand NAND2_3917 ( R1105_U88 , R1105_U166 , R1105_U165 );
and AND2_3918 ( R1105_U89 , R1105_U262 , R1105_U261 );
nand NAND2_3919 ( R1105_U90 , R1105_U162 , R1105_U161 );
and AND2_3920 ( R1105_U91 , R1105_U269 , R1105_U268 );
nand NAND2_3921 ( R1105_U92 , R1105_U158 , R1105_U157 );
and AND2_3922 ( R1105_U93 , R1105_U276 , R1105_U275 );
nand NAND2_3923 ( R1105_U94 , R1105_U154 , R1105_U153 );
and AND2_3924 ( R1105_U95 , R1105_U283 , R1105_U282 );
nand NAND2_3925 ( R1105_U96 , R1105_U150 , R1105_U149 );
and AND2_3926 ( R1105_U97 , R1105_U290 , R1105_U289 );
nand NAND2_3927 ( R1105_U98 , R1105_U146 , R1105_U145 );
and AND2_3928 ( R1105_U99 , R1105_U297 , R1105_U296 );
nand NAND2_3929 ( R1105_U100 , R1105_U142 , R1105_U141 );
and AND2_3930 ( R1105_U101 , R1105_U304 , R1105_U303 );
nand NAND2_3931 ( R1105_U102 , R1105_U138 , R1105_U137 );
not NOT1_3932 ( R1105_U103 , R1105_U82 );
not NOT1_3933 ( R1105_U104 , R1105_U9 );
nand NAND2_3934 ( R1105_U105 , R1105_U10 , R1105_U9 );
nand NAND2_3935 ( R1105_U106 , REG2_REG_1_ , R1105_U105 );
not NOT1_3936 ( R1105_U107 , R1105_U81 );
or OR2_3937 ( R1105_U108 , REG2_REG_2_ , U3442 );
nand NAND2_3938 ( R1105_U109 , R1105_U108 , R1105_U81 );
nand NAND2_3939 ( R1105_U110 , U3442 , REG2_REG_2_ );
not NOT1_3940 ( R1105_U111 , R1105_U79 );
or OR2_3941 ( R1105_U112 , REG2_REG_3_ , U3441 );
nand NAND2_3942 ( R1105_U113 , R1105_U112 , R1105_U79 );
nand NAND2_3943 ( R1105_U114 , U3441 , REG2_REG_3_ );
not NOT1_3944 ( R1105_U115 , R1105_U77 );
or OR2_3945 ( R1105_U116 , REG2_REG_4_ , U3440 );
nand NAND2_3946 ( R1105_U117 , R1105_U116 , R1105_U77 );
nand NAND2_3947 ( R1105_U118 , U3440 , REG2_REG_4_ );
not NOT1_3948 ( R1105_U119 , R1105_U75 );
or OR2_3949 ( R1105_U120 , REG2_REG_5_ , U3439 );
nand NAND2_3950 ( R1105_U121 , R1105_U120 , R1105_U75 );
nand NAND2_3951 ( R1105_U122 , U3439 , REG2_REG_5_ );
not NOT1_3952 ( R1105_U123 , R1105_U73 );
or OR2_3953 ( R1105_U124 , REG2_REG_6_ , U3438 );
nand NAND2_3954 ( R1105_U125 , R1105_U124 , R1105_U73 );
nand NAND2_3955 ( R1105_U126 , U3438 , REG2_REG_6_ );
not NOT1_3956 ( R1105_U127 , R1105_U71 );
or OR2_3957 ( R1105_U128 , REG2_REG_7_ , U3437 );
nand NAND2_3958 ( R1105_U129 , R1105_U128 , R1105_U71 );
nand NAND2_3959 ( R1105_U130 , U3437 , REG2_REG_7_ );
not NOT1_3960 ( R1105_U131 , R1105_U69 );
or OR2_3961 ( R1105_U132 , REG2_REG_8_ , U3436 );
nand NAND2_3962 ( R1105_U133 , R1105_U132 , R1105_U69 );
nand NAND2_3963 ( R1105_U134 , U3436 , REG2_REG_8_ );
not NOT1_3964 ( R1105_U135 , R1105_U67 );
or OR2_3965 ( R1105_U136 , REG2_REG_9_ , U3435 );
nand NAND2_3966 ( R1105_U137 , R1105_U136 , R1105_U67 );
nand NAND2_3967 ( R1105_U138 , REG2_REG_9_ , U3435 );
not NOT1_3968 ( R1105_U139 , R1105_U102 );
or OR2_3969 ( R1105_U140 , REG2_REG_10_ , U3452 );
nand NAND2_3970 ( R1105_U141 , R1105_U140 , R1105_U102 );
nand NAND2_3971 ( R1105_U142 , U3452 , REG2_REG_10_ );
not NOT1_3972 ( R1105_U143 , R1105_U100 );
or OR2_3973 ( R1105_U144 , REG2_REG_11_ , U3451 );
nand NAND2_3974 ( R1105_U145 , R1105_U144 , R1105_U100 );
nand NAND2_3975 ( R1105_U146 , U3451 , REG2_REG_11_ );
not NOT1_3976 ( R1105_U147 , R1105_U98 );
or OR2_3977 ( R1105_U148 , REG2_REG_12_ , U3450 );
nand NAND2_3978 ( R1105_U149 , R1105_U148 , R1105_U98 );
nand NAND2_3979 ( R1105_U150 , U3450 , REG2_REG_12_ );
not NOT1_3980 ( R1105_U151 , R1105_U96 );
or OR2_3981 ( R1105_U152 , REG2_REG_13_ , U3449 );
nand NAND2_3982 ( R1105_U153 , R1105_U152 , R1105_U96 );
nand NAND2_3983 ( R1105_U154 , U3449 , REG2_REG_13_ );
not NOT1_3984 ( R1105_U155 , R1105_U94 );
or OR2_3985 ( R1105_U156 , REG2_REG_14_ , U3448 );
nand NAND2_3986 ( R1105_U157 , R1105_U156 , R1105_U94 );
nand NAND2_3987 ( R1105_U158 , U3448 , REG2_REG_14_ );
not NOT1_3988 ( R1105_U159 , R1105_U92 );
or OR2_3989 ( R1105_U160 , REG2_REG_15_ , U3447 );
nand NAND2_3990 ( R1105_U161 , R1105_U160 , R1105_U92 );
nand NAND2_3991 ( R1105_U162 , U3447 , REG2_REG_15_ );
not NOT1_3992 ( R1105_U163 , R1105_U90 );
or OR2_3993 ( R1105_U164 , REG2_REG_16_ , U3446 );
nand NAND2_3994 ( R1105_U165 , R1105_U164 , R1105_U90 );
nand NAND2_3995 ( R1105_U166 , U3446 , REG2_REG_16_ );
not NOT1_3996 ( R1105_U167 , R1105_U88 );
or OR2_3997 ( R1105_U168 , REG2_REG_17_ , U3445 );
nand NAND2_3998 ( R1105_U169 , R1105_U168 , R1105_U88 );
nand NAND2_3999 ( R1105_U170 , U3445 , REG2_REG_17_ );
not NOT1_4000 ( R1105_U171 , R1105_U45 );
or OR2_4001 ( R1105_U172 , REG2_REG_18_ , U3444 );
nand NAND2_4002 ( R1105_U173 , R1105_U172 , R1105_U45 );
nand NAND2_4003 ( R1105_U174 , U3444 , REG2_REG_18_ );
nand NAND2_4004 ( R1105_U175 , R1105_U64 , R1105_U173 );
nand NAND2_4005 ( R1105_U176 , U3444 , REG2_REG_18_ );
nand NAND2_4006 ( R1105_U177 , R1105_U171 , R1105_U176 );
or OR2_4007 ( R1105_U178 , U3444 , REG2_REG_18_ );
nand NAND2_4008 ( R1105_U179 , R1105_U65 , R1105_U177 );
nand NAND2_4009 ( R1105_U180 , R1105_U239 , R1105_U10 );
nand NAND2_4010 ( R1105_U181 , U3435 , R1105_U26 );
nand NAND2_4011 ( R1105_U182 , REG2_REG_9_ , R1105_U25 );
nand NAND2_4012 ( R1105_U183 , U3435 , R1105_U26 );
nand NAND2_4013 ( R1105_U184 , REG2_REG_9_ , R1105_U25 );
nand NAND2_4014 ( R1105_U185 , R1105_U184 , R1105_U183 );
nand NAND2_4015 ( R1105_U186 , R1105_U66 , R1105_U67 );
nand NAND2_4016 ( R1105_U187 , R1105_U135 , R1105_U185 );
nand NAND2_4017 ( R1105_U188 , U3436 , R1105_U23 );
nand NAND2_4018 ( R1105_U189 , REG2_REG_8_ , R1105_U24 );
nand NAND2_4019 ( R1105_U190 , U3436 , R1105_U23 );
nand NAND2_4020 ( R1105_U191 , REG2_REG_8_ , R1105_U24 );
nand NAND2_4021 ( R1105_U192 , R1105_U191 , R1105_U190 );
nand NAND2_4022 ( R1105_U193 , R1105_U68 , R1105_U69 );
nand NAND2_4023 ( R1105_U194 , R1105_U131 , R1105_U192 );
nand NAND2_4024 ( R1105_U195 , U3437 , R1105_U21 );
nand NAND2_4025 ( R1105_U196 , REG2_REG_7_ , R1105_U22 );
nand NAND2_4026 ( R1105_U197 , U3437 , R1105_U21 );
nand NAND2_4027 ( R1105_U198 , REG2_REG_7_ , R1105_U22 );
nand NAND2_4028 ( R1105_U199 , R1105_U198 , R1105_U197 );
nand NAND2_4029 ( R1105_U200 , R1105_U70 , R1105_U71 );
nand NAND2_4030 ( R1105_U201 , R1105_U127 , R1105_U199 );
nand NAND2_4031 ( R1105_U202 , U3438 , R1105_U19 );
nand NAND2_4032 ( R1105_U203 , REG2_REG_6_ , R1105_U20 );
nand NAND2_4033 ( R1105_U204 , U3438 , R1105_U19 );
nand NAND2_4034 ( R1105_U205 , REG2_REG_6_ , R1105_U20 );
nand NAND2_4035 ( R1105_U206 , R1105_U205 , R1105_U204 );
nand NAND2_4036 ( R1105_U207 , R1105_U72 , R1105_U73 );
nand NAND2_4037 ( R1105_U208 , R1105_U123 , R1105_U206 );
nand NAND2_4038 ( R1105_U209 , U3439 , R1105_U17 );
nand NAND2_4039 ( R1105_U210 , REG2_REG_5_ , R1105_U18 );
nand NAND2_4040 ( R1105_U211 , U3439 , R1105_U17 );
nand NAND2_4041 ( R1105_U212 , REG2_REG_5_ , R1105_U18 );
nand NAND2_4042 ( R1105_U213 , R1105_U212 , R1105_U211 );
nand NAND2_4043 ( R1105_U214 , R1105_U74 , R1105_U75 );
nand NAND2_4044 ( R1105_U215 , R1105_U119 , R1105_U213 );
nand NAND2_4045 ( R1105_U216 , U3440 , R1105_U15 );
nand NAND2_4046 ( R1105_U217 , REG2_REG_4_ , R1105_U16 );
nand NAND2_4047 ( R1105_U218 , U3440 , R1105_U15 );
nand NAND2_4048 ( R1105_U219 , REG2_REG_4_ , R1105_U16 );
nand NAND2_4049 ( R1105_U220 , R1105_U219 , R1105_U218 );
nand NAND2_4050 ( R1105_U221 , R1105_U76 , R1105_U77 );
nand NAND2_4051 ( R1105_U222 , R1105_U115 , R1105_U220 );
nand NAND2_4052 ( R1105_U223 , U3441 , R1105_U13 );
nand NAND2_4053 ( R1105_U224 , REG2_REG_3_ , R1105_U14 );
nand NAND2_4054 ( R1105_U225 , U3441 , R1105_U13 );
nand NAND2_4055 ( R1105_U226 , REG2_REG_3_ , R1105_U14 );
nand NAND2_4056 ( R1105_U227 , R1105_U226 , R1105_U225 );
nand NAND2_4057 ( R1105_U228 , R1105_U78 , R1105_U79 );
nand NAND2_4058 ( R1105_U229 , R1105_U111 , R1105_U227 );
nand NAND2_4059 ( R1105_U230 , U3442 , R1105_U11 );
nand NAND2_4060 ( R1105_U231 , REG2_REG_2_ , R1105_U12 );
nand NAND2_4061 ( R1105_U232 , U3442 , R1105_U11 );
nand NAND2_4062 ( R1105_U233 , REG2_REG_2_ , R1105_U12 );
nand NAND2_4063 ( R1105_U234 , R1105_U233 , R1105_U232 );
nand NAND2_4064 ( R1105_U235 , R1105_U80 , R1105_U81 );
nand NAND2_4065 ( R1105_U236 , R1105_U107 , R1105_U234 );
nand NAND2_4066 ( R1105_U237 , REG2_REG_1_ , R1105_U9 );
nand NAND2_4067 ( R1105_U238 , R1105_U104 , R1105_U8 );
nand NAND2_4068 ( R1105_U239 , R1105_U238 , R1105_U237 );
nand NAND3_4069 ( R1105_U240 , U3443 , R1105_U9 , R1105_U8 );
nand NAND2_4070 ( R1105_U241 , R1105_U103 , REG2_REG_1_ );
nand NAND2_4071 ( R1105_U242 , U3461 , R1105_U85 );
nand NAND2_4072 ( R1105_U243 , REG2_REG_19_ , R1105_U84 );
nand NAND2_4073 ( R1105_U244 , U3461 , R1105_U85 );
nand NAND2_4074 ( R1105_U245 , REG2_REG_19_ , R1105_U84 );
nand NAND2_4075 ( R1105_U246 , R1105_U245 , R1105_U244 );
nand NAND2_4076 ( R1105_U247 , U3444 , R1105_U43 );
nand NAND2_4077 ( R1105_U248 , REG2_REG_18_ , R1105_U44 );
nand NAND2_4078 ( R1105_U249 , U3444 , R1105_U43 );
nand NAND2_4079 ( R1105_U250 , REG2_REG_18_ , R1105_U44 );
nand NAND2_4080 ( R1105_U251 , R1105_U250 , R1105_U249 );
nand NAND2_4081 ( R1105_U252 , R1105_U86 , R1105_U45 );
nand NAND2_4082 ( R1105_U253 , R1105_U251 , R1105_U171 );
nand NAND2_4083 ( R1105_U254 , U3445 , R1105_U41 );
nand NAND2_4084 ( R1105_U255 , REG2_REG_17_ , R1105_U42 );
nand NAND2_4085 ( R1105_U256 , U3445 , R1105_U41 );
nand NAND2_4086 ( R1105_U257 , REG2_REG_17_ , R1105_U42 );
nand NAND2_4087 ( R1105_U258 , R1105_U257 , R1105_U256 );
nand NAND2_4088 ( R1105_U259 , R1105_U87 , R1105_U88 );
nand NAND2_4089 ( R1105_U260 , R1105_U167 , R1105_U258 );
nand NAND2_4090 ( R1105_U261 , U3446 , R1105_U39 );
nand NAND2_4091 ( R1105_U262 , REG2_REG_16_ , R1105_U40 );
nand NAND2_4092 ( R1105_U263 , U3446 , R1105_U39 );
nand NAND2_4093 ( R1105_U264 , REG2_REG_16_ , R1105_U40 );
nand NAND2_4094 ( R1105_U265 , R1105_U264 , R1105_U263 );
nand NAND2_4095 ( R1105_U266 , R1105_U89 , R1105_U90 );
nand NAND2_4096 ( R1105_U267 , R1105_U163 , R1105_U265 );
nand NAND2_4097 ( R1105_U268 , U3447 , R1105_U37 );
nand NAND2_4098 ( R1105_U269 , REG2_REG_15_ , R1105_U38 );
nand NAND2_4099 ( R1105_U270 , U3447 , R1105_U37 );
nand NAND2_4100 ( R1105_U271 , REG2_REG_15_ , R1105_U38 );
nand NAND2_4101 ( R1105_U272 , R1105_U271 , R1105_U270 );
nand NAND2_4102 ( R1105_U273 , R1105_U91 , R1105_U92 );
nand NAND2_4103 ( R1105_U274 , R1105_U159 , R1105_U272 );
nand NAND2_4104 ( R1105_U275 , U3448 , R1105_U35 );
nand NAND2_4105 ( R1105_U276 , REG2_REG_14_ , R1105_U36 );
nand NAND2_4106 ( R1105_U277 , U3448 , R1105_U35 );
nand NAND2_4107 ( R1105_U278 , REG2_REG_14_ , R1105_U36 );
nand NAND2_4108 ( R1105_U279 , R1105_U278 , R1105_U277 );
nand NAND2_4109 ( R1105_U280 , R1105_U93 , R1105_U94 );
nand NAND2_4110 ( R1105_U281 , R1105_U155 , R1105_U279 );
nand NAND2_4111 ( R1105_U282 , U3449 , R1105_U33 );
nand NAND2_4112 ( R1105_U283 , REG2_REG_13_ , R1105_U34 );
nand NAND2_4113 ( R1105_U284 , U3449 , R1105_U33 );
nand NAND2_4114 ( R1105_U285 , REG2_REG_13_ , R1105_U34 );
nand NAND2_4115 ( R1105_U286 , R1105_U285 , R1105_U284 );
nand NAND2_4116 ( R1105_U287 , R1105_U95 , R1105_U96 );
nand NAND2_4117 ( R1105_U288 , R1105_U151 , R1105_U286 );
nand NAND2_4118 ( R1105_U289 , U3450 , R1105_U31 );
nand NAND2_4119 ( R1105_U290 , REG2_REG_12_ , R1105_U32 );
nand NAND2_4120 ( R1105_U291 , U3450 , R1105_U31 );
nand NAND2_4121 ( R1105_U292 , REG2_REG_12_ , R1105_U32 );
nand NAND2_4122 ( R1105_U293 , R1105_U292 , R1105_U291 );
nand NAND2_4123 ( R1105_U294 , R1105_U97 , R1105_U98 );
nand NAND2_4124 ( R1105_U295 , R1105_U147 , R1105_U293 );
nand NAND2_4125 ( R1105_U296 , U3451 , R1105_U29 );
nand NAND2_4126 ( R1105_U297 , REG2_REG_11_ , R1105_U30 );
nand NAND2_4127 ( R1105_U298 , U3451 , R1105_U29 );
nand NAND2_4128 ( R1105_U299 , REG2_REG_11_ , R1105_U30 );
nand NAND2_4129 ( R1105_U300 , R1105_U299 , R1105_U298 );
nand NAND2_4130 ( R1105_U301 , R1105_U99 , R1105_U100 );
nand NAND2_4131 ( R1105_U302 , R1105_U143 , R1105_U300 );
nand NAND2_4132 ( R1105_U303 , U3452 , R1105_U27 );
nand NAND2_4133 ( R1105_U304 , REG2_REG_10_ , R1105_U28 );
nand NAND2_4134 ( R1105_U305 , U3452 , R1105_U27 );
nand NAND2_4135 ( R1105_U306 , REG2_REG_10_ , R1105_U28 );
nand NAND2_4136 ( R1105_U307 , R1105_U306 , R1105_U305 );
nand NAND2_4137 ( R1105_U308 , R1105_U101 , R1105_U102 );
nand NAND2_4138 ( R1105_U309 , R1105_U139 , R1105_U307 );
nand NAND2_4139 ( R1105_U310 , U3453 , R1105_U6 );
nand NAND2_4140 ( R1105_U311 , REG2_REG_0_ , R1105_U7 );
not NOT1_4141 ( R1309_U6 , U3056 );
not NOT1_4142 ( R1309_U7 , U3053 );
and AND2_4143 ( R1309_U8 , R1309_U10 , R1309_U9 );
nand NAND2_4144 ( R1309_U9 , U3053 , R1309_U6 );
nand NAND2_4145 ( R1309_U10 , U3056 , R1309_U7 );
and AND2_4146 ( R1282_U6 , R1282_U130 , R1282_U12 );
and AND2_4147 ( R1282_U7 , R1282_U106 , R1282_U96 );
and AND2_4148 ( R1282_U8 , R1282_U105 , R1282_U13 );
and AND2_4149 ( R1282_U9 , R1282_U104 , R1282_U98 );
and AND2_4150 ( R1282_U10 , R1282_U103 , R1282_U14 );
and AND2_4151 ( R1282_U11 , R1282_U102 , R1282_U35 );
or OR3_4152 ( R1282_U12 , U3468 , U3464 , U3470 );
nand NAND3_4153 ( R1282_U13 , R1282_U19 , R1282_U20 , R1282_U95 );
nand NAND3_4154 ( R1282_U14 , R1282_U17 , R1282_U18 , R1282_U97 );
nand NAND3_4155 ( R1282_U15 , R1282_U34 , R1282_U16 , R1282_U99 );
not NOT1_4156 ( R1282_U16 , U3480 );
not NOT1_4157 ( R1282_U17 , U3478 );
not NOT1_4158 ( R1282_U18 , U3476 );
not NOT1_4159 ( R1282_U19 , U3474 );
not NOT1_4160 ( R1282_U20 , U3472 );
nand NAND3_4161 ( R1282_U21 , R1282_U32 , R1282_U92 , R1282_U101 );
nand NAND3_4162 ( R1282_U22 , R1282_U87 , R1282_U90 , R1282_U108 );
nand NAND3_4163 ( R1282_U23 , R1282_U82 , R1282_U85 , R1282_U110 );
nand NAND3_4164 ( R1282_U24 , R1282_U77 , R1282_U80 , R1282_U112 );
nand NAND3_4165 ( R1282_U25 , R1282_U72 , R1282_U75 , R1282_U114 );
nand NAND3_4166 ( R1282_U26 , R1282_U65 , R1282_U70 , R1282_U116 );
nand NAND3_4167 ( R1282_U27 , R1282_U60 , R1282_U63 , R1282_U118 );
nand NAND3_4168 ( R1282_U28 , R1282_U55 , R1282_U58 , R1282_U120 );
nand NAND3_4169 ( R1282_U29 , R1282_U50 , R1282_U53 , R1282_U122 );
nand NAND3_4170 ( R1282_U30 , R1282_U45 , R1282_U48 , R1282_U124 );
nand NAND2_4171 ( R1282_U31 , R1282_U160 , R1282_U159 );
not NOT1_4172 ( R1282_U32 , U3484 );
and AND2_4173 ( R1282_U33 , R1282_U132 , R1282_U131 );
not NOT1_4174 ( R1282_U34 , U3482 );
nand NAND2_4175 ( R1282_U35 , R1282_U99 , R1282_U16 );
and AND2_4176 ( R1282_U36 , R1282_U134 , R1282_U133 );
not NOT1_4177 ( R1282_U37 , U4038 );
nand NAND3_4178 ( R1282_U38 , R1282_U40 , R1282_U43 , R1282_U126 );
and AND2_4179 ( R1282_U39 , R1282_U136 , R1282_U135 );
not NOT1_4180 ( R1282_U40 , U4039 );
nand NAND2_4181 ( R1282_U41 , R1282_U126 , R1282_U43 );
and AND2_4182 ( R1282_U42 , R1282_U138 , R1282_U137 );
not NOT1_4183 ( R1282_U43 , U4040 );
and AND2_4184 ( R1282_U44 , R1282_U140 , R1282_U139 );
not NOT1_4185 ( R1282_U45 , U4029 );
nand NAND2_4186 ( R1282_U46 , R1282_U124 , R1282_U48 );
and AND2_4187 ( R1282_U47 , R1282_U142 , R1282_U141 );
not NOT1_4188 ( R1282_U48 , U4030 );
and AND2_4189 ( R1282_U49 , R1282_U144 , R1282_U143 );
not NOT1_4190 ( R1282_U50 , U4031 );
nand NAND2_4191 ( R1282_U51 , R1282_U122 , R1282_U53 );
and AND2_4192 ( R1282_U52 , R1282_U146 , R1282_U145 );
not NOT1_4193 ( R1282_U53 , U4032 );
and AND2_4194 ( R1282_U54 , R1282_U148 , R1282_U147 );
not NOT1_4195 ( R1282_U55 , U4033 );
nand NAND2_4196 ( R1282_U56 , R1282_U120 , R1282_U58 );
and AND2_4197 ( R1282_U57 , R1282_U150 , R1282_U149 );
not NOT1_4198 ( R1282_U58 , U4034 );
and AND2_4199 ( R1282_U59 , R1282_U152 , R1282_U151 );
not NOT1_4200 ( R1282_U60 , U4035 );
nand NAND2_4201 ( R1282_U61 , R1282_U118 , R1282_U63 );
and AND2_4202 ( R1282_U62 , R1282_U154 , R1282_U153 );
not NOT1_4203 ( R1282_U63 , U4036 );
and AND2_4204 ( R1282_U64 , R1282_U156 , R1282_U155 );
not NOT1_4205 ( R1282_U65 , U4037 );
nand NAND2_4206 ( R1282_U66 , R1282_U116 , R1282_U70 );
and AND2_4207 ( R1282_U67 , R1282_U158 , R1282_U157 );
not NOT1_4208 ( R1282_U68 , U3468 );
not NOT1_4209 ( R1282_U69 , U3464 );
not NOT1_4210 ( R1282_U70 , U3504 );
and AND2_4211 ( R1282_U71 , R1282_U162 , R1282_U161 );
not NOT1_4212 ( R1282_U72 , U3502 );
nand NAND2_4213 ( R1282_U73 , R1282_U114 , R1282_U75 );
and AND2_4214 ( R1282_U74 , R1282_U164 , R1282_U163 );
not NOT1_4215 ( R1282_U75 , U3500 );
and AND2_4216 ( R1282_U76 , R1282_U166 , R1282_U165 );
not NOT1_4217 ( R1282_U77 , U3498 );
nand NAND2_4218 ( R1282_U78 , R1282_U112 , R1282_U80 );
and AND2_4219 ( R1282_U79 , R1282_U168 , R1282_U167 );
not NOT1_4220 ( R1282_U80 , U3496 );
and AND2_4221 ( R1282_U81 , R1282_U170 , R1282_U169 );
not NOT1_4222 ( R1282_U82 , U3494 );
nand NAND2_4223 ( R1282_U83 , R1282_U110 , R1282_U85 );
and AND2_4224 ( R1282_U84 , R1282_U172 , R1282_U171 );
not NOT1_4225 ( R1282_U85 , U3492 );
and AND2_4226 ( R1282_U86 , R1282_U174 , R1282_U173 );
not NOT1_4227 ( R1282_U87 , U3490 );
nand NAND2_4228 ( R1282_U88 , R1282_U108 , R1282_U90 );
and AND2_4229 ( R1282_U89 , R1282_U176 , R1282_U175 );
not NOT1_4230 ( R1282_U90 , U3488 );
and AND2_4231 ( R1282_U91 , R1282_U178 , R1282_U177 );
not NOT1_4232 ( R1282_U92 , U3486 );
nand NAND2_4233 ( R1282_U93 , R1282_U101 , R1282_U32 );
and AND2_4234 ( R1282_U94 , R1282_U180 , R1282_U179 );
not NOT1_4235 ( R1282_U95 , R1282_U12 );
nand NAND2_4236 ( R1282_U96 , R1282_U95 , R1282_U20 );
not NOT1_4237 ( R1282_U97 , R1282_U13 );
nand NAND2_4238 ( R1282_U98 , R1282_U97 , R1282_U18 );
not NOT1_4239 ( R1282_U99 , R1282_U14 );
not NOT1_4240 ( R1282_U100 , R1282_U35 );
not NOT1_4241 ( R1282_U101 , R1282_U15 );
nand NAND2_4242 ( R1282_U102 , U3480 , R1282_U14 );
nand NAND2_4243 ( R1282_U103 , U3478 , R1282_U98 );
nand NAND2_4244 ( R1282_U104 , U3476 , R1282_U13 );
nand NAND2_4245 ( R1282_U105 , U3474 , R1282_U96 );
nand NAND2_4246 ( R1282_U106 , U3472 , R1282_U12 );
not NOT1_4247 ( R1282_U107 , R1282_U93 );
not NOT1_4248 ( R1282_U108 , R1282_U21 );
not NOT1_4249 ( R1282_U109 , R1282_U88 );
not NOT1_4250 ( R1282_U110 , R1282_U22 );
not NOT1_4251 ( R1282_U111 , R1282_U83 );
not NOT1_4252 ( R1282_U112 , R1282_U23 );
not NOT1_4253 ( R1282_U113 , R1282_U78 );
not NOT1_4254 ( R1282_U114 , R1282_U24 );
not NOT1_4255 ( R1282_U115 , R1282_U73 );
not NOT1_4256 ( R1282_U116 , R1282_U25 );
not NOT1_4257 ( R1282_U117 , R1282_U66 );
not NOT1_4258 ( R1282_U118 , R1282_U26 );
not NOT1_4259 ( R1282_U119 , R1282_U61 );
not NOT1_4260 ( R1282_U120 , R1282_U27 );
not NOT1_4261 ( R1282_U121 , R1282_U56 );
not NOT1_4262 ( R1282_U122 , R1282_U28 );
not NOT1_4263 ( R1282_U123 , R1282_U51 );
not NOT1_4264 ( R1282_U124 , R1282_U29 );
not NOT1_4265 ( R1282_U125 , R1282_U46 );
not NOT1_4266 ( R1282_U126 , R1282_U30 );
not NOT1_4267 ( R1282_U127 , R1282_U41 );
not NOT1_4268 ( R1282_U128 , R1282_U38 );
or OR2_4269 ( R1282_U129 , U3468 , U3464 );
nand NAND2_4270 ( R1282_U130 , U3470 , R1282_U129 );
nand NAND2_4271 ( R1282_U131 , U3484 , R1282_U15 );
nand NAND2_4272 ( R1282_U132 , R1282_U101 , R1282_U32 );
nand NAND2_4273 ( R1282_U133 , U3482 , R1282_U35 );
nand NAND2_4274 ( R1282_U134 , R1282_U100 , R1282_U34 );
nand NAND2_4275 ( R1282_U135 , U4038 , R1282_U38 );
nand NAND2_4276 ( R1282_U136 , R1282_U128 , R1282_U37 );
nand NAND2_4277 ( R1282_U137 , U4039 , R1282_U41 );
nand NAND2_4278 ( R1282_U138 , R1282_U127 , R1282_U40 );
nand NAND2_4279 ( R1282_U139 , U4040 , R1282_U30 );
nand NAND2_4280 ( R1282_U140 , R1282_U126 , R1282_U43 );
nand NAND2_4281 ( R1282_U141 , U4029 , R1282_U46 );
nand NAND2_4282 ( R1282_U142 , R1282_U125 , R1282_U45 );
nand NAND2_4283 ( R1282_U143 , U4030 , R1282_U29 );
nand NAND2_4284 ( R1282_U144 , R1282_U124 , R1282_U48 );
nand NAND2_4285 ( R1282_U145 , U4031 , R1282_U51 );
nand NAND2_4286 ( R1282_U146 , R1282_U123 , R1282_U50 );
nand NAND2_4287 ( R1282_U147 , U4032 , R1282_U28 );
nand NAND2_4288 ( R1282_U148 , R1282_U122 , R1282_U53 );
nand NAND2_4289 ( R1282_U149 , U4033 , R1282_U56 );
nand NAND2_4290 ( R1282_U150 , R1282_U121 , R1282_U55 );
nand NAND2_4291 ( R1282_U151 , U4034 , R1282_U27 );
nand NAND2_4292 ( R1282_U152 , R1282_U120 , R1282_U58 );
nand NAND2_4293 ( R1282_U153 , U4035 , R1282_U61 );
nand NAND2_4294 ( R1282_U154 , R1282_U119 , R1282_U60 );
nand NAND2_4295 ( R1282_U155 , U4036 , R1282_U26 );
nand NAND2_4296 ( R1282_U156 , R1282_U118 , R1282_U63 );
nand NAND2_4297 ( R1282_U157 , U4037 , R1282_U66 );
nand NAND2_4298 ( R1282_U158 , R1282_U117 , R1282_U65 );
nand NAND2_4299 ( R1282_U159 , U3468 , R1282_U69 );
nand NAND2_4300 ( R1282_U160 , U3464 , R1282_U68 );
nand NAND2_4301 ( R1282_U161 , U3504 , R1282_U25 );
nand NAND2_4302 ( R1282_U162 , R1282_U116 , R1282_U70 );
nand NAND2_4303 ( R1282_U163 , U3502 , R1282_U73 );
nand NAND2_4304 ( R1282_U164 , R1282_U115 , R1282_U72 );
nand NAND2_4305 ( R1282_U165 , U3500 , R1282_U24 );
nand NAND2_4306 ( R1282_U166 , R1282_U114 , R1282_U75 );
nand NAND2_4307 ( R1282_U167 , U3498 , R1282_U78 );
nand NAND2_4308 ( R1282_U168 , R1282_U113 , R1282_U77 );
nand NAND2_4309 ( R1282_U169 , U3496 , R1282_U23 );
nand NAND2_4310 ( R1282_U170 , R1282_U112 , R1282_U80 );
nand NAND2_4311 ( R1282_U171 , U3494 , R1282_U83 );
nand NAND2_4312 ( R1282_U172 , R1282_U111 , R1282_U82 );
nand NAND2_4313 ( R1282_U173 , U3492 , R1282_U22 );
nand NAND2_4314 ( R1282_U174 , R1282_U110 , R1282_U85 );
nand NAND2_4315 ( R1282_U175 , U3490 , R1282_U88 );
nand NAND2_4316 ( R1282_U176 , R1282_U109 , R1282_U87 );
nand NAND2_4317 ( R1282_U177 , U3488 , R1282_U21 );
nand NAND2_4318 ( R1282_U178 , R1282_U108 , R1282_U90 );
nand NAND2_4319 ( R1282_U179 , U3486 , R1282_U93 );
nand NAND2_4320 ( R1282_U180 , R1282_U107 , R1282_U92 );
and AND2_4321 ( R1240_U4 , R1240_U196 , R1240_U195 );
and AND2_4322 ( R1240_U5 , R1240_U197 , R1240_U198 );
and AND2_4323 ( R1240_U6 , R1240_U210 , R1240_U209 );
and AND2_4324 ( R1240_U7 , R1240_U250 , R1240_U249 );
and AND2_4325 ( R1240_U8 , R1240_U258 , R1240_U257 );
and AND2_4326 ( R1240_U9 , R1240_U274 , R1240_U273 );
and AND2_4327 ( R1240_U10 , R1240_U282 , R1240_U281 );
and AND2_4328 ( R1240_U11 , R1240_U10 , R1240_U283 );
and AND2_4329 ( R1240_U12 , R1240_U7 , R1240_U217 );
and AND2_4330 ( R1240_U13 , R1240_U8 , R1240_U262 );
and AND2_4331 ( R1240_U14 , R1240_U11 , R1240_U292 );
and AND2_4332 ( R1240_U15 , R1240_U13 , R1240_U267 );
and AND2_4333 ( R1240_U16 , R1240_U9 , R1240_U14 );
and AND2_4334 ( R1240_U17 , R1240_U299 , R1240_U305 );
and AND2_4335 ( R1240_U18 , R1240_U359 , R1240_U356 );
and AND2_4336 ( R1240_U19 , R1240_U352 , R1240_U349 );
and AND2_4337 ( R1240_U20 , R1240_U343 , R1240_U340 );
and AND2_4338 ( R1240_U21 , R1240_U334 , R1240_U331 );
and AND2_4339 ( R1240_U22 , R1240_U328 , R1240_U326 );
and AND2_4340 ( R1240_U23 , R1240_U321 , R1240_U318 );
and AND2_4341 ( R1240_U24 , R1240_U248 , R1240_U245 );
and AND2_4342 ( R1240_U25 , R1240_U240 , R1240_U237 );
and AND2_4343 ( R1240_U26 , R1240_U226 , R1240_U223 );
not NOT1_4344 ( R1240_U27 , U3470 );
not NOT1_4345 ( R1240_U28 , U3065 );
not NOT1_4346 ( R1240_U29 , U3472 );
not NOT1_4347 ( R1240_U30 , U3061 );
not NOT1_4348 ( R1240_U31 , U3474 );
not NOT1_4349 ( R1240_U32 , U3057 );
not NOT1_4350 ( R1240_U33 , U3064 );
nand NAND2_4351 ( R1240_U34 , U3057 , U3474 );
not NOT1_4352 ( R1240_U35 , U3476 );
nand NAND2_4353 ( R1240_U36 , U3468 , U3075 );
not NOT1_4354 ( R1240_U37 , U3464 );
not NOT1_4355 ( R1240_U38 , U3074 );
nand NAND2_4356 ( R1240_U39 , R1240_U131 , R1240_U200 );
not NOT1_4357 ( R1240_U40 , U3478 );
not NOT1_4358 ( R1240_U41 , U3068 );
not NOT1_4359 ( R1240_U42 , U3067 );
nand NAND2_4360 ( R1240_U43 , U3068 , U3478 );
not NOT1_4361 ( R1240_U44 , U3480 );
nand NAND2_4362 ( R1240_U45 , R1240_U214 , R1240_U213 );
not NOT1_4363 ( R1240_U46 , U3482 );
not NOT1_4364 ( R1240_U47 , U3081 );
not NOT1_4365 ( R1240_U48 , U3080 );
not NOT1_4366 ( R1240_U49 , U3484 );
nand NAND2_4367 ( R1240_U50 , R1240_U65 , R1240_U218 );
nand NAND2_4368 ( R1240_U51 , R1240_U133 , R1240_U132 );
nand NAND2_4369 ( R1240_U52 , R1240_U136 , R1240_U232 );
nand NAND2_4370 ( R1240_U53 , R1240_U229 , R1240_U228 );
not NOT1_4371 ( R1240_U54 , U4030 );
not NOT1_4372 ( R1240_U55 , U3050 );
not NOT1_4373 ( R1240_U56 , U3054 );
not NOT1_4374 ( R1240_U57 , U4031 );
not NOT1_4375 ( R1240_U58 , U4033 );
not NOT1_4376 ( R1240_U59 , U3062 );
nand NAND2_4377 ( R1240_U60 , U3062 , U4033 );
not NOT1_4378 ( R1240_U61 , U4035 );
not NOT1_4379 ( R1240_U62 , U3058 );
not NOT1_4380 ( R1240_U63 , U3496 );
not NOT1_4381 ( R1240_U64 , U3071 );
nand NAND2_4382 ( R1240_U65 , U3081 , U3482 );
not NOT1_4383 ( R1240_U66 , U3486 );
not NOT1_4384 ( R1240_U67 , U3059 );
not NOT1_4385 ( R1240_U68 , U3490 );
not NOT1_4386 ( R1240_U69 , U3069 );
not NOT1_4387 ( R1240_U70 , U3488 );
not NOT1_4388 ( R1240_U71 , U3060 );
nand NAND2_4389 ( R1240_U72 , U3060 , U3488 );
not NOT1_4390 ( R1240_U73 , U3492 );
not NOT1_4391 ( R1240_U74 , U3077 );
not NOT1_4392 ( R1240_U75 , U3494 );
not NOT1_4393 ( R1240_U76 , U3076 );
nand NAND2_4394 ( R1240_U77 , R1240_U380 , R1240_U267 );
not NOT1_4395 ( R1240_U78 , U3504 );
not NOT1_4396 ( R1240_U79 , U3078 );
nand NAND2_4397 ( R1240_U80 , U3078 , U3504 );
not NOT1_4398 ( R1240_U81 , U4037 );
not NOT1_4399 ( R1240_U82 , U3502 );
not NOT1_4400 ( R1240_U83 , U3079 );
nand NAND2_4401 ( R1240_U84 , U3079 , U3502 );
not NOT1_4402 ( R1240_U85 , U4036 );
not NOT1_4403 ( R1240_U86 , U3072 );
not NOT1_4404 ( R1240_U87 , U3498 );
not NOT1_4405 ( R1240_U88 , U3070 );
not NOT1_4406 ( R1240_U89 , U3066 );
nand NAND2_4407 ( R1240_U90 , U3070 , U3498 );
not NOT1_4408 ( R1240_U91 , U3500 );
not NOT1_4409 ( R1240_U92 , U4034 );
not NOT1_4410 ( R1240_U93 , U3063 );
nand NAND2_4411 ( R1240_U94 , R1240_U146 , R1240_U388 );
not NOT1_4412 ( R1240_U95 , U4032 );
not NOT1_4413 ( R1240_U96 , U3055 );
nand NAND3_4414 ( R1240_U97 , R1240_U396 , R1240_U306 , R1240_U397 );
not NOT1_4415 ( R1240_U98 , U3051 );
not NOT1_4416 ( R1240_U99 , U4029 );
nand NAND2_4417 ( R1240_U100 , R1240_U60 , R1240_U314 );
nand NAND2_4418 ( R1240_U101 , R1240_U385 , R1240_U294 );
nand NAND2_4419 ( R1240_U102 , R1240_U278 , R1240_U277 );
not NOT1_4420 ( R1240_U103 , U3073 );
nand NAND2_4421 ( R1240_U104 , R1240_U84 , R1240_U323 );
nand NAND3_4422 ( R1240_U105 , R1240_U383 , R1240_U271 , R1240_U382 );
nand NAND2_4423 ( R1240_U106 , R1240_U72 , R1240_U345 );
nand NAND2_4424 ( R1240_U107 , R1240_U484 , R1240_U483 );
nand NAND2_4425 ( R1240_U108 , R1240_U531 , R1240_U530 );
nand NAND2_4426 ( R1240_U109 , R1240_U402 , R1240_U401 );
nand NAND2_4427 ( R1240_U110 , R1240_U407 , R1240_U406 );
nand NAND2_4428 ( R1240_U111 , R1240_U414 , R1240_U413 );
nand NAND2_4429 ( R1240_U112 , R1240_U421 , R1240_U420 );
nand NAND2_4430 ( R1240_U113 , R1240_U426 , R1240_U425 );
nand NAND2_4431 ( R1240_U114 , R1240_U435 , R1240_U434 );
nand NAND2_4432 ( R1240_U115 , R1240_U442 , R1240_U441 );
nand NAND2_4433 ( R1240_U116 , R1240_U449 , R1240_U448 );
nand NAND2_4434 ( R1240_U117 , R1240_U456 , R1240_U455 );
nand NAND2_4435 ( R1240_U118 , R1240_U461 , R1240_U460 );
nand NAND2_4436 ( R1240_U119 , R1240_U468 , R1240_U467 );
nand NAND2_4437 ( R1240_U120 , R1240_U475 , R1240_U474 );
nand NAND2_4438 ( R1240_U121 , R1240_U489 , R1240_U488 );
nand NAND2_4439 ( R1240_U122 , R1240_U494 , R1240_U493 );
nand NAND2_4440 ( R1240_U123 , R1240_U501 , R1240_U500 );
nand NAND2_4441 ( R1240_U124 , R1240_U508 , R1240_U507 );
nand NAND2_4442 ( R1240_U125 , R1240_U515 , R1240_U514 );
nand NAND2_4443 ( R1240_U126 , R1240_U522 , R1240_U521 );
nand NAND2_4444 ( R1240_U127 , R1240_U527 , R1240_U526 );
and AND2_4445 ( R1240_U128 , R1240_U129 , R1240_U197 );
and AND2_4446 ( R1240_U129 , U3065 , U3470 );
and AND2_4447 ( R1240_U130 , U3472 , U3061 );
and AND2_4448 ( R1240_U131 , U3464 , U3074 );
and AND3_4449 ( R1240_U132 , R1240_U204 , R1240_U206 , R1240_U203 );
and AND3_4450 ( R1240_U133 , R1240_U373 , R1240_U207 , R1240_U374 );
and AND3_4451 ( R1240_U134 , R1240_U409 , R1240_U408 , R1240_U43 );
and AND2_4452 ( R1240_U135 , R1240_U225 , R1240_U6 );
and AND2_4453 ( R1240_U136 , R1240_U233 , R1240_U231 );
and AND3_4454 ( R1240_U137 , R1240_U416 , R1240_U415 , R1240_U34 );
and AND2_4455 ( R1240_U138 , R1240_U239 , R1240_U4 );
and AND2_4456 ( R1240_U139 , R1240_U247 , R1240_U198 );
and AND2_4457 ( R1240_U140 , R1240_U252 , R1240_U188 );
and AND2_4458 ( R1240_U141 , R1240_U6 , R1240_U12 );
and AND2_4459 ( R1240_U142 , R1240_U378 , R1240_U255 );
and AND2_4460 ( R1240_U143 , R1240_U270 , R1240_U15 );
and AND2_4461 ( R1240_U144 , R1240_U260 , R1240_U189 );
and AND2_4462 ( R1240_U145 , R1240_U296 , R1240_U16 );
and AND2_4463 ( R1240_U146 , R1240_U389 , R1240_U297 );
and AND2_4464 ( R1240_U147 , R1240_U309 , R1240_U185 );
and AND3_4465 ( R1240_U148 , R1240_U393 , R1240_U310 , R1240_U395 );
and AND2_4466 ( R1240_U149 , R1240_U17 , R1240_U185 );
and AND2_4467 ( R1240_U150 , R1240_U97 , R1240_U304 );
and AND3_4468 ( R1240_U151 , R1240_U451 , R1240_U450 , R1240_U190 );
and AND2_4469 ( R1240_U152 , R1240_U320 , R1240_U185 );
and AND2_4470 ( R1240_U153 , R1240_U176 , R1240_U288 );
and AND3_4471 ( R1240_U154 , R1240_U482 , R1240_U481 , R1240_U80 );
and AND2_4472 ( R1240_U155 , R1240_U333 , R1240_U10 );
and AND3_4473 ( R1240_U156 , R1240_U496 , R1240_U495 , R1240_U90 );
and AND2_4474 ( R1240_U157 , R1240_U342 , R1240_U9 );
and AND3_4475 ( R1240_U158 , R1240_U517 , R1240_U516 , R1240_U189 );
and AND2_4476 ( R1240_U159 , R1240_U351 , R1240_U8 );
and AND3_4477 ( R1240_U160 , R1240_U529 , R1240_U528 , R1240_U188 );
and AND2_4478 ( R1240_U161 , R1240_U358 , R1240_U7 );
nand NAND2_4479 ( R1240_U162 , R1240_U375 , R1240_U215 );
nand NAND2_4480 ( R1240_U163 , R1240_U230 , R1240_U242 );
not NOT1_4481 ( R1240_U164 , U3052 );
not NOT1_4482 ( R1240_U165 , U4040 );
and AND2_4483 ( R1240_U166 , R1240_U430 , R1240_U429 );
nand NAND3_4484 ( R1240_U167 , R1240_U312 , R1240_U186 , R1240_U372 );
and AND2_4485 ( R1240_U168 , R1240_U437 , R1240_U436 );
nand NAND2_4486 ( R1240_U169 , R1240_U148 , R1240_U394 );
and AND2_4487 ( R1240_U170 , R1240_U444 , R1240_U443 );
nand NAND2_4488 ( R1240_U171 , R1240_U150 , R1240_U307 );
nand NAND2_4489 ( R1240_U172 , R1240_U301 , R1240_U300 );
and AND2_4490 ( R1240_U173 , R1240_U463 , R1240_U462 );
and AND2_4491 ( R1240_U174 , R1240_U470 , R1240_U469 );
nand NAND2_4492 ( R1240_U175 , R1240_U386 , R1240_U384 );
and AND2_4493 ( R1240_U176 , R1240_U477 , R1240_U476 );
nand NAND2_4494 ( R1240_U177 , U3074 , U3464 );
nand NAND2_4495 ( R1240_U178 , R1240_U36 , R1240_U335 );
nand NAND2_4496 ( R1240_U179 , R1240_U376 , R1240_U279 );
and AND2_4497 ( R1240_U180 , R1240_U503 , R1240_U502 );
nand NAND2_4498 ( R1240_U181 , R1240_U77 , R1240_U379 );
and AND2_4499 ( R1240_U182 , R1240_U510 , R1240_U509 );
nand NAND2_4500 ( R1240_U183 , R1240_U265 , R1240_U264 );
nand NAND2_4501 ( R1240_U184 , R1240_U142 , R1240_U377 );
nand NAND2_4502 ( R1240_U185 , R1240_U391 , R1240_U390 );
nand NAND2_4503 ( R1240_U186 , U3051 , R1240_U169 );
not NOT1_4504 ( R1240_U187 , R1240_U34 );
nand NAND2_4505 ( R1240_U188 , U3484 , U3080 );
nand NAND2_4506 ( R1240_U189 , U3069 , U3490 );
nand NAND2_4507 ( R1240_U190 , U3055 , U4032 );
not NOT1_4508 ( R1240_U191 , R1240_U72 );
not NOT1_4509 ( R1240_U192 , R1240_U84 );
not NOT1_4510 ( R1240_U193 , R1240_U60 );
not NOT1_4511 ( R1240_U194 , R1240_U65 );
or OR2_4512 ( R1240_U195 , U3064 , U3476 );
or OR2_4513 ( R1240_U196 , U3057 , U3474 );
or OR2_4514 ( R1240_U197 , U3472 , U3061 );
or OR2_4515 ( R1240_U198 , U3470 , U3065 );
not NOT1_4516 ( R1240_U199 , R1240_U177 );
or OR2_4517 ( R1240_U200 , U3468 , U3075 );
not NOT1_4518 ( R1240_U201 , R1240_U39 );
not NOT1_4519 ( R1240_U202 , R1240_U36 );
nand NAND2_4520 ( R1240_U203 , R1240_U4 , R1240_U128 );
nand NAND2_4521 ( R1240_U204 , R1240_U130 , R1240_U4 );
nand NAND2_4522 ( R1240_U205 , R1240_U35 , R1240_U34 );
nand NAND2_4523 ( R1240_U206 , U3064 , R1240_U205 );
nand NAND2_4524 ( R1240_U207 , U3476 , R1240_U187 );
not NOT1_4525 ( R1240_U208 , R1240_U51 );
or OR2_4526 ( R1240_U209 , U3067 , U3480 );
or OR2_4527 ( R1240_U210 , U3068 , U3478 );
not NOT1_4528 ( R1240_U211 , R1240_U43 );
nand NAND2_4529 ( R1240_U212 , R1240_U44 , R1240_U43 );
nand NAND2_4530 ( R1240_U213 , U3067 , R1240_U212 );
nand NAND2_4531 ( R1240_U214 , U3480 , R1240_U211 );
nand NAND2_4532 ( R1240_U215 , R1240_U6 , R1240_U51 );
not NOT1_4533 ( R1240_U216 , R1240_U162 );
or OR2_4534 ( R1240_U217 , U3482 , U3081 );
nand NAND2_4535 ( R1240_U218 , R1240_U217 , R1240_U162 );
not NOT1_4536 ( R1240_U219 , R1240_U50 );
or OR2_4537 ( R1240_U220 , U3080 , U3484 );
or OR2_4538 ( R1240_U221 , U3478 , U3068 );
nand NAND2_4539 ( R1240_U222 , R1240_U221 , R1240_U51 );
nand NAND2_4540 ( R1240_U223 , R1240_U134 , R1240_U222 );
nand NAND2_4541 ( R1240_U224 , R1240_U208 , R1240_U43 );
nand NAND2_4542 ( R1240_U225 , U3480 , U3067 );
nand NAND2_4543 ( R1240_U226 , R1240_U135 , R1240_U224 );
or OR2_4544 ( R1240_U227 , U3068 , U3478 );
nand NAND2_4545 ( R1240_U228 , R1240_U202 , R1240_U198 );
nand NAND2_4546 ( R1240_U229 , U3065 , U3470 );
not NOT1_4547 ( R1240_U230 , R1240_U53 );
nand NAND2_4548 ( R1240_U231 , R1240_U201 , R1240_U5 );
nand NAND2_4549 ( R1240_U232 , R1240_U53 , R1240_U197 );
nand NAND2_4550 ( R1240_U233 , U3061 , U3472 );
not NOT1_4551 ( R1240_U234 , R1240_U52 );
or OR2_4552 ( R1240_U235 , U3474 , U3057 );
nand NAND2_4553 ( R1240_U236 , R1240_U235 , R1240_U52 );
nand NAND2_4554 ( R1240_U237 , R1240_U137 , R1240_U236 );
nand NAND2_4555 ( R1240_U238 , R1240_U234 , R1240_U34 );
nand NAND2_4556 ( R1240_U239 , U3476 , U3064 );
nand NAND2_4557 ( R1240_U240 , R1240_U138 , R1240_U238 );
or OR2_4558 ( R1240_U241 , U3057 , U3474 );
nand NAND2_4559 ( R1240_U242 , R1240_U201 , R1240_U198 );
not NOT1_4560 ( R1240_U243 , R1240_U163 );
nand NAND2_4561 ( R1240_U244 , U3061 , U3472 );
nand NAND4_4562 ( R1240_U245 , R1240_U428 , R1240_U427 , R1240_U36 , R1240_U39 );
nand NAND2_4563 ( R1240_U246 , R1240_U36 , R1240_U39 );
nand NAND2_4564 ( R1240_U247 , U3065 , U3470 );
nand NAND2_4565 ( R1240_U248 , R1240_U139 , R1240_U246 );
or OR2_4566 ( R1240_U249 , U3080 , U3484 );
or OR2_4567 ( R1240_U250 , U3059 , U3486 );
nand NAND2_4568 ( R1240_U251 , R1240_U194 , R1240_U7 );
nand NAND2_4569 ( R1240_U252 , U3059 , U3486 );
nand NAND2_4570 ( R1240_U253 , R1240_U140 , R1240_U251 );
or OR2_4571 ( R1240_U254 , U3486 , U3059 );
nand NAND2_4572 ( R1240_U255 , R1240_U254 , R1240_U253 );
not NOT1_4573 ( R1240_U256 , R1240_U184 );
or OR2_4574 ( R1240_U257 , U3077 , U3492 );
or OR2_4575 ( R1240_U258 , U3069 , U3490 );
nand NAND2_4576 ( R1240_U259 , R1240_U191 , R1240_U8 );
nand NAND2_4577 ( R1240_U260 , U3077 , U3492 );
nand NAND2_4578 ( R1240_U261 , R1240_U144 , R1240_U259 );
or OR2_4579 ( R1240_U262 , U3488 , U3060 );
or OR2_4580 ( R1240_U263 , U3492 , U3077 );
nand NAND2_4581 ( R1240_U264 , R1240_U13 , R1240_U184 );
nand NAND2_4582 ( R1240_U265 , R1240_U263 , R1240_U261 );
not NOT1_4583 ( R1240_U266 , R1240_U183 );
or OR2_4584 ( R1240_U267 , U3494 , U3076 );
nand NAND2_4585 ( R1240_U268 , U3076 , U3494 );
not NOT1_4586 ( R1240_U269 , R1240_U181 );
or OR2_4587 ( R1240_U270 , U3496 , U3071 );
nand NAND2_4588 ( R1240_U271 , U3071 , U3496 );
not NOT1_4589 ( R1240_U272 , R1240_U105 );
or OR2_4590 ( R1240_U273 , U3066 , U3500 );
or OR2_4591 ( R1240_U274 , U3070 , U3498 );
not NOT1_4592 ( R1240_U275 , R1240_U90 );
nand NAND2_4593 ( R1240_U276 , R1240_U91 , R1240_U90 );
nand NAND2_4594 ( R1240_U277 , U3066 , R1240_U276 );
nand NAND2_4595 ( R1240_U278 , U3500 , R1240_U275 );
nand NAND2_4596 ( R1240_U279 , R1240_U9 , R1240_U105 );
not NOT1_4597 ( R1240_U280 , R1240_U179 );
or OR2_4598 ( R1240_U281 , U3073 , U4037 );
or OR2_4599 ( R1240_U282 , U3078 , U3504 );
or OR2_4600 ( R1240_U283 , U3072 , U4036 );
not NOT1_4601 ( R1240_U284 , R1240_U80 );
nand NAND2_4602 ( R1240_U285 , U4037 , R1240_U284 );
nand NAND2_4603 ( R1240_U286 , R1240_U285 , R1240_U103 );
nand NAND2_4604 ( R1240_U287 , R1240_U80 , R1240_U81 );
nand NAND2_4605 ( R1240_U288 , R1240_U287 , R1240_U286 );
nand NAND2_4606 ( R1240_U289 , R1240_U192 , R1240_U11 );
nand NAND2_4607 ( R1240_U290 , U3072 , U4036 );
nand NAND3_4608 ( R1240_U291 , R1240_U289 , R1240_U288 , R1240_U290 );
or OR2_4609 ( R1240_U292 , U3502 , U3079 );
or OR2_4610 ( R1240_U293 , U4036 , U3072 );
nand NAND2_4611 ( R1240_U294 , R1240_U293 , R1240_U291 );
not NOT1_4612 ( R1240_U295 , R1240_U175 );
or OR2_4613 ( R1240_U296 , U4035 , U3058 );
nand NAND2_4614 ( R1240_U297 , U3058 , U4035 );
not NOT1_4615 ( R1240_U298 , R1240_U94 );
or OR2_4616 ( R1240_U299 , U4034 , U3063 );
nand NAND2_4617 ( R1240_U300 , R1240_U299 , R1240_U94 );
nand NAND2_4618 ( R1240_U301 , U3063 , U4034 );
not NOT1_4619 ( R1240_U302 , R1240_U172 );
or OR2_4620 ( R1240_U303 , U3055 , U4032 );
nand NAND2_4621 ( R1240_U304 , R1240_U193 , R1240_U185 );
or OR2_4622 ( R1240_U305 , U4033 , U3062 );
or OR2_4623 ( R1240_U306 , U4031 , U3054 );
nand NAND2_4624 ( R1240_U307 , R1240_U149 , R1240_U392 );
not NOT1_4625 ( R1240_U308 , R1240_U171 );
or OR2_4626 ( R1240_U309 , U4030 , U3050 );
nand NAND2_4627 ( R1240_U310 , U3050 , U4030 );
not NOT1_4628 ( R1240_U311 , R1240_U169 );
nand NAND2_4629 ( R1240_U312 , U4029 , R1240_U169 );
not NOT1_4630 ( R1240_U313 , R1240_U167 );
nand NAND2_4631 ( R1240_U314 , R1240_U305 , R1240_U172 );
not NOT1_4632 ( R1240_U315 , R1240_U100 );
or OR2_4633 ( R1240_U316 , U4032 , U3055 );
nand NAND2_4634 ( R1240_U317 , R1240_U316 , R1240_U100 );
nand NAND2_4635 ( R1240_U318 , R1240_U151 , R1240_U317 );
nand NAND2_4636 ( R1240_U319 , R1240_U315 , R1240_U190 );
nand NAND2_4637 ( R1240_U320 , U4031 , U3054 );
nand NAND2_4638 ( R1240_U321 , R1240_U152 , R1240_U319 );
or OR2_4639 ( R1240_U322 , U3055 , U4032 );
nand NAND2_4640 ( R1240_U323 , R1240_U292 , R1240_U179 );
not NOT1_4641 ( R1240_U324 , R1240_U104 );
nand NAND2_4642 ( R1240_U325 , R1240_U10 , R1240_U104 );
nand NAND2_4643 ( R1240_U326 , R1240_U153 , R1240_U325 );
nand NAND2_4644 ( R1240_U327 , R1240_U325 , R1240_U288 );
nand NAND2_4645 ( R1240_U328 , R1240_U480 , R1240_U327 );
or OR2_4646 ( R1240_U329 , U3504 , U3078 );
nand NAND2_4647 ( R1240_U330 , R1240_U329 , R1240_U104 );
nand NAND2_4648 ( R1240_U331 , R1240_U154 , R1240_U330 );
nand NAND2_4649 ( R1240_U332 , R1240_U324 , R1240_U80 );
nand NAND2_4650 ( R1240_U333 , U3073 , U4037 );
nand NAND2_4651 ( R1240_U334 , R1240_U155 , R1240_U332 );
or OR2_4652 ( R1240_U335 , U3468 , U3075 );
not NOT1_4653 ( R1240_U336 , R1240_U178 );
or OR2_4654 ( R1240_U337 , U3078 , U3504 );
or OR2_4655 ( R1240_U338 , U3498 , U3070 );
nand NAND2_4656 ( R1240_U339 , R1240_U338 , R1240_U105 );
nand NAND2_4657 ( R1240_U340 , R1240_U156 , R1240_U339 );
nand NAND2_4658 ( R1240_U341 , R1240_U272 , R1240_U90 );
nand NAND2_4659 ( R1240_U342 , U3500 , U3066 );
nand NAND2_4660 ( R1240_U343 , R1240_U157 , R1240_U341 );
or OR2_4661 ( R1240_U344 , U3070 , U3498 );
nand NAND2_4662 ( R1240_U345 , R1240_U262 , R1240_U184 );
not NOT1_4663 ( R1240_U346 , R1240_U106 );
or OR2_4664 ( R1240_U347 , U3490 , U3069 );
nand NAND2_4665 ( R1240_U348 , R1240_U347 , R1240_U106 );
nand NAND2_4666 ( R1240_U349 , R1240_U158 , R1240_U348 );
nand NAND2_4667 ( R1240_U350 , R1240_U346 , R1240_U189 );
nand NAND2_4668 ( R1240_U351 , U3077 , U3492 );
nand NAND2_4669 ( R1240_U352 , R1240_U159 , R1240_U350 );
or OR2_4670 ( R1240_U353 , U3069 , U3490 );
or OR2_4671 ( R1240_U354 , U3484 , U3080 );
nand NAND2_4672 ( R1240_U355 , R1240_U354 , R1240_U50 );
nand NAND2_4673 ( R1240_U356 , R1240_U160 , R1240_U355 );
nand NAND2_4674 ( R1240_U357 , R1240_U219 , R1240_U188 );
nand NAND2_4675 ( R1240_U358 , U3059 , U3486 );
nand NAND2_4676 ( R1240_U359 , R1240_U161 , R1240_U357 );
nand NAND2_4677 ( R1240_U360 , R1240_U220 , R1240_U188 );
nand NAND2_4678 ( R1240_U361 , R1240_U217 , R1240_U65 );
nand NAND2_4679 ( R1240_U362 , R1240_U227 , R1240_U43 );
nand NAND2_4680 ( R1240_U363 , R1240_U241 , R1240_U34 );
nand NAND2_4681 ( R1240_U364 , R1240_U244 , R1240_U197 );
nand NAND2_4682 ( R1240_U365 , R1240_U322 , R1240_U190 );
nand NAND2_4683 ( R1240_U366 , R1240_U305 , R1240_U60 );
nand NAND2_4684 ( R1240_U367 , R1240_U337 , R1240_U80 );
nand NAND2_4685 ( R1240_U368 , R1240_U292 , R1240_U84 );
nand NAND2_4686 ( R1240_U369 , R1240_U344 , R1240_U90 );
nand NAND2_4687 ( R1240_U370 , R1240_U353 , R1240_U189 );
nand NAND2_4688 ( R1240_U371 , R1240_U262 , R1240_U72 );
nand NAND2_4689 ( R1240_U372 , U4029 , U3051 );
nand NAND3_4690 ( R1240_U373 , R1240_U202 , R1240_U4 , R1240_U5 );
nand NAND3_4691 ( R1240_U374 , R1240_U5 , R1240_U4 , R1240_U201 );
not NOT1_4692 ( R1240_U375 , R1240_U45 );
not NOT1_4693 ( R1240_U376 , R1240_U102 );
nand NAND2_4694 ( R1240_U377 , R1240_U141 , R1240_U51 );
nand NAND2_4695 ( R1240_U378 , R1240_U12 , R1240_U45 );
nand NAND2_4696 ( R1240_U379 , R1240_U15 , R1240_U184 );
nand NAND2_4697 ( R1240_U380 , R1240_U268 , R1240_U265 );
not NOT1_4698 ( R1240_U381 , R1240_U77 );
nand NAND2_4699 ( R1240_U382 , R1240_U143 , R1240_U184 );
nand NAND2_4700 ( R1240_U383 , R1240_U381 , R1240_U270 );
nand NAND2_4701 ( R1240_U384 , R1240_U16 , R1240_U105 );
nand NAND2_4702 ( R1240_U385 , R1240_U14 , R1240_U102 );
not NOT1_4703 ( R1240_U386 , R1240_U101 );
not NOT1_4704 ( R1240_U387 , R1240_U97 );
nand NAND2_4705 ( R1240_U388 , R1240_U145 , R1240_U105 );
nand NAND2_4706 ( R1240_U389 , R1240_U101 , R1240_U296 );
nand NAND2_4707 ( R1240_U390 , U3054 , R1240_U303 );
nand NAND2_4708 ( R1240_U391 , U4031 , R1240_U303 );
nand NAND2_4709 ( R1240_U392 , R1240_U298 , R1240_U301 );
nand NAND3_4710 ( R1240_U393 , R1240_U193 , R1240_U185 , R1240_U309 );
nand NAND3_4711 ( R1240_U394 , R1240_U17 , R1240_U392 , R1240_U147 );
nand NAND2_4712 ( R1240_U395 , R1240_U387 , R1240_U309 );
nand NAND2_4713 ( R1240_U396 , R1240_U57 , R1240_U190 );
nand NAND2_4714 ( R1240_U397 , R1240_U56 , R1240_U190 );
nand NAND2_4715 ( R1240_U398 , U3080 , R1240_U49 );
nand NAND2_4716 ( R1240_U399 , U3484 , R1240_U48 );
nand NAND2_4717 ( R1240_U400 , R1240_U399 , R1240_U398 );
nand NAND2_4718 ( R1240_U401 , R1240_U360 , R1240_U50 );
nand NAND2_4719 ( R1240_U402 , R1240_U400 , R1240_U219 );
nand NAND2_4720 ( R1240_U403 , U3081 , R1240_U46 );
nand NAND2_4721 ( R1240_U404 , U3482 , R1240_U47 );
nand NAND2_4722 ( R1240_U405 , R1240_U404 , R1240_U403 );
nand NAND2_4723 ( R1240_U406 , R1240_U361 , R1240_U162 );
nand NAND2_4724 ( R1240_U407 , R1240_U216 , R1240_U405 );
nand NAND2_4725 ( R1240_U408 , U3067 , R1240_U44 );
nand NAND2_4726 ( R1240_U409 , U3480 , R1240_U42 );
nand NAND2_4727 ( R1240_U410 , U3068 , R1240_U40 );
nand NAND2_4728 ( R1240_U411 , U3478 , R1240_U41 );
nand NAND2_4729 ( R1240_U412 , R1240_U411 , R1240_U410 );
nand NAND2_4730 ( R1240_U413 , R1240_U362 , R1240_U51 );
nand NAND2_4731 ( R1240_U414 , R1240_U412 , R1240_U208 );
nand NAND2_4732 ( R1240_U415 , U3064 , R1240_U35 );
nand NAND2_4733 ( R1240_U416 , U3476 , R1240_U33 );
nand NAND2_4734 ( R1240_U417 , U3057 , R1240_U31 );
nand NAND2_4735 ( R1240_U418 , U3474 , R1240_U32 );
nand NAND2_4736 ( R1240_U419 , R1240_U418 , R1240_U417 );
nand NAND2_4737 ( R1240_U420 , R1240_U363 , R1240_U52 );
nand NAND2_4738 ( R1240_U421 , R1240_U419 , R1240_U234 );
nand NAND2_4739 ( R1240_U422 , U3061 , R1240_U29 );
nand NAND2_4740 ( R1240_U423 , U3472 , R1240_U30 );
nand NAND2_4741 ( R1240_U424 , R1240_U423 , R1240_U422 );
nand NAND2_4742 ( R1240_U425 , R1240_U364 , R1240_U163 );
nand NAND2_4743 ( R1240_U426 , R1240_U243 , R1240_U424 );
nand NAND2_4744 ( R1240_U427 , U3065 , R1240_U27 );
nand NAND2_4745 ( R1240_U428 , U3470 , R1240_U28 );
nand NAND2_4746 ( R1240_U429 , U3052 , R1240_U165 );
nand NAND2_4747 ( R1240_U430 , U4040 , R1240_U164 );
nand NAND2_4748 ( R1240_U431 , U3052 , R1240_U165 );
nand NAND2_4749 ( R1240_U432 , U4040 , R1240_U164 );
nand NAND2_4750 ( R1240_U433 , R1240_U432 , R1240_U431 );
nand NAND2_4751 ( R1240_U434 , R1240_U166 , R1240_U167 );
nand NAND2_4752 ( R1240_U435 , R1240_U313 , R1240_U433 );
nand NAND2_4753 ( R1240_U436 , U3051 , R1240_U99 );
nand NAND2_4754 ( R1240_U437 , U4029 , R1240_U98 );
nand NAND2_4755 ( R1240_U438 , U3051 , R1240_U99 );
nand NAND2_4756 ( R1240_U439 , U4029 , R1240_U98 );
nand NAND2_4757 ( R1240_U440 , R1240_U439 , R1240_U438 );
nand NAND2_4758 ( R1240_U441 , R1240_U168 , R1240_U169 );
nand NAND2_4759 ( R1240_U442 , R1240_U311 , R1240_U440 );
nand NAND2_4760 ( R1240_U443 , U3050 , R1240_U54 );
nand NAND2_4761 ( R1240_U444 , U4030 , R1240_U55 );
nand NAND2_4762 ( R1240_U445 , U3050 , R1240_U54 );
nand NAND2_4763 ( R1240_U446 , U4030 , R1240_U55 );
nand NAND2_4764 ( R1240_U447 , R1240_U446 , R1240_U445 );
nand NAND2_4765 ( R1240_U448 , R1240_U170 , R1240_U171 );
nand NAND2_4766 ( R1240_U449 , R1240_U308 , R1240_U447 );
nand NAND2_4767 ( R1240_U450 , U3054 , R1240_U57 );
nand NAND2_4768 ( R1240_U451 , U4031 , R1240_U56 );
nand NAND2_4769 ( R1240_U452 , U3055 , R1240_U95 );
nand NAND2_4770 ( R1240_U453 , U4032 , R1240_U96 );
nand NAND2_4771 ( R1240_U454 , R1240_U453 , R1240_U452 );
nand NAND2_4772 ( R1240_U455 , R1240_U365 , R1240_U100 );
nand NAND2_4773 ( R1240_U456 , R1240_U454 , R1240_U315 );
nand NAND2_4774 ( R1240_U457 , U3062 , R1240_U58 );
nand NAND2_4775 ( R1240_U458 , U4033 , R1240_U59 );
nand NAND2_4776 ( R1240_U459 , R1240_U458 , R1240_U457 );
nand NAND2_4777 ( R1240_U460 , R1240_U366 , R1240_U172 );
nand NAND2_4778 ( R1240_U461 , R1240_U302 , R1240_U459 );
nand NAND2_4779 ( R1240_U462 , U3063 , R1240_U92 );
nand NAND2_4780 ( R1240_U463 , U4034 , R1240_U93 );
nand NAND2_4781 ( R1240_U464 , U3063 , R1240_U92 );
nand NAND2_4782 ( R1240_U465 , U4034 , R1240_U93 );
nand NAND2_4783 ( R1240_U466 , R1240_U465 , R1240_U464 );
nand NAND2_4784 ( R1240_U467 , R1240_U173 , R1240_U94 );
nand NAND2_4785 ( R1240_U468 , R1240_U466 , R1240_U298 );
nand NAND2_4786 ( R1240_U469 , U3058 , R1240_U61 );
nand NAND2_4787 ( R1240_U470 , U4035 , R1240_U62 );
nand NAND2_4788 ( R1240_U471 , U3058 , R1240_U61 );
nand NAND2_4789 ( R1240_U472 , U4035 , R1240_U62 );
nand NAND2_4790 ( R1240_U473 , R1240_U472 , R1240_U471 );
nand NAND2_4791 ( R1240_U474 , R1240_U174 , R1240_U175 );
nand NAND2_4792 ( R1240_U475 , R1240_U295 , R1240_U473 );
nand NAND2_4793 ( R1240_U476 , U3072 , R1240_U85 );
nand NAND2_4794 ( R1240_U477 , U4036 , R1240_U86 );
nand NAND2_4795 ( R1240_U478 , U3072 , R1240_U85 );
nand NAND2_4796 ( R1240_U479 , U4036 , R1240_U86 );
nand NAND2_4797 ( R1240_U480 , R1240_U479 , R1240_U478 );
nand NAND2_4798 ( R1240_U481 , U3073 , R1240_U81 );
nand NAND2_4799 ( R1240_U482 , U4037 , R1240_U103 );
nand NAND2_4800 ( R1240_U483 , R1240_U199 , R1240_U178 );
nand NAND2_4801 ( R1240_U484 , R1240_U336 , R1240_U177 );
nand NAND2_4802 ( R1240_U485 , U3078 , R1240_U78 );
nand NAND2_4803 ( R1240_U486 , U3504 , R1240_U79 );
nand NAND2_4804 ( R1240_U487 , R1240_U486 , R1240_U485 );
nand NAND2_4805 ( R1240_U488 , R1240_U367 , R1240_U104 );
nand NAND2_4806 ( R1240_U489 , R1240_U487 , R1240_U324 );
nand NAND2_4807 ( R1240_U490 , U3079 , R1240_U82 );
nand NAND2_4808 ( R1240_U491 , U3502 , R1240_U83 );
nand NAND2_4809 ( R1240_U492 , R1240_U491 , R1240_U490 );
nand NAND2_4810 ( R1240_U493 , R1240_U368 , R1240_U179 );
nand NAND2_4811 ( R1240_U494 , R1240_U280 , R1240_U492 );
nand NAND2_4812 ( R1240_U495 , U3066 , R1240_U91 );
nand NAND2_4813 ( R1240_U496 , U3500 , R1240_U89 );
nand NAND2_4814 ( R1240_U497 , U3070 , R1240_U87 );
nand NAND2_4815 ( R1240_U498 , U3498 , R1240_U88 );
nand NAND2_4816 ( R1240_U499 , R1240_U498 , R1240_U497 );
nand NAND2_4817 ( R1240_U500 , R1240_U369 , R1240_U105 );
nand NAND2_4818 ( R1240_U501 , R1240_U499 , R1240_U272 );
nand NAND2_4819 ( R1240_U502 , U3071 , R1240_U63 );
nand NAND2_4820 ( R1240_U503 , U3496 , R1240_U64 );
nand NAND2_4821 ( R1240_U504 , U3071 , R1240_U63 );
nand NAND2_4822 ( R1240_U505 , U3496 , R1240_U64 );
nand NAND2_4823 ( R1240_U506 , R1240_U505 , R1240_U504 );
nand NAND2_4824 ( R1240_U507 , R1240_U180 , R1240_U181 );
nand NAND2_4825 ( R1240_U508 , R1240_U269 , R1240_U506 );
nand NAND2_4826 ( R1240_U509 , U3076 , R1240_U75 );
nand NAND2_4827 ( R1240_U510 , U3494 , R1240_U76 );
nand NAND2_4828 ( R1240_U511 , U3076 , R1240_U75 );
nand NAND2_4829 ( R1240_U512 , U3494 , R1240_U76 );
nand NAND2_4830 ( R1240_U513 , R1240_U512 , R1240_U511 );
nand NAND2_4831 ( R1240_U514 , R1240_U182 , R1240_U183 );
nand NAND2_4832 ( R1240_U515 , R1240_U266 , R1240_U513 );
nand NAND2_4833 ( R1240_U516 , U3077 , R1240_U73 );
nand NAND2_4834 ( R1240_U517 , U3492 , R1240_U74 );
nand NAND2_4835 ( R1240_U518 , U3069 , R1240_U68 );
nand NAND2_4836 ( R1240_U519 , U3490 , R1240_U69 );
nand NAND2_4837 ( R1240_U520 , R1240_U519 , R1240_U518 );
nand NAND2_4838 ( R1240_U521 , R1240_U370 , R1240_U106 );
nand NAND2_4839 ( R1240_U522 , R1240_U520 , R1240_U346 );
nand NAND2_4840 ( R1240_U523 , U3060 , R1240_U70 );
nand NAND2_4841 ( R1240_U524 , U3488 , R1240_U71 );
nand NAND2_4842 ( R1240_U525 , R1240_U524 , R1240_U523 );
nand NAND2_4843 ( R1240_U526 , R1240_U371 , R1240_U184 );
nand NAND2_4844 ( R1240_U527 , R1240_U256 , R1240_U525 );
nand NAND2_4845 ( R1240_U528 , U3059 , R1240_U66 );
nand NAND2_4846 ( R1240_U529 , U3486 , R1240_U67 );
nand NAND2_4847 ( R1240_U530 , U3074 , R1240_U37 );
nand NAND2_4848 ( R1240_U531 , U3464 , R1240_U38 );
and AND2_4849 ( R1162_U4 , R1162_U165 , R1162_U161 );
nand NAND2_4850 ( R1162_U5 , R1162_U84 , R1162_U166 );
not NOT1_4851 ( R1162_U6 , REG1_REG_0_ );
not NOT1_4852 ( R1162_U7 , U3453 );
not NOT1_4853 ( R1162_U8 , U3443 );
nand NAND2_4854 ( R1162_U9 , U3453 , REG1_REG_0_ );
not NOT1_4855 ( R1162_U10 , REG1_REG_1_ );
not NOT1_4856 ( R1162_U11 , REG1_REG_2_ );
not NOT1_4857 ( R1162_U12 , U3442 );
nand NAND2_4858 ( R1162_U13 , R1162_U103 , R1162_U102 );
not NOT1_4859 ( R1162_U14 , U3441 );
not NOT1_4860 ( R1162_U15 , REG1_REG_3_ );
not NOT1_4861 ( R1162_U16 , REG1_REG_4_ );
not NOT1_4862 ( R1162_U17 , U3440 );
nand NAND2_4863 ( R1162_U18 , R1162_U110 , R1162_U109 );
not NOT1_4864 ( R1162_U19 , U3439 );
not NOT1_4865 ( R1162_U20 , REG1_REG_5_ );
not NOT1_4866 ( R1162_U21 , REG1_REG_6_ );
not NOT1_4867 ( R1162_U22 , U3438 );
not NOT1_4868 ( R1162_U23 , REG1_REG_7_ );
not NOT1_4869 ( R1162_U24 , U3437 );
nand NAND2_4870 ( R1162_U25 , R1162_U121 , R1162_U120 );
not NOT1_4871 ( R1162_U26 , U3436 );
not NOT1_4872 ( R1162_U27 , REG1_REG_8_ );
not NOT1_4873 ( R1162_U28 , U3435 );
not NOT1_4874 ( R1162_U29 , REG1_REG_9_ );
nand NAND2_4875 ( R1162_U30 , R1162_U128 , R1162_U127 );
not NOT1_4876 ( R1162_U31 , U3452 );
not NOT1_4877 ( R1162_U32 , REG1_REG_10_ );
not NOT1_4878 ( R1162_U33 , REG1_REG_11_ );
not NOT1_4879 ( R1162_U34 , U3451 );
not NOT1_4880 ( R1162_U35 , REG1_REG_12_ );
not NOT1_4881 ( R1162_U36 , U3450 );
nand NAND2_4882 ( R1162_U37 , R1162_U139 , R1162_U138 );
not NOT1_4883 ( R1162_U38 , U3449 );
not NOT1_4884 ( R1162_U39 , REG1_REG_13_ );
nand NAND2_4885 ( R1162_U40 , R1162_U142 , R1162_U141 );
not NOT1_4886 ( R1162_U41 , U3448 );
not NOT1_4887 ( R1162_U42 , REG1_REG_14_ );
nand NAND2_4888 ( R1162_U43 , R1162_U145 , R1162_U144 );
not NOT1_4889 ( R1162_U44 , U3447 );
not NOT1_4890 ( R1162_U45 , REG1_REG_15_ );
not NOT1_4891 ( R1162_U46 , REG1_REG_16_ );
not NOT1_4892 ( R1162_U47 , U3446 );
not NOT1_4893 ( R1162_U48 , REG1_REG_17_ );
not NOT1_4894 ( R1162_U49 , U3445 );
not NOT1_4895 ( R1162_U50 , REG1_REG_18_ );
not NOT1_4896 ( R1162_U51 , U3444 );
nand NAND2_4897 ( R1162_U52 , R1162_U156 , R1162_U155 );
nand NAND2_4898 ( R1162_U53 , R1162_U290 , R1162_U289 );
nand NAND2_4899 ( R1162_U54 , R1162_U173 , R1162_U172 );
nand NAND2_4900 ( R1162_U55 , R1162_U179 , R1162_U178 );
nand NAND2_4901 ( R1162_U56 , R1162_U186 , R1162_U185 );
nand NAND2_4902 ( R1162_U57 , R1162_U193 , R1162_U192 );
nand NAND2_4903 ( R1162_U58 , R1162_U199 , R1162_U198 );
nand NAND2_4904 ( R1162_U59 , R1162_U206 , R1162_U205 );
nand NAND2_4905 ( R1162_U60 , R1162_U212 , R1162_U211 );
nand NAND2_4906 ( R1162_U61 , R1162_U219 , R1162_U218 );
nand NAND2_4907 ( R1162_U62 , R1162_U236 , R1162_U235 );
nand NAND2_4908 ( R1162_U63 , R1162_U243 , R1162_U242 );
nand NAND2_4909 ( R1162_U64 , R1162_U250 , R1162_U249 );
nand NAND2_4910 ( R1162_U65 , R1162_U256 , R1162_U255 );
nand NAND2_4911 ( R1162_U66 , R1162_U262 , R1162_U261 );
nand NAND2_4912 ( R1162_U67 , R1162_U268 , R1162_U267 );
nand NAND2_4913 ( R1162_U68 , R1162_U275 , R1162_U274 );
nand NAND2_4914 ( R1162_U69 , R1162_U282 , R1162_U281 );
nand NAND2_4915 ( R1162_U70 , R1162_U288 , R1162_U287 );
and AND3_4916 ( R1162_U71 , R1162_U226 , R1162_U225 , R1162_U160 );
and AND2_4917 ( R1162_U72 , R1162_U164 , R1162_U229 );
and AND2_4918 ( R1162_U73 , R1162_U168 , R1162_U167 );
nand NAND2_4919 ( R1162_U74 , R1162_U124 , R1162_U123 );
and AND2_4920 ( R1162_U75 , R1162_U181 , R1162_U180 );
nand NAND2_4921 ( R1162_U76 , R1162_U117 , R1162_U116 );
and AND2_4922 ( R1162_U77 , R1162_U188 , R1162_U187 );
nand NAND2_4923 ( R1162_U78 , R1162_U113 , R1162_U112 );
and AND2_4924 ( R1162_U79 , R1162_U201 , R1162_U200 );
nand NAND2_4925 ( R1162_U80 , R1162_U106 , R1162_U105 );
and AND2_4926 ( R1162_U81 , R1162_U214 , R1162_U213 );
nand NAND2_4927 ( R1162_U82 , R1162_U83 , R1162_U99 );
nand NAND2_4928 ( R1162_U83 , REG1_REG_1_ , R1162_U97 );
and AND2_4929 ( R1162_U84 , R1162_U224 , R1162_U223 );
not NOT1_4930 ( R1162_U85 , U3461 );
not NOT1_4931 ( R1162_U86 , REG1_REG_19_ );
and AND2_4932 ( R1162_U87 , R1162_U231 , R1162_U230 );
and AND2_4933 ( R1162_U88 , R1162_U238 , R1162_U237 );
nand NAND2_4934 ( R1162_U89 , R1162_U152 , R1162_U151 );
and AND2_4935 ( R1162_U90 , R1162_U245 , R1162_U244 );
nand NAND2_4936 ( R1162_U91 , R1162_U148 , R1162_U147 );
and AND2_4937 ( R1162_U92 , R1162_U270 , R1162_U269 );
nand NAND2_4938 ( R1162_U93 , R1162_U135 , R1162_U134 );
and AND2_4939 ( R1162_U94 , R1162_U277 , R1162_U276 );
nand NAND2_4940 ( R1162_U95 , R1162_U131 , R1162_U130 );
not NOT1_4941 ( R1162_U96 , R1162_U83 );
not NOT1_4942 ( R1162_U97 , R1162_U9 );
nand NAND2_4943 ( R1162_U98 , R1162_U10 , R1162_U9 );
nand NAND2_4944 ( R1162_U99 , U3443 , R1162_U98 );
not NOT1_4945 ( R1162_U100 , R1162_U82 );
or OR2_4946 ( R1162_U101 , REG1_REG_2_ , U3442 );
nand NAND2_4947 ( R1162_U102 , R1162_U101 , R1162_U82 );
nand NAND2_4948 ( R1162_U103 , U3442 , REG1_REG_2_ );
not NOT1_4949 ( R1162_U104 , R1162_U13 );
nand NAND2_4950 ( R1162_U105 , U3441 , R1162_U208 );
nand NAND2_4951 ( R1162_U106 , REG1_REG_3_ , R1162_U13 );
not NOT1_4952 ( R1162_U107 , R1162_U80 );
or OR2_4953 ( R1162_U108 , REG1_REG_4_ , U3440 );
nand NAND2_4954 ( R1162_U109 , R1162_U108 , R1162_U80 );
nand NAND2_4955 ( R1162_U110 , U3440 , REG1_REG_4_ );
not NOT1_4956 ( R1162_U111 , R1162_U18 );
nand NAND2_4957 ( R1162_U112 , U3439 , R1162_U195 );
nand NAND2_4958 ( R1162_U113 , REG1_REG_5_ , R1162_U18 );
not NOT1_4959 ( R1162_U114 , R1162_U78 );
or OR2_4960 ( R1162_U115 , REG1_REG_6_ , U3438 );
nand NAND2_4961 ( R1162_U116 , R1162_U115 , R1162_U78 );
nand NAND2_4962 ( R1162_U117 , U3438 , REG1_REG_6_ );
not NOT1_4963 ( R1162_U118 , R1162_U76 );
or OR2_4964 ( R1162_U119 , REG1_REG_7_ , U3437 );
nand NAND2_4965 ( R1162_U120 , R1162_U119 , R1162_U76 );
nand NAND2_4966 ( R1162_U121 , U3437 , REG1_REG_7_ );
not NOT1_4967 ( R1162_U122 , R1162_U25 );
nand NAND2_4968 ( R1162_U123 , U3436 , R1162_U175 );
nand NAND2_4969 ( R1162_U124 , REG1_REG_8_ , R1162_U25 );
not NOT1_4970 ( R1162_U125 , R1162_U74 );
or OR2_4971 ( R1162_U126 , REG1_REG_9_ , U3435 );
nand NAND2_4972 ( R1162_U127 , R1162_U126 , R1162_U74 );
nand NAND2_4973 ( R1162_U128 , REG1_REG_9_ , U3435 );
not NOT1_4974 ( R1162_U129 , R1162_U30 );
nand NAND2_4975 ( R1162_U130 , U3452 , R1162_U284 );
nand NAND2_4976 ( R1162_U131 , REG1_REG_10_ , R1162_U30 );
not NOT1_4977 ( R1162_U132 , R1162_U95 );
or OR2_4978 ( R1162_U133 , REG1_REG_11_ , U3451 );
nand NAND2_4979 ( R1162_U134 , R1162_U133 , R1162_U95 );
nand NAND2_4980 ( R1162_U135 , U3451 , REG1_REG_11_ );
not NOT1_4981 ( R1162_U136 , R1162_U93 );
or OR2_4982 ( R1162_U137 , REG1_REG_12_ , U3450 );
nand NAND2_4983 ( R1162_U138 , R1162_U137 , R1162_U93 );
nand NAND2_4984 ( R1162_U139 , U3450 , REG1_REG_12_ );
not NOT1_4985 ( R1162_U140 , R1162_U37 );
nand NAND2_4986 ( R1162_U141 , U3449 , R1162_U264 );
nand NAND2_4987 ( R1162_U142 , REG1_REG_13_ , R1162_U37 );
not NOT1_4988 ( R1162_U143 , R1162_U40 );
nand NAND2_4989 ( R1162_U144 , U3448 , R1162_U258 );
nand NAND2_4990 ( R1162_U145 , REG1_REG_14_ , R1162_U40 );
not NOT1_4991 ( R1162_U146 , R1162_U43 );
nand NAND2_4992 ( R1162_U147 , U3447 , R1162_U252 );
nand NAND2_4993 ( R1162_U148 , REG1_REG_15_ , R1162_U43 );
not NOT1_4994 ( R1162_U149 , R1162_U91 );
or OR2_4995 ( R1162_U150 , REG1_REG_16_ , U3446 );
nand NAND2_4996 ( R1162_U151 , R1162_U150 , R1162_U91 );
nand NAND2_4997 ( R1162_U152 , U3446 , REG1_REG_16_ );
not NOT1_4998 ( R1162_U153 , R1162_U89 );
or OR2_4999 ( R1162_U154 , REG1_REG_17_ , U3445 );
nand NAND2_5000 ( R1162_U155 , R1162_U154 , R1162_U89 );
nand NAND2_5001 ( R1162_U156 , U3445 , REG1_REG_17_ );
not NOT1_5002 ( R1162_U157 , R1162_U52 );
or OR2_5003 ( R1162_U158 , REG1_REG_18_ , U3444 );
nand NAND2_5004 ( R1162_U159 , R1162_U158 , R1162_U52 );
nand NAND2_5005 ( R1162_U160 , U3444 , REG1_REG_18_ );
nand NAND2_5006 ( R1162_U161 , R1162_U71 , R1162_U159 );
nand NAND2_5007 ( R1162_U162 , U3444 , REG1_REG_18_ );
nand NAND2_5008 ( R1162_U163 , R1162_U157 , R1162_U162 );
or OR2_5009 ( R1162_U164 , U3444 , REG1_REG_18_ );
nand NAND2_5010 ( R1162_U165 , R1162_U72 , R1162_U163 );
nand NAND2_5011 ( R1162_U166 , R1162_U222 , R1162_U10 );
nand NAND2_5012 ( R1162_U167 , U3435 , R1162_U29 );
nand NAND2_5013 ( R1162_U168 , REG1_REG_9_ , R1162_U28 );
nand NAND2_5014 ( R1162_U169 , U3435 , R1162_U29 );
nand NAND2_5015 ( R1162_U170 , REG1_REG_9_ , R1162_U28 );
nand NAND2_5016 ( R1162_U171 , R1162_U170 , R1162_U169 );
nand NAND2_5017 ( R1162_U172 , R1162_U73 , R1162_U74 );
nand NAND2_5018 ( R1162_U173 , R1162_U125 , R1162_U171 );
nand NAND2_5019 ( R1162_U174 , REG1_REG_8_ , R1162_U25 );
nand NAND2_5020 ( R1162_U175 , R1162_U122 , R1162_U27 );
nand NAND2_5021 ( R1162_U176 , REG1_REG_8_ , R1162_U25 );
nand NAND2_5022 ( R1162_U177 , R1162_U175 , R1162_U176 );
nand NAND3_5023 ( R1162_U178 , R1162_U175 , R1162_U174 , R1162_U26 );
nand NAND2_5024 ( R1162_U179 , R1162_U177 , U3436 );
nand NAND2_5025 ( R1162_U180 , U3437 , R1162_U23 );
nand NAND2_5026 ( R1162_U181 , REG1_REG_7_ , R1162_U24 );
nand NAND2_5027 ( R1162_U182 , U3437 , R1162_U23 );
nand NAND2_5028 ( R1162_U183 , REG1_REG_7_ , R1162_U24 );
nand NAND2_5029 ( R1162_U184 , R1162_U183 , R1162_U182 );
nand NAND2_5030 ( R1162_U185 , R1162_U75 , R1162_U76 );
nand NAND2_5031 ( R1162_U186 , R1162_U118 , R1162_U184 );
nand NAND2_5032 ( R1162_U187 , U3438 , R1162_U21 );
nand NAND2_5033 ( R1162_U188 , REG1_REG_6_ , R1162_U22 );
nand NAND2_5034 ( R1162_U189 , U3438 , R1162_U21 );
nand NAND2_5035 ( R1162_U190 , REG1_REG_6_ , R1162_U22 );
nand NAND2_5036 ( R1162_U191 , R1162_U190 , R1162_U189 );
nand NAND2_5037 ( R1162_U192 , R1162_U77 , R1162_U78 );
nand NAND2_5038 ( R1162_U193 , R1162_U114 , R1162_U191 );
nand NAND2_5039 ( R1162_U194 , REG1_REG_5_ , R1162_U18 );
nand NAND2_5040 ( R1162_U195 , R1162_U111 , R1162_U20 );
nand NAND2_5041 ( R1162_U196 , REG1_REG_5_ , R1162_U18 );
nand NAND2_5042 ( R1162_U197 , R1162_U195 , R1162_U196 );
nand NAND3_5043 ( R1162_U198 , R1162_U195 , R1162_U194 , R1162_U19 );
nand NAND2_5044 ( R1162_U199 , R1162_U197 , U3439 );
nand NAND2_5045 ( R1162_U200 , U3440 , R1162_U16 );
nand NAND2_5046 ( R1162_U201 , REG1_REG_4_ , R1162_U17 );
nand NAND2_5047 ( R1162_U202 , U3440 , R1162_U16 );
nand NAND2_5048 ( R1162_U203 , REG1_REG_4_ , R1162_U17 );
nand NAND2_5049 ( R1162_U204 , R1162_U203 , R1162_U202 );
nand NAND2_5050 ( R1162_U205 , R1162_U79 , R1162_U80 );
nand NAND2_5051 ( R1162_U206 , R1162_U107 , R1162_U204 );
nand NAND2_5052 ( R1162_U207 , REG1_REG_3_ , R1162_U13 );
nand NAND2_5053 ( R1162_U208 , R1162_U104 , R1162_U15 );
nand NAND2_5054 ( R1162_U209 , REG1_REG_3_ , R1162_U13 );
nand NAND2_5055 ( R1162_U210 , R1162_U208 , R1162_U209 );
nand NAND3_5056 ( R1162_U211 , R1162_U208 , R1162_U207 , R1162_U14 );
nand NAND2_5057 ( R1162_U212 , R1162_U210 , U3441 );
nand NAND2_5058 ( R1162_U213 , U3442 , R1162_U11 );
nand NAND2_5059 ( R1162_U214 , REG1_REG_2_ , R1162_U12 );
nand NAND2_5060 ( R1162_U215 , U3442 , R1162_U11 );
nand NAND2_5061 ( R1162_U216 , REG1_REG_2_ , R1162_U12 );
nand NAND2_5062 ( R1162_U217 , R1162_U216 , R1162_U215 );
nand NAND2_5063 ( R1162_U218 , R1162_U81 , R1162_U82 );
nand NAND2_5064 ( R1162_U219 , R1162_U100 , R1162_U217 );
nand NAND2_5065 ( R1162_U220 , U3443 , R1162_U9 );
nand NAND2_5066 ( R1162_U221 , R1162_U97 , R1162_U8 );
nand NAND2_5067 ( R1162_U222 , R1162_U221 , R1162_U220 );
nand NAND3_5068 ( R1162_U223 , REG1_REG_1_ , R1162_U9 , R1162_U8 );
nand NAND2_5069 ( R1162_U224 , R1162_U96 , U3443 );
nand NAND2_5070 ( R1162_U225 , U3461 , R1162_U86 );
nand NAND2_5071 ( R1162_U226 , REG1_REG_19_ , R1162_U85 );
nand NAND2_5072 ( R1162_U227 , U3461 , R1162_U86 );
nand NAND2_5073 ( R1162_U228 , REG1_REG_19_ , R1162_U85 );
nand NAND2_5074 ( R1162_U229 , R1162_U228 , R1162_U227 );
nand NAND2_5075 ( R1162_U230 , U3444 , R1162_U50 );
nand NAND2_5076 ( R1162_U231 , REG1_REG_18_ , R1162_U51 );
nand NAND2_5077 ( R1162_U232 , U3444 , R1162_U50 );
nand NAND2_5078 ( R1162_U233 , REG1_REG_18_ , R1162_U51 );
nand NAND2_5079 ( R1162_U234 , R1162_U233 , R1162_U232 );
nand NAND2_5080 ( R1162_U235 , R1162_U87 , R1162_U52 );
nand NAND2_5081 ( R1162_U236 , R1162_U234 , R1162_U157 );
nand NAND2_5082 ( R1162_U237 , U3445 , R1162_U48 );
nand NAND2_5083 ( R1162_U238 , REG1_REG_17_ , R1162_U49 );
nand NAND2_5084 ( R1162_U239 , U3445 , R1162_U48 );
nand NAND2_5085 ( R1162_U240 , REG1_REG_17_ , R1162_U49 );
nand NAND2_5086 ( R1162_U241 , R1162_U240 , R1162_U239 );
nand NAND2_5087 ( R1162_U242 , R1162_U88 , R1162_U89 );
nand NAND2_5088 ( R1162_U243 , R1162_U153 , R1162_U241 );
nand NAND2_5089 ( R1162_U244 , U3446 , R1162_U46 );
nand NAND2_5090 ( R1162_U245 , REG1_REG_16_ , R1162_U47 );
nand NAND2_5091 ( R1162_U246 , U3446 , R1162_U46 );
nand NAND2_5092 ( R1162_U247 , REG1_REG_16_ , R1162_U47 );
nand NAND2_5093 ( R1162_U248 , R1162_U247 , R1162_U246 );
nand NAND2_5094 ( R1162_U249 , R1162_U90 , R1162_U91 );
nand NAND2_5095 ( R1162_U250 , R1162_U149 , R1162_U248 );
nand NAND2_5096 ( R1162_U251 , REG1_REG_15_ , R1162_U43 );
nand NAND2_5097 ( R1162_U252 , R1162_U146 , R1162_U45 );
nand NAND2_5098 ( R1162_U253 , REG1_REG_15_ , R1162_U43 );
nand NAND2_5099 ( R1162_U254 , R1162_U252 , R1162_U253 );
nand NAND3_5100 ( R1162_U255 , R1162_U252 , R1162_U251 , R1162_U44 );
nand NAND2_5101 ( R1162_U256 , R1162_U254 , U3447 );
nand NAND2_5102 ( R1162_U257 , REG1_REG_14_ , R1162_U40 );
nand NAND2_5103 ( R1162_U258 , R1162_U143 , R1162_U42 );
nand NAND2_5104 ( R1162_U259 , REG1_REG_14_ , R1162_U40 );
nand NAND2_5105 ( R1162_U260 , R1162_U258 , R1162_U259 );
nand NAND3_5106 ( R1162_U261 , R1162_U258 , R1162_U257 , R1162_U41 );
nand NAND2_5107 ( R1162_U262 , R1162_U260 , U3448 );
nand NAND2_5108 ( R1162_U263 , REG1_REG_13_ , R1162_U37 );
nand NAND2_5109 ( R1162_U264 , R1162_U140 , R1162_U39 );
nand NAND2_5110 ( R1162_U265 , REG1_REG_13_ , R1162_U37 );
nand NAND2_5111 ( R1162_U266 , R1162_U264 , R1162_U265 );
nand NAND3_5112 ( R1162_U267 , R1162_U264 , R1162_U263 , R1162_U38 );
nand NAND2_5113 ( R1162_U268 , R1162_U266 , U3449 );
nand NAND2_5114 ( R1162_U269 , U3450 , R1162_U35 );
nand NAND2_5115 ( R1162_U270 , REG1_REG_12_ , R1162_U36 );
nand NAND2_5116 ( R1162_U271 , U3450 , R1162_U35 );
nand NAND2_5117 ( R1162_U272 , REG1_REG_12_ , R1162_U36 );
nand NAND2_5118 ( R1162_U273 , R1162_U272 , R1162_U271 );
nand NAND2_5119 ( R1162_U274 , R1162_U92 , R1162_U93 );
nand NAND2_5120 ( R1162_U275 , R1162_U136 , R1162_U273 );
nand NAND2_5121 ( R1162_U276 , U3451 , R1162_U33 );
nand NAND2_5122 ( R1162_U277 , REG1_REG_11_ , R1162_U34 );
nand NAND2_5123 ( R1162_U278 , U3451 , R1162_U33 );
nand NAND2_5124 ( R1162_U279 , REG1_REG_11_ , R1162_U34 );
nand NAND2_5125 ( R1162_U280 , R1162_U279 , R1162_U278 );
nand NAND2_5126 ( R1162_U281 , R1162_U94 , R1162_U95 );
nand NAND2_5127 ( R1162_U282 , R1162_U132 , R1162_U280 );
nand NAND2_5128 ( R1162_U283 , REG1_REG_10_ , R1162_U30 );
nand NAND2_5129 ( R1162_U284 , R1162_U129 , R1162_U32 );
nand NAND2_5130 ( R1162_U285 , REG1_REG_10_ , R1162_U30 );
nand NAND2_5131 ( R1162_U286 , R1162_U284 , R1162_U285 );
nand NAND3_5132 ( R1162_U287 , R1162_U284 , R1162_U283 , R1162_U31 );
nand NAND2_5133 ( R1162_U288 , R1162_U286 , U3452 );
nand NAND2_5134 ( R1162_U289 , U3453 , R1162_U6 );
nand NAND2_5135 ( R1162_U290 , REG1_REG_0_ , R1162_U7 );
and AND2_5136 ( R1117_U6 , R1117_U228 , R1117_U227 );
and AND2_5137 ( R1117_U7 , R1117_U208 , R1117_U261 );
and AND2_5138 ( R1117_U8 , R1117_U263 , R1117_U262 );
and AND2_5139 ( R1117_U9 , R1117_U209 , R1117_U272 );
and AND2_5140 ( R1117_U10 , R1117_U274 , R1117_U273 );
and AND2_5141 ( R1117_U11 , R1117_U186 , R1117_U290 );
and AND2_5142 ( R1117_U12 , R1117_U292 , R1117_U291 );
and AND2_5143 ( R1117_U13 , R1117_U304 , R1117_U211 );
and AND3_5144 ( R1117_U14 , R1117_U226 , R1117_U213 , R1117_U231 );
and AND2_5145 ( R1117_U15 , R1117_U236 , R1117_U214 );
and AND2_5146 ( R1117_U16 , R1117_U7 , R1117_U241 );
and AND2_5147 ( R1117_U17 , R1117_U9 , R1117_U277 );
and AND2_5148 ( R1117_U18 , R1117_U11 , R1117_U295 );
and AND2_5149 ( R1117_U19 , R1117_U16 , R1117_U268 );
and AND2_5150 ( R1117_U20 , R1117_U288 , R1117_U286 );
and AND2_5151 ( R1117_U21 , R1117_U20 , R1117_U18 );
and AND2_5152 ( R1117_U22 , R1117_U421 , R1117_U420 );
nand NAND2_5153 ( R1117_U23 , R1117_U328 , R1117_U331 );
nand NAND2_5154 ( R1117_U24 , R1117_U319 , R1117_U322 );
nand NAND4_5155 ( R1117_U25 , R1117_U383 , R1117_U382 , R1117_U454 , R1117_U453 );
nand NAND2_5156 ( R1117_U26 , R1117_U150 , R1117_U203 );
nand NAND2_5157 ( R1117_U27 , R1117_U259 , R1117_U371 );
nand NAND2_5158 ( R1117_U28 , R1117_U252 , R1117_U255 );
nand NAND2_5159 ( R1117_U29 , R1117_U244 , R1117_U246 );
nand NAND2_5160 ( R1117_U30 , R1117_U192 , R1117_U334 );
and AND2_5161 ( R1117_U31 , R1117_U373 , R1117_U379 );
not NOT1_5162 ( R1117_U32 , U3067 );
nand NAND2_5163 ( R1117_U33 , U3067 , R1117_U38 );
not NOT1_5164 ( R1117_U34 , U3081 );
not NOT1_5165 ( R1117_U35 , U3476 );
not NOT1_5166 ( R1117_U36 , U3478 );
not NOT1_5167 ( R1117_U37 , U3474 );
not NOT1_5168 ( R1117_U38 , U3480 );
not NOT1_5169 ( R1117_U39 , U3482 );
not NOT1_5170 ( R1117_U40 , U3065 );
nand NAND2_5171 ( R1117_U41 , U3065 , R1117_U43 );
not NOT1_5172 ( R1117_U42 , U3061 );
not NOT1_5173 ( R1117_U43 , U3470 );
not NOT1_5174 ( R1117_U44 , U3464 );
not NOT1_5175 ( R1117_U45 , U3075 );
not NOT1_5176 ( R1117_U46 , U3472 );
not NOT1_5177 ( R1117_U47 , U3068 );
not NOT1_5178 ( R1117_U48 , U3064 );
not NOT1_5179 ( R1117_U49 , U3057 );
nand NAND2_5180 ( R1117_U50 , U3057 , R1117_U37 );
nand NAND2_5181 ( R1117_U51 , R1117_U232 , R1117_U230 );
not NOT1_5182 ( R1117_U52 , U3484 );
not NOT1_5183 ( R1117_U53 , U3080 );
nand NAND2_5184 ( R1117_U54 , R1117_U51 , R1117_U233 );
nand NAND2_5185 ( R1117_U55 , R1117_U50 , R1117_U248 );
nand NAND3_5186 ( R1117_U56 , R1117_U220 , R1117_U204 , R1117_U335 );
not NOT1_5187 ( R1117_U57 , U4029 );
not NOT1_5188 ( R1117_U58 , U3054 );
nand NAND2_5189 ( R1117_U59 , U3054 , R1117_U99 );
not NOT1_5190 ( R1117_U60 , U3050 );
not NOT1_5191 ( R1117_U61 , U3062 );
not NOT1_5192 ( R1117_U62 , U4033 );
not NOT1_5193 ( R1117_U63 , U3063 );
not NOT1_5194 ( R1117_U64 , U3058 );
not NOT1_5195 ( R1117_U65 , U3072 );
not NOT1_5196 ( R1117_U66 , U4034 );
not NOT1_5197 ( R1117_U67 , U4035 );
nand NAND2_5198 ( R1117_U68 , U3072 , R1117_U69 );
not NOT1_5199 ( R1117_U69 , U4036 );
not NOT1_5200 ( R1117_U70 , U3073 );
not NOT1_5201 ( R1117_U71 , U3078 );
not NOT1_5202 ( R1117_U72 , U4037 );
nand NAND2_5203 ( R1117_U73 , U3078 , R1117_U74 );
not NOT1_5204 ( R1117_U74 , U3504 );
not NOT1_5205 ( R1117_U75 , U3079 );
not NOT1_5206 ( R1117_U76 , U3066 );
not NOT1_5207 ( R1117_U77 , U3500 );
not NOT1_5208 ( R1117_U78 , U3498 );
not NOT1_5209 ( R1117_U79 , U3496 );
not NOT1_5210 ( R1117_U80 , U3494 );
not NOT1_5211 ( R1117_U81 , U3077 );
not NOT1_5212 ( R1117_U82 , U3492 );
not NOT1_5213 ( R1117_U83 , U3490 );
not NOT1_5214 ( R1117_U84 , U3060 );
not NOT1_5215 ( R1117_U85 , U3059 );
not NOT1_5216 ( R1117_U86 , U3488 );
not NOT1_5217 ( R1117_U87 , U3486 );
nand NAND2_5218 ( R1117_U88 , U3080 , R1117_U52 );
not NOT1_5219 ( R1117_U89 , U3069 );
nand NAND2_5220 ( R1117_U90 , R1117_U339 , R1117_U268 );
not NOT1_5221 ( R1117_U91 , U3070 );
not NOT1_5222 ( R1117_U92 , U3071 );
not NOT1_5223 ( R1117_U93 , U3076 );
nand NAND2_5224 ( R1117_U94 , U3076 , R1117_U80 );
nand NAND2_5225 ( R1117_U95 , R1117_U278 , R1117_U276 );
not NOT1_5226 ( R1117_U96 , U3502 );
not NOT1_5227 ( R1117_U97 , U4032 );
not NOT1_5228 ( R1117_U98 , U3055 );
not NOT1_5229 ( R1117_U99 , U4031 );
not NOT1_5230 ( R1117_U100 , U4030 );
not NOT1_5231 ( R1117_U101 , U3051 );
nand NAND2_5232 ( R1117_U102 , R1117_U431 , R1117_U211 );
nand NAND2_5233 ( R1117_U103 , R1117_U346 , R1117_U297 );
nand NAND2_5234 ( R1117_U104 , R1117_U157 , R1117_U356 );
nand NAND2_5235 ( R1117_U105 , R1117_U344 , R1117_U289 );
nand NAND2_5236 ( R1117_U106 , R1117_U94 , R1117_U315 );
nand NAND2_5237 ( R1117_U107 , R1117_U360 , R1117_U88 );
not NOT1_5238 ( R1117_U108 , U3074 );
nand NAND2_5239 ( R1117_U109 , R1117_U428 , R1117_U427 );
nand NAND2_5240 ( R1117_U110 , R1117_U444 , R1117_U443 );
nand NAND2_5241 ( R1117_U111 , R1117_U449 , R1117_U448 );
nand NAND2_5242 ( R1117_U112 , R1117_U467 , R1117_U466 );
nand NAND2_5243 ( R1117_U113 , R1117_U472 , R1117_U471 );
nand NAND2_5244 ( R1117_U114 , R1117_U477 , R1117_U476 );
nand NAND2_5245 ( R1117_U115 , R1117_U482 , R1117_U481 );
nand NAND2_5246 ( R1117_U116 , R1117_U487 , R1117_U486 );
nand NAND2_5247 ( R1117_U117 , R1117_U503 , R1117_U502 );
nand NAND2_5248 ( R1117_U118 , R1117_U508 , R1117_U507 );
nand NAND2_5249 ( R1117_U119 , R1117_U387 , R1117_U386 );
nand NAND2_5250 ( R1117_U120 , R1117_U396 , R1117_U395 );
nand NAND2_5251 ( R1117_U121 , R1117_U403 , R1117_U402 );
nand NAND2_5252 ( R1117_U122 , R1117_U407 , R1117_U406 );
nand NAND2_5253 ( R1117_U123 , R1117_U416 , R1117_U415 );
nand NAND2_5254 ( R1117_U124 , R1117_U439 , R1117_U438 );
nand NAND2_5255 ( R1117_U125 , R1117_U458 , R1117_U457 );
nand NAND2_5256 ( R1117_U126 , R1117_U462 , R1117_U461 );
nand NAND2_5257 ( R1117_U127 , R1117_U494 , R1117_U493 );
nand NAND2_5258 ( R1117_U128 , R1117_U498 , R1117_U497 );
nand NAND2_5259 ( R1117_U129 , R1117_U515 , R1117_U514 );
and AND2_5260 ( R1117_U130 , R1117_U222 , R1117_U212 );
and AND2_5261 ( R1117_U131 , R1117_U225 , R1117_U224 );
and AND2_5262 ( R1117_U132 , R1117_U15 , R1117_U14 );
and AND2_5263 ( R1117_U133 , R1117_U239 , R1117_U238 );
and AND2_5264 ( R1117_U134 , R1117_U338 , R1117_U133 );
and AND3_5265 ( R1117_U135 , R1117_U389 , R1117_U388 , R1117_U33 );
and AND2_5266 ( R1117_U136 , R1117_U392 , R1117_U214 );
and AND2_5267 ( R1117_U137 , R1117_U254 , R1117_U6 );
and AND2_5268 ( R1117_U138 , R1117_U399 , R1117_U213 );
and AND3_5269 ( R1117_U139 , R1117_U409 , R1117_U408 , R1117_U41 );
and AND2_5270 ( R1117_U140 , R1117_U412 , R1117_U212 );
and AND2_5271 ( R1117_U141 , R1117_U270 , R1117_U19 );
and AND2_5272 ( R1117_U142 , R1117_U17 , R1117_U282 );
and AND2_5273 ( R1117_U143 , R1117_U343 , R1117_U283 );
and AND2_5274 ( R1117_U144 , R1117_U21 , R1117_U298 );
and AND2_5275 ( R1117_U145 , R1117_U348 , R1117_U299 );
and AND2_5276 ( R1117_U146 , R1117_U307 , R1117_U306 );
and AND2_5277 ( R1117_U147 , R1117_U419 , R1117_U308 );
and AND2_5278 ( R1117_U148 , R1117_U307 , R1117_U22 );
and AND3_5279 ( R1117_U149 , R1117_U148 , R1117_U306 , R1117_U309 );
and AND2_5280 ( R1117_U150 , R1117_U375 , R1117_U179 );
nand NAND2_5281 ( R1117_U151 , R1117_U425 , R1117_U424 );
and AND2_5282 ( R1117_U152 , R1117_U211 , R1117_U102 );
nand NAND2_5283 ( R1117_U153 , R1117_U441 , R1117_U440 );
nand NAND2_5284 ( R1117_U154 , R1117_U446 , R1117_U445 );
and AND2_5285 ( R1117_U155 , U3058 , R1117_U67 );
and AND2_5286 ( R1117_U156 , R1117_U20 , R1117_U295 );
and AND2_5287 ( R1117_U157 , R1117_U349 , R1117_U68 );
and AND2_5288 ( R1117_U158 , R1117_U12 , R1117_U311 );
nand NAND2_5289 ( R1117_U159 , R1117_U464 , R1117_U463 );
nand NAND2_5290 ( R1117_U160 , R1117_U469 , R1117_U468 );
nand NAND2_5291 ( R1117_U161 , R1117_U474 , R1117_U473 );
nand NAND2_5292 ( R1117_U162 , R1117_U479 , R1117_U478 );
nand NAND2_5293 ( R1117_U163 , R1117_U484 , R1117_U483 );
and AND2_5294 ( R1117_U164 , R1117_U321 , R1117_U10 );
and AND2_5295 ( R1117_U165 , R1117_U490 , R1117_U209 );
nand NAND2_5296 ( R1117_U166 , R1117_U500 , R1117_U499 );
nand NAND2_5297 ( R1117_U167 , R1117_U505 , R1117_U504 );
and AND2_5298 ( R1117_U168 , R1117_U330 , R1117_U8 );
and AND2_5299 ( R1117_U169 , R1117_U511 , R1117_U208 );
and AND2_5300 ( R1117_U170 , R1117_U385 , R1117_U384 );
nand NAND2_5301 ( R1117_U171 , R1117_U134 , R1117_U337 );
and AND2_5302 ( R1117_U172 , R1117_U394 , R1117_U393 );
and AND2_5303 ( R1117_U173 , R1117_U401 , R1117_U400 );
and AND2_5304 ( R1117_U174 , R1117_U405 , R1117_U404 );
nand NAND2_5305 ( R1117_U175 , R1117_U131 , R1117_U368 );
and AND2_5306 ( R1117_U176 , R1117_U414 , R1117_U413 );
not NOT1_5307 ( R1117_U177 , U4040 );
not NOT1_5308 ( R1117_U178 , U3052 );
and AND2_5309 ( R1117_U179 , R1117_U423 , R1117_U422 );
nand NAND2_5310 ( R1117_U180 , R1117_U146 , R1117_U376 );
and AND2_5311 ( R1117_U181 , R1117_U435 , R1117_U434 );
and AND2_5312 ( R1117_U182 , R1117_U437 , R1117_U436 );
nand NAND2_5313 ( R1117_U183 , R1117_U302 , R1117_U301 );
nand NAND2_5314 ( R1117_U184 , R1117_U145 , R1117_U358 );
nand NAND2_5315 ( R1117_U185 , R1117_U347 , R1117_U354 );
nand NAND2_5316 ( R1117_U186 , U4035 , R1117_U64 );
and AND2_5317 ( R1117_U187 , R1117_U456 , R1117_U455 );
and AND2_5318 ( R1117_U188 , R1117_U460 , R1117_U459 );
nand NAND2_5319 ( R1117_U189 , R1117_U345 , R1117_U352 );
nand NAND2_5320 ( R1117_U190 , R1117_U350 , R1117_U73 );
not NOT1_5321 ( R1117_U191 , U3468 );
nand NAND2_5322 ( R1117_U192 , U3464 , R1117_U108 );
nand NAND2_5323 ( R1117_U193 , R1117_U380 , R1117_U336 );
nand NAND2_5324 ( R1117_U194 , R1117_U143 , R1117_U342 );
nand NAND2_5325 ( R1117_U195 , R1117_U95 , R1117_U279 );
and AND2_5326 ( R1117_U196 , R1117_U492 , R1117_U491 );
and AND2_5327 ( R1117_U197 , R1117_U496 , R1117_U495 );
nand NAND3_5328 ( R1117_U198 , R1117_U341 , R1117_U271 , R1117_U366 );
nand NAND2_5329 ( R1117_U199 , R1117_U364 , R1117_U90 );
nand NAND2_5330 ( R1117_U200 , R1117_U362 , R1117_U267 );
and AND2_5331 ( R1117_U201 , R1117_U513 , R1117_U512 );
not NOT1_5332 ( R1117_U202 , R1117_U102 );
nand NAND2_5333 ( R1117_U203 , R1117_U147 , R1117_U180 );
nand NAND2_5334 ( R1117_U204 , R1117_U192 , R1117_U191 );
not NOT1_5335 ( R1117_U205 , R1117_U59 );
not NOT1_5336 ( R1117_U206 , R1117_U41 );
not NOT1_5337 ( R1117_U207 , R1117_U33 );
nand NAND2_5338 ( R1117_U208 , U3486 , R1117_U85 );
nand NAND2_5339 ( R1117_U209 , U3496 , R1117_U92 );
not NOT1_5340 ( R1117_U210 , R1117_U186 );
nand NAND2_5341 ( R1117_U211 , U4031 , R1117_U58 );
nand NAND2_5342 ( R1117_U212 , U3470 , R1117_U40 );
nand NAND2_5343 ( R1117_U213 , U3476 , R1117_U48 );
nand NAND2_5344 ( R1117_U214 , U3480 , R1117_U32 );
not NOT1_5345 ( R1117_U215 , R1117_U94 );
not NOT1_5346 ( R1117_U216 , R1117_U68 );
not NOT1_5347 ( R1117_U217 , R1117_U50 );
not NOT1_5348 ( R1117_U218 , R1117_U88 );
not NOT1_5349 ( R1117_U219 , R1117_U192 );
nand NAND2_5350 ( R1117_U220 , U3075 , R1117_U192 );
not NOT1_5351 ( R1117_U221 , R1117_U56 );
nand NAND2_5352 ( R1117_U222 , U3472 , R1117_U42 );
nand NAND2_5353 ( R1117_U223 , R1117_U42 , R1117_U41 );
nand NAND2_5354 ( R1117_U224 , R1117_U223 , R1117_U46 );
nand NAND2_5355 ( R1117_U225 , U3061 , R1117_U206 );
nand NAND2_5356 ( R1117_U226 , U3478 , R1117_U47 );
nand NAND2_5357 ( R1117_U227 , U3068 , R1117_U36 );
nand NAND2_5358 ( R1117_U228 , U3064 , R1117_U35 );
nand NAND2_5359 ( R1117_U229 , R1117_U217 , R1117_U213 );
nand NAND2_5360 ( R1117_U230 , R1117_U6 , R1117_U229 );
nand NAND2_5361 ( R1117_U231 , U3474 , R1117_U49 );
nand NAND2_5362 ( R1117_U232 , U3478 , R1117_U47 );
nand NAND2_5363 ( R1117_U233 , R1117_U14 , R1117_U175 );
not NOT1_5364 ( R1117_U234 , R1117_U51 );
not NOT1_5365 ( R1117_U235 , R1117_U54 );
nand NAND2_5366 ( R1117_U236 , U3482 , R1117_U34 );
nand NAND2_5367 ( R1117_U237 , R1117_U34 , R1117_U33 );
nand NAND2_5368 ( R1117_U238 , R1117_U237 , R1117_U39 );
nand NAND2_5369 ( R1117_U239 , U3081 , R1117_U207 );
not NOT1_5370 ( R1117_U240 , R1117_U171 );
nand NAND2_5371 ( R1117_U241 , U3484 , R1117_U53 );
nand NAND2_5372 ( R1117_U242 , R1117_U241 , R1117_U88 );
nand NAND2_5373 ( R1117_U243 , R1117_U235 , R1117_U33 );
nand NAND2_5374 ( R1117_U244 , R1117_U136 , R1117_U243 );
nand NAND2_5375 ( R1117_U245 , R1117_U54 , R1117_U214 );
nand NAND2_5376 ( R1117_U246 , R1117_U135 , R1117_U245 );
nand NAND2_5377 ( R1117_U247 , R1117_U33 , R1117_U214 );
nand NAND2_5378 ( R1117_U248 , R1117_U231 , R1117_U175 );
not NOT1_5379 ( R1117_U249 , R1117_U55 );
nand NAND2_5380 ( R1117_U250 , U3064 , R1117_U35 );
nand NAND2_5381 ( R1117_U251 , R1117_U249 , R1117_U250 );
nand NAND2_5382 ( R1117_U252 , R1117_U138 , R1117_U251 );
nand NAND2_5383 ( R1117_U253 , R1117_U55 , R1117_U213 );
nand NAND2_5384 ( R1117_U254 , U3478 , R1117_U47 );
nand NAND2_5385 ( R1117_U255 , R1117_U137 , R1117_U253 );
nand NAND2_5386 ( R1117_U256 , U3064 , R1117_U35 );
nand NAND2_5387 ( R1117_U257 , R1117_U213 , R1117_U256 );
nand NAND2_5388 ( R1117_U258 , R1117_U231 , R1117_U50 );
nand NAND2_5389 ( R1117_U259 , R1117_U140 , R1117_U372 );
nand NAND2_5390 ( R1117_U260 , R1117_U41 , R1117_U212 );
nand NAND2_5391 ( R1117_U261 , U3488 , R1117_U84 );
nand NAND2_5392 ( R1117_U262 , U3060 , R1117_U86 );
nand NAND2_5393 ( R1117_U263 , U3059 , R1117_U87 );
nand NAND2_5394 ( R1117_U264 , R1117_U218 , R1117_U7 );
nand NAND2_5395 ( R1117_U265 , R1117_U8 , R1117_U264 );
nand NAND2_5396 ( R1117_U266 , U3488 , R1117_U84 );
nand NAND2_5397 ( R1117_U267 , R1117_U266 , R1117_U265 );
nand NAND2_5398 ( R1117_U268 , U3490 , R1117_U89 );
nand NAND2_5399 ( R1117_U269 , U3069 , R1117_U83 );
nand NAND2_5400 ( R1117_U270 , U3492 , R1117_U81 );
nand NAND2_5401 ( R1117_U271 , U3077 , R1117_U82 );
nand NAND2_5402 ( R1117_U272 , U3498 , R1117_U91 );
nand NAND2_5403 ( R1117_U273 , U3070 , R1117_U78 );
nand NAND2_5404 ( R1117_U274 , U3071 , R1117_U79 );
nand NAND2_5405 ( R1117_U275 , R1117_U215 , R1117_U9 );
nand NAND2_5406 ( R1117_U276 , R1117_U10 , R1117_U275 );
nand NAND2_5407 ( R1117_U277 , U3494 , R1117_U93 );
nand NAND2_5408 ( R1117_U278 , U3498 , R1117_U91 );
nand NAND2_5409 ( R1117_U279 , R1117_U17 , R1117_U198 );
not NOT1_5410 ( R1117_U280 , R1117_U95 );
not NOT1_5411 ( R1117_U281 , R1117_U195 );
nand NAND2_5412 ( R1117_U282 , U3500 , R1117_U76 );
nand NAND2_5413 ( R1117_U283 , U3066 , R1117_U77 );
not NOT1_5414 ( R1117_U284 , R1117_U194 );
nand NAND2_5415 ( R1117_U285 , U3502 , R1117_U75 );
nand NAND2_5416 ( R1117_U286 , U3504 , R1117_U71 );
not NOT1_5417 ( R1117_U287 , R1117_U73 );
nand NAND2_5418 ( R1117_U288 , U4037 , R1117_U70 );
nand NAND2_5419 ( R1117_U289 , U3073 , R1117_U72 );
nand NAND2_5420 ( R1117_U290 , U4034 , R1117_U63 );
nand NAND2_5421 ( R1117_U291 , U3063 , R1117_U66 );
nand NAND2_5422 ( R1117_U292 , U3058 , R1117_U67 );
nand NAND2_5423 ( R1117_U293 , R1117_U216 , R1117_U11 );
nand NAND2_5424 ( R1117_U294 , R1117_U12 , R1117_U293 );
nand NAND2_5425 ( R1117_U295 , U4036 , R1117_U65 );
nand NAND2_5426 ( R1117_U296 , U4034 , R1117_U63 );
nand NAND2_5427 ( R1117_U297 , R1117_U296 , R1117_U294 );
nand NAND2_5428 ( R1117_U298 , U4033 , R1117_U61 );
nand NAND2_5429 ( R1117_U299 , U3062 , R1117_U62 );
nand NAND2_5430 ( R1117_U300 , U4032 , R1117_U98 );
nand NAND2_5431 ( R1117_U301 , R1117_U300 , R1117_U184 );
nand NAND2_5432 ( R1117_U302 , U3055 , R1117_U97 );
not NOT1_5433 ( R1117_U303 , R1117_U183 );
nand NAND2_5434 ( R1117_U304 , U4030 , R1117_U60 );
nand NAND2_5435 ( R1117_U305 , R1117_U60 , R1117_U59 );
nand NAND2_5436 ( R1117_U306 , R1117_U305 , R1117_U100 );
nand NAND2_5437 ( R1117_U307 , U3050 , R1117_U205 );
nand NAND2_5438 ( R1117_U308 , U4029 , R1117_U101 );
nand NAND2_5439 ( R1117_U309 , U3051 , R1117_U57 );
nand NAND2_5440 ( R1117_U310 , R1117_U59 , R1117_U211 );
nand NAND2_5441 ( R1117_U311 , U4034 , R1117_U63 );
nand NAND2_5442 ( R1117_U312 , U3058 , R1117_U67 );
nand NAND2_5443 ( R1117_U313 , R1117_U186 , R1117_U312 );
nand NAND2_5444 ( R1117_U314 , R1117_U295 , R1117_U68 );
nand NAND2_5445 ( R1117_U315 , R1117_U277 , R1117_U198 );
not NOT1_5446 ( R1117_U316 , R1117_U106 );
nand NAND2_5447 ( R1117_U317 , U3071 , R1117_U79 );
nand NAND2_5448 ( R1117_U318 , R1117_U316 , R1117_U317 );
nand NAND2_5449 ( R1117_U319 , R1117_U165 , R1117_U318 );
nand NAND2_5450 ( R1117_U320 , R1117_U106 , R1117_U209 );
nand NAND2_5451 ( R1117_U321 , U3498 , R1117_U91 );
nand NAND2_5452 ( R1117_U322 , R1117_U164 , R1117_U320 );
nand NAND2_5453 ( R1117_U323 , U3071 , R1117_U79 );
nand NAND2_5454 ( R1117_U324 , R1117_U209 , R1117_U323 );
nand NAND2_5455 ( R1117_U325 , R1117_U277 , R1117_U94 );
nand NAND2_5456 ( R1117_U326 , U3059 , R1117_U87 );
nand NAND2_5457 ( R1117_U327 , R1117_U361 , R1117_U326 );
nand NAND2_5458 ( R1117_U328 , R1117_U169 , R1117_U327 );
nand NAND2_5459 ( R1117_U329 , R1117_U107 , R1117_U208 );
nand NAND2_5460 ( R1117_U330 , U3488 , R1117_U84 );
nand NAND2_5461 ( R1117_U331 , R1117_U168 , R1117_U329 );
nand NAND2_5462 ( R1117_U332 , U3059 , R1117_U87 );
nand NAND2_5463 ( R1117_U333 , R1117_U208 , R1117_U332 );
nand NAND2_5464 ( R1117_U334 , U3074 , R1117_U44 );
nand NAND2_5465 ( R1117_U335 , U3075 , R1117_U191 );
nand NAND2_5466 ( R1117_U336 , U3079 , R1117_U96 );
nand NAND2_5467 ( R1117_U337 , R1117_U132 , R1117_U175 );
nand NAND2_5468 ( R1117_U338 , R1117_U234 , R1117_U15 );
nand NAND2_5469 ( R1117_U339 , R1117_U269 , R1117_U267 );
not NOT1_5470 ( R1117_U340 , R1117_U90 );
nand NAND2_5471 ( R1117_U341 , R1117_U340 , R1117_U270 );
nand NAND2_5472 ( R1117_U342 , R1117_U142 , R1117_U198 );
nand NAND2_5473 ( R1117_U343 , R1117_U280 , R1117_U282 );
nand NAND2_5474 ( R1117_U344 , R1117_U287 , R1117_U288 );
not NOT1_5475 ( R1117_U345 , R1117_U105 );
nand NAND2_5476 ( R1117_U346 , R1117_U18 , R1117_U105 );
not NOT1_5477 ( R1117_U347 , R1117_U103 );
nand NAND2_5478 ( R1117_U348 , R1117_U103 , R1117_U298 );
nand NAND2_5479 ( R1117_U349 , R1117_U105 , R1117_U295 );
nand NAND2_5480 ( R1117_U350 , R1117_U286 , R1117_U193 );
not NOT1_5481 ( R1117_U351 , R1117_U190 );
nand NAND2_5482 ( R1117_U352 , R1117_U20 , R1117_U193 );
not NOT1_5483 ( R1117_U353 , R1117_U189 );
nand NAND2_5484 ( R1117_U354 , R1117_U21 , R1117_U193 );
not NOT1_5485 ( R1117_U355 , R1117_U185 );
nand NAND2_5486 ( R1117_U356 , R1117_U156 , R1117_U193 );
not NOT1_5487 ( R1117_U357 , R1117_U104 );
nand NAND2_5488 ( R1117_U358 , R1117_U144 , R1117_U193 );
not NOT1_5489 ( R1117_U359 , R1117_U184 );
nand NAND2_5490 ( R1117_U360 , R1117_U241 , R1117_U171 );
not NOT1_5491 ( R1117_U361 , R1117_U107 );
nand NAND2_5492 ( R1117_U362 , R1117_U16 , R1117_U171 );
not NOT1_5493 ( R1117_U363 , R1117_U200 );
nand NAND2_5494 ( R1117_U364 , R1117_U19 , R1117_U171 );
not NOT1_5495 ( R1117_U365 , R1117_U199 );
nand NAND2_5496 ( R1117_U366 , R1117_U141 , R1117_U171 );
not NOT1_5497 ( R1117_U367 , R1117_U198 );
nand NAND2_5498 ( R1117_U368 , R1117_U130 , R1117_U56 );
not NOT1_5499 ( R1117_U369 , R1117_U175 );
nand NAND2_5500 ( R1117_U370 , R1117_U212 , R1117_U56 );
nand NAND2_5501 ( R1117_U371 , R1117_U139 , R1117_U370 );
nand NAND2_5502 ( R1117_U372 , R1117_U221 , R1117_U41 );
nand NAND2_5503 ( R1117_U373 , R1117_U152 , R1117_U183 );
nand NAND2_5504 ( R1117_U374 , R1117_U13 , R1117_U183 );
nand NAND2_5505 ( R1117_U375 , R1117_U149 , R1117_U374 );
nand NAND2_5506 ( R1117_U376 , R1117_U13 , R1117_U183 );
not NOT1_5507 ( R1117_U377 , R1117_U180 );
nand NAND2_5508 ( R1117_U378 , R1117_U202 , R1117_U183 );
nand NAND2_5509 ( R1117_U379 , R1117_U181 , R1117_U378 );
nand NAND2_5510 ( R1117_U380 , R1117_U285 , R1117_U194 );
not NOT1_5511 ( R1117_U381 , R1117_U193 );
nand NAND2_5512 ( R1117_U382 , R1117_U155 , R1117_U452 );
nand NAND2_5513 ( R1117_U383 , R1117_U158 , R1117_U357 );
nand NAND2_5514 ( R1117_U384 , U3484 , R1117_U53 );
nand NAND2_5515 ( R1117_U385 , U3080 , R1117_U52 );
nand NAND2_5516 ( R1117_U386 , R1117_U242 , R1117_U171 );
nand NAND2_5517 ( R1117_U387 , R1117_U240 , R1117_U170 );
nand NAND2_5518 ( R1117_U388 , U3482 , R1117_U34 );
nand NAND2_5519 ( R1117_U389 , U3081 , R1117_U39 );
nand NAND2_5520 ( R1117_U390 , U3482 , R1117_U34 );
nand NAND2_5521 ( R1117_U391 , U3081 , R1117_U39 );
nand NAND2_5522 ( R1117_U392 , R1117_U391 , R1117_U390 );
nand NAND2_5523 ( R1117_U393 , U3480 , R1117_U32 );
nand NAND2_5524 ( R1117_U394 , U3067 , R1117_U38 );
nand NAND2_5525 ( R1117_U395 , R1117_U247 , R1117_U54 );
nand NAND2_5526 ( R1117_U396 , R1117_U172 , R1117_U235 );
nand NAND2_5527 ( R1117_U397 , U3478 , R1117_U47 );
nand NAND2_5528 ( R1117_U398 , U3068 , R1117_U36 );
nand NAND2_5529 ( R1117_U399 , R1117_U398 , R1117_U397 );
nand NAND2_5530 ( R1117_U400 , U3476 , R1117_U48 );
nand NAND2_5531 ( R1117_U401 , U3064 , R1117_U35 );
nand NAND2_5532 ( R1117_U402 , R1117_U257 , R1117_U55 );
nand NAND2_5533 ( R1117_U403 , R1117_U173 , R1117_U249 );
nand NAND2_5534 ( R1117_U404 , U3474 , R1117_U49 );
nand NAND2_5535 ( R1117_U405 , U3057 , R1117_U37 );
nand NAND2_5536 ( R1117_U406 , R1117_U175 , R1117_U258 );
nand NAND2_5537 ( R1117_U407 , R1117_U369 , R1117_U174 );
nand NAND2_5538 ( R1117_U408 , U3472 , R1117_U42 );
nand NAND2_5539 ( R1117_U409 , U3061 , R1117_U46 );
nand NAND2_5540 ( R1117_U410 , U3472 , R1117_U42 );
nand NAND2_5541 ( R1117_U411 , U3061 , R1117_U46 );
nand NAND2_5542 ( R1117_U412 , R1117_U411 , R1117_U410 );
nand NAND2_5543 ( R1117_U413 , U3470 , R1117_U40 );
nand NAND2_5544 ( R1117_U414 , U3065 , R1117_U43 );
nand NAND2_5545 ( R1117_U415 , R1117_U260 , R1117_U56 );
nand NAND2_5546 ( R1117_U416 , R1117_U176 , R1117_U221 );
nand NAND2_5547 ( R1117_U417 , U4040 , R1117_U178 );
nand NAND2_5548 ( R1117_U418 , U3052 , R1117_U177 );
nand NAND2_5549 ( R1117_U419 , R1117_U418 , R1117_U417 );
nand NAND2_5550 ( R1117_U420 , U4040 , R1117_U178 );
nand NAND2_5551 ( R1117_U421 , U3052 , R1117_U177 );
nand NAND3_5552 ( R1117_U422 , U3051 , R1117_U419 , R1117_U57 );
nand NAND3_5553 ( R1117_U423 , R1117_U22 , R1117_U101 , U4029 );
nand NAND2_5554 ( R1117_U424 , U4029 , R1117_U101 );
nand NAND2_5555 ( R1117_U425 , U3051 , R1117_U57 );
not NOT1_5556 ( R1117_U426 , R1117_U151 );
nand NAND2_5557 ( R1117_U427 , R1117_U377 , R1117_U426 );
nand NAND2_5558 ( R1117_U428 , R1117_U151 , R1117_U180 );
nand NAND2_5559 ( R1117_U429 , U4030 , R1117_U60 );
nand NAND2_5560 ( R1117_U430 , U3050 , R1117_U100 );
nand NAND2_5561 ( R1117_U431 , R1117_U430 , R1117_U429 );
nand NAND2_5562 ( R1117_U432 , U4030 , R1117_U60 );
nand NAND2_5563 ( R1117_U433 , U3050 , R1117_U100 );
nand NAND3_5564 ( R1117_U434 , R1117_U433 , R1117_U432 , R1117_U59 );
nand NAND2_5565 ( R1117_U435 , R1117_U431 , R1117_U205 );
nand NAND2_5566 ( R1117_U436 , U4031 , R1117_U58 );
nand NAND2_5567 ( R1117_U437 , U3054 , R1117_U99 );
nand NAND2_5568 ( R1117_U438 , R1117_U310 , R1117_U183 );
nand NAND2_5569 ( R1117_U439 , R1117_U303 , R1117_U182 );
nand NAND2_5570 ( R1117_U440 , U4032 , R1117_U98 );
nand NAND2_5571 ( R1117_U441 , U3055 , R1117_U97 );
not NOT1_5572 ( R1117_U442 , R1117_U153 );
nand NAND2_5573 ( R1117_U443 , R1117_U359 , R1117_U442 );
nand NAND2_5574 ( R1117_U444 , R1117_U153 , R1117_U184 );
nand NAND2_5575 ( R1117_U445 , U4033 , R1117_U61 );
nand NAND2_5576 ( R1117_U446 , U3062 , R1117_U62 );
not NOT1_5577 ( R1117_U447 , R1117_U154 );
nand NAND2_5578 ( R1117_U448 , R1117_U355 , R1117_U447 );
nand NAND2_5579 ( R1117_U449 , R1117_U154 , R1117_U185 );
nand NAND2_5580 ( R1117_U450 , U4034 , R1117_U63 );
nand NAND2_5581 ( R1117_U451 , U3063 , R1117_U66 );
nand NAND2_5582 ( R1117_U452 , R1117_U451 , R1117_U450 );
nand NAND3_5583 ( R1117_U453 , R1117_U452 , R1117_U104 , R1117_U186 );
nand NAND3_5584 ( R1117_U454 , R1117_U12 , R1117_U311 , R1117_U210 );
nand NAND2_5585 ( R1117_U455 , U4035 , R1117_U64 );
nand NAND2_5586 ( R1117_U456 , U3058 , R1117_U67 );
nand NAND2_5587 ( R1117_U457 , R1117_U104 , R1117_U313 );
nand NAND2_5588 ( R1117_U458 , R1117_U187 , R1117_U357 );
nand NAND2_5589 ( R1117_U459 , U4036 , R1117_U65 );
nand NAND2_5590 ( R1117_U460 , U3072 , R1117_U69 );
nand NAND2_5591 ( R1117_U461 , R1117_U189 , R1117_U314 );
nand NAND2_5592 ( R1117_U462 , R1117_U353 , R1117_U188 );
nand NAND2_5593 ( R1117_U463 , U4037 , R1117_U70 );
nand NAND2_5594 ( R1117_U464 , U3073 , R1117_U72 );
not NOT1_5595 ( R1117_U465 , R1117_U159 );
nand NAND2_5596 ( R1117_U466 , R1117_U351 , R1117_U465 );
nand NAND2_5597 ( R1117_U467 , R1117_U159 , R1117_U190 );
nand NAND2_5598 ( R1117_U468 , U3468 , R1117_U45 );
nand NAND2_5599 ( R1117_U469 , U3075 , R1117_U191 );
not NOT1_5600 ( R1117_U470 , R1117_U160 );
nand NAND2_5601 ( R1117_U471 , R1117_U219 , R1117_U470 );
nand NAND2_5602 ( R1117_U472 , R1117_U160 , R1117_U192 );
nand NAND2_5603 ( R1117_U473 , U3504 , R1117_U71 );
nand NAND2_5604 ( R1117_U474 , U3078 , R1117_U74 );
not NOT1_5605 ( R1117_U475 , R1117_U161 );
nand NAND2_5606 ( R1117_U476 , R1117_U381 , R1117_U475 );
nand NAND2_5607 ( R1117_U477 , R1117_U161 , R1117_U193 );
nand NAND2_5608 ( R1117_U478 , U3502 , R1117_U75 );
nand NAND2_5609 ( R1117_U479 , U3079 , R1117_U96 );
not NOT1_5610 ( R1117_U480 , R1117_U162 );
nand NAND2_5611 ( R1117_U481 , R1117_U284 , R1117_U480 );
nand NAND2_5612 ( R1117_U482 , R1117_U162 , R1117_U194 );
nand NAND2_5613 ( R1117_U483 , U3500 , R1117_U76 );
nand NAND2_5614 ( R1117_U484 , U3066 , R1117_U77 );
not NOT1_5615 ( R1117_U485 , R1117_U163 );
nand NAND2_5616 ( R1117_U486 , R1117_U281 , R1117_U485 );
nand NAND2_5617 ( R1117_U487 , R1117_U163 , R1117_U195 );
nand NAND2_5618 ( R1117_U488 , U3498 , R1117_U91 );
nand NAND2_5619 ( R1117_U489 , U3070 , R1117_U78 );
nand NAND2_5620 ( R1117_U490 , R1117_U489 , R1117_U488 );
nand NAND2_5621 ( R1117_U491 , U3496 , R1117_U92 );
nand NAND2_5622 ( R1117_U492 , U3071 , R1117_U79 );
nand NAND2_5623 ( R1117_U493 , R1117_U324 , R1117_U106 );
nand NAND2_5624 ( R1117_U494 , R1117_U196 , R1117_U316 );
nand NAND2_5625 ( R1117_U495 , U3494 , R1117_U93 );
nand NAND2_5626 ( R1117_U496 , U3076 , R1117_U80 );
nand NAND2_5627 ( R1117_U497 , R1117_U198 , R1117_U325 );
nand NAND2_5628 ( R1117_U498 , R1117_U367 , R1117_U197 );
nand NAND2_5629 ( R1117_U499 , U3492 , R1117_U81 );
nand NAND2_5630 ( R1117_U500 , U3077 , R1117_U82 );
not NOT1_5631 ( R1117_U501 , R1117_U166 );
nand NAND2_5632 ( R1117_U502 , R1117_U365 , R1117_U501 );
nand NAND2_5633 ( R1117_U503 , R1117_U166 , R1117_U199 );
nand NAND2_5634 ( R1117_U504 , U3490 , R1117_U89 );
nand NAND2_5635 ( R1117_U505 , U3069 , R1117_U83 );
not NOT1_5636 ( R1117_U506 , R1117_U167 );
nand NAND2_5637 ( R1117_U507 , R1117_U363 , R1117_U506 );
nand NAND2_5638 ( R1117_U508 , R1117_U167 , R1117_U200 );
nand NAND2_5639 ( R1117_U509 , U3488 , R1117_U84 );
nand NAND2_5640 ( R1117_U510 , U3060 , R1117_U86 );
nand NAND2_5641 ( R1117_U511 , R1117_U510 , R1117_U509 );
nand NAND2_5642 ( R1117_U512 , U3486 , R1117_U85 );
nand NAND2_5643 ( R1117_U513 , U3059 , R1117_U87 );
nand NAND2_5644 ( R1117_U514 , R1117_U107 , R1117_U333 );
nand NAND2_5645 ( R1117_U515 , R1117_U201 , R1117_U361 );
and AND2_5646 ( R1375_U6 , R1375_U164 , R1375_U163 );
and AND2_5647 ( R1375_U7 , R1375_U172 , R1375_U173 );
and AND4_5648 ( R1375_U8 , R1375_U7 , R1375_U174 , R1375_U96 , R1375_U171 );
and AND2_5649 ( R1375_U9 , R1375_U97 , R1375_U8 );
and AND2_5650 ( R1375_U10 , R1375_U98 , R1375_U9 );
and AND2_5651 ( R1375_U11 , R1375_U181 , R1375_U182 );
and AND2_5652 ( R1375_U12 , R1375_U23 , R1375_U183 );
and AND3_5653 ( R1375_U13 , R1375_U185 , R1375_U184 , R1375_U186 );
and AND4_5654 ( R1375_U14 , R1375_U13 , R1375_U191 , R1375_U103 , R1375_U152 );
and AND4_5655 ( R1375_U15 , R1375_U154 , R1375_U153 , R1375_U155 , R1375_U157 );
and AND5_5656 ( R1375_U16 , R1375_U165 , R1375_U168 , R1375_U158 , R1375_U24 , R1375_U169 );
and AND4_5657 ( R1375_U17 , R1375_U10 , R1375_U179 , R1375_U24 , R1375_U109 );
and AND2_5658 ( R1375_U18 , R1375_U100 , R1375_U22 );
and AND2_5659 ( R1375_U19 , R1375_U10 , R1375_U165 );
and AND4_5660 ( R1375_U20 , U4030 , R1375_U155 , R1375_U154 , R1375_U34 );
and AND4_5661 ( R1375_U21 , U4029 , R1375_U154 , R1375_U155 , R1375_U27 );
and AND3_5662 ( R1375_U22 , R1375_U10 , R1375_U12 , R1375_U99 );
and AND4_5663 ( R1375_U23 , R1375_U11 , R1375_U180 , R1375_U179 , R1375_U178 );
and AND3_5664 ( R1375_U24 , R1375_U162 , R1375_U160 , R1375_U161 );
and AND2_5665 ( R1375_U25 , R1375_U100 , R1375_U165 );
nand NAND5_5666 ( R1375_U26 , R1375_U147 , R1375_U146 , R1375_U149 , R1375_U144 , R1375_U141 );
not NOT1_5667 ( R1375_U27 , U3051 );
not NOT1_5668 ( R1375_U28 , U3054 );
not NOT1_5669 ( R1375_U29 , U4032 );
not NOT1_5670 ( R1375_U30 , U4031 );
not NOT1_5671 ( R1375_U31 , U4038 );
not NOT1_5672 ( R1375_U32 , U3056 );
not NOT1_5673 ( R1375_U33 , U3052 );
not NOT1_5674 ( R1375_U34 , U3050 );
not NOT1_5675 ( R1375_U35 , U3057 );
not NOT1_5676 ( R1375_U36 , U3061 );
not NOT1_5677 ( R1375_U37 , U3065 );
not NOT1_5678 ( R1375_U38 , U3478 );
not NOT1_5679 ( R1375_U39 , U3064 );
not NOT1_5680 ( R1375_U40 , U4034 );
not NOT1_5681 ( R1375_U41 , U4033 );
not NOT1_5682 ( R1375_U42 , U3058 );
not NOT1_5683 ( R1375_U43 , U3077 );
not NOT1_5684 ( R1375_U44 , U3071 );
not NOT1_5685 ( R1375_U45 , U3073 );
not NOT1_5686 ( R1375_U46 , U3072 );
not NOT1_5687 ( R1375_U47 , U3502 );
not NOT1_5688 ( R1375_U48 , U3066 );
not NOT1_5689 ( R1375_U49 , U3079 );
not NOT1_5690 ( R1375_U50 , U3078 );
not NOT1_5691 ( R1375_U51 , U3070 );
not NOT1_5692 ( R1375_U52 , U3076 );
not NOT1_5693 ( R1375_U53 , U3069 );
not NOT1_5694 ( R1375_U54 , U3068 );
not NOT1_5695 ( R1375_U55 , U3490 );
not NOT1_5696 ( R1375_U56 , U3060 );
not NOT1_5697 ( R1375_U57 , U3059 );
not NOT1_5698 ( R1375_U58 , U3067 );
not NOT1_5699 ( R1375_U59 , U3081 );
not NOT1_5700 ( R1375_U60 , U3080 );
not NOT1_5701 ( R1375_U61 , U3063 );
not NOT1_5702 ( R1375_U62 , U3055 );
not NOT1_5703 ( R1375_U63 , U3062 );
not NOT1_5704 ( R1375_U64 , U3468 );
not NOT1_5705 ( R1375_U65 , U3075 );
not NOT1_5706 ( R1375_U66 , U3053 );
not NOT1_5707 ( R1375_U67 , U3488 );
not NOT1_5708 ( R1375_U68 , U3484 );
not NOT1_5709 ( R1375_U69 , U3496 );
not NOT1_5710 ( R1375_U70 , U3476 );
not NOT1_5711 ( R1375_U71 , U3472 );
not NOT1_5712 ( R1375_U72 , U3504 );
not NOT1_5713 ( R1375_U73 , U3492 );
not NOT1_5714 ( R1375_U74 , U3480 );
not NOT1_5715 ( R1375_U75 , U4037 );
not NOT1_5716 ( R1375_U76 , U3498 );
not NOT1_5717 ( R1375_U77 , U3494 );
not NOT1_5718 ( R1375_U78 , U3486 );
not NOT1_5719 ( R1375_U79 , U3482 );
not NOT1_5720 ( R1375_U80 , U3474 );
not NOT1_5721 ( R1375_U81 , U3470 );
not NOT1_5722 ( R1375_U82 , U4036 );
not NOT1_5723 ( R1375_U83 , U4035 );
not NOT1_5724 ( R1375_U84 , U3500 );
not NOT1_5725 ( R1375_U85 , U4030 );
not NOT1_5726 ( R1375_U86 , U4029 );
not NOT1_5727 ( R1375_U87 , U4040 );
not NOT1_5728 ( R1375_U88 , U4039 );
nand NAND2_5729 ( R1375_U89 , R1375_U198 , R1375_U197 );
and AND2_5730 ( R1375_U90 , U4032 , R1375_U62 );
and AND2_5731 ( R1375_U91 , U3063 , R1375_U40 );
and AND2_5732 ( R1375_U92 , U3064 , R1375_U70 );
and AND2_5733 ( R1375_U93 , U3058 , R1375_U83 );
and AND2_5734 ( R1375_U94 , U3060 , R1375_U67 );
and AND2_5735 ( R1375_U95 , U3066 , R1375_U84 );
and AND2_5736 ( R1375_U96 , R1375_U169 , R1375_U168 );
and AND2_5737 ( R1375_U97 , R1375_U175 , R1375_U167 );
and AND2_5738 ( R1375_U98 , R1375_U176 , R1375_U166 );
and AND2_5739 ( R1375_U99 , R1375_U165 , R1375_U152 );
and AND2_5740 ( R1375_U100 , R1375_U24 , R1375_U158 );
and AND2_5741 ( R1375_U101 , R1375_U15 , R1375_U65 );
and AND2_5742 ( R1375_U102 , R1375_U13 , U3468 );
and AND2_5743 ( R1375_U103 , R1375_U189 , R1375_U190 );
and AND2_5744 ( R1375_U104 , R1375_U192 , R1375_U156 );
and AND5_5745 ( R1375_U105 , R1375_U14 , R1375_U10 , R1375_U100 , R1375_U12 , R1375_U15 );
and AND2_5746 ( R1375_U106 , R1375_U156 , R1375_U53 );
and AND2_5747 ( R1375_U107 , R1375_U15 , R1375_U166 );
and AND2_5748 ( R1375_U108 , R1375_U15 , R1375_U56 );
and AND3_5749 ( R1375_U109 , R1375_U165 , R1375_U178 , R1375_U158 );
and AND2_5750 ( R1375_U110 , R1375_U15 , R1375_U60 );
and AND2_5751 ( R1375_U111 , R1375_U15 , R1375_U44 );
and AND2_5752 ( R1375_U112 , U3496 , R1375_U8 );
and AND2_5753 ( R1375_U113 , R1375_U156 , R1375_U54 );
and AND2_5754 ( R1375_U114 , U3478 , R1375_U15 );
and AND2_5755 ( R1375_U115 , R1375_U156 , R1375_U39 );
and AND5_5756 ( R1375_U116 , R1375_U19 , U3476 , R1375_U100 , R1375_U12 , R1375_U15 );
and AND3_5757 ( R1375_U117 , R1375_U184 , R1375_U36 , R1375_U156 );
and AND2_5758 ( R1375_U118 , R1375_U15 , R1375_U50 );
and AND2_5759 ( R1375_U119 , R1375_U15 , R1375_U43 );
and AND2_5760 ( R1375_U120 , R1375_U15 , R1375_U58 );
and AND2_5761 ( R1375_U121 , U3480 , R1375_U11 );
and AND3_5762 ( R1375_U122 , R1375_U169 , R1375_U45 , R1375_U156 );
and AND2_5763 ( R1375_U123 , R1375_U156 , R1375_U51 );
and AND2_5764 ( R1375_U124 , R1375_U15 , R1375_U171 );
and AND2_5765 ( R1375_U125 , U3498 , R1375_U7 );
and AND2_5766 ( R1375_U126 , R1375_U156 , R1375_U52 );
and AND2_5767 ( R1375_U127 , R1375_U15 , R1375_U167 );
and AND2_5768 ( R1375_U128 , U3494 , R1375_U8 );
and AND2_5769 ( R1375_U129 , R1375_U156 , R1375_U57 );
and AND5_5770 ( R1375_U130 , R1375_U19 , U3486 , R1375_U100 , R1375_U178 , R1375_U15 );
and AND3_5771 ( R1375_U131 , R1375_U181 , R1375_U59 , R1375_U156 );
and AND2_5772 ( R1375_U132 , R1375_U15 , R1375_U35 );
and AND4_5773 ( R1375_U133 , R1375_U185 , R1375_U184 , R1375_U37 , R1375_U156 );
and AND2_5774 ( R1375_U134 , R1375_U218 , R1375_U217 );
and AND2_5775 ( R1375_U135 , R1375_U219 , R1375_U156 );
and AND3_5776 ( R1375_U136 , R1375_U172 , R1375_U49 , R1375_U156 );
and AND2_5777 ( R1375_U137 , R1375_U15 , R1375_U48 );
and AND2_5778 ( R1375_U138 , U3500 , R1375_U7 );
and AND2_5779 ( R1375_U139 , R1375_U199 , R1375_U193 );
and AND3_5780 ( R1375_U140 , R1375_U201 , R1375_U202 , R1375_U200 );
and AND4_5781 ( R1375_U141 , R1375_U187 , R1375_U150 , R1375_U139 , R1375_U140 );
and AND2_5782 ( R1375_U142 , R1375_U204 , R1375_U203 );
and AND2_5783 ( R1375_U143 , R1375_U208 , R1375_U207 );
and AND5_5784 ( R1375_U144 , R1375_U206 , R1375_U205 , R1375_U142 , R1375_U143 , R1375_U209 );
and AND2_5785 ( R1375_U145 , R1375_U211 , R1375_U210 );
and AND3_5786 ( R1375_U146 , R1375_U213 , R1375_U212 , R1375_U145 );
and AND3_5787 ( R1375_U147 , R1375_U215 , R1375_U214 , R1375_U216 );
and AND3_5788 ( R1375_U148 , R1375_U224 , R1375_U225 , R1375_U223 );
and AND4_5789 ( R1375_U149 , R1375_U221 , R1375_U220 , R1375_U222 , R1375_U148 );
nand NAND3_5790 ( R1375_U150 , R1375_U196 , R1375_U15 , R1375_U156 );
nand NAND2_5791 ( R1375_U151 , U3478 , R1375_U54 );
nand NAND2_5792 ( R1375_U152 , R1375_U92 , R1375_U151 );
nand NAND2_5793 ( R1375_U153 , U4038 , R1375_U66 );
nand NAND2_5794 ( R1375_U154 , U3056 , R1375_U88 );
nand NAND2_5795 ( R1375_U155 , U3052 , R1375_U87 );
nand NAND2_5796 ( R1375_U156 , U3051 , R1375_U86 );
nand NAND2_5797 ( R1375_U157 , U3050 , R1375_U85 );
nand NAND2_5798 ( R1375_U158 , U3054 , R1375_U30 );
nand NAND2_5799 ( R1375_U159 , U4033 , R1375_U63 );
nand NAND2_5800 ( R1375_U160 , R1375_U91 , R1375_U159 );
nand NAND2_5801 ( R1375_U161 , U3055 , R1375_U29 );
nand NAND2_5802 ( R1375_U162 , U3062 , R1375_U41 );
nand NAND2_5803 ( R1375_U163 , U4034 , R1375_U61 );
nand NAND2_5804 ( R1375_U164 , U4033 , R1375_U63 );
nand NAND2_5805 ( R1375_U165 , R1375_U93 , R1375_U6 );
nand NAND2_5806 ( R1375_U166 , U3077 , R1375_U73 );
nand NAND2_5807 ( R1375_U167 , U3071 , R1375_U69 );
nand NAND2_5808 ( R1375_U168 , U3073 , R1375_U75 );
nand NAND2_5809 ( R1375_U169 , U3072 , R1375_U82 );
nand NAND2_5810 ( R1375_U170 , U3502 , R1375_U49 );
nand NAND2_5811 ( R1375_U171 , R1375_U95 , R1375_U170 );
nand NAND2_5812 ( R1375_U172 , U3078 , R1375_U72 );
nand NAND2_5813 ( R1375_U173 , U3079 , R1375_U47 );
nand NAND2_5814 ( R1375_U174 , U3070 , R1375_U76 );
nand NAND2_5815 ( R1375_U175 , U3076 , R1375_U77 );
nand NAND2_5816 ( R1375_U176 , U3069 , R1375_U55 );
nand NAND2_5817 ( R1375_U177 , U3490 , R1375_U53 );
nand NAND2_5818 ( R1375_U178 , R1375_U94 , R1375_U177 );
nand NAND2_5819 ( R1375_U179 , U3059 , R1375_U78 );
nand NAND2_5820 ( R1375_U180 , U3067 , R1375_U74 );
nand NAND2_5821 ( R1375_U181 , U3080 , R1375_U68 );
nand NAND2_5822 ( R1375_U182 , U3081 , R1375_U79 );
nand NAND2_5823 ( R1375_U183 , U3068 , R1375_U38 );
nand NAND2_5824 ( R1375_U184 , U3057 , R1375_U80 );
nand NAND2_5825 ( R1375_U185 , U3061 , R1375_U71 );
nand NAND2_5826 ( R1375_U186 , U3065 , R1375_U81 );
nand NAND4_5827 ( R1375_U187 , R1375_U102 , R1375_U18 , R1375_U156 , R1375_U101 );
nand NAND2_5828 ( R1375_U188 , U3464 , U3147 );
nand NAND2_5829 ( R1375_U189 , U3074 , R1375_U188 );
nand NAND2_5830 ( R1375_U190 , U3075 , R1375_U64 );
or OR2_5831 ( R1375_U191 , U3464 , U3147 );
nand NAND2_5832 ( R1375_U192 , U3058 , R1375_U83 );
nand NAND2_5833 ( R1375_U193 , R1375_U104 , R1375_U105 );
nand NAND2_5834 ( R1375_U194 , R1375_U90 , R1375_U158 );
nand NAND2_5835 ( R1375_U195 , U4031 , R1375_U28 );
nand NAND2_5836 ( R1375_U196 , R1375_U195 , R1375_U194 );
nand NAND3_5837 ( R1375_U197 , R1375_U154 , U4040 , R1375_U33 );
nand NAND2_5838 ( R1375_U198 , U4039 , R1375_U32 );
nand NAND2_5839 ( R1375_U199 , U3053 , R1375_U31 );
nand NAND5_5840 ( R1375_U200 , U3490 , R1375_U9 , R1375_U25 , R1375_U107 , R1375_U106 );
nand NAND5_5841 ( R1375_U201 , R1375_U19 , U3488 , R1375_U100 , R1375_U156 , R1375_U108 );
nand NAND4_5842 ( R1375_U202 , U3484 , R1375_U17 , R1375_U156 , R1375_U110 );
nand NAND4_5843 ( R1375_U203 , R1375_U112 , R1375_U25 , R1375_U156 , R1375_U111 );
nand NAND5_5844 ( R1375_U204 , R1375_U10 , R1375_U23 , R1375_U25 , R1375_U114 , R1375_U113 );
nand NAND2_5845 ( R1375_U205 , R1375_U115 , R1375_U116 );
nand NAND4_5846 ( R1375_U206 , R1375_U18 , U3472 , R1375_U15 , R1375_U117 );
nand NAND4_5847 ( R1375_U207 , U3504 , R1375_U16 , R1375_U156 , R1375_U118 );
nand NAND5_5848 ( R1375_U208 , U3492 , R1375_U9 , R1375_U25 , R1375_U156 , R1375_U119 );
nand NAND4_5849 ( R1375_U209 , R1375_U121 , R1375_U17 , R1375_U156 , R1375_U120 );
nand NAND4_5850 ( R1375_U210 , R1375_U25 , U4037 , R1375_U15 , R1375_U122 );
nand NAND4_5851 ( R1375_U211 , R1375_U125 , R1375_U16 , R1375_U124 , R1375_U123 );
nand NAND4_5852 ( R1375_U212 , R1375_U128 , R1375_U25 , R1375_U127 , R1375_U126 );
nand NAND2_5853 ( R1375_U213 , R1375_U129 , R1375_U130 );
nand NAND4_5854 ( R1375_U214 , R1375_U17 , U3482 , R1375_U15 , R1375_U131 );
nand NAND4_5855 ( R1375_U215 , U3474 , R1375_U18 , R1375_U156 , R1375_U132 );
nand NAND5_5856 ( R1375_U216 , U3470 , R1375_U22 , R1375_U100 , R1375_U15 , R1375_U133 );
nand NAND2_5857 ( R1375_U217 , U4036 , R1375_U46 );
nand NAND2_5858 ( R1375_U218 , U4035 , R1375_U42 );
nand NAND2_5859 ( R1375_U219 , R1375_U134 , R1375_U6 );
nand NAND3_5860 ( R1375_U220 , R1375_U25 , R1375_U15 , R1375_U135 );
nand NAND4_5861 ( R1375_U221 , U3502 , R1375_U16 , R1375_U15 , R1375_U136 );
nand NAND4_5862 ( R1375_U222 , R1375_U138 , R1375_U16 , R1375_U156 , R1375_U137 );
nand NAND3_5863 ( R1375_U223 , R1375_U20 , R1375_U153 , R1375_U156 );
nand NAND2_5864 ( R1375_U224 , R1375_U21 , R1375_U153 );
nand NAND2_5865 ( R1375_U225 , R1375_U89 , R1375_U153 );
and AND2_5866 ( R1352_U6 , U3056 , R1352_U7 );
not NOT1_5867 ( R1352_U7 , U3053 );
and AND2_5868 ( R1207_U6 , R1207_U231 , R1207_U230 );
and AND2_5869 ( R1207_U7 , R1207_U211 , R1207_U264 );
and AND2_5870 ( R1207_U8 , R1207_U266 , R1207_U265 );
and AND2_5871 ( R1207_U9 , R1207_U212 , R1207_U275 );
and AND2_5872 ( R1207_U10 , R1207_U277 , R1207_U276 );
and AND2_5873 ( R1207_U11 , R1207_U106 , R1207_U293 );
and AND2_5874 ( R1207_U12 , R1207_U295 , R1207_U294 );
and AND3_5875 ( R1207_U13 , R1207_U229 , R1207_U216 , R1207_U234 );
and AND2_5876 ( R1207_U14 , R1207_U239 , R1207_U217 );
and AND2_5877 ( R1207_U15 , R1207_U7 , R1207_U244 );
and AND2_5878 ( R1207_U16 , R1207_U9 , R1207_U280 );
and AND2_5879 ( R1207_U17 , R1207_U11 , R1207_U298 );
and AND2_5880 ( R1207_U18 , R1207_U15 , R1207_U271 );
and AND2_5881 ( R1207_U19 , R1207_U291 , R1207_U289 );
and AND2_5882 ( R1207_U20 , R1207_U19 , R1207_U17 );
and AND2_5883 ( R1207_U21 , R1207_U20 , R1207_U301 );
and AND2_5884 ( R1207_U22 , R1207_U457 , R1207_U106 );
and AND2_5885 ( R1207_U23 , R1207_U423 , R1207_U422 );
nand NAND2_5886 ( R1207_U24 , R1207_U334 , R1207_U337 );
nand NAND2_5887 ( R1207_U25 , R1207_U325 , R1207_U328 );
nand NAND5_5888 ( R1207_U26 , R1207_U459 , R1207_U458 , R1207_U388 , R1207_U387 , R1207_U359 );
and AND2_5889 ( R1207_U27 , R1207_U344 , R1207_U313 );
nand NAND3_5890 ( R1207_U28 , R1207_U182 , R1207_U206 , R1207_U343 );
nand NAND2_5891 ( R1207_U29 , R1207_U262 , R1207_U383 );
nand NAND2_5892 ( R1207_U30 , R1207_U255 , R1207_U258 );
nand NAND2_5893 ( R1207_U31 , R1207_U247 , R1207_U249 );
nand NAND2_5894 ( R1207_U32 , R1207_U195 , R1207_U340 );
not NOT1_5895 ( R1207_U33 , U3067 );
nand NAND2_5896 ( R1207_U34 , U3067 , R1207_U39 );
not NOT1_5897 ( R1207_U35 , U3081 );
not NOT1_5898 ( R1207_U36 , U3476 );
not NOT1_5899 ( R1207_U37 , U3478 );
not NOT1_5900 ( R1207_U38 , U3474 );
not NOT1_5901 ( R1207_U39 , U3480 );
not NOT1_5902 ( R1207_U40 , U3482 );
not NOT1_5903 ( R1207_U41 , U3065 );
nand NAND2_5904 ( R1207_U42 , U3065 , R1207_U44 );
not NOT1_5905 ( R1207_U43 , U3061 );
not NOT1_5906 ( R1207_U44 , U3470 );
not NOT1_5907 ( R1207_U45 , U3464 );
not NOT1_5908 ( R1207_U46 , U3075 );
not NOT1_5909 ( R1207_U47 , U3472 );
not NOT1_5910 ( R1207_U48 , U3068 );
not NOT1_5911 ( R1207_U49 , U3064 );
not NOT1_5912 ( R1207_U50 , U3057 );
nand NAND2_5913 ( R1207_U51 , U3057 , R1207_U38 );
nand NAND2_5914 ( R1207_U52 , R1207_U235 , R1207_U233 );
not NOT1_5915 ( R1207_U53 , U3484 );
not NOT1_5916 ( R1207_U54 , U3080 );
nand NAND2_5917 ( R1207_U55 , R1207_U52 , R1207_U236 );
nand NAND2_5918 ( R1207_U56 , R1207_U51 , R1207_U251 );
nand NAND3_5919 ( R1207_U57 , R1207_U223 , R1207_U207 , R1207_U341 );
not NOT1_5920 ( R1207_U58 , U4031 );
not NOT1_5921 ( R1207_U59 , U4030 );
not NOT1_5922 ( R1207_U60 , U3055 );
not NOT1_5923 ( R1207_U61 , U4032 );
not NOT1_5924 ( R1207_U62 , U3062 );
not NOT1_5925 ( R1207_U63 , U4033 );
not NOT1_5926 ( R1207_U64 , U3063 );
not NOT1_5927 ( R1207_U65 , U3058 );
not NOT1_5928 ( R1207_U66 , U3072 );
not NOT1_5929 ( R1207_U67 , U4034 );
not NOT1_5930 ( R1207_U68 , U4035 );
nand NAND2_5931 ( R1207_U69 , U3072 , R1207_U70 );
not NOT1_5932 ( R1207_U70 , U4036 );
not NOT1_5933 ( R1207_U71 , U3073 );
not NOT1_5934 ( R1207_U72 , U3078 );
not NOT1_5935 ( R1207_U73 , U4037 );
nand NAND2_5936 ( R1207_U74 , U3078 , R1207_U75 );
not NOT1_5937 ( R1207_U75 , U3504 );
not NOT1_5938 ( R1207_U76 , U3079 );
not NOT1_5939 ( R1207_U77 , U3066 );
not NOT1_5940 ( R1207_U78 , U3500 );
not NOT1_5941 ( R1207_U79 , U3498 );
not NOT1_5942 ( R1207_U80 , U3496 );
not NOT1_5943 ( R1207_U81 , U3494 );
not NOT1_5944 ( R1207_U82 , U3077 );
not NOT1_5945 ( R1207_U83 , U3492 );
not NOT1_5946 ( R1207_U84 , U3490 );
not NOT1_5947 ( R1207_U85 , U3060 );
not NOT1_5948 ( R1207_U86 , U3059 );
not NOT1_5949 ( R1207_U87 , U3488 );
not NOT1_5950 ( R1207_U88 , U3486 );
nand NAND2_5951 ( R1207_U89 , U3080 , R1207_U53 );
not NOT1_5952 ( R1207_U90 , U3069 );
nand NAND2_5953 ( R1207_U91 , R1207_U347 , R1207_U271 );
not NOT1_5954 ( R1207_U92 , U3070 );
not NOT1_5955 ( R1207_U93 , U3071 );
not NOT1_5956 ( R1207_U94 , U3076 );
nand NAND2_5957 ( R1207_U95 , U3076 , R1207_U81 );
nand NAND2_5958 ( R1207_U96 , R1207_U281 , R1207_U279 );
not NOT1_5959 ( R1207_U97 , U3502 );
not NOT1_5960 ( R1207_U98 , U3054 );
nand NAND2_5961 ( R1207_U99 , U3054 , R1207_U58 );
not NOT1_5962 ( R1207_U100 , U3050 );
not NOT1_5963 ( R1207_U101 , U4029 );
not NOT1_5964 ( R1207_U102 , U3051 );
nand NAND2_5965 ( R1207_U103 , R1207_U356 , R1207_U302 );
nand NAND2_5966 ( R1207_U104 , R1207_U354 , R1207_U300 );
nand NAND2_5967 ( R1207_U105 , R1207_U352 , R1207_U292 );
nand NAND2_5968 ( R1207_U106 , U4035 , R1207_U65 );
nand NAND2_5969 ( R1207_U107 , R1207_U95 , R1207_U321 );
nand NAND2_5970 ( R1207_U108 , R1207_U372 , R1207_U89 );
not NOT1_5971 ( R1207_U109 , U3074 );
nand NAND2_5972 ( R1207_U110 , R1207_U433 , R1207_U432 );
nand NAND2_5973 ( R1207_U111 , R1207_U449 , R1207_U448 );
nand NAND2_5974 ( R1207_U112 , R1207_U454 , R1207_U453 );
nand NAND2_5975 ( R1207_U113 , R1207_U472 , R1207_U471 );
nand NAND2_5976 ( R1207_U114 , R1207_U477 , R1207_U476 );
nand NAND2_5977 ( R1207_U115 , R1207_U482 , R1207_U481 );
nand NAND2_5978 ( R1207_U116 , R1207_U487 , R1207_U486 );
nand NAND2_5979 ( R1207_U117 , R1207_U492 , R1207_U491 );
nand NAND2_5980 ( R1207_U118 , R1207_U508 , R1207_U507 );
nand NAND2_5981 ( R1207_U119 , R1207_U513 , R1207_U512 );
nand NAND2_5982 ( R1207_U120 , R1207_U392 , R1207_U391 );
nand NAND2_5983 ( R1207_U121 , R1207_U401 , R1207_U400 );
nand NAND2_5984 ( R1207_U122 , R1207_U408 , R1207_U407 );
nand NAND2_5985 ( R1207_U123 , R1207_U412 , R1207_U411 );
nand NAND2_5986 ( R1207_U124 , R1207_U421 , R1207_U420 );
nand NAND2_5987 ( R1207_U125 , R1207_U444 , R1207_U443 );
nand NAND2_5988 ( R1207_U126 , R1207_U463 , R1207_U462 );
nand NAND2_5989 ( R1207_U127 , R1207_U467 , R1207_U466 );
nand NAND2_5990 ( R1207_U128 , R1207_U499 , R1207_U498 );
nand NAND2_5991 ( R1207_U129 , R1207_U503 , R1207_U502 );
nand NAND2_5992 ( R1207_U130 , R1207_U520 , R1207_U519 );
and AND2_5993 ( R1207_U131 , R1207_U225 , R1207_U215 );
and AND2_5994 ( R1207_U132 , R1207_U228 , R1207_U227 );
and AND2_5995 ( R1207_U133 , R1207_U14 , R1207_U13 );
and AND2_5996 ( R1207_U134 , R1207_U242 , R1207_U241 );
and AND2_5997 ( R1207_U135 , R1207_U346 , R1207_U134 );
and AND3_5998 ( R1207_U136 , R1207_U394 , R1207_U393 , R1207_U34 );
and AND2_5999 ( R1207_U137 , R1207_U397 , R1207_U217 );
and AND2_6000 ( R1207_U138 , R1207_U257 , R1207_U6 );
and AND2_6001 ( R1207_U139 , R1207_U404 , R1207_U216 );
and AND3_6002 ( R1207_U140 , R1207_U414 , R1207_U413 , R1207_U42 );
and AND2_6003 ( R1207_U141 , R1207_U417 , R1207_U215 );
and AND2_6004 ( R1207_U142 , R1207_U273 , R1207_U18 );
and AND2_6005 ( R1207_U143 , R1207_U16 , R1207_U285 );
and AND2_6006 ( R1207_U144 , R1207_U351 , R1207_U286 );
and AND2_6007 ( R1207_U145 , R1207_U21 , R1207_U303 );
and AND2_6008 ( R1207_U146 , R1207_U358 , R1207_U304 );
and AND2_6009 ( R1207_U147 , R1207_U305 , R1207_U214 );
and AND2_6010 ( R1207_U148 , R1207_U308 , R1207_U309 );
and AND2_6011 ( R1207_U149 , R1207_U311 , R1207_U426 );
and AND2_6012 ( R1207_U150 , R1207_U308 , R1207_U309 );
and AND2_6013 ( R1207_U151 , R1207_U23 , R1207_U312 );
nand NAND2_6014 ( R1207_U152 , R1207_U430 , R1207_U429 );
and AND2_6015 ( R1207_U153 , R1207_U436 , R1207_U214 );
and AND2_6016 ( R1207_U154 , R1207_U214 , R1207_U186 );
nand NAND2_6017 ( R1207_U155 , R1207_U446 , R1207_U445 );
nand NAND2_6018 ( R1207_U156 , R1207_U451 , R1207_U450 );
and AND2_6019 ( R1207_U157 , R1207_U22 , R1207_U298 );
and AND2_6020 ( R1207_U158 , R1207_U213 , R1207_U317 );
and AND2_6021 ( R1207_U159 , U3058 , R1207_U68 );
and AND2_6022 ( R1207_U160 , R1207_U19 , R1207_U298 );
and AND3_6023 ( R1207_U161 , R1207_U360 , R1207_U317 , R1207_U12 );
nand NAND2_6024 ( R1207_U162 , R1207_U469 , R1207_U468 );
nand NAND2_6025 ( R1207_U163 , R1207_U474 , R1207_U473 );
nand NAND2_6026 ( R1207_U164 , R1207_U479 , R1207_U478 );
nand NAND2_6027 ( R1207_U165 , R1207_U484 , R1207_U483 );
nand NAND2_6028 ( R1207_U166 , R1207_U489 , R1207_U488 );
and AND2_6029 ( R1207_U167 , R1207_U327 , R1207_U10 );
and AND2_6030 ( R1207_U168 , R1207_U495 , R1207_U212 );
nand NAND2_6031 ( R1207_U169 , R1207_U505 , R1207_U504 );
nand NAND2_6032 ( R1207_U170 , R1207_U510 , R1207_U509 );
and AND2_6033 ( R1207_U171 , R1207_U336 , R1207_U8 );
and AND2_6034 ( R1207_U172 , R1207_U516 , R1207_U211 );
and AND2_6035 ( R1207_U173 , R1207_U390 , R1207_U389 );
nand NAND2_6036 ( R1207_U174 , R1207_U135 , R1207_U345 );
and AND2_6037 ( R1207_U175 , R1207_U399 , R1207_U398 );
and AND2_6038 ( R1207_U176 , R1207_U406 , R1207_U405 );
and AND2_6039 ( R1207_U177 , R1207_U410 , R1207_U409 );
nand NAND2_6040 ( R1207_U178 , R1207_U132 , R1207_U380 );
and AND2_6041 ( R1207_U179 , R1207_U419 , R1207_U418 );
not NOT1_6042 ( R1207_U180 , U4040 );
not NOT1_6043 ( R1207_U181 , U3052 );
and AND2_6044 ( R1207_U182 , R1207_U428 , R1207_U427 );
nand NAND2_6045 ( R1207_U183 , R1207_U148 , R1207_U306 );
and AND2_6046 ( R1207_U184 , R1207_U440 , R1207_U439 );
and AND2_6047 ( R1207_U185 , R1207_U442 , R1207_U441 );
nand NAND2_6048 ( R1207_U186 , R1207_U146 , R1207_U370 );
nand NAND2_6049 ( R1207_U187 , R1207_U357 , R1207_U367 );
nand NAND2_6050 ( R1207_U188 , R1207_U355 , R1207_U365 );
and AND2_6051 ( R1207_U189 , R1207_U461 , R1207_U460 );
nand NAND2_6052 ( R1207_U190 , R1207_U69 , R1207_U315 );
and AND2_6053 ( R1207_U191 , R1207_U465 , R1207_U464 );
nand NAND2_6054 ( R1207_U192 , R1207_U353 , R1207_U363 );
nand NAND2_6055 ( R1207_U193 , R1207_U361 , R1207_U74 );
not NOT1_6056 ( R1207_U194 , U3468 );
nand NAND2_6057 ( R1207_U195 , U3464 , R1207_U109 );
nand NAND2_6058 ( R1207_U196 , R1207_U385 , R1207_U342 );
nand NAND2_6059 ( R1207_U197 , R1207_U144 , R1207_U350 );
nand NAND2_6060 ( R1207_U198 , R1207_U96 , R1207_U282 );
and AND2_6061 ( R1207_U199 , R1207_U497 , R1207_U496 );
and AND2_6062 ( R1207_U200 , R1207_U501 , R1207_U500 );
nand NAND3_6063 ( R1207_U201 , R1207_U349 , R1207_U274 , R1207_U378 );
nand NAND2_6064 ( R1207_U202 , R1207_U376 , R1207_U91 );
nand NAND2_6065 ( R1207_U203 , R1207_U374 , R1207_U270 );
and AND2_6066 ( R1207_U204 , R1207_U518 , R1207_U517 );
nand NAND2_6067 ( R1207_U205 , R1207_U153 , R1207_U186 );
nand NAND2_6068 ( R1207_U206 , R1207_U149 , R1207_U183 );
nand NAND2_6069 ( R1207_U207 , R1207_U195 , R1207_U194 );
not NOT1_6070 ( R1207_U208 , R1207_U99 );
not NOT1_6071 ( R1207_U209 , R1207_U42 );
not NOT1_6072 ( R1207_U210 , R1207_U34 );
nand NAND2_6073 ( R1207_U211 , U3486 , R1207_U86 );
nand NAND2_6074 ( R1207_U212 , U3496 , R1207_U93 );
not NOT1_6075 ( R1207_U213 , R1207_U106 );
nand NAND2_6076 ( R1207_U214 , U4031 , R1207_U98 );
nand NAND2_6077 ( R1207_U215 , U3470 , R1207_U41 );
nand NAND2_6078 ( R1207_U216 , U3476 , R1207_U49 );
nand NAND2_6079 ( R1207_U217 , U3480 , R1207_U33 );
not NOT1_6080 ( R1207_U218 , R1207_U95 );
not NOT1_6081 ( R1207_U219 , R1207_U69 );
not NOT1_6082 ( R1207_U220 , R1207_U51 );
not NOT1_6083 ( R1207_U221 , R1207_U89 );
not NOT1_6084 ( R1207_U222 , R1207_U195 );
nand NAND2_6085 ( R1207_U223 , U3075 , R1207_U195 );
not NOT1_6086 ( R1207_U224 , R1207_U57 );
nand NAND2_6087 ( R1207_U225 , U3472 , R1207_U43 );
nand NAND2_6088 ( R1207_U226 , R1207_U43 , R1207_U42 );
nand NAND2_6089 ( R1207_U227 , R1207_U226 , R1207_U47 );
nand NAND2_6090 ( R1207_U228 , U3061 , R1207_U209 );
nand NAND2_6091 ( R1207_U229 , U3478 , R1207_U48 );
nand NAND2_6092 ( R1207_U230 , U3068 , R1207_U37 );
nand NAND2_6093 ( R1207_U231 , U3064 , R1207_U36 );
nand NAND2_6094 ( R1207_U232 , R1207_U220 , R1207_U216 );
nand NAND2_6095 ( R1207_U233 , R1207_U6 , R1207_U232 );
nand NAND2_6096 ( R1207_U234 , U3474 , R1207_U50 );
nand NAND2_6097 ( R1207_U235 , U3478 , R1207_U48 );
nand NAND2_6098 ( R1207_U236 , R1207_U13 , R1207_U178 );
not NOT1_6099 ( R1207_U237 , R1207_U52 );
not NOT1_6100 ( R1207_U238 , R1207_U55 );
nand NAND2_6101 ( R1207_U239 , U3482 , R1207_U35 );
nand NAND2_6102 ( R1207_U240 , R1207_U35 , R1207_U34 );
nand NAND2_6103 ( R1207_U241 , R1207_U240 , R1207_U40 );
nand NAND2_6104 ( R1207_U242 , U3081 , R1207_U210 );
not NOT1_6105 ( R1207_U243 , R1207_U174 );
nand NAND2_6106 ( R1207_U244 , U3484 , R1207_U54 );
nand NAND2_6107 ( R1207_U245 , R1207_U244 , R1207_U89 );
nand NAND2_6108 ( R1207_U246 , R1207_U238 , R1207_U34 );
nand NAND2_6109 ( R1207_U247 , R1207_U137 , R1207_U246 );
nand NAND2_6110 ( R1207_U248 , R1207_U55 , R1207_U217 );
nand NAND2_6111 ( R1207_U249 , R1207_U136 , R1207_U248 );
nand NAND2_6112 ( R1207_U250 , R1207_U34 , R1207_U217 );
nand NAND2_6113 ( R1207_U251 , R1207_U234 , R1207_U178 );
not NOT1_6114 ( R1207_U252 , R1207_U56 );
nand NAND2_6115 ( R1207_U253 , U3064 , R1207_U36 );
nand NAND2_6116 ( R1207_U254 , R1207_U252 , R1207_U253 );
nand NAND2_6117 ( R1207_U255 , R1207_U139 , R1207_U254 );
nand NAND2_6118 ( R1207_U256 , R1207_U56 , R1207_U216 );
nand NAND2_6119 ( R1207_U257 , U3478 , R1207_U48 );
nand NAND2_6120 ( R1207_U258 , R1207_U138 , R1207_U256 );
nand NAND2_6121 ( R1207_U259 , U3064 , R1207_U36 );
nand NAND2_6122 ( R1207_U260 , R1207_U216 , R1207_U259 );
nand NAND2_6123 ( R1207_U261 , R1207_U234 , R1207_U51 );
nand NAND2_6124 ( R1207_U262 , R1207_U141 , R1207_U384 );
nand NAND2_6125 ( R1207_U263 , R1207_U42 , R1207_U215 );
nand NAND2_6126 ( R1207_U264 , U3488 , R1207_U85 );
nand NAND2_6127 ( R1207_U265 , U3060 , R1207_U87 );
nand NAND2_6128 ( R1207_U266 , U3059 , R1207_U88 );
nand NAND2_6129 ( R1207_U267 , R1207_U221 , R1207_U7 );
nand NAND2_6130 ( R1207_U268 , R1207_U8 , R1207_U267 );
nand NAND2_6131 ( R1207_U269 , U3488 , R1207_U85 );
nand NAND2_6132 ( R1207_U270 , R1207_U269 , R1207_U268 );
nand NAND2_6133 ( R1207_U271 , U3490 , R1207_U90 );
nand NAND2_6134 ( R1207_U272 , U3069 , R1207_U84 );
nand NAND2_6135 ( R1207_U273 , U3492 , R1207_U82 );
nand NAND2_6136 ( R1207_U274 , U3077 , R1207_U83 );
nand NAND2_6137 ( R1207_U275 , U3498 , R1207_U92 );
nand NAND2_6138 ( R1207_U276 , U3070 , R1207_U79 );
nand NAND2_6139 ( R1207_U277 , U3071 , R1207_U80 );
nand NAND2_6140 ( R1207_U278 , R1207_U218 , R1207_U9 );
nand NAND2_6141 ( R1207_U279 , R1207_U10 , R1207_U278 );
nand NAND2_6142 ( R1207_U280 , U3494 , R1207_U94 );
nand NAND2_6143 ( R1207_U281 , U3498 , R1207_U92 );
nand NAND2_6144 ( R1207_U282 , R1207_U16 , R1207_U201 );
not NOT1_6145 ( R1207_U283 , R1207_U96 );
not NOT1_6146 ( R1207_U284 , R1207_U198 );
nand NAND2_6147 ( R1207_U285 , U3500 , R1207_U77 );
nand NAND2_6148 ( R1207_U286 , U3066 , R1207_U78 );
not NOT1_6149 ( R1207_U287 , R1207_U197 );
nand NAND2_6150 ( R1207_U288 , U3502 , R1207_U76 );
nand NAND2_6151 ( R1207_U289 , U3504 , R1207_U72 );
not NOT1_6152 ( R1207_U290 , R1207_U74 );
nand NAND2_6153 ( R1207_U291 , U4037 , R1207_U71 );
nand NAND2_6154 ( R1207_U292 , U3073 , R1207_U73 );
nand NAND2_6155 ( R1207_U293 , U4034 , R1207_U64 );
nand NAND2_6156 ( R1207_U294 , U3063 , R1207_U67 );
nand NAND2_6157 ( R1207_U295 , U3058 , R1207_U68 );
nand NAND2_6158 ( R1207_U296 , R1207_U219 , R1207_U11 );
nand NAND2_6159 ( R1207_U297 , R1207_U12 , R1207_U296 );
nand NAND2_6160 ( R1207_U298 , U4036 , R1207_U66 );
nand NAND2_6161 ( R1207_U299 , U4034 , R1207_U64 );
nand NAND2_6162 ( R1207_U300 , R1207_U299 , R1207_U297 );
nand NAND2_6163 ( R1207_U301 , U4033 , R1207_U62 );
nand NAND2_6164 ( R1207_U302 , U3062 , R1207_U63 );
nand NAND2_6165 ( R1207_U303 , U4032 , R1207_U60 );
nand NAND2_6166 ( R1207_U304 , U3055 , R1207_U61 );
nand NAND2_6167 ( R1207_U305 , U4030 , R1207_U100 );
nand NAND2_6168 ( R1207_U306 , R1207_U147 , R1207_U186 );
nand NAND2_6169 ( R1207_U307 , R1207_U100 , R1207_U99 );
nand NAND2_6170 ( R1207_U308 , R1207_U307 , R1207_U59 );
nand NAND2_6171 ( R1207_U309 , U3050 , R1207_U208 );
not NOT1_6172 ( R1207_U310 , R1207_U183 );
nand NAND2_6173 ( R1207_U311 , U4029 , R1207_U102 );
nand NAND2_6174 ( R1207_U312 , U3051 , R1207_U101 );
nand NAND2_6175 ( R1207_U313 , R1207_U154 , R1207_U205 );
nand NAND2_6176 ( R1207_U314 , R1207_U99 , R1207_U214 );
nand NAND2_6177 ( R1207_U315 , R1207_U298 , R1207_U192 );
not NOT1_6178 ( R1207_U316 , R1207_U190 );
nand NAND2_6179 ( R1207_U317 , U4034 , R1207_U64 );
nand NAND2_6180 ( R1207_U318 , U3058 , R1207_U68 );
nand NAND2_6181 ( R1207_U319 , R1207_U106 , R1207_U318 );
nand NAND2_6182 ( R1207_U320 , R1207_U298 , R1207_U69 );
nand NAND2_6183 ( R1207_U321 , R1207_U280 , R1207_U201 );
not NOT1_6184 ( R1207_U322 , R1207_U107 );
nand NAND2_6185 ( R1207_U323 , U3071 , R1207_U80 );
nand NAND2_6186 ( R1207_U324 , R1207_U322 , R1207_U323 );
nand NAND2_6187 ( R1207_U325 , R1207_U168 , R1207_U324 );
nand NAND2_6188 ( R1207_U326 , R1207_U107 , R1207_U212 );
nand NAND2_6189 ( R1207_U327 , U3498 , R1207_U92 );
nand NAND2_6190 ( R1207_U328 , R1207_U167 , R1207_U326 );
nand NAND2_6191 ( R1207_U329 , U3071 , R1207_U80 );
nand NAND2_6192 ( R1207_U330 , R1207_U212 , R1207_U329 );
nand NAND2_6193 ( R1207_U331 , R1207_U280 , R1207_U95 );
nand NAND2_6194 ( R1207_U332 , U3059 , R1207_U88 );
nand NAND2_6195 ( R1207_U333 , R1207_U373 , R1207_U332 );
nand NAND2_6196 ( R1207_U334 , R1207_U172 , R1207_U333 );
nand NAND2_6197 ( R1207_U335 , R1207_U108 , R1207_U211 );
nand NAND2_6198 ( R1207_U336 , U3488 , R1207_U85 );
nand NAND2_6199 ( R1207_U337 , R1207_U171 , R1207_U335 );
nand NAND2_6200 ( R1207_U338 , U3059 , R1207_U88 );
nand NAND2_6201 ( R1207_U339 , R1207_U211 , R1207_U338 );
nand NAND2_6202 ( R1207_U340 , U3074 , R1207_U45 );
nand NAND2_6203 ( R1207_U341 , U3075 , R1207_U194 );
nand NAND2_6204 ( R1207_U342 , U3079 , R1207_U97 );
nand NAND3_6205 ( R1207_U343 , R1207_U150 , R1207_U306 , R1207_U151 );
nand NAND2_6206 ( R1207_U344 , R1207_U184 , R1207_U205 );
nand NAND2_6207 ( R1207_U345 , R1207_U133 , R1207_U178 );
nand NAND2_6208 ( R1207_U346 , R1207_U237 , R1207_U14 );
nand NAND2_6209 ( R1207_U347 , R1207_U272 , R1207_U270 );
not NOT1_6210 ( R1207_U348 , R1207_U91 );
nand NAND2_6211 ( R1207_U349 , R1207_U348 , R1207_U273 );
nand NAND2_6212 ( R1207_U350 , R1207_U143 , R1207_U201 );
nand NAND2_6213 ( R1207_U351 , R1207_U283 , R1207_U285 );
nand NAND2_6214 ( R1207_U352 , R1207_U290 , R1207_U291 );
not NOT1_6215 ( R1207_U353 , R1207_U105 );
nand NAND2_6216 ( R1207_U354 , R1207_U17 , R1207_U105 );
not NOT1_6217 ( R1207_U355 , R1207_U104 );
nand NAND2_6218 ( R1207_U356 , R1207_U104 , R1207_U301 );
not NOT1_6219 ( R1207_U357 , R1207_U103 );
nand NAND2_6220 ( R1207_U358 , R1207_U103 , R1207_U303 );
nand NAND2_6221 ( R1207_U359 , R1207_U157 , R1207_U192 );
nand NAND2_6222 ( R1207_U360 , R1207_U105 , R1207_U298 );
nand NAND2_6223 ( R1207_U361 , R1207_U289 , R1207_U196 );
not NOT1_6224 ( R1207_U362 , R1207_U193 );
nand NAND2_6225 ( R1207_U363 , R1207_U19 , R1207_U196 );
not NOT1_6226 ( R1207_U364 , R1207_U192 );
nand NAND2_6227 ( R1207_U365 , R1207_U20 , R1207_U196 );
not NOT1_6228 ( R1207_U366 , R1207_U188 );
nand NAND2_6229 ( R1207_U367 , R1207_U21 , R1207_U196 );
not NOT1_6230 ( R1207_U368 , R1207_U187 );
nand NAND2_6231 ( R1207_U369 , R1207_U160 , R1207_U196 );
nand NAND2_6232 ( R1207_U370 , R1207_U145 , R1207_U196 );
not NOT1_6233 ( R1207_U371 , R1207_U186 );
nand NAND2_6234 ( R1207_U372 , R1207_U244 , R1207_U174 );
not NOT1_6235 ( R1207_U373 , R1207_U108 );
nand NAND2_6236 ( R1207_U374 , R1207_U15 , R1207_U174 );
not NOT1_6237 ( R1207_U375 , R1207_U203 );
nand NAND2_6238 ( R1207_U376 , R1207_U18 , R1207_U174 );
not NOT1_6239 ( R1207_U377 , R1207_U202 );
nand NAND2_6240 ( R1207_U378 , R1207_U142 , R1207_U174 );
not NOT1_6241 ( R1207_U379 , R1207_U201 );
nand NAND2_6242 ( R1207_U380 , R1207_U131 , R1207_U57 );
not NOT1_6243 ( R1207_U381 , R1207_U178 );
nand NAND2_6244 ( R1207_U382 , R1207_U215 , R1207_U57 );
nand NAND2_6245 ( R1207_U383 , R1207_U140 , R1207_U382 );
nand NAND2_6246 ( R1207_U384 , R1207_U224 , R1207_U42 );
nand NAND2_6247 ( R1207_U385 , R1207_U288 , R1207_U197 );
not NOT1_6248 ( R1207_U386 , R1207_U196 );
nand NAND2_6249 ( R1207_U387 , R1207_U158 , R1207_U12 );
nand NAND2_6250 ( R1207_U388 , R1207_U159 , R1207_U457 );
nand NAND2_6251 ( R1207_U389 , U3484 , R1207_U54 );
nand NAND2_6252 ( R1207_U390 , U3080 , R1207_U53 );
nand NAND2_6253 ( R1207_U391 , R1207_U245 , R1207_U174 );
nand NAND2_6254 ( R1207_U392 , R1207_U243 , R1207_U173 );
nand NAND2_6255 ( R1207_U393 , U3482 , R1207_U35 );
nand NAND2_6256 ( R1207_U394 , U3081 , R1207_U40 );
nand NAND2_6257 ( R1207_U395 , U3482 , R1207_U35 );
nand NAND2_6258 ( R1207_U396 , U3081 , R1207_U40 );
nand NAND2_6259 ( R1207_U397 , R1207_U396 , R1207_U395 );
nand NAND2_6260 ( R1207_U398 , U3480 , R1207_U33 );
nand NAND2_6261 ( R1207_U399 , U3067 , R1207_U39 );
nand NAND2_6262 ( R1207_U400 , R1207_U250 , R1207_U55 );
nand NAND2_6263 ( R1207_U401 , R1207_U175 , R1207_U238 );
nand NAND2_6264 ( R1207_U402 , U3478 , R1207_U48 );
nand NAND2_6265 ( R1207_U403 , U3068 , R1207_U37 );
nand NAND2_6266 ( R1207_U404 , R1207_U403 , R1207_U402 );
nand NAND2_6267 ( R1207_U405 , U3476 , R1207_U49 );
nand NAND2_6268 ( R1207_U406 , U3064 , R1207_U36 );
nand NAND2_6269 ( R1207_U407 , R1207_U260 , R1207_U56 );
nand NAND2_6270 ( R1207_U408 , R1207_U176 , R1207_U252 );
nand NAND2_6271 ( R1207_U409 , U3474 , R1207_U50 );
nand NAND2_6272 ( R1207_U410 , U3057 , R1207_U38 );
nand NAND2_6273 ( R1207_U411 , R1207_U178 , R1207_U261 );
nand NAND2_6274 ( R1207_U412 , R1207_U381 , R1207_U177 );
nand NAND2_6275 ( R1207_U413 , U3472 , R1207_U43 );
nand NAND2_6276 ( R1207_U414 , U3061 , R1207_U47 );
nand NAND2_6277 ( R1207_U415 , U3472 , R1207_U43 );
nand NAND2_6278 ( R1207_U416 , U3061 , R1207_U47 );
nand NAND2_6279 ( R1207_U417 , R1207_U416 , R1207_U415 );
nand NAND2_6280 ( R1207_U418 , U3470 , R1207_U41 );
nand NAND2_6281 ( R1207_U419 , U3065 , R1207_U44 );
nand NAND2_6282 ( R1207_U420 , R1207_U263 , R1207_U57 );
nand NAND2_6283 ( R1207_U421 , R1207_U179 , R1207_U224 );
nand NAND2_6284 ( R1207_U422 , U4040 , R1207_U181 );
nand NAND2_6285 ( R1207_U423 , U3052 , R1207_U180 );
nand NAND2_6286 ( R1207_U424 , U4040 , R1207_U181 );
nand NAND2_6287 ( R1207_U425 , U3052 , R1207_U180 );
nand NAND2_6288 ( R1207_U426 , R1207_U425 , R1207_U424 );
nand NAND3_6289 ( R1207_U427 , U4029 , R1207_U23 , R1207_U102 );
nand NAND3_6290 ( R1207_U428 , R1207_U426 , R1207_U101 , U3051 );
nand NAND2_6291 ( R1207_U429 , U4029 , R1207_U102 );
nand NAND2_6292 ( R1207_U430 , U3051 , R1207_U101 );
not NOT1_6293 ( R1207_U431 , R1207_U152 );
nand NAND2_6294 ( R1207_U432 , R1207_U310 , R1207_U431 );
nand NAND2_6295 ( R1207_U433 , R1207_U152 , R1207_U183 );
nand NAND2_6296 ( R1207_U434 , U4030 , R1207_U100 );
nand NAND2_6297 ( R1207_U435 , U3050 , R1207_U59 );
nand NAND2_6298 ( R1207_U436 , R1207_U435 , R1207_U434 );
nand NAND2_6299 ( R1207_U437 , U4030 , R1207_U100 );
nand NAND2_6300 ( R1207_U438 , U3050 , R1207_U59 );
nand NAND3_6301 ( R1207_U439 , R1207_U438 , R1207_U437 , R1207_U99 );
nand NAND2_6302 ( R1207_U440 , R1207_U436 , R1207_U208 );
nand NAND2_6303 ( R1207_U441 , U4031 , R1207_U98 );
nand NAND2_6304 ( R1207_U442 , U3054 , R1207_U58 );
nand NAND2_6305 ( R1207_U443 , R1207_U186 , R1207_U314 );
nand NAND2_6306 ( R1207_U444 , R1207_U371 , R1207_U185 );
nand NAND2_6307 ( R1207_U445 , U4032 , R1207_U60 );
nand NAND2_6308 ( R1207_U446 , U3055 , R1207_U61 );
not NOT1_6309 ( R1207_U447 , R1207_U155 );
nand NAND2_6310 ( R1207_U448 , R1207_U368 , R1207_U447 );
nand NAND2_6311 ( R1207_U449 , R1207_U155 , R1207_U187 );
nand NAND2_6312 ( R1207_U450 , U4033 , R1207_U62 );
nand NAND2_6313 ( R1207_U451 , U3062 , R1207_U63 );
not NOT1_6314 ( R1207_U452 , R1207_U156 );
nand NAND2_6315 ( R1207_U453 , R1207_U366 , R1207_U452 );
nand NAND2_6316 ( R1207_U454 , R1207_U156 , R1207_U188 );
nand NAND2_6317 ( R1207_U455 , U4034 , R1207_U64 );
nand NAND2_6318 ( R1207_U456 , U3063 , R1207_U67 );
nand NAND2_6319 ( R1207_U457 , R1207_U456 , R1207_U455 );
nand NAND3_6320 ( R1207_U458 , R1207_U161 , R1207_U369 , R1207_U69 );
nand NAND2_6321 ( R1207_U459 , R1207_U22 , R1207_U219 );
nand NAND2_6322 ( R1207_U460 , U4035 , R1207_U65 );
nand NAND2_6323 ( R1207_U461 , U3058 , R1207_U68 );
nand NAND2_6324 ( R1207_U462 , R1207_U319 , R1207_U190 );
nand NAND2_6325 ( R1207_U463 , R1207_U316 , R1207_U189 );
nand NAND2_6326 ( R1207_U464 , U4036 , R1207_U66 );
nand NAND2_6327 ( R1207_U465 , U3072 , R1207_U70 );
nand NAND2_6328 ( R1207_U466 , R1207_U192 , R1207_U320 );
nand NAND2_6329 ( R1207_U467 , R1207_U364 , R1207_U191 );
nand NAND2_6330 ( R1207_U468 , U4037 , R1207_U71 );
nand NAND2_6331 ( R1207_U469 , U3073 , R1207_U73 );
not NOT1_6332 ( R1207_U470 , R1207_U162 );
nand NAND2_6333 ( R1207_U471 , R1207_U362 , R1207_U470 );
nand NAND2_6334 ( R1207_U472 , R1207_U162 , R1207_U193 );
nand NAND2_6335 ( R1207_U473 , U3468 , R1207_U46 );
nand NAND2_6336 ( R1207_U474 , U3075 , R1207_U194 );
not NOT1_6337 ( R1207_U475 , R1207_U163 );
nand NAND2_6338 ( R1207_U476 , R1207_U222 , R1207_U475 );
nand NAND2_6339 ( R1207_U477 , R1207_U163 , R1207_U195 );
nand NAND2_6340 ( R1207_U478 , U3504 , R1207_U72 );
nand NAND2_6341 ( R1207_U479 , U3078 , R1207_U75 );
not NOT1_6342 ( R1207_U480 , R1207_U164 );
nand NAND2_6343 ( R1207_U481 , R1207_U386 , R1207_U480 );
nand NAND2_6344 ( R1207_U482 , R1207_U164 , R1207_U196 );
nand NAND2_6345 ( R1207_U483 , U3502 , R1207_U76 );
nand NAND2_6346 ( R1207_U484 , U3079 , R1207_U97 );
not NOT1_6347 ( R1207_U485 , R1207_U165 );
nand NAND2_6348 ( R1207_U486 , R1207_U287 , R1207_U485 );
nand NAND2_6349 ( R1207_U487 , R1207_U165 , R1207_U197 );
nand NAND2_6350 ( R1207_U488 , U3500 , R1207_U77 );
nand NAND2_6351 ( R1207_U489 , U3066 , R1207_U78 );
not NOT1_6352 ( R1207_U490 , R1207_U166 );
nand NAND2_6353 ( R1207_U491 , R1207_U284 , R1207_U490 );
nand NAND2_6354 ( R1207_U492 , R1207_U166 , R1207_U198 );
nand NAND2_6355 ( R1207_U493 , U3498 , R1207_U92 );
nand NAND2_6356 ( R1207_U494 , U3070 , R1207_U79 );
nand NAND2_6357 ( R1207_U495 , R1207_U494 , R1207_U493 );
nand NAND2_6358 ( R1207_U496 , U3496 , R1207_U93 );
nand NAND2_6359 ( R1207_U497 , U3071 , R1207_U80 );
nand NAND2_6360 ( R1207_U498 , R1207_U330 , R1207_U107 );
nand NAND2_6361 ( R1207_U499 , R1207_U199 , R1207_U322 );
nand NAND2_6362 ( R1207_U500 , U3494 , R1207_U94 );
nand NAND2_6363 ( R1207_U501 , U3076 , R1207_U81 );
nand NAND2_6364 ( R1207_U502 , R1207_U201 , R1207_U331 );
nand NAND2_6365 ( R1207_U503 , R1207_U379 , R1207_U200 );
nand NAND2_6366 ( R1207_U504 , U3492 , R1207_U82 );
nand NAND2_6367 ( R1207_U505 , U3077 , R1207_U83 );
not NOT1_6368 ( R1207_U506 , R1207_U169 );
nand NAND2_6369 ( R1207_U507 , R1207_U377 , R1207_U506 );
nand NAND2_6370 ( R1207_U508 , R1207_U169 , R1207_U202 );
nand NAND2_6371 ( R1207_U509 , U3490 , R1207_U90 );
nand NAND2_6372 ( R1207_U510 , U3069 , R1207_U84 );
not NOT1_6373 ( R1207_U511 , R1207_U170 );
nand NAND2_6374 ( R1207_U512 , R1207_U375 , R1207_U511 );
nand NAND2_6375 ( R1207_U513 , R1207_U170 , R1207_U203 );
nand NAND2_6376 ( R1207_U514 , U3488 , R1207_U85 );
nand NAND2_6377 ( R1207_U515 , U3060 , R1207_U87 );
nand NAND2_6378 ( R1207_U516 , R1207_U515 , R1207_U514 );
nand NAND2_6379 ( R1207_U517 , U3486 , R1207_U86 );
nand NAND2_6380 ( R1207_U518 , U3059 , R1207_U88 );
nand NAND2_6381 ( R1207_U519 , R1207_U108 , R1207_U339 );
nand NAND2_6382 ( R1207_U520 , R1207_U204 , R1207_U373 );
and AND2_6383 ( R1165_U4 , R1165_U216 , R1165_U215 );
and AND2_6384 ( R1165_U5 , R1165_U226 , R1165_U225 );
and AND2_6385 ( R1165_U6 , R1165_U252 , R1165_U251 );
and AND2_6386 ( R1165_U7 , R1165_U268 , R1165_U267 );
and AND2_6387 ( R1165_U8 , R1165_U280 , R1165_U279 );
and AND2_6388 ( R1165_U9 , R1165_U298 , R1165_U297 );
and AND2_6389 ( R1165_U10 , R1165_U6 , R1165_U256 );
and AND2_6390 ( R1165_U11 , R1165_U5 , R1165_U223 );
and AND2_6391 ( R1165_U12 , R1165_U343 , R1165_U340 );
and AND2_6392 ( R1165_U13 , R1165_U334 , R1165_U331 );
and AND2_6393 ( R1165_U14 , R1165_U327 , R1165_U324 );
and AND2_6394 ( R1165_U15 , R1165_U318 , R1165_U315 );
and AND2_6395 ( R1165_U16 , R1165_U245 , R1165_U242 );
and AND2_6396 ( R1165_U17 , R1165_U238 , R1165_U235 );
not NOT1_6397 ( R1165_U18 , U3208 );
not NOT1_6398 ( R1165_U19 , U3170 );
not NOT1_6399 ( R1165_U20 , U3172 );
nand NAND2_6400 ( R1165_U21 , U3172 , R1165_U64 );
not NOT1_6401 ( R1165_U22 , U3171 );
not NOT1_6402 ( R1165_U23 , U3173 );
nand NAND2_6403 ( R1165_U24 , U3173 , R1165_U66 );
not NOT1_6404 ( R1165_U25 , U3174 );
not NOT1_6405 ( R1165_U26 , U3176 );
nand NAND2_6406 ( R1165_U27 , U3176 , R1165_U68 );
not NOT1_6407 ( R1165_U28 , U3175 );
not NOT1_6408 ( R1165_U29 , U3177 );
not NOT1_6409 ( R1165_U30 , U3178 );
nand NAND2_6410 ( R1165_U31 , U3178 , U3208 );
not NOT1_6411 ( R1165_U32 , U3169 );
nand NAND3_6412 ( R1165_U33 , R1165_U230 , R1165_U229 , R1165_U360 );
nand NAND2_6413 ( R1165_U34 , R1165_U364 , R1165_U24 );
nand NAND3_6414 ( R1165_U35 , R1165_U358 , R1165_U213 , R1165_U357 );
not NOT1_6415 ( R1165_U36 , U3162 );
nand NAND2_6416 ( R1165_U37 , U3162 , R1165_U72 );
not NOT1_6417 ( R1165_U38 , U3161 );
not NOT1_6418 ( R1165_U39 , U3166 );
not NOT1_6419 ( R1165_U40 , U3167 );
nand NAND2_6420 ( R1165_U41 , U3167 , R1165_U76 );
not NOT1_6421 ( R1165_U42 , U3165 );
not NOT1_6422 ( R1165_U43 , U3168 );
nand NAND2_6423 ( R1165_U44 , U3168 , R1165_U77 );
not NOT1_6424 ( R1165_U45 , U3164 );
not NOT1_6425 ( R1165_U46 , U3163 );
not NOT1_6426 ( R1165_U47 , U3160 );
not NOT1_6427 ( R1165_U48 , U3158 );
not NOT1_6428 ( R1165_U49 , U3159 );
nand NAND2_6429 ( R1165_U50 , U3159 , R1165_U81 );
not NOT1_6430 ( R1165_U51 , U3157 );
not NOT1_6431 ( R1165_U52 , U3156 );
not NOT1_6432 ( R1165_U53 , U3155 );
not NOT1_6433 ( R1165_U54 , U3153 );
not NOT1_6434 ( R1165_U55 , U3154 );
nand NAND2_6435 ( R1165_U56 , U3154 , R1165_U86 );
not NOT1_6436 ( R1165_U57 , U3152 );
not NOT1_6437 ( R1165_U58 , U3151 );
nand NAND2_6438 ( R1165_U59 , R1165_U50 , R1165_U320 );
nand NAND2_6439 ( R1165_U60 , R1165_U265 , R1165_U264 );
nand NAND2_6440 ( R1165_U61 , R1165_U41 , R1165_U336 );
nand NAND2_6441 ( R1165_U62 , R1165_U377 , R1165_U376 );
nand NAND2_6442 ( R1165_U63 , R1165_U400 , R1165_U399 );
nand NAND2_6443 ( R1165_U64 , R1165_U409 , R1165_U408 );
nand NAND2_6444 ( R1165_U65 , R1165_U406 , R1165_U405 );
nand NAND2_6445 ( R1165_U66 , R1165_U403 , R1165_U402 );
nand NAND2_6446 ( R1165_U67 , R1165_U385 , R1165_U384 );
nand NAND2_6447 ( R1165_U68 , R1165_U397 , R1165_U396 );
nand NAND2_6448 ( R1165_U69 , R1165_U394 , R1165_U393 );
nand NAND2_6449 ( R1165_U70 , R1165_U388 , R1165_U387 );
nand NAND2_6450 ( R1165_U71 , R1165_U391 , R1165_U390 );
nand NAND2_6451 ( R1165_U72 , R1165_U473 , R1165_U472 );
nand NAND2_6452 ( R1165_U73 , R1165_U470 , R1165_U469 );
nand NAND2_6453 ( R1165_U74 , R1165_U458 , R1165_U457 );
nand NAND2_6454 ( R1165_U75 , R1165_U455 , R1165_U454 );
nand NAND2_6455 ( R1165_U76 , R1165_U452 , R1165_U451 );
nand NAND2_6456 ( R1165_U77 , R1165_U461 , R1165_U460 );
nand NAND2_6457 ( R1165_U78 , R1165_U464 , R1165_U463 );
nand NAND2_6458 ( R1165_U79 , R1165_U467 , R1165_U466 );
nand NAND2_6459 ( R1165_U80 , R1165_U476 , R1165_U475 );
nand NAND2_6460 ( R1165_U81 , R1165_U485 , R1165_U484 );
nand NAND2_6461 ( R1165_U82 , R1165_U479 , R1165_U478 );
nand NAND2_6462 ( R1165_U83 , R1165_U482 , R1165_U481 );
nand NAND2_6463 ( R1165_U84 , R1165_U488 , R1165_U487 );
nand NAND2_6464 ( R1165_U85 , R1165_U491 , R1165_U490 );
nand NAND2_6465 ( R1165_U86 , R1165_U500 , R1165_U499 );
nand NAND2_6466 ( R1165_U87 , R1165_U494 , R1165_U493 );
nand NAND2_6467 ( R1165_U88 , R1165_U497 , R1165_U496 );
nand NAND2_6468 ( R1165_U89 , R1165_U449 , R1165_U448 );
nand NAND2_6469 ( R1165_U90 , R1165_U506 , R1165_U505 );
nand NAND2_6470 ( R1165_U91 , R1165_U613 , R1165_U612 );
nand NAND2_6471 ( R1165_U92 , R1165_U412 , R1165_U411 );
nand NAND2_6472 ( R1165_U93 , R1165_U419 , R1165_U418 );
nand NAND2_6473 ( R1165_U94 , R1165_U426 , R1165_U425 );
nand NAND2_6474 ( R1165_U95 , R1165_U433 , R1165_U432 );
nand NAND2_6475 ( R1165_U96 , R1165_U440 , R1165_U439 );
nand NAND2_6476 ( R1165_U97 , R1165_U447 , R1165_U446 );
nand NAND2_6477 ( R1165_U98 , R1165_U509 , R1165_U508 );
nand NAND2_6478 ( R1165_U99 , R1165_U516 , R1165_U515 );
nand NAND2_6479 ( R1165_U100 , R1165_U523 , R1165_U522 );
nand NAND2_6480 ( R1165_U101 , R1165_U528 , R1165_U527 );
nand NAND2_6481 ( R1165_U102 , R1165_U535 , R1165_U534 );
nand NAND2_6482 ( R1165_U103 , R1165_U542 , R1165_U541 );
nand NAND2_6483 ( R1165_U104 , R1165_U549 , R1165_U548 );
nand NAND2_6484 ( R1165_U105 , R1165_U556 , R1165_U555 );
nand NAND2_6485 ( R1165_U106 , R1165_U561 , R1165_U560 );
nand NAND2_6486 ( R1165_U107 , R1165_U568 , R1165_U567 );
nand NAND2_6487 ( R1165_U108 , R1165_U575 , R1165_U574 );
nand NAND2_6488 ( R1165_U109 , R1165_U582 , R1165_U581 );
nand NAND2_6489 ( R1165_U110 , R1165_U589 , R1165_U588 );
nand NAND2_6490 ( R1165_U111 , R1165_U596 , R1165_U595 );
nand NAND2_6491 ( R1165_U112 , R1165_U601 , R1165_U600 );
nand NAND2_6492 ( R1165_U113 , R1165_U608 , R1165_U607 );
and AND2_6493 ( R1165_U114 , R1165_U71 , R1165_U209 );
and AND2_6494 ( R1165_U115 , R1165_U219 , R1165_U218 );
and AND2_6495 ( R1165_U116 , R1165_U11 , R1165_U231 );
and AND2_6496 ( R1165_U117 , R1165_U362 , R1165_U232 );
and AND3_6497 ( R1165_U118 , R1165_U421 , R1165_U420 , R1165_U21 );
and AND2_6498 ( R1165_U119 , R1165_U237 , R1165_U5 );
and AND3_6499 ( R1165_U120 , R1165_U442 , R1165_U441 , R1165_U27 );
and AND2_6500 ( R1165_U121 , R1165_U244 , R1165_U4 );
and AND2_6501 ( R1165_U122 , R1165_U254 , R1165_U203 );
and AND2_6502 ( R1165_U123 , R1165_U249 , R1165_U10 );
and AND2_6503 ( R1165_U124 , R1165_U363 , R1165_U258 );
and AND2_6504 ( R1165_U125 , R1165_U272 , R1165_U271 );
and AND2_6505 ( R1165_U126 , R1165_U284 , R1165_U8 );
and AND2_6506 ( R1165_U127 , R1165_U282 , R1165_U204 );
and AND2_6507 ( R1165_U128 , R1165_U302 , R1165_U9 );
and AND2_6508 ( R1165_U129 , R1165_U300 , R1165_U205 );
and AND2_6509 ( R1165_U130 , R1165_U305 , R1165_U308 );
nand NAND2_6510 ( R1165_U131 , R1165_U503 , R1165_U502 );
and AND3_6511 ( R1165_U132 , R1165_U518 , R1165_U517 , R1165_U205 );
and AND2_6512 ( R1165_U133 , R1165_U56 , R1165_U205 );
and AND2_6513 ( R1165_U134 , R1165_U317 , R1165_U9 );
and AND3_6514 ( R1165_U135 , R1165_U544 , R1165_U543 , R1165_U204 );
and AND2_6515 ( R1165_U136 , R1165_U326 , R1165_U8 );
and AND3_6516 ( R1165_U137 , R1165_U570 , R1165_U569 , R1165_U37 );
and AND2_6517 ( R1165_U138 , R1165_U333 , R1165_U7 );
and AND3_6518 ( R1165_U139 , R1165_U591 , R1165_U590 , R1165_U203 );
and AND2_6519 ( R1165_U140 , R1165_U342 , R1165_U6 );
nand NAND2_6520 ( R1165_U141 , R1165_U610 , R1165_U609 );
not NOT1_6521 ( R1165_U142 , U3198 );
and AND2_6522 ( R1165_U143 , R1165_U380 , R1165_U379 );
not NOT1_6523 ( R1165_U144 , U3203 );
not NOT1_6524 ( R1165_U145 , U3206 );
not NOT1_6525 ( R1165_U146 , U3207 );
not NOT1_6526 ( R1165_U147 , U3204 );
not NOT1_6527 ( R1165_U148 , U3205 );
not NOT1_6528 ( R1165_U149 , U3199 );
not NOT1_6529 ( R1165_U150 , U3202 );
not NOT1_6530 ( R1165_U151 , U3200 );
not NOT1_6531 ( R1165_U152 , U3201 );
nand NAND2_6532 ( R1165_U153 , R1165_U117 , R1165_U368 );
and AND2_6533 ( R1165_U154 , R1165_U414 , R1165_U413 );
nand NAND2_6534 ( R1165_U155 , R1165_U361 , R1165_U366 );
and AND2_6535 ( R1165_U156 , R1165_U428 , R1165_U427 );
nand NAND2_6536 ( R1165_U157 , R1165_U370 , R1165_U354 );
and AND2_6537 ( R1165_U158 , R1165_U435 , R1165_U434 );
nand NAND2_6538 ( R1165_U159 , R1165_U115 , R1165_U220 );
not NOT1_6539 ( R1165_U160 , U3180 );
not NOT1_6540 ( R1165_U161 , U3196 );
not NOT1_6541 ( R1165_U162 , U3194 );
not NOT1_6542 ( R1165_U163 , U3195 );
not NOT1_6543 ( R1165_U164 , U3197 );
not NOT1_6544 ( R1165_U165 , U3193 );
not NOT1_6545 ( R1165_U166 , U3192 );
not NOT1_6546 ( R1165_U167 , U3190 );
not NOT1_6547 ( R1165_U168 , U3191 );
not NOT1_6548 ( R1165_U169 , U3189 );
not NOT1_6549 ( R1165_U170 , U3186 );
not NOT1_6550 ( R1165_U171 , U3187 );
not NOT1_6551 ( R1165_U172 , U3188 );
not NOT1_6552 ( R1165_U173 , U3185 );
not NOT1_6553 ( R1165_U174 , U3184 );
not NOT1_6554 ( R1165_U175 , U3181 );
not NOT1_6555 ( R1165_U176 , U3182 );
not NOT1_6556 ( R1165_U177 , U3183 );
not NOT1_6557 ( R1165_U178 , U3150 );
not NOT1_6558 ( R1165_U179 , U3179 );
and AND2_6559 ( R1165_U180 , R1165_U511 , R1165_U510 );
nand NAND2_6560 ( R1165_U181 , R1165_U305 , R1165_U304 );
nand NAND2_6561 ( R1165_U182 , R1165_U56 , R1165_U311 );
nand NAND2_6562 ( R1165_U183 , R1165_U295 , R1165_U294 );
and AND2_6563 ( R1165_U184 , R1165_U530 , R1165_U529 );
nand NAND2_6564 ( R1165_U185 , R1165_U291 , R1165_U290 );
and AND2_6565 ( R1165_U186 , R1165_U537 , R1165_U536 );
nand NAND2_6566 ( R1165_U187 , R1165_U287 , R1165_U286 );
and AND2_6567 ( R1165_U188 , R1165_U551 , R1165_U550 );
nand NAND2_6568 ( R1165_U189 , R1165_U31 , R1165_U210 );
nand NAND2_6569 ( R1165_U190 , R1165_U277 , R1165_U276 );
and AND2_6570 ( R1165_U191 , R1165_U563 , R1165_U562 );
nand NAND2_6571 ( R1165_U192 , R1165_U125 , R1165_U273 );
and AND2_6572 ( R1165_U193 , R1165_U577 , R1165_U576 );
nand NAND2_6573 ( R1165_U194 , R1165_U261 , R1165_U260 );
and AND2_6574 ( R1165_U195 , R1165_U584 , R1165_U583 );
nand NAND2_6575 ( R1165_U196 , R1165_U124 , R1165_U374 );
nand NAND2_6576 ( R1165_U197 , R1165_U372 , R1165_U44 );
and AND2_6577 ( R1165_U198 , R1165_U603 , R1165_U602 );
nand NAND3_6578 ( R1165_U199 , R1165_U247 , R1165_U201 , R1165_U355 );
nand NAND2_6579 ( R1165_U200 , R1165_U310 , R1165_U181 );
nand NAND2_6580 ( R1165_U201 , R1165_U62 , R1165_U153 );
not NOT1_6581 ( R1165_U202 , R1165_U27 );
nand NAND2_6582 ( R1165_U203 , U3166 , R1165_U74 );
nand NAND2_6583 ( R1165_U204 , U3158 , R1165_U83 );
nand NAND2_6584 ( R1165_U205 , U3153 , R1165_U88 );
not NOT1_6585 ( R1165_U206 , R1165_U41 );
not NOT1_6586 ( R1165_U207 , R1165_U50 );
not NOT1_6587 ( R1165_U208 , R1165_U56 );
or OR2_6588 ( R1165_U209 , U3208 , U3178 );
nand NAND2_6589 ( R1165_U210 , R1165_U71 , R1165_U209 );
not NOT1_6590 ( R1165_U211 , R1165_U31 );
not NOT1_6591 ( R1165_U212 , R1165_U189 );
nand NAND2_6592 ( R1165_U213 , U3177 , R1165_U70 );
not NOT1_6593 ( R1165_U214 , R1165_U35 );
nand NAND2_6594 ( R1165_U215 , R1165_U395 , R1165_U28 );
nand NAND2_6595 ( R1165_U216 , R1165_U398 , R1165_U26 );
nand NAND2_6596 ( R1165_U217 , R1165_U28 , R1165_U27 );
nand NAND2_6597 ( R1165_U218 , R1165_U69 , R1165_U217 );
nand NAND2_6598 ( R1165_U219 , U3175 , R1165_U202 );
nand NAND2_6599 ( R1165_U220 , R1165_U4 , R1165_U35 );
not NOT1_6600 ( R1165_U221 , R1165_U159 );
nand NAND2_6601 ( R1165_U222 , R1165_U386 , R1165_U25 );
nand NAND2_6602 ( R1165_U223 , R1165_U404 , R1165_U23 );
not NOT1_6603 ( R1165_U224 , R1165_U24 );
nand NAND2_6604 ( R1165_U225 , R1165_U407 , R1165_U22 );
nand NAND2_6605 ( R1165_U226 , R1165_U410 , R1165_U20 );
not NOT1_6606 ( R1165_U227 , R1165_U21 );
nand NAND2_6607 ( R1165_U228 , R1165_U22 , R1165_U21 );
nand NAND2_6608 ( R1165_U229 , R1165_U65 , R1165_U228 );
nand NAND2_6609 ( R1165_U230 , U3171 , R1165_U227 );
nand NAND2_6610 ( R1165_U231 , R1165_U401 , R1165_U19 );
nand NAND2_6611 ( R1165_U232 , U3170 , R1165_U63 );
nand NAND2_6612 ( R1165_U233 , R1165_U410 , R1165_U20 );
nand NAND2_6613 ( R1165_U234 , R1165_U233 , R1165_U34 );
nand NAND2_6614 ( R1165_U235 , R1165_U118 , R1165_U234 );
nand NAND2_6615 ( R1165_U236 , R1165_U365 , R1165_U21 );
nand NAND2_6616 ( R1165_U237 , U3171 , R1165_U65 );
nand NAND2_6617 ( R1165_U238 , R1165_U119 , R1165_U236 );
nand NAND2_6618 ( R1165_U239 , R1165_U410 , R1165_U20 );
nand NAND2_6619 ( R1165_U240 , R1165_U398 , R1165_U26 );
nand NAND2_6620 ( R1165_U241 , R1165_U240 , R1165_U35 );
nand NAND2_6621 ( R1165_U242 , R1165_U120 , R1165_U241 );
nand NAND2_6622 ( R1165_U243 , R1165_U214 , R1165_U27 );
nand NAND2_6623 ( R1165_U244 , U3175 , R1165_U69 );
nand NAND2_6624 ( R1165_U245 , R1165_U121 , R1165_U243 );
nand NAND2_6625 ( R1165_U246 , R1165_U398 , R1165_U26 );
nand NAND2_6626 ( R1165_U247 , U3169 , R1165_U153 );
not NOT1_6627 ( R1165_U248 , R1165_U199 );
nand NAND2_6628 ( R1165_U249 , R1165_U462 , R1165_U43 );
not NOT1_6629 ( R1165_U250 , R1165_U44 );
nand NAND2_6630 ( R1165_U251 , R1165_U456 , R1165_U42 );
nand NAND2_6631 ( R1165_U252 , R1165_U459 , R1165_U39 );
nand NAND2_6632 ( R1165_U253 , R1165_U206 , R1165_U6 );
nand NAND2_6633 ( R1165_U254 , U3165 , R1165_U75 );
nand NAND2_6634 ( R1165_U255 , R1165_U122 , R1165_U253 );
nand NAND2_6635 ( R1165_U256 , R1165_U453 , R1165_U40 );
nand NAND2_6636 ( R1165_U257 , R1165_U456 , R1165_U42 );
nand NAND2_6637 ( R1165_U258 , R1165_U257 , R1165_U255 );
nand NAND2_6638 ( R1165_U259 , R1165_U465 , R1165_U45 );
nand NAND2_6639 ( R1165_U260 , R1165_U259 , R1165_U196 );
nand NAND2_6640 ( R1165_U261 , U3164 , R1165_U78 );
not NOT1_6641 ( R1165_U262 , R1165_U194 );
nand NAND2_6642 ( R1165_U263 , R1165_U468 , R1165_U46 );
nand NAND2_6643 ( R1165_U264 , R1165_U263 , R1165_U194 );
nand NAND2_6644 ( R1165_U265 , U3163 , R1165_U79 );
not NOT1_6645 ( R1165_U266 , R1165_U60 );
nand NAND2_6646 ( R1165_U267 , R1165_U471 , R1165_U38 );
nand NAND2_6647 ( R1165_U268 , R1165_U474 , R1165_U36 );
not NOT1_6648 ( R1165_U269 , R1165_U37 );
nand NAND2_6649 ( R1165_U270 , R1165_U38 , R1165_U37 );
nand NAND2_6650 ( R1165_U271 , R1165_U73 , R1165_U270 );
nand NAND2_6651 ( R1165_U272 , U3161 , R1165_U269 );
nand NAND2_6652 ( R1165_U273 , R1165_U7 , R1165_U60 );
not NOT1_6653 ( R1165_U274 , R1165_U192 );
nand NAND2_6654 ( R1165_U275 , R1165_U477 , R1165_U47 );
nand NAND2_6655 ( R1165_U276 , R1165_U275 , R1165_U192 );
nand NAND2_6656 ( R1165_U277 , U3160 , R1165_U80 );
not NOT1_6657 ( R1165_U278 , R1165_U190 );
nand NAND2_6658 ( R1165_U279 , R1165_U480 , R1165_U51 );
nand NAND2_6659 ( R1165_U280 , R1165_U483 , R1165_U48 );
nand NAND2_6660 ( R1165_U281 , R1165_U207 , R1165_U8 );
nand NAND2_6661 ( R1165_U282 , U3157 , R1165_U82 );
nand NAND2_6662 ( R1165_U283 , R1165_U127 , R1165_U281 );
nand NAND2_6663 ( R1165_U284 , R1165_U486 , R1165_U49 );
nand NAND2_6664 ( R1165_U285 , R1165_U480 , R1165_U51 );
nand NAND2_6665 ( R1165_U286 , R1165_U126 , R1165_U190 );
nand NAND2_6666 ( R1165_U287 , R1165_U285 , R1165_U283 );
not NOT1_6667 ( R1165_U288 , R1165_U187 );
nand NAND2_6668 ( R1165_U289 , R1165_U489 , R1165_U52 );
nand NAND2_6669 ( R1165_U290 , R1165_U289 , R1165_U187 );
nand NAND2_6670 ( R1165_U291 , U3156 , R1165_U84 );
not NOT1_6671 ( R1165_U292 , R1165_U185 );
nand NAND2_6672 ( R1165_U293 , R1165_U492 , R1165_U53 );
nand NAND2_6673 ( R1165_U294 , R1165_U293 , R1165_U185 );
nand NAND2_6674 ( R1165_U295 , U3155 , R1165_U85 );
not NOT1_6675 ( R1165_U296 , R1165_U183 );
nand NAND2_6676 ( R1165_U297 , R1165_U495 , R1165_U57 );
nand NAND2_6677 ( R1165_U298 , R1165_U498 , R1165_U54 );
nand NAND2_6678 ( R1165_U299 , R1165_U208 , R1165_U9 );
nand NAND2_6679 ( R1165_U300 , U3152 , R1165_U87 );
nand NAND2_6680 ( R1165_U301 , R1165_U129 , R1165_U299 );
nand NAND2_6681 ( R1165_U302 , R1165_U501 , R1165_U55 );
nand NAND2_6682 ( R1165_U303 , R1165_U495 , R1165_U57 );
nand NAND2_6683 ( R1165_U304 , R1165_U128 , R1165_U183 );
nand NAND2_6684 ( R1165_U305 , R1165_U303 , R1165_U301 );
not NOT1_6685 ( R1165_U306 , R1165_U181 );
nand NAND2_6686 ( R1165_U307 , R1165_U450 , R1165_U58 );
nand NAND2_6687 ( R1165_U308 , U3151 , R1165_U89 );
nand NAND2_6688 ( R1165_U309 , U3151 , R1165_U89 );
nand NAND2_6689 ( R1165_U310 , R1165_U450 , R1165_U58 );
nand NAND2_6690 ( R1165_U311 , R1165_U302 , R1165_U183 );
not NOT1_6691 ( R1165_U312 , R1165_U182 );
nand NAND2_6692 ( R1165_U313 , R1165_U498 , R1165_U54 );
nand NAND2_6693 ( R1165_U314 , R1165_U313 , R1165_U182 );
nand NAND2_6694 ( R1165_U315 , R1165_U132 , R1165_U314 );
nand NAND2_6695 ( R1165_U316 , R1165_U133 , R1165_U311 );
nand NAND2_6696 ( R1165_U317 , U3152 , R1165_U87 );
nand NAND2_6697 ( R1165_U318 , R1165_U134 , R1165_U316 );
nand NAND2_6698 ( R1165_U319 , R1165_U498 , R1165_U54 );
nand NAND2_6699 ( R1165_U320 , R1165_U284 , R1165_U190 );
not NOT1_6700 ( R1165_U321 , R1165_U59 );
nand NAND2_6701 ( R1165_U322 , R1165_U483 , R1165_U48 );
nand NAND2_6702 ( R1165_U323 , R1165_U322 , R1165_U59 );
nand NAND2_6703 ( R1165_U324 , R1165_U135 , R1165_U323 );
nand NAND2_6704 ( R1165_U325 , R1165_U321 , R1165_U204 );
nand NAND2_6705 ( R1165_U326 , U3157 , R1165_U82 );
nand NAND2_6706 ( R1165_U327 , R1165_U136 , R1165_U325 );
nand NAND2_6707 ( R1165_U328 , R1165_U483 , R1165_U48 );
nand NAND2_6708 ( R1165_U329 , R1165_U474 , R1165_U36 );
nand NAND2_6709 ( R1165_U330 , R1165_U329 , R1165_U60 );
nand NAND2_6710 ( R1165_U331 , R1165_U137 , R1165_U330 );
nand NAND2_6711 ( R1165_U332 , R1165_U266 , R1165_U37 );
nand NAND2_6712 ( R1165_U333 , U3161 , R1165_U73 );
nand NAND2_6713 ( R1165_U334 , R1165_U138 , R1165_U332 );
nand NAND2_6714 ( R1165_U335 , R1165_U474 , R1165_U36 );
nand NAND2_6715 ( R1165_U336 , R1165_U256 , R1165_U197 );
not NOT1_6716 ( R1165_U337 , R1165_U61 );
nand NAND2_6717 ( R1165_U338 , R1165_U459 , R1165_U39 );
nand NAND2_6718 ( R1165_U339 , R1165_U338 , R1165_U61 );
nand NAND2_6719 ( R1165_U340 , R1165_U139 , R1165_U339 );
nand NAND2_6720 ( R1165_U341 , R1165_U337 , R1165_U203 );
nand NAND2_6721 ( R1165_U342 , U3165 , R1165_U75 );
nand NAND2_6722 ( R1165_U343 , R1165_U140 , R1165_U341 );
nand NAND2_6723 ( R1165_U344 , R1165_U459 , R1165_U39 );
nand NAND2_6724 ( R1165_U345 , R1165_U239 , R1165_U21 );
nand NAND2_6725 ( R1165_U346 , R1165_U246 , R1165_U27 );
nand NAND2_6726 ( R1165_U347 , R1165_U319 , R1165_U205 );
nand NAND2_6727 ( R1165_U348 , R1165_U302 , R1165_U56 );
nand NAND2_6728 ( R1165_U349 , R1165_U328 , R1165_U204 );
nand NAND2_6729 ( R1165_U350 , R1165_U284 , R1165_U50 );
nand NAND2_6730 ( R1165_U351 , R1165_U335 , R1165_U37 );
nand NAND2_6731 ( R1165_U352 , R1165_U344 , R1165_U203 );
nand NAND2_6732 ( R1165_U353 , R1165_U256 , R1165_U41 );
nand NAND2_6733 ( R1165_U354 , U3174 , R1165_U67 );
nand NAND2_6734 ( R1165_U355 , U3169 , R1165_U62 );
nand NAND2_6735 ( R1165_U356 , R1165_U130 , R1165_U304 );
nand NAND2_6736 ( R1165_U357 , R1165_U114 , R1165_U359 );
nand NAND2_6737 ( R1165_U358 , R1165_U211 , R1165_U359 );
nand NAND2_6738 ( R1165_U359 , R1165_U389 , R1165_U29 );
nand NAND2_6739 ( R1165_U360 , R1165_U224 , R1165_U5 );
not NOT1_6740 ( R1165_U361 , R1165_U33 );
nand NAND2_6741 ( R1165_U362 , R1165_U33 , R1165_U231 );
nand NAND2_6742 ( R1165_U363 , R1165_U250 , R1165_U10 );
nand NAND2_6743 ( R1165_U364 , R1165_U223 , R1165_U157 );
not NOT1_6744 ( R1165_U365 , R1165_U34 );
nand NAND2_6745 ( R1165_U366 , R1165_U11 , R1165_U157 );
not NOT1_6746 ( R1165_U367 , R1165_U155 );
nand NAND2_6747 ( R1165_U368 , R1165_U116 , R1165_U157 );
not NOT1_6748 ( R1165_U369 , R1165_U153 );
nand NAND2_6749 ( R1165_U370 , R1165_U222 , R1165_U159 );
not NOT1_6750 ( R1165_U371 , R1165_U157 );
nand NAND2_6751 ( R1165_U372 , R1165_U249 , R1165_U199 );
not NOT1_6752 ( R1165_U373 , R1165_U197 );
nand NAND2_6753 ( R1165_U374 , R1165_U123 , R1165_U199 );
not NOT1_6754 ( R1165_U375 , R1165_U196 );
nand NAND2_6755 ( R1165_U376 , U3208 , R1165_U142 );
nand NAND2_6756 ( R1165_U377 , U3198 , R1165_U18 );
not NOT1_6757 ( R1165_U378 , R1165_U62 );
nand NAND2_6758 ( R1165_U379 , R1165_U378 , U3169 );
nand NAND2_6759 ( R1165_U380 , R1165_U62 , R1165_U32 );
nand NAND2_6760 ( R1165_U381 , R1165_U378 , U3169 );
nand NAND2_6761 ( R1165_U382 , R1165_U62 , R1165_U32 );
nand NAND2_6762 ( R1165_U383 , R1165_U382 , R1165_U381 );
nand NAND2_6763 ( R1165_U384 , U3208 , R1165_U144 );
nand NAND2_6764 ( R1165_U385 , U3203 , R1165_U18 );
not NOT1_6765 ( R1165_U386 , R1165_U67 );
nand NAND2_6766 ( R1165_U387 , U3208 , R1165_U145 );
nand NAND2_6767 ( R1165_U388 , U3206 , R1165_U18 );
not NOT1_6768 ( R1165_U389 , R1165_U70 );
nand NAND2_6769 ( R1165_U390 , U3208 , R1165_U146 );
nand NAND2_6770 ( R1165_U391 , U3207 , R1165_U18 );
not NOT1_6771 ( R1165_U392 , R1165_U71 );
nand NAND2_6772 ( R1165_U393 , U3208 , R1165_U147 );
nand NAND2_6773 ( R1165_U394 , U3204 , R1165_U18 );
not NOT1_6774 ( R1165_U395 , R1165_U69 );
nand NAND2_6775 ( R1165_U396 , U3208 , R1165_U148 );
nand NAND2_6776 ( R1165_U397 , U3205 , R1165_U18 );
not NOT1_6777 ( R1165_U398 , R1165_U68 );
nand NAND2_6778 ( R1165_U399 , U3208 , R1165_U149 );
nand NAND2_6779 ( R1165_U400 , U3199 , R1165_U18 );
not NOT1_6780 ( R1165_U401 , R1165_U63 );
nand NAND2_6781 ( R1165_U402 , U3208 , R1165_U150 );
nand NAND2_6782 ( R1165_U403 , U3202 , R1165_U18 );
not NOT1_6783 ( R1165_U404 , R1165_U66 );
nand NAND2_6784 ( R1165_U405 , U3208 , R1165_U151 );
nand NAND2_6785 ( R1165_U406 , U3200 , R1165_U18 );
not NOT1_6786 ( R1165_U407 , R1165_U65 );
nand NAND2_6787 ( R1165_U408 , U3208 , R1165_U152 );
nand NAND2_6788 ( R1165_U409 , U3201 , R1165_U18 );
not NOT1_6789 ( R1165_U410 , R1165_U64 );
nand NAND2_6790 ( R1165_U411 , R1165_U143 , R1165_U153 );
nand NAND2_6791 ( R1165_U412 , R1165_U369 , R1165_U383 );
nand NAND2_6792 ( R1165_U413 , R1165_U401 , U3170 );
nand NAND2_6793 ( R1165_U414 , R1165_U63 , R1165_U19 );
nand NAND2_6794 ( R1165_U415 , R1165_U401 , U3170 );
nand NAND2_6795 ( R1165_U416 , R1165_U63 , R1165_U19 );
nand NAND2_6796 ( R1165_U417 , R1165_U416 , R1165_U415 );
nand NAND2_6797 ( R1165_U418 , R1165_U154 , R1165_U155 );
nand NAND2_6798 ( R1165_U419 , R1165_U367 , R1165_U417 );
nand NAND2_6799 ( R1165_U420 , R1165_U407 , U3171 );
nand NAND2_6800 ( R1165_U421 , R1165_U65 , R1165_U22 );
nand NAND2_6801 ( R1165_U422 , R1165_U410 , U3172 );
nand NAND2_6802 ( R1165_U423 , R1165_U64 , R1165_U20 );
nand NAND2_6803 ( R1165_U424 , R1165_U423 , R1165_U422 );
nand NAND2_6804 ( R1165_U425 , R1165_U34 , R1165_U345 );
nand NAND2_6805 ( R1165_U426 , R1165_U424 , R1165_U365 );
nand NAND2_6806 ( R1165_U427 , R1165_U404 , U3173 );
nand NAND2_6807 ( R1165_U428 , R1165_U66 , R1165_U23 );
nand NAND2_6808 ( R1165_U429 , R1165_U404 , U3173 );
nand NAND2_6809 ( R1165_U430 , R1165_U66 , R1165_U23 );
nand NAND2_6810 ( R1165_U431 , R1165_U430 , R1165_U429 );
nand NAND2_6811 ( R1165_U432 , R1165_U156 , R1165_U157 );
nand NAND2_6812 ( R1165_U433 , R1165_U371 , R1165_U431 );
nand NAND2_6813 ( R1165_U434 , R1165_U386 , U3174 );
nand NAND2_6814 ( R1165_U435 , R1165_U67 , R1165_U25 );
nand NAND2_6815 ( R1165_U436 , R1165_U386 , U3174 );
nand NAND2_6816 ( R1165_U437 , R1165_U67 , R1165_U25 );
nand NAND2_6817 ( R1165_U438 , R1165_U437 , R1165_U436 );
nand NAND2_6818 ( R1165_U439 , R1165_U158 , R1165_U159 );
nand NAND2_6819 ( R1165_U440 , R1165_U221 , R1165_U438 );
nand NAND2_6820 ( R1165_U441 , R1165_U395 , U3175 );
nand NAND2_6821 ( R1165_U442 , R1165_U69 , R1165_U28 );
nand NAND2_6822 ( R1165_U443 , R1165_U398 , U3176 );
nand NAND2_6823 ( R1165_U444 , R1165_U68 , R1165_U26 );
nand NAND2_6824 ( R1165_U445 , R1165_U444 , R1165_U443 );
nand NAND2_6825 ( R1165_U446 , R1165_U346 , R1165_U35 );
nand NAND2_6826 ( R1165_U447 , R1165_U445 , R1165_U214 );
nand NAND2_6827 ( R1165_U448 , U3208 , R1165_U160 );
nand NAND2_6828 ( R1165_U449 , U3180 , R1165_U18 );
not NOT1_6829 ( R1165_U450 , R1165_U89 );
nand NAND2_6830 ( R1165_U451 , U3208 , R1165_U161 );
nand NAND2_6831 ( R1165_U452 , U3196 , R1165_U18 );
not NOT1_6832 ( R1165_U453 , R1165_U76 );
nand NAND2_6833 ( R1165_U454 , U3208 , R1165_U162 );
nand NAND2_6834 ( R1165_U455 , U3194 , R1165_U18 );
not NOT1_6835 ( R1165_U456 , R1165_U75 );
nand NAND2_6836 ( R1165_U457 , U3208 , R1165_U163 );
nand NAND2_6837 ( R1165_U458 , U3195 , R1165_U18 );
not NOT1_6838 ( R1165_U459 , R1165_U74 );
nand NAND2_6839 ( R1165_U460 , U3208 , R1165_U164 );
nand NAND2_6840 ( R1165_U461 , U3197 , R1165_U18 );
not NOT1_6841 ( R1165_U462 , R1165_U77 );
nand NAND2_6842 ( R1165_U463 , U3208 , R1165_U165 );
nand NAND2_6843 ( R1165_U464 , U3193 , R1165_U18 );
not NOT1_6844 ( R1165_U465 , R1165_U78 );
nand NAND2_6845 ( R1165_U466 , U3208 , R1165_U166 );
nand NAND2_6846 ( R1165_U467 , U3192 , R1165_U18 );
not NOT1_6847 ( R1165_U468 , R1165_U79 );
nand NAND2_6848 ( R1165_U469 , U3208 , R1165_U167 );
nand NAND2_6849 ( R1165_U470 , U3190 , R1165_U18 );
not NOT1_6850 ( R1165_U471 , R1165_U73 );
nand NAND2_6851 ( R1165_U472 , U3208 , R1165_U168 );
nand NAND2_6852 ( R1165_U473 , U3191 , R1165_U18 );
not NOT1_6853 ( R1165_U474 , R1165_U72 );
nand NAND2_6854 ( R1165_U475 , U3208 , R1165_U169 );
nand NAND2_6855 ( R1165_U476 , U3189 , R1165_U18 );
not NOT1_6856 ( R1165_U477 , R1165_U80 );
nand NAND2_6857 ( R1165_U478 , U3208 , R1165_U170 );
nand NAND2_6858 ( R1165_U479 , U3186 , R1165_U18 );
not NOT1_6859 ( R1165_U480 , R1165_U82 );
nand NAND2_6860 ( R1165_U481 , U3208 , R1165_U171 );
nand NAND2_6861 ( R1165_U482 , U3187 , R1165_U18 );
not NOT1_6862 ( R1165_U483 , R1165_U83 );
nand NAND2_6863 ( R1165_U484 , U3208 , R1165_U172 );
nand NAND2_6864 ( R1165_U485 , U3188 , R1165_U18 );
not NOT1_6865 ( R1165_U486 , R1165_U81 );
nand NAND2_6866 ( R1165_U487 , U3208 , R1165_U173 );
nand NAND2_6867 ( R1165_U488 , U3185 , R1165_U18 );
not NOT1_6868 ( R1165_U489 , R1165_U84 );
nand NAND2_6869 ( R1165_U490 , U3208 , R1165_U174 );
nand NAND2_6870 ( R1165_U491 , U3184 , R1165_U18 );
not NOT1_6871 ( R1165_U492 , R1165_U85 );
nand NAND2_6872 ( R1165_U493 , U3208 , R1165_U175 );
nand NAND2_6873 ( R1165_U494 , U3181 , R1165_U18 );
not NOT1_6874 ( R1165_U495 , R1165_U87 );
nand NAND2_6875 ( R1165_U496 , U3208 , R1165_U176 );
nand NAND2_6876 ( R1165_U497 , U3182 , R1165_U18 );
not NOT1_6877 ( R1165_U498 , R1165_U88 );
nand NAND2_6878 ( R1165_U499 , U3208 , R1165_U177 );
nand NAND2_6879 ( R1165_U500 , U3183 , R1165_U18 );
not NOT1_6880 ( R1165_U501 , R1165_U86 );
nand NAND2_6881 ( R1165_U502 , U3208 , R1165_U178 );
nand NAND2_6882 ( R1165_U503 , U3150 , R1165_U18 );
not NOT1_6883 ( R1165_U504 , R1165_U131 );
nand NAND2_6884 ( R1165_U505 , U3179 , R1165_U504 );
nand NAND2_6885 ( R1165_U506 , R1165_U131 , R1165_U179 );
not NOT1_6886 ( R1165_U507 , R1165_U90 );
nand NAND3_6887 ( R1165_U508 , R1165_U356 , R1165_U307 , R1165_U507 );
nand NAND3_6888 ( R1165_U509 , R1165_U309 , R1165_U200 , R1165_U90 );
nand NAND2_6889 ( R1165_U510 , R1165_U450 , U3151 );
nand NAND2_6890 ( R1165_U511 , R1165_U89 , R1165_U58 );
nand NAND2_6891 ( R1165_U512 , R1165_U450 , U3151 );
nand NAND2_6892 ( R1165_U513 , R1165_U89 , R1165_U58 );
nand NAND2_6893 ( R1165_U514 , R1165_U513 , R1165_U512 );
nand NAND2_6894 ( R1165_U515 , R1165_U180 , R1165_U181 );
nand NAND2_6895 ( R1165_U516 , R1165_U306 , R1165_U514 );
nand NAND2_6896 ( R1165_U517 , R1165_U495 , U3152 );
nand NAND2_6897 ( R1165_U518 , R1165_U87 , R1165_U57 );
nand NAND2_6898 ( R1165_U519 , R1165_U498 , U3153 );
nand NAND2_6899 ( R1165_U520 , R1165_U88 , R1165_U54 );
nand NAND2_6900 ( R1165_U521 , R1165_U520 , R1165_U519 );
nand NAND2_6901 ( R1165_U522 , R1165_U347 , R1165_U182 );
nand NAND2_6902 ( R1165_U523 , R1165_U312 , R1165_U521 );
nand NAND2_6903 ( R1165_U524 , R1165_U501 , U3154 );
nand NAND2_6904 ( R1165_U525 , R1165_U86 , R1165_U55 );
nand NAND2_6905 ( R1165_U526 , R1165_U525 , R1165_U524 );
nand NAND2_6906 ( R1165_U527 , R1165_U348 , R1165_U183 );
nand NAND2_6907 ( R1165_U528 , R1165_U296 , R1165_U526 );
nand NAND2_6908 ( R1165_U529 , R1165_U492 , U3155 );
nand NAND2_6909 ( R1165_U530 , R1165_U85 , R1165_U53 );
nand NAND2_6910 ( R1165_U531 , R1165_U492 , U3155 );
nand NAND2_6911 ( R1165_U532 , R1165_U85 , R1165_U53 );
nand NAND2_6912 ( R1165_U533 , R1165_U532 , R1165_U531 );
nand NAND2_6913 ( R1165_U534 , R1165_U184 , R1165_U185 );
nand NAND2_6914 ( R1165_U535 , R1165_U292 , R1165_U533 );
nand NAND2_6915 ( R1165_U536 , R1165_U489 , U3156 );
nand NAND2_6916 ( R1165_U537 , R1165_U84 , R1165_U52 );
nand NAND2_6917 ( R1165_U538 , R1165_U489 , U3156 );
nand NAND2_6918 ( R1165_U539 , R1165_U84 , R1165_U52 );
nand NAND2_6919 ( R1165_U540 , R1165_U539 , R1165_U538 );
nand NAND2_6920 ( R1165_U541 , R1165_U186 , R1165_U187 );
nand NAND2_6921 ( R1165_U542 , R1165_U288 , R1165_U540 );
nand NAND2_6922 ( R1165_U543 , R1165_U480 , U3157 );
nand NAND2_6923 ( R1165_U544 , R1165_U82 , R1165_U51 );
nand NAND2_6924 ( R1165_U545 , R1165_U483 , U3158 );
nand NAND2_6925 ( R1165_U546 , R1165_U83 , R1165_U48 );
nand NAND2_6926 ( R1165_U547 , R1165_U546 , R1165_U545 );
nand NAND2_6927 ( R1165_U548 , R1165_U349 , R1165_U59 );
nand NAND2_6928 ( R1165_U549 , R1165_U547 , R1165_U321 );
nand NAND2_6929 ( R1165_U550 , R1165_U389 , U3177 );
nand NAND2_6930 ( R1165_U551 , R1165_U70 , R1165_U29 );
nand NAND2_6931 ( R1165_U552 , R1165_U389 , U3177 );
nand NAND2_6932 ( R1165_U553 , R1165_U70 , R1165_U29 );
nand NAND2_6933 ( R1165_U554 , R1165_U553 , R1165_U552 );
nand NAND2_6934 ( R1165_U555 , R1165_U188 , R1165_U189 );
nand NAND2_6935 ( R1165_U556 , R1165_U212 , R1165_U554 );
nand NAND2_6936 ( R1165_U557 , R1165_U486 , U3159 );
nand NAND2_6937 ( R1165_U558 , R1165_U81 , R1165_U49 );
nand NAND2_6938 ( R1165_U559 , R1165_U558 , R1165_U557 );
nand NAND2_6939 ( R1165_U560 , R1165_U350 , R1165_U190 );
nand NAND2_6940 ( R1165_U561 , R1165_U278 , R1165_U559 );
nand NAND2_6941 ( R1165_U562 , R1165_U477 , U3160 );
nand NAND2_6942 ( R1165_U563 , R1165_U80 , R1165_U47 );
nand NAND2_6943 ( R1165_U564 , R1165_U477 , U3160 );
nand NAND2_6944 ( R1165_U565 , R1165_U80 , R1165_U47 );
nand NAND2_6945 ( R1165_U566 , R1165_U565 , R1165_U564 );
nand NAND2_6946 ( R1165_U567 , R1165_U191 , R1165_U192 );
nand NAND2_6947 ( R1165_U568 , R1165_U274 , R1165_U566 );
nand NAND2_6948 ( R1165_U569 , R1165_U471 , U3161 );
nand NAND2_6949 ( R1165_U570 , R1165_U73 , R1165_U38 );
nand NAND2_6950 ( R1165_U571 , R1165_U474 , U3162 );
nand NAND2_6951 ( R1165_U572 , R1165_U72 , R1165_U36 );
nand NAND2_6952 ( R1165_U573 , R1165_U572 , R1165_U571 );
nand NAND2_6953 ( R1165_U574 , R1165_U351 , R1165_U60 );
nand NAND2_6954 ( R1165_U575 , R1165_U573 , R1165_U266 );
nand NAND2_6955 ( R1165_U576 , R1165_U468 , U3163 );
nand NAND2_6956 ( R1165_U577 , R1165_U79 , R1165_U46 );
nand NAND2_6957 ( R1165_U578 , R1165_U468 , U3163 );
nand NAND2_6958 ( R1165_U579 , R1165_U79 , R1165_U46 );
nand NAND2_6959 ( R1165_U580 , R1165_U579 , R1165_U578 );
nand NAND2_6960 ( R1165_U581 , R1165_U193 , R1165_U194 );
nand NAND2_6961 ( R1165_U582 , R1165_U262 , R1165_U580 );
nand NAND2_6962 ( R1165_U583 , R1165_U465 , U3164 );
nand NAND2_6963 ( R1165_U584 , R1165_U78 , R1165_U45 );
nand NAND2_6964 ( R1165_U585 , R1165_U465 , U3164 );
nand NAND2_6965 ( R1165_U586 , R1165_U78 , R1165_U45 );
nand NAND2_6966 ( R1165_U587 , R1165_U586 , R1165_U585 );
nand NAND2_6967 ( R1165_U588 , R1165_U195 , R1165_U196 );
nand NAND2_6968 ( R1165_U589 , R1165_U375 , R1165_U587 );
nand NAND2_6969 ( R1165_U590 , R1165_U456 , U3165 );
nand NAND2_6970 ( R1165_U591 , R1165_U75 , R1165_U42 );
nand NAND2_6971 ( R1165_U592 , R1165_U459 , U3166 );
nand NAND2_6972 ( R1165_U593 , R1165_U74 , R1165_U39 );
nand NAND2_6973 ( R1165_U594 , R1165_U593 , R1165_U592 );
nand NAND2_6974 ( R1165_U595 , R1165_U352 , R1165_U61 );
nand NAND2_6975 ( R1165_U596 , R1165_U594 , R1165_U337 );
nand NAND2_6976 ( R1165_U597 , R1165_U453 , U3167 );
nand NAND2_6977 ( R1165_U598 , R1165_U76 , R1165_U40 );
nand NAND2_6978 ( R1165_U599 , R1165_U598 , R1165_U597 );
nand NAND2_6979 ( R1165_U600 , R1165_U197 , R1165_U353 );
nand NAND2_6980 ( R1165_U601 , R1165_U373 , R1165_U599 );
nand NAND2_6981 ( R1165_U602 , R1165_U462 , U3168 );
nand NAND2_6982 ( R1165_U603 , R1165_U77 , R1165_U43 );
nand NAND2_6983 ( R1165_U604 , R1165_U462 , U3168 );
nand NAND2_6984 ( R1165_U605 , R1165_U77 , R1165_U43 );
nand NAND2_6985 ( R1165_U606 , R1165_U605 , R1165_U604 );
nand NAND2_6986 ( R1165_U607 , R1165_U198 , R1165_U199 );
nand NAND2_6987 ( R1165_U608 , R1165_U248 , R1165_U606 );
nand NAND2_6988 ( R1165_U609 , U3178 , R1165_U18 );
nand NAND2_6989 ( R1165_U610 , U3208 , R1165_U30 );
not NOT1_6990 ( R1165_U611 , R1165_U141 );
nand NAND2_6991 ( R1165_U612 , R1165_U71 , R1165_U611 );
nand NAND2_6992 ( R1165_U613 , R1165_U141 , R1165_U392 );
and AND2_6993 ( R1150_U6 , R1150_U224 , R1150_U223 );
and AND2_6994 ( R1150_U7 , R1150_U204 , R1150_U257 );
and AND2_6995 ( R1150_U8 , R1150_U259 , R1150_U258 );
and AND2_6996 ( R1150_U9 , R1150_U205 , R1150_U268 );
and AND2_6997 ( R1150_U10 , R1150_U270 , R1150_U269 );
and AND2_6998 ( R1150_U11 , R1150_U206 , R1150_U286 );
and AND2_6999 ( R1150_U12 , R1150_U288 , R1150_U287 );
and AND3_7000 ( R1150_U13 , R1150_U222 , R1150_U209 , R1150_U227 );
and AND2_7001 ( R1150_U14 , R1150_U232 , R1150_U210 );
and AND2_7002 ( R1150_U15 , R1150_U7 , R1150_U237 );
and AND2_7003 ( R1150_U16 , R1150_U9 , R1150_U273 );
and AND2_7004 ( R1150_U17 , R1150_U11 , R1150_U291 );
and AND2_7005 ( R1150_U18 , R1150_U15 , R1150_U264 );
and AND2_7006 ( R1150_U19 , R1150_U284 , R1150_U282 );
and AND2_7007 ( R1150_U20 , R1150_U19 , R1150_U17 );
and AND2_7008 ( R1150_U21 , R1150_U20 , R1150_U294 );
and AND2_7009 ( R1150_U22 , R1150_U418 , R1150_U417 );
nand NAND2_7010 ( R1150_U23 , R1150_U335 , R1150_U338 );
nand NAND2_7011 ( R1150_U24 , R1150_U326 , R1150_U329 );
nand NAND2_7012 ( R1150_U25 , R1150_U315 , R1150_U318 );
nand NAND2_7013 ( R1150_U26 , R1150_U307 , R1150_U309 );
nand NAND3_7014 ( R1150_U27 , R1150_U179 , R1150_U199 , R1150_U344 );
nand NAND2_7015 ( R1150_U28 , R1150_U255 , R1150_U380 );
nand NAND2_7016 ( R1150_U29 , R1150_U248 , R1150_U251 );
nand NAND2_7017 ( R1150_U30 , R1150_U240 , R1150_U242 );
nand NAND2_7018 ( R1150_U31 , R1150_U189 , R1150_U341 );
not NOT1_7019 ( R1150_U32 , U3067 );
nand NAND2_7020 ( R1150_U33 , U3067 , R1150_U38 );
not NOT1_7021 ( R1150_U34 , U3081 );
not NOT1_7022 ( R1150_U35 , U3476 );
not NOT1_7023 ( R1150_U36 , U3478 );
not NOT1_7024 ( R1150_U37 , U3474 );
not NOT1_7025 ( R1150_U38 , U3480 );
not NOT1_7026 ( R1150_U39 , U3482 );
not NOT1_7027 ( R1150_U40 , U3065 );
nand NAND2_7028 ( R1150_U41 , U3065 , R1150_U43 );
not NOT1_7029 ( R1150_U42 , U3061 );
not NOT1_7030 ( R1150_U43 , U3470 );
not NOT1_7031 ( R1150_U44 , U3464 );
not NOT1_7032 ( R1150_U45 , U3075 );
not NOT1_7033 ( R1150_U46 , U3472 );
not NOT1_7034 ( R1150_U47 , U3068 );
not NOT1_7035 ( R1150_U48 , U3064 );
not NOT1_7036 ( R1150_U49 , U3057 );
nand NAND2_7037 ( R1150_U50 , U3057 , R1150_U37 );
nand NAND2_7038 ( R1150_U51 , R1150_U228 , R1150_U226 );
not NOT1_7039 ( R1150_U52 , U3484 );
not NOT1_7040 ( R1150_U53 , U3080 );
nand NAND2_7041 ( R1150_U54 , R1150_U51 , R1150_U229 );
nand NAND2_7042 ( R1150_U55 , R1150_U50 , R1150_U244 );
nand NAND3_7043 ( R1150_U56 , R1150_U216 , R1150_U200 , R1150_U342 );
not NOT1_7044 ( R1150_U57 , U4031 );
not NOT1_7045 ( R1150_U58 , U4030 );
not NOT1_7046 ( R1150_U59 , U3055 );
not NOT1_7047 ( R1150_U60 , U4032 );
not NOT1_7048 ( R1150_U61 , U3062 );
not NOT1_7049 ( R1150_U62 , U4033 );
not NOT1_7050 ( R1150_U63 , U3063 );
not NOT1_7051 ( R1150_U64 , U3058 );
not NOT1_7052 ( R1150_U65 , U3072 );
not NOT1_7053 ( R1150_U66 , U4034 );
not NOT1_7054 ( R1150_U67 , U4035 );
nand NAND2_7055 ( R1150_U68 , U3072 , R1150_U69 );
not NOT1_7056 ( R1150_U69 , U4036 );
not NOT1_7057 ( R1150_U70 , U3073 );
not NOT1_7058 ( R1150_U71 , U3078 );
not NOT1_7059 ( R1150_U72 , U4037 );
nand NAND2_7060 ( R1150_U73 , U3078 , R1150_U74 );
not NOT1_7061 ( R1150_U74 , U3504 );
not NOT1_7062 ( R1150_U75 , U3079 );
not NOT1_7063 ( R1150_U76 , U3066 );
not NOT1_7064 ( R1150_U77 , U3500 );
not NOT1_7065 ( R1150_U78 , U3498 );
not NOT1_7066 ( R1150_U79 , U3496 );
not NOT1_7067 ( R1150_U80 , U3494 );
not NOT1_7068 ( R1150_U81 , U3077 );
not NOT1_7069 ( R1150_U82 , U3492 );
not NOT1_7070 ( R1150_U83 , U3490 );
not NOT1_7071 ( R1150_U84 , U3060 );
not NOT1_7072 ( R1150_U85 , U3059 );
not NOT1_7073 ( R1150_U86 , U3488 );
not NOT1_7074 ( R1150_U87 , U3486 );
nand NAND2_7075 ( R1150_U88 , U3080 , R1150_U52 );
not NOT1_7076 ( R1150_U89 , U3069 );
nand NAND2_7077 ( R1150_U90 , R1150_U347 , R1150_U264 );
not NOT1_7078 ( R1150_U91 , U3070 );
not NOT1_7079 ( R1150_U92 , U3071 );
not NOT1_7080 ( R1150_U93 , U3076 );
nand NAND2_7081 ( R1150_U94 , U3076 , R1150_U80 );
nand NAND2_7082 ( R1150_U95 , R1150_U274 , R1150_U272 );
not NOT1_7083 ( R1150_U96 , U3502 );
not NOT1_7084 ( R1150_U97 , U3054 );
nand NAND2_7085 ( R1150_U98 , U3054 , R1150_U57 );
not NOT1_7086 ( R1150_U99 , U3050 );
not NOT1_7087 ( R1150_U100 , U4029 );
not NOT1_7088 ( R1150_U101 , U3051 );
nand NAND2_7089 ( R1150_U102 , R1150_U146 , R1150_U367 );
nand NAND2_7090 ( R1150_U103 , R1150_U356 , R1150_U295 );
nand NAND2_7091 ( R1150_U104 , R1150_U354 , R1150_U293 );
nand NAND2_7092 ( R1150_U105 , R1150_U352 , R1150_U285 );
nand NAND2_7093 ( R1150_U106 , R1150_U68 , R1150_U311 );
nand NAND2_7094 ( R1150_U107 , R1150_U94 , R1150_U322 );
nand NAND2_7095 ( R1150_U108 , R1150_U369 , R1150_U88 );
not NOT1_7096 ( R1150_U109 , U3074 );
nand NAND2_7097 ( R1150_U110 , R1150_U428 , R1150_U427 );
nand NAND2_7098 ( R1150_U111 , R1150_U442 , R1150_U441 );
nand NAND2_7099 ( R1150_U112 , R1150_U447 , R1150_U446 );
nand NAND2_7100 ( R1150_U113 , R1150_U463 , R1150_U462 );
nand NAND2_7101 ( R1150_U114 , R1150_U468 , R1150_U467 );
nand NAND2_7102 ( R1150_U115 , R1150_U473 , R1150_U472 );
nand NAND2_7103 ( R1150_U116 , R1150_U478 , R1150_U477 );
nand NAND2_7104 ( R1150_U117 , R1150_U483 , R1150_U482 );
nand NAND2_7105 ( R1150_U118 , R1150_U499 , R1150_U498 );
nand NAND2_7106 ( R1150_U119 , R1150_U504 , R1150_U503 );
nand NAND2_7107 ( R1150_U120 , R1150_U387 , R1150_U386 );
nand NAND2_7108 ( R1150_U121 , R1150_U396 , R1150_U395 );
nand NAND2_7109 ( R1150_U122 , R1150_U403 , R1150_U402 );
nand NAND2_7110 ( R1150_U123 , R1150_U407 , R1150_U406 );
nand NAND2_7111 ( R1150_U124 , R1150_U416 , R1150_U415 );
nand NAND2_7112 ( R1150_U125 , R1150_U437 , R1150_U436 );
nand NAND2_7113 ( R1150_U126 , R1150_U454 , R1150_U453 );
nand NAND2_7114 ( R1150_U127 , R1150_U458 , R1150_U457 );
nand NAND2_7115 ( R1150_U128 , R1150_U490 , R1150_U489 );
nand NAND2_7116 ( R1150_U129 , R1150_U494 , R1150_U493 );
nand NAND2_7117 ( R1150_U130 , R1150_U511 , R1150_U510 );
and AND2_7118 ( R1150_U131 , R1150_U218 , R1150_U208 );
and AND2_7119 ( R1150_U132 , R1150_U221 , R1150_U220 );
and AND2_7120 ( R1150_U133 , R1150_U14 , R1150_U13 );
and AND2_7121 ( R1150_U134 , R1150_U235 , R1150_U234 );
and AND2_7122 ( R1150_U135 , R1150_U346 , R1150_U134 );
and AND3_7123 ( R1150_U136 , R1150_U389 , R1150_U388 , R1150_U33 );
and AND2_7124 ( R1150_U137 , R1150_U392 , R1150_U210 );
and AND2_7125 ( R1150_U138 , R1150_U250 , R1150_U6 );
and AND2_7126 ( R1150_U139 , R1150_U399 , R1150_U209 );
and AND3_7127 ( R1150_U140 , R1150_U409 , R1150_U408 , R1150_U41 );
and AND2_7128 ( R1150_U141 , R1150_U412 , R1150_U208 );
and AND2_7129 ( R1150_U142 , R1150_U266 , R1150_U18 );
and AND2_7130 ( R1150_U143 , R1150_U16 , R1150_U278 );
and AND2_7131 ( R1150_U144 , R1150_U351 , R1150_U279 );
and AND2_7132 ( R1150_U145 , R1150_U21 , R1150_U296 );
and AND2_7133 ( R1150_U146 , R1150_U358 , R1150_U297 );
and AND2_7134 ( R1150_U147 , R1150_U298 , R1150_U207 );
and AND2_7135 ( R1150_U148 , R1150_U301 , R1150_U302 );
and AND2_7136 ( R1150_U149 , R1150_U304 , R1150_U421 );
and AND2_7137 ( R1150_U150 , R1150_U301 , R1150_U302 );
and AND2_7138 ( R1150_U151 , R1150_U22 , R1150_U305 );
nand NAND2_7139 ( R1150_U152 , R1150_U425 , R1150_U424 );
and AND3_7140 ( R1150_U153 , R1150_U430 , R1150_U429 , R1150_U98 );
and AND2_7141 ( R1150_U154 , R1150_U433 , R1150_U207 );
nand NAND2_7142 ( R1150_U155 , R1150_U439 , R1150_U438 );
nand NAND2_7143 ( R1150_U156 , R1150_U444 , R1150_U443 );
and AND2_7144 ( R1150_U157 , R1150_U317 , R1150_U12 );
and AND2_7145 ( R1150_U158 , R1150_U450 , R1150_U206 );
nand NAND2_7146 ( R1150_U159 , R1150_U460 , R1150_U459 );
nand NAND2_7147 ( R1150_U160 , R1150_U465 , R1150_U464 );
nand NAND2_7148 ( R1150_U161 , R1150_U470 , R1150_U469 );
nand NAND2_7149 ( R1150_U162 , R1150_U475 , R1150_U474 );
nand NAND2_7150 ( R1150_U163 , R1150_U480 , R1150_U479 );
and AND2_7151 ( R1150_U164 , R1150_U328 , R1150_U10 );
and AND2_7152 ( R1150_U165 , R1150_U486 , R1150_U205 );
nand NAND2_7153 ( R1150_U166 , R1150_U496 , R1150_U495 );
nand NAND2_7154 ( R1150_U167 , R1150_U501 , R1150_U500 );
and AND2_7155 ( R1150_U168 , R1150_U337 , R1150_U8 );
and AND2_7156 ( R1150_U169 , R1150_U507 , R1150_U204 );
and AND2_7157 ( R1150_U170 , R1150_U385 , R1150_U384 );
nand NAND2_7158 ( R1150_U171 , R1150_U135 , R1150_U345 );
and AND2_7159 ( R1150_U172 , R1150_U394 , R1150_U393 );
and AND2_7160 ( R1150_U173 , R1150_U401 , R1150_U400 );
and AND2_7161 ( R1150_U174 , R1150_U405 , R1150_U404 );
nand NAND2_7162 ( R1150_U175 , R1150_U132 , R1150_U377 );
and AND2_7163 ( R1150_U176 , R1150_U414 , R1150_U413 );
not NOT1_7164 ( R1150_U177 , U4040 );
not NOT1_7165 ( R1150_U178 , U3052 );
and AND2_7166 ( R1150_U179 , R1150_U423 , R1150_U422 );
nand NAND2_7167 ( R1150_U180 , R1150_U148 , R1150_U299 );
and AND2_7168 ( R1150_U181 , R1150_U435 , R1150_U434 );
nand NAND2_7169 ( R1150_U182 , R1150_U357 , R1150_U365 );
nand NAND2_7170 ( R1150_U183 , R1150_U355 , R1150_U363 );
and AND2_7171 ( R1150_U184 , R1150_U452 , R1150_U451 );
and AND2_7172 ( R1150_U185 , R1150_U456 , R1150_U455 );
nand NAND2_7173 ( R1150_U186 , R1150_U353 , R1150_U361 );
nand NAND2_7174 ( R1150_U187 , R1150_U359 , R1150_U73 );
not NOT1_7175 ( R1150_U188 , U3468 );
nand NAND2_7176 ( R1150_U189 , U3464 , R1150_U109 );
nand NAND2_7177 ( R1150_U190 , R1150_U382 , R1150_U343 );
nand NAND2_7178 ( R1150_U191 , R1150_U144 , R1150_U350 );
nand NAND2_7179 ( R1150_U192 , R1150_U95 , R1150_U275 );
and AND2_7180 ( R1150_U193 , R1150_U488 , R1150_U487 );
and AND2_7181 ( R1150_U194 , R1150_U492 , R1150_U491 );
nand NAND3_7182 ( R1150_U195 , R1150_U349 , R1150_U267 , R1150_U375 );
nand NAND2_7183 ( R1150_U196 , R1150_U373 , R1150_U90 );
nand NAND2_7184 ( R1150_U197 , R1150_U371 , R1150_U263 );
and AND2_7185 ( R1150_U198 , R1150_U509 , R1150_U508 );
nand NAND2_7186 ( R1150_U199 , R1150_U149 , R1150_U180 );
nand NAND2_7187 ( R1150_U200 , R1150_U189 , R1150_U188 );
not NOT1_7188 ( R1150_U201 , R1150_U98 );
not NOT1_7189 ( R1150_U202 , R1150_U41 );
not NOT1_7190 ( R1150_U203 , R1150_U33 );
nand NAND2_7191 ( R1150_U204 , U3486 , R1150_U85 );
nand NAND2_7192 ( R1150_U205 , U3496 , R1150_U92 );
nand NAND2_7193 ( R1150_U206 , U4035 , R1150_U64 );
nand NAND2_7194 ( R1150_U207 , U4031 , R1150_U97 );
nand NAND2_7195 ( R1150_U208 , U3470 , R1150_U40 );
nand NAND2_7196 ( R1150_U209 , U3476 , R1150_U48 );
nand NAND2_7197 ( R1150_U210 , U3480 , R1150_U32 );
not NOT1_7198 ( R1150_U211 , R1150_U94 );
not NOT1_7199 ( R1150_U212 , R1150_U68 );
not NOT1_7200 ( R1150_U213 , R1150_U50 );
not NOT1_7201 ( R1150_U214 , R1150_U88 );
not NOT1_7202 ( R1150_U215 , R1150_U189 );
nand NAND2_7203 ( R1150_U216 , U3075 , R1150_U189 );
not NOT1_7204 ( R1150_U217 , R1150_U56 );
nand NAND2_7205 ( R1150_U218 , U3472 , R1150_U42 );
nand NAND2_7206 ( R1150_U219 , R1150_U42 , R1150_U41 );
nand NAND2_7207 ( R1150_U220 , R1150_U219 , R1150_U46 );
nand NAND2_7208 ( R1150_U221 , U3061 , R1150_U202 );
nand NAND2_7209 ( R1150_U222 , U3478 , R1150_U47 );
nand NAND2_7210 ( R1150_U223 , U3068 , R1150_U36 );
nand NAND2_7211 ( R1150_U224 , U3064 , R1150_U35 );
nand NAND2_7212 ( R1150_U225 , R1150_U213 , R1150_U209 );
nand NAND2_7213 ( R1150_U226 , R1150_U6 , R1150_U225 );
nand NAND2_7214 ( R1150_U227 , U3474 , R1150_U49 );
nand NAND2_7215 ( R1150_U228 , U3478 , R1150_U47 );
nand NAND2_7216 ( R1150_U229 , R1150_U13 , R1150_U175 );
not NOT1_7217 ( R1150_U230 , R1150_U51 );
not NOT1_7218 ( R1150_U231 , R1150_U54 );
nand NAND2_7219 ( R1150_U232 , U3482 , R1150_U34 );
nand NAND2_7220 ( R1150_U233 , R1150_U34 , R1150_U33 );
nand NAND2_7221 ( R1150_U234 , R1150_U233 , R1150_U39 );
nand NAND2_7222 ( R1150_U235 , U3081 , R1150_U203 );
not NOT1_7223 ( R1150_U236 , R1150_U171 );
nand NAND2_7224 ( R1150_U237 , U3484 , R1150_U53 );
nand NAND2_7225 ( R1150_U238 , R1150_U237 , R1150_U88 );
nand NAND2_7226 ( R1150_U239 , R1150_U231 , R1150_U33 );
nand NAND2_7227 ( R1150_U240 , R1150_U137 , R1150_U239 );
nand NAND2_7228 ( R1150_U241 , R1150_U54 , R1150_U210 );
nand NAND2_7229 ( R1150_U242 , R1150_U136 , R1150_U241 );
nand NAND2_7230 ( R1150_U243 , R1150_U33 , R1150_U210 );
nand NAND2_7231 ( R1150_U244 , R1150_U227 , R1150_U175 );
not NOT1_7232 ( R1150_U245 , R1150_U55 );
nand NAND2_7233 ( R1150_U246 , U3064 , R1150_U35 );
nand NAND2_7234 ( R1150_U247 , R1150_U245 , R1150_U246 );
nand NAND2_7235 ( R1150_U248 , R1150_U139 , R1150_U247 );
nand NAND2_7236 ( R1150_U249 , R1150_U55 , R1150_U209 );
nand NAND2_7237 ( R1150_U250 , U3478 , R1150_U47 );
nand NAND2_7238 ( R1150_U251 , R1150_U138 , R1150_U249 );
nand NAND2_7239 ( R1150_U252 , U3064 , R1150_U35 );
nand NAND2_7240 ( R1150_U253 , R1150_U209 , R1150_U252 );
nand NAND2_7241 ( R1150_U254 , R1150_U227 , R1150_U50 );
nand NAND2_7242 ( R1150_U255 , R1150_U141 , R1150_U381 );
nand NAND2_7243 ( R1150_U256 , R1150_U41 , R1150_U208 );
nand NAND2_7244 ( R1150_U257 , U3488 , R1150_U84 );
nand NAND2_7245 ( R1150_U258 , U3060 , R1150_U86 );
nand NAND2_7246 ( R1150_U259 , U3059 , R1150_U87 );
nand NAND2_7247 ( R1150_U260 , R1150_U214 , R1150_U7 );
nand NAND2_7248 ( R1150_U261 , R1150_U8 , R1150_U260 );
nand NAND2_7249 ( R1150_U262 , U3488 , R1150_U84 );
nand NAND2_7250 ( R1150_U263 , R1150_U262 , R1150_U261 );
nand NAND2_7251 ( R1150_U264 , U3490 , R1150_U89 );
nand NAND2_7252 ( R1150_U265 , U3069 , R1150_U83 );
nand NAND2_7253 ( R1150_U266 , U3492 , R1150_U81 );
nand NAND2_7254 ( R1150_U267 , U3077 , R1150_U82 );
nand NAND2_7255 ( R1150_U268 , U3498 , R1150_U91 );
nand NAND2_7256 ( R1150_U269 , U3070 , R1150_U78 );
nand NAND2_7257 ( R1150_U270 , U3071 , R1150_U79 );
nand NAND2_7258 ( R1150_U271 , R1150_U211 , R1150_U9 );
nand NAND2_7259 ( R1150_U272 , R1150_U10 , R1150_U271 );
nand NAND2_7260 ( R1150_U273 , U3494 , R1150_U93 );
nand NAND2_7261 ( R1150_U274 , U3498 , R1150_U91 );
nand NAND2_7262 ( R1150_U275 , R1150_U16 , R1150_U195 );
not NOT1_7263 ( R1150_U276 , R1150_U95 );
not NOT1_7264 ( R1150_U277 , R1150_U192 );
nand NAND2_7265 ( R1150_U278 , U3500 , R1150_U76 );
nand NAND2_7266 ( R1150_U279 , U3066 , R1150_U77 );
not NOT1_7267 ( R1150_U280 , R1150_U191 );
nand NAND2_7268 ( R1150_U281 , U3502 , R1150_U75 );
nand NAND2_7269 ( R1150_U282 , U3504 , R1150_U71 );
not NOT1_7270 ( R1150_U283 , R1150_U73 );
nand NAND2_7271 ( R1150_U284 , U4037 , R1150_U70 );
nand NAND2_7272 ( R1150_U285 , U3073 , R1150_U72 );
nand NAND2_7273 ( R1150_U286 , U4034 , R1150_U63 );
nand NAND2_7274 ( R1150_U287 , U3063 , R1150_U66 );
nand NAND2_7275 ( R1150_U288 , U3058 , R1150_U67 );
nand NAND2_7276 ( R1150_U289 , R1150_U212 , R1150_U11 );
nand NAND2_7277 ( R1150_U290 , R1150_U12 , R1150_U289 );
nand NAND2_7278 ( R1150_U291 , U4036 , R1150_U65 );
nand NAND2_7279 ( R1150_U292 , U4034 , R1150_U63 );
nand NAND2_7280 ( R1150_U293 , R1150_U292 , R1150_U290 );
nand NAND2_7281 ( R1150_U294 , U4033 , R1150_U61 );
nand NAND2_7282 ( R1150_U295 , U3062 , R1150_U62 );
nand NAND2_7283 ( R1150_U296 , U4032 , R1150_U59 );
nand NAND2_7284 ( R1150_U297 , U3055 , R1150_U60 );
nand NAND2_7285 ( R1150_U298 , U4030 , R1150_U99 );
nand NAND2_7286 ( R1150_U299 , R1150_U147 , R1150_U102 );
nand NAND2_7287 ( R1150_U300 , R1150_U99 , R1150_U98 );
nand NAND2_7288 ( R1150_U301 , R1150_U300 , R1150_U58 );
nand NAND2_7289 ( R1150_U302 , U3050 , R1150_U201 );
not NOT1_7290 ( R1150_U303 , R1150_U180 );
nand NAND2_7291 ( R1150_U304 , U4029 , R1150_U101 );
nand NAND2_7292 ( R1150_U305 , U3051 , R1150_U100 );
nand NAND2_7293 ( R1150_U306 , R1150_U368 , R1150_U98 );
nand NAND2_7294 ( R1150_U307 , R1150_U154 , R1150_U306 );
nand NAND2_7295 ( R1150_U308 , R1150_U102 , R1150_U207 );
nand NAND2_7296 ( R1150_U309 , R1150_U153 , R1150_U308 );
nand NAND2_7297 ( R1150_U310 , R1150_U98 , R1150_U207 );
nand NAND2_7298 ( R1150_U311 , R1150_U291 , R1150_U186 );
not NOT1_7299 ( R1150_U312 , R1150_U106 );
nand NAND2_7300 ( R1150_U313 , U3058 , R1150_U67 );
nand NAND2_7301 ( R1150_U314 , R1150_U312 , R1150_U313 );
nand NAND2_7302 ( R1150_U315 , R1150_U158 , R1150_U314 );
nand NAND2_7303 ( R1150_U316 , R1150_U106 , R1150_U206 );
nand NAND2_7304 ( R1150_U317 , U4034 , R1150_U63 );
nand NAND2_7305 ( R1150_U318 , R1150_U157 , R1150_U316 );
nand NAND2_7306 ( R1150_U319 , U3058 , R1150_U67 );
nand NAND2_7307 ( R1150_U320 , R1150_U206 , R1150_U319 );
nand NAND2_7308 ( R1150_U321 , R1150_U291 , R1150_U68 );
nand NAND2_7309 ( R1150_U322 , R1150_U273 , R1150_U195 );
not NOT1_7310 ( R1150_U323 , R1150_U107 );
nand NAND2_7311 ( R1150_U324 , U3071 , R1150_U79 );
nand NAND2_7312 ( R1150_U325 , R1150_U323 , R1150_U324 );
nand NAND2_7313 ( R1150_U326 , R1150_U165 , R1150_U325 );
nand NAND2_7314 ( R1150_U327 , R1150_U107 , R1150_U205 );
nand NAND2_7315 ( R1150_U328 , U3498 , R1150_U91 );
nand NAND2_7316 ( R1150_U329 , R1150_U164 , R1150_U327 );
nand NAND2_7317 ( R1150_U330 , U3071 , R1150_U79 );
nand NAND2_7318 ( R1150_U331 , R1150_U205 , R1150_U330 );
nand NAND2_7319 ( R1150_U332 , R1150_U273 , R1150_U94 );
nand NAND2_7320 ( R1150_U333 , U3059 , R1150_U87 );
nand NAND2_7321 ( R1150_U334 , R1150_U370 , R1150_U333 );
nand NAND2_7322 ( R1150_U335 , R1150_U169 , R1150_U334 );
nand NAND2_7323 ( R1150_U336 , R1150_U108 , R1150_U204 );
nand NAND2_7324 ( R1150_U337 , U3488 , R1150_U84 );
nand NAND2_7325 ( R1150_U338 , R1150_U168 , R1150_U336 );
nand NAND2_7326 ( R1150_U339 , U3059 , R1150_U87 );
nand NAND2_7327 ( R1150_U340 , R1150_U204 , R1150_U339 );
nand NAND2_7328 ( R1150_U341 , U3074 , R1150_U44 );
nand NAND2_7329 ( R1150_U342 , U3075 , R1150_U188 );
nand NAND2_7330 ( R1150_U343 , U3079 , R1150_U96 );
nand NAND3_7331 ( R1150_U344 , R1150_U150 , R1150_U299 , R1150_U151 );
nand NAND2_7332 ( R1150_U345 , R1150_U133 , R1150_U175 );
nand NAND2_7333 ( R1150_U346 , R1150_U230 , R1150_U14 );
nand NAND2_7334 ( R1150_U347 , R1150_U265 , R1150_U263 );
not NOT1_7335 ( R1150_U348 , R1150_U90 );
nand NAND2_7336 ( R1150_U349 , R1150_U348 , R1150_U266 );
nand NAND2_7337 ( R1150_U350 , R1150_U143 , R1150_U195 );
nand NAND2_7338 ( R1150_U351 , R1150_U276 , R1150_U278 );
nand NAND2_7339 ( R1150_U352 , R1150_U283 , R1150_U284 );
not NOT1_7340 ( R1150_U353 , R1150_U105 );
nand NAND2_7341 ( R1150_U354 , R1150_U17 , R1150_U105 );
not NOT1_7342 ( R1150_U355 , R1150_U104 );
nand NAND2_7343 ( R1150_U356 , R1150_U104 , R1150_U294 );
not NOT1_7344 ( R1150_U357 , R1150_U103 );
nand NAND2_7345 ( R1150_U358 , R1150_U103 , R1150_U296 );
nand NAND2_7346 ( R1150_U359 , R1150_U282 , R1150_U190 );
not NOT1_7347 ( R1150_U360 , R1150_U187 );
nand NAND2_7348 ( R1150_U361 , R1150_U19 , R1150_U190 );
not NOT1_7349 ( R1150_U362 , R1150_U186 );
nand NAND2_7350 ( R1150_U363 , R1150_U20 , R1150_U190 );
not NOT1_7351 ( R1150_U364 , R1150_U183 );
nand NAND2_7352 ( R1150_U365 , R1150_U21 , R1150_U190 );
not NOT1_7353 ( R1150_U366 , R1150_U182 );
nand NAND2_7354 ( R1150_U367 , R1150_U145 , R1150_U190 );
not NOT1_7355 ( R1150_U368 , R1150_U102 );
nand NAND2_7356 ( R1150_U369 , R1150_U237 , R1150_U171 );
not NOT1_7357 ( R1150_U370 , R1150_U108 );
nand NAND2_7358 ( R1150_U371 , R1150_U15 , R1150_U171 );
not NOT1_7359 ( R1150_U372 , R1150_U197 );
nand NAND2_7360 ( R1150_U373 , R1150_U18 , R1150_U171 );
not NOT1_7361 ( R1150_U374 , R1150_U196 );
nand NAND2_7362 ( R1150_U375 , R1150_U142 , R1150_U171 );
not NOT1_7363 ( R1150_U376 , R1150_U195 );
nand NAND2_7364 ( R1150_U377 , R1150_U131 , R1150_U56 );
not NOT1_7365 ( R1150_U378 , R1150_U175 );
nand NAND2_7366 ( R1150_U379 , R1150_U208 , R1150_U56 );
nand NAND2_7367 ( R1150_U380 , R1150_U140 , R1150_U379 );
nand NAND2_7368 ( R1150_U381 , R1150_U217 , R1150_U41 );
nand NAND2_7369 ( R1150_U382 , R1150_U281 , R1150_U191 );
not NOT1_7370 ( R1150_U383 , R1150_U190 );
nand NAND2_7371 ( R1150_U384 , U3484 , R1150_U53 );
nand NAND2_7372 ( R1150_U385 , U3080 , R1150_U52 );
nand NAND2_7373 ( R1150_U386 , R1150_U238 , R1150_U171 );
nand NAND2_7374 ( R1150_U387 , R1150_U236 , R1150_U170 );
nand NAND2_7375 ( R1150_U388 , U3482 , R1150_U34 );
nand NAND2_7376 ( R1150_U389 , U3081 , R1150_U39 );
nand NAND2_7377 ( R1150_U390 , U3482 , R1150_U34 );
nand NAND2_7378 ( R1150_U391 , U3081 , R1150_U39 );
nand NAND2_7379 ( R1150_U392 , R1150_U391 , R1150_U390 );
nand NAND2_7380 ( R1150_U393 , U3480 , R1150_U32 );
nand NAND2_7381 ( R1150_U394 , U3067 , R1150_U38 );
nand NAND2_7382 ( R1150_U395 , R1150_U243 , R1150_U54 );
nand NAND2_7383 ( R1150_U396 , R1150_U172 , R1150_U231 );
nand NAND2_7384 ( R1150_U397 , U3478 , R1150_U47 );
nand NAND2_7385 ( R1150_U398 , U3068 , R1150_U36 );
nand NAND2_7386 ( R1150_U399 , R1150_U398 , R1150_U397 );
nand NAND2_7387 ( R1150_U400 , U3476 , R1150_U48 );
nand NAND2_7388 ( R1150_U401 , U3064 , R1150_U35 );
nand NAND2_7389 ( R1150_U402 , R1150_U253 , R1150_U55 );
nand NAND2_7390 ( R1150_U403 , R1150_U173 , R1150_U245 );
nand NAND2_7391 ( R1150_U404 , U3474 , R1150_U49 );
nand NAND2_7392 ( R1150_U405 , U3057 , R1150_U37 );
nand NAND2_7393 ( R1150_U406 , R1150_U175 , R1150_U254 );
nand NAND2_7394 ( R1150_U407 , R1150_U378 , R1150_U174 );
nand NAND2_7395 ( R1150_U408 , U3472 , R1150_U42 );
nand NAND2_7396 ( R1150_U409 , U3061 , R1150_U46 );
nand NAND2_7397 ( R1150_U410 , U3472 , R1150_U42 );
nand NAND2_7398 ( R1150_U411 , U3061 , R1150_U46 );
nand NAND2_7399 ( R1150_U412 , R1150_U411 , R1150_U410 );
nand NAND2_7400 ( R1150_U413 , U3470 , R1150_U40 );
nand NAND2_7401 ( R1150_U414 , U3065 , R1150_U43 );
nand NAND2_7402 ( R1150_U415 , R1150_U256 , R1150_U56 );
nand NAND2_7403 ( R1150_U416 , R1150_U176 , R1150_U217 );
nand NAND2_7404 ( R1150_U417 , U4040 , R1150_U178 );
nand NAND2_7405 ( R1150_U418 , U3052 , R1150_U177 );
nand NAND2_7406 ( R1150_U419 , U4040 , R1150_U178 );
nand NAND2_7407 ( R1150_U420 , U3052 , R1150_U177 );
nand NAND2_7408 ( R1150_U421 , R1150_U420 , R1150_U419 );
nand NAND3_7409 ( R1150_U422 , U3051 , R1150_U421 , R1150_U100 );
nand NAND3_7410 ( R1150_U423 , R1150_U22 , R1150_U101 , U4029 );
nand NAND2_7411 ( R1150_U424 , U4029 , R1150_U101 );
nand NAND2_7412 ( R1150_U425 , U3051 , R1150_U100 );
not NOT1_7413 ( R1150_U426 , R1150_U152 );
nand NAND2_7414 ( R1150_U427 , R1150_U303 , R1150_U426 );
nand NAND2_7415 ( R1150_U428 , R1150_U152 , R1150_U180 );
nand NAND2_7416 ( R1150_U429 , U4030 , R1150_U99 );
nand NAND2_7417 ( R1150_U430 , U3050 , R1150_U58 );
nand NAND2_7418 ( R1150_U431 , U4030 , R1150_U99 );
nand NAND2_7419 ( R1150_U432 , U3050 , R1150_U58 );
nand NAND2_7420 ( R1150_U433 , R1150_U432 , R1150_U431 );
nand NAND2_7421 ( R1150_U434 , U4031 , R1150_U97 );
nand NAND2_7422 ( R1150_U435 , U3054 , R1150_U57 );
nand NAND2_7423 ( R1150_U436 , R1150_U102 , R1150_U310 );
nand NAND2_7424 ( R1150_U437 , R1150_U181 , R1150_U368 );
nand NAND2_7425 ( R1150_U438 , U4032 , R1150_U59 );
nand NAND2_7426 ( R1150_U439 , U3055 , R1150_U60 );
not NOT1_7427 ( R1150_U440 , R1150_U155 );
nand NAND2_7428 ( R1150_U441 , R1150_U366 , R1150_U440 );
nand NAND2_7429 ( R1150_U442 , R1150_U155 , R1150_U182 );
nand NAND2_7430 ( R1150_U443 , U4033 , R1150_U61 );
nand NAND2_7431 ( R1150_U444 , U3062 , R1150_U62 );
not NOT1_7432 ( R1150_U445 , R1150_U156 );
nand NAND2_7433 ( R1150_U446 , R1150_U364 , R1150_U445 );
nand NAND2_7434 ( R1150_U447 , R1150_U156 , R1150_U183 );
nand NAND2_7435 ( R1150_U448 , U4034 , R1150_U63 );
nand NAND2_7436 ( R1150_U449 , U3063 , R1150_U66 );
nand NAND2_7437 ( R1150_U450 , R1150_U449 , R1150_U448 );
nand NAND2_7438 ( R1150_U451 , U4035 , R1150_U64 );
nand NAND2_7439 ( R1150_U452 , U3058 , R1150_U67 );
nand NAND2_7440 ( R1150_U453 , R1150_U320 , R1150_U106 );
nand NAND2_7441 ( R1150_U454 , R1150_U184 , R1150_U312 );
nand NAND2_7442 ( R1150_U455 , U4036 , R1150_U65 );
nand NAND2_7443 ( R1150_U456 , U3072 , R1150_U69 );
nand NAND2_7444 ( R1150_U457 , R1150_U186 , R1150_U321 );
nand NAND2_7445 ( R1150_U458 , R1150_U362 , R1150_U185 );
nand NAND2_7446 ( R1150_U459 , U4037 , R1150_U70 );
nand NAND2_7447 ( R1150_U460 , U3073 , R1150_U72 );
not NOT1_7448 ( R1150_U461 , R1150_U159 );
nand NAND2_7449 ( R1150_U462 , R1150_U360 , R1150_U461 );
nand NAND2_7450 ( R1150_U463 , R1150_U159 , R1150_U187 );
nand NAND2_7451 ( R1150_U464 , U3468 , R1150_U45 );
nand NAND2_7452 ( R1150_U465 , U3075 , R1150_U188 );
not NOT1_7453 ( R1150_U466 , R1150_U160 );
nand NAND2_7454 ( R1150_U467 , R1150_U215 , R1150_U466 );
nand NAND2_7455 ( R1150_U468 , R1150_U160 , R1150_U189 );
nand NAND2_7456 ( R1150_U469 , U3504 , R1150_U71 );
nand NAND2_7457 ( R1150_U470 , U3078 , R1150_U74 );
not NOT1_7458 ( R1150_U471 , R1150_U161 );
nand NAND2_7459 ( R1150_U472 , R1150_U383 , R1150_U471 );
nand NAND2_7460 ( R1150_U473 , R1150_U161 , R1150_U190 );
nand NAND2_7461 ( R1150_U474 , U3502 , R1150_U75 );
nand NAND2_7462 ( R1150_U475 , U3079 , R1150_U96 );
not NOT1_7463 ( R1150_U476 , R1150_U162 );
nand NAND2_7464 ( R1150_U477 , R1150_U280 , R1150_U476 );
nand NAND2_7465 ( R1150_U478 , R1150_U162 , R1150_U191 );
nand NAND2_7466 ( R1150_U479 , U3500 , R1150_U76 );
nand NAND2_7467 ( R1150_U480 , U3066 , R1150_U77 );
not NOT1_7468 ( R1150_U481 , R1150_U163 );
nand NAND2_7469 ( R1150_U482 , R1150_U277 , R1150_U481 );
nand NAND2_7470 ( R1150_U483 , R1150_U163 , R1150_U192 );
nand NAND2_7471 ( R1150_U484 , U3498 , R1150_U91 );
nand NAND2_7472 ( R1150_U485 , U3070 , R1150_U78 );
nand NAND2_7473 ( R1150_U486 , R1150_U485 , R1150_U484 );
nand NAND2_7474 ( R1150_U487 , U3496 , R1150_U92 );
nand NAND2_7475 ( R1150_U488 , U3071 , R1150_U79 );
nand NAND2_7476 ( R1150_U489 , R1150_U331 , R1150_U107 );
nand NAND2_7477 ( R1150_U490 , R1150_U193 , R1150_U323 );
nand NAND2_7478 ( R1150_U491 , U3494 , R1150_U93 );
nand NAND2_7479 ( R1150_U492 , U3076 , R1150_U80 );
nand NAND2_7480 ( R1150_U493 , R1150_U195 , R1150_U332 );
nand NAND2_7481 ( R1150_U494 , R1150_U376 , R1150_U194 );
nand NAND2_7482 ( R1150_U495 , U3492 , R1150_U81 );
nand NAND2_7483 ( R1150_U496 , U3077 , R1150_U82 );
not NOT1_7484 ( R1150_U497 , R1150_U166 );
nand NAND2_7485 ( R1150_U498 , R1150_U374 , R1150_U497 );
nand NAND2_7486 ( R1150_U499 , R1150_U166 , R1150_U196 );
nand NAND2_7487 ( R1150_U500 , U3490 , R1150_U89 );
nand NAND2_7488 ( R1150_U501 , U3069 , R1150_U83 );
not NOT1_7489 ( R1150_U502 , R1150_U167 );
nand NAND2_7490 ( R1150_U503 , R1150_U372 , R1150_U502 );
nand NAND2_7491 ( R1150_U504 , R1150_U167 , R1150_U197 );
nand NAND2_7492 ( R1150_U505 , U3488 , R1150_U84 );
nand NAND2_7493 ( R1150_U506 , U3060 , R1150_U86 );
nand NAND2_7494 ( R1150_U507 , R1150_U506 , R1150_U505 );
nand NAND2_7495 ( R1150_U508 , U3486 , R1150_U85 );
nand NAND2_7496 ( R1150_U509 , U3059 , R1150_U87 );
nand NAND2_7497 ( R1150_U510 , R1150_U108 , R1150_U340 );
nand NAND2_7498 ( R1150_U511 , R1150_U198 , R1150_U370 );
and AND2_7499 ( R1192_U6 , R1192_U231 , R1192_U230 );
and AND2_7500 ( R1192_U7 , R1192_U211 , R1192_U264 );
and AND2_7501 ( R1192_U8 , R1192_U266 , R1192_U265 );
and AND2_7502 ( R1192_U9 , R1192_U212 , R1192_U275 );
and AND2_7503 ( R1192_U10 , R1192_U277 , R1192_U276 );
and AND2_7504 ( R1192_U11 , R1192_U106 , R1192_U293 );
and AND2_7505 ( R1192_U12 , R1192_U295 , R1192_U294 );
and AND3_7506 ( R1192_U13 , R1192_U229 , R1192_U216 , R1192_U234 );
and AND2_7507 ( R1192_U14 , R1192_U239 , R1192_U217 );
and AND2_7508 ( R1192_U15 , R1192_U7 , R1192_U244 );
and AND2_7509 ( R1192_U16 , R1192_U9 , R1192_U280 );
and AND2_7510 ( R1192_U17 , R1192_U11 , R1192_U298 );
and AND2_7511 ( R1192_U18 , R1192_U15 , R1192_U271 );
and AND2_7512 ( R1192_U19 , R1192_U291 , R1192_U289 );
and AND2_7513 ( R1192_U20 , R1192_U19 , R1192_U17 );
and AND2_7514 ( R1192_U21 , R1192_U20 , R1192_U301 );
and AND2_7515 ( R1192_U22 , R1192_U457 , R1192_U106 );
and AND2_7516 ( R1192_U23 , R1192_U423 , R1192_U422 );
nand NAND2_7517 ( R1192_U24 , R1192_U334 , R1192_U337 );
nand NAND2_7518 ( R1192_U25 , R1192_U325 , R1192_U328 );
nand NAND5_7519 ( R1192_U26 , R1192_U459 , R1192_U458 , R1192_U388 , R1192_U387 , R1192_U359 );
and AND2_7520 ( R1192_U27 , R1192_U344 , R1192_U313 );
nand NAND3_7521 ( R1192_U28 , R1192_U182 , R1192_U206 , R1192_U343 );
nand NAND2_7522 ( R1192_U29 , R1192_U262 , R1192_U383 );
nand NAND2_7523 ( R1192_U30 , R1192_U255 , R1192_U258 );
nand NAND2_7524 ( R1192_U31 , R1192_U247 , R1192_U249 );
nand NAND2_7525 ( R1192_U32 , R1192_U195 , R1192_U340 );
not NOT1_7526 ( R1192_U33 , U3067 );
nand NAND2_7527 ( R1192_U34 , U3067 , R1192_U39 );
not NOT1_7528 ( R1192_U35 , U3081 );
not NOT1_7529 ( R1192_U36 , U3476 );
not NOT1_7530 ( R1192_U37 , U3478 );
not NOT1_7531 ( R1192_U38 , U3474 );
not NOT1_7532 ( R1192_U39 , U3480 );
not NOT1_7533 ( R1192_U40 , U3482 );
not NOT1_7534 ( R1192_U41 , U3065 );
nand NAND2_7535 ( R1192_U42 , U3065 , R1192_U44 );
not NOT1_7536 ( R1192_U43 , U3061 );
not NOT1_7537 ( R1192_U44 , U3470 );
not NOT1_7538 ( R1192_U45 , U3464 );
not NOT1_7539 ( R1192_U46 , U3075 );
not NOT1_7540 ( R1192_U47 , U3472 );
not NOT1_7541 ( R1192_U48 , U3068 );
not NOT1_7542 ( R1192_U49 , U3064 );
not NOT1_7543 ( R1192_U50 , U3057 );
nand NAND2_7544 ( R1192_U51 , U3057 , R1192_U38 );
nand NAND2_7545 ( R1192_U52 , R1192_U235 , R1192_U233 );
not NOT1_7546 ( R1192_U53 , U3484 );
not NOT1_7547 ( R1192_U54 , U3080 );
nand NAND2_7548 ( R1192_U55 , R1192_U52 , R1192_U236 );
nand NAND2_7549 ( R1192_U56 , R1192_U51 , R1192_U251 );
nand NAND3_7550 ( R1192_U57 , R1192_U223 , R1192_U207 , R1192_U341 );
not NOT1_7551 ( R1192_U58 , U4031 );
not NOT1_7552 ( R1192_U59 , U4030 );
not NOT1_7553 ( R1192_U60 , U3055 );
not NOT1_7554 ( R1192_U61 , U4032 );
not NOT1_7555 ( R1192_U62 , U3062 );
not NOT1_7556 ( R1192_U63 , U4033 );
not NOT1_7557 ( R1192_U64 , U3063 );
not NOT1_7558 ( R1192_U65 , U3058 );
not NOT1_7559 ( R1192_U66 , U3072 );
not NOT1_7560 ( R1192_U67 , U4034 );
not NOT1_7561 ( R1192_U68 , U4035 );
nand NAND2_7562 ( R1192_U69 , U3072 , R1192_U70 );
not NOT1_7563 ( R1192_U70 , U4036 );
not NOT1_7564 ( R1192_U71 , U3073 );
not NOT1_7565 ( R1192_U72 , U3078 );
not NOT1_7566 ( R1192_U73 , U4037 );
nand NAND2_7567 ( R1192_U74 , U3078 , R1192_U75 );
not NOT1_7568 ( R1192_U75 , U3504 );
not NOT1_7569 ( R1192_U76 , U3079 );
not NOT1_7570 ( R1192_U77 , U3066 );
not NOT1_7571 ( R1192_U78 , U3500 );
not NOT1_7572 ( R1192_U79 , U3498 );
not NOT1_7573 ( R1192_U80 , U3496 );
not NOT1_7574 ( R1192_U81 , U3494 );
not NOT1_7575 ( R1192_U82 , U3077 );
not NOT1_7576 ( R1192_U83 , U3492 );
not NOT1_7577 ( R1192_U84 , U3490 );
not NOT1_7578 ( R1192_U85 , U3060 );
not NOT1_7579 ( R1192_U86 , U3059 );
not NOT1_7580 ( R1192_U87 , U3488 );
not NOT1_7581 ( R1192_U88 , U3486 );
nand NAND2_7582 ( R1192_U89 , U3080 , R1192_U53 );
not NOT1_7583 ( R1192_U90 , U3069 );
nand NAND2_7584 ( R1192_U91 , R1192_U347 , R1192_U271 );
not NOT1_7585 ( R1192_U92 , U3070 );
not NOT1_7586 ( R1192_U93 , U3071 );
not NOT1_7587 ( R1192_U94 , U3076 );
nand NAND2_7588 ( R1192_U95 , U3076 , R1192_U81 );
nand NAND2_7589 ( R1192_U96 , R1192_U281 , R1192_U279 );
not NOT1_7590 ( R1192_U97 , U3502 );
not NOT1_7591 ( R1192_U98 , U3054 );
nand NAND2_7592 ( R1192_U99 , U3054 , R1192_U58 );
not NOT1_7593 ( R1192_U100 , U3050 );
not NOT1_7594 ( R1192_U101 , U4029 );
not NOT1_7595 ( R1192_U102 , U3051 );
nand NAND2_7596 ( R1192_U103 , R1192_U356 , R1192_U302 );
nand NAND2_7597 ( R1192_U104 , R1192_U354 , R1192_U300 );
nand NAND2_7598 ( R1192_U105 , R1192_U352 , R1192_U292 );
nand NAND2_7599 ( R1192_U106 , U4035 , R1192_U65 );
nand NAND2_7600 ( R1192_U107 , R1192_U95 , R1192_U321 );
nand NAND2_7601 ( R1192_U108 , R1192_U372 , R1192_U89 );
not NOT1_7602 ( R1192_U109 , U3074 );
nand NAND2_7603 ( R1192_U110 , R1192_U433 , R1192_U432 );
nand NAND2_7604 ( R1192_U111 , R1192_U449 , R1192_U448 );
nand NAND2_7605 ( R1192_U112 , R1192_U454 , R1192_U453 );
nand NAND2_7606 ( R1192_U113 , R1192_U472 , R1192_U471 );
nand NAND2_7607 ( R1192_U114 , R1192_U477 , R1192_U476 );
nand NAND2_7608 ( R1192_U115 , R1192_U482 , R1192_U481 );
nand NAND2_7609 ( R1192_U116 , R1192_U487 , R1192_U486 );
nand NAND2_7610 ( R1192_U117 , R1192_U492 , R1192_U491 );
nand NAND2_7611 ( R1192_U118 , R1192_U508 , R1192_U507 );
nand NAND2_7612 ( R1192_U119 , R1192_U513 , R1192_U512 );
nand NAND2_7613 ( R1192_U120 , R1192_U392 , R1192_U391 );
nand NAND2_7614 ( R1192_U121 , R1192_U401 , R1192_U400 );
nand NAND2_7615 ( R1192_U122 , R1192_U408 , R1192_U407 );
nand NAND2_7616 ( R1192_U123 , R1192_U412 , R1192_U411 );
nand NAND2_7617 ( R1192_U124 , R1192_U421 , R1192_U420 );
nand NAND2_7618 ( R1192_U125 , R1192_U444 , R1192_U443 );
nand NAND2_7619 ( R1192_U126 , R1192_U463 , R1192_U462 );
nand NAND2_7620 ( R1192_U127 , R1192_U467 , R1192_U466 );
nand NAND2_7621 ( R1192_U128 , R1192_U499 , R1192_U498 );
nand NAND2_7622 ( R1192_U129 , R1192_U503 , R1192_U502 );
nand NAND2_7623 ( R1192_U130 , R1192_U520 , R1192_U519 );
and AND2_7624 ( R1192_U131 , R1192_U225 , R1192_U215 );
and AND2_7625 ( R1192_U132 , R1192_U228 , R1192_U227 );
and AND2_7626 ( R1192_U133 , R1192_U14 , R1192_U13 );
and AND2_7627 ( R1192_U134 , R1192_U242 , R1192_U241 );
and AND2_7628 ( R1192_U135 , R1192_U346 , R1192_U134 );
and AND3_7629 ( R1192_U136 , R1192_U394 , R1192_U393 , R1192_U34 );
and AND2_7630 ( R1192_U137 , R1192_U397 , R1192_U217 );
and AND2_7631 ( R1192_U138 , R1192_U257 , R1192_U6 );
and AND2_7632 ( R1192_U139 , R1192_U404 , R1192_U216 );
and AND3_7633 ( R1192_U140 , R1192_U414 , R1192_U413 , R1192_U42 );
and AND2_7634 ( R1192_U141 , R1192_U417 , R1192_U215 );
and AND2_7635 ( R1192_U142 , R1192_U273 , R1192_U18 );
and AND2_7636 ( R1192_U143 , R1192_U16 , R1192_U285 );
and AND2_7637 ( R1192_U144 , R1192_U351 , R1192_U286 );
and AND2_7638 ( R1192_U145 , R1192_U21 , R1192_U303 );
and AND2_7639 ( R1192_U146 , R1192_U358 , R1192_U304 );
and AND2_7640 ( R1192_U147 , R1192_U305 , R1192_U214 );
and AND2_7641 ( R1192_U148 , R1192_U308 , R1192_U309 );
and AND2_7642 ( R1192_U149 , R1192_U311 , R1192_U426 );
and AND2_7643 ( R1192_U150 , R1192_U308 , R1192_U309 );
and AND2_7644 ( R1192_U151 , R1192_U23 , R1192_U312 );
nand NAND2_7645 ( R1192_U152 , R1192_U430 , R1192_U429 );
and AND2_7646 ( R1192_U153 , R1192_U436 , R1192_U214 );
and AND2_7647 ( R1192_U154 , R1192_U214 , R1192_U186 );
nand NAND2_7648 ( R1192_U155 , R1192_U446 , R1192_U445 );
nand NAND2_7649 ( R1192_U156 , R1192_U451 , R1192_U450 );
and AND2_7650 ( R1192_U157 , R1192_U22 , R1192_U298 );
and AND2_7651 ( R1192_U158 , R1192_U213 , R1192_U317 );
and AND2_7652 ( R1192_U159 , U3058 , R1192_U68 );
and AND2_7653 ( R1192_U160 , R1192_U19 , R1192_U298 );
and AND3_7654 ( R1192_U161 , R1192_U360 , R1192_U317 , R1192_U12 );
nand NAND2_7655 ( R1192_U162 , R1192_U469 , R1192_U468 );
nand NAND2_7656 ( R1192_U163 , R1192_U474 , R1192_U473 );
nand NAND2_7657 ( R1192_U164 , R1192_U479 , R1192_U478 );
nand NAND2_7658 ( R1192_U165 , R1192_U484 , R1192_U483 );
nand NAND2_7659 ( R1192_U166 , R1192_U489 , R1192_U488 );
and AND2_7660 ( R1192_U167 , R1192_U327 , R1192_U10 );
and AND2_7661 ( R1192_U168 , R1192_U495 , R1192_U212 );
nand NAND2_7662 ( R1192_U169 , R1192_U505 , R1192_U504 );
nand NAND2_7663 ( R1192_U170 , R1192_U510 , R1192_U509 );
and AND2_7664 ( R1192_U171 , R1192_U336 , R1192_U8 );
and AND2_7665 ( R1192_U172 , R1192_U516 , R1192_U211 );
and AND2_7666 ( R1192_U173 , R1192_U390 , R1192_U389 );
nand NAND2_7667 ( R1192_U174 , R1192_U135 , R1192_U345 );
and AND2_7668 ( R1192_U175 , R1192_U399 , R1192_U398 );
and AND2_7669 ( R1192_U176 , R1192_U406 , R1192_U405 );
and AND2_7670 ( R1192_U177 , R1192_U410 , R1192_U409 );
nand NAND2_7671 ( R1192_U178 , R1192_U132 , R1192_U380 );
and AND2_7672 ( R1192_U179 , R1192_U419 , R1192_U418 );
not NOT1_7673 ( R1192_U180 , U4040 );
not NOT1_7674 ( R1192_U181 , U3052 );
and AND2_7675 ( R1192_U182 , R1192_U428 , R1192_U427 );
nand NAND2_7676 ( R1192_U183 , R1192_U148 , R1192_U306 );
and AND2_7677 ( R1192_U184 , R1192_U440 , R1192_U439 );
and AND2_7678 ( R1192_U185 , R1192_U442 , R1192_U441 );
nand NAND2_7679 ( R1192_U186 , R1192_U146 , R1192_U370 );
nand NAND2_7680 ( R1192_U187 , R1192_U357 , R1192_U367 );
nand NAND2_7681 ( R1192_U188 , R1192_U355 , R1192_U365 );
and AND2_7682 ( R1192_U189 , R1192_U461 , R1192_U460 );
nand NAND2_7683 ( R1192_U190 , R1192_U69 , R1192_U315 );
and AND2_7684 ( R1192_U191 , R1192_U465 , R1192_U464 );
nand NAND2_7685 ( R1192_U192 , R1192_U353 , R1192_U363 );
nand NAND2_7686 ( R1192_U193 , R1192_U361 , R1192_U74 );
not NOT1_7687 ( R1192_U194 , U3468 );
nand NAND2_7688 ( R1192_U195 , U3464 , R1192_U109 );
nand NAND2_7689 ( R1192_U196 , R1192_U385 , R1192_U342 );
nand NAND2_7690 ( R1192_U197 , R1192_U144 , R1192_U350 );
nand NAND2_7691 ( R1192_U198 , R1192_U96 , R1192_U282 );
and AND2_7692 ( R1192_U199 , R1192_U497 , R1192_U496 );
and AND2_7693 ( R1192_U200 , R1192_U501 , R1192_U500 );
nand NAND3_7694 ( R1192_U201 , R1192_U349 , R1192_U274 , R1192_U378 );
nand NAND2_7695 ( R1192_U202 , R1192_U376 , R1192_U91 );
nand NAND2_7696 ( R1192_U203 , R1192_U374 , R1192_U270 );
and AND2_7697 ( R1192_U204 , R1192_U518 , R1192_U517 );
nand NAND2_7698 ( R1192_U205 , R1192_U153 , R1192_U186 );
nand NAND2_7699 ( R1192_U206 , R1192_U149 , R1192_U183 );
nand NAND2_7700 ( R1192_U207 , R1192_U195 , R1192_U194 );
not NOT1_7701 ( R1192_U208 , R1192_U99 );
not NOT1_7702 ( R1192_U209 , R1192_U42 );
not NOT1_7703 ( R1192_U210 , R1192_U34 );
nand NAND2_7704 ( R1192_U211 , U3486 , R1192_U86 );
nand NAND2_7705 ( R1192_U212 , U3496 , R1192_U93 );
not NOT1_7706 ( R1192_U213 , R1192_U106 );
nand NAND2_7707 ( R1192_U214 , U4031 , R1192_U98 );
nand NAND2_7708 ( R1192_U215 , U3470 , R1192_U41 );
nand NAND2_7709 ( R1192_U216 , U3476 , R1192_U49 );
nand NAND2_7710 ( R1192_U217 , U3480 , R1192_U33 );
not NOT1_7711 ( R1192_U218 , R1192_U95 );
not NOT1_7712 ( R1192_U219 , R1192_U69 );
not NOT1_7713 ( R1192_U220 , R1192_U51 );
not NOT1_7714 ( R1192_U221 , R1192_U89 );
not NOT1_7715 ( R1192_U222 , R1192_U195 );
nand NAND2_7716 ( R1192_U223 , U3075 , R1192_U195 );
not NOT1_7717 ( R1192_U224 , R1192_U57 );
nand NAND2_7718 ( R1192_U225 , U3472 , R1192_U43 );
nand NAND2_7719 ( R1192_U226 , R1192_U43 , R1192_U42 );
nand NAND2_7720 ( R1192_U227 , R1192_U226 , R1192_U47 );
nand NAND2_7721 ( R1192_U228 , U3061 , R1192_U209 );
nand NAND2_7722 ( R1192_U229 , U3478 , R1192_U48 );
nand NAND2_7723 ( R1192_U230 , U3068 , R1192_U37 );
nand NAND2_7724 ( R1192_U231 , U3064 , R1192_U36 );
nand NAND2_7725 ( R1192_U232 , R1192_U220 , R1192_U216 );
nand NAND2_7726 ( R1192_U233 , R1192_U6 , R1192_U232 );
nand NAND2_7727 ( R1192_U234 , U3474 , R1192_U50 );
nand NAND2_7728 ( R1192_U235 , U3478 , R1192_U48 );
nand NAND2_7729 ( R1192_U236 , R1192_U13 , R1192_U178 );
not NOT1_7730 ( R1192_U237 , R1192_U52 );
not NOT1_7731 ( R1192_U238 , R1192_U55 );
nand NAND2_7732 ( R1192_U239 , U3482 , R1192_U35 );
nand NAND2_7733 ( R1192_U240 , R1192_U35 , R1192_U34 );
nand NAND2_7734 ( R1192_U241 , R1192_U240 , R1192_U40 );
nand NAND2_7735 ( R1192_U242 , U3081 , R1192_U210 );
not NOT1_7736 ( R1192_U243 , R1192_U174 );
nand NAND2_7737 ( R1192_U244 , U3484 , R1192_U54 );
nand NAND2_7738 ( R1192_U245 , R1192_U244 , R1192_U89 );
nand NAND2_7739 ( R1192_U246 , R1192_U238 , R1192_U34 );
nand NAND2_7740 ( R1192_U247 , R1192_U137 , R1192_U246 );
nand NAND2_7741 ( R1192_U248 , R1192_U55 , R1192_U217 );
nand NAND2_7742 ( R1192_U249 , R1192_U136 , R1192_U248 );
nand NAND2_7743 ( R1192_U250 , R1192_U34 , R1192_U217 );
nand NAND2_7744 ( R1192_U251 , R1192_U234 , R1192_U178 );
not NOT1_7745 ( R1192_U252 , R1192_U56 );
nand NAND2_7746 ( R1192_U253 , U3064 , R1192_U36 );
nand NAND2_7747 ( R1192_U254 , R1192_U252 , R1192_U253 );
nand NAND2_7748 ( R1192_U255 , R1192_U139 , R1192_U254 );
nand NAND2_7749 ( R1192_U256 , R1192_U56 , R1192_U216 );
nand NAND2_7750 ( R1192_U257 , U3478 , R1192_U48 );
nand NAND2_7751 ( R1192_U258 , R1192_U138 , R1192_U256 );
nand NAND2_7752 ( R1192_U259 , U3064 , R1192_U36 );
nand NAND2_7753 ( R1192_U260 , R1192_U216 , R1192_U259 );
nand NAND2_7754 ( R1192_U261 , R1192_U234 , R1192_U51 );
nand NAND2_7755 ( R1192_U262 , R1192_U141 , R1192_U384 );
nand NAND2_7756 ( R1192_U263 , R1192_U42 , R1192_U215 );
nand NAND2_7757 ( R1192_U264 , U3488 , R1192_U85 );
nand NAND2_7758 ( R1192_U265 , U3060 , R1192_U87 );
nand NAND2_7759 ( R1192_U266 , U3059 , R1192_U88 );
nand NAND2_7760 ( R1192_U267 , R1192_U221 , R1192_U7 );
nand NAND2_7761 ( R1192_U268 , R1192_U8 , R1192_U267 );
nand NAND2_7762 ( R1192_U269 , U3488 , R1192_U85 );
nand NAND2_7763 ( R1192_U270 , R1192_U269 , R1192_U268 );
nand NAND2_7764 ( R1192_U271 , U3490 , R1192_U90 );
nand NAND2_7765 ( R1192_U272 , U3069 , R1192_U84 );
nand NAND2_7766 ( R1192_U273 , U3492 , R1192_U82 );
nand NAND2_7767 ( R1192_U274 , U3077 , R1192_U83 );
nand NAND2_7768 ( R1192_U275 , U3498 , R1192_U92 );
nand NAND2_7769 ( R1192_U276 , U3070 , R1192_U79 );
nand NAND2_7770 ( R1192_U277 , U3071 , R1192_U80 );
nand NAND2_7771 ( R1192_U278 , R1192_U218 , R1192_U9 );
nand NAND2_7772 ( R1192_U279 , R1192_U10 , R1192_U278 );
nand NAND2_7773 ( R1192_U280 , U3494 , R1192_U94 );
nand NAND2_7774 ( R1192_U281 , U3498 , R1192_U92 );
nand NAND2_7775 ( R1192_U282 , R1192_U16 , R1192_U201 );
not NOT1_7776 ( R1192_U283 , R1192_U96 );
not NOT1_7777 ( R1192_U284 , R1192_U198 );
nand NAND2_7778 ( R1192_U285 , U3500 , R1192_U77 );
nand NAND2_7779 ( R1192_U286 , U3066 , R1192_U78 );
not NOT1_7780 ( R1192_U287 , R1192_U197 );
nand NAND2_7781 ( R1192_U288 , U3502 , R1192_U76 );
nand NAND2_7782 ( R1192_U289 , U3504 , R1192_U72 );
not NOT1_7783 ( R1192_U290 , R1192_U74 );
nand NAND2_7784 ( R1192_U291 , U4037 , R1192_U71 );
nand NAND2_7785 ( R1192_U292 , U3073 , R1192_U73 );
nand NAND2_7786 ( R1192_U293 , U4034 , R1192_U64 );
nand NAND2_7787 ( R1192_U294 , U3063 , R1192_U67 );
nand NAND2_7788 ( R1192_U295 , U3058 , R1192_U68 );
nand NAND2_7789 ( R1192_U296 , R1192_U219 , R1192_U11 );
nand NAND2_7790 ( R1192_U297 , R1192_U12 , R1192_U296 );
nand NAND2_7791 ( R1192_U298 , U4036 , R1192_U66 );
nand NAND2_7792 ( R1192_U299 , U4034 , R1192_U64 );
nand NAND2_7793 ( R1192_U300 , R1192_U299 , R1192_U297 );
nand NAND2_7794 ( R1192_U301 , U4033 , R1192_U62 );
nand NAND2_7795 ( R1192_U302 , U3062 , R1192_U63 );
nand NAND2_7796 ( R1192_U303 , U4032 , R1192_U60 );
nand NAND2_7797 ( R1192_U304 , U3055 , R1192_U61 );
nand NAND2_7798 ( R1192_U305 , U4030 , R1192_U100 );
nand NAND2_7799 ( R1192_U306 , R1192_U147 , R1192_U186 );
nand NAND2_7800 ( R1192_U307 , R1192_U100 , R1192_U99 );
nand NAND2_7801 ( R1192_U308 , R1192_U307 , R1192_U59 );
nand NAND2_7802 ( R1192_U309 , U3050 , R1192_U208 );
not NOT1_7803 ( R1192_U310 , R1192_U183 );
nand NAND2_7804 ( R1192_U311 , U4029 , R1192_U102 );
nand NAND2_7805 ( R1192_U312 , U3051 , R1192_U101 );
nand NAND2_7806 ( R1192_U313 , R1192_U154 , R1192_U205 );
nand NAND2_7807 ( R1192_U314 , R1192_U99 , R1192_U214 );
nand NAND2_7808 ( R1192_U315 , R1192_U298 , R1192_U192 );
not NOT1_7809 ( R1192_U316 , R1192_U190 );
nand NAND2_7810 ( R1192_U317 , U4034 , R1192_U64 );
nand NAND2_7811 ( R1192_U318 , U3058 , R1192_U68 );
nand NAND2_7812 ( R1192_U319 , R1192_U106 , R1192_U318 );
nand NAND2_7813 ( R1192_U320 , R1192_U298 , R1192_U69 );
nand NAND2_7814 ( R1192_U321 , R1192_U280 , R1192_U201 );
not NOT1_7815 ( R1192_U322 , R1192_U107 );
nand NAND2_7816 ( R1192_U323 , U3071 , R1192_U80 );
nand NAND2_7817 ( R1192_U324 , R1192_U322 , R1192_U323 );
nand NAND2_7818 ( R1192_U325 , R1192_U168 , R1192_U324 );
nand NAND2_7819 ( R1192_U326 , R1192_U107 , R1192_U212 );
nand NAND2_7820 ( R1192_U327 , U3498 , R1192_U92 );
nand NAND2_7821 ( R1192_U328 , R1192_U167 , R1192_U326 );
nand NAND2_7822 ( R1192_U329 , U3071 , R1192_U80 );
nand NAND2_7823 ( R1192_U330 , R1192_U212 , R1192_U329 );
nand NAND2_7824 ( R1192_U331 , R1192_U280 , R1192_U95 );
nand NAND2_7825 ( R1192_U332 , U3059 , R1192_U88 );
nand NAND2_7826 ( R1192_U333 , R1192_U373 , R1192_U332 );
nand NAND2_7827 ( R1192_U334 , R1192_U172 , R1192_U333 );
nand NAND2_7828 ( R1192_U335 , R1192_U108 , R1192_U211 );
nand NAND2_7829 ( R1192_U336 , U3488 , R1192_U85 );
nand NAND2_7830 ( R1192_U337 , R1192_U171 , R1192_U335 );
nand NAND2_7831 ( R1192_U338 , U3059 , R1192_U88 );
nand NAND2_7832 ( R1192_U339 , R1192_U211 , R1192_U338 );
nand NAND2_7833 ( R1192_U340 , U3074 , R1192_U45 );
nand NAND2_7834 ( R1192_U341 , U3075 , R1192_U194 );
nand NAND2_7835 ( R1192_U342 , U3079 , R1192_U97 );
nand NAND3_7836 ( R1192_U343 , R1192_U150 , R1192_U306 , R1192_U151 );
nand NAND2_7837 ( R1192_U344 , R1192_U184 , R1192_U205 );
nand NAND2_7838 ( R1192_U345 , R1192_U133 , R1192_U178 );
nand NAND2_7839 ( R1192_U346 , R1192_U237 , R1192_U14 );
nand NAND2_7840 ( R1192_U347 , R1192_U272 , R1192_U270 );
not NOT1_7841 ( R1192_U348 , R1192_U91 );
nand NAND2_7842 ( R1192_U349 , R1192_U348 , R1192_U273 );
nand NAND2_7843 ( R1192_U350 , R1192_U143 , R1192_U201 );
nand NAND2_7844 ( R1192_U351 , R1192_U283 , R1192_U285 );
nand NAND2_7845 ( R1192_U352 , R1192_U290 , R1192_U291 );
not NOT1_7846 ( R1192_U353 , R1192_U105 );
nand NAND2_7847 ( R1192_U354 , R1192_U17 , R1192_U105 );
not NOT1_7848 ( R1192_U355 , R1192_U104 );
nand NAND2_7849 ( R1192_U356 , R1192_U104 , R1192_U301 );
not NOT1_7850 ( R1192_U357 , R1192_U103 );
nand NAND2_7851 ( R1192_U358 , R1192_U103 , R1192_U303 );
nand NAND2_7852 ( R1192_U359 , R1192_U157 , R1192_U192 );
nand NAND2_7853 ( R1192_U360 , R1192_U105 , R1192_U298 );
nand NAND2_7854 ( R1192_U361 , R1192_U289 , R1192_U196 );
not NOT1_7855 ( R1192_U362 , R1192_U193 );
nand NAND2_7856 ( R1192_U363 , R1192_U19 , R1192_U196 );
not NOT1_7857 ( R1192_U364 , R1192_U192 );
nand NAND2_7858 ( R1192_U365 , R1192_U20 , R1192_U196 );
not NOT1_7859 ( R1192_U366 , R1192_U188 );
nand NAND2_7860 ( R1192_U367 , R1192_U21 , R1192_U196 );
not NOT1_7861 ( R1192_U368 , R1192_U187 );
nand NAND2_7862 ( R1192_U369 , R1192_U160 , R1192_U196 );
nand NAND2_7863 ( R1192_U370 , R1192_U145 , R1192_U196 );
not NOT1_7864 ( R1192_U371 , R1192_U186 );
nand NAND2_7865 ( R1192_U372 , R1192_U244 , R1192_U174 );
not NOT1_7866 ( R1192_U373 , R1192_U108 );
nand NAND2_7867 ( R1192_U374 , R1192_U15 , R1192_U174 );
not NOT1_7868 ( R1192_U375 , R1192_U203 );
nand NAND2_7869 ( R1192_U376 , R1192_U18 , R1192_U174 );
not NOT1_7870 ( R1192_U377 , R1192_U202 );
nand NAND2_7871 ( R1192_U378 , R1192_U142 , R1192_U174 );
not NOT1_7872 ( R1192_U379 , R1192_U201 );
nand NAND2_7873 ( R1192_U380 , R1192_U131 , R1192_U57 );
not NOT1_7874 ( R1192_U381 , R1192_U178 );
nand NAND2_7875 ( R1192_U382 , R1192_U215 , R1192_U57 );
nand NAND2_7876 ( R1192_U383 , R1192_U140 , R1192_U382 );
nand NAND2_7877 ( R1192_U384 , R1192_U224 , R1192_U42 );
nand NAND2_7878 ( R1192_U385 , R1192_U288 , R1192_U197 );
not NOT1_7879 ( R1192_U386 , R1192_U196 );
nand NAND2_7880 ( R1192_U387 , R1192_U158 , R1192_U12 );
nand NAND2_7881 ( R1192_U388 , R1192_U159 , R1192_U457 );
nand NAND2_7882 ( R1192_U389 , U3484 , R1192_U54 );
nand NAND2_7883 ( R1192_U390 , U3080 , R1192_U53 );
nand NAND2_7884 ( R1192_U391 , R1192_U245 , R1192_U174 );
nand NAND2_7885 ( R1192_U392 , R1192_U243 , R1192_U173 );
nand NAND2_7886 ( R1192_U393 , U3482 , R1192_U35 );
nand NAND2_7887 ( R1192_U394 , U3081 , R1192_U40 );
nand NAND2_7888 ( R1192_U395 , U3482 , R1192_U35 );
nand NAND2_7889 ( R1192_U396 , U3081 , R1192_U40 );
nand NAND2_7890 ( R1192_U397 , R1192_U396 , R1192_U395 );
nand NAND2_7891 ( R1192_U398 , U3480 , R1192_U33 );
nand NAND2_7892 ( R1192_U399 , U3067 , R1192_U39 );
nand NAND2_7893 ( R1192_U400 , R1192_U250 , R1192_U55 );
nand NAND2_7894 ( R1192_U401 , R1192_U175 , R1192_U238 );
nand NAND2_7895 ( R1192_U402 , U3478 , R1192_U48 );
nand NAND2_7896 ( R1192_U403 , U3068 , R1192_U37 );
nand NAND2_7897 ( R1192_U404 , R1192_U403 , R1192_U402 );
nand NAND2_7898 ( R1192_U405 , U3476 , R1192_U49 );
nand NAND2_7899 ( R1192_U406 , U3064 , R1192_U36 );
nand NAND2_7900 ( R1192_U407 , R1192_U260 , R1192_U56 );
nand NAND2_7901 ( R1192_U408 , R1192_U176 , R1192_U252 );
nand NAND2_7902 ( R1192_U409 , U3474 , R1192_U50 );
nand NAND2_7903 ( R1192_U410 , U3057 , R1192_U38 );
nand NAND2_7904 ( R1192_U411 , R1192_U178 , R1192_U261 );
nand NAND2_7905 ( R1192_U412 , R1192_U381 , R1192_U177 );
nand NAND2_7906 ( R1192_U413 , U3472 , R1192_U43 );
nand NAND2_7907 ( R1192_U414 , U3061 , R1192_U47 );
nand NAND2_7908 ( R1192_U415 , U3472 , R1192_U43 );
nand NAND2_7909 ( R1192_U416 , U3061 , R1192_U47 );
nand NAND2_7910 ( R1192_U417 , R1192_U416 , R1192_U415 );
nand NAND2_7911 ( R1192_U418 , U3470 , R1192_U41 );
nand NAND2_7912 ( R1192_U419 , U3065 , R1192_U44 );
nand NAND2_7913 ( R1192_U420 , R1192_U263 , R1192_U57 );
nand NAND2_7914 ( R1192_U421 , R1192_U179 , R1192_U224 );
nand NAND2_7915 ( R1192_U422 , U4040 , R1192_U181 );
nand NAND2_7916 ( R1192_U423 , U3052 , R1192_U180 );
nand NAND2_7917 ( R1192_U424 , U4040 , R1192_U181 );
nand NAND2_7918 ( R1192_U425 , U3052 , R1192_U180 );
nand NAND2_7919 ( R1192_U426 , R1192_U425 , R1192_U424 );
nand NAND3_7920 ( R1192_U427 , U4029 , R1192_U23 , R1192_U102 );
nand NAND3_7921 ( R1192_U428 , R1192_U426 , R1192_U101 , U3051 );
nand NAND2_7922 ( R1192_U429 , U4029 , R1192_U102 );
nand NAND2_7923 ( R1192_U430 , U3051 , R1192_U101 );
not NOT1_7924 ( R1192_U431 , R1192_U152 );
nand NAND2_7925 ( R1192_U432 , R1192_U310 , R1192_U431 );
nand NAND2_7926 ( R1192_U433 , R1192_U152 , R1192_U183 );
nand NAND2_7927 ( R1192_U434 , U4030 , R1192_U100 );
nand NAND2_7928 ( R1192_U435 , U3050 , R1192_U59 );
nand NAND2_7929 ( R1192_U436 , R1192_U435 , R1192_U434 );
nand NAND2_7930 ( R1192_U437 , U4030 , R1192_U100 );
nand NAND2_7931 ( R1192_U438 , U3050 , R1192_U59 );
nand NAND3_7932 ( R1192_U439 , R1192_U438 , R1192_U437 , R1192_U99 );
nand NAND2_7933 ( R1192_U440 , R1192_U436 , R1192_U208 );
nand NAND2_7934 ( R1192_U441 , U4031 , R1192_U98 );
nand NAND2_7935 ( R1192_U442 , U3054 , R1192_U58 );
nand NAND2_7936 ( R1192_U443 , R1192_U186 , R1192_U314 );
nand NAND2_7937 ( R1192_U444 , R1192_U371 , R1192_U185 );
nand NAND2_7938 ( R1192_U445 , U4032 , R1192_U60 );
nand NAND2_7939 ( R1192_U446 , U3055 , R1192_U61 );
not NOT1_7940 ( R1192_U447 , R1192_U155 );
nand NAND2_7941 ( R1192_U448 , R1192_U368 , R1192_U447 );
nand NAND2_7942 ( R1192_U449 , R1192_U155 , R1192_U187 );
nand NAND2_7943 ( R1192_U450 , U4033 , R1192_U62 );
nand NAND2_7944 ( R1192_U451 , U3062 , R1192_U63 );
not NOT1_7945 ( R1192_U452 , R1192_U156 );
nand NAND2_7946 ( R1192_U453 , R1192_U366 , R1192_U452 );
nand NAND2_7947 ( R1192_U454 , R1192_U156 , R1192_U188 );
nand NAND2_7948 ( R1192_U455 , U4034 , R1192_U64 );
nand NAND2_7949 ( R1192_U456 , U3063 , R1192_U67 );
nand NAND2_7950 ( R1192_U457 , R1192_U456 , R1192_U455 );
nand NAND3_7951 ( R1192_U458 , R1192_U161 , R1192_U369 , R1192_U69 );
nand NAND2_7952 ( R1192_U459 , R1192_U22 , R1192_U219 );
nand NAND2_7953 ( R1192_U460 , U4035 , R1192_U65 );
nand NAND2_7954 ( R1192_U461 , U3058 , R1192_U68 );
nand NAND2_7955 ( R1192_U462 , R1192_U319 , R1192_U190 );
nand NAND2_7956 ( R1192_U463 , R1192_U316 , R1192_U189 );
nand NAND2_7957 ( R1192_U464 , U4036 , R1192_U66 );
nand NAND2_7958 ( R1192_U465 , U3072 , R1192_U70 );
nand NAND2_7959 ( R1192_U466 , R1192_U192 , R1192_U320 );
nand NAND2_7960 ( R1192_U467 , R1192_U364 , R1192_U191 );
nand NAND2_7961 ( R1192_U468 , U4037 , R1192_U71 );
nand NAND2_7962 ( R1192_U469 , U3073 , R1192_U73 );
not NOT1_7963 ( R1192_U470 , R1192_U162 );
nand NAND2_7964 ( R1192_U471 , R1192_U362 , R1192_U470 );
nand NAND2_7965 ( R1192_U472 , R1192_U162 , R1192_U193 );
nand NAND2_7966 ( R1192_U473 , U3468 , R1192_U46 );
nand NAND2_7967 ( R1192_U474 , U3075 , R1192_U194 );
not NOT1_7968 ( R1192_U475 , R1192_U163 );
nand NAND2_7969 ( R1192_U476 , R1192_U222 , R1192_U475 );
nand NAND2_7970 ( R1192_U477 , R1192_U163 , R1192_U195 );
nand NAND2_7971 ( R1192_U478 , U3504 , R1192_U72 );
nand NAND2_7972 ( R1192_U479 , U3078 , R1192_U75 );
not NOT1_7973 ( R1192_U480 , R1192_U164 );
nand NAND2_7974 ( R1192_U481 , R1192_U386 , R1192_U480 );
nand NAND2_7975 ( R1192_U482 , R1192_U164 , R1192_U196 );
nand NAND2_7976 ( R1192_U483 , U3502 , R1192_U76 );
nand NAND2_7977 ( R1192_U484 , U3079 , R1192_U97 );
not NOT1_7978 ( R1192_U485 , R1192_U165 );
nand NAND2_7979 ( R1192_U486 , R1192_U287 , R1192_U485 );
nand NAND2_7980 ( R1192_U487 , R1192_U165 , R1192_U197 );
nand NAND2_7981 ( R1192_U488 , U3500 , R1192_U77 );
nand NAND2_7982 ( R1192_U489 , U3066 , R1192_U78 );
not NOT1_7983 ( R1192_U490 , R1192_U166 );
nand NAND2_7984 ( R1192_U491 , R1192_U284 , R1192_U490 );
nand NAND2_7985 ( R1192_U492 , R1192_U166 , R1192_U198 );
nand NAND2_7986 ( R1192_U493 , U3498 , R1192_U92 );
nand NAND2_7987 ( R1192_U494 , U3070 , R1192_U79 );
nand NAND2_7988 ( R1192_U495 , R1192_U494 , R1192_U493 );
nand NAND2_7989 ( R1192_U496 , U3496 , R1192_U93 );
nand NAND2_7990 ( R1192_U497 , U3071 , R1192_U80 );
nand NAND2_7991 ( R1192_U498 , R1192_U330 , R1192_U107 );
nand NAND2_7992 ( R1192_U499 , R1192_U199 , R1192_U322 );
nand NAND2_7993 ( R1192_U500 , U3494 , R1192_U94 );
nand NAND2_7994 ( R1192_U501 , U3076 , R1192_U81 );
nand NAND2_7995 ( R1192_U502 , R1192_U201 , R1192_U331 );
nand NAND2_7996 ( R1192_U503 , R1192_U379 , R1192_U200 );
nand NAND2_7997 ( R1192_U504 , U3492 , R1192_U82 );
nand NAND2_7998 ( R1192_U505 , U3077 , R1192_U83 );
not NOT1_7999 ( R1192_U506 , R1192_U169 );
nand NAND2_8000 ( R1192_U507 , R1192_U377 , R1192_U506 );
nand NAND2_8001 ( R1192_U508 , R1192_U169 , R1192_U202 );
nand NAND2_8002 ( R1192_U509 , U3490 , R1192_U90 );
nand NAND2_8003 ( R1192_U510 , U3069 , R1192_U84 );
not NOT1_8004 ( R1192_U511 , R1192_U170 );
nand NAND2_8005 ( R1192_U512 , R1192_U375 , R1192_U511 );
nand NAND2_8006 ( R1192_U513 , R1192_U170 , R1192_U203 );
nand NAND2_8007 ( R1192_U514 , U3488 , R1192_U85 );
nand NAND2_8008 ( R1192_U515 , U3060 , R1192_U87 );
nand NAND2_8009 ( R1192_U516 , R1192_U515 , R1192_U514 );
nand NAND2_8010 ( R1192_U517 , U3486 , R1192_U86 );
nand NAND2_8011 ( R1192_U518 , U3059 , R1192_U88 );
nand NAND2_8012 ( R1192_U519 , R1192_U108 , R1192_U339 );
nand NAND2_8013 ( R1192_U520 , R1192_U204 , R1192_U373 );
and AND4_8014 ( R1347_U6 , R1347_U143 , R1347_U142 , R1347_U141 , R1347_U139 );
and AND2_8015 ( R1347_U7 , R1347_U84 , R1347_U6 );
and AND2_8016 ( R1347_U8 , R1347_U7 , R1347_U147 );
and AND2_8017 ( R1347_U9 , R1347_U181 , R1347_U180 );
and AND2_8018 ( R1347_U10 , R1347_U83 , R1347_U11 );
and AND3_8019 ( R1347_U11 , R1347_U78 , R1347_U183 , R1347_U79 );
and AND2_8020 ( R1347_U12 , R1347_U209 , R1347_U132 );
and AND2_8021 ( R1347_U13 , R1347_U198 , R1347_U118 );
not NOT1_8022 ( R1347_U14 , U3596 );
not NOT1_8023 ( R1347_U15 , U3486 );
not NOT1_8024 ( R1347_U16 , U3484 );
not NOT1_8025 ( R1347_U17 , U3480 );
not NOT1_8026 ( R1347_U18 , U3482 );
not NOT1_8027 ( R1347_U19 , U3478 );
not NOT1_8028 ( R1347_U20 , U3476 );
not NOT1_8029 ( R1347_U21 , U3474 );
not NOT1_8030 ( R1347_U22 , U3472 );
not NOT1_8031 ( R1347_U23 , U3612 );
not NOT1_8032 ( R1347_U24 , U3470 );
not NOT1_8033 ( R1347_U25 , U3468 );
not NOT1_8034 ( R1347_U26 , U3498 );
not NOT1_8035 ( R1347_U27 , U3496 );
not NOT1_8036 ( R1347_U28 , U3608 );
not NOT1_8037 ( R1347_U29 , U3490 );
not NOT1_8038 ( R1347_U30 , U3609 );
nand NAND2_8039 ( R1347_U31 , R1347_U153 , R1347_U152 );
not NOT1_8040 ( R1347_U32 , U3488 );
not NOT1_8041 ( R1347_U33 , U3492 );
not NOT1_8042 ( R1347_U34 , U3494 );
not NOT1_8043 ( R1347_U35 , U4036 );
not NOT1_8044 ( R1347_U36 , U4035 );
not NOT1_8045 ( R1347_U37 , U3602 );
not NOT1_8046 ( R1347_U38 , U3502 );
not NOT1_8047 ( R1347_U39 , U3603 );
nand NAND2_8048 ( R1347_U40 , R1347_U135 , R1347_U136 );
not NOT1_8049 ( R1347_U41 , U3500 );
not NOT1_8050 ( R1347_U42 , U3504 );
not NOT1_8051 ( R1347_U43 , U4037 );
not NOT1_8052 ( R1347_U44 , U3601 );
not NOT1_8053 ( R1347_U45 , U3590 );
not NOT1_8054 ( R1347_U46 , U3587 );
not NOT1_8055 ( R1347_U47 , U3586 );
not NOT1_8056 ( R1347_U48 , U3585 );
not NOT1_8057 ( R1347_U49 , U3584 );
not NOT1_8058 ( R1347_U50 , U3583 );
not NOT1_8059 ( R1347_U51 , U3582 );
not NOT1_8060 ( R1347_U52 , U3611 );
not NOT1_8061 ( R1347_U53 , U3610 );
not NOT1_8062 ( R1347_U54 , U3607 );
not NOT1_8063 ( R1347_U55 , U3606 );
not NOT1_8064 ( R1347_U56 , U3605 );
not NOT1_8065 ( R1347_U57 , U3604 );
not NOT1_8066 ( R1347_U58 , U3600 );
not NOT1_8067 ( R1347_U59 , U3599 );
not NOT1_8068 ( R1347_U60 , U3598 );
not NOT1_8069 ( R1347_U61 , U3597 );
not NOT1_8070 ( R1347_U62 , U4034 );
not NOT1_8071 ( R1347_U63 , U4033 );
not NOT1_8072 ( R1347_U64 , U4031 );
not NOT1_8073 ( R1347_U65 , U4030 );
not NOT1_8074 ( R1347_U66 , U3588 );
not NOT1_8075 ( R1347_U67 , U4039 );
not NOT1_8076 ( R1347_U68 , U3589 );
not NOT1_8077 ( R1347_U69 , U4038 );
not NOT1_8078 ( R1347_U70 , U3592 );
not NOT1_8079 ( R1347_U71 , U3593 );
not NOT1_8080 ( R1347_U72 , U3594 );
and AND2_8081 ( R1347_U73 , U3464 , R1347_U121 );
and AND2_8082 ( R1347_U74 , U3490 , R1347_U30 );
and AND2_8083 ( R1347_U75 , U3488 , R1347_U53 );
and AND2_8084 ( R1347_U76 , U3502 , R1347_U39 );
and AND2_8085 ( R1347_U77 , U3500 , R1347_U57 );
and AND2_8086 ( R1347_U78 , R1347_U184 , R1347_U182 );
and AND2_8087 ( R1347_U79 , R1347_U9 , R1347_U185 );
and AND2_8088 ( R1347_U80 , R1347_U138 , R1347_U134 );
and AND2_8089 ( R1347_U81 , R1347_U80 , R1347_U172 );
and AND2_8090 ( R1347_U82 , R1347_U175 , R1347_U174 );
and AND3_8091 ( R1347_U83 , R1347_U81 , R1347_U173 , R1347_U82 );
and AND3_8092 ( R1347_U84 , R1347_U145 , R1347_U144 , R1347_U146 );
and AND2_8093 ( R1347_U85 , R1347_U149 , R1347_U150 );
and AND2_8094 ( R1347_U86 , R1347_U85 , R1347_U148 );
and AND2_8095 ( R1347_U87 , U3590 , R1347_U22 );
and AND2_8096 ( R1347_U88 , R1347_U7 , R1347_U87 );
and AND2_8097 ( R1347_U89 , R1347_U145 , R1347_U144 );
and AND2_8098 ( R1347_U90 , R1347_U162 , R1347_U163 );
and AND2_8099 ( R1347_U91 , R1347_U6 , R1347_U164 );
and AND2_8100 ( R1347_U92 , R1347_U141 , R1347_U139 );
and AND2_8101 ( R1347_U93 , R1347_U92 , R1347_U157 );
and AND2_8102 ( R1347_U94 , U3611 , R1347_U15 );
and AND2_8103 ( R1347_U95 , U3610 , R1347_U32 );
and AND4_8104 ( R1347_U96 , R1347_U134 , R1347_U34 , U3607 , R1347_U138 );
and AND2_8105 ( R1347_U97 , U3606 , R1347_U27 );
and AND2_8106 ( R1347_U98 , R1347_U134 , R1347_U97 );
and AND2_8107 ( R1347_U99 , U3605 , R1347_U26 );
and AND2_8108 ( R1347_U100 , U3604 , R1347_U41 );
and AND2_8109 ( R1347_U101 , U3600 , R1347_U43 );
and AND2_8110 ( R1347_U102 , U3599 , R1347_U35 );
and AND3_8111 ( R1347_U103 , R1347_U151 , R1347_U133 , R1347_U165 );
and AND2_8112 ( R1347_U104 , R1347_U167 , R1347_U166 );
and AND4_8113 ( R1347_U105 , R1347_U176 , R1347_U170 , R1347_U169 , R1347_U168 );
and AND2_8114 ( R1347_U106 , R1347_U178 , R1347_U177 );
and AND2_8115 ( R1347_U107 , R1347_U108 , R1347_U179 );
and AND2_8116 ( R1347_U108 , R1347_U188 , R1347_U186 );
and AND2_8117 ( R1347_U109 , R1347_U190 , R1347_U189 );
and AND2_8118 ( R1347_U110 , R1347_U109 , R1347_U206 );
and AND4_8119 ( R1347_U111 , R1347_U110 , R1347_U207 , R1347_U106 , R1347_U107 );
and AND2_8120 ( R1347_U112 , U4034 , R1347_U61 );
and AND2_8121 ( R1347_U113 , R1347_U192 , R1347_U193 );
and AND2_8122 ( R1347_U114 , R1347_U132 , R1347_U123 );
and AND2_8123 ( R1347_U115 , R1347_U12 , R1347_U197 );
and AND2_8124 ( R1347_U116 , R1347_U115 , R1347_U210 );
and AND2_8125 ( R1347_U117 , U3589 , R1347_U67 );
and AND2_8126 ( R1347_U118 , R1347_U212 , R1347_U120 );
and AND3_8127 ( R1347_U119 , R1347_U199 , R1347_U201 , R1347_U204 );
and AND2_8128 ( R1347_U120 , R1347_U119 , R1347_U205 );
not NOT1_8129 ( R1347_U121 , U3613 );
not NOT1_8130 ( R1347_U122 , U4040 );
not NOT1_8131 ( R1347_U123 , U4029 );
not NOT1_8132 ( R1347_U124 , U3595 );
nand NAND2_8133 ( R1347_U125 , R1347_U203 , R1347_U202 );
nand NAND2_8134 ( R1347_U126 , R1347_U208 , R1347_U131 );
nand NAND2_8135 ( R1347_U127 , U4032 , R1347_U194 );
nand NAND2_8136 ( R1347_U128 , U3588 , R1347_U69 );
nand NAND3_8137 ( R1347_U129 , R1347_U130 , R1347_U122 , R1347_U128 );
nand NAND2_8138 ( R1347_U130 , U4039 , R1347_U68 );
nand NAND2_8139 ( R1347_U131 , R1347_U114 , R1347_U209 );
nand NAND2_8140 ( R1347_U132 , U4030 , R1347_U71 );
nand NAND2_8141 ( R1347_U133 , U3596 , R1347_U63 );
nand NAND2_8142 ( R1347_U134 , U3498 , R1347_U56 );
nand NAND2_8143 ( R1347_U135 , U3602 , R1347_U42 );
nand NAND2_8144 ( R1347_U136 , U3603 , R1347_U38 );
not NOT1_8145 ( R1347_U137 , R1347_U40 );
nand NAND2_8146 ( R1347_U138 , U3496 , R1347_U55 );
nand NAND2_8147 ( R1347_U139 , U3486 , R1347_U52 );
nand NAND2_8148 ( R1347_U140 , U3612 , R1347_U25 );
nand NAND2_8149 ( R1347_U141 , U3484 , R1347_U51 );
nand NAND2_8150 ( R1347_U142 , U3480 , R1347_U49 );
nand NAND2_8151 ( R1347_U143 , U3482 , R1347_U50 );
nand NAND2_8152 ( R1347_U144 , U3478 , R1347_U48 );
nand NAND2_8153 ( R1347_U145 , U3476 , R1347_U47 );
nand NAND2_8154 ( R1347_U146 , U3474 , R1347_U46 );
nand NAND2_8155 ( R1347_U147 , U3472 , R1347_U45 );
nand NAND2_8156 ( R1347_U148 , R1347_U73 , R1347_U140 );
nand NAND2_8157 ( R1347_U149 , U3470 , R1347_U44 );
nand NAND2_8158 ( R1347_U150 , U3468 , R1347_U23 );
nand NAND3_8159 ( R1347_U151 , R1347_U8 , R1347_U86 , R1347_U10 );
nand NAND2_8160 ( R1347_U152 , U3609 , R1347_U29 );
nand NAND2_8161 ( R1347_U153 , U3608 , R1347_U33 );
not NOT1_8162 ( R1347_U154 , R1347_U31 );
nand NAND2_8163 ( R1347_U155 , U3583 , R1347_U18 );
nand NAND2_8164 ( R1347_U156 , U3582 , R1347_U16 );
nand NAND2_8165 ( R1347_U157 , R1347_U156 , R1347_U155 );
nand NAND2_8166 ( R1347_U158 , U3587 , R1347_U21 );
nand NAND2_8167 ( R1347_U159 , U3586 , R1347_U20 );
nand NAND2_8168 ( R1347_U160 , R1347_U159 , R1347_U158 );
nand NAND2_8169 ( R1347_U161 , R1347_U89 , R1347_U160 );
nand NAND2_8170 ( R1347_U162 , U3585 , R1347_U19 );
nand NAND2_8171 ( R1347_U163 , U3584 , R1347_U17 );
nand NAND2_8172 ( R1347_U164 , R1347_U90 , R1347_U161 );
nand NAND4_8173 ( R1347_U165 , U3601 , R1347_U8 , R1347_U10 , R1347_U24 );
nand NAND2_8174 ( R1347_U166 , R1347_U88 , R1347_U10 );
nand NAND2_8175 ( R1347_U167 , R1347_U91 , R1347_U10 );
nand NAND2_8176 ( R1347_U168 , R1347_U93 , R1347_U10 );
nand NAND2_8177 ( R1347_U169 , R1347_U94 , R1347_U10 );
nand NAND2_8178 ( R1347_U170 , R1347_U95 , R1347_U10 );
nand NAND2_8179 ( R1347_U171 , U3608 , R1347_U33 );
nand NAND2_8180 ( R1347_U172 , R1347_U74 , R1347_U171 );
nand NAND2_8181 ( R1347_U173 , R1347_U75 , R1347_U154 );
nand NAND2_8182 ( R1347_U174 , U3492 , R1347_U28 );
nand NAND2_8183 ( R1347_U175 , U3494 , R1347_U54 );
nand NAND2_8184 ( R1347_U176 , R1347_U96 , R1347_U11 );
nand NAND2_8185 ( R1347_U177 , R1347_U98 , R1347_U11 );
nand NAND2_8186 ( R1347_U178 , R1347_U99 , R1347_U11 );
nand NAND2_8187 ( R1347_U179 , R1347_U100 , R1347_U11 );
nand NAND2_8188 ( R1347_U180 , U4036 , R1347_U59 );
nand NAND2_8189 ( R1347_U181 , U4035 , R1347_U60 );
nand NAND2_8190 ( R1347_U182 , R1347_U76 , R1347_U135 );
nand NAND2_8191 ( R1347_U183 , R1347_U77 , R1347_U137 );
nand NAND2_8192 ( R1347_U184 , U3504 , R1347_U37 );
nand NAND2_8193 ( R1347_U185 , U4037 , R1347_U58 );
nand NAND2_8194 ( R1347_U186 , R1347_U101 , R1347_U9 );
nand NAND2_8195 ( R1347_U187 , U4035 , R1347_U60 );
nand NAND2_8196 ( R1347_U188 , R1347_U102 , R1347_U187 );
nand NAND2_8197 ( R1347_U189 , U3598 , R1347_U36 );
nand NAND2_8198 ( R1347_U190 , U3597 , R1347_U62 );
nand NAND4_8199 ( R1347_U191 , R1347_U104 , R1347_U103 , R1347_U105 , R1347_U111 );
nand NAND2_8200 ( R1347_U192 , R1347_U112 , R1347_U133 );
nand NAND2_8201 ( R1347_U193 , U4033 , R1347_U14 );
nand NAND2_8202 ( R1347_U194 , R1347_U113 , R1347_U191 );
nand NAND2_8203 ( R1347_U195 , U4032 , R1347_U124 );
nand NAND2_8204 ( R1347_U196 , R1347_U194 , R1347_U124 );
nand NAND2_8205 ( R1347_U197 , U4031 , R1347_U72 );
nand NAND4_8206 ( R1347_U198 , R1347_U195 , R1347_U127 , R1347_U116 , R1347_U196 );
nand NAND2_8207 ( R1347_U199 , R1347_U117 , R1347_U128 );
nand NAND2_8208 ( R1347_U200 , U4039 , R1347_U68 );
nand NAND4_8209 ( R1347_U201 , R1347_U200 , R1347_U122 , R1347_U128 , U3591 );
nand NAND2_8210 ( R1347_U202 , U3593 , R1347_U65 );
nand NAND2_8211 ( R1347_U203 , U3594 , R1347_U64 );
nand NAND2_8212 ( R1347_U204 , U4038 , R1347_U66 );
nand NAND3_8213 ( R1347_U205 , R1347_U209 , R1347_U123 , U3592 );
nand NAND2_8214 ( R1347_U206 , R1347_U11 , R1347_U40 );
nand NAND2_8215 ( R1347_U207 , R1347_U10 , R1347_U31 );
nand NAND2_8216 ( R1347_U208 , U3592 , R1347_U12 );
nand NAND2_8217 ( R1347_U209 , R1347_U129 , R1347_U211 );
nand NAND2_8218 ( R1347_U210 , R1347_U131 , R1347_U70 );
nand NAND3_8219 ( R1347_U211 , R1347_U130 , R1347_U128 , U3591 );
nand NAND2_8220 ( R1347_U212 , R1347_U126 , R1347_U125 );
and AND2_8221 ( R1171_U4 , R1171_U196 , R1171_U195 );
and AND2_8222 ( R1171_U5 , R1171_U197 , R1171_U198 );
and AND2_8223 ( R1171_U6 , R1171_U210 , R1171_U209 );
and AND2_8224 ( R1171_U7 , R1171_U250 , R1171_U249 );
and AND2_8225 ( R1171_U8 , R1171_U258 , R1171_U257 );
and AND2_8226 ( R1171_U9 , R1171_U274 , R1171_U273 );
and AND2_8227 ( R1171_U10 , R1171_U282 , R1171_U281 );
and AND2_8228 ( R1171_U11 , R1171_U10 , R1171_U283 );
and AND2_8229 ( R1171_U12 , R1171_U7 , R1171_U217 );
and AND2_8230 ( R1171_U13 , R1171_U8 , R1171_U262 );
and AND2_8231 ( R1171_U14 , R1171_U11 , R1171_U292 );
and AND2_8232 ( R1171_U15 , R1171_U13 , R1171_U267 );
and AND2_8233 ( R1171_U16 , R1171_U9 , R1171_U14 );
and AND2_8234 ( R1171_U17 , R1171_U299 , R1171_U305 );
and AND2_8235 ( R1171_U18 , R1171_U359 , R1171_U356 );
and AND2_8236 ( R1171_U19 , R1171_U352 , R1171_U349 );
and AND2_8237 ( R1171_U20 , R1171_U343 , R1171_U340 );
and AND2_8238 ( R1171_U21 , R1171_U334 , R1171_U331 );
and AND2_8239 ( R1171_U22 , R1171_U328 , R1171_U326 );
and AND2_8240 ( R1171_U23 , R1171_U321 , R1171_U318 );
and AND2_8241 ( R1171_U24 , R1171_U248 , R1171_U245 );
and AND2_8242 ( R1171_U25 , R1171_U240 , R1171_U237 );
and AND2_8243 ( R1171_U26 , R1171_U226 , R1171_U223 );
not NOT1_8244 ( R1171_U27 , U3470 );
not NOT1_8245 ( R1171_U28 , U3065 );
not NOT1_8246 ( R1171_U29 , U3472 );
not NOT1_8247 ( R1171_U30 , U3061 );
not NOT1_8248 ( R1171_U31 , U3474 );
not NOT1_8249 ( R1171_U32 , U3057 );
not NOT1_8250 ( R1171_U33 , U3064 );
nand NAND2_8251 ( R1171_U34 , U3057 , U3474 );
not NOT1_8252 ( R1171_U35 , U3476 );
nand NAND2_8253 ( R1171_U36 , U3468 , U3075 );
not NOT1_8254 ( R1171_U37 , U3464 );
not NOT1_8255 ( R1171_U38 , U3074 );
nand NAND2_8256 ( R1171_U39 , R1171_U131 , R1171_U200 );
not NOT1_8257 ( R1171_U40 , U3478 );
not NOT1_8258 ( R1171_U41 , U3068 );
not NOT1_8259 ( R1171_U42 , U3067 );
nand NAND2_8260 ( R1171_U43 , U3068 , U3478 );
not NOT1_8261 ( R1171_U44 , U3480 );
nand NAND2_8262 ( R1171_U45 , R1171_U214 , R1171_U213 );
not NOT1_8263 ( R1171_U46 , U3482 );
not NOT1_8264 ( R1171_U47 , U3081 );
not NOT1_8265 ( R1171_U48 , U3080 );
not NOT1_8266 ( R1171_U49 , U3484 );
nand NAND2_8267 ( R1171_U50 , R1171_U65 , R1171_U218 );
nand NAND2_8268 ( R1171_U51 , R1171_U133 , R1171_U132 );
nand NAND2_8269 ( R1171_U52 , R1171_U136 , R1171_U232 );
nand NAND2_8270 ( R1171_U53 , R1171_U229 , R1171_U228 );
not NOT1_8271 ( R1171_U54 , U4030 );
not NOT1_8272 ( R1171_U55 , U3050 );
not NOT1_8273 ( R1171_U56 , U3054 );
not NOT1_8274 ( R1171_U57 , U4031 );
not NOT1_8275 ( R1171_U58 , U4033 );
not NOT1_8276 ( R1171_U59 , U3062 );
nand NAND2_8277 ( R1171_U60 , U3062 , U4033 );
not NOT1_8278 ( R1171_U61 , U4035 );
not NOT1_8279 ( R1171_U62 , U3058 );
not NOT1_8280 ( R1171_U63 , U3496 );
not NOT1_8281 ( R1171_U64 , U3071 );
nand NAND2_8282 ( R1171_U65 , U3081 , U3482 );
not NOT1_8283 ( R1171_U66 , U3486 );
not NOT1_8284 ( R1171_U67 , U3059 );
not NOT1_8285 ( R1171_U68 , U3490 );
not NOT1_8286 ( R1171_U69 , U3069 );
not NOT1_8287 ( R1171_U70 , U3488 );
not NOT1_8288 ( R1171_U71 , U3060 );
nand NAND2_8289 ( R1171_U72 , U3060 , U3488 );
not NOT1_8290 ( R1171_U73 , U3492 );
not NOT1_8291 ( R1171_U74 , U3077 );
not NOT1_8292 ( R1171_U75 , U3494 );
not NOT1_8293 ( R1171_U76 , U3076 );
nand NAND2_8294 ( R1171_U77 , R1171_U380 , R1171_U267 );
not NOT1_8295 ( R1171_U78 , U3504 );
not NOT1_8296 ( R1171_U79 , U3078 );
nand NAND2_8297 ( R1171_U80 , U3078 , U3504 );
not NOT1_8298 ( R1171_U81 , U4037 );
not NOT1_8299 ( R1171_U82 , U3502 );
not NOT1_8300 ( R1171_U83 , U3079 );
nand NAND2_8301 ( R1171_U84 , U3079 , U3502 );
not NOT1_8302 ( R1171_U85 , U4036 );
not NOT1_8303 ( R1171_U86 , U3072 );
not NOT1_8304 ( R1171_U87 , U3498 );
not NOT1_8305 ( R1171_U88 , U3070 );
not NOT1_8306 ( R1171_U89 , U3066 );
nand NAND2_8307 ( R1171_U90 , U3070 , U3498 );
not NOT1_8308 ( R1171_U91 , U3500 );
not NOT1_8309 ( R1171_U92 , U4034 );
not NOT1_8310 ( R1171_U93 , U3063 );
nand NAND2_8311 ( R1171_U94 , R1171_U146 , R1171_U388 );
not NOT1_8312 ( R1171_U95 , U4032 );
not NOT1_8313 ( R1171_U96 , U3055 );
nand NAND3_8314 ( R1171_U97 , R1171_U396 , R1171_U306 , R1171_U397 );
not NOT1_8315 ( R1171_U98 , U3051 );
not NOT1_8316 ( R1171_U99 , U4029 );
nand NAND2_8317 ( R1171_U100 , R1171_U60 , R1171_U314 );
nand NAND2_8318 ( R1171_U101 , R1171_U385 , R1171_U294 );
nand NAND2_8319 ( R1171_U102 , R1171_U278 , R1171_U277 );
not NOT1_8320 ( R1171_U103 , U3073 );
nand NAND2_8321 ( R1171_U104 , R1171_U84 , R1171_U323 );
nand NAND3_8322 ( R1171_U105 , R1171_U383 , R1171_U271 , R1171_U382 );
nand NAND2_8323 ( R1171_U106 , R1171_U72 , R1171_U345 );
nand NAND2_8324 ( R1171_U107 , R1171_U484 , R1171_U483 );
nand NAND2_8325 ( R1171_U108 , R1171_U531 , R1171_U530 );
nand NAND2_8326 ( R1171_U109 , R1171_U402 , R1171_U401 );
nand NAND2_8327 ( R1171_U110 , R1171_U407 , R1171_U406 );
nand NAND2_8328 ( R1171_U111 , R1171_U414 , R1171_U413 );
nand NAND2_8329 ( R1171_U112 , R1171_U421 , R1171_U420 );
nand NAND2_8330 ( R1171_U113 , R1171_U426 , R1171_U425 );
nand NAND2_8331 ( R1171_U114 , R1171_U435 , R1171_U434 );
nand NAND2_8332 ( R1171_U115 , R1171_U442 , R1171_U441 );
nand NAND2_8333 ( R1171_U116 , R1171_U449 , R1171_U448 );
nand NAND2_8334 ( R1171_U117 , R1171_U456 , R1171_U455 );
nand NAND2_8335 ( R1171_U118 , R1171_U461 , R1171_U460 );
nand NAND2_8336 ( R1171_U119 , R1171_U468 , R1171_U467 );
nand NAND2_8337 ( R1171_U120 , R1171_U475 , R1171_U474 );
nand NAND2_8338 ( R1171_U121 , R1171_U489 , R1171_U488 );
nand NAND2_8339 ( R1171_U122 , R1171_U494 , R1171_U493 );
nand NAND2_8340 ( R1171_U123 , R1171_U501 , R1171_U500 );
nand NAND2_8341 ( R1171_U124 , R1171_U508 , R1171_U507 );
nand NAND2_8342 ( R1171_U125 , R1171_U515 , R1171_U514 );
nand NAND2_8343 ( R1171_U126 , R1171_U522 , R1171_U521 );
nand NAND2_8344 ( R1171_U127 , R1171_U527 , R1171_U526 );
and AND2_8345 ( R1171_U128 , R1171_U129 , R1171_U197 );
and AND2_8346 ( R1171_U129 , U3065 , U3470 );
and AND2_8347 ( R1171_U130 , U3472 , U3061 );
and AND2_8348 ( R1171_U131 , U3464 , U3074 );
and AND3_8349 ( R1171_U132 , R1171_U204 , R1171_U206 , R1171_U203 );
and AND3_8350 ( R1171_U133 , R1171_U373 , R1171_U207 , R1171_U374 );
and AND3_8351 ( R1171_U134 , R1171_U409 , R1171_U408 , R1171_U43 );
and AND2_8352 ( R1171_U135 , R1171_U225 , R1171_U6 );
and AND2_8353 ( R1171_U136 , R1171_U233 , R1171_U231 );
and AND3_8354 ( R1171_U137 , R1171_U416 , R1171_U415 , R1171_U34 );
and AND2_8355 ( R1171_U138 , R1171_U239 , R1171_U4 );
and AND2_8356 ( R1171_U139 , R1171_U247 , R1171_U198 );
and AND2_8357 ( R1171_U140 , R1171_U252 , R1171_U188 );
and AND2_8358 ( R1171_U141 , R1171_U6 , R1171_U12 );
and AND2_8359 ( R1171_U142 , R1171_U378 , R1171_U255 );
and AND2_8360 ( R1171_U143 , R1171_U270 , R1171_U15 );
and AND2_8361 ( R1171_U144 , R1171_U260 , R1171_U189 );
and AND2_8362 ( R1171_U145 , R1171_U296 , R1171_U16 );
and AND2_8363 ( R1171_U146 , R1171_U389 , R1171_U297 );
and AND2_8364 ( R1171_U147 , R1171_U309 , R1171_U185 );
and AND3_8365 ( R1171_U148 , R1171_U393 , R1171_U310 , R1171_U395 );
and AND2_8366 ( R1171_U149 , R1171_U17 , R1171_U185 );
and AND2_8367 ( R1171_U150 , R1171_U97 , R1171_U304 );
and AND3_8368 ( R1171_U151 , R1171_U451 , R1171_U450 , R1171_U190 );
and AND2_8369 ( R1171_U152 , R1171_U320 , R1171_U185 );
and AND2_8370 ( R1171_U153 , R1171_U176 , R1171_U288 );
and AND3_8371 ( R1171_U154 , R1171_U482 , R1171_U481 , R1171_U80 );
and AND2_8372 ( R1171_U155 , R1171_U333 , R1171_U10 );
and AND3_8373 ( R1171_U156 , R1171_U496 , R1171_U495 , R1171_U90 );
and AND2_8374 ( R1171_U157 , R1171_U342 , R1171_U9 );
and AND3_8375 ( R1171_U158 , R1171_U517 , R1171_U516 , R1171_U189 );
and AND2_8376 ( R1171_U159 , R1171_U351 , R1171_U8 );
and AND3_8377 ( R1171_U160 , R1171_U529 , R1171_U528 , R1171_U188 );
and AND2_8378 ( R1171_U161 , R1171_U358 , R1171_U7 );
nand NAND2_8379 ( R1171_U162 , R1171_U375 , R1171_U215 );
nand NAND2_8380 ( R1171_U163 , R1171_U230 , R1171_U242 );
not NOT1_8381 ( R1171_U164 , U3052 );
not NOT1_8382 ( R1171_U165 , U4040 );
and AND2_8383 ( R1171_U166 , R1171_U430 , R1171_U429 );
nand NAND3_8384 ( R1171_U167 , R1171_U312 , R1171_U186 , R1171_U372 );
and AND2_8385 ( R1171_U168 , R1171_U437 , R1171_U436 );
nand NAND2_8386 ( R1171_U169 , R1171_U148 , R1171_U394 );
and AND2_8387 ( R1171_U170 , R1171_U444 , R1171_U443 );
nand NAND2_8388 ( R1171_U171 , R1171_U150 , R1171_U307 );
nand NAND2_8389 ( R1171_U172 , R1171_U301 , R1171_U300 );
and AND2_8390 ( R1171_U173 , R1171_U463 , R1171_U462 );
and AND2_8391 ( R1171_U174 , R1171_U470 , R1171_U469 );
nand NAND2_8392 ( R1171_U175 , R1171_U386 , R1171_U384 );
and AND2_8393 ( R1171_U176 , R1171_U477 , R1171_U476 );
nand NAND2_8394 ( R1171_U177 , U3074 , U3464 );
nand NAND2_8395 ( R1171_U178 , R1171_U36 , R1171_U335 );
nand NAND2_8396 ( R1171_U179 , R1171_U376 , R1171_U279 );
and AND2_8397 ( R1171_U180 , R1171_U503 , R1171_U502 );
nand NAND2_8398 ( R1171_U181 , R1171_U77 , R1171_U379 );
and AND2_8399 ( R1171_U182 , R1171_U510 , R1171_U509 );
nand NAND2_8400 ( R1171_U183 , R1171_U265 , R1171_U264 );
nand NAND2_8401 ( R1171_U184 , R1171_U142 , R1171_U377 );
nand NAND2_8402 ( R1171_U185 , R1171_U391 , R1171_U390 );
nand NAND2_8403 ( R1171_U186 , U3051 , R1171_U169 );
not NOT1_8404 ( R1171_U187 , R1171_U34 );
nand NAND2_8405 ( R1171_U188 , U3484 , U3080 );
nand NAND2_8406 ( R1171_U189 , U3069 , U3490 );
nand NAND2_8407 ( R1171_U190 , U3055 , U4032 );
not NOT1_8408 ( R1171_U191 , R1171_U72 );
not NOT1_8409 ( R1171_U192 , R1171_U84 );
not NOT1_8410 ( R1171_U193 , R1171_U60 );
not NOT1_8411 ( R1171_U194 , R1171_U65 );
or OR2_8412 ( R1171_U195 , U3064 , U3476 );
or OR2_8413 ( R1171_U196 , U3057 , U3474 );
or OR2_8414 ( R1171_U197 , U3472 , U3061 );
or OR2_8415 ( R1171_U198 , U3470 , U3065 );
not NOT1_8416 ( R1171_U199 , R1171_U177 );
or OR2_8417 ( R1171_U200 , U3468 , U3075 );
not NOT1_8418 ( R1171_U201 , R1171_U39 );
not NOT1_8419 ( R1171_U202 , R1171_U36 );
nand NAND2_8420 ( R1171_U203 , R1171_U4 , R1171_U128 );
nand NAND2_8421 ( R1171_U204 , R1171_U130 , R1171_U4 );
nand NAND2_8422 ( R1171_U205 , R1171_U35 , R1171_U34 );
nand NAND2_8423 ( R1171_U206 , U3064 , R1171_U205 );
nand NAND2_8424 ( R1171_U207 , U3476 , R1171_U187 );
not NOT1_8425 ( R1171_U208 , R1171_U51 );
or OR2_8426 ( R1171_U209 , U3067 , U3480 );
or OR2_8427 ( R1171_U210 , U3068 , U3478 );
not NOT1_8428 ( R1171_U211 , R1171_U43 );
nand NAND2_8429 ( R1171_U212 , R1171_U44 , R1171_U43 );
nand NAND2_8430 ( R1171_U213 , U3067 , R1171_U212 );
nand NAND2_8431 ( R1171_U214 , U3480 , R1171_U211 );
nand NAND2_8432 ( R1171_U215 , R1171_U6 , R1171_U51 );
not NOT1_8433 ( R1171_U216 , R1171_U162 );
or OR2_8434 ( R1171_U217 , U3482 , U3081 );
nand NAND2_8435 ( R1171_U218 , R1171_U217 , R1171_U162 );
not NOT1_8436 ( R1171_U219 , R1171_U50 );
or OR2_8437 ( R1171_U220 , U3080 , U3484 );
or OR2_8438 ( R1171_U221 , U3478 , U3068 );
nand NAND2_8439 ( R1171_U222 , R1171_U221 , R1171_U51 );
nand NAND2_8440 ( R1171_U223 , R1171_U134 , R1171_U222 );
nand NAND2_8441 ( R1171_U224 , R1171_U208 , R1171_U43 );
nand NAND2_8442 ( R1171_U225 , U3480 , U3067 );
nand NAND2_8443 ( R1171_U226 , R1171_U135 , R1171_U224 );
or OR2_8444 ( R1171_U227 , U3068 , U3478 );
nand NAND2_8445 ( R1171_U228 , R1171_U202 , R1171_U198 );
nand NAND2_8446 ( R1171_U229 , U3065 , U3470 );
not NOT1_8447 ( R1171_U230 , R1171_U53 );
nand NAND2_8448 ( R1171_U231 , R1171_U201 , R1171_U5 );
nand NAND2_8449 ( R1171_U232 , R1171_U53 , R1171_U197 );
nand NAND2_8450 ( R1171_U233 , U3061 , U3472 );
not NOT1_8451 ( R1171_U234 , R1171_U52 );
or OR2_8452 ( R1171_U235 , U3474 , U3057 );
nand NAND2_8453 ( R1171_U236 , R1171_U235 , R1171_U52 );
nand NAND2_8454 ( R1171_U237 , R1171_U137 , R1171_U236 );
nand NAND2_8455 ( R1171_U238 , R1171_U234 , R1171_U34 );
nand NAND2_8456 ( R1171_U239 , U3476 , U3064 );
nand NAND2_8457 ( R1171_U240 , R1171_U138 , R1171_U238 );
or OR2_8458 ( R1171_U241 , U3057 , U3474 );
nand NAND2_8459 ( R1171_U242 , R1171_U201 , R1171_U198 );
not NOT1_8460 ( R1171_U243 , R1171_U163 );
nand NAND2_8461 ( R1171_U244 , U3061 , U3472 );
nand NAND4_8462 ( R1171_U245 , R1171_U428 , R1171_U427 , R1171_U36 , R1171_U39 );
nand NAND2_8463 ( R1171_U246 , R1171_U36 , R1171_U39 );
nand NAND2_8464 ( R1171_U247 , U3065 , U3470 );
nand NAND2_8465 ( R1171_U248 , R1171_U139 , R1171_U246 );
or OR2_8466 ( R1171_U249 , U3080 , U3484 );
or OR2_8467 ( R1171_U250 , U3059 , U3486 );
nand NAND2_8468 ( R1171_U251 , R1171_U194 , R1171_U7 );
nand NAND2_8469 ( R1171_U252 , U3059 , U3486 );
nand NAND2_8470 ( R1171_U253 , R1171_U140 , R1171_U251 );
or OR2_8471 ( R1171_U254 , U3486 , U3059 );
nand NAND2_8472 ( R1171_U255 , R1171_U254 , R1171_U253 );
not NOT1_8473 ( R1171_U256 , R1171_U184 );
or OR2_8474 ( R1171_U257 , U3077 , U3492 );
or OR2_8475 ( R1171_U258 , U3069 , U3490 );
nand NAND2_8476 ( R1171_U259 , R1171_U191 , R1171_U8 );
nand NAND2_8477 ( R1171_U260 , U3077 , U3492 );
nand NAND2_8478 ( R1171_U261 , R1171_U144 , R1171_U259 );
or OR2_8479 ( R1171_U262 , U3488 , U3060 );
or OR2_8480 ( R1171_U263 , U3492 , U3077 );
nand NAND2_8481 ( R1171_U264 , R1171_U13 , R1171_U184 );
nand NAND2_8482 ( R1171_U265 , R1171_U263 , R1171_U261 );
not NOT1_8483 ( R1171_U266 , R1171_U183 );
or OR2_8484 ( R1171_U267 , U3494 , U3076 );
nand NAND2_8485 ( R1171_U268 , U3076 , U3494 );
not NOT1_8486 ( R1171_U269 , R1171_U181 );
or OR2_8487 ( R1171_U270 , U3496 , U3071 );
nand NAND2_8488 ( R1171_U271 , U3071 , U3496 );
not NOT1_8489 ( R1171_U272 , R1171_U105 );
or OR2_8490 ( R1171_U273 , U3066 , U3500 );
or OR2_8491 ( R1171_U274 , U3070 , U3498 );
not NOT1_8492 ( R1171_U275 , R1171_U90 );
nand NAND2_8493 ( R1171_U276 , R1171_U91 , R1171_U90 );
nand NAND2_8494 ( R1171_U277 , U3066 , R1171_U276 );
nand NAND2_8495 ( R1171_U278 , U3500 , R1171_U275 );
nand NAND2_8496 ( R1171_U279 , R1171_U9 , R1171_U105 );
not NOT1_8497 ( R1171_U280 , R1171_U179 );
or OR2_8498 ( R1171_U281 , U3073 , U4037 );
or OR2_8499 ( R1171_U282 , U3078 , U3504 );
or OR2_8500 ( R1171_U283 , U3072 , U4036 );
not NOT1_8501 ( R1171_U284 , R1171_U80 );
nand NAND2_8502 ( R1171_U285 , U4037 , R1171_U284 );
nand NAND2_8503 ( R1171_U286 , R1171_U285 , R1171_U103 );
nand NAND2_8504 ( R1171_U287 , R1171_U80 , R1171_U81 );
nand NAND2_8505 ( R1171_U288 , R1171_U287 , R1171_U286 );
nand NAND2_8506 ( R1171_U289 , R1171_U192 , R1171_U11 );
nand NAND2_8507 ( R1171_U290 , U3072 , U4036 );
nand NAND3_8508 ( R1171_U291 , R1171_U289 , R1171_U288 , R1171_U290 );
or OR2_8509 ( R1171_U292 , U3502 , U3079 );
or OR2_8510 ( R1171_U293 , U4036 , U3072 );
nand NAND2_8511 ( R1171_U294 , R1171_U293 , R1171_U291 );
not NOT1_8512 ( R1171_U295 , R1171_U175 );
or OR2_8513 ( R1171_U296 , U4035 , U3058 );
nand NAND2_8514 ( R1171_U297 , U3058 , U4035 );
not NOT1_8515 ( R1171_U298 , R1171_U94 );
or OR2_8516 ( R1171_U299 , U4034 , U3063 );
nand NAND2_8517 ( R1171_U300 , R1171_U299 , R1171_U94 );
nand NAND2_8518 ( R1171_U301 , U3063 , U4034 );
not NOT1_8519 ( R1171_U302 , R1171_U172 );
or OR2_8520 ( R1171_U303 , U3055 , U4032 );
nand NAND2_8521 ( R1171_U304 , R1171_U193 , R1171_U185 );
or OR2_8522 ( R1171_U305 , U4033 , U3062 );
or OR2_8523 ( R1171_U306 , U4031 , U3054 );
nand NAND2_8524 ( R1171_U307 , R1171_U149 , R1171_U392 );
not NOT1_8525 ( R1171_U308 , R1171_U171 );
or OR2_8526 ( R1171_U309 , U4030 , U3050 );
nand NAND2_8527 ( R1171_U310 , U3050 , U4030 );
not NOT1_8528 ( R1171_U311 , R1171_U169 );
nand NAND2_8529 ( R1171_U312 , U4029 , R1171_U169 );
not NOT1_8530 ( R1171_U313 , R1171_U167 );
nand NAND2_8531 ( R1171_U314 , R1171_U305 , R1171_U172 );
not NOT1_8532 ( R1171_U315 , R1171_U100 );
or OR2_8533 ( R1171_U316 , U4032 , U3055 );
nand NAND2_8534 ( R1171_U317 , R1171_U316 , R1171_U100 );
nand NAND2_8535 ( R1171_U318 , R1171_U151 , R1171_U317 );
nand NAND2_8536 ( R1171_U319 , R1171_U315 , R1171_U190 );
nand NAND2_8537 ( R1171_U320 , U4031 , U3054 );
nand NAND2_8538 ( R1171_U321 , R1171_U152 , R1171_U319 );
or OR2_8539 ( R1171_U322 , U3055 , U4032 );
nand NAND2_8540 ( R1171_U323 , R1171_U292 , R1171_U179 );
not NOT1_8541 ( R1171_U324 , R1171_U104 );
nand NAND2_8542 ( R1171_U325 , R1171_U10 , R1171_U104 );
nand NAND2_8543 ( R1171_U326 , R1171_U153 , R1171_U325 );
nand NAND2_8544 ( R1171_U327 , R1171_U325 , R1171_U288 );
nand NAND2_8545 ( R1171_U328 , R1171_U480 , R1171_U327 );
or OR2_8546 ( R1171_U329 , U3504 , U3078 );
nand NAND2_8547 ( R1171_U330 , R1171_U329 , R1171_U104 );
nand NAND2_8548 ( R1171_U331 , R1171_U154 , R1171_U330 );
nand NAND2_8549 ( R1171_U332 , R1171_U324 , R1171_U80 );
nand NAND2_8550 ( R1171_U333 , U3073 , U4037 );
nand NAND2_8551 ( R1171_U334 , R1171_U155 , R1171_U332 );
or OR2_8552 ( R1171_U335 , U3468 , U3075 );
not NOT1_8553 ( R1171_U336 , R1171_U178 );
or OR2_8554 ( R1171_U337 , U3078 , U3504 );
or OR2_8555 ( R1171_U338 , U3498 , U3070 );
nand NAND2_8556 ( R1171_U339 , R1171_U338 , R1171_U105 );
nand NAND2_8557 ( R1171_U340 , R1171_U156 , R1171_U339 );
nand NAND2_8558 ( R1171_U341 , R1171_U272 , R1171_U90 );
nand NAND2_8559 ( R1171_U342 , U3500 , U3066 );
nand NAND2_8560 ( R1171_U343 , R1171_U157 , R1171_U341 );
or OR2_8561 ( R1171_U344 , U3070 , U3498 );
nand NAND2_8562 ( R1171_U345 , R1171_U262 , R1171_U184 );
not NOT1_8563 ( R1171_U346 , R1171_U106 );
or OR2_8564 ( R1171_U347 , U3490 , U3069 );
nand NAND2_8565 ( R1171_U348 , R1171_U347 , R1171_U106 );
nand NAND2_8566 ( R1171_U349 , R1171_U158 , R1171_U348 );
nand NAND2_8567 ( R1171_U350 , R1171_U346 , R1171_U189 );
nand NAND2_8568 ( R1171_U351 , U3077 , U3492 );
nand NAND2_8569 ( R1171_U352 , R1171_U159 , R1171_U350 );
or OR2_8570 ( R1171_U353 , U3069 , U3490 );
or OR2_8571 ( R1171_U354 , U3484 , U3080 );
nand NAND2_8572 ( R1171_U355 , R1171_U354 , R1171_U50 );
nand NAND2_8573 ( R1171_U356 , R1171_U160 , R1171_U355 );
nand NAND2_8574 ( R1171_U357 , R1171_U219 , R1171_U188 );
nand NAND2_8575 ( R1171_U358 , U3059 , U3486 );
nand NAND2_8576 ( R1171_U359 , R1171_U161 , R1171_U357 );
nand NAND2_8577 ( R1171_U360 , R1171_U220 , R1171_U188 );
nand NAND2_8578 ( R1171_U361 , R1171_U217 , R1171_U65 );
nand NAND2_8579 ( R1171_U362 , R1171_U227 , R1171_U43 );
nand NAND2_8580 ( R1171_U363 , R1171_U241 , R1171_U34 );
nand NAND2_8581 ( R1171_U364 , R1171_U244 , R1171_U197 );
nand NAND2_8582 ( R1171_U365 , R1171_U322 , R1171_U190 );
nand NAND2_8583 ( R1171_U366 , R1171_U305 , R1171_U60 );
nand NAND2_8584 ( R1171_U367 , R1171_U337 , R1171_U80 );
nand NAND2_8585 ( R1171_U368 , R1171_U292 , R1171_U84 );
nand NAND2_8586 ( R1171_U369 , R1171_U344 , R1171_U90 );
nand NAND2_8587 ( R1171_U370 , R1171_U353 , R1171_U189 );
nand NAND2_8588 ( R1171_U371 , R1171_U262 , R1171_U72 );
nand NAND2_8589 ( R1171_U372 , U4029 , U3051 );
nand NAND3_8590 ( R1171_U373 , R1171_U202 , R1171_U4 , R1171_U5 );
nand NAND3_8591 ( R1171_U374 , R1171_U5 , R1171_U4 , R1171_U201 );
not NOT1_8592 ( R1171_U375 , R1171_U45 );
not NOT1_8593 ( R1171_U376 , R1171_U102 );
nand NAND2_8594 ( R1171_U377 , R1171_U141 , R1171_U51 );
nand NAND2_8595 ( R1171_U378 , R1171_U12 , R1171_U45 );
nand NAND2_8596 ( R1171_U379 , R1171_U15 , R1171_U184 );
nand NAND2_8597 ( R1171_U380 , R1171_U268 , R1171_U265 );
not NOT1_8598 ( R1171_U381 , R1171_U77 );
nand NAND2_8599 ( R1171_U382 , R1171_U143 , R1171_U184 );
nand NAND2_8600 ( R1171_U383 , R1171_U381 , R1171_U270 );
nand NAND2_8601 ( R1171_U384 , R1171_U16 , R1171_U105 );
nand NAND2_8602 ( R1171_U385 , R1171_U14 , R1171_U102 );
not NOT1_8603 ( R1171_U386 , R1171_U101 );
not NOT1_8604 ( R1171_U387 , R1171_U97 );
nand NAND2_8605 ( R1171_U388 , R1171_U145 , R1171_U105 );
nand NAND2_8606 ( R1171_U389 , R1171_U101 , R1171_U296 );
nand NAND2_8607 ( R1171_U390 , U3054 , R1171_U303 );
nand NAND2_8608 ( R1171_U391 , U4031 , R1171_U303 );
nand NAND2_8609 ( R1171_U392 , R1171_U298 , R1171_U301 );
nand NAND3_8610 ( R1171_U393 , R1171_U193 , R1171_U185 , R1171_U309 );
nand NAND3_8611 ( R1171_U394 , R1171_U17 , R1171_U392 , R1171_U147 );
nand NAND2_8612 ( R1171_U395 , R1171_U387 , R1171_U309 );
nand NAND2_8613 ( R1171_U396 , R1171_U57 , R1171_U190 );
nand NAND2_8614 ( R1171_U397 , R1171_U56 , R1171_U190 );
nand NAND2_8615 ( R1171_U398 , U3080 , R1171_U49 );
nand NAND2_8616 ( R1171_U399 , U3484 , R1171_U48 );
nand NAND2_8617 ( R1171_U400 , R1171_U399 , R1171_U398 );
nand NAND2_8618 ( R1171_U401 , R1171_U360 , R1171_U50 );
nand NAND2_8619 ( R1171_U402 , R1171_U400 , R1171_U219 );
nand NAND2_8620 ( R1171_U403 , U3081 , R1171_U46 );
nand NAND2_8621 ( R1171_U404 , U3482 , R1171_U47 );
nand NAND2_8622 ( R1171_U405 , R1171_U404 , R1171_U403 );
nand NAND2_8623 ( R1171_U406 , R1171_U361 , R1171_U162 );
nand NAND2_8624 ( R1171_U407 , R1171_U216 , R1171_U405 );
nand NAND2_8625 ( R1171_U408 , U3067 , R1171_U44 );
nand NAND2_8626 ( R1171_U409 , U3480 , R1171_U42 );
nand NAND2_8627 ( R1171_U410 , U3068 , R1171_U40 );
nand NAND2_8628 ( R1171_U411 , U3478 , R1171_U41 );
nand NAND2_8629 ( R1171_U412 , R1171_U411 , R1171_U410 );
nand NAND2_8630 ( R1171_U413 , R1171_U362 , R1171_U51 );
nand NAND2_8631 ( R1171_U414 , R1171_U412 , R1171_U208 );
nand NAND2_8632 ( R1171_U415 , U3064 , R1171_U35 );
nand NAND2_8633 ( R1171_U416 , U3476 , R1171_U33 );
nand NAND2_8634 ( R1171_U417 , U3057 , R1171_U31 );
nand NAND2_8635 ( R1171_U418 , U3474 , R1171_U32 );
nand NAND2_8636 ( R1171_U419 , R1171_U418 , R1171_U417 );
nand NAND2_8637 ( R1171_U420 , R1171_U363 , R1171_U52 );
nand NAND2_8638 ( R1171_U421 , R1171_U419 , R1171_U234 );
nand NAND2_8639 ( R1171_U422 , U3061 , R1171_U29 );
nand NAND2_8640 ( R1171_U423 , U3472 , R1171_U30 );
nand NAND2_8641 ( R1171_U424 , R1171_U423 , R1171_U422 );
nand NAND2_8642 ( R1171_U425 , R1171_U364 , R1171_U163 );
nand NAND2_8643 ( R1171_U426 , R1171_U243 , R1171_U424 );
nand NAND2_8644 ( R1171_U427 , U3065 , R1171_U27 );
nand NAND2_8645 ( R1171_U428 , U3470 , R1171_U28 );
nand NAND2_8646 ( R1171_U429 , U3052 , R1171_U165 );
nand NAND2_8647 ( R1171_U430 , U4040 , R1171_U164 );
nand NAND2_8648 ( R1171_U431 , U3052 , R1171_U165 );
nand NAND2_8649 ( R1171_U432 , U4040 , R1171_U164 );
nand NAND2_8650 ( R1171_U433 , R1171_U432 , R1171_U431 );
nand NAND2_8651 ( R1171_U434 , R1171_U166 , R1171_U167 );
nand NAND2_8652 ( R1171_U435 , R1171_U313 , R1171_U433 );
nand NAND2_8653 ( R1171_U436 , U3051 , R1171_U99 );
nand NAND2_8654 ( R1171_U437 , U4029 , R1171_U98 );
nand NAND2_8655 ( R1171_U438 , U3051 , R1171_U99 );
nand NAND2_8656 ( R1171_U439 , U4029 , R1171_U98 );
nand NAND2_8657 ( R1171_U440 , R1171_U439 , R1171_U438 );
nand NAND2_8658 ( R1171_U441 , R1171_U168 , R1171_U169 );
nand NAND2_8659 ( R1171_U442 , R1171_U311 , R1171_U440 );
nand NAND2_8660 ( R1171_U443 , U3050 , R1171_U54 );
nand NAND2_8661 ( R1171_U444 , U4030 , R1171_U55 );
nand NAND2_8662 ( R1171_U445 , U3050 , R1171_U54 );
nand NAND2_8663 ( R1171_U446 , U4030 , R1171_U55 );
nand NAND2_8664 ( R1171_U447 , R1171_U446 , R1171_U445 );
nand NAND2_8665 ( R1171_U448 , R1171_U170 , R1171_U171 );
nand NAND2_8666 ( R1171_U449 , R1171_U308 , R1171_U447 );
nand NAND2_8667 ( R1171_U450 , U3054 , R1171_U57 );
nand NAND2_8668 ( R1171_U451 , U4031 , R1171_U56 );
nand NAND2_8669 ( R1171_U452 , U3055 , R1171_U95 );
nand NAND2_8670 ( R1171_U453 , U4032 , R1171_U96 );
nand NAND2_8671 ( R1171_U454 , R1171_U453 , R1171_U452 );
nand NAND2_8672 ( R1171_U455 , R1171_U365 , R1171_U100 );
nand NAND2_8673 ( R1171_U456 , R1171_U454 , R1171_U315 );
nand NAND2_8674 ( R1171_U457 , U3062 , R1171_U58 );
nand NAND2_8675 ( R1171_U458 , U4033 , R1171_U59 );
nand NAND2_8676 ( R1171_U459 , R1171_U458 , R1171_U457 );
nand NAND2_8677 ( R1171_U460 , R1171_U366 , R1171_U172 );
nand NAND2_8678 ( R1171_U461 , R1171_U302 , R1171_U459 );
nand NAND2_8679 ( R1171_U462 , U3063 , R1171_U92 );
nand NAND2_8680 ( R1171_U463 , U4034 , R1171_U93 );
nand NAND2_8681 ( R1171_U464 , U3063 , R1171_U92 );
nand NAND2_8682 ( R1171_U465 , U4034 , R1171_U93 );
nand NAND2_8683 ( R1171_U466 , R1171_U465 , R1171_U464 );
nand NAND2_8684 ( R1171_U467 , R1171_U173 , R1171_U94 );
nand NAND2_8685 ( R1171_U468 , R1171_U466 , R1171_U298 );
nand NAND2_8686 ( R1171_U469 , U3058 , R1171_U61 );
nand NAND2_8687 ( R1171_U470 , U4035 , R1171_U62 );
nand NAND2_8688 ( R1171_U471 , U3058 , R1171_U61 );
nand NAND2_8689 ( R1171_U472 , U4035 , R1171_U62 );
nand NAND2_8690 ( R1171_U473 , R1171_U472 , R1171_U471 );
nand NAND2_8691 ( R1171_U474 , R1171_U174 , R1171_U175 );
nand NAND2_8692 ( R1171_U475 , R1171_U295 , R1171_U473 );
nand NAND2_8693 ( R1171_U476 , U3072 , R1171_U85 );
nand NAND2_8694 ( R1171_U477 , U4036 , R1171_U86 );
nand NAND2_8695 ( R1171_U478 , U3072 , R1171_U85 );
nand NAND2_8696 ( R1171_U479 , U4036 , R1171_U86 );
nand NAND2_8697 ( R1171_U480 , R1171_U479 , R1171_U478 );
nand NAND2_8698 ( R1171_U481 , U3073 , R1171_U81 );
nand NAND2_8699 ( R1171_U482 , U4037 , R1171_U103 );
nand NAND2_8700 ( R1171_U483 , R1171_U199 , R1171_U178 );
nand NAND2_8701 ( R1171_U484 , R1171_U336 , R1171_U177 );
nand NAND2_8702 ( R1171_U485 , U3078 , R1171_U78 );
nand NAND2_8703 ( R1171_U486 , U3504 , R1171_U79 );
nand NAND2_8704 ( R1171_U487 , R1171_U486 , R1171_U485 );
nand NAND2_8705 ( R1171_U488 , R1171_U367 , R1171_U104 );
nand NAND2_8706 ( R1171_U489 , R1171_U487 , R1171_U324 );
nand NAND2_8707 ( R1171_U490 , U3079 , R1171_U82 );
nand NAND2_8708 ( R1171_U491 , U3502 , R1171_U83 );
nand NAND2_8709 ( R1171_U492 , R1171_U491 , R1171_U490 );
nand NAND2_8710 ( R1171_U493 , R1171_U368 , R1171_U179 );
nand NAND2_8711 ( R1171_U494 , R1171_U280 , R1171_U492 );
nand NAND2_8712 ( R1171_U495 , U3066 , R1171_U91 );
nand NAND2_8713 ( R1171_U496 , U3500 , R1171_U89 );
nand NAND2_8714 ( R1171_U497 , U3070 , R1171_U87 );
nand NAND2_8715 ( R1171_U498 , U3498 , R1171_U88 );
nand NAND2_8716 ( R1171_U499 , R1171_U498 , R1171_U497 );
nand NAND2_8717 ( R1171_U500 , R1171_U369 , R1171_U105 );
nand NAND2_8718 ( R1171_U501 , R1171_U499 , R1171_U272 );
nand NAND2_8719 ( R1171_U502 , U3071 , R1171_U63 );
nand NAND2_8720 ( R1171_U503 , U3496 , R1171_U64 );
nand NAND2_8721 ( R1171_U504 , U3071 , R1171_U63 );
nand NAND2_8722 ( R1171_U505 , U3496 , R1171_U64 );
nand NAND2_8723 ( R1171_U506 , R1171_U505 , R1171_U504 );
nand NAND2_8724 ( R1171_U507 , R1171_U180 , R1171_U181 );
nand NAND2_8725 ( R1171_U508 , R1171_U269 , R1171_U506 );
nand NAND2_8726 ( R1171_U509 , U3076 , R1171_U75 );
nand NAND2_8727 ( R1171_U510 , U3494 , R1171_U76 );
nand NAND2_8728 ( R1171_U511 , U3076 , R1171_U75 );
nand NAND2_8729 ( R1171_U512 , U3494 , R1171_U76 );
nand NAND2_8730 ( R1171_U513 , R1171_U512 , R1171_U511 );
nand NAND2_8731 ( R1171_U514 , R1171_U182 , R1171_U183 );
nand NAND2_8732 ( R1171_U515 , R1171_U266 , R1171_U513 );
nand NAND2_8733 ( R1171_U516 , U3077 , R1171_U73 );
nand NAND2_8734 ( R1171_U517 , U3492 , R1171_U74 );
nand NAND2_8735 ( R1171_U518 , U3069 , R1171_U68 );
nand NAND2_8736 ( R1171_U519 , U3490 , R1171_U69 );
nand NAND2_8737 ( R1171_U520 , R1171_U519 , R1171_U518 );
nand NAND2_8738 ( R1171_U521 , R1171_U370 , R1171_U106 );
nand NAND2_8739 ( R1171_U522 , R1171_U520 , R1171_U346 );
nand NAND2_8740 ( R1171_U523 , U3060 , R1171_U70 );
nand NAND2_8741 ( R1171_U524 , U3488 , R1171_U71 );
nand NAND2_8742 ( R1171_U525 , R1171_U524 , R1171_U523 );
nand NAND2_8743 ( R1171_U526 , R1171_U371 , R1171_U184 );
nand NAND2_8744 ( R1171_U527 , R1171_U256 , R1171_U525 );
nand NAND2_8745 ( R1171_U528 , U3059 , R1171_U66 );
nand NAND2_8746 ( R1171_U529 , U3486 , R1171_U67 );
nand NAND2_8747 ( R1171_U530 , U3074 , R1171_U37 );
nand NAND2_8748 ( R1171_U531 , U3464 , R1171_U38 );
and AND2_8749 ( R1138_U4 , R1138_U196 , R1138_U195 );
and AND2_8750 ( R1138_U5 , R1138_U197 , R1138_U198 );
and AND2_8751 ( R1138_U6 , R1138_U210 , R1138_U209 );
and AND2_8752 ( R1138_U7 , R1138_U250 , R1138_U249 );
and AND2_8753 ( R1138_U8 , R1138_U258 , R1138_U257 );
and AND2_8754 ( R1138_U9 , R1138_U274 , R1138_U273 );
and AND2_8755 ( R1138_U10 , R1138_U282 , R1138_U281 );
and AND2_8756 ( R1138_U11 , R1138_U10 , R1138_U283 );
and AND2_8757 ( R1138_U12 , R1138_U7 , R1138_U217 );
and AND2_8758 ( R1138_U13 , R1138_U8 , R1138_U262 );
and AND2_8759 ( R1138_U14 , R1138_U11 , R1138_U292 );
and AND2_8760 ( R1138_U15 , R1138_U13 , R1138_U267 );
and AND2_8761 ( R1138_U16 , R1138_U9 , R1138_U14 );
and AND2_8762 ( R1138_U17 , R1138_U299 , R1138_U305 );
and AND2_8763 ( R1138_U18 , R1138_U359 , R1138_U356 );
and AND2_8764 ( R1138_U19 , R1138_U352 , R1138_U349 );
and AND2_8765 ( R1138_U20 , R1138_U343 , R1138_U340 );
and AND2_8766 ( R1138_U21 , R1138_U334 , R1138_U331 );
and AND2_8767 ( R1138_U22 , R1138_U328 , R1138_U326 );
and AND2_8768 ( R1138_U23 , R1138_U321 , R1138_U318 );
and AND2_8769 ( R1138_U24 , R1138_U248 , R1138_U245 );
and AND2_8770 ( R1138_U25 , R1138_U240 , R1138_U237 );
and AND2_8771 ( R1138_U26 , R1138_U226 , R1138_U223 );
not NOT1_8772 ( R1138_U27 , U3470 );
not NOT1_8773 ( R1138_U28 , U3065 );
not NOT1_8774 ( R1138_U29 , U3472 );
not NOT1_8775 ( R1138_U30 , U3061 );
not NOT1_8776 ( R1138_U31 , U3474 );
not NOT1_8777 ( R1138_U32 , U3057 );
not NOT1_8778 ( R1138_U33 , U3064 );
nand NAND2_8779 ( R1138_U34 , U3057 , U3474 );
not NOT1_8780 ( R1138_U35 , U3476 );
nand NAND2_8781 ( R1138_U36 , U3468 , U3075 );
not NOT1_8782 ( R1138_U37 , U3464 );
not NOT1_8783 ( R1138_U38 , U3074 );
nand NAND2_8784 ( R1138_U39 , R1138_U131 , R1138_U200 );
not NOT1_8785 ( R1138_U40 , U3478 );
not NOT1_8786 ( R1138_U41 , U3068 );
not NOT1_8787 ( R1138_U42 , U3067 );
nand NAND2_8788 ( R1138_U43 , U3068 , U3478 );
not NOT1_8789 ( R1138_U44 , U3480 );
nand NAND2_8790 ( R1138_U45 , R1138_U214 , R1138_U213 );
not NOT1_8791 ( R1138_U46 , U3482 );
not NOT1_8792 ( R1138_U47 , U3081 );
not NOT1_8793 ( R1138_U48 , U3080 );
not NOT1_8794 ( R1138_U49 , U3484 );
nand NAND2_8795 ( R1138_U50 , R1138_U65 , R1138_U218 );
nand NAND2_8796 ( R1138_U51 , R1138_U133 , R1138_U132 );
nand NAND2_8797 ( R1138_U52 , R1138_U136 , R1138_U232 );
nand NAND2_8798 ( R1138_U53 , R1138_U229 , R1138_U228 );
not NOT1_8799 ( R1138_U54 , U4030 );
not NOT1_8800 ( R1138_U55 , U3050 );
not NOT1_8801 ( R1138_U56 , U3054 );
not NOT1_8802 ( R1138_U57 , U4031 );
not NOT1_8803 ( R1138_U58 , U4033 );
not NOT1_8804 ( R1138_U59 , U3062 );
nand NAND2_8805 ( R1138_U60 , U3062 , U4033 );
not NOT1_8806 ( R1138_U61 , U4035 );
not NOT1_8807 ( R1138_U62 , U3058 );
not NOT1_8808 ( R1138_U63 , U3496 );
not NOT1_8809 ( R1138_U64 , U3071 );
nand NAND2_8810 ( R1138_U65 , U3081 , U3482 );
not NOT1_8811 ( R1138_U66 , U3486 );
not NOT1_8812 ( R1138_U67 , U3059 );
not NOT1_8813 ( R1138_U68 , U3490 );
not NOT1_8814 ( R1138_U69 , U3069 );
not NOT1_8815 ( R1138_U70 , U3488 );
not NOT1_8816 ( R1138_U71 , U3060 );
nand NAND2_8817 ( R1138_U72 , U3060 , U3488 );
not NOT1_8818 ( R1138_U73 , U3492 );
not NOT1_8819 ( R1138_U74 , U3077 );
not NOT1_8820 ( R1138_U75 , U3494 );
not NOT1_8821 ( R1138_U76 , U3076 );
nand NAND2_8822 ( R1138_U77 , R1138_U380 , R1138_U267 );
not NOT1_8823 ( R1138_U78 , U3504 );
not NOT1_8824 ( R1138_U79 , U3078 );
nand NAND2_8825 ( R1138_U80 , U3078 , U3504 );
not NOT1_8826 ( R1138_U81 , U4037 );
not NOT1_8827 ( R1138_U82 , U3502 );
not NOT1_8828 ( R1138_U83 , U3079 );
nand NAND2_8829 ( R1138_U84 , U3079 , U3502 );
not NOT1_8830 ( R1138_U85 , U4036 );
not NOT1_8831 ( R1138_U86 , U3072 );
not NOT1_8832 ( R1138_U87 , U3498 );
not NOT1_8833 ( R1138_U88 , U3070 );
not NOT1_8834 ( R1138_U89 , U3066 );
nand NAND2_8835 ( R1138_U90 , U3070 , U3498 );
not NOT1_8836 ( R1138_U91 , U3500 );
not NOT1_8837 ( R1138_U92 , U4034 );
not NOT1_8838 ( R1138_U93 , U3063 );
nand NAND2_8839 ( R1138_U94 , R1138_U146 , R1138_U388 );
not NOT1_8840 ( R1138_U95 , U4032 );
not NOT1_8841 ( R1138_U96 , U3055 );
nand NAND3_8842 ( R1138_U97 , R1138_U396 , R1138_U306 , R1138_U397 );
not NOT1_8843 ( R1138_U98 , U3051 );
not NOT1_8844 ( R1138_U99 , U4029 );
nand NAND2_8845 ( R1138_U100 , R1138_U60 , R1138_U314 );
nand NAND2_8846 ( R1138_U101 , R1138_U385 , R1138_U294 );
nand NAND2_8847 ( R1138_U102 , R1138_U278 , R1138_U277 );
not NOT1_8848 ( R1138_U103 , U3073 );
nand NAND2_8849 ( R1138_U104 , R1138_U84 , R1138_U323 );
nand NAND3_8850 ( R1138_U105 , R1138_U383 , R1138_U271 , R1138_U382 );
nand NAND2_8851 ( R1138_U106 , R1138_U72 , R1138_U345 );
nand NAND2_8852 ( R1138_U107 , R1138_U484 , R1138_U483 );
nand NAND2_8853 ( R1138_U108 , R1138_U531 , R1138_U530 );
nand NAND2_8854 ( R1138_U109 , R1138_U402 , R1138_U401 );
nand NAND2_8855 ( R1138_U110 , R1138_U407 , R1138_U406 );
nand NAND2_8856 ( R1138_U111 , R1138_U414 , R1138_U413 );
nand NAND2_8857 ( R1138_U112 , R1138_U421 , R1138_U420 );
nand NAND2_8858 ( R1138_U113 , R1138_U426 , R1138_U425 );
nand NAND2_8859 ( R1138_U114 , R1138_U435 , R1138_U434 );
nand NAND2_8860 ( R1138_U115 , R1138_U442 , R1138_U441 );
nand NAND2_8861 ( R1138_U116 , R1138_U449 , R1138_U448 );
nand NAND2_8862 ( R1138_U117 , R1138_U456 , R1138_U455 );
nand NAND2_8863 ( R1138_U118 , R1138_U461 , R1138_U460 );
nand NAND2_8864 ( R1138_U119 , R1138_U468 , R1138_U467 );
nand NAND2_8865 ( R1138_U120 , R1138_U475 , R1138_U474 );
nand NAND2_8866 ( R1138_U121 , R1138_U489 , R1138_U488 );
nand NAND2_8867 ( R1138_U122 , R1138_U494 , R1138_U493 );
nand NAND2_8868 ( R1138_U123 , R1138_U501 , R1138_U500 );
nand NAND2_8869 ( R1138_U124 , R1138_U508 , R1138_U507 );
nand NAND2_8870 ( R1138_U125 , R1138_U515 , R1138_U514 );
nand NAND2_8871 ( R1138_U126 , R1138_U522 , R1138_U521 );
nand NAND2_8872 ( R1138_U127 , R1138_U527 , R1138_U526 );
and AND2_8873 ( R1138_U128 , R1138_U129 , R1138_U197 );
and AND2_8874 ( R1138_U129 , U3065 , U3470 );
and AND2_8875 ( R1138_U130 , U3472 , U3061 );
and AND2_8876 ( R1138_U131 , U3464 , U3074 );
and AND3_8877 ( R1138_U132 , R1138_U204 , R1138_U206 , R1138_U203 );
and AND3_8878 ( R1138_U133 , R1138_U373 , R1138_U207 , R1138_U374 );
and AND3_8879 ( R1138_U134 , R1138_U409 , R1138_U408 , R1138_U43 );
and AND2_8880 ( R1138_U135 , R1138_U225 , R1138_U6 );
and AND2_8881 ( R1138_U136 , R1138_U233 , R1138_U231 );
and AND3_8882 ( R1138_U137 , R1138_U416 , R1138_U415 , R1138_U34 );
and AND2_8883 ( R1138_U138 , R1138_U239 , R1138_U4 );
and AND2_8884 ( R1138_U139 , R1138_U247 , R1138_U198 );
and AND2_8885 ( R1138_U140 , R1138_U252 , R1138_U188 );
and AND2_8886 ( R1138_U141 , R1138_U6 , R1138_U12 );
and AND2_8887 ( R1138_U142 , R1138_U378 , R1138_U255 );
and AND2_8888 ( R1138_U143 , R1138_U270 , R1138_U15 );
and AND2_8889 ( R1138_U144 , R1138_U260 , R1138_U189 );
and AND2_8890 ( R1138_U145 , R1138_U296 , R1138_U16 );
and AND2_8891 ( R1138_U146 , R1138_U389 , R1138_U297 );
and AND2_8892 ( R1138_U147 , R1138_U309 , R1138_U185 );
and AND3_8893 ( R1138_U148 , R1138_U393 , R1138_U310 , R1138_U395 );
and AND2_8894 ( R1138_U149 , R1138_U17 , R1138_U185 );
and AND2_8895 ( R1138_U150 , R1138_U97 , R1138_U304 );
and AND3_8896 ( R1138_U151 , R1138_U451 , R1138_U450 , R1138_U190 );
and AND2_8897 ( R1138_U152 , R1138_U320 , R1138_U185 );
and AND2_8898 ( R1138_U153 , R1138_U176 , R1138_U288 );
and AND3_8899 ( R1138_U154 , R1138_U482 , R1138_U481 , R1138_U80 );
and AND2_8900 ( R1138_U155 , R1138_U333 , R1138_U10 );
and AND3_8901 ( R1138_U156 , R1138_U496 , R1138_U495 , R1138_U90 );
and AND2_8902 ( R1138_U157 , R1138_U342 , R1138_U9 );
and AND3_8903 ( R1138_U158 , R1138_U517 , R1138_U516 , R1138_U189 );
and AND2_8904 ( R1138_U159 , R1138_U351 , R1138_U8 );
and AND3_8905 ( R1138_U160 , R1138_U529 , R1138_U528 , R1138_U188 );
and AND2_8906 ( R1138_U161 , R1138_U358 , R1138_U7 );
nand NAND2_8907 ( R1138_U162 , R1138_U375 , R1138_U215 );
nand NAND2_8908 ( R1138_U163 , R1138_U230 , R1138_U242 );
not NOT1_8909 ( R1138_U164 , U3052 );
not NOT1_8910 ( R1138_U165 , U4040 );
and AND2_8911 ( R1138_U166 , R1138_U430 , R1138_U429 );
nand NAND3_8912 ( R1138_U167 , R1138_U312 , R1138_U186 , R1138_U372 );
and AND2_8913 ( R1138_U168 , R1138_U437 , R1138_U436 );
nand NAND2_8914 ( R1138_U169 , R1138_U148 , R1138_U394 );
and AND2_8915 ( R1138_U170 , R1138_U444 , R1138_U443 );
nand NAND2_8916 ( R1138_U171 , R1138_U150 , R1138_U307 );
nand NAND2_8917 ( R1138_U172 , R1138_U301 , R1138_U300 );
and AND2_8918 ( R1138_U173 , R1138_U463 , R1138_U462 );
and AND2_8919 ( R1138_U174 , R1138_U470 , R1138_U469 );
nand NAND2_8920 ( R1138_U175 , R1138_U386 , R1138_U384 );
and AND2_8921 ( R1138_U176 , R1138_U477 , R1138_U476 );
nand NAND2_8922 ( R1138_U177 , U3074 , U3464 );
nand NAND2_8923 ( R1138_U178 , R1138_U36 , R1138_U335 );
nand NAND2_8924 ( R1138_U179 , R1138_U376 , R1138_U279 );
and AND2_8925 ( R1138_U180 , R1138_U503 , R1138_U502 );
nand NAND2_8926 ( R1138_U181 , R1138_U77 , R1138_U379 );
and AND2_8927 ( R1138_U182 , R1138_U510 , R1138_U509 );
nand NAND2_8928 ( R1138_U183 , R1138_U265 , R1138_U264 );
nand NAND2_8929 ( R1138_U184 , R1138_U142 , R1138_U377 );
nand NAND2_8930 ( R1138_U185 , R1138_U391 , R1138_U390 );
nand NAND2_8931 ( R1138_U186 , U3051 , R1138_U169 );
not NOT1_8932 ( R1138_U187 , R1138_U34 );
nand NAND2_8933 ( R1138_U188 , U3484 , U3080 );
nand NAND2_8934 ( R1138_U189 , U3069 , U3490 );
nand NAND2_8935 ( R1138_U190 , U3055 , U4032 );
not NOT1_8936 ( R1138_U191 , R1138_U72 );
not NOT1_8937 ( R1138_U192 , R1138_U84 );
not NOT1_8938 ( R1138_U193 , R1138_U60 );
not NOT1_8939 ( R1138_U194 , R1138_U65 );
or OR2_8940 ( R1138_U195 , U3064 , U3476 );
or OR2_8941 ( R1138_U196 , U3057 , U3474 );
or OR2_8942 ( R1138_U197 , U3472 , U3061 );
or OR2_8943 ( R1138_U198 , U3470 , U3065 );
not NOT1_8944 ( R1138_U199 , R1138_U177 );
or OR2_8945 ( R1138_U200 , U3468 , U3075 );
not NOT1_8946 ( R1138_U201 , R1138_U39 );
not NOT1_8947 ( R1138_U202 , R1138_U36 );
nand NAND2_8948 ( R1138_U203 , R1138_U4 , R1138_U128 );
nand NAND2_8949 ( R1138_U204 , R1138_U130 , R1138_U4 );
nand NAND2_8950 ( R1138_U205 , R1138_U35 , R1138_U34 );
nand NAND2_8951 ( R1138_U206 , U3064 , R1138_U205 );
nand NAND2_8952 ( R1138_U207 , U3476 , R1138_U187 );
not NOT1_8953 ( R1138_U208 , R1138_U51 );
or OR2_8954 ( R1138_U209 , U3067 , U3480 );
or OR2_8955 ( R1138_U210 , U3068 , U3478 );
not NOT1_8956 ( R1138_U211 , R1138_U43 );
nand NAND2_8957 ( R1138_U212 , R1138_U44 , R1138_U43 );
nand NAND2_8958 ( R1138_U213 , U3067 , R1138_U212 );
nand NAND2_8959 ( R1138_U214 , U3480 , R1138_U211 );
nand NAND2_8960 ( R1138_U215 , R1138_U6 , R1138_U51 );
not NOT1_8961 ( R1138_U216 , R1138_U162 );
or OR2_8962 ( R1138_U217 , U3482 , U3081 );
nand NAND2_8963 ( R1138_U218 , R1138_U217 , R1138_U162 );
not NOT1_8964 ( R1138_U219 , R1138_U50 );
or OR2_8965 ( R1138_U220 , U3080 , U3484 );
or OR2_8966 ( R1138_U221 , U3478 , U3068 );
nand NAND2_8967 ( R1138_U222 , R1138_U221 , R1138_U51 );
nand NAND2_8968 ( R1138_U223 , R1138_U134 , R1138_U222 );
nand NAND2_8969 ( R1138_U224 , R1138_U208 , R1138_U43 );
nand NAND2_8970 ( R1138_U225 , U3480 , U3067 );
nand NAND2_8971 ( R1138_U226 , R1138_U135 , R1138_U224 );
or OR2_8972 ( R1138_U227 , U3068 , U3478 );
nand NAND2_8973 ( R1138_U228 , R1138_U202 , R1138_U198 );
nand NAND2_8974 ( R1138_U229 , U3065 , U3470 );
not NOT1_8975 ( R1138_U230 , R1138_U53 );
nand NAND2_8976 ( R1138_U231 , R1138_U201 , R1138_U5 );
nand NAND2_8977 ( R1138_U232 , R1138_U53 , R1138_U197 );
nand NAND2_8978 ( R1138_U233 , U3061 , U3472 );
not NOT1_8979 ( R1138_U234 , R1138_U52 );
or OR2_8980 ( R1138_U235 , U3474 , U3057 );
nand NAND2_8981 ( R1138_U236 , R1138_U235 , R1138_U52 );
nand NAND2_8982 ( R1138_U237 , R1138_U137 , R1138_U236 );
nand NAND2_8983 ( R1138_U238 , R1138_U234 , R1138_U34 );
nand NAND2_8984 ( R1138_U239 , U3476 , U3064 );
nand NAND2_8985 ( R1138_U240 , R1138_U138 , R1138_U238 );
or OR2_8986 ( R1138_U241 , U3057 , U3474 );
nand NAND2_8987 ( R1138_U242 , R1138_U201 , R1138_U198 );
not NOT1_8988 ( R1138_U243 , R1138_U163 );
nand NAND2_8989 ( R1138_U244 , U3061 , U3472 );
nand NAND4_8990 ( R1138_U245 , R1138_U428 , R1138_U427 , R1138_U36 , R1138_U39 );
nand NAND2_8991 ( R1138_U246 , R1138_U36 , R1138_U39 );
nand NAND2_8992 ( R1138_U247 , U3065 , U3470 );
nand NAND2_8993 ( R1138_U248 , R1138_U139 , R1138_U246 );
or OR2_8994 ( R1138_U249 , U3080 , U3484 );
or OR2_8995 ( R1138_U250 , U3059 , U3486 );
nand NAND2_8996 ( R1138_U251 , R1138_U194 , R1138_U7 );
nand NAND2_8997 ( R1138_U252 , U3059 , U3486 );
nand NAND2_8998 ( R1138_U253 , R1138_U140 , R1138_U251 );
or OR2_8999 ( R1138_U254 , U3486 , U3059 );
nand NAND2_9000 ( R1138_U255 , R1138_U254 , R1138_U253 );
not NOT1_9001 ( R1138_U256 , R1138_U184 );
or OR2_9002 ( R1138_U257 , U3077 , U3492 );
or OR2_9003 ( R1138_U258 , U3069 , U3490 );
nand NAND2_9004 ( R1138_U259 , R1138_U191 , R1138_U8 );
nand NAND2_9005 ( R1138_U260 , U3077 , U3492 );
nand NAND2_9006 ( R1138_U261 , R1138_U144 , R1138_U259 );
or OR2_9007 ( R1138_U262 , U3488 , U3060 );
or OR2_9008 ( R1138_U263 , U3492 , U3077 );
nand NAND2_9009 ( R1138_U264 , R1138_U13 , R1138_U184 );
nand NAND2_9010 ( R1138_U265 , R1138_U263 , R1138_U261 );
not NOT1_9011 ( R1138_U266 , R1138_U183 );
or OR2_9012 ( R1138_U267 , U3494 , U3076 );
nand NAND2_9013 ( R1138_U268 , U3076 , U3494 );
not NOT1_9014 ( R1138_U269 , R1138_U181 );
or OR2_9015 ( R1138_U270 , U3496 , U3071 );
nand NAND2_9016 ( R1138_U271 , U3071 , U3496 );
not NOT1_9017 ( R1138_U272 , R1138_U105 );
or OR2_9018 ( R1138_U273 , U3066 , U3500 );
or OR2_9019 ( R1138_U274 , U3070 , U3498 );
not NOT1_9020 ( R1138_U275 , R1138_U90 );
nand NAND2_9021 ( R1138_U276 , R1138_U91 , R1138_U90 );
nand NAND2_9022 ( R1138_U277 , U3066 , R1138_U276 );
nand NAND2_9023 ( R1138_U278 , U3500 , R1138_U275 );
nand NAND2_9024 ( R1138_U279 , R1138_U9 , R1138_U105 );
not NOT1_9025 ( R1138_U280 , R1138_U179 );
or OR2_9026 ( R1138_U281 , U3073 , U4037 );
or OR2_9027 ( R1138_U282 , U3078 , U3504 );
or OR2_9028 ( R1138_U283 , U3072 , U4036 );
not NOT1_9029 ( R1138_U284 , R1138_U80 );
nand NAND2_9030 ( R1138_U285 , U4037 , R1138_U284 );
nand NAND2_9031 ( R1138_U286 , R1138_U285 , R1138_U103 );
nand NAND2_9032 ( R1138_U287 , R1138_U80 , R1138_U81 );
nand NAND2_9033 ( R1138_U288 , R1138_U287 , R1138_U286 );
nand NAND2_9034 ( R1138_U289 , R1138_U192 , R1138_U11 );
nand NAND2_9035 ( R1138_U290 , U3072 , U4036 );
nand NAND3_9036 ( R1138_U291 , R1138_U289 , R1138_U288 , R1138_U290 );
or OR2_9037 ( R1138_U292 , U3502 , U3079 );
or OR2_9038 ( R1138_U293 , U4036 , U3072 );
nand NAND2_9039 ( R1138_U294 , R1138_U293 , R1138_U291 );
not NOT1_9040 ( R1138_U295 , R1138_U175 );
or OR2_9041 ( R1138_U296 , U4035 , U3058 );
nand NAND2_9042 ( R1138_U297 , U3058 , U4035 );
not NOT1_9043 ( R1138_U298 , R1138_U94 );
or OR2_9044 ( R1138_U299 , U4034 , U3063 );
nand NAND2_9045 ( R1138_U300 , R1138_U299 , R1138_U94 );
nand NAND2_9046 ( R1138_U301 , U3063 , U4034 );
not NOT1_9047 ( R1138_U302 , R1138_U172 );
or OR2_9048 ( R1138_U303 , U3055 , U4032 );
nand NAND2_9049 ( R1138_U304 , R1138_U193 , R1138_U185 );
or OR2_9050 ( R1138_U305 , U4033 , U3062 );
or OR2_9051 ( R1138_U306 , U4031 , U3054 );
nand NAND2_9052 ( R1138_U307 , R1138_U149 , R1138_U392 );
not NOT1_9053 ( R1138_U308 , R1138_U171 );
or OR2_9054 ( R1138_U309 , U4030 , U3050 );
nand NAND2_9055 ( R1138_U310 , U3050 , U4030 );
not NOT1_9056 ( R1138_U311 , R1138_U169 );
nand NAND2_9057 ( R1138_U312 , U4029 , R1138_U169 );
not NOT1_9058 ( R1138_U313 , R1138_U167 );
nand NAND2_9059 ( R1138_U314 , R1138_U305 , R1138_U172 );
not NOT1_9060 ( R1138_U315 , R1138_U100 );
or OR2_9061 ( R1138_U316 , U4032 , U3055 );
nand NAND2_9062 ( R1138_U317 , R1138_U316 , R1138_U100 );
nand NAND2_9063 ( R1138_U318 , R1138_U151 , R1138_U317 );
nand NAND2_9064 ( R1138_U319 , R1138_U315 , R1138_U190 );
nand NAND2_9065 ( R1138_U320 , U4031 , U3054 );
nand NAND2_9066 ( R1138_U321 , R1138_U152 , R1138_U319 );
or OR2_9067 ( R1138_U322 , U3055 , U4032 );
nand NAND2_9068 ( R1138_U323 , R1138_U292 , R1138_U179 );
not NOT1_9069 ( R1138_U324 , R1138_U104 );
nand NAND2_9070 ( R1138_U325 , R1138_U10 , R1138_U104 );
nand NAND2_9071 ( R1138_U326 , R1138_U153 , R1138_U325 );
nand NAND2_9072 ( R1138_U327 , R1138_U325 , R1138_U288 );
nand NAND2_9073 ( R1138_U328 , R1138_U480 , R1138_U327 );
or OR2_9074 ( R1138_U329 , U3504 , U3078 );
nand NAND2_9075 ( R1138_U330 , R1138_U329 , R1138_U104 );
nand NAND2_9076 ( R1138_U331 , R1138_U154 , R1138_U330 );
nand NAND2_9077 ( R1138_U332 , R1138_U324 , R1138_U80 );
nand NAND2_9078 ( R1138_U333 , U3073 , U4037 );
nand NAND2_9079 ( R1138_U334 , R1138_U155 , R1138_U332 );
or OR2_9080 ( R1138_U335 , U3468 , U3075 );
not NOT1_9081 ( R1138_U336 , R1138_U178 );
or OR2_9082 ( R1138_U337 , U3078 , U3504 );
or OR2_9083 ( R1138_U338 , U3498 , U3070 );
nand NAND2_9084 ( R1138_U339 , R1138_U338 , R1138_U105 );
nand NAND2_9085 ( R1138_U340 , R1138_U156 , R1138_U339 );
nand NAND2_9086 ( R1138_U341 , R1138_U272 , R1138_U90 );
nand NAND2_9087 ( R1138_U342 , U3500 , U3066 );
nand NAND2_9088 ( R1138_U343 , R1138_U157 , R1138_U341 );
or OR2_9089 ( R1138_U344 , U3070 , U3498 );
nand NAND2_9090 ( R1138_U345 , R1138_U262 , R1138_U184 );
not NOT1_9091 ( R1138_U346 , R1138_U106 );
or OR2_9092 ( R1138_U347 , U3490 , U3069 );
nand NAND2_9093 ( R1138_U348 , R1138_U347 , R1138_U106 );
nand NAND2_9094 ( R1138_U349 , R1138_U158 , R1138_U348 );
nand NAND2_9095 ( R1138_U350 , R1138_U346 , R1138_U189 );
nand NAND2_9096 ( R1138_U351 , U3077 , U3492 );
nand NAND2_9097 ( R1138_U352 , R1138_U159 , R1138_U350 );
or OR2_9098 ( R1138_U353 , U3069 , U3490 );
or OR2_9099 ( R1138_U354 , U3484 , U3080 );
nand NAND2_9100 ( R1138_U355 , R1138_U354 , R1138_U50 );
nand NAND2_9101 ( R1138_U356 , R1138_U160 , R1138_U355 );
nand NAND2_9102 ( R1138_U357 , R1138_U219 , R1138_U188 );
nand NAND2_9103 ( R1138_U358 , U3059 , U3486 );
nand NAND2_9104 ( R1138_U359 , R1138_U161 , R1138_U357 );
nand NAND2_9105 ( R1138_U360 , R1138_U220 , R1138_U188 );
nand NAND2_9106 ( R1138_U361 , R1138_U217 , R1138_U65 );
nand NAND2_9107 ( R1138_U362 , R1138_U227 , R1138_U43 );
nand NAND2_9108 ( R1138_U363 , R1138_U241 , R1138_U34 );
nand NAND2_9109 ( R1138_U364 , R1138_U244 , R1138_U197 );
nand NAND2_9110 ( R1138_U365 , R1138_U322 , R1138_U190 );
nand NAND2_9111 ( R1138_U366 , R1138_U305 , R1138_U60 );
nand NAND2_9112 ( R1138_U367 , R1138_U337 , R1138_U80 );
nand NAND2_9113 ( R1138_U368 , R1138_U292 , R1138_U84 );
nand NAND2_9114 ( R1138_U369 , R1138_U344 , R1138_U90 );
nand NAND2_9115 ( R1138_U370 , R1138_U353 , R1138_U189 );
nand NAND2_9116 ( R1138_U371 , R1138_U262 , R1138_U72 );
nand NAND2_9117 ( R1138_U372 , U4029 , U3051 );
nand NAND3_9118 ( R1138_U373 , R1138_U202 , R1138_U4 , R1138_U5 );
nand NAND3_9119 ( R1138_U374 , R1138_U5 , R1138_U4 , R1138_U201 );
not NOT1_9120 ( R1138_U375 , R1138_U45 );
not NOT1_9121 ( R1138_U376 , R1138_U102 );
nand NAND2_9122 ( R1138_U377 , R1138_U141 , R1138_U51 );
nand NAND2_9123 ( R1138_U378 , R1138_U12 , R1138_U45 );
nand NAND2_9124 ( R1138_U379 , R1138_U15 , R1138_U184 );
nand NAND2_9125 ( R1138_U380 , R1138_U268 , R1138_U265 );
not NOT1_9126 ( R1138_U381 , R1138_U77 );
nand NAND2_9127 ( R1138_U382 , R1138_U143 , R1138_U184 );
nand NAND2_9128 ( R1138_U383 , R1138_U381 , R1138_U270 );
nand NAND2_9129 ( R1138_U384 , R1138_U16 , R1138_U105 );
nand NAND2_9130 ( R1138_U385 , R1138_U14 , R1138_U102 );
not NOT1_9131 ( R1138_U386 , R1138_U101 );
not NOT1_9132 ( R1138_U387 , R1138_U97 );
nand NAND2_9133 ( R1138_U388 , R1138_U145 , R1138_U105 );
nand NAND2_9134 ( R1138_U389 , R1138_U101 , R1138_U296 );
nand NAND2_9135 ( R1138_U390 , U3054 , R1138_U303 );
nand NAND2_9136 ( R1138_U391 , U4031 , R1138_U303 );
nand NAND2_9137 ( R1138_U392 , R1138_U298 , R1138_U301 );
nand NAND3_9138 ( R1138_U393 , R1138_U193 , R1138_U185 , R1138_U309 );
nand NAND3_9139 ( R1138_U394 , R1138_U17 , R1138_U392 , R1138_U147 );
nand NAND2_9140 ( R1138_U395 , R1138_U387 , R1138_U309 );
nand NAND2_9141 ( R1138_U396 , R1138_U57 , R1138_U190 );
nand NAND2_9142 ( R1138_U397 , R1138_U56 , R1138_U190 );
nand NAND2_9143 ( R1138_U398 , U3080 , R1138_U49 );
nand NAND2_9144 ( R1138_U399 , U3484 , R1138_U48 );
nand NAND2_9145 ( R1138_U400 , R1138_U399 , R1138_U398 );
nand NAND2_9146 ( R1138_U401 , R1138_U360 , R1138_U50 );
nand NAND2_9147 ( R1138_U402 , R1138_U400 , R1138_U219 );
nand NAND2_9148 ( R1138_U403 , U3081 , R1138_U46 );
nand NAND2_9149 ( R1138_U404 , U3482 , R1138_U47 );
nand NAND2_9150 ( R1138_U405 , R1138_U404 , R1138_U403 );
nand NAND2_9151 ( R1138_U406 , R1138_U361 , R1138_U162 );
nand NAND2_9152 ( R1138_U407 , R1138_U216 , R1138_U405 );
nand NAND2_9153 ( R1138_U408 , U3067 , R1138_U44 );
nand NAND2_9154 ( R1138_U409 , U3480 , R1138_U42 );
nand NAND2_9155 ( R1138_U410 , U3068 , R1138_U40 );
nand NAND2_9156 ( R1138_U411 , U3478 , R1138_U41 );
nand NAND2_9157 ( R1138_U412 , R1138_U411 , R1138_U410 );
nand NAND2_9158 ( R1138_U413 , R1138_U362 , R1138_U51 );
nand NAND2_9159 ( R1138_U414 , R1138_U412 , R1138_U208 );
nand NAND2_9160 ( R1138_U415 , U3064 , R1138_U35 );
nand NAND2_9161 ( R1138_U416 , U3476 , R1138_U33 );
nand NAND2_9162 ( R1138_U417 , U3057 , R1138_U31 );
nand NAND2_9163 ( R1138_U418 , U3474 , R1138_U32 );
nand NAND2_9164 ( R1138_U419 , R1138_U418 , R1138_U417 );
nand NAND2_9165 ( R1138_U420 , R1138_U363 , R1138_U52 );
nand NAND2_9166 ( R1138_U421 , R1138_U419 , R1138_U234 );
nand NAND2_9167 ( R1138_U422 , U3061 , R1138_U29 );
nand NAND2_9168 ( R1138_U423 , U3472 , R1138_U30 );
nand NAND2_9169 ( R1138_U424 , R1138_U423 , R1138_U422 );
nand NAND2_9170 ( R1138_U425 , R1138_U364 , R1138_U163 );
nand NAND2_9171 ( R1138_U426 , R1138_U243 , R1138_U424 );
nand NAND2_9172 ( R1138_U427 , U3065 , R1138_U27 );
nand NAND2_9173 ( R1138_U428 , U3470 , R1138_U28 );
nand NAND2_9174 ( R1138_U429 , U3052 , R1138_U165 );
nand NAND2_9175 ( R1138_U430 , U4040 , R1138_U164 );
nand NAND2_9176 ( R1138_U431 , U3052 , R1138_U165 );
nand NAND2_9177 ( R1138_U432 , U4040 , R1138_U164 );
nand NAND2_9178 ( R1138_U433 , R1138_U432 , R1138_U431 );
nand NAND2_9179 ( R1138_U434 , R1138_U166 , R1138_U167 );
nand NAND2_9180 ( R1138_U435 , R1138_U313 , R1138_U433 );
nand NAND2_9181 ( R1138_U436 , U3051 , R1138_U99 );
nand NAND2_9182 ( R1138_U437 , U4029 , R1138_U98 );
nand NAND2_9183 ( R1138_U438 , U3051 , R1138_U99 );
nand NAND2_9184 ( R1138_U439 , U4029 , R1138_U98 );
nand NAND2_9185 ( R1138_U440 , R1138_U439 , R1138_U438 );
nand NAND2_9186 ( R1138_U441 , R1138_U168 , R1138_U169 );
nand NAND2_9187 ( R1138_U442 , R1138_U311 , R1138_U440 );
nand NAND2_9188 ( R1138_U443 , U3050 , R1138_U54 );
nand NAND2_9189 ( R1138_U444 , U4030 , R1138_U55 );
nand NAND2_9190 ( R1138_U445 , U3050 , R1138_U54 );
nand NAND2_9191 ( R1138_U446 , U4030 , R1138_U55 );
nand NAND2_9192 ( R1138_U447 , R1138_U446 , R1138_U445 );
nand NAND2_9193 ( R1138_U448 , R1138_U170 , R1138_U171 );
nand NAND2_9194 ( R1138_U449 , R1138_U308 , R1138_U447 );
nand NAND2_9195 ( R1138_U450 , U3054 , R1138_U57 );
nand NAND2_9196 ( R1138_U451 , U4031 , R1138_U56 );
nand NAND2_9197 ( R1138_U452 , U3055 , R1138_U95 );
nand NAND2_9198 ( R1138_U453 , U4032 , R1138_U96 );
nand NAND2_9199 ( R1138_U454 , R1138_U453 , R1138_U452 );
nand NAND2_9200 ( R1138_U455 , R1138_U365 , R1138_U100 );
nand NAND2_9201 ( R1138_U456 , R1138_U454 , R1138_U315 );
nand NAND2_9202 ( R1138_U457 , U3062 , R1138_U58 );
nand NAND2_9203 ( R1138_U458 , U4033 , R1138_U59 );
nand NAND2_9204 ( R1138_U459 , R1138_U458 , R1138_U457 );
nand NAND2_9205 ( R1138_U460 , R1138_U366 , R1138_U172 );
nand NAND2_9206 ( R1138_U461 , R1138_U302 , R1138_U459 );
nand NAND2_9207 ( R1138_U462 , U3063 , R1138_U92 );
nand NAND2_9208 ( R1138_U463 , U4034 , R1138_U93 );
nand NAND2_9209 ( R1138_U464 , U3063 , R1138_U92 );
nand NAND2_9210 ( R1138_U465 , U4034 , R1138_U93 );
nand NAND2_9211 ( R1138_U466 , R1138_U465 , R1138_U464 );
nand NAND2_9212 ( R1138_U467 , R1138_U173 , R1138_U94 );
nand NAND2_9213 ( R1138_U468 , R1138_U466 , R1138_U298 );
nand NAND2_9214 ( R1138_U469 , U3058 , R1138_U61 );
nand NAND2_9215 ( R1138_U470 , U4035 , R1138_U62 );
nand NAND2_9216 ( R1138_U471 , U3058 , R1138_U61 );
nand NAND2_9217 ( R1138_U472 , U4035 , R1138_U62 );
nand NAND2_9218 ( R1138_U473 , R1138_U472 , R1138_U471 );
nand NAND2_9219 ( R1138_U474 , R1138_U174 , R1138_U175 );
nand NAND2_9220 ( R1138_U475 , R1138_U295 , R1138_U473 );
nand NAND2_9221 ( R1138_U476 , U3072 , R1138_U85 );
nand NAND2_9222 ( R1138_U477 , U4036 , R1138_U86 );
nand NAND2_9223 ( R1138_U478 , U3072 , R1138_U85 );
nand NAND2_9224 ( R1138_U479 , U4036 , R1138_U86 );
nand NAND2_9225 ( R1138_U480 , R1138_U479 , R1138_U478 );
nand NAND2_9226 ( R1138_U481 , U3073 , R1138_U81 );
nand NAND2_9227 ( R1138_U482 , U4037 , R1138_U103 );
nand NAND2_9228 ( R1138_U483 , R1138_U199 , R1138_U178 );
nand NAND2_9229 ( R1138_U484 , R1138_U336 , R1138_U177 );
nand NAND2_9230 ( R1138_U485 , U3078 , R1138_U78 );
nand NAND2_9231 ( R1138_U486 , U3504 , R1138_U79 );
nand NAND2_9232 ( R1138_U487 , R1138_U486 , R1138_U485 );
nand NAND2_9233 ( R1138_U488 , R1138_U367 , R1138_U104 );
nand NAND2_9234 ( R1138_U489 , R1138_U487 , R1138_U324 );
nand NAND2_9235 ( R1138_U490 , U3079 , R1138_U82 );
nand NAND2_9236 ( R1138_U491 , U3502 , R1138_U83 );
nand NAND2_9237 ( R1138_U492 , R1138_U491 , R1138_U490 );
nand NAND2_9238 ( R1138_U493 , R1138_U368 , R1138_U179 );
nand NAND2_9239 ( R1138_U494 , R1138_U280 , R1138_U492 );
nand NAND2_9240 ( R1138_U495 , U3066 , R1138_U91 );
nand NAND2_9241 ( R1138_U496 , U3500 , R1138_U89 );
nand NAND2_9242 ( R1138_U497 , U3070 , R1138_U87 );
nand NAND2_9243 ( R1138_U498 , U3498 , R1138_U88 );
nand NAND2_9244 ( R1138_U499 , R1138_U498 , R1138_U497 );
nand NAND2_9245 ( R1138_U500 , R1138_U369 , R1138_U105 );
nand NAND2_9246 ( R1138_U501 , R1138_U499 , R1138_U272 );
nand NAND2_9247 ( R1138_U502 , U3071 , R1138_U63 );
nand NAND2_9248 ( R1138_U503 , U3496 , R1138_U64 );
nand NAND2_9249 ( R1138_U504 , U3071 , R1138_U63 );
nand NAND2_9250 ( R1138_U505 , U3496 , R1138_U64 );
nand NAND2_9251 ( R1138_U506 , R1138_U505 , R1138_U504 );
nand NAND2_9252 ( R1138_U507 , R1138_U180 , R1138_U181 );
nand NAND2_9253 ( R1138_U508 , R1138_U269 , R1138_U506 );
nand NAND2_9254 ( R1138_U509 , U3076 , R1138_U75 );
nand NAND2_9255 ( R1138_U510 , U3494 , R1138_U76 );
nand NAND2_9256 ( R1138_U511 , U3076 , R1138_U75 );
nand NAND2_9257 ( R1138_U512 , U3494 , R1138_U76 );
nand NAND2_9258 ( R1138_U513 , R1138_U512 , R1138_U511 );
nand NAND2_9259 ( R1138_U514 , R1138_U182 , R1138_U183 );
nand NAND2_9260 ( R1138_U515 , R1138_U266 , R1138_U513 );
nand NAND2_9261 ( R1138_U516 , U3077 , R1138_U73 );
nand NAND2_9262 ( R1138_U517 , U3492 , R1138_U74 );
nand NAND2_9263 ( R1138_U518 , U3069 , R1138_U68 );
nand NAND2_9264 ( R1138_U519 , U3490 , R1138_U69 );
nand NAND2_9265 ( R1138_U520 , R1138_U519 , R1138_U518 );
nand NAND2_9266 ( R1138_U521 , R1138_U370 , R1138_U106 );
nand NAND2_9267 ( R1138_U522 , R1138_U520 , R1138_U346 );
nand NAND2_9268 ( R1138_U523 , U3060 , R1138_U70 );
nand NAND2_9269 ( R1138_U524 , U3488 , R1138_U71 );
nand NAND2_9270 ( R1138_U525 , R1138_U524 , R1138_U523 );
nand NAND2_9271 ( R1138_U526 , R1138_U371 , R1138_U184 );
nand NAND2_9272 ( R1138_U527 , R1138_U256 , R1138_U525 );
nand NAND2_9273 ( R1138_U528 , U3059 , R1138_U66 );
nand NAND2_9274 ( R1138_U529 , U3486 , R1138_U67 );
nand NAND2_9275 ( R1138_U530 , U3074 , R1138_U37 );
nand NAND2_9276 ( R1138_U531 , U3464 , R1138_U38 );
and AND2_9277 ( R1222_U4 , R1222_U190 , R1222_U189 );
and AND2_9278 ( R1222_U5 , R1222_U191 , R1222_U192 );
and AND2_9279 ( R1222_U6 , R1222_U204 , R1222_U203 );
and AND2_9280 ( R1222_U7 , R1222_U239 , R1222_U238 );
and AND2_9281 ( R1222_U8 , R1222_U246 , R1222_U245 );
and AND2_9282 ( R1222_U9 , R1222_U262 , R1222_U261 );
and AND2_9283 ( R1222_U10 , R1222_U268 , R1222_U267 );
and AND2_9284 ( R1222_U11 , R1222_U10 , R1222_U269 );
and AND2_9285 ( R1222_U12 , R1222_U290 , R1222_U289 );
and AND2_9286 ( R1222_U13 , R1222_U7 , R1222_U209 );
and AND2_9287 ( R1222_U14 , R1222_U8 , R1222_U250 );
and AND2_9288 ( R1222_U15 , R1222_U11 , R1222_U278 );
and AND2_9289 ( R1222_U16 , R1222_U14 , R1222_U255 );
and AND2_9290 ( R1222_U17 , R1222_U347 , R1222_U344 );
and AND2_9291 ( R1222_U18 , R1222_U340 , R1222_U337 );
and AND2_9292 ( R1222_U19 , R1222_U331 , R1222_U383 );
and AND2_9293 ( R1222_U20 , R1222_U325 , R1222_U322 );
and AND2_9294 ( R1222_U21 , R1222_U319 , R1222_U317 );
and AND2_9295 ( R1222_U22 , R1222_U312 , R1222_U309 );
and AND2_9296 ( R1222_U23 , R1222_U237 , R1222_U234 );
and AND2_9297 ( R1222_U24 , R1222_U229 , R1222_U226 );
and AND2_9298 ( R1222_U25 , R1222_U215 , R1222_U376 );
not NOT1_9299 ( R1222_U26 , U3478 );
not NOT1_9300 ( R1222_U27 , U3068 );
not NOT1_9301 ( R1222_U28 , U3067 );
nand NAND2_9302 ( R1222_U29 , U3068 , U3478 );
not NOT1_9303 ( R1222_U30 , U3480 );
not NOT1_9304 ( R1222_U31 , U3470 );
not NOT1_9305 ( R1222_U32 , U3065 );
not NOT1_9306 ( R1222_U33 , U3472 );
not NOT1_9307 ( R1222_U34 , U3061 );
not NOT1_9308 ( R1222_U35 , U3474 );
not NOT1_9309 ( R1222_U36 , U3057 );
not NOT1_9310 ( R1222_U37 , U3064 );
nand NAND2_9311 ( R1222_U38 , U3057 , U3474 );
not NOT1_9312 ( R1222_U39 , U3476 );
nand NAND2_9313 ( R1222_U40 , U3468 , U3075 );
not NOT1_9314 ( R1222_U41 , U3464 );
not NOT1_9315 ( R1222_U42 , U3074 );
nand NAND2_9316 ( R1222_U43 , R1222_U127 , R1222_U194 );
nand NAND2_9317 ( R1222_U44 , R1222_U208 , R1222_U207 );
not NOT1_9318 ( R1222_U45 , U3482 );
not NOT1_9319 ( R1222_U46 , U3081 );
not NOT1_9320 ( R1222_U47 , U3080 );
not NOT1_9321 ( R1222_U48 , U3484 );
nand NAND2_9322 ( R1222_U49 , R1222_U69 , R1222_U210 );
nand NAND2_9323 ( R1222_U50 , R1222_U129 , R1222_U128 );
nand NAND2_9324 ( R1222_U51 , R1222_U132 , R1222_U221 );
nand NAND2_9325 ( R1222_U52 , R1222_U218 , R1222_U217 );
not NOT1_9326 ( R1222_U53 , U3504 );
not NOT1_9327 ( R1222_U54 , U3078 );
nand NAND2_9328 ( R1222_U55 , U3078 , U3504 );
not NOT1_9329 ( R1222_U56 , U4037 );
not NOT1_9330 ( R1222_U57 , U3502 );
not NOT1_9331 ( R1222_U58 , U3079 );
nand NAND2_9332 ( R1222_U59 , U3079 , U3502 );
not NOT1_9333 ( R1222_U60 , U4036 );
not NOT1_9334 ( R1222_U61 , U3072 );
not NOT1_9335 ( R1222_U62 , U3498 );
not NOT1_9336 ( R1222_U63 , U3070 );
not NOT1_9337 ( R1222_U64 , U3066 );
nand NAND2_9338 ( R1222_U65 , U3070 , U3498 );
not NOT1_9339 ( R1222_U66 , U3500 );
not NOT1_9340 ( R1222_U67 , U3496 );
not NOT1_9341 ( R1222_U68 , U3071 );
nand NAND2_9342 ( R1222_U69 , U3081 , U3482 );
not NOT1_9343 ( R1222_U70 , U3486 );
not NOT1_9344 ( R1222_U71 , U3059 );
not NOT1_9345 ( R1222_U72 , U3490 );
not NOT1_9346 ( R1222_U73 , U3069 );
not NOT1_9347 ( R1222_U74 , U3488 );
not NOT1_9348 ( R1222_U75 , U3060 );
nand NAND2_9349 ( R1222_U76 , U3060 , U3488 );
not NOT1_9350 ( R1222_U77 , U3492 );
not NOT1_9351 ( R1222_U78 , U3077 );
not NOT1_9352 ( R1222_U79 , U3494 );
not NOT1_9353 ( R1222_U80 , U3076 );
nand NAND2_9354 ( R1222_U81 , R1222_U367 , R1222_U255 );
not NOT1_9355 ( R1222_U82 , U4035 );
not NOT1_9356 ( R1222_U83 , U3058 );
not NOT1_9357 ( R1222_U84 , U4034 );
not NOT1_9358 ( R1222_U85 , U3063 );
not NOT1_9359 ( R1222_U86 , U4032 );
not NOT1_9360 ( R1222_U87 , U3055 );
not NOT1_9361 ( R1222_U88 , U4033 );
not NOT1_9362 ( R1222_U89 , U3062 );
nand NAND2_9363 ( R1222_U90 , U3062 , U4033 );
not NOT1_9364 ( R1222_U91 , U4031 );
not NOT1_9365 ( R1222_U92 , U3054 );
not NOT1_9366 ( R1222_U93 , U4030 );
not NOT1_9367 ( R1222_U94 , U3050 );
not NOT1_9368 ( R1222_U95 , U3051 );
not NOT1_9369 ( R1222_U96 , U4029 );
nand NAND2_9370 ( R1222_U97 , R1222_U90 , R1222_U305 );
nand NAND2_9371 ( R1222_U98 , R1222_U266 , R1222_U265 );
not NOT1_9372 ( R1222_U99 , U3073 );
nand NAND2_9373 ( R1222_U100 , R1222_U59 , R1222_U314 );
nand NAND3_9374 ( R1222_U101 , R1222_U370 , R1222_U259 , R1222_U369 );
nand NAND2_9375 ( R1222_U102 , R1222_U76 , R1222_U333 );
nand NAND2_9376 ( R1222_U103 , R1222_U472 , R1222_U471 );
nand NAND2_9377 ( R1222_U104 , R1222_U519 , R1222_U518 );
nand NAND2_9378 ( R1222_U105 , R1222_U390 , R1222_U389 );
nand NAND2_9379 ( R1222_U106 , R1222_U395 , R1222_U394 );
nand NAND2_9380 ( R1222_U107 , R1222_U402 , R1222_U401 );
nand NAND2_9381 ( R1222_U108 , R1222_U409 , R1222_U408 );
nand NAND2_9382 ( R1222_U109 , R1222_U414 , R1222_U413 );
nand NAND2_9383 ( R1222_U110 , R1222_U423 , R1222_U422 );
nand NAND2_9384 ( R1222_U111 , R1222_U430 , R1222_U429 );
nand NAND2_9385 ( R1222_U112 , R1222_U437 , R1222_U436 );
nand NAND2_9386 ( R1222_U113 , R1222_U444 , R1222_U443 );
nand NAND2_9387 ( R1222_U114 , R1222_U449 , R1222_U448 );
nand NAND2_9388 ( R1222_U115 , R1222_U456 , R1222_U455 );
nand NAND2_9389 ( R1222_U116 , R1222_U463 , R1222_U462 );
nand NAND2_9390 ( R1222_U117 , R1222_U477 , R1222_U476 );
nand NAND2_9391 ( R1222_U118 , R1222_U482 , R1222_U481 );
nand NAND2_9392 ( R1222_U119 , R1222_U489 , R1222_U488 );
nand NAND2_9393 ( R1222_U120 , R1222_U496 , R1222_U495 );
nand NAND2_9394 ( R1222_U121 , R1222_U503 , R1222_U502 );
nand NAND2_9395 ( R1222_U122 , R1222_U510 , R1222_U509 );
nand NAND2_9396 ( R1222_U123 , R1222_U515 , R1222_U514 );
and AND2_9397 ( R1222_U124 , R1222_U125 , R1222_U191 );
and AND2_9398 ( R1222_U125 , U3065 , U3470 );
and AND2_9399 ( R1222_U126 , U3472 , U3061 );
and AND2_9400 ( R1222_U127 , U3464 , U3074 );
and AND3_9401 ( R1222_U128 , R1222_U198 , R1222_U200 , R1222_U197 );
and AND3_9402 ( R1222_U129 , R1222_U361 , R1222_U201 , R1222_U362 );
and AND3_9403 ( R1222_U130 , R1222_U397 , R1222_U396 , R1222_U29 );
and AND2_9404 ( R1222_U131 , R1222_U6 , R1222_U214 );
and AND2_9405 ( R1222_U132 , R1222_U222 , R1222_U220 );
and AND3_9406 ( R1222_U133 , R1222_U404 , R1222_U403 , R1222_U38 );
and AND2_9407 ( R1222_U134 , R1222_U228 , R1222_U4 );
and AND2_9408 ( R1222_U135 , R1222_U236 , R1222_U192 );
and AND2_9409 ( R1222_U136 , R1222_U241 , R1222_U182 );
and AND2_9410 ( R1222_U137 , R1222_U6 , R1222_U13 );
and AND2_9411 ( R1222_U138 , R1222_U365 , R1222_U244 );
and AND2_9412 ( R1222_U139 , R1222_U16 , R1222_U258 );
and AND2_9413 ( R1222_U140 , R1222_U248 , R1222_U183 );
and AND2_9414 ( R1222_U141 , R1222_U15 , R1222_U9 );
and AND2_9415 ( R1222_U142 , R1222_U371 , R1222_U280 );
and AND2_9416 ( R1222_U143 , R1222_U294 , R1222_U12 );
and AND2_9417 ( R1222_U144 , R1222_U292 , R1222_U184 );
and AND3_9418 ( R1222_U145 , R1222_U439 , R1222_U438 , R1222_U184 );
and AND2_9419 ( R1222_U146 , R1222_U311 , R1222_U12 );
and AND2_9420 ( R1222_U147 , R1222_U171 , R1222_U274 );
and AND3_9421 ( R1222_U148 , R1222_U470 , R1222_U469 , R1222_U55 );
and AND2_9422 ( R1222_U149 , R1222_U324 , R1222_U10 );
and AND3_9423 ( R1222_U150 , R1222_U484 , R1222_U483 , R1222_U65 );
and AND2_9424 ( R1222_U151 , R1222_U9 , R1222_U330 );
and AND3_9425 ( R1222_U152 , R1222_U505 , R1222_U504 , R1222_U183 );
and AND2_9426 ( R1222_U153 , R1222_U339 , R1222_U8 );
and AND3_9427 ( R1222_U154 , R1222_U517 , R1222_U516 , R1222_U182 );
and AND2_9428 ( R1222_U155 , R1222_U346 , R1222_U7 );
nand NAND2_9429 ( R1222_U156 , R1222_U363 , R1222_U373 );
nand NAND2_9430 ( R1222_U157 , R1222_U219 , R1222_U231 );
not NOT1_9431 ( R1222_U158 , U3052 );
not NOT1_9432 ( R1222_U159 , U4040 );
and AND2_9433 ( R1222_U160 , R1222_U418 , R1222_U417 );
nand NAND3_9434 ( R1222_U161 , R1222_U303 , R1222_U180 , R1222_U360 );
and AND2_9435 ( R1222_U162 , R1222_U425 , R1222_U424 );
nand NAND2_9436 ( R1222_U163 , R1222_U301 , R1222_U300 );
and AND2_9437 ( R1222_U164 , R1222_U432 , R1222_U431 );
nand NAND2_9438 ( R1222_U165 , R1222_U297 , R1222_U296 );
nand NAND2_9439 ( R1222_U166 , R1222_U287 , R1222_U286 );
and AND2_9440 ( R1222_U167 , R1222_U451 , R1222_U450 );
nand NAND2_9441 ( R1222_U168 , R1222_U283 , R1222_U282 );
and AND2_9442 ( R1222_U169 , R1222_U458 , R1222_U457 );
nand NAND2_9443 ( R1222_U170 , R1222_U142 , R1222_U384 );
and AND2_9444 ( R1222_U171 , R1222_U465 , R1222_U464 );
nand NAND2_9445 ( R1222_U172 , U3074 , U3464 );
nand NAND2_9446 ( R1222_U173 , R1222_U40 , R1222_U326 );
nand NAND2_9447 ( R1222_U174 , R1222_U364 , R1222_U380 );
and AND2_9448 ( R1222_U175 , R1222_U491 , R1222_U490 );
nand NAND2_9449 ( R1222_U176 , R1222_U81 , R1222_U366 );
and AND2_9450 ( R1222_U177 , R1222_U498 , R1222_U497 );
nand NAND2_9451 ( R1222_U178 , R1222_U253 , R1222_U252 );
nand NAND2_9452 ( R1222_U179 , R1222_U138 , R1222_U377 );
nand NAND2_9453 ( R1222_U180 , U3051 , R1222_U163 );
not NOT1_9454 ( R1222_U181 , R1222_U38 );
nand NAND2_9455 ( R1222_U182 , U3484 , U3080 );
nand NAND2_9456 ( R1222_U183 , U3069 , U3490 );
nand NAND2_9457 ( R1222_U184 , U3055 , U4032 );
not NOT1_9458 ( R1222_U185 , R1222_U76 );
not NOT1_9459 ( R1222_U186 , R1222_U59 );
not NOT1_9460 ( R1222_U187 , R1222_U90 );
not NOT1_9461 ( R1222_U188 , R1222_U69 );
or OR2_9462 ( R1222_U189 , U3064 , U3476 );
or OR2_9463 ( R1222_U190 , U3057 , U3474 );
or OR2_9464 ( R1222_U191 , U3472 , U3061 );
or OR2_9465 ( R1222_U192 , U3470 , U3065 );
not NOT1_9466 ( R1222_U193 , R1222_U172 );
or OR2_9467 ( R1222_U194 , U3468 , U3075 );
not NOT1_9468 ( R1222_U195 , R1222_U43 );
not NOT1_9469 ( R1222_U196 , R1222_U40 );
nand NAND2_9470 ( R1222_U197 , R1222_U4 , R1222_U124 );
nand NAND2_9471 ( R1222_U198 , R1222_U126 , R1222_U4 );
nand NAND2_9472 ( R1222_U199 , R1222_U39 , R1222_U38 );
nand NAND2_9473 ( R1222_U200 , U3064 , R1222_U199 );
nand NAND2_9474 ( R1222_U201 , U3476 , R1222_U181 );
not NOT1_9475 ( R1222_U202 , R1222_U50 );
or OR2_9476 ( R1222_U203 , U3067 , U3480 );
or OR2_9477 ( R1222_U204 , U3068 , U3478 );
not NOT1_9478 ( R1222_U205 , R1222_U29 );
nand NAND2_9479 ( R1222_U206 , R1222_U30 , R1222_U29 );
nand NAND2_9480 ( R1222_U207 , U3067 , R1222_U206 );
nand NAND2_9481 ( R1222_U208 , U3480 , R1222_U205 );
or OR2_9482 ( R1222_U209 , U3482 , U3081 );
nand NAND2_9483 ( R1222_U210 , R1222_U209 , R1222_U156 );
not NOT1_9484 ( R1222_U211 , R1222_U49 );
or OR2_9485 ( R1222_U212 , U3080 , U3484 );
or OR2_9486 ( R1222_U213 , U3478 , U3068 );
nand NAND2_9487 ( R1222_U214 , U3480 , U3067 );
nand NAND2_9488 ( R1222_U215 , R1222_U131 , R1222_U372 );
or OR2_9489 ( R1222_U216 , U3068 , U3478 );
nand NAND2_9490 ( R1222_U217 , R1222_U196 , R1222_U192 );
nand NAND2_9491 ( R1222_U218 , U3065 , U3470 );
not NOT1_9492 ( R1222_U219 , R1222_U52 );
nand NAND2_9493 ( R1222_U220 , R1222_U195 , R1222_U5 );
nand NAND2_9494 ( R1222_U221 , R1222_U52 , R1222_U191 );
nand NAND2_9495 ( R1222_U222 , U3061 , U3472 );
not NOT1_9496 ( R1222_U223 , R1222_U51 );
or OR2_9497 ( R1222_U224 , U3474 , U3057 );
nand NAND2_9498 ( R1222_U225 , R1222_U224 , R1222_U51 );
nand NAND2_9499 ( R1222_U226 , R1222_U133 , R1222_U225 );
nand NAND2_9500 ( R1222_U227 , R1222_U223 , R1222_U38 );
nand NAND2_9501 ( R1222_U228 , U3476 , U3064 );
nand NAND2_9502 ( R1222_U229 , R1222_U134 , R1222_U227 );
or OR2_9503 ( R1222_U230 , U3057 , U3474 );
nand NAND2_9504 ( R1222_U231 , R1222_U195 , R1222_U192 );
not NOT1_9505 ( R1222_U232 , R1222_U157 );
nand NAND2_9506 ( R1222_U233 , U3061 , U3472 );
nand NAND4_9507 ( R1222_U234 , R1222_U416 , R1222_U415 , R1222_U40 , R1222_U43 );
nand NAND2_9508 ( R1222_U235 , R1222_U40 , R1222_U43 );
nand NAND2_9509 ( R1222_U236 , U3065 , U3470 );
nand NAND2_9510 ( R1222_U237 , R1222_U135 , R1222_U235 );
or OR2_9511 ( R1222_U238 , U3080 , U3484 );
or OR2_9512 ( R1222_U239 , U3059 , U3486 );
nand NAND2_9513 ( R1222_U240 , R1222_U188 , R1222_U7 );
nand NAND2_9514 ( R1222_U241 , U3059 , U3486 );
nand NAND2_9515 ( R1222_U242 , R1222_U136 , R1222_U240 );
or OR2_9516 ( R1222_U243 , U3486 , U3059 );
nand NAND2_9517 ( R1222_U244 , R1222_U243 , R1222_U242 );
or OR2_9518 ( R1222_U245 , U3077 , U3492 );
or OR2_9519 ( R1222_U246 , U3069 , U3490 );
nand NAND2_9520 ( R1222_U247 , R1222_U185 , R1222_U8 );
nand NAND2_9521 ( R1222_U248 , U3077 , U3492 );
nand NAND2_9522 ( R1222_U249 , R1222_U140 , R1222_U247 );
or OR2_9523 ( R1222_U250 , U3488 , U3060 );
or OR2_9524 ( R1222_U251 , U3492 , U3077 );
nand NAND2_9525 ( R1222_U252 , R1222_U14 , R1222_U179 );
nand NAND2_9526 ( R1222_U253 , R1222_U251 , R1222_U249 );
not NOT1_9527 ( R1222_U254 , R1222_U178 );
or OR2_9528 ( R1222_U255 , U3494 , U3076 );
nand NAND2_9529 ( R1222_U256 , U3076 , U3494 );
not NOT1_9530 ( R1222_U257 , R1222_U176 );
or OR2_9531 ( R1222_U258 , U3496 , U3071 );
nand NAND2_9532 ( R1222_U259 , U3071 , U3496 );
not NOT1_9533 ( R1222_U260 , R1222_U101 );
or OR2_9534 ( R1222_U261 , U3066 , U3500 );
or OR2_9535 ( R1222_U262 , U3070 , U3498 );
not NOT1_9536 ( R1222_U263 , R1222_U65 );
nand NAND2_9537 ( R1222_U264 , R1222_U66 , R1222_U65 );
nand NAND2_9538 ( R1222_U265 , U3066 , R1222_U264 );
nand NAND2_9539 ( R1222_U266 , U3500 , R1222_U263 );
or OR2_9540 ( R1222_U267 , U3073 , U4037 );
or OR2_9541 ( R1222_U268 , U3078 , U3504 );
or OR2_9542 ( R1222_U269 , U3072 , U4036 );
not NOT1_9543 ( R1222_U270 , R1222_U55 );
nand NAND2_9544 ( R1222_U271 , U4037 , R1222_U270 );
nand NAND2_9545 ( R1222_U272 , R1222_U271 , R1222_U99 );
nand NAND2_9546 ( R1222_U273 , R1222_U55 , R1222_U56 );
nand NAND2_9547 ( R1222_U274 , R1222_U273 , R1222_U272 );
nand NAND2_9548 ( R1222_U275 , R1222_U186 , R1222_U11 );
nand NAND2_9549 ( R1222_U276 , U3072 , U4036 );
nand NAND3_9550 ( R1222_U277 , R1222_U275 , R1222_U274 , R1222_U276 );
or OR2_9551 ( R1222_U278 , U3502 , U3079 );
or OR2_9552 ( R1222_U279 , U4036 , U3072 );
nand NAND2_9553 ( R1222_U280 , R1222_U279 , R1222_U277 );
or OR2_9554 ( R1222_U281 , U4035 , U3058 );
nand NAND2_9555 ( R1222_U282 , R1222_U281 , R1222_U170 );
nand NAND2_9556 ( R1222_U283 , U3058 , U4035 );
not NOT1_9557 ( R1222_U284 , R1222_U168 );
or OR2_9558 ( R1222_U285 , U4034 , U3063 );
nand NAND2_9559 ( R1222_U286 , R1222_U285 , R1222_U168 );
nand NAND2_9560 ( R1222_U287 , U3063 , U4034 );
not NOT1_9561 ( R1222_U288 , R1222_U166 );
or OR2_9562 ( R1222_U289 , U3054 , U4031 );
or OR2_9563 ( R1222_U290 , U3055 , U4032 );
nand NAND2_9564 ( R1222_U291 , R1222_U187 , R1222_U12 );
nand NAND2_9565 ( R1222_U292 , U3054 , U4031 );
nand NAND2_9566 ( R1222_U293 , R1222_U144 , R1222_U291 );
or OR2_9567 ( R1222_U294 , U4033 , U3062 );
or OR2_9568 ( R1222_U295 , U4031 , U3054 );
nand NAND2_9569 ( R1222_U296 , R1222_U143 , R1222_U166 );
nand NAND2_9570 ( R1222_U297 , R1222_U295 , R1222_U293 );
not NOT1_9571 ( R1222_U298 , R1222_U165 );
or OR2_9572 ( R1222_U299 , U4030 , U3050 );
nand NAND2_9573 ( R1222_U300 , R1222_U299 , R1222_U165 );
nand NAND2_9574 ( R1222_U301 , U3050 , U4030 );
not NOT1_9575 ( R1222_U302 , R1222_U163 );
nand NAND2_9576 ( R1222_U303 , U4029 , R1222_U163 );
not NOT1_9577 ( R1222_U304 , R1222_U161 );
nand NAND2_9578 ( R1222_U305 , R1222_U294 , R1222_U166 );
not NOT1_9579 ( R1222_U306 , R1222_U97 );
or OR2_9580 ( R1222_U307 , U4032 , U3055 );
nand NAND2_9581 ( R1222_U308 , R1222_U307 , R1222_U97 );
nand NAND2_9582 ( R1222_U309 , R1222_U145 , R1222_U308 );
nand NAND2_9583 ( R1222_U310 , R1222_U306 , R1222_U184 );
nand NAND2_9584 ( R1222_U311 , U3054 , U4031 );
nand NAND2_9585 ( R1222_U312 , R1222_U146 , R1222_U310 );
or OR2_9586 ( R1222_U313 , U3055 , U4032 );
nand NAND2_9587 ( R1222_U314 , R1222_U278 , R1222_U174 );
not NOT1_9588 ( R1222_U315 , R1222_U100 );
nand NAND2_9589 ( R1222_U316 , R1222_U10 , R1222_U100 );
nand NAND2_9590 ( R1222_U317 , R1222_U147 , R1222_U316 );
nand NAND2_9591 ( R1222_U318 , R1222_U316 , R1222_U274 );
nand NAND2_9592 ( R1222_U319 , R1222_U468 , R1222_U318 );
or OR2_9593 ( R1222_U320 , U3504 , U3078 );
nand NAND2_9594 ( R1222_U321 , R1222_U320 , R1222_U100 );
nand NAND2_9595 ( R1222_U322 , R1222_U148 , R1222_U321 );
nand NAND2_9596 ( R1222_U323 , R1222_U315 , R1222_U55 );
nand NAND2_9597 ( R1222_U324 , U3073 , U4037 );
nand NAND2_9598 ( R1222_U325 , R1222_U149 , R1222_U323 );
or OR2_9599 ( R1222_U326 , U3468 , U3075 );
not NOT1_9600 ( R1222_U327 , R1222_U173 );
or OR2_9601 ( R1222_U328 , U3078 , U3504 );
or OR2_9602 ( R1222_U329 , U3498 , U3070 );
nand NAND2_9603 ( R1222_U330 , U3500 , U3066 );
nand NAND2_9604 ( R1222_U331 , R1222_U151 , R1222_U379 );
or OR2_9605 ( R1222_U332 , U3070 , U3498 );
nand NAND2_9606 ( R1222_U333 , R1222_U250 , R1222_U179 );
not NOT1_9607 ( R1222_U334 , R1222_U102 );
or OR2_9608 ( R1222_U335 , U3490 , U3069 );
nand NAND2_9609 ( R1222_U336 , R1222_U335 , R1222_U102 );
nand NAND2_9610 ( R1222_U337 , R1222_U152 , R1222_U336 );
nand NAND2_9611 ( R1222_U338 , R1222_U334 , R1222_U183 );
nand NAND2_9612 ( R1222_U339 , U3077 , U3492 );
nand NAND2_9613 ( R1222_U340 , R1222_U153 , R1222_U338 );
or OR2_9614 ( R1222_U341 , U3069 , U3490 );
or OR2_9615 ( R1222_U342 , U3484 , U3080 );
nand NAND2_9616 ( R1222_U343 , R1222_U342 , R1222_U49 );
nand NAND2_9617 ( R1222_U344 , R1222_U154 , R1222_U343 );
nand NAND2_9618 ( R1222_U345 , R1222_U211 , R1222_U182 );
nand NAND2_9619 ( R1222_U346 , U3059 , U3486 );
nand NAND2_9620 ( R1222_U347 , R1222_U155 , R1222_U345 );
nand NAND2_9621 ( R1222_U348 , R1222_U212 , R1222_U182 );
nand NAND2_9622 ( R1222_U349 , R1222_U209 , R1222_U69 );
nand NAND2_9623 ( R1222_U350 , R1222_U216 , R1222_U29 );
nand NAND2_9624 ( R1222_U351 , R1222_U230 , R1222_U38 );
nand NAND2_9625 ( R1222_U352 , R1222_U233 , R1222_U191 );
nand NAND2_9626 ( R1222_U353 , R1222_U313 , R1222_U184 );
nand NAND2_9627 ( R1222_U354 , R1222_U294 , R1222_U90 );
nand NAND2_9628 ( R1222_U355 , R1222_U328 , R1222_U55 );
nand NAND2_9629 ( R1222_U356 , R1222_U278 , R1222_U59 );
nand NAND2_9630 ( R1222_U357 , R1222_U332 , R1222_U65 );
nand NAND2_9631 ( R1222_U358 , R1222_U341 , R1222_U183 );
nand NAND2_9632 ( R1222_U359 , R1222_U250 , R1222_U76 );
nand NAND2_9633 ( R1222_U360 , U4029 , U3051 );
nand NAND3_9634 ( R1222_U361 , R1222_U196 , R1222_U4 , R1222_U5 );
nand NAND3_9635 ( R1222_U362 , R1222_U5 , R1222_U4 , R1222_U195 );
not NOT1_9636 ( R1222_U363 , R1222_U44 );
not NOT1_9637 ( R1222_U364 , R1222_U98 );
nand NAND2_9638 ( R1222_U365 , R1222_U13 , R1222_U44 );
nand NAND2_9639 ( R1222_U366 , R1222_U16 , R1222_U179 );
nand NAND2_9640 ( R1222_U367 , R1222_U256 , R1222_U253 );
not NOT1_9641 ( R1222_U368 , R1222_U81 );
nand NAND2_9642 ( R1222_U369 , R1222_U139 , R1222_U179 );
nand NAND2_9643 ( R1222_U370 , R1222_U368 , R1222_U258 );
nand NAND2_9644 ( R1222_U371 , R1222_U15 , R1222_U98 );
nand NAND2_9645 ( R1222_U372 , R1222_U202 , R1222_U29 );
nand NAND2_9646 ( R1222_U373 , R1222_U6 , R1222_U50 );
not NOT1_9647 ( R1222_U374 , R1222_U156 );
nand NAND2_9648 ( R1222_U375 , R1222_U213 , R1222_U50 );
nand NAND2_9649 ( R1222_U376 , R1222_U130 , R1222_U375 );
nand NAND2_9650 ( R1222_U377 , R1222_U137 , R1222_U50 );
not NOT1_9651 ( R1222_U378 , R1222_U179 );
nand NAND2_9652 ( R1222_U379 , R1222_U260 , R1222_U65 );
nand NAND2_9653 ( R1222_U380 , R1222_U9 , R1222_U101 );
not NOT1_9654 ( R1222_U381 , R1222_U174 );
nand NAND2_9655 ( R1222_U382 , R1222_U329 , R1222_U101 );
nand NAND2_9656 ( R1222_U383 , R1222_U150 , R1222_U382 );
nand NAND2_9657 ( R1222_U384 , R1222_U141 , R1222_U101 );
not NOT1_9658 ( R1222_U385 , R1222_U170 );
nand NAND2_9659 ( R1222_U386 , U3080 , R1222_U48 );
nand NAND2_9660 ( R1222_U387 , U3484 , R1222_U47 );
nand NAND2_9661 ( R1222_U388 , R1222_U387 , R1222_U386 );
nand NAND2_9662 ( R1222_U389 , R1222_U348 , R1222_U49 );
nand NAND2_9663 ( R1222_U390 , R1222_U388 , R1222_U211 );
nand NAND2_9664 ( R1222_U391 , U3081 , R1222_U45 );
nand NAND2_9665 ( R1222_U392 , U3482 , R1222_U46 );
nand NAND2_9666 ( R1222_U393 , R1222_U392 , R1222_U391 );
nand NAND2_9667 ( R1222_U394 , R1222_U156 , R1222_U349 );
nand NAND2_9668 ( R1222_U395 , R1222_U374 , R1222_U393 );
nand NAND2_9669 ( R1222_U396 , U3067 , R1222_U30 );
nand NAND2_9670 ( R1222_U397 , U3480 , R1222_U28 );
nand NAND2_9671 ( R1222_U398 , U3068 , R1222_U26 );
nand NAND2_9672 ( R1222_U399 , U3478 , R1222_U27 );
nand NAND2_9673 ( R1222_U400 , R1222_U399 , R1222_U398 );
nand NAND2_9674 ( R1222_U401 , R1222_U350 , R1222_U50 );
nand NAND2_9675 ( R1222_U402 , R1222_U400 , R1222_U202 );
nand NAND2_9676 ( R1222_U403 , U3064 , R1222_U39 );
nand NAND2_9677 ( R1222_U404 , U3476 , R1222_U37 );
nand NAND2_9678 ( R1222_U405 , U3057 , R1222_U35 );
nand NAND2_9679 ( R1222_U406 , U3474 , R1222_U36 );
nand NAND2_9680 ( R1222_U407 , R1222_U406 , R1222_U405 );
nand NAND2_9681 ( R1222_U408 , R1222_U351 , R1222_U51 );
nand NAND2_9682 ( R1222_U409 , R1222_U407 , R1222_U223 );
nand NAND2_9683 ( R1222_U410 , U3061 , R1222_U33 );
nand NAND2_9684 ( R1222_U411 , U3472 , R1222_U34 );
nand NAND2_9685 ( R1222_U412 , R1222_U411 , R1222_U410 );
nand NAND2_9686 ( R1222_U413 , R1222_U352 , R1222_U157 );
nand NAND2_9687 ( R1222_U414 , R1222_U232 , R1222_U412 );
nand NAND2_9688 ( R1222_U415 , U3065 , R1222_U31 );
nand NAND2_9689 ( R1222_U416 , U3470 , R1222_U32 );
nand NAND2_9690 ( R1222_U417 , U3052 , R1222_U159 );
nand NAND2_9691 ( R1222_U418 , U4040 , R1222_U158 );
nand NAND2_9692 ( R1222_U419 , U3052 , R1222_U159 );
nand NAND2_9693 ( R1222_U420 , U4040 , R1222_U158 );
nand NAND2_9694 ( R1222_U421 , R1222_U420 , R1222_U419 );
nand NAND2_9695 ( R1222_U422 , R1222_U160 , R1222_U161 );
nand NAND2_9696 ( R1222_U423 , R1222_U304 , R1222_U421 );
nand NAND2_9697 ( R1222_U424 , U3051 , R1222_U96 );
nand NAND2_9698 ( R1222_U425 , U4029 , R1222_U95 );
nand NAND2_9699 ( R1222_U426 , U3051 , R1222_U96 );
nand NAND2_9700 ( R1222_U427 , U4029 , R1222_U95 );
nand NAND2_9701 ( R1222_U428 , R1222_U427 , R1222_U426 );
nand NAND2_9702 ( R1222_U429 , R1222_U162 , R1222_U163 );
nand NAND2_9703 ( R1222_U430 , R1222_U302 , R1222_U428 );
nand NAND2_9704 ( R1222_U431 , U3050 , R1222_U93 );
nand NAND2_9705 ( R1222_U432 , U4030 , R1222_U94 );
nand NAND2_9706 ( R1222_U433 , U3050 , R1222_U93 );
nand NAND2_9707 ( R1222_U434 , U4030 , R1222_U94 );
nand NAND2_9708 ( R1222_U435 , R1222_U434 , R1222_U433 );
nand NAND2_9709 ( R1222_U436 , R1222_U164 , R1222_U165 );
nand NAND2_9710 ( R1222_U437 , R1222_U298 , R1222_U435 );
nand NAND2_9711 ( R1222_U438 , U3054 , R1222_U91 );
nand NAND2_9712 ( R1222_U439 , U4031 , R1222_U92 );
nand NAND2_9713 ( R1222_U440 , U3055 , R1222_U86 );
nand NAND2_9714 ( R1222_U441 , U4032 , R1222_U87 );
nand NAND2_9715 ( R1222_U442 , R1222_U441 , R1222_U440 );
nand NAND2_9716 ( R1222_U443 , R1222_U353 , R1222_U97 );
nand NAND2_9717 ( R1222_U444 , R1222_U442 , R1222_U306 );
nand NAND2_9718 ( R1222_U445 , U3062 , R1222_U88 );
nand NAND2_9719 ( R1222_U446 , U4033 , R1222_U89 );
nand NAND2_9720 ( R1222_U447 , R1222_U446 , R1222_U445 );
nand NAND2_9721 ( R1222_U448 , R1222_U354 , R1222_U166 );
nand NAND2_9722 ( R1222_U449 , R1222_U288 , R1222_U447 );
nand NAND2_9723 ( R1222_U450 , U3063 , R1222_U84 );
nand NAND2_9724 ( R1222_U451 , U4034 , R1222_U85 );
nand NAND2_9725 ( R1222_U452 , U3063 , R1222_U84 );
nand NAND2_9726 ( R1222_U453 , U4034 , R1222_U85 );
nand NAND2_9727 ( R1222_U454 , R1222_U453 , R1222_U452 );
nand NAND2_9728 ( R1222_U455 , R1222_U167 , R1222_U168 );
nand NAND2_9729 ( R1222_U456 , R1222_U284 , R1222_U454 );
nand NAND2_9730 ( R1222_U457 , U3058 , R1222_U82 );
nand NAND2_9731 ( R1222_U458 , U4035 , R1222_U83 );
nand NAND2_9732 ( R1222_U459 , U3058 , R1222_U82 );
nand NAND2_9733 ( R1222_U460 , U4035 , R1222_U83 );
nand NAND2_9734 ( R1222_U461 , R1222_U460 , R1222_U459 );
nand NAND2_9735 ( R1222_U462 , R1222_U169 , R1222_U170 );
nand NAND2_9736 ( R1222_U463 , R1222_U385 , R1222_U461 );
nand NAND2_9737 ( R1222_U464 , U3072 , R1222_U60 );
nand NAND2_9738 ( R1222_U465 , U4036 , R1222_U61 );
nand NAND2_9739 ( R1222_U466 , U3072 , R1222_U60 );
nand NAND2_9740 ( R1222_U467 , U4036 , R1222_U61 );
nand NAND2_9741 ( R1222_U468 , R1222_U467 , R1222_U466 );
nand NAND2_9742 ( R1222_U469 , U3073 , R1222_U56 );
nand NAND2_9743 ( R1222_U470 , U4037 , R1222_U99 );
nand NAND2_9744 ( R1222_U471 , R1222_U193 , R1222_U173 );
nand NAND2_9745 ( R1222_U472 , R1222_U327 , R1222_U172 );
nand NAND2_9746 ( R1222_U473 , U3078 , R1222_U53 );
nand NAND2_9747 ( R1222_U474 , U3504 , R1222_U54 );
nand NAND2_9748 ( R1222_U475 , R1222_U474 , R1222_U473 );
nand NAND2_9749 ( R1222_U476 , R1222_U355 , R1222_U100 );
nand NAND2_9750 ( R1222_U477 , R1222_U475 , R1222_U315 );
nand NAND2_9751 ( R1222_U478 , U3079 , R1222_U57 );
nand NAND2_9752 ( R1222_U479 , U3502 , R1222_U58 );
nand NAND2_9753 ( R1222_U480 , R1222_U479 , R1222_U478 );
nand NAND2_9754 ( R1222_U481 , R1222_U174 , R1222_U356 );
nand NAND2_9755 ( R1222_U482 , R1222_U381 , R1222_U480 );
nand NAND2_9756 ( R1222_U483 , U3066 , R1222_U66 );
nand NAND2_9757 ( R1222_U484 , U3500 , R1222_U64 );
nand NAND2_9758 ( R1222_U485 , U3070 , R1222_U62 );
nand NAND2_9759 ( R1222_U486 , U3498 , R1222_U63 );
nand NAND2_9760 ( R1222_U487 , R1222_U486 , R1222_U485 );
nand NAND2_9761 ( R1222_U488 , R1222_U357 , R1222_U101 );
nand NAND2_9762 ( R1222_U489 , R1222_U487 , R1222_U260 );
nand NAND2_9763 ( R1222_U490 , U3071 , R1222_U67 );
nand NAND2_9764 ( R1222_U491 , U3496 , R1222_U68 );
nand NAND2_9765 ( R1222_U492 , U3071 , R1222_U67 );
nand NAND2_9766 ( R1222_U493 , U3496 , R1222_U68 );
nand NAND2_9767 ( R1222_U494 , R1222_U493 , R1222_U492 );

// 54 Additional buffers.
buf add_BUF1_1 ( ADDR_REG_19_ , ADDR_REG_19__EXTRA );
buf add_BUF1_2 ( ADDR_REG_18_ , ADDR_REG_18__EXTRA );
buf add_BUF1_3 ( ADDR_REG_17_ , ADDR_REG_17__EXTRA );
buf add_BUF1_4 ( ADDR_REG_16_ , ADDR_REG_16__EXTRA );
buf add_BUF1_5 ( ADDR_REG_15_ , ADDR_REG_15__EXTRA );
buf add_BUF1_6 ( ADDR_REG_14_ , ADDR_REG_14__EXTRA );
buf add_BUF1_7 ( ADDR_REG_13_ , ADDR_REG_13__EXTRA );
buf add_BUF1_8 ( ADDR_REG_12_ , ADDR_REG_12__EXTRA );
buf add_BUF1_9 ( ADDR_REG_11_ , ADDR_REG_11__EXTRA );
buf add_BUF1_10 ( ADDR_REG_10_ , ADDR_REG_10__EXTRA );
buf add_BUF1_11 ( ADDR_REG_9_ , ADDR_REG_9__EXTRA );
buf add_BUF1_12 ( ADDR_REG_8_ , ADDR_REG_8__EXTRA );
buf add_BUF1_13 ( ADDR_REG_7_ , ADDR_REG_7__EXTRA );
buf add_BUF1_14 ( ADDR_REG_6_ , ADDR_REG_6__EXTRA );
buf add_BUF1_15 ( ADDR_REG_5_ , ADDR_REG_5__EXTRA );
buf add_BUF1_16 ( ADDR_REG_4_ , ADDR_REG_4__EXTRA );
buf add_BUF1_17 ( ADDR_REG_3_ , ADDR_REG_3__EXTRA );
buf add_BUF1_18 ( ADDR_REG_2_ , ADDR_REG_2__EXTRA );
buf add_BUF1_19 ( ADDR_REG_1_ , ADDR_REG_1__EXTRA );
buf add_BUF1_20 ( ADDR_REG_0_ , ADDR_REG_0__EXTRA );
buf add_BUF1_21 ( DATAO_REG_0_ , DATAO_REG_0__EXTRA );
buf add_BUF1_22 ( DATAO_REG_1_ , DATAO_REG_1__EXTRA );
buf add_BUF1_23 ( DATAO_REG_2_ , DATAO_REG_2__EXTRA );
buf add_BUF1_24 ( DATAO_REG_3_ , DATAO_REG_3__EXTRA );
buf add_BUF1_25 ( DATAO_REG_4_ , DATAO_REG_4__EXTRA );
buf add_BUF1_26 ( DATAO_REG_5_ , DATAO_REG_5__EXTRA );
buf add_BUF1_27 ( DATAO_REG_6_ , DATAO_REG_6__EXTRA );
buf add_BUF1_28 ( DATAO_REG_7_ , DATAO_REG_7__EXTRA );
buf add_BUF1_29 ( DATAO_REG_8_ , DATAO_REG_8__EXTRA );
buf add_BUF1_30 ( DATAO_REG_9_ , DATAO_REG_9__EXTRA );
buf add_BUF1_31 ( DATAO_REG_10_ , DATAO_REG_10__EXTRA );
buf add_BUF1_32 ( DATAO_REG_11_ , DATAO_REG_11__EXTRA );
buf add_BUF1_33 ( DATAO_REG_12_ , DATAO_REG_12__EXTRA );
buf add_BUF1_34 ( DATAO_REG_13_ , DATAO_REG_13__EXTRA );
buf add_BUF1_35 ( DATAO_REG_14_ , DATAO_REG_14__EXTRA );
buf add_BUF1_36 ( DATAO_REG_15_ , DATAO_REG_15__EXTRA );
buf add_BUF1_37 ( DATAO_REG_16_ , DATAO_REG_16__EXTRA );
buf add_BUF1_38 ( DATAO_REG_17_ , DATAO_REG_17__EXTRA );
buf add_BUF1_39 ( DATAO_REG_18_ , DATAO_REG_18__EXTRA );
buf add_BUF1_40 ( DATAO_REG_19_ , DATAO_REG_19__EXTRA );
buf add_BUF1_41 ( DATAO_REG_20_ , DATAO_REG_20__EXTRA );
buf add_BUF1_42 ( DATAO_REG_21_ , DATAO_REG_21__EXTRA );
buf add_BUF1_43 ( DATAO_REG_22_ , DATAO_REG_22__EXTRA );
buf add_BUF1_44 ( DATAO_REG_23_ , DATAO_REG_23__EXTRA );
buf add_BUF1_45 ( DATAO_REG_24_ , DATAO_REG_24__EXTRA );
buf add_BUF1_46 ( DATAO_REG_25_ , DATAO_REG_25__EXTRA );
buf add_BUF1_47 ( DATAO_REG_26_ , DATAO_REG_26__EXTRA );
buf add_BUF1_48 ( DATAO_REG_27_ , DATAO_REG_27__EXTRA );
buf add_BUF1_49 ( DATAO_REG_28_ , DATAO_REG_28__EXTRA );
buf add_BUF1_50 ( DATAO_REG_29_ , DATAO_REG_29__EXTRA );
buf add_BUF1_51 ( DATAO_REG_30_ , DATAO_REG_30__EXTRA );
buf add_BUF1_52 ( DATAO_REG_31_ , DATAO_REG_31__EXTRA );
buf add_BUF1_53 ( RD_REG , RD_REG_EXTRA );
buf add_BUF1_54 ( WR_REG , WR_REG_EXTRA );

endmodule
