`timescale 1ns/10ps

`define cycle 10.0
`define terminate_cycle 400000//200000 // Modify your terminate ycle here

module b21_ras_testfixture;

`define in_file "b21_ras/rand_input_vector_b21_ras_0.out"
`define out_file "b21_ras/rand_output_vector_b21_ras_0.out"

parameter vec_width = 522;
parameter vec_length = 1;

reg clk = 0;


reg [vec_width-1:0] input_vec_mem [0:vec_length-1];
reg [vec_width-1:0] vec;

wire add_1071_u4, add_1071_u55, add_1071_u56, add_1071_u57, add_1071_u58, add_1071_u59, add_1071_u60, add_1071_u61, add_1071_u62, add_1071_u63, add_1071_u47, add_1071_u48, add_1071_u49, add_1071_u50, add_1071_u51, add_1071_u52, add_1071_u53, add_1071_u54, add_1071_u5, add_1071_u46, u126, u123, p1_u3353, p1_u3352, p1_u3351, p1_u3350, p1_u3349, p1_u3348, p1_u3347, p1_u3346, p1_u3345, p1_u3344, p1_u3343, p1_u3342, p1_u3341, p1_u3340, p1_u3339, p1_u3338, p1_u3337, p1_u3336, p1_u3335, p1_u3334, p1_u3333, p1_u3332, p1_u3331, p1_u3330, p1_u3329, p1_u3328, p1_u3327, p1_u3326, p1_u3325, p1_u3324, p1_u3323, p1_u3322, p1_u3440, p1_u3441, p1_u3321, p1_u3320, p1_u3319, p1_u3318, p1_u3317, p1_u3316, p1_u3315, p1_u3314, p1_u3313, p1_u3312, p1_u3311, p1_u3310, p1_u3309, p1_u3308, p1_u3307, p1_u3306, p1_u3305, p1_u3304, p1_u3303, p1_u3302, p1_u3301, p1_u3300, p1_u3299, p1_u3298, p1_u3297, p1_u3296, p1_u3295, p1_u3294, p1_u3293, p1_u3292, p1_u3454, p1_u3457, p1_u3460, p1_u3463, p1_u3466, p1_u3469, p1_u3472, p1_u3475, p1_u3478, p1_u3481, p1_u3484, p1_u3487, p1_u3490, p1_u3493, p1_u3496, p1_u3499, p1_u3502, p1_u3505, p1_u3508, p1_u3510, p1_u3511, p1_u3512, p1_u3513, p1_u3514, p1_u3515, p1_u3516, p1_u3517, p1_u3518, p1_u3519, p1_u3520, p1_u3521, p1_u3522, p1_u3523, p1_u3524, p1_u3525, p1_u3526, p1_u3527, p1_u3528, p1_u3529, p1_u3530, p1_u3531, p1_u3532, p1_u3533, p1_u3534, p1_u3535, p1_u3536, p1_u3537, p1_u3538, p1_u3539, p1_u3540, p1_u3541, p1_u3542, p1_u3543, p1_u3544, p1_u3545, p1_u3546, p1_u3547, p1_u3548, p1_u3549, p1_u3550, p1_u3551, p1_u3552, p1_u3553, p1_u3554, p1_u3291, p1_u3290, p1_u3289, p1_u3288, p1_u3287, p1_u3286, p1_u3285, p1_u3284, p1_u3283, p1_u3282, p1_u3281, p1_u3280, p1_u3279, p1_u3278, p1_u3277, p1_u3276, p1_u3275, p1_u3274, p1_u3273, p1_u3272, p1_u3271, p1_u3270, p1_u3269, p1_u3268, p1_u3267, p1_u3266, p1_u3265, p1_u3264, p1_u3263, p1_u3355, p1_u3262, p1_u3261, p1_u3260, p1_u3259, p1_u3258, p1_u3257, p1_u3256, p1_u3255, p1_u3254, p1_u3253, p1_u3252, p1_u3251, p1_u3250, p1_u3249, p1_u3248, p1_u3247, p1_u3246, p1_u3245, p1_u3244, p1_u3243, p1_u3242, p1_u3241, p1_u3555, p1_u3556, p1_u3557, p1_u3558, p1_u3559, p1_u3560, p1_u3561, p1_u3562, p1_u3563, p1_u3564, p1_u3565, p1_u3566, p1_u3567, p1_u3568, p1_u3569, p1_u3570, p1_u3571, p1_u3572, p1_u3573, p1_u3574, p1_u3575, p1_u3576, p1_u3577, p1_u3578, p1_u3579, p1_u3580, p1_u3581, p1_u3582, p1_u3583, p1_u3584, p1_u3585, p1_u3586, p1_u3240, p1_u3239, p1_u3238, p1_u3237, p1_u3236, p1_u3235, p1_u3234, p1_u3233, p1_u3232, p1_u3231, p1_u3230, p1_u3229, p1_u3228, p1_u3227, p1_u3226, p1_u3225, p1_u3224, p1_u3223, p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218, p1_u3217, p1_u3216, p1_u3215, p1_u3214, p1_u3213, p1_u3212, p1_u3211, p1_u3084, p1_u3083, p1_u4006, p2_u3358, p2_u3357, p2_u3356, p2_u3355, p2_u3354, p2_u3353, p2_u3352, p2_u3351, p2_u3350, p2_u3349, p2_u3348, p2_u3347, p2_u3346, p2_u3345, p2_u3344, p2_u3343, p2_u3342, p2_u3341, p2_u3340, p2_u3339, p2_u3338, p2_u3337, p2_u3336, p2_u3335, p2_u3334, p2_u3333, p2_u3332, p2_u3331, p2_u3330, p2_u3329, p2_u3328, p2_u3327, p2_u3437, p2_u3438, p2_u3326, p2_u3325, p2_u3324, p2_u3323, p2_u3322, p2_u3321, p2_u3320, p2_u3319, p2_u3318, p2_u3317, p2_u3316, p2_u3315, p2_u3314, p2_u3313, p2_u3312, p2_u3311, p2_u3310, p2_u3309, p2_u3308, p2_u3307, p2_u3306, p2_u3305, p2_u3304, p2_u3303, p2_u3302, p2_u3301, p2_u3300, p2_u3299, p2_u3298, p2_u3297, p2_u3451, p2_u3454, p2_u3457, p2_u3460, p2_u3463, p2_u3466, p2_u3469, p2_u3472, p2_u3475, p2_u3478, p2_u3481, p2_u3484, p2_u3487, p2_u3490, p2_u3493, p2_u3496, p2_u3499, p2_u3502, p2_u3505, p2_u3507, p2_u3508, p2_u3509, p2_u3510, p2_u3511, p2_u3512, p2_u3513, p2_u3514, p2_u3515, p2_u3516, p2_u3517, p2_u3518, p2_u3519, p2_u3520, p2_u3521, p2_u3522, p2_u3523, p2_u3524, p2_u3525, p2_u3526, p2_u3527, p2_u3528, p2_u3529, p2_u3530, p2_u3531, p2_u3532, p2_u3533, p2_u3534, p2_u3535, p2_u3536, p2_u3537, p2_u3538, p2_u3539, p2_u3540, p2_u3541, p2_u3542, p2_u3543, p2_u3544, p2_u3545, p2_u3546, p2_u3547, p2_u3548, p2_u3549, p2_u3550, p2_u3551, p2_u3296, p2_u3295, p2_u3294, p2_u3293, p2_u3292, p2_u3291, p2_u3290, p2_u3289, p2_u3288, p2_u3287, p2_u3286, p2_u3285, p2_u3284, p2_u3283, p2_u3282, p2_u3281, p2_u3280, p2_u3279, p2_u3278, p2_u3277, p2_u3276, p2_u3275, p2_u3274, p2_u3273, p2_u3272, p2_u3271, p2_u3270, p2_u3269, p2_u3268, p2_u3267, p2_u3266, p2_u3265, p2_u3264, p2_u3263, p2_u3262, p2_u3261, p2_u3260, p2_u3259, p2_u3258, p2_u3257, p2_u3256, p2_u3255, p2_u3254, p2_u3253, p2_u3252, p2_u3251, p2_u3250, p2_u3249, p2_u3248, p2_u3247, p2_u3246, p2_u3245, p2_u3552, p2_u3553, p2_u3554, p2_u3555, p2_u3556, p2_u3557, p2_u3558, p2_u3559, p2_u3560, p2_u3561, p2_u3562, p2_u3563, p2_u3564, p2_u3565, p2_u3566, p2_u3567, p2_u3568, p2_u3569, p2_u3570, p2_u3571, p2_u3572, p2_u3573, p2_u3574, p2_u3575, p2_u3576, p2_u3577, p2_u3578, p2_u3579, p2_u3580, p2_u3581, p2_u3582, p2_u3583, p2_u3244, p2_u3243, p2_u3242, p2_u3241, p2_u3240, p2_u3239, p2_u3238, p2_u3237, p2_u3236, p2_u3235, p2_u3234, p2_u3233, p2_u3232, p2_u3231, p2_u3230, p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225, p2_u3224, p2_u3223, p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218, p2_u3217, p2_u3216, p2_u3215, p2_u3152, p2_u3151, p2_u3966;
initial begin
	$readmemb(`in_file, input_vec_mem );
end

always #(`cycle/2) clk = ~clk;

b21_ras cc (.SI_31_(vec[521]), .SI_30_(vec[520]), .SI_29_(vec[519]), .SI_28_(vec[518]), .SI_27_(vec[517]), .SI_26_(vec[516]), .SI_25_(vec[515]), .SI_24_(vec[514]), .SI_23_(vec[513]), .SI_22_(vec[512]), .SI_21_(vec[511]), .SI_20_(vec[510]), .SI_19_(vec[509]), .SI_18_(vec[508]), .SI_17_(vec[507]), .SI_16_(vec[506]), .SI_15_(vec[505]), .SI_14_(vec[504]), .SI_13_(vec[503]), .SI_12_(vec[502]), .SI_11_(vec[501]), .SI_10_(vec[500]), .SI_9_(vec[499]), .SI_8_(vec[498]), .SI_7_(vec[497]), .SI_6_(vec[496]), .SI_5_(vec[495]), .SI_4_(vec[494]), .SI_3_(vec[493]), .SI_2_(vec[492]), .SI_1_(vec[491]), .SI_0_(vec[490]), .P1_IR_REG_0_(vec[489]), .P1_IR_REG_1_(vec[488]), .P1_IR_REG_2_(vec[487]), .P1_IR_REG_3_(vec[486]), .P1_IR_REG_4_(vec[485]), .P1_IR_REG_5_(vec[484]), .P1_IR_REG_6_(vec[483]), .P1_IR_REG_7_(vec[482]), .P1_IR_REG_8_(vec[481]), .P1_IR_REG_9_(vec[480]), .P1_IR_REG_10_(vec[479]), .P1_IR_REG_11_(vec[478]), .P1_IR_REG_12_(vec[477]), .P1_IR_REG_13_(vec[476]), .P1_IR_REG_14_(vec[475]), .P1_IR_REG_15_(vec[474]), .P1_IR_REG_16_(vec[473]), .P1_IR_REG_17_(vec[472]), .P1_IR_REG_18_(vec[471]), .P1_IR_REG_19_(vec[470]), .P1_IR_REG_20_(vec[469]), .P1_IR_REG_21_(vec[468]), .P1_IR_REG_22_(vec[467]), .P1_IR_REG_23_(vec[466]), .P1_IR_REG_24_(vec[465]), .P1_IR_REG_25_(vec[464]), .P1_IR_REG_26_(vec[463]), .P1_IR_REG_27_(vec[462]), .P1_IR_REG_28_(vec[461]), .P1_IR_REG_29_(vec[460]), .P1_IR_REG_30_(vec[459]), .P1_IR_REG_31_(vec[458]), .P1_D_REG_0_(vec[457]), .P1_D_REG_1_(vec[456]), .P1_D_REG_2_(vec[455]), .P1_D_REG_3_(vec[454]), .P1_D_REG_4_(vec[453]), .P1_D_REG_5_(vec[452]), .P1_D_REG_6_(vec[451]), .P1_D_REG_7_(vec[450]), .P1_D_REG_8_(vec[449]), .P1_D_REG_9_(vec[448]), .P1_D_REG_10_(vec[447]), .P1_D_REG_11_(vec[446]), .P1_D_REG_12_(vec[445]), .P1_D_REG_13_(vec[444]), .P1_D_REG_14_(vec[443]), .P1_D_REG_15_(vec[442]), .P1_D_REG_16_(vec[441]), .P1_D_REG_17_(vec[440]), .P1_D_REG_18_(vec[439]), .P1_D_REG_19_(vec[438]), .P1_D_REG_20_(vec[437]), .P1_D_REG_21_(vec[436]), .P1_D_REG_22_(vec[435]), .P1_D_REG_23_(vec[434]), .P1_D_REG_24_(vec[433]), .P1_D_REG_25_(vec[432]), .P1_D_REG_26_(vec[431]), .P1_D_REG_27_(vec[430]), .P1_D_REG_28_(vec[429]), .P1_D_REG_29_(vec[428]), .P1_D_REG_30_(vec[427]), .P1_D_REG_31_(vec[426]), .P1_REG0_REG_0_(vec[425]), .P1_REG0_REG_1_(vec[424]), .P1_REG0_REG_2_(vec[423]), .P1_REG0_REG_3_(vec[422]), .P1_REG0_REG_4_(vec[421]), .P1_REG0_REG_5_(vec[420]), .P1_REG0_REG_6_(vec[419]), .P1_REG0_REG_7_(vec[418]), .P1_REG0_REG_8_(vec[417]), .P1_REG0_REG_9_(vec[416]), .P1_REG0_REG_10_(vec[415]), .P1_REG0_REG_11_(vec[414]), .P1_REG0_REG_12_(vec[413]), .P1_REG0_REG_13_(vec[412]), .P1_REG0_REG_14_(vec[411]), .P1_REG0_REG_15_(vec[410]), .P1_REG0_REG_16_(vec[409]), .P1_REG0_REG_17_(vec[408]), .P1_REG0_REG_18_(vec[407]), .P1_REG0_REG_19_(vec[406]), .P1_REG0_REG_20_(vec[405]), .P1_REG0_REG_21_(vec[404]), .P1_REG0_REG_22_(vec[403]), .P1_REG0_REG_23_(vec[402]), .P1_REG0_REG_24_(vec[401]), .P1_REG0_REG_25_(vec[400]), .P1_REG0_REG_26_(vec[399]), .P1_REG0_REG_27_(vec[398]), .P1_REG0_REG_28_(vec[397]), .P1_REG0_REG_29_(vec[396]), .P1_REG0_REG_30_(vec[395]), .P1_REG0_REG_31_(vec[394]), .P1_REG1_REG_0_(vec[393]), .P1_REG1_REG_1_(vec[392]), .P1_REG1_REG_2_(vec[391]), .P1_REG1_REG_3_(vec[390]), .P1_REG1_REG_4_(vec[389]), .P1_REG1_REG_5_(vec[388]), .P1_REG1_REG_6_(vec[387]), .P1_REG1_REG_7_(vec[386]), .P1_REG1_REG_8_(vec[385]), .P1_REG1_REG_9_(vec[384]), .P1_REG1_REG_10_(vec[383]), .P1_REG1_REG_11_(vec[382]), .P1_REG1_REG_12_(vec[381]), .P1_REG1_REG_13_(vec[380]), .P1_REG1_REG_14_(vec[379]), .P1_REG1_REG_15_(vec[378]), .P1_REG1_REG_16_(vec[377]), .P1_REG1_REG_17_(vec[376]), .P1_REG1_REG_18_(vec[375]), .P1_REG1_REG_19_(vec[374]), .P1_REG1_REG_20_(vec[373]), .P1_REG1_REG_21_(vec[372]), .P1_REG1_REG_22_(vec[371]), .P1_REG1_REG_23_(vec[370]), .P1_REG1_REG_24_(vec[369]), .P1_REG1_REG_25_(vec[368]), .P1_REG1_REG_26_(vec[367]), .P1_REG1_REG_27_(vec[366]), .P1_REG1_REG_28_(vec[365]), .P1_REG1_REG_29_(vec[364]), .P1_REG1_REG_30_(vec[363]), .P1_REG1_REG_31_(vec[362]), .P1_REG2_REG_0_(vec[361]), .P1_REG2_REG_1_(vec[360]), .P1_REG2_REG_2_(vec[359]), .P1_REG2_REG_3_(vec[358]), .P1_REG2_REG_4_(vec[357]), .P1_REG2_REG_5_(vec[356]), .P1_REG2_REG_6_(vec[355]), .P1_REG2_REG_7_(vec[354]), .P1_REG2_REG_8_(vec[353]), .P1_REG2_REG_9_(vec[352]), .P1_REG2_REG_10_(vec[351]), .P1_REG2_REG_11_(vec[350]), .P1_REG2_REG_12_(vec[349]), .P1_REG2_REG_13_(vec[348]), .P1_REG2_REG_14_(vec[347]), .P1_REG2_REG_15_(vec[346]), .P1_REG2_REG_16_(vec[345]), .P1_REG2_REG_17_(vec[344]), .P1_REG2_REG_18_(vec[343]), .P1_REG2_REG_19_(vec[342]), .P1_REG2_REG_20_(vec[341]), .P1_REG2_REG_21_(vec[340]), .P1_REG2_REG_22_(vec[339]), .P1_REG2_REG_23_(vec[338]), .P1_REG2_REG_24_(vec[337]), .P1_REG2_REG_25_(vec[336]), .P1_REG2_REG_26_(vec[335]), .P1_REG2_REG_27_(vec[334]), .P1_REG2_REG_28_(vec[333]), .P1_REG2_REG_29_(vec[332]), .P1_REG2_REG_30_(vec[331]), .P1_REG2_REG_31_(vec[330]), .P1_ADDR_REG_19_(vec[329]), .P1_ADDR_REG_18_(vec[328]), .P1_ADDR_REG_17_(vec[327]), .P1_ADDR_REG_16_(vec[326]), .P1_ADDR_REG_15_(vec[325]), .P1_ADDR_REG_14_(vec[324]), .P1_ADDR_REG_13_(vec[323]), .P1_ADDR_REG_12_(vec[322]), .P1_ADDR_REG_11_(vec[321]), .P1_ADDR_REG_10_(vec[320]), .P1_ADDR_REG_9_(vec[319]), .P1_ADDR_REG_8_(vec[318]), .P1_ADDR_REG_7_(vec[317]), .P1_ADDR_REG_6_(vec[316]), .P1_ADDR_REG_5_(vec[315]), .P1_ADDR_REG_4_(vec[314]), .P1_ADDR_REG_3_(vec[313]), .P1_ADDR_REG_2_(vec[312]), .P1_ADDR_REG_1_(vec[311]), .P1_ADDR_REG_0_(vec[310]), .P1_DATAO_REG_0_(vec[309]), .P1_DATAO_REG_1_(vec[308]), .P1_DATAO_REG_2_(vec[307]), .P1_DATAO_REG_3_(vec[306]), .P1_DATAO_REG_4_(vec[305]), .P1_DATAO_REG_5_(vec[304]), .P1_DATAO_REG_6_(vec[303]), .P1_DATAO_REG_7_(vec[302]), .P1_DATAO_REG_8_(vec[301]), .P1_DATAO_REG_9_(vec[300]), .P1_DATAO_REG_10_(vec[299]), .P1_DATAO_REG_11_(vec[298]), .P1_DATAO_REG_12_(vec[297]), .P1_DATAO_REG_13_(vec[296]), .P1_DATAO_REG_14_(vec[295]), .P1_DATAO_REG_15_(vec[294]), .P1_DATAO_REG_16_(vec[293]), .P1_DATAO_REG_17_(vec[292]), .P1_DATAO_REG_18_(vec[291]), .P1_DATAO_REG_19_(vec[290]), .P1_DATAO_REG_20_(vec[289]), .P1_DATAO_REG_21_(vec[288]), .P1_DATAO_REG_22_(vec[287]), .P1_DATAO_REG_23_(vec[286]), .P1_DATAO_REG_24_(vec[285]), .P1_DATAO_REG_25_(vec[284]), .P1_DATAO_REG_26_(vec[283]), .P1_DATAO_REG_27_(vec[282]), .P1_DATAO_REG_28_(vec[281]), .P1_DATAO_REG_29_(vec[280]), .P1_DATAO_REG_30_(vec[279]), .P1_DATAO_REG_31_(vec[278]), .P1_B_REG(vec[277]), .P1_REG3_REG_15_(vec[276]), .P1_REG3_REG_26_(vec[275]), .P1_REG3_REG_6_(vec[274]), .P1_REG3_REG_18_(vec[273]), .P1_REG3_REG_2_(vec[272]), .P1_REG3_REG_11_(vec[271]), .P1_REG3_REG_22_(vec[270]), .P1_REG3_REG_13_(vec[269]), .P1_REG3_REG_20_(vec[268]), .P1_REG3_REG_0_(vec[267]), .P1_REG3_REG_9_(vec[266]), .P1_REG3_REG_4_(vec[265]), .P1_REG3_REG_24_(vec[264]), .P1_REG3_REG_17_(vec[263]), .P1_REG3_REG_5_(vec[262]), .P1_REG3_REG_16_(vec[261]), .P1_REG3_REG_25_(vec[260]), .P1_REG3_REG_12_(vec[259]), .P1_REG3_REG_21_(vec[258]), .P1_REG3_REG_1_(vec[257]), .P1_REG3_REG_8_(vec[256]), .P1_REG3_REG_28_(vec[255]), .P1_REG3_REG_19_(vec[254]), .P1_REG3_REG_3_(vec[253]), .P1_REG3_REG_10_(vec[252]), .P1_REG3_REG_23_(vec[251]), .P1_REG3_REG_14_(vec[250]), .P1_REG3_REG_27_(vec[249]), .P1_REG3_REG_7_(vec[248]), .P1_STATE_REG(vec[247]), .P1_RD_REG(vec[246]), .P1_WR_REG(vec[245]), .P2_IR_REG_0_(vec[244]), .P2_IR_REG_1_(vec[243]), .P2_IR_REG_2_(vec[242]), .P2_IR_REG_3_(vec[241]), .P2_IR_REG_4_(vec[240]), .P2_IR_REG_5_(vec[239]), .P2_IR_REG_6_(vec[238]), .P2_IR_REG_7_(vec[237]), .P2_IR_REG_8_(vec[236]), .P2_IR_REG_9_(vec[235]), .P2_IR_REG_10_(vec[234]), .P2_IR_REG_11_(vec[233]), .P2_IR_REG_12_(vec[232]), .P2_IR_REG_13_(vec[231]), .P2_IR_REG_14_(vec[230]), .P2_IR_REG_15_(vec[229]), .P2_IR_REG_16_(vec[228]), .P2_IR_REG_17_(vec[227]), .P2_IR_REG_18_(vec[226]), .P2_IR_REG_19_(vec[225]), .P2_IR_REG_20_(vec[224]), .P2_IR_REG_21_(vec[223]), .P2_IR_REG_22_(vec[222]), .P2_IR_REG_23_(vec[221]), .P2_IR_REG_24_(vec[220]), .P2_IR_REG_25_(vec[219]), .P2_IR_REG_26_(vec[218]), .P2_IR_REG_27_(vec[217]), .P2_IR_REG_28_(vec[216]), .P2_IR_REG_29_(vec[215]), .P2_IR_REG_30_(vec[214]), .P2_IR_REG_31_(vec[213]), .P2_D_REG_0_(vec[212]), .P2_D_REG_1_(vec[211]), .P2_D_REG_2_(vec[210]), .P2_D_REG_3_(vec[209]), .P2_D_REG_4_(vec[208]), .P2_D_REG_5_(vec[207]), .P2_D_REG_6_(vec[206]), .P2_D_REG_7_(vec[205]), .P2_D_REG_8_(vec[204]), .P2_D_REG_9_(vec[203]), .P2_D_REG_10_(vec[202]), .P2_D_REG_11_(vec[201]), .P2_D_REG_12_(vec[200]), .P2_D_REG_13_(vec[199]), .P2_D_REG_14_(vec[198]), .P2_D_REG_15_(vec[197]), .P2_D_REG_16_(vec[196]), .P2_D_REG_17_(vec[195]), .P2_D_REG_18_(vec[194]), .P2_D_REG_19_(vec[193]), .P2_D_REG_20_(vec[192]), .P2_D_REG_21_(vec[191]), .P2_D_REG_22_(vec[190]), .P2_D_REG_23_(vec[189]), .P2_D_REG_24_(vec[188]), .P2_D_REG_25_(vec[187]), .P2_D_REG_26_(vec[186]), .P2_D_REG_27_(vec[185]), .P2_D_REG_28_(vec[184]), .P2_D_REG_29_(vec[183]), .P2_D_REG_30_(vec[182]), .P2_D_REG_31_(vec[181]), .P2_REG0_REG_0_(vec[180]), .P2_REG0_REG_1_(vec[179]), .P2_REG0_REG_2_(vec[178]), .P2_REG0_REG_3_(vec[177]), .P2_REG0_REG_4_(vec[176]), .P2_REG0_REG_5_(vec[175]), .P2_REG0_REG_6_(vec[174]), .P2_REG0_REG_7_(vec[173]), .P2_REG0_REG_8_(vec[172]), .P2_REG0_REG_9_(vec[171]), .P2_REG0_REG_10_(vec[170]), .P2_REG0_REG_11_(vec[169]), .P2_REG0_REG_12_(vec[168]), .P2_REG0_REG_13_(vec[167]), .P2_REG0_REG_14_(vec[166]), .P2_REG0_REG_15_(vec[165]), .P2_REG0_REG_16_(vec[164]), .P2_REG0_REG_17_(vec[163]), .P2_REG0_REG_18_(vec[162]), .P2_REG0_REG_19_(vec[161]), .P2_REG0_REG_20_(vec[160]), .P2_REG0_REG_21_(vec[159]), .P2_REG0_REG_22_(vec[158]), .P2_REG0_REG_23_(vec[157]), .P2_REG0_REG_24_(vec[156]), .P2_REG0_REG_25_(vec[155]), .P2_REG0_REG_26_(vec[154]), .P2_REG0_REG_27_(vec[153]), .P2_REG0_REG_28_(vec[152]), .P2_REG0_REG_29_(vec[151]), .P2_REG0_REG_30_(vec[150]), .P2_REG0_REG_31_(vec[149]), .P2_REG1_REG_0_(vec[148]), .P2_REG1_REG_1_(vec[147]), .P2_REG1_REG_2_(vec[146]), .P2_REG1_REG_3_(vec[145]), .P2_REG1_REG_4_(vec[144]), .P2_REG1_REG_5_(vec[143]), .P2_REG1_REG_6_(vec[142]), .P2_REG1_REG_7_(vec[141]), .P2_REG1_REG_8_(vec[140]), .P2_REG1_REG_9_(vec[139]), .P2_REG1_REG_10_(vec[138]), .P2_REG1_REG_11_(vec[137]), .P2_REG1_REG_12_(vec[136]), .P2_REG1_REG_13_(vec[135]), .P2_REG1_REG_14_(vec[134]), .P2_REG1_REG_15_(vec[133]), .P2_REG1_REG_16_(vec[132]), .P2_REG1_REG_17_(vec[131]), .P2_REG1_REG_18_(vec[130]), .P2_REG1_REG_19_(vec[129]), .P2_REG1_REG_20_(vec[128]), .P2_REG1_REG_21_(vec[127]), .P2_REG1_REG_22_(vec[126]), .P2_REG1_REG_23_(vec[125]), .P2_REG1_REG_24_(vec[124]), .P2_REG1_REG_25_(vec[123]), .P2_REG1_REG_26_(vec[122]), .P2_REG1_REG_27_(vec[121]), .P2_REG1_REG_28_(vec[120]), .P2_REG1_REG_29_(vec[119]), .P2_REG1_REG_30_(vec[118]), .P2_REG1_REG_31_(vec[117]), .P2_REG2_REG_0_(vec[116]), .P2_REG2_REG_1_(vec[115]), .P2_REG2_REG_2_(vec[114]), .P2_REG2_REG_3_(vec[113]), .P2_REG2_REG_4_(vec[112]), .P2_REG2_REG_5_(vec[111]), .P2_REG2_REG_6_(vec[110]), .P2_REG2_REG_7_(vec[109]), .P2_REG2_REG_8_(vec[108]), .P2_REG2_REG_9_(vec[107]), .P2_REG2_REG_10_(vec[106]), .P2_REG2_REG_11_(vec[105]), .P2_REG2_REG_12_(vec[104]), .P2_REG2_REG_13_(vec[103]), .P2_REG2_REG_14_(vec[102]), .P2_REG2_REG_15_(vec[101]), .P2_REG2_REG_16_(vec[100]), .P2_REG2_REG_17_(vec[99]), .P2_REG2_REG_18_(vec[98]), .P2_REG2_REG_19_(vec[97]), .P2_REG2_REG_20_(vec[96]), .P2_REG2_REG_21_(vec[95]), .P2_REG2_REG_22_(vec[94]), .P2_REG2_REG_23_(vec[93]), .P2_REG2_REG_24_(vec[92]), .P2_REG2_REG_25_(vec[91]), .P2_REG2_REG_26_(vec[90]), .P2_REG2_REG_27_(vec[89]), .P2_REG2_REG_28_(vec[88]), .P2_REG2_REG_29_(vec[87]), .P2_REG2_REG_30_(vec[86]), .P2_REG2_REG_31_(vec[85]), .P2_ADDR_REG_19_(vec[84]), .P2_ADDR_REG_18_(vec[83]), .P2_ADDR_REG_17_(vec[82]), .P2_ADDR_REG_16_(vec[81]), .P2_ADDR_REG_15_(vec[80]), .P2_ADDR_REG_14_(vec[79]), .P2_ADDR_REG_13_(vec[78]), .P2_ADDR_REG_12_(vec[77]), .P2_ADDR_REG_11_(vec[76]), .P2_ADDR_REG_10_(vec[75]), .P2_ADDR_REG_9_(vec[74]), .P2_ADDR_REG_8_(vec[73]), .P2_ADDR_REG_7_(vec[72]), .P2_ADDR_REG_6_(vec[71]), .P2_ADDR_REG_5_(vec[70]), .P2_ADDR_REG_4_(vec[69]), .P2_ADDR_REG_3_(vec[68]), .P2_ADDR_REG_2_(vec[67]), .P2_ADDR_REG_1_(vec[66]), .P2_ADDR_REG_0_(vec[65]), .P2_DATAO_REG_0_(vec[64]), .P2_DATAO_REG_1_(vec[63]), .P2_DATAO_REG_2_(vec[62]), .P2_DATAO_REG_3_(vec[61]), .P2_DATAO_REG_4_(vec[60]), .P2_DATAO_REG_5_(vec[59]), .P2_DATAO_REG_6_(vec[58]), .P2_DATAO_REG_7_(vec[57]), .P2_DATAO_REG_8_(vec[56]), .P2_DATAO_REG_9_(vec[55]), .P2_DATAO_REG_10_(vec[54]), .P2_DATAO_REG_11_(vec[53]), .P2_DATAO_REG_12_(vec[52]), .P2_DATAO_REG_13_(vec[51]), .P2_DATAO_REG_14_(vec[50]), .P2_DATAO_REG_15_(vec[49]), .P2_DATAO_REG_16_(vec[48]), .P2_DATAO_REG_17_(vec[47]), .P2_DATAO_REG_18_(vec[46]), .P2_DATAO_REG_19_(vec[45]), .P2_DATAO_REG_20_(vec[44]), .P2_DATAO_REG_21_(vec[43]), .P2_DATAO_REG_22_(vec[42]), .P2_DATAO_REG_23_(vec[41]), .P2_DATAO_REG_24_(vec[40]), .P2_DATAO_REG_25_(vec[39]), .P2_DATAO_REG_26_(vec[38]), .P2_DATAO_REG_27_(vec[37]), .P2_DATAO_REG_28_(vec[36]), .P2_DATAO_REG_29_(vec[35]), .P2_DATAO_REG_30_(vec[34]), .P2_DATAO_REG_31_(vec[33]), .P2_B_REG(vec[32]), .P2_REG3_REG_15_(vec[31]), .P2_REG3_REG_26_(vec[30]), .P2_REG3_REG_6_(vec[29]), .P2_REG3_REG_18_(vec[28]), .P2_REG3_REG_2_(vec[27]), .P2_REG3_REG_11_(vec[26]), .P2_REG3_REG_22_(vec[25]), .P2_REG3_REG_13_(vec[24]), .P2_REG3_REG_20_(vec[23]), .P2_REG3_REG_0_(vec[22]), .P2_REG3_REG_9_(vec[21]), .P2_REG3_REG_4_(vec[20]), .P2_REG3_REG_24_(vec[19]), .P2_REG3_REG_17_(vec[18]), .P2_REG3_REG_5_(vec[17]), .P2_REG3_REG_16_(vec[16]), .P2_REG3_REG_25_(vec[15]), .P2_REG3_REG_12_(vec[14]), .P2_REG3_REG_21_(vec[13]), .P2_REG3_REG_1_(vec[12]), .P2_REG3_REG_8_(vec[11]), .P2_REG3_REG_28_(vec[10]), .P2_REG3_REG_19_(vec[9]), .P2_REG3_REG_3_(vec[8]), .P2_REG3_REG_10_(vec[7]), .P2_REG3_REG_23_(vec[6]), .P2_REG3_REG_14_(vec[5]), .P2_REG3_REG_27_(vec[4]), .P2_REG3_REG_7_(vec[3]), .P2_STATE_REG(vec[2]), .P2_RD_REG(vec[1]), .P2_WR_REG(vec[0]), .ADD_1071_U4(add_1071_u4), .ADD_1071_U55(add_1071_u55), .ADD_1071_U56(add_1071_u56), .ADD_1071_U57(add_1071_u57), .ADD_1071_U58(add_1071_u58), .ADD_1071_U59(add_1071_u59), .ADD_1071_U60(add_1071_u60), .ADD_1071_U61(add_1071_u61), .ADD_1071_U62(add_1071_u62), .ADD_1071_U63(add_1071_u63), .ADD_1071_U47(add_1071_u47), .ADD_1071_U48(add_1071_u48), .ADD_1071_U49(add_1071_u49), .ADD_1071_U50(add_1071_u50), .ADD_1071_U51(add_1071_u51), .ADD_1071_U52(add_1071_u52), .ADD_1071_U53(add_1071_u53), .ADD_1071_U54(add_1071_u54), .ADD_1071_U5(add_1071_u5), .ADD_1071_U46(add_1071_u46), .U126(u126), .U123(u123), .P1_U3353(p1_u3353), .P1_U3352(p1_u3352), .P1_U3351(p1_u3351), .P1_U3350(p1_u3350), .P1_U3349(p1_u3349), .P1_U3348(p1_u3348), .P1_U3347(p1_u3347), .P1_U3346(p1_u3346), .P1_U3345(p1_u3345), .P1_U3344(p1_u3344), .P1_U3343(p1_u3343), .P1_U3342(p1_u3342), .P1_U3341(p1_u3341), .P1_U3340(p1_u3340), .P1_U3339(p1_u3339), .P1_U3338(p1_u3338), .P1_U3337(p1_u3337), .P1_U3336(p1_u3336), .P1_U3335(p1_u3335), .P1_U3334(p1_u3334), .P1_U3333(p1_u3333), .P1_U3332(p1_u3332), .P1_U3331(p1_u3331), .P1_U3330(p1_u3330), .P1_U3329(p1_u3329), .P1_U3328(p1_u3328), .P1_U3327(p1_u3327), .P1_U3326(p1_u3326), .P1_U3325(p1_u3325), .P1_U3324(p1_u3324), .P1_U3323(p1_u3323), .P1_U3322(p1_u3322), .P1_U3440(p1_u3440), .P1_U3441(p1_u3441), .P1_U3321(p1_u3321), .P1_U3320(p1_u3320), .P1_U3319(p1_u3319), .P1_U3318(p1_u3318), .P1_U3317(p1_u3317), .P1_U3316(p1_u3316), .P1_U3315(p1_u3315), .P1_U3314(p1_u3314), .P1_U3313(p1_u3313), .P1_U3312(p1_u3312), .P1_U3311(p1_u3311), .P1_U3310(p1_u3310), .P1_U3309(p1_u3309), .P1_U3308(p1_u3308), .P1_U3307(p1_u3307), .P1_U3306(p1_u3306), .P1_U3305(p1_u3305), .P1_U3304(p1_u3304), .P1_U3303(p1_u3303), .P1_U3302(p1_u3302), .P1_U3301(p1_u3301), .P1_U3300(p1_u3300), .P1_U3299(p1_u3299), .P1_U3298(p1_u3298), .P1_U3297(p1_u3297), .P1_U3296(p1_u3296), .P1_U3295(p1_u3295), .P1_U3294(p1_u3294), .P1_U3293(p1_u3293), .P1_U3292(p1_u3292), .P1_U3454(p1_u3454), .P1_U3457(p1_u3457), .P1_U3460(p1_u3460), .P1_U3463(p1_u3463), .P1_U3466(p1_u3466), .P1_U3469(p1_u3469), .P1_U3472(p1_u3472), .P1_U3475(p1_u3475), .P1_U3478(p1_u3478), .P1_U3481(p1_u3481), .P1_U3484(p1_u3484), .P1_U3487(p1_u3487), .P1_U3490(p1_u3490), .P1_U3493(p1_u3493), .P1_U3496(p1_u3496), .P1_U3499(p1_u3499), .P1_U3502(p1_u3502), .P1_U3505(p1_u3505), .P1_U3508(p1_u3508), .P1_U3510(p1_u3510), .P1_U3511(p1_u3511), .P1_U3512(p1_u3512), .P1_U3513(p1_u3513), .P1_U3514(p1_u3514), .P1_U3515(p1_u3515), .P1_U3516(p1_u3516), .P1_U3517(p1_u3517), .P1_U3518(p1_u3518), .P1_U3519(p1_u3519), .P1_U3520(p1_u3520), .P1_U3521(p1_u3521), .P1_U3522(p1_u3522), .P1_U3523(p1_u3523), .P1_U3524(p1_u3524), .P1_U3525(p1_u3525), .P1_U3526(p1_u3526), .P1_U3527(p1_u3527), .P1_U3528(p1_u3528), .P1_U3529(p1_u3529), .P1_U3530(p1_u3530), .P1_U3531(p1_u3531), .P1_U3532(p1_u3532), .P1_U3533(p1_u3533), .P1_U3534(p1_u3534), .P1_U3535(p1_u3535), .P1_U3536(p1_u3536), .P1_U3537(p1_u3537), .P1_U3538(p1_u3538), .P1_U3539(p1_u3539), .P1_U3540(p1_u3540), .P1_U3541(p1_u3541), .P1_U3542(p1_u3542), .P1_U3543(p1_u3543), .P1_U3544(p1_u3544), .P1_U3545(p1_u3545), .P1_U3546(p1_u3546), .P1_U3547(p1_u3547), .P1_U3548(p1_u3548), .P1_U3549(p1_u3549), .P1_U3550(p1_u3550), .P1_U3551(p1_u3551), .P1_U3552(p1_u3552), .P1_U3553(p1_u3553), .P1_U3554(p1_u3554), .P1_U3291(p1_u3291), .P1_U3290(p1_u3290), .P1_U3289(p1_u3289), .P1_U3288(p1_u3288), .P1_U3287(p1_u3287), .P1_U3286(p1_u3286), .P1_U3285(p1_u3285), .P1_U3284(p1_u3284), .P1_U3283(p1_u3283), .P1_U3282(p1_u3282), .P1_U3281(p1_u3281), .P1_U3280(p1_u3280), .P1_U3279(p1_u3279), .P1_U3278(p1_u3278), .P1_U3277(p1_u3277), .P1_U3276(p1_u3276), .P1_U3275(p1_u3275), .P1_U3274(p1_u3274), .P1_U3273(p1_u3273), .P1_U3272(p1_u3272), .P1_U3271(p1_u3271), .P1_U3270(p1_u3270), .P1_U3269(p1_u3269), .P1_U3268(p1_u3268), .P1_U3267(p1_u3267), .P1_U3266(p1_u3266), .P1_U3265(p1_u3265), .P1_U3264(p1_u3264), .P1_U3263(p1_u3263), .P1_U3355(p1_u3355), .P1_U3262(p1_u3262), .P1_U3261(p1_u3261), .P1_U3260(p1_u3260), .P1_U3259(p1_u3259), .P1_U3258(p1_u3258), .P1_U3257(p1_u3257), .P1_U3256(p1_u3256), .P1_U3255(p1_u3255), .P1_U3254(p1_u3254), .P1_U3253(p1_u3253), .P1_U3252(p1_u3252), .P1_U3251(p1_u3251), .P1_U3250(p1_u3250), .P1_U3249(p1_u3249), .P1_U3248(p1_u3248), .P1_U3247(p1_u3247), .P1_U3246(p1_u3246), .P1_U3245(p1_u3245), .P1_U3244(p1_u3244), .P1_U3243(p1_u3243), .P1_U3242(p1_u3242), .P1_U3241(p1_u3241), .P1_U3555(p1_u3555), .P1_U3556(p1_u3556), .P1_U3557(p1_u3557), .P1_U3558(p1_u3558), .P1_U3559(p1_u3559), .P1_U3560(p1_u3560), .P1_U3561(p1_u3561), .P1_U3562(p1_u3562), .P1_U3563(p1_u3563), .P1_U3564(p1_u3564), .P1_U3565(p1_u3565), .P1_U3566(p1_u3566), .P1_U3567(p1_u3567), .P1_U3568(p1_u3568), .P1_U3569(p1_u3569), .P1_U3570(p1_u3570), .P1_U3571(p1_u3571), .P1_U3572(p1_u3572), .P1_U3573(p1_u3573), .P1_U3574(p1_u3574), .P1_U3575(p1_u3575), .P1_U3576(p1_u3576), .P1_U3577(p1_u3577), .P1_U3578(p1_u3578), .P1_U3579(p1_u3579), .P1_U3580(p1_u3580), .P1_U3581(p1_u3581), .P1_U3582(p1_u3582), .P1_U3583(p1_u3583), .P1_U3584(p1_u3584), .P1_U3585(p1_u3585), .P1_U3586(p1_u3586), .P1_U3240(p1_u3240), .P1_U3239(p1_u3239), .P1_U3238(p1_u3238), .P1_U3237(p1_u3237), .P1_U3236(p1_u3236), .P1_U3235(p1_u3235), .P1_U3234(p1_u3234), .P1_U3233(p1_u3233), .P1_U3232(p1_u3232), .P1_U3231(p1_u3231), .P1_U3230(p1_u3230), .P1_U3229(p1_u3229), .P1_U3228(p1_u3228), .P1_U3227(p1_u3227), .P1_U3226(p1_u3226), .P1_U3225(p1_u3225), .P1_U3224(p1_u3224), .P1_U3223(p1_u3223), .P1_U3222(p1_u3222), .P1_U3221(p1_u3221), .P1_U3220(p1_u3220), .P1_U3219(p1_u3219), .P1_U3218(p1_u3218), .P1_U3217(p1_u3217), .P1_U3216(p1_u3216), .P1_U3215(p1_u3215), .P1_U3214(p1_u3214), .P1_U3213(p1_u3213), .P1_U3212(p1_u3212), .P1_U3211(p1_u3211), .P1_U3084(p1_u3084), .P1_U3083(p1_u3083), .P1_U4006(p1_u4006), .P2_U3358(p2_u3358), .P2_U3357(p2_u3357), .P2_U3356(p2_u3356), .P2_U3355(p2_u3355), .P2_U3354(p2_u3354), .P2_U3353(p2_u3353), .P2_U3352(p2_u3352), .P2_U3351(p2_u3351), .P2_U3350(p2_u3350), .P2_U3349(p2_u3349), .P2_U3348(p2_u3348), .P2_U3347(p2_u3347), .P2_U3346(p2_u3346), .P2_U3345(p2_u3345), .P2_U3344(p2_u3344), .P2_U3343(p2_u3343), .P2_U3342(p2_u3342), .P2_U3341(p2_u3341), .P2_U3340(p2_u3340), .P2_U3339(p2_u3339), .P2_U3338(p2_u3338), .P2_U3337(p2_u3337), .P2_U3336(p2_u3336), .P2_U3335(p2_u3335), .P2_U3334(p2_u3334), .P2_U3333(p2_u3333), .P2_U3332(p2_u3332), .P2_U3331(p2_u3331), .P2_U3330(p2_u3330), .P2_U3329(p2_u3329), .P2_U3328(p2_u3328), .P2_U3327(p2_u3327), .P2_U3437(p2_u3437), .P2_U3438(p2_u3438), .P2_U3326(p2_u3326), .P2_U3325(p2_u3325), .P2_U3324(p2_u3324), .P2_U3323(p2_u3323), .P2_U3322(p2_u3322), .P2_U3321(p2_u3321), .P2_U3320(p2_u3320), .P2_U3319(p2_u3319), .P2_U3318(p2_u3318), .P2_U3317(p2_u3317), .P2_U3316(p2_u3316), .P2_U3315(p2_u3315), .P2_U3314(p2_u3314), .P2_U3313(p2_u3313), .P2_U3312(p2_u3312), .P2_U3311(p2_u3311), .P2_U3310(p2_u3310), .P2_U3309(p2_u3309), .P2_U3308(p2_u3308), .P2_U3307(p2_u3307), .P2_U3306(p2_u3306), .P2_U3305(p2_u3305), .P2_U3304(p2_u3304), .P2_U3303(p2_u3303), .P2_U3302(p2_u3302), .P2_U3301(p2_u3301), .P2_U3300(p2_u3300), .P2_U3299(p2_u3299), .P2_U3298(p2_u3298), .P2_U3297(p2_u3297), .P2_U3451(p2_u3451), .P2_U3454(p2_u3454), .P2_U3457(p2_u3457), .P2_U3460(p2_u3460), .P2_U3463(p2_u3463), .P2_U3466(p2_u3466), .P2_U3469(p2_u3469), .P2_U3472(p2_u3472), .P2_U3475(p2_u3475), .P2_U3478(p2_u3478), .P2_U3481(p2_u3481), .P2_U3484(p2_u3484), .P2_U3487(p2_u3487), .P2_U3490(p2_u3490), .P2_U3493(p2_u3493), .P2_U3496(p2_u3496), .P2_U3499(p2_u3499), .P2_U3502(p2_u3502), .P2_U3505(p2_u3505), .P2_U3507(p2_u3507), .P2_U3508(p2_u3508), .P2_U3509(p2_u3509), .P2_U3510(p2_u3510), .P2_U3511(p2_u3511), .P2_U3512(p2_u3512), .P2_U3513(p2_u3513), .P2_U3514(p2_u3514), .P2_U3515(p2_u3515), .P2_U3516(p2_u3516), .P2_U3517(p2_u3517), .P2_U3518(p2_u3518), .P2_U3519(p2_u3519), .P2_U3520(p2_u3520), .P2_U3521(p2_u3521), .P2_U3522(p2_u3522), .P2_U3523(p2_u3523), .P2_U3524(p2_u3524), .P2_U3525(p2_u3525), .P2_U3526(p2_u3526), .P2_U3527(p2_u3527), .P2_U3528(p2_u3528), .P2_U3529(p2_u3529), .P2_U3530(p2_u3530), .P2_U3531(p2_u3531), .P2_U3532(p2_u3532), .P2_U3533(p2_u3533), .P2_U3534(p2_u3534), .P2_U3535(p2_u3535), .P2_U3536(p2_u3536), .P2_U3537(p2_u3537), .P2_U3538(p2_u3538), .P2_U3539(p2_u3539), .P2_U3540(p2_u3540), .P2_U3541(p2_u3541), .P2_U3542(p2_u3542), .P2_U3543(p2_u3543), .P2_U3544(p2_u3544), .P2_U3545(p2_u3545), .P2_U3546(p2_u3546), .P2_U3547(p2_u3547), .P2_U3548(p2_u3548), .P2_U3549(p2_u3549), .P2_U3550(p2_u3550), .P2_U3551(p2_u3551), .P2_U3296(p2_u3296), .P2_U3295(p2_u3295), .P2_U3294(p2_u3294), .P2_U3293(p2_u3293), .P2_U3292(p2_u3292), .P2_U3291(p2_u3291), .P2_U3290(p2_u3290), .P2_U3289(p2_u3289), .P2_U3288(p2_u3288), .P2_U3287(p2_u3287), .P2_U3286(p2_u3286), .P2_U3285(p2_u3285), .P2_U3284(p2_u3284), .P2_U3283(p2_u3283), .P2_U3282(p2_u3282), .P2_U3281(p2_u3281), .P2_U3280(p2_u3280), .P2_U3279(p2_u3279), .P2_U3278(p2_u3278), .P2_U3277(p2_u3277), .P2_U3276(p2_u3276), .P2_U3275(p2_u3275), .P2_U3274(p2_u3274), .P2_U3273(p2_u3273), .P2_U3272(p2_u3272), .P2_U3271(p2_u3271), .P2_U3270(p2_u3270), .P2_U3269(p2_u3269), .P2_U3268(p2_u3268), .P2_U3267(p2_u3267), .P2_U3266(p2_u3266), .P2_U3265(p2_u3265), .P2_U3264(p2_u3264), .P2_U3263(p2_u3263), .P2_U3262(p2_u3262), .P2_U3261(p2_u3261), .P2_U3260(p2_u3260), .P2_U3259(p2_u3259), .P2_U3258(p2_u3258), .P2_U3257(p2_u3257), .P2_U3256(p2_u3256), .P2_U3255(p2_u3255), .P2_U3254(p2_u3254), .P2_U3253(p2_u3253), .P2_U3252(p2_u3252), .P2_U3251(p2_u3251), .P2_U3250(p2_u3250), .P2_U3249(p2_u3249), .P2_U3248(p2_u3248), .P2_U3247(p2_u3247), .P2_U3246(p2_u3246), .P2_U3245(p2_u3245), .P2_U3552(p2_u3552), .P2_U3553(p2_u3553), .P2_U3554(p2_u3554), .P2_U3555(p2_u3555), .P2_U3556(p2_u3556), .P2_U3557(p2_u3557), .P2_U3558(p2_u3558), .P2_U3559(p2_u3559), .P2_U3560(p2_u3560), .P2_U3561(p2_u3561), .P2_U3562(p2_u3562), .P2_U3563(p2_u3563), .P2_U3564(p2_u3564), .P2_U3565(p2_u3565), .P2_U3566(p2_u3566), .P2_U3567(p2_u3567), .P2_U3568(p2_u3568), .P2_U3569(p2_u3569), .P2_U3570(p2_u3570), .P2_U3571(p2_u3571), .P2_U3572(p2_u3572), .P2_U3573(p2_u3573), .P2_U3574(p2_u3574), .P2_U3575(p2_u3575), .P2_U3576(p2_u3576), .P2_U3577(p2_u3577), .P2_U3578(p2_u3578), .P2_U3579(p2_u3579), .P2_U3580(p2_u3580), .P2_U3581(p2_u3581), .P2_U3582(p2_u3582), .P2_U3583(p2_u3583), .P2_U3244(p2_u3244), .P2_U3243(p2_u3243), .P2_U3242(p2_u3242), .P2_U3241(p2_u3241), .P2_U3240(p2_u3240), .P2_U3239(p2_u3239), .P2_U3238(p2_u3238), .P2_U3237(p2_u3237), .P2_U3236(p2_u3236), .P2_U3235(p2_u3235), .P2_U3234(p2_u3234), .P2_U3233(p2_u3233), .P2_U3232(p2_u3232), .P2_U3231(p2_u3231), .P2_U3230(p2_u3230), .P2_U3229(p2_u3229), .P2_U3228(p2_u3228), .P2_U3227(p2_u3227), .P2_U3226(p2_u3226), .P2_U3225(p2_u3225), .P2_U3224(p2_u3224), .P2_U3223(p2_u3223), .P2_U3222(p2_u3222), .P2_U3221(p2_u3221), .P2_U3220(p2_u3220), .P2_U3219(p2_u3219), .P2_U3218(p2_u3218), .P2_U3217(p2_u3217), .P2_U3216(p2_u3216), .P2_U3215(p2_u3215), .P2_U3152(p2_u3152), .P2_U3151(p2_u3151), .P2_U3966(p2_u3966));

integer i=0;
always @ (posedge clk) begin
	vec = input_vec_mem[i];
	$monitor(vec);
	i = i + 1;

end

always @ (negedge clk)begin
	$fdisplay ( fh_w, add_1071_u4, add_1071_u55, add_1071_u56, add_1071_u57, add_1071_u58, add_1071_u59, add_1071_u60, add_1071_u61, add_1071_u62, add_1071_u63, add_1071_u47, add_1071_u48, add_1071_u49, add_1071_u50, add_1071_u51, add_1071_u52, add_1071_u53, add_1071_u54, add_1071_u5, add_1071_u46, u126, u123, p1_u3353, p1_u3352, p1_u3351, p1_u3350, p1_u3349, p1_u3348, p1_u3347, p1_u3346, p1_u3345, p1_u3344, p1_u3343, p1_u3342, p1_u3341, p1_u3340, p1_u3339, p1_u3338, p1_u3337, p1_u3336, p1_u3335, p1_u3334, p1_u3333, p1_u3332, p1_u3331, p1_u3330, p1_u3329, p1_u3328, p1_u3327, p1_u3326, p1_u3325, p1_u3324, p1_u3323, p1_u3322, p1_u3440, p1_u3441, p1_u3321, p1_u3320, p1_u3319, p1_u3318, p1_u3317, p1_u3316, p1_u3315, p1_u3314, p1_u3313, p1_u3312, p1_u3311, p1_u3310, p1_u3309, p1_u3308, p1_u3307, p1_u3306, p1_u3305, p1_u3304, p1_u3303, p1_u3302, p1_u3301, p1_u3300, p1_u3299, p1_u3298, p1_u3297, p1_u3296, p1_u3295, p1_u3294, p1_u3293, p1_u3292, p1_u3454, p1_u3457, p1_u3460, p1_u3463, p1_u3466, p1_u3469, p1_u3472, p1_u3475, p1_u3478, p1_u3481, p1_u3484, p1_u3487, p1_u3490, p1_u3493, p1_u3496, p1_u3499, p1_u3502, p1_u3505, p1_u3508, p1_u3510, p1_u3511, p1_u3512, p1_u3513, p1_u3514, p1_u3515, p1_u3516, p1_u3517, p1_u3518, p1_u3519, p1_u3520, p1_u3521, p1_u3522, p1_u3523, p1_u3524, p1_u3525, p1_u3526, p1_u3527, p1_u3528, p1_u3529, p1_u3530, p1_u3531, p1_u3532, p1_u3533, p1_u3534, p1_u3535, p1_u3536, p1_u3537, p1_u3538, p1_u3539, p1_u3540, p1_u3541, p1_u3542, p1_u3543, p1_u3544, p1_u3545, p1_u3546, p1_u3547, p1_u3548, p1_u3549, p1_u3550, p1_u3551, p1_u3552, p1_u3553, p1_u3554, p1_u3291, p1_u3290, p1_u3289, p1_u3288, p1_u3287, p1_u3286, p1_u3285, p1_u3284, p1_u3283, p1_u3282, p1_u3281, p1_u3280, p1_u3279, p1_u3278, p1_u3277, p1_u3276, p1_u3275, p1_u3274, p1_u3273, p1_u3272, p1_u3271, p1_u3270, p1_u3269, p1_u3268, p1_u3267, p1_u3266, p1_u3265, p1_u3264, p1_u3263, p1_u3355, p1_u3262, p1_u3261, p1_u3260, p1_u3259, p1_u3258, p1_u3257, p1_u3256, p1_u3255, p1_u3254, p1_u3253, p1_u3252, p1_u3251, p1_u3250, p1_u3249, p1_u3248, p1_u3247, p1_u3246, p1_u3245, p1_u3244, p1_u3243, p1_u3242, p1_u3241, p1_u3555, p1_u3556, p1_u3557, p1_u3558, p1_u3559, p1_u3560, p1_u3561, p1_u3562, p1_u3563, p1_u3564, p1_u3565, p1_u3566, p1_u3567, p1_u3568, p1_u3569, p1_u3570, p1_u3571, p1_u3572, p1_u3573, p1_u3574, p1_u3575, p1_u3576, p1_u3577, p1_u3578, p1_u3579, p1_u3580, p1_u3581, p1_u3582, p1_u3583, p1_u3584, p1_u3585, p1_u3586, p1_u3240, p1_u3239, p1_u3238, p1_u3237, p1_u3236, p1_u3235, p1_u3234, p1_u3233, p1_u3232, p1_u3231, p1_u3230, p1_u3229, p1_u3228, p1_u3227, p1_u3226, p1_u3225, p1_u3224, p1_u3223, p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218, p1_u3217, p1_u3216, p1_u3215, p1_u3214, p1_u3213, p1_u3212, p1_u3211, p1_u3084, p1_u3083, p1_u4006, p2_u3358, p2_u3357, p2_u3356, p2_u3355, p2_u3354, p2_u3353, p2_u3352, p2_u3351, p2_u3350, p2_u3349, p2_u3348, p2_u3347, p2_u3346, p2_u3345, p2_u3344, p2_u3343, p2_u3342, p2_u3341, p2_u3340, p2_u3339, p2_u3338, p2_u3337, p2_u3336, p2_u3335, p2_u3334, p2_u3333, p2_u3332, p2_u3331, p2_u3330, p2_u3329, p2_u3328, p2_u3327, p2_u3437, p2_u3438, p2_u3326, p2_u3325, p2_u3324, p2_u3323, p2_u3322, p2_u3321, p2_u3320, p2_u3319, p2_u3318, p2_u3317, p2_u3316, p2_u3315, p2_u3314, p2_u3313, p2_u3312, p2_u3311, p2_u3310, p2_u3309, p2_u3308, p2_u3307, p2_u3306, p2_u3305, p2_u3304, p2_u3303, p2_u3302, p2_u3301, p2_u3300, p2_u3299, p2_u3298, p2_u3297, p2_u3451, p2_u3454, p2_u3457, p2_u3460, p2_u3463, p2_u3466, p2_u3469, p2_u3472, p2_u3475, p2_u3478, p2_u3481, p2_u3484, p2_u3487, p2_u3490, p2_u3493, p2_u3496, p2_u3499, p2_u3502, p2_u3505, p2_u3507, p2_u3508, p2_u3509, p2_u3510, p2_u3511, p2_u3512, p2_u3513, p2_u3514, p2_u3515, p2_u3516, p2_u3517, p2_u3518, p2_u3519, p2_u3520, p2_u3521, p2_u3522, p2_u3523, p2_u3524, p2_u3525, p2_u3526, p2_u3527, p2_u3528, p2_u3529, p2_u3530, p2_u3531, p2_u3532, p2_u3533, p2_u3534, p2_u3535, p2_u3536, p2_u3537, p2_u3538, p2_u3539, p2_u3540, p2_u3541, p2_u3542, p2_u3543, p2_u3544, p2_u3545, p2_u3546, p2_u3547, p2_u3548, p2_u3549, p2_u3550, p2_u3551, p2_u3296, p2_u3295, p2_u3294, p2_u3293, p2_u3292, p2_u3291, p2_u3290, p2_u3289, p2_u3288, p2_u3287, p2_u3286, p2_u3285, p2_u3284, p2_u3283, p2_u3282, p2_u3281, p2_u3280, p2_u3279, p2_u3278, p2_u3277, p2_u3276, p2_u3275, p2_u3274, p2_u3273, p2_u3272, p2_u3271, p2_u3270, p2_u3269, p2_u3268, p2_u3267, p2_u3266, p2_u3265, p2_u3264, p2_u3263, p2_u3262, p2_u3261, p2_u3260, p2_u3259, p2_u3258, p2_u3257, p2_u3256, p2_u3255, p2_u3254, p2_u3253, p2_u3252, p2_u3251, p2_u3250, p2_u3249, p2_u3248, p2_u3247, p2_u3246, p2_u3245, p2_u3552, p2_u3553, p2_u3554, p2_u3555, p2_u3556, p2_u3557, p2_u3558, p2_u3559, p2_u3560, p2_u3561, p2_u3562, p2_u3563, p2_u3564, p2_u3565, p2_u3566, p2_u3567, p2_u3568, p2_u3569, p2_u3570, p2_u3571, p2_u3572, p2_u3573, p2_u3574, p2_u3575, p2_u3576, p2_u3577, p2_u3578, p2_u3579, p2_u3580, p2_u3581, p2_u3582, p2_u3583, p2_u3244, p2_u3243, p2_u3242, p2_u3241, p2_u3240, p2_u3239, p2_u3238, p2_u3237, p2_u3236, p2_u3235, p2_u3234, p2_u3233, p2_u3232, p2_u3231, p2_u3230, p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225, p2_u3224, p2_u3223, p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218, p2_u3217, p2_u3216, p2_u3215, p2_u3152, p2_u3151, p2_u3966);
	if(i == vec_length)begin
		$finish;
	end
end

integer fh_w;
initial begin
	fh_w = $fopen(`out_file, "w");
end
 
initial begin
	//$fsdbDumpfile("SET.fsdb");
	//$fsdbDumpvars;
	//$fsdbDumpMDA;
	$dumpfile("test_result.vcd");
    $dumpvars;

end
endmodule
