`timescale 1ns/10ps

`define cycle 10.0
`define terminate_cycle 400000//200000 // Modify your terminate ycle here

module b15_ras_testfixture;

`define in_file "b15_ras/rand_input_vector_b15_ras_0.out"
`define out_file "b15_ras/rand_output_vector_b15_ras_0.out"

parameter vec_width = 485;
parameter vec_length = 7;

reg clk = 0;


reg [vec_width-1:0] input_vec_mem [0:vec_length-1];
reg [vec_width-1:0] vec;

wire u3445, u3446, u3447, u3448, u3213, u3212, u3211, u3210, u3209, u3208, u3207, u3206, u3205, u3204, u3203, u3202, u3201, u3200, u3199, u3198, u3197, u3196, u3195, u3194, u3193, u3192, u3191, u3190, u3189, u3188, u3187, u3186, u3185, u3184, u3183, u3182, u3181, u3451, u3452, u3180, u3179, u3178, u3177, u3176, u3175, u3174, u3173, u3172, u3171, u3170, u3169, u3168, u3167, u3166, u3165, u3164, u3163, u3162, u3161, u3160, u3159, u3158, u3157, u3156, u3155, u3154, u3153, u3152, u3151, u3453, u3150, u3149, u3148, u3147, u3146, u3145, u3144, u3143, u3142, u3141, u3140, u3139, u3138, u3137, u3136, u3135, u3134, u3133, u3132, u3131, u3130, u3129, u3128, u3127, u3126, u3125, u3124, u3123, u3122, u3121, u3120, u3119, u3118, u3117, u3116, u3115, u3114, u3113, u3112, u3111, u3110, u3109, u3108, u3107, u3106, u3105, u3104, u3103, u3102, u3101, u3100, u3099, u3098, u3097, u3096, u3095, u3094, u3093, u3092, u3091, u3090, u3089, u3088, u3087, u3086, u3085, u3084, u3083, u3082, u3081, u3080, u3079, u3078, u3077, u3076, u3075, u3074, u3073, u3072, u3071, u3070, u3069, u3068, u3067, u3066, u3065, u3064, u3063, u3062, u3061, u3060, u3059, u3058, u3057, u3056, u3055, u3054, u3053, u3052, u3051, u3050, u3049, u3048, u3047, u3046, u3045, u3044, u3043, u3042, u3041, u3040, u3039, u3038, u3037, u3036, u3035, u3034, u3033, u3032, u3031, u3030, u3029, u3028, u3027, u3026, u3025, u3024, u3023, u3022, u3021, u3020, u3455, u3456, u3459, u3460, u3461, u3019, u3462, u3463, u3464, u3465, u3018, u3017, u3016, u3015, u3014, u3013, u3012, u3011, u3010, u3009, u3008, u3007, u3006, u3005, u3004, u3003, u3002, u3001, u3000, u2999, u2998, u2997, u2996, u2995, u2994, u2993, u2992, u2991, u2990, u2989, u2988, u2987, u2986, u2985, u2984, u2983, u2982, u2981, u2980, u2979, u2978, u2977, u2976, u2975, u2974, u2973, u2972, u2971, u2970, u2969, u2968, u2967, u2966, u2965, u2964, u2963, u2962, u2961, u2960, u2959, u2958, u2957, u2956, u2955, u2954, u2953, u2952, u2951, u2950, u2949, u2948, u2947, u2946, u2945, u2944, u2943, u2942, u2941, u2940, u2939, u2938, u2937, u2936, u2935, u2934, u2933, u2932, u2931, u2930, u2929, u2928, u2927, u2926, u2925, u2924, u2923, u2922, u2921, u2920, u2919, u2918, u2917, u2916, u2915, u2914, u2913, u2912, u2911, u2910, u2909, u2908, u2907, u2906, u2905, u2904, u2903, u2902, u2901, u2900, u2899, u2898, u2897, u2896, u2895, u2894, u2893, u2892, u2891, u2890, u2889, u2888, u2887, u2886, u2885, u2884, u2883, u2882, u2881, u2880, u2879, u2878, u2877, u2876, u2875, u2874, u2873, u2872, u2871, u2870, u2869, u2868, u2867, u2866, u2865, u2864, u2863, u2862, u2861, u2860, u2859, u2858, u2857, u2856, u2855, u2854, u2853, u2852, u2851, u2850, u2849, u2848, u2847, u2846, u2845, u2844, u2843, u2842, u2841, u2840, u2839, u2838, u2837, u2836, u2835, u2834, u2833, u2832, u2831, u2830, u2829, u2828, u2827, u2826, u2825, u2824, u2823, u2822, u2821, u2820, u2819, u2818, u2817, u2816, u2815, u2814, u2813, u2812, u2811, u2810, u2809, u2808, u2807, u2806, u2805, u2804, u2803, u2802, u2801, u2800, u2799, u2798, u2797, u2796, u2795, u3468, u2794, u3469, u3470, u2793, u3471, u2792, u3472, u2791, u3473, u2790, u2789, u3474, u2788, be_n_reg_3_, be_n_reg_2_, be_n_reg_1_, be_n_reg_0_, address_reg_29_, address_reg_28_, address_reg_27_, address_reg_26_, address_reg_25_, address_reg_24_, address_reg_23_, address_reg_22_, address_reg_21_, address_reg_20_, address_reg_19_, address_reg_18_, address_reg_17_, address_reg_16_, address_reg_15_, address_reg_14_, address_reg_13_, address_reg_12_, address_reg_11_, address_reg_10_, address_reg_9_, address_reg_8_, address_reg_7_, address_reg_6_, address_reg_5_, address_reg_4_, address_reg_3_, address_reg_2_, address_reg_1_, address_reg_0_, w_r_n_reg, d_c_n_reg, m_io_n_reg, ads_n_reg, datao_reg_31_, datao_reg_30_, datao_reg_29_, datao_reg_28_, datao_reg_27_, datao_reg_26_, datao_reg_25_, datao_reg_24_, datao_reg_23_, datao_reg_22_, datao_reg_21_, datao_reg_20_, datao_reg_19_, datao_reg_18_, datao_reg_17_, datao_reg_16_, datao_reg_15_, datao_reg_14_, datao_reg_13_, datao_reg_12_, datao_reg_11_, datao_reg_10_, datao_reg_9_, datao_reg_8_, datao_reg_7_, datao_reg_6_, datao_reg_5_, datao_reg_4_, datao_reg_3_, datao_reg_2_, datao_reg_1_, datao_reg_0_;
initial begin
	$readmemb(`in_file, input_vec_mem );
end

always #(`cycle/2) clk = ~clk;

b15_ras cc (.BE_N_REG_3__EXTRA(vec[484]), .BE_N_REG_2__EXTRA(vec[483]), .BE_N_REG_1__EXTRA(vec[482]), .BE_N_REG_0__EXTRA(vec[481]), .ADDRESS_REG_29__EXTRA(vec[480]), .ADDRESS_REG_28__EXTRA(vec[479]), .ADDRESS_REG_27__EXTRA(vec[478]), .ADDRESS_REG_26__EXTRA(vec[477]), .ADDRESS_REG_25__EXTRA(vec[476]), .ADDRESS_REG_24__EXTRA(vec[475]), .ADDRESS_REG_23__EXTRA(vec[474]), .ADDRESS_REG_22__EXTRA(vec[473]), .ADDRESS_REG_21__EXTRA(vec[472]), .ADDRESS_REG_20__EXTRA(vec[471]), .ADDRESS_REG_19__EXTRA(vec[470]), .ADDRESS_REG_18__EXTRA(vec[469]), .ADDRESS_REG_17__EXTRA(vec[468]), .ADDRESS_REG_16__EXTRA(vec[467]), .ADDRESS_REG_15__EXTRA(vec[466]), .ADDRESS_REG_14__EXTRA(vec[465]), .ADDRESS_REG_13__EXTRA(vec[464]), .ADDRESS_REG_12__EXTRA(vec[463]), .ADDRESS_REG_11__EXTRA(vec[462]), .ADDRESS_REG_10__EXTRA(vec[461]), .ADDRESS_REG_9__EXTRA(vec[460]), .ADDRESS_REG_8__EXTRA(vec[459]), .ADDRESS_REG_7__EXTRA(vec[458]), .ADDRESS_REG_6__EXTRA(vec[457]), .ADDRESS_REG_5__EXTRA(vec[456]), .ADDRESS_REG_4__EXTRA(vec[455]), .ADDRESS_REG_3__EXTRA(vec[454]), .ADDRESS_REG_2__EXTRA(vec[453]), .ADDRESS_REG_1__EXTRA(vec[452]), .ADDRESS_REG_0__EXTRA(vec[451]), .STATE_REG_2_(vec[450]), .STATE_REG_1_(vec[449]), .STATE_REG_0_(vec[448]), .DATAWIDTH_REG_0_(vec[447]), .DATAWIDTH_REG_1_(vec[446]), .DATAWIDTH_REG_2_(vec[445]), .DATAWIDTH_REG_3_(vec[444]), .DATAWIDTH_REG_4_(vec[443]), .DATAWIDTH_REG_5_(vec[442]), .DATAWIDTH_REG_6_(vec[441]), .DATAWIDTH_REG_7_(vec[440]), .DATAWIDTH_REG_8_(vec[439]), .DATAWIDTH_REG_9_(vec[438]), .DATAWIDTH_REG_10_(vec[437]), .DATAWIDTH_REG_11_(vec[436]), .DATAWIDTH_REG_12_(vec[435]), .DATAWIDTH_REG_13_(vec[434]), .DATAWIDTH_REG_14_(vec[433]), .DATAWIDTH_REG_15_(vec[432]), .DATAWIDTH_REG_16_(vec[431]), .DATAWIDTH_REG_17_(vec[430]), .DATAWIDTH_REG_18_(vec[429]), .DATAWIDTH_REG_19_(vec[428]), .DATAWIDTH_REG_20_(vec[427]), .DATAWIDTH_REG_21_(vec[426]), .DATAWIDTH_REG_22_(vec[425]), .DATAWIDTH_REG_23_(vec[424]), .DATAWIDTH_REG_24_(vec[423]), .DATAWIDTH_REG_25_(vec[422]), .DATAWIDTH_REG_26_(vec[421]), .DATAWIDTH_REG_27_(vec[420]), .DATAWIDTH_REG_28_(vec[419]), .DATAWIDTH_REG_29_(vec[418]), .DATAWIDTH_REG_30_(vec[417]), .DATAWIDTH_REG_31_(vec[416]), .STATE2_REG_3_(vec[415]), .STATE2_REG_2_(vec[414]), .STATE2_REG_1_(vec[413]), .STATE2_REG_0_(vec[412]), .INSTQUEUE_REG_15__7_(vec[411]), .INSTQUEUE_REG_15__6_(vec[410]), .INSTQUEUE_REG_15__5_(vec[409]), .INSTQUEUE_REG_15__4_(vec[408]), .INSTQUEUE_REG_15__3_(vec[407]), .INSTQUEUE_REG_15__2_(vec[406]), .INSTQUEUE_REG_15__1_(vec[405]), .INSTQUEUE_REG_15__0_(vec[404]), .INSTQUEUE_REG_14__7_(vec[403]), .INSTQUEUE_REG_14__6_(vec[402]), .INSTQUEUE_REG_14__5_(vec[401]), .INSTQUEUE_REG_14__4_(vec[400]), .INSTQUEUE_REG_14__3_(vec[399]), .INSTQUEUE_REG_14__2_(vec[398]), .INSTQUEUE_REG_14__1_(vec[397]), .INSTQUEUE_REG_14__0_(vec[396]), .INSTQUEUE_REG_13__7_(vec[395]), .INSTQUEUE_REG_13__6_(vec[394]), .INSTQUEUE_REG_13__5_(vec[393]), .INSTQUEUE_REG_13__4_(vec[392]), .INSTQUEUE_REG_13__3_(vec[391]), .INSTQUEUE_REG_13__2_(vec[390]), .INSTQUEUE_REG_13__1_(vec[389]), .INSTQUEUE_REG_13__0_(vec[388]), .INSTQUEUE_REG_12__7_(vec[387]), .INSTQUEUE_REG_12__6_(vec[386]), .INSTQUEUE_REG_12__5_(vec[385]), .INSTQUEUE_REG_12__4_(vec[384]), .INSTQUEUE_REG_12__3_(vec[383]), .INSTQUEUE_REG_12__2_(vec[382]), .INSTQUEUE_REG_12__1_(vec[381]), .INSTQUEUE_REG_12__0_(vec[380]), .INSTQUEUE_REG_11__7_(vec[379]), .INSTQUEUE_REG_11__6_(vec[378]), .INSTQUEUE_REG_11__5_(vec[377]), .INSTQUEUE_REG_11__4_(vec[376]), .INSTQUEUE_REG_11__3_(vec[375]), .INSTQUEUE_REG_11__2_(vec[374]), .INSTQUEUE_REG_11__1_(vec[373]), .INSTQUEUE_REG_11__0_(vec[372]), .INSTQUEUE_REG_10__7_(vec[371]), .INSTQUEUE_REG_10__6_(vec[370]), .INSTQUEUE_REG_10__5_(vec[369]), .INSTQUEUE_REG_10__4_(vec[368]), .INSTQUEUE_REG_10__3_(vec[367]), .INSTQUEUE_REG_10__2_(vec[366]), .INSTQUEUE_REG_10__1_(vec[365]), .INSTQUEUE_REG_10__0_(vec[364]), .INSTQUEUE_REG_9__7_(vec[363]), .INSTQUEUE_REG_9__6_(vec[362]), .INSTQUEUE_REG_9__5_(vec[361]), .INSTQUEUE_REG_9__4_(vec[360]), .INSTQUEUE_REG_9__3_(vec[359]), .INSTQUEUE_REG_9__2_(vec[358]), .INSTQUEUE_REG_9__1_(vec[357]), .INSTQUEUE_REG_9__0_(vec[356]), .INSTQUEUE_REG_8__7_(vec[355]), .INSTQUEUE_REG_8__6_(vec[354]), .INSTQUEUE_REG_8__5_(vec[353]), .INSTQUEUE_REG_8__4_(vec[352]), .INSTQUEUE_REG_8__3_(vec[351]), .INSTQUEUE_REG_8__2_(vec[350]), .INSTQUEUE_REG_8__1_(vec[349]), .INSTQUEUE_REG_8__0_(vec[348]), .INSTQUEUE_REG_7__7_(vec[347]), .INSTQUEUE_REG_7__6_(vec[346]), .INSTQUEUE_REG_7__5_(vec[345]), .INSTQUEUE_REG_7__4_(vec[344]), .INSTQUEUE_REG_7__3_(vec[343]), .INSTQUEUE_REG_7__2_(vec[342]), .INSTQUEUE_REG_7__1_(vec[341]), .INSTQUEUE_REG_7__0_(vec[340]), .INSTQUEUE_REG_6__7_(vec[339]), .INSTQUEUE_REG_6__6_(vec[338]), .INSTQUEUE_REG_6__5_(vec[337]), .INSTQUEUE_REG_6__4_(vec[336]), .INSTQUEUE_REG_6__3_(vec[335]), .INSTQUEUE_REG_6__2_(vec[334]), .INSTQUEUE_REG_6__1_(vec[333]), .INSTQUEUE_REG_6__0_(vec[332]), .INSTQUEUE_REG_5__7_(vec[331]), .INSTQUEUE_REG_5__6_(vec[330]), .INSTQUEUE_REG_5__5_(vec[329]), .INSTQUEUE_REG_5__4_(vec[328]), .INSTQUEUE_REG_5__3_(vec[327]), .INSTQUEUE_REG_5__2_(vec[326]), .INSTQUEUE_REG_5__1_(vec[325]), .INSTQUEUE_REG_5__0_(vec[324]), .INSTQUEUE_REG_4__7_(vec[323]), .INSTQUEUE_REG_4__6_(vec[322]), .INSTQUEUE_REG_4__5_(vec[321]), .INSTQUEUE_REG_4__4_(vec[320]), .INSTQUEUE_REG_4__3_(vec[319]), .INSTQUEUE_REG_4__2_(vec[318]), .INSTQUEUE_REG_4__1_(vec[317]), .INSTQUEUE_REG_4__0_(vec[316]), .INSTQUEUE_REG_3__7_(vec[315]), .INSTQUEUE_REG_3__6_(vec[314]), .INSTQUEUE_REG_3__5_(vec[313]), .INSTQUEUE_REG_3__4_(vec[312]), .INSTQUEUE_REG_3__3_(vec[311]), .INSTQUEUE_REG_3__2_(vec[310]), .INSTQUEUE_REG_3__1_(vec[309]), .INSTQUEUE_REG_3__0_(vec[308]), .INSTQUEUE_REG_2__7_(vec[307]), .INSTQUEUE_REG_2__6_(vec[306]), .INSTQUEUE_REG_2__5_(vec[305]), .INSTQUEUE_REG_2__4_(vec[304]), .INSTQUEUE_REG_2__3_(vec[303]), .INSTQUEUE_REG_2__2_(vec[302]), .INSTQUEUE_REG_2__1_(vec[301]), .INSTQUEUE_REG_2__0_(vec[300]), .INSTQUEUE_REG_1__7_(vec[299]), .INSTQUEUE_REG_1__6_(vec[298]), .INSTQUEUE_REG_1__5_(vec[297]), .INSTQUEUE_REG_1__4_(vec[296]), .INSTQUEUE_REG_1__3_(vec[295]), .INSTQUEUE_REG_1__2_(vec[294]), .INSTQUEUE_REG_1__1_(vec[293]), .INSTQUEUE_REG_1__0_(vec[292]), .INSTQUEUE_REG_0__7_(vec[291]), .INSTQUEUE_REG_0__6_(vec[290]), .INSTQUEUE_REG_0__5_(vec[289]), .INSTQUEUE_REG_0__4_(vec[288]), .INSTQUEUE_REG_0__3_(vec[287]), .INSTQUEUE_REG_0__2_(vec[286]), .INSTQUEUE_REG_0__1_(vec[285]), .INSTQUEUE_REG_0__0_(vec[284]), .INSTQUEUERD_ADDR_REG_4_(vec[283]), .INSTQUEUERD_ADDR_REG_3_(vec[282]), .INSTQUEUERD_ADDR_REG_2_(vec[281]), .INSTQUEUERD_ADDR_REG_1_(vec[280]), .INSTQUEUERD_ADDR_REG_0_(vec[279]), .INSTQUEUEWR_ADDR_REG_4_(vec[278]), .INSTQUEUEWR_ADDR_REG_3_(vec[277]), .INSTQUEUEWR_ADDR_REG_2_(vec[276]), .INSTQUEUEWR_ADDR_REG_1_(vec[275]), .INSTQUEUEWR_ADDR_REG_0_(vec[274]), .INSTADDRPOINTER_REG_0_(vec[273]), .INSTADDRPOINTER_REG_1_(vec[272]), .INSTADDRPOINTER_REG_2_(vec[271]), .INSTADDRPOINTER_REG_3_(vec[270]), .INSTADDRPOINTER_REG_4_(vec[269]), .INSTADDRPOINTER_REG_5_(vec[268]), .INSTADDRPOINTER_REG_6_(vec[267]), .INSTADDRPOINTER_REG_7_(vec[266]), .INSTADDRPOINTER_REG_8_(vec[265]), .INSTADDRPOINTER_REG_9_(vec[264]), .INSTADDRPOINTER_REG_10_(vec[263]), .INSTADDRPOINTER_REG_11_(vec[262]), .INSTADDRPOINTER_REG_12_(vec[261]), .INSTADDRPOINTER_REG_13_(vec[260]), .INSTADDRPOINTER_REG_14_(vec[259]), .INSTADDRPOINTER_REG_15_(vec[258]), .INSTADDRPOINTER_REG_16_(vec[257]), .INSTADDRPOINTER_REG_17_(vec[256]), .INSTADDRPOINTER_REG_18_(vec[255]), .INSTADDRPOINTER_REG_19_(vec[254]), .INSTADDRPOINTER_REG_20_(vec[253]), .INSTADDRPOINTER_REG_21_(vec[252]), .INSTADDRPOINTER_REG_22_(vec[251]), .INSTADDRPOINTER_REG_23_(vec[250]), .INSTADDRPOINTER_REG_24_(vec[249]), .INSTADDRPOINTER_REG_25_(vec[248]), .INSTADDRPOINTER_REG_26_(vec[247]), .INSTADDRPOINTER_REG_27_(vec[246]), .INSTADDRPOINTER_REG_28_(vec[245]), .INSTADDRPOINTER_REG_29_(vec[244]), .INSTADDRPOINTER_REG_30_(vec[243]), .INSTADDRPOINTER_REG_31_(vec[242]), .PHYADDRPOINTER_REG_0_(vec[241]), .PHYADDRPOINTER_REG_1_(vec[240]), .PHYADDRPOINTER_REG_2_(vec[239]), .PHYADDRPOINTER_REG_3_(vec[238]), .PHYADDRPOINTER_REG_4_(vec[237]), .PHYADDRPOINTER_REG_5_(vec[236]), .PHYADDRPOINTER_REG_6_(vec[235]), .PHYADDRPOINTER_REG_7_(vec[234]), .PHYADDRPOINTER_REG_8_(vec[233]), .PHYADDRPOINTER_REG_9_(vec[232]), .PHYADDRPOINTER_REG_10_(vec[231]), .PHYADDRPOINTER_REG_11_(vec[230]), .PHYADDRPOINTER_REG_12_(vec[229]), .PHYADDRPOINTER_REG_13_(vec[228]), .PHYADDRPOINTER_REG_14_(vec[227]), .PHYADDRPOINTER_REG_15_(vec[226]), .PHYADDRPOINTER_REG_16_(vec[225]), .PHYADDRPOINTER_REG_17_(vec[224]), .PHYADDRPOINTER_REG_18_(vec[223]), .PHYADDRPOINTER_REG_19_(vec[222]), .PHYADDRPOINTER_REG_20_(vec[221]), .PHYADDRPOINTER_REG_21_(vec[220]), .PHYADDRPOINTER_REG_22_(vec[219]), .PHYADDRPOINTER_REG_23_(vec[218]), .PHYADDRPOINTER_REG_24_(vec[217]), .PHYADDRPOINTER_REG_25_(vec[216]), .PHYADDRPOINTER_REG_26_(vec[215]), .PHYADDRPOINTER_REG_27_(vec[214]), .PHYADDRPOINTER_REG_28_(vec[213]), .PHYADDRPOINTER_REG_29_(vec[212]), .PHYADDRPOINTER_REG_30_(vec[211]), .PHYADDRPOINTER_REG_31_(vec[210]), .LWORD_REG_15_(vec[209]), .LWORD_REG_14_(vec[208]), .LWORD_REG_13_(vec[207]), .LWORD_REG_12_(vec[206]), .LWORD_REG_11_(vec[205]), .LWORD_REG_10_(vec[204]), .LWORD_REG_9_(vec[203]), .LWORD_REG_8_(vec[202]), .LWORD_REG_7_(vec[201]), .LWORD_REG_6_(vec[200]), .LWORD_REG_5_(vec[199]), .LWORD_REG_4_(vec[198]), .LWORD_REG_3_(vec[197]), .LWORD_REG_2_(vec[196]), .LWORD_REG_1_(vec[195]), .LWORD_REG_0_(vec[194]), .UWORD_REG_14_(vec[193]), .UWORD_REG_13_(vec[192]), .UWORD_REG_12_(vec[191]), .UWORD_REG_11_(vec[190]), .UWORD_REG_10_(vec[189]), .UWORD_REG_9_(vec[188]), .UWORD_REG_8_(vec[187]), .UWORD_REG_7_(vec[186]), .UWORD_REG_6_(vec[185]), .UWORD_REG_5_(vec[184]), .UWORD_REG_4_(vec[183]), .UWORD_REG_3_(vec[182]), .UWORD_REG_2_(vec[181]), .UWORD_REG_1_(vec[180]), .UWORD_REG_0_(vec[179]), .DATAO_REG_0__EXTRA(vec[178]), .DATAO_REG_1__EXTRA(vec[177]), .DATAO_REG_2__EXTRA(vec[176]), .DATAO_REG_3__EXTRA(vec[175]), .DATAO_REG_4__EXTRA(vec[174]), .DATAO_REG_5__EXTRA(vec[173]), .DATAO_REG_6__EXTRA(vec[172]), .DATAO_REG_7__EXTRA(vec[171]), .DATAO_REG_8__EXTRA(vec[170]), .DATAO_REG_9__EXTRA(vec[169]), .DATAO_REG_10__EXTRA(vec[168]), .DATAO_REG_11__EXTRA(vec[167]), .DATAO_REG_12__EXTRA(vec[166]), .DATAO_REG_13__EXTRA(vec[165]), .DATAO_REG_14__EXTRA(vec[164]), .DATAO_REG_15__EXTRA(vec[163]), .DATAO_REG_16__EXTRA(vec[162]), .DATAO_REG_17__EXTRA(vec[161]), .DATAO_REG_18__EXTRA(vec[160]), .DATAO_REG_19__EXTRA(vec[159]), .DATAO_REG_20__EXTRA(vec[158]), .DATAO_REG_21__EXTRA(vec[157]), .DATAO_REG_22__EXTRA(vec[156]), .DATAO_REG_23__EXTRA(vec[155]), .DATAO_REG_24__EXTRA(vec[154]), .DATAO_REG_25__EXTRA(vec[153]), .DATAO_REG_26__EXTRA(vec[152]), .DATAO_REG_27__EXTRA(vec[151]), .DATAO_REG_28__EXTRA(vec[150]), .DATAO_REG_29__EXTRA(vec[149]), .DATAO_REG_30__EXTRA(vec[148]), .DATAO_REG_31__EXTRA(vec[147]), .EAX_REG_0_(vec[146]), .EAX_REG_1_(vec[145]), .EAX_REG_2_(vec[144]), .EAX_REG_3_(vec[143]), .EAX_REG_4_(vec[142]), .EAX_REG_5_(vec[141]), .EAX_REG_6_(vec[140]), .EAX_REG_7_(vec[139]), .EAX_REG_8_(vec[138]), .EAX_REG_9_(vec[137]), .EAX_REG_10_(vec[136]), .EAX_REG_11_(vec[135]), .EAX_REG_12_(vec[134]), .EAX_REG_13_(vec[133]), .EAX_REG_14_(vec[132]), .EAX_REG_15_(vec[131]), .EAX_REG_16_(vec[130]), .EAX_REG_17_(vec[129]), .EAX_REG_18_(vec[128]), .EAX_REG_19_(vec[127]), .EAX_REG_20_(vec[126]), .EAX_REG_21_(vec[125]), .EAX_REG_22_(vec[124]), .EAX_REG_23_(vec[123]), .EAX_REG_24_(vec[122]), .EAX_REG_25_(vec[121]), .EAX_REG_26_(vec[120]), .EAX_REG_27_(vec[119]), .EAX_REG_28_(vec[118]), .EAX_REG_29_(vec[117]), .EAX_REG_30_(vec[116]), .EAX_REG_31_(vec[115]), .EBX_REG_0_(vec[114]), .EBX_REG_1_(vec[113]), .EBX_REG_2_(vec[112]), .EBX_REG_3_(vec[111]), .EBX_REG_4_(vec[110]), .EBX_REG_5_(vec[109]), .EBX_REG_6_(vec[108]), .EBX_REG_7_(vec[107]), .EBX_REG_8_(vec[106]), .EBX_REG_9_(vec[105]), .EBX_REG_10_(vec[104]), .EBX_REG_11_(vec[103]), .EBX_REG_12_(vec[102]), .EBX_REG_13_(vec[101]), .EBX_REG_14_(vec[100]), .EBX_REG_15_(vec[99]), .EBX_REG_16_(vec[98]), .EBX_REG_17_(vec[97]), .EBX_REG_18_(vec[96]), .EBX_REG_19_(vec[95]), .EBX_REG_20_(vec[94]), .EBX_REG_21_(vec[93]), .EBX_REG_22_(vec[92]), .EBX_REG_23_(vec[91]), .EBX_REG_24_(vec[90]), .EBX_REG_25_(vec[89]), .EBX_REG_26_(vec[88]), .EBX_REG_27_(vec[87]), .EBX_REG_28_(vec[86]), .EBX_REG_29_(vec[85]), .EBX_REG_30_(vec[84]), .EBX_REG_31_(vec[83]), .REIP_REG_0_(vec[82]), .REIP_REG_1_(vec[81]), .REIP_REG_2_(vec[80]), .REIP_REG_3_(vec[79]), .REIP_REG_4_(vec[78]), .REIP_REG_5_(vec[77]), .REIP_REG_6_(vec[76]), .REIP_REG_7_(vec[75]), .REIP_REG_8_(vec[74]), .REIP_REG_9_(vec[73]), .REIP_REG_10_(vec[72]), .REIP_REG_11_(vec[71]), .REIP_REG_12_(vec[70]), .REIP_REG_13_(vec[69]), .REIP_REG_14_(vec[68]), .REIP_REG_15_(vec[67]), .REIP_REG_16_(vec[66]), .REIP_REG_17_(vec[65]), .REIP_REG_18_(vec[64]), .REIP_REG_19_(vec[63]), .REIP_REG_20_(vec[62]), .REIP_REG_21_(vec[61]), .REIP_REG_22_(vec[60]), .REIP_REG_23_(vec[59]), .REIP_REG_24_(vec[58]), .REIP_REG_25_(vec[57]), .REIP_REG_26_(vec[56]), .REIP_REG_27_(vec[55]), .REIP_REG_28_(vec[54]), .REIP_REG_29_(vec[53]), .REIP_REG_30_(vec[52]), .REIP_REG_31_(vec[51]), .BYTEENABLE_REG_3_(vec[50]), .BYTEENABLE_REG_2_(vec[49]), .BYTEENABLE_REG_1_(vec[48]), .BYTEENABLE_REG_0_(vec[47]), .W_R_N_REG_EXTRA(vec[46]), .FLUSH_REG(vec[45]), .MORE_REG(vec[44]), .STATEBS16_REG(vec[43]), .REQUESTPENDING_REG(vec[42]), .D_C_N_REG_EXTRA(vec[41]), .M_IO_N_REG_EXTRA(vec[40]), .CODEFETCH_REG(vec[39]), .ADS_N_REG_EXTRA(vec[38]), .READREQUEST_REG(vec[37]), .MEMORYFETCH_REG(vec[36]), .DATAI_31_(vec[35]), .DATAI_30_(vec[34]), .DATAI_29_(vec[33]), .DATAI_28_(vec[32]), .DATAI_27_(vec[31]), .DATAI_26_(vec[30]), .DATAI_25_(vec[29]), .DATAI_24_(vec[28]), .DATAI_23_(vec[27]), .DATAI_22_(vec[26]), .DATAI_21_(vec[25]), .DATAI_20_(vec[24]), .DATAI_19_(vec[23]), .DATAI_18_(vec[22]), .DATAI_17_(vec[21]), .DATAI_16_(vec[20]), .DATAI_15_(vec[19]), .DATAI_14_(vec[18]), .DATAI_13_(vec[17]), .DATAI_12_(vec[16]), .DATAI_11_(vec[15]), .DATAI_10_(vec[14]), .DATAI_9_(vec[13]), .DATAI_8_(vec[12]), .DATAI_7_(vec[11]), .DATAI_6_(vec[10]), .DATAI_5_(vec[9]), .DATAI_4_(vec[8]), .DATAI_3_(vec[7]), .DATAI_2_(vec[6]), .DATAI_1_(vec[5]), .DATAI_0_(vec[4]), .NA_N(vec[3]), .BS16_N(vec[2]), .READY_N(vec[1]), .HOLD(vec[0]), .U3445(u3445), .U3446(u3446), .U3447(u3447), .U3448(u3448), .U3213(u3213), .U3212(u3212), .U3211(u3211), .U3210(u3210), .U3209(u3209), .U3208(u3208), .U3207(u3207), .U3206(u3206), .U3205(u3205), .U3204(u3204), .U3203(u3203), .U3202(u3202), .U3201(u3201), .U3200(u3200), .U3199(u3199), .U3198(u3198), .U3197(u3197), .U3196(u3196), .U3195(u3195), .U3194(u3194), .U3193(u3193), .U3192(u3192), .U3191(u3191), .U3190(u3190), .U3189(u3189), .U3188(u3188), .U3187(u3187), .U3186(u3186), .U3185(u3185), .U3184(u3184), .U3183(u3183), .U3182(u3182), .U3181(u3181), .U3451(u3451), .U3452(u3452), .U3180(u3180), .U3179(u3179), .U3178(u3178), .U3177(u3177), .U3176(u3176), .U3175(u3175), .U3174(u3174), .U3173(u3173), .U3172(u3172), .U3171(u3171), .U3170(u3170), .U3169(u3169), .U3168(u3168), .U3167(u3167), .U3166(u3166), .U3165(u3165), .U3164(u3164), .U3163(u3163), .U3162(u3162), .U3161(u3161), .U3160(u3160), .U3159(u3159), .U3158(u3158), .U3157(u3157), .U3156(u3156), .U3155(u3155), .U3154(u3154), .U3153(u3153), .U3152(u3152), .U3151(u3151), .U3453(u3453), .U3150(u3150), .U3149(u3149), .U3148(u3148), .U3147(u3147), .U3146(u3146), .U3145(u3145), .U3144(u3144), .U3143(u3143), .U3142(u3142), .U3141(u3141), .U3140(u3140), .U3139(u3139), .U3138(u3138), .U3137(u3137), .U3136(u3136), .U3135(u3135), .U3134(u3134), .U3133(u3133), .U3132(u3132), .U3131(u3131), .U3130(u3130), .U3129(u3129), .U3128(u3128), .U3127(u3127), .U3126(u3126), .U3125(u3125), .U3124(u3124), .U3123(u3123), .U3122(u3122), .U3121(u3121), .U3120(u3120), .U3119(u3119), .U3118(u3118), .U3117(u3117), .U3116(u3116), .U3115(u3115), .U3114(u3114), .U3113(u3113), .U3112(u3112), .U3111(u3111), .U3110(u3110), .U3109(u3109), .U3108(u3108), .U3107(u3107), .U3106(u3106), .U3105(u3105), .U3104(u3104), .U3103(u3103), .U3102(u3102), .U3101(u3101), .U3100(u3100), .U3099(u3099), .U3098(u3098), .U3097(u3097), .U3096(u3096), .U3095(u3095), .U3094(u3094), .U3093(u3093), .U3092(u3092), .U3091(u3091), .U3090(u3090), .U3089(u3089), .U3088(u3088), .U3087(u3087), .U3086(u3086), .U3085(u3085), .U3084(u3084), .U3083(u3083), .U3082(u3082), .U3081(u3081), .U3080(u3080), .U3079(u3079), .U3078(u3078), .U3077(u3077), .U3076(u3076), .U3075(u3075), .U3074(u3074), .U3073(u3073), .U3072(u3072), .U3071(u3071), .U3070(u3070), .U3069(u3069), .U3068(u3068), .U3067(u3067), .U3066(u3066), .U3065(u3065), .U3064(u3064), .U3063(u3063), .U3062(u3062), .U3061(u3061), .U3060(u3060), .U3059(u3059), .U3058(u3058), .U3057(u3057), .U3056(u3056), .U3055(u3055), .U3054(u3054), .U3053(u3053), .U3052(u3052), .U3051(u3051), .U3050(u3050), .U3049(u3049), .U3048(u3048), .U3047(u3047), .U3046(u3046), .U3045(u3045), .U3044(u3044), .U3043(u3043), .U3042(u3042), .U3041(u3041), .U3040(u3040), .U3039(u3039), .U3038(u3038), .U3037(u3037), .U3036(u3036), .U3035(u3035), .U3034(u3034), .U3033(u3033), .U3032(u3032), .U3031(u3031), .U3030(u3030), .U3029(u3029), .U3028(u3028), .U3027(u3027), .U3026(u3026), .U3025(u3025), .U3024(u3024), .U3023(u3023), .U3022(u3022), .U3021(u3021), .U3020(u3020), .U3455(u3455), .U3456(u3456), .U3459(u3459), .U3460(u3460), .U3461(u3461), .U3019(u3019), .U3462(u3462), .U3463(u3463), .U3464(u3464), .U3465(u3465), .U3018(u3018), .U3017(u3017), .U3016(u3016), .U3015(u3015), .U3014(u3014), .U3013(u3013), .U3012(u3012), .U3011(u3011), .U3010(u3010), .U3009(u3009), .U3008(u3008), .U3007(u3007), .U3006(u3006), .U3005(u3005), .U3004(u3004), .U3003(u3003), .U3002(u3002), .U3001(u3001), .U3000(u3000), .U2999(u2999), .U2998(u2998), .U2997(u2997), .U2996(u2996), .U2995(u2995), .U2994(u2994), .U2993(u2993), .U2992(u2992), .U2991(u2991), .U2990(u2990), .U2989(u2989), .U2988(u2988), .U2987(u2987), .U2986(u2986), .U2985(u2985), .U2984(u2984), .U2983(u2983), .U2982(u2982), .U2981(u2981), .U2980(u2980), .U2979(u2979), .U2978(u2978), .U2977(u2977), .U2976(u2976), .U2975(u2975), .U2974(u2974), .U2973(u2973), .U2972(u2972), .U2971(u2971), .U2970(u2970), .U2969(u2969), .U2968(u2968), .U2967(u2967), .U2966(u2966), .U2965(u2965), .U2964(u2964), .U2963(u2963), .U2962(u2962), .U2961(u2961), .U2960(u2960), .U2959(u2959), .U2958(u2958), .U2957(u2957), .U2956(u2956), .U2955(u2955), .U2954(u2954), .U2953(u2953), .U2952(u2952), .U2951(u2951), .U2950(u2950), .U2949(u2949), .U2948(u2948), .U2947(u2947), .U2946(u2946), .U2945(u2945), .U2944(u2944), .U2943(u2943), .U2942(u2942), .U2941(u2941), .U2940(u2940), .U2939(u2939), .U2938(u2938), .U2937(u2937), .U2936(u2936), .U2935(u2935), .U2934(u2934), .U2933(u2933), .U2932(u2932), .U2931(u2931), .U2930(u2930), .U2929(u2929), .U2928(u2928), .U2927(u2927), .U2926(u2926), .U2925(u2925), .U2924(u2924), .U2923(u2923), .U2922(u2922), .U2921(u2921), .U2920(u2920), .U2919(u2919), .U2918(u2918), .U2917(u2917), .U2916(u2916), .U2915(u2915), .U2914(u2914), .U2913(u2913), .U2912(u2912), .U2911(u2911), .U2910(u2910), .U2909(u2909), .U2908(u2908), .U2907(u2907), .U2906(u2906), .U2905(u2905), .U2904(u2904), .U2903(u2903), .U2902(u2902), .U2901(u2901), .U2900(u2900), .U2899(u2899), .U2898(u2898), .U2897(u2897), .U2896(u2896), .U2895(u2895), .U2894(u2894), .U2893(u2893), .U2892(u2892), .U2891(u2891), .U2890(u2890), .U2889(u2889), .U2888(u2888), .U2887(u2887), .U2886(u2886), .U2885(u2885), .U2884(u2884), .U2883(u2883), .U2882(u2882), .U2881(u2881), .U2880(u2880), .U2879(u2879), .U2878(u2878), .U2877(u2877), .U2876(u2876), .U2875(u2875), .U2874(u2874), .U2873(u2873), .U2872(u2872), .U2871(u2871), .U2870(u2870), .U2869(u2869), .U2868(u2868), .U2867(u2867), .U2866(u2866), .U2865(u2865), .U2864(u2864), .U2863(u2863), .U2862(u2862), .U2861(u2861), .U2860(u2860), .U2859(u2859), .U2858(u2858), .U2857(u2857), .U2856(u2856), .U2855(u2855), .U2854(u2854), .U2853(u2853), .U2852(u2852), .U2851(u2851), .U2850(u2850), .U2849(u2849), .U2848(u2848), .U2847(u2847), .U2846(u2846), .U2845(u2845), .U2844(u2844), .U2843(u2843), .U2842(u2842), .U2841(u2841), .U2840(u2840), .U2839(u2839), .U2838(u2838), .U2837(u2837), .U2836(u2836), .U2835(u2835), .U2834(u2834), .U2833(u2833), .U2832(u2832), .U2831(u2831), .U2830(u2830), .U2829(u2829), .U2828(u2828), .U2827(u2827), .U2826(u2826), .U2825(u2825), .U2824(u2824), .U2823(u2823), .U2822(u2822), .U2821(u2821), .U2820(u2820), .U2819(u2819), .U2818(u2818), .U2817(u2817), .U2816(u2816), .U2815(u2815), .U2814(u2814), .U2813(u2813), .U2812(u2812), .U2811(u2811), .U2810(u2810), .U2809(u2809), .U2808(u2808), .U2807(u2807), .U2806(u2806), .U2805(u2805), .U2804(u2804), .U2803(u2803), .U2802(u2802), .U2801(u2801), .U2800(u2800), .U2799(u2799), .U2798(u2798), .U2797(u2797), .U2796(u2796), .U2795(u2795), .U3468(u3468), .U2794(u2794), .U3469(u3469), .U3470(u3470), .U2793(u2793), .U3471(u3471), .U2792(u2792), .U3472(u3472), .U2791(u2791), .U3473(u3473), .U2790(u2790), .U2789(u2789), .U3474(u3474), .U2788(u2788), .BE_N_REG_3_(be_n_reg_3_), .BE_N_REG_2_(be_n_reg_2_), .BE_N_REG_1_(be_n_reg_1_), .BE_N_REG_0_(be_n_reg_0_), .ADDRESS_REG_29_(address_reg_29_), .ADDRESS_REG_28_(address_reg_28_), .ADDRESS_REG_27_(address_reg_27_), .ADDRESS_REG_26_(address_reg_26_), .ADDRESS_REG_25_(address_reg_25_), .ADDRESS_REG_24_(address_reg_24_), .ADDRESS_REG_23_(address_reg_23_), .ADDRESS_REG_22_(address_reg_22_), .ADDRESS_REG_21_(address_reg_21_), .ADDRESS_REG_20_(address_reg_20_), .ADDRESS_REG_19_(address_reg_19_), .ADDRESS_REG_18_(address_reg_18_), .ADDRESS_REG_17_(address_reg_17_), .ADDRESS_REG_16_(address_reg_16_), .ADDRESS_REG_15_(address_reg_15_), .ADDRESS_REG_14_(address_reg_14_), .ADDRESS_REG_13_(address_reg_13_), .ADDRESS_REG_12_(address_reg_12_), .ADDRESS_REG_11_(address_reg_11_), .ADDRESS_REG_10_(address_reg_10_), .ADDRESS_REG_9_(address_reg_9_), .ADDRESS_REG_8_(address_reg_8_), .ADDRESS_REG_7_(address_reg_7_), .ADDRESS_REG_6_(address_reg_6_), .ADDRESS_REG_5_(address_reg_5_), .ADDRESS_REG_4_(address_reg_4_), .ADDRESS_REG_3_(address_reg_3_), .ADDRESS_REG_2_(address_reg_2_), .ADDRESS_REG_1_(address_reg_1_), .ADDRESS_REG_0_(address_reg_0_), .W_R_N_REG(w_r_n_reg), .D_C_N_REG(d_c_n_reg), .M_IO_N_REG(m_io_n_reg), .ADS_N_REG(ads_n_reg), .DATAO_REG_31_(datao_reg_31_), .DATAO_REG_30_(datao_reg_30_), .DATAO_REG_29_(datao_reg_29_), .DATAO_REG_28_(datao_reg_28_), .DATAO_REG_27_(datao_reg_27_), .DATAO_REG_26_(datao_reg_26_), .DATAO_REG_25_(datao_reg_25_), .DATAO_REG_24_(datao_reg_24_), .DATAO_REG_23_(datao_reg_23_), .DATAO_REG_22_(datao_reg_22_), .DATAO_REG_21_(datao_reg_21_), .DATAO_REG_20_(datao_reg_20_), .DATAO_REG_19_(datao_reg_19_), .DATAO_REG_18_(datao_reg_18_), .DATAO_REG_17_(datao_reg_17_), .DATAO_REG_16_(datao_reg_16_), .DATAO_REG_15_(datao_reg_15_), .DATAO_REG_14_(datao_reg_14_), .DATAO_REG_13_(datao_reg_13_), .DATAO_REG_12_(datao_reg_12_), .DATAO_REG_11_(datao_reg_11_), .DATAO_REG_10_(datao_reg_10_), .DATAO_REG_9_(datao_reg_9_), .DATAO_REG_8_(datao_reg_8_), .DATAO_REG_7_(datao_reg_7_), .DATAO_REG_6_(datao_reg_6_), .DATAO_REG_5_(datao_reg_5_), .DATAO_REG_4_(datao_reg_4_), .DATAO_REG_3_(datao_reg_3_), .DATAO_REG_2_(datao_reg_2_), .DATAO_REG_1_(datao_reg_1_), .DATAO_REG_0_(datao_reg_0_));

integer i=0;
always @ (posedge clk) begin
	vec = input_vec_mem[i];
	$monitor(vec);
	i = i + 1;

end

always @ (negedge clk)begin
	$fdisplay ( fh_w, u3445, u3446, u3447, u3448, u3213, u3212, u3211, u3210, u3209, u3208, u3207, u3206, u3205, u3204, u3203, u3202, u3201, u3200, u3199, u3198, u3197, u3196, u3195, u3194, u3193, u3192, u3191, u3190, u3189, u3188, u3187, u3186, u3185, u3184, u3183, u3182, u3181, u3451, u3452, u3180, u3179, u3178, u3177, u3176, u3175, u3174, u3173, u3172, u3171, u3170, u3169, u3168, u3167, u3166, u3165, u3164, u3163, u3162, u3161, u3160, u3159, u3158, u3157, u3156, u3155, u3154, u3153, u3152, u3151, u3453, u3150, u3149, u3148, u3147, u3146, u3145, u3144, u3143, u3142, u3141, u3140, u3139, u3138, u3137, u3136, u3135, u3134, u3133, u3132, u3131, u3130, u3129, u3128, u3127, u3126, u3125, u3124, u3123, u3122, u3121, u3120, u3119, u3118, u3117, u3116, u3115, u3114, u3113, u3112, u3111, u3110, u3109, u3108, u3107, u3106, u3105, u3104, u3103, u3102, u3101, u3100, u3099, u3098, u3097, u3096, u3095, u3094, u3093, u3092, u3091, u3090, u3089, u3088, u3087, u3086, u3085, u3084, u3083, u3082, u3081, u3080, u3079, u3078, u3077, u3076, u3075, u3074, u3073, u3072, u3071, u3070, u3069, u3068, u3067, u3066, u3065, u3064, u3063, u3062, u3061, u3060, u3059, u3058, u3057, u3056, u3055, u3054, u3053, u3052, u3051, u3050, u3049, u3048, u3047, u3046, u3045, u3044, u3043, u3042, u3041, u3040, u3039, u3038, u3037, u3036, u3035, u3034, u3033, u3032, u3031, u3030, u3029, u3028, u3027, u3026, u3025, u3024, u3023, u3022, u3021, u3020, u3455, u3456, u3459, u3460, u3461, u3019, u3462, u3463, u3464, u3465, u3018, u3017, u3016, u3015, u3014, u3013, u3012, u3011, u3010, u3009, u3008, u3007, u3006, u3005, u3004, u3003, u3002, u3001, u3000, u2999, u2998, u2997, u2996, u2995, u2994, u2993, u2992, u2991, u2990, u2989, u2988, u2987, u2986, u2985, u2984, u2983, u2982, u2981, u2980, u2979, u2978, u2977, u2976, u2975, u2974, u2973, u2972, u2971, u2970, u2969, u2968, u2967, u2966, u2965, u2964, u2963, u2962, u2961, u2960, u2959, u2958, u2957, u2956, u2955, u2954, u2953, u2952, u2951, u2950, u2949, u2948, u2947, u2946, u2945, u2944, u2943, u2942, u2941, u2940, u2939, u2938, u2937, u2936, u2935, u2934, u2933, u2932, u2931, u2930, u2929, u2928, u2927, u2926, u2925, u2924, u2923, u2922, u2921, u2920, u2919, u2918, u2917, u2916, u2915, u2914, u2913, u2912, u2911, u2910, u2909, u2908, u2907, u2906, u2905, u2904, u2903, u2902, u2901, u2900, u2899, u2898, u2897, u2896, u2895, u2894, u2893, u2892, u2891, u2890, u2889, u2888, u2887, u2886, u2885, u2884, u2883, u2882, u2881, u2880, u2879, u2878, u2877, u2876, u2875, u2874, u2873, u2872, u2871, u2870, u2869, u2868, u2867, u2866, u2865, u2864, u2863, u2862, u2861, u2860, u2859, u2858, u2857, u2856, u2855, u2854, u2853, u2852, u2851, u2850, u2849, u2848, u2847, u2846, u2845, u2844, u2843, u2842, u2841, u2840, u2839, u2838, u2837, u2836, u2835, u2834, u2833, u2832, u2831, u2830, u2829, u2828, u2827, u2826, u2825, u2824, u2823, u2822, u2821, u2820, u2819, u2818, u2817, u2816, u2815, u2814, u2813, u2812, u2811, u2810, u2809, u2808, u2807, u2806, u2805, u2804, u2803, u2802, u2801, u2800, u2799, u2798, u2797, u2796, u2795, u3468, u2794, u3469, u3470, u2793, u3471, u2792, u3472, u2791, u3473, u2790, u2789, u3474, u2788, be_n_reg_3_, be_n_reg_2_, be_n_reg_1_, be_n_reg_0_, address_reg_29_, address_reg_28_, address_reg_27_, address_reg_26_, address_reg_25_, address_reg_24_, address_reg_23_, address_reg_22_, address_reg_21_, address_reg_20_, address_reg_19_, address_reg_18_, address_reg_17_, address_reg_16_, address_reg_15_, address_reg_14_, address_reg_13_, address_reg_12_, address_reg_11_, address_reg_10_, address_reg_9_, address_reg_8_, address_reg_7_, address_reg_6_, address_reg_5_, address_reg_4_, address_reg_3_, address_reg_2_, address_reg_1_, address_reg_0_, w_r_n_reg, d_c_n_reg, m_io_n_reg, ads_n_reg, datao_reg_31_, datao_reg_30_, datao_reg_29_, datao_reg_28_, datao_reg_27_, datao_reg_26_, datao_reg_25_, datao_reg_24_, datao_reg_23_, datao_reg_22_, datao_reg_21_, datao_reg_20_, datao_reg_19_, datao_reg_18_, datao_reg_17_, datao_reg_16_, datao_reg_15_, datao_reg_14_, datao_reg_13_, datao_reg_12_, datao_reg_11_, datao_reg_10_, datao_reg_9_, datao_reg_8_, datao_reg_7_, datao_reg_6_, datao_reg_5_, datao_reg_4_, datao_reg_3_, datao_reg_2_, datao_reg_1_, datao_reg_0_);
	if(i == vec_length)begin
		$finish;
	end
end

integer fh_w;
initial begin
	fh_w = $fopen(`out_file, "w");
end
 
initial begin
	//$fsdbDumpfile("SET.fsdb");
	//$fsdbDumpvars;
	//$fsdbDumpMDA;
	$dumpfile("test_result.vcd");
    $dumpvars;

end
endmodule
