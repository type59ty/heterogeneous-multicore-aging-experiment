// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module c499d (N11,  N15,  N19,  N113, N117, N121, N125, N129, N133, N137,
             N141, N145, N149, N153, N157, N161, N165, N169, N173, N177,
             N181, N185, N189, N193, N197, N1101,N1105,N1109,N1113,N1117,
             N1121,N1125,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,
             N1137,N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,
             N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,
             N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,
             N1753,N1754,N1755,
             N21,  N25,  N29,  N213, N217, N221, N225, N229, N233, N237,
             N241, N245, N249, N253, N257, N261, N265, N269, N273, N277,
             N281, N285, N289, N293, N297, N2101,N2105,N2109,N2113,N2117,
             N2121,N2125,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,
             N2137,N2724,N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,
             N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,
             N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,
             N2753,N2754,N2755);

input N11,N15,N19,N113,N117,N121,N125,N129,N133,N137,
      N141,N145,N149,N153,N157,N161,N165,N169,N173,N177,
      N181,N185,N189,N193,N197,N1101,N1105,N1109,N1113,N1117,
      N1121,N1125,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,
      N1137,
      N21,N25,N29,N213,N217,N221,N225,N229,N233,N237,
      N241,N245,N249,N253,N257,N261,N265,N269,N273,N277,
      N281,N285,N289,N293,N297,N2101,N2105,N2109,N2113,N2117,
      N2121,N2125,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,
      N2137;

output N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,
       N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,
       N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,
       N1754,N1755,
       N2724,N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,
       N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,
       N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,
       N2754,N2755;

wire N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,
     N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,
     N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,
     N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
     N1290,N1293,N1296,N1299,N1302,N1305,N1308,N1311,N1314,N1315,
     N1316,N1317,N1318,N1319,N1320,N1321,N1338,N1339,N1340,N1341,
     N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,
     N1352,N1353,N1354,N1367,N1380,N1393,N1406,N1419,N1432,N1445,
     N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,
     N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,
     N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,
     N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,
     N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1607,
     N1620,N1625,N1630,N1635,N1640,N1645,N1650,N1655,N1692,N1693,
     N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,
     N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,
     N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,

     N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,
     N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,
     N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278,N2279,
     N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,
     N2290,N2293,N2296,N2299,N2302,N2305,N2308,N2311,N2314,N2315,
     N2316,N2317,N2318,N2319,N2320,N2321,N2338,N2339,N2340,N2341,
     N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,
     N2352,N2353,N2354,N2367,N2380,N2393,N2406,N2419,N2432,N2445,
     N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,
     N2564,N2565,N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,
     N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,
     N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,
     N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2607,
     N2620,N2625,N2630,N2635,N2640,N2645,N2650,N2655,N2692,N2693,
     N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,
     N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,
     N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723;

xor XOR2_11 (N1250, N11, N15);
xor XOR2_12 (N1251, N19, N113);
xor XOR2_13 (N1252, N117, N121);
xor XOR2_14 (N1253, N125, N129);
xor XOR2_15 (N1254, N133, N137);
xor XOR2_16 (N1255, N141, N145);
xor XOR2_17 (N1256, N149, N153);
xor XOR2_18 (N1257, N157, N161);
xor XOR2_19 (N1258, N165, N169);
xor XOR2_110 (N1259, N173, N177);
xor XOR2_111 (N1260, N181, N185);
xor XOR2_112 (N1261, N189, N193);
xor XOR2_113 (N1262, N197, N1101);
xor XOR2_114 (N1263, N1105, N1109);
xor XOR2_115 (N1264, N1113, N1117);
xor XOR2_116 (N1265, N1121, N1125);
and AND2_117 (N1266, N1129, N1137);
and AND2_118 (N1267, N1130, N1137);
and AND2_119 (N1268, N1131, N1137);
and AND2_120 (N1269, N1132, N1137);
and AND2_121 (N1270, N1133, N1137);
and AND2_122 (N1271, N1134, N1137);
and AND2_123 (N1272, N1135, N1137);
and AND2_124 (N1273, N1136, N1137);
xor XOR2_125 (N1274, N11, N117);
xor XOR2_126 (N1275, N133, N149);
xor XOR2_127 (N1276, N15, N121);
xor XOR2_128 (N1277, N137, N153);
xor XOR2_129 (N1278, N19, N125);
xor XOR2_130 (N1279, N141, N157);
xor XOR2_131 (N1280, N113, N129);
xor XOR2_132 (N1281, N145, N161);
xor XOR2_133 (N1282, N165, N181);
xor XOR2_134 (N1283, N197, N1113);
xor XOR2_135 (N1284, N169, N185);
xor XOR2_136 (N1285, N1101, N1117);
xor XOR2_137 (N1286, N173, N189);
xor XOR2_138 (N1287, N1105, N1121);
xor XOR2_139 (N1288, N177, N193);
xor XOR2_140 (N1289, N1109, N1125);
xor XOR2_141 (N1290, N1250, N1251);
xor XOR2_142 (N1293, N1252, N1253);
xor XOR2_143 (N1296, N1254, N1255);
xor XOR2_144 (N1299, N1256, N1257);
xor XOR2_145 (N1302, N1258, N1259);
xor XOR2_146 (N1305, N1260, N1261);
xor XOR2_147 (N1308, N1262, N1263);
xor XOR2_148 (N1311, N1264, N1265);
xor XOR2_149 (N1314, N1274, N1275);
xor XOR2_150 (N1315, N1276, N1277);
xor XOR2_151 (N1316, N1278, N1279);
xor XOR2_152 (N1317, N1280, N1281);
xor XOR2_153 (N1318, N1282, N1283);
xor XOR2_154 (N1319, N1284, N1285);
xor XOR2_155 (N1320, N1286, N1287);
xor XOR2_156 (N1321, N1288, N1289);
xor XOR2_157 (N1338, N1290, N1293);
xor XOR2_158 (N1339, N1296, N1299);
xor XOR2_159 (N1340, N1290, N1296);
xor XOR2_160 (N1341, N1293, N1299);
xor XOR2_161 (N1342, N1302, N1305);
xor XOR2_162 (N1343, N1308, N1311);
xor XOR2_163 (N1344, N1302, N1308);
xor XOR2_164 (N1345, N1305, N1311);
xor XOR2_165 (N1346, N1266, N1342);
xor XOR2_166 (N1347, N1267, N1343);
xor XOR2_167 (N1348, N1268, N1344);
xor XOR2_168 (N1349, N1269, N1345);
xor XOR2_169 (N1350, N1270, N1338);
xor XOR2_170 (N1351, N1271, N1339);
xor XOR2_171 (N1352, N1272, N1340);
xor XOR2_172 (N1353, N1273, N1341);
xor XOR2_173 (N1354, N1314, N1346);
xor XOR2_174 (N1367, N1315, N1347);
xor XOR2_175 (N1380, N1316, N1348);
xor XOR2_176 (N1393, N1317, N1349);
xor XOR2_177 (N1406, N1318, N1350);
xor XOR2_178 (N1419, N1319, N1351);
xor XOR2_179 (N1432, N1320, N1352);
xor XOR2_180 (N1445, N1321, N1353);
not NOT1_181 (N1554, N1354);
not NOT1_182 (N1555, N1367);
not NOT1_183 (N1556, N1380);
not NOT1_184 (N1557, N1354);
not NOT1_185 (N1558, N1367);
not NOT1_186 (N1559, N1393);
not NOT1_187 (N1560, N1354);
not NOT1_188 (N1561, N1380);
not NOT1_189 (N1562, N1393);
not NOT1_190 (N1563, N1367);
not NOT1_191 (N1564, N1380);
not NOT1_192 (N1565, N1393);
not NOT1_193 (N1566, N1419);
not NOT1_194 (N1567, N1445);
not NOT1_195 (N1568, N1419);
not NOT1_196 (N1569, N1432);
not NOT1_197 (N1570, N1406);
not NOT1_198 (N1571, N1445);
not NOT1_199 (N1572, N1406);
not NOT1_1100 (N1573, N1432);
not NOT1_1101 (N1574, N1406);
not NOT1_1102 (N1575, N1419);
not NOT1_1103 (N1576, N1432);
not NOT1_1104 (N1577, N1406);
not NOT1_1105 (N1578, N1419);
not NOT1_1106 (N1579, N1445);
not NOT1_1107 (N1580, N1406);
not NOT1_1108 (N1581, N1432);
not NOT1_1109 (N1582, N1445);
not NOT1_1110 (N1583, N1419);
not NOT1_1111 (N1584, N1432);
not NOT1_1112 (N1585, N1445);
not NOT1_1113 (N1586, N1367);
not NOT1_1114 (N1587, N1393);
not NOT1_1115 (N1588, N1367);
not NOT1_1116 (N1589, N1380);
not NOT1_1117 (N1590, N1354);
not NOT1_1118 (N1591, N1393);
not NOT1_1119 (N1592, N1354);
not NOT1_1120 (N1593, N1380);
and AND4_1121 (N1594, N1554, N1555, N1556, N1393);
and AND4_1122 (N1595, N1557, N1558, N1380, N1559);
and AND4_1123 (N1596, N1560, N1367, N1561, N1562);
and AND4_1124 (N1597, N1354, N1563, N1564, N1565);
and AND4_1125 (N1598, N1574, N1575, N1576, N1445);
and AND4_1126 (N1599, N1577, N1578, N1432, N1579);
and AND4_1127 (N1600, N1580, N1419, N1581, N1582);
and AND4_1128 (N1601, N1406, N1583, N1584, N1585);
or OR4_1129 (N1602, N1594, N1595, N1596, N1597);
or OR4_1130 (N1607, N1598, N1599, N1600, N1601);
and AND5_1131 (N1620, N1406, N1566, N1432, N1567, N1602);
and AND5_1132 (N1625, N1406, N1568, N1569, N1445, N1602);
and AND5_1133 (N1630, N1570, N1419, N1432, N1571, N1602);
and AND5_1134 (N1635, N1572, N1419, N1573, N1445, N1602);
and AND5_1135 (N1640, N1354, N1586, N1380, N1587, N1607);
and AND5_1136 (N1645, N1354, N1588, N1589, N1393, N1607);
and AND5_1137 (N1650, N1590, N1367, N1380, N1591, N1607);
and AND5_1138 (N1655, N1592, N1367, N1593, N1393, N1607);
and AND2_1139 (N1692, N1354, N1620);
and AND2_1140 (N1693, N1367, N1620);
and AND2_1141 (N1694, N1380, N1620);
and AND2_1142 (N1695, N1393, N1620);
and AND2_1143 (N1696, N1354, N1625);
and AND2_1144 (N1697, N1367, N1625);
and AND2_1145 (N1698, N1380, N1625);
and AND2_1146 (N1699, N1393, N1625);
and AND2_1147 (N1700, N1354, N1630);
and AND2_1148 (N1701, N1367, N1630);
and AND2_1149 (N1702, N1380, N1630);
and AND2_1150 (N1703, N1393, N1630);
and AND2_1151 (N1704, N1354, N1635);
and AND2_1152 (N1705, N1367, N1635);
and AND2_1153 (N1706, N1380, N1635);
and AND2_1154 (N1707, N1393, N1635);
and AND2_1155 (N1708, N1406, N1640);
and AND2_1156 (N1709, N1419, N1640);
and AND2_1157 (N1710, N1432, N1640);
and AND2_1158 (N1711, N1445, N1640);
and AND2_1159 (N1712, N1406, N1645);
and AND2_1160 (N1713, N1419, N1645);
and AND2_1161 (N1714, N1432, N1645);
and AND2_1162 (N1715, N1445, N1645);
and AND2_1163 (N1716, N1406, N1650);
and AND2_1164 (N1717, N1419, N1650);
and AND2_1165 (N1718, N1432, N1650);
and AND2_1166 (N1719, N1445, N1650);
and AND2_1167 (N1720, N1406, N1655);
and AND2_1168 (N1721, N1419, N1655);
and AND2_1169 (N1722, N1432, N1655);
and AND2_1170 (N1723, N1445, N1655);
xor XOR2_1171 (N1724, N11, N1692);
xor XOR2_1172 (N1725, N15, N1693);
xor XOR2_1173 (N1726, N19, N1694);
xor XOR2_1174 (N1727, N113, N1695);
xor XOR2_1175 (N1728, N117, N1696);
xor XOR2_1176 (N1729, N121, N1697);
xor XOR2_1177 (N1730, N125, N1698);
xor XOR2_1178 (N1731, N129, N1699);
xor XOR2_1179 (N1732, N133, N1700);
xor XOR2_1180 (N1733, N137, N1701);
xor XOR2_1181 (N1734, N141, N1702);
xor XOR2_1182 (N1735, N145, N1703);
xor XOR2_1183 (N1736, N149, N1704);
xor XOR2_1184 (N1737, N153, N1705);
xor XOR2_1185 (N1738, N157, N1706);
xor XOR2_1186 (N1739, N161, N1707);
xor XOR2_1187 (N1740, N165, N1708);
xor XOR2_1188 (N1741, N169, N1709);
xor XOR2_1189 (N1742, N173, N1710);
xor XOR2_1190 (N1743, N177, N1711);
xor XOR2_1191 (N1744, N181, N1712);
xor XOR2_1192 (N1745, N185, N1713);
xor XOR2_1193 (N1746, N189, N1714);
xor XOR2_1194 (N1747, N193, N1715);
xor XOR2_1195 (N1748, N197, N1716);
xor XOR2_1196 (N1749, N1101, N1717);
xor XOR2_1197 (N1750, N1105, N1718);
xor XOR2_1198 (N1751, N1109, N1719);
xor XOR2_1199 (N1752, N1113, N1720);
xor XOR2_1200 (N1753, N1117, N1721);
xor XOR2_1201 (N1754, N1121, N1722);
xor XOR2_1202 (N1755, N1125, N1723);

xor XOR2_21 (N2250, N21, N25);
xor XOR2_22 (N2251, N29, N213);
xor XOR2_23 (N2252, N217, N221);
xor XOR2_24 (N2253, N225, N229);
xor XOR2_25 (N2254, N233, N237);
xor XOR2_26 (N2255, N241, N245);
xor XOR2_27 (N2256, N249, N253);
xor XOR2_28 (N2257, N257, N261);
xor XOR2_29 (N2258, N265, N269);
xor XOR2_210 (N2259, N273, N277);
xor XOR2_211 (N2260, N281, N285);
xor XOR2_212 (N2261, N289, N293);
xor XOR2_213 (N2262, N297, N2101);
xor XOR2_214 (N2263, N2105, N2109);
xor XOR2_215 (N2264, N2113, N2117);
xor XOR2_216 (N2265, N2121, N2125);
and AND2_217 (N2266, N2129, N2137);
and AND2_218 (N2267, N2130, N2137);
and AND2_219 (N2268, N2131, N2137);
and AND2_220 (N2269, N2132, N2137);
and AND2_221 (N2270, N2133, N2137);
and AND2_222 (N2271, N2134, N2137);
and AND2_223 (N2272, N2135, N2137);
and AND2_224 (N2273, N2136, N2137);
xor XOR2_225 (N2274, N21, N217);
xor XOR2_226 (N2275, N233, N249);
xor XOR2_227 (N2276, N25, N221);
xor XOR2_228 (N2277, N237, N253);
xor XOR2_229 (N2278, N29, N225);
xor XOR2_230 (N2279, N241, N257);
xor XOR2_231 (N2280, N213, N229);
xor XOR2_232 (N2281, N245, N261);
xor XOR2_233 (N2282, N265, N281);
xor XOR2_234 (N2283, N297, N2113);
xor XOR2_235 (N2284, N269, N285);
xor XOR2_236 (N2285, N2101, N2117);
xor XOR2_237 (N2286, N273, N289);
xor XOR2_238 (N2287, N2105, N2121);
xor XOR2_239 (N2288, N277, N293);
xor XOR2_240 (N2289, N2109, N2125);
xor XOR2_241 (N2290, N2250, N2251);
xor XOR2_242 (N2293, N2252, N2253);
xor XOR2_243 (N2296, N2254, N2255);
xor XOR2_244 (N2299, N2256, N2257);
xor XOR2_245 (N2302, N2258, N2259);
xor XOR2_246 (N2305, N2260, N2261);
xor XOR2_247 (N2308, N2262, N2263);
xor XOR2_248 (N2311, N2264, N2265);
xor XOR2_249 (N2314, N2274, N2275);
xor XOR2_250 (N2315, N2276, N2277);
xor XOR2_251 (N2316, N2278, N2279);
xor XOR2_252 (N2317, N2280, N2281);
xor XOR2_253 (N2318, N2282, N2283);
xor XOR2_254 (N2319, N2284, N2285);
xor XOR2_255 (N2320, N2286, N2287);
xor XOR2_256 (N2321, N2288, N2289);
xor XOR2_257 (N2338, N2290, N2293);
xor XOR2_258 (N2339, N2296, N2299);
xor XOR2_259 (N2340, N2290, N2296);
xor XOR2_260 (N2341, N2293, N2299);
xor XOR2_261 (N2342, N2302, N2305);
xor XOR2_262 (N2343, N2308, N2311);
xor XOR2_263 (N2344, N2302, N2308);
xor XOR2_264 (N2345, N2305, N2311);
xor XOR2_265 (N2346, N2266, N2342);
xor XOR2_266 (N2347, N2267, N2343);
xor XOR2_267 (N2348, N2268, N2344);
xor XOR2_268 (N2349, N2269, N2345);
xor XOR2_269 (N2350, N2270, N2338);
xor XOR2_270 (N2351, N2271, N2339);
xor XOR2_271 (N2352, N2272, N2340);
xor XOR2_272 (N2353, N2273, N2341);
xor XOR2_273 (N2354, N2314, N2346);
xor XOR2_274 (N2367, N2315, N2347);
xor XOR2_275 (N2380, N2316, N2348);
xor XOR2_276 (N2393, N2317, N2349);
xor XOR2_277 (N2406, N2318, N2350);
xor XOR2_278 (N2419, N2319, N2351);
xor XOR2_279 (N2432, N2320, N2352);
xor XOR2_280 (N2445, N2321, N2353);
not NOT1_281 (N2554, N2354);
not NOT1_282 (N2555, N2367);
not NOT1_283 (N2556, N2380);
not NOT1_284 (N2557, N2354);
not NOT1_285 (N2558, N2367);
not NOT1_286 (N2559, N2393);
not NOT1_287 (N2560, N2354);
not NOT1_288 (N2561, N2380);
not NOT1_289 (N2562, N2393);
not NOT1_290 (N2563, N2367);
not NOT1_291 (N2564, N2380);
not NOT1_292 (N2565, N2393);
not NOT1_293 (N2566, N2419);
not NOT1_294 (N2567, N2445);
not NOT1_295 (N2568, N2419);
not NOT1_296 (N2569, N2432);
not NOT1_297 (N2570, N2406);
not NOT1_298 (N2571, N2445);
not NOT1_299 (N2572, N2406);
not NOT1_2100 (N2573, N2432);
not NOT1_2101 (N2574, N2406);
not NOT1_2102 (N2575, N2419);
not NOT1_2103 (N2576, N2432);
not NOT1_2104 (N2577, N2406);
not NOT1_2105 (N2578, N2419);
not NOT1_2106 (N2579, N2445);
not NOT1_2107 (N2580, N2406);
not NOT1_2108 (N2581, N2432);
not NOT1_2109 (N2582, N2445);
not NOT1_2110 (N2583, N2419);
not NOT1_2111 (N2584, N2432);
not NOT1_2112 (N2585, N2445);
not NOT1_2113 (N2586, N2367);
not NOT1_2114 (N2587, N2393);
not NOT1_2115 (N2588, N2367);
not NOT1_2116 (N2589, N2380);
not NOT1_2117 (N2590, N2354);
not NOT1_2118 (N2591, N2393);
not NOT1_2119 (N2592, N2354);
not NOT1_2120 (N2593, N2380);
and AND4_2121 (N2594, N2554, N2555, N2556, N2393);
and AND4_2122 (N2595, N2557, N2558, N2380, N2559);
and AND4_2123 (N2596, N2560, N2367, N2561, N2562);
and AND4_2124 (N2597, N2354, N2563, N2564, N2565);
and AND4_2125 (N2598, N2574, N2575, N2576, N2445);
and AND4_2126 (N2599, N2577, N2578, N2432, N2579);
and AND4_2127 (N2600, N2580, N2419, N2581, N2582);
and AND4_2128 (N2601, N2406, N2583, N2584, N2585);
or OR4_2129 (N2602, N2594, N2595, N2596, N2597);
or OR4_2130 (N2607, N2598, N2599, N2600, N2601);
and AND5_2131 (N2620, N2406, N2566, N2432, N2567, N2602);
and AND5_2132 (N2625, N2406, N2568, N2569, N2445, N2602);
and AND5_2133 (N2630, N2570, N2419, N2432, N2571, N2602);
and AND5_2134 (N2635, N2572, N2419, N2573, N2445, N2602);
and AND5_2135 (N2640, N2354, N2586, N2380, N2587, N2607);
and AND5_2136 (N2645, N2354, N2588, N2589, N2393, N2607);
and AND5_2137 (N2650, N2590, N2367, N2380, N2591, N2607);
and AND5_2138 (N2655, N2592, N2367, N2593, N2393, N2607);
and AND2_2139 (N2692, N2354, N2620);
and AND2_2140 (N2693, N2367, N2620);
and AND2_2141 (N2694, N2380, N2620);
and AND2_2142 (N2695, N2393, N2620);
and AND2_2143 (N2696, N2354, N2625);
and AND2_2144 (N2697, N2367, N2625);
and AND2_2145 (N2698, N2380, N2625);
and AND2_2146 (N2699, N2393, N2625);
and AND2_2147 (N2700, N2354, N2630);
and AND2_2148 (N2701, N2367, N2630);
and AND2_2149 (N2702, N2380, N2630);
and AND2_2150 (N2703, N2393, N2630);
and AND2_2151 (N2704, N2354, N2635);
and AND2_2152 (N2705, N2367, N2635);
and AND2_2153 (N2706, N2380, N2635);
and AND2_2154 (N2707, N2393, N2635);
and AND2_2155 (N2708, N2406, N2640);
and AND2_2156 (N2709, N2419, N2640);
and AND2_2157 (N2710, N2432, N2640);
and AND2_2158 (N2711, N2445, N2640);
and AND2_2159 (N2712, N2406, N2645);
and AND2_2160 (N2713, N2419, N2645);
and AND2_2161 (N2714, N2432, N2645);
and AND2_2162 (N2715, N2445, N2645);
and AND2_2163 (N2716, N2406, N2650);
and AND2_2164 (N2717, N2419, N2650);
and AND2_2165 (N2718, N2432, N2650);
and AND2_2166 (N2719, N2445, N2650);
and AND2_2167 (N2720, N2406, N2655);
and AND2_2168 (N2721, N2419, N2655);
and AND2_2169 (N2722, N2432, N2655);
and AND2_2170 (N2723, N2445, N2655);
xor XOR2_2171 (N2724, N21, N2692);
xor XOR2_2172 (N2725, N25, N2693);
xor XOR2_2173 (N2726, N29, N2694);
xor XOR2_2174 (N2727, N213, N2695);
xor XOR2_2175 (N2728, N217, N2696);
xor XOR2_2176 (N2729, N221, N2697);
xor XOR2_2177 (N2730, N225, N2698);
xor XOR2_2178 (N2731, N229, N2699);
xor XOR2_2179 (N2732, N233, N2700);
xor XOR2_2180 (N2733, N237, N2701);
xor XOR2_2181 (N2734, N241, N2702);
xor XOR2_2182 (N2735, N245, N2703);
xor XOR2_2183 (N2736, N249, N2704);
xor XOR2_2184 (N2737, N253, N2705);
xor XOR2_2185 (N2738, N257, N2706);
xor XOR2_2186 (N2739, N261, N2707);
xor XOR2_2187 (N2740, N265, N2708);
xor XOR2_2188 (N2741, N269, N2709);
xor XOR2_2189 (N2742, N273, N2710);
xor XOR2_2190 (N2743, N277, N2711);
xor XOR2_2191 (N2744, N281, N2712);
xor XOR2_2192 (N2745, N285, N2713);
xor XOR2_2193 (N2746, N289, N2714);
xor XOR2_2194 (N2747, N293, N2715);
xor XOR2_2195 (N2748, N297, N2716);
xor XOR2_2196 (N2749, N2101, N2717);
xor XOR2_2197 (N2750, N2105, N2718);
xor XOR2_2198 (N2751, N2109, N2719);
xor XOR2_2199 (N2752, N2113, N2720);
xor XOR2_2200 (N2753, N2117, N2721);
xor XOR2_2201 (N2754, N2121, N2722);
xor XOR2_2202 (N2755, N2125, N2723);

endmodule
