`timescale 1ns/10ps

`define cycle 10.0
`define terminate_cycle 400000//200000 // Modify your terminate ycle here

module b14_ras_testfixture;

`define in_file "b14_ras/rand_input_vector_b14_ras_0.out"
`define out_file "b14_ras/rand_output_vector_b14_ras_0.out"

parameter vec_width = 277;
parameter vec_length = 2;

reg clk = 0;


reg [vec_width-1:0] input_vec_mem [0:vec_length-1];
reg [vec_width-1:0] vec;

wire u3352, u3351, u3350, u3349, u3348, u3347, u3346, u3345, u3344, u3343, u3342, u3341, u3340, u3339, u3338, u3337, u3336, u3335, u3334, u3333, u3332, u3331, u3330, u3329, u3328, u3327, u3326, u3325, u3324, u3323, u3322, u3321, u3458, u3459, u3320, u3319, u3318, u3317, u3316, u3315, u3314, u3313, u3312, u3311, u3310, u3309, u3308, u3307, u3306, u3305, u3304, u3303, u3302, u3301, u3300, u3299, u3298, u3297, u3296, u3295, u3294, u3293, u3292, u3291, u3467, u3469, u3471, u3473, u3475, u3477, u3479, u3481, u3483, u3485, u3487, u3489, u3491, u3493, u3495, u3497, u3499, u3501, u3503, u3505, u3506, u3507, u3508, u3509, u3510, u3511, u3512, u3513, u3514, u3515, u3516, u3517, u3518, u3519, u3520, u3521, u3522, u3523, u3524, u3525, u3526, u3527, u3528, u3529, u3530, u3531, u3532, u3533, u3534, u3535, u3536, u3537, u3538, u3539, u3540, u3541, u3542, u3543, u3544, u3545, u3546, u3547, u3548, u3549, u3290, u3289, u3288, u3287, u3286, u3285, u3284, u3283, u3282, u3281, u3280, u3279, u3278, u3277, u3276, u3275, u3274, u3273, u3272, u3271, u3270, u3269, u3268, u3267, u3266, u3265, u3264, u3263, u3262, u3354, u3261, u3260, u3259, u3258, u3257, u3256, u3255, u3254, u3253, u3252, u3251, u3250, u3249, u3248, u3247, u3246, u3245, u3244, u3243, u3242, u3241, u3240, u3550, u3551, u3552, u3553, u3554, u3555, u3556, u3557, u3558, u3559, u3560, u3561, u3562, u3563, u3564, u3565, u3566, u3567, u3568, u3569, u3570, u3571, u3572, u3573, u3574, u3575, u3576, u3577, u3578, u3579, u3580, u3581, u3239, u3238, u3237, u3236, u3235, u3234, u3233, u3232, u3231, u3230, u3229, u3228, u3227, u3226, u3225, u3224, u3223, u3222, u3221, u3220, u3219, u3218, u3217, u3216, u3215, u3214, u3213, u3212, u3211, u3210, u3149, u3148, u4043, addr_reg_19_, addr_reg_18_, addr_reg_17_, addr_reg_16_, addr_reg_15_, addr_reg_14_, addr_reg_13_, addr_reg_12_, addr_reg_11_, addr_reg_10_, addr_reg_9_, addr_reg_8_, addr_reg_7_, addr_reg_6_, addr_reg_5_, addr_reg_4_, addr_reg_3_, addr_reg_2_, addr_reg_1_, addr_reg_0_, datao_reg_31_, datao_reg_30_, datao_reg_29_, datao_reg_28_, datao_reg_27_, datao_reg_26_, datao_reg_25_, datao_reg_24_, datao_reg_23_, datao_reg_22_, datao_reg_21_, datao_reg_20_, datao_reg_19_, datao_reg_18_, datao_reg_17_, datao_reg_16_, datao_reg_15_, datao_reg_14_, datao_reg_13_, datao_reg_12_, datao_reg_11_, datao_reg_10_, datao_reg_9_, datao_reg_8_, datao_reg_7_, datao_reg_6_, datao_reg_5_, datao_reg_4_, datao_reg_3_, datao_reg_2_, datao_reg_1_, datao_reg_0_, rd_reg, wr_reg;
initial begin
	$readmemb(`in_file, input_vec_mem );
end

always #(`cycle/2) clk = ~clk;

b14_ras cc (.IR_REG_0_(vec[276]), .IR_REG_1_(vec[275]), .IR_REG_2_(vec[274]), .IR_REG_3_(vec[273]), .IR_REG_4_(vec[272]), .IR_REG_5_(vec[271]), .IR_REG_6_(vec[270]), .IR_REG_7_(vec[269]), .IR_REG_8_(vec[268]), .IR_REG_9_(vec[267]), .IR_REG_10_(vec[266]), .IR_REG_11_(vec[265]), .IR_REG_12_(vec[264]), .IR_REG_13_(vec[263]), .IR_REG_14_(vec[262]), .IR_REG_15_(vec[261]), .IR_REG_16_(vec[260]), .IR_REG_17_(vec[259]), .IR_REG_18_(vec[258]), .IR_REG_19_(vec[257]), .IR_REG_20_(vec[256]), .IR_REG_21_(vec[255]), .IR_REG_22_(vec[254]), .IR_REG_23_(vec[253]), .IR_REG_24_(vec[252]), .IR_REG_25_(vec[251]), .IR_REG_26_(vec[250]), .IR_REG_27_(vec[249]), .IR_REG_28_(vec[248]), .IR_REG_29_(vec[247]), .IR_REG_30_(vec[246]), .IR_REG_31_(vec[245]), .D_REG_0_(vec[244]), .D_REG_1_(vec[243]), .D_REG_2_(vec[242]), .D_REG_3_(vec[241]), .D_REG_4_(vec[240]), .D_REG_5_(vec[239]), .D_REG_6_(vec[238]), .D_REG_7_(vec[237]), .D_REG_8_(vec[236]), .D_REG_9_(vec[235]), .D_REG_10_(vec[234]), .D_REG_11_(vec[233]), .D_REG_12_(vec[232]), .D_REG_13_(vec[231]), .D_REG_14_(vec[230]), .D_REG_15_(vec[229]), .D_REG_16_(vec[228]), .D_REG_17_(vec[227]), .D_REG_18_(vec[226]), .D_REG_19_(vec[225]), .D_REG_20_(vec[224]), .D_REG_21_(vec[223]), .D_REG_22_(vec[222]), .D_REG_23_(vec[221]), .D_REG_24_(vec[220]), .D_REG_25_(vec[219]), .D_REG_26_(vec[218]), .D_REG_27_(vec[217]), .D_REG_28_(vec[216]), .D_REG_29_(vec[215]), .D_REG_30_(vec[214]), .D_REG_31_(vec[213]), .REG0_REG_0_(vec[212]), .REG0_REG_1_(vec[211]), .REG0_REG_2_(vec[210]), .REG0_REG_3_(vec[209]), .REG0_REG_4_(vec[208]), .REG0_REG_5_(vec[207]), .REG0_REG_6_(vec[206]), .REG0_REG_7_(vec[205]), .REG0_REG_8_(vec[204]), .REG0_REG_9_(vec[203]), .REG0_REG_10_(vec[202]), .REG0_REG_11_(vec[201]), .REG0_REG_12_(vec[200]), .REG0_REG_13_(vec[199]), .REG0_REG_14_(vec[198]), .REG0_REG_15_(vec[197]), .REG0_REG_16_(vec[196]), .REG0_REG_17_(vec[195]), .REG0_REG_18_(vec[194]), .REG0_REG_19_(vec[193]), .REG0_REG_20_(vec[192]), .REG0_REG_21_(vec[191]), .REG0_REG_22_(vec[190]), .REG0_REG_23_(vec[189]), .REG0_REG_24_(vec[188]), .REG0_REG_25_(vec[187]), .REG0_REG_26_(vec[186]), .REG0_REG_27_(vec[185]), .REG0_REG_28_(vec[184]), .REG0_REG_29_(vec[183]), .REG0_REG_30_(vec[182]), .REG0_REG_31_(vec[181]), .REG1_REG_0_(vec[180]), .REG1_REG_1_(vec[179]), .REG1_REG_2_(vec[178]), .REG1_REG_3_(vec[177]), .REG1_REG_4_(vec[176]), .REG1_REG_5_(vec[175]), .REG1_REG_6_(vec[174]), .REG1_REG_7_(vec[173]), .REG1_REG_8_(vec[172]), .REG1_REG_9_(vec[171]), .REG1_REG_10_(vec[170]), .REG1_REG_11_(vec[169]), .REG1_REG_12_(vec[168]), .REG1_REG_13_(vec[167]), .REG1_REG_14_(vec[166]), .REG1_REG_15_(vec[165]), .REG1_REG_16_(vec[164]), .REG1_REG_17_(vec[163]), .REG1_REG_18_(vec[162]), .REG1_REG_19_(vec[161]), .REG1_REG_20_(vec[160]), .REG1_REG_21_(vec[159]), .REG1_REG_22_(vec[158]), .REG1_REG_23_(vec[157]), .REG1_REG_24_(vec[156]), .REG1_REG_25_(vec[155]), .REG1_REG_26_(vec[154]), .REG1_REG_27_(vec[153]), .REG1_REG_28_(vec[152]), .REG1_REG_29_(vec[151]), .REG1_REG_30_(vec[150]), .REG1_REG_31_(vec[149]), .REG2_REG_0_(vec[148]), .REG2_REG_1_(vec[147]), .REG2_REG_2_(vec[146]), .REG2_REG_3_(vec[145]), .REG2_REG_4_(vec[144]), .REG2_REG_5_(vec[143]), .REG2_REG_6_(vec[142]), .REG2_REG_7_(vec[141]), .REG2_REG_8_(vec[140]), .REG2_REG_9_(vec[139]), .REG2_REG_10_(vec[138]), .REG2_REG_11_(vec[137]), .REG2_REG_12_(vec[136]), .REG2_REG_13_(vec[135]), .REG2_REG_14_(vec[134]), .REG2_REG_15_(vec[133]), .REG2_REG_16_(vec[132]), .REG2_REG_17_(vec[131]), .REG2_REG_18_(vec[130]), .REG2_REG_19_(vec[129]), .REG2_REG_20_(vec[128]), .REG2_REG_21_(vec[127]), .REG2_REG_22_(vec[126]), .REG2_REG_23_(vec[125]), .REG2_REG_24_(vec[124]), .REG2_REG_25_(vec[123]), .REG2_REG_26_(vec[122]), .REG2_REG_27_(vec[121]), .REG2_REG_28_(vec[120]), .REG2_REG_29_(vec[119]), .REG2_REG_30_(vec[118]), .REG2_REG_31_(vec[117]), .ADDR_REG_19__EXTRA(vec[116]), .ADDR_REG_18__EXTRA(vec[115]), .ADDR_REG_17__EXTRA(vec[114]), .ADDR_REG_16__EXTRA(vec[113]), .ADDR_REG_15__EXTRA(vec[112]), .ADDR_REG_14__EXTRA(vec[111]), .ADDR_REG_13__EXTRA(vec[110]), .ADDR_REG_12__EXTRA(vec[109]), .ADDR_REG_11__EXTRA(vec[108]), .ADDR_REG_10__EXTRA(vec[107]), .ADDR_REG_9__EXTRA(vec[106]), .ADDR_REG_8__EXTRA(vec[105]), .ADDR_REG_7__EXTRA(vec[104]), .ADDR_REG_6__EXTRA(vec[103]), .ADDR_REG_5__EXTRA(vec[102]), .ADDR_REG_4__EXTRA(vec[101]), .ADDR_REG_3__EXTRA(vec[100]), .ADDR_REG_2__EXTRA(vec[99]), .ADDR_REG_1__EXTRA(vec[98]), .ADDR_REG_0__EXTRA(vec[97]), .DATAO_REG_0__EXTRA(vec[96]), .DATAO_REG_1__EXTRA(vec[95]), .DATAO_REG_2__EXTRA(vec[94]), .DATAO_REG_3__EXTRA(vec[93]), .DATAO_REG_4__EXTRA(vec[92]), .DATAO_REG_5__EXTRA(vec[91]), .DATAO_REG_6__EXTRA(vec[90]), .DATAO_REG_7__EXTRA(vec[89]), .DATAO_REG_8__EXTRA(vec[88]), .DATAO_REG_9__EXTRA(vec[87]), .DATAO_REG_10__EXTRA(vec[86]), .DATAO_REG_11__EXTRA(vec[85]), .DATAO_REG_12__EXTRA(vec[84]), .DATAO_REG_13__EXTRA(vec[83]), .DATAO_REG_14__EXTRA(vec[82]), .DATAO_REG_15__EXTRA(vec[81]), .DATAO_REG_16__EXTRA(vec[80]), .DATAO_REG_17__EXTRA(vec[79]), .DATAO_REG_18__EXTRA(vec[78]), .DATAO_REG_19__EXTRA(vec[77]), .DATAO_REG_20__EXTRA(vec[76]), .DATAO_REG_21__EXTRA(vec[75]), .DATAO_REG_22__EXTRA(vec[74]), .DATAO_REG_23__EXTRA(vec[73]), .DATAO_REG_24__EXTRA(vec[72]), .DATAO_REG_25__EXTRA(vec[71]), .DATAO_REG_26__EXTRA(vec[70]), .DATAO_REG_27__EXTRA(vec[69]), .DATAO_REG_28__EXTRA(vec[68]), .DATAO_REG_29__EXTRA(vec[67]), .DATAO_REG_30__EXTRA(vec[66]), .DATAO_REG_31__EXTRA(vec[65]), .B_REG(vec[64]), .REG3_REG_15_(vec[63]), .REG3_REG_26_(vec[62]), .REG3_REG_6_(vec[61]), .REG3_REG_18_(vec[60]), .REG3_REG_2_(vec[59]), .REG3_REG_11_(vec[58]), .REG3_REG_22_(vec[57]), .REG3_REG_13_(vec[56]), .REG3_REG_20_(vec[55]), .REG3_REG_0_(vec[54]), .REG3_REG_9_(vec[53]), .REG3_REG_4_(vec[52]), .REG3_REG_24_(vec[51]), .REG3_REG_17_(vec[50]), .REG3_REG_5_(vec[49]), .REG3_REG_16_(vec[48]), .REG3_REG_25_(vec[47]), .REG3_REG_12_(vec[46]), .REG3_REG_21_(vec[45]), .REG3_REG_1_(vec[44]), .REG3_REG_8_(vec[43]), .REG3_REG_28_(vec[42]), .REG3_REG_19_(vec[41]), .REG3_REG_3_(vec[40]), .REG3_REG_10_(vec[39]), .REG3_REG_23_(vec[38]), .REG3_REG_14_(vec[37]), .REG3_REG_27_(vec[36]), .REG3_REG_7_(vec[35]), .STATE_REG(vec[34]), .RD_REG_EXTRA(vec[33]), .WR_REG_EXTRA(vec[32]), .DATAI_31_(vec[31]), .DATAI_30_(vec[30]), .DATAI_29_(vec[29]), .DATAI_28_(vec[28]), .DATAI_27_(vec[27]), .DATAI_26_(vec[26]), .DATAI_25_(vec[25]), .DATAI_24_(vec[24]), .DATAI_23_(vec[23]), .DATAI_22_(vec[22]), .DATAI_21_(vec[21]), .DATAI_20_(vec[20]), .DATAI_19_(vec[19]), .DATAI_18_(vec[18]), .DATAI_17_(vec[17]), .DATAI_16_(vec[16]), .DATAI_15_(vec[15]), .DATAI_14_(vec[14]), .DATAI_13_(vec[13]), .DATAI_12_(vec[12]), .DATAI_11_(vec[11]), .DATAI_10_(vec[10]), .DATAI_9_(vec[9]), .DATAI_8_(vec[8]), .DATAI_7_(vec[7]), .DATAI_6_(vec[6]), .DATAI_5_(vec[5]), .DATAI_4_(vec[4]), .DATAI_3_(vec[3]), .DATAI_2_(vec[2]), .DATAI_1_(vec[1]), .DATAI_0_(vec[0]), .U3352(u3352), .U3351(u3351), .U3350(u3350), .U3349(u3349), .U3348(u3348), .U3347(u3347), .U3346(u3346), .U3345(u3345), .U3344(u3344), .U3343(u3343), .U3342(u3342), .U3341(u3341), .U3340(u3340), .U3339(u3339), .U3338(u3338), .U3337(u3337), .U3336(u3336), .U3335(u3335), .U3334(u3334), .U3333(u3333), .U3332(u3332), .U3331(u3331), .U3330(u3330), .U3329(u3329), .U3328(u3328), .U3327(u3327), .U3326(u3326), .U3325(u3325), .U3324(u3324), .U3323(u3323), .U3322(u3322), .U3321(u3321), .U3458(u3458), .U3459(u3459), .U3320(u3320), .U3319(u3319), .U3318(u3318), .U3317(u3317), .U3316(u3316), .U3315(u3315), .U3314(u3314), .U3313(u3313), .U3312(u3312), .U3311(u3311), .U3310(u3310), .U3309(u3309), .U3308(u3308), .U3307(u3307), .U3306(u3306), .U3305(u3305), .U3304(u3304), .U3303(u3303), .U3302(u3302), .U3301(u3301), .U3300(u3300), .U3299(u3299), .U3298(u3298), .U3297(u3297), .U3296(u3296), .U3295(u3295), .U3294(u3294), .U3293(u3293), .U3292(u3292), .U3291(u3291), .U3467(u3467), .U3469(u3469), .U3471(u3471), .U3473(u3473), .U3475(u3475), .U3477(u3477), .U3479(u3479), .U3481(u3481), .U3483(u3483), .U3485(u3485), .U3487(u3487), .U3489(u3489), .U3491(u3491), .U3493(u3493), .U3495(u3495), .U3497(u3497), .U3499(u3499), .U3501(u3501), .U3503(u3503), .U3505(u3505), .U3506(u3506), .U3507(u3507), .U3508(u3508), .U3509(u3509), .U3510(u3510), .U3511(u3511), .U3512(u3512), .U3513(u3513), .U3514(u3514), .U3515(u3515), .U3516(u3516), .U3517(u3517), .U3518(u3518), .U3519(u3519), .U3520(u3520), .U3521(u3521), .U3522(u3522), .U3523(u3523), .U3524(u3524), .U3525(u3525), .U3526(u3526), .U3527(u3527), .U3528(u3528), .U3529(u3529), .U3530(u3530), .U3531(u3531), .U3532(u3532), .U3533(u3533), .U3534(u3534), .U3535(u3535), .U3536(u3536), .U3537(u3537), .U3538(u3538), .U3539(u3539), .U3540(u3540), .U3541(u3541), .U3542(u3542), .U3543(u3543), .U3544(u3544), .U3545(u3545), .U3546(u3546), .U3547(u3547), .U3548(u3548), .U3549(u3549), .U3290(u3290), .U3289(u3289), .U3288(u3288), .U3287(u3287), .U3286(u3286), .U3285(u3285), .U3284(u3284), .U3283(u3283), .U3282(u3282), .U3281(u3281), .U3280(u3280), .U3279(u3279), .U3278(u3278), .U3277(u3277), .U3276(u3276), .U3275(u3275), .U3274(u3274), .U3273(u3273), .U3272(u3272), .U3271(u3271), .U3270(u3270), .U3269(u3269), .U3268(u3268), .U3267(u3267), .U3266(u3266), .U3265(u3265), .U3264(u3264), .U3263(u3263), .U3262(u3262), .U3354(u3354), .U3261(u3261), .U3260(u3260), .U3259(u3259), .U3258(u3258), .U3257(u3257), .U3256(u3256), .U3255(u3255), .U3254(u3254), .U3253(u3253), .U3252(u3252), .U3251(u3251), .U3250(u3250), .U3249(u3249), .U3248(u3248), .U3247(u3247), .U3246(u3246), .U3245(u3245), .U3244(u3244), .U3243(u3243), .U3242(u3242), .U3241(u3241), .U3240(u3240), .U3550(u3550), .U3551(u3551), .U3552(u3552), .U3553(u3553), .U3554(u3554), .U3555(u3555), .U3556(u3556), .U3557(u3557), .U3558(u3558), .U3559(u3559), .U3560(u3560), .U3561(u3561), .U3562(u3562), .U3563(u3563), .U3564(u3564), .U3565(u3565), .U3566(u3566), .U3567(u3567), .U3568(u3568), .U3569(u3569), .U3570(u3570), .U3571(u3571), .U3572(u3572), .U3573(u3573), .U3574(u3574), .U3575(u3575), .U3576(u3576), .U3577(u3577), .U3578(u3578), .U3579(u3579), .U3580(u3580), .U3581(u3581), .U3239(u3239), .U3238(u3238), .U3237(u3237), .U3236(u3236), .U3235(u3235), .U3234(u3234), .U3233(u3233), .U3232(u3232), .U3231(u3231), .U3230(u3230), .U3229(u3229), .U3228(u3228), .U3227(u3227), .U3226(u3226), .U3225(u3225), .U3224(u3224), .U3223(u3223), .U3222(u3222), .U3221(u3221), .U3220(u3220), .U3219(u3219), .U3218(u3218), .U3217(u3217), .U3216(u3216), .U3215(u3215), .U3214(u3214), .U3213(u3213), .U3212(u3212), .U3211(u3211), .U3210(u3210), .U3149(u3149), .U3148(u3148), .U4043(u4043), .ADDR_REG_19_(addr_reg_19_), .ADDR_REG_18_(addr_reg_18_), .ADDR_REG_17_(addr_reg_17_), .ADDR_REG_16_(addr_reg_16_), .ADDR_REG_15_(addr_reg_15_), .ADDR_REG_14_(addr_reg_14_), .ADDR_REG_13_(addr_reg_13_), .ADDR_REG_12_(addr_reg_12_), .ADDR_REG_11_(addr_reg_11_), .ADDR_REG_10_(addr_reg_10_), .ADDR_REG_9_(addr_reg_9_), .ADDR_REG_8_(addr_reg_8_), .ADDR_REG_7_(addr_reg_7_), .ADDR_REG_6_(addr_reg_6_), .ADDR_REG_5_(addr_reg_5_), .ADDR_REG_4_(addr_reg_4_), .ADDR_REG_3_(addr_reg_3_), .ADDR_REG_2_(addr_reg_2_), .ADDR_REG_1_(addr_reg_1_), .ADDR_REG_0_(addr_reg_0_), .DATAO_REG_31_(datao_reg_31_), .DATAO_REG_30_(datao_reg_30_), .DATAO_REG_29_(datao_reg_29_), .DATAO_REG_28_(datao_reg_28_), .DATAO_REG_27_(datao_reg_27_), .DATAO_REG_26_(datao_reg_26_), .DATAO_REG_25_(datao_reg_25_), .DATAO_REG_24_(datao_reg_24_), .DATAO_REG_23_(datao_reg_23_), .DATAO_REG_22_(datao_reg_22_), .DATAO_REG_21_(datao_reg_21_), .DATAO_REG_20_(datao_reg_20_), .DATAO_REG_19_(datao_reg_19_), .DATAO_REG_18_(datao_reg_18_), .DATAO_REG_17_(datao_reg_17_), .DATAO_REG_16_(datao_reg_16_), .DATAO_REG_15_(datao_reg_15_), .DATAO_REG_14_(datao_reg_14_), .DATAO_REG_13_(datao_reg_13_), .DATAO_REG_12_(datao_reg_12_), .DATAO_REG_11_(datao_reg_11_), .DATAO_REG_10_(datao_reg_10_), .DATAO_REG_9_(datao_reg_9_), .DATAO_REG_8_(datao_reg_8_), .DATAO_REG_7_(datao_reg_7_), .DATAO_REG_6_(datao_reg_6_), .DATAO_REG_5_(datao_reg_5_), .DATAO_REG_4_(datao_reg_4_), .DATAO_REG_3_(datao_reg_3_), .DATAO_REG_2_(datao_reg_2_), .DATAO_REG_1_(datao_reg_1_), .DATAO_REG_0_(datao_reg_0_), .RD_REG(rd_reg), .WR_REG(wr_reg));

integer i=0;
always @ (posedge clk) begin
	vec = input_vec_mem[i];
	$monitor(vec);
	i = i + 1;

end

always @ (negedge clk)begin
	$fdisplay ( fh_w, u3352, u3351, u3350, u3349, u3348, u3347, u3346, u3345, u3344, u3343, u3342, u3341, u3340, u3339, u3338, u3337, u3336, u3335, u3334, u3333, u3332, u3331, u3330, u3329, u3328, u3327, u3326, u3325, u3324, u3323, u3322, u3321, u3458, u3459, u3320, u3319, u3318, u3317, u3316, u3315, u3314, u3313, u3312, u3311, u3310, u3309, u3308, u3307, u3306, u3305, u3304, u3303, u3302, u3301, u3300, u3299, u3298, u3297, u3296, u3295, u3294, u3293, u3292, u3291, u3467, u3469, u3471, u3473, u3475, u3477, u3479, u3481, u3483, u3485, u3487, u3489, u3491, u3493, u3495, u3497, u3499, u3501, u3503, u3505, u3506, u3507, u3508, u3509, u3510, u3511, u3512, u3513, u3514, u3515, u3516, u3517, u3518, u3519, u3520, u3521, u3522, u3523, u3524, u3525, u3526, u3527, u3528, u3529, u3530, u3531, u3532, u3533, u3534, u3535, u3536, u3537, u3538, u3539, u3540, u3541, u3542, u3543, u3544, u3545, u3546, u3547, u3548, u3549, u3290, u3289, u3288, u3287, u3286, u3285, u3284, u3283, u3282, u3281, u3280, u3279, u3278, u3277, u3276, u3275, u3274, u3273, u3272, u3271, u3270, u3269, u3268, u3267, u3266, u3265, u3264, u3263, u3262, u3354, u3261, u3260, u3259, u3258, u3257, u3256, u3255, u3254, u3253, u3252, u3251, u3250, u3249, u3248, u3247, u3246, u3245, u3244, u3243, u3242, u3241, u3240, u3550, u3551, u3552, u3553, u3554, u3555, u3556, u3557, u3558, u3559, u3560, u3561, u3562, u3563, u3564, u3565, u3566, u3567, u3568, u3569, u3570, u3571, u3572, u3573, u3574, u3575, u3576, u3577, u3578, u3579, u3580, u3581, u3239, u3238, u3237, u3236, u3235, u3234, u3233, u3232, u3231, u3230, u3229, u3228, u3227, u3226, u3225, u3224, u3223, u3222, u3221, u3220, u3219, u3218, u3217, u3216, u3215, u3214, u3213, u3212, u3211, u3210, u3149, u3148, u4043, addr_reg_19_, addr_reg_18_, addr_reg_17_, addr_reg_16_, addr_reg_15_, addr_reg_14_, addr_reg_13_, addr_reg_12_, addr_reg_11_, addr_reg_10_, addr_reg_9_, addr_reg_8_, addr_reg_7_, addr_reg_6_, addr_reg_5_, addr_reg_4_, addr_reg_3_, addr_reg_2_, addr_reg_1_, addr_reg_0_, datao_reg_31_, datao_reg_30_, datao_reg_29_, datao_reg_28_, datao_reg_27_, datao_reg_26_, datao_reg_25_, datao_reg_24_, datao_reg_23_, datao_reg_22_, datao_reg_21_, datao_reg_20_, datao_reg_19_, datao_reg_18_, datao_reg_17_, datao_reg_16_, datao_reg_15_, datao_reg_14_, datao_reg_13_, datao_reg_12_, datao_reg_11_, datao_reg_10_, datao_reg_9_, datao_reg_8_, datao_reg_7_, datao_reg_6_, datao_reg_5_, datao_reg_4_, datao_reg_3_, datao_reg_2_, datao_reg_1_, datao_reg_0_, rd_reg, wr_reg);
	if(i == vec_length)begin
		$finish;
	end
end

integer fh_w;
initial begin
	fh_w = $fopen(`out_file, "w");
end
 
initial begin
	//$fsdbDumpfile("SET.fsdb");
	//$fsdbDumpvars;
	//$fsdbDumpMDA;
	$dumpfile("test_result.vcd");
    $dumpvars;

end
endmodule
