`timescale 1ns/10ps

`define cycle 10.0
`define terminate_cycle 400000//200000 // Modify your terminate ycle here

module b17_ras_testfixture;

`define in_file "b17_ras/rand_input_vector_b17_ras_0.out"
`define out_file "b17_ras/rand_output_vector_b17_ras_0.out"

parameter vec_width = 1452;
parameter vec_length = 7;

reg clk = 0;


reg [vec_width-1:0] input_vec_mem [0:vec_length-1];
reg [vec_width-1:0] vec;

wire p3_datao_reg_31_, p3_datao_reg_30_, p3_datao_reg_29_, p3_datao_reg_28_, p3_datao_reg_27_, p3_datao_reg_26_, p3_datao_reg_25_, p3_datao_reg_24_, p3_datao_reg_23_, p3_datao_reg_22_, p3_datao_reg_21_, p3_datao_reg_20_, p3_datao_reg_19_, p3_datao_reg_18_, p3_datao_reg_17_, p3_datao_reg_16_, p3_datao_reg_15_, p3_datao_reg_14_, p3_datao_reg_13_, p3_datao_reg_12_, p3_datao_reg_11_, p3_datao_reg_10_, p3_datao_reg_9_, p3_datao_reg_8_, p3_datao_reg_7_, p3_datao_reg_6_, p3_datao_reg_5_, p3_datao_reg_4_, p3_datao_reg_3_, p3_datao_reg_2_, p3_datao_reg_1_, p3_datao_reg_0_, p1_address_reg_29_, p1_address_reg_28_, p1_address_reg_27_, p1_address_reg_26_, p1_address_reg_25_, p1_address_reg_24_, p1_address_reg_23_, p1_address_reg_22_, p1_address_reg_21_, p1_address_reg_20_, p1_address_reg_19_, p1_address_reg_18_, p1_address_reg_17_, p1_address_reg_16_, p1_address_reg_15_, p1_address_reg_14_, p1_address_reg_13_, p1_address_reg_12_, p1_address_reg_11_, p1_address_reg_10_, p1_address_reg_9_, p1_address_reg_8_, p1_address_reg_7_, p1_address_reg_6_, p1_address_reg_5_, p1_address_reg_4_, p1_address_reg_3_, p1_address_reg_2_, p1_address_reg_1_, p1_address_reg_0_, u355, u356, u357, u358, u359, u360, u361, u362, u363, u364, u366, u367, u368, u369, u370, u371, u372, u373, u374, u375, u347, u348, u349, u350, u351, u352, u353, u354, u365, u376, p3_w_r_n_reg, p3_d_c_n_reg, p3_m_io_n_reg, p1_ads_n_reg, p3_ads_n_reg, u247, u246, u245, u244, u243, u242, u241, u240, u239, u238, u237, u236, u235, u234, u233, u232, u231, u230, u229, u228, u227, u226, u225, u224, u223, u222, u221, u220, u219, u218, u217, u216, u251, u252, u253, u254, u255, u256, u257, u258, u259, u260, u261, u262, u263, u264, u265, u266, u267, u268, u269, u270, u271, u272, u273, u274, u275, u276, u277, u278, u279, u280, u281, u282, u212, u215, u213, u214, p3_u3274, p3_u3275, p3_u3276, p3_u3277, p3_u3061, p3_u3060, p3_u3059, p3_u3058, p3_u3057, p3_u3056, p3_u3055, p3_u3054, p3_u3053, p3_u3052, p3_u3051, p3_u3050, p3_u3049, p3_u3048, p3_u3047, p3_u3046, p3_u3045, p3_u3044, p3_u3043, p3_u3042, p3_u3041, p3_u3040, p3_u3039, p3_u3038, p3_u3037, p3_u3036, p3_u3035, p3_u3034, p3_u3033, p3_u3032, p3_u3031, p3_u3030, p3_u3029, p3_u3280, p3_u3281, p3_u3028, p3_u3027, p3_u3026, p3_u3025, p3_u3024, p3_u3023, p3_u3022, p3_u3021, p3_u3020, p3_u3019, p3_u3018, p3_u3017, p3_u3016, p3_u3015, p3_u3014, p3_u3013, p3_u3012, p3_u3011, p3_u3010, p3_u3009, p3_u3008, p3_u3007, p3_u3006, p3_u3005, p3_u3004, p3_u3003, p3_u3002, p3_u3001, p3_u3000, p3_u2999, p3_u3282, p3_u2998, p3_u2997, p3_u2996, p3_u2995, p3_u2994, p3_u2993, p3_u2992, p3_u2991, p3_u2990, p3_u2989, p3_u2988, p3_u2987, p3_u2986, p3_u2985, p3_u2984, p3_u2983, p3_u2982, p3_u2981, p3_u2980, p3_u2979, p3_u2978, p3_u2977, p3_u2976, p3_u2975, p3_u2974, p3_u2973, p3_u2972, p3_u2971, p3_u2970, p3_u2969, p3_u2968, p3_u2967, p3_u2966, p3_u2965, p3_u2964, p3_u2963, p3_u2962, p3_u2961, p3_u2960, p3_u2959, p3_u2958, p3_u2957, p3_u2956, p3_u2955, p3_u2954, p3_u2953, p3_u2952, p3_u2951, p3_u2950, p3_u2949, p3_u2948, p3_u2947, p3_u2946, p3_u2945, p3_u2944, p3_u2943, p3_u2942, p3_u2941, p3_u2940, p3_u2939, p3_u2938, p3_u2937, p3_u2936, p3_u2935, p3_u2934, p3_u2933, p3_u2932, p3_u2931, p3_u2930, p3_u2929, p3_u2928, p3_u2927, p3_u2926, p3_u2925, p3_u2924, p3_u2923, p3_u2922, p3_u2921, p3_u2920, p3_u2919, p3_u2918, p3_u2917, p3_u2916, p3_u2915, p3_u2914, p3_u2913, p3_u2912, p3_u2911, p3_u2910, p3_u2909, p3_u2908, p3_u2907, p3_u2906, p3_u2905, p3_u2904, p3_u2903, p3_u2902, p3_u2901, p3_u2900, p3_u2899, p3_u2898, p3_u2897, p3_u2896, p3_u2895, p3_u2894, p3_u2893, p3_u2892, p3_u2891, p3_u2890, p3_u2889, p3_u2888, p3_u2887, p3_u2886, p3_u2885, p3_u2884, p3_u2883, p3_u2882, p3_u2881, p3_u2880, p3_u2879, p3_u2878, p3_u2877, p3_u2876, p3_u2875, p3_u2874, p3_u2873, p3_u2872, p3_u2871, p3_u2870, p3_u2869, p3_u2868, p3_u3284, p3_u3285, p3_u3288, p3_u3289, p3_u3290, p3_u2867, p3_u2866, p3_u2865, p3_u2864, p3_u2863, p3_u2862, p3_u2861, p3_u2860, p3_u2859, p3_u2858, p3_u2857, p3_u2856, p3_u2855, p3_u2854, p3_u2853, p3_u2852, p3_u2851, p3_u2850, p3_u2849, p3_u2848, p3_u2847, p3_u2846, p3_u2845, p3_u2844, p3_u2843, p3_u2842, p3_u2841, p3_u2840, p3_u2839, p3_u2838, p3_u2837, p3_u2836, p3_u2835, p3_u2834, p3_u2833, p3_u2832, p3_u2831, p3_u2830, p3_u2829, p3_u2828, p3_u2827, p3_u2826, p3_u2825, p3_u2824, p3_u2823, p3_u2822, p3_u2821, p3_u2820, p3_u2819, p3_u2818, p3_u2817, p3_u2816, p3_u2815, p3_u2814, p3_u2813, p3_u2812, p3_u2811, p3_u2810, p3_u2809, p3_u2808, p3_u2807, p3_u2806, p3_u2805, p3_u2804, p3_u2803, p3_u2802, p3_u2801, p3_u2800, p3_u2799, p3_u2798, p3_u2797, p3_u2796, p3_u2795, p3_u2794, p3_u2793, p3_u2792, p3_u2791, p3_u2790, p3_u2789, p3_u2788, p3_u2787, p3_u2786, p3_u2785, p3_u2784, p3_u2783, p3_u2782, p3_u2781, p3_u2780, p3_u2779, p3_u2778, p3_u2777, p3_u2776, p3_u2775, p3_u2774, p3_u2773, p3_u2772, p3_u2771, p3_u2770, p3_u2769, p3_u2768, p3_u2767, p3_u2766, p3_u2765, p3_u2764, p3_u2763, p3_u2762, p3_u2761, p3_u2760, p3_u2759, p3_u2758, p3_u2757, p3_u2756, p3_u2755, p3_u2754, p3_u2753, p3_u2752, p3_u2751, p3_u2750, p3_u2749, p3_u2748, p3_u2747, p3_u2746, p3_u2745, p3_u2744, p3_u2743, p3_u2742, p3_u2741, p3_u2740, p3_u2739, p3_u2738, p3_u2737, p3_u2736, p3_u2735, p3_u2734, p3_u2733, p3_u2732, p3_u2731, p3_u2730, p3_u2729, p3_u2728, p3_u2727, p3_u2726, p3_u2725, p3_u2724, p3_u2723, p3_u2722, p3_u2721, p3_u2720, p3_u2719, p3_u2718, p3_u2717, p3_u2716, p3_u2715, p3_u2714, p3_u2713, p3_u2712, p3_u2711, p3_u2710, p3_u2709, p3_u2708, p3_u2707, p3_u2706, p3_u2705, p3_u2704, p3_u2703, p3_u2702, p3_u2701, p3_u2700, p3_u2699, p3_u2698, p3_u2697, p3_u2696, p3_u2695, p3_u2694, p3_u2693, p3_u2692, p3_u2691, p3_u2690, p3_u2689, p3_u2688, p3_u2687, p3_u2686, p3_u2685, p3_u2684, p3_u2683, p3_u2682, p3_u2681, p3_u2680, p3_u2679, p3_u2678, p3_u2677, p3_u2676, p3_u2675, p3_u2674, p3_u2673, p3_u2672, p3_u2671, p3_u2670, p3_u2669, p3_u2668, p3_u2667, p3_u2666, p3_u2665, p3_u2664, p3_u2663, p3_u2662, p3_u2661, p3_u2660, p3_u2659, p3_u2658, p3_u2657, p3_u2656, p3_u2655, p3_u2654, p3_u2653, p3_u2652, p3_u2651, p3_u2650, p3_u2649, p3_u2648, p3_u2647, p3_u2646, p3_u2645, p3_u2644, p3_u2643, p3_u2642, p3_u2641, p3_u2640, p3_u2639, p3_u3292, p3_u2638, p3_u3293, p3_u3294, p3_u2637, p3_u3295, p3_u2636, p3_u3296, p3_u2635, p3_u3297, p3_u2634, p3_u2633, p3_u3298, p3_u3299, p2_u3585, p2_u3586, p2_u3587, p2_u3588, p2_u3241, p2_u3240, p2_u3239, p2_u3238, p2_u3237, p2_u3236, p2_u3235, p2_u3234, p2_u3233, p2_u3232, p2_u3231, p2_u3230, p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225, p2_u3224, p2_u3223, p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218, p2_u3217, p2_u3216, p2_u3215, p2_u3214, p2_u3213, p2_u3212, p2_u3211, p2_u3210, p2_u3209, p2_u3591, p2_u3592, p2_u3208, p2_u3207, p2_u3206, p2_u3205, p2_u3204, p2_u3203, p2_u3202, p2_u3201, p2_u3200, p2_u3199, p2_u3198, p2_u3197, p2_u3196, p2_u3195, p2_u3194, p2_u3193, p2_u3192, p2_u3191, p2_u3190, p2_u3189, p2_u3188, p2_u3187, p2_u3186, p2_u3185, p2_u3184, p2_u3183, p2_u3182, p2_u3181, p2_u3180, p2_u3179, p2_u3593, p2_u3178, p2_u3177, p2_u3176, p2_u3175, p2_u3174, p2_u3173, p2_u3172, p2_u3171, p2_u3170, p2_u3169, p2_u3168, p2_u3167, p2_u3166, p2_u3165, p2_u3164, p2_u3163, p2_u3162, p2_u3161, p2_u3160, p2_u3159, p2_u3158, p2_u3157, p2_u3156, p2_u3155, p2_u3154, p2_u3153, p2_u3152, p2_u3151, p2_u3150, p2_u3149, p2_u3148, p2_u3147, p2_u3146, p2_u3145, p2_u3144, p2_u3143, p2_u3142, p2_u3141, p2_u3140, p2_u3139, p2_u3138, p2_u3137, p2_u3136, p2_u3135, p2_u3134, p2_u3133, p2_u3132, p2_u3131, p2_u3130, p2_u3129, p2_u3128, p2_u3127, p2_u3126, p2_u3125, p2_u3124, p2_u3123, p2_u3122, p2_u3121, p2_u3120, p2_u3119, p2_u3118, p2_u3117, p2_u3116, p2_u3115, p2_u3114, p2_u3113, p2_u3112, p2_u3111, p2_u3110, p2_u3109, p2_u3108, p2_u3107, p2_u3106, p2_u3105, p2_u3104, p2_u3103, p2_u3102, p2_u3101, p2_u3100, p2_u3099, p2_u3098, p2_u3097, p2_u3096, p2_u3095, p2_u3094, p2_u3093, p2_u3092, p2_u3091, p2_u3090, p2_u3089, p2_u3088, p2_u3087, p2_u3086, p2_u3085, p2_u3084, p2_u3083, p2_u3082, p2_u3081, p2_u3080, p2_u3079, p2_u3078, p2_u3077, p2_u3076, p2_u3075, p2_u3074, p2_u3073, p2_u3072, p2_u3071, p2_u3070, p2_u3069, p2_u3068, p2_u3067, p2_u3066, p2_u3065, p2_u3064, p2_u3063, p2_u3062, p2_u3061, p2_u3060, p2_u3059, p2_u3058, p2_u3057, p2_u3056, p2_u3055, p2_u3054, p2_u3053, p2_u3052, p2_u3051, p2_u3050, p2_u3049, p2_u3048, p2_u3595, p2_u3596, p2_u3599, p2_u3600, p2_u3601, p2_u3047, p2_u3602, p2_u3603, p2_u3604, p2_u3605, p2_u3046, p2_u3045, p2_u3044, p2_u3043, p2_u3042, p2_u3041, p2_u3040, p2_u3039, p2_u3038, p2_u3037, p2_u3036, p2_u3035, p2_u3034, p2_u3033, p2_u3032, p2_u3031, p2_u3030, p2_u3029, p2_u3028, p2_u3027, p2_u3026, p2_u3025, p2_u3024, p2_u3023, p2_u3022, p2_u3021, p2_u3020, p2_u3019, p2_u3018, p2_u3017, p2_u3016, p2_u3015, p2_u3014, p2_u3013, p2_u3012, p2_u3011, p2_u3010, p2_u3009, p2_u3008, p2_u3007, p2_u3006, p2_u3005, p2_u3004, p2_u3003, p2_u3002, p2_u3001, p2_u3000, p2_u2999, p2_u2998, p2_u2997, p2_u2996, p2_u2995, p2_u2994, p2_u2993, p2_u2992, p2_u2991, p2_u2990, p2_u2989, p2_u2988, p2_u2987, p2_u2986, p2_u2985, p2_u2984, p2_u2983, p2_u2982, p2_u2981, p2_u2980, p2_u2979, p2_u2978, p2_u2977, p2_u2976, p2_u2975, p2_u2974, p2_u2973, p2_u2972, p2_u2971, p2_u2970, p2_u2969, p2_u2968, p2_u2967, p2_u2966, p2_u2965, p2_u2964, p2_u2963, p2_u2962, p2_u2961, p2_u2960, p2_u2959, p2_u2958, p2_u2957, p2_u2956, p2_u2955, p2_u2954, p2_u2953, p2_u2952, p2_u2951, p2_u2950, p2_u2949, p2_u2948, p2_u2947, p2_u2946, p2_u2945, p2_u2944, p2_u2943, p2_u2942, p2_u2941, p2_u2940, p2_u2939, p2_u2938, p2_u2937, p2_u2936, p2_u2935, p2_u2934, p2_u2933, p2_u2932, p2_u2931, p2_u2930, p2_u2929, p2_u2928, p2_u2927, p2_u2926, p2_u2925, p2_u2924, p2_u2923, p2_u2922, p2_u2921, p2_u2920, p2_u2919, p2_u2918, p2_u2917, p2_u2916, p2_u2915, p2_u2914, p2_u2913, p2_u2912, p2_u2911, p2_u2910, p2_u2909, p2_u2908, p2_u2907, p2_u2906, p2_u2905, p2_u2904, p2_u2903, p2_u2902, p2_u2901, p2_u2900, p2_u2899, p2_u2898, p2_u2897, p2_u2896, p2_u2895, p2_u2894, p2_u2893, p2_u2892, p2_u2891, p2_u2890, p2_u2889, p2_u2888, p2_u2887, p2_u2886, p2_u2885, p2_u2884, p2_u2883, p2_u2882, p2_u2881, p2_u2880, p2_u2879, p2_u2878, p2_u2877, p2_u2876, p2_u2875, p2_u2874, p2_u2873, p2_u2872, p2_u2871, p2_u2870, p2_u2869, p2_u2868, p2_u2867, p2_u2866, p2_u2865, p2_u2864, p2_u2863, p2_u2862, p2_u2861, p2_u2860, p2_u2859, p2_u2858, p2_u2857, p2_u2856, p2_u2855, p2_u2854, p2_u2853, p2_u2852, p2_u2851, p2_u2850, p2_u2849, p2_u2848, p2_u2847, p2_u2846, p2_u2845, p2_u2844, p2_u2843, p2_u2842, p2_u2841, p2_u2840, p2_u2839, p2_u2838, p2_u2837, p2_u2836, p2_u2835, p2_u2834, p2_u2833, p2_u2832, p2_u2831, p2_u2830, p2_u2829, p2_u2828, p2_u2827, p2_u2826, p2_u2825, p2_u2824, p2_u2823, p2_u2822, p2_u2821, p2_u2820, p2_u3608, p2_u2819, p2_u3609, p2_u2818, p2_u3610, p2_u2817, p2_u3611, p2_u2816, p2_u2815, p2_u3612, p2_u2814, p1_u3458, p1_u3459, p1_u3460, p1_u3461, p1_u3226, p1_u3225, p1_u3224, p1_u3223, p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218, p1_u3217, p1_u3216, p1_u3215, p1_u3214, p1_u3213, p1_u3212, p1_u3211, p1_u3210, p1_u3209, p1_u3208, p1_u3207, p1_u3206, p1_u3205, p1_u3204, p1_u3203, p1_u3202, p1_u3201, p1_u3200, p1_u3199, p1_u3198, p1_u3197, p1_u3196, p1_u3195, p1_u3194, p1_u3464, p1_u3465, p1_u3193, p1_u3192, p1_u3191, p1_u3190, p1_u3189, p1_u3188, p1_u3187, p1_u3186, p1_u3185, p1_u3184, p1_u3183, p1_u3182, p1_u3181, p1_u3180, p1_u3179, p1_u3178, p1_u3177, p1_u3176, p1_u3175, p1_u3174, p1_u3173, p1_u3172, p1_u3171, p1_u3170, p1_u3169, p1_u3168, p1_u3167, p1_u3166, p1_u3165, p1_u3164, p1_u3466, p1_u3163, p1_u3162, p1_u3161, p1_u3160, p1_u3159, p1_u3158, p1_u3157, p1_u3156, p1_u3155, p1_u3154, p1_u3153, p1_u3152, p1_u3151, p1_u3150, p1_u3149, p1_u3148, p1_u3147, p1_u3146, p1_u3145, p1_u3144, p1_u3143, p1_u3142, p1_u3141, p1_u3140, p1_u3139, p1_u3138, p1_u3137, p1_u3136, p1_u3135, p1_u3134, p1_u3133, p1_u3132, p1_u3131, p1_u3130, p1_u3129, p1_u3128, p1_u3127, p1_u3126, p1_u3125, p1_u3124, p1_u3123, p1_u3122, p1_u3121, p1_u3120, p1_u3119, p1_u3118, p1_u3117, p1_u3116, p1_u3115, p1_u3114, p1_u3113, p1_u3112, p1_u3111, p1_u3110, p1_u3109, p1_u3108, p1_u3107, p1_u3106, p1_u3105, p1_u3104, p1_u3103, p1_u3102, p1_u3101, p1_u3100, p1_u3099, p1_u3098, p1_u3097, p1_u3096, p1_u3095, p1_u3094, p1_u3093, p1_u3092, p1_u3091, p1_u3090, p1_u3089, p1_u3088, p1_u3087, p1_u3086, p1_u3085, p1_u3084, p1_u3083, p1_u3082, p1_u3081, p1_u3080, p1_u3079, p1_u3078, p1_u3077, p1_u3076, p1_u3075, p1_u3074, p1_u3073, p1_u3072, p1_u3071, p1_u3070, p1_u3069, p1_u3068, p1_u3067, p1_u3066, p1_u3065, p1_u3064, p1_u3063, p1_u3062, p1_u3061, p1_u3060, p1_u3059, p1_u3058, p1_u3057, p1_u3056, p1_u3055, p1_u3054, p1_u3053, p1_u3052, p1_u3051, p1_u3050, p1_u3049, p1_u3048, p1_u3047, p1_u3046, p1_u3045, p1_u3044, p1_u3043, p1_u3042, p1_u3041, p1_u3040, p1_u3039, p1_u3038, p1_u3037, p1_u3036, p1_u3035, p1_u3034, p1_u3033, p1_u3468, p1_u3469, p1_u3472, p1_u3473, p1_u3474, p1_u3032, p1_u3475, p1_u3476, p1_u3477, p1_u3478, p1_u3031, p1_u3030, p1_u3029, p1_u3028, p1_u3027, p1_u3026, p1_u3025, p1_u3024, p1_u3023, p1_u3022, p1_u3021, p1_u3020, p1_u3019, p1_u3018, p1_u3017, p1_u3016, p1_u3015, p1_u3014, p1_u3013, p1_u3012, p1_u3011, p1_u3010, p1_u3009, p1_u3008, p1_u3007, p1_u3006, p1_u3005, p1_u3004, p1_u3003, p1_u3002, p1_u3001, p1_u3000, p1_u2999, p1_u2998, p1_u2997, p1_u2996, p1_u2995, p1_u2994, p1_u2993, p1_u2992, p1_u2991, p1_u2990, p1_u2989, p1_u2988, p1_u2987, p1_u2986, p1_u2985, p1_u2984, p1_u2983, p1_u2982, p1_u2981, p1_u2980, p1_u2979, p1_u2978, p1_u2977, p1_u2976, p1_u2975, p1_u2974, p1_u2973, p1_u2972, p1_u2971, p1_u2970, p1_u2969, p1_u2968, p1_u2967, p1_u2966, p1_u2965, p1_u2964, p1_u2963, p1_u2962, p1_u2961, p1_u2960, p1_u2959, p1_u2958, p1_u2957, p1_u2956, p1_u2955, p1_u2954, p1_u2953, p1_u2952, p1_u2951, p1_u2950, p1_u2949, p1_u2948, p1_u2947, p1_u2946, p1_u2945, p1_u2944, p1_u2943, p1_u2942, p1_u2941, p1_u2940, p1_u2939, p1_u2938, p1_u2937, p1_u2936, p1_u2935, p1_u2934, p1_u2933, p1_u2932, p1_u2931, p1_u2930, p1_u2929, p1_u2928, p1_u2927, p1_u2926, p1_u2925, p1_u2924, p1_u2923, p1_u2922, p1_u2921, p1_u2920, p1_u2919, p1_u2918, p1_u2917, p1_u2916, p1_u2915, p1_u2914, p1_u2913, p1_u2912, p1_u2911, p1_u2910, p1_u2909, p1_u2908, p1_u2907, p1_u2906, p1_u2905, p1_u2904, p1_u2903, p1_u2902, p1_u2901, p1_u2900, p1_u2899, p1_u2898, p1_u2897, p1_u2896, p1_u2895, p1_u2894, p1_u2893, p1_u2892, p1_u2891, p1_u2890, p1_u2889, p1_u2888, p1_u2887, p1_u2886, p1_u2885, p1_u2884, p1_u2883, p1_u2882, p1_u2881, p1_u2880, p1_u2879, p1_u2878, p1_u2877, p1_u2876, p1_u2875, p1_u2874, p1_u2873, p1_u2872, p1_u2871, p1_u2870, p1_u2869, p1_u2868, p1_u2867, p1_u2866, p1_u2865, p1_u2864, p1_u2863, p1_u2862, p1_u2861, p1_u2860, p1_u2859, p1_u2858, p1_u2857, p1_u2856, p1_u2855, p1_u2854, p1_u2853, p1_u2852, p1_u2851, p1_u2850, p1_u2849, p1_u2848, p1_u2847, p1_u2846, p1_u2845, p1_u2844, p1_u2843, p1_u2842, p1_u2841, p1_u2840, p1_u2839, p1_u2838, p1_u2837, p1_u2836, p1_u2835, p1_u2834, p1_u2833, p1_u2832, p1_u2831, p1_u2830, p1_u2829, p1_u2828, p1_u2827, p1_u2826, p1_u2825, p1_u2824, p1_u2823, p1_u2822, p1_u2821, p1_u2820, p1_u2819, p1_u2818, p1_u2817, p1_u2816, p1_u2815, p1_u2814, p1_u2813, p1_u2812, p1_u2811, p1_u2810, p1_u2809, p1_u2808, p1_u3481, p1_u2807, p1_u3482, p1_u3483, p1_u2806, p1_u3484, p1_u2805, p1_u3485, p1_u2804, p1_u3486, p1_u2803, p1_u2802, p1_u3487, p1_u2801;
initial begin
	$readmemb(`in_file, input_vec_mem );
end

always #(`cycle/2) clk = ~clk;

b17_ras cc (.DATAI_31_(vec[1451]), .DATAI_30_(vec[1450]), .DATAI_29_(vec[1449]), .DATAI_28_(vec[1448]), .DATAI_27_(vec[1447]), .DATAI_26_(vec[1446]), .DATAI_25_(vec[1445]), .DATAI_24_(vec[1444]), .DATAI_23_(vec[1443]), .DATAI_22_(vec[1442]), .DATAI_21_(vec[1441]), .DATAI_20_(vec[1440]), .DATAI_19_(vec[1439]), .DATAI_18_(vec[1438]), .DATAI_17_(vec[1437]), .DATAI_16_(vec[1436]), .DATAI_15_(vec[1435]), .DATAI_14_(vec[1434]), .DATAI_13_(vec[1433]), .DATAI_12_(vec[1432]), .DATAI_11_(vec[1431]), .DATAI_10_(vec[1430]), .DATAI_9_(vec[1429]), .DATAI_8_(vec[1428]), .DATAI_7_(vec[1427]), .DATAI_6_(vec[1426]), .DATAI_5_(vec[1425]), .DATAI_4_(vec[1424]), .DATAI_3_(vec[1423]), .DATAI_2_(vec[1422]), .DATAI_1_(vec[1421]), .DATAI_0_(vec[1420]), .HOLD(vec[1419]), .NA(vec[1418]), .BS16(vec[1417]), .READY1(vec[1416]), .READY2(vec[1415]), .BUF1_REG_0_(vec[1414]), .BUF1_REG_1_(vec[1413]), .BUF1_REG_2_(vec[1412]), .BUF1_REG_3_(vec[1411]), .BUF1_REG_4_(vec[1410]), .BUF1_REG_5_(vec[1409]), .BUF1_REG_6_(vec[1408]), .BUF1_REG_7_(vec[1407]), .BUF1_REG_8_(vec[1406]), .BUF1_REG_9_(vec[1405]), .BUF1_REG_10_(vec[1404]), .BUF1_REG_11_(vec[1403]), .BUF1_REG_12_(vec[1402]), .BUF1_REG_13_(vec[1401]), .BUF1_REG_14_(vec[1400]), .BUF1_REG_15_(vec[1399]), .BUF1_REG_16_(vec[1398]), .BUF1_REG_17_(vec[1397]), .BUF1_REG_18_(vec[1396]), .BUF1_REG_19_(vec[1395]), .BUF1_REG_20_(vec[1394]), .BUF1_REG_21_(vec[1393]), .BUF1_REG_22_(vec[1392]), .BUF1_REG_23_(vec[1391]), .BUF1_REG_24_(vec[1390]), .BUF1_REG_25_(vec[1389]), .BUF1_REG_26_(vec[1388]), .BUF1_REG_27_(vec[1387]), .BUF1_REG_28_(vec[1386]), .BUF1_REG_29_(vec[1385]), .BUF1_REG_30_(vec[1384]), .BUF1_REG_31_(vec[1383]), .BUF2_REG_0_(vec[1382]), .BUF2_REG_1_(vec[1381]), .BUF2_REG_2_(vec[1380]), .BUF2_REG_3_(vec[1379]), .BUF2_REG_4_(vec[1378]), .BUF2_REG_5_(vec[1377]), .BUF2_REG_6_(vec[1376]), .BUF2_REG_7_(vec[1375]), .BUF2_REG_8_(vec[1374]), .BUF2_REG_9_(vec[1373]), .BUF2_REG_10_(vec[1372]), .BUF2_REG_11_(vec[1371]), .BUF2_REG_12_(vec[1370]), .BUF2_REG_13_(vec[1369]), .BUF2_REG_14_(vec[1368]), .BUF2_REG_15_(vec[1367]), .BUF2_REG_16_(vec[1366]), .BUF2_REG_17_(vec[1365]), .BUF2_REG_18_(vec[1364]), .BUF2_REG_19_(vec[1363]), .BUF2_REG_20_(vec[1362]), .BUF2_REG_21_(vec[1361]), .BUF2_REG_22_(vec[1360]), .BUF2_REG_23_(vec[1359]), .BUF2_REG_24_(vec[1358]), .BUF2_REG_25_(vec[1357]), .BUF2_REG_26_(vec[1356]), .BUF2_REG_27_(vec[1355]), .BUF2_REG_28_(vec[1354]), .BUF2_REG_29_(vec[1353]), .BUF2_REG_30_(vec[1352]), .BUF2_REG_31_(vec[1351]), .READY12_REG(vec[1350]), .READY21_REG(vec[1349]), .READY22_REG(vec[1348]), .READY11_REG(vec[1347]), .P3_BE_N_REG_3_(vec[1346]), .P3_BE_N_REG_2_(vec[1345]), .P3_BE_N_REG_1_(vec[1344]), .P3_BE_N_REG_0_(vec[1343]), .P3_ADDRESS_REG_29_(vec[1342]), .P3_ADDRESS_REG_28_(vec[1341]), .P3_ADDRESS_REG_27_(vec[1340]), .P3_ADDRESS_REG_26_(vec[1339]), .P3_ADDRESS_REG_25_(vec[1338]), .P3_ADDRESS_REG_24_(vec[1337]), .P3_ADDRESS_REG_23_(vec[1336]), .P3_ADDRESS_REG_22_(vec[1335]), .P3_ADDRESS_REG_21_(vec[1334]), .P3_ADDRESS_REG_20_(vec[1333]), .P3_ADDRESS_REG_19_(vec[1332]), .P3_ADDRESS_REG_18_(vec[1331]), .P3_ADDRESS_REG_17_(vec[1330]), .P3_ADDRESS_REG_16_(vec[1329]), .P3_ADDRESS_REG_15_(vec[1328]), .P3_ADDRESS_REG_14_(vec[1327]), .P3_ADDRESS_REG_13_(vec[1326]), .P3_ADDRESS_REG_12_(vec[1325]), .P3_ADDRESS_REG_11_(vec[1324]), .P3_ADDRESS_REG_10_(vec[1323]), .P3_ADDRESS_REG_9_(vec[1322]), .P3_ADDRESS_REG_8_(vec[1321]), .P3_ADDRESS_REG_7_(vec[1320]), .P3_ADDRESS_REG_6_(vec[1319]), .P3_ADDRESS_REG_5_(vec[1318]), .P3_ADDRESS_REG_4_(vec[1317]), .P3_ADDRESS_REG_3_(vec[1316]), .P3_ADDRESS_REG_2_(vec[1315]), .P3_ADDRESS_REG_1_(vec[1314]), .P3_ADDRESS_REG_0_(vec[1313]), .P3_STATE_REG_2_(vec[1312]), .P3_STATE_REG_1_(vec[1311]), .P3_STATE_REG_0_(vec[1310]), .P3_DATAWIDTH_REG_0_(vec[1309]), .P3_DATAWIDTH_REG_1_(vec[1308]), .P3_DATAWIDTH_REG_2_(vec[1307]), .P3_DATAWIDTH_REG_3_(vec[1306]), .P3_DATAWIDTH_REG_4_(vec[1305]), .P3_DATAWIDTH_REG_5_(vec[1304]), .P3_DATAWIDTH_REG_6_(vec[1303]), .P3_DATAWIDTH_REG_7_(vec[1302]), .P3_DATAWIDTH_REG_8_(vec[1301]), .P3_DATAWIDTH_REG_9_(vec[1300]), .P3_DATAWIDTH_REG_10_(vec[1299]), .P3_DATAWIDTH_REG_11_(vec[1298]), .P3_DATAWIDTH_REG_12_(vec[1297]), .P3_DATAWIDTH_REG_13_(vec[1296]), .P3_DATAWIDTH_REG_14_(vec[1295]), .P3_DATAWIDTH_REG_15_(vec[1294]), .P3_DATAWIDTH_REG_16_(vec[1293]), .P3_DATAWIDTH_REG_17_(vec[1292]), .P3_DATAWIDTH_REG_18_(vec[1291]), .P3_DATAWIDTH_REG_19_(vec[1290]), .P3_DATAWIDTH_REG_20_(vec[1289]), .P3_DATAWIDTH_REG_21_(vec[1288]), .P3_DATAWIDTH_REG_22_(vec[1287]), .P3_DATAWIDTH_REG_23_(vec[1286]), .P3_DATAWIDTH_REG_24_(vec[1285]), .P3_DATAWIDTH_REG_25_(vec[1284]), .P3_DATAWIDTH_REG_26_(vec[1283]), .P3_DATAWIDTH_REG_27_(vec[1282]), .P3_DATAWIDTH_REG_28_(vec[1281]), .P3_DATAWIDTH_REG_29_(vec[1280]), .P3_DATAWIDTH_REG_30_(vec[1279]), .P3_DATAWIDTH_REG_31_(vec[1278]), .P3_STATE2_REG_3_(vec[1277]), .P3_STATE2_REG_2_(vec[1276]), .P3_STATE2_REG_1_(vec[1275]), .P3_STATE2_REG_0_(vec[1274]), .P3_INSTQUEUE_REG_15__7_(vec[1273]), .P3_INSTQUEUE_REG_15__6_(vec[1272]), .P3_INSTQUEUE_REG_15__5_(vec[1271]), .P3_INSTQUEUE_REG_15__4_(vec[1270]), .P3_INSTQUEUE_REG_15__3_(vec[1269]), .P3_INSTQUEUE_REG_15__2_(vec[1268]), .P3_INSTQUEUE_REG_15__1_(vec[1267]), .P3_INSTQUEUE_REG_15__0_(vec[1266]), .P3_INSTQUEUE_REG_14__7_(vec[1265]), .P3_INSTQUEUE_REG_14__6_(vec[1264]), .P3_INSTQUEUE_REG_14__5_(vec[1263]), .P3_INSTQUEUE_REG_14__4_(vec[1262]), .P3_INSTQUEUE_REG_14__3_(vec[1261]), .P3_INSTQUEUE_REG_14__2_(vec[1260]), .P3_INSTQUEUE_REG_14__1_(vec[1259]), .P3_INSTQUEUE_REG_14__0_(vec[1258]), .P3_INSTQUEUE_REG_13__7_(vec[1257]), .P3_INSTQUEUE_REG_13__6_(vec[1256]), .P3_INSTQUEUE_REG_13__5_(vec[1255]), .P3_INSTQUEUE_REG_13__4_(vec[1254]), .P3_INSTQUEUE_REG_13__3_(vec[1253]), .P3_INSTQUEUE_REG_13__2_(vec[1252]), .P3_INSTQUEUE_REG_13__1_(vec[1251]), .P3_INSTQUEUE_REG_13__0_(vec[1250]), .P3_INSTQUEUE_REG_12__7_(vec[1249]), .P3_INSTQUEUE_REG_12__6_(vec[1248]), .P3_INSTQUEUE_REG_12__5_(vec[1247]), .P3_INSTQUEUE_REG_12__4_(vec[1246]), .P3_INSTQUEUE_REG_12__3_(vec[1245]), .P3_INSTQUEUE_REG_12__2_(vec[1244]), .P3_INSTQUEUE_REG_12__1_(vec[1243]), .P3_INSTQUEUE_REG_12__0_(vec[1242]), .P3_INSTQUEUE_REG_11__7_(vec[1241]), .P3_INSTQUEUE_REG_11__6_(vec[1240]), .P3_INSTQUEUE_REG_11__5_(vec[1239]), .P3_INSTQUEUE_REG_11__4_(vec[1238]), .P3_INSTQUEUE_REG_11__3_(vec[1237]), .P3_INSTQUEUE_REG_11__2_(vec[1236]), .P3_INSTQUEUE_REG_11__1_(vec[1235]), .P3_INSTQUEUE_REG_11__0_(vec[1234]), .P3_INSTQUEUE_REG_10__7_(vec[1233]), .P3_INSTQUEUE_REG_10__6_(vec[1232]), .P3_INSTQUEUE_REG_10__5_(vec[1231]), .P3_INSTQUEUE_REG_10__4_(vec[1230]), .P3_INSTQUEUE_REG_10__3_(vec[1229]), .P3_INSTQUEUE_REG_10__2_(vec[1228]), .P3_INSTQUEUE_REG_10__1_(vec[1227]), .P3_INSTQUEUE_REG_10__0_(vec[1226]), .P3_INSTQUEUE_REG_9__7_(vec[1225]), .P3_INSTQUEUE_REG_9__6_(vec[1224]), .P3_INSTQUEUE_REG_9__5_(vec[1223]), .P3_INSTQUEUE_REG_9__4_(vec[1222]), .P3_INSTQUEUE_REG_9__3_(vec[1221]), .P3_INSTQUEUE_REG_9__2_(vec[1220]), .P3_INSTQUEUE_REG_9__1_(vec[1219]), .P3_INSTQUEUE_REG_9__0_(vec[1218]), .P3_INSTQUEUE_REG_8__7_(vec[1217]), .P3_INSTQUEUE_REG_8__6_(vec[1216]), .P3_INSTQUEUE_REG_8__5_(vec[1215]), .P3_INSTQUEUE_REG_8__4_(vec[1214]), .P3_INSTQUEUE_REG_8__3_(vec[1213]), .P3_INSTQUEUE_REG_8__2_(vec[1212]), .P3_INSTQUEUE_REG_8__1_(vec[1211]), .P3_INSTQUEUE_REG_8__0_(vec[1210]), .P3_INSTQUEUE_REG_7__7_(vec[1209]), .P3_INSTQUEUE_REG_7__6_(vec[1208]), .P3_INSTQUEUE_REG_7__5_(vec[1207]), .P3_INSTQUEUE_REG_7__4_(vec[1206]), .P3_INSTQUEUE_REG_7__3_(vec[1205]), .P3_INSTQUEUE_REG_7__2_(vec[1204]), .P3_INSTQUEUE_REG_7__1_(vec[1203]), .P3_INSTQUEUE_REG_7__0_(vec[1202]), .P3_INSTQUEUE_REG_6__7_(vec[1201]), .P3_INSTQUEUE_REG_6__6_(vec[1200]), .P3_INSTQUEUE_REG_6__5_(vec[1199]), .P3_INSTQUEUE_REG_6__4_(vec[1198]), .P3_INSTQUEUE_REG_6__3_(vec[1197]), .P3_INSTQUEUE_REG_6__2_(vec[1196]), .P3_INSTQUEUE_REG_6__1_(vec[1195]), .P3_INSTQUEUE_REG_6__0_(vec[1194]), .P3_INSTQUEUE_REG_5__7_(vec[1193]), .P3_INSTQUEUE_REG_5__6_(vec[1192]), .P3_INSTQUEUE_REG_5__5_(vec[1191]), .P3_INSTQUEUE_REG_5__4_(vec[1190]), .P3_INSTQUEUE_REG_5__3_(vec[1189]), .P3_INSTQUEUE_REG_5__2_(vec[1188]), .P3_INSTQUEUE_REG_5__1_(vec[1187]), .P3_INSTQUEUE_REG_5__0_(vec[1186]), .P3_INSTQUEUE_REG_4__7_(vec[1185]), .P3_INSTQUEUE_REG_4__6_(vec[1184]), .P3_INSTQUEUE_REG_4__5_(vec[1183]), .P3_INSTQUEUE_REG_4__4_(vec[1182]), .P3_INSTQUEUE_REG_4__3_(vec[1181]), .P3_INSTQUEUE_REG_4__2_(vec[1180]), .P3_INSTQUEUE_REG_4__1_(vec[1179]), .P3_INSTQUEUE_REG_4__0_(vec[1178]), .P3_INSTQUEUE_REG_3__7_(vec[1177]), .P3_INSTQUEUE_REG_3__6_(vec[1176]), .P3_INSTQUEUE_REG_3__5_(vec[1175]), .P3_INSTQUEUE_REG_3__4_(vec[1174]), .P3_INSTQUEUE_REG_3__3_(vec[1173]), .P3_INSTQUEUE_REG_3__2_(vec[1172]), .P3_INSTQUEUE_REG_3__1_(vec[1171]), .P3_INSTQUEUE_REG_3__0_(vec[1170]), .P3_INSTQUEUE_REG_2__7_(vec[1169]), .P3_INSTQUEUE_REG_2__6_(vec[1168]), .P3_INSTQUEUE_REG_2__5_(vec[1167]), .P3_INSTQUEUE_REG_2__4_(vec[1166]), .P3_INSTQUEUE_REG_2__3_(vec[1165]), .P3_INSTQUEUE_REG_2__2_(vec[1164]), .P3_INSTQUEUE_REG_2__1_(vec[1163]), .P3_INSTQUEUE_REG_2__0_(vec[1162]), .P3_INSTQUEUE_REG_1__7_(vec[1161]), .P3_INSTQUEUE_REG_1__6_(vec[1160]), .P3_INSTQUEUE_REG_1__5_(vec[1159]), .P3_INSTQUEUE_REG_1__4_(vec[1158]), .P3_INSTQUEUE_REG_1__3_(vec[1157]), .P3_INSTQUEUE_REG_1__2_(vec[1156]), .P3_INSTQUEUE_REG_1__1_(vec[1155]), .P3_INSTQUEUE_REG_1__0_(vec[1154]), .P3_INSTQUEUE_REG_0__7_(vec[1153]), .P3_INSTQUEUE_REG_0__6_(vec[1152]), .P3_INSTQUEUE_REG_0__5_(vec[1151]), .P3_INSTQUEUE_REG_0__4_(vec[1150]), .P3_INSTQUEUE_REG_0__3_(vec[1149]), .P3_INSTQUEUE_REG_0__2_(vec[1148]), .P3_INSTQUEUE_REG_0__1_(vec[1147]), .P3_INSTQUEUE_REG_0__0_(vec[1146]), .P3_INSTQUEUERD_ADDR_REG_4_(vec[1145]), .P3_INSTQUEUERD_ADDR_REG_3_(vec[1144]), .P3_INSTQUEUERD_ADDR_REG_2_(vec[1143]), .P3_INSTQUEUERD_ADDR_REG_1_(vec[1142]), .P3_INSTQUEUERD_ADDR_REG_0_(vec[1141]), .P3_INSTQUEUEWR_ADDR_REG_4_(vec[1140]), .P3_INSTQUEUEWR_ADDR_REG_3_(vec[1139]), .P3_INSTQUEUEWR_ADDR_REG_2_(vec[1138]), .P3_INSTQUEUEWR_ADDR_REG_1_(vec[1137]), .P3_INSTQUEUEWR_ADDR_REG_0_(vec[1136]), .P3_INSTADDRPOINTER_REG_0_(vec[1135]), .P3_INSTADDRPOINTER_REG_1_(vec[1134]), .P3_INSTADDRPOINTER_REG_2_(vec[1133]), .P3_INSTADDRPOINTER_REG_3_(vec[1132]), .P3_INSTADDRPOINTER_REG_4_(vec[1131]), .P3_INSTADDRPOINTER_REG_5_(vec[1130]), .P3_INSTADDRPOINTER_REG_6_(vec[1129]), .P3_INSTADDRPOINTER_REG_7_(vec[1128]), .P3_INSTADDRPOINTER_REG_8_(vec[1127]), .P3_INSTADDRPOINTER_REG_9_(vec[1126]), .P3_INSTADDRPOINTER_REG_10_(vec[1125]), .P3_INSTADDRPOINTER_REG_11_(vec[1124]), .P3_INSTADDRPOINTER_REG_12_(vec[1123]), .P3_INSTADDRPOINTER_REG_13_(vec[1122]), .P3_INSTADDRPOINTER_REG_14_(vec[1121]), .P3_INSTADDRPOINTER_REG_15_(vec[1120]), .P3_INSTADDRPOINTER_REG_16_(vec[1119]), .P3_INSTADDRPOINTER_REG_17_(vec[1118]), .P3_INSTADDRPOINTER_REG_18_(vec[1117]), .P3_INSTADDRPOINTER_REG_19_(vec[1116]), .P3_INSTADDRPOINTER_REG_20_(vec[1115]), .P3_INSTADDRPOINTER_REG_21_(vec[1114]), .P3_INSTADDRPOINTER_REG_22_(vec[1113]), .P3_INSTADDRPOINTER_REG_23_(vec[1112]), .P3_INSTADDRPOINTER_REG_24_(vec[1111]), .P3_INSTADDRPOINTER_REG_25_(vec[1110]), .P3_INSTADDRPOINTER_REG_26_(vec[1109]), .P3_INSTADDRPOINTER_REG_27_(vec[1108]), .P3_INSTADDRPOINTER_REG_28_(vec[1107]), .P3_INSTADDRPOINTER_REG_29_(vec[1106]), .P3_INSTADDRPOINTER_REG_30_(vec[1105]), .P3_INSTADDRPOINTER_REG_31_(vec[1104]), .P3_PHYADDRPOINTER_REG_0_(vec[1103]), .P3_PHYADDRPOINTER_REG_1_(vec[1102]), .P3_PHYADDRPOINTER_REG_2_(vec[1101]), .P3_PHYADDRPOINTER_REG_3_(vec[1100]), .P3_PHYADDRPOINTER_REG_4_(vec[1099]), .P3_PHYADDRPOINTER_REG_5_(vec[1098]), .P3_PHYADDRPOINTER_REG_6_(vec[1097]), .P3_PHYADDRPOINTER_REG_7_(vec[1096]), .P3_PHYADDRPOINTER_REG_8_(vec[1095]), .P3_PHYADDRPOINTER_REG_9_(vec[1094]), .P3_PHYADDRPOINTER_REG_10_(vec[1093]), .P3_PHYADDRPOINTER_REG_11_(vec[1092]), .P3_PHYADDRPOINTER_REG_12_(vec[1091]), .P3_PHYADDRPOINTER_REG_13_(vec[1090]), .P3_PHYADDRPOINTER_REG_14_(vec[1089]), .P3_PHYADDRPOINTER_REG_15_(vec[1088]), .P3_PHYADDRPOINTER_REG_16_(vec[1087]), .P3_PHYADDRPOINTER_REG_17_(vec[1086]), .P3_PHYADDRPOINTER_REG_18_(vec[1085]), .P3_PHYADDRPOINTER_REG_19_(vec[1084]), .P3_PHYADDRPOINTER_REG_20_(vec[1083]), .P3_PHYADDRPOINTER_REG_21_(vec[1082]), .P3_PHYADDRPOINTER_REG_22_(vec[1081]), .P3_PHYADDRPOINTER_REG_23_(vec[1080]), .P3_PHYADDRPOINTER_REG_24_(vec[1079]), .P3_PHYADDRPOINTER_REG_25_(vec[1078]), .P3_PHYADDRPOINTER_REG_26_(vec[1077]), .P3_PHYADDRPOINTER_REG_27_(vec[1076]), .P3_PHYADDRPOINTER_REG_28_(vec[1075]), .P3_PHYADDRPOINTER_REG_29_(vec[1074]), .P3_PHYADDRPOINTER_REG_30_(vec[1073]), .P3_PHYADDRPOINTER_REG_31_(vec[1072]), .P3_LWORD_REG_15_(vec[1071]), .P3_LWORD_REG_14_(vec[1070]), .P3_LWORD_REG_13_(vec[1069]), .P3_LWORD_REG_12_(vec[1068]), .P3_LWORD_REG_11_(vec[1067]), .P3_LWORD_REG_10_(vec[1066]), .P3_LWORD_REG_9_(vec[1065]), .P3_LWORD_REG_8_(vec[1064]), .P3_LWORD_REG_7_(vec[1063]), .P3_LWORD_REG_6_(vec[1062]), .P3_LWORD_REG_5_(vec[1061]), .P3_LWORD_REG_4_(vec[1060]), .P3_LWORD_REG_3_(vec[1059]), .P3_LWORD_REG_2_(vec[1058]), .P3_LWORD_REG_1_(vec[1057]), .P3_LWORD_REG_0_(vec[1056]), .P3_UWORD_REG_14_(vec[1055]), .P3_UWORD_REG_13_(vec[1054]), .P3_UWORD_REG_12_(vec[1053]), .P3_UWORD_REG_11_(vec[1052]), .P3_UWORD_REG_10_(vec[1051]), .P3_UWORD_REG_9_(vec[1050]), .P3_UWORD_REG_8_(vec[1049]), .P3_UWORD_REG_7_(vec[1048]), .P3_UWORD_REG_6_(vec[1047]), .P3_UWORD_REG_5_(vec[1046]), .P3_UWORD_REG_4_(vec[1045]), .P3_UWORD_REG_3_(vec[1044]), .P3_UWORD_REG_2_(vec[1043]), .P3_UWORD_REG_1_(vec[1042]), .P3_UWORD_REG_0_(vec[1041]), .P3_DATAO_REG_0__EXTRA(vec[1040]), .P3_DATAO_REG_1__EXTRA(vec[1039]), .P3_DATAO_REG_2__EXTRA(vec[1038]), .P3_DATAO_REG_3__EXTRA(vec[1037]), .P3_DATAO_REG_4__EXTRA(vec[1036]), .P3_DATAO_REG_5__EXTRA(vec[1035]), .P3_DATAO_REG_6__EXTRA(vec[1034]), .P3_DATAO_REG_7__EXTRA(vec[1033]), .P3_DATAO_REG_8__EXTRA(vec[1032]), .P3_DATAO_REG_9__EXTRA(vec[1031]), .P3_DATAO_REG_10__EXTRA(vec[1030]), .P3_DATAO_REG_11__EXTRA(vec[1029]), .P3_DATAO_REG_12__EXTRA(vec[1028]), .P3_DATAO_REG_13__EXTRA(vec[1027]), .P3_DATAO_REG_14__EXTRA(vec[1026]), .P3_DATAO_REG_15__EXTRA(vec[1025]), .P3_DATAO_REG_16__EXTRA(vec[1024]), .P3_DATAO_REG_17__EXTRA(vec[1023]), .P3_DATAO_REG_18__EXTRA(vec[1022]), .P3_DATAO_REG_19__EXTRA(vec[1021]), .P3_DATAO_REG_20__EXTRA(vec[1020]), .P3_DATAO_REG_21__EXTRA(vec[1019]), .P3_DATAO_REG_22__EXTRA(vec[1018]), .P3_DATAO_REG_23__EXTRA(vec[1017]), .P3_DATAO_REG_24__EXTRA(vec[1016]), .P3_DATAO_REG_25__EXTRA(vec[1015]), .P3_DATAO_REG_26__EXTRA(vec[1014]), .P3_DATAO_REG_27__EXTRA(vec[1013]), .P3_DATAO_REG_28__EXTRA(vec[1012]), .P3_DATAO_REG_29__EXTRA(vec[1011]), .P3_DATAO_REG_30__EXTRA(vec[1010]), .P3_DATAO_REG_31__EXTRA(vec[1009]), .P3_EAX_REG_0_(vec[1008]), .P3_EAX_REG_1_(vec[1007]), .P3_EAX_REG_2_(vec[1006]), .P3_EAX_REG_3_(vec[1005]), .P3_EAX_REG_4_(vec[1004]), .P3_EAX_REG_5_(vec[1003]), .P3_EAX_REG_6_(vec[1002]), .P3_EAX_REG_7_(vec[1001]), .P3_EAX_REG_8_(vec[1000]), .P3_EAX_REG_9_(vec[999]), .P3_EAX_REG_10_(vec[998]), .P3_EAX_REG_11_(vec[997]), .P3_EAX_REG_12_(vec[996]), .P3_EAX_REG_13_(vec[995]), .P3_EAX_REG_14_(vec[994]), .P3_EAX_REG_15_(vec[993]), .P3_EAX_REG_16_(vec[992]), .P3_EAX_REG_17_(vec[991]), .P3_EAX_REG_18_(vec[990]), .P3_EAX_REG_19_(vec[989]), .P3_EAX_REG_20_(vec[988]), .P3_EAX_REG_21_(vec[987]), .P3_EAX_REG_22_(vec[986]), .P3_EAX_REG_23_(vec[985]), .P3_EAX_REG_24_(vec[984]), .P3_EAX_REG_25_(vec[983]), .P3_EAX_REG_26_(vec[982]), .P3_EAX_REG_27_(vec[981]), .P3_EAX_REG_28_(vec[980]), .P3_EAX_REG_29_(vec[979]), .P3_EAX_REG_30_(vec[978]), .P3_EAX_REG_31_(vec[977]), .P3_EBX_REG_0_(vec[976]), .P3_EBX_REG_1_(vec[975]), .P3_EBX_REG_2_(vec[974]), .P3_EBX_REG_3_(vec[973]), .P3_EBX_REG_4_(vec[972]), .P3_EBX_REG_5_(vec[971]), .P3_EBX_REG_6_(vec[970]), .P3_EBX_REG_7_(vec[969]), .P3_EBX_REG_8_(vec[968]), .P3_EBX_REG_9_(vec[967]), .P3_EBX_REG_10_(vec[966]), .P3_EBX_REG_11_(vec[965]), .P3_EBX_REG_12_(vec[964]), .P3_EBX_REG_13_(vec[963]), .P3_EBX_REG_14_(vec[962]), .P3_EBX_REG_15_(vec[961]), .P3_EBX_REG_16_(vec[960]), .P3_EBX_REG_17_(vec[959]), .P3_EBX_REG_18_(vec[958]), .P3_EBX_REG_19_(vec[957]), .P3_EBX_REG_20_(vec[956]), .P3_EBX_REG_21_(vec[955]), .P3_EBX_REG_22_(vec[954]), .P3_EBX_REG_23_(vec[953]), .P3_EBX_REG_24_(vec[952]), .P3_EBX_REG_25_(vec[951]), .P3_EBX_REG_26_(vec[950]), .P3_EBX_REG_27_(vec[949]), .P3_EBX_REG_28_(vec[948]), .P3_EBX_REG_29_(vec[947]), .P3_EBX_REG_30_(vec[946]), .P3_EBX_REG_31_(vec[945]), .P3_REIP_REG_0_(vec[944]), .P3_REIP_REG_1_(vec[943]), .P3_REIP_REG_2_(vec[942]), .P3_REIP_REG_3_(vec[941]), .P3_REIP_REG_4_(vec[940]), .P3_REIP_REG_5_(vec[939]), .P3_REIP_REG_6_(vec[938]), .P3_REIP_REG_7_(vec[937]), .P3_REIP_REG_8_(vec[936]), .P3_REIP_REG_9_(vec[935]), .P3_REIP_REG_10_(vec[934]), .P3_REIP_REG_11_(vec[933]), .P3_REIP_REG_12_(vec[932]), .P3_REIP_REG_13_(vec[931]), .P3_REIP_REG_14_(vec[930]), .P3_REIP_REG_15_(vec[929]), .P3_REIP_REG_16_(vec[928]), .P3_REIP_REG_17_(vec[927]), .P3_REIP_REG_18_(vec[926]), .P3_REIP_REG_19_(vec[925]), .P3_REIP_REG_20_(vec[924]), .P3_REIP_REG_21_(vec[923]), .P3_REIP_REG_22_(vec[922]), .P3_REIP_REG_23_(vec[921]), .P3_REIP_REG_24_(vec[920]), .P3_REIP_REG_25_(vec[919]), .P3_REIP_REG_26_(vec[918]), .P3_REIP_REG_27_(vec[917]), .P3_REIP_REG_28_(vec[916]), .P3_REIP_REG_29_(vec[915]), .P3_REIP_REG_30_(vec[914]), .P3_REIP_REG_31_(vec[913]), .P3_BYTEENABLE_REG_3_(vec[912]), .P3_BYTEENABLE_REG_2_(vec[911]), .P3_BYTEENABLE_REG_1_(vec[910]), .P3_BYTEENABLE_REG_0_(vec[909]), .P3_W_R_N_REG_EXTRA(vec[908]), .P3_FLUSH_REG(vec[907]), .P3_MORE_REG(vec[906]), .P3_STATEBS16_REG(vec[905]), .P3_REQUESTPENDING_REG(vec[904]), .P3_D_C_N_REG_EXTRA(vec[903]), .P3_M_IO_N_REG_EXTRA(vec[902]), .P3_CODEFETCH_REG(vec[901]), .P3_ADS_N_REG_EXTRA(vec[900]), .P3_READREQUEST_REG(vec[899]), .P3_MEMORYFETCH_REG(vec[898]), .P2_BE_N_REG_3_(vec[897]), .P2_BE_N_REG_2_(vec[896]), .P2_BE_N_REG_1_(vec[895]), .P2_BE_N_REG_0_(vec[894]), .P2_ADDRESS_REG_29_(vec[893]), .P2_ADDRESS_REG_28_(vec[892]), .P2_ADDRESS_REG_27_(vec[891]), .P2_ADDRESS_REG_26_(vec[890]), .P2_ADDRESS_REG_25_(vec[889]), .P2_ADDRESS_REG_24_(vec[888]), .P2_ADDRESS_REG_23_(vec[887]), .P2_ADDRESS_REG_22_(vec[886]), .P2_ADDRESS_REG_21_(vec[885]), .P2_ADDRESS_REG_20_(vec[884]), .P2_ADDRESS_REG_19_(vec[883]), .P2_ADDRESS_REG_18_(vec[882]), .P2_ADDRESS_REG_17_(vec[881]), .P2_ADDRESS_REG_16_(vec[880]), .P2_ADDRESS_REG_15_(vec[879]), .P2_ADDRESS_REG_14_(vec[878]), .P2_ADDRESS_REG_13_(vec[877]), .P2_ADDRESS_REG_12_(vec[876]), .P2_ADDRESS_REG_11_(vec[875]), .P2_ADDRESS_REG_10_(vec[874]), .P2_ADDRESS_REG_9_(vec[873]), .P2_ADDRESS_REG_8_(vec[872]), .P2_ADDRESS_REG_7_(vec[871]), .P2_ADDRESS_REG_6_(vec[870]), .P2_ADDRESS_REG_5_(vec[869]), .P2_ADDRESS_REG_4_(vec[868]), .P2_ADDRESS_REG_3_(vec[867]), .P2_ADDRESS_REG_2_(vec[866]), .P2_ADDRESS_REG_1_(vec[865]), .P2_ADDRESS_REG_0_(vec[864]), .P2_STATE_REG_2_(vec[863]), .P2_STATE_REG_1_(vec[862]), .P2_STATE_REG_0_(vec[861]), .P2_DATAWIDTH_REG_0_(vec[860]), .P2_DATAWIDTH_REG_1_(vec[859]), .P2_DATAWIDTH_REG_2_(vec[858]), .P2_DATAWIDTH_REG_3_(vec[857]), .P2_DATAWIDTH_REG_4_(vec[856]), .P2_DATAWIDTH_REG_5_(vec[855]), .P2_DATAWIDTH_REG_6_(vec[854]), .P2_DATAWIDTH_REG_7_(vec[853]), .P2_DATAWIDTH_REG_8_(vec[852]), .P2_DATAWIDTH_REG_9_(vec[851]), .P2_DATAWIDTH_REG_10_(vec[850]), .P2_DATAWIDTH_REG_11_(vec[849]), .P2_DATAWIDTH_REG_12_(vec[848]), .P2_DATAWIDTH_REG_13_(vec[847]), .P2_DATAWIDTH_REG_14_(vec[846]), .P2_DATAWIDTH_REG_15_(vec[845]), .P2_DATAWIDTH_REG_16_(vec[844]), .P2_DATAWIDTH_REG_17_(vec[843]), .P2_DATAWIDTH_REG_18_(vec[842]), .P2_DATAWIDTH_REG_19_(vec[841]), .P2_DATAWIDTH_REG_20_(vec[840]), .P2_DATAWIDTH_REG_21_(vec[839]), .P2_DATAWIDTH_REG_22_(vec[838]), .P2_DATAWIDTH_REG_23_(vec[837]), .P2_DATAWIDTH_REG_24_(vec[836]), .P2_DATAWIDTH_REG_25_(vec[835]), .P2_DATAWIDTH_REG_26_(vec[834]), .P2_DATAWIDTH_REG_27_(vec[833]), .P2_DATAWIDTH_REG_28_(vec[832]), .P2_DATAWIDTH_REG_29_(vec[831]), .P2_DATAWIDTH_REG_30_(vec[830]), .P2_DATAWIDTH_REG_31_(vec[829]), .P2_STATE2_REG_3_(vec[828]), .P2_STATE2_REG_2_(vec[827]), .P2_STATE2_REG_1_(vec[826]), .P2_STATE2_REG_0_(vec[825]), .P2_INSTQUEUE_REG_15__7_(vec[824]), .P2_INSTQUEUE_REG_15__6_(vec[823]), .P2_INSTQUEUE_REG_15__5_(vec[822]), .P2_INSTQUEUE_REG_15__4_(vec[821]), .P2_INSTQUEUE_REG_15__3_(vec[820]), .P2_INSTQUEUE_REG_15__2_(vec[819]), .P2_INSTQUEUE_REG_15__1_(vec[818]), .P2_INSTQUEUE_REG_15__0_(vec[817]), .P2_INSTQUEUE_REG_14__7_(vec[816]), .P2_INSTQUEUE_REG_14__6_(vec[815]), .P2_INSTQUEUE_REG_14__5_(vec[814]), .P2_INSTQUEUE_REG_14__4_(vec[813]), .P2_INSTQUEUE_REG_14__3_(vec[812]), .P2_INSTQUEUE_REG_14__2_(vec[811]), .P2_INSTQUEUE_REG_14__1_(vec[810]), .P2_INSTQUEUE_REG_14__0_(vec[809]), .P2_INSTQUEUE_REG_13__7_(vec[808]), .P2_INSTQUEUE_REG_13__6_(vec[807]), .P2_INSTQUEUE_REG_13__5_(vec[806]), .P2_INSTQUEUE_REG_13__4_(vec[805]), .P2_INSTQUEUE_REG_13__3_(vec[804]), .P2_INSTQUEUE_REG_13__2_(vec[803]), .P2_INSTQUEUE_REG_13__1_(vec[802]), .P2_INSTQUEUE_REG_13__0_(vec[801]), .P2_INSTQUEUE_REG_12__7_(vec[800]), .P2_INSTQUEUE_REG_12__6_(vec[799]), .P2_INSTQUEUE_REG_12__5_(vec[798]), .P2_INSTQUEUE_REG_12__4_(vec[797]), .P2_INSTQUEUE_REG_12__3_(vec[796]), .P2_INSTQUEUE_REG_12__2_(vec[795]), .P2_INSTQUEUE_REG_12__1_(vec[794]), .P2_INSTQUEUE_REG_12__0_(vec[793]), .P2_INSTQUEUE_REG_11__7_(vec[792]), .P2_INSTQUEUE_REG_11__6_(vec[791]), .P2_INSTQUEUE_REG_11__5_(vec[790]), .P2_INSTQUEUE_REG_11__4_(vec[789]), .P2_INSTQUEUE_REG_11__3_(vec[788]), .P2_INSTQUEUE_REG_11__2_(vec[787]), .P2_INSTQUEUE_REG_11__1_(vec[786]), .P2_INSTQUEUE_REG_11__0_(vec[785]), .P2_INSTQUEUE_REG_10__7_(vec[784]), .P2_INSTQUEUE_REG_10__6_(vec[783]), .P2_INSTQUEUE_REG_10__5_(vec[782]), .P2_INSTQUEUE_REG_10__4_(vec[781]), .P2_INSTQUEUE_REG_10__3_(vec[780]), .P2_INSTQUEUE_REG_10__2_(vec[779]), .P2_INSTQUEUE_REG_10__1_(vec[778]), .P2_INSTQUEUE_REG_10__0_(vec[777]), .P2_INSTQUEUE_REG_9__7_(vec[776]), .P2_INSTQUEUE_REG_9__6_(vec[775]), .P2_INSTQUEUE_REG_9__5_(vec[774]), .P2_INSTQUEUE_REG_9__4_(vec[773]), .P2_INSTQUEUE_REG_9__3_(vec[772]), .P2_INSTQUEUE_REG_9__2_(vec[771]), .P2_INSTQUEUE_REG_9__1_(vec[770]), .P2_INSTQUEUE_REG_9__0_(vec[769]), .P2_INSTQUEUE_REG_8__7_(vec[768]), .P2_INSTQUEUE_REG_8__6_(vec[767]), .P2_INSTQUEUE_REG_8__5_(vec[766]), .P2_INSTQUEUE_REG_8__4_(vec[765]), .P2_INSTQUEUE_REG_8__3_(vec[764]), .P2_INSTQUEUE_REG_8__2_(vec[763]), .P2_INSTQUEUE_REG_8__1_(vec[762]), .P2_INSTQUEUE_REG_8__0_(vec[761]), .P2_INSTQUEUE_REG_7__7_(vec[760]), .P2_INSTQUEUE_REG_7__6_(vec[759]), .P2_INSTQUEUE_REG_7__5_(vec[758]), .P2_INSTQUEUE_REG_7__4_(vec[757]), .P2_INSTQUEUE_REG_7__3_(vec[756]), .P2_INSTQUEUE_REG_7__2_(vec[755]), .P2_INSTQUEUE_REG_7__1_(vec[754]), .P2_INSTQUEUE_REG_7__0_(vec[753]), .P2_INSTQUEUE_REG_6__7_(vec[752]), .P2_INSTQUEUE_REG_6__6_(vec[751]), .P2_INSTQUEUE_REG_6__5_(vec[750]), .P2_INSTQUEUE_REG_6__4_(vec[749]), .P2_INSTQUEUE_REG_6__3_(vec[748]), .P2_INSTQUEUE_REG_6__2_(vec[747]), .P2_INSTQUEUE_REG_6__1_(vec[746]), .P2_INSTQUEUE_REG_6__0_(vec[745]), .P2_INSTQUEUE_REG_5__7_(vec[744]), .P2_INSTQUEUE_REG_5__6_(vec[743]), .P2_INSTQUEUE_REG_5__5_(vec[742]), .P2_INSTQUEUE_REG_5__4_(vec[741]), .P2_INSTQUEUE_REG_5__3_(vec[740]), .P2_INSTQUEUE_REG_5__2_(vec[739]), .P2_INSTQUEUE_REG_5__1_(vec[738]), .P2_INSTQUEUE_REG_5__0_(vec[737]), .P2_INSTQUEUE_REG_4__7_(vec[736]), .P2_INSTQUEUE_REG_4__6_(vec[735]), .P2_INSTQUEUE_REG_4__5_(vec[734]), .P2_INSTQUEUE_REG_4__4_(vec[733]), .P2_INSTQUEUE_REG_4__3_(vec[732]), .P2_INSTQUEUE_REG_4__2_(vec[731]), .P2_INSTQUEUE_REG_4__1_(vec[730]), .P2_INSTQUEUE_REG_4__0_(vec[729]), .P2_INSTQUEUE_REG_3__7_(vec[728]), .P2_INSTQUEUE_REG_3__6_(vec[727]), .P2_INSTQUEUE_REG_3__5_(vec[726]), .P2_INSTQUEUE_REG_3__4_(vec[725]), .P2_INSTQUEUE_REG_3__3_(vec[724]), .P2_INSTQUEUE_REG_3__2_(vec[723]), .P2_INSTQUEUE_REG_3__1_(vec[722]), .P2_INSTQUEUE_REG_3__0_(vec[721]), .P2_INSTQUEUE_REG_2__7_(vec[720]), .P2_INSTQUEUE_REG_2__6_(vec[719]), .P2_INSTQUEUE_REG_2__5_(vec[718]), .P2_INSTQUEUE_REG_2__4_(vec[717]), .P2_INSTQUEUE_REG_2__3_(vec[716]), .P2_INSTQUEUE_REG_2__2_(vec[715]), .P2_INSTQUEUE_REG_2__1_(vec[714]), .P2_INSTQUEUE_REG_2__0_(vec[713]), .P2_INSTQUEUE_REG_1__7_(vec[712]), .P2_INSTQUEUE_REG_1__6_(vec[711]), .P2_INSTQUEUE_REG_1__5_(vec[710]), .P2_INSTQUEUE_REG_1__4_(vec[709]), .P2_INSTQUEUE_REG_1__3_(vec[708]), .P2_INSTQUEUE_REG_1__2_(vec[707]), .P2_INSTQUEUE_REG_1__1_(vec[706]), .P2_INSTQUEUE_REG_1__0_(vec[705]), .P2_INSTQUEUE_REG_0__7_(vec[704]), .P2_INSTQUEUE_REG_0__6_(vec[703]), .P2_INSTQUEUE_REG_0__5_(vec[702]), .P2_INSTQUEUE_REG_0__4_(vec[701]), .P2_INSTQUEUE_REG_0__3_(vec[700]), .P2_INSTQUEUE_REG_0__2_(vec[699]), .P2_INSTQUEUE_REG_0__1_(vec[698]), .P2_INSTQUEUE_REG_0__0_(vec[697]), .P2_INSTQUEUERD_ADDR_REG_4_(vec[696]), .P2_INSTQUEUERD_ADDR_REG_3_(vec[695]), .P2_INSTQUEUERD_ADDR_REG_2_(vec[694]), .P2_INSTQUEUERD_ADDR_REG_1_(vec[693]), .P2_INSTQUEUERD_ADDR_REG_0_(vec[692]), .P2_INSTQUEUEWR_ADDR_REG_4_(vec[691]), .P2_INSTQUEUEWR_ADDR_REG_3_(vec[690]), .P2_INSTQUEUEWR_ADDR_REG_2_(vec[689]), .P2_INSTQUEUEWR_ADDR_REG_1_(vec[688]), .P2_INSTQUEUEWR_ADDR_REG_0_(vec[687]), .P2_INSTADDRPOINTER_REG_0_(vec[686]), .P2_INSTADDRPOINTER_REG_1_(vec[685]), .P2_INSTADDRPOINTER_REG_2_(vec[684]), .P2_INSTADDRPOINTER_REG_3_(vec[683]), .P2_INSTADDRPOINTER_REG_4_(vec[682]), .P2_INSTADDRPOINTER_REG_5_(vec[681]), .P2_INSTADDRPOINTER_REG_6_(vec[680]), .P2_INSTADDRPOINTER_REG_7_(vec[679]), .P2_INSTADDRPOINTER_REG_8_(vec[678]), .P2_INSTADDRPOINTER_REG_9_(vec[677]), .P2_INSTADDRPOINTER_REG_10_(vec[676]), .P2_INSTADDRPOINTER_REG_11_(vec[675]), .P2_INSTADDRPOINTER_REG_12_(vec[674]), .P2_INSTADDRPOINTER_REG_13_(vec[673]), .P2_INSTADDRPOINTER_REG_14_(vec[672]), .P2_INSTADDRPOINTER_REG_15_(vec[671]), .P2_INSTADDRPOINTER_REG_16_(vec[670]), .P2_INSTADDRPOINTER_REG_17_(vec[669]), .P2_INSTADDRPOINTER_REG_18_(vec[668]), .P2_INSTADDRPOINTER_REG_19_(vec[667]), .P2_INSTADDRPOINTER_REG_20_(vec[666]), .P2_INSTADDRPOINTER_REG_21_(vec[665]), .P2_INSTADDRPOINTER_REG_22_(vec[664]), .P2_INSTADDRPOINTER_REG_23_(vec[663]), .P2_INSTADDRPOINTER_REG_24_(vec[662]), .P2_INSTADDRPOINTER_REG_25_(vec[661]), .P2_INSTADDRPOINTER_REG_26_(vec[660]), .P2_INSTADDRPOINTER_REG_27_(vec[659]), .P2_INSTADDRPOINTER_REG_28_(vec[658]), .P2_INSTADDRPOINTER_REG_29_(vec[657]), .P2_INSTADDRPOINTER_REG_30_(vec[656]), .P2_INSTADDRPOINTER_REG_31_(vec[655]), .P2_PHYADDRPOINTER_REG_0_(vec[654]), .P2_PHYADDRPOINTER_REG_1_(vec[653]), .P2_PHYADDRPOINTER_REG_2_(vec[652]), .P2_PHYADDRPOINTER_REG_3_(vec[651]), .P2_PHYADDRPOINTER_REG_4_(vec[650]), .P2_PHYADDRPOINTER_REG_5_(vec[649]), .P2_PHYADDRPOINTER_REG_6_(vec[648]), .P2_PHYADDRPOINTER_REG_7_(vec[647]), .P2_PHYADDRPOINTER_REG_8_(vec[646]), .P2_PHYADDRPOINTER_REG_9_(vec[645]), .P2_PHYADDRPOINTER_REG_10_(vec[644]), .P2_PHYADDRPOINTER_REG_11_(vec[643]), .P2_PHYADDRPOINTER_REG_12_(vec[642]), .P2_PHYADDRPOINTER_REG_13_(vec[641]), .P2_PHYADDRPOINTER_REG_14_(vec[640]), .P2_PHYADDRPOINTER_REG_15_(vec[639]), .P2_PHYADDRPOINTER_REG_16_(vec[638]), .P2_PHYADDRPOINTER_REG_17_(vec[637]), .P2_PHYADDRPOINTER_REG_18_(vec[636]), .P2_PHYADDRPOINTER_REG_19_(vec[635]), .P2_PHYADDRPOINTER_REG_20_(vec[634]), .P2_PHYADDRPOINTER_REG_21_(vec[633]), .P2_PHYADDRPOINTER_REG_22_(vec[632]), .P2_PHYADDRPOINTER_REG_23_(vec[631]), .P2_PHYADDRPOINTER_REG_24_(vec[630]), .P2_PHYADDRPOINTER_REG_25_(vec[629]), .P2_PHYADDRPOINTER_REG_26_(vec[628]), .P2_PHYADDRPOINTER_REG_27_(vec[627]), .P2_PHYADDRPOINTER_REG_28_(vec[626]), .P2_PHYADDRPOINTER_REG_29_(vec[625]), .P2_PHYADDRPOINTER_REG_30_(vec[624]), .P2_PHYADDRPOINTER_REG_31_(vec[623]), .P2_LWORD_REG_15_(vec[622]), .P2_LWORD_REG_14_(vec[621]), .P2_LWORD_REG_13_(vec[620]), .P2_LWORD_REG_12_(vec[619]), .P2_LWORD_REG_11_(vec[618]), .P2_LWORD_REG_10_(vec[617]), .P2_LWORD_REG_9_(vec[616]), .P2_LWORD_REG_8_(vec[615]), .P2_LWORD_REG_7_(vec[614]), .P2_LWORD_REG_6_(vec[613]), .P2_LWORD_REG_5_(vec[612]), .P2_LWORD_REG_4_(vec[611]), .P2_LWORD_REG_3_(vec[610]), .P2_LWORD_REG_2_(vec[609]), .P2_LWORD_REG_1_(vec[608]), .P2_LWORD_REG_0_(vec[607]), .P2_UWORD_REG_14_(vec[606]), .P2_UWORD_REG_13_(vec[605]), .P2_UWORD_REG_12_(vec[604]), .P2_UWORD_REG_11_(vec[603]), .P2_UWORD_REG_10_(vec[602]), .P2_UWORD_REG_9_(vec[601]), .P2_UWORD_REG_8_(vec[600]), .P2_UWORD_REG_7_(vec[599]), .P2_UWORD_REG_6_(vec[598]), .P2_UWORD_REG_5_(vec[597]), .P2_UWORD_REG_4_(vec[596]), .P2_UWORD_REG_3_(vec[595]), .P2_UWORD_REG_2_(vec[594]), .P2_UWORD_REG_1_(vec[593]), .P2_UWORD_REG_0_(vec[592]), .P2_DATAO_REG_0_(vec[591]), .P2_DATAO_REG_1_(vec[590]), .P2_DATAO_REG_2_(vec[589]), .P2_DATAO_REG_3_(vec[588]), .P2_DATAO_REG_4_(vec[587]), .P2_DATAO_REG_5_(vec[586]), .P2_DATAO_REG_6_(vec[585]), .P2_DATAO_REG_7_(vec[584]), .P2_DATAO_REG_8_(vec[583]), .P2_DATAO_REG_9_(vec[582]), .P2_DATAO_REG_10_(vec[581]), .P2_DATAO_REG_11_(vec[580]), .P2_DATAO_REG_12_(vec[579]), .P2_DATAO_REG_13_(vec[578]), .P2_DATAO_REG_14_(vec[577]), .P2_DATAO_REG_15_(vec[576]), .P2_DATAO_REG_16_(vec[575]), .P2_DATAO_REG_17_(vec[574]), .P2_DATAO_REG_18_(vec[573]), .P2_DATAO_REG_19_(vec[572]), .P2_DATAO_REG_20_(vec[571]), .P2_DATAO_REG_21_(vec[570]), .P2_DATAO_REG_22_(vec[569]), .P2_DATAO_REG_23_(vec[568]), .P2_DATAO_REG_24_(vec[567]), .P2_DATAO_REG_25_(vec[566]), .P2_DATAO_REG_26_(vec[565]), .P2_DATAO_REG_27_(vec[564]), .P2_DATAO_REG_28_(vec[563]), .P2_DATAO_REG_29_(vec[562]), .P2_DATAO_REG_30_(vec[561]), .P2_DATAO_REG_31_(vec[560]), .P2_EAX_REG_0_(vec[559]), .P2_EAX_REG_1_(vec[558]), .P2_EAX_REG_2_(vec[557]), .P2_EAX_REG_3_(vec[556]), .P2_EAX_REG_4_(vec[555]), .P2_EAX_REG_5_(vec[554]), .P2_EAX_REG_6_(vec[553]), .P2_EAX_REG_7_(vec[552]), .P2_EAX_REG_8_(vec[551]), .P2_EAX_REG_9_(vec[550]), .P2_EAX_REG_10_(vec[549]), .P2_EAX_REG_11_(vec[548]), .P2_EAX_REG_12_(vec[547]), .P2_EAX_REG_13_(vec[546]), .P2_EAX_REG_14_(vec[545]), .P2_EAX_REG_15_(vec[544]), .P2_EAX_REG_16_(vec[543]), .P2_EAX_REG_17_(vec[542]), .P2_EAX_REG_18_(vec[541]), .P2_EAX_REG_19_(vec[540]), .P2_EAX_REG_20_(vec[539]), .P2_EAX_REG_21_(vec[538]), .P2_EAX_REG_22_(vec[537]), .P2_EAX_REG_23_(vec[536]), .P2_EAX_REG_24_(vec[535]), .P2_EAX_REG_25_(vec[534]), .P2_EAX_REG_26_(vec[533]), .P2_EAX_REG_27_(vec[532]), .P2_EAX_REG_28_(vec[531]), .P2_EAX_REG_29_(vec[530]), .P2_EAX_REG_30_(vec[529]), .P2_EAX_REG_31_(vec[528]), .P2_EBX_REG_0_(vec[527]), .P2_EBX_REG_1_(vec[526]), .P2_EBX_REG_2_(vec[525]), .P2_EBX_REG_3_(vec[524]), .P2_EBX_REG_4_(vec[523]), .P2_EBX_REG_5_(vec[522]), .P2_EBX_REG_6_(vec[521]), .P2_EBX_REG_7_(vec[520]), .P2_EBX_REG_8_(vec[519]), .P2_EBX_REG_9_(vec[518]), .P2_EBX_REG_10_(vec[517]), .P2_EBX_REG_11_(vec[516]), .P2_EBX_REG_12_(vec[515]), .P2_EBX_REG_13_(vec[514]), .P2_EBX_REG_14_(vec[513]), .P2_EBX_REG_15_(vec[512]), .P2_EBX_REG_16_(vec[511]), .P2_EBX_REG_17_(vec[510]), .P2_EBX_REG_18_(vec[509]), .P2_EBX_REG_19_(vec[508]), .P2_EBX_REG_20_(vec[507]), .P2_EBX_REG_21_(vec[506]), .P2_EBX_REG_22_(vec[505]), .P2_EBX_REG_23_(vec[504]), .P2_EBX_REG_24_(vec[503]), .P2_EBX_REG_25_(vec[502]), .P2_EBX_REG_26_(vec[501]), .P2_EBX_REG_27_(vec[500]), .P2_EBX_REG_28_(vec[499]), .P2_EBX_REG_29_(vec[498]), .P2_EBX_REG_30_(vec[497]), .P2_EBX_REG_31_(vec[496]), .P2_REIP_REG_0_(vec[495]), .P2_REIP_REG_1_(vec[494]), .P2_REIP_REG_2_(vec[493]), .P2_REIP_REG_3_(vec[492]), .P2_REIP_REG_4_(vec[491]), .P2_REIP_REG_5_(vec[490]), .P2_REIP_REG_6_(vec[489]), .P2_REIP_REG_7_(vec[488]), .P2_REIP_REG_8_(vec[487]), .P2_REIP_REG_9_(vec[486]), .P2_REIP_REG_10_(vec[485]), .P2_REIP_REG_11_(vec[484]), .P2_REIP_REG_12_(vec[483]), .P2_REIP_REG_13_(vec[482]), .P2_REIP_REG_14_(vec[481]), .P2_REIP_REG_15_(vec[480]), .P2_REIP_REG_16_(vec[479]), .P2_REIP_REG_17_(vec[478]), .P2_REIP_REG_18_(vec[477]), .P2_REIP_REG_19_(vec[476]), .P2_REIP_REG_20_(vec[475]), .P2_REIP_REG_21_(vec[474]), .P2_REIP_REG_22_(vec[473]), .P2_REIP_REG_23_(vec[472]), .P2_REIP_REG_24_(vec[471]), .P2_REIP_REG_25_(vec[470]), .P2_REIP_REG_26_(vec[469]), .P2_REIP_REG_27_(vec[468]), .P2_REIP_REG_28_(vec[467]), .P2_REIP_REG_29_(vec[466]), .P2_REIP_REG_30_(vec[465]), .P2_REIP_REG_31_(vec[464]), .P2_BYTEENABLE_REG_3_(vec[463]), .P2_BYTEENABLE_REG_2_(vec[462]), .P2_BYTEENABLE_REG_1_(vec[461]), .P2_BYTEENABLE_REG_0_(vec[460]), .P2_W_R_N_REG(vec[459]), .P2_FLUSH_REG(vec[458]), .P2_MORE_REG(vec[457]), .P2_STATEBS16_REG(vec[456]), .P2_REQUESTPENDING_REG(vec[455]), .P2_D_C_N_REG(vec[454]), .P2_M_IO_N_REG(vec[453]), .P2_CODEFETCH_REG(vec[452]), .P2_ADS_N_REG(vec[451]), .P2_READREQUEST_REG(vec[450]), .P2_MEMORYFETCH_REG(vec[449]), .P1_BE_N_REG_3_(vec[448]), .P1_BE_N_REG_2_(vec[447]), .P1_BE_N_REG_1_(vec[446]), .P1_BE_N_REG_0_(vec[445]), .P1_ADDRESS_REG_29__EXTRA(vec[444]), .P1_ADDRESS_REG_28__EXTRA(vec[443]), .P1_ADDRESS_REG_27__EXTRA(vec[442]), .P1_ADDRESS_REG_26__EXTRA(vec[441]), .P1_ADDRESS_REG_25__EXTRA(vec[440]), .P1_ADDRESS_REG_24__EXTRA(vec[439]), .P1_ADDRESS_REG_23__EXTRA(vec[438]), .P1_ADDRESS_REG_22__EXTRA(vec[437]), .P1_ADDRESS_REG_21__EXTRA(vec[436]), .P1_ADDRESS_REG_20__EXTRA(vec[435]), .P1_ADDRESS_REG_19__EXTRA(vec[434]), .P1_ADDRESS_REG_18__EXTRA(vec[433]), .P1_ADDRESS_REG_17__EXTRA(vec[432]), .P1_ADDRESS_REG_16__EXTRA(vec[431]), .P1_ADDRESS_REG_15__EXTRA(vec[430]), .P1_ADDRESS_REG_14__EXTRA(vec[429]), .P1_ADDRESS_REG_13__EXTRA(vec[428]), .P1_ADDRESS_REG_12__EXTRA(vec[427]), .P1_ADDRESS_REG_11__EXTRA(vec[426]), .P1_ADDRESS_REG_10__EXTRA(vec[425]), .P1_ADDRESS_REG_9__EXTRA(vec[424]), .P1_ADDRESS_REG_8__EXTRA(vec[423]), .P1_ADDRESS_REG_7__EXTRA(vec[422]), .P1_ADDRESS_REG_6__EXTRA(vec[421]), .P1_ADDRESS_REG_5__EXTRA(vec[420]), .P1_ADDRESS_REG_4__EXTRA(vec[419]), .P1_ADDRESS_REG_3__EXTRA(vec[418]), .P1_ADDRESS_REG_2__EXTRA(vec[417]), .P1_ADDRESS_REG_1__EXTRA(vec[416]), .P1_ADDRESS_REG_0__EXTRA(vec[415]), .P1_STATE_REG_2_(vec[414]), .P1_STATE_REG_1_(vec[413]), .P1_STATE_REG_0_(vec[412]), .P1_DATAWIDTH_REG_0_(vec[411]), .P1_DATAWIDTH_REG_1_(vec[410]), .P1_DATAWIDTH_REG_2_(vec[409]), .P1_DATAWIDTH_REG_3_(vec[408]), .P1_DATAWIDTH_REG_4_(vec[407]), .P1_DATAWIDTH_REG_5_(vec[406]), .P1_DATAWIDTH_REG_6_(vec[405]), .P1_DATAWIDTH_REG_7_(vec[404]), .P1_DATAWIDTH_REG_8_(vec[403]), .P1_DATAWIDTH_REG_9_(vec[402]), .P1_DATAWIDTH_REG_10_(vec[401]), .P1_DATAWIDTH_REG_11_(vec[400]), .P1_DATAWIDTH_REG_12_(vec[399]), .P1_DATAWIDTH_REG_13_(vec[398]), .P1_DATAWIDTH_REG_14_(vec[397]), .P1_DATAWIDTH_REG_15_(vec[396]), .P1_DATAWIDTH_REG_16_(vec[395]), .P1_DATAWIDTH_REG_17_(vec[394]), .P1_DATAWIDTH_REG_18_(vec[393]), .P1_DATAWIDTH_REG_19_(vec[392]), .P1_DATAWIDTH_REG_20_(vec[391]), .P1_DATAWIDTH_REG_21_(vec[390]), .P1_DATAWIDTH_REG_22_(vec[389]), .P1_DATAWIDTH_REG_23_(vec[388]), .P1_DATAWIDTH_REG_24_(vec[387]), .P1_DATAWIDTH_REG_25_(vec[386]), .P1_DATAWIDTH_REG_26_(vec[385]), .P1_DATAWIDTH_REG_27_(vec[384]), .P1_DATAWIDTH_REG_28_(vec[383]), .P1_DATAWIDTH_REG_29_(vec[382]), .P1_DATAWIDTH_REG_30_(vec[381]), .P1_DATAWIDTH_REG_31_(vec[380]), .P1_STATE2_REG_3_(vec[379]), .P1_STATE2_REG_2_(vec[378]), .P1_STATE2_REG_1_(vec[377]), .P1_STATE2_REG_0_(vec[376]), .P1_INSTQUEUE_REG_15__7_(vec[375]), .P1_INSTQUEUE_REG_15__6_(vec[374]), .P1_INSTQUEUE_REG_15__5_(vec[373]), .P1_INSTQUEUE_REG_15__4_(vec[372]), .P1_INSTQUEUE_REG_15__3_(vec[371]), .P1_INSTQUEUE_REG_15__2_(vec[370]), .P1_INSTQUEUE_REG_15__1_(vec[369]), .P1_INSTQUEUE_REG_15__0_(vec[368]), .P1_INSTQUEUE_REG_14__7_(vec[367]), .P1_INSTQUEUE_REG_14__6_(vec[366]), .P1_INSTQUEUE_REG_14__5_(vec[365]), .P1_INSTQUEUE_REG_14__4_(vec[364]), .P1_INSTQUEUE_REG_14__3_(vec[363]), .P1_INSTQUEUE_REG_14__2_(vec[362]), .P1_INSTQUEUE_REG_14__1_(vec[361]), .P1_INSTQUEUE_REG_14__0_(vec[360]), .P1_INSTQUEUE_REG_13__7_(vec[359]), .P1_INSTQUEUE_REG_13__6_(vec[358]), .P1_INSTQUEUE_REG_13__5_(vec[357]), .P1_INSTQUEUE_REG_13__4_(vec[356]), .P1_INSTQUEUE_REG_13__3_(vec[355]), .P1_INSTQUEUE_REG_13__2_(vec[354]), .P1_INSTQUEUE_REG_13__1_(vec[353]), .P1_INSTQUEUE_REG_13__0_(vec[352]), .P1_INSTQUEUE_REG_12__7_(vec[351]), .P1_INSTQUEUE_REG_12__6_(vec[350]), .P1_INSTQUEUE_REG_12__5_(vec[349]), .P1_INSTQUEUE_REG_12__4_(vec[348]), .P1_INSTQUEUE_REG_12__3_(vec[347]), .P1_INSTQUEUE_REG_12__2_(vec[346]), .P1_INSTQUEUE_REG_12__1_(vec[345]), .P1_INSTQUEUE_REG_12__0_(vec[344]), .P1_INSTQUEUE_REG_11__7_(vec[343]), .P1_INSTQUEUE_REG_11__6_(vec[342]), .P1_INSTQUEUE_REG_11__5_(vec[341]), .P1_INSTQUEUE_REG_11__4_(vec[340]), .P1_INSTQUEUE_REG_11__3_(vec[339]), .P1_INSTQUEUE_REG_11__2_(vec[338]), .P1_INSTQUEUE_REG_11__1_(vec[337]), .P1_INSTQUEUE_REG_11__0_(vec[336]), .P1_INSTQUEUE_REG_10__7_(vec[335]), .P1_INSTQUEUE_REG_10__6_(vec[334]), .P1_INSTQUEUE_REG_10__5_(vec[333]), .P1_INSTQUEUE_REG_10__4_(vec[332]), .P1_INSTQUEUE_REG_10__3_(vec[331]), .P1_INSTQUEUE_REG_10__2_(vec[330]), .P1_INSTQUEUE_REG_10__1_(vec[329]), .P1_INSTQUEUE_REG_10__0_(vec[328]), .P1_INSTQUEUE_REG_9__7_(vec[327]), .P1_INSTQUEUE_REG_9__6_(vec[326]), .P1_INSTQUEUE_REG_9__5_(vec[325]), .P1_INSTQUEUE_REG_9__4_(vec[324]), .P1_INSTQUEUE_REG_9__3_(vec[323]), .P1_INSTQUEUE_REG_9__2_(vec[322]), .P1_INSTQUEUE_REG_9__1_(vec[321]), .P1_INSTQUEUE_REG_9__0_(vec[320]), .P1_INSTQUEUE_REG_8__7_(vec[319]), .P1_INSTQUEUE_REG_8__6_(vec[318]), .P1_INSTQUEUE_REG_8__5_(vec[317]), .P1_INSTQUEUE_REG_8__4_(vec[316]), .P1_INSTQUEUE_REG_8__3_(vec[315]), .P1_INSTQUEUE_REG_8__2_(vec[314]), .P1_INSTQUEUE_REG_8__1_(vec[313]), .P1_INSTQUEUE_REG_8__0_(vec[312]), .P1_INSTQUEUE_REG_7__7_(vec[311]), .P1_INSTQUEUE_REG_7__6_(vec[310]), .P1_INSTQUEUE_REG_7__5_(vec[309]), .P1_INSTQUEUE_REG_7__4_(vec[308]), .P1_INSTQUEUE_REG_7__3_(vec[307]), .P1_INSTQUEUE_REG_7__2_(vec[306]), .P1_INSTQUEUE_REG_7__1_(vec[305]), .P1_INSTQUEUE_REG_7__0_(vec[304]), .P1_INSTQUEUE_REG_6__7_(vec[303]), .P1_INSTQUEUE_REG_6__6_(vec[302]), .P1_INSTQUEUE_REG_6__5_(vec[301]), .P1_INSTQUEUE_REG_6__4_(vec[300]), .P1_INSTQUEUE_REG_6__3_(vec[299]), .P1_INSTQUEUE_REG_6__2_(vec[298]), .P1_INSTQUEUE_REG_6__1_(vec[297]), .P1_INSTQUEUE_REG_6__0_(vec[296]), .P1_INSTQUEUE_REG_5__7_(vec[295]), .P1_INSTQUEUE_REG_5__6_(vec[294]), .P1_INSTQUEUE_REG_5__5_(vec[293]), .P1_INSTQUEUE_REG_5__4_(vec[292]), .P1_INSTQUEUE_REG_5__3_(vec[291]), .P1_INSTQUEUE_REG_5__2_(vec[290]), .P1_INSTQUEUE_REG_5__1_(vec[289]), .P1_INSTQUEUE_REG_5__0_(vec[288]), .P1_INSTQUEUE_REG_4__7_(vec[287]), .P1_INSTQUEUE_REG_4__6_(vec[286]), .P1_INSTQUEUE_REG_4__5_(vec[285]), .P1_INSTQUEUE_REG_4__4_(vec[284]), .P1_INSTQUEUE_REG_4__3_(vec[283]), .P1_INSTQUEUE_REG_4__2_(vec[282]), .P1_INSTQUEUE_REG_4__1_(vec[281]), .P1_INSTQUEUE_REG_4__0_(vec[280]), .P1_INSTQUEUE_REG_3__7_(vec[279]), .P1_INSTQUEUE_REG_3__6_(vec[278]), .P1_INSTQUEUE_REG_3__5_(vec[277]), .P1_INSTQUEUE_REG_3__4_(vec[276]), .P1_INSTQUEUE_REG_3__3_(vec[275]), .P1_INSTQUEUE_REG_3__2_(vec[274]), .P1_INSTQUEUE_REG_3__1_(vec[273]), .P1_INSTQUEUE_REG_3__0_(vec[272]), .P1_INSTQUEUE_REG_2__7_(vec[271]), .P1_INSTQUEUE_REG_2__6_(vec[270]), .P1_INSTQUEUE_REG_2__5_(vec[269]), .P1_INSTQUEUE_REG_2__4_(vec[268]), .P1_INSTQUEUE_REG_2__3_(vec[267]), .P1_INSTQUEUE_REG_2__2_(vec[266]), .P1_INSTQUEUE_REG_2__1_(vec[265]), .P1_INSTQUEUE_REG_2__0_(vec[264]), .P1_INSTQUEUE_REG_1__7_(vec[263]), .P1_INSTQUEUE_REG_1__6_(vec[262]), .P1_INSTQUEUE_REG_1__5_(vec[261]), .P1_INSTQUEUE_REG_1__4_(vec[260]), .P1_INSTQUEUE_REG_1__3_(vec[259]), .P1_INSTQUEUE_REG_1__2_(vec[258]), .P1_INSTQUEUE_REG_1__1_(vec[257]), .P1_INSTQUEUE_REG_1__0_(vec[256]), .P1_INSTQUEUE_REG_0__7_(vec[255]), .P1_INSTQUEUE_REG_0__6_(vec[254]), .P1_INSTQUEUE_REG_0__5_(vec[253]), .P1_INSTQUEUE_REG_0__4_(vec[252]), .P1_INSTQUEUE_REG_0__3_(vec[251]), .P1_INSTQUEUE_REG_0__2_(vec[250]), .P1_INSTQUEUE_REG_0__1_(vec[249]), .P1_INSTQUEUE_REG_0__0_(vec[248]), .P1_INSTQUEUERD_ADDR_REG_4_(vec[247]), .P1_INSTQUEUERD_ADDR_REG_3_(vec[246]), .P1_INSTQUEUERD_ADDR_REG_2_(vec[245]), .P1_INSTQUEUERD_ADDR_REG_1_(vec[244]), .P1_INSTQUEUERD_ADDR_REG_0_(vec[243]), .P1_INSTQUEUEWR_ADDR_REG_4_(vec[242]), .P1_INSTQUEUEWR_ADDR_REG_3_(vec[241]), .P1_INSTQUEUEWR_ADDR_REG_2_(vec[240]), .P1_INSTQUEUEWR_ADDR_REG_1_(vec[239]), .P1_INSTQUEUEWR_ADDR_REG_0_(vec[238]), .P1_INSTADDRPOINTER_REG_0_(vec[237]), .P1_INSTADDRPOINTER_REG_1_(vec[236]), .P1_INSTADDRPOINTER_REG_2_(vec[235]), .P1_INSTADDRPOINTER_REG_3_(vec[234]), .P1_INSTADDRPOINTER_REG_4_(vec[233]), .P1_INSTADDRPOINTER_REG_5_(vec[232]), .P1_INSTADDRPOINTER_REG_6_(vec[231]), .P1_INSTADDRPOINTER_REG_7_(vec[230]), .P1_INSTADDRPOINTER_REG_8_(vec[229]), .P1_INSTADDRPOINTER_REG_9_(vec[228]), .P1_INSTADDRPOINTER_REG_10_(vec[227]), .P1_INSTADDRPOINTER_REG_11_(vec[226]), .P1_INSTADDRPOINTER_REG_12_(vec[225]), .P1_INSTADDRPOINTER_REG_13_(vec[224]), .P1_INSTADDRPOINTER_REG_14_(vec[223]), .P1_INSTADDRPOINTER_REG_15_(vec[222]), .P1_INSTADDRPOINTER_REG_16_(vec[221]), .P1_INSTADDRPOINTER_REG_17_(vec[220]), .P1_INSTADDRPOINTER_REG_18_(vec[219]), .P1_INSTADDRPOINTER_REG_19_(vec[218]), .P1_INSTADDRPOINTER_REG_20_(vec[217]), .P1_INSTADDRPOINTER_REG_21_(vec[216]), .P1_INSTADDRPOINTER_REG_22_(vec[215]), .P1_INSTADDRPOINTER_REG_23_(vec[214]), .P1_INSTADDRPOINTER_REG_24_(vec[213]), .P1_INSTADDRPOINTER_REG_25_(vec[212]), .P1_INSTADDRPOINTER_REG_26_(vec[211]), .P1_INSTADDRPOINTER_REG_27_(vec[210]), .P1_INSTADDRPOINTER_REG_28_(vec[209]), .P1_INSTADDRPOINTER_REG_29_(vec[208]), .P1_INSTADDRPOINTER_REG_30_(vec[207]), .P1_INSTADDRPOINTER_REG_31_(vec[206]), .P1_PHYADDRPOINTER_REG_0_(vec[205]), .P1_PHYADDRPOINTER_REG_1_(vec[204]), .P1_PHYADDRPOINTER_REG_2_(vec[203]), .P1_PHYADDRPOINTER_REG_3_(vec[202]), .P1_PHYADDRPOINTER_REG_4_(vec[201]), .P1_PHYADDRPOINTER_REG_5_(vec[200]), .P1_PHYADDRPOINTER_REG_6_(vec[199]), .P1_PHYADDRPOINTER_REG_7_(vec[198]), .P1_PHYADDRPOINTER_REG_8_(vec[197]), .P1_PHYADDRPOINTER_REG_9_(vec[196]), .P1_PHYADDRPOINTER_REG_10_(vec[195]), .P1_PHYADDRPOINTER_REG_11_(vec[194]), .P1_PHYADDRPOINTER_REG_12_(vec[193]), .P1_PHYADDRPOINTER_REG_13_(vec[192]), .P1_PHYADDRPOINTER_REG_14_(vec[191]), .P1_PHYADDRPOINTER_REG_15_(vec[190]), .P1_PHYADDRPOINTER_REG_16_(vec[189]), .P1_PHYADDRPOINTER_REG_17_(vec[188]), .P1_PHYADDRPOINTER_REG_18_(vec[187]), .P1_PHYADDRPOINTER_REG_19_(vec[186]), .P1_PHYADDRPOINTER_REG_20_(vec[185]), .P1_PHYADDRPOINTER_REG_21_(vec[184]), .P1_PHYADDRPOINTER_REG_22_(vec[183]), .P1_PHYADDRPOINTER_REG_23_(vec[182]), .P1_PHYADDRPOINTER_REG_24_(vec[181]), .P1_PHYADDRPOINTER_REG_25_(vec[180]), .P1_PHYADDRPOINTER_REG_26_(vec[179]), .P1_PHYADDRPOINTER_REG_27_(vec[178]), .P1_PHYADDRPOINTER_REG_28_(vec[177]), .P1_PHYADDRPOINTER_REG_29_(vec[176]), .P1_PHYADDRPOINTER_REG_30_(vec[175]), .P1_PHYADDRPOINTER_REG_31_(vec[174]), .P1_LWORD_REG_15_(vec[173]), .P1_LWORD_REG_14_(vec[172]), .P1_LWORD_REG_13_(vec[171]), .P1_LWORD_REG_12_(vec[170]), .P1_LWORD_REG_11_(vec[169]), .P1_LWORD_REG_10_(vec[168]), .P1_LWORD_REG_9_(vec[167]), .P1_LWORD_REG_8_(vec[166]), .P1_LWORD_REG_7_(vec[165]), .P1_LWORD_REG_6_(vec[164]), .P1_LWORD_REG_5_(vec[163]), .P1_LWORD_REG_4_(vec[162]), .P1_LWORD_REG_3_(vec[161]), .P1_LWORD_REG_2_(vec[160]), .P1_LWORD_REG_1_(vec[159]), .P1_LWORD_REG_0_(vec[158]), .P1_UWORD_REG_14_(vec[157]), .P1_UWORD_REG_13_(vec[156]), .P1_UWORD_REG_12_(vec[155]), .P1_UWORD_REG_11_(vec[154]), .P1_UWORD_REG_10_(vec[153]), .P1_UWORD_REG_9_(vec[152]), .P1_UWORD_REG_8_(vec[151]), .P1_UWORD_REG_7_(vec[150]), .P1_UWORD_REG_6_(vec[149]), .P1_UWORD_REG_5_(vec[148]), .P1_UWORD_REG_4_(vec[147]), .P1_UWORD_REG_3_(vec[146]), .P1_UWORD_REG_2_(vec[145]), .P1_UWORD_REG_1_(vec[144]), .P1_UWORD_REG_0_(vec[143]), .P1_DATAO_REG_0_(vec[142]), .P1_DATAO_REG_1_(vec[141]), .P1_DATAO_REG_2_(vec[140]), .P1_DATAO_REG_3_(vec[139]), .P1_DATAO_REG_4_(vec[138]), .P1_DATAO_REG_5_(vec[137]), .P1_DATAO_REG_6_(vec[136]), .P1_DATAO_REG_7_(vec[135]), .P1_DATAO_REG_8_(vec[134]), .P1_DATAO_REG_9_(vec[133]), .P1_DATAO_REG_10_(vec[132]), .P1_DATAO_REG_11_(vec[131]), .P1_DATAO_REG_12_(vec[130]), .P1_DATAO_REG_13_(vec[129]), .P1_DATAO_REG_14_(vec[128]), .P1_DATAO_REG_15_(vec[127]), .P1_DATAO_REG_16_(vec[126]), .P1_DATAO_REG_17_(vec[125]), .P1_DATAO_REG_18_(vec[124]), .P1_DATAO_REG_19_(vec[123]), .P1_DATAO_REG_20_(vec[122]), .P1_DATAO_REG_21_(vec[121]), .P1_DATAO_REG_22_(vec[120]), .P1_DATAO_REG_23_(vec[119]), .P1_DATAO_REG_24_(vec[118]), .P1_DATAO_REG_25_(vec[117]), .P1_DATAO_REG_26_(vec[116]), .P1_DATAO_REG_27_(vec[115]), .P1_DATAO_REG_28_(vec[114]), .P1_DATAO_REG_29_(vec[113]), .P1_DATAO_REG_30_(vec[112]), .P1_DATAO_REG_31_(vec[111]), .P1_EAX_REG_0_(vec[110]), .P1_EAX_REG_1_(vec[109]), .P1_EAX_REG_2_(vec[108]), .P1_EAX_REG_3_(vec[107]), .P1_EAX_REG_4_(vec[106]), .P1_EAX_REG_5_(vec[105]), .P1_EAX_REG_6_(vec[104]), .P1_EAX_REG_7_(vec[103]), .P1_EAX_REG_8_(vec[102]), .P1_EAX_REG_9_(vec[101]), .P1_EAX_REG_10_(vec[100]), .P1_EAX_REG_11_(vec[99]), .P1_EAX_REG_12_(vec[98]), .P1_EAX_REG_13_(vec[97]), .P1_EAX_REG_14_(vec[96]), .P1_EAX_REG_15_(vec[95]), .P1_EAX_REG_16_(vec[94]), .P1_EAX_REG_17_(vec[93]), .P1_EAX_REG_18_(vec[92]), .P1_EAX_REG_19_(vec[91]), .P1_EAX_REG_20_(vec[90]), .P1_EAX_REG_21_(vec[89]), .P1_EAX_REG_22_(vec[88]), .P1_EAX_REG_23_(vec[87]), .P1_EAX_REG_24_(vec[86]), .P1_EAX_REG_25_(vec[85]), .P1_EAX_REG_26_(vec[84]), .P1_EAX_REG_27_(vec[83]), .P1_EAX_REG_28_(vec[82]), .P1_EAX_REG_29_(vec[81]), .P1_EAX_REG_30_(vec[80]), .P1_EAX_REG_31_(vec[79]), .P1_EBX_REG_0_(vec[78]), .P1_EBX_REG_1_(vec[77]), .P1_EBX_REG_2_(vec[76]), .P1_EBX_REG_3_(vec[75]), .P1_EBX_REG_4_(vec[74]), .P1_EBX_REG_5_(vec[73]), .P1_EBX_REG_6_(vec[72]), .P1_EBX_REG_7_(vec[71]), .P1_EBX_REG_8_(vec[70]), .P1_EBX_REG_9_(vec[69]), .P1_EBX_REG_10_(vec[68]), .P1_EBX_REG_11_(vec[67]), .P1_EBX_REG_12_(vec[66]), .P1_EBX_REG_13_(vec[65]), .P1_EBX_REG_14_(vec[64]), .P1_EBX_REG_15_(vec[63]), .P1_EBX_REG_16_(vec[62]), .P1_EBX_REG_17_(vec[61]), .P1_EBX_REG_18_(vec[60]), .P1_EBX_REG_19_(vec[59]), .P1_EBX_REG_20_(vec[58]), .P1_EBX_REG_21_(vec[57]), .P1_EBX_REG_22_(vec[56]), .P1_EBX_REG_23_(vec[55]), .P1_EBX_REG_24_(vec[54]), .P1_EBX_REG_25_(vec[53]), .P1_EBX_REG_26_(vec[52]), .P1_EBX_REG_27_(vec[51]), .P1_EBX_REG_28_(vec[50]), .P1_EBX_REG_29_(vec[49]), .P1_EBX_REG_30_(vec[48]), .P1_EBX_REG_31_(vec[47]), .P1_REIP_REG_0_(vec[46]), .P1_REIP_REG_1_(vec[45]), .P1_REIP_REG_2_(vec[44]), .P1_REIP_REG_3_(vec[43]), .P1_REIP_REG_4_(vec[42]), .P1_REIP_REG_5_(vec[41]), .P1_REIP_REG_6_(vec[40]), .P1_REIP_REG_7_(vec[39]), .P1_REIP_REG_8_(vec[38]), .P1_REIP_REG_9_(vec[37]), .P1_REIP_REG_10_(vec[36]), .P1_REIP_REG_11_(vec[35]), .P1_REIP_REG_12_(vec[34]), .P1_REIP_REG_13_(vec[33]), .P1_REIP_REG_14_(vec[32]), .P1_REIP_REG_15_(vec[31]), .P1_REIP_REG_16_(vec[30]), .P1_REIP_REG_17_(vec[29]), .P1_REIP_REG_18_(vec[28]), .P1_REIP_REG_19_(vec[27]), .P1_REIP_REG_20_(vec[26]), .P1_REIP_REG_21_(vec[25]), .P1_REIP_REG_22_(vec[24]), .P1_REIP_REG_23_(vec[23]), .P1_REIP_REG_24_(vec[22]), .P1_REIP_REG_25_(vec[21]), .P1_REIP_REG_26_(vec[20]), .P1_REIP_REG_27_(vec[19]), .P1_REIP_REG_28_(vec[18]), .P1_REIP_REG_29_(vec[17]), .P1_REIP_REG_30_(vec[16]), .P1_REIP_REG_31_(vec[15]), .P1_BYTEENABLE_REG_3_(vec[14]), .P1_BYTEENABLE_REG_2_(vec[13]), .P1_BYTEENABLE_REG_1_(vec[12]), .P1_BYTEENABLE_REG_0_(vec[11]), .P1_W_R_N_REG(vec[10]), .P1_FLUSH_REG(vec[9]), .P1_MORE_REG(vec[8]), .P1_STATEBS16_REG(vec[7]), .P1_REQUESTPENDING_REG(vec[6]), .P1_D_C_N_REG(vec[5]), .P1_M_IO_N_REG(vec[4]), .P1_CODEFETCH_REG(vec[3]), .P1_ADS_N_REG_EXTRA(vec[2]), .P1_READREQUEST_REG(vec[1]), .P1_MEMORYFETCH_REG(vec[0]), .P3_DATAO_REG_31_(p3_datao_reg_31_), .P3_DATAO_REG_30_(p3_datao_reg_30_), .P3_DATAO_REG_29_(p3_datao_reg_29_), .P3_DATAO_REG_28_(p3_datao_reg_28_), .P3_DATAO_REG_27_(p3_datao_reg_27_), .P3_DATAO_REG_26_(p3_datao_reg_26_), .P3_DATAO_REG_25_(p3_datao_reg_25_), .P3_DATAO_REG_24_(p3_datao_reg_24_), .P3_DATAO_REG_23_(p3_datao_reg_23_), .P3_DATAO_REG_22_(p3_datao_reg_22_), .P3_DATAO_REG_21_(p3_datao_reg_21_), .P3_DATAO_REG_20_(p3_datao_reg_20_), .P3_DATAO_REG_19_(p3_datao_reg_19_), .P3_DATAO_REG_18_(p3_datao_reg_18_), .P3_DATAO_REG_17_(p3_datao_reg_17_), .P3_DATAO_REG_16_(p3_datao_reg_16_), .P3_DATAO_REG_15_(p3_datao_reg_15_), .P3_DATAO_REG_14_(p3_datao_reg_14_), .P3_DATAO_REG_13_(p3_datao_reg_13_), .P3_DATAO_REG_12_(p3_datao_reg_12_), .P3_DATAO_REG_11_(p3_datao_reg_11_), .P3_DATAO_REG_10_(p3_datao_reg_10_), .P3_DATAO_REG_9_(p3_datao_reg_9_), .P3_DATAO_REG_8_(p3_datao_reg_8_), .P3_DATAO_REG_7_(p3_datao_reg_7_), .P3_DATAO_REG_6_(p3_datao_reg_6_), .P3_DATAO_REG_5_(p3_datao_reg_5_), .P3_DATAO_REG_4_(p3_datao_reg_4_), .P3_DATAO_REG_3_(p3_datao_reg_3_), .P3_DATAO_REG_2_(p3_datao_reg_2_), .P3_DATAO_REG_1_(p3_datao_reg_1_), .P3_DATAO_REG_0_(p3_datao_reg_0_), .P1_ADDRESS_REG_29_(p1_address_reg_29_), .P1_ADDRESS_REG_28_(p1_address_reg_28_), .P1_ADDRESS_REG_27_(p1_address_reg_27_), .P1_ADDRESS_REG_26_(p1_address_reg_26_), .P1_ADDRESS_REG_25_(p1_address_reg_25_), .P1_ADDRESS_REG_24_(p1_address_reg_24_), .P1_ADDRESS_REG_23_(p1_address_reg_23_), .P1_ADDRESS_REG_22_(p1_address_reg_22_), .P1_ADDRESS_REG_21_(p1_address_reg_21_), .P1_ADDRESS_REG_20_(p1_address_reg_20_), .P1_ADDRESS_REG_19_(p1_address_reg_19_), .P1_ADDRESS_REG_18_(p1_address_reg_18_), .P1_ADDRESS_REG_17_(p1_address_reg_17_), .P1_ADDRESS_REG_16_(p1_address_reg_16_), .P1_ADDRESS_REG_15_(p1_address_reg_15_), .P1_ADDRESS_REG_14_(p1_address_reg_14_), .P1_ADDRESS_REG_13_(p1_address_reg_13_), .P1_ADDRESS_REG_12_(p1_address_reg_12_), .P1_ADDRESS_REG_11_(p1_address_reg_11_), .P1_ADDRESS_REG_10_(p1_address_reg_10_), .P1_ADDRESS_REG_9_(p1_address_reg_9_), .P1_ADDRESS_REG_8_(p1_address_reg_8_), .P1_ADDRESS_REG_7_(p1_address_reg_7_), .P1_ADDRESS_REG_6_(p1_address_reg_6_), .P1_ADDRESS_REG_5_(p1_address_reg_5_), .P1_ADDRESS_REG_4_(p1_address_reg_4_), .P1_ADDRESS_REG_3_(p1_address_reg_3_), .P1_ADDRESS_REG_2_(p1_address_reg_2_), .P1_ADDRESS_REG_1_(p1_address_reg_1_), .P1_ADDRESS_REG_0_(p1_address_reg_0_), .U355(u355), .U356(u356), .U357(u357), .U358(u358), .U359(u359), .U360(u360), .U361(u361), .U362(u362), .U363(u363), .U364(u364), .U366(u366), .U367(u367), .U368(u368), .U369(u369), .U370(u370), .U371(u371), .U372(u372), .U373(u373), .U374(u374), .U375(u375), .U347(u347), .U348(u348), .U349(u349), .U350(u350), .U351(u351), .U352(u352), .U353(u353), .U354(u354), .U365(u365), .U376(u376), .P3_W_R_N_REG(p3_w_r_n_reg), .P3_D_C_N_REG(p3_d_c_n_reg), .P3_M_IO_N_REG(p3_m_io_n_reg), .P1_ADS_N_REG(p1_ads_n_reg), .P3_ADS_N_REG(p3_ads_n_reg), .U247(u247), .U246(u246), .U245(u245), .U244(u244), .U243(u243), .U242(u242), .U241(u241), .U240(u240), .U239(u239), .U238(u238), .U237(u237), .U236(u236), .U235(u235), .U234(u234), .U233(u233), .U232(u232), .U231(u231), .U230(u230), .U229(u229), .U228(u228), .U227(u227), .U226(u226), .U225(u225), .U224(u224), .U223(u223), .U222(u222), .U221(u221), .U220(u220), .U219(u219), .U218(u218), .U217(u217), .U216(u216), .U251(u251), .U252(u252), .U253(u253), .U254(u254), .U255(u255), .U256(u256), .U257(u257), .U258(u258), .U259(u259), .U260(u260), .U261(u261), .U262(u262), .U263(u263), .U264(u264), .U265(u265), .U266(u266), .U267(u267), .U268(u268), .U269(u269), .U270(u270), .U271(u271), .U272(u272), .U273(u273), .U274(u274), .U275(u275), .U276(u276), .U277(u277), .U278(u278), .U279(u279), .U280(u280), .U281(u281), .U282(u282), .U212(u212), .U215(u215), .U213(u213), .U214(u214), .P3_U3274(p3_u3274), .P3_U3275(p3_u3275), .P3_U3276(p3_u3276), .P3_U3277(p3_u3277), .P3_U3061(p3_u3061), .P3_U3060(p3_u3060), .P3_U3059(p3_u3059), .P3_U3058(p3_u3058), .P3_U3057(p3_u3057), .P3_U3056(p3_u3056), .P3_U3055(p3_u3055), .P3_U3054(p3_u3054), .P3_U3053(p3_u3053), .P3_U3052(p3_u3052), .P3_U3051(p3_u3051), .P3_U3050(p3_u3050), .P3_U3049(p3_u3049), .P3_U3048(p3_u3048), .P3_U3047(p3_u3047), .P3_U3046(p3_u3046), .P3_U3045(p3_u3045), .P3_U3044(p3_u3044), .P3_U3043(p3_u3043), .P3_U3042(p3_u3042), .P3_U3041(p3_u3041), .P3_U3040(p3_u3040), .P3_U3039(p3_u3039), .P3_U3038(p3_u3038), .P3_U3037(p3_u3037), .P3_U3036(p3_u3036), .P3_U3035(p3_u3035), .P3_U3034(p3_u3034), .P3_U3033(p3_u3033), .P3_U3032(p3_u3032), .P3_U3031(p3_u3031), .P3_U3030(p3_u3030), .P3_U3029(p3_u3029), .P3_U3280(p3_u3280), .P3_U3281(p3_u3281), .P3_U3028(p3_u3028), .P3_U3027(p3_u3027), .P3_U3026(p3_u3026), .P3_U3025(p3_u3025), .P3_U3024(p3_u3024), .P3_U3023(p3_u3023), .P3_U3022(p3_u3022), .P3_U3021(p3_u3021), .P3_U3020(p3_u3020), .P3_U3019(p3_u3019), .P3_U3018(p3_u3018), .P3_U3017(p3_u3017), .P3_U3016(p3_u3016), .P3_U3015(p3_u3015), .P3_U3014(p3_u3014), .P3_U3013(p3_u3013), .P3_U3012(p3_u3012), .P3_U3011(p3_u3011), .P3_U3010(p3_u3010), .P3_U3009(p3_u3009), .P3_U3008(p3_u3008), .P3_U3007(p3_u3007), .P3_U3006(p3_u3006), .P3_U3005(p3_u3005), .P3_U3004(p3_u3004), .P3_U3003(p3_u3003), .P3_U3002(p3_u3002), .P3_U3001(p3_u3001), .P3_U3000(p3_u3000), .P3_U2999(p3_u2999), .P3_U3282(p3_u3282), .P3_U2998(p3_u2998), .P3_U2997(p3_u2997), .P3_U2996(p3_u2996), .P3_U2995(p3_u2995), .P3_U2994(p3_u2994), .P3_U2993(p3_u2993), .P3_U2992(p3_u2992), .P3_U2991(p3_u2991), .P3_U2990(p3_u2990), .P3_U2989(p3_u2989), .P3_U2988(p3_u2988), .P3_U2987(p3_u2987), .P3_U2986(p3_u2986), .P3_U2985(p3_u2985), .P3_U2984(p3_u2984), .P3_U2983(p3_u2983), .P3_U2982(p3_u2982), .P3_U2981(p3_u2981), .P3_U2980(p3_u2980), .P3_U2979(p3_u2979), .P3_U2978(p3_u2978), .P3_U2977(p3_u2977), .P3_U2976(p3_u2976), .P3_U2975(p3_u2975), .P3_U2974(p3_u2974), .P3_U2973(p3_u2973), .P3_U2972(p3_u2972), .P3_U2971(p3_u2971), .P3_U2970(p3_u2970), .P3_U2969(p3_u2969), .P3_U2968(p3_u2968), .P3_U2967(p3_u2967), .P3_U2966(p3_u2966), .P3_U2965(p3_u2965), .P3_U2964(p3_u2964), .P3_U2963(p3_u2963), .P3_U2962(p3_u2962), .P3_U2961(p3_u2961), .P3_U2960(p3_u2960), .P3_U2959(p3_u2959), .P3_U2958(p3_u2958), .P3_U2957(p3_u2957), .P3_U2956(p3_u2956), .P3_U2955(p3_u2955), .P3_U2954(p3_u2954), .P3_U2953(p3_u2953), .P3_U2952(p3_u2952), .P3_U2951(p3_u2951), .P3_U2950(p3_u2950), .P3_U2949(p3_u2949), .P3_U2948(p3_u2948), .P3_U2947(p3_u2947), .P3_U2946(p3_u2946), .P3_U2945(p3_u2945), .P3_U2944(p3_u2944), .P3_U2943(p3_u2943), .P3_U2942(p3_u2942), .P3_U2941(p3_u2941), .P3_U2940(p3_u2940), .P3_U2939(p3_u2939), .P3_U2938(p3_u2938), .P3_U2937(p3_u2937), .P3_U2936(p3_u2936), .P3_U2935(p3_u2935), .P3_U2934(p3_u2934), .P3_U2933(p3_u2933), .P3_U2932(p3_u2932), .P3_U2931(p3_u2931), .P3_U2930(p3_u2930), .P3_U2929(p3_u2929), .P3_U2928(p3_u2928), .P3_U2927(p3_u2927), .P3_U2926(p3_u2926), .P3_U2925(p3_u2925), .P3_U2924(p3_u2924), .P3_U2923(p3_u2923), .P3_U2922(p3_u2922), .P3_U2921(p3_u2921), .P3_U2920(p3_u2920), .P3_U2919(p3_u2919), .P3_U2918(p3_u2918), .P3_U2917(p3_u2917), .P3_U2916(p3_u2916), .P3_U2915(p3_u2915), .P3_U2914(p3_u2914), .P3_U2913(p3_u2913), .P3_U2912(p3_u2912), .P3_U2911(p3_u2911), .P3_U2910(p3_u2910), .P3_U2909(p3_u2909), .P3_U2908(p3_u2908), .P3_U2907(p3_u2907), .P3_U2906(p3_u2906), .P3_U2905(p3_u2905), .P3_U2904(p3_u2904), .P3_U2903(p3_u2903), .P3_U2902(p3_u2902), .P3_U2901(p3_u2901), .P3_U2900(p3_u2900), .P3_U2899(p3_u2899), .P3_U2898(p3_u2898), .P3_U2897(p3_u2897), .P3_U2896(p3_u2896), .P3_U2895(p3_u2895), .P3_U2894(p3_u2894), .P3_U2893(p3_u2893), .P3_U2892(p3_u2892), .P3_U2891(p3_u2891), .P3_U2890(p3_u2890), .P3_U2889(p3_u2889), .P3_U2888(p3_u2888), .P3_U2887(p3_u2887), .P3_U2886(p3_u2886), .P3_U2885(p3_u2885), .P3_U2884(p3_u2884), .P3_U2883(p3_u2883), .P3_U2882(p3_u2882), .P3_U2881(p3_u2881), .P3_U2880(p3_u2880), .P3_U2879(p3_u2879), .P3_U2878(p3_u2878), .P3_U2877(p3_u2877), .P3_U2876(p3_u2876), .P3_U2875(p3_u2875), .P3_U2874(p3_u2874), .P3_U2873(p3_u2873), .P3_U2872(p3_u2872), .P3_U2871(p3_u2871), .P3_U2870(p3_u2870), .P3_U2869(p3_u2869), .P3_U2868(p3_u2868), .P3_U3284(p3_u3284), .P3_U3285(p3_u3285), .P3_U3288(p3_u3288), .P3_U3289(p3_u3289), .P3_U3290(p3_u3290), .P3_U2867(p3_u2867), .P3_U2866(p3_u2866), .P3_U2865(p3_u2865), .P3_U2864(p3_u2864), .P3_U2863(p3_u2863), .P3_U2862(p3_u2862), .P3_U2861(p3_u2861), .P3_U2860(p3_u2860), .P3_U2859(p3_u2859), .P3_U2858(p3_u2858), .P3_U2857(p3_u2857), .P3_U2856(p3_u2856), .P3_U2855(p3_u2855), .P3_U2854(p3_u2854), .P3_U2853(p3_u2853), .P3_U2852(p3_u2852), .P3_U2851(p3_u2851), .P3_U2850(p3_u2850), .P3_U2849(p3_u2849), .P3_U2848(p3_u2848), .P3_U2847(p3_u2847), .P3_U2846(p3_u2846), .P3_U2845(p3_u2845), .P3_U2844(p3_u2844), .P3_U2843(p3_u2843), .P3_U2842(p3_u2842), .P3_U2841(p3_u2841), .P3_U2840(p3_u2840), .P3_U2839(p3_u2839), .P3_U2838(p3_u2838), .P3_U2837(p3_u2837), .P3_U2836(p3_u2836), .P3_U2835(p3_u2835), .P3_U2834(p3_u2834), .P3_U2833(p3_u2833), .P3_U2832(p3_u2832), .P3_U2831(p3_u2831), .P3_U2830(p3_u2830), .P3_U2829(p3_u2829), .P3_U2828(p3_u2828), .P3_U2827(p3_u2827), .P3_U2826(p3_u2826), .P3_U2825(p3_u2825), .P3_U2824(p3_u2824), .P3_U2823(p3_u2823), .P3_U2822(p3_u2822), .P3_U2821(p3_u2821), .P3_U2820(p3_u2820), .P3_U2819(p3_u2819), .P3_U2818(p3_u2818), .P3_U2817(p3_u2817), .P3_U2816(p3_u2816), .P3_U2815(p3_u2815), .P3_U2814(p3_u2814), .P3_U2813(p3_u2813), .P3_U2812(p3_u2812), .P3_U2811(p3_u2811), .P3_U2810(p3_u2810), .P3_U2809(p3_u2809), .P3_U2808(p3_u2808), .P3_U2807(p3_u2807), .P3_U2806(p3_u2806), .P3_U2805(p3_u2805), .P3_U2804(p3_u2804), .P3_U2803(p3_u2803), .P3_U2802(p3_u2802), .P3_U2801(p3_u2801), .P3_U2800(p3_u2800), .P3_U2799(p3_u2799), .P3_U2798(p3_u2798), .P3_U2797(p3_u2797), .P3_U2796(p3_u2796), .P3_U2795(p3_u2795), .P3_U2794(p3_u2794), .P3_U2793(p3_u2793), .P3_U2792(p3_u2792), .P3_U2791(p3_u2791), .P3_U2790(p3_u2790), .P3_U2789(p3_u2789), .P3_U2788(p3_u2788), .P3_U2787(p3_u2787), .P3_U2786(p3_u2786), .P3_U2785(p3_u2785), .P3_U2784(p3_u2784), .P3_U2783(p3_u2783), .P3_U2782(p3_u2782), .P3_U2781(p3_u2781), .P3_U2780(p3_u2780), .P3_U2779(p3_u2779), .P3_U2778(p3_u2778), .P3_U2777(p3_u2777), .P3_U2776(p3_u2776), .P3_U2775(p3_u2775), .P3_U2774(p3_u2774), .P3_U2773(p3_u2773), .P3_U2772(p3_u2772), .P3_U2771(p3_u2771), .P3_U2770(p3_u2770), .P3_U2769(p3_u2769), .P3_U2768(p3_u2768), .P3_U2767(p3_u2767), .P3_U2766(p3_u2766), .P3_U2765(p3_u2765), .P3_U2764(p3_u2764), .P3_U2763(p3_u2763), .P3_U2762(p3_u2762), .P3_U2761(p3_u2761), .P3_U2760(p3_u2760), .P3_U2759(p3_u2759), .P3_U2758(p3_u2758), .P3_U2757(p3_u2757), .P3_U2756(p3_u2756), .P3_U2755(p3_u2755), .P3_U2754(p3_u2754), .P3_U2753(p3_u2753), .P3_U2752(p3_u2752), .P3_U2751(p3_u2751), .P3_U2750(p3_u2750), .P3_U2749(p3_u2749), .P3_U2748(p3_u2748), .P3_U2747(p3_u2747), .P3_U2746(p3_u2746), .P3_U2745(p3_u2745), .P3_U2744(p3_u2744), .P3_U2743(p3_u2743), .P3_U2742(p3_u2742), .P3_U2741(p3_u2741), .P3_U2740(p3_u2740), .P3_U2739(p3_u2739), .P3_U2738(p3_u2738), .P3_U2737(p3_u2737), .P3_U2736(p3_u2736), .P3_U2735(p3_u2735), .P3_U2734(p3_u2734), .P3_U2733(p3_u2733), .P3_U2732(p3_u2732), .P3_U2731(p3_u2731), .P3_U2730(p3_u2730), .P3_U2729(p3_u2729), .P3_U2728(p3_u2728), .P3_U2727(p3_u2727), .P3_U2726(p3_u2726), .P3_U2725(p3_u2725), .P3_U2724(p3_u2724), .P3_U2723(p3_u2723), .P3_U2722(p3_u2722), .P3_U2721(p3_u2721), .P3_U2720(p3_u2720), .P3_U2719(p3_u2719), .P3_U2718(p3_u2718), .P3_U2717(p3_u2717), .P3_U2716(p3_u2716), .P3_U2715(p3_u2715), .P3_U2714(p3_u2714), .P3_U2713(p3_u2713), .P3_U2712(p3_u2712), .P3_U2711(p3_u2711), .P3_U2710(p3_u2710), .P3_U2709(p3_u2709), .P3_U2708(p3_u2708), .P3_U2707(p3_u2707), .P3_U2706(p3_u2706), .P3_U2705(p3_u2705), .P3_U2704(p3_u2704), .P3_U2703(p3_u2703), .P3_U2702(p3_u2702), .P3_U2701(p3_u2701), .P3_U2700(p3_u2700), .P3_U2699(p3_u2699), .P3_U2698(p3_u2698), .P3_U2697(p3_u2697), .P3_U2696(p3_u2696), .P3_U2695(p3_u2695), .P3_U2694(p3_u2694), .P3_U2693(p3_u2693), .P3_U2692(p3_u2692), .P3_U2691(p3_u2691), .P3_U2690(p3_u2690), .P3_U2689(p3_u2689), .P3_U2688(p3_u2688), .P3_U2687(p3_u2687), .P3_U2686(p3_u2686), .P3_U2685(p3_u2685), .P3_U2684(p3_u2684), .P3_U2683(p3_u2683), .P3_U2682(p3_u2682), .P3_U2681(p3_u2681), .P3_U2680(p3_u2680), .P3_U2679(p3_u2679), .P3_U2678(p3_u2678), .P3_U2677(p3_u2677), .P3_U2676(p3_u2676), .P3_U2675(p3_u2675), .P3_U2674(p3_u2674), .P3_U2673(p3_u2673), .P3_U2672(p3_u2672), .P3_U2671(p3_u2671), .P3_U2670(p3_u2670), .P3_U2669(p3_u2669), .P3_U2668(p3_u2668), .P3_U2667(p3_u2667), .P3_U2666(p3_u2666), .P3_U2665(p3_u2665), .P3_U2664(p3_u2664), .P3_U2663(p3_u2663), .P3_U2662(p3_u2662), .P3_U2661(p3_u2661), .P3_U2660(p3_u2660), .P3_U2659(p3_u2659), .P3_U2658(p3_u2658), .P3_U2657(p3_u2657), .P3_U2656(p3_u2656), .P3_U2655(p3_u2655), .P3_U2654(p3_u2654), .P3_U2653(p3_u2653), .P3_U2652(p3_u2652), .P3_U2651(p3_u2651), .P3_U2650(p3_u2650), .P3_U2649(p3_u2649), .P3_U2648(p3_u2648), .P3_U2647(p3_u2647), .P3_U2646(p3_u2646), .P3_U2645(p3_u2645), .P3_U2644(p3_u2644), .P3_U2643(p3_u2643), .P3_U2642(p3_u2642), .P3_U2641(p3_u2641), .P3_U2640(p3_u2640), .P3_U2639(p3_u2639), .P3_U3292(p3_u3292), .P3_U2638(p3_u2638), .P3_U3293(p3_u3293), .P3_U3294(p3_u3294), .P3_U2637(p3_u2637), .P3_U3295(p3_u3295), .P3_U2636(p3_u2636), .P3_U3296(p3_u3296), .P3_U2635(p3_u2635), .P3_U3297(p3_u3297), .P3_U2634(p3_u2634), .P3_U2633(p3_u2633), .P3_U3298(p3_u3298), .P3_U3299(p3_u3299), .P2_U3585(p2_u3585), .P2_U3586(p2_u3586), .P2_U3587(p2_u3587), .P2_U3588(p2_u3588), .P2_U3241(p2_u3241), .P2_U3240(p2_u3240), .P2_U3239(p2_u3239), .P2_U3238(p2_u3238), .P2_U3237(p2_u3237), .P2_U3236(p2_u3236), .P2_U3235(p2_u3235), .P2_U3234(p2_u3234), .P2_U3233(p2_u3233), .P2_U3232(p2_u3232), .P2_U3231(p2_u3231), .P2_U3230(p2_u3230), .P2_U3229(p2_u3229), .P2_U3228(p2_u3228), .P2_U3227(p2_u3227), .P2_U3226(p2_u3226), .P2_U3225(p2_u3225), .P2_U3224(p2_u3224), .P2_U3223(p2_u3223), .P2_U3222(p2_u3222), .P2_U3221(p2_u3221), .P2_U3220(p2_u3220), .P2_U3219(p2_u3219), .P2_U3218(p2_u3218), .P2_U3217(p2_u3217), .P2_U3216(p2_u3216), .P2_U3215(p2_u3215), .P2_U3214(p2_u3214), .P2_U3213(p2_u3213), .P2_U3212(p2_u3212), .P2_U3211(p2_u3211), .P2_U3210(p2_u3210), .P2_U3209(p2_u3209), .P2_U3591(p2_u3591), .P2_U3592(p2_u3592), .P2_U3208(p2_u3208), .P2_U3207(p2_u3207), .P2_U3206(p2_u3206), .P2_U3205(p2_u3205), .P2_U3204(p2_u3204), .P2_U3203(p2_u3203), .P2_U3202(p2_u3202), .P2_U3201(p2_u3201), .P2_U3200(p2_u3200), .P2_U3199(p2_u3199), .P2_U3198(p2_u3198), .P2_U3197(p2_u3197), .P2_U3196(p2_u3196), .P2_U3195(p2_u3195), .P2_U3194(p2_u3194), .P2_U3193(p2_u3193), .P2_U3192(p2_u3192), .P2_U3191(p2_u3191), .P2_U3190(p2_u3190), .P2_U3189(p2_u3189), .P2_U3188(p2_u3188), .P2_U3187(p2_u3187), .P2_U3186(p2_u3186), .P2_U3185(p2_u3185), .P2_U3184(p2_u3184), .P2_U3183(p2_u3183), .P2_U3182(p2_u3182), .P2_U3181(p2_u3181), .P2_U3180(p2_u3180), .P2_U3179(p2_u3179), .P2_U3593(p2_u3593), .P2_U3178(p2_u3178), .P2_U3177(p2_u3177), .P2_U3176(p2_u3176), .P2_U3175(p2_u3175), .P2_U3174(p2_u3174), .P2_U3173(p2_u3173), .P2_U3172(p2_u3172), .P2_U3171(p2_u3171), .P2_U3170(p2_u3170), .P2_U3169(p2_u3169), .P2_U3168(p2_u3168), .P2_U3167(p2_u3167), .P2_U3166(p2_u3166), .P2_U3165(p2_u3165), .P2_U3164(p2_u3164), .P2_U3163(p2_u3163), .P2_U3162(p2_u3162), .P2_U3161(p2_u3161), .P2_U3160(p2_u3160), .P2_U3159(p2_u3159), .P2_U3158(p2_u3158), .P2_U3157(p2_u3157), .P2_U3156(p2_u3156), .P2_U3155(p2_u3155), .P2_U3154(p2_u3154), .P2_U3153(p2_u3153), .P2_U3152(p2_u3152), .P2_U3151(p2_u3151), .P2_U3150(p2_u3150), .P2_U3149(p2_u3149), .P2_U3148(p2_u3148), .P2_U3147(p2_u3147), .P2_U3146(p2_u3146), .P2_U3145(p2_u3145), .P2_U3144(p2_u3144), .P2_U3143(p2_u3143), .P2_U3142(p2_u3142), .P2_U3141(p2_u3141), .P2_U3140(p2_u3140), .P2_U3139(p2_u3139), .P2_U3138(p2_u3138), .P2_U3137(p2_u3137), .P2_U3136(p2_u3136), .P2_U3135(p2_u3135), .P2_U3134(p2_u3134), .P2_U3133(p2_u3133), .P2_U3132(p2_u3132), .P2_U3131(p2_u3131), .P2_U3130(p2_u3130), .P2_U3129(p2_u3129), .P2_U3128(p2_u3128), .P2_U3127(p2_u3127), .P2_U3126(p2_u3126), .P2_U3125(p2_u3125), .P2_U3124(p2_u3124), .P2_U3123(p2_u3123), .P2_U3122(p2_u3122), .P2_U3121(p2_u3121), .P2_U3120(p2_u3120), .P2_U3119(p2_u3119), .P2_U3118(p2_u3118), .P2_U3117(p2_u3117), .P2_U3116(p2_u3116), .P2_U3115(p2_u3115), .P2_U3114(p2_u3114), .P2_U3113(p2_u3113), .P2_U3112(p2_u3112), .P2_U3111(p2_u3111), .P2_U3110(p2_u3110), .P2_U3109(p2_u3109), .P2_U3108(p2_u3108), .P2_U3107(p2_u3107), .P2_U3106(p2_u3106), .P2_U3105(p2_u3105), .P2_U3104(p2_u3104), .P2_U3103(p2_u3103), .P2_U3102(p2_u3102), .P2_U3101(p2_u3101), .P2_U3100(p2_u3100), .P2_U3099(p2_u3099), .P2_U3098(p2_u3098), .P2_U3097(p2_u3097), .P2_U3096(p2_u3096), .P2_U3095(p2_u3095), .P2_U3094(p2_u3094), .P2_U3093(p2_u3093), .P2_U3092(p2_u3092), .P2_U3091(p2_u3091), .P2_U3090(p2_u3090), .P2_U3089(p2_u3089), .P2_U3088(p2_u3088), .P2_U3087(p2_u3087), .P2_U3086(p2_u3086), .P2_U3085(p2_u3085), .P2_U3084(p2_u3084), .P2_U3083(p2_u3083), .P2_U3082(p2_u3082), .P2_U3081(p2_u3081), .P2_U3080(p2_u3080), .P2_U3079(p2_u3079), .P2_U3078(p2_u3078), .P2_U3077(p2_u3077), .P2_U3076(p2_u3076), .P2_U3075(p2_u3075), .P2_U3074(p2_u3074), .P2_U3073(p2_u3073), .P2_U3072(p2_u3072), .P2_U3071(p2_u3071), .P2_U3070(p2_u3070), .P2_U3069(p2_u3069), .P2_U3068(p2_u3068), .P2_U3067(p2_u3067), .P2_U3066(p2_u3066), .P2_U3065(p2_u3065), .P2_U3064(p2_u3064), .P2_U3063(p2_u3063), .P2_U3062(p2_u3062), .P2_U3061(p2_u3061), .P2_U3060(p2_u3060), .P2_U3059(p2_u3059), .P2_U3058(p2_u3058), .P2_U3057(p2_u3057), .P2_U3056(p2_u3056), .P2_U3055(p2_u3055), .P2_U3054(p2_u3054), .P2_U3053(p2_u3053), .P2_U3052(p2_u3052), .P2_U3051(p2_u3051), .P2_U3050(p2_u3050), .P2_U3049(p2_u3049), .P2_U3048(p2_u3048), .P2_U3595(p2_u3595), .P2_U3596(p2_u3596), .P2_U3599(p2_u3599), .P2_U3600(p2_u3600), .P2_U3601(p2_u3601), .P2_U3047(p2_u3047), .P2_U3602(p2_u3602), .P2_U3603(p2_u3603), .P2_U3604(p2_u3604), .P2_U3605(p2_u3605), .P2_U3046(p2_u3046), .P2_U3045(p2_u3045), .P2_U3044(p2_u3044), .P2_U3043(p2_u3043), .P2_U3042(p2_u3042), .P2_U3041(p2_u3041), .P2_U3040(p2_u3040), .P2_U3039(p2_u3039), .P2_U3038(p2_u3038), .P2_U3037(p2_u3037), .P2_U3036(p2_u3036), .P2_U3035(p2_u3035), .P2_U3034(p2_u3034), .P2_U3033(p2_u3033), .P2_U3032(p2_u3032), .P2_U3031(p2_u3031), .P2_U3030(p2_u3030), .P2_U3029(p2_u3029), .P2_U3028(p2_u3028), .P2_U3027(p2_u3027), .P2_U3026(p2_u3026), .P2_U3025(p2_u3025), .P2_U3024(p2_u3024), .P2_U3023(p2_u3023), .P2_U3022(p2_u3022), .P2_U3021(p2_u3021), .P2_U3020(p2_u3020), .P2_U3019(p2_u3019), .P2_U3018(p2_u3018), .P2_U3017(p2_u3017), .P2_U3016(p2_u3016), .P2_U3015(p2_u3015), .P2_U3014(p2_u3014), .P2_U3013(p2_u3013), .P2_U3012(p2_u3012), .P2_U3011(p2_u3011), .P2_U3010(p2_u3010), .P2_U3009(p2_u3009), .P2_U3008(p2_u3008), .P2_U3007(p2_u3007), .P2_U3006(p2_u3006), .P2_U3005(p2_u3005), .P2_U3004(p2_u3004), .P2_U3003(p2_u3003), .P2_U3002(p2_u3002), .P2_U3001(p2_u3001), .P2_U3000(p2_u3000), .P2_U2999(p2_u2999), .P2_U2998(p2_u2998), .P2_U2997(p2_u2997), .P2_U2996(p2_u2996), .P2_U2995(p2_u2995), .P2_U2994(p2_u2994), .P2_U2993(p2_u2993), .P2_U2992(p2_u2992), .P2_U2991(p2_u2991), .P2_U2990(p2_u2990), .P2_U2989(p2_u2989), .P2_U2988(p2_u2988), .P2_U2987(p2_u2987), .P2_U2986(p2_u2986), .P2_U2985(p2_u2985), .P2_U2984(p2_u2984), .P2_U2983(p2_u2983), .P2_U2982(p2_u2982), .P2_U2981(p2_u2981), .P2_U2980(p2_u2980), .P2_U2979(p2_u2979), .P2_U2978(p2_u2978), .P2_U2977(p2_u2977), .P2_U2976(p2_u2976), .P2_U2975(p2_u2975), .P2_U2974(p2_u2974), .P2_U2973(p2_u2973), .P2_U2972(p2_u2972), .P2_U2971(p2_u2971), .P2_U2970(p2_u2970), .P2_U2969(p2_u2969), .P2_U2968(p2_u2968), .P2_U2967(p2_u2967), .P2_U2966(p2_u2966), .P2_U2965(p2_u2965), .P2_U2964(p2_u2964), .P2_U2963(p2_u2963), .P2_U2962(p2_u2962), .P2_U2961(p2_u2961), .P2_U2960(p2_u2960), .P2_U2959(p2_u2959), .P2_U2958(p2_u2958), .P2_U2957(p2_u2957), .P2_U2956(p2_u2956), .P2_U2955(p2_u2955), .P2_U2954(p2_u2954), .P2_U2953(p2_u2953), .P2_U2952(p2_u2952), .P2_U2951(p2_u2951), .P2_U2950(p2_u2950), .P2_U2949(p2_u2949), .P2_U2948(p2_u2948), .P2_U2947(p2_u2947), .P2_U2946(p2_u2946), .P2_U2945(p2_u2945), .P2_U2944(p2_u2944), .P2_U2943(p2_u2943), .P2_U2942(p2_u2942), .P2_U2941(p2_u2941), .P2_U2940(p2_u2940), .P2_U2939(p2_u2939), .P2_U2938(p2_u2938), .P2_U2937(p2_u2937), .P2_U2936(p2_u2936), .P2_U2935(p2_u2935), .P2_U2934(p2_u2934), .P2_U2933(p2_u2933), .P2_U2932(p2_u2932), .P2_U2931(p2_u2931), .P2_U2930(p2_u2930), .P2_U2929(p2_u2929), .P2_U2928(p2_u2928), .P2_U2927(p2_u2927), .P2_U2926(p2_u2926), .P2_U2925(p2_u2925), .P2_U2924(p2_u2924), .P2_U2923(p2_u2923), .P2_U2922(p2_u2922), .P2_U2921(p2_u2921), .P2_U2920(p2_u2920), .P2_U2919(p2_u2919), .P2_U2918(p2_u2918), .P2_U2917(p2_u2917), .P2_U2916(p2_u2916), .P2_U2915(p2_u2915), .P2_U2914(p2_u2914), .P2_U2913(p2_u2913), .P2_U2912(p2_u2912), .P2_U2911(p2_u2911), .P2_U2910(p2_u2910), .P2_U2909(p2_u2909), .P2_U2908(p2_u2908), .P2_U2907(p2_u2907), .P2_U2906(p2_u2906), .P2_U2905(p2_u2905), .P2_U2904(p2_u2904), .P2_U2903(p2_u2903), .P2_U2902(p2_u2902), .P2_U2901(p2_u2901), .P2_U2900(p2_u2900), .P2_U2899(p2_u2899), .P2_U2898(p2_u2898), .P2_U2897(p2_u2897), .P2_U2896(p2_u2896), .P2_U2895(p2_u2895), .P2_U2894(p2_u2894), .P2_U2893(p2_u2893), .P2_U2892(p2_u2892), .P2_U2891(p2_u2891), .P2_U2890(p2_u2890), .P2_U2889(p2_u2889), .P2_U2888(p2_u2888), .P2_U2887(p2_u2887), .P2_U2886(p2_u2886), .P2_U2885(p2_u2885), .P2_U2884(p2_u2884), .P2_U2883(p2_u2883), .P2_U2882(p2_u2882), .P2_U2881(p2_u2881), .P2_U2880(p2_u2880), .P2_U2879(p2_u2879), .P2_U2878(p2_u2878), .P2_U2877(p2_u2877), .P2_U2876(p2_u2876), .P2_U2875(p2_u2875), .P2_U2874(p2_u2874), .P2_U2873(p2_u2873), .P2_U2872(p2_u2872), .P2_U2871(p2_u2871), .P2_U2870(p2_u2870), .P2_U2869(p2_u2869), .P2_U2868(p2_u2868), .P2_U2867(p2_u2867), .P2_U2866(p2_u2866), .P2_U2865(p2_u2865), .P2_U2864(p2_u2864), .P2_U2863(p2_u2863), .P2_U2862(p2_u2862), .P2_U2861(p2_u2861), .P2_U2860(p2_u2860), .P2_U2859(p2_u2859), .P2_U2858(p2_u2858), .P2_U2857(p2_u2857), .P2_U2856(p2_u2856), .P2_U2855(p2_u2855), .P2_U2854(p2_u2854), .P2_U2853(p2_u2853), .P2_U2852(p2_u2852), .P2_U2851(p2_u2851), .P2_U2850(p2_u2850), .P2_U2849(p2_u2849), .P2_U2848(p2_u2848), .P2_U2847(p2_u2847), .P2_U2846(p2_u2846), .P2_U2845(p2_u2845), .P2_U2844(p2_u2844), .P2_U2843(p2_u2843), .P2_U2842(p2_u2842), .P2_U2841(p2_u2841), .P2_U2840(p2_u2840), .P2_U2839(p2_u2839), .P2_U2838(p2_u2838), .P2_U2837(p2_u2837), .P2_U2836(p2_u2836), .P2_U2835(p2_u2835), .P2_U2834(p2_u2834), .P2_U2833(p2_u2833), .P2_U2832(p2_u2832), .P2_U2831(p2_u2831), .P2_U2830(p2_u2830), .P2_U2829(p2_u2829), .P2_U2828(p2_u2828), .P2_U2827(p2_u2827), .P2_U2826(p2_u2826), .P2_U2825(p2_u2825), .P2_U2824(p2_u2824), .P2_U2823(p2_u2823), .P2_U2822(p2_u2822), .P2_U2821(p2_u2821), .P2_U2820(p2_u2820), .P2_U3608(p2_u3608), .P2_U2819(p2_u2819), .P2_U3609(p2_u3609), .P2_U2818(p2_u2818), .P2_U3610(p2_u3610), .P2_U2817(p2_u2817), .P2_U3611(p2_u3611), .P2_U2816(p2_u2816), .P2_U2815(p2_u2815), .P2_U3612(p2_u3612), .P2_U2814(p2_u2814), .P1_U3458(p1_u3458), .P1_U3459(p1_u3459), .P1_U3460(p1_u3460), .P1_U3461(p1_u3461), .P1_U3226(p1_u3226), .P1_U3225(p1_u3225), .P1_U3224(p1_u3224), .P1_U3223(p1_u3223), .P1_U3222(p1_u3222), .P1_U3221(p1_u3221), .P1_U3220(p1_u3220), .P1_U3219(p1_u3219), .P1_U3218(p1_u3218), .P1_U3217(p1_u3217), .P1_U3216(p1_u3216), .P1_U3215(p1_u3215), .P1_U3214(p1_u3214), .P1_U3213(p1_u3213), .P1_U3212(p1_u3212), .P1_U3211(p1_u3211), .P1_U3210(p1_u3210), .P1_U3209(p1_u3209), .P1_U3208(p1_u3208), .P1_U3207(p1_u3207), .P1_U3206(p1_u3206), .P1_U3205(p1_u3205), .P1_U3204(p1_u3204), .P1_U3203(p1_u3203), .P1_U3202(p1_u3202), .P1_U3201(p1_u3201), .P1_U3200(p1_u3200), .P1_U3199(p1_u3199), .P1_U3198(p1_u3198), .P1_U3197(p1_u3197), .P1_U3196(p1_u3196), .P1_U3195(p1_u3195), .P1_U3194(p1_u3194), .P1_U3464(p1_u3464), .P1_U3465(p1_u3465), .P1_U3193(p1_u3193), .P1_U3192(p1_u3192), .P1_U3191(p1_u3191), .P1_U3190(p1_u3190), .P1_U3189(p1_u3189), .P1_U3188(p1_u3188), .P1_U3187(p1_u3187), .P1_U3186(p1_u3186), .P1_U3185(p1_u3185), .P1_U3184(p1_u3184), .P1_U3183(p1_u3183), .P1_U3182(p1_u3182), .P1_U3181(p1_u3181), .P1_U3180(p1_u3180), .P1_U3179(p1_u3179), .P1_U3178(p1_u3178), .P1_U3177(p1_u3177), .P1_U3176(p1_u3176), .P1_U3175(p1_u3175), .P1_U3174(p1_u3174), .P1_U3173(p1_u3173), .P1_U3172(p1_u3172), .P1_U3171(p1_u3171), .P1_U3170(p1_u3170), .P1_U3169(p1_u3169), .P1_U3168(p1_u3168), .P1_U3167(p1_u3167), .P1_U3166(p1_u3166), .P1_U3165(p1_u3165), .P1_U3164(p1_u3164), .P1_U3466(p1_u3466), .P1_U3163(p1_u3163), .P1_U3162(p1_u3162), .P1_U3161(p1_u3161), .P1_U3160(p1_u3160), .P1_U3159(p1_u3159), .P1_U3158(p1_u3158), .P1_U3157(p1_u3157), .P1_U3156(p1_u3156), .P1_U3155(p1_u3155), .P1_U3154(p1_u3154), .P1_U3153(p1_u3153), .P1_U3152(p1_u3152), .P1_U3151(p1_u3151), .P1_U3150(p1_u3150), .P1_U3149(p1_u3149), .P1_U3148(p1_u3148), .P1_U3147(p1_u3147), .P1_U3146(p1_u3146), .P1_U3145(p1_u3145), .P1_U3144(p1_u3144), .P1_U3143(p1_u3143), .P1_U3142(p1_u3142), .P1_U3141(p1_u3141), .P1_U3140(p1_u3140), .P1_U3139(p1_u3139), .P1_U3138(p1_u3138), .P1_U3137(p1_u3137), .P1_U3136(p1_u3136), .P1_U3135(p1_u3135), .P1_U3134(p1_u3134), .P1_U3133(p1_u3133), .P1_U3132(p1_u3132), .P1_U3131(p1_u3131), .P1_U3130(p1_u3130), .P1_U3129(p1_u3129), .P1_U3128(p1_u3128), .P1_U3127(p1_u3127), .P1_U3126(p1_u3126), .P1_U3125(p1_u3125), .P1_U3124(p1_u3124), .P1_U3123(p1_u3123), .P1_U3122(p1_u3122), .P1_U3121(p1_u3121), .P1_U3120(p1_u3120), .P1_U3119(p1_u3119), .P1_U3118(p1_u3118), .P1_U3117(p1_u3117), .P1_U3116(p1_u3116), .P1_U3115(p1_u3115), .P1_U3114(p1_u3114), .P1_U3113(p1_u3113), .P1_U3112(p1_u3112), .P1_U3111(p1_u3111), .P1_U3110(p1_u3110), .P1_U3109(p1_u3109), .P1_U3108(p1_u3108), .P1_U3107(p1_u3107), .P1_U3106(p1_u3106), .P1_U3105(p1_u3105), .P1_U3104(p1_u3104), .P1_U3103(p1_u3103), .P1_U3102(p1_u3102), .P1_U3101(p1_u3101), .P1_U3100(p1_u3100), .P1_U3099(p1_u3099), .P1_U3098(p1_u3098), .P1_U3097(p1_u3097), .P1_U3096(p1_u3096), .P1_U3095(p1_u3095), .P1_U3094(p1_u3094), .P1_U3093(p1_u3093), .P1_U3092(p1_u3092), .P1_U3091(p1_u3091), .P1_U3090(p1_u3090), .P1_U3089(p1_u3089), .P1_U3088(p1_u3088), .P1_U3087(p1_u3087), .P1_U3086(p1_u3086), .P1_U3085(p1_u3085), .P1_U3084(p1_u3084), .P1_U3083(p1_u3083), .P1_U3082(p1_u3082), .P1_U3081(p1_u3081), .P1_U3080(p1_u3080), .P1_U3079(p1_u3079), .P1_U3078(p1_u3078), .P1_U3077(p1_u3077), .P1_U3076(p1_u3076), .P1_U3075(p1_u3075), .P1_U3074(p1_u3074), .P1_U3073(p1_u3073), .P1_U3072(p1_u3072), .P1_U3071(p1_u3071), .P1_U3070(p1_u3070), .P1_U3069(p1_u3069), .P1_U3068(p1_u3068), .P1_U3067(p1_u3067), .P1_U3066(p1_u3066), .P1_U3065(p1_u3065), .P1_U3064(p1_u3064), .P1_U3063(p1_u3063), .P1_U3062(p1_u3062), .P1_U3061(p1_u3061), .P1_U3060(p1_u3060), .P1_U3059(p1_u3059), .P1_U3058(p1_u3058), .P1_U3057(p1_u3057), .P1_U3056(p1_u3056), .P1_U3055(p1_u3055), .P1_U3054(p1_u3054), .P1_U3053(p1_u3053), .P1_U3052(p1_u3052), .P1_U3051(p1_u3051), .P1_U3050(p1_u3050), .P1_U3049(p1_u3049), .P1_U3048(p1_u3048), .P1_U3047(p1_u3047), .P1_U3046(p1_u3046), .P1_U3045(p1_u3045), .P1_U3044(p1_u3044), .P1_U3043(p1_u3043), .P1_U3042(p1_u3042), .P1_U3041(p1_u3041), .P1_U3040(p1_u3040), .P1_U3039(p1_u3039), .P1_U3038(p1_u3038), .P1_U3037(p1_u3037), .P1_U3036(p1_u3036), .P1_U3035(p1_u3035), .P1_U3034(p1_u3034), .P1_U3033(p1_u3033), .P1_U3468(p1_u3468), .P1_U3469(p1_u3469), .P1_U3472(p1_u3472), .P1_U3473(p1_u3473), .P1_U3474(p1_u3474), .P1_U3032(p1_u3032), .P1_U3475(p1_u3475), .P1_U3476(p1_u3476), .P1_U3477(p1_u3477), .P1_U3478(p1_u3478), .P1_U3031(p1_u3031), .P1_U3030(p1_u3030), .P1_U3029(p1_u3029), .P1_U3028(p1_u3028), .P1_U3027(p1_u3027), .P1_U3026(p1_u3026), .P1_U3025(p1_u3025), .P1_U3024(p1_u3024), .P1_U3023(p1_u3023), .P1_U3022(p1_u3022), .P1_U3021(p1_u3021), .P1_U3020(p1_u3020), .P1_U3019(p1_u3019), .P1_U3018(p1_u3018), .P1_U3017(p1_u3017), .P1_U3016(p1_u3016), .P1_U3015(p1_u3015), .P1_U3014(p1_u3014), .P1_U3013(p1_u3013), .P1_U3012(p1_u3012), .P1_U3011(p1_u3011), .P1_U3010(p1_u3010), .P1_U3009(p1_u3009), .P1_U3008(p1_u3008), .P1_U3007(p1_u3007), .P1_U3006(p1_u3006), .P1_U3005(p1_u3005), .P1_U3004(p1_u3004), .P1_U3003(p1_u3003), .P1_U3002(p1_u3002), .P1_U3001(p1_u3001), .P1_U3000(p1_u3000), .P1_U2999(p1_u2999), .P1_U2998(p1_u2998), .P1_U2997(p1_u2997), .P1_U2996(p1_u2996), .P1_U2995(p1_u2995), .P1_U2994(p1_u2994), .P1_U2993(p1_u2993), .P1_U2992(p1_u2992), .P1_U2991(p1_u2991), .P1_U2990(p1_u2990), .P1_U2989(p1_u2989), .P1_U2988(p1_u2988), .P1_U2987(p1_u2987), .P1_U2986(p1_u2986), .P1_U2985(p1_u2985), .P1_U2984(p1_u2984), .P1_U2983(p1_u2983), .P1_U2982(p1_u2982), .P1_U2981(p1_u2981), .P1_U2980(p1_u2980), .P1_U2979(p1_u2979), .P1_U2978(p1_u2978), .P1_U2977(p1_u2977), .P1_U2976(p1_u2976), .P1_U2975(p1_u2975), .P1_U2974(p1_u2974), .P1_U2973(p1_u2973), .P1_U2972(p1_u2972), .P1_U2971(p1_u2971), .P1_U2970(p1_u2970), .P1_U2969(p1_u2969), .P1_U2968(p1_u2968), .P1_U2967(p1_u2967), .P1_U2966(p1_u2966), .P1_U2965(p1_u2965), .P1_U2964(p1_u2964), .P1_U2963(p1_u2963), .P1_U2962(p1_u2962), .P1_U2961(p1_u2961), .P1_U2960(p1_u2960), .P1_U2959(p1_u2959), .P1_U2958(p1_u2958), .P1_U2957(p1_u2957), .P1_U2956(p1_u2956), .P1_U2955(p1_u2955), .P1_U2954(p1_u2954), .P1_U2953(p1_u2953), .P1_U2952(p1_u2952), .P1_U2951(p1_u2951), .P1_U2950(p1_u2950), .P1_U2949(p1_u2949), .P1_U2948(p1_u2948), .P1_U2947(p1_u2947), .P1_U2946(p1_u2946), .P1_U2945(p1_u2945), .P1_U2944(p1_u2944), .P1_U2943(p1_u2943), .P1_U2942(p1_u2942), .P1_U2941(p1_u2941), .P1_U2940(p1_u2940), .P1_U2939(p1_u2939), .P1_U2938(p1_u2938), .P1_U2937(p1_u2937), .P1_U2936(p1_u2936), .P1_U2935(p1_u2935), .P1_U2934(p1_u2934), .P1_U2933(p1_u2933), .P1_U2932(p1_u2932), .P1_U2931(p1_u2931), .P1_U2930(p1_u2930), .P1_U2929(p1_u2929), .P1_U2928(p1_u2928), .P1_U2927(p1_u2927), .P1_U2926(p1_u2926), .P1_U2925(p1_u2925), .P1_U2924(p1_u2924), .P1_U2923(p1_u2923), .P1_U2922(p1_u2922), .P1_U2921(p1_u2921), .P1_U2920(p1_u2920), .P1_U2919(p1_u2919), .P1_U2918(p1_u2918), .P1_U2917(p1_u2917), .P1_U2916(p1_u2916), .P1_U2915(p1_u2915), .P1_U2914(p1_u2914), .P1_U2913(p1_u2913), .P1_U2912(p1_u2912), .P1_U2911(p1_u2911), .P1_U2910(p1_u2910), .P1_U2909(p1_u2909), .P1_U2908(p1_u2908), .P1_U2907(p1_u2907), .P1_U2906(p1_u2906), .P1_U2905(p1_u2905), .P1_U2904(p1_u2904), .P1_U2903(p1_u2903), .P1_U2902(p1_u2902), .P1_U2901(p1_u2901), .P1_U2900(p1_u2900), .P1_U2899(p1_u2899), .P1_U2898(p1_u2898), .P1_U2897(p1_u2897), .P1_U2896(p1_u2896), .P1_U2895(p1_u2895), .P1_U2894(p1_u2894), .P1_U2893(p1_u2893), .P1_U2892(p1_u2892), .P1_U2891(p1_u2891), .P1_U2890(p1_u2890), .P1_U2889(p1_u2889), .P1_U2888(p1_u2888), .P1_U2887(p1_u2887), .P1_U2886(p1_u2886), .P1_U2885(p1_u2885), .P1_U2884(p1_u2884), .P1_U2883(p1_u2883), .P1_U2882(p1_u2882), .P1_U2881(p1_u2881), .P1_U2880(p1_u2880), .P1_U2879(p1_u2879), .P1_U2878(p1_u2878), .P1_U2877(p1_u2877), .P1_U2876(p1_u2876), .P1_U2875(p1_u2875), .P1_U2874(p1_u2874), .P1_U2873(p1_u2873), .P1_U2872(p1_u2872), .P1_U2871(p1_u2871), .P1_U2870(p1_u2870), .P1_U2869(p1_u2869), .P1_U2868(p1_u2868), .P1_U2867(p1_u2867), .P1_U2866(p1_u2866), .P1_U2865(p1_u2865), .P1_U2864(p1_u2864), .P1_U2863(p1_u2863), .P1_U2862(p1_u2862), .P1_U2861(p1_u2861), .P1_U2860(p1_u2860), .P1_U2859(p1_u2859), .P1_U2858(p1_u2858), .P1_U2857(p1_u2857), .P1_U2856(p1_u2856), .P1_U2855(p1_u2855), .P1_U2854(p1_u2854), .P1_U2853(p1_u2853), .P1_U2852(p1_u2852), .P1_U2851(p1_u2851), .P1_U2850(p1_u2850), .P1_U2849(p1_u2849), .P1_U2848(p1_u2848), .P1_U2847(p1_u2847), .P1_U2846(p1_u2846), .P1_U2845(p1_u2845), .P1_U2844(p1_u2844), .P1_U2843(p1_u2843), .P1_U2842(p1_u2842), .P1_U2841(p1_u2841), .P1_U2840(p1_u2840), .P1_U2839(p1_u2839), .P1_U2838(p1_u2838), .P1_U2837(p1_u2837), .P1_U2836(p1_u2836), .P1_U2835(p1_u2835), .P1_U2834(p1_u2834), .P1_U2833(p1_u2833), .P1_U2832(p1_u2832), .P1_U2831(p1_u2831), .P1_U2830(p1_u2830), .P1_U2829(p1_u2829), .P1_U2828(p1_u2828), .P1_U2827(p1_u2827), .P1_U2826(p1_u2826), .P1_U2825(p1_u2825), .P1_U2824(p1_u2824), .P1_U2823(p1_u2823), .P1_U2822(p1_u2822), .P1_U2821(p1_u2821), .P1_U2820(p1_u2820), .P1_U2819(p1_u2819), .P1_U2818(p1_u2818), .P1_U2817(p1_u2817), .P1_U2816(p1_u2816), .P1_U2815(p1_u2815), .P1_U2814(p1_u2814), .P1_U2813(p1_u2813), .P1_U2812(p1_u2812), .P1_U2811(p1_u2811), .P1_U2810(p1_u2810), .P1_U2809(p1_u2809), .P1_U2808(p1_u2808), .P1_U3481(p1_u3481), .P1_U2807(p1_u2807), .P1_U3482(p1_u3482), .P1_U3483(p1_u3483), .P1_U2806(p1_u2806), .P1_U3484(p1_u3484), .P1_U2805(p1_u2805), .P1_U3485(p1_u3485), .P1_U2804(p1_u2804), .P1_U3486(p1_u3486), .P1_U2803(p1_u2803), .P1_U2802(p1_u2802), .P1_U3487(p1_u3487), .P1_U2801(p1_u2801));

integer i=0;
always @ (posedge clk) begin
	vec = input_vec_mem[i];
	$monitor(vec);
	i = i + 1;

end

always @ (negedge clk)begin
	$fdisplay ( fh_w, p3_datao_reg_31_, p3_datao_reg_30_, p3_datao_reg_29_, p3_datao_reg_28_, p3_datao_reg_27_, p3_datao_reg_26_, p3_datao_reg_25_, p3_datao_reg_24_, p3_datao_reg_23_, p3_datao_reg_22_, p3_datao_reg_21_, p3_datao_reg_20_, p3_datao_reg_19_, p3_datao_reg_18_, p3_datao_reg_17_, p3_datao_reg_16_, p3_datao_reg_15_, p3_datao_reg_14_, p3_datao_reg_13_, p3_datao_reg_12_, p3_datao_reg_11_, p3_datao_reg_10_, p3_datao_reg_9_, p3_datao_reg_8_, p3_datao_reg_7_, p3_datao_reg_6_, p3_datao_reg_5_, p3_datao_reg_4_, p3_datao_reg_3_, p3_datao_reg_2_, p3_datao_reg_1_, p3_datao_reg_0_, p1_address_reg_29_, p1_address_reg_28_, p1_address_reg_27_, p1_address_reg_26_, p1_address_reg_25_, p1_address_reg_24_, p1_address_reg_23_, p1_address_reg_22_, p1_address_reg_21_, p1_address_reg_20_, p1_address_reg_19_, p1_address_reg_18_, p1_address_reg_17_, p1_address_reg_16_, p1_address_reg_15_, p1_address_reg_14_, p1_address_reg_13_, p1_address_reg_12_, p1_address_reg_11_, p1_address_reg_10_, p1_address_reg_9_, p1_address_reg_8_, p1_address_reg_7_, p1_address_reg_6_, p1_address_reg_5_, p1_address_reg_4_, p1_address_reg_3_, p1_address_reg_2_, p1_address_reg_1_, p1_address_reg_0_, u355, u356, u357, u358, u359, u360, u361, u362, u363, u364, u366, u367, u368, u369, u370, u371, u372, u373, u374, u375, u347, u348, u349, u350, u351, u352, u353, u354, u365, u376, p3_w_r_n_reg, p3_d_c_n_reg, p3_m_io_n_reg, p1_ads_n_reg, p3_ads_n_reg, u247, u246, u245, u244, u243, u242, u241, u240, u239, u238, u237, u236, u235, u234, u233, u232, u231, u230, u229, u228, u227, u226, u225, u224, u223, u222, u221, u220, u219, u218, u217, u216, u251, u252, u253, u254, u255, u256, u257, u258, u259, u260, u261, u262, u263, u264, u265, u266, u267, u268, u269, u270, u271, u272, u273, u274, u275, u276, u277, u278, u279, u280, u281, u282, u212, u215, u213, u214, p3_u3274, p3_u3275, p3_u3276, p3_u3277, p3_u3061, p3_u3060, p3_u3059, p3_u3058, p3_u3057, p3_u3056, p3_u3055, p3_u3054, p3_u3053, p3_u3052, p3_u3051, p3_u3050, p3_u3049, p3_u3048, p3_u3047, p3_u3046, p3_u3045, p3_u3044, p3_u3043, p3_u3042, p3_u3041, p3_u3040, p3_u3039, p3_u3038, p3_u3037, p3_u3036, p3_u3035, p3_u3034, p3_u3033, p3_u3032, p3_u3031, p3_u3030, p3_u3029, p3_u3280, p3_u3281, p3_u3028, p3_u3027, p3_u3026, p3_u3025, p3_u3024, p3_u3023, p3_u3022, p3_u3021, p3_u3020, p3_u3019, p3_u3018, p3_u3017, p3_u3016, p3_u3015, p3_u3014, p3_u3013, p3_u3012, p3_u3011, p3_u3010, p3_u3009, p3_u3008, p3_u3007, p3_u3006, p3_u3005, p3_u3004, p3_u3003, p3_u3002, p3_u3001, p3_u3000, p3_u2999, p3_u3282, p3_u2998, p3_u2997, p3_u2996, p3_u2995, p3_u2994, p3_u2993, p3_u2992, p3_u2991, p3_u2990, p3_u2989, p3_u2988, p3_u2987, p3_u2986, p3_u2985, p3_u2984, p3_u2983, p3_u2982, p3_u2981, p3_u2980, p3_u2979, p3_u2978, p3_u2977, p3_u2976, p3_u2975, p3_u2974, p3_u2973, p3_u2972, p3_u2971, p3_u2970, p3_u2969, p3_u2968, p3_u2967, p3_u2966, p3_u2965, p3_u2964, p3_u2963, p3_u2962, p3_u2961, p3_u2960, p3_u2959, p3_u2958, p3_u2957, p3_u2956, p3_u2955, p3_u2954, p3_u2953, p3_u2952, p3_u2951, p3_u2950, p3_u2949, p3_u2948, p3_u2947, p3_u2946, p3_u2945, p3_u2944, p3_u2943, p3_u2942, p3_u2941, p3_u2940, p3_u2939, p3_u2938, p3_u2937, p3_u2936, p3_u2935, p3_u2934, p3_u2933, p3_u2932, p3_u2931, p3_u2930, p3_u2929, p3_u2928, p3_u2927, p3_u2926, p3_u2925, p3_u2924, p3_u2923, p3_u2922, p3_u2921, p3_u2920, p3_u2919, p3_u2918, p3_u2917, p3_u2916, p3_u2915, p3_u2914, p3_u2913, p3_u2912, p3_u2911, p3_u2910, p3_u2909, p3_u2908, p3_u2907, p3_u2906, p3_u2905, p3_u2904, p3_u2903, p3_u2902, p3_u2901, p3_u2900, p3_u2899, p3_u2898, p3_u2897, p3_u2896, p3_u2895, p3_u2894, p3_u2893, p3_u2892, p3_u2891, p3_u2890, p3_u2889, p3_u2888, p3_u2887, p3_u2886, p3_u2885, p3_u2884, p3_u2883, p3_u2882, p3_u2881, p3_u2880, p3_u2879, p3_u2878, p3_u2877, p3_u2876, p3_u2875, p3_u2874, p3_u2873, p3_u2872, p3_u2871, p3_u2870, p3_u2869, p3_u2868, p3_u3284, p3_u3285, p3_u3288, p3_u3289, p3_u3290, p3_u2867, p3_u2866, p3_u2865, p3_u2864, p3_u2863, p3_u2862, p3_u2861, p3_u2860, p3_u2859, p3_u2858, p3_u2857, p3_u2856, p3_u2855, p3_u2854, p3_u2853, p3_u2852, p3_u2851, p3_u2850, p3_u2849, p3_u2848, p3_u2847, p3_u2846, p3_u2845, p3_u2844, p3_u2843, p3_u2842, p3_u2841, p3_u2840, p3_u2839, p3_u2838, p3_u2837, p3_u2836, p3_u2835, p3_u2834, p3_u2833, p3_u2832, p3_u2831, p3_u2830, p3_u2829, p3_u2828, p3_u2827, p3_u2826, p3_u2825, p3_u2824, p3_u2823, p3_u2822, p3_u2821, p3_u2820, p3_u2819, p3_u2818, p3_u2817, p3_u2816, p3_u2815, p3_u2814, p3_u2813, p3_u2812, p3_u2811, p3_u2810, p3_u2809, p3_u2808, p3_u2807, p3_u2806, p3_u2805, p3_u2804, p3_u2803, p3_u2802, p3_u2801, p3_u2800, p3_u2799, p3_u2798, p3_u2797, p3_u2796, p3_u2795, p3_u2794, p3_u2793, p3_u2792, p3_u2791, p3_u2790, p3_u2789, p3_u2788, p3_u2787, p3_u2786, p3_u2785, p3_u2784, p3_u2783, p3_u2782, p3_u2781, p3_u2780, p3_u2779, p3_u2778, p3_u2777, p3_u2776, p3_u2775, p3_u2774, p3_u2773, p3_u2772, p3_u2771, p3_u2770, p3_u2769, p3_u2768, p3_u2767, p3_u2766, p3_u2765, p3_u2764, p3_u2763, p3_u2762, p3_u2761, p3_u2760, p3_u2759, p3_u2758, p3_u2757, p3_u2756, p3_u2755, p3_u2754, p3_u2753, p3_u2752, p3_u2751, p3_u2750, p3_u2749, p3_u2748, p3_u2747, p3_u2746, p3_u2745, p3_u2744, p3_u2743, p3_u2742, p3_u2741, p3_u2740, p3_u2739, p3_u2738, p3_u2737, p3_u2736, p3_u2735, p3_u2734, p3_u2733, p3_u2732, p3_u2731, p3_u2730, p3_u2729, p3_u2728, p3_u2727, p3_u2726, p3_u2725, p3_u2724, p3_u2723, p3_u2722, p3_u2721, p3_u2720, p3_u2719, p3_u2718, p3_u2717, p3_u2716, p3_u2715, p3_u2714, p3_u2713, p3_u2712, p3_u2711, p3_u2710, p3_u2709, p3_u2708, p3_u2707, p3_u2706, p3_u2705, p3_u2704, p3_u2703, p3_u2702, p3_u2701, p3_u2700, p3_u2699, p3_u2698, p3_u2697, p3_u2696, p3_u2695, p3_u2694, p3_u2693, p3_u2692, p3_u2691, p3_u2690, p3_u2689, p3_u2688, p3_u2687, p3_u2686, p3_u2685, p3_u2684, p3_u2683, p3_u2682, p3_u2681, p3_u2680, p3_u2679, p3_u2678, p3_u2677, p3_u2676, p3_u2675, p3_u2674, p3_u2673, p3_u2672, p3_u2671, p3_u2670, p3_u2669, p3_u2668, p3_u2667, p3_u2666, p3_u2665, p3_u2664, p3_u2663, p3_u2662, p3_u2661, p3_u2660, p3_u2659, p3_u2658, p3_u2657, p3_u2656, p3_u2655, p3_u2654, p3_u2653, p3_u2652, p3_u2651, p3_u2650, p3_u2649, p3_u2648, p3_u2647, p3_u2646, p3_u2645, p3_u2644, p3_u2643, p3_u2642, p3_u2641, p3_u2640, p3_u2639, p3_u3292, p3_u2638, p3_u3293, p3_u3294, p3_u2637, p3_u3295, p3_u2636, p3_u3296, p3_u2635, p3_u3297, p3_u2634, p3_u2633, p3_u3298, p3_u3299, p2_u3585, p2_u3586, p2_u3587, p2_u3588, p2_u3241, p2_u3240, p2_u3239, p2_u3238, p2_u3237, p2_u3236, p2_u3235, p2_u3234, p2_u3233, p2_u3232, p2_u3231, p2_u3230, p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225, p2_u3224, p2_u3223, p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218, p2_u3217, p2_u3216, p2_u3215, p2_u3214, p2_u3213, p2_u3212, p2_u3211, p2_u3210, p2_u3209, p2_u3591, p2_u3592, p2_u3208, p2_u3207, p2_u3206, p2_u3205, p2_u3204, p2_u3203, p2_u3202, p2_u3201, p2_u3200, p2_u3199, p2_u3198, p2_u3197, p2_u3196, p2_u3195, p2_u3194, p2_u3193, p2_u3192, p2_u3191, p2_u3190, p2_u3189, p2_u3188, p2_u3187, p2_u3186, p2_u3185, p2_u3184, p2_u3183, p2_u3182, p2_u3181, p2_u3180, p2_u3179, p2_u3593, p2_u3178, p2_u3177, p2_u3176, p2_u3175, p2_u3174, p2_u3173, p2_u3172, p2_u3171, p2_u3170, p2_u3169, p2_u3168, p2_u3167, p2_u3166, p2_u3165, p2_u3164, p2_u3163, p2_u3162, p2_u3161, p2_u3160, p2_u3159, p2_u3158, p2_u3157, p2_u3156, p2_u3155, p2_u3154, p2_u3153, p2_u3152, p2_u3151, p2_u3150, p2_u3149, p2_u3148, p2_u3147, p2_u3146, p2_u3145, p2_u3144, p2_u3143, p2_u3142, p2_u3141, p2_u3140, p2_u3139, p2_u3138, p2_u3137, p2_u3136, p2_u3135, p2_u3134, p2_u3133, p2_u3132, p2_u3131, p2_u3130, p2_u3129, p2_u3128, p2_u3127, p2_u3126, p2_u3125, p2_u3124, p2_u3123, p2_u3122, p2_u3121, p2_u3120, p2_u3119, p2_u3118, p2_u3117, p2_u3116, p2_u3115, p2_u3114, p2_u3113, p2_u3112, p2_u3111, p2_u3110, p2_u3109, p2_u3108, p2_u3107, p2_u3106, p2_u3105, p2_u3104, p2_u3103, p2_u3102, p2_u3101, p2_u3100, p2_u3099, p2_u3098, p2_u3097, p2_u3096, p2_u3095, p2_u3094, p2_u3093, p2_u3092, p2_u3091, p2_u3090, p2_u3089, p2_u3088, p2_u3087, p2_u3086, p2_u3085, p2_u3084, p2_u3083, p2_u3082, p2_u3081, p2_u3080, p2_u3079, p2_u3078, p2_u3077, p2_u3076, p2_u3075, p2_u3074, p2_u3073, p2_u3072, p2_u3071, p2_u3070, p2_u3069, p2_u3068, p2_u3067, p2_u3066, p2_u3065, p2_u3064, p2_u3063, p2_u3062, p2_u3061, p2_u3060, p2_u3059, p2_u3058, p2_u3057, p2_u3056, p2_u3055, p2_u3054, p2_u3053, p2_u3052, p2_u3051, p2_u3050, p2_u3049, p2_u3048, p2_u3595, p2_u3596, p2_u3599, p2_u3600, p2_u3601, p2_u3047, p2_u3602, p2_u3603, p2_u3604, p2_u3605, p2_u3046, p2_u3045, p2_u3044, p2_u3043, p2_u3042, p2_u3041, p2_u3040, p2_u3039, p2_u3038, p2_u3037, p2_u3036, p2_u3035, p2_u3034, p2_u3033, p2_u3032, p2_u3031, p2_u3030, p2_u3029, p2_u3028, p2_u3027, p2_u3026, p2_u3025, p2_u3024, p2_u3023, p2_u3022, p2_u3021, p2_u3020, p2_u3019, p2_u3018, p2_u3017, p2_u3016, p2_u3015, p2_u3014, p2_u3013, p2_u3012, p2_u3011, p2_u3010, p2_u3009, p2_u3008, p2_u3007, p2_u3006, p2_u3005, p2_u3004, p2_u3003, p2_u3002, p2_u3001, p2_u3000, p2_u2999, p2_u2998, p2_u2997, p2_u2996, p2_u2995, p2_u2994, p2_u2993, p2_u2992, p2_u2991, p2_u2990, p2_u2989, p2_u2988, p2_u2987, p2_u2986, p2_u2985, p2_u2984, p2_u2983, p2_u2982, p2_u2981, p2_u2980, p2_u2979, p2_u2978, p2_u2977, p2_u2976, p2_u2975, p2_u2974, p2_u2973, p2_u2972, p2_u2971, p2_u2970, p2_u2969, p2_u2968, p2_u2967, p2_u2966, p2_u2965, p2_u2964, p2_u2963, p2_u2962, p2_u2961, p2_u2960, p2_u2959, p2_u2958, p2_u2957, p2_u2956, p2_u2955, p2_u2954, p2_u2953, p2_u2952, p2_u2951, p2_u2950, p2_u2949, p2_u2948, p2_u2947, p2_u2946, p2_u2945, p2_u2944, p2_u2943, p2_u2942, p2_u2941, p2_u2940, p2_u2939, p2_u2938, p2_u2937, p2_u2936, p2_u2935, p2_u2934, p2_u2933, p2_u2932, p2_u2931, p2_u2930, p2_u2929, p2_u2928, p2_u2927, p2_u2926, p2_u2925, p2_u2924, p2_u2923, p2_u2922, p2_u2921, p2_u2920, p2_u2919, p2_u2918, p2_u2917, p2_u2916, p2_u2915, p2_u2914, p2_u2913, p2_u2912, p2_u2911, p2_u2910, p2_u2909, p2_u2908, p2_u2907, p2_u2906, p2_u2905, p2_u2904, p2_u2903, p2_u2902, p2_u2901, p2_u2900, p2_u2899, p2_u2898, p2_u2897, p2_u2896, p2_u2895, p2_u2894, p2_u2893, p2_u2892, p2_u2891, p2_u2890, p2_u2889, p2_u2888, p2_u2887, p2_u2886, p2_u2885, p2_u2884, p2_u2883, p2_u2882, p2_u2881, p2_u2880, p2_u2879, p2_u2878, p2_u2877, p2_u2876, p2_u2875, p2_u2874, p2_u2873, p2_u2872, p2_u2871, p2_u2870, p2_u2869, p2_u2868, p2_u2867, p2_u2866, p2_u2865, p2_u2864, p2_u2863, p2_u2862, p2_u2861, p2_u2860, p2_u2859, p2_u2858, p2_u2857, p2_u2856, p2_u2855, p2_u2854, p2_u2853, p2_u2852, p2_u2851, p2_u2850, p2_u2849, p2_u2848, p2_u2847, p2_u2846, p2_u2845, p2_u2844, p2_u2843, p2_u2842, p2_u2841, p2_u2840, p2_u2839, p2_u2838, p2_u2837, p2_u2836, p2_u2835, p2_u2834, p2_u2833, p2_u2832, p2_u2831, p2_u2830, p2_u2829, p2_u2828, p2_u2827, p2_u2826, p2_u2825, p2_u2824, p2_u2823, p2_u2822, p2_u2821, p2_u2820, p2_u3608, p2_u2819, p2_u3609, p2_u2818, p2_u3610, p2_u2817, p2_u3611, p2_u2816, p2_u2815, p2_u3612, p2_u2814, p1_u3458, p1_u3459, p1_u3460, p1_u3461, p1_u3226, p1_u3225, p1_u3224, p1_u3223, p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218, p1_u3217, p1_u3216, p1_u3215, p1_u3214, p1_u3213, p1_u3212, p1_u3211, p1_u3210, p1_u3209, p1_u3208, p1_u3207, p1_u3206, p1_u3205, p1_u3204, p1_u3203, p1_u3202, p1_u3201, p1_u3200, p1_u3199, p1_u3198, p1_u3197, p1_u3196, p1_u3195, p1_u3194, p1_u3464, p1_u3465, p1_u3193, p1_u3192, p1_u3191, p1_u3190, p1_u3189, p1_u3188, p1_u3187, p1_u3186, p1_u3185, p1_u3184, p1_u3183, p1_u3182, p1_u3181, p1_u3180, p1_u3179, p1_u3178, p1_u3177, p1_u3176, p1_u3175, p1_u3174, p1_u3173, p1_u3172, p1_u3171, p1_u3170, p1_u3169, p1_u3168, p1_u3167, p1_u3166, p1_u3165, p1_u3164, p1_u3466, p1_u3163, p1_u3162, p1_u3161, p1_u3160, p1_u3159, p1_u3158, p1_u3157, p1_u3156, p1_u3155, p1_u3154, p1_u3153, p1_u3152, p1_u3151, p1_u3150, p1_u3149, p1_u3148, p1_u3147, p1_u3146, p1_u3145, p1_u3144, p1_u3143, p1_u3142, p1_u3141, p1_u3140, p1_u3139, p1_u3138, p1_u3137, p1_u3136, p1_u3135, p1_u3134, p1_u3133, p1_u3132, p1_u3131, p1_u3130, p1_u3129, p1_u3128, p1_u3127, p1_u3126, p1_u3125, p1_u3124, p1_u3123, p1_u3122, p1_u3121, p1_u3120, p1_u3119, p1_u3118, p1_u3117, p1_u3116, p1_u3115, p1_u3114, p1_u3113, p1_u3112, p1_u3111, p1_u3110, p1_u3109, p1_u3108, p1_u3107, p1_u3106, p1_u3105, p1_u3104, p1_u3103, p1_u3102, p1_u3101, p1_u3100, p1_u3099, p1_u3098, p1_u3097, p1_u3096, p1_u3095, p1_u3094, p1_u3093, p1_u3092, p1_u3091, p1_u3090, p1_u3089, p1_u3088, p1_u3087, p1_u3086, p1_u3085, p1_u3084, p1_u3083, p1_u3082, p1_u3081, p1_u3080, p1_u3079, p1_u3078, p1_u3077, p1_u3076, p1_u3075, p1_u3074, p1_u3073, p1_u3072, p1_u3071, p1_u3070, p1_u3069, p1_u3068, p1_u3067, p1_u3066, p1_u3065, p1_u3064, p1_u3063, p1_u3062, p1_u3061, p1_u3060, p1_u3059, p1_u3058, p1_u3057, p1_u3056, p1_u3055, p1_u3054, p1_u3053, p1_u3052, p1_u3051, p1_u3050, p1_u3049, p1_u3048, p1_u3047, p1_u3046, p1_u3045, p1_u3044, p1_u3043, p1_u3042, p1_u3041, p1_u3040, p1_u3039, p1_u3038, p1_u3037, p1_u3036, p1_u3035, p1_u3034, p1_u3033, p1_u3468, p1_u3469, p1_u3472, p1_u3473, p1_u3474, p1_u3032, p1_u3475, p1_u3476, p1_u3477, p1_u3478, p1_u3031, p1_u3030, p1_u3029, p1_u3028, p1_u3027, p1_u3026, p1_u3025, p1_u3024, p1_u3023, p1_u3022, p1_u3021, p1_u3020, p1_u3019, p1_u3018, p1_u3017, p1_u3016, p1_u3015, p1_u3014, p1_u3013, p1_u3012, p1_u3011, p1_u3010, p1_u3009, p1_u3008, p1_u3007, p1_u3006, p1_u3005, p1_u3004, p1_u3003, p1_u3002, p1_u3001, p1_u3000, p1_u2999, p1_u2998, p1_u2997, p1_u2996, p1_u2995, p1_u2994, p1_u2993, p1_u2992, p1_u2991, p1_u2990, p1_u2989, p1_u2988, p1_u2987, p1_u2986, p1_u2985, p1_u2984, p1_u2983, p1_u2982, p1_u2981, p1_u2980, p1_u2979, p1_u2978, p1_u2977, p1_u2976, p1_u2975, p1_u2974, p1_u2973, p1_u2972, p1_u2971, p1_u2970, p1_u2969, p1_u2968, p1_u2967, p1_u2966, p1_u2965, p1_u2964, p1_u2963, p1_u2962, p1_u2961, p1_u2960, p1_u2959, p1_u2958, p1_u2957, p1_u2956, p1_u2955, p1_u2954, p1_u2953, p1_u2952, p1_u2951, p1_u2950, p1_u2949, p1_u2948, p1_u2947, p1_u2946, p1_u2945, p1_u2944, p1_u2943, p1_u2942, p1_u2941, p1_u2940, p1_u2939, p1_u2938, p1_u2937, p1_u2936, p1_u2935, p1_u2934, p1_u2933, p1_u2932, p1_u2931, p1_u2930, p1_u2929, p1_u2928, p1_u2927, p1_u2926, p1_u2925, p1_u2924, p1_u2923, p1_u2922, p1_u2921, p1_u2920, p1_u2919, p1_u2918, p1_u2917, p1_u2916, p1_u2915, p1_u2914, p1_u2913, p1_u2912, p1_u2911, p1_u2910, p1_u2909, p1_u2908, p1_u2907, p1_u2906, p1_u2905, p1_u2904, p1_u2903, p1_u2902, p1_u2901, p1_u2900, p1_u2899, p1_u2898, p1_u2897, p1_u2896, p1_u2895, p1_u2894, p1_u2893, p1_u2892, p1_u2891, p1_u2890, p1_u2889, p1_u2888, p1_u2887, p1_u2886, p1_u2885, p1_u2884, p1_u2883, p1_u2882, p1_u2881, p1_u2880, p1_u2879, p1_u2878, p1_u2877, p1_u2876, p1_u2875, p1_u2874, p1_u2873, p1_u2872, p1_u2871, p1_u2870, p1_u2869, p1_u2868, p1_u2867, p1_u2866, p1_u2865, p1_u2864, p1_u2863, p1_u2862, p1_u2861, p1_u2860, p1_u2859, p1_u2858, p1_u2857, p1_u2856, p1_u2855, p1_u2854, p1_u2853, p1_u2852, p1_u2851, p1_u2850, p1_u2849, p1_u2848, p1_u2847, p1_u2846, p1_u2845, p1_u2844, p1_u2843, p1_u2842, p1_u2841, p1_u2840, p1_u2839, p1_u2838, p1_u2837, p1_u2836, p1_u2835, p1_u2834, p1_u2833, p1_u2832, p1_u2831, p1_u2830, p1_u2829, p1_u2828, p1_u2827, p1_u2826, p1_u2825, p1_u2824, p1_u2823, p1_u2822, p1_u2821, p1_u2820, p1_u2819, p1_u2818, p1_u2817, p1_u2816, p1_u2815, p1_u2814, p1_u2813, p1_u2812, p1_u2811, p1_u2810, p1_u2809, p1_u2808, p1_u3481, p1_u2807, p1_u3482, p1_u3483, p1_u2806, p1_u3484, p1_u2805, p1_u3485, p1_u2804, p1_u3486, p1_u2803, p1_u2802, p1_u3487, p1_u2801);
	if(i == vec_length)begin
		$finish;
	end
end

integer fh_w;
initial begin
	fh_w = $fopen(`out_file, "w");
end
 
initial begin
	//$fsdbDumpfile("SET.fsdb");
	//$fsdbDumpvars;
	//$fsdbDumpMDA;
	$dumpfile("test_result.vcd");
    $dumpvars;

end
endmodule
