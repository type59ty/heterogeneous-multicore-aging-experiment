// Verilog
// c1908
// Ninputs 33
// Noutputs 25
// NtotalGates 880
// NOT1 277
// NAND2 347
// BUFF1 162
// AND2 30
// AND3 12
// NAND4 2
// NAND3 1
// NAND8 3
// AND4 2
// NAND5 24
// AND5 16
// AND8 3
// NOR2 1

module c1908d (N11,N14,N17,N110,N113,N116,N119,N122,N125,N128,
              N131,N134,N137,N140,N143,N146,N149,N153,N156,N160,
              N163,N166,N169,N172,N176,N179,N182,N185,N188,N191,
              N194,N199,N1104,N12753,N12754,N12755,N12756,N12762,N12767,N12768,
              N12779,N12780,N12781,N12782,N12783,N12784,N12785,N12786,N12787,N12811,
              N12886,N12887,N12888,N12889,N12890,N12891,N12892,N12899,
              N21,N24,N27,N210,N213,N216,N219,N222,N225,N228,
              N231,N234,N237,N240,N243,N246,N249,N253,N256,N260,
              N263,N266,N269,N272,N276,N279,N282,N285,N288,N291,
              N294,N299,N2104,N22753,N22754,N22755,N22756,N22762,N22767,N22768,
              N22779,N22780,N22781,N22782,N22783,N22784,N22785,N22786,N22787,N22811,
              N22886,N22887,N22888,N22889,N22890,N22891,N22892,N22899);

input N11,N14,N17,N110,N113,N116,N119,N122,N125,N128,
      N131,N134,N137,N140,N143,N146,N149,N153,N156,N160,
      N163,N166,N169,N172,N176,N179,N182,N185,N188,N191,
      N194,N199,N1104,
      N21,N24,N27,N210,N213,N216,N219,N222,N225,N228,
      N231,N234,N237,N240,N243,N246,N249,N253,N256,N260,
      N263,N266,N269,N272,N276,N279,N282,N285,N288,N291,
      N294,N299,N2104;

output N12753,N12754,N12755,N12756,N12762,N12767,N12768,N12779,N12780,N12781,
       N12782,N12783,N12784,N12785,N12786,N12787,N12811,N12886,N12887,N12888,
       N12889,N12890,N12891,N12892,N12899,
       N22753,N22754,N22755,N22756,N22762,N22767,N22768,N22779,N22780,N22781,
       N22782,N22783,N22784,N22785,N22786,N22787,N22811,N22886,N22887,N22888,
       N22889,N22890,N22891,N22892,N22899;

wire N1190,N1194,N1197,N1201,N1206,N1209,N1212,N1216,N1220,N1225,
     N1229,N1232,N1235,N1239,N1243,N1247,N1251,N1252,N1253,N1256,
     N1257,N1260,N1263,N1266,N1269,N1272,N1275,N1276,N1277,N1280,
     N1283,N1290,N1297,N1300,N1303,N1306,N1313,N1316,N1319,N1326,
     N1331,N1338,N1343,N1346,N1349,N1352,N1355,N1358,N1361,N1364,
     N1367,N1370,N1373,N1376,N1379,N1382,N1385,N1388,N1534,N1535,
     N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,
     N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,
     N1556,N1559,N1562,N1565,N1568,N1571,N1574,N1577,N1580,N1583,
     N1586,N1589,N1592,N1595,N1598,N1601,N1602,N1603,N1608,N1612,
     N1616,N1619,N1622,N1625,N1628,N1631,N1634,N1637,N1640,N1643,
     N1646,N1649,N1652,N1655,N1658,N1661,N1664,N1667,N1670,N1673,
     N1676,N1679,N1682,N1685,N1688,N1691,N1694,N1697,N1700,N1703,
     N1706,N1709,N1712,N1715,N1718,N1721,N1724,N1727,N1730,N1733,
     N1736,N1739,N1742,N1745,N1748,N1751,N1886,N1887,N1888,N1889,
     N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,
     N1903,N1907,N1910,N1913,N1914,N1915,N1916,N1917,N1918,N1919,
     N1920,N1921,N1922,N1923,N1926,N1935,N1938,N1939,N1942,N1943,
     N1946,N1947,N1950,N1951,N1954,N1955,N1958,N1959,N1962,N1965,
     N1968,N1969,N1972,N1973,N1976,N1977,N1980,N1981,N1984,N1985,
     N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1997,N1998,N11001,
     N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11009,N11010,N11013,
     N11016,N11019,N11022,N11025,N11028,N11031,N11034,N11037,N11040,N11043,
     N11046,N11049,N11054,N11055,N11063,N11064,N11067,N11068,N11119,N11120,
     N11121,N11122,N11128,N11129,N11130,N11131,N11132,N11133,N11148,N11149,
     N11150,N11151,N11152,N11153,N11154,N11155,N11156,N11157,N11158,N11159,
     N11160,N11161,N11162,N11163,N11164,N11167,N11168,N11171,N11188,N11205,
     N11206,N11207,N11208,N11209,N11210,N11211,N11212,N11213,N11214,N11215,
     N11216,N11217,N11218,N11219,N11220,N11221,N11222,N11223,N11224,N11225,
     N11226,N11227,N11228,N11229,N11230,N11231,N11232,N11235,N11238,N11239,
     N11240,N11241,N11242,N11243,N11246,N11249,N11252,N11255,N11258,N11261,
     N11264,N11267,N11309,N11310,N11311,N11312,N11313,N11314,N11315,N11316,
     N11317,N11318,N11319,N11322,N11327,N11328,N11334,N11344,N11345,N11346,
     N11348,N11349,N11350,N11351,N11352,N11355,N11358,N11361,N11364,N11367,
     N11370,N11373,N11376,N11379,N11383,N11386,N11387,N11388,N11389,N11390,
     N11393,N11396,N11397,N11398,N11399,N11409,N11412,N11413,N11416,N11419,
     N11433,N11434,N11438,N11439,N11440,N11443,N11444,N11445,N11446,N11447,
     N11448,N11451,N11452,N11453,N11454,N11455,N11456,N11457,N11458,N11459,
     N11460,N11461,N11462,N11463,N11464,N11468,N11469,N11470,N11471,N11472,
     N11475,N11476,N11478,N11481,N11484,N11487,N11488,N11489,N11490,N11491,
     N11492,N11493,N11494,N11495,N11496,N11498,N11499,N11500,N11501,N11504,
     N11510,N11513,N11514,N11517,N11520,N11521,N11522,N11526,N11527,N11528,
     N11529,N11530,N11531,N11532,N11534,N11537,N11540,N11546,N11554,N11557,
     N11561,N11567,N11568,N11569,N11571,N11576,N11588,N11591,N11593,N11594,
     N11595,N11596,N11600,N11603,N11606,N11609,N11612,N11615,N11620,N11623,
     N11635,N11636,N11638,N11639,N11640,N11643,N11647,N11651,N11658,N11661,
     N11664,N11671,N11672,N11675,N11677,N11678,N11679,N11680,N11681,N11682,
     N11683,N11685,N11688,N11697,N11701,N11706,N11707,N11708,N11709,N11710,
     N11711,N11712,N11713,N11714,N11717,N11720,N11721,N11723,N11727,N11728,
     N11730,N11731,N11734,N11740,N11741,N11742,N11746,N11747,N11748,N11751,
     N11759,N11761,N11762,N11763,N11764,N11768,N11769,N11772,N11773,N11774,
     N11777,N11783,N11784,N11785,N11786,N11787,N11788,N11791,N11792,N11795,
     N11796,N11798,N11801,N11802,N11807,N11808,N11809,N11810,N11812,N11815,
     N11818,N11821,N11822,N11823,N11824,N11825,N11826,N11827,N11830,N11837,
     N11838,N11841,N11848,N11849,N11850,N11852,N11855,N11856,N11857,N11858,
     N11864,N11865,N11866,N11869,N11872,N11875,N11878,N11879,N11882,N11883,
     N11884,N11885,N11889,N11895,N11896,N11897,N11898,N11902,N11910,N11911,
     N11912,N11913,N11915,N11919,N11920,N11921,N11922,N11923,N11924,N11927,
     N11930,N11933,N11936,N11937,N11938,N11941,N11942,N11944,N11947,N11950,
     N11953,N11958,N11961,N11965,N11968,N11975,N11976,N11977,N11978,N11979,
     N11980,N11985,N11987,N11999,N12000,N12002,N12003,N12004,N12005,N12006,
     N12007,N12008,N12009,N12012,N12013,N12014,N12015,N12016,N12018,N12019,
     N12020,N12021,N12022,N12023,N12024,N12025,N12026,N12027,N12030,N12033,
     N12036,N12037,N12038,N12039,N12040,N12041,N12042,N12047,N12052,N12055,
     N12060,N12061,N12062,N12067,N12068,N12071,N12076,N12077,N12078,N12081,
     N12086,N12089,N12104,N12119,N12129,N12143,N12148,N12151,N12196,N12199,
     N12202,N12205,N12214,N12215,N12216,N12217,N12222,N12223,N12224,N12225,
     N12226,N12227,N12228,N12229,N12230,N12231,N12232,N12233,N12234,N12235,
     N12236,N12237,N12240,N12241,N12244,N12245,N12250,N12253,N12256,N12257,
     N12260,N12263,N12266,N12269,N12272,N12279,N12286,N12297,N12315,N12326,
     N12340,N12353,N12361,N12375,N12384,N12385,N12386,N12426,N12427,N12537,
     N12540,N12543,N12546,N12549,N12552,N12555,N12558,N12561,N12564,N12567,
     N12570,N12573,N12576,N12594,N12597,N12600,N12603,N12606,N12611,N12614,
     N12617,N12620,N12627,N12628,N12629,N12630,N12631,N12632,N12633,N12634,
     N12639,N12642,N12645,N12648,N12651,N12655,N12658,N12661,N12664,N12669,
     N12670,N12671,N12672,N12673,N12674,N12675,N12676,N12682,N12683,N12688,
     N12689,N12690,N12691,N12710,N12720,N12721,N12722,N12723,N12724,N12725,
     N12726,N12727,N12728,N12729,N12730,N12731,N12732,N12733,N12734,N12735,
     N12736,N12737,N12738,N12739,N12740,N12741,N12742,N12743,N12744,N12745,
     N12746,N12747,N12750,N12757,N12758,N12759,N12760,N12761,N12763,N12764,
     N12765,N12766,N12773,N12776,N12788,N12789,N12800,N12807,N12808,N12809,
     N12810,N12812,N12815,N12818,N12821,N12824,N12827,N12828,N12829,N12843,
     N12846,N12850,N12851,N12852,N12853,N12854,N12857,N12858,N12859,N12860,
     N12861,N12862,N12863,N12866,N12867,N12868,N12869,N12870,N12871,N12872,
     N12873,N12874,N12875,N12876,N12877,N12878,N12879,N12880,N12881,N12882,
     N12883,N12895,N12896,N12897,N12898,

     N2190,N2194,N2197,N2201,N2206,N2209,N2212,N2216,N2220,N2225,
     N2229,N2232,N2235,N2239,N2243,N2247,N2251,N2252,N2253,N2256,
     N2257,N2260,N2263,N2266,N2269,N2272,N2275,N2276,N2277,N2280,
     N2283,N2290,N2297,N2300,N2303,N2306,N2313,N2316,N2319,N2326,
     N2331,N2338,N2343,N2346,N2349,N2352,N2355,N2358,N2361,N2364,
     N2367,N2370,N2373,N2376,N2379,N2382,N2385,N2388,N2534,N2535,
     N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,N2545,
     N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,
     N2556,N2559,N2562,N2565,N2568,N2571,N2574,N2577,N2580,N2583,
     N2586,N2589,N2592,N2595,N2598,N2601,N2602,N2603,N2608,N2612,
     N2616,N2619,N2622,N2625,N2628,N2631,N2634,N2637,N2640,N2643,
     N2646,N2649,N2652,N2655,N2658,N2661,N2664,N2667,N2670,N2673,
     N2676,N2679,N2682,N2685,N2688,N2691,N2694,N2697,N2700,N2703,
     N2706,N2709,N2712,N2715,N2718,N2721,N2724,N2727,N2730,N2733,
     N2736,N2739,N2742,N2745,N2748,N2751,N2886,N2887,N2888,N2889,
     N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,
     N2903,N2907,N2910,N2913,N2914,N2915,N2916,N2917,N2918,N2919,
     N2920,N2921,N2922,N2923,N2926,N2935,N2938,N2939,N2942,N2943,
     N2946,N2947,N2950,N2951,N2954,N2955,N2958,N2959,N2962,N2965,
     N2968,N2969,N2972,N2973,N2976,N2977,N2980,N2981,N2984,N2985,
     N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2997,N2998,N21001,
     N21002,N21003,N21004,N21005,N21006,N21007,N21008,N21009,N21010,N21013,
     N21016,N21019,N21022,N21025,N21028,N21031,N21034,N21037,N21040,N21043,
     N21046,N21049,N21054,N21055,N21063,N21064,N21067,N21068,N21119,N21120,
     N21121,N21122,N21128,N21129,N21130,N21131,N21132,N21133,N21148,N21149,
     N21150,N21151,N21152,N21153,N21154,N21155,N21156,N21157,N21158,N21159,
     N21160,N21161,N21162,N21163,N21164,N21167,N21168,N21171,N21188,N21205,
     N21206,N21207,N21208,N21209,N21210,N21211,N21212,N21213,N21214,N21215,
     N21216,N21217,N21218,N21219,N21220,N21221,N21222,N21223,N21224,N21225,
     N21226,N21227,N21228,N21229,N21230,N21231,N21232,N21235,N21238,N21239,
     N21240,N21241,N21242,N21243,N21246,N21249,N21252,N21255,N21258,N21261,
     N21264,N21267,N21309,N21310,N21311,N21312,N21313,N21314,N21315,N21316,
     N21317,N21318,N21319,N21322,N21327,N21328,N21334,N21344,N21345,N21346,
     N21348,N21349,N21350,N21351,N21352,N21355,N21358,N21361,N21364,N21367,
     N21370,N21373,N21376,N21379,N21383,N21386,N21387,N21388,N21389,N21390,
     N21393,N21396,N21397,N21398,N21399,N21409,N21412,N21413,N21416,N21419,
     N21433,N21434,N21438,N21439,N21440,N21443,N21444,N21445,N21446,N21447,
     N21448,N21451,N21452,N21453,N21454,N21455,N21456,N21457,N21458,N21459,
     N21460,N21461,N21462,N21463,N21464,N21468,N21469,N21470,N21471,N21472,
     N21475,N21476,N21478,N21481,N21484,N21487,N21488,N21489,N21490,N21491,
     N21492,N21493,N21494,N21495,N21496,N21498,N21499,N21500,N21501,N21504,
     N21510,N21513,N21514,N21517,N21520,N21521,N21522,N21526,N21527,N21528,
     N21529,N21530,N21531,N21532,N21534,N21537,N21540,N21546,N21554,N21557,
     N21561,N21567,N21568,N21569,N21571,N21576,N21588,N21591,N21593,N21594,
     N21595,N21596,N21600,N21603,N21606,N21609,N21612,N21615,N21620,N21623,
     N21635,N21636,N21638,N21639,N21640,N21643,N21647,N21651,N21658,N21661,
     N21664,N21671,N21672,N21675,N21677,N21678,N21679,N21680,N21681,N21682,
     N21683,N21685,N21688,N21697,N21701,N21706,N21707,N21708,N21709,N21710,
     N21711,N21712,N21713,N21714,N21717,N21720,N21721,N21723,N21727,N21728,
     N21730,N21731,N21734,N21740,N21741,N21742,N21746,N21747,N21748,N21751,
     N21759,N21761,N21762,N21763,N21764,N21768,N21769,N21772,N21773,N21774,
     N21777,N21783,N21784,N21785,N21786,N21787,N21788,N21791,N21792,N21795,
     N21796,N21798,N21801,N21802,N21807,N21808,N21809,N21810,N21812,N21815,
     N21818,N21821,N21822,N21823,N21824,N21825,N21826,N21827,N21830,N21837,
     N21838,N21841,N21848,N21849,N21850,N21852,N21855,N21856,N21857,N21858,
     N21864,N21865,N21866,N21869,N21872,N21875,N21878,N21879,N21882,N21883,
     N21884,N21885,N21889,N21895,N21896,N21897,N21898,N21902,N21910,N21911,
     N21912,N21913,N21915,N21919,N21920,N21921,N21922,N21923,N21924,N21927,
     N21930,N21933,N21936,N21937,N21938,N21941,N21942,N21944,N21947,N21950,
     N21953,N21958,N21961,N21965,N21968,N21975,N21976,N21977,N21978,N21979,
     N21980,N21985,N21987,N21999,N22000,N22002,N22003,N22004,N22005,N22006,
     N22007,N22008,N22009,N22012,N22013,N22014,N22015,N22016,N22018,N22019,
     N22020,N22021,N22022,N22023,N22024,N22025,N22026,N22027,N22030,N22033,
     N22036,N22037,N22038,N22039,N22040,N22041,N22042,N22047,N22052,N22055,
     N22060,N22061,N22062,N22067,N22068,N22071,N22076,N22077,N22078,N22081,
     N22086,N22089,N22104,N22119,N22129,N22143,N22148,N22151,N22196,N22199,
     N22202,N22205,N22214,N22215,N22216,N22217,N22222,N22223,N22224,N22225,
     N22226,N22227,N22228,N22229,N22230,N22231,N22232,N22233,N22234,N22235,
     N22236,N22237,N22240,N22241,N22244,N22245,N22250,N22253,N22256,N22257,
     N22260,N22263,N22266,N22269,N22272,N22279,N22286,N22297,N22315,N22326,
     N22340,N22353,N22361,N22375,N22384,N22385,N22386,N22426,N22427,N22537,
     N22540,N22543,N22546,N22549,N22552,N22555,N22558,N22561,N22564,N22567,
     N22570,N22573,N22576,N22594,N22597,N22600,N22603,N22606,N22611,N22614,
     N22617,N22620,N22627,N22628,N22629,N22630,N22631,N22632,N22633,N22634,
     N22639,N22642,N22645,N22648,N22651,N22655,N22658,N22661,N22664,N22669,
     N22670,N22671,N22672,N22673,N22674,N22675,N22676,N22682,N22683,N22688,
     N22689,N22690,N22691,N22710,N22720,N22721,N22722,N22723,N22724,N22725,
     N22726,N22727,N22728,N22729,N22730,N22731,N22732,N22733,N22734,N22735,
     N22736,N22737,N22738,N22739,N22740,N22741,N22742,N22743,N22744,N22745,
     N22746,N22747,N22750,N22757,N22758,N22759,N22760,N22761,N22763,N22764,
     N22765,N22766,N22773,N22776,N22788,N22789,N22800,N22807,N22808,N22809,
     N22810,N22812,N22815,N22818,N22821,N22824,N22827,N22828,N22829,N22843,
     N22846,N22850,N22851,N22852,N22853,N22854,N22857,N22858,N22859,N22860,
     N22861,N22862,N22863,N22866,N22867,N22868,N22869,N22870,N22871,N22872,
     N22873,N22874,N22875,N22876,N22877,N22878,N22879,N22880,N22881,N22882,
     N22883,N22895,N22896,N22897,N22898;


not NOT1_11 (N1190, N11);
not NOT1_12 (N1194, N14);
not NOT1_13 (N1197, N17);
not NOT1_14 (N1201, N110);
not NOT1_15 (N1206, N113);
not NOT1_16 (N1209, N116);
not NOT1_17 (N1212, N119);
not NOT1_18 (N1216, N122);
not NOT1_19 (N1220, N125);
not NOT1_110 (N1225, N128);
not NOT1_111 (N1229, N131);
not NOT1_112 (N1232, N134);
not NOT1_113 (N1235, N137);
not NOT1_114 (N1239, N140);
not NOT1_115 (N1243, N143);
not NOT1_116 (N1247, N146);
nand NAND2_117 (N1251, N163, N188);
nand NAND2_118 (N1252, N166, N191);
not NOT1_119 (N1253, N172);
not NOT1_120 (N1256, N172);
buf BUFF1_121 (N1257, N169);
buf BUFF1_122 (N1260, N169);
not NOT1_123 (N1263, N176);
not NOT1_124 (N1266, N179);
not NOT1_125 (N1269, N182);
not NOT1_126 (N1272, N185);
not NOT1_127 (N1275, N1104);
not NOT1_128 (N1276, N1104);
not NOT1_129 (N1277, N188);
not NOT1_130 (N1280, N191);
buf BUFF1_131 (N1283, N194);
not NOT1_132 (N1290, N194);
buf BUFF1_133 (N1297, N194);
not NOT1_134 (N1300, N194);
buf BUFF1_135 (N1303, N199);
not NOT1_136 (N1306, N199);
not NOT1_137 (N1313, N199);
buf BUFF1_138 (N1316, N1104);
not NOT1_139 (N1319, N1104);
buf BUFF1_140 (N1326, N1104);
buf BUFF1_141 (N1331, N1104);
not NOT1_142 (N1338, N1104);
buf BUFF1_143 (N1343, N11);
buf BUFF1_144 (N1346, N14);
buf BUFF1_145 (N1349, N17);
buf BUFF1_146 (N1352, N110);
buf BUFF1_147 (N1355, N113);
buf BUFF1_148 (N1358, N116);
buf BUFF1_149 (N1361, N119);
buf BUFF1_150 (N1364, N122);
buf BUFF1_151 (N1367, N125);
buf BUFF1_152 (N1370, N128);
buf BUFF1_153 (N1373, N131);
buf BUFF1_154 (N1376, N134);
buf BUFF1_155 (N1379, N137);
buf BUFF1_156 (N1382, N140);
buf BUFF1_157 (N1385, N143);
buf BUFF1_158 (N1388, N146);
not NOT1_159 (N1534, N1343);
not NOT1_160 (N1535, N1346);
not NOT1_161 (N1536, N1349);
not NOT1_162 (N1537, N1352);
not NOT1_163 (N1538, N1355);
not NOT1_164 (N1539, N1358);
not NOT1_165 (N1540, N1361);
not NOT1_166 (N1541, N1364);
not NOT1_167 (N1542, N1367);
not NOT1_168 (N1543, N1370);
not NOT1_169 (N1544, N1373);
not NOT1_170 (N1545, N1376);
not NOT1_171 (N1546, N1379);
not NOT1_172 (N1547, N1382);
not NOT1_173 (N1548, N1385);
not NOT1_174 (N1549, N1388);
nand NAND2_175 (N1550, N1306, N1331);
nand NAND2_176 (N1551, N1306, N1331);
nand NAND2_177 (N1552, N1306, N1331);
nand NAND2_178 (N1553, N1306, N1331);
nand NAND2_179 (N1554, N1306, N1331);
nand NAND2_180 (N1555, N1306, N1331);
buf BUFF1_181 (N1556, N1190);
buf BUFF1_182 (N1559, N1194);
buf BUFF1_183 (N1562, N1206);
buf BUFF1_184 (N1565, N1209);
buf BUFF1_185 (N1568, N1225);
buf BUFF1_186 (N1571, N1243);
and AND2_187 (N1574, N163, N1319);
buf BUFF1_188 (N1577, N1220);
buf BUFF1_189 (N1580, N1229);
buf BUFF1_190 (N1583, N1232);
and AND2_191 (N1586, N166, N1319);
buf BUFF1_192 (N1589, N1239);
and AND3_193 (N1592, N149, N1253, N1319);
buf BUFF1_194 (N1595, N1247);
buf BUFF1_195 (N1598, N1239);
nand NAND2_196 (N1601, N1326, N1277);
nand NAND2_197 (N1602, N1326, N1280);
nand NAND2_198 (N1603, N1260, N172);
nand NAND2_199 (N1608, N1260, N1300);
nand NAND2_1100 (N1612, N1256, N1300);
buf BUFF1_1101 (N1616, N1201);
buf BUFF1_1102 (N1619, N1216);
buf BUFF1_1103 (N1622, N1220);
buf BUFF1_1104 (N1625, N1239);
buf BUFF1_1105 (N1628, N1190);
buf BUFF1_1106 (N1631, N1190);
buf BUFF1_1107 (N1634, N1194);
buf BUFF1_1108 (N1637, N1229);
buf BUFF1_1109 (N1640, N1197);
and AND3_1110 (N1643, N156, N1257, N1319);
buf BUFF1_1111 (N1646, N1232);
buf BUFF1_1112 (N1649, N1201);
buf BUFF1_1113 (N1652, N1235);
and AND3_1114 (N1655, N160, N1257, N1319);
buf BUFF1_1115 (N1658, N1263);
buf BUFF1_1116 (N1661, N1263);
buf BUFF1_1117 (N1664, N1266);
buf BUFF1_1118 (N1667, N1266);
buf BUFF1_1119 (N1670, N1269);
buf BUFF1_1120 (N1673, N1269);
buf BUFF1_1121 (N1676, N1272);
buf BUFF1_1122 (N1679, N1272);
and AND2_1123 (N1682, N1251, N1316);
and AND2_1124 (N1685, N1252, N1316);
buf BUFF1_1125 (N1688, N1197);
buf BUFF1_1126 (N1691, N1197);
buf BUFF1_1127 (N1694, N1212);
buf BUFF1_1128 (N1697, N1212);
buf BUFF1_1129 (N1700, N1247);
buf BUFF1_1130 (N1703, N1247);
buf BUFF1_1131 (N1706, N1235);
buf BUFF1_1132 (N1709, N1235);
buf BUFF1_1133 (N1712, N1201);
buf BUFF1_1134 (N1715, N1201);
buf BUFF1_1135 (N1718, N1206);
buf BUFF1_1136 (N1721, N1216);
and AND3_1137 (N1724, N153, N1253, N1319);
buf BUFF1_1138 (N1727, N1243);
buf BUFF1_1139 (N1730, N1220);
buf BUFF1_1140 (N1733, N1220);
buf BUFF1_1141 (N1736, N1209);
buf BUFF1_1142 (N1739, N1216);
buf BUFF1_1143 (N1742, N1225);
buf BUFF1_1144 (N1745, N1243);
buf BUFF1_1145 (N1748, N1212);
buf BUFF1_1146 (N1751, N1225);
not NOT1_1147 (N1886, N1682);
not NOT1_1148 (N1887, N1685);
not NOT1_1149 (N1888, N1616);
not NOT1_1150 (N1889, N1619);
not NOT1_1151 (N1890, N1622);
not NOT1_1152 (N1891, N1625);
not NOT1_1153 (N1892, N1631);
not NOT1_1154 (N1893, N1643);
not NOT1_1155 (N1894, N1649);
not NOT1_1156 (N1895, N1652);
not NOT1_1157 (N1896, N1655);
and AND2_1158 (N1897, N149, N1612);
and AND2_1159 (N1898, N156, N1608);
nand NAND2_1160 (N1899, N153, N1612);
nand NAND2_1161 (N1903, N160, N1608);
nand NAND2_1162 (N1907, N149, N1612);
nand NAND2_1163 (N1910, N156, N1608);
not NOT1_1164 (N1913, N1661);
not NOT1_1165 (N1914, N1658);
not NOT1_1166 (N1915, N1667);
not NOT1_1167 (N1916, N1664);
not NOT1_1168 (N1917, N1673);
not NOT1_1169 (N1918, N1670);
not NOT1_1170 (N1919, N1679);
not NOT1_1171 (N1920, N1676);
nand NAND4_1172 (N1921, N1277, N1297, N1326, N1603);
nand NAND4_1173 (N1922, N1280, N1297, N1326, N1603);
nand NAND3_1174 (N1923, N1303, N1338, N1603);
and AND3_1175 (N1926, N1303, N1338, N1603);
buf BUFF1_1176 (N1935, N1556);
not NOT1_1177 (N1938, N1688);
buf BUFF1_1178 (N1939, N1556);
not NOT1_1179 (N1942, N1691);
buf BUFF1_1180 (N1943, N1562);
not NOT1_1181 (N1946, N1694);
buf BUFF1_1182 (N1947, N1562);
not NOT1_1183 (N1950, N1697);
buf BUFF1_1184 (N1951, N1568);
not NOT1_1185 (N1954, N1700);
buf BUFF1_1186 (N1955, N1568);
not NOT1_1187 (N1958, N1703);
buf BUFF1_1188 (N1959, N1574);
buf BUFF1_1189 (N1962, N1574);
buf BUFF1_1190 (N1965, N1580);
not NOT1_1191 (N1968, N1706);
buf BUFF1_1192 (N1969, N1580);
not NOT1_1193 (N1972, N1709);
buf BUFF1_1194 (N1973, N1586);
not NOT1_1195 (N1976, N1712);
buf BUFF1_1196 (N1977, N1586);
not NOT1_1197 (N1980, N1715);
buf BUFF1_1198 (N1981, N1592);
not NOT1_1199 (N1984, N1628);
buf BUFF1_1200 (N1985, N1592);
not NOT1_1201 (N1988, N1718);
not NOT1_1202 (N1989, N1721);
not NOT1_1203 (N1990, N1634);
not NOT1_1204 (N1991, N1724);
not NOT1_1205 (N1992, N1727);
not NOT1_1206 (N1993, N1637);
buf BUFF1_1207 (N1994, N1595);
not NOT1_1208 (N1997, N1730);
buf BUFF1_1209 (N1998, N1595);
not NOT1_1210 (N11001, N1733);
not NOT1_1211 (N11002, N1736);
not NOT1_1212 (N11003, N1739);
not NOT1_1213 (N11004, N1640);
not NOT1_1214 (N11005, N1742);
not NOT1_1215 (N11006, N1745);
not NOT1_1216 (N11007, N1646);
not NOT1_1217 (N11008, N1748);
not NOT1_1218 (N11009, N1751);
buf BUFF1_1219 (N11010, N1559);
buf BUFF1_1220 (N11013, N1559);
buf BUFF1_1221 (N11016, N1565);
buf BUFF1_1222 (N11019, N1565);
buf BUFF1_1223 (N11022, N1571);
buf BUFF1_1224 (N11025, N1571);
buf BUFF1_1225 (N11028, N1577);
buf BUFF1_1226 (N11031, N1577);
buf BUFF1_1227 (N11034, N1583);
buf BUFF1_1228 (N11037, N1583);
buf BUFF1_1229 (N11040, N1589);
buf BUFF1_1230 (N11043, N1589);
buf BUFF1_1231 (N11046, N1598);
buf BUFF1_1232 (N11049, N1598);
nand NAND2_1233 (N11054, N1619, N1888);
nand NAND2_1234 (N11055, N1616, N1889);
nand NAND2_1235 (N11063, N1625, N1890);
nand NAND2_1236 (N11064, N1622, N1891);
nand NAND2_1237 (N11067, N1655, N1895);
nand NAND2_1238 (N11068, N1652, N1896);
nand NAND2_1239 (N11119, N1721, N1988);
nand NAND2_1240 (N11120, N1718, N1989);
nand NAND2_1241 (N11121, N1727, N1991);
nand NAND2_1242 (N11122, N1724, N1992);
nand NAND2_1243 (N11128, N1739, N11002);
nand NAND2_1244 (N11129, N1736, N11003);
nand NAND2_1245 (N11130, N1745, N11005);
nand NAND2_1246 (N11131, N1742, N11006);
nand NAND2_1247 (N11132, N1751, N11008);
nand NAND2_1248 (N11133, N1748, N11009);
not NOT1_1249 (N11148, N1939);
not NOT1_1250 (N11149, N1935);
nand NAND2_1251 (N11150, N11054, N11055);
not NOT1_1252 (N11151, N1943);
not NOT1_1253 (N11152, N1947);
not NOT1_1254 (N11153, N1955);
not NOT1_1255 (N11154, N1951);
not NOT1_1256 (N11155, N1962);
not NOT1_1257 (N11156, N1969);
not NOT1_1258 (N11157, N1977);
nand NAND2_1259 (N11158, N11063, N11064);
not NOT1_1260 (N11159, N1985);
nand NAND2_1261 (N11160, N1985, N1892);
not NOT1_1262 (N11161, N1998);
nand NAND2_1263 (N11162, N11067, N11068);
not NOT1_1264 (N11163, N1899);
buf BUFF1_1265 (N11164, N1899);
not NOT1_1266 (N11167, N1903);
buf BUFF1_1267 (N11168, N1903);
nand NAND2_1268 (N11171, N1921, N1923);
nand NAND2_1269 (N11188, N1922, N1923);
not NOT1_1270 (N11205, N11010);
nand NAND2_1271 (N11206, N11010, N1938);
not NOT1_1272 (N11207, N11013);
nand NAND2_1273 (N11208, N11013, N1942);
not NOT1_1274 (N11209, N11016);
nand NAND2_1275 (N11210, N11016, N1946);
not NOT1_1276 (N11211, N11019);
nand NAND2_1277 (N11212, N11019, N1950);
not NOT1_1278 (N11213, N11022);
nand NAND2_1279 (N11214, N11022, N1954);
not NOT1_1280 (N11215, N11025);
nand NAND2_1281 (N11216, N11025, N1958);
not NOT1_1282 (N11217, N11028);
not NOT1_1283 (N11218, N1959);
not NOT1_1284 (N11219, N11031);
not NOT1_1285 (N11220, N11034);
nand NAND2_1286 (N11221, N11034, N1968);
not NOT1_1287 (N11222, N1965);
not NOT1_1288 (N11223, N11037);
nand NAND2_1289 (N11224, N11037, N1972);
not NOT1_1290 (N11225, N11040);
nand NAND2_1291 (N11226, N11040, N1976);
not NOT1_1292 (N11227, N1973);
not NOT1_1293 (N11228, N11043);
nand NAND2_1294 (N11229, N11043, N1980);
not NOT1_1295 (N11230, N1981);
nand NAND2_1296 (N11231, N1981, N1984);
nand NAND2_1297 (N11232, N11119, N11120);
nand NAND2_1298 (N11235, N11121, N11122);
not NOT1_1299 (N11238, N11046);
nand NAND2_1300 (N11239, N11046, N1997);
not NOT1_1301 (N11240, N1994);
not NOT1_1302 (N11241, N11049);
nand NAND2_1303 (N11242, N11049, N11001);
nand NAND2_1304 (N11243, N11128, N11129);
nand NAND2_1305 (N11246, N11130, N11131);
nand NAND2_1306 (N11249, N11132, N11133);
buf BUFF1_1307 (N11252, N1907);
buf BUFF1_1308 (N11255, N1907);
buf BUFF1_1309 (N11258, N1910);
buf BUFF1_1310 (N11261, N1910);
not NOT1_1311 (N11264, N11150);
nand NAND2_1312 (N11267, N1631, N11159);
nand NAND2_1313 (N11309, N1688, N11205);
nand NAND2_1314 (N11310, N1691, N11207);
nand NAND2_1315 (N11311, N1694, N11209);
nand NAND2_1316 (N11312, N1697, N11211);
nand NAND2_1317 (N11313, N1700, N11213);
nand NAND2_1318 (N11314, N1703, N11215);
nand NAND2_1319 (N11315, N1706, N11220);
nand NAND2_1320 (N11316, N1709, N11223);
nand NAND2_1321 (N11317, N1712, N11225);
nand NAND2_1322 (N11318, N1715, N11228);
not NOT1_1323 (N11319, N11158);
nand NAND2_1324 (N11322, N1628, N11230);
nand NAND2_1325 (N11327, N1730, N11238);
nand NAND2_1326 (N11328, N1733, N11241);
not NOT1_1327 (N11334, N11162);
nand NAND2_1328 (N11344, N11267, N11160);
nand NAND2_1329 (N11345, N11249, N1894);
not NOT1_1330 (N11346, N11249);
not NOT1_1331 (N11348, N11255);
not NOT1_1332 (N11349, N11252);
not NOT1_1333 (N11350, N11261);
not NOT1_1334 (N11351, N11258);
nand NAND2_1335 (N11352, N11309, N11206);
nand NAND2_1336 (N11355, N11310, N11208);
nand NAND2_1337 (N11358, N11311, N11210);
nand NAND2_1338 (N11361, N11312, N11212);
nand NAND2_1339 (N11364, N11313, N11214);
nand NAND2_1340 (N11367, N11314, N11216);
nand NAND2_1341 (N11370, N11315, N11221);
nand NAND2_1342 (N11373, N11316, N11224);
nand NAND2_1343 (N11376, N11317, N11226);
nand NAND2_1344 (N11379, N11318, N11229);
nand NAND2_1345 (N11383, N11322, N11231);
not NOT1_1346 (N11386, N11232);
nand NAND2_1347 (N11387, N11232, N1990);
not NOT1_1348 (N11388, N11235);
nand NAND2_1349 (N11389, N11235, N1993);
nand NAND2_1350 (N11390, N11327, N11239);
nand NAND2_1351 (N11393, N11328, N11242);
not NOT1_1352 (N11396, N11243);
nand NAND2_1353 (N11397, N11243, N11004);
not NOT1_1354 (N11398, N11246);
nand NAND2_1355 (N11399, N11246, N11007);
not NOT1_1356 (N11409, N11319);
nand NAND2_1357 (N11412, N1649, N11346);
not NOT1_1358 (N11413, N11334);
buf BUFF1_1359 (N11416, N11264);
buf BUFF1_1360 (N11419, N11264);
nand NAND2_1361 (N11433, N1634, N11386);
nand NAND2_1362 (N11434, N1637, N11388);
nand NAND2_1363 (N11438, N1640, N11396);
nand NAND2_1364 (N11439, N1646, N11398);
not NOT1_1365 (N11440, N11344);
nand NAND2_1366 (N11443, N11355, N11148);
not NOT1_1367 (N11444, N11355);
nand NAND2_1368 (N11445, N11352, N11149);
not NOT1_1369 (N11446, N11352);
nand NAND2_1370 (N11447, N11358, N11151);
not NOT1_1371 (N11448, N11358);
nand NAND2_1372 (N11451, N11361, N11152);
not NOT1_1373 (N11452, N11361);
nand NAND2_1374 (N11453, N11367, N11153);
not NOT1_1375 (N11454, N11367);
nand NAND2_1376 (N11455, N11364, N11154);
not NOT1_1377 (N11456, N11364);
nand NAND2_1378 (N11457, N11373, N11156);
not NOT1_1379 (N11458, N11373);
nand NAND2_1380 (N11459, N11379, N11157);
not NOT1_1381 (N11460, N11379);
not NOT1_1382 (N11461, N11383);
nand NAND2_1383 (N11462, N11393, N11161);
not NOT1_1384 (N11463, N11393);
nand NAND2_1385 (N11464, N11345, N11412);
not NOT1_1386 (N11468, N11370);
nand NAND2_1387 (N11469, N11370, N11222);
not NOT1_1388 (N11470, N11376);
nand NAND2_1389 (N11471, N11376, N11227);
nand NAND2_1390 (N11472, N11387, N11433);
not NOT1_1391 (N11475, N11390);
nand NAND2_1392 (N11476, N11390, N11240);
nand NAND2_1393 (N11478, N11389, N11434);
nand NAND2_1394 (N11481, N11399, N11439);
nand NAND2_1395 (N11484, N11397, N11438);
nand NAND2_1396 (N11487, N1939, N11444);
nand NAND2_1397 (N11488, N1935, N11446);
nand NAND2_1398 (N11489, N1943, N11448);
not NOT1_1399 (N11490, N11419);
not NOT1_1400 (N11491, N11416);
nand NAND2_1401 (N11492, N1947, N11452);
nand NAND2_1402 (N11493, N1955, N11454);
nand NAND2_1403 (N11494, N1951, N11456);
nand NAND2_1404 (N11495, N1969, N11458);
nand NAND2_1405 (N11496, N1977, N11460);
nand NAND2_1406 (N11498, N1998, N11463);
not NOT1_1407 (N11499, N11440);
nand NAND2_1408 (N11500, N1965, N11468);
nand NAND2_1409 (N11501, N1973, N11470);
nand NAND2_1410 (N11504, N1994, N11475);
not NOT1_1411 (N11510, N11464);
nand NAND2_1412 (N11513, N11443, N11487);
nand NAND2_1413 (N11514, N11445, N11488);
nand NAND2_1414 (N11517, N11447, N11489);
nand NAND2_1415 (N11520, N11451, N11492);
nand NAND2_1416 (N11521, N11453, N11493);
nand NAND2_1417 (N11522, N11455, N11494);
nand NAND2_1418 (N11526, N11457, N11495);
nand NAND2_1419 (N11527, N11459, N11496);
not NOT1_1420 (N11528, N11472);
nand NAND2_1421 (N11529, N11462, N11498);
not NOT1_1422 (N11530, N11478);
not NOT1_1423 (N11531, N11481);
not NOT1_1424 (N11532, N11484);
nand NAND2_1425 (N11534, N11471, N11501);
nand NAND2_1426 (N11537, N11469, N11500);
nand NAND2_1427 (N11540, N11476, N11504);
not NOT1_1428 (N11546, N11513);
not NOT1_1429 (N11554, N11521);
not NOT1_1430 (N11557, N11526);
not NOT1_1431 (N11561, N11520);
nand NAND2_1432 (N11567, N11484, N11531);
nand NAND2_1433 (N11568, N11481, N11532);
not NOT1_1434 (N11569, N11510);
not NOT1_1435 (N11571, N11527);
not NOT1_1436 (N11576, N11529);
buf BUFF1_1437 (N11588, N11522);
not NOT1_1438 (N11591, N11534);
not NOT1_1439 (N11593, N11537);
nand NAND2_1440 (N11594, N11540, N11530);
not NOT1_1441 (N11595, N11540);
nand NAND2_1442 (N11596, N11567, N11568);
buf BUFF1_1443 (N11600, N11517);
buf BUFF1_1444 (N11603, N11517);
buf BUFF1_1445 (N11606, N11522);
buf BUFF1_1446 (N11609, N11522);
buf BUFF1_1447 (N11612, N11514);
buf BUFF1_1448 (N11615, N11514);
buf BUFF1_1449 (N11620, N11557);
buf BUFF1_1450 (N11623, N11554);
not NOT1_1451 (N11635, N11571);
nand NAND2_1452 (N11636, N11478, N11595);
nand NAND2_1453 (N11638, N11576, N11569);
not NOT1_1454 (N11639, N11576);
buf BUFF1_1455 (N11640, N11561);
buf BUFF1_1456 (N11643, N11561);
buf BUFF1_1457 (N11647, N11546);
buf BUFF1_1458 (N11651, N11546);
buf BUFF1_1459 (N11658, N11554);
buf BUFF1_1460 (N11661, N11557);
buf BUFF1_1461 (N11664, N11557);
nand NAND2_1462 (N11671, N11596, N1893);
not NOT1_1463 (N11672, N11596);
not NOT1_1464 (N11675, N11600);
not NOT1_1465 (N11677, N11603);
nand NAND2_1466 (N11678, N11606, N11217);
not NOT1_1467 (N11679, N11606);
nand NAND2_1468 (N11680, N11609, N11219);
not NOT1_1469 (N11681, N11609);
not NOT1_1470 (N11682, N11612);
not NOT1_1471 (N11683, N11615);
nand NAND2_1472 (N11685, N11594, N11636);
nand NAND2_1473 (N11688, N11510, N11639);
buf BUFF1_1474 (N11697, N11588);
buf BUFF1_1475 (N11701, N11588);
nand NAND2_1476 (N11706, N1643, N11672);
not NOT1_1477 (N11707, N11643);
nand NAND2_1478 (N11708, N11647, N11675);
not NOT1_1479 (N11709, N11647);
nand NAND2_1480 (N11710, N11651, N11677);
not NOT1_1481 (N11711, N11651);
nand NAND2_1482 (N11712, N11028, N11679);
nand NAND2_1483 (N11713, N11031, N11681);
buf BUFF1_1484 (N11714, N11620);
buf BUFF1_1485 (N11717, N11620);
nand NAND2_1486 (N11720, N11658, N11593);
not NOT1_1487 (N11721, N11658);
nand NAND2_1488 (N11723, N11638, N11688);
not NOT1_1489 (N11727, N11661);
not NOT1_1490 (N11728, N11640);
not NOT1_1491 (N11730, N11664);
buf BUFF1_1492 (N11731, N11623);
buf BUFF1_1493 (N11734, N11623);
nand NAND2_1494 (N11740, N11685, N11528);
not NOT1_1495 (N11741, N11685);
nand NAND2_1496 (N11742, N11671, N11706);
nand NAND2_1497 (N11746, N11600, N11709);
nand NAND2_1498 (N11747, N11603, N11711);
nand NAND2_1499 (N11748, N11678, N11712);
nand NAND2_1500 (N11751, N11680, N11713);
nand NAND2_1501 (N11759, N11537, N11721);
not NOT1_1502 (N11761, N11697);
nand NAND2_1503 (N11762, N11697, N11727);
not NOT1_1504 (N11763, N11701);
nand NAND2_1505 (N11764, N11701, N11730);
not NOT1_1506 (N11768, N11717);
nand NAND2_1507 (N11769, N11472, N11741);
nand NAND2_1508 (N11772, N11723, N11413);
not NOT1_1509 (N11773, N11723);
nand NAND2_1510 (N11774, N11708, N11746);
nand NAND2_1511 (N11777, N11710, N11747);
not NOT1_1512 (N11783, N11731);
nand NAND2_1513 (N11784, N11731, N11682);
not NOT1_1514 (N11785, N11714);
not NOT1_1515 (N11786, N11734);
nand NAND2_1516 (N11787, N11734, N11683);
nand NAND2_1517 (N11788, N11720, N11759);
nand NAND2_1518 (N11791, N11661, N11761);
nand NAND2_1519 (N11792, N11664, N11763);
nand NAND2_1520 (N11795, N11751, N11155);
not NOT1_1521 (N11796, N11751);
nand NAND2_1522 (N11798, N11740, N11769);
nand NAND2_1523 (N11801, N11334, N11773);
nand NAND2_1524 (N11802, N11742, N1290);
not NOT1_1525 (N11807, N11748);
nand NAND2_1526 (N11808, N11748, N11218);
nand NAND2_1527 (N11809, N11612, N11783);
nand NAND2_1528 (N11810, N11615, N11786);
nand NAND2_1529 (N11812, N11791, N11762);
nand NAND2_1530 (N11815, N11792, N11764);
buf BUFF1_1531 (N11818, N11742);
nand NAND2_1532 (N11821, N11777, N11490);
not NOT1_1533 (N11822, N11777);
nand NAND2_1534 (N11823, N11774, N11491);
not NOT1_1535 (N11824, N11774);
nand NAND2_1536 (N11825, N1962, N11796);
nand NAND2_1537 (N11826, N11788, N11409);
not NOT1_1538 (N11827, N11788);
nand NAND2_1539 (N11830, N11772, N11801);
nand NAND2_1540 (N11837, N1959, N11807);
nand NAND2_1541 (N11838, N11809, N11784);
nand NAND2_1542 (N11841, N11810, N11787);
nand NAND2_1543 (N11848, N11419, N11822);
nand NAND2_1544 (N11849, N11416, N11824);
nand NAND2_1545 (N11850, N11795, N11825);
nand NAND2_1546 (N11852, N11319, N11827);
nand NAND2_1547 (N11855, N11815, N11707);
not NOT1_1548 (N11856, N11815);
not NOT1_1549 (N11857, N11818);
nand NAND2_1550 (N11858, N11798, N1290);
not NOT1_1551 (N11864, N11812);
nand NAND2_1552 (N11865, N11812, N11728);
buf BUFF1_1553 (N11866, N11798);
buf BUFF1_1554 (N11869, N11802);
buf BUFF1_1555 (N11872, N11802);
nand NAND2_1556 (N11875, N11808, N11837);
nand NAND2_1557 (N11878, N11821, N11848);
nand NAND2_1558 (N11879, N11823, N11849);
nand NAND2_1559 (N11882, N11841, N11768);
not NOT1_1560 (N11883, N11841);
nand NAND2_1561 (N11884, N11826, N11852);
nand NAND2_1562 (N11885, N11643, N11856);
nand NAND2_1563 (N11889, N11830, N1290);
not NOT1_1564 (N11895, N11838);
nand NAND2_1565 (N11896, N11838, N11785);
nand NAND2_1566 (N11897, N11640, N11864);
not NOT1_1567 (N11898, N11850);
buf BUFF1_1568 (N11902, N11830);
not NOT1_1569 (N11910, N11878);
nand NAND2_1570 (N11911, N11717, N11883);
not NOT1_1571 (N11912, N11884);
nand NAND2_1572 (N11913, N11855, N11885);
not NOT1_1573 (N11915, N11866);
nand NAND2_1574 (N11919, N11872, N1919);
not NOT1_1575 (N11920, N11872);
nand NAND2_1576 (N11921, N11869, N1920);
not NOT1_1577 (N11922, N11869);
not NOT1_1578 (N11923, N11875);
nand NAND2_1579 (N11924, N11714, N11895);
buf BUFF1_1580 (N11927, N11858);
buf BUFF1_1581 (N11930, N11858);
nand NAND2_1582 (N11933, N11865, N11897);
nand NAND2_1583 (N11936, N11882, N11911);
not NOT1_1584 (N11937, N11898);
not NOT1_1585 (N11938, N11902);
nand NAND2_1586 (N11941, N1679, N11920);
nand NAND2_1587 (N11942, N1676, N11922);
buf BUFF1_1588 (N11944, N11879);
not NOT1_1589 (N11947, N11913);
buf BUFF1_1590 (N11950, N11889);
buf BUFF1_1591 (N11953, N11889);
buf BUFF1_1592 (N11958, N11879);
nand NAND2_1593 (N11961, N11896, N11924);
and AND2_1594 (N11965, N11910, N1601);
and AND2_1595 (N11968, N1602, N11912);
nand NAND2_1596 (N11975, N11930, N1917);
not NOT1_1597 (N11976, N11930);
nand NAND2_1598 (N11977, N11927, N1918);
not NOT1_1599 (N11978, N11927);
nand NAND2_1600 (N11979, N11919, N11941);
nand NAND2_1601 (N11980, N11921, N11942);
not NOT1_1602 (N11985, N11933);
not NOT1_1603 (N11987, N11936);
not NOT1_1604 (N11999, N11944);
nand NAND2_1605 (N12000, N11944, N11937);
not NOT1_1606 (N12002, N11947);
nand NAND2_1607 (N12003, N11947, N11499);
nand NAND2_1608 (N12004, N11953, N11350);
not NOT1_1609 (N12005, N11953);
nand NAND2_1610 (N12006, N11950, N11351);
not NOT1_1611 (N12007, N11950);
nand NAND2_1612 (N12008, N1673, N11976);
nand NAND2_1613 (N12009, N1670, N11978);
not NOT1_1614 (N12012, N11979);
not NOT1_1615 (N12013, N11958);
nand NAND2_1616 (N12014, N11958, N11923);
not NOT1_1617 (N12015, N11961);
nand NAND2_1618 (N12016, N11961, N11635);
not NOT1_1619 (N12018, N11965);
not NOT1_1620 (N12019, N11968);
nand NAND2_1621 (N12020, N11898, N11999);
not NOT1_1622 (N12021, N11987);
nand NAND2_1623 (N12022, N11987, N11591);
nand NAND2_1624 (N12023, N11440, N12002);
nand NAND2_1625 (N12024, N11261, N12005);
nand NAND2_1626 (N12025, N11258, N12007);
nand NAND2_1627 (N12026, N11975, N12008);
nand NAND2_1628 (N12027, N11977, N12009);
not NOT1_1629 (N12030, N11980);
buf BUFF1_1630 (N12033, N11980);
nand NAND2_1631 (N12036, N11875, N12013);
nand NAND2_1632 (N12037, N11571, N12015);
nand NAND2_1633 (N12038, N12020, N12000);
nand NAND2_1634 (N12039, N11534, N12021);
nand NAND2_1635 (N12040, N12023, N12003);
nand NAND2_1636 (N12041, N12004, N12024);
nand NAND2_1637 (N12042, N12006, N12025);
not NOT1_1638 (N12047, N12026);
nand NAND2_1639 (N12052, N12036, N12014);
nand NAND2_1640 (N12055, N12037, N12016);
not NOT1_1641 (N12060, N12038);
nand NAND2_1642 (N12061, N12039, N12022);
nand NAND2_1643 (N12062, N12040, N1290);
not NOT1_1644 (N12067, N12041);
not NOT1_1645 (N12068, N12027);
buf BUFF1_1646 (N12071, N12027);
not NOT1_1647 (N12076, N12052);
not NOT1_1648 (N12077, N12055);
nand NAND2_1649 (N12078, N12060, N1290);
nand NAND2_1650 (N12081, N12061, N1290);
not NOT1_1651 (N12086, N12042);
buf BUFF1_1652 (N12089, N12042);
and AND2_1653 (N12104, N12030, N12068);
and AND2_1654 (N12119, N12033, N12068);
and AND2_1655 (N12129, N12030, N12071);
and AND2_1656 (N12143, N12033, N12071);
buf BUFF1_1657 (N12148, N12062);
buf BUFF1_1658 (N12151, N12062);
buf BUFF1_1659 (N12196, N12078);
buf BUFF1_1660 (N12199, N12078);
buf BUFF1_1661 (N12202, N12081);
buf BUFF1_1662 (N12205, N12081);
nand NAND2_1663 (N12214, N12151, N1915);
not NOT1_1664 (N12215, N12151);
nand NAND2_1665 (N12216, N12148, N1916);
not NOT1_1666 (N12217, N12148);
nand NAND2_1667 (N12222, N12199, N11348);
not NOT1_1668 (N12223, N12199);
nand NAND2_1669 (N12224, N12196, N11349);
not NOT1_1670 (N12225, N12196);
nand NAND2_1671 (N12226, N12205, N1913);
not NOT1_1672 (N12227, N12205);
nand NAND2_1673 (N12228, N12202, N1914);
not NOT1_1674 (N12229, N12202);
nand NAND2_1675 (N12230, N1667, N12215);
nand NAND2_1676 (N12231, N1664, N12217);
nand NAND2_1677 (N12232, N11255, N12223);
nand NAND2_1678 (N12233, N11252, N12225);
nand NAND2_1679 (N12234, N1661, N12227);
nand NAND2_1680 (N12235, N1658, N12229);
nand NAND2_1681 (N12236, N12214, N12230);
nand NAND2_1682 (N12237, N12216, N12231);
nand NAND2_1683 (N12240, N12222, N12232);
nand NAND2_1684 (N12241, N12224, N12233);
nand NAND2_1685 (N12244, N12226, N12234);
nand NAND2_1686 (N12245, N12228, N12235);
not NOT1_1687 (N12250, N12236);
not NOT1_1688 (N12253, N12240);
not NOT1_1689 (N12256, N12244);
not NOT1_1690 (N12257, N12237);
buf BUFF1_1691 (N12260, N12237);
not NOT1_1692 (N12263, N12241);
and AND2_1693 (N12266, N11164, N12241);
not NOT1_1694 (N12269, N12245);
and AND2_1695 (N12272, N11168, N12245);
nand NAND8_1696 (N12279, N12067, N12012, N12047, N12250, N1899, N12256, N12253, N1903);
buf BUFF1_1697 (N12286, N12266);
buf BUFF1_1698 (N12297, N12266);
buf BUFF1_1699 (N12315, N12272);
buf BUFF1_1700 (N12326, N12272);
and AND2_1701 (N12340, N12086, N12257);
and AND2_1702 (N12353, N12089, N12257);
and AND2_1703 (N12361, N12086, N12260);
and AND2_1704 (N12375, N12089, N12260);
and AND4_1705 (N12384, N1338, N12279, N1313, N1313);
and AND2_1706 (N12385, N11163, N12263);
and AND2_1707 (N12386, N11164, N12263);
and AND2_1708 (N12426, N11167, N12269);
and AND2_1709 (N12427, N11168, N12269);
nand NAND5_1710 (N12537, N12286, N12315, N12361, N12104, N11171);
nand NAND5_1711 (N12540, N12286, N12315, N12340, N12129, N11171);
nand NAND5_1712 (N12543, N12286, N12315, N12340, N12119, N11171);
nand NAND5_1713 (N12546, N12286, N12315, N12353, N12104, N11171);
nand NAND5_1714 (N12549, N12297, N12315, N12375, N12119, N11188);
nand NAND5_1715 (N12552, N12297, N12326, N12361, N12143, N11188);
nand NAND5_1716 (N12555, N12297, N12326, N12375, N12129, N11188);
and AND5_1717 (N12558, N12286, N12315, N12361, N12104, N11171);
and AND5_1718 (N12561, N12286, N12315, N12340, N12129, N11171);
and AND5_1719 (N12564, N12286, N12315, N12340, N12119, N11171);
and AND5_1720 (N12567, N12286, N12315, N12353, N12104, N11171);
and AND5_1721 (N12570, N12297, N12315, N12375, N12119, N11188);
and AND5_1722 (N12573, N12297, N12326, N12361, N12143, N11188);
and AND5_1723 (N12576, N12297, N12326, N12375, N12129, N11188);
nand NAND5_1724 (N12594, N12286, N12427, N12361, N12129, N11171);
nand NAND5_1725 (N12597, N12297, N12427, N12361, N12119, N11171);
nand NAND5_1726 (N12600, N12297, N12427, N12375, N12104, N11171);
nand NAND5_1727 (N12603, N12297, N12427, N12340, N12143, N11171);
nand NAND5_1728 (N12606, N12297, N12427, N12353, N12129, N11188);
nand NAND5_1729 (N12611, N12386, N12326, N12361, N12129, N11188);
nand NAND5_1730 (N12614, N12386, N12326, N12361, N12119, N11188);
nand NAND5_1731 (N12617, N12386, N12326, N12375, N12104, N11188);
nand NAND5_1732 (N12620, N12386, N12326, N12353, N12129, N11188);
nand NAND5_1733 (N12627, N12297, N12427, N12340, N12104, N1926);
nand NAND5_1734 (N12628, N12386, N12326, N12340, N12104, N1926);
nand NAND5_1735 (N12629, N12386, N12427, N12361, N12104, N1926);
nand NAND5_1736 (N12630, N12386, N12427, N12340, N12129, N1926);
nand NAND5_1737 (N12631, N12386, N12427, N12340, N12119, N1926);
nand NAND5_1738 (N12632, N12386, N12427, N12353, N12104, N1926);
nand NAND5_1739 (N12633, N12386, N12426, N12340, N12104, N1926);
nand NAND5_1740 (N12634, N12385, N12427, N12340, N12104, N1926);
and AND5_1741 (N12639, N12286, N12427, N12361, N12129, N11171);
and AND5_1742 (N12642, N12297, N12427, N12361, N12119, N11171);
and AND5_1743 (N12645, N12297, N12427, N12375, N12104, N11171);
and AND5_1744 (N12648, N12297, N12427, N12340, N12143, N11171);
and AND5_1745 (N12651, N12297, N12427, N12353, N12129, N11188);
and AND5_1746 (N12655, N12386, N12326, N12361, N12129, N11188);
and AND5_1747 (N12658, N12386, N12326, N12361, N12119, N11188);
and AND5_1748 (N12661, N12386, N12326, N12375, N12104, N11188);
and AND5_1749 (N12664, N12386, N12326, N12353, N12129, N11188);
nand NAND2_1750 (N12669, N12558, N1534);
not NOT1_1751 (N12670, N12558);
nand NAND2_1752 (N12671, N12561, N1535);
not NOT1_1753 (N12672, N12561);
nand NAND2_1754 (N12673, N12564, N1536);
not NOT1_1755 (N12674, N12564);
nand NAND2_1756 (N12675, N12567, N1537);
not NOT1_1757 (N12676, N12567);
nand NAND2_1758 (N12682, N12570, N1543);
not NOT1_1759 (N12683, N12570);
nand NAND2_1760 (N12688, N12573, N1548);
not NOT1_1761 (N12689, N12573);
nand NAND2_1762 (N12690, N12576, N1549);
not NOT1_1763 (N12691, N12576);
and AND8_1764 (N12710, N12627, N12628, N12629, N12630, N12631, N12632, N12633, N12634);
nand NAND2_1765 (N12720, N1343, N12670);
nand NAND2_1766 (N12721, N1346, N12672);
nand NAND2_1767 (N12722, N1349, N12674);
nand NAND2_1768 (N12723, N1352, N12676);
nand NAND2_1769 (N12724, N12639, N1538);
not NOT1_1770 (N12725, N12639);
nand NAND2_1771 (N12726, N12642, N1539);
not NOT1_1772 (N12727, N12642);
nand NAND2_1773 (N12728, N12645, N1540);
not NOT1_1774 (N12729, N12645);
nand NAND2_1775 (N12730, N12648, N1541);
not NOT1_1776 (N12731, N12648);
nand NAND2_1777 (N12732, N12651, N1542);
not NOT1_1778 (N12733, N12651);
nand NAND2_1779 (N12734, N1370, N12683);
nand NAND2_1780 (N12735, N12655, N1544);
not NOT1_1781 (N12736, N12655);
nand NAND2_1782 (N12737, N12658, N1545);
not NOT1_1783 (N12738, N12658);
nand NAND2_1784 (N12739, N12661, N1546);
not NOT1_1785 (N12740, N12661);
nand NAND2_1786 (N12741, N12664, N1547);
not NOT1_1787 (N12742, N12664);
nand NAND2_1788 (N12743, N1385, N12689);
nand NAND2_1789 (N12744, N1388, N12691);
nand NAND8_1790 (N12745, N12537, N12540, N12543, N12546, N12594, N12597, N12600, N12603);
nand NAND8_1791 (N12746, N12606, N12549, N12611, N12614, N12617, N12620, N12552, N12555);
and AND8_1792 (N12747, N12537, N12540, N12543, N12546, N12594, N12597, N12600, N12603);
and AND8_1793 (N12750, N12606, N12549, N12611, N12614, N12617, N12620, N12552, N12555);
nand NAND2_1794 (N12753, N12669, N12720);
nand NAND2_1795 (N12754, N12671, N12721);
nand NAND2_1796 (N12755, N12673, N12722);
nand NAND2_1797 (N12756, N12675, N12723);
nand NAND2_1798 (N12757, N1355, N12725);
nand NAND2_1799 (N12758, N1358, N12727);
nand NAND2_1800 (N12759, N1361, N12729);
nand NAND2_1801 (N12760, N1364, N12731);
nand NAND2_1802 (N12761, N1367, N12733);
nand NAND2_1803 (N12762, N12682, N12734);
nand NAND2_1804 (N12763, N1373, N12736);
nand NAND2_1805 (N12764, N1376, N12738);
nand NAND2_1806 (N12765, N1379, N12740);
nand NAND2_1807 (N12766, N1382, N12742);
nand NAND2_1808 (N12767, N12688, N12743);
nand NAND2_1809 (N12768, N12690, N12744);
and AND2_1810 (N12773, N12745, N1275);
and AND2_1811 (N12776, N12746, N1276);
nand NAND2_1812 (N12779, N12724, N12757);
nand NAND2_1813 (N12780, N12726, N12758);
nand NAND2_1814 (N12781, N12728, N12759);
nand NAND2_1815 (N12782, N12730, N12760);
nand NAND2_1816 (N12783, N12732, N12761);
nand NAND2_1817 (N12784, N12735, N12763);
nand NAND2_1818 (N12785, N12737, N12764);
nand NAND2_1819 (N12786, N12739, N12765);
nand NAND2_1820 (N12787, N12741, N12766);
and AND3_1821 (N12788, N12747, N12750, N12710);
nand NAND2_1822 (N12789, N12747, N12750);
and AND4_1823 (N12800, N1338, N12279, N199, N12788);
nand NAND2_1824 (N12807, N12773, N12018);
not NOT1_1825 (N12808, N12773);
nand NAND2_1826 (N12809, N12776, N12019);
not NOT1_1827 (N12810, N12776);
nor N1OR2_1828 (N12811, N12384, N12800);
and AND3_1829 (N12812, N1897, N1283, N12789);
and AND3_1830 (N12815, N176, N1283, N12789);
and AND3_1831 (N12818, N182, N1283, N12789);
and AND3_1832 (N12821, N185, N1283, N12789);
and AND3_1833 (N12824, N1898, N1283, N12789);
nand NAND2_1834 (N12827, N11965, N12808);
nand NAND2_1835 (N12828, N11968, N12810);
and AND3_1836 (N12829, N179, N1283, N12789);
nand NAND2_1837 (N12843, N12807, N12827);
nand NAND2_1838 (N12846, N12809, N12828);
nand NAND2_1839 (N12850, N12812, N12076);
nand NAND2_1840 (N12851, N12815, N12077);
nand NAND2_1841 (N12852, N12818, N11915);
nand NAND2_1842 (N12853, N12821, N11857);
nand NAND2_1843 (N12854, N12824, N11938);
not NOT1_1844 (N12857, N12812);
not NOT1_1845 (N12858, N12815);
not NOT1_1846 (N12859, N12818);
not NOT1_1847 (N12860, N12821);
not NOT1_1848 (N12861, N12824);
not NOT1_1849 (N12862, N12829);
nand NAND2_1850 (N12863, N12829, N11985);
nand NAND2_1851 (N12866, N12052, N12857);
nand NAND2_1852 (N12867, N12055, N12858);
nand NAND2_1853 (N12868, N11866, N12859);
nand NAND2_1854 (N12869, N11818, N12860);
nand NAND2_1855 (N12870, N11902, N12861);
nand NAND2_1856 (N12871, N12843, N1886);
not NOT1_1857 (N12872, N12843);
nand NAND2_1858 (N12873, N12846, N1887);
not NOT1_1859 (N12874, N12846);
nand NAND2_1860 (N12875, N11933, N12862);
nand NAND2_1861 (N12876, N12866, N12850);
nand NAND2_1862 (N12877, N12867, N12851);
nand NAND2_1863 (N12878, N12868, N12852);
nand NAND2_1864 (N12879, N12869, N12853);
nand NAND2_1865 (N12880, N12870, N12854);
nand NAND2_1866 (N12881, N1682, N12872);
nand NAND2_1867 (N12882, N1685, N12874);
nand NAND2_1868 (N12883, N12875, N12863);
and AND2_1869 (N12886, N12876, N1550);
and AND2_1870 (N12887, N1551, N12877);
and AND2_1871 (N12888, N1553, N12878);
and AND2_1872 (N12889, N12879, N1554);
and AND2_1873 (N12890, N1555, N12880);
nand NAND2_1874 (N12891, N12871, N12881);
nand NAND2_1875 (N12892, N12873, N12882);
nand NAND2_1876 (N12895, N12883, N11461);
not NOT1_1877 (N12896, N12883);
nand NAND2_1878 (N12897, N11383, N12896);
nand NAND2_1879 (N12898, N12895, N12897);
and AND2_1880 (N12899, N12898, N1552);

not NOT1_21 (N2190, N21);
not NOT1_22 (N2194, N24);
not NOT1_23 (N2197, N27);
not NOT1_24 (N2201, N210);
not NOT1_25 (N2206, N213);
not NOT1_26 (N2209, N216);
not NOT1_27 (N2212, N219);
not NOT1_28 (N2216, N222);
not NOT1_29 (N2220, N225);
not NOT1_210 (N2225, N228);
not NOT1_211 (N2229, N231);
not NOT1_212 (N2232, N234);
not NOT1_213 (N2235, N237);
not NOT1_214 (N2239, N240);
not NOT1_215 (N2243, N243);
not NOT1_216 (N2247, N246);
nand NAND2_217 (N2251, N263, N288);
nand NAND2_218 (N2252, N266, N291);
not NOT1_219 (N2253, N272);
not NOT1_220 (N2256, N272);
buf BUFF1_221 (N2257, N269);
buf BUFF1_222 (N2260, N269);
not NOT1_223 (N2263, N276);
not NOT1_224 (N2266, N279);
not NOT1_225 (N2269, N282);
not NOT1_226 (N2272, N285);
not NOT1_227 (N2275, N2104);
not NOT1_228 (N2276, N2104);
not NOT1_229 (N2277, N288);
not NOT1_230 (N2280, N291);
buf BUFF1_231 (N2283, N294);
not NOT1_232 (N2290, N294);
buf BUFF1_233 (N2297, N294);
not NOT1_234 (N2300, N294);
buf BUFF1_235 (N2303, N299);
not NOT1_236 (N2306, N299);
not NOT1_237 (N2313, N299);
buf BUFF1_238 (N2316, N2104);
not NOT1_239 (N2319, N2104);
buf BUFF1_240 (N2326, N2104);
buf BUFF1_241 (N2331, N2104);
not NOT1_242 (N2338, N2104);
buf BUFF1_243 (N2343, N21);
buf BUFF1_244 (N2346, N24);
buf BUFF1_245 (N2349, N27);
buf BUFF1_246 (N2352, N210);
buf BUFF1_247 (N2355, N213);
buf BUFF1_248 (N2358, N216);
buf BUFF1_249 (N2361, N219);
buf BUFF1_250 (N2364, N222);
buf BUFF1_251 (N2367, N225);
buf BUFF1_252 (N2370, N228);
buf BUFF1_253 (N2373, N231);
buf BUFF1_254 (N2376, N234);
buf BUFF1_255 (N2379, N237);
buf BUFF1_256 (N2382, N240);
buf BUFF1_257 (N2385, N243);
buf BUFF1_258 (N2388, N246);
not NOT1_259 (N2534, N2343);
not NOT1_260 (N2535, N2346);
not NOT1_261 (N2536, N2349);
not NOT1_262 (N2537, N2352);
not NOT1_263 (N2538, N2355);
not NOT1_264 (N2539, N2358);
not NOT1_265 (N2540, N2361);
not NOT1_266 (N2541, N2364);
not NOT1_267 (N2542, N2367);
not NOT1_268 (N2543, N2370);
not NOT1_269 (N2544, N2373);
not NOT1_270 (N2545, N2376);
not NOT1_271 (N2546, N2379);
not NOT1_272 (N2547, N2382);
not NOT1_273 (N2548, N2385);
not NOT1_274 (N2549, N2388);
nand NAND2_275 (N2550, N2306, N2331);
nand NAND2_276 (N2551, N2306, N2331);
nand NAND2_277 (N2552, N2306, N2331);
nand NAND2_278 (N2553, N2306, N2331);
nand NAND2_279 (N2554, N2306, N2331);
nand NAND2_280 (N2555, N2306, N2331);
buf BUFF1_281 (N2556, N2190);
buf BUFF1_282 (N2559, N2194);
buf BUFF1_283 (N2562, N2206);
buf BUFF1_284 (N2565, N2209);
buf BUFF1_285 (N2568, N2225);
buf BUFF1_286 (N2571, N2243);
and AND2_287 (N2574, N263, N2319);
buf BUFF1_288 (N2577, N2220);
buf BUFF1_289 (N2580, N2229);
buf BUFF1_290 (N2583, N2232);
and AND2_291 (N2586, N266, N2319);
buf BUFF1_292 (N2589, N2239);
and AND3_293 (N2592, N249, N2253, N2319);
buf BUFF1_294 (N2595, N2247);
buf BUFF1_295 (N2598, N2239);
nand NAND2_296 (N2601, N2326, N2277);
nand NAND2_297 (N2602, N2326, N2280);
nand NAND2_298 (N2603, N2260, N272);
nand NAND2_299 (N2608, N2260, N2300);
nand NAND2_2100 (N2612, N2256, N2300);
buf BUFF1_2101 (N2616, N2201);
buf BUFF1_2102 (N2619, N2216);
buf BUFF1_2103 (N2622, N2220);
buf BUFF1_2104 (N2625, N2239);
buf BUFF1_2105 (N2628, N2190);
buf BUFF1_2106 (N2631, N2190);
buf BUFF1_2107 (N2634, N2194);
buf BUFF1_2108 (N2637, N2229);
buf BUFF1_2109 (N2640, N2197);
and AND3_2110 (N2643, N256, N2257, N2319);
buf BUFF1_2111 (N2646, N2232);
buf BUFF1_2112 (N2649, N2201);
buf BUFF1_2113 (N2652, N2235);
and AND3_2114 (N2655, N260, N2257, N2319);
buf BUFF1_2115 (N2658, N2263);
buf BUFF1_2116 (N2661, N2263);
buf BUFF1_2117 (N2664, N2266);
buf BUFF1_2118 (N2667, N2266);
buf BUFF1_2119 (N2670, N2269);
buf BUFF1_2120 (N2673, N2269);
buf BUFF1_2121 (N2676, N2272);
buf BUFF1_2122 (N2679, N2272);
and AND2_2123 (N2682, N2251, N2316);
and AND2_2124 (N2685, N2252, N2316);
buf BUFF1_2125 (N2688, N2197);
buf BUFF1_2126 (N2691, N2197);
buf BUFF1_2127 (N2694, N2212);
buf BUFF1_2128 (N2697, N2212);
buf BUFF1_2129 (N2700, N2247);
buf BUFF1_2130 (N2703, N2247);
buf BUFF1_2131 (N2706, N2235);
buf BUFF1_2132 (N2709, N2235);
buf BUFF1_2133 (N2712, N2201);
buf BUFF1_2134 (N2715, N2201);
buf BUFF1_2135 (N2718, N2206);
buf BUFF1_2136 (N2721, N2216);
and AND3_2137 (N2724, N253, N2253, N2319);
buf BUFF1_2138 (N2727, N2243);
buf BUFF1_2139 (N2730, N2220);
buf BUFF1_2140 (N2733, N2220);
buf BUFF1_2141 (N2736, N2209);
buf BUFF1_2142 (N2739, N2216);
buf BUFF1_2143 (N2742, N2225);
buf BUFF1_2144 (N2745, N2243);
buf BUFF1_2145 (N2748, N2212);
buf BUFF1_2146 (N2751, N2225);
not NOT1_2147 (N2886, N2682);
not NOT1_2148 (N2887, N2685);
not NOT1_2149 (N2888, N2616);
not NOT1_2150 (N2889, N2619);
not NOT1_2151 (N2890, N2622);
not NOT1_2152 (N2891, N2625);
not NOT1_2153 (N2892, N2631);
not NOT1_2154 (N2893, N2643);
not NOT1_2155 (N2894, N2649);
not NOT1_2156 (N2895, N2652);
not NOT1_2157 (N2896, N2655);
and AND2_2158 (N2897, N249, N2612);
and AND2_2159 (N2898, N256, N2608);
nand NAND2_2160 (N2899, N253, N2612);
nand NAND2_2161 (N2903, N260, N2608);
nand NAND2_2162 (N2907, N249, N2612);
nand NAND2_2163 (N2910, N256, N2608);
not NOT1_2164 (N2913, N2661);
not NOT1_2165 (N2914, N2658);
not NOT1_2166 (N2915, N2667);
not NOT1_2167 (N2916, N2664);
not NOT1_2168 (N2917, N2673);
not NOT1_2169 (N2918, N2670);
not NOT1_2170 (N2919, N2679);
not NOT1_2171 (N2920, N2676);
nand NAND4_2172 (N2921, N2277, N2297, N2326, N2603);
nand NAND4_2173 (N2922, N2280, N2297, N2326, N2603);
nand NAND3_2174 (N2923, N2303, N2338, N2603);
and AND3_2175 (N2926, N2303, N2338, N2603);
buf BUFF1_2176 (N2935, N2556);
not NOT1_2177 (N2938, N2688);
buf BUFF1_2178 (N2939, N2556);
not NOT1_2179 (N2942, N2691);
buf BUFF1_2180 (N2943, N2562);
not NOT1_2181 (N2946, N2694);
buf BUFF1_2182 (N2947, N2562);
not NOT1_2183 (N2950, N2697);
buf BUFF1_2184 (N2951, N2568);
not NOT1_2185 (N2954, N2700);
buf BUFF1_2186 (N2955, N2568);
not NOT1_2187 (N2958, N2703);
buf BUFF1_2188 (N2959, N2574);
buf BUFF1_2189 (N2962, N2574);
buf BUFF1_2190 (N2965, N2580);
not NOT1_2191 (N2968, N2706);
buf BUFF1_2192 (N2969, N2580);
not NOT1_2193 (N2972, N2709);
buf BUFF1_2194 (N2973, N2586);
not NOT1_2195 (N2976, N2712);
buf BUFF1_2196 (N2977, N2586);
not NOT1_2197 (N2980, N2715);
buf BUFF1_2198 (N2981, N2592);
not NOT1_2199 (N2984, N2628);
buf BUFF1_2200 (N2985, N2592);
not NOT1_2201 (N2988, N2718);
not NOT1_2202 (N2989, N2721);
not NOT1_2203 (N2990, N2634);
not NOT1_2204 (N2991, N2724);
not NOT1_2205 (N2992, N2727);
not NOT1_2206 (N2993, N2637);
buf BUFF1_2207 (N2994, N2595);
not NOT1_2208 (N2997, N2730);
buf BUFF1_2209 (N2998, N2595);
not NOT1_2210 (N21001, N2733);
not NOT1_2211 (N21002, N2736);
not NOT1_2212 (N21003, N2739);
not NOT1_2213 (N21004, N2640);
not NOT1_2214 (N21005, N2742);
not NOT1_2215 (N21006, N2745);
not NOT1_2216 (N21007, N2646);
not NOT1_2217 (N21008, N2748);
not NOT1_2218 (N21009, N2751);
buf BUFF1_2219 (N21010, N2559);
buf BUFF1_2220 (N21013, N2559);
buf BUFF1_2221 (N21016, N2565);
buf BUFF1_2222 (N21019, N2565);
buf BUFF1_2223 (N21022, N2571);
buf BUFF1_2224 (N21025, N2571);
buf BUFF1_2225 (N21028, N2577);
buf BUFF1_2226 (N21031, N2577);
buf BUFF1_2227 (N21034, N2583);
buf BUFF1_2228 (N21037, N2583);
buf BUFF1_2229 (N21040, N2589);
buf BUFF1_2230 (N21043, N2589);
buf BUFF1_2231 (N21046, N2598);
buf BUFF1_2232 (N21049, N2598);
nand NAND2_2233 (N21054, N2619, N2888);
nand NAND2_2234 (N21055, N2616, N2889);
nand NAND2_2235 (N21063, N2625, N2890);
nand NAND2_2236 (N21064, N2622, N2891);
nand NAND2_2237 (N21067, N2655, N2895);
nand NAND2_2238 (N21068, N2652, N2896);
nand NAND2_2239 (N21119, N2721, N2988);
nand NAND2_2240 (N21120, N2718, N2989);
nand NAND2_2241 (N21121, N2727, N2991);
nand NAND2_2242 (N21122, N2724, N2992);
nand NAND2_2243 (N21128, N2739, N21002);
nand NAND2_2244 (N21129, N2736, N21003);
nand NAND2_2245 (N21130, N2745, N21005);
nand NAND2_2246 (N21131, N2742, N21006);
nand NAND2_2247 (N21132, N2751, N21008);
nand NAND2_2248 (N21133, N2748, N21009);
not NOT1_2249 (N21148, N2939);
not NOT1_2250 (N21149, N2935);
nand NAND2_2251 (N21150, N21054, N21055);
not NOT1_2252 (N21151, N2943);
not NOT1_2253 (N21152, N2947);
not NOT1_2254 (N21153, N2955);
not NOT1_2255 (N21154, N2951);
not NOT1_2256 (N21155, N2962);
not NOT1_2257 (N21156, N2969);
not NOT1_2258 (N21157, N2977);
nand NAND2_2259 (N21158, N21063, N21064);
not NOT1_2260 (N21159, N2985);
nand NAND2_2261 (N21160, N2985, N2892);
not NOT1_2262 (N21161, N2998);
nand NAND2_2263 (N21162, N21067, N21068);
not NOT1_2264 (N21163, N2899);
buf BUFF1_2265 (N21164, N2899);
not NOT1_2266 (N21167, N2903);
buf BUFF1_2267 (N21168, N2903);
nand NAND2_2268 (N21171, N2921, N2923);
nand NAND2_2269 (N21188, N2922, N2923);
not NOT1_2270 (N21205, N21010);
nand NAND2_2271 (N21206, N21010, N2938);
not NOT1_2272 (N21207, N21013);
nand NAND2_2273 (N21208, N21013, N2942);
not NOT1_2274 (N21209, N21016);
nand NAND2_2275 (N21210, N21016, N2946);
not NOT1_2276 (N21211, N21019);
nand NAND2_2277 (N21212, N21019, N2950);
not NOT1_2278 (N21213, N21022);
nand NAND2_2279 (N21214, N21022, N2954);
not NOT1_2280 (N21215, N21025);
nand NAND2_2281 (N21216, N21025, N2958);
not NOT1_2282 (N21217, N21028);
not NOT1_2283 (N21218, N2959);
not NOT1_2284 (N21219, N21031);
not NOT1_2285 (N21220, N21034);
nand NAND2_2286 (N21221, N21034, N2968);
not NOT1_2287 (N21222, N2965);
not NOT1_2288 (N21223, N21037);
nand NAND2_2289 (N21224, N21037, N2972);
not NOT1_2290 (N21225, N21040);
nand NAND2_2291 (N21226, N21040, N2976);
not NOT1_2292 (N21227, N2973);
not NOT1_2293 (N21228, N21043);
nand NAND2_2294 (N21229, N21043, N2980);
not NOT1_2295 (N21230, N2981);
nand NAND2_2296 (N21231, N2981, N2984);
nand NAND2_2297 (N21232, N21119, N21120);
nand NAND2_2298 (N21235, N21121, N21122);
not NOT1_2299 (N21238, N21046);
nand NAND2_2300 (N21239, N21046, N2997);
not NOT1_2301 (N21240, N2994);
not NOT1_2302 (N21241, N21049);
nand NAND2_2303 (N21242, N21049, N21001);
nand NAND2_2304 (N21243, N21128, N21129);
nand NAND2_2305 (N21246, N21130, N21131);
nand NAND2_2306 (N21249, N21132, N21133);
buf BUFF1_2307 (N21252, N2907);
buf BUFF1_2308 (N21255, N2907);
buf BUFF1_2309 (N21258, N2910);
buf BUFF1_2310 (N21261, N2910);
not NOT1_2311 (N21264, N21150);
nand NAND2_2312 (N21267, N2631, N21159);
nand NAND2_2313 (N21309, N2688, N21205);
nand NAND2_2314 (N21310, N2691, N21207);
nand NAND2_2315 (N21311, N2694, N21209);
nand NAND2_2316 (N21312, N2697, N21211);
nand NAND2_2317 (N21313, N2700, N21213);
nand NAND2_2318 (N21314, N2703, N21215);
nand NAND2_2319 (N21315, N2706, N21220);
nand NAND2_2320 (N21316, N2709, N21223);
nand NAND2_2321 (N21317, N2712, N21225);
nand NAND2_2322 (N21318, N2715, N21228);
not NOT1_2323 (N21319, N21158);
nand NAND2_2324 (N21322, N2628, N21230);
nand NAND2_2325 (N21327, N2730, N21238);
nand NAND2_2326 (N21328, N2733, N21241);
not NOT1_2327 (N21334, N21162);
nand NAND2_2328 (N21344, N21267, N21160);
nand NAND2_2329 (N21345, N21249, N2894);
not NOT1_2330 (N21346, N21249);
not NOT1_2331 (N21348, N21255);
not NOT1_2332 (N21349, N21252);
not NOT1_2333 (N21350, N21261);
not NOT1_2334 (N21351, N21258);
nand NAND2_2335 (N21352, N21309, N21206);
nand NAND2_2336 (N21355, N21310, N21208);
nand NAND2_2337 (N21358, N21311, N21210);
nand NAND2_2338 (N21361, N21312, N21212);
nand NAND2_2339 (N21364, N21313, N21214);
nand NAND2_2340 (N21367, N21314, N21216);
nand NAND2_2341 (N21370, N21315, N21221);
nand NAND2_2342 (N21373, N21316, N21224);
nand NAND2_2343 (N21376, N21317, N21226);
nand NAND2_2344 (N21379, N21318, N21229);
nand NAND2_2345 (N21383, N21322, N21231);
not NOT1_2346 (N21386, N21232);
nand NAND2_2347 (N21387, N21232, N2990);
not NOT1_2348 (N21388, N21235);
nand NAND2_2349 (N21389, N21235, N2993);
nand NAND2_2350 (N21390, N21327, N21239);
nand NAND2_2351 (N21393, N21328, N21242);
not NOT1_2352 (N21396, N21243);
nand NAND2_2353 (N21397, N21243, N21004);
not NOT1_2354 (N21398, N21246);
nand NAND2_2355 (N21399, N21246, N21007);
not NOT1_2356 (N21409, N21319);
nand NAND2_2357 (N21412, N2649, N21346);
not NOT1_2358 (N21413, N21334);
buf BUFF1_2359 (N21416, N21264);
buf BUFF1_2360 (N21419, N21264);
nand NAND2_2361 (N21433, N2634, N21386);
nand NAND2_2362 (N21434, N2637, N21388);
nand NAND2_2363 (N21438, N2640, N21396);
nand NAND2_2364 (N21439, N2646, N21398);
not NOT1_2365 (N21440, N21344);
nand NAND2_2366 (N21443, N21355, N21148);
not NOT1_2367 (N21444, N21355);
nand NAND2_2368 (N21445, N21352, N21149);
not NOT1_2369 (N21446, N21352);
nand NAND2_2370 (N21447, N21358, N21151);
not NOT1_2371 (N21448, N21358);
nand NAND2_2372 (N21451, N21361, N21152);
not NOT1_2373 (N21452, N21361);
nand NAND2_2374 (N21453, N21367, N21153);
not NOT1_2375 (N21454, N21367);
nand NAND2_2376 (N21455, N21364, N21154);
not NOT1_2377 (N21456, N21364);
nand NAND2_2378 (N21457, N21373, N21156);
not NOT1_2379 (N21458, N21373);
nand NAND2_2380 (N21459, N21379, N21157);
not NOT1_2381 (N21460, N21379);
not NOT1_2382 (N21461, N21383);
nand NAND2_2383 (N21462, N21393, N21161);
not NOT1_2384 (N21463, N21393);
nand NAND2_2385 (N21464, N21345, N21412);
not NOT1_2386 (N21468, N21370);
nand NAND2_2387 (N21469, N21370, N21222);
not NOT1_2388 (N21470, N21376);
nand NAND2_2389 (N21471, N21376, N21227);
nand NAND2_2390 (N21472, N21387, N21433);
not NOT1_2391 (N21475, N21390);
nand NAND2_2392 (N21476, N21390, N21240);
nand NAND2_2393 (N21478, N21389, N21434);
nand NAND2_2394 (N21481, N21399, N21439);
nand NAND2_2395 (N21484, N21397, N21438);
nand NAND2_2396 (N21487, N2939, N21444);
nand NAND2_2397 (N21488, N2935, N21446);
nand NAND2_2398 (N21489, N2943, N21448);
not NOT1_2399 (N21490, N21419);
not NOT1_2400 (N21491, N21416);
nand NAND2_2401 (N21492, N2947, N21452);
nand NAND2_2402 (N21493, N2955, N21454);
nand NAND2_2403 (N21494, N2951, N21456);
nand NAND2_2404 (N21495, N2969, N21458);
nand NAND2_2405 (N21496, N2977, N21460);
nand NAND2_2406 (N21498, N2998, N21463);
not NOT1_2407 (N21499, N21440);
nand NAND2_2408 (N21500, N2965, N21468);
nand NAND2_2409 (N21501, N2973, N21470);
nand NAND2_2410 (N21504, N2994, N21475);
not NOT1_2411 (N21510, N21464);
nand NAND2_2412 (N21513, N21443, N21487);
nand NAND2_2413 (N21514, N21445, N21488);
nand NAND2_2414 (N21517, N21447, N21489);
nand NAND2_2415 (N21520, N21451, N21492);
nand NAND2_2416 (N21521, N21453, N21493);
nand NAND2_2417 (N21522, N21455, N21494);
nand NAND2_2418 (N21526, N21457, N21495);
nand NAND2_2419 (N21527, N21459, N21496);
not NOT1_2420 (N21528, N21472);
nand NAND2_2421 (N21529, N21462, N21498);
not NOT1_2422 (N21530, N21478);
not NOT1_2423 (N21531, N21481);
not NOT1_2424 (N21532, N21484);
nand NAND2_2425 (N21534, N21471, N21501);
nand NAND2_2426 (N21537, N21469, N21500);
nand NAND2_2427 (N21540, N21476, N21504);
not NOT1_2428 (N21546, N21513);
not NOT1_2429 (N21554, N21521);
not NOT1_2430 (N21557, N21526);
not NOT1_2431 (N21561, N21520);
nand NAND2_2432 (N21567, N21484, N21531);
nand NAND2_2433 (N21568, N21481, N21532);
not NOT1_2434 (N21569, N21510);
not NOT1_2435 (N21571, N21527);
not NOT1_2436 (N21576, N21529);
buf BUFF1_2437 (N21588, N21522);
not NOT1_2438 (N21591, N21534);
not NOT1_2439 (N21593, N21537);
nand NAND2_2440 (N21594, N21540, N21530);
not NOT1_2441 (N21595, N21540);
nand NAND2_2442 (N21596, N21567, N21568);
buf BUFF1_2443 (N21600, N21517);
buf BUFF1_2444 (N21603, N21517);
buf BUFF1_2445 (N21606, N21522);
buf BUFF1_2446 (N21609, N21522);
buf BUFF1_2447 (N21612, N21514);
buf BUFF1_2448 (N21615, N21514);
buf BUFF1_2449 (N21620, N21557);
buf BUFF1_2450 (N21623, N21554);
not NOT1_2451 (N21635, N21571);
nand NAND2_2452 (N21636, N21478, N21595);
nand NAND2_2453 (N21638, N21576, N21569);
not NOT1_2454 (N21639, N21576);
buf BUFF1_2455 (N21640, N21561);
buf BUFF1_2456 (N21643, N21561);
buf BUFF1_2457 (N21647, N21546);
buf BUFF1_2458 (N21651, N21546);
buf BUFF1_2459 (N21658, N21554);
buf BUFF1_2460 (N21661, N21557);
buf BUFF1_2461 (N21664, N21557);
nand NAND2_2462 (N21671, N21596, N2893);
not NOT1_2463 (N21672, N21596);
not NOT1_2464 (N21675, N21600);
not NOT1_2465 (N21677, N21603);
nand NAND2_2466 (N21678, N21606, N21217);
not NOT1_2467 (N21679, N21606);
nand NAND2_2468 (N21680, N21609, N21219);
not NOT1_2469 (N21681, N21609);
not NOT1_2470 (N21682, N21612);
not NOT1_2471 (N21683, N21615);
nand NAND2_2472 (N21685, N21594, N21636);
nand NAND2_2473 (N21688, N21510, N21639);
buf BUFF1_2474 (N21697, N21588);
buf BUFF1_2475 (N21701, N21588);
nand NAND2_2476 (N21706, N2643, N21672);
not NOT1_2477 (N21707, N21643);
nand NAND2_2478 (N21708, N21647, N21675);
not NOT1_2479 (N21709, N21647);
nand NAND2_2480 (N21710, N21651, N21677);
not NOT1_2481 (N21711, N21651);
nand NAND2_2482 (N21712, N21028, N21679);
nand NAND2_2483 (N21713, N21031, N21681);
buf BUFF1_2484 (N21714, N21620);
buf BUFF1_2485 (N21717, N21620);
nand NAND2_2486 (N21720, N21658, N21593);
not NOT1_2487 (N21721, N21658);
nand NAND2_2488 (N21723, N21638, N21688);
not NOT1_2489 (N21727, N21661);
not NOT1_2490 (N21728, N21640);
not NOT1_2491 (N21730, N21664);
buf BUFF1_2492 (N21731, N21623);
buf BUFF1_2493 (N21734, N21623);
nand NAND2_2494 (N21740, N21685, N21528);
not NOT1_2495 (N21741, N21685);
nand NAND2_2496 (N21742, N21671, N21706);
nand NAND2_2497 (N21746, N21600, N21709);
nand NAND2_2498 (N21747, N21603, N21711);
nand NAND2_2499 (N21748, N21678, N21712);
nand NAND2_2500 (N21751, N21680, N21713);
nand NAND2_2501 (N21759, N21537, N21721);
not NOT1_2502 (N21761, N21697);
nand NAND2_2503 (N21762, N21697, N21727);
not NOT1_2504 (N21763, N21701);
nand NAND2_2505 (N21764, N21701, N21730);
not NOT1_2506 (N21768, N21717);
nand NAND2_2507 (N21769, N21472, N21741);
nand NAND2_2508 (N21772, N21723, N21413);
not NOT1_2509 (N21773, N21723);
nand NAND2_2510 (N21774, N21708, N21746);
nand NAND2_2511 (N21777, N21710, N21747);
not NOT1_2512 (N21783, N21731);
nand NAND2_2513 (N21784, N21731, N21682);
not NOT1_2514 (N21785, N21714);
not NOT1_2515 (N21786, N21734);
nand NAND2_2516 (N21787, N21734, N21683);
nand NAND2_2517 (N21788, N21720, N21759);
nand NAND2_2518 (N21791, N21661, N21761);
nand NAND2_2519 (N21792, N21664, N21763);
nand NAND2_2520 (N21795, N21751, N21155);
not NOT1_2521 (N21796, N21751);
nand NAND2_2522 (N21798, N21740, N21769);
nand NAND2_2523 (N21801, N21334, N21773);
nand NAND2_2524 (N21802, N21742, N2290);
not NOT1_2525 (N21807, N21748);
nand NAND2_2526 (N21808, N21748, N21218);
nand NAND2_2527 (N21809, N21612, N21783);
nand NAND2_2528 (N21810, N21615, N21786);
nand NAND2_2529 (N21812, N21791, N21762);
nand NAND2_2530 (N21815, N21792, N21764);
buf BUFF1_2531 (N21818, N21742);
nand NAND2_2532 (N21821, N21777, N21490);
not NOT1_2533 (N21822, N21777);
nand NAND2_2534 (N21823, N21774, N21491);
not NOT1_2535 (N21824, N21774);
nand NAND2_2536 (N21825, N2962, N21796);
nand NAND2_2537 (N21826, N21788, N21409);
not NOT1_2538 (N21827, N21788);
nand NAND2_2539 (N21830, N21772, N21801);
nand NAND2_2540 (N21837, N2959, N21807);
nand NAND2_2541 (N21838, N21809, N21784);
nand NAND2_2542 (N21841, N21810, N21787);
nand NAND2_2543 (N21848, N21419, N21822);
nand NAND2_2544 (N21849, N21416, N21824);
nand NAND2_2545 (N21850, N21795, N21825);
nand NAND2_2546 (N21852, N21319, N21827);
nand NAND2_2547 (N21855, N21815, N21707);
not NOT1_2548 (N21856, N21815);
not NOT1_2549 (N21857, N21818);
nand NAND2_2550 (N21858, N21798, N2290);
not NOT1_2551 (N21864, N21812);
nand NAND2_2552 (N21865, N21812, N21728);
buf BUFF1_2553 (N21866, N21798);
buf BUFF1_2554 (N21869, N21802);
buf BUFF1_2555 (N21872, N21802);
nand NAND2_2556 (N21875, N21808, N21837);
nand NAND2_2557 (N21878, N21821, N21848);
nand NAND2_2558 (N21879, N21823, N21849);
nand NAND2_2559 (N21882, N21841, N21768);
not NOT1_2560 (N21883, N21841);
nand NAND2_2561 (N21884, N21826, N21852);
nand NAND2_2562 (N21885, N21643, N21856);
nand NAND2_2563 (N21889, N21830, N2290);
not NOT1_2564 (N21895, N21838);
nand NAND2_2565 (N21896, N21838, N21785);
nand NAND2_2566 (N21897, N21640, N21864);
not NOT1_2567 (N21898, N21850);
buf BUFF1_2568 (N21902, N21830);
not NOT1_2569 (N21910, N21878);
nand NAND2_2570 (N21911, N21717, N21883);
not NOT1_2571 (N21912, N21884);
nand NAND2_2572 (N21913, N21855, N21885);
not NOT1_2573 (N21915, N21866);
nand NAND2_2574 (N21919, N21872, N2919);
not NOT1_2575 (N21920, N21872);
nand NAND2_2576 (N21921, N21869, N2920);
not NOT1_2577 (N21922, N21869);
not NOT1_2578 (N21923, N21875);
nand NAND2_2579 (N21924, N21714, N21895);
buf BUFF1_2580 (N21927, N21858);
buf BUFF1_2581 (N21930, N21858);
nand NAND2_2582 (N21933, N21865, N21897);
nand NAND2_2583 (N21936, N21882, N21911);
not NOT1_2584 (N21937, N21898);
not NOT1_2585 (N21938, N21902);
nand NAND2_2586 (N21941, N2679, N21920);
nand NAND2_2587 (N21942, N2676, N21922);
buf BUFF1_2588 (N21944, N21879);
not NOT1_2589 (N21947, N21913);
buf BUFF1_2590 (N21950, N21889);
buf BUFF1_2591 (N21953, N21889);
buf BUFF1_2592 (N21958, N21879);
nand NAND2_2593 (N21961, N21896, N21924);
and AND2_2594 (N21965, N21910, N2601);
and AND2_2595 (N21968, N2602, N21912);
nand NAND2_2596 (N21975, N21930, N2917);
not NOT1_2597 (N21976, N21930);
nand NAND2_2598 (N21977, N21927, N2918);
not NOT1_2599 (N21978, N21927);
nand NAND2_2600 (N21979, N21919, N21941);
nand NAND2_2601 (N21980, N21921, N21942);
not NOT1_2602 (N21985, N21933);
not NOT1_2603 (N21987, N21936);
not NOT1_2604 (N21999, N21944);
nand NAND2_2605 (N22000, N21944, N21937);
not NOT1_2606 (N22002, N21947);
nand NAND2_2607 (N22003, N21947, N21499);
nand NAND2_2608 (N22004, N21953, N21350);
not NOT1_2609 (N22005, N21953);
nand NAND2_2610 (N22006, N21950, N21351);
not NOT1_2611 (N22007, N21950);
nand NAND2_2612 (N22008, N2673, N21976);
nand NAND2_2613 (N22009, N2670, N21978);
not NOT1_2614 (N22012, N21979);
not NOT1_2615 (N22013, N21958);
nand NAND2_2616 (N22014, N21958, N21923);
not NOT1_2617 (N22015, N21961);
nand NAND2_2618 (N22016, N21961, N21635);
not NOT1_2619 (N22018, N21965);
not NOT1_2620 (N22019, N21968);
nand NAND2_2621 (N22020, N21898, N21999);
not NOT1_2622 (N22021, N21987);
nand NAND2_2623 (N22022, N21987, N21591);
nand NAND2_2624 (N22023, N21440, N22002);
nand NAND2_2625 (N22024, N21261, N22005);
nand NAND2_2626 (N22025, N21258, N22007);
nand NAND2_2627 (N22026, N21975, N22008);
nand NAND2_2628 (N22027, N21977, N22009);
not NOT1_2629 (N22030, N21980);
buf BUFF1_2630 (N22033, N21980);
nand NAND2_2631 (N22036, N21875, N22013);
nand NAND2_2632 (N22037, N21571, N22015);
nand NAND2_2633 (N22038, N22020, N22000);
nand NAND2_2634 (N22039, N21534, N22021);
nand NAND2_2635 (N22040, N22023, N22003);
nand NAND2_2636 (N22041, N22004, N22024);
nand NAND2_2637 (N22042, N22006, N22025);
not NOT1_2638 (N22047, N22026);
nand NAND2_2639 (N22052, N22036, N22014);
nand NAND2_2640 (N22055, N22037, N22016);
not NOT1_2641 (N22060, N22038);
nand NAND2_2642 (N22061, N22039, N22022);
nand NAND2_2643 (N22062, N22040, N2290);
not NOT1_2644 (N22067, N22041);
not NOT1_2645 (N22068, N22027);
buf BUFF1_2646 (N22071, N22027);
not NOT1_2647 (N22076, N22052);
not NOT1_2648 (N22077, N22055);
nand NAND2_2649 (N22078, N22060, N2290);
nand NAND2_2650 (N22081, N22061, N2290);
not NOT1_2651 (N22086, N22042);
buf BUFF1_2652 (N22089, N22042);
and AND2_2653 (N22104, N22030, N22068);
and AND2_2654 (N22119, N22033, N22068);
and AND2_2655 (N22129, N22030, N22071);
and AND2_2656 (N22143, N22033, N22071);
buf BUFF1_2657 (N22148, N22062);
buf BUFF1_2658 (N22151, N22062);
buf BUFF1_2659 (N22196, N22078);
buf BUFF1_2660 (N22199, N22078);
buf BUFF1_2661 (N22202, N22081);
buf BUFF1_2662 (N22205, N22081);
nand NAND2_2663 (N22214, N22151, N2915);
not NOT1_2664 (N22215, N22151);
nand NAND2_2665 (N22216, N22148, N2916);
not NOT1_2666 (N22217, N22148);
nand NAND2_2667 (N22222, N22199, N21348);
not NOT1_2668 (N22223, N22199);
nand NAND2_2669 (N22224, N22196, N21349);
not NOT1_2670 (N22225, N22196);
nand NAND2_2671 (N22226, N22205, N2913);
not NOT1_2672 (N22227, N22205);
nand NAND2_2673 (N22228, N22202, N2914);
not NOT1_2674 (N22229, N22202);
nand NAND2_2675 (N22230, N2667, N22215);
nand NAND2_2676 (N22231, N2664, N22217);
nand NAND2_2677 (N22232, N21255, N22223);
nand NAND2_2678 (N22233, N21252, N22225);
nand NAND2_2679 (N22234, N2661, N22227);
nand NAND2_2680 (N22235, N2658, N22229);
nand NAND2_2681 (N22236, N22214, N22230);
nand NAND2_2682 (N22237, N22216, N22231);
nand NAND2_2683 (N22240, N22222, N22232);
nand NAND2_2684 (N22241, N22224, N22233);
nand NAND2_2685 (N22244, N22226, N22234);
nand NAND2_2686 (N22245, N22228, N22235);
not NOT1_2687 (N22250, N22236);
not NOT1_2688 (N22253, N22240);
not NOT1_2689 (N22256, N22244);
not NOT1_2690 (N22257, N22237);
buf BUFF1_2691 (N22260, N22237);
not NOT1_2692 (N22263, N22241);
and AND2_2693 (N22266, N21164, N22241);
not NOT1_2694 (N22269, N22245);
and AND2_2695 (N22272, N21168, N22245);
nand NAND8_2696 (N22279, N22067, N22012, N22047, N22250, N2899, N22256, N22253, N2903);
buf BUFF1_2697 (N22286, N22266);
buf BUFF1_2698 (N22297, N22266);
buf BUFF1_2699 (N22315, N22272);
buf BUFF1_2700 (N22326, N22272);
and AND2_2701 (N22340, N22086, N22257);
and AND2_2702 (N22353, N22089, N22257);
and AND2_2703 (N22361, N22086, N22260);
and AND2_2704 (N22375, N22089, N22260);
and AND4_2705 (N22384, N2338, N22279, N2313, N2313);
and AND2_2706 (N22385, N21163, N22263);
and AND2_2707 (N22386, N21164, N22263);
and AND2_2708 (N22426, N21167, N22269);
and AND2_2709 (N22427, N21168, N22269);
nand NAND5_2710 (N22537, N22286, N22315, N22361, N22104, N21171);
nand NAND5_2711 (N22540, N22286, N22315, N22340, N22129, N21171);
nand NAND5_2712 (N22543, N22286, N22315, N22340, N22119, N21171);
nand NAND5_2713 (N22546, N22286, N22315, N22353, N22104, N21171);
nand NAND5_2714 (N22549, N22297, N22315, N22375, N22119, N21188);
nand NAND5_2715 (N22552, N22297, N22326, N22361, N22143, N21188);
nand NAND5_2716 (N22555, N22297, N22326, N22375, N22129, N21188);
and AND5_2717 (N22558, N22286, N22315, N22361, N22104, N21171);
and AND5_2718 (N22561, N22286, N22315, N22340, N22129, N21171);
and AND5_2719 (N22564, N22286, N22315, N22340, N22119, N21171);
and AND5_2720 (N22567, N22286, N22315, N22353, N22104, N21171);
and AND5_2721 (N22570, N22297, N22315, N22375, N22119, N21188);
and AND5_2722 (N22573, N22297, N22326, N22361, N22143, N21188);
and AND5_2723 (N22576, N22297, N22326, N22375, N22129, N21188);
nand NAND5_2724 (N22594, N22286, N22427, N22361, N22129, N21171);
nand NAND5_2725 (N22597, N22297, N22427, N22361, N22119, N21171);
nand NAND5_2726 (N22600, N22297, N22427, N22375, N22104, N21171);
nand NAND5_2727 (N22603, N22297, N22427, N22340, N22143, N21171);
nand NAND5_2728 (N22606, N22297, N22427, N22353, N22129, N21188);
nand NAND5_2729 (N22611, N22386, N22326, N22361, N22129, N21188);
nand NAND5_2730 (N22614, N22386, N22326, N22361, N22119, N21188);
nand NAND5_2731 (N22617, N22386, N22326, N22375, N22104, N21188);
nand NAND5_2732 (N22620, N22386, N22326, N22353, N22129, N21188);
nand NAND5_2733 (N22627, N22297, N22427, N22340, N22104, N2926);
nand NAND5_2734 (N22628, N22386, N22326, N22340, N22104, N2926);
nand NAND5_2735 (N22629, N22386, N22427, N22361, N22104, N2926);
nand NAND5_2736 (N22630, N22386, N22427, N22340, N22129, N2926);
nand NAND5_2737 (N22631, N22386, N22427, N22340, N22119, N2926);
nand NAND5_2738 (N22632, N22386, N22427, N22353, N22104, N2926);
nand NAND5_2739 (N22633, N22386, N22426, N22340, N22104, N2926);
nand NAND5_2740 (N22634, N22385, N22427, N22340, N22104, N2926);
and AND5_2741 (N22639, N22286, N22427, N22361, N22129, N21171);
and AND5_2742 (N22642, N22297, N22427, N22361, N22119, N21171);
and AND5_2743 (N22645, N22297, N22427, N22375, N22104, N21171);
and AND5_2744 (N22648, N22297, N22427, N22340, N22143, N21171);
and AND5_2745 (N22651, N22297, N22427, N22353, N22129, N21188);
and AND5_2746 (N22655, N22386, N22326, N22361, N22129, N21188);
and AND5_2747 (N22658, N22386, N22326, N22361, N22119, N21188);
and AND5_2748 (N22661, N22386, N22326, N22375, N22104, N21188);
and AND5_2749 (N22664, N22386, N22326, N22353, N22129, N21188);
nand NAND2_2750 (N22669, N22558, N2534);
not NOT1_2751 (N22670, N22558);
nand NAND2_2752 (N22671, N22561, N2535);
not NOT1_2753 (N22672, N22561);
nand NAND2_2754 (N22673, N22564, N2536);
not NOT1_2755 (N22674, N22564);
nand NAND2_2756 (N22675, N22567, N2537);
not NOT1_2757 (N22676, N22567);
nand NAND2_2758 (N22682, N22570, N2543);
not NOT1_2759 (N22683, N22570);
nand NAND2_2760 (N22688, N22573, N2548);
not NOT1_2761 (N22689, N22573);
nand NAND2_2762 (N22690, N22576, N2549);
not NOT1_2763 (N22691, N22576);
and AND8_2764 (N22710, N22627, N22628, N22629, N22630, N22631, N22632, N22633, N22634);
nand NAND2_2765 (N22720, N2343, N22670);
nand NAND2_2766 (N22721, N2346, N22672);
nand NAND2_2767 (N22722, N2349, N22674);
nand NAND2_2768 (N22723, N2352, N22676);
nand NAND2_2769 (N22724, N22639, N2538);
not NOT1_2770 (N22725, N22639);
nand NAND2_2771 (N22726, N22642, N2539);
not NOT1_2772 (N22727, N22642);
nand NAND2_2773 (N22728, N22645, N2540);
not NOT1_2774 (N22729, N22645);
nand NAND2_2775 (N22730, N22648, N2541);
not NOT1_2776 (N22731, N22648);
nand NAND2_2777 (N22732, N22651, N2542);
not NOT1_2778 (N22733, N22651);
nand NAND2_2779 (N22734, N2370, N22683);
nand NAND2_2780 (N22735, N22655, N2544);
not NOT1_2781 (N22736, N22655);
nand NAND2_2782 (N22737, N22658, N2545);
not NOT1_2783 (N22738, N22658);
nand NAND2_2784 (N22739, N22661, N2546);
not NOT1_2785 (N22740, N22661);
nand NAND2_2786 (N22741, N22664, N2547);
not NOT1_2787 (N22742, N22664);
nand NAND2_2788 (N22743, N2385, N22689);
nand NAND2_2789 (N22744, N2388, N22691);
nand NAND8_2790 (N22745, N22537, N22540, N22543, N22546, N22594, N22597, N22600, N22603);
nand NAND8_2791 (N22746, N22606, N22549, N22611, N22614, N22617, N22620, N22552, N22555);
and AND8_2792 (N22747, N22537, N22540, N22543, N22546, N22594, N22597, N22600, N22603);
and AND8_2793 (N22750, N22606, N22549, N22611, N22614, N22617, N22620, N22552, N22555);
nand NAND2_2794 (N22753, N22669, N22720);
nand NAND2_2795 (N22754, N22671, N22721);
nand NAND2_2796 (N22755, N22673, N22722);
nand NAND2_2797 (N22756, N22675, N22723);
nand NAND2_2798 (N22757, N2355, N22725);
nand NAND2_2799 (N22758, N2358, N22727);
nand NAND2_2800 (N22759, N2361, N22729);
nand NAND2_2801 (N22760, N2364, N22731);
nand NAND2_2802 (N22761, N2367, N22733);
nand NAND2_2803 (N22762, N22682, N22734);
nand NAND2_2804 (N22763, N2373, N22736);
nand NAND2_2805 (N22764, N2376, N22738);
nand NAND2_2806 (N22765, N2379, N22740);
nand NAND2_2807 (N22766, N2382, N22742);
nand NAND2_2808 (N22767, N22688, N22743);
nand NAND2_2809 (N22768, N22690, N22744);
and AND2_2810 (N22773, N22745, N2275);
and AND2_2811 (N22776, N22746, N2276);
nand NAND2_2812 (N22779, N22724, N22757);
nand NAND2_2813 (N22780, N22726, N22758);
nand NAND2_2814 (N22781, N22728, N22759);
nand NAND2_2815 (N22782, N22730, N22760);
nand NAND2_2816 (N22783, N22732, N22761);
nand NAND2_2817 (N22784, N22735, N22763);
nand NAND2_2818 (N22785, N22737, N22764);
nand NAND2_2819 (N22786, N22739, N22765);
nand NAND2_2820 (N22787, N22741, N22766);
and AND3_2821 (N22788, N22747, N22750, N22710);
nand NAND2_2822 (N22789, N22747, N22750);
and AND4_2823 (N22800, N2338, N22279, N299, N22788);
nand NAND2_2824 (N22807, N22773, N22018);
not NOT1_2825 (N22808, N22773);
nand NAND2_2826 (N22809, N22776, N22019);
not NOT1_2827 (N22810, N22776);
nor N2OR2_2828 (N22811, N22384, N22800);
and AND3_2829 (N22812, N2897, N2283, N22789);
and AND3_2830 (N22815, N276, N2283, N22789);
and AND3_2831 (N22818, N282, N2283, N22789);
and AND3_2832 (N22821, N285, N2283, N22789);
and AND3_2833 (N22824, N2898, N2283, N22789);
nand NAND2_2834 (N22827, N21965, N22808);
nand NAND2_2835 (N22828, N21968, N22810);
and AND3_2836 (N22829, N279, N2283, N22789);
nand NAND2_2837 (N22843, N22807, N22827);
nand NAND2_2838 (N22846, N22809, N22828);
nand NAND2_2839 (N22850, N22812, N22076);
nand NAND2_2840 (N22851, N22815, N22077);
nand NAND2_2841 (N22852, N22818, N21915);
nand NAND2_2842 (N22853, N22821, N21857);
nand NAND2_2843 (N22854, N22824, N21938);
not NOT1_2844 (N22857, N22812);
not NOT1_2845 (N22858, N22815);
not NOT1_2846 (N22859, N22818);
not NOT1_2847 (N22860, N22821);
not NOT1_2848 (N22861, N22824);
not NOT1_2849 (N22862, N22829);
nand NAND2_2850 (N22863, N22829, N21985);
nand NAND2_2851 (N22866, N22052, N22857);
nand NAND2_2852 (N22867, N22055, N22858);
nand NAND2_2853 (N22868, N21866, N22859);
nand NAND2_2854 (N22869, N21818, N22860);
nand NAND2_2855 (N22870, N21902, N22861);
nand NAND2_2856 (N22871, N22843, N2886);
not NOT1_2857 (N22872, N22843);
nand NAND2_2858 (N22873, N22846, N2887);
not NOT1_2859 (N22874, N22846);
nand NAND2_2860 (N22875, N21933, N22862);
nand NAND2_2861 (N22876, N22866, N22850);
nand NAND2_2862 (N22877, N22867, N22851);
nand NAND2_2863 (N22878, N22868, N22852);
nand NAND2_2864 (N22879, N22869, N22853);
nand NAND2_2865 (N22880, N22870, N22854);
nand NAND2_2866 (N22881, N2682, N22872);
nand NAND2_2867 (N22882, N2685, N22874);
nand NAND2_2868 (N22883, N22875, N22863);
and AND2_2869 (N22886, N22876, N2550);
and AND2_2870 (N22887, N2551, N22877);
and AND2_2871 (N22888, N2553, N22878);
and AND2_2872 (N22889, N22879, N2554);
and AND2_2873 (N22890, N2555, N22880);
nand NAND2_2874 (N22891, N22871, N22881);
nand NAND2_2875 (N22892, N22873, N22882);
nand NAND2_2876 (N22895, N22883, N21461);
not NOT1_2877 (N22896, N22883);
nand NAND2_2878 (N22897, N21383, N22896);
nand NAND2_2879 (N22898, N22895, N22897);
and AND2_2880 (N22899, N22898, N2552);

endmodule
