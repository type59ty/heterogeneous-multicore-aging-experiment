`timescale 1ns/10ps

`define cycle 10.0
`define terminate_cycle 400000//200000 // Modify your terminate ycle here

module b18_ras_testfixture;

`define in_file "b18_ras/rand_input_vector_b18_ras_0.out"
`define out_file "b18_ras/rand_output_vector_b18_ras_0.out"

parameter vec_width = 3357;
parameter vec_length = 7;

reg clk = 0;


reg [vec_width-1:0] input_vec_mem [0:vec_length-1];
reg [vec_width-1:0] vec;

wire logic0_po_extra, mul_1411_u378, mul_1411_u438, mul_1411_u10, mul_1411_u439, mul_1411_u9, mul_1411_u440, mul_1411_u8, mul_1411_u441, mul_1411_u7, mul_1411_u385, mul_1411_u14, mul_1411_u386, mul_1411_u13, mul_1411_u387, mul_1411_u12, mul_1411_u388, mul_1411_u11, mul_1411_u15, mul_1411_u5_po_extra, mul_1421_a1_u5, u154, u39_po_extra, p1_u247, p1_u246, p1_u245, p1_u244, p1_u243, p1_u242, p1_u241, p1_u240, p1_u239, p1_u238, p1_u237, p1_u236, p1_u235, p1_u234, p1_u233, p1_u232, p1_u231, p1_u230, p1_u229, p1_u228, p1_u227, p1_u226, p1_u225, p1_u224, p1_u223, p1_u222, p1_u221, p1_u220, p1_u219, p1_u218, p1_u217, p1_u216, p1_u251, p1_u252, p1_u253, p1_u254, p1_u255, p1_u256, p1_u257, p1_u258, p1_u259, p1_u260, p1_u261, p1_u262, p1_u263, p1_u264, p1_u265, p1_u266, p1_u267, p1_u268, p1_u269, p1_u270, p1_u271, p1_u272, p1_u273, p1_u274, p1_u275, p1_u276, p1_u277, p1_u278, p1_u279, p1_u280, p1_u281, p1_u282, p1_u212, p1_u215, p1_u213, p1_u214, p2_u247, p2_u246, p2_u245, p2_u244, p2_u243, p2_u242, p2_u241, p2_u240, p2_u239, p2_u238, p2_u237, p2_u236, p2_u235, p2_u234, p2_u233, p2_u232, p2_u231, p2_u230, p2_u229, p2_u228, p2_u227, p2_u226, p2_u225, p2_u224, p2_u223, p2_u222, p2_u221, p2_u220, p2_u219, p2_u218, p2_u217, p2_u216, p2_u251, p2_u252, p2_u253, p2_u254, p2_u255, p2_u256, p2_u257, p2_u258, p2_u259, p2_u260, p2_u261, p2_u262, p2_u263, p2_u264, p2_u265, p2_u266, p2_u267, p2_u268, p2_u269, p2_u270, p2_u271, p2_u272, p2_u273, p2_u274, p2_u275, p2_u276, p2_u277, p2_u278, p2_u279, p2_u280, p2_u281, p2_u282, p2_u212, p2_u215, p2_u213, p2_u214, p3_u3354, p3_u3353, p3_u3352, p3_u3351, p3_u3350, p3_u3349, p3_u3348, p3_u3347, p3_u3346, p3_u3345, p3_u3344, p3_u3343, p3_u3342, p3_u3341, p3_u3340, p3_u3339, p3_u3338, p3_u3337, p3_u3336, p3_u3335, p3_u3334, p3_u3333, p3_u3332, p3_u3331, p3_u3330, p3_u3329, p3_u3328, p3_u3327, p3_u3326, p3_u3325, p3_u3324, p3_u3323, p3_u3442, p3_u3443, p3_u3322, p3_u3321, p3_u3320, p3_u3319, p3_u3318, p3_u3317, p3_u3316, p3_u3315, p3_u3314, p3_u3313, p3_u3312, p3_u3311, p3_u3310, p3_u3309, p3_u3308, p3_u3307, p3_u3306, p3_u3305, p3_u3304, p3_u3303, p3_u3302, p3_u3301, p3_u3300, p3_u3299, p3_u3298, p3_u3297, p3_u3296, p3_u3295, p3_u3294, p3_u3293, p3_u3456, p3_u3459, p3_u3462, p3_u3465, p3_u3468, p3_u3471, p3_u3474, p3_u3477, p3_u3480, p3_u3483, p3_u3486, p3_u3489, p3_u3492, p3_u3495, p3_u3498, p3_u3501, p3_u3504, p3_u3507, p3_u3510, p3_u3512, p3_u3513, p3_u3514, p3_u3515, p3_u3516, p3_u3517, p3_u3518, p3_u3519, p3_u3520, p3_u3521, p3_u3522, p3_u3523, p3_u3524, p3_u3525, p3_u3526, p3_u3527, p3_u3528, p3_u3529, p3_u3530, p3_u3531, p3_u3532, p3_u3533, p3_u3534, p3_u3535, p3_u3536, p3_u3537, p3_u3538, p3_u3539, p3_u3540, p3_u3541, p3_u3542, p3_u3543, p3_u3544, p3_u3545, p3_u3546, p3_u3547, p3_u3548, p3_u3549, p3_u3550, p3_u3551, p3_u3552, p3_u3553, p3_u3554, p3_u3555, p3_u3556, p3_u3292, p3_u3291, p3_u3290, p3_u3289, p3_u3288, p3_u3287, p3_u3286, p3_u3285, p3_u3284, p3_u3283, p3_u3282, p3_u3281, p3_u3280, p3_u3279, p3_u3278, p3_u3277, p3_u3276, p3_u3275, p3_u3274, p3_u3273, p3_u3272, p3_u3271, p3_u3270, p3_u3269, p3_u3268, p3_u3267, p3_u3266, p3_u3265, p3_u3264, p3_u3263, p3_u3262, p3_u3261, p3_u3260, p3_u3259, p3_u3258, p3_u3257, p3_u3256, p3_u3255, p3_u3254, p3_u3253, p3_u3252, p3_u3251, p3_u3250, p3_u3249, p3_u3248, p3_u3247, p3_u3246, p3_u3245, p3_u3244, p3_u3243, p3_u3242, p3_u3241, p3_u3557, p3_u3558, p3_u3559, p3_u3560, p3_u3561, p3_u3562, p3_u3563, p3_u3564, p3_u3565, p3_u3566, p3_u3567, p3_u3568, p3_u3569, p3_u3570, p3_u3571, p3_u3572, p3_u3573, p3_u3574, p3_u3575, p3_u3576, p3_u3577, p3_u3578, p3_u3579, p3_u3580, p3_u3581, p3_u3582, p3_u3583, p3_u3584, p3_u3585, p3_u3586, p3_u3587, p3_u3588, p3_u3240, p3_u3239, p3_u3238, p3_u3237, p3_u3236, p3_u3235, p3_u3234, p3_u3233, p3_u3232, p3_u3231, p3_u3230, p3_u3229, p3_u3228, p3_u3227, p3_u3226, p3_u3225, p3_u3224, p3_u3223, p3_u3222, p3_u3221, p3_u3220, p3_u3219, p3_u3218, p3_u3217, p3_u3216, p3_u3215, p3_u3214, p3_u3213, p3_u3212, p3_u3211, p3_u3084, p3_u3083, p3_u4038, p4_u3351, p4_u3350, p4_u3349, p4_u3348, p4_u3347, p4_u3346, p4_u3345, p4_u3344, p4_u3343, p4_u3342, p4_u3341, p4_u3340, p4_u3339, p4_u3338, p4_u3337, p4_u3336, p4_u3335, p4_u3334, p4_u3333, p4_u3332, p4_u3331, p4_u3330, p4_u3329, p4_u3328, p4_u3327, p4_u3326, p4_u3325, p4_u3324, p4_u3323, p4_u3322, p4_u3321, p4_u3320, p4_u3437, p4_u3438, p4_u3319, p4_u3318, p4_u3317, p4_u3316, p4_u3315, p4_u3314, p4_u3313, p4_u3312, p4_u3311, p4_u3310, p4_u3309, p4_u3308, p4_u3307, p4_u3306, p4_u3305, p4_u3304, p4_u3303, p4_u3302, p4_u3301, p4_u3300, p4_u3299, p4_u3298, p4_u3297, p4_u3296, p4_u3295, p4_u3294, p4_u3293, p4_u3292, p4_u3291, p4_u3290, p4_u3451, p4_u3454, p4_u3457, p4_u3460, p4_u3463, p4_u3466, p4_u3469, p4_u3472, p4_u3475, p4_u3478, p4_u3481, p4_u3484, p4_u3487, p4_u3490, p4_u3493, p4_u3496, p4_u3499, p4_u3502, p4_u3505, p4_u3507, p4_u3508, p4_u3509, p4_u3510, p4_u3511, p4_u3512, p4_u3513, p4_u3514, p4_u3515, p4_u3516, p4_u3517, p4_u3518, p4_u3519, p4_u3520, p4_u3521, p4_u3522, p4_u3523, p4_u3524, p4_u3525, p4_u3526, p4_u3527, p4_u3528, p4_u3529, p4_u3530, p4_u3531, p4_u3532, p4_u3533, p4_u3534, p4_u3535, p4_u3536, p4_u3537, p4_u3538, p4_u3539, p4_u3540, p4_u3541, p4_u3542, p4_u3543, p4_u3544, p4_u3545, p4_u3546, p4_u3547, p4_u3548, p4_u3549, p4_u3550, p4_u3551, p4_u3289, p4_u3288, p4_u3287, p4_u3286, p4_u3285, p4_u3284, p4_u3283, p4_u3282, p4_u3281, p4_u3280, p4_u3279, p4_u3278, p4_u3277, p4_u3276, p4_u3275, p4_u3274, p4_u3273, p4_u3272, p4_u3271, p4_u3270, p4_u3269, p4_u3268, p4_u3267, p4_u3266, p4_u3265, p4_u3264, p4_u3263, p4_u3262, p4_u3261, p4_u3260, p4_u3259, p4_u3258, p4_u3257, p4_u3256, p4_u3255, p4_u3254, p4_u3253, p4_u3252, p4_u3251, p4_u3250, p4_u3249, p4_u3248, p4_u3247, p4_u3246, p4_u3245, p4_u3244, p4_u3243, p4_u3242, p4_u3241, p4_u3240, p4_u3239, p4_u3238, p4_u3552, p4_u3553, p4_u3554, p4_u3555, p4_u3556, p4_u3557, p4_u3558, p4_u3559, p4_u3560, p4_u3561, p4_u3562, p4_u3563, p4_u3564, p4_u3565, p4_u3566, p4_u3567, p4_u3568, p4_u3569, p4_u3570, p4_u3571, p4_u3572, p4_u3573, p4_u3574, p4_u3575, p4_u3576, p4_u3577, p4_u3578, p4_u3579, p4_u3580, p4_u3581, p4_u3582, p4_u3583, p4_u3237, p4_u3236, p4_u3235, p4_u3234, p4_u3233, p4_u3232, p4_u3231, p4_u3230, p4_u3229, p4_u3228, p4_u3227, p4_u3226, p4_u3225, p4_u3224, p4_u3223, p4_u3222, p4_u3221, p4_u3220, p4_u3219, p4_u3218, p4_u3217, p4_u3216, p4_u3215, p4_u3214, p4_u3213, p4_u3212, p4_u3211, p4_u3210, p4_u3209, p4_u3208, p4_u3147, p4_u3146, p4_u4028, p1_p3_u3274, p1_p3_u3275, p1_p3_u3276, p1_p3_u3277, p1_p3_u3061, p1_p3_u3060, p1_p3_u3059, p1_p3_u3058, p1_p3_u3057, p1_p3_u3056, p1_p3_u3055, p1_p3_u3054, p1_p3_u3053, p1_p3_u3052, p1_p3_u3051, p1_p3_u3050, p1_p3_u3049, p1_p3_u3048, p1_p3_u3047, p1_p3_u3046, p1_p3_u3045, p1_p3_u3044, p1_p3_u3043, p1_p3_u3042, p1_p3_u3041, p1_p3_u3040, p1_p3_u3039, p1_p3_u3038, p1_p3_u3037, p1_p3_u3036, p1_p3_u3035, p1_p3_u3034, p1_p3_u3033, p1_p3_u3032, p1_p3_u3031, p1_p3_u3030, p1_p3_u3029, p1_p3_u3280, p1_p3_u3281, p1_p3_u3028, p1_p3_u3027, p1_p3_u3026, p1_p3_u3025, p1_p3_u3024, p1_p3_u3023, p1_p3_u3022, p1_p3_u3021, p1_p3_u3020, p1_p3_u3019, p1_p3_u3018, p1_p3_u3017, p1_p3_u3016, p1_p3_u3015, p1_p3_u3014, p1_p3_u3013, p1_p3_u3012, p1_p3_u3011, p1_p3_u3010, p1_p3_u3009, p1_p3_u3008, p1_p3_u3007, p1_p3_u3006, p1_p3_u3005, p1_p3_u3004, p1_p3_u3003, p1_p3_u3002, p1_p3_u3001, p1_p3_u3000, p1_p3_u2999, p1_p3_u3282, p1_p3_u2998, p1_p3_u2997, p1_p3_u2996, p1_p3_u2995, p1_p3_u2994, p1_p3_u2993, p1_p3_u2992, p1_p3_u2991, p1_p3_u2990, p1_p3_u2989, p1_p3_u2988, p1_p3_u2987, p1_p3_u2986, p1_p3_u2985, p1_p3_u2984, p1_p3_u2983, p1_p3_u2982, p1_p3_u2981, p1_p3_u2980, p1_p3_u2979, p1_p3_u2978, p1_p3_u2977, p1_p3_u2976, p1_p3_u2975, p1_p3_u2974, p1_p3_u2973, p1_p3_u2972, p1_p3_u2971, p1_p3_u2970, p1_p3_u2969, p1_p3_u2968, p1_p3_u2967, p1_p3_u2966, p1_p3_u2965, p1_p3_u2964, p1_p3_u2963, p1_p3_u2962, p1_p3_u2961, p1_p3_u2960, p1_p3_u2959, p1_p3_u2958, p1_p3_u2957, p1_p3_u2956, p1_p3_u2955, p1_p3_u2954, p1_p3_u2953, p1_p3_u2952, p1_p3_u2951, p1_p3_u2950, p1_p3_u2949, p1_p3_u2948, p1_p3_u2947, p1_p3_u2946, p1_p3_u2945, p1_p3_u2944, p1_p3_u2943, p1_p3_u2942, p1_p3_u2941, p1_p3_u2940, p1_p3_u2939, p1_p3_u2938, p1_p3_u2937, p1_p3_u2936, p1_p3_u2935, p1_p3_u2934, p1_p3_u2933, p1_p3_u2932, p1_p3_u2931, p1_p3_u2930, p1_p3_u2929, p1_p3_u2928, p1_p3_u2927, p1_p3_u2926, p1_p3_u2925, p1_p3_u2924, p1_p3_u2923, p1_p3_u2922, p1_p3_u2921, p1_p3_u2920, p1_p3_u2919, p1_p3_u2918, p1_p3_u2917, p1_p3_u2916, p1_p3_u2915, p1_p3_u2914, p1_p3_u2913, p1_p3_u2912, p1_p3_u2911, p1_p3_u2910, p1_p3_u2909, p1_p3_u2908, p1_p3_u2907, p1_p3_u2906, p1_p3_u2905, p1_p3_u2904, p1_p3_u2903, p1_p3_u2902, p1_p3_u2901, p1_p3_u2900, p1_p3_u2899, p1_p3_u2898, p1_p3_u2897, p1_p3_u2896, p1_p3_u2895, p1_p3_u2894, p1_p3_u2893, p1_p3_u2892, p1_p3_u2891, p1_p3_u2890, p1_p3_u2889, p1_p3_u2888, p1_p3_u2887, p1_p3_u2886, p1_p3_u2885, p1_p3_u2884, p1_p3_u2883, p1_p3_u2882, p1_p3_u2881, p1_p3_u2880, p1_p3_u2879, p1_p3_u2878, p1_p3_u2877, p1_p3_u2876, p1_p3_u2875, p1_p3_u2874, p1_p3_u2873, p1_p3_u2872, p1_p3_u2871, p1_p3_u2870, p1_p3_u2869, p1_p3_u2868, p1_p3_u3284, p1_p3_u3285, p1_p3_u3288, p1_p3_u3289, p1_p3_u3290, p1_p3_u2867, p1_p3_u2866, p1_p3_u2865, p1_p3_u2864, p1_p3_u2863, p1_p3_u2862, p1_p3_u2861, p1_p3_u2860, p1_p3_u2859, p1_p3_u2858, p1_p3_u2857, p1_p3_u2856, p1_p3_u2855, p1_p3_u2854, p1_p3_u2853, p1_p3_u2852, p1_p3_u2851, p1_p3_u2850, p1_p3_u2849, p1_p3_u2848, p1_p3_u2847, p1_p3_u2846, p1_p3_u2845, p1_p3_u2844, p1_p3_u2843, p1_p3_u2842, p1_p3_u2841, p1_p3_u2840, p1_p3_u2839, p1_p3_u2838, p1_p3_u2837, p1_p3_u2836, p1_p3_u2835, p1_p3_u2834, p1_p3_u2833, p1_p3_u2832, p1_p3_u2831, p1_p3_u2830, p1_p3_u2829, p1_p3_u2828, p1_p3_u2827, p1_p3_u2826, p1_p3_u2825, p1_p3_u2824, p1_p3_u2823, p1_p3_u2822, p1_p3_u2821, p1_p3_u2820, p1_p3_u2819, p1_p3_u2818, p1_p3_u2817, p1_p3_u2816, p1_p3_u2815, p1_p3_u2814, p1_p3_u2813, p1_p3_u2812, p1_p3_u2811, p1_p3_u2810, p1_p3_u2809, p1_p3_u2808, p1_p3_u2807, p1_p3_u2806, p1_p3_u2805, p1_p3_u2804, p1_p3_u2803, p1_p3_u2802, p1_p3_u2801, p1_p3_u2800, p1_p3_u2799, p1_p3_u2798, p1_p3_u2797, p1_p3_u2796, p1_p3_u2795, p1_p3_u2794, p1_p3_u2793, p1_p3_u2792, p1_p3_u2791, p1_p3_u2790, p1_p3_u2789, p1_p3_u2788, p1_p3_u2787, p1_p3_u2786, p1_p3_u2785, p1_p3_u2784, p1_p3_u2783, p1_p3_u2782, p1_p3_u2781, p1_p3_u2780, p1_p3_u2779, p1_p3_u2778, p1_p3_u2777, p1_p3_u2776, p1_p3_u2775, p1_p3_u2774, p1_p3_u2773, p1_p3_u2772, p1_p3_u2771, p1_p3_u2770, p1_p3_u2769, p1_p3_u2768, p1_p3_u2767, p1_p3_u2766, p1_p3_u2765, p1_p3_u2764, p1_p3_u2763, p1_p3_u2762, p1_p3_u2761, p1_p3_u2760, p1_p3_u2759, p1_p3_u2758, p1_p3_u2757, p1_p3_u2756, p1_p3_u2755, p1_p3_u2754, p1_p3_u2753, p1_p3_u2752, p1_p3_u2751, p1_p3_u2750, p1_p3_u2749, p1_p3_u2748, p1_p3_u2747, p1_p3_u2746, p1_p3_u2745, p1_p3_u2744, p1_p3_u2743, p1_p3_u2742, p1_p3_u2741, p1_p3_u2740, p1_p3_u2739, p1_p3_u2738, p1_p3_u2737, p1_p3_u2736, p1_p3_u2735, p1_p3_u2734, p1_p3_u2733, p1_p3_u2732, p1_p3_u2731, p1_p3_u2730, p1_p3_u2729, p1_p3_u2728, p1_p3_u2727, p1_p3_u2726, p1_p3_u2725, p1_p3_u2724, p1_p3_u2723, p1_p3_u2722, p1_p3_u2721, p1_p3_u2720, p1_p3_u2719, p1_p3_u2718, p1_p3_u2717, p1_p3_u2716, p1_p3_u2715, p1_p3_u2714, p1_p3_u2713, p1_p3_u2712, p1_p3_u2711, p1_p3_u2710, p1_p3_u2709, p1_p3_u2708, p1_p3_u2707, p1_p3_u2706, p1_p3_u2705, p1_p3_u2704, p1_p3_u2703, p1_p3_u2702, p1_p3_u2701, p1_p3_u2700, p1_p3_u2699, p1_p3_u2698, p1_p3_u2697, p1_p3_u2696, p1_p3_u2695, p1_p3_u2694, p1_p3_u2693, p1_p3_u2692, p1_p3_u2691, p1_p3_u2690, p1_p3_u2689, p1_p3_u2688, p1_p3_u2687, p1_p3_u2686, p1_p3_u2685, p1_p3_u2684, p1_p3_u2683, p1_p3_u2682, p1_p3_u2681, p1_p3_u2680, p1_p3_u2679, p1_p3_u2678, p1_p3_u2677, p1_p3_u2676, p1_p3_u2675, p1_p3_u2674, p1_p3_u2673, p1_p3_u2672, p1_p3_u2671, p1_p3_u2670, p1_p3_u2669, p1_p3_u2668, p1_p3_u2667, p1_p3_u2666, p1_p3_u2665, p1_p3_u2664, p1_p3_u2663, p1_p3_u2662, p1_p3_u2661, p1_p3_u2660, p1_p3_u2659, p1_p3_u2658, p1_p3_u2657, p1_p3_u2656, p1_p3_u2655, p1_p3_u2654, p1_p3_u2653, p1_p3_u2652, p1_p3_u2651, p1_p3_u2650, p1_p3_u2649, p1_p3_u2648, p1_p3_u2647, p1_p3_u2646, p1_p3_u2645, p1_p3_u2644, p1_p3_u2643, p1_p3_u2642, p1_p3_u2641, p1_p3_u2640, p1_p3_u2639, p1_p3_u3292, p1_p3_u2638, p1_p3_u3293, p1_p3_u3294, p1_p3_u2637, p1_p3_u3295, p1_p3_u2636, p1_p3_u3296, p1_p3_u2635, p1_p3_u3297, p1_p3_u2634, p1_p3_u2633, p1_p3_u3298, p1_p3_u3299, p1_p2_u3274, p1_p2_u3275, p1_p2_u3276, p1_p2_u3277, p1_p2_u3061, p1_p2_u3060, p1_p2_u3059, p1_p2_u3058, p1_p2_u3057, p1_p2_u3056, p1_p2_u3055, p1_p2_u3054, p1_p2_u3053, p1_p2_u3052, p1_p2_u3051, p1_p2_u3050, p1_p2_u3049, p1_p2_u3048, p1_p2_u3047, p1_p2_u3046, p1_p2_u3045, p1_p2_u3044, p1_p2_u3043, p1_p2_u3042, p1_p2_u3041, p1_p2_u3040, p1_p2_u3039, p1_p2_u3038, p1_p2_u3037, p1_p2_u3036, p1_p2_u3035, p1_p2_u3034, p1_p2_u3033, p1_p2_u3032, p1_p2_u3031, p1_p2_u3030, p1_p2_u3029, p1_p2_u3280, p1_p2_u3281, p1_p2_u3028, p1_p2_u3027, p1_p2_u3026, p1_p2_u3025, p1_p2_u3024, p1_p2_u3023, p1_p2_u3022, p1_p2_u3021, p1_p2_u3020, p1_p2_u3019, p1_p2_u3018, p1_p2_u3017, p1_p2_u3016, p1_p2_u3015, p1_p2_u3014, p1_p2_u3013, p1_p2_u3012, p1_p2_u3011, p1_p2_u3010, p1_p2_u3009, p1_p2_u3008, p1_p2_u3007, p1_p2_u3006, p1_p2_u3005, p1_p2_u3004, p1_p2_u3003, p1_p2_u3002, p1_p2_u3001, p1_p2_u3000, p1_p2_u2999, p1_p2_u3282, p1_p2_u2998, p1_p2_u2997, p1_p2_u2996, p1_p2_u2995, p1_p2_u2994, p1_p2_u2993, p1_p2_u2992, p1_p2_u2991, p1_p2_u2990, p1_p2_u2989, p1_p2_u2988, p1_p2_u2987, p1_p2_u2986, p1_p2_u2985, p1_p2_u2984, p1_p2_u2983, p1_p2_u2982, p1_p2_u2981, p1_p2_u2980, p1_p2_u2979, p1_p2_u2978, p1_p2_u2977, p1_p2_u2976, p1_p2_u2975, p1_p2_u2974, p1_p2_u2973, p1_p2_u2972, p1_p2_u2971, p1_p2_u2970, p1_p2_u2969, p1_p2_u2968, p1_p2_u2967, p1_p2_u2966, p1_p2_u2965, p1_p2_u2964, p1_p2_u2963, p1_p2_u2962, p1_p2_u2961, p1_p2_u2960, p1_p2_u2959, p1_p2_u2958, p1_p2_u2957, p1_p2_u2956, p1_p2_u2955, p1_p2_u2954, p1_p2_u2953, p1_p2_u2952, p1_p2_u2951, p1_p2_u2950, p1_p2_u2949, p1_p2_u2948, p1_p2_u2947, p1_p2_u2946, p1_p2_u2945, p1_p2_u2944, p1_p2_u2943, p1_p2_u2942, p1_p2_u2941, p1_p2_u2940, p1_p2_u2939, p1_p2_u2938, p1_p2_u2937, p1_p2_u2936, p1_p2_u2935, p1_p2_u2934, p1_p2_u2933, p1_p2_u2932, p1_p2_u2931, p1_p2_u2930, p1_p2_u2929, p1_p2_u2928, p1_p2_u2927, p1_p2_u2926, p1_p2_u2925, p1_p2_u2924, p1_p2_u2923, p1_p2_u2922, p1_p2_u2921, p1_p2_u2920, p1_p2_u2919, p1_p2_u2918, p1_p2_u2917, p1_p2_u2916, p1_p2_u2915, p1_p2_u2914, p1_p2_u2913, p1_p2_u2912, p1_p2_u2911, p1_p2_u2910, p1_p2_u2909, p1_p2_u2908, p1_p2_u2907, p1_p2_u2906, p1_p2_u2905, p1_p2_u2904, p1_p2_u2903, p1_p2_u2902, p1_p2_u2901, p1_p2_u2900, p1_p2_u2899, p1_p2_u2898, p1_p2_u2897, p1_p2_u2896, p1_p2_u2895, p1_p2_u2894, p1_p2_u2893, p1_p2_u2892, p1_p2_u2891, p1_p2_u2890, p1_p2_u2889, p1_p2_u2888, p1_p2_u2887, p1_p2_u2886, p1_p2_u2885, p1_p2_u2884, p1_p2_u2883, p1_p2_u2882, p1_p2_u2881, p1_p2_u2880, p1_p2_u2879, p1_p2_u2878, p1_p2_u2877, p1_p2_u2876, p1_p2_u2875, p1_p2_u2874, p1_p2_u2873, p1_p2_u2872, p1_p2_u2871, p1_p2_u2870, p1_p2_u2869, p1_p2_u2868, p1_p2_u3284, p1_p2_u3285, p1_p2_u3288, p1_p2_u3289, p1_p2_u3290, p1_p2_u2867, p1_p2_u2866, p1_p2_u2865, p1_p2_u2864, p1_p2_u2863, p1_p2_u2862, p1_p2_u2861, p1_p2_u2860, p1_p2_u2859, p1_p2_u2858, p1_p2_u2857, p1_p2_u2856, p1_p2_u2855, p1_p2_u2854, p1_p2_u2853, p1_p2_u2852, p1_p2_u2851, p1_p2_u2850, p1_p2_u2849, p1_p2_u2848, p1_p2_u2847, p1_p2_u2846, p1_p2_u2845, p1_p2_u2844, p1_p2_u2843, p1_p2_u2842, p1_p2_u2841, p1_p2_u2840, p1_p2_u2839, p1_p2_u2838, p1_p2_u2837, p1_p2_u2836, p1_p2_u2835, p1_p2_u2834, p1_p2_u2833, p1_p2_u2832, p1_p2_u2831, p1_p2_u2830, p1_p2_u2829, p1_p2_u2828, p1_p2_u2827, p1_p2_u2826, p1_p2_u2825, p1_p2_u2824, p1_p2_u2823, p1_p2_u2822, p1_p2_u2821, p1_p2_u2820, p1_p2_u2819, p1_p2_u2818, p1_p2_u2817, p1_p2_u2816, p1_p2_u2815, p1_p2_u2814, p1_p2_u2813, p1_p2_u2812, p1_p2_u2811, p1_p2_u2810, p1_p2_u2809, p1_p2_u2808, p1_p2_u2807, p1_p2_u2806, p1_p2_u2805, p1_p2_u2804, p1_p2_u2803, p1_p2_u2802, p1_p2_u2801, p1_p2_u2800, p1_p2_u2799, p1_p2_u2798, p1_p2_u2797, p1_p2_u2796, p1_p2_u2795, p1_p2_u2794, p1_p2_u2793, p1_p2_u2792, p1_p2_u2791, p1_p2_u2790, p1_p2_u2789, p1_p2_u2788, p1_p2_u2787, p1_p2_u2786, p1_p2_u2785, p1_p2_u2784, p1_p2_u2783, p1_p2_u2782, p1_p2_u2781, p1_p2_u2780, p1_p2_u2779, p1_p2_u2778, p1_p2_u2777, p1_p2_u2776, p1_p2_u2775, p1_p2_u2774, p1_p2_u2773, p1_p2_u2772, p1_p2_u2771, p1_p2_u2770, p1_p2_u2769, p1_p2_u2768, p1_p2_u2767, p1_p2_u2766, p1_p2_u2765, p1_p2_u2764, p1_p2_u2763, p1_p2_u2762, p1_p2_u2761, p1_p2_u2760, p1_p2_u2759, p1_p2_u2758, p1_p2_u2757, p1_p2_u2756, p1_p2_u2755, p1_p2_u2754, p1_p2_u2753, p1_p2_u2752, p1_p2_u2751, p1_p2_u2750, p1_p2_u2749, p1_p2_u2748, p1_p2_u2747, p1_p2_u2746, p1_p2_u2745, p1_p2_u2744, p1_p2_u2743, p1_p2_u2742, p1_p2_u2741, p1_p2_u2740, p1_p2_u2739, p1_p2_u2738, p1_p2_u2737, p1_p2_u2736, p1_p2_u2735, p1_p2_u2734, p1_p2_u2733, p1_p2_u2732, p1_p2_u2731, p1_p2_u2730, p1_p2_u2729, p1_p2_u2728, p1_p2_u2727, p1_p2_u2726, p1_p2_u2725, p1_p2_u2724, p1_p2_u2723, p1_p2_u2722, p1_p2_u2721, p1_p2_u2720, p1_p2_u2719, p1_p2_u2718, p1_p2_u2717, p1_p2_u2716, p1_p2_u2715, p1_p2_u2714, p1_p2_u2713, p1_p2_u2712, p1_p2_u2711, p1_p2_u2710, p1_p2_u2709, p1_p2_u2708, p1_p2_u2707, p1_p2_u2706, p1_p2_u2705, p1_p2_u2704, p1_p2_u2703, p1_p2_u2702, p1_p2_u2701, p1_p2_u2700, p1_p2_u2699, p1_p2_u2698, p1_p2_u2697, p1_p2_u2696, p1_p2_u2695, p1_p2_u2694, p1_p2_u2693, p1_p2_u2692, p1_p2_u2691, p1_p2_u2690, p1_p2_u2689, p1_p2_u2688, p1_p2_u2687, p1_p2_u2686, p1_p2_u2685, p1_p2_u2684, p1_p2_u2683, p1_p2_u2682, p1_p2_u2681, p1_p2_u2680, p1_p2_u2679, p1_p2_u2678, p1_p2_u2677, p1_p2_u2676, p1_p2_u2675, p1_p2_u2674, p1_p2_u2673, p1_p2_u2672, p1_p2_u2671, p1_p2_u2670, p1_p2_u2669, p1_p2_u2668, p1_p2_u2667, p1_p2_u2666, p1_p2_u2665, p1_p2_u2664, p1_p2_u2663, p1_p2_u2662, p1_p2_u2661, p1_p2_u2660, p1_p2_u2659, p1_p2_u2658, p1_p2_u2657, p1_p2_u2656, p1_p2_u2655, p1_p2_u2654, p1_p2_u2653, p1_p2_u2652, p1_p2_u2651, p1_p2_u2650, p1_p2_u2649, p1_p2_u2648, p1_p2_u2647, p1_p2_u2646, p1_p2_u2645, p1_p2_u2644, p1_p2_u2643, p1_p2_u2642, p1_p2_u2641, p1_p2_u2640, p1_p2_u2639, p1_p2_u3292, p1_p2_u2638, p1_p2_u3293, p1_p2_u3294, p1_p2_u2637, p1_p2_u3295, p1_p2_u2636, p1_p2_u3296, p1_p2_u2635, p1_p2_u3297, p1_p2_u2634, p1_p2_u2633, p1_p2_u3298, p1_p2_u3299, p1_p1_u3288, p1_p1_u3289, p1_p1_u3290, p1_p1_u3291, p1_p1_u3077, p1_p1_u3076, p1_p1_u3075, p1_p1_u3074, p1_p1_u3073, p1_p1_u3072, p1_p1_u3071, p1_p1_u3070, p1_p1_u3069, p1_p1_u3068, p1_p1_u3067, p1_p1_u3066, p1_p1_u3065, p1_p1_u3064, p1_p1_u3063, p1_p1_u3062, p1_p1_u3061, p1_p1_u3060, p1_p1_u3059, p1_p1_u3058, p1_p1_u3057, p1_p1_u3056, p1_p1_u3055, p1_p1_u3054, p1_p1_u3053, p1_p1_u3052, p1_p1_u3051, p1_p1_u3050, p1_p1_u3049, p1_p1_u3048, p1_p1_u3047, p1_p1_u3046, p1_p1_u3045, p1_p1_u3294, p1_p1_u3295, p1_p1_u3044, p1_p1_u3043, p1_p1_u3042, p1_p1_u3041, p1_p1_u3040, p1_p1_u3039, p1_p1_u3038, p1_p1_u3037, p1_p1_u3036, p1_p1_u3035, p1_p1_u3034, p1_p1_u3033, p1_p1_u3032, p1_p1_u3031, p1_p1_u3030, p1_p1_u3029, p1_p1_u3028, p1_p1_u3027, p1_p1_u3026, p1_p1_u3025, p1_p1_u3024, p1_p1_u3023, p1_p1_u3022, p1_p1_u3021, p1_p1_u3020, p1_p1_u3019, p1_p1_u3018, p1_p1_u3017, p1_p1_u3016, p1_p1_u3015, p1_p1_u3296, p1_p1_u3014, p1_p1_u3013, p1_p1_u3012, p1_p1_u3011, p1_p1_u3010, p1_p1_u3009, p1_p1_u3008, p1_p1_u3007, p1_p1_u3006, p1_p1_u3005, p1_p1_u3004, p1_p1_u3003, p1_p1_u3002, p1_p1_u3001, p1_p1_u3000, p1_p1_u2999, p1_p1_u2998, p1_p1_u2997, p1_p1_u2996, p1_p1_u2995, p1_p1_u2994, p1_p1_u2993, p1_p1_u2992, p1_p1_u2991, p1_p1_u2990, p1_p1_u2989, p1_p1_u2988, p1_p1_u2987, p1_p1_u2986, p1_p1_u2985, p1_p1_u2984, p1_p1_u2983, p1_p1_u2982, p1_p1_u2981, p1_p1_u2980, p1_p1_u2979, p1_p1_u2978, p1_p1_u2977, p1_p1_u2976, p1_p1_u2975, p1_p1_u2974, p1_p1_u2973, p1_p1_u2972, p1_p1_u2971, p1_p1_u2970, p1_p1_u2969, p1_p1_u2968, p1_p1_u2967, p1_p1_u2966, p1_p1_u2965, p1_p1_u2964, p1_p1_u2963, p1_p1_u2962, p1_p1_u2961, p1_p1_u2960, p1_p1_u2959, p1_p1_u2958, p1_p1_u2957, p1_p1_u2956, p1_p1_u2955, p1_p1_u2954, p1_p1_u2953, p1_p1_u2952, p1_p1_u2951, p1_p1_u2950, p1_p1_u2949, p1_p1_u2948, p1_p1_u2947, p1_p1_u2946, p1_p1_u2945, p1_p1_u2944, p1_p1_u2943, p1_p1_u2942, p1_p1_u2941, p1_p1_u2940, p1_p1_u2939, p1_p1_u2938, p1_p1_u2937, p1_p1_u2936, p1_p1_u2935, p1_p1_u2934, p1_p1_u2933, p1_p1_u2932, p1_p1_u2931, p1_p1_u2930, p1_p1_u2929, p1_p1_u2928, p1_p1_u2927, p1_p1_u2926, p1_p1_u2925, p1_p1_u2924, p1_p1_u2923, p1_p1_u2922, p1_p1_u2921, p1_p1_u2920, p1_p1_u2919, p1_p1_u2918, p1_p1_u2917, p1_p1_u2916, p1_p1_u2915, p1_p1_u2914, p1_p1_u2913, p1_p1_u2912, p1_p1_u2911, p1_p1_u2910, p1_p1_u2909, p1_p1_u2908, p1_p1_u2907, p1_p1_u2906, p1_p1_u2905, p1_p1_u2904, p1_p1_u2903, p1_p1_u2902, p1_p1_u2901, p1_p1_u2900, p1_p1_u2899, p1_p1_u2898, p1_p1_u2897, p1_p1_u2896, p1_p1_u2895, p1_p1_u2894, p1_p1_u2893, p1_p1_u2892, p1_p1_u2891, p1_p1_u2890, p1_p1_u2889, p1_p1_u2888, p1_p1_u2887, p1_p1_u2886, p1_p1_u2885, p1_p1_u2884, p1_p1_u3298, p1_p1_u3299, p1_p1_u3302, p1_p1_u3303, p1_p1_u3304, p1_p1_u2883, p1_p1_u2882, p1_p1_u2881, p1_p1_u2880, p1_p1_u2879, p1_p1_u2878, p1_p1_u2877, p1_p1_u2876, p1_p1_u2875, p1_p1_u2874, p1_p1_u2873, p1_p1_u2872, p1_p1_u2871, p1_p1_u2870, p1_p1_u2869, p1_p1_u2868, p1_p1_u2867, p1_p1_u2866, p1_p1_u2865, p1_p1_u2864, p1_p1_u2863, p1_p1_u2862, p1_p1_u2861, p1_p1_u2860, p1_p1_u2859, p1_p1_u2858, p1_p1_u2857, p1_p1_u2856, p1_p1_u2855, p1_p1_u2854, p1_p1_u2853, p1_p1_u2852, p1_p1_u2851, p1_p1_u2850, p1_p1_u2849, p1_p1_u2848, p1_p1_u2847, p1_p1_u2846, p1_p1_u2845, p1_p1_u2844, p1_p1_u2843, p1_p1_u2842, p1_p1_u2841, p1_p1_u2840, p1_p1_u2839, p1_p1_u2838, p1_p1_u2837, p1_p1_u2836, p1_p1_u2835, p1_p1_u2834, p1_p1_u2833, p1_p1_u2832, p1_p1_u2831, p1_p1_u2830, p1_p1_u2829, p1_p1_u2828, p1_p1_u2827, p1_p1_u2826, p1_p1_u2825, p1_p1_u2824, p1_p1_u2823, p1_p1_u2822, p1_p1_u2821, p1_p1_u2820, p1_p1_u2819, p1_p1_u2818, p1_p1_u2817, p1_p1_u2816, p1_p1_u2815, p1_p1_u2814, p1_p1_u2813, p1_p1_u2812, p1_p1_u2811, p1_p1_u2810, p1_p1_u2809, p1_p1_u2808, p1_p1_u2807, p1_p1_u2806, p1_p1_u2805, p1_p1_u2804, p1_p1_u2803, p1_p1_u2802, p1_p1_u2801, p1_p1_u2800, p1_p1_u2799, p1_p1_u2798, p1_p1_u2797, p1_p1_u2796, p1_p1_u2795, p1_p1_u2794, p1_p1_u2793, p1_p1_u2792, p1_p1_u2791, p1_p1_u2790, p1_p1_u2789, p1_p1_u2788, p1_p1_u2787, p1_p1_u2786, p1_p1_u2785, p1_p1_u2784, p1_p1_u2783, p1_p1_u2782, p1_p1_u2781, p1_p1_u2780, p1_p1_u2779, p1_p1_u2778, p1_p1_u2777, p1_p1_u2776, p1_p1_u2775, p1_p1_u2774, p1_p1_u2773, p1_p1_u2772, p1_p1_u2771, p1_p1_u2770, p1_p1_u2769, p1_p1_u2768, p1_p1_u2767, p1_p1_u2766, p1_p1_u2765, p1_p1_u2764, p1_p1_u2763, p1_p1_u2762, p1_p1_u2761, p1_p1_u2760, p1_p1_u2759, p1_p1_u2758, p1_p1_u2757, p1_p1_u2756, p1_p1_u2755, p1_p1_u2754, p1_p1_u2753, p1_p1_u2752, p1_p1_u2751, p1_p1_u2750, p1_p1_u2749, p1_p1_u2748, p1_p1_u2747, p1_p1_u2746, p1_p1_u2745, p1_p1_u2744, p1_p1_u2743, p1_p1_u2742, p1_p1_u2741, p1_p1_u2740, p1_p1_u2739, p1_p1_u2738, p1_p1_u2737, p1_p1_u2736, p1_p1_u2735, p1_p1_u2734, p1_p1_u2733, p1_p1_u2732, p1_p1_u2731, p1_p1_u2730, p1_p1_u2729, p1_p1_u2728, p1_p1_u2727, p1_p1_u2726, p1_p1_u2725, p1_p1_u2724, p1_p1_u2723, p1_p1_u2722, p1_p1_u2721, p1_p1_u2720, p1_p1_u2719, p1_p1_u2718, p1_p1_u2717, p1_p1_u2716, p1_p1_u2715, p1_p1_u2714, p1_p1_u2713, p1_p1_u2712, p1_p1_u2711, p1_p1_u2710, p1_p1_u2709, p1_p1_u2708, p1_p1_u2707, p1_p1_u2706, p1_p1_u2705, p1_p1_u2704, p1_p1_u2703, p1_p1_u2702, p1_p1_u2701, p1_p1_u2700, p1_p1_u2699, p1_p1_u2698, p1_p1_u2697, p1_p1_u2696, p1_p1_u2695, p1_p1_u2694, p1_p1_u2693, p1_p1_u2692, p1_p1_u2691, p1_p1_u2690, p1_p1_u2689, p1_p1_u2688, p1_p1_u2687, p1_p1_u2686, p1_p1_u2685, p1_p1_u2684, p1_p1_u2683, p1_p1_u2682, p1_p1_u2681, p1_p1_u2680, p1_p1_u2679, p1_p1_u2678, p1_p1_u2677, p1_p1_u2676, p1_p1_u2675, p1_p1_u2674, p1_p1_u2673, p1_p1_u2672, p1_p1_u2671, p1_p1_u2670, p1_p1_u2669, p1_p1_u2668, p1_p1_u2667, p1_p1_u2666, p1_p1_u2665, p1_p1_u2664, p1_p1_u2663, p1_p1_u2662, p1_p1_u2661, p1_p1_u2660, p1_p1_u2659, p1_p1_u2658, p1_p1_u2657, p1_p1_u2656, p1_p1_u2655, p1_p1_u3306, p1_p1_u2654, p1_p1_u3307, p1_p1_u3308, p1_p1_u2653, p1_p1_u3309, p1_p1_u2652, p1_p1_u3310, p1_p1_u2651, p1_p1_u3311, p1_p1_u2650, p1_p1_u2649, p1_p1_u3312, p1_p1_u3313, p2_p3_u3274, p2_p3_u3275, p2_p3_u3276, p2_p3_u3277, p2_p3_u3061, p2_p3_u3060, p2_p3_u3059, p2_p3_u3058, p2_p3_u3057, p2_p3_u3056, p2_p3_u3055, p2_p3_u3054, p2_p3_u3053, p2_p3_u3052, p2_p3_u3051, p2_p3_u3050, p2_p3_u3049, p2_p3_u3048, p2_p3_u3047, p2_p3_u3046, p2_p3_u3045, p2_p3_u3044, p2_p3_u3043, p2_p3_u3042, p2_p3_u3041, p2_p3_u3040, p2_p3_u3039, p2_p3_u3038, p2_p3_u3037, p2_p3_u3036, p2_p3_u3035, p2_p3_u3034, p2_p3_u3033, p2_p3_u3032, p2_p3_u3031, p2_p3_u3030, p2_p3_u3029, p2_p3_u3280, p2_p3_u3281, p2_p3_u3028, p2_p3_u3027, p2_p3_u3026, p2_p3_u3025, p2_p3_u3024, p2_p3_u3023, p2_p3_u3022, p2_p3_u3021, p2_p3_u3020, p2_p3_u3019, p2_p3_u3018, p2_p3_u3017, p2_p3_u3016, p2_p3_u3015, p2_p3_u3014, p2_p3_u3013, p2_p3_u3012, p2_p3_u3011, p2_p3_u3010, p2_p3_u3009, p2_p3_u3008, p2_p3_u3007, p2_p3_u3006, p2_p3_u3005, p2_p3_u3004, p2_p3_u3003, p2_p3_u3002, p2_p3_u3001, p2_p3_u3000, p2_p3_u2999, p2_p3_u3282, p2_p3_u2998, p2_p3_u2997, p2_p3_u2996, p2_p3_u2995, p2_p3_u2994, p2_p3_u2993, p2_p3_u2992, p2_p3_u2991, p2_p3_u2990, p2_p3_u2989, p2_p3_u2988, p2_p3_u2987, p2_p3_u2986, p2_p3_u2985, p2_p3_u2984, p2_p3_u2983, p2_p3_u2982, p2_p3_u2981, p2_p3_u2980, p2_p3_u2979, p2_p3_u2978, p2_p3_u2977, p2_p3_u2976, p2_p3_u2975, p2_p3_u2974, p2_p3_u2973, p2_p3_u2972, p2_p3_u2971, p2_p3_u2970, p2_p3_u2969, p2_p3_u2968, p2_p3_u2967, p2_p3_u2966, p2_p3_u2965, p2_p3_u2964, p2_p3_u2963, p2_p3_u2962, p2_p3_u2961, p2_p3_u2960, p2_p3_u2959, p2_p3_u2958, p2_p3_u2957, p2_p3_u2956, p2_p3_u2955, p2_p3_u2954, p2_p3_u2953, p2_p3_u2952, p2_p3_u2951, p2_p3_u2950, p2_p3_u2949, p2_p3_u2948, p2_p3_u2947, p2_p3_u2946, p2_p3_u2945, p2_p3_u2944, p2_p3_u2943, p2_p3_u2942, p2_p3_u2941, p2_p3_u2940, p2_p3_u2939, p2_p3_u2938, p2_p3_u2937, p2_p3_u2936, p2_p3_u2935, p2_p3_u2934, p2_p3_u2933, p2_p3_u2932, p2_p3_u2931, p2_p3_u2930, p2_p3_u2929, p2_p3_u2928, p2_p3_u2927, p2_p3_u2926, p2_p3_u2925, p2_p3_u2924, p2_p3_u2923, p2_p3_u2922, p2_p3_u2921, p2_p3_u2920, p2_p3_u2919, p2_p3_u2918, p2_p3_u2917, p2_p3_u2916, p2_p3_u2915, p2_p3_u2914, p2_p3_u2913, p2_p3_u2912, p2_p3_u2911, p2_p3_u2910, p2_p3_u2909, p2_p3_u2908, p2_p3_u2907, p2_p3_u2906, p2_p3_u2905, p2_p3_u2904, p2_p3_u2903, p2_p3_u2902, p2_p3_u2901, p2_p3_u2900, p2_p3_u2899, p2_p3_u2898, p2_p3_u2897, p2_p3_u2896, p2_p3_u2895, p2_p3_u2894, p2_p3_u2893, p2_p3_u2892, p2_p3_u2891, p2_p3_u2890, p2_p3_u2889, p2_p3_u2888, p2_p3_u2887, p2_p3_u2886, p2_p3_u2885, p2_p3_u2884, p2_p3_u2883, p2_p3_u2882, p2_p3_u2881, p2_p3_u2880, p2_p3_u2879, p2_p3_u2878, p2_p3_u2877, p2_p3_u2876, p2_p3_u2875, p2_p3_u2874, p2_p3_u2873, p2_p3_u2872, p2_p3_u2871, p2_p3_u2870, p2_p3_u2869, p2_p3_u2868, p2_p3_u3284, p2_p3_u3285, p2_p3_u3288, p2_p3_u3289, p2_p3_u3290, p2_p3_u2867, p2_p3_u2866, p2_p3_u2865, p2_p3_u2864, p2_p3_u2863, p2_p3_u2862, p2_p3_u2861, p2_p3_u2860, p2_p3_u2859, p2_p3_u2858, p2_p3_u2857, p2_p3_u2856, p2_p3_u2855, p2_p3_u2854, p2_p3_u2853, p2_p3_u2852, p2_p3_u2851, p2_p3_u2850, p2_p3_u2849, p2_p3_u2848, p2_p3_u2847, p2_p3_u2846, p2_p3_u2845, p2_p3_u2844, p2_p3_u2843, p2_p3_u2842, p2_p3_u2841, p2_p3_u2840, p2_p3_u2839, p2_p3_u2838, p2_p3_u2837, p2_p3_u2836, p2_p3_u2835, p2_p3_u2834, p2_p3_u2833, p2_p3_u2832, p2_p3_u2831, p2_p3_u2830, p2_p3_u2829, p2_p3_u2828, p2_p3_u2827, p2_p3_u2826, p2_p3_u2825, p2_p3_u2824, p2_p3_u2823, p2_p3_u2822, p2_p3_u2821, p2_p3_u2820, p2_p3_u2819, p2_p3_u2818, p2_p3_u2817, p2_p3_u2816, p2_p3_u2815, p2_p3_u2814, p2_p3_u2813, p2_p3_u2812, p2_p3_u2811, p2_p3_u2810, p2_p3_u2809, p2_p3_u2808, p2_p3_u2807, p2_p3_u2806, p2_p3_u2805, p2_p3_u2804, p2_p3_u2803, p2_p3_u2802, p2_p3_u2801, p2_p3_u2800, p2_p3_u2799, p2_p3_u2798, p2_p3_u2797, p2_p3_u2796, p2_p3_u2795, p2_p3_u2794, p2_p3_u2793, p2_p3_u2792, p2_p3_u2791, p2_p3_u2790, p2_p3_u2789, p2_p3_u2788, p2_p3_u2787, p2_p3_u2786, p2_p3_u2785, p2_p3_u2784, p2_p3_u2783, p2_p3_u2782, p2_p3_u2781, p2_p3_u2780, p2_p3_u2779, p2_p3_u2778, p2_p3_u2777, p2_p3_u2776, p2_p3_u2775, p2_p3_u2774, p2_p3_u2773, p2_p3_u2772, p2_p3_u2771, p2_p3_u2770, p2_p3_u2769, p2_p3_u2768, p2_p3_u2767, p2_p3_u2766, p2_p3_u2765, p2_p3_u2764, p2_p3_u2763, p2_p3_u2762, p2_p3_u2761, p2_p3_u2760, p2_p3_u2759, p2_p3_u2758, p2_p3_u2757, p2_p3_u2756, p2_p3_u2755, p2_p3_u2754, p2_p3_u2753, p2_p3_u2752, p2_p3_u2751, p2_p3_u2750, p2_p3_u2749, p2_p3_u2748, p2_p3_u2747, p2_p3_u2746, p2_p3_u2745, p2_p3_u2744, p2_p3_u2743, p2_p3_u2742, p2_p3_u2741, p2_p3_u2740, p2_p3_u2739, p2_p3_u2738, p2_p3_u2737, p2_p3_u2736, p2_p3_u2735, p2_p3_u2734, p2_p3_u2733, p2_p3_u2732, p2_p3_u2731, p2_p3_u2730, p2_p3_u2729, p2_p3_u2728, p2_p3_u2727, p2_p3_u2726, p2_p3_u2725, p2_p3_u2724, p2_p3_u2723, p2_p3_u2722, p2_p3_u2721, p2_p3_u2720, p2_p3_u2719, p2_p3_u2718, p2_p3_u2717, p2_p3_u2716, p2_p3_u2715, p2_p3_u2714, p2_p3_u2713, p2_p3_u2712, p2_p3_u2711, p2_p3_u2710, p2_p3_u2709, p2_p3_u2708, p2_p3_u2707, p2_p3_u2706, p2_p3_u2705, p2_p3_u2704, p2_p3_u2703, p2_p3_u2702, p2_p3_u2701, p2_p3_u2700, p2_p3_u2699, p2_p3_u2698, p2_p3_u2697, p2_p3_u2696, p2_p3_u2695, p2_p3_u2694, p2_p3_u2693, p2_p3_u2692, p2_p3_u2691, p2_p3_u2690, p2_p3_u2689, p2_p3_u2688, p2_p3_u2687, p2_p3_u2686, p2_p3_u2685, p2_p3_u2684, p2_p3_u2683, p2_p3_u2682, p2_p3_u2681, p2_p3_u2680, p2_p3_u2679, p2_p3_u2678, p2_p3_u2677, p2_p3_u2676, p2_p3_u2675, p2_p3_u2674, p2_p3_u2673, p2_p3_u2672, p2_p3_u2671, p2_p3_u2670, p2_p3_u2669, p2_p3_u2668, p2_p3_u2667, p2_p3_u2666, p2_p3_u2665, p2_p3_u2664, p2_p3_u2663, p2_p3_u2662, p2_p3_u2661, p2_p3_u2660, p2_p3_u2659, p2_p3_u2658, p2_p3_u2657, p2_p3_u2656, p2_p3_u2655, p2_p3_u2654, p2_p3_u2653, p2_p3_u2652, p2_p3_u2651, p2_p3_u2650, p2_p3_u2649, p2_p3_u2648, p2_p3_u2647, p2_p3_u2646, p2_p3_u2645, p2_p3_u2644, p2_p3_u2643, p2_p3_u2642, p2_p3_u2641, p2_p3_u2640, p2_p3_u2639, p2_p3_u3292, p2_p3_u2638, p2_p3_u3293, p2_p3_u3294, p2_p3_u2637, p2_p3_u3295, p2_p3_u2636, p2_p3_u3296, p2_p3_u2635, p2_p3_u3297, p2_p3_u2634, p2_p3_u2633, p2_p3_u3298, p2_p3_u3299, p2_p2_u3274, p2_p2_u3275, p2_p2_u3276, p2_p2_u3277, p2_p2_u3061, p2_p2_u3060, p2_p2_u3059, p2_p2_u3058, p2_p2_u3057, p2_p2_u3056, p2_p2_u3055, p2_p2_u3054, p2_p2_u3053, p2_p2_u3052, p2_p2_u3051, p2_p2_u3050, p2_p2_u3049, p2_p2_u3048, p2_p2_u3047, p2_p2_u3046, p2_p2_u3045, p2_p2_u3044, p2_p2_u3043, p2_p2_u3042, p2_p2_u3041, p2_p2_u3040, p2_p2_u3039, p2_p2_u3038, p2_p2_u3037, p2_p2_u3036, p2_p2_u3035, p2_p2_u3034, p2_p2_u3033, p2_p2_u3032, p2_p2_u3031, p2_p2_u3030, p2_p2_u3029, p2_p2_u3280, p2_p2_u3281, p2_p2_u3028, p2_p2_u3027, p2_p2_u3026, p2_p2_u3025, p2_p2_u3024, p2_p2_u3023, p2_p2_u3022, p2_p2_u3021, p2_p2_u3020, p2_p2_u3019, p2_p2_u3018, p2_p2_u3017, p2_p2_u3016, p2_p2_u3015, p2_p2_u3014, p2_p2_u3013, p2_p2_u3012, p2_p2_u3011, p2_p2_u3010, p2_p2_u3009, p2_p2_u3008, p2_p2_u3007, p2_p2_u3006, p2_p2_u3005, p2_p2_u3004, p2_p2_u3003, p2_p2_u3002, p2_p2_u3001, p2_p2_u3000, p2_p2_u2999, p2_p2_u3282, p2_p2_u2998, p2_p2_u2997, p2_p2_u2996, p2_p2_u2995, p2_p2_u2994, p2_p2_u2993, p2_p2_u2992, p2_p2_u2991, p2_p2_u2990, p2_p2_u2989, p2_p2_u2988, p2_p2_u2987, p2_p2_u2986, p2_p2_u2985, p2_p2_u2984, p2_p2_u2983, p2_p2_u2982, p2_p2_u2981, p2_p2_u2980, p2_p2_u2979, p2_p2_u2978, p2_p2_u2977, p2_p2_u2976, p2_p2_u2975, p2_p2_u2974, p2_p2_u2973, p2_p2_u2972, p2_p2_u2971, p2_p2_u2970, p2_p2_u2969, p2_p2_u2968, p2_p2_u2967, p2_p2_u2966, p2_p2_u2965, p2_p2_u2964, p2_p2_u2963, p2_p2_u2962, p2_p2_u2961, p2_p2_u2960, p2_p2_u2959, p2_p2_u2958, p2_p2_u2957, p2_p2_u2956, p2_p2_u2955, p2_p2_u2954, p2_p2_u2953, p2_p2_u2952, p2_p2_u2951, p2_p2_u2950, p2_p2_u2949, p2_p2_u2948, p2_p2_u2947, p2_p2_u2946, p2_p2_u2945, p2_p2_u2944, p2_p2_u2943, p2_p2_u2942, p2_p2_u2941, p2_p2_u2940, p2_p2_u2939, p2_p2_u2938, p2_p2_u2937, p2_p2_u2936, p2_p2_u2935, p2_p2_u2934, p2_p2_u2933, p2_p2_u2932, p2_p2_u2931, p2_p2_u2930, p2_p2_u2929, p2_p2_u2928, p2_p2_u2927, p2_p2_u2926, p2_p2_u2925, p2_p2_u2924, p2_p2_u2923, p2_p2_u2922, p2_p2_u2921, p2_p2_u2920, p2_p2_u2919, p2_p2_u2918, p2_p2_u2917, p2_p2_u2916, p2_p2_u2915, p2_p2_u2914, p2_p2_u2913, p2_p2_u2912, p2_p2_u2911, p2_p2_u2910, p2_p2_u2909, p2_p2_u2908, p2_p2_u2907, p2_p2_u2906, p2_p2_u2905, p2_p2_u2904, p2_p2_u2903, p2_p2_u2902, p2_p2_u2901, p2_p2_u2900, p2_p2_u2899, p2_p2_u2898, p2_p2_u2897, p2_p2_u2896, p2_p2_u2895, p2_p2_u2894, p2_p2_u2893, p2_p2_u2892, p2_p2_u2891, p2_p2_u2890, p2_p2_u2889, p2_p2_u2888, p2_p2_u2887, p2_p2_u2886, p2_p2_u2885, p2_p2_u2884, p2_p2_u2883, p2_p2_u2882, p2_p2_u2881, p2_p2_u2880, p2_p2_u2879, p2_p2_u2878, p2_p2_u2877, p2_p2_u2876, p2_p2_u2875, p2_p2_u2874, p2_p2_u2873, p2_p2_u2872, p2_p2_u2871, p2_p2_u2870, p2_p2_u2869, p2_p2_u2868, p2_p2_u3284, p2_p2_u3285, p2_p2_u3288, p2_p2_u3289, p2_p2_u3290, p2_p2_u2867, p2_p2_u2866, p2_p2_u2865, p2_p2_u2864, p2_p2_u2863, p2_p2_u2862, p2_p2_u2861, p2_p2_u2860, p2_p2_u2859, p2_p2_u2858, p2_p2_u2857, p2_p2_u2856, p2_p2_u2855, p2_p2_u2854, p2_p2_u2853, p2_p2_u2852, p2_p2_u2851, p2_p2_u2850, p2_p2_u2849, p2_p2_u2848, p2_p2_u2847, p2_p2_u2846, p2_p2_u2845, p2_p2_u2844, p2_p2_u2843, p2_p2_u2842, p2_p2_u2841, p2_p2_u2840, p2_p2_u2839, p2_p2_u2838, p2_p2_u2837, p2_p2_u2836, p2_p2_u2835, p2_p2_u2834, p2_p2_u2833, p2_p2_u2832, p2_p2_u2831, p2_p2_u2830, p2_p2_u2829, p2_p2_u2828, p2_p2_u2827, p2_p2_u2826, p2_p2_u2825, p2_p2_u2824, p2_p2_u2823, p2_p2_u2822, p2_p2_u2821, p2_p2_u2820, p2_p2_u2819, p2_p2_u2818, p2_p2_u2817, p2_p2_u2816, p2_p2_u2815, p2_p2_u2814, p2_p2_u2813, p2_p2_u2812, p2_p2_u2811, p2_p2_u2810, p2_p2_u2809, p2_p2_u2808, p2_p2_u2807, p2_p2_u2806, p2_p2_u2805, p2_p2_u2804, p2_p2_u2803, p2_p2_u2802, p2_p2_u2801, p2_p2_u2800, p2_p2_u2799, p2_p2_u2798, p2_p2_u2797, p2_p2_u2796, p2_p2_u2795, p2_p2_u2794, p2_p2_u2793, p2_p2_u2792, p2_p2_u2791, p2_p2_u2790, p2_p2_u2789, p2_p2_u2788, p2_p2_u2787, p2_p2_u2786, p2_p2_u2785, p2_p2_u2784, p2_p2_u2783, p2_p2_u2782, p2_p2_u2781, p2_p2_u2780, p2_p2_u2779, p2_p2_u2778, p2_p2_u2777, p2_p2_u2776, p2_p2_u2775, p2_p2_u2774, p2_p2_u2773, p2_p2_u2772, p2_p2_u2771, p2_p2_u2770, p2_p2_u2769, p2_p2_u2768, p2_p2_u2767, p2_p2_u2766, p2_p2_u2765, p2_p2_u2764, p2_p2_u2763, p2_p2_u2762, p2_p2_u2761, p2_p2_u2760, p2_p2_u2759, p2_p2_u2758, p2_p2_u2757, p2_p2_u2756, p2_p2_u2755, p2_p2_u2754, p2_p2_u2753, p2_p2_u2752, p2_p2_u2751, p2_p2_u2750, p2_p2_u2749, p2_p2_u2748, p2_p2_u2747, p2_p2_u2746, p2_p2_u2745, p2_p2_u2744, p2_p2_u2743, p2_p2_u2742, p2_p2_u2741, p2_p2_u2740, p2_p2_u2739, p2_p2_u2738, p2_p2_u2737, p2_p2_u2736, p2_p2_u2735, p2_p2_u2734, p2_p2_u2733, p2_p2_u2732, p2_p2_u2731, p2_p2_u2730, p2_p2_u2729, p2_p2_u2728, p2_p2_u2727, p2_p2_u2726, p2_p2_u2725, p2_p2_u2724, p2_p2_u2723, p2_p2_u2722, p2_p2_u2721, p2_p2_u2720, p2_p2_u2719, p2_p2_u2718, p2_p2_u2717, p2_p2_u2716, p2_p2_u2715, p2_p2_u2714, p2_p2_u2713, p2_p2_u2712, p2_p2_u2711, p2_p2_u2710, p2_p2_u2709, p2_p2_u2708, p2_p2_u2707, p2_p2_u2706, p2_p2_u2705, p2_p2_u2704, p2_p2_u2703, p2_p2_u2702, p2_p2_u2701, p2_p2_u2700, p2_p2_u2699, p2_p2_u2698, p2_p2_u2697, p2_p2_u2696, p2_p2_u2695, p2_p2_u2694, p2_p2_u2693, p2_p2_u2692, p2_p2_u2691, p2_p2_u2690, p2_p2_u2689, p2_p2_u2688, p2_p2_u2687, p2_p2_u2686, p2_p2_u2685, p2_p2_u2684, p2_p2_u2683, p2_p2_u2682, p2_p2_u2681, p2_p2_u2680, p2_p2_u2679, p2_p2_u2678, p2_p2_u2677, p2_p2_u2676, p2_p2_u2675, p2_p2_u2674, p2_p2_u2673, p2_p2_u2672, p2_p2_u2671, p2_p2_u2670, p2_p2_u2669, p2_p2_u2668, p2_p2_u2667, p2_p2_u2666, p2_p2_u2665, p2_p2_u2664, p2_p2_u2663, p2_p2_u2662, p2_p2_u2661, p2_p2_u2660, p2_p2_u2659, p2_p2_u2658, p2_p2_u2657, p2_p2_u2656, p2_p2_u2655, p2_p2_u2654, p2_p2_u2653, p2_p2_u2652, p2_p2_u2651, p2_p2_u2650, p2_p2_u2649, p2_p2_u2648, p2_p2_u2647, p2_p2_u2646, p2_p2_u2645, p2_p2_u2644, p2_p2_u2643, p2_p2_u2642, p2_p2_u2641, p2_p2_u2640, p2_p2_u2639, p2_p2_u3292, p2_p2_u2638, p2_p2_u3293, p2_p2_u3294, p2_p2_u2637, p2_p2_u3295, p2_p2_u2636, p2_p2_u3296, p2_p2_u2635, p2_p2_u3297, p2_p2_u2634, p2_p2_u2633, p2_p2_u3298, p2_p2_u3299, p2_p1_u3288, p2_p1_u3289, p2_p1_u3290, p2_p1_u3291, p2_p1_u3077, p2_p1_u3076, p2_p1_u3075, p2_p1_u3074, p2_p1_u3073, p2_p1_u3072, p2_p1_u3071, p2_p1_u3070, p2_p1_u3069, p2_p1_u3068, p2_p1_u3067, p2_p1_u3066, p2_p1_u3065, p2_p1_u3064, p2_p1_u3063, p2_p1_u3062, p2_p1_u3061, p2_p1_u3060, p2_p1_u3059, p2_p1_u3058, p2_p1_u3057, p2_p1_u3056, p2_p1_u3055, p2_p1_u3054, p2_p1_u3053, p2_p1_u3052, p2_p1_u3051, p2_p1_u3050, p2_p1_u3049, p2_p1_u3048, p2_p1_u3047, p2_p1_u3046, p2_p1_u3045, p2_p1_u3294, p2_p1_u3295, p2_p1_u3044, p2_p1_u3043, p2_p1_u3042, p2_p1_u3041, p2_p1_u3040, p2_p1_u3039, p2_p1_u3038, p2_p1_u3037, p2_p1_u3036, p2_p1_u3035, p2_p1_u3034, p2_p1_u3033, p2_p1_u3032, p2_p1_u3031, p2_p1_u3030, p2_p1_u3029, p2_p1_u3028, p2_p1_u3027, p2_p1_u3026, p2_p1_u3025, p2_p1_u3024, p2_p1_u3023, p2_p1_u3022, p2_p1_u3021, p2_p1_u3020, p2_p1_u3019, p2_p1_u3018, p2_p1_u3017, p2_p1_u3016, p2_p1_u3015, p2_p1_u3296, p2_p1_u3014, p2_p1_u3013, p2_p1_u3012, p2_p1_u3011, p2_p1_u3010, p2_p1_u3009, p2_p1_u3008, p2_p1_u3007, p2_p1_u3006, p2_p1_u3005, p2_p1_u3004, p2_p1_u3003, p2_p1_u3002, p2_p1_u3001, p2_p1_u3000, p2_p1_u2999, p2_p1_u2998, p2_p1_u2997, p2_p1_u2996, p2_p1_u2995, p2_p1_u2994, p2_p1_u2993, p2_p1_u2992, p2_p1_u2991, p2_p1_u2990, p2_p1_u2989, p2_p1_u2988, p2_p1_u2987, p2_p1_u2986, p2_p1_u2985, p2_p1_u2984, p2_p1_u2983, p2_p1_u2982, p2_p1_u2981, p2_p1_u2980, p2_p1_u2979, p2_p1_u2978, p2_p1_u2977, p2_p1_u2976, p2_p1_u2975, p2_p1_u2974, p2_p1_u2973, p2_p1_u2972, p2_p1_u2971, p2_p1_u2970, p2_p1_u2969, p2_p1_u2968, p2_p1_u2967, p2_p1_u2966, p2_p1_u2965, p2_p1_u2964, p2_p1_u2963, p2_p1_u2962, p2_p1_u2961, p2_p1_u2960, p2_p1_u2959, p2_p1_u2958, p2_p1_u2957, p2_p1_u2956, p2_p1_u2955, p2_p1_u2954, p2_p1_u2953, p2_p1_u2952, p2_p1_u2951, p2_p1_u2950, p2_p1_u2949, p2_p1_u2948, p2_p1_u2947, p2_p1_u2946, p2_p1_u2945, p2_p1_u2944, p2_p1_u2943, p2_p1_u2942, p2_p1_u2941, p2_p1_u2940, p2_p1_u2939, p2_p1_u2938, p2_p1_u2937, p2_p1_u2936, p2_p1_u2935, p2_p1_u2934, p2_p1_u2933, p2_p1_u2932, p2_p1_u2931, p2_p1_u2930, p2_p1_u2929, p2_p1_u2928, p2_p1_u2927, p2_p1_u2926, p2_p1_u2925, p2_p1_u2924, p2_p1_u2923, p2_p1_u2922, p2_p1_u2921, p2_p1_u2920, p2_p1_u2919, p2_p1_u2918, p2_p1_u2917, p2_p1_u2916, p2_p1_u2915, p2_p1_u2914, p2_p1_u2913, p2_p1_u2912, p2_p1_u2911, p2_p1_u2910, p2_p1_u2909, p2_p1_u2908, p2_p1_u2907, p2_p1_u2906, p2_p1_u2905, p2_p1_u2904, p2_p1_u2903, p2_p1_u2902, p2_p1_u2901, p2_p1_u2900, p2_p1_u2899, p2_p1_u2898, p2_p1_u2897, p2_p1_u2896, p2_p1_u2895, p2_p1_u2894, p2_p1_u2893, p2_p1_u2892, p2_p1_u2891, p2_p1_u2890, p2_p1_u2889, p2_p1_u2888, p2_p1_u2887, p2_p1_u2886, p2_p1_u2885, p2_p1_u2884, p2_p1_u3298, p2_p1_u3299, p2_p1_u3302, p2_p1_u3303, p2_p1_u3304, p2_p1_u2883, p2_p1_u2882, p2_p1_u2881, p2_p1_u2880, p2_p1_u2879, p2_p1_u2878, p2_p1_u2877, p2_p1_u2876, p2_p1_u2875, p2_p1_u2874, p2_p1_u2873, p2_p1_u2872, p2_p1_u2871, p2_p1_u2870, p2_p1_u2869, p2_p1_u2868, p2_p1_u2867, p2_p1_u2866, p2_p1_u2865, p2_p1_u2864, p2_p1_u2863, p2_p1_u2862, p2_p1_u2861, p2_p1_u2860, p2_p1_u2859, p2_p1_u2858, p2_p1_u2857, p2_p1_u2856, p2_p1_u2855, p2_p1_u2854, p2_p1_u2853, p2_p1_u2852, p2_p1_u2851, p2_p1_u2850, p2_p1_u2849, p2_p1_u2848, p2_p1_u2847, p2_p1_u2846, p2_p1_u2845, p2_p1_u2844, p2_p1_u2843, p2_p1_u2842, p2_p1_u2841, p2_p1_u2840, p2_p1_u2839, p2_p1_u2838, p2_p1_u2837, p2_p1_u2836, p2_p1_u2835, p2_p1_u2834, p2_p1_u2833, p2_p1_u2832, p2_p1_u2831, p2_p1_u2830, p2_p1_u2829, p2_p1_u2828, p2_p1_u2827, p2_p1_u2826, p2_p1_u2825, p2_p1_u2824, p2_p1_u2823, p2_p1_u2822, p2_p1_u2821, p2_p1_u2820, p2_p1_u2819, p2_p1_u2818, p2_p1_u2817, p2_p1_u2816, p2_p1_u2815, p2_p1_u2814, p2_p1_u2813, p2_p1_u2812, p2_p1_u2811, p2_p1_u2810, p2_p1_u2809, p2_p1_u2808, p2_p1_u2807, p2_p1_u2806, p2_p1_u2805, p2_p1_u2804, p2_p1_u2803, p2_p1_u2802, p2_p1_u2801, p2_p1_u2800, p2_p1_u2799, p2_p1_u2798, p2_p1_u2797, p2_p1_u2796, p2_p1_u2795, p2_p1_u2794, p2_p1_u2793, p2_p1_u2792, p2_p1_u2791, p2_p1_u2790, p2_p1_u2789, p2_p1_u2788, p2_p1_u2787, p2_p1_u2786, p2_p1_u2785, p2_p1_u2784, p2_p1_u2783, p2_p1_u2782, p2_p1_u2781, p2_p1_u2780, p2_p1_u2779, p2_p1_u2778, p2_p1_u2777, p2_p1_u2776, p2_p1_u2775, p2_p1_u2774, p2_p1_u2773, p2_p1_u2772, p2_p1_u2771, p2_p1_u2770, p2_p1_u2769, p2_p1_u2768, p2_p1_u2767, p2_p1_u2766, p2_p1_u2765, p2_p1_u2764, p2_p1_u2763, p2_p1_u2762, p2_p1_u2761, p2_p1_u2760, p2_p1_u2759, p2_p1_u2758, p2_p1_u2757, p2_p1_u2756, p2_p1_u2755, p2_p1_u2754, p2_p1_u2753, p2_p1_u2752, p2_p1_u2751, p2_p1_u2750, p2_p1_u2749, p2_p1_u2748, p2_p1_u2747, p2_p1_u2746, p2_p1_u2745, p2_p1_u2744, p2_p1_u2743, p2_p1_u2742, p2_p1_u2741, p2_p1_u2740, p2_p1_u2739, p2_p1_u2738, p2_p1_u2737, p2_p1_u2736, p2_p1_u2735, p2_p1_u2734, p2_p1_u2733, p2_p1_u2732, p2_p1_u2731, p2_p1_u2730, p2_p1_u2729, p2_p1_u2728, p2_p1_u2727, p2_p1_u2726, p2_p1_u2725, p2_p1_u2724, p2_p1_u2723, p2_p1_u2722, p2_p1_u2721, p2_p1_u2720, p2_p1_u2719, p2_p1_u2718, p2_p1_u2717, p2_p1_u2716, p2_p1_u2715, p2_p1_u2714, p2_p1_u2713, p2_p1_u2712, p2_p1_u2711, p2_p1_u2710, p2_p1_u2709, p2_p1_u2708, p2_p1_u2707, p2_p1_u2706, p2_p1_u2705, p2_p1_u2704, p2_p1_u2703, p2_p1_u2702, p2_p1_u2701, p2_p1_u2700, p2_p1_u2699, p2_p1_u2698, p2_p1_u2697, p2_p1_u2696, p2_p1_u2695, p2_p1_u2694, p2_p1_u2693, p2_p1_u2692, p2_p1_u2691, p2_p1_u2690, p2_p1_u2689, p2_p1_u2688, p2_p1_u2687, p2_p1_u2686, p2_p1_u2685, p2_p1_u2684, p2_p1_u2683, p2_p1_u2682, p2_p1_u2681, p2_p1_u2680, p2_p1_u2679, p2_p1_u2678, p2_p1_u2677, p2_p1_u2676, p2_p1_u2675, p2_p1_u2674, p2_p1_u2673, p2_p1_u2672, p2_p1_u2671, p2_p1_u2670, p2_p1_u2669, p2_p1_u2668, p2_p1_u2667, p2_p1_u2666, p2_p1_u2665, p2_p1_u2664, p2_p1_u2663, p2_p1_u2662, p2_p1_u2661, p2_p1_u2660, p2_p1_u2659, p2_p1_u2658, p2_p1_u2657, p2_p1_u2656, p2_p1_u2655, p2_p1_u3306, p2_p1_u2654, p2_p1_u3307, p2_p1_u3308, p2_p1_u2653, p2_p1_u3309, p2_p1_u2652, p2_p1_u3310, p2_p1_u2651, p2_p1_u3311, p2_p1_u2650, p2_p1_u2649, p2_p1_u3312, p2_p1_u3313;
initial begin
	$readmemb(`in_file, input_vec_mem );
end

always #(`cycle/2) clk = ~clk;

b18_ras cc (.HOLD(vec[3356]), .NA(vec[3355]), .BS(vec[3354]), .SEL(vec[3353]), .DIN_31_(vec[3352]), .DIN_30_(vec[3351]), .DIN_29_(vec[3350]), .DIN_28_(vec[3349]), .DIN_27_(vec[3348]), .DIN_26_(vec[3347]), .DIN_25_(vec[3346]), .DIN_24_(vec[3345]), .DIN_23_(vec[3344]), .DIN_22_(vec[3343]), .DIN_21_(vec[3342]), .DIN_20_(vec[3341]), .DIN_19_(vec[3340]), .DIN_18_(vec[3339]), .DIN_17_(vec[3338]), .DIN_16_(vec[3337]), .DIN_15_(vec[3336]), .DIN_14_(vec[3335]), .DIN_13_(vec[3334]), .DIN_12_(vec[3333]), .DIN_11_(vec[3332]), .DIN_10_(vec[3331]), .DIN_9_(vec[3330]), .DIN_8_(vec[3329]), .DIN_7_(vec[3328]), .DIN_6_(vec[3327]), .DIN_5_(vec[3326]), .DIN_4_(vec[3325]), .DIN_3_(vec[3324]), .DIN_2_(vec[3323]), .DIN_1_(vec[3322]), .DIN_0_(vec[3321]), .LOGIC0(vec[3320]), .P1_BUF1_REG_0_(vec[3319]), .P1_BUF1_REG_1_(vec[3318]), .P1_BUF1_REG_2_(vec[3317]), .P1_BUF1_REG_3_(vec[3316]), .P1_BUF1_REG_4_(vec[3315]), .P1_BUF1_REG_5_(vec[3314]), .P1_BUF1_REG_6_(vec[3313]), .P1_BUF1_REG_7_(vec[3312]), .P1_BUF1_REG_8_(vec[3311]), .P1_BUF1_REG_9_(vec[3310]), .P1_BUF1_REG_10_(vec[3309]), .P1_BUF1_REG_11_(vec[3308]), .P1_BUF1_REG_12_(vec[3307]), .P1_BUF1_REG_13_(vec[3306]), .P1_BUF1_REG_14_(vec[3305]), .P1_BUF1_REG_15_(vec[3304]), .P1_BUF1_REG_16_(vec[3303]), .P1_BUF1_REG_17_(vec[3302]), .P1_BUF1_REG_18_(vec[3301]), .P1_BUF1_REG_19_(vec[3300]), .P1_BUF1_REG_20_(vec[3299]), .P1_BUF1_REG_21_(vec[3298]), .P1_BUF1_REG_22_(vec[3297]), .P1_BUF1_REG_23_(vec[3296]), .P1_BUF1_REG_24_(vec[3295]), .P1_BUF1_REG_25_(vec[3294]), .P1_BUF1_REG_26_(vec[3293]), .P1_BUF1_REG_27_(vec[3292]), .P1_BUF1_REG_28_(vec[3291]), .P1_BUF1_REG_29_(vec[3290]), .P1_BUF1_REG_30_(vec[3289]), .P1_BUF1_REG_31_(vec[3288]), .P1_BUF2_REG_0_(vec[3287]), .P1_BUF2_REG_1_(vec[3286]), .P1_BUF2_REG_2_(vec[3285]), .P1_BUF2_REG_3_(vec[3284]), .P1_BUF2_REG_4_(vec[3283]), .P1_BUF2_REG_5_(vec[3282]), .P1_BUF2_REG_6_(vec[3281]), .P1_BUF2_REG_7_(vec[3280]), .P1_BUF2_REG_8_(vec[3279]), .P1_BUF2_REG_9_(vec[3278]), .P1_BUF2_REG_10_(vec[3277]), .P1_BUF2_REG_11_(vec[3276]), .P1_BUF2_REG_12_(vec[3275]), .P1_BUF2_REG_13_(vec[3274]), .P1_BUF2_REG_14_(vec[3273]), .P1_BUF2_REG_15_(vec[3272]), .P1_BUF2_REG_16_(vec[3271]), .P1_BUF2_REG_17_(vec[3270]), .P1_BUF2_REG_18_(vec[3269]), .P1_BUF2_REG_19_(vec[3268]), .P1_BUF2_REG_20_(vec[3267]), .P1_BUF2_REG_21_(vec[3266]), .P1_BUF2_REG_22_(vec[3265]), .P1_BUF2_REG_23_(vec[3264]), .P1_BUF2_REG_24_(vec[3263]), .P1_BUF2_REG_25_(vec[3262]), .P1_BUF2_REG_26_(vec[3261]), .P1_BUF2_REG_27_(vec[3260]), .P1_BUF2_REG_28_(vec[3259]), .P1_BUF2_REG_29_(vec[3258]), .P1_BUF2_REG_30_(vec[3257]), .P1_BUF2_REG_31_(vec[3256]), .P1_READY12_REG(vec[3255]), .P1_READY21_REG(vec[3254]), .P1_READY22_REG(vec[3253]), .P1_READY11_REG(vec[3252]), .P2_BUF1_REG_0_(vec[3251]), .P2_BUF1_REG_1_(vec[3250]), .P2_BUF1_REG_2_(vec[3249]), .P2_BUF1_REG_3_(vec[3248]), .P2_BUF1_REG_4_(vec[3247]), .P2_BUF1_REG_5_(vec[3246]), .P2_BUF1_REG_6_(vec[3245]), .P2_BUF1_REG_7_(vec[3244]), .P2_BUF1_REG_8_(vec[3243]), .P2_BUF1_REG_9_(vec[3242]), .P2_BUF1_REG_10_(vec[3241]), .P2_BUF1_REG_11_(vec[3240]), .P2_BUF1_REG_12_(vec[3239]), .P2_BUF1_REG_13_(vec[3238]), .P2_BUF1_REG_14_(vec[3237]), .P2_BUF1_REG_15_(vec[3236]), .P2_BUF1_REG_16_(vec[3235]), .P2_BUF1_REG_17_(vec[3234]), .P2_BUF1_REG_18_(vec[3233]), .P2_BUF1_REG_19_(vec[3232]), .P2_BUF1_REG_20_(vec[3231]), .P2_BUF1_REG_21_(vec[3230]), .P2_BUF1_REG_22_(vec[3229]), .P2_BUF1_REG_23_(vec[3228]), .P2_BUF1_REG_24_(vec[3227]), .P2_BUF1_REG_25_(vec[3226]), .P2_BUF1_REG_26_(vec[3225]), .P2_BUF1_REG_27_(vec[3224]), .P2_BUF1_REG_28_(vec[3223]), .P2_BUF1_REG_29_(vec[3222]), .P2_BUF1_REG_30_(vec[3221]), .P2_BUF1_REG_31_(vec[3220]), .P2_BUF2_REG_0_(vec[3219]), .P2_BUF2_REG_1_(vec[3218]), .P2_BUF2_REG_2_(vec[3217]), .P2_BUF2_REG_3_(vec[3216]), .P2_BUF2_REG_4_(vec[3215]), .P2_BUF2_REG_5_(vec[3214]), .P2_BUF2_REG_6_(vec[3213]), .P2_BUF2_REG_7_(vec[3212]), .P2_BUF2_REG_8_(vec[3211]), .P2_BUF2_REG_9_(vec[3210]), .P2_BUF2_REG_10_(vec[3209]), .P2_BUF2_REG_11_(vec[3208]), .P2_BUF2_REG_12_(vec[3207]), .P2_BUF2_REG_13_(vec[3206]), .P2_BUF2_REG_14_(vec[3205]), .P2_BUF2_REG_15_(vec[3204]), .P2_BUF2_REG_16_(vec[3203]), .P2_BUF2_REG_17_(vec[3202]), .P2_BUF2_REG_18_(vec[3201]), .P2_BUF2_REG_19_(vec[3200]), .P2_BUF2_REG_20_(vec[3199]), .P2_BUF2_REG_21_(vec[3198]), .P2_BUF2_REG_22_(vec[3197]), .P2_BUF2_REG_23_(vec[3196]), .P2_BUF2_REG_24_(vec[3195]), .P2_BUF2_REG_25_(vec[3194]), .P2_BUF2_REG_26_(vec[3193]), .P2_BUF2_REG_27_(vec[3192]), .P2_BUF2_REG_28_(vec[3191]), .P2_BUF2_REG_29_(vec[3190]), .P2_BUF2_REG_30_(vec[3189]), .P2_BUF2_REG_31_(vec[3188]), .P2_READY12_REG(vec[3187]), .P2_READY21_REG(vec[3186]), .P2_READY22_REG(vec[3185]), .P2_READY11_REG(vec[3184]), .P3_IR_REG_0_(vec[3183]), .P3_IR_REG_1_(vec[3182]), .P3_IR_REG_2_(vec[3181]), .P3_IR_REG_3_(vec[3180]), .P3_IR_REG_4_(vec[3179]), .P3_IR_REG_5_(vec[3178]), .P3_IR_REG_6_(vec[3177]), .P3_IR_REG_7_(vec[3176]), .P3_IR_REG_8_(vec[3175]), .P3_IR_REG_9_(vec[3174]), .P3_IR_REG_10_(vec[3173]), .P3_IR_REG_11_(vec[3172]), .P3_IR_REG_12_(vec[3171]), .P3_IR_REG_13_(vec[3170]), .P3_IR_REG_14_(vec[3169]), .P3_IR_REG_15_(vec[3168]), .P3_IR_REG_16_(vec[3167]), .P3_IR_REG_17_(vec[3166]), .P3_IR_REG_18_(vec[3165]), .P3_IR_REG_19_(vec[3164]), .P3_IR_REG_20_(vec[3163]), .P3_IR_REG_21_(vec[3162]), .P3_IR_REG_22_(vec[3161]), .P3_IR_REG_23_(vec[3160]), .P3_IR_REG_24_(vec[3159]), .P3_IR_REG_25_(vec[3158]), .P3_IR_REG_26_(vec[3157]), .P3_IR_REG_27_(vec[3156]), .P3_IR_REG_28_(vec[3155]), .P3_IR_REG_29_(vec[3154]), .P3_IR_REG_30_(vec[3153]), .P3_IR_REG_31_(vec[3152]), .P3_D_REG_0_(vec[3151]), .P3_D_REG_1_(vec[3150]), .P3_D_REG_2_(vec[3149]), .P3_D_REG_3_(vec[3148]), .P3_D_REG_4_(vec[3147]), .P3_D_REG_5_(vec[3146]), .P3_D_REG_6_(vec[3145]), .P3_D_REG_7_(vec[3144]), .P3_D_REG_8_(vec[3143]), .P3_D_REG_9_(vec[3142]), .P3_D_REG_10_(vec[3141]), .P3_D_REG_11_(vec[3140]), .P3_D_REG_12_(vec[3139]), .P3_D_REG_13_(vec[3138]), .P3_D_REG_14_(vec[3137]), .P3_D_REG_15_(vec[3136]), .P3_D_REG_16_(vec[3135]), .P3_D_REG_17_(vec[3134]), .P3_D_REG_18_(vec[3133]), .P3_D_REG_19_(vec[3132]), .P3_D_REG_20_(vec[3131]), .P3_D_REG_21_(vec[3130]), .P3_D_REG_22_(vec[3129]), .P3_D_REG_23_(vec[3128]), .P3_D_REG_24_(vec[3127]), .P3_D_REG_25_(vec[3126]), .P3_D_REG_26_(vec[3125]), .P3_D_REG_27_(vec[3124]), .P3_D_REG_28_(vec[3123]), .P3_D_REG_29_(vec[3122]), .P3_D_REG_30_(vec[3121]), .P3_D_REG_31_(vec[3120]), .P3_REG0_REG_0_(vec[3119]), .P3_REG0_REG_1_(vec[3118]), .P3_REG0_REG_2_(vec[3117]), .P3_REG0_REG_3_(vec[3116]), .P3_REG0_REG_4_(vec[3115]), .P3_REG0_REG_5_(vec[3114]), .P3_REG0_REG_6_(vec[3113]), .P3_REG0_REG_7_(vec[3112]), .P3_REG0_REG_8_(vec[3111]), .P3_REG0_REG_9_(vec[3110]), .P3_REG0_REG_10_(vec[3109]), .P3_REG0_REG_11_(vec[3108]), .P3_REG0_REG_12_(vec[3107]), .P3_REG0_REG_13_(vec[3106]), .P3_REG0_REG_14_(vec[3105]), .P3_REG0_REG_15_(vec[3104]), .P3_REG0_REG_16_(vec[3103]), .P3_REG0_REG_17_(vec[3102]), .P3_REG0_REG_18_(vec[3101]), .P3_REG0_REG_19_(vec[3100]), .P3_REG0_REG_20_(vec[3099]), .P3_REG0_REG_21_(vec[3098]), .P3_REG0_REG_22_(vec[3097]), .P3_REG0_REG_23_(vec[3096]), .P3_REG0_REG_24_(vec[3095]), .P3_REG0_REG_25_(vec[3094]), .P3_REG0_REG_26_(vec[3093]), .P3_REG0_REG_27_(vec[3092]), .P3_REG0_REG_28_(vec[3091]), .P3_REG0_REG_29_(vec[3090]), .P3_REG0_REG_30_(vec[3089]), .P3_REG0_REG_31_(vec[3088]), .P3_REG1_REG_0_(vec[3087]), .P3_REG1_REG_1_(vec[3086]), .P3_REG1_REG_2_(vec[3085]), .P3_REG1_REG_3_(vec[3084]), .P3_REG1_REG_4_(vec[3083]), .P3_REG1_REG_5_(vec[3082]), .P3_REG1_REG_6_(vec[3081]), .P3_REG1_REG_7_(vec[3080]), .P3_REG1_REG_8_(vec[3079]), .P3_REG1_REG_9_(vec[3078]), .P3_REG1_REG_10_(vec[3077]), .P3_REG1_REG_11_(vec[3076]), .P3_REG1_REG_12_(vec[3075]), .P3_REG1_REG_13_(vec[3074]), .P3_REG1_REG_14_(vec[3073]), .P3_REG1_REG_15_(vec[3072]), .P3_REG1_REG_16_(vec[3071]), .P3_REG1_REG_17_(vec[3070]), .P3_REG1_REG_18_(vec[3069]), .P3_REG1_REG_19_(vec[3068]), .P3_REG1_REG_20_(vec[3067]), .P3_REG1_REG_21_(vec[3066]), .P3_REG1_REG_22_(vec[3065]), .P3_REG1_REG_23_(vec[3064]), .P3_REG1_REG_24_(vec[3063]), .P3_REG1_REG_25_(vec[3062]), .P3_REG1_REG_26_(vec[3061]), .P3_REG1_REG_27_(vec[3060]), .P3_REG1_REG_28_(vec[3059]), .P3_REG1_REG_29_(vec[3058]), .P3_REG1_REG_30_(vec[3057]), .P3_REG1_REG_31_(vec[3056]), .P3_REG2_REG_0_(vec[3055]), .P3_REG2_REG_1_(vec[3054]), .P3_REG2_REG_2_(vec[3053]), .P3_REG2_REG_3_(vec[3052]), .P3_REG2_REG_4_(vec[3051]), .P3_REG2_REG_5_(vec[3050]), .P3_REG2_REG_6_(vec[3049]), .P3_REG2_REG_7_(vec[3048]), .P3_REG2_REG_8_(vec[3047]), .P3_REG2_REG_9_(vec[3046]), .P3_REG2_REG_10_(vec[3045]), .P3_REG2_REG_11_(vec[3044]), .P3_REG2_REG_12_(vec[3043]), .P3_REG2_REG_13_(vec[3042]), .P3_REG2_REG_14_(vec[3041]), .P3_REG2_REG_15_(vec[3040]), .P3_REG2_REG_16_(vec[3039]), .P3_REG2_REG_17_(vec[3038]), .P3_REG2_REG_18_(vec[3037]), .P3_REG2_REG_19_(vec[3036]), .P3_REG2_REG_20_(vec[3035]), .P3_REG2_REG_21_(vec[3034]), .P3_REG2_REG_22_(vec[3033]), .P3_REG2_REG_23_(vec[3032]), .P3_REG2_REG_24_(vec[3031]), .P3_REG2_REG_25_(vec[3030]), .P3_REG2_REG_26_(vec[3029]), .P3_REG2_REG_27_(vec[3028]), .P3_REG2_REG_28_(vec[3027]), .P3_REG2_REG_29_(vec[3026]), .P3_REG2_REG_30_(vec[3025]), .P3_REG2_REG_31_(vec[3024]), .P3_ADDR_REG_19_(vec[3023]), .P3_ADDR_REG_18_(vec[3022]), .P3_ADDR_REG_17_(vec[3021]), .P3_ADDR_REG_16_(vec[3020]), .P3_ADDR_REG_15_(vec[3019]), .P3_ADDR_REG_14_(vec[3018]), .P3_ADDR_REG_13_(vec[3017]), .P3_ADDR_REG_12_(vec[3016]), .P3_ADDR_REG_11_(vec[3015]), .P3_ADDR_REG_10_(vec[3014]), .P3_ADDR_REG_9_(vec[3013]), .P3_ADDR_REG_8_(vec[3012]), .P3_ADDR_REG_7_(vec[3011]), .P3_ADDR_REG_6_(vec[3010]), .P3_ADDR_REG_5_(vec[3009]), .P3_ADDR_REG_4_(vec[3008]), .P3_ADDR_REG_3_(vec[3007]), .P3_ADDR_REG_2_(vec[3006]), .P3_ADDR_REG_1_(vec[3005]), .P3_ADDR_REG_0_(vec[3004]), .P3_DATAO_REG_0_(vec[3003]), .P3_DATAO_REG_1_(vec[3002]), .P3_DATAO_REG_2_(vec[3001]), .P3_DATAO_REG_3_(vec[3000]), .P3_DATAO_REG_4_(vec[2999]), .P3_DATAO_REG_5_(vec[2998]), .P3_DATAO_REG_6_(vec[2997]), .P3_DATAO_REG_7_(vec[2996]), .P3_DATAO_REG_8_(vec[2995]), .P3_DATAO_REG_9_(vec[2994]), .P3_DATAO_REG_10_(vec[2993]), .P3_DATAO_REG_11_(vec[2992]), .P3_DATAO_REG_12_(vec[2991]), .P3_DATAO_REG_13_(vec[2990]), .P3_DATAO_REG_14_(vec[2989]), .P3_DATAO_REG_15_(vec[2988]), .P3_DATAO_REG_16_(vec[2987]), .P3_DATAO_REG_17_(vec[2986]), .P3_DATAO_REG_18_(vec[2985]), .P3_DATAO_REG_19_(vec[2984]), .P3_DATAO_REG_20_(vec[2983]), .P3_DATAO_REG_21_(vec[2982]), .P3_DATAO_REG_22_(vec[2981]), .P3_DATAO_REG_23_(vec[2980]), .P3_DATAO_REG_24_(vec[2979]), .P3_DATAO_REG_25_(vec[2978]), .P3_DATAO_REG_26_(vec[2977]), .P3_DATAO_REG_27_(vec[2976]), .P3_DATAO_REG_28_(vec[2975]), .P3_DATAO_REG_29_(vec[2974]), .P3_DATAO_REG_30_(vec[2973]), .P3_DATAO_REG_31_(vec[2972]), .P3_B_REG(vec[2971]), .P3_REG3_REG_15_(vec[2970]), .P3_REG3_REG_26_(vec[2969]), .P3_REG3_REG_6_(vec[2968]), .P3_REG3_REG_18_(vec[2967]), .P3_REG3_REG_2_(vec[2966]), .P3_REG3_REG_11_(vec[2965]), .P3_REG3_REG_22_(vec[2964]), .P3_REG3_REG_13_(vec[2963]), .P3_REG3_REG_20_(vec[2962]), .P3_REG3_REG_0_(vec[2961]), .P3_REG3_REG_9_(vec[2960]), .P3_REG3_REG_4_(vec[2959]), .P3_REG3_REG_24_(vec[2958]), .P3_REG3_REG_17_(vec[2957]), .P3_REG3_REG_5_(vec[2956]), .P3_REG3_REG_16_(vec[2955]), .P3_REG3_REG_25_(vec[2954]), .P3_REG3_REG_12_(vec[2953]), .P3_REG3_REG_21_(vec[2952]), .P3_REG3_REG_1_(vec[2951]), .P3_REG3_REG_8_(vec[2950]), .P3_REG3_REG_28_(vec[2949]), .P3_REG3_REG_19_(vec[2948]), .P3_REG3_REG_3_(vec[2947]), .P3_REG3_REG_10_(vec[2946]), .P3_REG3_REG_23_(vec[2945]), .P3_REG3_REG_14_(vec[2944]), .P3_REG3_REG_27_(vec[2943]), .P3_REG3_REG_7_(vec[2942]), .P3_STATE_REG(vec[2941]), .P3_RD_REG(vec[2940]), .P3_WR_REG(vec[2939]), .P4_IR_REG_0_(vec[2938]), .P4_IR_REG_1_(vec[2937]), .P4_IR_REG_2_(vec[2936]), .P4_IR_REG_3_(vec[2935]), .P4_IR_REG_4_(vec[2934]), .P4_IR_REG_5_(vec[2933]), .P4_IR_REG_6_(vec[2932]), .P4_IR_REG_7_(vec[2931]), .P4_IR_REG_8_(vec[2930]), .P4_IR_REG_9_(vec[2929]), .P4_IR_REG_10_(vec[2928]), .P4_IR_REG_11_(vec[2927]), .P4_IR_REG_12_(vec[2926]), .P4_IR_REG_13_(vec[2925]), .P4_IR_REG_14_(vec[2924]), .P4_IR_REG_15_(vec[2923]), .P4_IR_REG_16_(vec[2922]), .P4_IR_REG_17_(vec[2921]), .P4_IR_REG_18_(vec[2920]), .P4_IR_REG_19_(vec[2919]), .P4_IR_REG_20_(vec[2918]), .P4_IR_REG_21_(vec[2917]), .P4_IR_REG_22_(vec[2916]), .P4_IR_REG_23_(vec[2915]), .P4_IR_REG_24_(vec[2914]), .P4_IR_REG_25_(vec[2913]), .P4_IR_REG_26_(vec[2912]), .P4_IR_REG_27_(vec[2911]), .P4_IR_REG_28_(vec[2910]), .P4_IR_REG_29_(vec[2909]), .P4_IR_REG_30_(vec[2908]), .P4_IR_REG_31_(vec[2907]), .P4_D_REG_0_(vec[2906]), .P4_D_REG_1_(vec[2905]), .P4_D_REG_2_(vec[2904]), .P4_D_REG_3_(vec[2903]), .P4_D_REG_4_(vec[2902]), .P4_D_REG_5_(vec[2901]), .P4_D_REG_6_(vec[2900]), .P4_D_REG_7_(vec[2899]), .P4_D_REG_8_(vec[2898]), .P4_D_REG_9_(vec[2897]), .P4_D_REG_10_(vec[2896]), .P4_D_REG_11_(vec[2895]), .P4_D_REG_12_(vec[2894]), .P4_D_REG_13_(vec[2893]), .P4_D_REG_14_(vec[2892]), .P4_D_REG_15_(vec[2891]), .P4_D_REG_16_(vec[2890]), .P4_D_REG_17_(vec[2889]), .P4_D_REG_18_(vec[2888]), .P4_D_REG_19_(vec[2887]), .P4_D_REG_20_(vec[2886]), .P4_D_REG_21_(vec[2885]), .P4_D_REG_22_(vec[2884]), .P4_D_REG_23_(vec[2883]), .P4_D_REG_24_(vec[2882]), .P4_D_REG_25_(vec[2881]), .P4_D_REG_26_(vec[2880]), .P4_D_REG_27_(vec[2879]), .P4_D_REG_28_(vec[2878]), .P4_D_REG_29_(vec[2877]), .P4_D_REG_30_(vec[2876]), .P4_D_REG_31_(vec[2875]), .P4_REG0_REG_0_(vec[2874]), .P4_REG0_REG_1_(vec[2873]), .P4_REG0_REG_2_(vec[2872]), .P4_REG0_REG_3_(vec[2871]), .P4_REG0_REG_4_(vec[2870]), .P4_REG0_REG_5_(vec[2869]), .P4_REG0_REG_6_(vec[2868]), .P4_REG0_REG_7_(vec[2867]), .P4_REG0_REG_8_(vec[2866]), .P4_REG0_REG_9_(vec[2865]), .P4_REG0_REG_10_(vec[2864]), .P4_REG0_REG_11_(vec[2863]), .P4_REG0_REG_12_(vec[2862]), .P4_REG0_REG_13_(vec[2861]), .P4_REG0_REG_14_(vec[2860]), .P4_REG0_REG_15_(vec[2859]), .P4_REG0_REG_16_(vec[2858]), .P4_REG0_REG_17_(vec[2857]), .P4_REG0_REG_18_(vec[2856]), .P4_REG0_REG_19_(vec[2855]), .P4_REG0_REG_20_(vec[2854]), .P4_REG0_REG_21_(vec[2853]), .P4_REG0_REG_22_(vec[2852]), .P4_REG0_REG_23_(vec[2851]), .P4_REG0_REG_24_(vec[2850]), .P4_REG0_REG_25_(vec[2849]), .P4_REG0_REG_26_(vec[2848]), .P4_REG0_REG_27_(vec[2847]), .P4_REG0_REG_28_(vec[2846]), .P4_REG0_REG_29_(vec[2845]), .P4_REG0_REG_30_(vec[2844]), .P4_REG0_REG_31_(vec[2843]), .P4_REG1_REG_0_(vec[2842]), .P4_REG1_REG_1_(vec[2841]), .P4_REG1_REG_2_(vec[2840]), .P4_REG1_REG_3_(vec[2839]), .P4_REG1_REG_4_(vec[2838]), .P4_REG1_REG_5_(vec[2837]), .P4_REG1_REG_6_(vec[2836]), .P4_REG1_REG_7_(vec[2835]), .P4_REG1_REG_8_(vec[2834]), .P4_REG1_REG_9_(vec[2833]), .P4_REG1_REG_10_(vec[2832]), .P4_REG1_REG_11_(vec[2831]), .P4_REG1_REG_12_(vec[2830]), .P4_REG1_REG_13_(vec[2829]), .P4_REG1_REG_14_(vec[2828]), .P4_REG1_REG_15_(vec[2827]), .P4_REG1_REG_16_(vec[2826]), .P4_REG1_REG_17_(vec[2825]), .P4_REG1_REG_18_(vec[2824]), .P4_REG1_REG_19_(vec[2823]), .P4_REG1_REG_20_(vec[2822]), .P4_REG1_REG_21_(vec[2821]), .P4_REG1_REG_22_(vec[2820]), .P4_REG1_REG_23_(vec[2819]), .P4_REG1_REG_24_(vec[2818]), .P4_REG1_REG_25_(vec[2817]), .P4_REG1_REG_26_(vec[2816]), .P4_REG1_REG_27_(vec[2815]), .P4_REG1_REG_28_(vec[2814]), .P4_REG1_REG_29_(vec[2813]), .P4_REG1_REG_30_(vec[2812]), .P4_REG1_REG_31_(vec[2811]), .P4_REG2_REG_0_(vec[2810]), .P4_REG2_REG_1_(vec[2809]), .P4_REG2_REG_2_(vec[2808]), .P4_REG2_REG_3_(vec[2807]), .P4_REG2_REG_4_(vec[2806]), .P4_REG2_REG_5_(vec[2805]), .P4_REG2_REG_6_(vec[2804]), .P4_REG2_REG_7_(vec[2803]), .P4_REG2_REG_8_(vec[2802]), .P4_REG2_REG_9_(vec[2801]), .P4_REG2_REG_10_(vec[2800]), .P4_REG2_REG_11_(vec[2799]), .P4_REG2_REG_12_(vec[2798]), .P4_REG2_REG_13_(vec[2797]), .P4_REG2_REG_14_(vec[2796]), .P4_REG2_REG_15_(vec[2795]), .P4_REG2_REG_16_(vec[2794]), .P4_REG2_REG_17_(vec[2793]), .P4_REG2_REG_18_(vec[2792]), .P4_REG2_REG_19_(vec[2791]), .P4_REG2_REG_20_(vec[2790]), .P4_REG2_REG_21_(vec[2789]), .P4_REG2_REG_22_(vec[2788]), .P4_REG2_REG_23_(vec[2787]), .P4_REG2_REG_24_(vec[2786]), .P4_REG2_REG_25_(vec[2785]), .P4_REG2_REG_26_(vec[2784]), .P4_REG2_REG_27_(vec[2783]), .P4_REG2_REG_28_(vec[2782]), .P4_REG2_REG_29_(vec[2781]), .P4_REG2_REG_30_(vec[2780]), .P4_REG2_REG_31_(vec[2779]), .P4_ADDR_REG_19_(vec[2778]), .P4_ADDR_REG_18_(vec[2777]), .P4_ADDR_REG_17_(vec[2776]), .P4_ADDR_REG_16_(vec[2775]), .P4_ADDR_REG_15_(vec[2774]), .P4_ADDR_REG_14_(vec[2773]), .P4_ADDR_REG_13_(vec[2772]), .P4_ADDR_REG_12_(vec[2771]), .P4_ADDR_REG_11_(vec[2770]), .P4_ADDR_REG_10_(vec[2769]), .P4_ADDR_REG_9_(vec[2768]), .P4_ADDR_REG_8_(vec[2767]), .P4_ADDR_REG_7_(vec[2766]), .P4_ADDR_REG_6_(vec[2765]), .P4_ADDR_REG_5_(vec[2764]), .P4_ADDR_REG_4_(vec[2763]), .P4_ADDR_REG_3_(vec[2762]), .P4_ADDR_REG_2_(vec[2761]), .P4_ADDR_REG_1_(vec[2760]), .P4_ADDR_REG_0_(vec[2759]), .P4_DATAO_REG_0_(vec[2758]), .P4_DATAO_REG_1_(vec[2757]), .P4_DATAO_REG_2_(vec[2756]), .P4_DATAO_REG_3_(vec[2755]), .P4_DATAO_REG_4_(vec[2754]), .P4_DATAO_REG_5_(vec[2753]), .P4_DATAO_REG_6_(vec[2752]), .P4_DATAO_REG_7_(vec[2751]), .P4_DATAO_REG_8_(vec[2750]), .P4_DATAO_REG_9_(vec[2749]), .P4_DATAO_REG_10_(vec[2748]), .P4_DATAO_REG_11_(vec[2747]), .P4_DATAO_REG_12_(vec[2746]), .P4_DATAO_REG_13_(vec[2745]), .P4_DATAO_REG_14_(vec[2744]), .P4_DATAO_REG_15_(vec[2743]), .P4_DATAO_REG_16_(vec[2742]), .P4_DATAO_REG_17_(vec[2741]), .P4_DATAO_REG_18_(vec[2740]), .P4_DATAO_REG_19_(vec[2739]), .P4_DATAO_REG_20_(vec[2738]), .P4_DATAO_REG_21_(vec[2737]), .P4_DATAO_REG_22_(vec[2736]), .P4_DATAO_REG_23_(vec[2735]), .P4_DATAO_REG_24_(vec[2734]), .P4_DATAO_REG_25_(vec[2733]), .P4_DATAO_REG_26_(vec[2732]), .P4_DATAO_REG_27_(vec[2731]), .P4_DATAO_REG_28_(vec[2730]), .P4_DATAO_REG_29_(vec[2729]), .P4_DATAO_REG_30_(vec[2728]), .P4_DATAO_REG_31_(vec[2727]), .P4_B_REG(vec[2726]), .P4_REG3_REG_15_(vec[2725]), .P4_REG3_REG_26_(vec[2724]), .P4_REG3_REG_6_(vec[2723]), .P4_REG3_REG_18_(vec[2722]), .P4_REG3_REG_2_(vec[2721]), .P4_REG3_REG_11_(vec[2720]), .P4_REG3_REG_22_(vec[2719]), .P4_REG3_REG_13_(vec[2718]), .P4_REG3_REG_20_(vec[2717]), .P4_REG3_REG_0_(vec[2716]), .P4_REG3_REG_9_(vec[2715]), .P4_REG3_REG_4_(vec[2714]), .P4_REG3_REG_24_(vec[2713]), .P4_REG3_REG_17_(vec[2712]), .P4_REG3_REG_5_(vec[2711]), .P4_REG3_REG_16_(vec[2710]), .P4_REG3_REG_25_(vec[2709]), .P4_REG3_REG_12_(vec[2708]), .P4_REG3_REG_21_(vec[2707]), .P4_REG3_REG_1_(vec[2706]), .P4_REG3_REG_8_(vec[2705]), .P4_REG3_REG_28_(vec[2704]), .P4_REG3_REG_19_(vec[2703]), .P4_REG3_REG_3_(vec[2702]), .P4_REG3_REG_10_(vec[2701]), .P4_REG3_REG_23_(vec[2700]), .P4_REG3_REG_14_(vec[2699]), .P4_REG3_REG_27_(vec[2698]), .P4_REG3_REG_7_(vec[2697]), .P4_STATE_REG(vec[2696]), .P4_RD_REG(vec[2695]), .P4_WR_REG(vec[2694]), .P1_P3_BE_N_REG_3_(vec[2693]), .P1_P3_BE_N_REG_2_(vec[2692]), .P1_P3_BE_N_REG_1_(vec[2691]), .P1_P3_BE_N_REG_0_(vec[2690]), .P1_P3_ADDRESS_REG_29_(vec[2689]), .P1_P3_ADDRESS_REG_28_(vec[2688]), .P1_P3_ADDRESS_REG_27_(vec[2687]), .P1_P3_ADDRESS_REG_26_(vec[2686]), .P1_P3_ADDRESS_REG_25_(vec[2685]), .P1_P3_ADDRESS_REG_24_(vec[2684]), .P1_P3_ADDRESS_REG_23_(vec[2683]), .P1_P3_ADDRESS_REG_22_(vec[2682]), .P1_P3_ADDRESS_REG_21_(vec[2681]), .P1_P3_ADDRESS_REG_20_(vec[2680]), .P1_P3_ADDRESS_REG_19_(vec[2679]), .P1_P3_ADDRESS_REG_18_(vec[2678]), .P1_P3_ADDRESS_REG_17_(vec[2677]), .P1_P3_ADDRESS_REG_16_(vec[2676]), .P1_P3_ADDRESS_REG_15_(vec[2675]), .P1_P3_ADDRESS_REG_14_(vec[2674]), .P1_P3_ADDRESS_REG_13_(vec[2673]), .P1_P3_ADDRESS_REG_12_(vec[2672]), .P1_P3_ADDRESS_REG_11_(vec[2671]), .P1_P3_ADDRESS_REG_10_(vec[2670]), .P1_P3_ADDRESS_REG_9_(vec[2669]), .P1_P3_ADDRESS_REG_8_(vec[2668]), .P1_P3_ADDRESS_REG_7_(vec[2667]), .P1_P3_ADDRESS_REG_6_(vec[2666]), .P1_P3_ADDRESS_REG_5_(vec[2665]), .P1_P3_ADDRESS_REG_4_(vec[2664]), .P1_P3_ADDRESS_REG_3_(vec[2663]), .P1_P3_ADDRESS_REG_2_(vec[2662]), .P1_P3_ADDRESS_REG_1_(vec[2661]), .P1_P3_ADDRESS_REG_0_(vec[2660]), .P1_P3_STATE_REG_2_(vec[2659]), .P1_P3_STATE_REG_1_(vec[2658]), .P1_P3_STATE_REG_0_(vec[2657]), .P1_P3_DATAWIDTH_REG_0_(vec[2656]), .P1_P3_DATAWIDTH_REG_1_(vec[2655]), .P1_P3_DATAWIDTH_REG_2_(vec[2654]), .P1_P3_DATAWIDTH_REG_3_(vec[2653]), .P1_P3_DATAWIDTH_REG_4_(vec[2652]), .P1_P3_DATAWIDTH_REG_5_(vec[2651]), .P1_P3_DATAWIDTH_REG_6_(vec[2650]), .P1_P3_DATAWIDTH_REG_7_(vec[2649]), .P1_P3_DATAWIDTH_REG_8_(vec[2648]), .P1_P3_DATAWIDTH_REG_9_(vec[2647]), .P1_P3_DATAWIDTH_REG_10_(vec[2646]), .P1_P3_DATAWIDTH_REG_11_(vec[2645]), .P1_P3_DATAWIDTH_REG_12_(vec[2644]), .P1_P3_DATAWIDTH_REG_13_(vec[2643]), .P1_P3_DATAWIDTH_REG_14_(vec[2642]), .P1_P3_DATAWIDTH_REG_15_(vec[2641]), .P1_P3_DATAWIDTH_REG_16_(vec[2640]), .P1_P3_DATAWIDTH_REG_17_(vec[2639]), .P1_P3_DATAWIDTH_REG_18_(vec[2638]), .P1_P3_DATAWIDTH_REG_19_(vec[2637]), .P1_P3_DATAWIDTH_REG_20_(vec[2636]), .P1_P3_DATAWIDTH_REG_21_(vec[2635]), .P1_P3_DATAWIDTH_REG_22_(vec[2634]), .P1_P3_DATAWIDTH_REG_23_(vec[2633]), .P1_P3_DATAWIDTH_REG_24_(vec[2632]), .P1_P3_DATAWIDTH_REG_25_(vec[2631]), .P1_P3_DATAWIDTH_REG_26_(vec[2630]), .P1_P3_DATAWIDTH_REG_27_(vec[2629]), .P1_P3_DATAWIDTH_REG_28_(vec[2628]), .P1_P3_DATAWIDTH_REG_29_(vec[2627]), .P1_P3_DATAWIDTH_REG_30_(vec[2626]), .P1_P3_DATAWIDTH_REG_31_(vec[2625]), .P1_P3_STATE2_REG_3_(vec[2624]), .P1_P3_STATE2_REG_2_(vec[2623]), .P1_P3_STATE2_REG_1_(vec[2622]), .P1_P3_STATE2_REG_0_(vec[2621]), .P1_P3_INSTQUEUE_REG_15__7_(vec[2620]), .P1_P3_INSTQUEUE_REG_15__6_(vec[2619]), .P1_P3_INSTQUEUE_REG_15__5_(vec[2618]), .P1_P3_INSTQUEUE_REG_15__4_(vec[2617]), .P1_P3_INSTQUEUE_REG_15__3_(vec[2616]), .P1_P3_INSTQUEUE_REG_15__2_(vec[2615]), .P1_P3_INSTQUEUE_REG_15__1_(vec[2614]), .P1_P3_INSTQUEUE_REG_15__0_(vec[2613]), .P1_P3_INSTQUEUE_REG_14__7_(vec[2612]), .P1_P3_INSTQUEUE_REG_14__6_(vec[2611]), .P1_P3_INSTQUEUE_REG_14__5_(vec[2610]), .P1_P3_INSTQUEUE_REG_14__4_(vec[2609]), .P1_P3_INSTQUEUE_REG_14__3_(vec[2608]), .P1_P3_INSTQUEUE_REG_14__2_(vec[2607]), .P1_P3_INSTQUEUE_REG_14__1_(vec[2606]), .P1_P3_INSTQUEUE_REG_14__0_(vec[2605]), .P1_P3_INSTQUEUE_REG_13__7_(vec[2604]), .P1_P3_INSTQUEUE_REG_13__6_(vec[2603]), .P1_P3_INSTQUEUE_REG_13__5_(vec[2602]), .P1_P3_INSTQUEUE_REG_13__4_(vec[2601]), .P1_P3_INSTQUEUE_REG_13__3_(vec[2600]), .P1_P3_INSTQUEUE_REG_13__2_(vec[2599]), .P1_P3_INSTQUEUE_REG_13__1_(vec[2598]), .P1_P3_INSTQUEUE_REG_13__0_(vec[2597]), .P1_P3_INSTQUEUE_REG_12__7_(vec[2596]), .P1_P3_INSTQUEUE_REG_12__6_(vec[2595]), .P1_P3_INSTQUEUE_REG_12__5_(vec[2594]), .P1_P3_INSTQUEUE_REG_12__4_(vec[2593]), .P1_P3_INSTQUEUE_REG_12__3_(vec[2592]), .P1_P3_INSTQUEUE_REG_12__2_(vec[2591]), .P1_P3_INSTQUEUE_REG_12__1_(vec[2590]), .P1_P3_INSTQUEUE_REG_12__0_(vec[2589]), .P1_P3_INSTQUEUE_REG_11__7_(vec[2588]), .P1_P3_INSTQUEUE_REG_11__6_(vec[2587]), .P1_P3_INSTQUEUE_REG_11__5_(vec[2586]), .P1_P3_INSTQUEUE_REG_11__4_(vec[2585]), .P1_P3_INSTQUEUE_REG_11__3_(vec[2584]), .P1_P3_INSTQUEUE_REG_11__2_(vec[2583]), .P1_P3_INSTQUEUE_REG_11__1_(vec[2582]), .P1_P3_INSTQUEUE_REG_11__0_(vec[2581]), .P1_P3_INSTQUEUE_REG_10__7_(vec[2580]), .P1_P3_INSTQUEUE_REG_10__6_(vec[2579]), .P1_P3_INSTQUEUE_REG_10__5_(vec[2578]), .P1_P3_INSTQUEUE_REG_10__4_(vec[2577]), .P1_P3_INSTQUEUE_REG_10__3_(vec[2576]), .P1_P3_INSTQUEUE_REG_10__2_(vec[2575]), .P1_P3_INSTQUEUE_REG_10__1_(vec[2574]), .P1_P3_INSTQUEUE_REG_10__0_(vec[2573]), .P1_P3_INSTQUEUE_REG_9__7_(vec[2572]), .P1_P3_INSTQUEUE_REG_9__6_(vec[2571]), .P1_P3_INSTQUEUE_REG_9__5_(vec[2570]), .P1_P3_INSTQUEUE_REG_9__4_(vec[2569]), .P1_P3_INSTQUEUE_REG_9__3_(vec[2568]), .P1_P3_INSTQUEUE_REG_9__2_(vec[2567]), .P1_P3_INSTQUEUE_REG_9__1_(vec[2566]), .P1_P3_INSTQUEUE_REG_9__0_(vec[2565]), .P1_P3_INSTQUEUE_REG_8__7_(vec[2564]), .P1_P3_INSTQUEUE_REG_8__6_(vec[2563]), .P1_P3_INSTQUEUE_REG_8__5_(vec[2562]), .P1_P3_INSTQUEUE_REG_8__4_(vec[2561]), .P1_P3_INSTQUEUE_REG_8__3_(vec[2560]), .P1_P3_INSTQUEUE_REG_8__2_(vec[2559]), .P1_P3_INSTQUEUE_REG_8__1_(vec[2558]), .P1_P3_INSTQUEUE_REG_8__0_(vec[2557]), .P1_P3_INSTQUEUE_REG_7__7_(vec[2556]), .P1_P3_INSTQUEUE_REG_7__6_(vec[2555]), .P1_P3_INSTQUEUE_REG_7__5_(vec[2554]), .P1_P3_INSTQUEUE_REG_7__4_(vec[2553]), .P1_P3_INSTQUEUE_REG_7__3_(vec[2552]), .P1_P3_INSTQUEUE_REG_7__2_(vec[2551]), .P1_P3_INSTQUEUE_REG_7__1_(vec[2550]), .P1_P3_INSTQUEUE_REG_7__0_(vec[2549]), .P1_P3_INSTQUEUE_REG_6__7_(vec[2548]), .P1_P3_INSTQUEUE_REG_6__6_(vec[2547]), .P1_P3_INSTQUEUE_REG_6__5_(vec[2546]), .P1_P3_INSTQUEUE_REG_6__4_(vec[2545]), .P1_P3_INSTQUEUE_REG_6__3_(vec[2544]), .P1_P3_INSTQUEUE_REG_6__2_(vec[2543]), .P1_P3_INSTQUEUE_REG_6__1_(vec[2542]), .P1_P3_INSTQUEUE_REG_6__0_(vec[2541]), .P1_P3_INSTQUEUE_REG_5__7_(vec[2540]), .P1_P3_INSTQUEUE_REG_5__6_(vec[2539]), .P1_P3_INSTQUEUE_REG_5__5_(vec[2538]), .P1_P3_INSTQUEUE_REG_5__4_(vec[2537]), .P1_P3_INSTQUEUE_REG_5__3_(vec[2536]), .P1_P3_INSTQUEUE_REG_5__2_(vec[2535]), .P1_P3_INSTQUEUE_REG_5__1_(vec[2534]), .P1_P3_INSTQUEUE_REG_5__0_(vec[2533]), .P1_P3_INSTQUEUE_REG_4__7_(vec[2532]), .P1_P3_INSTQUEUE_REG_4__6_(vec[2531]), .P1_P3_INSTQUEUE_REG_4__5_(vec[2530]), .P1_P3_INSTQUEUE_REG_4__4_(vec[2529]), .P1_P3_INSTQUEUE_REG_4__3_(vec[2528]), .P1_P3_INSTQUEUE_REG_4__2_(vec[2527]), .P1_P3_INSTQUEUE_REG_4__1_(vec[2526]), .P1_P3_INSTQUEUE_REG_4__0_(vec[2525]), .P1_P3_INSTQUEUE_REG_3__7_(vec[2524]), .P1_P3_INSTQUEUE_REG_3__6_(vec[2523]), .P1_P3_INSTQUEUE_REG_3__5_(vec[2522]), .P1_P3_INSTQUEUE_REG_3__4_(vec[2521]), .P1_P3_INSTQUEUE_REG_3__3_(vec[2520]), .P1_P3_INSTQUEUE_REG_3__2_(vec[2519]), .P1_P3_INSTQUEUE_REG_3__1_(vec[2518]), .P1_P3_INSTQUEUE_REG_3__0_(vec[2517]), .P1_P3_INSTQUEUE_REG_2__7_(vec[2516]), .P1_P3_INSTQUEUE_REG_2__6_(vec[2515]), .P1_P3_INSTQUEUE_REG_2__5_(vec[2514]), .P1_P3_INSTQUEUE_REG_2__4_(vec[2513]), .P1_P3_INSTQUEUE_REG_2__3_(vec[2512]), .P1_P3_INSTQUEUE_REG_2__2_(vec[2511]), .P1_P3_INSTQUEUE_REG_2__1_(vec[2510]), .P1_P3_INSTQUEUE_REG_2__0_(vec[2509]), .P1_P3_INSTQUEUE_REG_1__7_(vec[2508]), .P1_P3_INSTQUEUE_REG_1__6_(vec[2507]), .P1_P3_INSTQUEUE_REG_1__5_(vec[2506]), .P1_P3_INSTQUEUE_REG_1__4_(vec[2505]), .P1_P3_INSTQUEUE_REG_1__3_(vec[2504]), .P1_P3_INSTQUEUE_REG_1__2_(vec[2503]), .P1_P3_INSTQUEUE_REG_1__1_(vec[2502]), .P1_P3_INSTQUEUE_REG_1__0_(vec[2501]), .P1_P3_INSTQUEUE_REG_0__7_(vec[2500]), .P1_P3_INSTQUEUE_REG_0__6_(vec[2499]), .P1_P3_INSTQUEUE_REG_0__5_(vec[2498]), .P1_P3_INSTQUEUE_REG_0__4_(vec[2497]), .P1_P3_INSTQUEUE_REG_0__3_(vec[2496]), .P1_P3_INSTQUEUE_REG_0__2_(vec[2495]), .P1_P3_INSTQUEUE_REG_0__1_(vec[2494]), .P1_P3_INSTQUEUE_REG_0__0_(vec[2493]), .P1_P3_INSTQUEUERD_ADDR_REG_4_(vec[2492]), .P1_P3_INSTQUEUERD_ADDR_REG_3_(vec[2491]), .P1_P3_INSTQUEUERD_ADDR_REG_2_(vec[2490]), .P1_P3_INSTQUEUERD_ADDR_REG_1_(vec[2489]), .P1_P3_INSTQUEUERD_ADDR_REG_0_(vec[2488]), .P1_P3_INSTQUEUEWR_ADDR_REG_4_(vec[2487]), .P1_P3_INSTQUEUEWR_ADDR_REG_3_(vec[2486]), .P1_P3_INSTQUEUEWR_ADDR_REG_2_(vec[2485]), .P1_P3_INSTQUEUEWR_ADDR_REG_1_(vec[2484]), .P1_P3_INSTQUEUEWR_ADDR_REG_0_(vec[2483]), .P1_P3_INSTADDRPOINTER_REG_0_(vec[2482]), .P1_P3_INSTADDRPOINTER_REG_1_(vec[2481]), .P1_P3_INSTADDRPOINTER_REG_2_(vec[2480]), .P1_P3_INSTADDRPOINTER_REG_3_(vec[2479]), .P1_P3_INSTADDRPOINTER_REG_4_(vec[2478]), .P1_P3_INSTADDRPOINTER_REG_5_(vec[2477]), .P1_P3_INSTADDRPOINTER_REG_6_(vec[2476]), .P1_P3_INSTADDRPOINTER_REG_7_(vec[2475]), .P1_P3_INSTADDRPOINTER_REG_8_(vec[2474]), .P1_P3_INSTADDRPOINTER_REG_9_(vec[2473]), .P1_P3_INSTADDRPOINTER_REG_10_(vec[2472]), .P1_P3_INSTADDRPOINTER_REG_11_(vec[2471]), .P1_P3_INSTADDRPOINTER_REG_12_(vec[2470]), .P1_P3_INSTADDRPOINTER_REG_13_(vec[2469]), .P1_P3_INSTADDRPOINTER_REG_14_(vec[2468]), .P1_P3_INSTADDRPOINTER_REG_15_(vec[2467]), .P1_P3_INSTADDRPOINTER_REG_16_(vec[2466]), .P1_P3_INSTADDRPOINTER_REG_17_(vec[2465]), .P1_P3_INSTADDRPOINTER_REG_18_(vec[2464]), .P1_P3_INSTADDRPOINTER_REG_19_(vec[2463]), .P1_P3_INSTADDRPOINTER_REG_20_(vec[2462]), .P1_P3_INSTADDRPOINTER_REG_21_(vec[2461]), .P1_P3_INSTADDRPOINTER_REG_22_(vec[2460]), .P1_P3_INSTADDRPOINTER_REG_23_(vec[2459]), .P1_P3_INSTADDRPOINTER_REG_24_(vec[2458]), .P1_P3_INSTADDRPOINTER_REG_25_(vec[2457]), .P1_P3_INSTADDRPOINTER_REG_26_(vec[2456]), .P1_P3_INSTADDRPOINTER_REG_27_(vec[2455]), .P1_P3_INSTADDRPOINTER_REG_28_(vec[2454]), .P1_P3_INSTADDRPOINTER_REG_29_(vec[2453]), .P1_P3_INSTADDRPOINTER_REG_30_(vec[2452]), .P1_P3_INSTADDRPOINTER_REG_31_(vec[2451]), .P1_P3_PHYADDRPOINTER_REG_0_(vec[2450]), .P1_P3_PHYADDRPOINTER_REG_1_(vec[2449]), .P1_P3_PHYADDRPOINTER_REG_2_(vec[2448]), .P1_P3_PHYADDRPOINTER_REG_3_(vec[2447]), .P1_P3_PHYADDRPOINTER_REG_4_(vec[2446]), .P1_P3_PHYADDRPOINTER_REG_5_(vec[2445]), .P1_P3_PHYADDRPOINTER_REG_6_(vec[2444]), .P1_P3_PHYADDRPOINTER_REG_7_(vec[2443]), .P1_P3_PHYADDRPOINTER_REG_8_(vec[2442]), .P1_P3_PHYADDRPOINTER_REG_9_(vec[2441]), .P1_P3_PHYADDRPOINTER_REG_10_(vec[2440]), .P1_P3_PHYADDRPOINTER_REG_11_(vec[2439]), .P1_P3_PHYADDRPOINTER_REG_12_(vec[2438]), .P1_P3_PHYADDRPOINTER_REG_13_(vec[2437]), .P1_P3_PHYADDRPOINTER_REG_14_(vec[2436]), .P1_P3_PHYADDRPOINTER_REG_15_(vec[2435]), .P1_P3_PHYADDRPOINTER_REG_16_(vec[2434]), .P1_P3_PHYADDRPOINTER_REG_17_(vec[2433]), .P1_P3_PHYADDRPOINTER_REG_18_(vec[2432]), .P1_P3_PHYADDRPOINTER_REG_19_(vec[2431]), .P1_P3_PHYADDRPOINTER_REG_20_(vec[2430]), .P1_P3_PHYADDRPOINTER_REG_21_(vec[2429]), .P1_P3_PHYADDRPOINTER_REG_22_(vec[2428]), .P1_P3_PHYADDRPOINTER_REG_23_(vec[2427]), .P1_P3_PHYADDRPOINTER_REG_24_(vec[2426]), .P1_P3_PHYADDRPOINTER_REG_25_(vec[2425]), .P1_P3_PHYADDRPOINTER_REG_26_(vec[2424]), .P1_P3_PHYADDRPOINTER_REG_27_(vec[2423]), .P1_P3_PHYADDRPOINTER_REG_28_(vec[2422]), .P1_P3_PHYADDRPOINTER_REG_29_(vec[2421]), .P1_P3_PHYADDRPOINTER_REG_30_(vec[2420]), .P1_P3_PHYADDRPOINTER_REG_31_(vec[2419]), .P1_P3_LWORD_REG_15_(vec[2418]), .P1_P3_LWORD_REG_14_(vec[2417]), .P1_P3_LWORD_REG_13_(vec[2416]), .P1_P3_LWORD_REG_12_(vec[2415]), .P1_P3_LWORD_REG_11_(vec[2414]), .P1_P3_LWORD_REG_10_(vec[2413]), .P1_P3_LWORD_REG_9_(vec[2412]), .P1_P3_LWORD_REG_8_(vec[2411]), .P1_P3_LWORD_REG_7_(vec[2410]), .P1_P3_LWORD_REG_6_(vec[2409]), .P1_P3_LWORD_REG_5_(vec[2408]), .P1_P3_LWORD_REG_4_(vec[2407]), .P1_P3_LWORD_REG_3_(vec[2406]), .P1_P3_LWORD_REG_2_(vec[2405]), .P1_P3_LWORD_REG_1_(vec[2404]), .P1_P3_LWORD_REG_0_(vec[2403]), .P1_P3_UWORD_REG_14_(vec[2402]), .P1_P3_UWORD_REG_13_(vec[2401]), .P1_P3_UWORD_REG_12_(vec[2400]), .P1_P3_UWORD_REG_11_(vec[2399]), .P1_P3_UWORD_REG_10_(vec[2398]), .P1_P3_UWORD_REG_9_(vec[2397]), .P1_P3_UWORD_REG_8_(vec[2396]), .P1_P3_UWORD_REG_7_(vec[2395]), .P1_P3_UWORD_REG_6_(vec[2394]), .P1_P3_UWORD_REG_5_(vec[2393]), .P1_P3_UWORD_REG_4_(vec[2392]), .P1_P3_UWORD_REG_3_(vec[2391]), .P1_P3_UWORD_REG_2_(vec[2390]), .P1_P3_UWORD_REG_1_(vec[2389]), .P1_P3_UWORD_REG_0_(vec[2388]), .P1_P3_DATAO_REG_0_(vec[2387]), .P1_P3_DATAO_REG_1_(vec[2386]), .P1_P3_DATAO_REG_2_(vec[2385]), .P1_P3_DATAO_REG_3_(vec[2384]), .P1_P3_DATAO_REG_4_(vec[2383]), .P1_P3_DATAO_REG_5_(vec[2382]), .P1_P3_DATAO_REG_6_(vec[2381]), .P1_P3_DATAO_REG_7_(vec[2380]), .P1_P3_DATAO_REG_8_(vec[2379]), .P1_P3_DATAO_REG_9_(vec[2378]), .P1_P3_DATAO_REG_10_(vec[2377]), .P1_P3_DATAO_REG_11_(vec[2376]), .P1_P3_DATAO_REG_12_(vec[2375]), .P1_P3_DATAO_REG_13_(vec[2374]), .P1_P3_DATAO_REG_14_(vec[2373]), .P1_P3_DATAO_REG_15_(vec[2372]), .P1_P3_DATAO_REG_16_(vec[2371]), .P1_P3_DATAO_REG_17_(vec[2370]), .P1_P3_DATAO_REG_18_(vec[2369]), .P1_P3_DATAO_REG_19_(vec[2368]), .P1_P3_DATAO_REG_20_(vec[2367]), .P1_P3_DATAO_REG_21_(vec[2366]), .P1_P3_DATAO_REG_22_(vec[2365]), .P1_P3_DATAO_REG_23_(vec[2364]), .P1_P3_DATAO_REG_24_(vec[2363]), .P1_P3_DATAO_REG_25_(vec[2362]), .P1_P3_DATAO_REG_26_(vec[2361]), .P1_P3_DATAO_REG_27_(vec[2360]), .P1_P3_DATAO_REG_28_(vec[2359]), .P1_P3_DATAO_REG_29_(vec[2358]), .P1_P3_DATAO_REG_30_(vec[2357]), .P1_P3_DATAO_REG_31_(vec[2356]), .P1_P3_EAX_REG_0_(vec[2355]), .P1_P3_EAX_REG_1_(vec[2354]), .P1_P3_EAX_REG_2_(vec[2353]), .P1_P3_EAX_REG_3_(vec[2352]), .P1_P3_EAX_REG_4_(vec[2351]), .P1_P3_EAX_REG_5_(vec[2350]), .P1_P3_EAX_REG_6_(vec[2349]), .P1_P3_EAX_REG_7_(vec[2348]), .P1_P3_EAX_REG_8_(vec[2347]), .P1_P3_EAX_REG_9_(vec[2346]), .P1_P3_EAX_REG_10_(vec[2345]), .P1_P3_EAX_REG_11_(vec[2344]), .P1_P3_EAX_REG_12_(vec[2343]), .P1_P3_EAX_REG_13_(vec[2342]), .P1_P3_EAX_REG_14_(vec[2341]), .P1_P3_EAX_REG_15_(vec[2340]), .P1_P3_EAX_REG_16_(vec[2339]), .P1_P3_EAX_REG_17_(vec[2338]), .P1_P3_EAX_REG_18_(vec[2337]), .P1_P3_EAX_REG_19_(vec[2336]), .P1_P3_EAX_REG_20_(vec[2335]), .P1_P3_EAX_REG_21_(vec[2334]), .P1_P3_EAX_REG_22_(vec[2333]), .P1_P3_EAX_REG_23_(vec[2332]), .P1_P3_EAX_REG_24_(vec[2331]), .P1_P3_EAX_REG_25_(vec[2330]), .P1_P3_EAX_REG_26_(vec[2329]), .P1_P3_EAX_REG_27_(vec[2328]), .P1_P3_EAX_REG_28_(vec[2327]), .P1_P3_EAX_REG_29_(vec[2326]), .P1_P3_EAX_REG_30_(vec[2325]), .P1_P3_EAX_REG_31_(vec[2324]), .P1_P3_EBX_REG_0_(vec[2323]), .P1_P3_EBX_REG_1_(vec[2322]), .P1_P3_EBX_REG_2_(vec[2321]), .P1_P3_EBX_REG_3_(vec[2320]), .P1_P3_EBX_REG_4_(vec[2319]), .P1_P3_EBX_REG_5_(vec[2318]), .P1_P3_EBX_REG_6_(vec[2317]), .P1_P3_EBX_REG_7_(vec[2316]), .P1_P3_EBX_REG_8_(vec[2315]), .P1_P3_EBX_REG_9_(vec[2314]), .P1_P3_EBX_REG_10_(vec[2313]), .P1_P3_EBX_REG_11_(vec[2312]), .P1_P3_EBX_REG_12_(vec[2311]), .P1_P3_EBX_REG_13_(vec[2310]), .P1_P3_EBX_REG_14_(vec[2309]), .P1_P3_EBX_REG_15_(vec[2308]), .P1_P3_EBX_REG_16_(vec[2307]), .P1_P3_EBX_REG_17_(vec[2306]), .P1_P3_EBX_REG_18_(vec[2305]), .P1_P3_EBX_REG_19_(vec[2304]), .P1_P3_EBX_REG_20_(vec[2303]), .P1_P3_EBX_REG_21_(vec[2302]), .P1_P3_EBX_REG_22_(vec[2301]), .P1_P3_EBX_REG_23_(vec[2300]), .P1_P3_EBX_REG_24_(vec[2299]), .P1_P3_EBX_REG_25_(vec[2298]), .P1_P3_EBX_REG_26_(vec[2297]), .P1_P3_EBX_REG_27_(vec[2296]), .P1_P3_EBX_REG_28_(vec[2295]), .P1_P3_EBX_REG_29_(vec[2294]), .P1_P3_EBX_REG_30_(vec[2293]), .P1_P3_EBX_REG_31_(vec[2292]), .P1_P3_REIP_REG_0_(vec[2291]), .P1_P3_REIP_REG_1_(vec[2290]), .P1_P3_REIP_REG_2_(vec[2289]), .P1_P3_REIP_REG_3_(vec[2288]), .P1_P3_REIP_REG_4_(vec[2287]), .P1_P3_REIP_REG_5_(vec[2286]), .P1_P3_REIP_REG_6_(vec[2285]), .P1_P3_REIP_REG_7_(vec[2284]), .P1_P3_REIP_REG_8_(vec[2283]), .P1_P3_REIP_REG_9_(vec[2282]), .P1_P3_REIP_REG_10_(vec[2281]), .P1_P3_REIP_REG_11_(vec[2280]), .P1_P3_REIP_REG_12_(vec[2279]), .P1_P3_REIP_REG_13_(vec[2278]), .P1_P3_REIP_REG_14_(vec[2277]), .P1_P3_REIP_REG_15_(vec[2276]), .P1_P3_REIP_REG_16_(vec[2275]), .P1_P3_REIP_REG_17_(vec[2274]), .P1_P3_REIP_REG_18_(vec[2273]), .P1_P3_REIP_REG_19_(vec[2272]), .P1_P3_REIP_REG_20_(vec[2271]), .P1_P3_REIP_REG_21_(vec[2270]), .P1_P3_REIP_REG_22_(vec[2269]), .P1_P3_REIP_REG_23_(vec[2268]), .P1_P3_REIP_REG_24_(vec[2267]), .P1_P3_REIP_REG_25_(vec[2266]), .P1_P3_REIP_REG_26_(vec[2265]), .P1_P3_REIP_REG_27_(vec[2264]), .P1_P3_REIP_REG_28_(vec[2263]), .P1_P3_REIP_REG_29_(vec[2262]), .P1_P3_REIP_REG_30_(vec[2261]), .P1_P3_REIP_REG_31_(vec[2260]), .P1_P3_BYTEENABLE_REG_3_(vec[2259]), .P1_P3_BYTEENABLE_REG_2_(vec[2258]), .P1_P3_BYTEENABLE_REG_1_(vec[2257]), .P1_P3_BYTEENABLE_REG_0_(vec[2256]), .P1_P3_W_R_N_REG(vec[2255]), .P1_P3_FLUSH_REG(vec[2254]), .P1_P3_MORE_REG(vec[2253]), .P1_P3_STATEBS16_REG(vec[2252]), .P1_P3_REQUESTPENDING_REG(vec[2251]), .P1_P3_D_C_N_REG(vec[2250]), .P1_P3_M_IO_N_REG(vec[2249]), .P1_P3_CODEFETCH_REG(vec[2248]), .P1_P3_ADS_N_REG(vec[2247]), .P1_P3_READREQUEST_REG(vec[2246]), .P1_P3_MEMORYFETCH_REG(vec[2245]), .P1_P2_BE_N_REG_3_(vec[2244]), .P1_P2_BE_N_REG_2_(vec[2243]), .P1_P2_BE_N_REG_1_(vec[2242]), .P1_P2_BE_N_REG_0_(vec[2241]), .P1_P2_ADDRESS_REG_29_(vec[2240]), .P1_P2_ADDRESS_REG_28_(vec[2239]), .P1_P2_ADDRESS_REG_27_(vec[2238]), .P1_P2_ADDRESS_REG_26_(vec[2237]), .P1_P2_ADDRESS_REG_25_(vec[2236]), .P1_P2_ADDRESS_REG_24_(vec[2235]), .P1_P2_ADDRESS_REG_23_(vec[2234]), .P1_P2_ADDRESS_REG_22_(vec[2233]), .P1_P2_ADDRESS_REG_21_(vec[2232]), .P1_P2_ADDRESS_REG_20_(vec[2231]), .P1_P2_ADDRESS_REG_19_(vec[2230]), .P1_P2_ADDRESS_REG_18_(vec[2229]), .P1_P2_ADDRESS_REG_17_(vec[2228]), .P1_P2_ADDRESS_REG_16_(vec[2227]), .P1_P2_ADDRESS_REG_15_(vec[2226]), .P1_P2_ADDRESS_REG_14_(vec[2225]), .P1_P2_ADDRESS_REG_13_(vec[2224]), .P1_P2_ADDRESS_REG_12_(vec[2223]), .P1_P2_ADDRESS_REG_11_(vec[2222]), .P1_P2_ADDRESS_REG_10_(vec[2221]), .P1_P2_ADDRESS_REG_9_(vec[2220]), .P1_P2_ADDRESS_REG_8_(vec[2219]), .P1_P2_ADDRESS_REG_7_(vec[2218]), .P1_P2_ADDRESS_REG_6_(vec[2217]), .P1_P2_ADDRESS_REG_5_(vec[2216]), .P1_P2_ADDRESS_REG_4_(vec[2215]), .P1_P2_ADDRESS_REG_3_(vec[2214]), .P1_P2_ADDRESS_REG_2_(vec[2213]), .P1_P2_ADDRESS_REG_1_(vec[2212]), .P1_P2_ADDRESS_REG_0_(vec[2211]), .P1_P2_STATE_REG_2_(vec[2210]), .P1_P2_STATE_REG_1_(vec[2209]), .P1_P2_STATE_REG_0_(vec[2208]), .P1_P2_DATAWIDTH_REG_0_(vec[2207]), .P1_P2_DATAWIDTH_REG_1_(vec[2206]), .P1_P2_DATAWIDTH_REG_2_(vec[2205]), .P1_P2_DATAWIDTH_REG_3_(vec[2204]), .P1_P2_DATAWIDTH_REG_4_(vec[2203]), .P1_P2_DATAWIDTH_REG_5_(vec[2202]), .P1_P2_DATAWIDTH_REG_6_(vec[2201]), .P1_P2_DATAWIDTH_REG_7_(vec[2200]), .P1_P2_DATAWIDTH_REG_8_(vec[2199]), .P1_P2_DATAWIDTH_REG_9_(vec[2198]), .P1_P2_DATAWIDTH_REG_10_(vec[2197]), .P1_P2_DATAWIDTH_REG_11_(vec[2196]), .P1_P2_DATAWIDTH_REG_12_(vec[2195]), .P1_P2_DATAWIDTH_REG_13_(vec[2194]), .P1_P2_DATAWIDTH_REG_14_(vec[2193]), .P1_P2_DATAWIDTH_REG_15_(vec[2192]), .P1_P2_DATAWIDTH_REG_16_(vec[2191]), .P1_P2_DATAWIDTH_REG_17_(vec[2190]), .P1_P2_DATAWIDTH_REG_18_(vec[2189]), .P1_P2_DATAWIDTH_REG_19_(vec[2188]), .P1_P2_DATAWIDTH_REG_20_(vec[2187]), .P1_P2_DATAWIDTH_REG_21_(vec[2186]), .P1_P2_DATAWIDTH_REG_22_(vec[2185]), .P1_P2_DATAWIDTH_REG_23_(vec[2184]), .P1_P2_DATAWIDTH_REG_24_(vec[2183]), .P1_P2_DATAWIDTH_REG_25_(vec[2182]), .P1_P2_DATAWIDTH_REG_26_(vec[2181]), .P1_P2_DATAWIDTH_REG_27_(vec[2180]), .P1_P2_DATAWIDTH_REG_28_(vec[2179]), .P1_P2_DATAWIDTH_REG_29_(vec[2178]), .P1_P2_DATAWIDTH_REG_30_(vec[2177]), .P1_P2_DATAWIDTH_REG_31_(vec[2176]), .P1_P2_STATE2_REG_3_(vec[2175]), .P1_P2_STATE2_REG_2_(vec[2174]), .P1_P2_STATE2_REG_1_(vec[2173]), .P1_P2_STATE2_REG_0_(vec[2172]), .P1_P2_INSTQUEUE_REG_15__7_(vec[2171]), .P1_P2_INSTQUEUE_REG_15__6_(vec[2170]), .P1_P2_INSTQUEUE_REG_15__5_(vec[2169]), .P1_P2_INSTQUEUE_REG_15__4_(vec[2168]), .P1_P2_INSTQUEUE_REG_15__3_(vec[2167]), .P1_P2_INSTQUEUE_REG_15__2_(vec[2166]), .P1_P2_INSTQUEUE_REG_15__1_(vec[2165]), .P1_P2_INSTQUEUE_REG_15__0_(vec[2164]), .P1_P2_INSTQUEUE_REG_14__7_(vec[2163]), .P1_P2_INSTQUEUE_REG_14__6_(vec[2162]), .P1_P2_INSTQUEUE_REG_14__5_(vec[2161]), .P1_P2_INSTQUEUE_REG_14__4_(vec[2160]), .P1_P2_INSTQUEUE_REG_14__3_(vec[2159]), .P1_P2_INSTQUEUE_REG_14__2_(vec[2158]), .P1_P2_INSTQUEUE_REG_14__1_(vec[2157]), .P1_P2_INSTQUEUE_REG_14__0_(vec[2156]), .P1_P2_INSTQUEUE_REG_13__7_(vec[2155]), .P1_P2_INSTQUEUE_REG_13__6_(vec[2154]), .P1_P2_INSTQUEUE_REG_13__5_(vec[2153]), .P1_P2_INSTQUEUE_REG_13__4_(vec[2152]), .P1_P2_INSTQUEUE_REG_13__3_(vec[2151]), .P1_P2_INSTQUEUE_REG_13__2_(vec[2150]), .P1_P2_INSTQUEUE_REG_13__1_(vec[2149]), .P1_P2_INSTQUEUE_REG_13__0_(vec[2148]), .P1_P2_INSTQUEUE_REG_12__7_(vec[2147]), .P1_P2_INSTQUEUE_REG_12__6_(vec[2146]), .P1_P2_INSTQUEUE_REG_12__5_(vec[2145]), .P1_P2_INSTQUEUE_REG_12__4_(vec[2144]), .P1_P2_INSTQUEUE_REG_12__3_(vec[2143]), .P1_P2_INSTQUEUE_REG_12__2_(vec[2142]), .P1_P2_INSTQUEUE_REG_12__1_(vec[2141]), .P1_P2_INSTQUEUE_REG_12__0_(vec[2140]), .P1_P2_INSTQUEUE_REG_11__7_(vec[2139]), .P1_P2_INSTQUEUE_REG_11__6_(vec[2138]), .P1_P2_INSTQUEUE_REG_11__5_(vec[2137]), .P1_P2_INSTQUEUE_REG_11__4_(vec[2136]), .P1_P2_INSTQUEUE_REG_11__3_(vec[2135]), .P1_P2_INSTQUEUE_REG_11__2_(vec[2134]), .P1_P2_INSTQUEUE_REG_11__1_(vec[2133]), .P1_P2_INSTQUEUE_REG_11__0_(vec[2132]), .P1_P2_INSTQUEUE_REG_10__7_(vec[2131]), .P1_P2_INSTQUEUE_REG_10__6_(vec[2130]), .P1_P2_INSTQUEUE_REG_10__5_(vec[2129]), .P1_P2_INSTQUEUE_REG_10__4_(vec[2128]), .P1_P2_INSTQUEUE_REG_10__3_(vec[2127]), .P1_P2_INSTQUEUE_REG_10__2_(vec[2126]), .P1_P2_INSTQUEUE_REG_10__1_(vec[2125]), .P1_P2_INSTQUEUE_REG_10__0_(vec[2124]), .P1_P2_INSTQUEUE_REG_9__7_(vec[2123]), .P1_P2_INSTQUEUE_REG_9__6_(vec[2122]), .P1_P2_INSTQUEUE_REG_9__5_(vec[2121]), .P1_P2_INSTQUEUE_REG_9__4_(vec[2120]), .P1_P2_INSTQUEUE_REG_9__3_(vec[2119]), .P1_P2_INSTQUEUE_REG_9__2_(vec[2118]), .P1_P2_INSTQUEUE_REG_9__1_(vec[2117]), .P1_P2_INSTQUEUE_REG_9__0_(vec[2116]), .P1_P2_INSTQUEUE_REG_8__7_(vec[2115]), .P1_P2_INSTQUEUE_REG_8__6_(vec[2114]), .P1_P2_INSTQUEUE_REG_8__5_(vec[2113]), .P1_P2_INSTQUEUE_REG_8__4_(vec[2112]), .P1_P2_INSTQUEUE_REG_8__3_(vec[2111]), .P1_P2_INSTQUEUE_REG_8__2_(vec[2110]), .P1_P2_INSTQUEUE_REG_8__1_(vec[2109]), .P1_P2_INSTQUEUE_REG_8__0_(vec[2108]), .P1_P2_INSTQUEUE_REG_7__7_(vec[2107]), .P1_P2_INSTQUEUE_REG_7__6_(vec[2106]), .P1_P2_INSTQUEUE_REG_7__5_(vec[2105]), .P1_P2_INSTQUEUE_REG_7__4_(vec[2104]), .P1_P2_INSTQUEUE_REG_7__3_(vec[2103]), .P1_P2_INSTQUEUE_REG_7__2_(vec[2102]), .P1_P2_INSTQUEUE_REG_7__1_(vec[2101]), .P1_P2_INSTQUEUE_REG_7__0_(vec[2100]), .P1_P2_INSTQUEUE_REG_6__7_(vec[2099]), .P1_P2_INSTQUEUE_REG_6__6_(vec[2098]), .P1_P2_INSTQUEUE_REG_6__5_(vec[2097]), .P1_P2_INSTQUEUE_REG_6__4_(vec[2096]), .P1_P2_INSTQUEUE_REG_6__3_(vec[2095]), .P1_P2_INSTQUEUE_REG_6__2_(vec[2094]), .P1_P2_INSTQUEUE_REG_6__1_(vec[2093]), .P1_P2_INSTQUEUE_REG_6__0_(vec[2092]), .P1_P2_INSTQUEUE_REG_5__7_(vec[2091]), .P1_P2_INSTQUEUE_REG_5__6_(vec[2090]), .P1_P2_INSTQUEUE_REG_5__5_(vec[2089]), .P1_P2_INSTQUEUE_REG_5__4_(vec[2088]), .P1_P2_INSTQUEUE_REG_5__3_(vec[2087]), .P1_P2_INSTQUEUE_REG_5__2_(vec[2086]), .P1_P2_INSTQUEUE_REG_5__1_(vec[2085]), .P1_P2_INSTQUEUE_REG_5__0_(vec[2084]), .P1_P2_INSTQUEUE_REG_4__7_(vec[2083]), .P1_P2_INSTQUEUE_REG_4__6_(vec[2082]), .P1_P2_INSTQUEUE_REG_4__5_(vec[2081]), .P1_P2_INSTQUEUE_REG_4__4_(vec[2080]), .P1_P2_INSTQUEUE_REG_4__3_(vec[2079]), .P1_P2_INSTQUEUE_REG_4__2_(vec[2078]), .P1_P2_INSTQUEUE_REG_4__1_(vec[2077]), .P1_P2_INSTQUEUE_REG_4__0_(vec[2076]), .P1_P2_INSTQUEUE_REG_3__7_(vec[2075]), .P1_P2_INSTQUEUE_REG_3__6_(vec[2074]), .P1_P2_INSTQUEUE_REG_3__5_(vec[2073]), .P1_P2_INSTQUEUE_REG_3__4_(vec[2072]), .P1_P2_INSTQUEUE_REG_3__3_(vec[2071]), .P1_P2_INSTQUEUE_REG_3__2_(vec[2070]), .P1_P2_INSTQUEUE_REG_3__1_(vec[2069]), .P1_P2_INSTQUEUE_REG_3__0_(vec[2068]), .P1_P2_INSTQUEUE_REG_2__7_(vec[2067]), .P1_P2_INSTQUEUE_REG_2__6_(vec[2066]), .P1_P2_INSTQUEUE_REG_2__5_(vec[2065]), .P1_P2_INSTQUEUE_REG_2__4_(vec[2064]), .P1_P2_INSTQUEUE_REG_2__3_(vec[2063]), .P1_P2_INSTQUEUE_REG_2__2_(vec[2062]), .P1_P2_INSTQUEUE_REG_2__1_(vec[2061]), .P1_P2_INSTQUEUE_REG_2__0_(vec[2060]), .P1_P2_INSTQUEUE_REG_1__7_(vec[2059]), .P1_P2_INSTQUEUE_REG_1__6_(vec[2058]), .P1_P2_INSTQUEUE_REG_1__5_(vec[2057]), .P1_P2_INSTQUEUE_REG_1__4_(vec[2056]), .P1_P2_INSTQUEUE_REG_1__3_(vec[2055]), .P1_P2_INSTQUEUE_REG_1__2_(vec[2054]), .P1_P2_INSTQUEUE_REG_1__1_(vec[2053]), .P1_P2_INSTQUEUE_REG_1__0_(vec[2052]), .P1_P2_INSTQUEUE_REG_0__7_(vec[2051]), .P1_P2_INSTQUEUE_REG_0__6_(vec[2050]), .P1_P2_INSTQUEUE_REG_0__5_(vec[2049]), .P1_P2_INSTQUEUE_REG_0__4_(vec[2048]), .P1_P2_INSTQUEUE_REG_0__3_(vec[2047]), .P1_P2_INSTQUEUE_REG_0__2_(vec[2046]), .P1_P2_INSTQUEUE_REG_0__1_(vec[2045]), .P1_P2_INSTQUEUE_REG_0__0_(vec[2044]), .P1_P2_INSTQUEUERD_ADDR_REG_4_(vec[2043]), .P1_P2_INSTQUEUERD_ADDR_REG_3_(vec[2042]), .P1_P2_INSTQUEUERD_ADDR_REG_2_(vec[2041]), .P1_P2_INSTQUEUERD_ADDR_REG_1_(vec[2040]), .P1_P2_INSTQUEUERD_ADDR_REG_0_(vec[2039]), .P1_P2_INSTQUEUEWR_ADDR_REG_4_(vec[2038]), .P1_P2_INSTQUEUEWR_ADDR_REG_3_(vec[2037]), .P1_P2_INSTQUEUEWR_ADDR_REG_2_(vec[2036]), .P1_P2_INSTQUEUEWR_ADDR_REG_1_(vec[2035]), .P1_P2_INSTQUEUEWR_ADDR_REG_0_(vec[2034]), .P1_P2_INSTADDRPOINTER_REG_0_(vec[2033]), .P1_P2_INSTADDRPOINTER_REG_1_(vec[2032]), .P1_P2_INSTADDRPOINTER_REG_2_(vec[2031]), .P1_P2_INSTADDRPOINTER_REG_3_(vec[2030]), .P1_P2_INSTADDRPOINTER_REG_4_(vec[2029]), .P1_P2_INSTADDRPOINTER_REG_5_(vec[2028]), .P1_P2_INSTADDRPOINTER_REG_6_(vec[2027]), .P1_P2_INSTADDRPOINTER_REG_7_(vec[2026]), .P1_P2_INSTADDRPOINTER_REG_8_(vec[2025]), .P1_P2_INSTADDRPOINTER_REG_9_(vec[2024]), .P1_P2_INSTADDRPOINTER_REG_10_(vec[2023]), .P1_P2_INSTADDRPOINTER_REG_11_(vec[2022]), .P1_P2_INSTADDRPOINTER_REG_12_(vec[2021]), .P1_P2_INSTADDRPOINTER_REG_13_(vec[2020]), .P1_P2_INSTADDRPOINTER_REG_14_(vec[2019]), .P1_P2_INSTADDRPOINTER_REG_15_(vec[2018]), .P1_P2_INSTADDRPOINTER_REG_16_(vec[2017]), .P1_P2_INSTADDRPOINTER_REG_17_(vec[2016]), .P1_P2_INSTADDRPOINTER_REG_18_(vec[2015]), .P1_P2_INSTADDRPOINTER_REG_19_(vec[2014]), .P1_P2_INSTADDRPOINTER_REG_20_(vec[2013]), .P1_P2_INSTADDRPOINTER_REG_21_(vec[2012]), .P1_P2_INSTADDRPOINTER_REG_22_(vec[2011]), .P1_P2_INSTADDRPOINTER_REG_23_(vec[2010]), .P1_P2_INSTADDRPOINTER_REG_24_(vec[2009]), .P1_P2_INSTADDRPOINTER_REG_25_(vec[2008]), .P1_P2_INSTADDRPOINTER_REG_26_(vec[2007]), .P1_P2_INSTADDRPOINTER_REG_27_(vec[2006]), .P1_P2_INSTADDRPOINTER_REG_28_(vec[2005]), .P1_P2_INSTADDRPOINTER_REG_29_(vec[2004]), .P1_P2_INSTADDRPOINTER_REG_30_(vec[2003]), .P1_P2_INSTADDRPOINTER_REG_31_(vec[2002]), .P1_P2_PHYADDRPOINTER_REG_0_(vec[2001]), .P1_P2_PHYADDRPOINTER_REG_1_(vec[2000]), .P1_P2_PHYADDRPOINTER_REG_2_(vec[1999]), .P1_P2_PHYADDRPOINTER_REG_3_(vec[1998]), .P1_P2_PHYADDRPOINTER_REG_4_(vec[1997]), .P1_P2_PHYADDRPOINTER_REG_5_(vec[1996]), .P1_P2_PHYADDRPOINTER_REG_6_(vec[1995]), .P1_P2_PHYADDRPOINTER_REG_7_(vec[1994]), .P1_P2_PHYADDRPOINTER_REG_8_(vec[1993]), .P1_P2_PHYADDRPOINTER_REG_9_(vec[1992]), .P1_P2_PHYADDRPOINTER_REG_10_(vec[1991]), .P1_P2_PHYADDRPOINTER_REG_11_(vec[1990]), .P1_P2_PHYADDRPOINTER_REG_12_(vec[1989]), .P1_P2_PHYADDRPOINTER_REG_13_(vec[1988]), .P1_P2_PHYADDRPOINTER_REG_14_(vec[1987]), .P1_P2_PHYADDRPOINTER_REG_15_(vec[1986]), .P1_P2_PHYADDRPOINTER_REG_16_(vec[1985]), .P1_P2_PHYADDRPOINTER_REG_17_(vec[1984]), .P1_P2_PHYADDRPOINTER_REG_18_(vec[1983]), .P1_P2_PHYADDRPOINTER_REG_19_(vec[1982]), .P1_P2_PHYADDRPOINTER_REG_20_(vec[1981]), .P1_P2_PHYADDRPOINTER_REG_21_(vec[1980]), .P1_P2_PHYADDRPOINTER_REG_22_(vec[1979]), .P1_P2_PHYADDRPOINTER_REG_23_(vec[1978]), .P1_P2_PHYADDRPOINTER_REG_24_(vec[1977]), .P1_P2_PHYADDRPOINTER_REG_25_(vec[1976]), .P1_P2_PHYADDRPOINTER_REG_26_(vec[1975]), .P1_P2_PHYADDRPOINTER_REG_27_(vec[1974]), .P1_P2_PHYADDRPOINTER_REG_28_(vec[1973]), .P1_P2_PHYADDRPOINTER_REG_29_(vec[1972]), .P1_P2_PHYADDRPOINTER_REG_30_(vec[1971]), .P1_P2_PHYADDRPOINTER_REG_31_(vec[1970]), .P1_P2_LWORD_REG_15_(vec[1969]), .P1_P2_LWORD_REG_14_(vec[1968]), .P1_P2_LWORD_REG_13_(vec[1967]), .P1_P2_LWORD_REG_12_(vec[1966]), .P1_P2_LWORD_REG_11_(vec[1965]), .P1_P2_LWORD_REG_10_(vec[1964]), .P1_P2_LWORD_REG_9_(vec[1963]), .P1_P2_LWORD_REG_8_(vec[1962]), .P1_P2_LWORD_REG_7_(vec[1961]), .P1_P2_LWORD_REG_6_(vec[1960]), .P1_P2_LWORD_REG_5_(vec[1959]), .P1_P2_LWORD_REG_4_(vec[1958]), .P1_P2_LWORD_REG_3_(vec[1957]), .P1_P2_LWORD_REG_2_(vec[1956]), .P1_P2_LWORD_REG_1_(vec[1955]), .P1_P2_LWORD_REG_0_(vec[1954]), .P1_P2_UWORD_REG_14_(vec[1953]), .P1_P2_UWORD_REG_13_(vec[1952]), .P1_P2_UWORD_REG_12_(vec[1951]), .P1_P2_UWORD_REG_11_(vec[1950]), .P1_P2_UWORD_REG_10_(vec[1949]), .P1_P2_UWORD_REG_9_(vec[1948]), .P1_P2_UWORD_REG_8_(vec[1947]), .P1_P2_UWORD_REG_7_(vec[1946]), .P1_P2_UWORD_REG_6_(vec[1945]), .P1_P2_UWORD_REG_5_(vec[1944]), .P1_P2_UWORD_REG_4_(vec[1943]), .P1_P2_UWORD_REG_3_(vec[1942]), .P1_P2_UWORD_REG_2_(vec[1941]), .P1_P2_UWORD_REG_1_(vec[1940]), .P1_P2_UWORD_REG_0_(vec[1939]), .P1_P2_DATAO_REG_0_(vec[1938]), .P1_P2_DATAO_REG_1_(vec[1937]), .P1_P2_DATAO_REG_2_(vec[1936]), .P1_P2_DATAO_REG_3_(vec[1935]), .P1_P2_DATAO_REG_4_(vec[1934]), .P1_P2_DATAO_REG_5_(vec[1933]), .P1_P2_DATAO_REG_6_(vec[1932]), .P1_P2_DATAO_REG_7_(vec[1931]), .P1_P2_DATAO_REG_8_(vec[1930]), .P1_P2_DATAO_REG_9_(vec[1929]), .P1_P2_DATAO_REG_10_(vec[1928]), .P1_P2_DATAO_REG_11_(vec[1927]), .P1_P2_DATAO_REG_12_(vec[1926]), .P1_P2_DATAO_REG_13_(vec[1925]), .P1_P2_DATAO_REG_14_(vec[1924]), .P1_P2_DATAO_REG_15_(vec[1923]), .P1_P2_DATAO_REG_16_(vec[1922]), .P1_P2_DATAO_REG_17_(vec[1921]), .P1_P2_DATAO_REG_18_(vec[1920]), .P1_P2_DATAO_REG_19_(vec[1919]), .P1_P2_DATAO_REG_20_(vec[1918]), .P1_P2_DATAO_REG_21_(vec[1917]), .P1_P2_DATAO_REG_22_(vec[1916]), .P1_P2_DATAO_REG_23_(vec[1915]), .P1_P2_DATAO_REG_24_(vec[1914]), .P1_P2_DATAO_REG_25_(vec[1913]), .P1_P2_DATAO_REG_26_(vec[1912]), .P1_P2_DATAO_REG_27_(vec[1911]), .P1_P2_DATAO_REG_28_(vec[1910]), .P1_P2_DATAO_REG_29_(vec[1909]), .P1_P2_DATAO_REG_30_(vec[1908]), .P1_P2_DATAO_REG_31_(vec[1907]), .P1_P2_EAX_REG_0_(vec[1906]), .P1_P2_EAX_REG_1_(vec[1905]), .P1_P2_EAX_REG_2_(vec[1904]), .P1_P2_EAX_REG_3_(vec[1903]), .P1_P2_EAX_REG_4_(vec[1902]), .P1_P2_EAX_REG_5_(vec[1901]), .P1_P2_EAX_REG_6_(vec[1900]), .P1_P2_EAX_REG_7_(vec[1899]), .P1_P2_EAX_REG_8_(vec[1898]), .P1_P2_EAX_REG_9_(vec[1897]), .P1_P2_EAX_REG_10_(vec[1896]), .P1_P2_EAX_REG_11_(vec[1895]), .P1_P2_EAX_REG_12_(vec[1894]), .P1_P2_EAX_REG_13_(vec[1893]), .P1_P2_EAX_REG_14_(vec[1892]), .P1_P2_EAX_REG_15_(vec[1891]), .P1_P2_EAX_REG_16_(vec[1890]), .P1_P2_EAX_REG_17_(vec[1889]), .P1_P2_EAX_REG_18_(vec[1888]), .P1_P2_EAX_REG_19_(vec[1887]), .P1_P2_EAX_REG_20_(vec[1886]), .P1_P2_EAX_REG_21_(vec[1885]), .P1_P2_EAX_REG_22_(vec[1884]), .P1_P2_EAX_REG_23_(vec[1883]), .P1_P2_EAX_REG_24_(vec[1882]), .P1_P2_EAX_REG_25_(vec[1881]), .P1_P2_EAX_REG_26_(vec[1880]), .P1_P2_EAX_REG_27_(vec[1879]), .P1_P2_EAX_REG_28_(vec[1878]), .P1_P2_EAX_REG_29_(vec[1877]), .P1_P2_EAX_REG_30_(vec[1876]), .P1_P2_EAX_REG_31_(vec[1875]), .P1_P2_EBX_REG_0_(vec[1874]), .P1_P2_EBX_REG_1_(vec[1873]), .P1_P2_EBX_REG_2_(vec[1872]), .P1_P2_EBX_REG_3_(vec[1871]), .P1_P2_EBX_REG_4_(vec[1870]), .P1_P2_EBX_REG_5_(vec[1869]), .P1_P2_EBX_REG_6_(vec[1868]), .P1_P2_EBX_REG_7_(vec[1867]), .P1_P2_EBX_REG_8_(vec[1866]), .P1_P2_EBX_REG_9_(vec[1865]), .P1_P2_EBX_REG_10_(vec[1864]), .P1_P2_EBX_REG_11_(vec[1863]), .P1_P2_EBX_REG_12_(vec[1862]), .P1_P2_EBX_REG_13_(vec[1861]), .P1_P2_EBX_REG_14_(vec[1860]), .P1_P2_EBX_REG_15_(vec[1859]), .P1_P2_EBX_REG_16_(vec[1858]), .P1_P2_EBX_REG_17_(vec[1857]), .P1_P2_EBX_REG_18_(vec[1856]), .P1_P2_EBX_REG_19_(vec[1855]), .P1_P2_EBX_REG_20_(vec[1854]), .P1_P2_EBX_REG_21_(vec[1853]), .P1_P2_EBX_REG_22_(vec[1852]), .P1_P2_EBX_REG_23_(vec[1851]), .P1_P2_EBX_REG_24_(vec[1850]), .P1_P2_EBX_REG_25_(vec[1849]), .P1_P2_EBX_REG_26_(vec[1848]), .P1_P2_EBX_REG_27_(vec[1847]), .P1_P2_EBX_REG_28_(vec[1846]), .P1_P2_EBX_REG_29_(vec[1845]), .P1_P2_EBX_REG_30_(vec[1844]), .P1_P2_EBX_REG_31_(vec[1843]), .P1_P2_REIP_REG_0_(vec[1842]), .P1_P2_REIP_REG_1_(vec[1841]), .P1_P2_REIP_REG_2_(vec[1840]), .P1_P2_REIP_REG_3_(vec[1839]), .P1_P2_REIP_REG_4_(vec[1838]), .P1_P2_REIP_REG_5_(vec[1837]), .P1_P2_REIP_REG_6_(vec[1836]), .P1_P2_REIP_REG_7_(vec[1835]), .P1_P2_REIP_REG_8_(vec[1834]), .P1_P2_REIP_REG_9_(vec[1833]), .P1_P2_REIP_REG_10_(vec[1832]), .P1_P2_REIP_REG_11_(vec[1831]), .P1_P2_REIP_REG_12_(vec[1830]), .P1_P2_REIP_REG_13_(vec[1829]), .P1_P2_REIP_REG_14_(vec[1828]), .P1_P2_REIP_REG_15_(vec[1827]), .P1_P2_REIP_REG_16_(vec[1826]), .P1_P2_REIP_REG_17_(vec[1825]), .P1_P2_REIP_REG_18_(vec[1824]), .P1_P2_REIP_REG_19_(vec[1823]), .P1_P2_REIP_REG_20_(vec[1822]), .P1_P2_REIP_REG_21_(vec[1821]), .P1_P2_REIP_REG_22_(vec[1820]), .P1_P2_REIP_REG_23_(vec[1819]), .P1_P2_REIP_REG_24_(vec[1818]), .P1_P2_REIP_REG_25_(vec[1817]), .P1_P2_REIP_REG_26_(vec[1816]), .P1_P2_REIP_REG_27_(vec[1815]), .P1_P2_REIP_REG_28_(vec[1814]), .P1_P2_REIP_REG_29_(vec[1813]), .P1_P2_REIP_REG_30_(vec[1812]), .P1_P2_REIP_REG_31_(vec[1811]), .P1_P2_BYTEENABLE_REG_3_(vec[1810]), .P1_P2_BYTEENABLE_REG_2_(vec[1809]), .P1_P2_BYTEENABLE_REG_1_(vec[1808]), .P1_P2_BYTEENABLE_REG_0_(vec[1807]), .P1_P2_W_R_N_REG(vec[1806]), .P1_P2_FLUSH_REG(vec[1805]), .P1_P2_MORE_REG(vec[1804]), .P1_P2_STATEBS16_REG(vec[1803]), .P1_P2_REQUESTPENDING_REG(vec[1802]), .P1_P2_D_C_N_REG(vec[1801]), .P1_P2_M_IO_N_REG(vec[1800]), .P1_P2_CODEFETCH_REG(vec[1799]), .P1_P2_ADS_N_REG(vec[1798]), .P1_P2_READREQUEST_REG(vec[1797]), .P1_P2_MEMORYFETCH_REG(vec[1796]), .P1_P1_BE_N_REG_3_(vec[1795]), .P1_P1_BE_N_REG_2_(vec[1794]), .P1_P1_BE_N_REG_1_(vec[1793]), .P1_P1_BE_N_REG_0_(vec[1792]), .P1_P1_ADDRESS_REG_29_(vec[1791]), .P1_P1_ADDRESS_REG_28_(vec[1790]), .P1_P1_ADDRESS_REG_27_(vec[1789]), .P1_P1_ADDRESS_REG_26_(vec[1788]), .P1_P1_ADDRESS_REG_25_(vec[1787]), .P1_P1_ADDRESS_REG_24_(vec[1786]), .P1_P1_ADDRESS_REG_23_(vec[1785]), .P1_P1_ADDRESS_REG_22_(vec[1784]), .P1_P1_ADDRESS_REG_21_(vec[1783]), .P1_P1_ADDRESS_REG_20_(vec[1782]), .P1_P1_ADDRESS_REG_19_(vec[1781]), .P1_P1_ADDRESS_REG_18_(vec[1780]), .P1_P1_ADDRESS_REG_17_(vec[1779]), .P1_P1_ADDRESS_REG_16_(vec[1778]), .P1_P1_ADDRESS_REG_15_(vec[1777]), .P1_P1_ADDRESS_REG_14_(vec[1776]), .P1_P1_ADDRESS_REG_13_(vec[1775]), .P1_P1_ADDRESS_REG_12_(vec[1774]), .P1_P1_ADDRESS_REG_11_(vec[1773]), .P1_P1_ADDRESS_REG_10_(vec[1772]), .P1_P1_ADDRESS_REG_9_(vec[1771]), .P1_P1_ADDRESS_REG_8_(vec[1770]), .P1_P1_ADDRESS_REG_7_(vec[1769]), .P1_P1_ADDRESS_REG_6_(vec[1768]), .P1_P1_ADDRESS_REG_5_(vec[1767]), .P1_P1_ADDRESS_REG_4_(vec[1766]), .P1_P1_ADDRESS_REG_3_(vec[1765]), .P1_P1_ADDRESS_REG_2_(vec[1764]), .P1_P1_ADDRESS_REG_1_(vec[1763]), .P1_P1_ADDRESS_REG_0_(vec[1762]), .P1_P1_STATE_REG_2_(vec[1761]), .P1_P1_STATE_REG_1_(vec[1760]), .P1_P1_STATE_REG_0_(vec[1759]), .P1_P1_DATAWIDTH_REG_0_(vec[1758]), .P1_P1_DATAWIDTH_REG_1_(vec[1757]), .P1_P1_DATAWIDTH_REG_2_(vec[1756]), .P1_P1_DATAWIDTH_REG_3_(vec[1755]), .P1_P1_DATAWIDTH_REG_4_(vec[1754]), .P1_P1_DATAWIDTH_REG_5_(vec[1753]), .P1_P1_DATAWIDTH_REG_6_(vec[1752]), .P1_P1_DATAWIDTH_REG_7_(vec[1751]), .P1_P1_DATAWIDTH_REG_8_(vec[1750]), .P1_P1_DATAWIDTH_REG_9_(vec[1749]), .P1_P1_DATAWIDTH_REG_10_(vec[1748]), .P1_P1_DATAWIDTH_REG_11_(vec[1747]), .P1_P1_DATAWIDTH_REG_12_(vec[1746]), .P1_P1_DATAWIDTH_REG_13_(vec[1745]), .P1_P1_DATAWIDTH_REG_14_(vec[1744]), .P1_P1_DATAWIDTH_REG_15_(vec[1743]), .P1_P1_DATAWIDTH_REG_16_(vec[1742]), .P1_P1_DATAWIDTH_REG_17_(vec[1741]), .P1_P1_DATAWIDTH_REG_18_(vec[1740]), .P1_P1_DATAWIDTH_REG_19_(vec[1739]), .P1_P1_DATAWIDTH_REG_20_(vec[1738]), .P1_P1_DATAWIDTH_REG_21_(vec[1737]), .P1_P1_DATAWIDTH_REG_22_(vec[1736]), .P1_P1_DATAWIDTH_REG_23_(vec[1735]), .P1_P1_DATAWIDTH_REG_24_(vec[1734]), .P1_P1_DATAWIDTH_REG_25_(vec[1733]), .P1_P1_DATAWIDTH_REG_26_(vec[1732]), .P1_P1_DATAWIDTH_REG_27_(vec[1731]), .P1_P1_DATAWIDTH_REG_28_(vec[1730]), .P1_P1_DATAWIDTH_REG_29_(vec[1729]), .P1_P1_DATAWIDTH_REG_30_(vec[1728]), .P1_P1_DATAWIDTH_REG_31_(vec[1727]), .P1_P1_STATE2_REG_3_(vec[1726]), .P1_P1_STATE2_REG_2_(vec[1725]), .P1_P1_STATE2_REG_1_(vec[1724]), .P1_P1_STATE2_REG_0_(vec[1723]), .P1_P1_INSTQUEUE_REG_15__7_(vec[1722]), .P1_P1_INSTQUEUE_REG_15__6_(vec[1721]), .P1_P1_INSTQUEUE_REG_15__5_(vec[1720]), .P1_P1_INSTQUEUE_REG_15__4_(vec[1719]), .P1_P1_INSTQUEUE_REG_15__3_(vec[1718]), .P1_P1_INSTQUEUE_REG_15__2_(vec[1717]), .P1_P1_INSTQUEUE_REG_15__1_(vec[1716]), .P1_P1_INSTQUEUE_REG_15__0_(vec[1715]), .P1_P1_INSTQUEUE_REG_14__7_(vec[1714]), .P1_P1_INSTQUEUE_REG_14__6_(vec[1713]), .P1_P1_INSTQUEUE_REG_14__5_(vec[1712]), .P1_P1_INSTQUEUE_REG_14__4_(vec[1711]), .P1_P1_INSTQUEUE_REG_14__3_(vec[1710]), .P1_P1_INSTQUEUE_REG_14__2_(vec[1709]), .P1_P1_INSTQUEUE_REG_14__1_(vec[1708]), .P1_P1_INSTQUEUE_REG_14__0_(vec[1707]), .P1_P1_INSTQUEUE_REG_13__7_(vec[1706]), .P1_P1_INSTQUEUE_REG_13__6_(vec[1705]), .P1_P1_INSTQUEUE_REG_13__5_(vec[1704]), .P1_P1_INSTQUEUE_REG_13__4_(vec[1703]), .P1_P1_INSTQUEUE_REG_13__3_(vec[1702]), .P1_P1_INSTQUEUE_REG_13__2_(vec[1701]), .P1_P1_INSTQUEUE_REG_13__1_(vec[1700]), .P1_P1_INSTQUEUE_REG_13__0_(vec[1699]), .P1_P1_INSTQUEUE_REG_12__7_(vec[1698]), .P1_P1_INSTQUEUE_REG_12__6_(vec[1697]), .P1_P1_INSTQUEUE_REG_12__5_(vec[1696]), .P1_P1_INSTQUEUE_REG_12__4_(vec[1695]), .P1_P1_INSTQUEUE_REG_12__3_(vec[1694]), .P1_P1_INSTQUEUE_REG_12__2_(vec[1693]), .P1_P1_INSTQUEUE_REG_12__1_(vec[1692]), .P1_P1_INSTQUEUE_REG_12__0_(vec[1691]), .P1_P1_INSTQUEUE_REG_11__7_(vec[1690]), .P1_P1_INSTQUEUE_REG_11__6_(vec[1689]), .P1_P1_INSTQUEUE_REG_11__5_(vec[1688]), .P1_P1_INSTQUEUE_REG_11__4_(vec[1687]), .P1_P1_INSTQUEUE_REG_11__3_(vec[1686]), .P1_P1_INSTQUEUE_REG_11__2_(vec[1685]), .P1_P1_INSTQUEUE_REG_11__1_(vec[1684]), .P1_P1_INSTQUEUE_REG_11__0_(vec[1683]), .P1_P1_INSTQUEUE_REG_10__7_(vec[1682]), .P1_P1_INSTQUEUE_REG_10__6_(vec[1681]), .P1_P1_INSTQUEUE_REG_10__5_(vec[1680]), .P1_P1_INSTQUEUE_REG_10__4_(vec[1679]), .P1_P1_INSTQUEUE_REG_10__3_(vec[1678]), .P1_P1_INSTQUEUE_REG_10__2_(vec[1677]), .P1_P1_INSTQUEUE_REG_10__1_(vec[1676]), .P1_P1_INSTQUEUE_REG_10__0_(vec[1675]), .P1_P1_INSTQUEUE_REG_9__7_(vec[1674]), .P1_P1_INSTQUEUE_REG_9__6_(vec[1673]), .P1_P1_INSTQUEUE_REG_9__5_(vec[1672]), .P1_P1_INSTQUEUE_REG_9__4_(vec[1671]), .P1_P1_INSTQUEUE_REG_9__3_(vec[1670]), .P1_P1_INSTQUEUE_REG_9__2_(vec[1669]), .P1_P1_INSTQUEUE_REG_9__1_(vec[1668]), .P1_P1_INSTQUEUE_REG_9__0_(vec[1667]), .P1_P1_INSTQUEUE_REG_8__7_(vec[1666]), .P1_P1_INSTQUEUE_REG_8__6_(vec[1665]), .P1_P1_INSTQUEUE_REG_8__5_(vec[1664]), .P1_P1_INSTQUEUE_REG_8__4_(vec[1663]), .P1_P1_INSTQUEUE_REG_8__3_(vec[1662]), .P1_P1_INSTQUEUE_REG_8__2_(vec[1661]), .P1_P1_INSTQUEUE_REG_8__1_(vec[1660]), .P1_P1_INSTQUEUE_REG_8__0_(vec[1659]), .P1_P1_INSTQUEUE_REG_7__7_(vec[1658]), .P1_P1_INSTQUEUE_REG_7__6_(vec[1657]), .P1_P1_INSTQUEUE_REG_7__5_(vec[1656]), .P1_P1_INSTQUEUE_REG_7__4_(vec[1655]), .P1_P1_INSTQUEUE_REG_7__3_(vec[1654]), .P1_P1_INSTQUEUE_REG_7__2_(vec[1653]), .P1_P1_INSTQUEUE_REG_7__1_(vec[1652]), .P1_P1_INSTQUEUE_REG_7__0_(vec[1651]), .P1_P1_INSTQUEUE_REG_6__7_(vec[1650]), .P1_P1_INSTQUEUE_REG_6__6_(vec[1649]), .P1_P1_INSTQUEUE_REG_6__5_(vec[1648]), .P1_P1_INSTQUEUE_REG_6__4_(vec[1647]), .P1_P1_INSTQUEUE_REG_6__3_(vec[1646]), .P1_P1_INSTQUEUE_REG_6__2_(vec[1645]), .P1_P1_INSTQUEUE_REG_6__1_(vec[1644]), .P1_P1_INSTQUEUE_REG_6__0_(vec[1643]), .P1_P1_INSTQUEUE_REG_5__7_(vec[1642]), .P1_P1_INSTQUEUE_REG_5__6_(vec[1641]), .P1_P1_INSTQUEUE_REG_5__5_(vec[1640]), .P1_P1_INSTQUEUE_REG_5__4_(vec[1639]), .P1_P1_INSTQUEUE_REG_5__3_(vec[1638]), .P1_P1_INSTQUEUE_REG_5__2_(vec[1637]), .P1_P1_INSTQUEUE_REG_5__1_(vec[1636]), .P1_P1_INSTQUEUE_REG_5__0_(vec[1635]), .P1_P1_INSTQUEUE_REG_4__7_(vec[1634]), .P1_P1_INSTQUEUE_REG_4__6_(vec[1633]), .P1_P1_INSTQUEUE_REG_4__5_(vec[1632]), .P1_P1_INSTQUEUE_REG_4__4_(vec[1631]), .P1_P1_INSTQUEUE_REG_4__3_(vec[1630]), .P1_P1_INSTQUEUE_REG_4__2_(vec[1629]), .P1_P1_INSTQUEUE_REG_4__1_(vec[1628]), .P1_P1_INSTQUEUE_REG_4__0_(vec[1627]), .P1_P1_INSTQUEUE_REG_3__7_(vec[1626]), .P1_P1_INSTQUEUE_REG_3__6_(vec[1625]), .P1_P1_INSTQUEUE_REG_3__5_(vec[1624]), .P1_P1_INSTQUEUE_REG_3__4_(vec[1623]), .P1_P1_INSTQUEUE_REG_3__3_(vec[1622]), .P1_P1_INSTQUEUE_REG_3__2_(vec[1621]), .P1_P1_INSTQUEUE_REG_3__1_(vec[1620]), .P1_P1_INSTQUEUE_REG_3__0_(vec[1619]), .P1_P1_INSTQUEUE_REG_2__7_(vec[1618]), .P1_P1_INSTQUEUE_REG_2__6_(vec[1617]), .P1_P1_INSTQUEUE_REG_2__5_(vec[1616]), .P1_P1_INSTQUEUE_REG_2__4_(vec[1615]), .P1_P1_INSTQUEUE_REG_2__3_(vec[1614]), .P1_P1_INSTQUEUE_REG_2__2_(vec[1613]), .P1_P1_INSTQUEUE_REG_2__1_(vec[1612]), .P1_P1_INSTQUEUE_REG_2__0_(vec[1611]), .P1_P1_INSTQUEUE_REG_1__7_(vec[1610]), .P1_P1_INSTQUEUE_REG_1__6_(vec[1609]), .P1_P1_INSTQUEUE_REG_1__5_(vec[1608]), .P1_P1_INSTQUEUE_REG_1__4_(vec[1607]), .P1_P1_INSTQUEUE_REG_1__3_(vec[1606]), .P1_P1_INSTQUEUE_REG_1__2_(vec[1605]), .P1_P1_INSTQUEUE_REG_1__1_(vec[1604]), .P1_P1_INSTQUEUE_REG_1__0_(vec[1603]), .P1_P1_INSTQUEUE_REG_0__7_(vec[1602]), .P1_P1_INSTQUEUE_REG_0__6_(vec[1601]), .P1_P1_INSTQUEUE_REG_0__5_(vec[1600]), .P1_P1_INSTQUEUE_REG_0__4_(vec[1599]), .P1_P1_INSTQUEUE_REG_0__3_(vec[1598]), .P1_P1_INSTQUEUE_REG_0__2_(vec[1597]), .P1_P1_INSTQUEUE_REG_0__1_(vec[1596]), .P1_P1_INSTQUEUE_REG_0__0_(vec[1595]), .P1_P1_INSTQUEUERD_ADDR_REG_4_(vec[1594]), .P1_P1_INSTQUEUERD_ADDR_REG_3_(vec[1593]), .P1_P1_INSTQUEUERD_ADDR_REG_2_(vec[1592]), .P1_P1_INSTQUEUERD_ADDR_REG_1_(vec[1591]), .P1_P1_INSTQUEUERD_ADDR_REG_0_(vec[1590]), .P1_P1_INSTQUEUEWR_ADDR_REG_4_(vec[1589]), .P1_P1_INSTQUEUEWR_ADDR_REG_3_(vec[1588]), .P1_P1_INSTQUEUEWR_ADDR_REG_2_(vec[1587]), .P1_P1_INSTQUEUEWR_ADDR_REG_1_(vec[1586]), .P1_P1_INSTQUEUEWR_ADDR_REG_0_(vec[1585]), .P1_P1_INSTADDRPOINTER_REG_0_(vec[1584]), .P1_P1_INSTADDRPOINTER_REG_1_(vec[1583]), .P1_P1_INSTADDRPOINTER_REG_2_(vec[1582]), .P1_P1_INSTADDRPOINTER_REG_3_(vec[1581]), .P1_P1_INSTADDRPOINTER_REG_4_(vec[1580]), .P1_P1_INSTADDRPOINTER_REG_5_(vec[1579]), .P1_P1_INSTADDRPOINTER_REG_6_(vec[1578]), .P1_P1_INSTADDRPOINTER_REG_7_(vec[1577]), .P1_P1_INSTADDRPOINTER_REG_8_(vec[1576]), .P1_P1_INSTADDRPOINTER_REG_9_(vec[1575]), .P1_P1_INSTADDRPOINTER_REG_10_(vec[1574]), .P1_P1_INSTADDRPOINTER_REG_11_(vec[1573]), .P1_P1_INSTADDRPOINTER_REG_12_(vec[1572]), .P1_P1_INSTADDRPOINTER_REG_13_(vec[1571]), .P1_P1_INSTADDRPOINTER_REG_14_(vec[1570]), .P1_P1_INSTADDRPOINTER_REG_15_(vec[1569]), .P1_P1_INSTADDRPOINTER_REG_16_(vec[1568]), .P1_P1_INSTADDRPOINTER_REG_17_(vec[1567]), .P1_P1_INSTADDRPOINTER_REG_18_(vec[1566]), .P1_P1_INSTADDRPOINTER_REG_19_(vec[1565]), .P1_P1_INSTADDRPOINTER_REG_20_(vec[1564]), .P1_P1_INSTADDRPOINTER_REG_21_(vec[1563]), .P1_P1_INSTADDRPOINTER_REG_22_(vec[1562]), .P1_P1_INSTADDRPOINTER_REG_23_(vec[1561]), .P1_P1_INSTADDRPOINTER_REG_24_(vec[1560]), .P1_P1_INSTADDRPOINTER_REG_25_(vec[1559]), .P1_P1_INSTADDRPOINTER_REG_26_(vec[1558]), .P1_P1_INSTADDRPOINTER_REG_27_(vec[1557]), .P1_P1_INSTADDRPOINTER_REG_28_(vec[1556]), .P1_P1_INSTADDRPOINTER_REG_29_(vec[1555]), .P1_P1_INSTADDRPOINTER_REG_30_(vec[1554]), .P1_P1_INSTADDRPOINTER_REG_31_(vec[1553]), .P1_P1_PHYADDRPOINTER_REG_0_(vec[1552]), .P1_P1_PHYADDRPOINTER_REG_1_(vec[1551]), .P1_P1_PHYADDRPOINTER_REG_2_(vec[1550]), .P1_P1_PHYADDRPOINTER_REG_3_(vec[1549]), .P1_P1_PHYADDRPOINTER_REG_4_(vec[1548]), .P1_P1_PHYADDRPOINTER_REG_5_(vec[1547]), .P1_P1_PHYADDRPOINTER_REG_6_(vec[1546]), .P1_P1_PHYADDRPOINTER_REG_7_(vec[1545]), .P1_P1_PHYADDRPOINTER_REG_8_(vec[1544]), .P1_P1_PHYADDRPOINTER_REG_9_(vec[1543]), .P1_P1_PHYADDRPOINTER_REG_10_(vec[1542]), .P1_P1_PHYADDRPOINTER_REG_11_(vec[1541]), .P1_P1_PHYADDRPOINTER_REG_12_(vec[1540]), .P1_P1_PHYADDRPOINTER_REG_13_(vec[1539]), .P1_P1_PHYADDRPOINTER_REG_14_(vec[1538]), .P1_P1_PHYADDRPOINTER_REG_15_(vec[1537]), .P1_P1_PHYADDRPOINTER_REG_16_(vec[1536]), .P1_P1_PHYADDRPOINTER_REG_17_(vec[1535]), .P1_P1_PHYADDRPOINTER_REG_18_(vec[1534]), .P1_P1_PHYADDRPOINTER_REG_19_(vec[1533]), .P1_P1_PHYADDRPOINTER_REG_20_(vec[1532]), .P1_P1_PHYADDRPOINTER_REG_21_(vec[1531]), .P1_P1_PHYADDRPOINTER_REG_22_(vec[1530]), .P1_P1_PHYADDRPOINTER_REG_23_(vec[1529]), .P1_P1_PHYADDRPOINTER_REG_24_(vec[1528]), .P1_P1_PHYADDRPOINTER_REG_25_(vec[1527]), .P1_P1_PHYADDRPOINTER_REG_26_(vec[1526]), .P1_P1_PHYADDRPOINTER_REG_27_(vec[1525]), .P1_P1_PHYADDRPOINTER_REG_28_(vec[1524]), .P1_P1_PHYADDRPOINTER_REG_29_(vec[1523]), .P1_P1_PHYADDRPOINTER_REG_30_(vec[1522]), .P1_P1_PHYADDRPOINTER_REG_31_(vec[1521]), .P1_P1_LWORD_REG_15_(vec[1520]), .P1_P1_LWORD_REG_14_(vec[1519]), .P1_P1_LWORD_REG_13_(vec[1518]), .P1_P1_LWORD_REG_12_(vec[1517]), .P1_P1_LWORD_REG_11_(vec[1516]), .P1_P1_LWORD_REG_10_(vec[1515]), .P1_P1_LWORD_REG_9_(vec[1514]), .P1_P1_LWORD_REG_8_(vec[1513]), .P1_P1_LWORD_REG_7_(vec[1512]), .P1_P1_LWORD_REG_6_(vec[1511]), .P1_P1_LWORD_REG_5_(vec[1510]), .P1_P1_LWORD_REG_4_(vec[1509]), .P1_P1_LWORD_REG_3_(vec[1508]), .P1_P1_LWORD_REG_2_(vec[1507]), .P1_P1_LWORD_REG_1_(vec[1506]), .P1_P1_LWORD_REG_0_(vec[1505]), .P1_P1_UWORD_REG_14_(vec[1504]), .P1_P1_UWORD_REG_13_(vec[1503]), .P1_P1_UWORD_REG_12_(vec[1502]), .P1_P1_UWORD_REG_11_(vec[1501]), .P1_P1_UWORD_REG_10_(vec[1500]), .P1_P1_UWORD_REG_9_(vec[1499]), .P1_P1_UWORD_REG_8_(vec[1498]), .P1_P1_UWORD_REG_7_(vec[1497]), .P1_P1_UWORD_REG_6_(vec[1496]), .P1_P1_UWORD_REG_5_(vec[1495]), .P1_P1_UWORD_REG_4_(vec[1494]), .P1_P1_UWORD_REG_3_(vec[1493]), .P1_P1_UWORD_REG_2_(vec[1492]), .P1_P1_UWORD_REG_1_(vec[1491]), .P1_P1_UWORD_REG_0_(vec[1490]), .P1_P1_DATAO_REG_0_(vec[1489]), .P1_P1_DATAO_REG_1_(vec[1488]), .P1_P1_DATAO_REG_2_(vec[1487]), .P1_P1_DATAO_REG_3_(vec[1486]), .P1_P1_DATAO_REG_4_(vec[1485]), .P1_P1_DATAO_REG_5_(vec[1484]), .P1_P1_DATAO_REG_6_(vec[1483]), .P1_P1_DATAO_REG_7_(vec[1482]), .P1_P1_DATAO_REG_8_(vec[1481]), .P1_P1_DATAO_REG_9_(vec[1480]), .P1_P1_DATAO_REG_10_(vec[1479]), .P1_P1_DATAO_REG_11_(vec[1478]), .P1_P1_DATAO_REG_12_(vec[1477]), .P1_P1_DATAO_REG_13_(vec[1476]), .P1_P1_DATAO_REG_14_(vec[1475]), .P1_P1_DATAO_REG_15_(vec[1474]), .P1_P1_DATAO_REG_16_(vec[1473]), .P1_P1_DATAO_REG_17_(vec[1472]), .P1_P1_DATAO_REG_18_(vec[1471]), .P1_P1_DATAO_REG_19_(vec[1470]), .P1_P1_DATAO_REG_20_(vec[1469]), .P1_P1_DATAO_REG_21_(vec[1468]), .P1_P1_DATAO_REG_22_(vec[1467]), .P1_P1_DATAO_REG_23_(vec[1466]), .P1_P1_DATAO_REG_24_(vec[1465]), .P1_P1_DATAO_REG_25_(vec[1464]), .P1_P1_DATAO_REG_26_(vec[1463]), .P1_P1_DATAO_REG_27_(vec[1462]), .P1_P1_DATAO_REG_28_(vec[1461]), .P1_P1_DATAO_REG_29_(vec[1460]), .P1_P1_DATAO_REG_30_(vec[1459]), .P1_P1_DATAO_REG_31_(vec[1458]), .P1_P1_EAX_REG_0_(vec[1457]), .P1_P1_EAX_REG_1_(vec[1456]), .P1_P1_EAX_REG_2_(vec[1455]), .P1_P1_EAX_REG_3_(vec[1454]), .P1_P1_EAX_REG_4_(vec[1453]), .P1_P1_EAX_REG_5_(vec[1452]), .P1_P1_EAX_REG_6_(vec[1451]), .P1_P1_EAX_REG_7_(vec[1450]), .P1_P1_EAX_REG_8_(vec[1449]), .P1_P1_EAX_REG_9_(vec[1448]), .P1_P1_EAX_REG_10_(vec[1447]), .P1_P1_EAX_REG_11_(vec[1446]), .P1_P1_EAX_REG_12_(vec[1445]), .P1_P1_EAX_REG_13_(vec[1444]), .P1_P1_EAX_REG_14_(vec[1443]), .P1_P1_EAX_REG_15_(vec[1442]), .P1_P1_EAX_REG_16_(vec[1441]), .P1_P1_EAX_REG_17_(vec[1440]), .P1_P1_EAX_REG_18_(vec[1439]), .P1_P1_EAX_REG_19_(vec[1438]), .P1_P1_EAX_REG_20_(vec[1437]), .P1_P1_EAX_REG_21_(vec[1436]), .P1_P1_EAX_REG_22_(vec[1435]), .P1_P1_EAX_REG_23_(vec[1434]), .P1_P1_EAX_REG_24_(vec[1433]), .P1_P1_EAX_REG_25_(vec[1432]), .P1_P1_EAX_REG_26_(vec[1431]), .P1_P1_EAX_REG_27_(vec[1430]), .P1_P1_EAX_REG_28_(vec[1429]), .P1_P1_EAX_REG_29_(vec[1428]), .P1_P1_EAX_REG_30_(vec[1427]), .P1_P1_EAX_REG_31_(vec[1426]), .P1_P1_EBX_REG_0_(vec[1425]), .P1_P1_EBX_REG_1_(vec[1424]), .P1_P1_EBX_REG_2_(vec[1423]), .P1_P1_EBX_REG_3_(vec[1422]), .P1_P1_EBX_REG_4_(vec[1421]), .P1_P1_EBX_REG_5_(vec[1420]), .P1_P1_EBX_REG_6_(vec[1419]), .P1_P1_EBX_REG_7_(vec[1418]), .P1_P1_EBX_REG_8_(vec[1417]), .P1_P1_EBX_REG_9_(vec[1416]), .P1_P1_EBX_REG_10_(vec[1415]), .P1_P1_EBX_REG_11_(vec[1414]), .P1_P1_EBX_REG_12_(vec[1413]), .P1_P1_EBX_REG_13_(vec[1412]), .P1_P1_EBX_REG_14_(vec[1411]), .P1_P1_EBX_REG_15_(vec[1410]), .P1_P1_EBX_REG_16_(vec[1409]), .P1_P1_EBX_REG_17_(vec[1408]), .P1_P1_EBX_REG_18_(vec[1407]), .P1_P1_EBX_REG_19_(vec[1406]), .P1_P1_EBX_REG_20_(vec[1405]), .P1_P1_EBX_REG_21_(vec[1404]), .P1_P1_EBX_REG_22_(vec[1403]), .P1_P1_EBX_REG_23_(vec[1402]), .P1_P1_EBX_REG_24_(vec[1401]), .P1_P1_EBX_REG_25_(vec[1400]), .P1_P1_EBX_REG_26_(vec[1399]), .P1_P1_EBX_REG_27_(vec[1398]), .P1_P1_EBX_REG_28_(vec[1397]), .P1_P1_EBX_REG_29_(vec[1396]), .P1_P1_EBX_REG_30_(vec[1395]), .P1_P1_EBX_REG_31_(vec[1394]), .P1_P1_REIP_REG_0_(vec[1393]), .P1_P1_REIP_REG_1_(vec[1392]), .P1_P1_REIP_REG_2_(vec[1391]), .P1_P1_REIP_REG_3_(vec[1390]), .P1_P1_REIP_REG_4_(vec[1389]), .P1_P1_REIP_REG_5_(vec[1388]), .P1_P1_REIP_REG_6_(vec[1387]), .P1_P1_REIP_REG_7_(vec[1386]), .P1_P1_REIP_REG_8_(vec[1385]), .P1_P1_REIP_REG_9_(vec[1384]), .P1_P1_REIP_REG_10_(vec[1383]), .P1_P1_REIP_REG_11_(vec[1382]), .P1_P1_REIP_REG_12_(vec[1381]), .P1_P1_REIP_REG_13_(vec[1380]), .P1_P1_REIP_REG_14_(vec[1379]), .P1_P1_REIP_REG_15_(vec[1378]), .P1_P1_REIP_REG_16_(vec[1377]), .P1_P1_REIP_REG_17_(vec[1376]), .P1_P1_REIP_REG_18_(vec[1375]), .P1_P1_REIP_REG_19_(vec[1374]), .P1_P1_REIP_REG_20_(vec[1373]), .P1_P1_REIP_REG_21_(vec[1372]), .P1_P1_REIP_REG_22_(vec[1371]), .P1_P1_REIP_REG_23_(vec[1370]), .P1_P1_REIP_REG_24_(vec[1369]), .P1_P1_REIP_REG_25_(vec[1368]), .P1_P1_REIP_REG_26_(vec[1367]), .P1_P1_REIP_REG_27_(vec[1366]), .P1_P1_REIP_REG_28_(vec[1365]), .P1_P1_REIP_REG_29_(vec[1364]), .P1_P1_REIP_REG_30_(vec[1363]), .P1_P1_REIP_REG_31_(vec[1362]), .P1_P1_BYTEENABLE_REG_3_(vec[1361]), .P1_P1_BYTEENABLE_REG_2_(vec[1360]), .P1_P1_BYTEENABLE_REG_1_(vec[1359]), .P1_P1_BYTEENABLE_REG_0_(vec[1358]), .P1_P1_W_R_N_REG(vec[1357]), .P1_P1_FLUSH_REG(vec[1356]), .P1_P1_MORE_REG(vec[1355]), .P1_P1_STATEBS16_REG(vec[1354]), .P1_P1_REQUESTPENDING_REG(vec[1353]), .P1_P1_D_C_N_REG(vec[1352]), .P1_P1_M_IO_N_REG(vec[1351]), .P1_P1_CODEFETCH_REG(vec[1350]), .P1_P1_ADS_N_REG(vec[1349]), .P1_P1_READREQUEST_REG(vec[1348]), .P1_P1_MEMORYFETCH_REG(vec[1347]), .P2_P3_BE_N_REG_3_(vec[1346]), .P2_P3_BE_N_REG_2_(vec[1345]), .P2_P3_BE_N_REG_1_(vec[1344]), .P2_P3_BE_N_REG_0_(vec[1343]), .P2_P3_ADDRESS_REG_29_(vec[1342]), .P2_P3_ADDRESS_REG_28_(vec[1341]), .P2_P3_ADDRESS_REG_27_(vec[1340]), .P2_P3_ADDRESS_REG_26_(vec[1339]), .P2_P3_ADDRESS_REG_25_(vec[1338]), .P2_P3_ADDRESS_REG_24_(vec[1337]), .P2_P3_ADDRESS_REG_23_(vec[1336]), .P2_P3_ADDRESS_REG_22_(vec[1335]), .P2_P3_ADDRESS_REG_21_(vec[1334]), .P2_P3_ADDRESS_REG_20_(vec[1333]), .P2_P3_ADDRESS_REG_19_(vec[1332]), .P2_P3_ADDRESS_REG_18_(vec[1331]), .P2_P3_ADDRESS_REG_17_(vec[1330]), .P2_P3_ADDRESS_REG_16_(vec[1329]), .P2_P3_ADDRESS_REG_15_(vec[1328]), .P2_P3_ADDRESS_REG_14_(vec[1327]), .P2_P3_ADDRESS_REG_13_(vec[1326]), .P2_P3_ADDRESS_REG_12_(vec[1325]), .P2_P3_ADDRESS_REG_11_(vec[1324]), .P2_P3_ADDRESS_REG_10_(vec[1323]), .P2_P3_ADDRESS_REG_9_(vec[1322]), .P2_P3_ADDRESS_REG_8_(vec[1321]), .P2_P3_ADDRESS_REG_7_(vec[1320]), .P2_P3_ADDRESS_REG_6_(vec[1319]), .P2_P3_ADDRESS_REG_5_(vec[1318]), .P2_P3_ADDRESS_REG_4_(vec[1317]), .P2_P3_ADDRESS_REG_3_(vec[1316]), .P2_P3_ADDRESS_REG_2_(vec[1315]), .P2_P3_ADDRESS_REG_1_(vec[1314]), .P2_P3_ADDRESS_REG_0_(vec[1313]), .P2_P3_STATE_REG_2_(vec[1312]), .P2_P3_STATE_REG_1_(vec[1311]), .P2_P3_STATE_REG_0_(vec[1310]), .P2_P3_DATAWIDTH_REG_0_(vec[1309]), .P2_P3_DATAWIDTH_REG_1_(vec[1308]), .P2_P3_DATAWIDTH_REG_2_(vec[1307]), .P2_P3_DATAWIDTH_REG_3_(vec[1306]), .P2_P3_DATAWIDTH_REG_4_(vec[1305]), .P2_P3_DATAWIDTH_REG_5_(vec[1304]), .P2_P3_DATAWIDTH_REG_6_(vec[1303]), .P2_P3_DATAWIDTH_REG_7_(vec[1302]), .P2_P3_DATAWIDTH_REG_8_(vec[1301]), .P2_P3_DATAWIDTH_REG_9_(vec[1300]), .P2_P3_DATAWIDTH_REG_10_(vec[1299]), .P2_P3_DATAWIDTH_REG_11_(vec[1298]), .P2_P3_DATAWIDTH_REG_12_(vec[1297]), .P2_P3_DATAWIDTH_REG_13_(vec[1296]), .P2_P3_DATAWIDTH_REG_14_(vec[1295]), .P2_P3_DATAWIDTH_REG_15_(vec[1294]), .P2_P3_DATAWIDTH_REG_16_(vec[1293]), .P2_P3_DATAWIDTH_REG_17_(vec[1292]), .P2_P3_DATAWIDTH_REG_18_(vec[1291]), .P2_P3_DATAWIDTH_REG_19_(vec[1290]), .P2_P3_DATAWIDTH_REG_20_(vec[1289]), .P2_P3_DATAWIDTH_REG_21_(vec[1288]), .P2_P3_DATAWIDTH_REG_22_(vec[1287]), .P2_P3_DATAWIDTH_REG_23_(vec[1286]), .P2_P3_DATAWIDTH_REG_24_(vec[1285]), .P2_P3_DATAWIDTH_REG_25_(vec[1284]), .P2_P3_DATAWIDTH_REG_26_(vec[1283]), .P2_P3_DATAWIDTH_REG_27_(vec[1282]), .P2_P3_DATAWIDTH_REG_28_(vec[1281]), .P2_P3_DATAWIDTH_REG_29_(vec[1280]), .P2_P3_DATAWIDTH_REG_30_(vec[1279]), .P2_P3_DATAWIDTH_REG_31_(vec[1278]), .P2_P3_STATE2_REG_3_(vec[1277]), .P2_P3_STATE2_REG_2_(vec[1276]), .P2_P3_STATE2_REG_1_(vec[1275]), .P2_P3_STATE2_REG_0_(vec[1274]), .P2_P3_INSTQUEUE_REG_15__7_(vec[1273]), .P2_P3_INSTQUEUE_REG_15__6_(vec[1272]), .P2_P3_INSTQUEUE_REG_15__5_(vec[1271]), .P2_P3_INSTQUEUE_REG_15__4_(vec[1270]), .P2_P3_INSTQUEUE_REG_15__3_(vec[1269]), .P2_P3_INSTQUEUE_REG_15__2_(vec[1268]), .P2_P3_INSTQUEUE_REG_15__1_(vec[1267]), .P2_P3_INSTQUEUE_REG_15__0_(vec[1266]), .P2_P3_INSTQUEUE_REG_14__7_(vec[1265]), .P2_P3_INSTQUEUE_REG_14__6_(vec[1264]), .P2_P3_INSTQUEUE_REG_14__5_(vec[1263]), .P2_P3_INSTQUEUE_REG_14__4_(vec[1262]), .P2_P3_INSTQUEUE_REG_14__3_(vec[1261]), .P2_P3_INSTQUEUE_REG_14__2_(vec[1260]), .P2_P3_INSTQUEUE_REG_14__1_(vec[1259]), .P2_P3_INSTQUEUE_REG_14__0_(vec[1258]), .P2_P3_INSTQUEUE_REG_13__7_(vec[1257]), .P2_P3_INSTQUEUE_REG_13__6_(vec[1256]), .P2_P3_INSTQUEUE_REG_13__5_(vec[1255]), .P2_P3_INSTQUEUE_REG_13__4_(vec[1254]), .P2_P3_INSTQUEUE_REG_13__3_(vec[1253]), .P2_P3_INSTQUEUE_REG_13__2_(vec[1252]), .P2_P3_INSTQUEUE_REG_13__1_(vec[1251]), .P2_P3_INSTQUEUE_REG_13__0_(vec[1250]), .P2_P3_INSTQUEUE_REG_12__7_(vec[1249]), .P2_P3_INSTQUEUE_REG_12__6_(vec[1248]), .P2_P3_INSTQUEUE_REG_12__5_(vec[1247]), .P2_P3_INSTQUEUE_REG_12__4_(vec[1246]), .P2_P3_INSTQUEUE_REG_12__3_(vec[1245]), .P2_P3_INSTQUEUE_REG_12__2_(vec[1244]), .P2_P3_INSTQUEUE_REG_12__1_(vec[1243]), .P2_P3_INSTQUEUE_REG_12__0_(vec[1242]), .P2_P3_INSTQUEUE_REG_11__7_(vec[1241]), .P2_P3_INSTQUEUE_REG_11__6_(vec[1240]), .P2_P3_INSTQUEUE_REG_11__5_(vec[1239]), .P2_P3_INSTQUEUE_REG_11__4_(vec[1238]), .P2_P3_INSTQUEUE_REG_11__3_(vec[1237]), .P2_P3_INSTQUEUE_REG_11__2_(vec[1236]), .P2_P3_INSTQUEUE_REG_11__1_(vec[1235]), .P2_P3_INSTQUEUE_REG_11__0_(vec[1234]), .P2_P3_INSTQUEUE_REG_10__7_(vec[1233]), .P2_P3_INSTQUEUE_REG_10__6_(vec[1232]), .P2_P3_INSTQUEUE_REG_10__5_(vec[1231]), .P2_P3_INSTQUEUE_REG_10__4_(vec[1230]), .P2_P3_INSTQUEUE_REG_10__3_(vec[1229]), .P2_P3_INSTQUEUE_REG_10__2_(vec[1228]), .P2_P3_INSTQUEUE_REG_10__1_(vec[1227]), .P2_P3_INSTQUEUE_REG_10__0_(vec[1226]), .P2_P3_INSTQUEUE_REG_9__7_(vec[1225]), .P2_P3_INSTQUEUE_REG_9__6_(vec[1224]), .P2_P3_INSTQUEUE_REG_9__5_(vec[1223]), .P2_P3_INSTQUEUE_REG_9__4_(vec[1222]), .P2_P3_INSTQUEUE_REG_9__3_(vec[1221]), .P2_P3_INSTQUEUE_REG_9__2_(vec[1220]), .P2_P3_INSTQUEUE_REG_9__1_(vec[1219]), .P2_P3_INSTQUEUE_REG_9__0_(vec[1218]), .P2_P3_INSTQUEUE_REG_8__7_(vec[1217]), .P2_P3_INSTQUEUE_REG_8__6_(vec[1216]), .P2_P3_INSTQUEUE_REG_8__5_(vec[1215]), .P2_P3_INSTQUEUE_REG_8__4_(vec[1214]), .P2_P3_INSTQUEUE_REG_8__3_(vec[1213]), .P2_P3_INSTQUEUE_REG_8__2_(vec[1212]), .P2_P3_INSTQUEUE_REG_8__1_(vec[1211]), .P2_P3_INSTQUEUE_REG_8__0_(vec[1210]), .P2_P3_INSTQUEUE_REG_7__7_(vec[1209]), .P2_P3_INSTQUEUE_REG_7__6_(vec[1208]), .P2_P3_INSTQUEUE_REG_7__5_(vec[1207]), .P2_P3_INSTQUEUE_REG_7__4_(vec[1206]), .P2_P3_INSTQUEUE_REG_7__3_(vec[1205]), .P2_P3_INSTQUEUE_REG_7__2_(vec[1204]), .P2_P3_INSTQUEUE_REG_7__1_(vec[1203]), .P2_P3_INSTQUEUE_REG_7__0_(vec[1202]), .P2_P3_INSTQUEUE_REG_6__7_(vec[1201]), .P2_P3_INSTQUEUE_REG_6__6_(vec[1200]), .P2_P3_INSTQUEUE_REG_6__5_(vec[1199]), .P2_P3_INSTQUEUE_REG_6__4_(vec[1198]), .P2_P3_INSTQUEUE_REG_6__3_(vec[1197]), .P2_P3_INSTQUEUE_REG_6__2_(vec[1196]), .P2_P3_INSTQUEUE_REG_6__1_(vec[1195]), .P2_P3_INSTQUEUE_REG_6__0_(vec[1194]), .P2_P3_INSTQUEUE_REG_5__7_(vec[1193]), .P2_P3_INSTQUEUE_REG_5__6_(vec[1192]), .P2_P3_INSTQUEUE_REG_5__5_(vec[1191]), .P2_P3_INSTQUEUE_REG_5__4_(vec[1190]), .P2_P3_INSTQUEUE_REG_5__3_(vec[1189]), .P2_P3_INSTQUEUE_REG_5__2_(vec[1188]), .P2_P3_INSTQUEUE_REG_5__1_(vec[1187]), .P2_P3_INSTQUEUE_REG_5__0_(vec[1186]), .P2_P3_INSTQUEUE_REG_4__7_(vec[1185]), .P2_P3_INSTQUEUE_REG_4__6_(vec[1184]), .P2_P3_INSTQUEUE_REG_4__5_(vec[1183]), .P2_P3_INSTQUEUE_REG_4__4_(vec[1182]), .P2_P3_INSTQUEUE_REG_4__3_(vec[1181]), .P2_P3_INSTQUEUE_REG_4__2_(vec[1180]), .P2_P3_INSTQUEUE_REG_4__1_(vec[1179]), .P2_P3_INSTQUEUE_REG_4__0_(vec[1178]), .P2_P3_INSTQUEUE_REG_3__7_(vec[1177]), .P2_P3_INSTQUEUE_REG_3__6_(vec[1176]), .P2_P3_INSTQUEUE_REG_3__5_(vec[1175]), .P2_P3_INSTQUEUE_REG_3__4_(vec[1174]), .P2_P3_INSTQUEUE_REG_3__3_(vec[1173]), .P2_P3_INSTQUEUE_REG_3__2_(vec[1172]), .P2_P3_INSTQUEUE_REG_3__1_(vec[1171]), .P2_P3_INSTQUEUE_REG_3__0_(vec[1170]), .P2_P3_INSTQUEUE_REG_2__7_(vec[1169]), .P2_P3_INSTQUEUE_REG_2__6_(vec[1168]), .P2_P3_INSTQUEUE_REG_2__5_(vec[1167]), .P2_P3_INSTQUEUE_REG_2__4_(vec[1166]), .P2_P3_INSTQUEUE_REG_2__3_(vec[1165]), .P2_P3_INSTQUEUE_REG_2__2_(vec[1164]), .P2_P3_INSTQUEUE_REG_2__1_(vec[1163]), .P2_P3_INSTQUEUE_REG_2__0_(vec[1162]), .P2_P3_INSTQUEUE_REG_1__7_(vec[1161]), .P2_P3_INSTQUEUE_REG_1__6_(vec[1160]), .P2_P3_INSTQUEUE_REG_1__5_(vec[1159]), .P2_P3_INSTQUEUE_REG_1__4_(vec[1158]), .P2_P3_INSTQUEUE_REG_1__3_(vec[1157]), .P2_P3_INSTQUEUE_REG_1__2_(vec[1156]), .P2_P3_INSTQUEUE_REG_1__1_(vec[1155]), .P2_P3_INSTQUEUE_REG_1__0_(vec[1154]), .P2_P3_INSTQUEUE_REG_0__7_(vec[1153]), .P2_P3_INSTQUEUE_REG_0__6_(vec[1152]), .P2_P3_INSTQUEUE_REG_0__5_(vec[1151]), .P2_P3_INSTQUEUE_REG_0__4_(vec[1150]), .P2_P3_INSTQUEUE_REG_0__3_(vec[1149]), .P2_P3_INSTQUEUE_REG_0__2_(vec[1148]), .P2_P3_INSTQUEUE_REG_0__1_(vec[1147]), .P2_P3_INSTQUEUE_REG_0__0_(vec[1146]), .P2_P3_INSTQUEUERD_ADDR_REG_4_(vec[1145]), .P2_P3_INSTQUEUERD_ADDR_REG_3_(vec[1144]), .P2_P3_INSTQUEUERD_ADDR_REG_2_(vec[1143]), .P2_P3_INSTQUEUERD_ADDR_REG_1_(vec[1142]), .P2_P3_INSTQUEUERD_ADDR_REG_0_(vec[1141]), .P2_P3_INSTQUEUEWR_ADDR_REG_4_(vec[1140]), .P2_P3_INSTQUEUEWR_ADDR_REG_3_(vec[1139]), .P2_P3_INSTQUEUEWR_ADDR_REG_2_(vec[1138]), .P2_P3_INSTQUEUEWR_ADDR_REG_1_(vec[1137]), .P2_P3_INSTQUEUEWR_ADDR_REG_0_(vec[1136]), .P2_P3_INSTADDRPOINTER_REG_0_(vec[1135]), .P2_P3_INSTADDRPOINTER_REG_1_(vec[1134]), .P2_P3_INSTADDRPOINTER_REG_2_(vec[1133]), .P2_P3_INSTADDRPOINTER_REG_3_(vec[1132]), .P2_P3_INSTADDRPOINTER_REG_4_(vec[1131]), .P2_P3_INSTADDRPOINTER_REG_5_(vec[1130]), .P2_P3_INSTADDRPOINTER_REG_6_(vec[1129]), .P2_P3_INSTADDRPOINTER_REG_7_(vec[1128]), .P2_P3_INSTADDRPOINTER_REG_8_(vec[1127]), .P2_P3_INSTADDRPOINTER_REG_9_(vec[1126]), .P2_P3_INSTADDRPOINTER_REG_10_(vec[1125]), .P2_P3_INSTADDRPOINTER_REG_11_(vec[1124]), .P2_P3_INSTADDRPOINTER_REG_12_(vec[1123]), .P2_P3_INSTADDRPOINTER_REG_13_(vec[1122]), .P2_P3_INSTADDRPOINTER_REG_14_(vec[1121]), .P2_P3_INSTADDRPOINTER_REG_15_(vec[1120]), .P2_P3_INSTADDRPOINTER_REG_16_(vec[1119]), .P2_P3_INSTADDRPOINTER_REG_17_(vec[1118]), .P2_P3_INSTADDRPOINTER_REG_18_(vec[1117]), .P2_P3_INSTADDRPOINTER_REG_19_(vec[1116]), .P2_P3_INSTADDRPOINTER_REG_20_(vec[1115]), .P2_P3_INSTADDRPOINTER_REG_21_(vec[1114]), .P2_P3_INSTADDRPOINTER_REG_22_(vec[1113]), .P2_P3_INSTADDRPOINTER_REG_23_(vec[1112]), .P2_P3_INSTADDRPOINTER_REG_24_(vec[1111]), .P2_P3_INSTADDRPOINTER_REG_25_(vec[1110]), .P2_P3_INSTADDRPOINTER_REG_26_(vec[1109]), .P2_P3_INSTADDRPOINTER_REG_27_(vec[1108]), .P2_P3_INSTADDRPOINTER_REG_28_(vec[1107]), .P2_P3_INSTADDRPOINTER_REG_29_(vec[1106]), .P2_P3_INSTADDRPOINTER_REG_30_(vec[1105]), .P2_P3_INSTADDRPOINTER_REG_31_(vec[1104]), .P2_P3_PHYADDRPOINTER_REG_0_(vec[1103]), .P2_P3_PHYADDRPOINTER_REG_1_(vec[1102]), .P2_P3_PHYADDRPOINTER_REG_2_(vec[1101]), .P2_P3_PHYADDRPOINTER_REG_3_(vec[1100]), .P2_P3_PHYADDRPOINTER_REG_4_(vec[1099]), .P2_P3_PHYADDRPOINTER_REG_5_(vec[1098]), .P2_P3_PHYADDRPOINTER_REG_6_(vec[1097]), .P2_P3_PHYADDRPOINTER_REG_7_(vec[1096]), .P2_P3_PHYADDRPOINTER_REG_8_(vec[1095]), .P2_P3_PHYADDRPOINTER_REG_9_(vec[1094]), .P2_P3_PHYADDRPOINTER_REG_10_(vec[1093]), .P2_P3_PHYADDRPOINTER_REG_11_(vec[1092]), .P2_P3_PHYADDRPOINTER_REG_12_(vec[1091]), .P2_P3_PHYADDRPOINTER_REG_13_(vec[1090]), .P2_P3_PHYADDRPOINTER_REG_14_(vec[1089]), .P2_P3_PHYADDRPOINTER_REG_15_(vec[1088]), .P2_P3_PHYADDRPOINTER_REG_16_(vec[1087]), .P2_P3_PHYADDRPOINTER_REG_17_(vec[1086]), .P2_P3_PHYADDRPOINTER_REG_18_(vec[1085]), .P2_P3_PHYADDRPOINTER_REG_19_(vec[1084]), .P2_P3_PHYADDRPOINTER_REG_20_(vec[1083]), .P2_P3_PHYADDRPOINTER_REG_21_(vec[1082]), .P2_P3_PHYADDRPOINTER_REG_22_(vec[1081]), .P2_P3_PHYADDRPOINTER_REG_23_(vec[1080]), .P2_P3_PHYADDRPOINTER_REG_24_(vec[1079]), .P2_P3_PHYADDRPOINTER_REG_25_(vec[1078]), .P2_P3_PHYADDRPOINTER_REG_26_(vec[1077]), .P2_P3_PHYADDRPOINTER_REG_27_(vec[1076]), .P2_P3_PHYADDRPOINTER_REG_28_(vec[1075]), .P2_P3_PHYADDRPOINTER_REG_29_(vec[1074]), .P2_P3_PHYADDRPOINTER_REG_30_(vec[1073]), .P2_P3_PHYADDRPOINTER_REG_31_(vec[1072]), .P2_P3_LWORD_REG_15_(vec[1071]), .P2_P3_LWORD_REG_14_(vec[1070]), .P2_P3_LWORD_REG_13_(vec[1069]), .P2_P3_LWORD_REG_12_(vec[1068]), .P2_P3_LWORD_REG_11_(vec[1067]), .P2_P3_LWORD_REG_10_(vec[1066]), .P2_P3_LWORD_REG_9_(vec[1065]), .P2_P3_LWORD_REG_8_(vec[1064]), .P2_P3_LWORD_REG_7_(vec[1063]), .P2_P3_LWORD_REG_6_(vec[1062]), .P2_P3_LWORD_REG_5_(vec[1061]), .P2_P3_LWORD_REG_4_(vec[1060]), .P2_P3_LWORD_REG_3_(vec[1059]), .P2_P3_LWORD_REG_2_(vec[1058]), .P2_P3_LWORD_REG_1_(vec[1057]), .P2_P3_LWORD_REG_0_(vec[1056]), .P2_P3_UWORD_REG_14_(vec[1055]), .P2_P3_UWORD_REG_13_(vec[1054]), .P2_P3_UWORD_REG_12_(vec[1053]), .P2_P3_UWORD_REG_11_(vec[1052]), .P2_P3_UWORD_REG_10_(vec[1051]), .P2_P3_UWORD_REG_9_(vec[1050]), .P2_P3_UWORD_REG_8_(vec[1049]), .P2_P3_UWORD_REG_7_(vec[1048]), .P2_P3_UWORD_REG_6_(vec[1047]), .P2_P3_UWORD_REG_5_(vec[1046]), .P2_P3_UWORD_REG_4_(vec[1045]), .P2_P3_UWORD_REG_3_(vec[1044]), .P2_P3_UWORD_REG_2_(vec[1043]), .P2_P3_UWORD_REG_1_(vec[1042]), .P2_P3_UWORD_REG_0_(vec[1041]), .P2_P3_DATAO_REG_0_(vec[1040]), .P2_P3_DATAO_REG_1_(vec[1039]), .P2_P3_DATAO_REG_2_(vec[1038]), .P2_P3_DATAO_REG_3_(vec[1037]), .P2_P3_DATAO_REG_4_(vec[1036]), .P2_P3_DATAO_REG_5_(vec[1035]), .P2_P3_DATAO_REG_6_(vec[1034]), .P2_P3_DATAO_REG_7_(vec[1033]), .P2_P3_DATAO_REG_8_(vec[1032]), .P2_P3_DATAO_REG_9_(vec[1031]), .P2_P3_DATAO_REG_10_(vec[1030]), .P2_P3_DATAO_REG_11_(vec[1029]), .P2_P3_DATAO_REG_12_(vec[1028]), .P2_P3_DATAO_REG_13_(vec[1027]), .P2_P3_DATAO_REG_14_(vec[1026]), .P2_P3_DATAO_REG_15_(vec[1025]), .P2_P3_DATAO_REG_16_(vec[1024]), .P2_P3_DATAO_REG_17_(vec[1023]), .P2_P3_DATAO_REG_18_(vec[1022]), .P2_P3_DATAO_REG_19_(vec[1021]), .P2_P3_DATAO_REG_20_(vec[1020]), .P2_P3_DATAO_REG_21_(vec[1019]), .P2_P3_DATAO_REG_22_(vec[1018]), .P2_P3_DATAO_REG_23_(vec[1017]), .P2_P3_DATAO_REG_24_(vec[1016]), .P2_P3_DATAO_REG_25_(vec[1015]), .P2_P3_DATAO_REG_26_(vec[1014]), .P2_P3_DATAO_REG_27_(vec[1013]), .P2_P3_DATAO_REG_28_(vec[1012]), .P2_P3_DATAO_REG_29_(vec[1011]), .P2_P3_DATAO_REG_30_(vec[1010]), .P2_P3_DATAO_REG_31_(vec[1009]), .P2_P3_EAX_REG_0_(vec[1008]), .P2_P3_EAX_REG_1_(vec[1007]), .P2_P3_EAX_REG_2_(vec[1006]), .P2_P3_EAX_REG_3_(vec[1005]), .P2_P3_EAX_REG_4_(vec[1004]), .P2_P3_EAX_REG_5_(vec[1003]), .P2_P3_EAX_REG_6_(vec[1002]), .P2_P3_EAX_REG_7_(vec[1001]), .P2_P3_EAX_REG_8_(vec[1000]), .P2_P3_EAX_REG_9_(vec[999]), .P2_P3_EAX_REG_10_(vec[998]), .P2_P3_EAX_REG_11_(vec[997]), .P2_P3_EAX_REG_12_(vec[996]), .P2_P3_EAX_REG_13_(vec[995]), .P2_P3_EAX_REG_14_(vec[994]), .P2_P3_EAX_REG_15_(vec[993]), .P2_P3_EAX_REG_16_(vec[992]), .P2_P3_EAX_REG_17_(vec[991]), .P2_P3_EAX_REG_18_(vec[990]), .P2_P3_EAX_REG_19_(vec[989]), .P2_P3_EAX_REG_20_(vec[988]), .P2_P3_EAX_REG_21_(vec[987]), .P2_P3_EAX_REG_22_(vec[986]), .P2_P3_EAX_REG_23_(vec[985]), .P2_P3_EAX_REG_24_(vec[984]), .P2_P3_EAX_REG_25_(vec[983]), .P2_P3_EAX_REG_26_(vec[982]), .P2_P3_EAX_REG_27_(vec[981]), .P2_P3_EAX_REG_28_(vec[980]), .P2_P3_EAX_REG_29_(vec[979]), .P2_P3_EAX_REG_30_(vec[978]), .P2_P3_EAX_REG_31_(vec[977]), .P2_P3_EBX_REG_0_(vec[976]), .P2_P3_EBX_REG_1_(vec[975]), .P2_P3_EBX_REG_2_(vec[974]), .P2_P3_EBX_REG_3_(vec[973]), .P2_P3_EBX_REG_4_(vec[972]), .P2_P3_EBX_REG_5_(vec[971]), .P2_P3_EBX_REG_6_(vec[970]), .P2_P3_EBX_REG_7_(vec[969]), .P2_P3_EBX_REG_8_(vec[968]), .P2_P3_EBX_REG_9_(vec[967]), .P2_P3_EBX_REG_10_(vec[966]), .P2_P3_EBX_REG_11_(vec[965]), .P2_P3_EBX_REG_12_(vec[964]), .P2_P3_EBX_REG_13_(vec[963]), .P2_P3_EBX_REG_14_(vec[962]), .P2_P3_EBX_REG_15_(vec[961]), .P2_P3_EBX_REG_16_(vec[960]), .P2_P3_EBX_REG_17_(vec[959]), .P2_P3_EBX_REG_18_(vec[958]), .P2_P3_EBX_REG_19_(vec[957]), .P2_P3_EBX_REG_20_(vec[956]), .P2_P3_EBX_REG_21_(vec[955]), .P2_P3_EBX_REG_22_(vec[954]), .P2_P3_EBX_REG_23_(vec[953]), .P2_P3_EBX_REG_24_(vec[952]), .P2_P3_EBX_REG_25_(vec[951]), .P2_P3_EBX_REG_26_(vec[950]), .P2_P3_EBX_REG_27_(vec[949]), .P2_P3_EBX_REG_28_(vec[948]), .P2_P3_EBX_REG_29_(vec[947]), .P2_P3_EBX_REG_30_(vec[946]), .P2_P3_EBX_REG_31_(vec[945]), .P2_P3_REIP_REG_0_(vec[944]), .P2_P3_REIP_REG_1_(vec[943]), .P2_P3_REIP_REG_2_(vec[942]), .P2_P3_REIP_REG_3_(vec[941]), .P2_P3_REIP_REG_4_(vec[940]), .P2_P3_REIP_REG_5_(vec[939]), .P2_P3_REIP_REG_6_(vec[938]), .P2_P3_REIP_REG_7_(vec[937]), .P2_P3_REIP_REG_8_(vec[936]), .P2_P3_REIP_REG_9_(vec[935]), .P2_P3_REIP_REG_10_(vec[934]), .P2_P3_REIP_REG_11_(vec[933]), .P2_P3_REIP_REG_12_(vec[932]), .P2_P3_REIP_REG_13_(vec[931]), .P2_P3_REIP_REG_14_(vec[930]), .P2_P3_REIP_REG_15_(vec[929]), .P2_P3_REIP_REG_16_(vec[928]), .P2_P3_REIP_REG_17_(vec[927]), .P2_P3_REIP_REG_18_(vec[926]), .P2_P3_REIP_REG_19_(vec[925]), .P2_P3_REIP_REG_20_(vec[924]), .P2_P3_REIP_REG_21_(vec[923]), .P2_P3_REIP_REG_22_(vec[922]), .P2_P3_REIP_REG_23_(vec[921]), .P2_P3_REIP_REG_24_(vec[920]), .P2_P3_REIP_REG_25_(vec[919]), .P2_P3_REIP_REG_26_(vec[918]), .P2_P3_REIP_REG_27_(vec[917]), .P2_P3_REIP_REG_28_(vec[916]), .P2_P3_REIP_REG_29_(vec[915]), .P2_P3_REIP_REG_30_(vec[914]), .P2_P3_REIP_REG_31_(vec[913]), .P2_P3_BYTEENABLE_REG_3_(vec[912]), .P2_P3_BYTEENABLE_REG_2_(vec[911]), .P2_P3_BYTEENABLE_REG_1_(vec[910]), .P2_P3_BYTEENABLE_REG_0_(vec[909]), .P2_P3_W_R_N_REG(vec[908]), .P2_P3_FLUSH_REG(vec[907]), .P2_P3_MORE_REG(vec[906]), .P2_P3_STATEBS16_REG(vec[905]), .P2_P3_REQUESTPENDING_REG(vec[904]), .P2_P3_D_C_N_REG(vec[903]), .P2_P3_M_IO_N_REG(vec[902]), .P2_P3_CODEFETCH_REG(vec[901]), .P2_P3_ADS_N_REG(vec[900]), .P2_P3_READREQUEST_REG(vec[899]), .P2_P3_MEMORYFETCH_REG(vec[898]), .P2_P2_BE_N_REG_3_(vec[897]), .P2_P2_BE_N_REG_2_(vec[896]), .P2_P2_BE_N_REG_1_(vec[895]), .P2_P2_BE_N_REG_0_(vec[894]), .P2_P2_ADDRESS_REG_29_(vec[893]), .P2_P2_ADDRESS_REG_28_(vec[892]), .P2_P2_ADDRESS_REG_27_(vec[891]), .P2_P2_ADDRESS_REG_26_(vec[890]), .P2_P2_ADDRESS_REG_25_(vec[889]), .P2_P2_ADDRESS_REG_24_(vec[888]), .P2_P2_ADDRESS_REG_23_(vec[887]), .P2_P2_ADDRESS_REG_22_(vec[886]), .P2_P2_ADDRESS_REG_21_(vec[885]), .P2_P2_ADDRESS_REG_20_(vec[884]), .P2_P2_ADDRESS_REG_19_(vec[883]), .P2_P2_ADDRESS_REG_18_(vec[882]), .P2_P2_ADDRESS_REG_17_(vec[881]), .P2_P2_ADDRESS_REG_16_(vec[880]), .P2_P2_ADDRESS_REG_15_(vec[879]), .P2_P2_ADDRESS_REG_14_(vec[878]), .P2_P2_ADDRESS_REG_13_(vec[877]), .P2_P2_ADDRESS_REG_12_(vec[876]), .P2_P2_ADDRESS_REG_11_(vec[875]), .P2_P2_ADDRESS_REG_10_(vec[874]), .P2_P2_ADDRESS_REG_9_(vec[873]), .P2_P2_ADDRESS_REG_8_(vec[872]), .P2_P2_ADDRESS_REG_7_(vec[871]), .P2_P2_ADDRESS_REG_6_(vec[870]), .P2_P2_ADDRESS_REG_5_(vec[869]), .P2_P2_ADDRESS_REG_4_(vec[868]), .P2_P2_ADDRESS_REG_3_(vec[867]), .P2_P2_ADDRESS_REG_2_(vec[866]), .P2_P2_ADDRESS_REG_1_(vec[865]), .P2_P2_ADDRESS_REG_0_(vec[864]), .P2_P2_STATE_REG_2_(vec[863]), .P2_P2_STATE_REG_1_(vec[862]), .P2_P2_STATE_REG_0_(vec[861]), .P2_P2_DATAWIDTH_REG_0_(vec[860]), .P2_P2_DATAWIDTH_REG_1_(vec[859]), .P2_P2_DATAWIDTH_REG_2_(vec[858]), .P2_P2_DATAWIDTH_REG_3_(vec[857]), .P2_P2_DATAWIDTH_REG_4_(vec[856]), .P2_P2_DATAWIDTH_REG_5_(vec[855]), .P2_P2_DATAWIDTH_REG_6_(vec[854]), .P2_P2_DATAWIDTH_REG_7_(vec[853]), .P2_P2_DATAWIDTH_REG_8_(vec[852]), .P2_P2_DATAWIDTH_REG_9_(vec[851]), .P2_P2_DATAWIDTH_REG_10_(vec[850]), .P2_P2_DATAWIDTH_REG_11_(vec[849]), .P2_P2_DATAWIDTH_REG_12_(vec[848]), .P2_P2_DATAWIDTH_REG_13_(vec[847]), .P2_P2_DATAWIDTH_REG_14_(vec[846]), .P2_P2_DATAWIDTH_REG_15_(vec[845]), .P2_P2_DATAWIDTH_REG_16_(vec[844]), .P2_P2_DATAWIDTH_REG_17_(vec[843]), .P2_P2_DATAWIDTH_REG_18_(vec[842]), .P2_P2_DATAWIDTH_REG_19_(vec[841]), .P2_P2_DATAWIDTH_REG_20_(vec[840]), .P2_P2_DATAWIDTH_REG_21_(vec[839]), .P2_P2_DATAWIDTH_REG_22_(vec[838]), .P2_P2_DATAWIDTH_REG_23_(vec[837]), .P2_P2_DATAWIDTH_REG_24_(vec[836]), .P2_P2_DATAWIDTH_REG_25_(vec[835]), .P2_P2_DATAWIDTH_REG_26_(vec[834]), .P2_P2_DATAWIDTH_REG_27_(vec[833]), .P2_P2_DATAWIDTH_REG_28_(vec[832]), .P2_P2_DATAWIDTH_REG_29_(vec[831]), .P2_P2_DATAWIDTH_REG_30_(vec[830]), .P2_P2_DATAWIDTH_REG_31_(vec[829]), .P2_P2_STATE2_REG_3_(vec[828]), .P2_P2_STATE2_REG_2_(vec[827]), .P2_P2_STATE2_REG_1_(vec[826]), .P2_P2_STATE2_REG_0_(vec[825]), .P2_P2_INSTQUEUE_REG_15__7_(vec[824]), .P2_P2_INSTQUEUE_REG_15__6_(vec[823]), .P2_P2_INSTQUEUE_REG_15__5_(vec[822]), .P2_P2_INSTQUEUE_REG_15__4_(vec[821]), .P2_P2_INSTQUEUE_REG_15__3_(vec[820]), .P2_P2_INSTQUEUE_REG_15__2_(vec[819]), .P2_P2_INSTQUEUE_REG_15__1_(vec[818]), .P2_P2_INSTQUEUE_REG_15__0_(vec[817]), .P2_P2_INSTQUEUE_REG_14__7_(vec[816]), .P2_P2_INSTQUEUE_REG_14__6_(vec[815]), .P2_P2_INSTQUEUE_REG_14__5_(vec[814]), .P2_P2_INSTQUEUE_REG_14__4_(vec[813]), .P2_P2_INSTQUEUE_REG_14__3_(vec[812]), .P2_P2_INSTQUEUE_REG_14__2_(vec[811]), .P2_P2_INSTQUEUE_REG_14__1_(vec[810]), .P2_P2_INSTQUEUE_REG_14__0_(vec[809]), .P2_P2_INSTQUEUE_REG_13__7_(vec[808]), .P2_P2_INSTQUEUE_REG_13__6_(vec[807]), .P2_P2_INSTQUEUE_REG_13__5_(vec[806]), .P2_P2_INSTQUEUE_REG_13__4_(vec[805]), .P2_P2_INSTQUEUE_REG_13__3_(vec[804]), .P2_P2_INSTQUEUE_REG_13__2_(vec[803]), .P2_P2_INSTQUEUE_REG_13__1_(vec[802]), .P2_P2_INSTQUEUE_REG_13__0_(vec[801]), .P2_P2_INSTQUEUE_REG_12__7_(vec[800]), .P2_P2_INSTQUEUE_REG_12__6_(vec[799]), .P2_P2_INSTQUEUE_REG_12__5_(vec[798]), .P2_P2_INSTQUEUE_REG_12__4_(vec[797]), .P2_P2_INSTQUEUE_REG_12__3_(vec[796]), .P2_P2_INSTQUEUE_REG_12__2_(vec[795]), .P2_P2_INSTQUEUE_REG_12__1_(vec[794]), .P2_P2_INSTQUEUE_REG_12__0_(vec[793]), .P2_P2_INSTQUEUE_REG_11__7_(vec[792]), .P2_P2_INSTQUEUE_REG_11__6_(vec[791]), .P2_P2_INSTQUEUE_REG_11__5_(vec[790]), .P2_P2_INSTQUEUE_REG_11__4_(vec[789]), .P2_P2_INSTQUEUE_REG_11__3_(vec[788]), .P2_P2_INSTQUEUE_REG_11__2_(vec[787]), .P2_P2_INSTQUEUE_REG_11__1_(vec[786]), .P2_P2_INSTQUEUE_REG_11__0_(vec[785]), .P2_P2_INSTQUEUE_REG_10__7_(vec[784]), .P2_P2_INSTQUEUE_REG_10__6_(vec[783]), .P2_P2_INSTQUEUE_REG_10__5_(vec[782]), .P2_P2_INSTQUEUE_REG_10__4_(vec[781]), .P2_P2_INSTQUEUE_REG_10__3_(vec[780]), .P2_P2_INSTQUEUE_REG_10__2_(vec[779]), .P2_P2_INSTQUEUE_REG_10__1_(vec[778]), .P2_P2_INSTQUEUE_REG_10__0_(vec[777]), .P2_P2_INSTQUEUE_REG_9__7_(vec[776]), .P2_P2_INSTQUEUE_REG_9__6_(vec[775]), .P2_P2_INSTQUEUE_REG_9__5_(vec[774]), .P2_P2_INSTQUEUE_REG_9__4_(vec[773]), .P2_P2_INSTQUEUE_REG_9__3_(vec[772]), .P2_P2_INSTQUEUE_REG_9__2_(vec[771]), .P2_P2_INSTQUEUE_REG_9__1_(vec[770]), .P2_P2_INSTQUEUE_REG_9__0_(vec[769]), .P2_P2_INSTQUEUE_REG_8__7_(vec[768]), .P2_P2_INSTQUEUE_REG_8__6_(vec[767]), .P2_P2_INSTQUEUE_REG_8__5_(vec[766]), .P2_P2_INSTQUEUE_REG_8__4_(vec[765]), .P2_P2_INSTQUEUE_REG_8__3_(vec[764]), .P2_P2_INSTQUEUE_REG_8__2_(vec[763]), .P2_P2_INSTQUEUE_REG_8__1_(vec[762]), .P2_P2_INSTQUEUE_REG_8__0_(vec[761]), .P2_P2_INSTQUEUE_REG_7__7_(vec[760]), .P2_P2_INSTQUEUE_REG_7__6_(vec[759]), .P2_P2_INSTQUEUE_REG_7__5_(vec[758]), .P2_P2_INSTQUEUE_REG_7__4_(vec[757]), .P2_P2_INSTQUEUE_REG_7__3_(vec[756]), .P2_P2_INSTQUEUE_REG_7__2_(vec[755]), .P2_P2_INSTQUEUE_REG_7__1_(vec[754]), .P2_P2_INSTQUEUE_REG_7__0_(vec[753]), .P2_P2_INSTQUEUE_REG_6__7_(vec[752]), .P2_P2_INSTQUEUE_REG_6__6_(vec[751]), .P2_P2_INSTQUEUE_REG_6__5_(vec[750]), .P2_P2_INSTQUEUE_REG_6__4_(vec[749]), .P2_P2_INSTQUEUE_REG_6__3_(vec[748]), .P2_P2_INSTQUEUE_REG_6__2_(vec[747]), .P2_P2_INSTQUEUE_REG_6__1_(vec[746]), .P2_P2_INSTQUEUE_REG_6__0_(vec[745]), .P2_P2_INSTQUEUE_REG_5__7_(vec[744]), .P2_P2_INSTQUEUE_REG_5__6_(vec[743]), .P2_P2_INSTQUEUE_REG_5__5_(vec[742]), .P2_P2_INSTQUEUE_REG_5__4_(vec[741]), .P2_P2_INSTQUEUE_REG_5__3_(vec[740]), .P2_P2_INSTQUEUE_REG_5__2_(vec[739]), .P2_P2_INSTQUEUE_REG_5__1_(vec[738]), .P2_P2_INSTQUEUE_REG_5__0_(vec[737]), .P2_P2_INSTQUEUE_REG_4__7_(vec[736]), .P2_P2_INSTQUEUE_REG_4__6_(vec[735]), .P2_P2_INSTQUEUE_REG_4__5_(vec[734]), .P2_P2_INSTQUEUE_REG_4__4_(vec[733]), .P2_P2_INSTQUEUE_REG_4__3_(vec[732]), .P2_P2_INSTQUEUE_REG_4__2_(vec[731]), .P2_P2_INSTQUEUE_REG_4__1_(vec[730]), .P2_P2_INSTQUEUE_REG_4__0_(vec[729]), .P2_P2_INSTQUEUE_REG_3__7_(vec[728]), .P2_P2_INSTQUEUE_REG_3__6_(vec[727]), .P2_P2_INSTQUEUE_REG_3__5_(vec[726]), .P2_P2_INSTQUEUE_REG_3__4_(vec[725]), .P2_P2_INSTQUEUE_REG_3__3_(vec[724]), .P2_P2_INSTQUEUE_REG_3__2_(vec[723]), .P2_P2_INSTQUEUE_REG_3__1_(vec[722]), .P2_P2_INSTQUEUE_REG_3__0_(vec[721]), .P2_P2_INSTQUEUE_REG_2__7_(vec[720]), .P2_P2_INSTQUEUE_REG_2__6_(vec[719]), .P2_P2_INSTQUEUE_REG_2__5_(vec[718]), .P2_P2_INSTQUEUE_REG_2__4_(vec[717]), .P2_P2_INSTQUEUE_REG_2__3_(vec[716]), .P2_P2_INSTQUEUE_REG_2__2_(vec[715]), .P2_P2_INSTQUEUE_REG_2__1_(vec[714]), .P2_P2_INSTQUEUE_REG_2__0_(vec[713]), .P2_P2_INSTQUEUE_REG_1__7_(vec[712]), .P2_P2_INSTQUEUE_REG_1__6_(vec[711]), .P2_P2_INSTQUEUE_REG_1__5_(vec[710]), .P2_P2_INSTQUEUE_REG_1__4_(vec[709]), .P2_P2_INSTQUEUE_REG_1__3_(vec[708]), .P2_P2_INSTQUEUE_REG_1__2_(vec[707]), .P2_P2_INSTQUEUE_REG_1__1_(vec[706]), .P2_P2_INSTQUEUE_REG_1__0_(vec[705]), .P2_P2_INSTQUEUE_REG_0__7_(vec[704]), .P2_P2_INSTQUEUE_REG_0__6_(vec[703]), .P2_P2_INSTQUEUE_REG_0__5_(vec[702]), .P2_P2_INSTQUEUE_REG_0__4_(vec[701]), .P2_P2_INSTQUEUE_REG_0__3_(vec[700]), .P2_P2_INSTQUEUE_REG_0__2_(vec[699]), .P2_P2_INSTQUEUE_REG_0__1_(vec[698]), .P2_P2_INSTQUEUE_REG_0__0_(vec[697]), .P2_P2_INSTQUEUERD_ADDR_REG_4_(vec[696]), .P2_P2_INSTQUEUERD_ADDR_REG_3_(vec[695]), .P2_P2_INSTQUEUERD_ADDR_REG_2_(vec[694]), .P2_P2_INSTQUEUERD_ADDR_REG_1_(vec[693]), .P2_P2_INSTQUEUERD_ADDR_REG_0_(vec[692]), .P2_P2_INSTQUEUEWR_ADDR_REG_4_(vec[691]), .P2_P2_INSTQUEUEWR_ADDR_REG_3_(vec[690]), .P2_P2_INSTQUEUEWR_ADDR_REG_2_(vec[689]), .P2_P2_INSTQUEUEWR_ADDR_REG_1_(vec[688]), .P2_P2_INSTQUEUEWR_ADDR_REG_0_(vec[687]), .P2_P2_INSTADDRPOINTER_REG_0_(vec[686]), .P2_P2_INSTADDRPOINTER_REG_1_(vec[685]), .P2_P2_INSTADDRPOINTER_REG_2_(vec[684]), .P2_P2_INSTADDRPOINTER_REG_3_(vec[683]), .P2_P2_INSTADDRPOINTER_REG_4_(vec[682]), .P2_P2_INSTADDRPOINTER_REG_5_(vec[681]), .P2_P2_INSTADDRPOINTER_REG_6_(vec[680]), .P2_P2_INSTADDRPOINTER_REG_7_(vec[679]), .P2_P2_INSTADDRPOINTER_REG_8_(vec[678]), .P2_P2_INSTADDRPOINTER_REG_9_(vec[677]), .P2_P2_INSTADDRPOINTER_REG_10_(vec[676]), .P2_P2_INSTADDRPOINTER_REG_11_(vec[675]), .P2_P2_INSTADDRPOINTER_REG_12_(vec[674]), .P2_P2_INSTADDRPOINTER_REG_13_(vec[673]), .P2_P2_INSTADDRPOINTER_REG_14_(vec[672]), .P2_P2_INSTADDRPOINTER_REG_15_(vec[671]), .P2_P2_INSTADDRPOINTER_REG_16_(vec[670]), .P2_P2_INSTADDRPOINTER_REG_17_(vec[669]), .P2_P2_INSTADDRPOINTER_REG_18_(vec[668]), .P2_P2_INSTADDRPOINTER_REG_19_(vec[667]), .P2_P2_INSTADDRPOINTER_REG_20_(vec[666]), .P2_P2_INSTADDRPOINTER_REG_21_(vec[665]), .P2_P2_INSTADDRPOINTER_REG_22_(vec[664]), .P2_P2_INSTADDRPOINTER_REG_23_(vec[663]), .P2_P2_INSTADDRPOINTER_REG_24_(vec[662]), .P2_P2_INSTADDRPOINTER_REG_25_(vec[661]), .P2_P2_INSTADDRPOINTER_REG_26_(vec[660]), .P2_P2_INSTADDRPOINTER_REG_27_(vec[659]), .P2_P2_INSTADDRPOINTER_REG_28_(vec[658]), .P2_P2_INSTADDRPOINTER_REG_29_(vec[657]), .P2_P2_INSTADDRPOINTER_REG_30_(vec[656]), .P2_P2_INSTADDRPOINTER_REG_31_(vec[655]), .P2_P2_PHYADDRPOINTER_REG_0_(vec[654]), .P2_P2_PHYADDRPOINTER_REG_1_(vec[653]), .P2_P2_PHYADDRPOINTER_REG_2_(vec[652]), .P2_P2_PHYADDRPOINTER_REG_3_(vec[651]), .P2_P2_PHYADDRPOINTER_REG_4_(vec[650]), .P2_P2_PHYADDRPOINTER_REG_5_(vec[649]), .P2_P2_PHYADDRPOINTER_REG_6_(vec[648]), .P2_P2_PHYADDRPOINTER_REG_7_(vec[647]), .P2_P2_PHYADDRPOINTER_REG_8_(vec[646]), .P2_P2_PHYADDRPOINTER_REG_9_(vec[645]), .P2_P2_PHYADDRPOINTER_REG_10_(vec[644]), .P2_P2_PHYADDRPOINTER_REG_11_(vec[643]), .P2_P2_PHYADDRPOINTER_REG_12_(vec[642]), .P2_P2_PHYADDRPOINTER_REG_13_(vec[641]), .P2_P2_PHYADDRPOINTER_REG_14_(vec[640]), .P2_P2_PHYADDRPOINTER_REG_15_(vec[639]), .P2_P2_PHYADDRPOINTER_REG_16_(vec[638]), .P2_P2_PHYADDRPOINTER_REG_17_(vec[637]), .P2_P2_PHYADDRPOINTER_REG_18_(vec[636]), .P2_P2_PHYADDRPOINTER_REG_19_(vec[635]), .P2_P2_PHYADDRPOINTER_REG_20_(vec[634]), .P2_P2_PHYADDRPOINTER_REG_21_(vec[633]), .P2_P2_PHYADDRPOINTER_REG_22_(vec[632]), .P2_P2_PHYADDRPOINTER_REG_23_(vec[631]), .P2_P2_PHYADDRPOINTER_REG_24_(vec[630]), .P2_P2_PHYADDRPOINTER_REG_25_(vec[629]), .P2_P2_PHYADDRPOINTER_REG_26_(vec[628]), .P2_P2_PHYADDRPOINTER_REG_27_(vec[627]), .P2_P2_PHYADDRPOINTER_REG_28_(vec[626]), .P2_P2_PHYADDRPOINTER_REG_29_(vec[625]), .P2_P2_PHYADDRPOINTER_REG_30_(vec[624]), .P2_P2_PHYADDRPOINTER_REG_31_(vec[623]), .P2_P2_LWORD_REG_15_(vec[622]), .P2_P2_LWORD_REG_14_(vec[621]), .P2_P2_LWORD_REG_13_(vec[620]), .P2_P2_LWORD_REG_12_(vec[619]), .P2_P2_LWORD_REG_11_(vec[618]), .P2_P2_LWORD_REG_10_(vec[617]), .P2_P2_LWORD_REG_9_(vec[616]), .P2_P2_LWORD_REG_8_(vec[615]), .P2_P2_LWORD_REG_7_(vec[614]), .P2_P2_LWORD_REG_6_(vec[613]), .P2_P2_LWORD_REG_5_(vec[612]), .P2_P2_LWORD_REG_4_(vec[611]), .P2_P2_LWORD_REG_3_(vec[610]), .P2_P2_LWORD_REG_2_(vec[609]), .P2_P2_LWORD_REG_1_(vec[608]), .P2_P2_LWORD_REG_0_(vec[607]), .P2_P2_UWORD_REG_14_(vec[606]), .P2_P2_UWORD_REG_13_(vec[605]), .P2_P2_UWORD_REG_12_(vec[604]), .P2_P2_UWORD_REG_11_(vec[603]), .P2_P2_UWORD_REG_10_(vec[602]), .P2_P2_UWORD_REG_9_(vec[601]), .P2_P2_UWORD_REG_8_(vec[600]), .P2_P2_UWORD_REG_7_(vec[599]), .P2_P2_UWORD_REG_6_(vec[598]), .P2_P2_UWORD_REG_5_(vec[597]), .P2_P2_UWORD_REG_4_(vec[596]), .P2_P2_UWORD_REG_3_(vec[595]), .P2_P2_UWORD_REG_2_(vec[594]), .P2_P2_UWORD_REG_1_(vec[593]), .P2_P2_UWORD_REG_0_(vec[592]), .P2_P2_DATAO_REG_0_(vec[591]), .P2_P2_DATAO_REG_1_(vec[590]), .P2_P2_DATAO_REG_2_(vec[589]), .P2_P2_DATAO_REG_3_(vec[588]), .P2_P2_DATAO_REG_4_(vec[587]), .P2_P2_DATAO_REG_5_(vec[586]), .P2_P2_DATAO_REG_6_(vec[585]), .P2_P2_DATAO_REG_7_(vec[584]), .P2_P2_DATAO_REG_8_(vec[583]), .P2_P2_DATAO_REG_9_(vec[582]), .P2_P2_DATAO_REG_10_(vec[581]), .P2_P2_DATAO_REG_11_(vec[580]), .P2_P2_DATAO_REG_12_(vec[579]), .P2_P2_DATAO_REG_13_(vec[578]), .P2_P2_DATAO_REG_14_(vec[577]), .P2_P2_DATAO_REG_15_(vec[576]), .P2_P2_DATAO_REG_16_(vec[575]), .P2_P2_DATAO_REG_17_(vec[574]), .P2_P2_DATAO_REG_18_(vec[573]), .P2_P2_DATAO_REG_19_(vec[572]), .P2_P2_DATAO_REG_20_(vec[571]), .P2_P2_DATAO_REG_21_(vec[570]), .P2_P2_DATAO_REG_22_(vec[569]), .P2_P2_DATAO_REG_23_(vec[568]), .P2_P2_DATAO_REG_24_(vec[567]), .P2_P2_DATAO_REG_25_(vec[566]), .P2_P2_DATAO_REG_26_(vec[565]), .P2_P2_DATAO_REG_27_(vec[564]), .P2_P2_DATAO_REG_28_(vec[563]), .P2_P2_DATAO_REG_29_(vec[562]), .P2_P2_DATAO_REG_30_(vec[561]), .P2_P2_DATAO_REG_31_(vec[560]), .P2_P2_EAX_REG_0_(vec[559]), .P2_P2_EAX_REG_1_(vec[558]), .P2_P2_EAX_REG_2_(vec[557]), .P2_P2_EAX_REG_3_(vec[556]), .P2_P2_EAX_REG_4_(vec[555]), .P2_P2_EAX_REG_5_(vec[554]), .P2_P2_EAX_REG_6_(vec[553]), .P2_P2_EAX_REG_7_(vec[552]), .P2_P2_EAX_REG_8_(vec[551]), .P2_P2_EAX_REG_9_(vec[550]), .P2_P2_EAX_REG_10_(vec[549]), .P2_P2_EAX_REG_11_(vec[548]), .P2_P2_EAX_REG_12_(vec[547]), .P2_P2_EAX_REG_13_(vec[546]), .P2_P2_EAX_REG_14_(vec[545]), .P2_P2_EAX_REG_15_(vec[544]), .P2_P2_EAX_REG_16_(vec[543]), .P2_P2_EAX_REG_17_(vec[542]), .P2_P2_EAX_REG_18_(vec[541]), .P2_P2_EAX_REG_19_(vec[540]), .P2_P2_EAX_REG_20_(vec[539]), .P2_P2_EAX_REG_21_(vec[538]), .P2_P2_EAX_REG_22_(vec[537]), .P2_P2_EAX_REG_23_(vec[536]), .P2_P2_EAX_REG_24_(vec[535]), .P2_P2_EAX_REG_25_(vec[534]), .P2_P2_EAX_REG_26_(vec[533]), .P2_P2_EAX_REG_27_(vec[532]), .P2_P2_EAX_REG_28_(vec[531]), .P2_P2_EAX_REG_29_(vec[530]), .P2_P2_EAX_REG_30_(vec[529]), .P2_P2_EAX_REG_31_(vec[528]), .P2_P2_EBX_REG_0_(vec[527]), .P2_P2_EBX_REG_1_(vec[526]), .P2_P2_EBX_REG_2_(vec[525]), .P2_P2_EBX_REG_3_(vec[524]), .P2_P2_EBX_REG_4_(vec[523]), .P2_P2_EBX_REG_5_(vec[522]), .P2_P2_EBX_REG_6_(vec[521]), .P2_P2_EBX_REG_7_(vec[520]), .P2_P2_EBX_REG_8_(vec[519]), .P2_P2_EBX_REG_9_(vec[518]), .P2_P2_EBX_REG_10_(vec[517]), .P2_P2_EBX_REG_11_(vec[516]), .P2_P2_EBX_REG_12_(vec[515]), .P2_P2_EBX_REG_13_(vec[514]), .P2_P2_EBX_REG_14_(vec[513]), .P2_P2_EBX_REG_15_(vec[512]), .P2_P2_EBX_REG_16_(vec[511]), .P2_P2_EBX_REG_17_(vec[510]), .P2_P2_EBX_REG_18_(vec[509]), .P2_P2_EBX_REG_19_(vec[508]), .P2_P2_EBX_REG_20_(vec[507]), .P2_P2_EBX_REG_21_(vec[506]), .P2_P2_EBX_REG_22_(vec[505]), .P2_P2_EBX_REG_23_(vec[504]), .P2_P2_EBX_REG_24_(vec[503]), .P2_P2_EBX_REG_25_(vec[502]), .P2_P2_EBX_REG_26_(vec[501]), .P2_P2_EBX_REG_27_(vec[500]), .P2_P2_EBX_REG_28_(vec[499]), .P2_P2_EBX_REG_29_(vec[498]), .P2_P2_EBX_REG_30_(vec[497]), .P2_P2_EBX_REG_31_(vec[496]), .P2_P2_REIP_REG_0_(vec[495]), .P2_P2_REIP_REG_1_(vec[494]), .P2_P2_REIP_REG_2_(vec[493]), .P2_P2_REIP_REG_3_(vec[492]), .P2_P2_REIP_REG_4_(vec[491]), .P2_P2_REIP_REG_5_(vec[490]), .P2_P2_REIP_REG_6_(vec[489]), .P2_P2_REIP_REG_7_(vec[488]), .P2_P2_REIP_REG_8_(vec[487]), .P2_P2_REIP_REG_9_(vec[486]), .P2_P2_REIP_REG_10_(vec[485]), .P2_P2_REIP_REG_11_(vec[484]), .P2_P2_REIP_REG_12_(vec[483]), .P2_P2_REIP_REG_13_(vec[482]), .P2_P2_REIP_REG_14_(vec[481]), .P2_P2_REIP_REG_15_(vec[480]), .P2_P2_REIP_REG_16_(vec[479]), .P2_P2_REIP_REG_17_(vec[478]), .P2_P2_REIP_REG_18_(vec[477]), .P2_P2_REIP_REG_19_(vec[476]), .P2_P2_REIP_REG_20_(vec[475]), .P2_P2_REIP_REG_21_(vec[474]), .P2_P2_REIP_REG_22_(vec[473]), .P2_P2_REIP_REG_23_(vec[472]), .P2_P2_REIP_REG_24_(vec[471]), .P2_P2_REIP_REG_25_(vec[470]), .P2_P2_REIP_REG_26_(vec[469]), .P2_P2_REIP_REG_27_(vec[468]), .P2_P2_REIP_REG_28_(vec[467]), .P2_P2_REIP_REG_29_(vec[466]), .P2_P2_REIP_REG_30_(vec[465]), .P2_P2_REIP_REG_31_(vec[464]), .P2_P2_BYTEENABLE_REG_3_(vec[463]), .P2_P2_BYTEENABLE_REG_2_(vec[462]), .P2_P2_BYTEENABLE_REG_1_(vec[461]), .P2_P2_BYTEENABLE_REG_0_(vec[460]), .P2_P2_W_R_N_REG(vec[459]), .P2_P2_FLUSH_REG(vec[458]), .P2_P2_MORE_REG(vec[457]), .P2_P2_STATEBS16_REG(vec[456]), .P2_P2_REQUESTPENDING_REG(vec[455]), .P2_P2_D_C_N_REG(vec[454]), .P2_P2_M_IO_N_REG(vec[453]), .P2_P2_CODEFETCH_REG(vec[452]), .P2_P2_ADS_N_REG(vec[451]), .P2_P2_READREQUEST_REG(vec[450]), .P2_P2_MEMORYFETCH_REG(vec[449]), .P2_P1_BE_N_REG_3_(vec[448]), .P2_P1_BE_N_REG_2_(vec[447]), .P2_P1_BE_N_REG_1_(vec[446]), .P2_P1_BE_N_REG_0_(vec[445]), .P2_P1_ADDRESS_REG_29_(vec[444]), .P2_P1_ADDRESS_REG_28_(vec[443]), .P2_P1_ADDRESS_REG_27_(vec[442]), .P2_P1_ADDRESS_REG_26_(vec[441]), .P2_P1_ADDRESS_REG_25_(vec[440]), .P2_P1_ADDRESS_REG_24_(vec[439]), .P2_P1_ADDRESS_REG_23_(vec[438]), .P2_P1_ADDRESS_REG_22_(vec[437]), .P2_P1_ADDRESS_REG_21_(vec[436]), .P2_P1_ADDRESS_REG_20_(vec[435]), .P2_P1_ADDRESS_REG_19_(vec[434]), .P2_P1_ADDRESS_REG_18_(vec[433]), .P2_P1_ADDRESS_REG_17_(vec[432]), .P2_P1_ADDRESS_REG_16_(vec[431]), .P2_P1_ADDRESS_REG_15_(vec[430]), .P2_P1_ADDRESS_REG_14_(vec[429]), .P2_P1_ADDRESS_REG_13_(vec[428]), .P2_P1_ADDRESS_REG_12_(vec[427]), .P2_P1_ADDRESS_REG_11_(vec[426]), .P2_P1_ADDRESS_REG_10_(vec[425]), .P2_P1_ADDRESS_REG_9_(vec[424]), .P2_P1_ADDRESS_REG_8_(vec[423]), .P2_P1_ADDRESS_REG_7_(vec[422]), .P2_P1_ADDRESS_REG_6_(vec[421]), .P2_P1_ADDRESS_REG_5_(vec[420]), .P2_P1_ADDRESS_REG_4_(vec[419]), .P2_P1_ADDRESS_REG_3_(vec[418]), .P2_P1_ADDRESS_REG_2_(vec[417]), .P2_P1_ADDRESS_REG_1_(vec[416]), .P2_P1_ADDRESS_REG_0_(vec[415]), .P2_P1_STATE_REG_2_(vec[414]), .P2_P1_STATE_REG_1_(vec[413]), .P2_P1_STATE_REG_0_(vec[412]), .P2_P1_DATAWIDTH_REG_0_(vec[411]), .P2_P1_DATAWIDTH_REG_1_(vec[410]), .P2_P1_DATAWIDTH_REG_2_(vec[409]), .P2_P1_DATAWIDTH_REG_3_(vec[408]), .P2_P1_DATAWIDTH_REG_4_(vec[407]), .P2_P1_DATAWIDTH_REG_5_(vec[406]), .P2_P1_DATAWIDTH_REG_6_(vec[405]), .P2_P1_DATAWIDTH_REG_7_(vec[404]), .P2_P1_DATAWIDTH_REG_8_(vec[403]), .P2_P1_DATAWIDTH_REG_9_(vec[402]), .P2_P1_DATAWIDTH_REG_10_(vec[401]), .P2_P1_DATAWIDTH_REG_11_(vec[400]), .P2_P1_DATAWIDTH_REG_12_(vec[399]), .P2_P1_DATAWIDTH_REG_13_(vec[398]), .P2_P1_DATAWIDTH_REG_14_(vec[397]), .P2_P1_DATAWIDTH_REG_15_(vec[396]), .P2_P1_DATAWIDTH_REG_16_(vec[395]), .P2_P1_DATAWIDTH_REG_17_(vec[394]), .P2_P1_DATAWIDTH_REG_18_(vec[393]), .P2_P1_DATAWIDTH_REG_19_(vec[392]), .P2_P1_DATAWIDTH_REG_20_(vec[391]), .P2_P1_DATAWIDTH_REG_21_(vec[390]), .P2_P1_DATAWIDTH_REG_22_(vec[389]), .P2_P1_DATAWIDTH_REG_23_(vec[388]), .P2_P1_DATAWIDTH_REG_24_(vec[387]), .P2_P1_DATAWIDTH_REG_25_(vec[386]), .P2_P1_DATAWIDTH_REG_26_(vec[385]), .P2_P1_DATAWIDTH_REG_27_(vec[384]), .P2_P1_DATAWIDTH_REG_28_(vec[383]), .P2_P1_DATAWIDTH_REG_29_(vec[382]), .P2_P1_DATAWIDTH_REG_30_(vec[381]), .P2_P1_DATAWIDTH_REG_31_(vec[380]), .P2_P1_STATE2_REG_3_(vec[379]), .P2_P1_STATE2_REG_2_(vec[378]), .P2_P1_STATE2_REG_1_(vec[377]), .P2_P1_STATE2_REG_0_(vec[376]), .P2_P1_INSTQUEUE_REG_15__7_(vec[375]), .P2_P1_INSTQUEUE_REG_15__6_(vec[374]), .P2_P1_INSTQUEUE_REG_15__5_(vec[373]), .P2_P1_INSTQUEUE_REG_15__4_(vec[372]), .P2_P1_INSTQUEUE_REG_15__3_(vec[371]), .P2_P1_INSTQUEUE_REG_15__2_(vec[370]), .P2_P1_INSTQUEUE_REG_15__1_(vec[369]), .P2_P1_INSTQUEUE_REG_15__0_(vec[368]), .P2_P1_INSTQUEUE_REG_14__7_(vec[367]), .P2_P1_INSTQUEUE_REG_14__6_(vec[366]), .P2_P1_INSTQUEUE_REG_14__5_(vec[365]), .P2_P1_INSTQUEUE_REG_14__4_(vec[364]), .P2_P1_INSTQUEUE_REG_14__3_(vec[363]), .P2_P1_INSTQUEUE_REG_14__2_(vec[362]), .P2_P1_INSTQUEUE_REG_14__1_(vec[361]), .P2_P1_INSTQUEUE_REG_14__0_(vec[360]), .P2_P1_INSTQUEUE_REG_13__7_(vec[359]), .P2_P1_INSTQUEUE_REG_13__6_(vec[358]), .P2_P1_INSTQUEUE_REG_13__5_(vec[357]), .P2_P1_INSTQUEUE_REG_13__4_(vec[356]), .P2_P1_INSTQUEUE_REG_13__3_(vec[355]), .P2_P1_INSTQUEUE_REG_13__2_(vec[354]), .P2_P1_INSTQUEUE_REG_13__1_(vec[353]), .P2_P1_INSTQUEUE_REG_13__0_(vec[352]), .P2_P1_INSTQUEUE_REG_12__7_(vec[351]), .P2_P1_INSTQUEUE_REG_12__6_(vec[350]), .P2_P1_INSTQUEUE_REG_12__5_(vec[349]), .P2_P1_INSTQUEUE_REG_12__4_(vec[348]), .P2_P1_INSTQUEUE_REG_12__3_(vec[347]), .P2_P1_INSTQUEUE_REG_12__2_(vec[346]), .P2_P1_INSTQUEUE_REG_12__1_(vec[345]), .P2_P1_INSTQUEUE_REG_12__0_(vec[344]), .P2_P1_INSTQUEUE_REG_11__7_(vec[343]), .P2_P1_INSTQUEUE_REG_11__6_(vec[342]), .P2_P1_INSTQUEUE_REG_11__5_(vec[341]), .P2_P1_INSTQUEUE_REG_11__4_(vec[340]), .P2_P1_INSTQUEUE_REG_11__3_(vec[339]), .P2_P1_INSTQUEUE_REG_11__2_(vec[338]), .P2_P1_INSTQUEUE_REG_11__1_(vec[337]), .P2_P1_INSTQUEUE_REG_11__0_(vec[336]), .P2_P1_INSTQUEUE_REG_10__7_(vec[335]), .P2_P1_INSTQUEUE_REG_10__6_(vec[334]), .P2_P1_INSTQUEUE_REG_10__5_(vec[333]), .P2_P1_INSTQUEUE_REG_10__4_(vec[332]), .P2_P1_INSTQUEUE_REG_10__3_(vec[331]), .P2_P1_INSTQUEUE_REG_10__2_(vec[330]), .P2_P1_INSTQUEUE_REG_10__1_(vec[329]), .P2_P1_INSTQUEUE_REG_10__0_(vec[328]), .P2_P1_INSTQUEUE_REG_9__7_(vec[327]), .P2_P1_INSTQUEUE_REG_9__6_(vec[326]), .P2_P1_INSTQUEUE_REG_9__5_(vec[325]), .P2_P1_INSTQUEUE_REG_9__4_(vec[324]), .P2_P1_INSTQUEUE_REG_9__3_(vec[323]), .P2_P1_INSTQUEUE_REG_9__2_(vec[322]), .P2_P1_INSTQUEUE_REG_9__1_(vec[321]), .P2_P1_INSTQUEUE_REG_9__0_(vec[320]), .P2_P1_INSTQUEUE_REG_8__7_(vec[319]), .P2_P1_INSTQUEUE_REG_8__6_(vec[318]), .P2_P1_INSTQUEUE_REG_8__5_(vec[317]), .P2_P1_INSTQUEUE_REG_8__4_(vec[316]), .P2_P1_INSTQUEUE_REG_8__3_(vec[315]), .P2_P1_INSTQUEUE_REG_8__2_(vec[314]), .P2_P1_INSTQUEUE_REG_8__1_(vec[313]), .P2_P1_INSTQUEUE_REG_8__0_(vec[312]), .P2_P1_INSTQUEUE_REG_7__7_(vec[311]), .P2_P1_INSTQUEUE_REG_7__6_(vec[310]), .P2_P1_INSTQUEUE_REG_7__5_(vec[309]), .P2_P1_INSTQUEUE_REG_7__4_(vec[308]), .P2_P1_INSTQUEUE_REG_7__3_(vec[307]), .P2_P1_INSTQUEUE_REG_7__2_(vec[306]), .P2_P1_INSTQUEUE_REG_7__1_(vec[305]), .P2_P1_INSTQUEUE_REG_7__0_(vec[304]), .P2_P1_INSTQUEUE_REG_6__7_(vec[303]), .P2_P1_INSTQUEUE_REG_6__6_(vec[302]), .P2_P1_INSTQUEUE_REG_6__5_(vec[301]), .P2_P1_INSTQUEUE_REG_6__4_(vec[300]), .P2_P1_INSTQUEUE_REG_6__3_(vec[299]), .P2_P1_INSTQUEUE_REG_6__2_(vec[298]), .P2_P1_INSTQUEUE_REG_6__1_(vec[297]), .P2_P1_INSTQUEUE_REG_6__0_(vec[296]), .P2_P1_INSTQUEUE_REG_5__7_(vec[295]), .P2_P1_INSTQUEUE_REG_5__6_(vec[294]), .P2_P1_INSTQUEUE_REG_5__5_(vec[293]), .P2_P1_INSTQUEUE_REG_5__4_(vec[292]), .P2_P1_INSTQUEUE_REG_5__3_(vec[291]), .P2_P1_INSTQUEUE_REG_5__2_(vec[290]), .P2_P1_INSTQUEUE_REG_5__1_(vec[289]), .P2_P1_INSTQUEUE_REG_5__0_(vec[288]), .P2_P1_INSTQUEUE_REG_4__7_(vec[287]), .P2_P1_INSTQUEUE_REG_4__6_(vec[286]), .P2_P1_INSTQUEUE_REG_4__5_(vec[285]), .P2_P1_INSTQUEUE_REG_4__4_(vec[284]), .P2_P1_INSTQUEUE_REG_4__3_(vec[283]), .P2_P1_INSTQUEUE_REG_4__2_(vec[282]), .P2_P1_INSTQUEUE_REG_4__1_(vec[281]), .P2_P1_INSTQUEUE_REG_4__0_(vec[280]), .P2_P1_INSTQUEUE_REG_3__7_(vec[279]), .P2_P1_INSTQUEUE_REG_3__6_(vec[278]), .P2_P1_INSTQUEUE_REG_3__5_(vec[277]), .P2_P1_INSTQUEUE_REG_3__4_(vec[276]), .P2_P1_INSTQUEUE_REG_3__3_(vec[275]), .P2_P1_INSTQUEUE_REG_3__2_(vec[274]), .P2_P1_INSTQUEUE_REG_3__1_(vec[273]), .P2_P1_INSTQUEUE_REG_3__0_(vec[272]), .P2_P1_INSTQUEUE_REG_2__7_(vec[271]), .P2_P1_INSTQUEUE_REG_2__6_(vec[270]), .P2_P1_INSTQUEUE_REG_2__5_(vec[269]), .P2_P1_INSTQUEUE_REG_2__4_(vec[268]), .P2_P1_INSTQUEUE_REG_2__3_(vec[267]), .P2_P1_INSTQUEUE_REG_2__2_(vec[266]), .P2_P1_INSTQUEUE_REG_2__1_(vec[265]), .P2_P1_INSTQUEUE_REG_2__0_(vec[264]), .P2_P1_INSTQUEUE_REG_1__7_(vec[263]), .P2_P1_INSTQUEUE_REG_1__6_(vec[262]), .P2_P1_INSTQUEUE_REG_1__5_(vec[261]), .P2_P1_INSTQUEUE_REG_1__4_(vec[260]), .P2_P1_INSTQUEUE_REG_1__3_(vec[259]), .P2_P1_INSTQUEUE_REG_1__2_(vec[258]), .P2_P1_INSTQUEUE_REG_1__1_(vec[257]), .P2_P1_INSTQUEUE_REG_1__0_(vec[256]), .P2_P1_INSTQUEUE_REG_0__7_(vec[255]), .P2_P1_INSTQUEUE_REG_0__6_(vec[254]), .P2_P1_INSTQUEUE_REG_0__5_(vec[253]), .P2_P1_INSTQUEUE_REG_0__4_(vec[252]), .P2_P1_INSTQUEUE_REG_0__3_(vec[251]), .P2_P1_INSTQUEUE_REG_0__2_(vec[250]), .P2_P1_INSTQUEUE_REG_0__1_(vec[249]), .P2_P1_INSTQUEUE_REG_0__0_(vec[248]), .P2_P1_INSTQUEUERD_ADDR_REG_4_(vec[247]), .P2_P1_INSTQUEUERD_ADDR_REG_3_(vec[246]), .P2_P1_INSTQUEUERD_ADDR_REG_2_(vec[245]), .P2_P1_INSTQUEUERD_ADDR_REG_1_(vec[244]), .P2_P1_INSTQUEUERD_ADDR_REG_0_(vec[243]), .P2_P1_INSTQUEUEWR_ADDR_REG_4_(vec[242]), .P2_P1_INSTQUEUEWR_ADDR_REG_3_(vec[241]), .P2_P1_INSTQUEUEWR_ADDR_REG_2_(vec[240]), .P2_P1_INSTQUEUEWR_ADDR_REG_1_(vec[239]), .P2_P1_INSTQUEUEWR_ADDR_REG_0_(vec[238]), .P2_P1_INSTADDRPOINTER_REG_0_(vec[237]), .P2_P1_INSTADDRPOINTER_REG_1_(vec[236]), .P2_P1_INSTADDRPOINTER_REG_2_(vec[235]), .P2_P1_INSTADDRPOINTER_REG_3_(vec[234]), .P2_P1_INSTADDRPOINTER_REG_4_(vec[233]), .P2_P1_INSTADDRPOINTER_REG_5_(vec[232]), .P2_P1_INSTADDRPOINTER_REG_6_(vec[231]), .P2_P1_INSTADDRPOINTER_REG_7_(vec[230]), .P2_P1_INSTADDRPOINTER_REG_8_(vec[229]), .P2_P1_INSTADDRPOINTER_REG_9_(vec[228]), .P2_P1_INSTADDRPOINTER_REG_10_(vec[227]), .P2_P1_INSTADDRPOINTER_REG_11_(vec[226]), .P2_P1_INSTADDRPOINTER_REG_12_(vec[225]), .P2_P1_INSTADDRPOINTER_REG_13_(vec[224]), .P2_P1_INSTADDRPOINTER_REG_14_(vec[223]), .P2_P1_INSTADDRPOINTER_REG_15_(vec[222]), .P2_P1_INSTADDRPOINTER_REG_16_(vec[221]), .P2_P1_INSTADDRPOINTER_REG_17_(vec[220]), .P2_P1_INSTADDRPOINTER_REG_18_(vec[219]), .P2_P1_INSTADDRPOINTER_REG_19_(vec[218]), .P2_P1_INSTADDRPOINTER_REG_20_(vec[217]), .P2_P1_INSTADDRPOINTER_REG_21_(vec[216]), .P2_P1_INSTADDRPOINTER_REG_22_(vec[215]), .P2_P1_INSTADDRPOINTER_REG_23_(vec[214]), .P2_P1_INSTADDRPOINTER_REG_24_(vec[213]), .P2_P1_INSTADDRPOINTER_REG_25_(vec[212]), .P2_P1_INSTADDRPOINTER_REG_26_(vec[211]), .P2_P1_INSTADDRPOINTER_REG_27_(vec[210]), .P2_P1_INSTADDRPOINTER_REG_28_(vec[209]), .P2_P1_INSTADDRPOINTER_REG_29_(vec[208]), .P2_P1_INSTADDRPOINTER_REG_30_(vec[207]), .P2_P1_INSTADDRPOINTER_REG_31_(vec[206]), .P2_P1_PHYADDRPOINTER_REG_0_(vec[205]), .P2_P1_PHYADDRPOINTER_REG_1_(vec[204]), .P2_P1_PHYADDRPOINTER_REG_2_(vec[203]), .P2_P1_PHYADDRPOINTER_REG_3_(vec[202]), .P2_P1_PHYADDRPOINTER_REG_4_(vec[201]), .P2_P1_PHYADDRPOINTER_REG_5_(vec[200]), .P2_P1_PHYADDRPOINTER_REG_6_(vec[199]), .P2_P1_PHYADDRPOINTER_REG_7_(vec[198]), .P2_P1_PHYADDRPOINTER_REG_8_(vec[197]), .P2_P1_PHYADDRPOINTER_REG_9_(vec[196]), .P2_P1_PHYADDRPOINTER_REG_10_(vec[195]), .P2_P1_PHYADDRPOINTER_REG_11_(vec[194]), .P2_P1_PHYADDRPOINTER_REG_12_(vec[193]), .P2_P1_PHYADDRPOINTER_REG_13_(vec[192]), .P2_P1_PHYADDRPOINTER_REG_14_(vec[191]), .P2_P1_PHYADDRPOINTER_REG_15_(vec[190]), .P2_P1_PHYADDRPOINTER_REG_16_(vec[189]), .P2_P1_PHYADDRPOINTER_REG_17_(vec[188]), .P2_P1_PHYADDRPOINTER_REG_18_(vec[187]), .P2_P1_PHYADDRPOINTER_REG_19_(vec[186]), .P2_P1_PHYADDRPOINTER_REG_20_(vec[185]), .P2_P1_PHYADDRPOINTER_REG_21_(vec[184]), .P2_P1_PHYADDRPOINTER_REG_22_(vec[183]), .P2_P1_PHYADDRPOINTER_REG_23_(vec[182]), .P2_P1_PHYADDRPOINTER_REG_24_(vec[181]), .P2_P1_PHYADDRPOINTER_REG_25_(vec[180]), .P2_P1_PHYADDRPOINTER_REG_26_(vec[179]), .P2_P1_PHYADDRPOINTER_REG_27_(vec[178]), .P2_P1_PHYADDRPOINTER_REG_28_(vec[177]), .P2_P1_PHYADDRPOINTER_REG_29_(vec[176]), .P2_P1_PHYADDRPOINTER_REG_30_(vec[175]), .P2_P1_PHYADDRPOINTER_REG_31_(vec[174]), .P2_P1_LWORD_REG_15_(vec[173]), .P2_P1_LWORD_REG_14_(vec[172]), .P2_P1_LWORD_REG_13_(vec[171]), .P2_P1_LWORD_REG_12_(vec[170]), .P2_P1_LWORD_REG_11_(vec[169]), .P2_P1_LWORD_REG_10_(vec[168]), .P2_P1_LWORD_REG_9_(vec[167]), .P2_P1_LWORD_REG_8_(vec[166]), .P2_P1_LWORD_REG_7_(vec[165]), .P2_P1_LWORD_REG_6_(vec[164]), .P2_P1_LWORD_REG_5_(vec[163]), .P2_P1_LWORD_REG_4_(vec[162]), .P2_P1_LWORD_REG_3_(vec[161]), .P2_P1_LWORD_REG_2_(vec[160]), .P2_P1_LWORD_REG_1_(vec[159]), .P2_P1_LWORD_REG_0_(vec[158]), .P2_P1_UWORD_REG_14_(vec[157]), .P2_P1_UWORD_REG_13_(vec[156]), .P2_P1_UWORD_REG_12_(vec[155]), .P2_P1_UWORD_REG_11_(vec[154]), .P2_P1_UWORD_REG_10_(vec[153]), .P2_P1_UWORD_REG_9_(vec[152]), .P2_P1_UWORD_REG_8_(vec[151]), .P2_P1_UWORD_REG_7_(vec[150]), .P2_P1_UWORD_REG_6_(vec[149]), .P2_P1_UWORD_REG_5_(vec[148]), .P2_P1_UWORD_REG_4_(vec[147]), .P2_P1_UWORD_REG_3_(vec[146]), .P2_P1_UWORD_REG_2_(vec[145]), .P2_P1_UWORD_REG_1_(vec[144]), .P2_P1_UWORD_REG_0_(vec[143]), .P2_P1_DATAO_REG_0_(vec[142]), .P2_P1_DATAO_REG_1_(vec[141]), .P2_P1_DATAO_REG_2_(vec[140]), .P2_P1_DATAO_REG_3_(vec[139]), .P2_P1_DATAO_REG_4_(vec[138]), .P2_P1_DATAO_REG_5_(vec[137]), .P2_P1_DATAO_REG_6_(vec[136]), .P2_P1_DATAO_REG_7_(vec[135]), .P2_P1_DATAO_REG_8_(vec[134]), .P2_P1_DATAO_REG_9_(vec[133]), .P2_P1_DATAO_REG_10_(vec[132]), .P2_P1_DATAO_REG_11_(vec[131]), .P2_P1_DATAO_REG_12_(vec[130]), .P2_P1_DATAO_REG_13_(vec[129]), .P2_P1_DATAO_REG_14_(vec[128]), .P2_P1_DATAO_REG_15_(vec[127]), .P2_P1_DATAO_REG_16_(vec[126]), .P2_P1_DATAO_REG_17_(vec[125]), .P2_P1_DATAO_REG_18_(vec[124]), .P2_P1_DATAO_REG_19_(vec[123]), .P2_P1_DATAO_REG_20_(vec[122]), .P2_P1_DATAO_REG_21_(vec[121]), .P2_P1_DATAO_REG_22_(vec[120]), .P2_P1_DATAO_REG_23_(vec[119]), .P2_P1_DATAO_REG_24_(vec[118]), .P2_P1_DATAO_REG_25_(vec[117]), .P2_P1_DATAO_REG_26_(vec[116]), .P2_P1_DATAO_REG_27_(vec[115]), .P2_P1_DATAO_REG_28_(vec[114]), .P2_P1_DATAO_REG_29_(vec[113]), .P2_P1_DATAO_REG_30_(vec[112]), .P2_P1_DATAO_REG_31_(vec[111]), .P2_P1_EAX_REG_0_(vec[110]), .P2_P1_EAX_REG_1_(vec[109]), .P2_P1_EAX_REG_2_(vec[108]), .P2_P1_EAX_REG_3_(vec[107]), .P2_P1_EAX_REG_4_(vec[106]), .P2_P1_EAX_REG_5_(vec[105]), .P2_P1_EAX_REG_6_(vec[104]), .P2_P1_EAX_REG_7_(vec[103]), .P2_P1_EAX_REG_8_(vec[102]), .P2_P1_EAX_REG_9_(vec[101]), .P2_P1_EAX_REG_10_(vec[100]), .P2_P1_EAX_REG_11_(vec[99]), .P2_P1_EAX_REG_12_(vec[98]), .P2_P1_EAX_REG_13_(vec[97]), .P2_P1_EAX_REG_14_(vec[96]), .P2_P1_EAX_REG_15_(vec[95]), .P2_P1_EAX_REG_16_(vec[94]), .P2_P1_EAX_REG_17_(vec[93]), .P2_P1_EAX_REG_18_(vec[92]), .P2_P1_EAX_REG_19_(vec[91]), .P2_P1_EAX_REG_20_(vec[90]), .P2_P1_EAX_REG_21_(vec[89]), .P2_P1_EAX_REG_22_(vec[88]), .P2_P1_EAX_REG_23_(vec[87]), .P2_P1_EAX_REG_24_(vec[86]), .P2_P1_EAX_REG_25_(vec[85]), .P2_P1_EAX_REG_26_(vec[84]), .P2_P1_EAX_REG_27_(vec[83]), .P2_P1_EAX_REG_28_(vec[82]), .P2_P1_EAX_REG_29_(vec[81]), .P2_P1_EAX_REG_30_(vec[80]), .P2_P1_EAX_REG_31_(vec[79]), .P2_P1_EBX_REG_0_(vec[78]), .P2_P1_EBX_REG_1_(vec[77]), .P2_P1_EBX_REG_2_(vec[76]), .P2_P1_EBX_REG_3_(vec[75]), .P2_P1_EBX_REG_4_(vec[74]), .P2_P1_EBX_REG_5_(vec[73]), .P2_P1_EBX_REG_6_(vec[72]), .P2_P1_EBX_REG_7_(vec[71]), .P2_P1_EBX_REG_8_(vec[70]), .P2_P1_EBX_REG_9_(vec[69]), .P2_P1_EBX_REG_10_(vec[68]), .P2_P1_EBX_REG_11_(vec[67]), .P2_P1_EBX_REG_12_(vec[66]), .P2_P1_EBX_REG_13_(vec[65]), .P2_P1_EBX_REG_14_(vec[64]), .P2_P1_EBX_REG_15_(vec[63]), .P2_P1_EBX_REG_16_(vec[62]), .P2_P1_EBX_REG_17_(vec[61]), .P2_P1_EBX_REG_18_(vec[60]), .P2_P1_EBX_REG_19_(vec[59]), .P2_P1_EBX_REG_20_(vec[58]), .P2_P1_EBX_REG_21_(vec[57]), .P2_P1_EBX_REG_22_(vec[56]), .P2_P1_EBX_REG_23_(vec[55]), .P2_P1_EBX_REG_24_(vec[54]), .P2_P1_EBX_REG_25_(vec[53]), .P2_P1_EBX_REG_26_(vec[52]), .P2_P1_EBX_REG_27_(vec[51]), .P2_P1_EBX_REG_28_(vec[50]), .P2_P1_EBX_REG_29_(vec[49]), .P2_P1_EBX_REG_30_(vec[48]), .P2_P1_EBX_REG_31_(vec[47]), .P2_P1_REIP_REG_0_(vec[46]), .P2_P1_REIP_REG_1_(vec[45]), .P2_P1_REIP_REG_2_(vec[44]), .P2_P1_REIP_REG_3_(vec[43]), .P2_P1_REIP_REG_4_(vec[42]), .P2_P1_REIP_REG_5_(vec[41]), .P2_P1_REIP_REG_6_(vec[40]), .P2_P1_REIP_REG_7_(vec[39]), .P2_P1_REIP_REG_8_(vec[38]), .P2_P1_REIP_REG_9_(vec[37]), .P2_P1_REIP_REG_10_(vec[36]), .P2_P1_REIP_REG_11_(vec[35]), .P2_P1_REIP_REG_12_(vec[34]), .P2_P1_REIP_REG_13_(vec[33]), .P2_P1_REIP_REG_14_(vec[32]), .P2_P1_REIP_REG_15_(vec[31]), .P2_P1_REIP_REG_16_(vec[30]), .P2_P1_REIP_REG_17_(vec[29]), .P2_P1_REIP_REG_18_(vec[28]), .P2_P1_REIP_REG_19_(vec[27]), .P2_P1_REIP_REG_20_(vec[26]), .P2_P1_REIP_REG_21_(vec[25]), .P2_P1_REIP_REG_22_(vec[24]), .P2_P1_REIP_REG_23_(vec[23]), .P2_P1_REIP_REG_24_(vec[22]), .P2_P1_REIP_REG_25_(vec[21]), .P2_P1_REIP_REG_26_(vec[20]), .P2_P1_REIP_REG_27_(vec[19]), .P2_P1_REIP_REG_28_(vec[18]), .P2_P1_REIP_REG_29_(vec[17]), .P2_P1_REIP_REG_30_(vec[16]), .P2_P1_REIP_REG_31_(vec[15]), .P2_P1_BYTEENABLE_REG_3_(vec[14]), .P2_P1_BYTEENABLE_REG_2_(vec[13]), .P2_P1_BYTEENABLE_REG_1_(vec[12]), .P2_P1_BYTEENABLE_REG_0_(vec[11]), .P2_P1_W_R_N_REG(vec[10]), .P2_P1_FLUSH_REG(vec[9]), .P2_P1_MORE_REG(vec[8]), .P2_P1_STATEBS16_REG(vec[7]), .P2_P1_REQUESTPENDING_REG(vec[6]), .P2_P1_D_C_N_REG(vec[5]), .P2_P1_M_IO_N_REG(vec[4]), .P2_P1_CODEFETCH_REG(vec[3]), .P2_P1_ADS_N_REG(vec[2]), .P2_P1_READREQUEST_REG(vec[1]), .P2_P1_MEMORYFETCH_REG(vec[0]), .LOGIC0_PO_EXTRA(logic0_po_extra), .MUL_1411_U378(mul_1411_u378), .MUL_1411_U438(mul_1411_u438), .MUL_1411_U10(mul_1411_u10), .MUL_1411_U439(mul_1411_u439), .MUL_1411_U9(mul_1411_u9), .MUL_1411_U440(mul_1411_u440), .MUL_1411_U8(mul_1411_u8), .MUL_1411_U441(mul_1411_u441), .MUL_1411_U7(mul_1411_u7), .MUL_1411_U385(mul_1411_u385), .MUL_1411_U14(mul_1411_u14), .MUL_1411_U386(mul_1411_u386), .MUL_1411_U13(mul_1411_u13), .MUL_1411_U387(mul_1411_u387), .MUL_1411_U12(mul_1411_u12), .MUL_1411_U388(mul_1411_u388), .MUL_1411_U11(mul_1411_u11), .MUL_1411_U15(mul_1411_u15), .MUL_1411_U5_PO_EXTRA(mul_1411_u5_po_extra), .MUL_1421_A1_U5(mul_1421_a1_u5), .U154(u154), .U39_PO_EXTRA(u39_po_extra), .P1_U247(p1_u247), .P1_U246(p1_u246), .P1_U245(p1_u245), .P1_U244(p1_u244), .P1_U243(p1_u243), .P1_U242(p1_u242), .P1_U241(p1_u241), .P1_U240(p1_u240), .P1_U239(p1_u239), .P1_U238(p1_u238), .P1_U237(p1_u237), .P1_U236(p1_u236), .P1_U235(p1_u235), .P1_U234(p1_u234), .P1_U233(p1_u233), .P1_U232(p1_u232), .P1_U231(p1_u231), .P1_U230(p1_u230), .P1_U229(p1_u229), .P1_U228(p1_u228), .P1_U227(p1_u227), .P1_U226(p1_u226), .P1_U225(p1_u225), .P1_U224(p1_u224), .P1_U223(p1_u223), .P1_U222(p1_u222), .P1_U221(p1_u221), .P1_U220(p1_u220), .P1_U219(p1_u219), .P1_U218(p1_u218), .P1_U217(p1_u217), .P1_U216(p1_u216), .P1_U251(p1_u251), .P1_U252(p1_u252), .P1_U253(p1_u253), .P1_U254(p1_u254), .P1_U255(p1_u255), .P1_U256(p1_u256), .P1_U257(p1_u257), .P1_U258(p1_u258), .P1_U259(p1_u259), .P1_U260(p1_u260), .P1_U261(p1_u261), .P1_U262(p1_u262), .P1_U263(p1_u263), .P1_U264(p1_u264), .P1_U265(p1_u265), .P1_U266(p1_u266), .P1_U267(p1_u267), .P1_U268(p1_u268), .P1_U269(p1_u269), .P1_U270(p1_u270), .P1_U271(p1_u271), .P1_U272(p1_u272), .P1_U273(p1_u273), .P1_U274(p1_u274), .P1_U275(p1_u275), .P1_U276(p1_u276), .P1_U277(p1_u277), .P1_U278(p1_u278), .P1_U279(p1_u279), .P1_U280(p1_u280), .P1_U281(p1_u281), .P1_U282(p1_u282), .P1_U212(p1_u212), .P1_U215(p1_u215), .P1_U213(p1_u213), .P1_U214(p1_u214), .P2_U247(p2_u247), .P2_U246(p2_u246), .P2_U245(p2_u245), .P2_U244(p2_u244), .P2_U243(p2_u243), .P2_U242(p2_u242), .P2_U241(p2_u241), .P2_U240(p2_u240), .P2_U239(p2_u239), .P2_U238(p2_u238), .P2_U237(p2_u237), .P2_U236(p2_u236), .P2_U235(p2_u235), .P2_U234(p2_u234), .P2_U233(p2_u233), .P2_U232(p2_u232), .P2_U231(p2_u231), .P2_U230(p2_u230), .P2_U229(p2_u229), .P2_U228(p2_u228), .P2_U227(p2_u227), .P2_U226(p2_u226), .P2_U225(p2_u225), .P2_U224(p2_u224), .P2_U223(p2_u223), .P2_U222(p2_u222), .P2_U221(p2_u221), .P2_U220(p2_u220), .P2_U219(p2_u219), .P2_U218(p2_u218), .P2_U217(p2_u217), .P2_U216(p2_u216), .P2_U251(p2_u251), .P2_U252(p2_u252), .P2_U253(p2_u253), .P2_U254(p2_u254), .P2_U255(p2_u255), .P2_U256(p2_u256), .P2_U257(p2_u257), .P2_U258(p2_u258), .P2_U259(p2_u259), .P2_U260(p2_u260), .P2_U261(p2_u261), .P2_U262(p2_u262), .P2_U263(p2_u263), .P2_U264(p2_u264), .P2_U265(p2_u265), .P2_U266(p2_u266), .P2_U267(p2_u267), .P2_U268(p2_u268), .P2_U269(p2_u269), .P2_U270(p2_u270), .P2_U271(p2_u271), .P2_U272(p2_u272), .P2_U273(p2_u273), .P2_U274(p2_u274), .P2_U275(p2_u275), .P2_U276(p2_u276), .P2_U277(p2_u277), .P2_U278(p2_u278), .P2_U279(p2_u279), .P2_U280(p2_u280), .P2_U281(p2_u281), .P2_U282(p2_u282), .P2_U212(p2_u212), .P2_U215(p2_u215), .P2_U213(p2_u213), .P2_U214(p2_u214), .P3_U3354(p3_u3354), .P3_U3353(p3_u3353), .P3_U3352(p3_u3352), .P3_U3351(p3_u3351), .P3_U3350(p3_u3350), .P3_U3349(p3_u3349), .P3_U3348(p3_u3348), .P3_U3347(p3_u3347), .P3_U3346(p3_u3346), .P3_U3345(p3_u3345), .P3_U3344(p3_u3344), .P3_U3343(p3_u3343), .P3_U3342(p3_u3342), .P3_U3341(p3_u3341), .P3_U3340(p3_u3340), .P3_U3339(p3_u3339), .P3_U3338(p3_u3338), .P3_U3337(p3_u3337), .P3_U3336(p3_u3336), .P3_U3335(p3_u3335), .P3_U3334(p3_u3334), .P3_U3333(p3_u3333), .P3_U3332(p3_u3332), .P3_U3331(p3_u3331), .P3_U3330(p3_u3330), .P3_U3329(p3_u3329), .P3_U3328(p3_u3328), .P3_U3327(p3_u3327), .P3_U3326(p3_u3326), .P3_U3325(p3_u3325), .P3_U3324(p3_u3324), .P3_U3323(p3_u3323), .P3_U3442(p3_u3442), .P3_U3443(p3_u3443), .P3_U3322(p3_u3322), .P3_U3321(p3_u3321), .P3_U3320(p3_u3320), .P3_U3319(p3_u3319), .P3_U3318(p3_u3318), .P3_U3317(p3_u3317), .P3_U3316(p3_u3316), .P3_U3315(p3_u3315), .P3_U3314(p3_u3314), .P3_U3313(p3_u3313), .P3_U3312(p3_u3312), .P3_U3311(p3_u3311), .P3_U3310(p3_u3310), .P3_U3309(p3_u3309), .P3_U3308(p3_u3308), .P3_U3307(p3_u3307), .P3_U3306(p3_u3306), .P3_U3305(p3_u3305), .P3_U3304(p3_u3304), .P3_U3303(p3_u3303), .P3_U3302(p3_u3302), .P3_U3301(p3_u3301), .P3_U3300(p3_u3300), .P3_U3299(p3_u3299), .P3_U3298(p3_u3298), .P3_U3297(p3_u3297), .P3_U3296(p3_u3296), .P3_U3295(p3_u3295), .P3_U3294(p3_u3294), .P3_U3293(p3_u3293), .P3_U3456(p3_u3456), .P3_U3459(p3_u3459), .P3_U3462(p3_u3462), .P3_U3465(p3_u3465), .P3_U3468(p3_u3468), .P3_U3471(p3_u3471), .P3_U3474(p3_u3474), .P3_U3477(p3_u3477), .P3_U3480(p3_u3480), .P3_U3483(p3_u3483), .P3_U3486(p3_u3486), .P3_U3489(p3_u3489), .P3_U3492(p3_u3492), .P3_U3495(p3_u3495), .P3_U3498(p3_u3498), .P3_U3501(p3_u3501), .P3_U3504(p3_u3504), .P3_U3507(p3_u3507), .P3_U3510(p3_u3510), .P3_U3512(p3_u3512), .P3_U3513(p3_u3513), .P3_U3514(p3_u3514), .P3_U3515(p3_u3515), .P3_U3516(p3_u3516), .P3_U3517(p3_u3517), .P3_U3518(p3_u3518), .P3_U3519(p3_u3519), .P3_U3520(p3_u3520), .P3_U3521(p3_u3521), .P3_U3522(p3_u3522), .P3_U3523(p3_u3523), .P3_U3524(p3_u3524), .P3_U3525(p3_u3525), .P3_U3526(p3_u3526), .P3_U3527(p3_u3527), .P3_U3528(p3_u3528), .P3_U3529(p3_u3529), .P3_U3530(p3_u3530), .P3_U3531(p3_u3531), .P3_U3532(p3_u3532), .P3_U3533(p3_u3533), .P3_U3534(p3_u3534), .P3_U3535(p3_u3535), .P3_U3536(p3_u3536), .P3_U3537(p3_u3537), .P3_U3538(p3_u3538), .P3_U3539(p3_u3539), .P3_U3540(p3_u3540), .P3_U3541(p3_u3541), .P3_U3542(p3_u3542), .P3_U3543(p3_u3543), .P3_U3544(p3_u3544), .P3_U3545(p3_u3545), .P3_U3546(p3_u3546), .P3_U3547(p3_u3547), .P3_U3548(p3_u3548), .P3_U3549(p3_u3549), .P3_U3550(p3_u3550), .P3_U3551(p3_u3551), .P3_U3552(p3_u3552), .P3_U3553(p3_u3553), .P3_U3554(p3_u3554), .P3_U3555(p3_u3555), .P3_U3556(p3_u3556), .P3_U3292(p3_u3292), .P3_U3291(p3_u3291), .P3_U3290(p3_u3290), .P3_U3289(p3_u3289), .P3_U3288(p3_u3288), .P3_U3287(p3_u3287), .P3_U3286(p3_u3286), .P3_U3285(p3_u3285), .P3_U3284(p3_u3284), .P3_U3283(p3_u3283), .P3_U3282(p3_u3282), .P3_U3281(p3_u3281), .P3_U3280(p3_u3280), .P3_U3279(p3_u3279), .P3_U3278(p3_u3278), .P3_U3277(p3_u3277), .P3_U3276(p3_u3276), .P3_U3275(p3_u3275), .P3_U3274(p3_u3274), .P3_U3273(p3_u3273), .P3_U3272(p3_u3272), .P3_U3271(p3_u3271), .P3_U3270(p3_u3270), .P3_U3269(p3_u3269), .P3_U3268(p3_u3268), .P3_U3267(p3_u3267), .P3_U3266(p3_u3266), .P3_U3265(p3_u3265), .P3_U3264(p3_u3264), .P3_U3263(p3_u3263), .P3_U3262(p3_u3262), .P3_U3261(p3_u3261), .P3_U3260(p3_u3260), .P3_U3259(p3_u3259), .P3_U3258(p3_u3258), .P3_U3257(p3_u3257), .P3_U3256(p3_u3256), .P3_U3255(p3_u3255), .P3_U3254(p3_u3254), .P3_U3253(p3_u3253), .P3_U3252(p3_u3252), .P3_U3251(p3_u3251), .P3_U3250(p3_u3250), .P3_U3249(p3_u3249), .P3_U3248(p3_u3248), .P3_U3247(p3_u3247), .P3_U3246(p3_u3246), .P3_U3245(p3_u3245), .P3_U3244(p3_u3244), .P3_U3243(p3_u3243), .P3_U3242(p3_u3242), .P3_U3241(p3_u3241), .P3_U3557(p3_u3557), .P3_U3558(p3_u3558), .P3_U3559(p3_u3559), .P3_U3560(p3_u3560), .P3_U3561(p3_u3561), .P3_U3562(p3_u3562), .P3_U3563(p3_u3563), .P3_U3564(p3_u3564), .P3_U3565(p3_u3565), .P3_U3566(p3_u3566), .P3_U3567(p3_u3567), .P3_U3568(p3_u3568), .P3_U3569(p3_u3569), .P3_U3570(p3_u3570), .P3_U3571(p3_u3571), .P3_U3572(p3_u3572), .P3_U3573(p3_u3573), .P3_U3574(p3_u3574), .P3_U3575(p3_u3575), .P3_U3576(p3_u3576), .P3_U3577(p3_u3577), .P3_U3578(p3_u3578), .P3_U3579(p3_u3579), .P3_U3580(p3_u3580), .P3_U3581(p3_u3581), .P3_U3582(p3_u3582), .P3_U3583(p3_u3583), .P3_U3584(p3_u3584), .P3_U3585(p3_u3585), .P3_U3586(p3_u3586), .P3_U3587(p3_u3587), .P3_U3588(p3_u3588), .P3_U3240(p3_u3240), .P3_U3239(p3_u3239), .P3_U3238(p3_u3238), .P3_U3237(p3_u3237), .P3_U3236(p3_u3236), .P3_U3235(p3_u3235), .P3_U3234(p3_u3234), .P3_U3233(p3_u3233), .P3_U3232(p3_u3232), .P3_U3231(p3_u3231), .P3_U3230(p3_u3230), .P3_U3229(p3_u3229), .P3_U3228(p3_u3228), .P3_U3227(p3_u3227), .P3_U3226(p3_u3226), .P3_U3225(p3_u3225), .P3_U3224(p3_u3224), .P3_U3223(p3_u3223), .P3_U3222(p3_u3222), .P3_U3221(p3_u3221), .P3_U3220(p3_u3220), .P3_U3219(p3_u3219), .P3_U3218(p3_u3218), .P3_U3217(p3_u3217), .P3_U3216(p3_u3216), .P3_U3215(p3_u3215), .P3_U3214(p3_u3214), .P3_U3213(p3_u3213), .P3_U3212(p3_u3212), .P3_U3211(p3_u3211), .P3_U3084(p3_u3084), .P3_U3083(p3_u3083), .P3_U4038(p3_u4038), .P4_U3351(p4_u3351), .P4_U3350(p4_u3350), .P4_U3349(p4_u3349), .P4_U3348(p4_u3348), .P4_U3347(p4_u3347), .P4_U3346(p4_u3346), .P4_U3345(p4_u3345), .P4_U3344(p4_u3344), .P4_U3343(p4_u3343), .P4_U3342(p4_u3342), .P4_U3341(p4_u3341), .P4_U3340(p4_u3340), .P4_U3339(p4_u3339), .P4_U3338(p4_u3338), .P4_U3337(p4_u3337), .P4_U3336(p4_u3336), .P4_U3335(p4_u3335), .P4_U3334(p4_u3334), .P4_U3333(p4_u3333), .P4_U3332(p4_u3332), .P4_U3331(p4_u3331), .P4_U3330(p4_u3330), .P4_U3329(p4_u3329), .P4_U3328(p4_u3328), .P4_U3327(p4_u3327), .P4_U3326(p4_u3326), .P4_U3325(p4_u3325), .P4_U3324(p4_u3324), .P4_U3323(p4_u3323), .P4_U3322(p4_u3322), .P4_U3321(p4_u3321), .P4_U3320(p4_u3320), .P4_U3437(p4_u3437), .P4_U3438(p4_u3438), .P4_U3319(p4_u3319), .P4_U3318(p4_u3318), .P4_U3317(p4_u3317), .P4_U3316(p4_u3316), .P4_U3315(p4_u3315), .P4_U3314(p4_u3314), .P4_U3313(p4_u3313), .P4_U3312(p4_u3312), .P4_U3311(p4_u3311), .P4_U3310(p4_u3310), .P4_U3309(p4_u3309), .P4_U3308(p4_u3308), .P4_U3307(p4_u3307), .P4_U3306(p4_u3306), .P4_U3305(p4_u3305), .P4_U3304(p4_u3304), .P4_U3303(p4_u3303), .P4_U3302(p4_u3302), .P4_U3301(p4_u3301), .P4_U3300(p4_u3300), .P4_U3299(p4_u3299), .P4_U3298(p4_u3298), .P4_U3297(p4_u3297), .P4_U3296(p4_u3296), .P4_U3295(p4_u3295), .P4_U3294(p4_u3294), .P4_U3293(p4_u3293), .P4_U3292(p4_u3292), .P4_U3291(p4_u3291), .P4_U3290(p4_u3290), .P4_U3451(p4_u3451), .P4_U3454(p4_u3454), .P4_U3457(p4_u3457), .P4_U3460(p4_u3460), .P4_U3463(p4_u3463), .P4_U3466(p4_u3466), .P4_U3469(p4_u3469), .P4_U3472(p4_u3472), .P4_U3475(p4_u3475), .P4_U3478(p4_u3478), .P4_U3481(p4_u3481), .P4_U3484(p4_u3484), .P4_U3487(p4_u3487), .P4_U3490(p4_u3490), .P4_U3493(p4_u3493), .P4_U3496(p4_u3496), .P4_U3499(p4_u3499), .P4_U3502(p4_u3502), .P4_U3505(p4_u3505), .P4_U3507(p4_u3507), .P4_U3508(p4_u3508), .P4_U3509(p4_u3509), .P4_U3510(p4_u3510), .P4_U3511(p4_u3511), .P4_U3512(p4_u3512), .P4_U3513(p4_u3513), .P4_U3514(p4_u3514), .P4_U3515(p4_u3515), .P4_U3516(p4_u3516), .P4_U3517(p4_u3517), .P4_U3518(p4_u3518), .P4_U3519(p4_u3519), .P4_U3520(p4_u3520), .P4_U3521(p4_u3521), .P4_U3522(p4_u3522), .P4_U3523(p4_u3523), .P4_U3524(p4_u3524), .P4_U3525(p4_u3525), .P4_U3526(p4_u3526), .P4_U3527(p4_u3527), .P4_U3528(p4_u3528), .P4_U3529(p4_u3529), .P4_U3530(p4_u3530), .P4_U3531(p4_u3531), .P4_U3532(p4_u3532), .P4_U3533(p4_u3533), .P4_U3534(p4_u3534), .P4_U3535(p4_u3535), .P4_U3536(p4_u3536), .P4_U3537(p4_u3537), .P4_U3538(p4_u3538), .P4_U3539(p4_u3539), .P4_U3540(p4_u3540), .P4_U3541(p4_u3541), .P4_U3542(p4_u3542), .P4_U3543(p4_u3543), .P4_U3544(p4_u3544), .P4_U3545(p4_u3545), .P4_U3546(p4_u3546), .P4_U3547(p4_u3547), .P4_U3548(p4_u3548), .P4_U3549(p4_u3549), .P4_U3550(p4_u3550), .P4_U3551(p4_u3551), .P4_U3289(p4_u3289), .P4_U3288(p4_u3288), .P4_U3287(p4_u3287), .P4_U3286(p4_u3286), .P4_U3285(p4_u3285), .P4_U3284(p4_u3284), .P4_U3283(p4_u3283), .P4_U3282(p4_u3282), .P4_U3281(p4_u3281), .P4_U3280(p4_u3280), .P4_U3279(p4_u3279), .P4_U3278(p4_u3278), .P4_U3277(p4_u3277), .P4_U3276(p4_u3276), .P4_U3275(p4_u3275), .P4_U3274(p4_u3274), .P4_U3273(p4_u3273), .P4_U3272(p4_u3272), .P4_U3271(p4_u3271), .P4_U3270(p4_u3270), .P4_U3269(p4_u3269), .P4_U3268(p4_u3268), .P4_U3267(p4_u3267), .P4_U3266(p4_u3266), .P4_U3265(p4_u3265), .P4_U3264(p4_u3264), .P4_U3263(p4_u3263), .P4_U3262(p4_u3262), .P4_U3261(p4_u3261), .P4_U3260(p4_u3260), .P4_U3259(p4_u3259), .P4_U3258(p4_u3258), .P4_U3257(p4_u3257), .P4_U3256(p4_u3256), .P4_U3255(p4_u3255), .P4_U3254(p4_u3254), .P4_U3253(p4_u3253), .P4_U3252(p4_u3252), .P4_U3251(p4_u3251), .P4_U3250(p4_u3250), .P4_U3249(p4_u3249), .P4_U3248(p4_u3248), .P4_U3247(p4_u3247), .P4_U3246(p4_u3246), .P4_U3245(p4_u3245), .P4_U3244(p4_u3244), .P4_U3243(p4_u3243), .P4_U3242(p4_u3242), .P4_U3241(p4_u3241), .P4_U3240(p4_u3240), .P4_U3239(p4_u3239), .P4_U3238(p4_u3238), .P4_U3552(p4_u3552), .P4_U3553(p4_u3553), .P4_U3554(p4_u3554), .P4_U3555(p4_u3555), .P4_U3556(p4_u3556), .P4_U3557(p4_u3557), .P4_U3558(p4_u3558), .P4_U3559(p4_u3559), .P4_U3560(p4_u3560), .P4_U3561(p4_u3561), .P4_U3562(p4_u3562), .P4_U3563(p4_u3563), .P4_U3564(p4_u3564), .P4_U3565(p4_u3565), .P4_U3566(p4_u3566), .P4_U3567(p4_u3567), .P4_U3568(p4_u3568), .P4_U3569(p4_u3569), .P4_U3570(p4_u3570), .P4_U3571(p4_u3571), .P4_U3572(p4_u3572), .P4_U3573(p4_u3573), .P4_U3574(p4_u3574), .P4_U3575(p4_u3575), .P4_U3576(p4_u3576), .P4_U3577(p4_u3577), .P4_U3578(p4_u3578), .P4_U3579(p4_u3579), .P4_U3580(p4_u3580), .P4_U3581(p4_u3581), .P4_U3582(p4_u3582), .P4_U3583(p4_u3583), .P4_U3237(p4_u3237), .P4_U3236(p4_u3236), .P4_U3235(p4_u3235), .P4_U3234(p4_u3234), .P4_U3233(p4_u3233), .P4_U3232(p4_u3232), .P4_U3231(p4_u3231), .P4_U3230(p4_u3230), .P4_U3229(p4_u3229), .P4_U3228(p4_u3228), .P4_U3227(p4_u3227), .P4_U3226(p4_u3226), .P4_U3225(p4_u3225), .P4_U3224(p4_u3224), .P4_U3223(p4_u3223), .P4_U3222(p4_u3222), .P4_U3221(p4_u3221), .P4_U3220(p4_u3220), .P4_U3219(p4_u3219), .P4_U3218(p4_u3218), .P4_U3217(p4_u3217), .P4_U3216(p4_u3216), .P4_U3215(p4_u3215), .P4_U3214(p4_u3214), .P4_U3213(p4_u3213), .P4_U3212(p4_u3212), .P4_U3211(p4_u3211), .P4_U3210(p4_u3210), .P4_U3209(p4_u3209), .P4_U3208(p4_u3208), .P4_U3147(p4_u3147), .P4_U3146(p4_u3146), .P4_U4028(p4_u4028), .P1_P3_U3274(p1_p3_u3274), .P1_P3_U3275(p1_p3_u3275), .P1_P3_U3276(p1_p3_u3276), .P1_P3_U3277(p1_p3_u3277), .P1_P3_U3061(p1_p3_u3061), .P1_P3_U3060(p1_p3_u3060), .P1_P3_U3059(p1_p3_u3059), .P1_P3_U3058(p1_p3_u3058), .P1_P3_U3057(p1_p3_u3057), .P1_P3_U3056(p1_p3_u3056), .P1_P3_U3055(p1_p3_u3055), .P1_P3_U3054(p1_p3_u3054), .P1_P3_U3053(p1_p3_u3053), .P1_P3_U3052(p1_p3_u3052), .P1_P3_U3051(p1_p3_u3051), .P1_P3_U3050(p1_p3_u3050), .P1_P3_U3049(p1_p3_u3049), .P1_P3_U3048(p1_p3_u3048), .P1_P3_U3047(p1_p3_u3047), .P1_P3_U3046(p1_p3_u3046), .P1_P3_U3045(p1_p3_u3045), .P1_P3_U3044(p1_p3_u3044), .P1_P3_U3043(p1_p3_u3043), .P1_P3_U3042(p1_p3_u3042), .P1_P3_U3041(p1_p3_u3041), .P1_P3_U3040(p1_p3_u3040), .P1_P3_U3039(p1_p3_u3039), .P1_P3_U3038(p1_p3_u3038), .P1_P3_U3037(p1_p3_u3037), .P1_P3_U3036(p1_p3_u3036), .P1_P3_U3035(p1_p3_u3035), .P1_P3_U3034(p1_p3_u3034), .P1_P3_U3033(p1_p3_u3033), .P1_P3_U3032(p1_p3_u3032), .P1_P3_U3031(p1_p3_u3031), .P1_P3_U3030(p1_p3_u3030), .P1_P3_U3029(p1_p3_u3029), .P1_P3_U3280(p1_p3_u3280), .P1_P3_U3281(p1_p3_u3281), .P1_P3_U3028(p1_p3_u3028), .P1_P3_U3027(p1_p3_u3027), .P1_P3_U3026(p1_p3_u3026), .P1_P3_U3025(p1_p3_u3025), .P1_P3_U3024(p1_p3_u3024), .P1_P3_U3023(p1_p3_u3023), .P1_P3_U3022(p1_p3_u3022), .P1_P3_U3021(p1_p3_u3021), .P1_P3_U3020(p1_p3_u3020), .P1_P3_U3019(p1_p3_u3019), .P1_P3_U3018(p1_p3_u3018), .P1_P3_U3017(p1_p3_u3017), .P1_P3_U3016(p1_p3_u3016), .P1_P3_U3015(p1_p3_u3015), .P1_P3_U3014(p1_p3_u3014), .P1_P3_U3013(p1_p3_u3013), .P1_P3_U3012(p1_p3_u3012), .P1_P3_U3011(p1_p3_u3011), .P1_P3_U3010(p1_p3_u3010), .P1_P3_U3009(p1_p3_u3009), .P1_P3_U3008(p1_p3_u3008), .P1_P3_U3007(p1_p3_u3007), .P1_P3_U3006(p1_p3_u3006), .P1_P3_U3005(p1_p3_u3005), .P1_P3_U3004(p1_p3_u3004), .P1_P3_U3003(p1_p3_u3003), .P1_P3_U3002(p1_p3_u3002), .P1_P3_U3001(p1_p3_u3001), .P1_P3_U3000(p1_p3_u3000), .P1_P3_U2999(p1_p3_u2999), .P1_P3_U3282(p1_p3_u3282), .P1_P3_U2998(p1_p3_u2998), .P1_P3_U2997(p1_p3_u2997), .P1_P3_U2996(p1_p3_u2996), .P1_P3_U2995(p1_p3_u2995), .P1_P3_U2994(p1_p3_u2994), .P1_P3_U2993(p1_p3_u2993), .P1_P3_U2992(p1_p3_u2992), .P1_P3_U2991(p1_p3_u2991), .P1_P3_U2990(p1_p3_u2990), .P1_P3_U2989(p1_p3_u2989), .P1_P3_U2988(p1_p3_u2988), .P1_P3_U2987(p1_p3_u2987), .P1_P3_U2986(p1_p3_u2986), .P1_P3_U2985(p1_p3_u2985), .P1_P3_U2984(p1_p3_u2984), .P1_P3_U2983(p1_p3_u2983), .P1_P3_U2982(p1_p3_u2982), .P1_P3_U2981(p1_p3_u2981), .P1_P3_U2980(p1_p3_u2980), .P1_P3_U2979(p1_p3_u2979), .P1_P3_U2978(p1_p3_u2978), .P1_P3_U2977(p1_p3_u2977), .P1_P3_U2976(p1_p3_u2976), .P1_P3_U2975(p1_p3_u2975), .P1_P3_U2974(p1_p3_u2974), .P1_P3_U2973(p1_p3_u2973), .P1_P3_U2972(p1_p3_u2972), .P1_P3_U2971(p1_p3_u2971), .P1_P3_U2970(p1_p3_u2970), .P1_P3_U2969(p1_p3_u2969), .P1_P3_U2968(p1_p3_u2968), .P1_P3_U2967(p1_p3_u2967), .P1_P3_U2966(p1_p3_u2966), .P1_P3_U2965(p1_p3_u2965), .P1_P3_U2964(p1_p3_u2964), .P1_P3_U2963(p1_p3_u2963), .P1_P3_U2962(p1_p3_u2962), .P1_P3_U2961(p1_p3_u2961), .P1_P3_U2960(p1_p3_u2960), .P1_P3_U2959(p1_p3_u2959), .P1_P3_U2958(p1_p3_u2958), .P1_P3_U2957(p1_p3_u2957), .P1_P3_U2956(p1_p3_u2956), .P1_P3_U2955(p1_p3_u2955), .P1_P3_U2954(p1_p3_u2954), .P1_P3_U2953(p1_p3_u2953), .P1_P3_U2952(p1_p3_u2952), .P1_P3_U2951(p1_p3_u2951), .P1_P3_U2950(p1_p3_u2950), .P1_P3_U2949(p1_p3_u2949), .P1_P3_U2948(p1_p3_u2948), .P1_P3_U2947(p1_p3_u2947), .P1_P3_U2946(p1_p3_u2946), .P1_P3_U2945(p1_p3_u2945), .P1_P3_U2944(p1_p3_u2944), .P1_P3_U2943(p1_p3_u2943), .P1_P3_U2942(p1_p3_u2942), .P1_P3_U2941(p1_p3_u2941), .P1_P3_U2940(p1_p3_u2940), .P1_P3_U2939(p1_p3_u2939), .P1_P3_U2938(p1_p3_u2938), .P1_P3_U2937(p1_p3_u2937), .P1_P3_U2936(p1_p3_u2936), .P1_P3_U2935(p1_p3_u2935), .P1_P3_U2934(p1_p3_u2934), .P1_P3_U2933(p1_p3_u2933), .P1_P3_U2932(p1_p3_u2932), .P1_P3_U2931(p1_p3_u2931), .P1_P3_U2930(p1_p3_u2930), .P1_P3_U2929(p1_p3_u2929), .P1_P3_U2928(p1_p3_u2928), .P1_P3_U2927(p1_p3_u2927), .P1_P3_U2926(p1_p3_u2926), .P1_P3_U2925(p1_p3_u2925), .P1_P3_U2924(p1_p3_u2924), .P1_P3_U2923(p1_p3_u2923), .P1_P3_U2922(p1_p3_u2922), .P1_P3_U2921(p1_p3_u2921), .P1_P3_U2920(p1_p3_u2920), .P1_P3_U2919(p1_p3_u2919), .P1_P3_U2918(p1_p3_u2918), .P1_P3_U2917(p1_p3_u2917), .P1_P3_U2916(p1_p3_u2916), .P1_P3_U2915(p1_p3_u2915), .P1_P3_U2914(p1_p3_u2914), .P1_P3_U2913(p1_p3_u2913), .P1_P3_U2912(p1_p3_u2912), .P1_P3_U2911(p1_p3_u2911), .P1_P3_U2910(p1_p3_u2910), .P1_P3_U2909(p1_p3_u2909), .P1_P3_U2908(p1_p3_u2908), .P1_P3_U2907(p1_p3_u2907), .P1_P3_U2906(p1_p3_u2906), .P1_P3_U2905(p1_p3_u2905), .P1_P3_U2904(p1_p3_u2904), .P1_P3_U2903(p1_p3_u2903), .P1_P3_U2902(p1_p3_u2902), .P1_P3_U2901(p1_p3_u2901), .P1_P3_U2900(p1_p3_u2900), .P1_P3_U2899(p1_p3_u2899), .P1_P3_U2898(p1_p3_u2898), .P1_P3_U2897(p1_p3_u2897), .P1_P3_U2896(p1_p3_u2896), .P1_P3_U2895(p1_p3_u2895), .P1_P3_U2894(p1_p3_u2894), .P1_P3_U2893(p1_p3_u2893), .P1_P3_U2892(p1_p3_u2892), .P1_P3_U2891(p1_p3_u2891), .P1_P3_U2890(p1_p3_u2890), .P1_P3_U2889(p1_p3_u2889), .P1_P3_U2888(p1_p3_u2888), .P1_P3_U2887(p1_p3_u2887), .P1_P3_U2886(p1_p3_u2886), .P1_P3_U2885(p1_p3_u2885), .P1_P3_U2884(p1_p3_u2884), .P1_P3_U2883(p1_p3_u2883), .P1_P3_U2882(p1_p3_u2882), .P1_P3_U2881(p1_p3_u2881), .P1_P3_U2880(p1_p3_u2880), .P1_P3_U2879(p1_p3_u2879), .P1_P3_U2878(p1_p3_u2878), .P1_P3_U2877(p1_p3_u2877), .P1_P3_U2876(p1_p3_u2876), .P1_P3_U2875(p1_p3_u2875), .P1_P3_U2874(p1_p3_u2874), .P1_P3_U2873(p1_p3_u2873), .P1_P3_U2872(p1_p3_u2872), .P1_P3_U2871(p1_p3_u2871), .P1_P3_U2870(p1_p3_u2870), .P1_P3_U2869(p1_p3_u2869), .P1_P3_U2868(p1_p3_u2868), .P1_P3_U3284(p1_p3_u3284), .P1_P3_U3285(p1_p3_u3285), .P1_P3_U3288(p1_p3_u3288), .P1_P3_U3289(p1_p3_u3289), .P1_P3_U3290(p1_p3_u3290), .P1_P3_U2867(p1_p3_u2867), .P1_P3_U2866(p1_p3_u2866), .P1_P3_U2865(p1_p3_u2865), .P1_P3_U2864(p1_p3_u2864), .P1_P3_U2863(p1_p3_u2863), .P1_P3_U2862(p1_p3_u2862), .P1_P3_U2861(p1_p3_u2861), .P1_P3_U2860(p1_p3_u2860), .P1_P3_U2859(p1_p3_u2859), .P1_P3_U2858(p1_p3_u2858), .P1_P3_U2857(p1_p3_u2857), .P1_P3_U2856(p1_p3_u2856), .P1_P3_U2855(p1_p3_u2855), .P1_P3_U2854(p1_p3_u2854), .P1_P3_U2853(p1_p3_u2853), .P1_P3_U2852(p1_p3_u2852), .P1_P3_U2851(p1_p3_u2851), .P1_P3_U2850(p1_p3_u2850), .P1_P3_U2849(p1_p3_u2849), .P1_P3_U2848(p1_p3_u2848), .P1_P3_U2847(p1_p3_u2847), .P1_P3_U2846(p1_p3_u2846), .P1_P3_U2845(p1_p3_u2845), .P1_P3_U2844(p1_p3_u2844), .P1_P3_U2843(p1_p3_u2843), .P1_P3_U2842(p1_p3_u2842), .P1_P3_U2841(p1_p3_u2841), .P1_P3_U2840(p1_p3_u2840), .P1_P3_U2839(p1_p3_u2839), .P1_P3_U2838(p1_p3_u2838), .P1_P3_U2837(p1_p3_u2837), .P1_P3_U2836(p1_p3_u2836), .P1_P3_U2835(p1_p3_u2835), .P1_P3_U2834(p1_p3_u2834), .P1_P3_U2833(p1_p3_u2833), .P1_P3_U2832(p1_p3_u2832), .P1_P3_U2831(p1_p3_u2831), .P1_P3_U2830(p1_p3_u2830), .P1_P3_U2829(p1_p3_u2829), .P1_P3_U2828(p1_p3_u2828), .P1_P3_U2827(p1_p3_u2827), .P1_P3_U2826(p1_p3_u2826), .P1_P3_U2825(p1_p3_u2825), .P1_P3_U2824(p1_p3_u2824), .P1_P3_U2823(p1_p3_u2823), .P1_P3_U2822(p1_p3_u2822), .P1_P3_U2821(p1_p3_u2821), .P1_P3_U2820(p1_p3_u2820), .P1_P3_U2819(p1_p3_u2819), .P1_P3_U2818(p1_p3_u2818), .P1_P3_U2817(p1_p3_u2817), .P1_P3_U2816(p1_p3_u2816), .P1_P3_U2815(p1_p3_u2815), .P1_P3_U2814(p1_p3_u2814), .P1_P3_U2813(p1_p3_u2813), .P1_P3_U2812(p1_p3_u2812), .P1_P3_U2811(p1_p3_u2811), .P1_P3_U2810(p1_p3_u2810), .P1_P3_U2809(p1_p3_u2809), .P1_P3_U2808(p1_p3_u2808), .P1_P3_U2807(p1_p3_u2807), .P1_P3_U2806(p1_p3_u2806), .P1_P3_U2805(p1_p3_u2805), .P1_P3_U2804(p1_p3_u2804), .P1_P3_U2803(p1_p3_u2803), .P1_P3_U2802(p1_p3_u2802), .P1_P3_U2801(p1_p3_u2801), .P1_P3_U2800(p1_p3_u2800), .P1_P3_U2799(p1_p3_u2799), .P1_P3_U2798(p1_p3_u2798), .P1_P3_U2797(p1_p3_u2797), .P1_P3_U2796(p1_p3_u2796), .P1_P3_U2795(p1_p3_u2795), .P1_P3_U2794(p1_p3_u2794), .P1_P3_U2793(p1_p3_u2793), .P1_P3_U2792(p1_p3_u2792), .P1_P3_U2791(p1_p3_u2791), .P1_P3_U2790(p1_p3_u2790), .P1_P3_U2789(p1_p3_u2789), .P1_P3_U2788(p1_p3_u2788), .P1_P3_U2787(p1_p3_u2787), .P1_P3_U2786(p1_p3_u2786), .P1_P3_U2785(p1_p3_u2785), .P1_P3_U2784(p1_p3_u2784), .P1_P3_U2783(p1_p3_u2783), .P1_P3_U2782(p1_p3_u2782), .P1_P3_U2781(p1_p3_u2781), .P1_P3_U2780(p1_p3_u2780), .P1_P3_U2779(p1_p3_u2779), .P1_P3_U2778(p1_p3_u2778), .P1_P3_U2777(p1_p3_u2777), .P1_P3_U2776(p1_p3_u2776), .P1_P3_U2775(p1_p3_u2775), .P1_P3_U2774(p1_p3_u2774), .P1_P3_U2773(p1_p3_u2773), .P1_P3_U2772(p1_p3_u2772), .P1_P3_U2771(p1_p3_u2771), .P1_P3_U2770(p1_p3_u2770), .P1_P3_U2769(p1_p3_u2769), .P1_P3_U2768(p1_p3_u2768), .P1_P3_U2767(p1_p3_u2767), .P1_P3_U2766(p1_p3_u2766), .P1_P3_U2765(p1_p3_u2765), .P1_P3_U2764(p1_p3_u2764), .P1_P3_U2763(p1_p3_u2763), .P1_P3_U2762(p1_p3_u2762), .P1_P3_U2761(p1_p3_u2761), .P1_P3_U2760(p1_p3_u2760), .P1_P3_U2759(p1_p3_u2759), .P1_P3_U2758(p1_p3_u2758), .P1_P3_U2757(p1_p3_u2757), .P1_P3_U2756(p1_p3_u2756), .P1_P3_U2755(p1_p3_u2755), .P1_P3_U2754(p1_p3_u2754), .P1_P3_U2753(p1_p3_u2753), .P1_P3_U2752(p1_p3_u2752), .P1_P3_U2751(p1_p3_u2751), .P1_P3_U2750(p1_p3_u2750), .P1_P3_U2749(p1_p3_u2749), .P1_P3_U2748(p1_p3_u2748), .P1_P3_U2747(p1_p3_u2747), .P1_P3_U2746(p1_p3_u2746), .P1_P3_U2745(p1_p3_u2745), .P1_P3_U2744(p1_p3_u2744), .P1_P3_U2743(p1_p3_u2743), .P1_P3_U2742(p1_p3_u2742), .P1_P3_U2741(p1_p3_u2741), .P1_P3_U2740(p1_p3_u2740), .P1_P3_U2739(p1_p3_u2739), .P1_P3_U2738(p1_p3_u2738), .P1_P3_U2737(p1_p3_u2737), .P1_P3_U2736(p1_p3_u2736), .P1_P3_U2735(p1_p3_u2735), .P1_P3_U2734(p1_p3_u2734), .P1_P3_U2733(p1_p3_u2733), .P1_P3_U2732(p1_p3_u2732), .P1_P3_U2731(p1_p3_u2731), .P1_P3_U2730(p1_p3_u2730), .P1_P3_U2729(p1_p3_u2729), .P1_P3_U2728(p1_p3_u2728), .P1_P3_U2727(p1_p3_u2727), .P1_P3_U2726(p1_p3_u2726), .P1_P3_U2725(p1_p3_u2725), .P1_P3_U2724(p1_p3_u2724), .P1_P3_U2723(p1_p3_u2723), .P1_P3_U2722(p1_p3_u2722), .P1_P3_U2721(p1_p3_u2721), .P1_P3_U2720(p1_p3_u2720), .P1_P3_U2719(p1_p3_u2719), .P1_P3_U2718(p1_p3_u2718), .P1_P3_U2717(p1_p3_u2717), .P1_P3_U2716(p1_p3_u2716), .P1_P3_U2715(p1_p3_u2715), .P1_P3_U2714(p1_p3_u2714), .P1_P3_U2713(p1_p3_u2713), .P1_P3_U2712(p1_p3_u2712), .P1_P3_U2711(p1_p3_u2711), .P1_P3_U2710(p1_p3_u2710), .P1_P3_U2709(p1_p3_u2709), .P1_P3_U2708(p1_p3_u2708), .P1_P3_U2707(p1_p3_u2707), .P1_P3_U2706(p1_p3_u2706), .P1_P3_U2705(p1_p3_u2705), .P1_P3_U2704(p1_p3_u2704), .P1_P3_U2703(p1_p3_u2703), .P1_P3_U2702(p1_p3_u2702), .P1_P3_U2701(p1_p3_u2701), .P1_P3_U2700(p1_p3_u2700), .P1_P3_U2699(p1_p3_u2699), .P1_P3_U2698(p1_p3_u2698), .P1_P3_U2697(p1_p3_u2697), .P1_P3_U2696(p1_p3_u2696), .P1_P3_U2695(p1_p3_u2695), .P1_P3_U2694(p1_p3_u2694), .P1_P3_U2693(p1_p3_u2693), .P1_P3_U2692(p1_p3_u2692), .P1_P3_U2691(p1_p3_u2691), .P1_P3_U2690(p1_p3_u2690), .P1_P3_U2689(p1_p3_u2689), .P1_P3_U2688(p1_p3_u2688), .P1_P3_U2687(p1_p3_u2687), .P1_P3_U2686(p1_p3_u2686), .P1_P3_U2685(p1_p3_u2685), .P1_P3_U2684(p1_p3_u2684), .P1_P3_U2683(p1_p3_u2683), .P1_P3_U2682(p1_p3_u2682), .P1_P3_U2681(p1_p3_u2681), .P1_P3_U2680(p1_p3_u2680), .P1_P3_U2679(p1_p3_u2679), .P1_P3_U2678(p1_p3_u2678), .P1_P3_U2677(p1_p3_u2677), .P1_P3_U2676(p1_p3_u2676), .P1_P3_U2675(p1_p3_u2675), .P1_P3_U2674(p1_p3_u2674), .P1_P3_U2673(p1_p3_u2673), .P1_P3_U2672(p1_p3_u2672), .P1_P3_U2671(p1_p3_u2671), .P1_P3_U2670(p1_p3_u2670), .P1_P3_U2669(p1_p3_u2669), .P1_P3_U2668(p1_p3_u2668), .P1_P3_U2667(p1_p3_u2667), .P1_P3_U2666(p1_p3_u2666), .P1_P3_U2665(p1_p3_u2665), .P1_P3_U2664(p1_p3_u2664), .P1_P3_U2663(p1_p3_u2663), .P1_P3_U2662(p1_p3_u2662), .P1_P3_U2661(p1_p3_u2661), .P1_P3_U2660(p1_p3_u2660), .P1_P3_U2659(p1_p3_u2659), .P1_P3_U2658(p1_p3_u2658), .P1_P3_U2657(p1_p3_u2657), .P1_P3_U2656(p1_p3_u2656), .P1_P3_U2655(p1_p3_u2655), .P1_P3_U2654(p1_p3_u2654), .P1_P3_U2653(p1_p3_u2653), .P1_P3_U2652(p1_p3_u2652), .P1_P3_U2651(p1_p3_u2651), .P1_P3_U2650(p1_p3_u2650), .P1_P3_U2649(p1_p3_u2649), .P1_P3_U2648(p1_p3_u2648), .P1_P3_U2647(p1_p3_u2647), .P1_P3_U2646(p1_p3_u2646), .P1_P3_U2645(p1_p3_u2645), .P1_P3_U2644(p1_p3_u2644), .P1_P3_U2643(p1_p3_u2643), .P1_P3_U2642(p1_p3_u2642), .P1_P3_U2641(p1_p3_u2641), .P1_P3_U2640(p1_p3_u2640), .P1_P3_U2639(p1_p3_u2639), .P1_P3_U3292(p1_p3_u3292), .P1_P3_U2638(p1_p3_u2638), .P1_P3_U3293(p1_p3_u3293), .P1_P3_U3294(p1_p3_u3294), .P1_P3_U2637(p1_p3_u2637), .P1_P3_U3295(p1_p3_u3295), .P1_P3_U2636(p1_p3_u2636), .P1_P3_U3296(p1_p3_u3296), .P1_P3_U2635(p1_p3_u2635), .P1_P3_U3297(p1_p3_u3297), .P1_P3_U2634(p1_p3_u2634), .P1_P3_U2633(p1_p3_u2633), .P1_P3_U3298(p1_p3_u3298), .P1_P3_U3299(p1_p3_u3299), .P1_P2_U3274(p1_p2_u3274), .P1_P2_U3275(p1_p2_u3275), .P1_P2_U3276(p1_p2_u3276), .P1_P2_U3277(p1_p2_u3277), .P1_P2_U3061(p1_p2_u3061), .P1_P2_U3060(p1_p2_u3060), .P1_P2_U3059(p1_p2_u3059), .P1_P2_U3058(p1_p2_u3058), .P1_P2_U3057(p1_p2_u3057), .P1_P2_U3056(p1_p2_u3056), .P1_P2_U3055(p1_p2_u3055), .P1_P2_U3054(p1_p2_u3054), .P1_P2_U3053(p1_p2_u3053), .P1_P2_U3052(p1_p2_u3052), .P1_P2_U3051(p1_p2_u3051), .P1_P2_U3050(p1_p2_u3050), .P1_P2_U3049(p1_p2_u3049), .P1_P2_U3048(p1_p2_u3048), .P1_P2_U3047(p1_p2_u3047), .P1_P2_U3046(p1_p2_u3046), .P1_P2_U3045(p1_p2_u3045), .P1_P2_U3044(p1_p2_u3044), .P1_P2_U3043(p1_p2_u3043), .P1_P2_U3042(p1_p2_u3042), .P1_P2_U3041(p1_p2_u3041), .P1_P2_U3040(p1_p2_u3040), .P1_P2_U3039(p1_p2_u3039), .P1_P2_U3038(p1_p2_u3038), .P1_P2_U3037(p1_p2_u3037), .P1_P2_U3036(p1_p2_u3036), .P1_P2_U3035(p1_p2_u3035), .P1_P2_U3034(p1_p2_u3034), .P1_P2_U3033(p1_p2_u3033), .P1_P2_U3032(p1_p2_u3032), .P1_P2_U3031(p1_p2_u3031), .P1_P2_U3030(p1_p2_u3030), .P1_P2_U3029(p1_p2_u3029), .P1_P2_U3280(p1_p2_u3280), .P1_P2_U3281(p1_p2_u3281), .P1_P2_U3028(p1_p2_u3028), .P1_P2_U3027(p1_p2_u3027), .P1_P2_U3026(p1_p2_u3026), .P1_P2_U3025(p1_p2_u3025), .P1_P2_U3024(p1_p2_u3024), .P1_P2_U3023(p1_p2_u3023), .P1_P2_U3022(p1_p2_u3022), .P1_P2_U3021(p1_p2_u3021), .P1_P2_U3020(p1_p2_u3020), .P1_P2_U3019(p1_p2_u3019), .P1_P2_U3018(p1_p2_u3018), .P1_P2_U3017(p1_p2_u3017), .P1_P2_U3016(p1_p2_u3016), .P1_P2_U3015(p1_p2_u3015), .P1_P2_U3014(p1_p2_u3014), .P1_P2_U3013(p1_p2_u3013), .P1_P2_U3012(p1_p2_u3012), .P1_P2_U3011(p1_p2_u3011), .P1_P2_U3010(p1_p2_u3010), .P1_P2_U3009(p1_p2_u3009), .P1_P2_U3008(p1_p2_u3008), .P1_P2_U3007(p1_p2_u3007), .P1_P2_U3006(p1_p2_u3006), .P1_P2_U3005(p1_p2_u3005), .P1_P2_U3004(p1_p2_u3004), .P1_P2_U3003(p1_p2_u3003), .P1_P2_U3002(p1_p2_u3002), .P1_P2_U3001(p1_p2_u3001), .P1_P2_U3000(p1_p2_u3000), .P1_P2_U2999(p1_p2_u2999), .P1_P2_U3282(p1_p2_u3282), .P1_P2_U2998(p1_p2_u2998), .P1_P2_U2997(p1_p2_u2997), .P1_P2_U2996(p1_p2_u2996), .P1_P2_U2995(p1_p2_u2995), .P1_P2_U2994(p1_p2_u2994), .P1_P2_U2993(p1_p2_u2993), .P1_P2_U2992(p1_p2_u2992), .P1_P2_U2991(p1_p2_u2991), .P1_P2_U2990(p1_p2_u2990), .P1_P2_U2989(p1_p2_u2989), .P1_P2_U2988(p1_p2_u2988), .P1_P2_U2987(p1_p2_u2987), .P1_P2_U2986(p1_p2_u2986), .P1_P2_U2985(p1_p2_u2985), .P1_P2_U2984(p1_p2_u2984), .P1_P2_U2983(p1_p2_u2983), .P1_P2_U2982(p1_p2_u2982), .P1_P2_U2981(p1_p2_u2981), .P1_P2_U2980(p1_p2_u2980), .P1_P2_U2979(p1_p2_u2979), .P1_P2_U2978(p1_p2_u2978), .P1_P2_U2977(p1_p2_u2977), .P1_P2_U2976(p1_p2_u2976), .P1_P2_U2975(p1_p2_u2975), .P1_P2_U2974(p1_p2_u2974), .P1_P2_U2973(p1_p2_u2973), .P1_P2_U2972(p1_p2_u2972), .P1_P2_U2971(p1_p2_u2971), .P1_P2_U2970(p1_p2_u2970), .P1_P2_U2969(p1_p2_u2969), .P1_P2_U2968(p1_p2_u2968), .P1_P2_U2967(p1_p2_u2967), .P1_P2_U2966(p1_p2_u2966), .P1_P2_U2965(p1_p2_u2965), .P1_P2_U2964(p1_p2_u2964), .P1_P2_U2963(p1_p2_u2963), .P1_P2_U2962(p1_p2_u2962), .P1_P2_U2961(p1_p2_u2961), .P1_P2_U2960(p1_p2_u2960), .P1_P2_U2959(p1_p2_u2959), .P1_P2_U2958(p1_p2_u2958), .P1_P2_U2957(p1_p2_u2957), .P1_P2_U2956(p1_p2_u2956), .P1_P2_U2955(p1_p2_u2955), .P1_P2_U2954(p1_p2_u2954), .P1_P2_U2953(p1_p2_u2953), .P1_P2_U2952(p1_p2_u2952), .P1_P2_U2951(p1_p2_u2951), .P1_P2_U2950(p1_p2_u2950), .P1_P2_U2949(p1_p2_u2949), .P1_P2_U2948(p1_p2_u2948), .P1_P2_U2947(p1_p2_u2947), .P1_P2_U2946(p1_p2_u2946), .P1_P2_U2945(p1_p2_u2945), .P1_P2_U2944(p1_p2_u2944), .P1_P2_U2943(p1_p2_u2943), .P1_P2_U2942(p1_p2_u2942), .P1_P2_U2941(p1_p2_u2941), .P1_P2_U2940(p1_p2_u2940), .P1_P2_U2939(p1_p2_u2939), .P1_P2_U2938(p1_p2_u2938), .P1_P2_U2937(p1_p2_u2937), .P1_P2_U2936(p1_p2_u2936), .P1_P2_U2935(p1_p2_u2935), .P1_P2_U2934(p1_p2_u2934), .P1_P2_U2933(p1_p2_u2933), .P1_P2_U2932(p1_p2_u2932), .P1_P2_U2931(p1_p2_u2931), .P1_P2_U2930(p1_p2_u2930), .P1_P2_U2929(p1_p2_u2929), .P1_P2_U2928(p1_p2_u2928), .P1_P2_U2927(p1_p2_u2927), .P1_P2_U2926(p1_p2_u2926), .P1_P2_U2925(p1_p2_u2925), .P1_P2_U2924(p1_p2_u2924), .P1_P2_U2923(p1_p2_u2923), .P1_P2_U2922(p1_p2_u2922), .P1_P2_U2921(p1_p2_u2921), .P1_P2_U2920(p1_p2_u2920), .P1_P2_U2919(p1_p2_u2919), .P1_P2_U2918(p1_p2_u2918), .P1_P2_U2917(p1_p2_u2917), .P1_P2_U2916(p1_p2_u2916), .P1_P2_U2915(p1_p2_u2915), .P1_P2_U2914(p1_p2_u2914), .P1_P2_U2913(p1_p2_u2913), .P1_P2_U2912(p1_p2_u2912), .P1_P2_U2911(p1_p2_u2911), .P1_P2_U2910(p1_p2_u2910), .P1_P2_U2909(p1_p2_u2909), .P1_P2_U2908(p1_p2_u2908), .P1_P2_U2907(p1_p2_u2907), .P1_P2_U2906(p1_p2_u2906), .P1_P2_U2905(p1_p2_u2905), .P1_P2_U2904(p1_p2_u2904), .P1_P2_U2903(p1_p2_u2903), .P1_P2_U2902(p1_p2_u2902), .P1_P2_U2901(p1_p2_u2901), .P1_P2_U2900(p1_p2_u2900), .P1_P2_U2899(p1_p2_u2899), .P1_P2_U2898(p1_p2_u2898), .P1_P2_U2897(p1_p2_u2897), .P1_P2_U2896(p1_p2_u2896), .P1_P2_U2895(p1_p2_u2895), .P1_P2_U2894(p1_p2_u2894), .P1_P2_U2893(p1_p2_u2893), .P1_P2_U2892(p1_p2_u2892), .P1_P2_U2891(p1_p2_u2891), .P1_P2_U2890(p1_p2_u2890), .P1_P2_U2889(p1_p2_u2889), .P1_P2_U2888(p1_p2_u2888), .P1_P2_U2887(p1_p2_u2887), .P1_P2_U2886(p1_p2_u2886), .P1_P2_U2885(p1_p2_u2885), .P1_P2_U2884(p1_p2_u2884), .P1_P2_U2883(p1_p2_u2883), .P1_P2_U2882(p1_p2_u2882), .P1_P2_U2881(p1_p2_u2881), .P1_P2_U2880(p1_p2_u2880), .P1_P2_U2879(p1_p2_u2879), .P1_P2_U2878(p1_p2_u2878), .P1_P2_U2877(p1_p2_u2877), .P1_P2_U2876(p1_p2_u2876), .P1_P2_U2875(p1_p2_u2875), .P1_P2_U2874(p1_p2_u2874), .P1_P2_U2873(p1_p2_u2873), .P1_P2_U2872(p1_p2_u2872), .P1_P2_U2871(p1_p2_u2871), .P1_P2_U2870(p1_p2_u2870), .P1_P2_U2869(p1_p2_u2869), .P1_P2_U2868(p1_p2_u2868), .P1_P2_U3284(p1_p2_u3284), .P1_P2_U3285(p1_p2_u3285), .P1_P2_U3288(p1_p2_u3288), .P1_P2_U3289(p1_p2_u3289), .P1_P2_U3290(p1_p2_u3290), .P1_P2_U2867(p1_p2_u2867), .P1_P2_U2866(p1_p2_u2866), .P1_P2_U2865(p1_p2_u2865), .P1_P2_U2864(p1_p2_u2864), .P1_P2_U2863(p1_p2_u2863), .P1_P2_U2862(p1_p2_u2862), .P1_P2_U2861(p1_p2_u2861), .P1_P2_U2860(p1_p2_u2860), .P1_P2_U2859(p1_p2_u2859), .P1_P2_U2858(p1_p2_u2858), .P1_P2_U2857(p1_p2_u2857), .P1_P2_U2856(p1_p2_u2856), .P1_P2_U2855(p1_p2_u2855), .P1_P2_U2854(p1_p2_u2854), .P1_P2_U2853(p1_p2_u2853), .P1_P2_U2852(p1_p2_u2852), .P1_P2_U2851(p1_p2_u2851), .P1_P2_U2850(p1_p2_u2850), .P1_P2_U2849(p1_p2_u2849), .P1_P2_U2848(p1_p2_u2848), .P1_P2_U2847(p1_p2_u2847), .P1_P2_U2846(p1_p2_u2846), .P1_P2_U2845(p1_p2_u2845), .P1_P2_U2844(p1_p2_u2844), .P1_P2_U2843(p1_p2_u2843), .P1_P2_U2842(p1_p2_u2842), .P1_P2_U2841(p1_p2_u2841), .P1_P2_U2840(p1_p2_u2840), .P1_P2_U2839(p1_p2_u2839), .P1_P2_U2838(p1_p2_u2838), .P1_P2_U2837(p1_p2_u2837), .P1_P2_U2836(p1_p2_u2836), .P1_P2_U2835(p1_p2_u2835), .P1_P2_U2834(p1_p2_u2834), .P1_P2_U2833(p1_p2_u2833), .P1_P2_U2832(p1_p2_u2832), .P1_P2_U2831(p1_p2_u2831), .P1_P2_U2830(p1_p2_u2830), .P1_P2_U2829(p1_p2_u2829), .P1_P2_U2828(p1_p2_u2828), .P1_P2_U2827(p1_p2_u2827), .P1_P2_U2826(p1_p2_u2826), .P1_P2_U2825(p1_p2_u2825), .P1_P2_U2824(p1_p2_u2824), .P1_P2_U2823(p1_p2_u2823), .P1_P2_U2822(p1_p2_u2822), .P1_P2_U2821(p1_p2_u2821), .P1_P2_U2820(p1_p2_u2820), .P1_P2_U2819(p1_p2_u2819), .P1_P2_U2818(p1_p2_u2818), .P1_P2_U2817(p1_p2_u2817), .P1_P2_U2816(p1_p2_u2816), .P1_P2_U2815(p1_p2_u2815), .P1_P2_U2814(p1_p2_u2814), .P1_P2_U2813(p1_p2_u2813), .P1_P2_U2812(p1_p2_u2812), .P1_P2_U2811(p1_p2_u2811), .P1_P2_U2810(p1_p2_u2810), .P1_P2_U2809(p1_p2_u2809), .P1_P2_U2808(p1_p2_u2808), .P1_P2_U2807(p1_p2_u2807), .P1_P2_U2806(p1_p2_u2806), .P1_P2_U2805(p1_p2_u2805), .P1_P2_U2804(p1_p2_u2804), .P1_P2_U2803(p1_p2_u2803), .P1_P2_U2802(p1_p2_u2802), .P1_P2_U2801(p1_p2_u2801), .P1_P2_U2800(p1_p2_u2800), .P1_P2_U2799(p1_p2_u2799), .P1_P2_U2798(p1_p2_u2798), .P1_P2_U2797(p1_p2_u2797), .P1_P2_U2796(p1_p2_u2796), .P1_P2_U2795(p1_p2_u2795), .P1_P2_U2794(p1_p2_u2794), .P1_P2_U2793(p1_p2_u2793), .P1_P2_U2792(p1_p2_u2792), .P1_P2_U2791(p1_p2_u2791), .P1_P2_U2790(p1_p2_u2790), .P1_P2_U2789(p1_p2_u2789), .P1_P2_U2788(p1_p2_u2788), .P1_P2_U2787(p1_p2_u2787), .P1_P2_U2786(p1_p2_u2786), .P1_P2_U2785(p1_p2_u2785), .P1_P2_U2784(p1_p2_u2784), .P1_P2_U2783(p1_p2_u2783), .P1_P2_U2782(p1_p2_u2782), .P1_P2_U2781(p1_p2_u2781), .P1_P2_U2780(p1_p2_u2780), .P1_P2_U2779(p1_p2_u2779), .P1_P2_U2778(p1_p2_u2778), .P1_P2_U2777(p1_p2_u2777), .P1_P2_U2776(p1_p2_u2776), .P1_P2_U2775(p1_p2_u2775), .P1_P2_U2774(p1_p2_u2774), .P1_P2_U2773(p1_p2_u2773), .P1_P2_U2772(p1_p2_u2772), .P1_P2_U2771(p1_p2_u2771), .P1_P2_U2770(p1_p2_u2770), .P1_P2_U2769(p1_p2_u2769), .P1_P2_U2768(p1_p2_u2768), .P1_P2_U2767(p1_p2_u2767), .P1_P2_U2766(p1_p2_u2766), .P1_P2_U2765(p1_p2_u2765), .P1_P2_U2764(p1_p2_u2764), .P1_P2_U2763(p1_p2_u2763), .P1_P2_U2762(p1_p2_u2762), .P1_P2_U2761(p1_p2_u2761), .P1_P2_U2760(p1_p2_u2760), .P1_P2_U2759(p1_p2_u2759), .P1_P2_U2758(p1_p2_u2758), .P1_P2_U2757(p1_p2_u2757), .P1_P2_U2756(p1_p2_u2756), .P1_P2_U2755(p1_p2_u2755), .P1_P2_U2754(p1_p2_u2754), .P1_P2_U2753(p1_p2_u2753), .P1_P2_U2752(p1_p2_u2752), .P1_P2_U2751(p1_p2_u2751), .P1_P2_U2750(p1_p2_u2750), .P1_P2_U2749(p1_p2_u2749), .P1_P2_U2748(p1_p2_u2748), .P1_P2_U2747(p1_p2_u2747), .P1_P2_U2746(p1_p2_u2746), .P1_P2_U2745(p1_p2_u2745), .P1_P2_U2744(p1_p2_u2744), .P1_P2_U2743(p1_p2_u2743), .P1_P2_U2742(p1_p2_u2742), .P1_P2_U2741(p1_p2_u2741), .P1_P2_U2740(p1_p2_u2740), .P1_P2_U2739(p1_p2_u2739), .P1_P2_U2738(p1_p2_u2738), .P1_P2_U2737(p1_p2_u2737), .P1_P2_U2736(p1_p2_u2736), .P1_P2_U2735(p1_p2_u2735), .P1_P2_U2734(p1_p2_u2734), .P1_P2_U2733(p1_p2_u2733), .P1_P2_U2732(p1_p2_u2732), .P1_P2_U2731(p1_p2_u2731), .P1_P2_U2730(p1_p2_u2730), .P1_P2_U2729(p1_p2_u2729), .P1_P2_U2728(p1_p2_u2728), .P1_P2_U2727(p1_p2_u2727), .P1_P2_U2726(p1_p2_u2726), .P1_P2_U2725(p1_p2_u2725), .P1_P2_U2724(p1_p2_u2724), .P1_P2_U2723(p1_p2_u2723), .P1_P2_U2722(p1_p2_u2722), .P1_P2_U2721(p1_p2_u2721), .P1_P2_U2720(p1_p2_u2720), .P1_P2_U2719(p1_p2_u2719), .P1_P2_U2718(p1_p2_u2718), .P1_P2_U2717(p1_p2_u2717), .P1_P2_U2716(p1_p2_u2716), .P1_P2_U2715(p1_p2_u2715), .P1_P2_U2714(p1_p2_u2714), .P1_P2_U2713(p1_p2_u2713), .P1_P2_U2712(p1_p2_u2712), .P1_P2_U2711(p1_p2_u2711), .P1_P2_U2710(p1_p2_u2710), .P1_P2_U2709(p1_p2_u2709), .P1_P2_U2708(p1_p2_u2708), .P1_P2_U2707(p1_p2_u2707), .P1_P2_U2706(p1_p2_u2706), .P1_P2_U2705(p1_p2_u2705), .P1_P2_U2704(p1_p2_u2704), .P1_P2_U2703(p1_p2_u2703), .P1_P2_U2702(p1_p2_u2702), .P1_P2_U2701(p1_p2_u2701), .P1_P2_U2700(p1_p2_u2700), .P1_P2_U2699(p1_p2_u2699), .P1_P2_U2698(p1_p2_u2698), .P1_P2_U2697(p1_p2_u2697), .P1_P2_U2696(p1_p2_u2696), .P1_P2_U2695(p1_p2_u2695), .P1_P2_U2694(p1_p2_u2694), .P1_P2_U2693(p1_p2_u2693), .P1_P2_U2692(p1_p2_u2692), .P1_P2_U2691(p1_p2_u2691), .P1_P2_U2690(p1_p2_u2690), .P1_P2_U2689(p1_p2_u2689), .P1_P2_U2688(p1_p2_u2688), .P1_P2_U2687(p1_p2_u2687), .P1_P2_U2686(p1_p2_u2686), .P1_P2_U2685(p1_p2_u2685), .P1_P2_U2684(p1_p2_u2684), .P1_P2_U2683(p1_p2_u2683), .P1_P2_U2682(p1_p2_u2682), .P1_P2_U2681(p1_p2_u2681), .P1_P2_U2680(p1_p2_u2680), .P1_P2_U2679(p1_p2_u2679), .P1_P2_U2678(p1_p2_u2678), .P1_P2_U2677(p1_p2_u2677), .P1_P2_U2676(p1_p2_u2676), .P1_P2_U2675(p1_p2_u2675), .P1_P2_U2674(p1_p2_u2674), .P1_P2_U2673(p1_p2_u2673), .P1_P2_U2672(p1_p2_u2672), .P1_P2_U2671(p1_p2_u2671), .P1_P2_U2670(p1_p2_u2670), .P1_P2_U2669(p1_p2_u2669), .P1_P2_U2668(p1_p2_u2668), .P1_P2_U2667(p1_p2_u2667), .P1_P2_U2666(p1_p2_u2666), .P1_P2_U2665(p1_p2_u2665), .P1_P2_U2664(p1_p2_u2664), .P1_P2_U2663(p1_p2_u2663), .P1_P2_U2662(p1_p2_u2662), .P1_P2_U2661(p1_p2_u2661), .P1_P2_U2660(p1_p2_u2660), .P1_P2_U2659(p1_p2_u2659), .P1_P2_U2658(p1_p2_u2658), .P1_P2_U2657(p1_p2_u2657), .P1_P2_U2656(p1_p2_u2656), .P1_P2_U2655(p1_p2_u2655), .P1_P2_U2654(p1_p2_u2654), .P1_P2_U2653(p1_p2_u2653), .P1_P2_U2652(p1_p2_u2652), .P1_P2_U2651(p1_p2_u2651), .P1_P2_U2650(p1_p2_u2650), .P1_P2_U2649(p1_p2_u2649), .P1_P2_U2648(p1_p2_u2648), .P1_P2_U2647(p1_p2_u2647), .P1_P2_U2646(p1_p2_u2646), .P1_P2_U2645(p1_p2_u2645), .P1_P2_U2644(p1_p2_u2644), .P1_P2_U2643(p1_p2_u2643), .P1_P2_U2642(p1_p2_u2642), .P1_P2_U2641(p1_p2_u2641), .P1_P2_U2640(p1_p2_u2640), .P1_P2_U2639(p1_p2_u2639), .P1_P2_U3292(p1_p2_u3292), .P1_P2_U2638(p1_p2_u2638), .P1_P2_U3293(p1_p2_u3293), .P1_P2_U3294(p1_p2_u3294), .P1_P2_U2637(p1_p2_u2637), .P1_P2_U3295(p1_p2_u3295), .P1_P2_U2636(p1_p2_u2636), .P1_P2_U3296(p1_p2_u3296), .P1_P2_U2635(p1_p2_u2635), .P1_P2_U3297(p1_p2_u3297), .P1_P2_U2634(p1_p2_u2634), .P1_P2_U2633(p1_p2_u2633), .P1_P2_U3298(p1_p2_u3298), .P1_P2_U3299(p1_p2_u3299), .P1_P1_U3288(p1_p1_u3288), .P1_P1_U3289(p1_p1_u3289), .P1_P1_U3290(p1_p1_u3290), .P1_P1_U3291(p1_p1_u3291), .P1_P1_U3077(p1_p1_u3077), .P1_P1_U3076(p1_p1_u3076), .P1_P1_U3075(p1_p1_u3075), .P1_P1_U3074(p1_p1_u3074), .P1_P1_U3073(p1_p1_u3073), .P1_P1_U3072(p1_p1_u3072), .P1_P1_U3071(p1_p1_u3071), .P1_P1_U3070(p1_p1_u3070), .P1_P1_U3069(p1_p1_u3069), .P1_P1_U3068(p1_p1_u3068), .P1_P1_U3067(p1_p1_u3067), .P1_P1_U3066(p1_p1_u3066), .P1_P1_U3065(p1_p1_u3065), .P1_P1_U3064(p1_p1_u3064), .P1_P1_U3063(p1_p1_u3063), .P1_P1_U3062(p1_p1_u3062), .P1_P1_U3061(p1_p1_u3061), .P1_P1_U3060(p1_p1_u3060), .P1_P1_U3059(p1_p1_u3059), .P1_P1_U3058(p1_p1_u3058), .P1_P1_U3057(p1_p1_u3057), .P1_P1_U3056(p1_p1_u3056), .P1_P1_U3055(p1_p1_u3055), .P1_P1_U3054(p1_p1_u3054), .P1_P1_U3053(p1_p1_u3053), .P1_P1_U3052(p1_p1_u3052), .P1_P1_U3051(p1_p1_u3051), .P1_P1_U3050(p1_p1_u3050), .P1_P1_U3049(p1_p1_u3049), .P1_P1_U3048(p1_p1_u3048), .P1_P1_U3047(p1_p1_u3047), .P1_P1_U3046(p1_p1_u3046), .P1_P1_U3045(p1_p1_u3045), .P1_P1_U3294(p1_p1_u3294), .P1_P1_U3295(p1_p1_u3295), .P1_P1_U3044(p1_p1_u3044), .P1_P1_U3043(p1_p1_u3043), .P1_P1_U3042(p1_p1_u3042), .P1_P1_U3041(p1_p1_u3041), .P1_P1_U3040(p1_p1_u3040), .P1_P1_U3039(p1_p1_u3039), .P1_P1_U3038(p1_p1_u3038), .P1_P1_U3037(p1_p1_u3037), .P1_P1_U3036(p1_p1_u3036), .P1_P1_U3035(p1_p1_u3035), .P1_P1_U3034(p1_p1_u3034), .P1_P1_U3033(p1_p1_u3033), .P1_P1_U3032(p1_p1_u3032), .P1_P1_U3031(p1_p1_u3031), .P1_P1_U3030(p1_p1_u3030), .P1_P1_U3029(p1_p1_u3029), .P1_P1_U3028(p1_p1_u3028), .P1_P1_U3027(p1_p1_u3027), .P1_P1_U3026(p1_p1_u3026), .P1_P1_U3025(p1_p1_u3025), .P1_P1_U3024(p1_p1_u3024), .P1_P1_U3023(p1_p1_u3023), .P1_P1_U3022(p1_p1_u3022), .P1_P1_U3021(p1_p1_u3021), .P1_P1_U3020(p1_p1_u3020), .P1_P1_U3019(p1_p1_u3019), .P1_P1_U3018(p1_p1_u3018), .P1_P1_U3017(p1_p1_u3017), .P1_P1_U3016(p1_p1_u3016), .P1_P1_U3015(p1_p1_u3015), .P1_P1_U3296(p1_p1_u3296), .P1_P1_U3014(p1_p1_u3014), .P1_P1_U3013(p1_p1_u3013), .P1_P1_U3012(p1_p1_u3012), .P1_P1_U3011(p1_p1_u3011), .P1_P1_U3010(p1_p1_u3010), .P1_P1_U3009(p1_p1_u3009), .P1_P1_U3008(p1_p1_u3008), .P1_P1_U3007(p1_p1_u3007), .P1_P1_U3006(p1_p1_u3006), .P1_P1_U3005(p1_p1_u3005), .P1_P1_U3004(p1_p1_u3004), .P1_P1_U3003(p1_p1_u3003), .P1_P1_U3002(p1_p1_u3002), .P1_P1_U3001(p1_p1_u3001), .P1_P1_U3000(p1_p1_u3000), .P1_P1_U2999(p1_p1_u2999), .P1_P1_U2998(p1_p1_u2998), .P1_P1_U2997(p1_p1_u2997), .P1_P1_U2996(p1_p1_u2996), .P1_P1_U2995(p1_p1_u2995), .P1_P1_U2994(p1_p1_u2994), .P1_P1_U2993(p1_p1_u2993), .P1_P1_U2992(p1_p1_u2992), .P1_P1_U2991(p1_p1_u2991), .P1_P1_U2990(p1_p1_u2990), .P1_P1_U2989(p1_p1_u2989), .P1_P1_U2988(p1_p1_u2988), .P1_P1_U2987(p1_p1_u2987), .P1_P1_U2986(p1_p1_u2986), .P1_P1_U2985(p1_p1_u2985), .P1_P1_U2984(p1_p1_u2984), .P1_P1_U2983(p1_p1_u2983), .P1_P1_U2982(p1_p1_u2982), .P1_P1_U2981(p1_p1_u2981), .P1_P1_U2980(p1_p1_u2980), .P1_P1_U2979(p1_p1_u2979), .P1_P1_U2978(p1_p1_u2978), .P1_P1_U2977(p1_p1_u2977), .P1_P1_U2976(p1_p1_u2976), .P1_P1_U2975(p1_p1_u2975), .P1_P1_U2974(p1_p1_u2974), .P1_P1_U2973(p1_p1_u2973), .P1_P1_U2972(p1_p1_u2972), .P1_P1_U2971(p1_p1_u2971), .P1_P1_U2970(p1_p1_u2970), .P1_P1_U2969(p1_p1_u2969), .P1_P1_U2968(p1_p1_u2968), .P1_P1_U2967(p1_p1_u2967), .P1_P1_U2966(p1_p1_u2966), .P1_P1_U2965(p1_p1_u2965), .P1_P1_U2964(p1_p1_u2964), .P1_P1_U2963(p1_p1_u2963), .P1_P1_U2962(p1_p1_u2962), .P1_P1_U2961(p1_p1_u2961), .P1_P1_U2960(p1_p1_u2960), .P1_P1_U2959(p1_p1_u2959), .P1_P1_U2958(p1_p1_u2958), .P1_P1_U2957(p1_p1_u2957), .P1_P1_U2956(p1_p1_u2956), .P1_P1_U2955(p1_p1_u2955), .P1_P1_U2954(p1_p1_u2954), .P1_P1_U2953(p1_p1_u2953), .P1_P1_U2952(p1_p1_u2952), .P1_P1_U2951(p1_p1_u2951), .P1_P1_U2950(p1_p1_u2950), .P1_P1_U2949(p1_p1_u2949), .P1_P1_U2948(p1_p1_u2948), .P1_P1_U2947(p1_p1_u2947), .P1_P1_U2946(p1_p1_u2946), .P1_P1_U2945(p1_p1_u2945), .P1_P1_U2944(p1_p1_u2944), .P1_P1_U2943(p1_p1_u2943), .P1_P1_U2942(p1_p1_u2942), .P1_P1_U2941(p1_p1_u2941), .P1_P1_U2940(p1_p1_u2940), .P1_P1_U2939(p1_p1_u2939), .P1_P1_U2938(p1_p1_u2938), .P1_P1_U2937(p1_p1_u2937), .P1_P1_U2936(p1_p1_u2936), .P1_P1_U2935(p1_p1_u2935), .P1_P1_U2934(p1_p1_u2934), .P1_P1_U2933(p1_p1_u2933), .P1_P1_U2932(p1_p1_u2932), .P1_P1_U2931(p1_p1_u2931), .P1_P1_U2930(p1_p1_u2930), .P1_P1_U2929(p1_p1_u2929), .P1_P1_U2928(p1_p1_u2928), .P1_P1_U2927(p1_p1_u2927), .P1_P1_U2926(p1_p1_u2926), .P1_P1_U2925(p1_p1_u2925), .P1_P1_U2924(p1_p1_u2924), .P1_P1_U2923(p1_p1_u2923), .P1_P1_U2922(p1_p1_u2922), .P1_P1_U2921(p1_p1_u2921), .P1_P1_U2920(p1_p1_u2920), .P1_P1_U2919(p1_p1_u2919), .P1_P1_U2918(p1_p1_u2918), .P1_P1_U2917(p1_p1_u2917), .P1_P1_U2916(p1_p1_u2916), .P1_P1_U2915(p1_p1_u2915), .P1_P1_U2914(p1_p1_u2914), .P1_P1_U2913(p1_p1_u2913), .P1_P1_U2912(p1_p1_u2912), .P1_P1_U2911(p1_p1_u2911), .P1_P1_U2910(p1_p1_u2910), .P1_P1_U2909(p1_p1_u2909), .P1_P1_U2908(p1_p1_u2908), .P1_P1_U2907(p1_p1_u2907), .P1_P1_U2906(p1_p1_u2906), .P1_P1_U2905(p1_p1_u2905), .P1_P1_U2904(p1_p1_u2904), .P1_P1_U2903(p1_p1_u2903), .P1_P1_U2902(p1_p1_u2902), .P1_P1_U2901(p1_p1_u2901), .P1_P1_U2900(p1_p1_u2900), .P1_P1_U2899(p1_p1_u2899), .P1_P1_U2898(p1_p1_u2898), .P1_P1_U2897(p1_p1_u2897), .P1_P1_U2896(p1_p1_u2896), .P1_P1_U2895(p1_p1_u2895), .P1_P1_U2894(p1_p1_u2894), .P1_P1_U2893(p1_p1_u2893), .P1_P1_U2892(p1_p1_u2892), .P1_P1_U2891(p1_p1_u2891), .P1_P1_U2890(p1_p1_u2890), .P1_P1_U2889(p1_p1_u2889), .P1_P1_U2888(p1_p1_u2888), .P1_P1_U2887(p1_p1_u2887), .P1_P1_U2886(p1_p1_u2886), .P1_P1_U2885(p1_p1_u2885), .P1_P1_U2884(p1_p1_u2884), .P1_P1_U3298(p1_p1_u3298), .P1_P1_U3299(p1_p1_u3299), .P1_P1_U3302(p1_p1_u3302), .P1_P1_U3303(p1_p1_u3303), .P1_P1_U3304(p1_p1_u3304), .P1_P1_U2883(p1_p1_u2883), .P1_P1_U2882(p1_p1_u2882), .P1_P1_U2881(p1_p1_u2881), .P1_P1_U2880(p1_p1_u2880), .P1_P1_U2879(p1_p1_u2879), .P1_P1_U2878(p1_p1_u2878), .P1_P1_U2877(p1_p1_u2877), .P1_P1_U2876(p1_p1_u2876), .P1_P1_U2875(p1_p1_u2875), .P1_P1_U2874(p1_p1_u2874), .P1_P1_U2873(p1_p1_u2873), .P1_P1_U2872(p1_p1_u2872), .P1_P1_U2871(p1_p1_u2871), .P1_P1_U2870(p1_p1_u2870), .P1_P1_U2869(p1_p1_u2869), .P1_P1_U2868(p1_p1_u2868), .P1_P1_U2867(p1_p1_u2867), .P1_P1_U2866(p1_p1_u2866), .P1_P1_U2865(p1_p1_u2865), .P1_P1_U2864(p1_p1_u2864), .P1_P1_U2863(p1_p1_u2863), .P1_P1_U2862(p1_p1_u2862), .P1_P1_U2861(p1_p1_u2861), .P1_P1_U2860(p1_p1_u2860), .P1_P1_U2859(p1_p1_u2859), .P1_P1_U2858(p1_p1_u2858), .P1_P1_U2857(p1_p1_u2857), .P1_P1_U2856(p1_p1_u2856), .P1_P1_U2855(p1_p1_u2855), .P1_P1_U2854(p1_p1_u2854), .P1_P1_U2853(p1_p1_u2853), .P1_P1_U2852(p1_p1_u2852), .P1_P1_U2851(p1_p1_u2851), .P1_P1_U2850(p1_p1_u2850), .P1_P1_U2849(p1_p1_u2849), .P1_P1_U2848(p1_p1_u2848), .P1_P1_U2847(p1_p1_u2847), .P1_P1_U2846(p1_p1_u2846), .P1_P1_U2845(p1_p1_u2845), .P1_P1_U2844(p1_p1_u2844), .P1_P1_U2843(p1_p1_u2843), .P1_P1_U2842(p1_p1_u2842), .P1_P1_U2841(p1_p1_u2841), .P1_P1_U2840(p1_p1_u2840), .P1_P1_U2839(p1_p1_u2839), .P1_P1_U2838(p1_p1_u2838), .P1_P1_U2837(p1_p1_u2837), .P1_P1_U2836(p1_p1_u2836), .P1_P1_U2835(p1_p1_u2835), .P1_P1_U2834(p1_p1_u2834), .P1_P1_U2833(p1_p1_u2833), .P1_P1_U2832(p1_p1_u2832), .P1_P1_U2831(p1_p1_u2831), .P1_P1_U2830(p1_p1_u2830), .P1_P1_U2829(p1_p1_u2829), .P1_P1_U2828(p1_p1_u2828), .P1_P1_U2827(p1_p1_u2827), .P1_P1_U2826(p1_p1_u2826), .P1_P1_U2825(p1_p1_u2825), .P1_P1_U2824(p1_p1_u2824), .P1_P1_U2823(p1_p1_u2823), .P1_P1_U2822(p1_p1_u2822), .P1_P1_U2821(p1_p1_u2821), .P1_P1_U2820(p1_p1_u2820), .P1_P1_U2819(p1_p1_u2819), .P1_P1_U2818(p1_p1_u2818), .P1_P1_U2817(p1_p1_u2817), .P1_P1_U2816(p1_p1_u2816), .P1_P1_U2815(p1_p1_u2815), .P1_P1_U2814(p1_p1_u2814), .P1_P1_U2813(p1_p1_u2813), .P1_P1_U2812(p1_p1_u2812), .P1_P1_U2811(p1_p1_u2811), .P1_P1_U2810(p1_p1_u2810), .P1_P1_U2809(p1_p1_u2809), .P1_P1_U2808(p1_p1_u2808), .P1_P1_U2807(p1_p1_u2807), .P1_P1_U2806(p1_p1_u2806), .P1_P1_U2805(p1_p1_u2805), .P1_P1_U2804(p1_p1_u2804), .P1_P1_U2803(p1_p1_u2803), .P1_P1_U2802(p1_p1_u2802), .P1_P1_U2801(p1_p1_u2801), .P1_P1_U2800(p1_p1_u2800), .P1_P1_U2799(p1_p1_u2799), .P1_P1_U2798(p1_p1_u2798), .P1_P1_U2797(p1_p1_u2797), .P1_P1_U2796(p1_p1_u2796), .P1_P1_U2795(p1_p1_u2795), .P1_P1_U2794(p1_p1_u2794), .P1_P1_U2793(p1_p1_u2793), .P1_P1_U2792(p1_p1_u2792), .P1_P1_U2791(p1_p1_u2791), .P1_P1_U2790(p1_p1_u2790), .P1_P1_U2789(p1_p1_u2789), .P1_P1_U2788(p1_p1_u2788), .P1_P1_U2787(p1_p1_u2787), .P1_P1_U2786(p1_p1_u2786), .P1_P1_U2785(p1_p1_u2785), .P1_P1_U2784(p1_p1_u2784), .P1_P1_U2783(p1_p1_u2783), .P1_P1_U2782(p1_p1_u2782), .P1_P1_U2781(p1_p1_u2781), .P1_P1_U2780(p1_p1_u2780), .P1_P1_U2779(p1_p1_u2779), .P1_P1_U2778(p1_p1_u2778), .P1_P1_U2777(p1_p1_u2777), .P1_P1_U2776(p1_p1_u2776), .P1_P1_U2775(p1_p1_u2775), .P1_P1_U2774(p1_p1_u2774), .P1_P1_U2773(p1_p1_u2773), .P1_P1_U2772(p1_p1_u2772), .P1_P1_U2771(p1_p1_u2771), .P1_P1_U2770(p1_p1_u2770), .P1_P1_U2769(p1_p1_u2769), .P1_P1_U2768(p1_p1_u2768), .P1_P1_U2767(p1_p1_u2767), .P1_P1_U2766(p1_p1_u2766), .P1_P1_U2765(p1_p1_u2765), .P1_P1_U2764(p1_p1_u2764), .P1_P1_U2763(p1_p1_u2763), .P1_P1_U2762(p1_p1_u2762), .P1_P1_U2761(p1_p1_u2761), .P1_P1_U2760(p1_p1_u2760), .P1_P1_U2759(p1_p1_u2759), .P1_P1_U2758(p1_p1_u2758), .P1_P1_U2757(p1_p1_u2757), .P1_P1_U2756(p1_p1_u2756), .P1_P1_U2755(p1_p1_u2755), .P1_P1_U2754(p1_p1_u2754), .P1_P1_U2753(p1_p1_u2753), .P1_P1_U2752(p1_p1_u2752), .P1_P1_U2751(p1_p1_u2751), .P1_P1_U2750(p1_p1_u2750), .P1_P1_U2749(p1_p1_u2749), .P1_P1_U2748(p1_p1_u2748), .P1_P1_U2747(p1_p1_u2747), .P1_P1_U2746(p1_p1_u2746), .P1_P1_U2745(p1_p1_u2745), .P1_P1_U2744(p1_p1_u2744), .P1_P1_U2743(p1_p1_u2743), .P1_P1_U2742(p1_p1_u2742), .P1_P1_U2741(p1_p1_u2741), .P1_P1_U2740(p1_p1_u2740), .P1_P1_U2739(p1_p1_u2739), .P1_P1_U2738(p1_p1_u2738), .P1_P1_U2737(p1_p1_u2737), .P1_P1_U2736(p1_p1_u2736), .P1_P1_U2735(p1_p1_u2735), .P1_P1_U2734(p1_p1_u2734), .P1_P1_U2733(p1_p1_u2733), .P1_P1_U2732(p1_p1_u2732), .P1_P1_U2731(p1_p1_u2731), .P1_P1_U2730(p1_p1_u2730), .P1_P1_U2729(p1_p1_u2729), .P1_P1_U2728(p1_p1_u2728), .P1_P1_U2727(p1_p1_u2727), .P1_P1_U2726(p1_p1_u2726), .P1_P1_U2725(p1_p1_u2725), .P1_P1_U2724(p1_p1_u2724), .P1_P1_U2723(p1_p1_u2723), .P1_P1_U2722(p1_p1_u2722), .P1_P1_U2721(p1_p1_u2721), .P1_P1_U2720(p1_p1_u2720), .P1_P1_U2719(p1_p1_u2719), .P1_P1_U2718(p1_p1_u2718), .P1_P1_U2717(p1_p1_u2717), .P1_P1_U2716(p1_p1_u2716), .P1_P1_U2715(p1_p1_u2715), .P1_P1_U2714(p1_p1_u2714), .P1_P1_U2713(p1_p1_u2713), .P1_P1_U2712(p1_p1_u2712), .P1_P1_U2711(p1_p1_u2711), .P1_P1_U2710(p1_p1_u2710), .P1_P1_U2709(p1_p1_u2709), .P1_P1_U2708(p1_p1_u2708), .P1_P1_U2707(p1_p1_u2707), .P1_P1_U2706(p1_p1_u2706), .P1_P1_U2705(p1_p1_u2705), .P1_P1_U2704(p1_p1_u2704), .P1_P1_U2703(p1_p1_u2703), .P1_P1_U2702(p1_p1_u2702), .P1_P1_U2701(p1_p1_u2701), .P1_P1_U2700(p1_p1_u2700), .P1_P1_U2699(p1_p1_u2699), .P1_P1_U2698(p1_p1_u2698), .P1_P1_U2697(p1_p1_u2697), .P1_P1_U2696(p1_p1_u2696), .P1_P1_U2695(p1_p1_u2695), .P1_P1_U2694(p1_p1_u2694), .P1_P1_U2693(p1_p1_u2693), .P1_P1_U2692(p1_p1_u2692), .P1_P1_U2691(p1_p1_u2691), .P1_P1_U2690(p1_p1_u2690), .P1_P1_U2689(p1_p1_u2689), .P1_P1_U2688(p1_p1_u2688), .P1_P1_U2687(p1_p1_u2687), .P1_P1_U2686(p1_p1_u2686), .P1_P1_U2685(p1_p1_u2685), .P1_P1_U2684(p1_p1_u2684), .P1_P1_U2683(p1_p1_u2683), .P1_P1_U2682(p1_p1_u2682), .P1_P1_U2681(p1_p1_u2681), .P1_P1_U2680(p1_p1_u2680), .P1_P1_U2679(p1_p1_u2679), .P1_P1_U2678(p1_p1_u2678), .P1_P1_U2677(p1_p1_u2677), .P1_P1_U2676(p1_p1_u2676), .P1_P1_U2675(p1_p1_u2675), .P1_P1_U2674(p1_p1_u2674), .P1_P1_U2673(p1_p1_u2673), .P1_P1_U2672(p1_p1_u2672), .P1_P1_U2671(p1_p1_u2671), .P1_P1_U2670(p1_p1_u2670), .P1_P1_U2669(p1_p1_u2669), .P1_P1_U2668(p1_p1_u2668), .P1_P1_U2667(p1_p1_u2667), .P1_P1_U2666(p1_p1_u2666), .P1_P1_U2665(p1_p1_u2665), .P1_P1_U2664(p1_p1_u2664), .P1_P1_U2663(p1_p1_u2663), .P1_P1_U2662(p1_p1_u2662), .P1_P1_U2661(p1_p1_u2661), .P1_P1_U2660(p1_p1_u2660), .P1_P1_U2659(p1_p1_u2659), .P1_P1_U2658(p1_p1_u2658), .P1_P1_U2657(p1_p1_u2657), .P1_P1_U2656(p1_p1_u2656), .P1_P1_U2655(p1_p1_u2655), .P1_P1_U3306(p1_p1_u3306), .P1_P1_U2654(p1_p1_u2654), .P1_P1_U3307(p1_p1_u3307), .P1_P1_U3308(p1_p1_u3308), .P1_P1_U2653(p1_p1_u2653), .P1_P1_U3309(p1_p1_u3309), .P1_P1_U2652(p1_p1_u2652), .P1_P1_U3310(p1_p1_u3310), .P1_P1_U2651(p1_p1_u2651), .P1_P1_U3311(p1_p1_u3311), .P1_P1_U2650(p1_p1_u2650), .P1_P1_U2649(p1_p1_u2649), .P1_P1_U3312(p1_p1_u3312), .P1_P1_U3313(p1_p1_u3313), .P2_P3_U3274(p2_p3_u3274), .P2_P3_U3275(p2_p3_u3275), .P2_P3_U3276(p2_p3_u3276), .P2_P3_U3277(p2_p3_u3277), .P2_P3_U3061(p2_p3_u3061), .P2_P3_U3060(p2_p3_u3060), .P2_P3_U3059(p2_p3_u3059), .P2_P3_U3058(p2_p3_u3058), .P2_P3_U3057(p2_p3_u3057), .P2_P3_U3056(p2_p3_u3056), .P2_P3_U3055(p2_p3_u3055), .P2_P3_U3054(p2_p3_u3054), .P2_P3_U3053(p2_p3_u3053), .P2_P3_U3052(p2_p3_u3052), .P2_P3_U3051(p2_p3_u3051), .P2_P3_U3050(p2_p3_u3050), .P2_P3_U3049(p2_p3_u3049), .P2_P3_U3048(p2_p3_u3048), .P2_P3_U3047(p2_p3_u3047), .P2_P3_U3046(p2_p3_u3046), .P2_P3_U3045(p2_p3_u3045), .P2_P3_U3044(p2_p3_u3044), .P2_P3_U3043(p2_p3_u3043), .P2_P3_U3042(p2_p3_u3042), .P2_P3_U3041(p2_p3_u3041), .P2_P3_U3040(p2_p3_u3040), .P2_P3_U3039(p2_p3_u3039), .P2_P3_U3038(p2_p3_u3038), .P2_P3_U3037(p2_p3_u3037), .P2_P3_U3036(p2_p3_u3036), .P2_P3_U3035(p2_p3_u3035), .P2_P3_U3034(p2_p3_u3034), .P2_P3_U3033(p2_p3_u3033), .P2_P3_U3032(p2_p3_u3032), .P2_P3_U3031(p2_p3_u3031), .P2_P3_U3030(p2_p3_u3030), .P2_P3_U3029(p2_p3_u3029), .P2_P3_U3280(p2_p3_u3280), .P2_P3_U3281(p2_p3_u3281), .P2_P3_U3028(p2_p3_u3028), .P2_P3_U3027(p2_p3_u3027), .P2_P3_U3026(p2_p3_u3026), .P2_P3_U3025(p2_p3_u3025), .P2_P3_U3024(p2_p3_u3024), .P2_P3_U3023(p2_p3_u3023), .P2_P3_U3022(p2_p3_u3022), .P2_P3_U3021(p2_p3_u3021), .P2_P3_U3020(p2_p3_u3020), .P2_P3_U3019(p2_p3_u3019), .P2_P3_U3018(p2_p3_u3018), .P2_P3_U3017(p2_p3_u3017), .P2_P3_U3016(p2_p3_u3016), .P2_P3_U3015(p2_p3_u3015), .P2_P3_U3014(p2_p3_u3014), .P2_P3_U3013(p2_p3_u3013), .P2_P3_U3012(p2_p3_u3012), .P2_P3_U3011(p2_p3_u3011), .P2_P3_U3010(p2_p3_u3010), .P2_P3_U3009(p2_p3_u3009), .P2_P3_U3008(p2_p3_u3008), .P2_P3_U3007(p2_p3_u3007), .P2_P3_U3006(p2_p3_u3006), .P2_P3_U3005(p2_p3_u3005), .P2_P3_U3004(p2_p3_u3004), .P2_P3_U3003(p2_p3_u3003), .P2_P3_U3002(p2_p3_u3002), .P2_P3_U3001(p2_p3_u3001), .P2_P3_U3000(p2_p3_u3000), .P2_P3_U2999(p2_p3_u2999), .P2_P3_U3282(p2_p3_u3282), .P2_P3_U2998(p2_p3_u2998), .P2_P3_U2997(p2_p3_u2997), .P2_P3_U2996(p2_p3_u2996), .P2_P3_U2995(p2_p3_u2995), .P2_P3_U2994(p2_p3_u2994), .P2_P3_U2993(p2_p3_u2993), .P2_P3_U2992(p2_p3_u2992), .P2_P3_U2991(p2_p3_u2991), .P2_P3_U2990(p2_p3_u2990), .P2_P3_U2989(p2_p3_u2989), .P2_P3_U2988(p2_p3_u2988), .P2_P3_U2987(p2_p3_u2987), .P2_P3_U2986(p2_p3_u2986), .P2_P3_U2985(p2_p3_u2985), .P2_P3_U2984(p2_p3_u2984), .P2_P3_U2983(p2_p3_u2983), .P2_P3_U2982(p2_p3_u2982), .P2_P3_U2981(p2_p3_u2981), .P2_P3_U2980(p2_p3_u2980), .P2_P3_U2979(p2_p3_u2979), .P2_P3_U2978(p2_p3_u2978), .P2_P3_U2977(p2_p3_u2977), .P2_P3_U2976(p2_p3_u2976), .P2_P3_U2975(p2_p3_u2975), .P2_P3_U2974(p2_p3_u2974), .P2_P3_U2973(p2_p3_u2973), .P2_P3_U2972(p2_p3_u2972), .P2_P3_U2971(p2_p3_u2971), .P2_P3_U2970(p2_p3_u2970), .P2_P3_U2969(p2_p3_u2969), .P2_P3_U2968(p2_p3_u2968), .P2_P3_U2967(p2_p3_u2967), .P2_P3_U2966(p2_p3_u2966), .P2_P3_U2965(p2_p3_u2965), .P2_P3_U2964(p2_p3_u2964), .P2_P3_U2963(p2_p3_u2963), .P2_P3_U2962(p2_p3_u2962), .P2_P3_U2961(p2_p3_u2961), .P2_P3_U2960(p2_p3_u2960), .P2_P3_U2959(p2_p3_u2959), .P2_P3_U2958(p2_p3_u2958), .P2_P3_U2957(p2_p3_u2957), .P2_P3_U2956(p2_p3_u2956), .P2_P3_U2955(p2_p3_u2955), .P2_P3_U2954(p2_p3_u2954), .P2_P3_U2953(p2_p3_u2953), .P2_P3_U2952(p2_p3_u2952), .P2_P3_U2951(p2_p3_u2951), .P2_P3_U2950(p2_p3_u2950), .P2_P3_U2949(p2_p3_u2949), .P2_P3_U2948(p2_p3_u2948), .P2_P3_U2947(p2_p3_u2947), .P2_P3_U2946(p2_p3_u2946), .P2_P3_U2945(p2_p3_u2945), .P2_P3_U2944(p2_p3_u2944), .P2_P3_U2943(p2_p3_u2943), .P2_P3_U2942(p2_p3_u2942), .P2_P3_U2941(p2_p3_u2941), .P2_P3_U2940(p2_p3_u2940), .P2_P3_U2939(p2_p3_u2939), .P2_P3_U2938(p2_p3_u2938), .P2_P3_U2937(p2_p3_u2937), .P2_P3_U2936(p2_p3_u2936), .P2_P3_U2935(p2_p3_u2935), .P2_P3_U2934(p2_p3_u2934), .P2_P3_U2933(p2_p3_u2933), .P2_P3_U2932(p2_p3_u2932), .P2_P3_U2931(p2_p3_u2931), .P2_P3_U2930(p2_p3_u2930), .P2_P3_U2929(p2_p3_u2929), .P2_P3_U2928(p2_p3_u2928), .P2_P3_U2927(p2_p3_u2927), .P2_P3_U2926(p2_p3_u2926), .P2_P3_U2925(p2_p3_u2925), .P2_P3_U2924(p2_p3_u2924), .P2_P3_U2923(p2_p3_u2923), .P2_P3_U2922(p2_p3_u2922), .P2_P3_U2921(p2_p3_u2921), .P2_P3_U2920(p2_p3_u2920), .P2_P3_U2919(p2_p3_u2919), .P2_P3_U2918(p2_p3_u2918), .P2_P3_U2917(p2_p3_u2917), .P2_P3_U2916(p2_p3_u2916), .P2_P3_U2915(p2_p3_u2915), .P2_P3_U2914(p2_p3_u2914), .P2_P3_U2913(p2_p3_u2913), .P2_P3_U2912(p2_p3_u2912), .P2_P3_U2911(p2_p3_u2911), .P2_P3_U2910(p2_p3_u2910), .P2_P3_U2909(p2_p3_u2909), .P2_P3_U2908(p2_p3_u2908), .P2_P3_U2907(p2_p3_u2907), .P2_P3_U2906(p2_p3_u2906), .P2_P3_U2905(p2_p3_u2905), .P2_P3_U2904(p2_p3_u2904), .P2_P3_U2903(p2_p3_u2903), .P2_P3_U2902(p2_p3_u2902), .P2_P3_U2901(p2_p3_u2901), .P2_P3_U2900(p2_p3_u2900), .P2_P3_U2899(p2_p3_u2899), .P2_P3_U2898(p2_p3_u2898), .P2_P3_U2897(p2_p3_u2897), .P2_P3_U2896(p2_p3_u2896), .P2_P3_U2895(p2_p3_u2895), .P2_P3_U2894(p2_p3_u2894), .P2_P3_U2893(p2_p3_u2893), .P2_P3_U2892(p2_p3_u2892), .P2_P3_U2891(p2_p3_u2891), .P2_P3_U2890(p2_p3_u2890), .P2_P3_U2889(p2_p3_u2889), .P2_P3_U2888(p2_p3_u2888), .P2_P3_U2887(p2_p3_u2887), .P2_P3_U2886(p2_p3_u2886), .P2_P3_U2885(p2_p3_u2885), .P2_P3_U2884(p2_p3_u2884), .P2_P3_U2883(p2_p3_u2883), .P2_P3_U2882(p2_p3_u2882), .P2_P3_U2881(p2_p3_u2881), .P2_P3_U2880(p2_p3_u2880), .P2_P3_U2879(p2_p3_u2879), .P2_P3_U2878(p2_p3_u2878), .P2_P3_U2877(p2_p3_u2877), .P2_P3_U2876(p2_p3_u2876), .P2_P3_U2875(p2_p3_u2875), .P2_P3_U2874(p2_p3_u2874), .P2_P3_U2873(p2_p3_u2873), .P2_P3_U2872(p2_p3_u2872), .P2_P3_U2871(p2_p3_u2871), .P2_P3_U2870(p2_p3_u2870), .P2_P3_U2869(p2_p3_u2869), .P2_P3_U2868(p2_p3_u2868), .P2_P3_U3284(p2_p3_u3284), .P2_P3_U3285(p2_p3_u3285), .P2_P3_U3288(p2_p3_u3288), .P2_P3_U3289(p2_p3_u3289), .P2_P3_U3290(p2_p3_u3290), .P2_P3_U2867(p2_p3_u2867), .P2_P3_U2866(p2_p3_u2866), .P2_P3_U2865(p2_p3_u2865), .P2_P3_U2864(p2_p3_u2864), .P2_P3_U2863(p2_p3_u2863), .P2_P3_U2862(p2_p3_u2862), .P2_P3_U2861(p2_p3_u2861), .P2_P3_U2860(p2_p3_u2860), .P2_P3_U2859(p2_p3_u2859), .P2_P3_U2858(p2_p3_u2858), .P2_P3_U2857(p2_p3_u2857), .P2_P3_U2856(p2_p3_u2856), .P2_P3_U2855(p2_p3_u2855), .P2_P3_U2854(p2_p3_u2854), .P2_P3_U2853(p2_p3_u2853), .P2_P3_U2852(p2_p3_u2852), .P2_P3_U2851(p2_p3_u2851), .P2_P3_U2850(p2_p3_u2850), .P2_P3_U2849(p2_p3_u2849), .P2_P3_U2848(p2_p3_u2848), .P2_P3_U2847(p2_p3_u2847), .P2_P3_U2846(p2_p3_u2846), .P2_P3_U2845(p2_p3_u2845), .P2_P3_U2844(p2_p3_u2844), .P2_P3_U2843(p2_p3_u2843), .P2_P3_U2842(p2_p3_u2842), .P2_P3_U2841(p2_p3_u2841), .P2_P3_U2840(p2_p3_u2840), .P2_P3_U2839(p2_p3_u2839), .P2_P3_U2838(p2_p3_u2838), .P2_P3_U2837(p2_p3_u2837), .P2_P3_U2836(p2_p3_u2836), .P2_P3_U2835(p2_p3_u2835), .P2_P3_U2834(p2_p3_u2834), .P2_P3_U2833(p2_p3_u2833), .P2_P3_U2832(p2_p3_u2832), .P2_P3_U2831(p2_p3_u2831), .P2_P3_U2830(p2_p3_u2830), .P2_P3_U2829(p2_p3_u2829), .P2_P3_U2828(p2_p3_u2828), .P2_P3_U2827(p2_p3_u2827), .P2_P3_U2826(p2_p3_u2826), .P2_P3_U2825(p2_p3_u2825), .P2_P3_U2824(p2_p3_u2824), .P2_P3_U2823(p2_p3_u2823), .P2_P3_U2822(p2_p3_u2822), .P2_P3_U2821(p2_p3_u2821), .P2_P3_U2820(p2_p3_u2820), .P2_P3_U2819(p2_p3_u2819), .P2_P3_U2818(p2_p3_u2818), .P2_P3_U2817(p2_p3_u2817), .P2_P3_U2816(p2_p3_u2816), .P2_P3_U2815(p2_p3_u2815), .P2_P3_U2814(p2_p3_u2814), .P2_P3_U2813(p2_p3_u2813), .P2_P3_U2812(p2_p3_u2812), .P2_P3_U2811(p2_p3_u2811), .P2_P3_U2810(p2_p3_u2810), .P2_P3_U2809(p2_p3_u2809), .P2_P3_U2808(p2_p3_u2808), .P2_P3_U2807(p2_p3_u2807), .P2_P3_U2806(p2_p3_u2806), .P2_P3_U2805(p2_p3_u2805), .P2_P3_U2804(p2_p3_u2804), .P2_P3_U2803(p2_p3_u2803), .P2_P3_U2802(p2_p3_u2802), .P2_P3_U2801(p2_p3_u2801), .P2_P3_U2800(p2_p3_u2800), .P2_P3_U2799(p2_p3_u2799), .P2_P3_U2798(p2_p3_u2798), .P2_P3_U2797(p2_p3_u2797), .P2_P3_U2796(p2_p3_u2796), .P2_P3_U2795(p2_p3_u2795), .P2_P3_U2794(p2_p3_u2794), .P2_P3_U2793(p2_p3_u2793), .P2_P3_U2792(p2_p3_u2792), .P2_P3_U2791(p2_p3_u2791), .P2_P3_U2790(p2_p3_u2790), .P2_P3_U2789(p2_p3_u2789), .P2_P3_U2788(p2_p3_u2788), .P2_P3_U2787(p2_p3_u2787), .P2_P3_U2786(p2_p3_u2786), .P2_P3_U2785(p2_p3_u2785), .P2_P3_U2784(p2_p3_u2784), .P2_P3_U2783(p2_p3_u2783), .P2_P3_U2782(p2_p3_u2782), .P2_P3_U2781(p2_p3_u2781), .P2_P3_U2780(p2_p3_u2780), .P2_P3_U2779(p2_p3_u2779), .P2_P3_U2778(p2_p3_u2778), .P2_P3_U2777(p2_p3_u2777), .P2_P3_U2776(p2_p3_u2776), .P2_P3_U2775(p2_p3_u2775), .P2_P3_U2774(p2_p3_u2774), .P2_P3_U2773(p2_p3_u2773), .P2_P3_U2772(p2_p3_u2772), .P2_P3_U2771(p2_p3_u2771), .P2_P3_U2770(p2_p3_u2770), .P2_P3_U2769(p2_p3_u2769), .P2_P3_U2768(p2_p3_u2768), .P2_P3_U2767(p2_p3_u2767), .P2_P3_U2766(p2_p3_u2766), .P2_P3_U2765(p2_p3_u2765), .P2_P3_U2764(p2_p3_u2764), .P2_P3_U2763(p2_p3_u2763), .P2_P3_U2762(p2_p3_u2762), .P2_P3_U2761(p2_p3_u2761), .P2_P3_U2760(p2_p3_u2760), .P2_P3_U2759(p2_p3_u2759), .P2_P3_U2758(p2_p3_u2758), .P2_P3_U2757(p2_p3_u2757), .P2_P3_U2756(p2_p3_u2756), .P2_P3_U2755(p2_p3_u2755), .P2_P3_U2754(p2_p3_u2754), .P2_P3_U2753(p2_p3_u2753), .P2_P3_U2752(p2_p3_u2752), .P2_P3_U2751(p2_p3_u2751), .P2_P3_U2750(p2_p3_u2750), .P2_P3_U2749(p2_p3_u2749), .P2_P3_U2748(p2_p3_u2748), .P2_P3_U2747(p2_p3_u2747), .P2_P3_U2746(p2_p3_u2746), .P2_P3_U2745(p2_p3_u2745), .P2_P3_U2744(p2_p3_u2744), .P2_P3_U2743(p2_p3_u2743), .P2_P3_U2742(p2_p3_u2742), .P2_P3_U2741(p2_p3_u2741), .P2_P3_U2740(p2_p3_u2740), .P2_P3_U2739(p2_p3_u2739), .P2_P3_U2738(p2_p3_u2738), .P2_P3_U2737(p2_p3_u2737), .P2_P3_U2736(p2_p3_u2736), .P2_P3_U2735(p2_p3_u2735), .P2_P3_U2734(p2_p3_u2734), .P2_P3_U2733(p2_p3_u2733), .P2_P3_U2732(p2_p3_u2732), .P2_P3_U2731(p2_p3_u2731), .P2_P3_U2730(p2_p3_u2730), .P2_P3_U2729(p2_p3_u2729), .P2_P3_U2728(p2_p3_u2728), .P2_P3_U2727(p2_p3_u2727), .P2_P3_U2726(p2_p3_u2726), .P2_P3_U2725(p2_p3_u2725), .P2_P3_U2724(p2_p3_u2724), .P2_P3_U2723(p2_p3_u2723), .P2_P3_U2722(p2_p3_u2722), .P2_P3_U2721(p2_p3_u2721), .P2_P3_U2720(p2_p3_u2720), .P2_P3_U2719(p2_p3_u2719), .P2_P3_U2718(p2_p3_u2718), .P2_P3_U2717(p2_p3_u2717), .P2_P3_U2716(p2_p3_u2716), .P2_P3_U2715(p2_p3_u2715), .P2_P3_U2714(p2_p3_u2714), .P2_P3_U2713(p2_p3_u2713), .P2_P3_U2712(p2_p3_u2712), .P2_P3_U2711(p2_p3_u2711), .P2_P3_U2710(p2_p3_u2710), .P2_P3_U2709(p2_p3_u2709), .P2_P3_U2708(p2_p3_u2708), .P2_P3_U2707(p2_p3_u2707), .P2_P3_U2706(p2_p3_u2706), .P2_P3_U2705(p2_p3_u2705), .P2_P3_U2704(p2_p3_u2704), .P2_P3_U2703(p2_p3_u2703), .P2_P3_U2702(p2_p3_u2702), .P2_P3_U2701(p2_p3_u2701), .P2_P3_U2700(p2_p3_u2700), .P2_P3_U2699(p2_p3_u2699), .P2_P3_U2698(p2_p3_u2698), .P2_P3_U2697(p2_p3_u2697), .P2_P3_U2696(p2_p3_u2696), .P2_P3_U2695(p2_p3_u2695), .P2_P3_U2694(p2_p3_u2694), .P2_P3_U2693(p2_p3_u2693), .P2_P3_U2692(p2_p3_u2692), .P2_P3_U2691(p2_p3_u2691), .P2_P3_U2690(p2_p3_u2690), .P2_P3_U2689(p2_p3_u2689), .P2_P3_U2688(p2_p3_u2688), .P2_P3_U2687(p2_p3_u2687), .P2_P3_U2686(p2_p3_u2686), .P2_P3_U2685(p2_p3_u2685), .P2_P3_U2684(p2_p3_u2684), .P2_P3_U2683(p2_p3_u2683), .P2_P3_U2682(p2_p3_u2682), .P2_P3_U2681(p2_p3_u2681), .P2_P3_U2680(p2_p3_u2680), .P2_P3_U2679(p2_p3_u2679), .P2_P3_U2678(p2_p3_u2678), .P2_P3_U2677(p2_p3_u2677), .P2_P3_U2676(p2_p3_u2676), .P2_P3_U2675(p2_p3_u2675), .P2_P3_U2674(p2_p3_u2674), .P2_P3_U2673(p2_p3_u2673), .P2_P3_U2672(p2_p3_u2672), .P2_P3_U2671(p2_p3_u2671), .P2_P3_U2670(p2_p3_u2670), .P2_P3_U2669(p2_p3_u2669), .P2_P3_U2668(p2_p3_u2668), .P2_P3_U2667(p2_p3_u2667), .P2_P3_U2666(p2_p3_u2666), .P2_P3_U2665(p2_p3_u2665), .P2_P3_U2664(p2_p3_u2664), .P2_P3_U2663(p2_p3_u2663), .P2_P3_U2662(p2_p3_u2662), .P2_P3_U2661(p2_p3_u2661), .P2_P3_U2660(p2_p3_u2660), .P2_P3_U2659(p2_p3_u2659), .P2_P3_U2658(p2_p3_u2658), .P2_P3_U2657(p2_p3_u2657), .P2_P3_U2656(p2_p3_u2656), .P2_P3_U2655(p2_p3_u2655), .P2_P3_U2654(p2_p3_u2654), .P2_P3_U2653(p2_p3_u2653), .P2_P3_U2652(p2_p3_u2652), .P2_P3_U2651(p2_p3_u2651), .P2_P3_U2650(p2_p3_u2650), .P2_P3_U2649(p2_p3_u2649), .P2_P3_U2648(p2_p3_u2648), .P2_P3_U2647(p2_p3_u2647), .P2_P3_U2646(p2_p3_u2646), .P2_P3_U2645(p2_p3_u2645), .P2_P3_U2644(p2_p3_u2644), .P2_P3_U2643(p2_p3_u2643), .P2_P3_U2642(p2_p3_u2642), .P2_P3_U2641(p2_p3_u2641), .P2_P3_U2640(p2_p3_u2640), .P2_P3_U2639(p2_p3_u2639), .P2_P3_U3292(p2_p3_u3292), .P2_P3_U2638(p2_p3_u2638), .P2_P3_U3293(p2_p3_u3293), .P2_P3_U3294(p2_p3_u3294), .P2_P3_U2637(p2_p3_u2637), .P2_P3_U3295(p2_p3_u3295), .P2_P3_U2636(p2_p3_u2636), .P2_P3_U3296(p2_p3_u3296), .P2_P3_U2635(p2_p3_u2635), .P2_P3_U3297(p2_p3_u3297), .P2_P3_U2634(p2_p3_u2634), .P2_P3_U2633(p2_p3_u2633), .P2_P3_U3298(p2_p3_u3298), .P2_P3_U3299(p2_p3_u3299), .P2_P2_U3274(p2_p2_u3274), .P2_P2_U3275(p2_p2_u3275), .P2_P2_U3276(p2_p2_u3276), .P2_P2_U3277(p2_p2_u3277), .P2_P2_U3061(p2_p2_u3061), .P2_P2_U3060(p2_p2_u3060), .P2_P2_U3059(p2_p2_u3059), .P2_P2_U3058(p2_p2_u3058), .P2_P2_U3057(p2_p2_u3057), .P2_P2_U3056(p2_p2_u3056), .P2_P2_U3055(p2_p2_u3055), .P2_P2_U3054(p2_p2_u3054), .P2_P2_U3053(p2_p2_u3053), .P2_P2_U3052(p2_p2_u3052), .P2_P2_U3051(p2_p2_u3051), .P2_P2_U3050(p2_p2_u3050), .P2_P2_U3049(p2_p2_u3049), .P2_P2_U3048(p2_p2_u3048), .P2_P2_U3047(p2_p2_u3047), .P2_P2_U3046(p2_p2_u3046), .P2_P2_U3045(p2_p2_u3045), .P2_P2_U3044(p2_p2_u3044), .P2_P2_U3043(p2_p2_u3043), .P2_P2_U3042(p2_p2_u3042), .P2_P2_U3041(p2_p2_u3041), .P2_P2_U3040(p2_p2_u3040), .P2_P2_U3039(p2_p2_u3039), .P2_P2_U3038(p2_p2_u3038), .P2_P2_U3037(p2_p2_u3037), .P2_P2_U3036(p2_p2_u3036), .P2_P2_U3035(p2_p2_u3035), .P2_P2_U3034(p2_p2_u3034), .P2_P2_U3033(p2_p2_u3033), .P2_P2_U3032(p2_p2_u3032), .P2_P2_U3031(p2_p2_u3031), .P2_P2_U3030(p2_p2_u3030), .P2_P2_U3029(p2_p2_u3029), .P2_P2_U3280(p2_p2_u3280), .P2_P2_U3281(p2_p2_u3281), .P2_P2_U3028(p2_p2_u3028), .P2_P2_U3027(p2_p2_u3027), .P2_P2_U3026(p2_p2_u3026), .P2_P2_U3025(p2_p2_u3025), .P2_P2_U3024(p2_p2_u3024), .P2_P2_U3023(p2_p2_u3023), .P2_P2_U3022(p2_p2_u3022), .P2_P2_U3021(p2_p2_u3021), .P2_P2_U3020(p2_p2_u3020), .P2_P2_U3019(p2_p2_u3019), .P2_P2_U3018(p2_p2_u3018), .P2_P2_U3017(p2_p2_u3017), .P2_P2_U3016(p2_p2_u3016), .P2_P2_U3015(p2_p2_u3015), .P2_P2_U3014(p2_p2_u3014), .P2_P2_U3013(p2_p2_u3013), .P2_P2_U3012(p2_p2_u3012), .P2_P2_U3011(p2_p2_u3011), .P2_P2_U3010(p2_p2_u3010), .P2_P2_U3009(p2_p2_u3009), .P2_P2_U3008(p2_p2_u3008), .P2_P2_U3007(p2_p2_u3007), .P2_P2_U3006(p2_p2_u3006), .P2_P2_U3005(p2_p2_u3005), .P2_P2_U3004(p2_p2_u3004), .P2_P2_U3003(p2_p2_u3003), .P2_P2_U3002(p2_p2_u3002), .P2_P2_U3001(p2_p2_u3001), .P2_P2_U3000(p2_p2_u3000), .P2_P2_U2999(p2_p2_u2999), .P2_P2_U3282(p2_p2_u3282), .P2_P2_U2998(p2_p2_u2998), .P2_P2_U2997(p2_p2_u2997), .P2_P2_U2996(p2_p2_u2996), .P2_P2_U2995(p2_p2_u2995), .P2_P2_U2994(p2_p2_u2994), .P2_P2_U2993(p2_p2_u2993), .P2_P2_U2992(p2_p2_u2992), .P2_P2_U2991(p2_p2_u2991), .P2_P2_U2990(p2_p2_u2990), .P2_P2_U2989(p2_p2_u2989), .P2_P2_U2988(p2_p2_u2988), .P2_P2_U2987(p2_p2_u2987), .P2_P2_U2986(p2_p2_u2986), .P2_P2_U2985(p2_p2_u2985), .P2_P2_U2984(p2_p2_u2984), .P2_P2_U2983(p2_p2_u2983), .P2_P2_U2982(p2_p2_u2982), .P2_P2_U2981(p2_p2_u2981), .P2_P2_U2980(p2_p2_u2980), .P2_P2_U2979(p2_p2_u2979), .P2_P2_U2978(p2_p2_u2978), .P2_P2_U2977(p2_p2_u2977), .P2_P2_U2976(p2_p2_u2976), .P2_P2_U2975(p2_p2_u2975), .P2_P2_U2974(p2_p2_u2974), .P2_P2_U2973(p2_p2_u2973), .P2_P2_U2972(p2_p2_u2972), .P2_P2_U2971(p2_p2_u2971), .P2_P2_U2970(p2_p2_u2970), .P2_P2_U2969(p2_p2_u2969), .P2_P2_U2968(p2_p2_u2968), .P2_P2_U2967(p2_p2_u2967), .P2_P2_U2966(p2_p2_u2966), .P2_P2_U2965(p2_p2_u2965), .P2_P2_U2964(p2_p2_u2964), .P2_P2_U2963(p2_p2_u2963), .P2_P2_U2962(p2_p2_u2962), .P2_P2_U2961(p2_p2_u2961), .P2_P2_U2960(p2_p2_u2960), .P2_P2_U2959(p2_p2_u2959), .P2_P2_U2958(p2_p2_u2958), .P2_P2_U2957(p2_p2_u2957), .P2_P2_U2956(p2_p2_u2956), .P2_P2_U2955(p2_p2_u2955), .P2_P2_U2954(p2_p2_u2954), .P2_P2_U2953(p2_p2_u2953), .P2_P2_U2952(p2_p2_u2952), .P2_P2_U2951(p2_p2_u2951), .P2_P2_U2950(p2_p2_u2950), .P2_P2_U2949(p2_p2_u2949), .P2_P2_U2948(p2_p2_u2948), .P2_P2_U2947(p2_p2_u2947), .P2_P2_U2946(p2_p2_u2946), .P2_P2_U2945(p2_p2_u2945), .P2_P2_U2944(p2_p2_u2944), .P2_P2_U2943(p2_p2_u2943), .P2_P2_U2942(p2_p2_u2942), .P2_P2_U2941(p2_p2_u2941), .P2_P2_U2940(p2_p2_u2940), .P2_P2_U2939(p2_p2_u2939), .P2_P2_U2938(p2_p2_u2938), .P2_P2_U2937(p2_p2_u2937), .P2_P2_U2936(p2_p2_u2936), .P2_P2_U2935(p2_p2_u2935), .P2_P2_U2934(p2_p2_u2934), .P2_P2_U2933(p2_p2_u2933), .P2_P2_U2932(p2_p2_u2932), .P2_P2_U2931(p2_p2_u2931), .P2_P2_U2930(p2_p2_u2930), .P2_P2_U2929(p2_p2_u2929), .P2_P2_U2928(p2_p2_u2928), .P2_P2_U2927(p2_p2_u2927), .P2_P2_U2926(p2_p2_u2926), .P2_P2_U2925(p2_p2_u2925), .P2_P2_U2924(p2_p2_u2924), .P2_P2_U2923(p2_p2_u2923), .P2_P2_U2922(p2_p2_u2922), .P2_P2_U2921(p2_p2_u2921), .P2_P2_U2920(p2_p2_u2920), .P2_P2_U2919(p2_p2_u2919), .P2_P2_U2918(p2_p2_u2918), .P2_P2_U2917(p2_p2_u2917), .P2_P2_U2916(p2_p2_u2916), .P2_P2_U2915(p2_p2_u2915), .P2_P2_U2914(p2_p2_u2914), .P2_P2_U2913(p2_p2_u2913), .P2_P2_U2912(p2_p2_u2912), .P2_P2_U2911(p2_p2_u2911), .P2_P2_U2910(p2_p2_u2910), .P2_P2_U2909(p2_p2_u2909), .P2_P2_U2908(p2_p2_u2908), .P2_P2_U2907(p2_p2_u2907), .P2_P2_U2906(p2_p2_u2906), .P2_P2_U2905(p2_p2_u2905), .P2_P2_U2904(p2_p2_u2904), .P2_P2_U2903(p2_p2_u2903), .P2_P2_U2902(p2_p2_u2902), .P2_P2_U2901(p2_p2_u2901), .P2_P2_U2900(p2_p2_u2900), .P2_P2_U2899(p2_p2_u2899), .P2_P2_U2898(p2_p2_u2898), .P2_P2_U2897(p2_p2_u2897), .P2_P2_U2896(p2_p2_u2896), .P2_P2_U2895(p2_p2_u2895), .P2_P2_U2894(p2_p2_u2894), .P2_P2_U2893(p2_p2_u2893), .P2_P2_U2892(p2_p2_u2892), .P2_P2_U2891(p2_p2_u2891), .P2_P2_U2890(p2_p2_u2890), .P2_P2_U2889(p2_p2_u2889), .P2_P2_U2888(p2_p2_u2888), .P2_P2_U2887(p2_p2_u2887), .P2_P2_U2886(p2_p2_u2886), .P2_P2_U2885(p2_p2_u2885), .P2_P2_U2884(p2_p2_u2884), .P2_P2_U2883(p2_p2_u2883), .P2_P2_U2882(p2_p2_u2882), .P2_P2_U2881(p2_p2_u2881), .P2_P2_U2880(p2_p2_u2880), .P2_P2_U2879(p2_p2_u2879), .P2_P2_U2878(p2_p2_u2878), .P2_P2_U2877(p2_p2_u2877), .P2_P2_U2876(p2_p2_u2876), .P2_P2_U2875(p2_p2_u2875), .P2_P2_U2874(p2_p2_u2874), .P2_P2_U2873(p2_p2_u2873), .P2_P2_U2872(p2_p2_u2872), .P2_P2_U2871(p2_p2_u2871), .P2_P2_U2870(p2_p2_u2870), .P2_P2_U2869(p2_p2_u2869), .P2_P2_U2868(p2_p2_u2868), .P2_P2_U3284(p2_p2_u3284), .P2_P2_U3285(p2_p2_u3285), .P2_P2_U3288(p2_p2_u3288), .P2_P2_U3289(p2_p2_u3289), .P2_P2_U3290(p2_p2_u3290), .P2_P2_U2867(p2_p2_u2867), .P2_P2_U2866(p2_p2_u2866), .P2_P2_U2865(p2_p2_u2865), .P2_P2_U2864(p2_p2_u2864), .P2_P2_U2863(p2_p2_u2863), .P2_P2_U2862(p2_p2_u2862), .P2_P2_U2861(p2_p2_u2861), .P2_P2_U2860(p2_p2_u2860), .P2_P2_U2859(p2_p2_u2859), .P2_P2_U2858(p2_p2_u2858), .P2_P2_U2857(p2_p2_u2857), .P2_P2_U2856(p2_p2_u2856), .P2_P2_U2855(p2_p2_u2855), .P2_P2_U2854(p2_p2_u2854), .P2_P2_U2853(p2_p2_u2853), .P2_P2_U2852(p2_p2_u2852), .P2_P2_U2851(p2_p2_u2851), .P2_P2_U2850(p2_p2_u2850), .P2_P2_U2849(p2_p2_u2849), .P2_P2_U2848(p2_p2_u2848), .P2_P2_U2847(p2_p2_u2847), .P2_P2_U2846(p2_p2_u2846), .P2_P2_U2845(p2_p2_u2845), .P2_P2_U2844(p2_p2_u2844), .P2_P2_U2843(p2_p2_u2843), .P2_P2_U2842(p2_p2_u2842), .P2_P2_U2841(p2_p2_u2841), .P2_P2_U2840(p2_p2_u2840), .P2_P2_U2839(p2_p2_u2839), .P2_P2_U2838(p2_p2_u2838), .P2_P2_U2837(p2_p2_u2837), .P2_P2_U2836(p2_p2_u2836), .P2_P2_U2835(p2_p2_u2835), .P2_P2_U2834(p2_p2_u2834), .P2_P2_U2833(p2_p2_u2833), .P2_P2_U2832(p2_p2_u2832), .P2_P2_U2831(p2_p2_u2831), .P2_P2_U2830(p2_p2_u2830), .P2_P2_U2829(p2_p2_u2829), .P2_P2_U2828(p2_p2_u2828), .P2_P2_U2827(p2_p2_u2827), .P2_P2_U2826(p2_p2_u2826), .P2_P2_U2825(p2_p2_u2825), .P2_P2_U2824(p2_p2_u2824), .P2_P2_U2823(p2_p2_u2823), .P2_P2_U2822(p2_p2_u2822), .P2_P2_U2821(p2_p2_u2821), .P2_P2_U2820(p2_p2_u2820), .P2_P2_U2819(p2_p2_u2819), .P2_P2_U2818(p2_p2_u2818), .P2_P2_U2817(p2_p2_u2817), .P2_P2_U2816(p2_p2_u2816), .P2_P2_U2815(p2_p2_u2815), .P2_P2_U2814(p2_p2_u2814), .P2_P2_U2813(p2_p2_u2813), .P2_P2_U2812(p2_p2_u2812), .P2_P2_U2811(p2_p2_u2811), .P2_P2_U2810(p2_p2_u2810), .P2_P2_U2809(p2_p2_u2809), .P2_P2_U2808(p2_p2_u2808), .P2_P2_U2807(p2_p2_u2807), .P2_P2_U2806(p2_p2_u2806), .P2_P2_U2805(p2_p2_u2805), .P2_P2_U2804(p2_p2_u2804), .P2_P2_U2803(p2_p2_u2803), .P2_P2_U2802(p2_p2_u2802), .P2_P2_U2801(p2_p2_u2801), .P2_P2_U2800(p2_p2_u2800), .P2_P2_U2799(p2_p2_u2799), .P2_P2_U2798(p2_p2_u2798), .P2_P2_U2797(p2_p2_u2797), .P2_P2_U2796(p2_p2_u2796), .P2_P2_U2795(p2_p2_u2795), .P2_P2_U2794(p2_p2_u2794), .P2_P2_U2793(p2_p2_u2793), .P2_P2_U2792(p2_p2_u2792), .P2_P2_U2791(p2_p2_u2791), .P2_P2_U2790(p2_p2_u2790), .P2_P2_U2789(p2_p2_u2789), .P2_P2_U2788(p2_p2_u2788), .P2_P2_U2787(p2_p2_u2787), .P2_P2_U2786(p2_p2_u2786), .P2_P2_U2785(p2_p2_u2785), .P2_P2_U2784(p2_p2_u2784), .P2_P2_U2783(p2_p2_u2783), .P2_P2_U2782(p2_p2_u2782), .P2_P2_U2781(p2_p2_u2781), .P2_P2_U2780(p2_p2_u2780), .P2_P2_U2779(p2_p2_u2779), .P2_P2_U2778(p2_p2_u2778), .P2_P2_U2777(p2_p2_u2777), .P2_P2_U2776(p2_p2_u2776), .P2_P2_U2775(p2_p2_u2775), .P2_P2_U2774(p2_p2_u2774), .P2_P2_U2773(p2_p2_u2773), .P2_P2_U2772(p2_p2_u2772), .P2_P2_U2771(p2_p2_u2771), .P2_P2_U2770(p2_p2_u2770), .P2_P2_U2769(p2_p2_u2769), .P2_P2_U2768(p2_p2_u2768), .P2_P2_U2767(p2_p2_u2767), .P2_P2_U2766(p2_p2_u2766), .P2_P2_U2765(p2_p2_u2765), .P2_P2_U2764(p2_p2_u2764), .P2_P2_U2763(p2_p2_u2763), .P2_P2_U2762(p2_p2_u2762), .P2_P2_U2761(p2_p2_u2761), .P2_P2_U2760(p2_p2_u2760), .P2_P2_U2759(p2_p2_u2759), .P2_P2_U2758(p2_p2_u2758), .P2_P2_U2757(p2_p2_u2757), .P2_P2_U2756(p2_p2_u2756), .P2_P2_U2755(p2_p2_u2755), .P2_P2_U2754(p2_p2_u2754), .P2_P2_U2753(p2_p2_u2753), .P2_P2_U2752(p2_p2_u2752), .P2_P2_U2751(p2_p2_u2751), .P2_P2_U2750(p2_p2_u2750), .P2_P2_U2749(p2_p2_u2749), .P2_P2_U2748(p2_p2_u2748), .P2_P2_U2747(p2_p2_u2747), .P2_P2_U2746(p2_p2_u2746), .P2_P2_U2745(p2_p2_u2745), .P2_P2_U2744(p2_p2_u2744), .P2_P2_U2743(p2_p2_u2743), .P2_P2_U2742(p2_p2_u2742), .P2_P2_U2741(p2_p2_u2741), .P2_P2_U2740(p2_p2_u2740), .P2_P2_U2739(p2_p2_u2739), .P2_P2_U2738(p2_p2_u2738), .P2_P2_U2737(p2_p2_u2737), .P2_P2_U2736(p2_p2_u2736), .P2_P2_U2735(p2_p2_u2735), .P2_P2_U2734(p2_p2_u2734), .P2_P2_U2733(p2_p2_u2733), .P2_P2_U2732(p2_p2_u2732), .P2_P2_U2731(p2_p2_u2731), .P2_P2_U2730(p2_p2_u2730), .P2_P2_U2729(p2_p2_u2729), .P2_P2_U2728(p2_p2_u2728), .P2_P2_U2727(p2_p2_u2727), .P2_P2_U2726(p2_p2_u2726), .P2_P2_U2725(p2_p2_u2725), .P2_P2_U2724(p2_p2_u2724), .P2_P2_U2723(p2_p2_u2723), .P2_P2_U2722(p2_p2_u2722), .P2_P2_U2721(p2_p2_u2721), .P2_P2_U2720(p2_p2_u2720), .P2_P2_U2719(p2_p2_u2719), .P2_P2_U2718(p2_p2_u2718), .P2_P2_U2717(p2_p2_u2717), .P2_P2_U2716(p2_p2_u2716), .P2_P2_U2715(p2_p2_u2715), .P2_P2_U2714(p2_p2_u2714), .P2_P2_U2713(p2_p2_u2713), .P2_P2_U2712(p2_p2_u2712), .P2_P2_U2711(p2_p2_u2711), .P2_P2_U2710(p2_p2_u2710), .P2_P2_U2709(p2_p2_u2709), .P2_P2_U2708(p2_p2_u2708), .P2_P2_U2707(p2_p2_u2707), .P2_P2_U2706(p2_p2_u2706), .P2_P2_U2705(p2_p2_u2705), .P2_P2_U2704(p2_p2_u2704), .P2_P2_U2703(p2_p2_u2703), .P2_P2_U2702(p2_p2_u2702), .P2_P2_U2701(p2_p2_u2701), .P2_P2_U2700(p2_p2_u2700), .P2_P2_U2699(p2_p2_u2699), .P2_P2_U2698(p2_p2_u2698), .P2_P2_U2697(p2_p2_u2697), .P2_P2_U2696(p2_p2_u2696), .P2_P2_U2695(p2_p2_u2695), .P2_P2_U2694(p2_p2_u2694), .P2_P2_U2693(p2_p2_u2693), .P2_P2_U2692(p2_p2_u2692), .P2_P2_U2691(p2_p2_u2691), .P2_P2_U2690(p2_p2_u2690), .P2_P2_U2689(p2_p2_u2689), .P2_P2_U2688(p2_p2_u2688), .P2_P2_U2687(p2_p2_u2687), .P2_P2_U2686(p2_p2_u2686), .P2_P2_U2685(p2_p2_u2685), .P2_P2_U2684(p2_p2_u2684), .P2_P2_U2683(p2_p2_u2683), .P2_P2_U2682(p2_p2_u2682), .P2_P2_U2681(p2_p2_u2681), .P2_P2_U2680(p2_p2_u2680), .P2_P2_U2679(p2_p2_u2679), .P2_P2_U2678(p2_p2_u2678), .P2_P2_U2677(p2_p2_u2677), .P2_P2_U2676(p2_p2_u2676), .P2_P2_U2675(p2_p2_u2675), .P2_P2_U2674(p2_p2_u2674), .P2_P2_U2673(p2_p2_u2673), .P2_P2_U2672(p2_p2_u2672), .P2_P2_U2671(p2_p2_u2671), .P2_P2_U2670(p2_p2_u2670), .P2_P2_U2669(p2_p2_u2669), .P2_P2_U2668(p2_p2_u2668), .P2_P2_U2667(p2_p2_u2667), .P2_P2_U2666(p2_p2_u2666), .P2_P2_U2665(p2_p2_u2665), .P2_P2_U2664(p2_p2_u2664), .P2_P2_U2663(p2_p2_u2663), .P2_P2_U2662(p2_p2_u2662), .P2_P2_U2661(p2_p2_u2661), .P2_P2_U2660(p2_p2_u2660), .P2_P2_U2659(p2_p2_u2659), .P2_P2_U2658(p2_p2_u2658), .P2_P2_U2657(p2_p2_u2657), .P2_P2_U2656(p2_p2_u2656), .P2_P2_U2655(p2_p2_u2655), .P2_P2_U2654(p2_p2_u2654), .P2_P2_U2653(p2_p2_u2653), .P2_P2_U2652(p2_p2_u2652), .P2_P2_U2651(p2_p2_u2651), .P2_P2_U2650(p2_p2_u2650), .P2_P2_U2649(p2_p2_u2649), .P2_P2_U2648(p2_p2_u2648), .P2_P2_U2647(p2_p2_u2647), .P2_P2_U2646(p2_p2_u2646), .P2_P2_U2645(p2_p2_u2645), .P2_P2_U2644(p2_p2_u2644), .P2_P2_U2643(p2_p2_u2643), .P2_P2_U2642(p2_p2_u2642), .P2_P2_U2641(p2_p2_u2641), .P2_P2_U2640(p2_p2_u2640), .P2_P2_U2639(p2_p2_u2639), .P2_P2_U3292(p2_p2_u3292), .P2_P2_U2638(p2_p2_u2638), .P2_P2_U3293(p2_p2_u3293), .P2_P2_U3294(p2_p2_u3294), .P2_P2_U2637(p2_p2_u2637), .P2_P2_U3295(p2_p2_u3295), .P2_P2_U2636(p2_p2_u2636), .P2_P2_U3296(p2_p2_u3296), .P2_P2_U2635(p2_p2_u2635), .P2_P2_U3297(p2_p2_u3297), .P2_P2_U2634(p2_p2_u2634), .P2_P2_U2633(p2_p2_u2633), .P2_P2_U3298(p2_p2_u3298), .P2_P2_U3299(p2_p2_u3299), .P2_P1_U3288(p2_p1_u3288), .P2_P1_U3289(p2_p1_u3289), .P2_P1_U3290(p2_p1_u3290), .P2_P1_U3291(p2_p1_u3291), .P2_P1_U3077(p2_p1_u3077), .P2_P1_U3076(p2_p1_u3076), .P2_P1_U3075(p2_p1_u3075), .P2_P1_U3074(p2_p1_u3074), .P2_P1_U3073(p2_p1_u3073), .P2_P1_U3072(p2_p1_u3072), .P2_P1_U3071(p2_p1_u3071), .P2_P1_U3070(p2_p1_u3070), .P2_P1_U3069(p2_p1_u3069), .P2_P1_U3068(p2_p1_u3068), .P2_P1_U3067(p2_p1_u3067), .P2_P1_U3066(p2_p1_u3066), .P2_P1_U3065(p2_p1_u3065), .P2_P1_U3064(p2_p1_u3064), .P2_P1_U3063(p2_p1_u3063), .P2_P1_U3062(p2_p1_u3062), .P2_P1_U3061(p2_p1_u3061), .P2_P1_U3060(p2_p1_u3060), .P2_P1_U3059(p2_p1_u3059), .P2_P1_U3058(p2_p1_u3058), .P2_P1_U3057(p2_p1_u3057), .P2_P1_U3056(p2_p1_u3056), .P2_P1_U3055(p2_p1_u3055), .P2_P1_U3054(p2_p1_u3054), .P2_P1_U3053(p2_p1_u3053), .P2_P1_U3052(p2_p1_u3052), .P2_P1_U3051(p2_p1_u3051), .P2_P1_U3050(p2_p1_u3050), .P2_P1_U3049(p2_p1_u3049), .P2_P1_U3048(p2_p1_u3048), .P2_P1_U3047(p2_p1_u3047), .P2_P1_U3046(p2_p1_u3046), .P2_P1_U3045(p2_p1_u3045), .P2_P1_U3294(p2_p1_u3294), .P2_P1_U3295(p2_p1_u3295), .P2_P1_U3044(p2_p1_u3044), .P2_P1_U3043(p2_p1_u3043), .P2_P1_U3042(p2_p1_u3042), .P2_P1_U3041(p2_p1_u3041), .P2_P1_U3040(p2_p1_u3040), .P2_P1_U3039(p2_p1_u3039), .P2_P1_U3038(p2_p1_u3038), .P2_P1_U3037(p2_p1_u3037), .P2_P1_U3036(p2_p1_u3036), .P2_P1_U3035(p2_p1_u3035), .P2_P1_U3034(p2_p1_u3034), .P2_P1_U3033(p2_p1_u3033), .P2_P1_U3032(p2_p1_u3032), .P2_P1_U3031(p2_p1_u3031), .P2_P1_U3030(p2_p1_u3030), .P2_P1_U3029(p2_p1_u3029), .P2_P1_U3028(p2_p1_u3028), .P2_P1_U3027(p2_p1_u3027), .P2_P1_U3026(p2_p1_u3026), .P2_P1_U3025(p2_p1_u3025), .P2_P1_U3024(p2_p1_u3024), .P2_P1_U3023(p2_p1_u3023), .P2_P1_U3022(p2_p1_u3022), .P2_P1_U3021(p2_p1_u3021), .P2_P1_U3020(p2_p1_u3020), .P2_P1_U3019(p2_p1_u3019), .P2_P1_U3018(p2_p1_u3018), .P2_P1_U3017(p2_p1_u3017), .P2_P1_U3016(p2_p1_u3016), .P2_P1_U3015(p2_p1_u3015), .P2_P1_U3296(p2_p1_u3296), .P2_P1_U3014(p2_p1_u3014), .P2_P1_U3013(p2_p1_u3013), .P2_P1_U3012(p2_p1_u3012), .P2_P1_U3011(p2_p1_u3011), .P2_P1_U3010(p2_p1_u3010), .P2_P1_U3009(p2_p1_u3009), .P2_P1_U3008(p2_p1_u3008), .P2_P1_U3007(p2_p1_u3007), .P2_P1_U3006(p2_p1_u3006), .P2_P1_U3005(p2_p1_u3005), .P2_P1_U3004(p2_p1_u3004), .P2_P1_U3003(p2_p1_u3003), .P2_P1_U3002(p2_p1_u3002), .P2_P1_U3001(p2_p1_u3001), .P2_P1_U3000(p2_p1_u3000), .P2_P1_U2999(p2_p1_u2999), .P2_P1_U2998(p2_p1_u2998), .P2_P1_U2997(p2_p1_u2997), .P2_P1_U2996(p2_p1_u2996), .P2_P1_U2995(p2_p1_u2995), .P2_P1_U2994(p2_p1_u2994), .P2_P1_U2993(p2_p1_u2993), .P2_P1_U2992(p2_p1_u2992), .P2_P1_U2991(p2_p1_u2991), .P2_P1_U2990(p2_p1_u2990), .P2_P1_U2989(p2_p1_u2989), .P2_P1_U2988(p2_p1_u2988), .P2_P1_U2987(p2_p1_u2987), .P2_P1_U2986(p2_p1_u2986), .P2_P1_U2985(p2_p1_u2985), .P2_P1_U2984(p2_p1_u2984), .P2_P1_U2983(p2_p1_u2983), .P2_P1_U2982(p2_p1_u2982), .P2_P1_U2981(p2_p1_u2981), .P2_P1_U2980(p2_p1_u2980), .P2_P1_U2979(p2_p1_u2979), .P2_P1_U2978(p2_p1_u2978), .P2_P1_U2977(p2_p1_u2977), .P2_P1_U2976(p2_p1_u2976), .P2_P1_U2975(p2_p1_u2975), .P2_P1_U2974(p2_p1_u2974), .P2_P1_U2973(p2_p1_u2973), .P2_P1_U2972(p2_p1_u2972), .P2_P1_U2971(p2_p1_u2971), .P2_P1_U2970(p2_p1_u2970), .P2_P1_U2969(p2_p1_u2969), .P2_P1_U2968(p2_p1_u2968), .P2_P1_U2967(p2_p1_u2967), .P2_P1_U2966(p2_p1_u2966), .P2_P1_U2965(p2_p1_u2965), .P2_P1_U2964(p2_p1_u2964), .P2_P1_U2963(p2_p1_u2963), .P2_P1_U2962(p2_p1_u2962), .P2_P1_U2961(p2_p1_u2961), .P2_P1_U2960(p2_p1_u2960), .P2_P1_U2959(p2_p1_u2959), .P2_P1_U2958(p2_p1_u2958), .P2_P1_U2957(p2_p1_u2957), .P2_P1_U2956(p2_p1_u2956), .P2_P1_U2955(p2_p1_u2955), .P2_P1_U2954(p2_p1_u2954), .P2_P1_U2953(p2_p1_u2953), .P2_P1_U2952(p2_p1_u2952), .P2_P1_U2951(p2_p1_u2951), .P2_P1_U2950(p2_p1_u2950), .P2_P1_U2949(p2_p1_u2949), .P2_P1_U2948(p2_p1_u2948), .P2_P1_U2947(p2_p1_u2947), .P2_P1_U2946(p2_p1_u2946), .P2_P1_U2945(p2_p1_u2945), .P2_P1_U2944(p2_p1_u2944), .P2_P1_U2943(p2_p1_u2943), .P2_P1_U2942(p2_p1_u2942), .P2_P1_U2941(p2_p1_u2941), .P2_P1_U2940(p2_p1_u2940), .P2_P1_U2939(p2_p1_u2939), .P2_P1_U2938(p2_p1_u2938), .P2_P1_U2937(p2_p1_u2937), .P2_P1_U2936(p2_p1_u2936), .P2_P1_U2935(p2_p1_u2935), .P2_P1_U2934(p2_p1_u2934), .P2_P1_U2933(p2_p1_u2933), .P2_P1_U2932(p2_p1_u2932), .P2_P1_U2931(p2_p1_u2931), .P2_P1_U2930(p2_p1_u2930), .P2_P1_U2929(p2_p1_u2929), .P2_P1_U2928(p2_p1_u2928), .P2_P1_U2927(p2_p1_u2927), .P2_P1_U2926(p2_p1_u2926), .P2_P1_U2925(p2_p1_u2925), .P2_P1_U2924(p2_p1_u2924), .P2_P1_U2923(p2_p1_u2923), .P2_P1_U2922(p2_p1_u2922), .P2_P1_U2921(p2_p1_u2921), .P2_P1_U2920(p2_p1_u2920), .P2_P1_U2919(p2_p1_u2919), .P2_P1_U2918(p2_p1_u2918), .P2_P1_U2917(p2_p1_u2917), .P2_P1_U2916(p2_p1_u2916), .P2_P1_U2915(p2_p1_u2915), .P2_P1_U2914(p2_p1_u2914), .P2_P1_U2913(p2_p1_u2913), .P2_P1_U2912(p2_p1_u2912), .P2_P1_U2911(p2_p1_u2911), .P2_P1_U2910(p2_p1_u2910), .P2_P1_U2909(p2_p1_u2909), .P2_P1_U2908(p2_p1_u2908), .P2_P1_U2907(p2_p1_u2907), .P2_P1_U2906(p2_p1_u2906), .P2_P1_U2905(p2_p1_u2905), .P2_P1_U2904(p2_p1_u2904), .P2_P1_U2903(p2_p1_u2903), .P2_P1_U2902(p2_p1_u2902), .P2_P1_U2901(p2_p1_u2901), .P2_P1_U2900(p2_p1_u2900), .P2_P1_U2899(p2_p1_u2899), .P2_P1_U2898(p2_p1_u2898), .P2_P1_U2897(p2_p1_u2897), .P2_P1_U2896(p2_p1_u2896), .P2_P1_U2895(p2_p1_u2895), .P2_P1_U2894(p2_p1_u2894), .P2_P1_U2893(p2_p1_u2893), .P2_P1_U2892(p2_p1_u2892), .P2_P1_U2891(p2_p1_u2891), .P2_P1_U2890(p2_p1_u2890), .P2_P1_U2889(p2_p1_u2889), .P2_P1_U2888(p2_p1_u2888), .P2_P1_U2887(p2_p1_u2887), .P2_P1_U2886(p2_p1_u2886), .P2_P1_U2885(p2_p1_u2885), .P2_P1_U2884(p2_p1_u2884), .P2_P1_U3298(p2_p1_u3298), .P2_P1_U3299(p2_p1_u3299), .P2_P1_U3302(p2_p1_u3302), .P2_P1_U3303(p2_p1_u3303), .P2_P1_U3304(p2_p1_u3304), .P2_P1_U2883(p2_p1_u2883), .P2_P1_U2882(p2_p1_u2882), .P2_P1_U2881(p2_p1_u2881), .P2_P1_U2880(p2_p1_u2880), .P2_P1_U2879(p2_p1_u2879), .P2_P1_U2878(p2_p1_u2878), .P2_P1_U2877(p2_p1_u2877), .P2_P1_U2876(p2_p1_u2876), .P2_P1_U2875(p2_p1_u2875), .P2_P1_U2874(p2_p1_u2874), .P2_P1_U2873(p2_p1_u2873), .P2_P1_U2872(p2_p1_u2872), .P2_P1_U2871(p2_p1_u2871), .P2_P1_U2870(p2_p1_u2870), .P2_P1_U2869(p2_p1_u2869), .P2_P1_U2868(p2_p1_u2868), .P2_P1_U2867(p2_p1_u2867), .P2_P1_U2866(p2_p1_u2866), .P2_P1_U2865(p2_p1_u2865), .P2_P1_U2864(p2_p1_u2864), .P2_P1_U2863(p2_p1_u2863), .P2_P1_U2862(p2_p1_u2862), .P2_P1_U2861(p2_p1_u2861), .P2_P1_U2860(p2_p1_u2860), .P2_P1_U2859(p2_p1_u2859), .P2_P1_U2858(p2_p1_u2858), .P2_P1_U2857(p2_p1_u2857), .P2_P1_U2856(p2_p1_u2856), .P2_P1_U2855(p2_p1_u2855), .P2_P1_U2854(p2_p1_u2854), .P2_P1_U2853(p2_p1_u2853), .P2_P1_U2852(p2_p1_u2852), .P2_P1_U2851(p2_p1_u2851), .P2_P1_U2850(p2_p1_u2850), .P2_P1_U2849(p2_p1_u2849), .P2_P1_U2848(p2_p1_u2848), .P2_P1_U2847(p2_p1_u2847), .P2_P1_U2846(p2_p1_u2846), .P2_P1_U2845(p2_p1_u2845), .P2_P1_U2844(p2_p1_u2844), .P2_P1_U2843(p2_p1_u2843), .P2_P1_U2842(p2_p1_u2842), .P2_P1_U2841(p2_p1_u2841), .P2_P1_U2840(p2_p1_u2840), .P2_P1_U2839(p2_p1_u2839), .P2_P1_U2838(p2_p1_u2838), .P2_P1_U2837(p2_p1_u2837), .P2_P1_U2836(p2_p1_u2836), .P2_P1_U2835(p2_p1_u2835), .P2_P1_U2834(p2_p1_u2834), .P2_P1_U2833(p2_p1_u2833), .P2_P1_U2832(p2_p1_u2832), .P2_P1_U2831(p2_p1_u2831), .P2_P1_U2830(p2_p1_u2830), .P2_P1_U2829(p2_p1_u2829), .P2_P1_U2828(p2_p1_u2828), .P2_P1_U2827(p2_p1_u2827), .P2_P1_U2826(p2_p1_u2826), .P2_P1_U2825(p2_p1_u2825), .P2_P1_U2824(p2_p1_u2824), .P2_P1_U2823(p2_p1_u2823), .P2_P1_U2822(p2_p1_u2822), .P2_P1_U2821(p2_p1_u2821), .P2_P1_U2820(p2_p1_u2820), .P2_P1_U2819(p2_p1_u2819), .P2_P1_U2818(p2_p1_u2818), .P2_P1_U2817(p2_p1_u2817), .P2_P1_U2816(p2_p1_u2816), .P2_P1_U2815(p2_p1_u2815), .P2_P1_U2814(p2_p1_u2814), .P2_P1_U2813(p2_p1_u2813), .P2_P1_U2812(p2_p1_u2812), .P2_P1_U2811(p2_p1_u2811), .P2_P1_U2810(p2_p1_u2810), .P2_P1_U2809(p2_p1_u2809), .P2_P1_U2808(p2_p1_u2808), .P2_P1_U2807(p2_p1_u2807), .P2_P1_U2806(p2_p1_u2806), .P2_P1_U2805(p2_p1_u2805), .P2_P1_U2804(p2_p1_u2804), .P2_P1_U2803(p2_p1_u2803), .P2_P1_U2802(p2_p1_u2802), .P2_P1_U2801(p2_p1_u2801), .P2_P1_U2800(p2_p1_u2800), .P2_P1_U2799(p2_p1_u2799), .P2_P1_U2798(p2_p1_u2798), .P2_P1_U2797(p2_p1_u2797), .P2_P1_U2796(p2_p1_u2796), .P2_P1_U2795(p2_p1_u2795), .P2_P1_U2794(p2_p1_u2794), .P2_P1_U2793(p2_p1_u2793), .P2_P1_U2792(p2_p1_u2792), .P2_P1_U2791(p2_p1_u2791), .P2_P1_U2790(p2_p1_u2790), .P2_P1_U2789(p2_p1_u2789), .P2_P1_U2788(p2_p1_u2788), .P2_P1_U2787(p2_p1_u2787), .P2_P1_U2786(p2_p1_u2786), .P2_P1_U2785(p2_p1_u2785), .P2_P1_U2784(p2_p1_u2784), .P2_P1_U2783(p2_p1_u2783), .P2_P1_U2782(p2_p1_u2782), .P2_P1_U2781(p2_p1_u2781), .P2_P1_U2780(p2_p1_u2780), .P2_P1_U2779(p2_p1_u2779), .P2_P1_U2778(p2_p1_u2778), .P2_P1_U2777(p2_p1_u2777), .P2_P1_U2776(p2_p1_u2776), .P2_P1_U2775(p2_p1_u2775), .P2_P1_U2774(p2_p1_u2774), .P2_P1_U2773(p2_p1_u2773), .P2_P1_U2772(p2_p1_u2772), .P2_P1_U2771(p2_p1_u2771), .P2_P1_U2770(p2_p1_u2770), .P2_P1_U2769(p2_p1_u2769), .P2_P1_U2768(p2_p1_u2768), .P2_P1_U2767(p2_p1_u2767), .P2_P1_U2766(p2_p1_u2766), .P2_P1_U2765(p2_p1_u2765), .P2_P1_U2764(p2_p1_u2764), .P2_P1_U2763(p2_p1_u2763), .P2_P1_U2762(p2_p1_u2762), .P2_P1_U2761(p2_p1_u2761), .P2_P1_U2760(p2_p1_u2760), .P2_P1_U2759(p2_p1_u2759), .P2_P1_U2758(p2_p1_u2758), .P2_P1_U2757(p2_p1_u2757), .P2_P1_U2756(p2_p1_u2756), .P2_P1_U2755(p2_p1_u2755), .P2_P1_U2754(p2_p1_u2754), .P2_P1_U2753(p2_p1_u2753), .P2_P1_U2752(p2_p1_u2752), .P2_P1_U2751(p2_p1_u2751), .P2_P1_U2750(p2_p1_u2750), .P2_P1_U2749(p2_p1_u2749), .P2_P1_U2748(p2_p1_u2748), .P2_P1_U2747(p2_p1_u2747), .P2_P1_U2746(p2_p1_u2746), .P2_P1_U2745(p2_p1_u2745), .P2_P1_U2744(p2_p1_u2744), .P2_P1_U2743(p2_p1_u2743), .P2_P1_U2742(p2_p1_u2742), .P2_P1_U2741(p2_p1_u2741), .P2_P1_U2740(p2_p1_u2740), .P2_P1_U2739(p2_p1_u2739), .P2_P1_U2738(p2_p1_u2738), .P2_P1_U2737(p2_p1_u2737), .P2_P1_U2736(p2_p1_u2736), .P2_P1_U2735(p2_p1_u2735), .P2_P1_U2734(p2_p1_u2734), .P2_P1_U2733(p2_p1_u2733), .P2_P1_U2732(p2_p1_u2732), .P2_P1_U2731(p2_p1_u2731), .P2_P1_U2730(p2_p1_u2730), .P2_P1_U2729(p2_p1_u2729), .P2_P1_U2728(p2_p1_u2728), .P2_P1_U2727(p2_p1_u2727), .P2_P1_U2726(p2_p1_u2726), .P2_P1_U2725(p2_p1_u2725), .P2_P1_U2724(p2_p1_u2724), .P2_P1_U2723(p2_p1_u2723), .P2_P1_U2722(p2_p1_u2722), .P2_P1_U2721(p2_p1_u2721), .P2_P1_U2720(p2_p1_u2720), .P2_P1_U2719(p2_p1_u2719), .P2_P1_U2718(p2_p1_u2718), .P2_P1_U2717(p2_p1_u2717), .P2_P1_U2716(p2_p1_u2716), .P2_P1_U2715(p2_p1_u2715), .P2_P1_U2714(p2_p1_u2714), .P2_P1_U2713(p2_p1_u2713), .P2_P1_U2712(p2_p1_u2712), .P2_P1_U2711(p2_p1_u2711), .P2_P1_U2710(p2_p1_u2710), .P2_P1_U2709(p2_p1_u2709), .P2_P1_U2708(p2_p1_u2708), .P2_P1_U2707(p2_p1_u2707), .P2_P1_U2706(p2_p1_u2706), .P2_P1_U2705(p2_p1_u2705), .P2_P1_U2704(p2_p1_u2704), .P2_P1_U2703(p2_p1_u2703), .P2_P1_U2702(p2_p1_u2702), .P2_P1_U2701(p2_p1_u2701), .P2_P1_U2700(p2_p1_u2700), .P2_P1_U2699(p2_p1_u2699), .P2_P1_U2698(p2_p1_u2698), .P2_P1_U2697(p2_p1_u2697), .P2_P1_U2696(p2_p1_u2696), .P2_P1_U2695(p2_p1_u2695), .P2_P1_U2694(p2_p1_u2694), .P2_P1_U2693(p2_p1_u2693), .P2_P1_U2692(p2_p1_u2692), .P2_P1_U2691(p2_p1_u2691), .P2_P1_U2690(p2_p1_u2690), .P2_P1_U2689(p2_p1_u2689), .P2_P1_U2688(p2_p1_u2688), .P2_P1_U2687(p2_p1_u2687), .P2_P1_U2686(p2_p1_u2686), .P2_P1_U2685(p2_p1_u2685), .P2_P1_U2684(p2_p1_u2684), .P2_P1_U2683(p2_p1_u2683), .P2_P1_U2682(p2_p1_u2682), .P2_P1_U2681(p2_p1_u2681), .P2_P1_U2680(p2_p1_u2680), .P2_P1_U2679(p2_p1_u2679), .P2_P1_U2678(p2_p1_u2678), .P2_P1_U2677(p2_p1_u2677), .P2_P1_U2676(p2_p1_u2676), .P2_P1_U2675(p2_p1_u2675), .P2_P1_U2674(p2_p1_u2674), .P2_P1_U2673(p2_p1_u2673), .P2_P1_U2672(p2_p1_u2672), .P2_P1_U2671(p2_p1_u2671), .P2_P1_U2670(p2_p1_u2670), .P2_P1_U2669(p2_p1_u2669), .P2_P1_U2668(p2_p1_u2668), .P2_P1_U2667(p2_p1_u2667), .P2_P1_U2666(p2_p1_u2666), .P2_P1_U2665(p2_p1_u2665), .P2_P1_U2664(p2_p1_u2664), .P2_P1_U2663(p2_p1_u2663), .P2_P1_U2662(p2_p1_u2662), .P2_P1_U2661(p2_p1_u2661), .P2_P1_U2660(p2_p1_u2660), .P2_P1_U2659(p2_p1_u2659), .P2_P1_U2658(p2_p1_u2658), .P2_P1_U2657(p2_p1_u2657), .P2_P1_U2656(p2_p1_u2656), .P2_P1_U2655(p2_p1_u2655), .P2_P1_U3306(p2_p1_u3306), .P2_P1_U2654(p2_p1_u2654), .P2_P1_U3307(p2_p1_u3307), .P2_P1_U3308(p2_p1_u3308), .P2_P1_U2653(p2_p1_u2653), .P2_P1_U3309(p2_p1_u3309), .P2_P1_U2652(p2_p1_u2652), .P2_P1_U3310(p2_p1_u3310), .P2_P1_U2651(p2_p1_u2651), .P2_P1_U3311(p2_p1_u3311), .P2_P1_U2650(p2_p1_u2650), .P2_P1_U2649(p2_p1_u2649), .P2_P1_U3312(p2_p1_u3312), .P2_P1_U3313(p2_p1_u3313));

integer i=0;
always @ (posedge clk) begin
	vec = input_vec_mem[i];
	$monitor(vec);
	i = i + 1;

end

always @ (negedge clk)begin
	$fdisplay ( fh_w, logic0_po_extra, mul_1411_u378, mul_1411_u438, mul_1411_u10, mul_1411_u439, mul_1411_u9, mul_1411_u440, mul_1411_u8, mul_1411_u441, mul_1411_u7, mul_1411_u385, mul_1411_u14, mul_1411_u386, mul_1411_u13, mul_1411_u387, mul_1411_u12, mul_1411_u388, mul_1411_u11, mul_1411_u15, mul_1411_u5_po_extra, mul_1421_a1_u5, u154, u39_po_extra, p1_u247, p1_u246, p1_u245, p1_u244, p1_u243, p1_u242, p1_u241, p1_u240, p1_u239, p1_u238, p1_u237, p1_u236, p1_u235, p1_u234, p1_u233, p1_u232, p1_u231, p1_u230, p1_u229, p1_u228, p1_u227, p1_u226, p1_u225, p1_u224, p1_u223, p1_u222, p1_u221, p1_u220, p1_u219, p1_u218, p1_u217, p1_u216, p1_u251, p1_u252, p1_u253, p1_u254, p1_u255, p1_u256, p1_u257, p1_u258, p1_u259, p1_u260, p1_u261, p1_u262, p1_u263, p1_u264, p1_u265, p1_u266, p1_u267, p1_u268, p1_u269, p1_u270, p1_u271, p1_u272, p1_u273, p1_u274, p1_u275, p1_u276, p1_u277, p1_u278, p1_u279, p1_u280, p1_u281, p1_u282, p1_u212, p1_u215, p1_u213, p1_u214, p2_u247, p2_u246, p2_u245, p2_u244, p2_u243, p2_u242, p2_u241, p2_u240, p2_u239, p2_u238, p2_u237, p2_u236, p2_u235, p2_u234, p2_u233, p2_u232, p2_u231, p2_u230, p2_u229, p2_u228, p2_u227, p2_u226, p2_u225, p2_u224, p2_u223, p2_u222, p2_u221, p2_u220, p2_u219, p2_u218, p2_u217, p2_u216, p2_u251, p2_u252, p2_u253, p2_u254, p2_u255, p2_u256, p2_u257, p2_u258, p2_u259, p2_u260, p2_u261, p2_u262, p2_u263, p2_u264, p2_u265, p2_u266, p2_u267, p2_u268, p2_u269, p2_u270, p2_u271, p2_u272, p2_u273, p2_u274, p2_u275, p2_u276, p2_u277, p2_u278, p2_u279, p2_u280, p2_u281, p2_u282, p2_u212, p2_u215, p2_u213, p2_u214, p3_u3354, p3_u3353, p3_u3352, p3_u3351, p3_u3350, p3_u3349, p3_u3348, p3_u3347, p3_u3346, p3_u3345, p3_u3344, p3_u3343, p3_u3342, p3_u3341, p3_u3340, p3_u3339, p3_u3338, p3_u3337, p3_u3336, p3_u3335, p3_u3334, p3_u3333, p3_u3332, p3_u3331, p3_u3330, p3_u3329, p3_u3328, p3_u3327, p3_u3326, p3_u3325, p3_u3324, p3_u3323, p3_u3442, p3_u3443, p3_u3322, p3_u3321, p3_u3320, p3_u3319, p3_u3318, p3_u3317, p3_u3316, p3_u3315, p3_u3314, p3_u3313, p3_u3312, p3_u3311, p3_u3310, p3_u3309, p3_u3308, p3_u3307, p3_u3306, p3_u3305, p3_u3304, p3_u3303, p3_u3302, p3_u3301, p3_u3300, p3_u3299, p3_u3298, p3_u3297, p3_u3296, p3_u3295, p3_u3294, p3_u3293, p3_u3456, p3_u3459, p3_u3462, p3_u3465, p3_u3468, p3_u3471, p3_u3474, p3_u3477, p3_u3480, p3_u3483, p3_u3486, p3_u3489, p3_u3492, p3_u3495, p3_u3498, p3_u3501, p3_u3504, p3_u3507, p3_u3510, p3_u3512, p3_u3513, p3_u3514, p3_u3515, p3_u3516, p3_u3517, p3_u3518, p3_u3519, p3_u3520, p3_u3521, p3_u3522, p3_u3523, p3_u3524, p3_u3525, p3_u3526, p3_u3527, p3_u3528, p3_u3529, p3_u3530, p3_u3531, p3_u3532, p3_u3533, p3_u3534, p3_u3535, p3_u3536, p3_u3537, p3_u3538, p3_u3539, p3_u3540, p3_u3541, p3_u3542, p3_u3543, p3_u3544, p3_u3545, p3_u3546, p3_u3547, p3_u3548, p3_u3549, p3_u3550, p3_u3551, p3_u3552, p3_u3553, p3_u3554, p3_u3555, p3_u3556, p3_u3292, p3_u3291, p3_u3290, p3_u3289, p3_u3288, p3_u3287, p3_u3286, p3_u3285, p3_u3284, p3_u3283, p3_u3282, p3_u3281, p3_u3280, p3_u3279, p3_u3278, p3_u3277, p3_u3276, p3_u3275, p3_u3274, p3_u3273, p3_u3272, p3_u3271, p3_u3270, p3_u3269, p3_u3268, p3_u3267, p3_u3266, p3_u3265, p3_u3264, p3_u3263, p3_u3262, p3_u3261, p3_u3260, p3_u3259, p3_u3258, p3_u3257, p3_u3256, p3_u3255, p3_u3254, p3_u3253, p3_u3252, p3_u3251, p3_u3250, p3_u3249, p3_u3248, p3_u3247, p3_u3246, p3_u3245, p3_u3244, p3_u3243, p3_u3242, p3_u3241, p3_u3557, p3_u3558, p3_u3559, p3_u3560, p3_u3561, p3_u3562, p3_u3563, p3_u3564, p3_u3565, p3_u3566, p3_u3567, p3_u3568, p3_u3569, p3_u3570, p3_u3571, p3_u3572, p3_u3573, p3_u3574, p3_u3575, p3_u3576, p3_u3577, p3_u3578, p3_u3579, p3_u3580, p3_u3581, p3_u3582, p3_u3583, p3_u3584, p3_u3585, p3_u3586, p3_u3587, p3_u3588, p3_u3240, p3_u3239, p3_u3238, p3_u3237, p3_u3236, p3_u3235, p3_u3234, p3_u3233, p3_u3232, p3_u3231, p3_u3230, p3_u3229, p3_u3228, p3_u3227, p3_u3226, p3_u3225, p3_u3224, p3_u3223, p3_u3222, p3_u3221, p3_u3220, p3_u3219, p3_u3218, p3_u3217, p3_u3216, p3_u3215, p3_u3214, p3_u3213, p3_u3212, p3_u3211, p3_u3084, p3_u3083, p3_u4038, p4_u3351, p4_u3350, p4_u3349, p4_u3348, p4_u3347, p4_u3346, p4_u3345, p4_u3344, p4_u3343, p4_u3342, p4_u3341, p4_u3340, p4_u3339, p4_u3338, p4_u3337, p4_u3336, p4_u3335, p4_u3334, p4_u3333, p4_u3332, p4_u3331, p4_u3330, p4_u3329, p4_u3328, p4_u3327, p4_u3326, p4_u3325, p4_u3324, p4_u3323, p4_u3322, p4_u3321, p4_u3320, p4_u3437, p4_u3438, p4_u3319, p4_u3318, p4_u3317, p4_u3316, p4_u3315, p4_u3314, p4_u3313, p4_u3312, p4_u3311, p4_u3310, p4_u3309, p4_u3308, p4_u3307, p4_u3306, p4_u3305, p4_u3304, p4_u3303, p4_u3302, p4_u3301, p4_u3300, p4_u3299, p4_u3298, p4_u3297, p4_u3296, p4_u3295, p4_u3294, p4_u3293, p4_u3292, p4_u3291, p4_u3290, p4_u3451, p4_u3454, p4_u3457, p4_u3460, p4_u3463, p4_u3466, p4_u3469, p4_u3472, p4_u3475, p4_u3478, p4_u3481, p4_u3484, p4_u3487, p4_u3490, p4_u3493, p4_u3496, p4_u3499, p4_u3502, p4_u3505, p4_u3507, p4_u3508, p4_u3509, p4_u3510, p4_u3511, p4_u3512, p4_u3513, p4_u3514, p4_u3515, p4_u3516, p4_u3517, p4_u3518, p4_u3519, p4_u3520, p4_u3521, p4_u3522, p4_u3523, p4_u3524, p4_u3525, p4_u3526, p4_u3527, p4_u3528, p4_u3529, p4_u3530, p4_u3531, p4_u3532, p4_u3533, p4_u3534, p4_u3535, p4_u3536, p4_u3537, p4_u3538, p4_u3539, p4_u3540, p4_u3541, p4_u3542, p4_u3543, p4_u3544, p4_u3545, p4_u3546, p4_u3547, p4_u3548, p4_u3549, p4_u3550, p4_u3551, p4_u3289, p4_u3288, p4_u3287, p4_u3286, p4_u3285, p4_u3284, p4_u3283, p4_u3282, p4_u3281, p4_u3280, p4_u3279, p4_u3278, p4_u3277, p4_u3276, p4_u3275, p4_u3274, p4_u3273, p4_u3272, p4_u3271, p4_u3270, p4_u3269, p4_u3268, p4_u3267, p4_u3266, p4_u3265, p4_u3264, p4_u3263, p4_u3262, p4_u3261, p4_u3260, p4_u3259, p4_u3258, p4_u3257, p4_u3256, p4_u3255, p4_u3254, p4_u3253, p4_u3252, p4_u3251, p4_u3250, p4_u3249, p4_u3248, p4_u3247, p4_u3246, p4_u3245, p4_u3244, p4_u3243, p4_u3242, p4_u3241, p4_u3240, p4_u3239, p4_u3238, p4_u3552, p4_u3553, p4_u3554, p4_u3555, p4_u3556, p4_u3557, p4_u3558, p4_u3559, p4_u3560, p4_u3561, p4_u3562, p4_u3563, p4_u3564, p4_u3565, p4_u3566, p4_u3567, p4_u3568, p4_u3569, p4_u3570, p4_u3571, p4_u3572, p4_u3573, p4_u3574, p4_u3575, p4_u3576, p4_u3577, p4_u3578, p4_u3579, p4_u3580, p4_u3581, p4_u3582, p4_u3583, p4_u3237, p4_u3236, p4_u3235, p4_u3234, p4_u3233, p4_u3232, p4_u3231, p4_u3230, p4_u3229, p4_u3228, p4_u3227, p4_u3226, p4_u3225, p4_u3224, p4_u3223, p4_u3222, p4_u3221, p4_u3220, p4_u3219, p4_u3218, p4_u3217, p4_u3216, p4_u3215, p4_u3214, p4_u3213, p4_u3212, p4_u3211, p4_u3210, p4_u3209, p4_u3208, p4_u3147, p4_u3146, p4_u4028, p1_p3_u3274, p1_p3_u3275, p1_p3_u3276, p1_p3_u3277, p1_p3_u3061, p1_p3_u3060, p1_p3_u3059, p1_p3_u3058, p1_p3_u3057, p1_p3_u3056, p1_p3_u3055, p1_p3_u3054, p1_p3_u3053, p1_p3_u3052, p1_p3_u3051, p1_p3_u3050, p1_p3_u3049, p1_p3_u3048, p1_p3_u3047, p1_p3_u3046, p1_p3_u3045, p1_p3_u3044, p1_p3_u3043, p1_p3_u3042, p1_p3_u3041, p1_p3_u3040, p1_p3_u3039, p1_p3_u3038, p1_p3_u3037, p1_p3_u3036, p1_p3_u3035, p1_p3_u3034, p1_p3_u3033, p1_p3_u3032, p1_p3_u3031, p1_p3_u3030, p1_p3_u3029, p1_p3_u3280, p1_p3_u3281, p1_p3_u3028, p1_p3_u3027, p1_p3_u3026, p1_p3_u3025, p1_p3_u3024, p1_p3_u3023, p1_p3_u3022, p1_p3_u3021, p1_p3_u3020, p1_p3_u3019, p1_p3_u3018, p1_p3_u3017, p1_p3_u3016, p1_p3_u3015, p1_p3_u3014, p1_p3_u3013, p1_p3_u3012, p1_p3_u3011, p1_p3_u3010, p1_p3_u3009, p1_p3_u3008, p1_p3_u3007, p1_p3_u3006, p1_p3_u3005, p1_p3_u3004, p1_p3_u3003, p1_p3_u3002, p1_p3_u3001, p1_p3_u3000, p1_p3_u2999, p1_p3_u3282, p1_p3_u2998, p1_p3_u2997, p1_p3_u2996, p1_p3_u2995, p1_p3_u2994, p1_p3_u2993, p1_p3_u2992, p1_p3_u2991, p1_p3_u2990, p1_p3_u2989, p1_p3_u2988, p1_p3_u2987, p1_p3_u2986, p1_p3_u2985, p1_p3_u2984, p1_p3_u2983, p1_p3_u2982, p1_p3_u2981, p1_p3_u2980, p1_p3_u2979, p1_p3_u2978, p1_p3_u2977, p1_p3_u2976, p1_p3_u2975, p1_p3_u2974, p1_p3_u2973, p1_p3_u2972, p1_p3_u2971, p1_p3_u2970, p1_p3_u2969, p1_p3_u2968, p1_p3_u2967, p1_p3_u2966, p1_p3_u2965, p1_p3_u2964, p1_p3_u2963, p1_p3_u2962, p1_p3_u2961, p1_p3_u2960, p1_p3_u2959, p1_p3_u2958, p1_p3_u2957, p1_p3_u2956, p1_p3_u2955, p1_p3_u2954, p1_p3_u2953, p1_p3_u2952, p1_p3_u2951, p1_p3_u2950, p1_p3_u2949, p1_p3_u2948, p1_p3_u2947, p1_p3_u2946, p1_p3_u2945, p1_p3_u2944, p1_p3_u2943, p1_p3_u2942, p1_p3_u2941, p1_p3_u2940, p1_p3_u2939, p1_p3_u2938, p1_p3_u2937, p1_p3_u2936, p1_p3_u2935, p1_p3_u2934, p1_p3_u2933, p1_p3_u2932, p1_p3_u2931, p1_p3_u2930, p1_p3_u2929, p1_p3_u2928, p1_p3_u2927, p1_p3_u2926, p1_p3_u2925, p1_p3_u2924, p1_p3_u2923, p1_p3_u2922, p1_p3_u2921, p1_p3_u2920, p1_p3_u2919, p1_p3_u2918, p1_p3_u2917, p1_p3_u2916, p1_p3_u2915, p1_p3_u2914, p1_p3_u2913, p1_p3_u2912, p1_p3_u2911, p1_p3_u2910, p1_p3_u2909, p1_p3_u2908, p1_p3_u2907, p1_p3_u2906, p1_p3_u2905, p1_p3_u2904, p1_p3_u2903, p1_p3_u2902, p1_p3_u2901, p1_p3_u2900, p1_p3_u2899, p1_p3_u2898, p1_p3_u2897, p1_p3_u2896, p1_p3_u2895, p1_p3_u2894, p1_p3_u2893, p1_p3_u2892, p1_p3_u2891, p1_p3_u2890, p1_p3_u2889, p1_p3_u2888, p1_p3_u2887, p1_p3_u2886, p1_p3_u2885, p1_p3_u2884, p1_p3_u2883, p1_p3_u2882, p1_p3_u2881, p1_p3_u2880, p1_p3_u2879, p1_p3_u2878, p1_p3_u2877, p1_p3_u2876, p1_p3_u2875, p1_p3_u2874, p1_p3_u2873, p1_p3_u2872, p1_p3_u2871, p1_p3_u2870, p1_p3_u2869, p1_p3_u2868, p1_p3_u3284, p1_p3_u3285, p1_p3_u3288, p1_p3_u3289, p1_p3_u3290, p1_p3_u2867, p1_p3_u2866, p1_p3_u2865, p1_p3_u2864, p1_p3_u2863, p1_p3_u2862, p1_p3_u2861, p1_p3_u2860, p1_p3_u2859, p1_p3_u2858, p1_p3_u2857, p1_p3_u2856, p1_p3_u2855, p1_p3_u2854, p1_p3_u2853, p1_p3_u2852, p1_p3_u2851, p1_p3_u2850, p1_p3_u2849, p1_p3_u2848, p1_p3_u2847, p1_p3_u2846, p1_p3_u2845, p1_p3_u2844, p1_p3_u2843, p1_p3_u2842, p1_p3_u2841, p1_p3_u2840, p1_p3_u2839, p1_p3_u2838, p1_p3_u2837, p1_p3_u2836, p1_p3_u2835, p1_p3_u2834, p1_p3_u2833, p1_p3_u2832, p1_p3_u2831, p1_p3_u2830, p1_p3_u2829, p1_p3_u2828, p1_p3_u2827, p1_p3_u2826, p1_p3_u2825, p1_p3_u2824, p1_p3_u2823, p1_p3_u2822, p1_p3_u2821, p1_p3_u2820, p1_p3_u2819, p1_p3_u2818, p1_p3_u2817, p1_p3_u2816, p1_p3_u2815, p1_p3_u2814, p1_p3_u2813, p1_p3_u2812, p1_p3_u2811, p1_p3_u2810, p1_p3_u2809, p1_p3_u2808, p1_p3_u2807, p1_p3_u2806, p1_p3_u2805, p1_p3_u2804, p1_p3_u2803, p1_p3_u2802, p1_p3_u2801, p1_p3_u2800, p1_p3_u2799, p1_p3_u2798, p1_p3_u2797, p1_p3_u2796, p1_p3_u2795, p1_p3_u2794, p1_p3_u2793, p1_p3_u2792, p1_p3_u2791, p1_p3_u2790, p1_p3_u2789, p1_p3_u2788, p1_p3_u2787, p1_p3_u2786, p1_p3_u2785, p1_p3_u2784, p1_p3_u2783, p1_p3_u2782, p1_p3_u2781, p1_p3_u2780, p1_p3_u2779, p1_p3_u2778, p1_p3_u2777, p1_p3_u2776, p1_p3_u2775, p1_p3_u2774, p1_p3_u2773, p1_p3_u2772, p1_p3_u2771, p1_p3_u2770, p1_p3_u2769, p1_p3_u2768, p1_p3_u2767, p1_p3_u2766, p1_p3_u2765, p1_p3_u2764, p1_p3_u2763, p1_p3_u2762, p1_p3_u2761, p1_p3_u2760, p1_p3_u2759, p1_p3_u2758, p1_p3_u2757, p1_p3_u2756, p1_p3_u2755, p1_p3_u2754, p1_p3_u2753, p1_p3_u2752, p1_p3_u2751, p1_p3_u2750, p1_p3_u2749, p1_p3_u2748, p1_p3_u2747, p1_p3_u2746, p1_p3_u2745, p1_p3_u2744, p1_p3_u2743, p1_p3_u2742, p1_p3_u2741, p1_p3_u2740, p1_p3_u2739, p1_p3_u2738, p1_p3_u2737, p1_p3_u2736, p1_p3_u2735, p1_p3_u2734, p1_p3_u2733, p1_p3_u2732, p1_p3_u2731, p1_p3_u2730, p1_p3_u2729, p1_p3_u2728, p1_p3_u2727, p1_p3_u2726, p1_p3_u2725, p1_p3_u2724, p1_p3_u2723, p1_p3_u2722, p1_p3_u2721, p1_p3_u2720, p1_p3_u2719, p1_p3_u2718, p1_p3_u2717, p1_p3_u2716, p1_p3_u2715, p1_p3_u2714, p1_p3_u2713, p1_p3_u2712, p1_p3_u2711, p1_p3_u2710, p1_p3_u2709, p1_p3_u2708, p1_p3_u2707, p1_p3_u2706, p1_p3_u2705, p1_p3_u2704, p1_p3_u2703, p1_p3_u2702, p1_p3_u2701, p1_p3_u2700, p1_p3_u2699, p1_p3_u2698, p1_p3_u2697, p1_p3_u2696, p1_p3_u2695, p1_p3_u2694, p1_p3_u2693, p1_p3_u2692, p1_p3_u2691, p1_p3_u2690, p1_p3_u2689, p1_p3_u2688, p1_p3_u2687, p1_p3_u2686, p1_p3_u2685, p1_p3_u2684, p1_p3_u2683, p1_p3_u2682, p1_p3_u2681, p1_p3_u2680, p1_p3_u2679, p1_p3_u2678, p1_p3_u2677, p1_p3_u2676, p1_p3_u2675, p1_p3_u2674, p1_p3_u2673, p1_p3_u2672, p1_p3_u2671, p1_p3_u2670, p1_p3_u2669, p1_p3_u2668, p1_p3_u2667, p1_p3_u2666, p1_p3_u2665, p1_p3_u2664, p1_p3_u2663, p1_p3_u2662, p1_p3_u2661, p1_p3_u2660, p1_p3_u2659, p1_p3_u2658, p1_p3_u2657, p1_p3_u2656, p1_p3_u2655, p1_p3_u2654, p1_p3_u2653, p1_p3_u2652, p1_p3_u2651, p1_p3_u2650, p1_p3_u2649, p1_p3_u2648, p1_p3_u2647, p1_p3_u2646, p1_p3_u2645, p1_p3_u2644, p1_p3_u2643, p1_p3_u2642, p1_p3_u2641, p1_p3_u2640, p1_p3_u2639, p1_p3_u3292, p1_p3_u2638, p1_p3_u3293, p1_p3_u3294, p1_p3_u2637, p1_p3_u3295, p1_p3_u2636, p1_p3_u3296, p1_p3_u2635, p1_p3_u3297, p1_p3_u2634, p1_p3_u2633, p1_p3_u3298, p1_p3_u3299, p1_p2_u3274, p1_p2_u3275, p1_p2_u3276, p1_p2_u3277, p1_p2_u3061, p1_p2_u3060, p1_p2_u3059, p1_p2_u3058, p1_p2_u3057, p1_p2_u3056, p1_p2_u3055, p1_p2_u3054, p1_p2_u3053, p1_p2_u3052, p1_p2_u3051, p1_p2_u3050, p1_p2_u3049, p1_p2_u3048, p1_p2_u3047, p1_p2_u3046, p1_p2_u3045, p1_p2_u3044, p1_p2_u3043, p1_p2_u3042, p1_p2_u3041, p1_p2_u3040, p1_p2_u3039, p1_p2_u3038, p1_p2_u3037, p1_p2_u3036, p1_p2_u3035, p1_p2_u3034, p1_p2_u3033, p1_p2_u3032, p1_p2_u3031, p1_p2_u3030, p1_p2_u3029, p1_p2_u3280, p1_p2_u3281, p1_p2_u3028, p1_p2_u3027, p1_p2_u3026, p1_p2_u3025, p1_p2_u3024, p1_p2_u3023, p1_p2_u3022, p1_p2_u3021, p1_p2_u3020, p1_p2_u3019, p1_p2_u3018, p1_p2_u3017, p1_p2_u3016, p1_p2_u3015, p1_p2_u3014, p1_p2_u3013, p1_p2_u3012, p1_p2_u3011, p1_p2_u3010, p1_p2_u3009, p1_p2_u3008, p1_p2_u3007, p1_p2_u3006, p1_p2_u3005, p1_p2_u3004, p1_p2_u3003, p1_p2_u3002, p1_p2_u3001, p1_p2_u3000, p1_p2_u2999, p1_p2_u3282, p1_p2_u2998, p1_p2_u2997, p1_p2_u2996, p1_p2_u2995, p1_p2_u2994, p1_p2_u2993, p1_p2_u2992, p1_p2_u2991, p1_p2_u2990, p1_p2_u2989, p1_p2_u2988, p1_p2_u2987, p1_p2_u2986, p1_p2_u2985, p1_p2_u2984, p1_p2_u2983, p1_p2_u2982, p1_p2_u2981, p1_p2_u2980, p1_p2_u2979, p1_p2_u2978, p1_p2_u2977, p1_p2_u2976, p1_p2_u2975, p1_p2_u2974, p1_p2_u2973, p1_p2_u2972, p1_p2_u2971, p1_p2_u2970, p1_p2_u2969, p1_p2_u2968, p1_p2_u2967, p1_p2_u2966, p1_p2_u2965, p1_p2_u2964, p1_p2_u2963, p1_p2_u2962, p1_p2_u2961, p1_p2_u2960, p1_p2_u2959, p1_p2_u2958, p1_p2_u2957, p1_p2_u2956, p1_p2_u2955, p1_p2_u2954, p1_p2_u2953, p1_p2_u2952, p1_p2_u2951, p1_p2_u2950, p1_p2_u2949, p1_p2_u2948, p1_p2_u2947, p1_p2_u2946, p1_p2_u2945, p1_p2_u2944, p1_p2_u2943, p1_p2_u2942, p1_p2_u2941, p1_p2_u2940, p1_p2_u2939, p1_p2_u2938, p1_p2_u2937, p1_p2_u2936, p1_p2_u2935, p1_p2_u2934, p1_p2_u2933, p1_p2_u2932, p1_p2_u2931, p1_p2_u2930, p1_p2_u2929, p1_p2_u2928, p1_p2_u2927, p1_p2_u2926, p1_p2_u2925, p1_p2_u2924, p1_p2_u2923, p1_p2_u2922, p1_p2_u2921, p1_p2_u2920, p1_p2_u2919, p1_p2_u2918, p1_p2_u2917, p1_p2_u2916, p1_p2_u2915, p1_p2_u2914, p1_p2_u2913, p1_p2_u2912, p1_p2_u2911, p1_p2_u2910, p1_p2_u2909, p1_p2_u2908, p1_p2_u2907, p1_p2_u2906, p1_p2_u2905, p1_p2_u2904, p1_p2_u2903, p1_p2_u2902, p1_p2_u2901, p1_p2_u2900, p1_p2_u2899, p1_p2_u2898, p1_p2_u2897, p1_p2_u2896, p1_p2_u2895, p1_p2_u2894, p1_p2_u2893, p1_p2_u2892, p1_p2_u2891, p1_p2_u2890, p1_p2_u2889, p1_p2_u2888, p1_p2_u2887, p1_p2_u2886, p1_p2_u2885, p1_p2_u2884, p1_p2_u2883, p1_p2_u2882, p1_p2_u2881, p1_p2_u2880, p1_p2_u2879, p1_p2_u2878, p1_p2_u2877, p1_p2_u2876, p1_p2_u2875, p1_p2_u2874, p1_p2_u2873, p1_p2_u2872, p1_p2_u2871, p1_p2_u2870, p1_p2_u2869, p1_p2_u2868, p1_p2_u3284, p1_p2_u3285, p1_p2_u3288, p1_p2_u3289, p1_p2_u3290, p1_p2_u2867, p1_p2_u2866, p1_p2_u2865, p1_p2_u2864, p1_p2_u2863, p1_p2_u2862, p1_p2_u2861, p1_p2_u2860, p1_p2_u2859, p1_p2_u2858, p1_p2_u2857, p1_p2_u2856, p1_p2_u2855, p1_p2_u2854, p1_p2_u2853, p1_p2_u2852, p1_p2_u2851, p1_p2_u2850, p1_p2_u2849, p1_p2_u2848, p1_p2_u2847, p1_p2_u2846, p1_p2_u2845, p1_p2_u2844, p1_p2_u2843, p1_p2_u2842, p1_p2_u2841, p1_p2_u2840, p1_p2_u2839, p1_p2_u2838, p1_p2_u2837, p1_p2_u2836, p1_p2_u2835, p1_p2_u2834, p1_p2_u2833, p1_p2_u2832, p1_p2_u2831, p1_p2_u2830, p1_p2_u2829, p1_p2_u2828, p1_p2_u2827, p1_p2_u2826, p1_p2_u2825, p1_p2_u2824, p1_p2_u2823, p1_p2_u2822, p1_p2_u2821, p1_p2_u2820, p1_p2_u2819, p1_p2_u2818, p1_p2_u2817, p1_p2_u2816, p1_p2_u2815, p1_p2_u2814, p1_p2_u2813, p1_p2_u2812, p1_p2_u2811, p1_p2_u2810, p1_p2_u2809, p1_p2_u2808, p1_p2_u2807, p1_p2_u2806, p1_p2_u2805, p1_p2_u2804, p1_p2_u2803, p1_p2_u2802, p1_p2_u2801, p1_p2_u2800, p1_p2_u2799, p1_p2_u2798, p1_p2_u2797, p1_p2_u2796, p1_p2_u2795, p1_p2_u2794, p1_p2_u2793, p1_p2_u2792, p1_p2_u2791, p1_p2_u2790, p1_p2_u2789, p1_p2_u2788, p1_p2_u2787, p1_p2_u2786, p1_p2_u2785, p1_p2_u2784, p1_p2_u2783, p1_p2_u2782, p1_p2_u2781, p1_p2_u2780, p1_p2_u2779, p1_p2_u2778, p1_p2_u2777, p1_p2_u2776, p1_p2_u2775, p1_p2_u2774, p1_p2_u2773, p1_p2_u2772, p1_p2_u2771, p1_p2_u2770, p1_p2_u2769, p1_p2_u2768, p1_p2_u2767, p1_p2_u2766, p1_p2_u2765, p1_p2_u2764, p1_p2_u2763, p1_p2_u2762, p1_p2_u2761, p1_p2_u2760, p1_p2_u2759, p1_p2_u2758, p1_p2_u2757, p1_p2_u2756, p1_p2_u2755, p1_p2_u2754, p1_p2_u2753, p1_p2_u2752, p1_p2_u2751, p1_p2_u2750, p1_p2_u2749, p1_p2_u2748, p1_p2_u2747, p1_p2_u2746, p1_p2_u2745, p1_p2_u2744, p1_p2_u2743, p1_p2_u2742, p1_p2_u2741, p1_p2_u2740, p1_p2_u2739, p1_p2_u2738, p1_p2_u2737, p1_p2_u2736, p1_p2_u2735, p1_p2_u2734, p1_p2_u2733, p1_p2_u2732, p1_p2_u2731, p1_p2_u2730, p1_p2_u2729, p1_p2_u2728, p1_p2_u2727, p1_p2_u2726, p1_p2_u2725, p1_p2_u2724, p1_p2_u2723, p1_p2_u2722, p1_p2_u2721, p1_p2_u2720, p1_p2_u2719, p1_p2_u2718, p1_p2_u2717, p1_p2_u2716, p1_p2_u2715, p1_p2_u2714, p1_p2_u2713, p1_p2_u2712, p1_p2_u2711, p1_p2_u2710, p1_p2_u2709, p1_p2_u2708, p1_p2_u2707, p1_p2_u2706, p1_p2_u2705, p1_p2_u2704, p1_p2_u2703, p1_p2_u2702, p1_p2_u2701, p1_p2_u2700, p1_p2_u2699, p1_p2_u2698, p1_p2_u2697, p1_p2_u2696, p1_p2_u2695, p1_p2_u2694, p1_p2_u2693, p1_p2_u2692, p1_p2_u2691, p1_p2_u2690, p1_p2_u2689, p1_p2_u2688, p1_p2_u2687, p1_p2_u2686, p1_p2_u2685, p1_p2_u2684, p1_p2_u2683, p1_p2_u2682, p1_p2_u2681, p1_p2_u2680, p1_p2_u2679, p1_p2_u2678, p1_p2_u2677, p1_p2_u2676, p1_p2_u2675, p1_p2_u2674, p1_p2_u2673, p1_p2_u2672, p1_p2_u2671, p1_p2_u2670, p1_p2_u2669, p1_p2_u2668, p1_p2_u2667, p1_p2_u2666, p1_p2_u2665, p1_p2_u2664, p1_p2_u2663, p1_p2_u2662, p1_p2_u2661, p1_p2_u2660, p1_p2_u2659, p1_p2_u2658, p1_p2_u2657, p1_p2_u2656, p1_p2_u2655, p1_p2_u2654, p1_p2_u2653, p1_p2_u2652, p1_p2_u2651, p1_p2_u2650, p1_p2_u2649, p1_p2_u2648, p1_p2_u2647, p1_p2_u2646, p1_p2_u2645, p1_p2_u2644, p1_p2_u2643, p1_p2_u2642, p1_p2_u2641, p1_p2_u2640, p1_p2_u2639, p1_p2_u3292, p1_p2_u2638, p1_p2_u3293, p1_p2_u3294, p1_p2_u2637, p1_p2_u3295, p1_p2_u2636, p1_p2_u3296, p1_p2_u2635, p1_p2_u3297, p1_p2_u2634, p1_p2_u2633, p1_p2_u3298, p1_p2_u3299, p1_p1_u3288, p1_p1_u3289, p1_p1_u3290, p1_p1_u3291, p1_p1_u3077, p1_p1_u3076, p1_p1_u3075, p1_p1_u3074, p1_p1_u3073, p1_p1_u3072, p1_p1_u3071, p1_p1_u3070, p1_p1_u3069, p1_p1_u3068, p1_p1_u3067, p1_p1_u3066, p1_p1_u3065, p1_p1_u3064, p1_p1_u3063, p1_p1_u3062, p1_p1_u3061, p1_p1_u3060, p1_p1_u3059, p1_p1_u3058, p1_p1_u3057, p1_p1_u3056, p1_p1_u3055, p1_p1_u3054, p1_p1_u3053, p1_p1_u3052, p1_p1_u3051, p1_p1_u3050, p1_p1_u3049, p1_p1_u3048, p1_p1_u3047, p1_p1_u3046, p1_p1_u3045, p1_p1_u3294, p1_p1_u3295, p1_p1_u3044, p1_p1_u3043, p1_p1_u3042, p1_p1_u3041, p1_p1_u3040, p1_p1_u3039, p1_p1_u3038, p1_p1_u3037, p1_p1_u3036, p1_p1_u3035, p1_p1_u3034, p1_p1_u3033, p1_p1_u3032, p1_p1_u3031, p1_p1_u3030, p1_p1_u3029, p1_p1_u3028, p1_p1_u3027, p1_p1_u3026, p1_p1_u3025, p1_p1_u3024, p1_p1_u3023, p1_p1_u3022, p1_p1_u3021, p1_p1_u3020, p1_p1_u3019, p1_p1_u3018, p1_p1_u3017, p1_p1_u3016, p1_p1_u3015, p1_p1_u3296, p1_p1_u3014, p1_p1_u3013, p1_p1_u3012, p1_p1_u3011, p1_p1_u3010, p1_p1_u3009, p1_p1_u3008, p1_p1_u3007, p1_p1_u3006, p1_p1_u3005, p1_p1_u3004, p1_p1_u3003, p1_p1_u3002, p1_p1_u3001, p1_p1_u3000, p1_p1_u2999, p1_p1_u2998, p1_p1_u2997, p1_p1_u2996, p1_p1_u2995, p1_p1_u2994, p1_p1_u2993, p1_p1_u2992, p1_p1_u2991, p1_p1_u2990, p1_p1_u2989, p1_p1_u2988, p1_p1_u2987, p1_p1_u2986, p1_p1_u2985, p1_p1_u2984, p1_p1_u2983, p1_p1_u2982, p1_p1_u2981, p1_p1_u2980, p1_p1_u2979, p1_p1_u2978, p1_p1_u2977, p1_p1_u2976, p1_p1_u2975, p1_p1_u2974, p1_p1_u2973, p1_p1_u2972, p1_p1_u2971, p1_p1_u2970, p1_p1_u2969, p1_p1_u2968, p1_p1_u2967, p1_p1_u2966, p1_p1_u2965, p1_p1_u2964, p1_p1_u2963, p1_p1_u2962, p1_p1_u2961, p1_p1_u2960, p1_p1_u2959, p1_p1_u2958, p1_p1_u2957, p1_p1_u2956, p1_p1_u2955, p1_p1_u2954, p1_p1_u2953, p1_p1_u2952, p1_p1_u2951, p1_p1_u2950, p1_p1_u2949, p1_p1_u2948, p1_p1_u2947, p1_p1_u2946, p1_p1_u2945, p1_p1_u2944, p1_p1_u2943, p1_p1_u2942, p1_p1_u2941, p1_p1_u2940, p1_p1_u2939, p1_p1_u2938, p1_p1_u2937, p1_p1_u2936, p1_p1_u2935, p1_p1_u2934, p1_p1_u2933, p1_p1_u2932, p1_p1_u2931, p1_p1_u2930, p1_p1_u2929, p1_p1_u2928, p1_p1_u2927, p1_p1_u2926, p1_p1_u2925, p1_p1_u2924, p1_p1_u2923, p1_p1_u2922, p1_p1_u2921, p1_p1_u2920, p1_p1_u2919, p1_p1_u2918, p1_p1_u2917, p1_p1_u2916, p1_p1_u2915, p1_p1_u2914, p1_p1_u2913, p1_p1_u2912, p1_p1_u2911, p1_p1_u2910, p1_p1_u2909, p1_p1_u2908, p1_p1_u2907, p1_p1_u2906, p1_p1_u2905, p1_p1_u2904, p1_p1_u2903, p1_p1_u2902, p1_p1_u2901, p1_p1_u2900, p1_p1_u2899, p1_p1_u2898, p1_p1_u2897, p1_p1_u2896, p1_p1_u2895, p1_p1_u2894, p1_p1_u2893, p1_p1_u2892, p1_p1_u2891, p1_p1_u2890, p1_p1_u2889, p1_p1_u2888, p1_p1_u2887, p1_p1_u2886, p1_p1_u2885, p1_p1_u2884, p1_p1_u3298, p1_p1_u3299, p1_p1_u3302, p1_p1_u3303, p1_p1_u3304, p1_p1_u2883, p1_p1_u2882, p1_p1_u2881, p1_p1_u2880, p1_p1_u2879, p1_p1_u2878, p1_p1_u2877, p1_p1_u2876, p1_p1_u2875, p1_p1_u2874, p1_p1_u2873, p1_p1_u2872, p1_p1_u2871, p1_p1_u2870, p1_p1_u2869, p1_p1_u2868, p1_p1_u2867, p1_p1_u2866, p1_p1_u2865, p1_p1_u2864, p1_p1_u2863, p1_p1_u2862, p1_p1_u2861, p1_p1_u2860, p1_p1_u2859, p1_p1_u2858, p1_p1_u2857, p1_p1_u2856, p1_p1_u2855, p1_p1_u2854, p1_p1_u2853, p1_p1_u2852, p1_p1_u2851, p1_p1_u2850, p1_p1_u2849, p1_p1_u2848, p1_p1_u2847, p1_p1_u2846, p1_p1_u2845, p1_p1_u2844, p1_p1_u2843, p1_p1_u2842, p1_p1_u2841, p1_p1_u2840, p1_p1_u2839, p1_p1_u2838, p1_p1_u2837, p1_p1_u2836, p1_p1_u2835, p1_p1_u2834, p1_p1_u2833, p1_p1_u2832, p1_p1_u2831, p1_p1_u2830, p1_p1_u2829, p1_p1_u2828, p1_p1_u2827, p1_p1_u2826, p1_p1_u2825, p1_p1_u2824, p1_p1_u2823, p1_p1_u2822, p1_p1_u2821, p1_p1_u2820, p1_p1_u2819, p1_p1_u2818, p1_p1_u2817, p1_p1_u2816, p1_p1_u2815, p1_p1_u2814, p1_p1_u2813, p1_p1_u2812, p1_p1_u2811, p1_p1_u2810, p1_p1_u2809, p1_p1_u2808, p1_p1_u2807, p1_p1_u2806, p1_p1_u2805, p1_p1_u2804, p1_p1_u2803, p1_p1_u2802, p1_p1_u2801, p1_p1_u2800, p1_p1_u2799, p1_p1_u2798, p1_p1_u2797, p1_p1_u2796, p1_p1_u2795, p1_p1_u2794, p1_p1_u2793, p1_p1_u2792, p1_p1_u2791, p1_p1_u2790, p1_p1_u2789, p1_p1_u2788, p1_p1_u2787, p1_p1_u2786, p1_p1_u2785, p1_p1_u2784, p1_p1_u2783, p1_p1_u2782, p1_p1_u2781, p1_p1_u2780, p1_p1_u2779, p1_p1_u2778, p1_p1_u2777, p1_p1_u2776, p1_p1_u2775, p1_p1_u2774, p1_p1_u2773, p1_p1_u2772, p1_p1_u2771, p1_p1_u2770, p1_p1_u2769, p1_p1_u2768, p1_p1_u2767, p1_p1_u2766, p1_p1_u2765, p1_p1_u2764, p1_p1_u2763, p1_p1_u2762, p1_p1_u2761, p1_p1_u2760, p1_p1_u2759, p1_p1_u2758, p1_p1_u2757, p1_p1_u2756, p1_p1_u2755, p1_p1_u2754, p1_p1_u2753, p1_p1_u2752, p1_p1_u2751, p1_p1_u2750, p1_p1_u2749, p1_p1_u2748, p1_p1_u2747, p1_p1_u2746, p1_p1_u2745, p1_p1_u2744, p1_p1_u2743, p1_p1_u2742, p1_p1_u2741, p1_p1_u2740, p1_p1_u2739, p1_p1_u2738, p1_p1_u2737, p1_p1_u2736, p1_p1_u2735, p1_p1_u2734, p1_p1_u2733, p1_p1_u2732, p1_p1_u2731, p1_p1_u2730, p1_p1_u2729, p1_p1_u2728, p1_p1_u2727, p1_p1_u2726, p1_p1_u2725, p1_p1_u2724, p1_p1_u2723, p1_p1_u2722, p1_p1_u2721, p1_p1_u2720, p1_p1_u2719, p1_p1_u2718, p1_p1_u2717, p1_p1_u2716, p1_p1_u2715, p1_p1_u2714, p1_p1_u2713, p1_p1_u2712, p1_p1_u2711, p1_p1_u2710, p1_p1_u2709, p1_p1_u2708, p1_p1_u2707, p1_p1_u2706, p1_p1_u2705, p1_p1_u2704, p1_p1_u2703, p1_p1_u2702, p1_p1_u2701, p1_p1_u2700, p1_p1_u2699, p1_p1_u2698, p1_p1_u2697, p1_p1_u2696, p1_p1_u2695, p1_p1_u2694, p1_p1_u2693, p1_p1_u2692, p1_p1_u2691, p1_p1_u2690, p1_p1_u2689, p1_p1_u2688, p1_p1_u2687, p1_p1_u2686, p1_p1_u2685, p1_p1_u2684, p1_p1_u2683, p1_p1_u2682, p1_p1_u2681, p1_p1_u2680, p1_p1_u2679, p1_p1_u2678, p1_p1_u2677, p1_p1_u2676, p1_p1_u2675, p1_p1_u2674, p1_p1_u2673, p1_p1_u2672, p1_p1_u2671, p1_p1_u2670, p1_p1_u2669, p1_p1_u2668, p1_p1_u2667, p1_p1_u2666, p1_p1_u2665, p1_p1_u2664, p1_p1_u2663, p1_p1_u2662, p1_p1_u2661, p1_p1_u2660, p1_p1_u2659, p1_p1_u2658, p1_p1_u2657, p1_p1_u2656, p1_p1_u2655, p1_p1_u3306, p1_p1_u2654, p1_p1_u3307, p1_p1_u3308, p1_p1_u2653, p1_p1_u3309, p1_p1_u2652, p1_p1_u3310, p1_p1_u2651, p1_p1_u3311, p1_p1_u2650, p1_p1_u2649, p1_p1_u3312, p1_p1_u3313, p2_p3_u3274, p2_p3_u3275, p2_p3_u3276, p2_p3_u3277, p2_p3_u3061, p2_p3_u3060, p2_p3_u3059, p2_p3_u3058, p2_p3_u3057, p2_p3_u3056, p2_p3_u3055, p2_p3_u3054, p2_p3_u3053, p2_p3_u3052, p2_p3_u3051, p2_p3_u3050, p2_p3_u3049, p2_p3_u3048, p2_p3_u3047, p2_p3_u3046, p2_p3_u3045, p2_p3_u3044, p2_p3_u3043, p2_p3_u3042, p2_p3_u3041, p2_p3_u3040, p2_p3_u3039, p2_p3_u3038, p2_p3_u3037, p2_p3_u3036, p2_p3_u3035, p2_p3_u3034, p2_p3_u3033, p2_p3_u3032, p2_p3_u3031, p2_p3_u3030, p2_p3_u3029, p2_p3_u3280, p2_p3_u3281, p2_p3_u3028, p2_p3_u3027, p2_p3_u3026, p2_p3_u3025, p2_p3_u3024, p2_p3_u3023, p2_p3_u3022, p2_p3_u3021, p2_p3_u3020, p2_p3_u3019, p2_p3_u3018, p2_p3_u3017, p2_p3_u3016, p2_p3_u3015, p2_p3_u3014, p2_p3_u3013, p2_p3_u3012, p2_p3_u3011, p2_p3_u3010, p2_p3_u3009, p2_p3_u3008, p2_p3_u3007, p2_p3_u3006, p2_p3_u3005, p2_p3_u3004, p2_p3_u3003, p2_p3_u3002, p2_p3_u3001, p2_p3_u3000, p2_p3_u2999, p2_p3_u3282, p2_p3_u2998, p2_p3_u2997, p2_p3_u2996, p2_p3_u2995, p2_p3_u2994, p2_p3_u2993, p2_p3_u2992, p2_p3_u2991, p2_p3_u2990, p2_p3_u2989, p2_p3_u2988, p2_p3_u2987, p2_p3_u2986, p2_p3_u2985, p2_p3_u2984, p2_p3_u2983, p2_p3_u2982, p2_p3_u2981, p2_p3_u2980, p2_p3_u2979, p2_p3_u2978, p2_p3_u2977, p2_p3_u2976, p2_p3_u2975, p2_p3_u2974, p2_p3_u2973, p2_p3_u2972, p2_p3_u2971, p2_p3_u2970, p2_p3_u2969, p2_p3_u2968, p2_p3_u2967, p2_p3_u2966, p2_p3_u2965, p2_p3_u2964, p2_p3_u2963, p2_p3_u2962, p2_p3_u2961, p2_p3_u2960, p2_p3_u2959, p2_p3_u2958, p2_p3_u2957, p2_p3_u2956, p2_p3_u2955, p2_p3_u2954, p2_p3_u2953, p2_p3_u2952, p2_p3_u2951, p2_p3_u2950, p2_p3_u2949, p2_p3_u2948, p2_p3_u2947, p2_p3_u2946, p2_p3_u2945, p2_p3_u2944, p2_p3_u2943, p2_p3_u2942, p2_p3_u2941, p2_p3_u2940, p2_p3_u2939, p2_p3_u2938, p2_p3_u2937, p2_p3_u2936, p2_p3_u2935, p2_p3_u2934, p2_p3_u2933, p2_p3_u2932, p2_p3_u2931, p2_p3_u2930, p2_p3_u2929, p2_p3_u2928, p2_p3_u2927, p2_p3_u2926, p2_p3_u2925, p2_p3_u2924, p2_p3_u2923, p2_p3_u2922, p2_p3_u2921, p2_p3_u2920, p2_p3_u2919, p2_p3_u2918, p2_p3_u2917, p2_p3_u2916, p2_p3_u2915, p2_p3_u2914, p2_p3_u2913, p2_p3_u2912, p2_p3_u2911, p2_p3_u2910, p2_p3_u2909, p2_p3_u2908, p2_p3_u2907, p2_p3_u2906, p2_p3_u2905, p2_p3_u2904, p2_p3_u2903, p2_p3_u2902, p2_p3_u2901, p2_p3_u2900, p2_p3_u2899, p2_p3_u2898, p2_p3_u2897, p2_p3_u2896, p2_p3_u2895, p2_p3_u2894, p2_p3_u2893, p2_p3_u2892, p2_p3_u2891, p2_p3_u2890, p2_p3_u2889, p2_p3_u2888, p2_p3_u2887, p2_p3_u2886, p2_p3_u2885, p2_p3_u2884, p2_p3_u2883, p2_p3_u2882, p2_p3_u2881, p2_p3_u2880, p2_p3_u2879, p2_p3_u2878, p2_p3_u2877, p2_p3_u2876, p2_p3_u2875, p2_p3_u2874, p2_p3_u2873, p2_p3_u2872, p2_p3_u2871, p2_p3_u2870, p2_p3_u2869, p2_p3_u2868, p2_p3_u3284, p2_p3_u3285, p2_p3_u3288, p2_p3_u3289, p2_p3_u3290, p2_p3_u2867, p2_p3_u2866, p2_p3_u2865, p2_p3_u2864, p2_p3_u2863, p2_p3_u2862, p2_p3_u2861, p2_p3_u2860, p2_p3_u2859, p2_p3_u2858, p2_p3_u2857, p2_p3_u2856, p2_p3_u2855, p2_p3_u2854, p2_p3_u2853, p2_p3_u2852, p2_p3_u2851, p2_p3_u2850, p2_p3_u2849, p2_p3_u2848, p2_p3_u2847, p2_p3_u2846, p2_p3_u2845, p2_p3_u2844, p2_p3_u2843, p2_p3_u2842, p2_p3_u2841, p2_p3_u2840, p2_p3_u2839, p2_p3_u2838, p2_p3_u2837, p2_p3_u2836, p2_p3_u2835, p2_p3_u2834, p2_p3_u2833, p2_p3_u2832, p2_p3_u2831, p2_p3_u2830, p2_p3_u2829, p2_p3_u2828, p2_p3_u2827, p2_p3_u2826, p2_p3_u2825, p2_p3_u2824, p2_p3_u2823, p2_p3_u2822, p2_p3_u2821, p2_p3_u2820, p2_p3_u2819, p2_p3_u2818, p2_p3_u2817, p2_p3_u2816, p2_p3_u2815, p2_p3_u2814, p2_p3_u2813, p2_p3_u2812, p2_p3_u2811, p2_p3_u2810, p2_p3_u2809, p2_p3_u2808, p2_p3_u2807, p2_p3_u2806, p2_p3_u2805, p2_p3_u2804, p2_p3_u2803, p2_p3_u2802, p2_p3_u2801, p2_p3_u2800, p2_p3_u2799, p2_p3_u2798, p2_p3_u2797, p2_p3_u2796, p2_p3_u2795, p2_p3_u2794, p2_p3_u2793, p2_p3_u2792, p2_p3_u2791, p2_p3_u2790, p2_p3_u2789, p2_p3_u2788, p2_p3_u2787, p2_p3_u2786, p2_p3_u2785, p2_p3_u2784, p2_p3_u2783, p2_p3_u2782, p2_p3_u2781, p2_p3_u2780, p2_p3_u2779, p2_p3_u2778, p2_p3_u2777, p2_p3_u2776, p2_p3_u2775, p2_p3_u2774, p2_p3_u2773, p2_p3_u2772, p2_p3_u2771, p2_p3_u2770, p2_p3_u2769, p2_p3_u2768, p2_p3_u2767, p2_p3_u2766, p2_p3_u2765, p2_p3_u2764, p2_p3_u2763, p2_p3_u2762, p2_p3_u2761, p2_p3_u2760, p2_p3_u2759, p2_p3_u2758, p2_p3_u2757, p2_p3_u2756, p2_p3_u2755, p2_p3_u2754, p2_p3_u2753, p2_p3_u2752, p2_p3_u2751, p2_p3_u2750, p2_p3_u2749, p2_p3_u2748, p2_p3_u2747, p2_p3_u2746, p2_p3_u2745, p2_p3_u2744, p2_p3_u2743, p2_p3_u2742, p2_p3_u2741, p2_p3_u2740, p2_p3_u2739, p2_p3_u2738, p2_p3_u2737, p2_p3_u2736, p2_p3_u2735, p2_p3_u2734, p2_p3_u2733, p2_p3_u2732, p2_p3_u2731, p2_p3_u2730, p2_p3_u2729, p2_p3_u2728, p2_p3_u2727, p2_p3_u2726, p2_p3_u2725, p2_p3_u2724, p2_p3_u2723, p2_p3_u2722, p2_p3_u2721, p2_p3_u2720, p2_p3_u2719, p2_p3_u2718, p2_p3_u2717, p2_p3_u2716, p2_p3_u2715, p2_p3_u2714, p2_p3_u2713, p2_p3_u2712, p2_p3_u2711, p2_p3_u2710, p2_p3_u2709, p2_p3_u2708, p2_p3_u2707, p2_p3_u2706, p2_p3_u2705, p2_p3_u2704, p2_p3_u2703, p2_p3_u2702, p2_p3_u2701, p2_p3_u2700, p2_p3_u2699, p2_p3_u2698, p2_p3_u2697, p2_p3_u2696, p2_p3_u2695, p2_p3_u2694, p2_p3_u2693, p2_p3_u2692, p2_p3_u2691, p2_p3_u2690, p2_p3_u2689, p2_p3_u2688, p2_p3_u2687, p2_p3_u2686, p2_p3_u2685, p2_p3_u2684, p2_p3_u2683, p2_p3_u2682, p2_p3_u2681, p2_p3_u2680, p2_p3_u2679, p2_p3_u2678, p2_p3_u2677, p2_p3_u2676, p2_p3_u2675, p2_p3_u2674, p2_p3_u2673, p2_p3_u2672, p2_p3_u2671, p2_p3_u2670, p2_p3_u2669, p2_p3_u2668, p2_p3_u2667, p2_p3_u2666, p2_p3_u2665, p2_p3_u2664, p2_p3_u2663, p2_p3_u2662, p2_p3_u2661, p2_p3_u2660, p2_p3_u2659, p2_p3_u2658, p2_p3_u2657, p2_p3_u2656, p2_p3_u2655, p2_p3_u2654, p2_p3_u2653, p2_p3_u2652, p2_p3_u2651, p2_p3_u2650, p2_p3_u2649, p2_p3_u2648, p2_p3_u2647, p2_p3_u2646, p2_p3_u2645, p2_p3_u2644, p2_p3_u2643, p2_p3_u2642, p2_p3_u2641, p2_p3_u2640, p2_p3_u2639, p2_p3_u3292, p2_p3_u2638, p2_p3_u3293, p2_p3_u3294, p2_p3_u2637, p2_p3_u3295, p2_p3_u2636, p2_p3_u3296, p2_p3_u2635, p2_p3_u3297, p2_p3_u2634, p2_p3_u2633, p2_p3_u3298, p2_p3_u3299, p2_p2_u3274, p2_p2_u3275, p2_p2_u3276, p2_p2_u3277, p2_p2_u3061, p2_p2_u3060, p2_p2_u3059, p2_p2_u3058, p2_p2_u3057, p2_p2_u3056, p2_p2_u3055, p2_p2_u3054, p2_p2_u3053, p2_p2_u3052, p2_p2_u3051, p2_p2_u3050, p2_p2_u3049, p2_p2_u3048, p2_p2_u3047, p2_p2_u3046, p2_p2_u3045, p2_p2_u3044, p2_p2_u3043, p2_p2_u3042, p2_p2_u3041, p2_p2_u3040, p2_p2_u3039, p2_p2_u3038, p2_p2_u3037, p2_p2_u3036, p2_p2_u3035, p2_p2_u3034, p2_p2_u3033, p2_p2_u3032, p2_p2_u3031, p2_p2_u3030, p2_p2_u3029, p2_p2_u3280, p2_p2_u3281, p2_p2_u3028, p2_p2_u3027, p2_p2_u3026, p2_p2_u3025, p2_p2_u3024, p2_p2_u3023, p2_p2_u3022, p2_p2_u3021, p2_p2_u3020, p2_p2_u3019, p2_p2_u3018, p2_p2_u3017, p2_p2_u3016, p2_p2_u3015, p2_p2_u3014, p2_p2_u3013, p2_p2_u3012, p2_p2_u3011, p2_p2_u3010, p2_p2_u3009, p2_p2_u3008, p2_p2_u3007, p2_p2_u3006, p2_p2_u3005, p2_p2_u3004, p2_p2_u3003, p2_p2_u3002, p2_p2_u3001, p2_p2_u3000, p2_p2_u2999, p2_p2_u3282, p2_p2_u2998, p2_p2_u2997, p2_p2_u2996, p2_p2_u2995, p2_p2_u2994, p2_p2_u2993, p2_p2_u2992, p2_p2_u2991, p2_p2_u2990, p2_p2_u2989, p2_p2_u2988, p2_p2_u2987, p2_p2_u2986, p2_p2_u2985, p2_p2_u2984, p2_p2_u2983, p2_p2_u2982, p2_p2_u2981, p2_p2_u2980, p2_p2_u2979, p2_p2_u2978, p2_p2_u2977, p2_p2_u2976, p2_p2_u2975, p2_p2_u2974, p2_p2_u2973, p2_p2_u2972, p2_p2_u2971, p2_p2_u2970, p2_p2_u2969, p2_p2_u2968, p2_p2_u2967, p2_p2_u2966, p2_p2_u2965, p2_p2_u2964, p2_p2_u2963, p2_p2_u2962, p2_p2_u2961, p2_p2_u2960, p2_p2_u2959, p2_p2_u2958, p2_p2_u2957, p2_p2_u2956, p2_p2_u2955, p2_p2_u2954, p2_p2_u2953, p2_p2_u2952, p2_p2_u2951, p2_p2_u2950, p2_p2_u2949, p2_p2_u2948, p2_p2_u2947, p2_p2_u2946, p2_p2_u2945, p2_p2_u2944, p2_p2_u2943, p2_p2_u2942, p2_p2_u2941, p2_p2_u2940, p2_p2_u2939, p2_p2_u2938, p2_p2_u2937, p2_p2_u2936, p2_p2_u2935, p2_p2_u2934, p2_p2_u2933, p2_p2_u2932, p2_p2_u2931, p2_p2_u2930, p2_p2_u2929, p2_p2_u2928, p2_p2_u2927, p2_p2_u2926, p2_p2_u2925, p2_p2_u2924, p2_p2_u2923, p2_p2_u2922, p2_p2_u2921, p2_p2_u2920, p2_p2_u2919, p2_p2_u2918, p2_p2_u2917, p2_p2_u2916, p2_p2_u2915, p2_p2_u2914, p2_p2_u2913, p2_p2_u2912, p2_p2_u2911, p2_p2_u2910, p2_p2_u2909, p2_p2_u2908, p2_p2_u2907, p2_p2_u2906, p2_p2_u2905, p2_p2_u2904, p2_p2_u2903, p2_p2_u2902, p2_p2_u2901, p2_p2_u2900, p2_p2_u2899, p2_p2_u2898, p2_p2_u2897, p2_p2_u2896, p2_p2_u2895, p2_p2_u2894, p2_p2_u2893, p2_p2_u2892, p2_p2_u2891, p2_p2_u2890, p2_p2_u2889, p2_p2_u2888, p2_p2_u2887, p2_p2_u2886, p2_p2_u2885, p2_p2_u2884, p2_p2_u2883, p2_p2_u2882, p2_p2_u2881, p2_p2_u2880, p2_p2_u2879, p2_p2_u2878, p2_p2_u2877, p2_p2_u2876, p2_p2_u2875, p2_p2_u2874, p2_p2_u2873, p2_p2_u2872, p2_p2_u2871, p2_p2_u2870, p2_p2_u2869, p2_p2_u2868, p2_p2_u3284, p2_p2_u3285, p2_p2_u3288, p2_p2_u3289, p2_p2_u3290, p2_p2_u2867, p2_p2_u2866, p2_p2_u2865, p2_p2_u2864, p2_p2_u2863, p2_p2_u2862, p2_p2_u2861, p2_p2_u2860, p2_p2_u2859, p2_p2_u2858, p2_p2_u2857, p2_p2_u2856, p2_p2_u2855, p2_p2_u2854, p2_p2_u2853, p2_p2_u2852, p2_p2_u2851, p2_p2_u2850, p2_p2_u2849, p2_p2_u2848, p2_p2_u2847, p2_p2_u2846, p2_p2_u2845, p2_p2_u2844, p2_p2_u2843, p2_p2_u2842, p2_p2_u2841, p2_p2_u2840, p2_p2_u2839, p2_p2_u2838, p2_p2_u2837, p2_p2_u2836, p2_p2_u2835, p2_p2_u2834, p2_p2_u2833, p2_p2_u2832, p2_p2_u2831, p2_p2_u2830, p2_p2_u2829, p2_p2_u2828, p2_p2_u2827, p2_p2_u2826, p2_p2_u2825, p2_p2_u2824, p2_p2_u2823, p2_p2_u2822, p2_p2_u2821, p2_p2_u2820, p2_p2_u2819, p2_p2_u2818, p2_p2_u2817, p2_p2_u2816, p2_p2_u2815, p2_p2_u2814, p2_p2_u2813, p2_p2_u2812, p2_p2_u2811, p2_p2_u2810, p2_p2_u2809, p2_p2_u2808, p2_p2_u2807, p2_p2_u2806, p2_p2_u2805, p2_p2_u2804, p2_p2_u2803, p2_p2_u2802, p2_p2_u2801, p2_p2_u2800, p2_p2_u2799, p2_p2_u2798, p2_p2_u2797, p2_p2_u2796, p2_p2_u2795, p2_p2_u2794, p2_p2_u2793, p2_p2_u2792, p2_p2_u2791, p2_p2_u2790, p2_p2_u2789, p2_p2_u2788, p2_p2_u2787, p2_p2_u2786, p2_p2_u2785, p2_p2_u2784, p2_p2_u2783, p2_p2_u2782, p2_p2_u2781, p2_p2_u2780, p2_p2_u2779, p2_p2_u2778, p2_p2_u2777, p2_p2_u2776, p2_p2_u2775, p2_p2_u2774, p2_p2_u2773, p2_p2_u2772, p2_p2_u2771, p2_p2_u2770, p2_p2_u2769, p2_p2_u2768, p2_p2_u2767, p2_p2_u2766, p2_p2_u2765, p2_p2_u2764, p2_p2_u2763, p2_p2_u2762, p2_p2_u2761, p2_p2_u2760, p2_p2_u2759, p2_p2_u2758, p2_p2_u2757, p2_p2_u2756, p2_p2_u2755, p2_p2_u2754, p2_p2_u2753, p2_p2_u2752, p2_p2_u2751, p2_p2_u2750, p2_p2_u2749, p2_p2_u2748, p2_p2_u2747, p2_p2_u2746, p2_p2_u2745, p2_p2_u2744, p2_p2_u2743, p2_p2_u2742, p2_p2_u2741, p2_p2_u2740, p2_p2_u2739, p2_p2_u2738, p2_p2_u2737, p2_p2_u2736, p2_p2_u2735, p2_p2_u2734, p2_p2_u2733, p2_p2_u2732, p2_p2_u2731, p2_p2_u2730, p2_p2_u2729, p2_p2_u2728, p2_p2_u2727, p2_p2_u2726, p2_p2_u2725, p2_p2_u2724, p2_p2_u2723, p2_p2_u2722, p2_p2_u2721, p2_p2_u2720, p2_p2_u2719, p2_p2_u2718, p2_p2_u2717, p2_p2_u2716, p2_p2_u2715, p2_p2_u2714, p2_p2_u2713, p2_p2_u2712, p2_p2_u2711, p2_p2_u2710, p2_p2_u2709, p2_p2_u2708, p2_p2_u2707, p2_p2_u2706, p2_p2_u2705, p2_p2_u2704, p2_p2_u2703, p2_p2_u2702, p2_p2_u2701, p2_p2_u2700, p2_p2_u2699, p2_p2_u2698, p2_p2_u2697, p2_p2_u2696, p2_p2_u2695, p2_p2_u2694, p2_p2_u2693, p2_p2_u2692, p2_p2_u2691, p2_p2_u2690, p2_p2_u2689, p2_p2_u2688, p2_p2_u2687, p2_p2_u2686, p2_p2_u2685, p2_p2_u2684, p2_p2_u2683, p2_p2_u2682, p2_p2_u2681, p2_p2_u2680, p2_p2_u2679, p2_p2_u2678, p2_p2_u2677, p2_p2_u2676, p2_p2_u2675, p2_p2_u2674, p2_p2_u2673, p2_p2_u2672, p2_p2_u2671, p2_p2_u2670, p2_p2_u2669, p2_p2_u2668, p2_p2_u2667, p2_p2_u2666, p2_p2_u2665, p2_p2_u2664, p2_p2_u2663, p2_p2_u2662, p2_p2_u2661, p2_p2_u2660, p2_p2_u2659, p2_p2_u2658, p2_p2_u2657, p2_p2_u2656, p2_p2_u2655, p2_p2_u2654, p2_p2_u2653, p2_p2_u2652, p2_p2_u2651, p2_p2_u2650, p2_p2_u2649, p2_p2_u2648, p2_p2_u2647, p2_p2_u2646, p2_p2_u2645, p2_p2_u2644, p2_p2_u2643, p2_p2_u2642, p2_p2_u2641, p2_p2_u2640, p2_p2_u2639, p2_p2_u3292, p2_p2_u2638, p2_p2_u3293, p2_p2_u3294, p2_p2_u2637, p2_p2_u3295, p2_p2_u2636, p2_p2_u3296, p2_p2_u2635, p2_p2_u3297, p2_p2_u2634, p2_p2_u2633, p2_p2_u3298, p2_p2_u3299, p2_p1_u3288, p2_p1_u3289, p2_p1_u3290, p2_p1_u3291, p2_p1_u3077, p2_p1_u3076, p2_p1_u3075, p2_p1_u3074, p2_p1_u3073, p2_p1_u3072, p2_p1_u3071, p2_p1_u3070, p2_p1_u3069, p2_p1_u3068, p2_p1_u3067, p2_p1_u3066, p2_p1_u3065, p2_p1_u3064, p2_p1_u3063, p2_p1_u3062, p2_p1_u3061, p2_p1_u3060, p2_p1_u3059, p2_p1_u3058, p2_p1_u3057, p2_p1_u3056, p2_p1_u3055, p2_p1_u3054, p2_p1_u3053, p2_p1_u3052, p2_p1_u3051, p2_p1_u3050, p2_p1_u3049, p2_p1_u3048, p2_p1_u3047, p2_p1_u3046, p2_p1_u3045, p2_p1_u3294, p2_p1_u3295, p2_p1_u3044, p2_p1_u3043, p2_p1_u3042, p2_p1_u3041, p2_p1_u3040, p2_p1_u3039, p2_p1_u3038, p2_p1_u3037, p2_p1_u3036, p2_p1_u3035, p2_p1_u3034, p2_p1_u3033, p2_p1_u3032, p2_p1_u3031, p2_p1_u3030, p2_p1_u3029, p2_p1_u3028, p2_p1_u3027, p2_p1_u3026, p2_p1_u3025, p2_p1_u3024, p2_p1_u3023, p2_p1_u3022, p2_p1_u3021, p2_p1_u3020, p2_p1_u3019, p2_p1_u3018, p2_p1_u3017, p2_p1_u3016, p2_p1_u3015, p2_p1_u3296, p2_p1_u3014, p2_p1_u3013, p2_p1_u3012, p2_p1_u3011, p2_p1_u3010, p2_p1_u3009, p2_p1_u3008, p2_p1_u3007, p2_p1_u3006, p2_p1_u3005, p2_p1_u3004, p2_p1_u3003, p2_p1_u3002, p2_p1_u3001, p2_p1_u3000, p2_p1_u2999, p2_p1_u2998, p2_p1_u2997, p2_p1_u2996, p2_p1_u2995, p2_p1_u2994, p2_p1_u2993, p2_p1_u2992, p2_p1_u2991, p2_p1_u2990, p2_p1_u2989, p2_p1_u2988, p2_p1_u2987, p2_p1_u2986, p2_p1_u2985, p2_p1_u2984, p2_p1_u2983, p2_p1_u2982, p2_p1_u2981, p2_p1_u2980, p2_p1_u2979, p2_p1_u2978, p2_p1_u2977, p2_p1_u2976, p2_p1_u2975, p2_p1_u2974, p2_p1_u2973, p2_p1_u2972, p2_p1_u2971, p2_p1_u2970, p2_p1_u2969, p2_p1_u2968, p2_p1_u2967, p2_p1_u2966, p2_p1_u2965, p2_p1_u2964, p2_p1_u2963, p2_p1_u2962, p2_p1_u2961, p2_p1_u2960, p2_p1_u2959, p2_p1_u2958, p2_p1_u2957, p2_p1_u2956, p2_p1_u2955, p2_p1_u2954, p2_p1_u2953, p2_p1_u2952, p2_p1_u2951, p2_p1_u2950, p2_p1_u2949, p2_p1_u2948, p2_p1_u2947, p2_p1_u2946, p2_p1_u2945, p2_p1_u2944, p2_p1_u2943, p2_p1_u2942, p2_p1_u2941, p2_p1_u2940, p2_p1_u2939, p2_p1_u2938, p2_p1_u2937, p2_p1_u2936, p2_p1_u2935, p2_p1_u2934, p2_p1_u2933, p2_p1_u2932, p2_p1_u2931, p2_p1_u2930, p2_p1_u2929, p2_p1_u2928, p2_p1_u2927, p2_p1_u2926, p2_p1_u2925, p2_p1_u2924, p2_p1_u2923, p2_p1_u2922, p2_p1_u2921, p2_p1_u2920, p2_p1_u2919, p2_p1_u2918, p2_p1_u2917, p2_p1_u2916, p2_p1_u2915, p2_p1_u2914, p2_p1_u2913, p2_p1_u2912, p2_p1_u2911, p2_p1_u2910, p2_p1_u2909, p2_p1_u2908, p2_p1_u2907, p2_p1_u2906, p2_p1_u2905, p2_p1_u2904, p2_p1_u2903, p2_p1_u2902, p2_p1_u2901, p2_p1_u2900, p2_p1_u2899, p2_p1_u2898, p2_p1_u2897, p2_p1_u2896, p2_p1_u2895, p2_p1_u2894, p2_p1_u2893, p2_p1_u2892, p2_p1_u2891, p2_p1_u2890, p2_p1_u2889, p2_p1_u2888, p2_p1_u2887, p2_p1_u2886, p2_p1_u2885, p2_p1_u2884, p2_p1_u3298, p2_p1_u3299, p2_p1_u3302, p2_p1_u3303, p2_p1_u3304, p2_p1_u2883, p2_p1_u2882, p2_p1_u2881, p2_p1_u2880, p2_p1_u2879, p2_p1_u2878, p2_p1_u2877, p2_p1_u2876, p2_p1_u2875, p2_p1_u2874, p2_p1_u2873, p2_p1_u2872, p2_p1_u2871, p2_p1_u2870, p2_p1_u2869, p2_p1_u2868, p2_p1_u2867, p2_p1_u2866, p2_p1_u2865, p2_p1_u2864, p2_p1_u2863, p2_p1_u2862, p2_p1_u2861, p2_p1_u2860, p2_p1_u2859, p2_p1_u2858, p2_p1_u2857, p2_p1_u2856, p2_p1_u2855, p2_p1_u2854, p2_p1_u2853, p2_p1_u2852, p2_p1_u2851, p2_p1_u2850, p2_p1_u2849, p2_p1_u2848, p2_p1_u2847, p2_p1_u2846, p2_p1_u2845, p2_p1_u2844, p2_p1_u2843, p2_p1_u2842, p2_p1_u2841, p2_p1_u2840, p2_p1_u2839, p2_p1_u2838, p2_p1_u2837, p2_p1_u2836, p2_p1_u2835, p2_p1_u2834, p2_p1_u2833, p2_p1_u2832, p2_p1_u2831, p2_p1_u2830, p2_p1_u2829, p2_p1_u2828, p2_p1_u2827, p2_p1_u2826, p2_p1_u2825, p2_p1_u2824, p2_p1_u2823, p2_p1_u2822, p2_p1_u2821, p2_p1_u2820, p2_p1_u2819, p2_p1_u2818, p2_p1_u2817, p2_p1_u2816, p2_p1_u2815, p2_p1_u2814, p2_p1_u2813, p2_p1_u2812, p2_p1_u2811, p2_p1_u2810, p2_p1_u2809, p2_p1_u2808, p2_p1_u2807, p2_p1_u2806, p2_p1_u2805, p2_p1_u2804, p2_p1_u2803, p2_p1_u2802, p2_p1_u2801, p2_p1_u2800, p2_p1_u2799, p2_p1_u2798, p2_p1_u2797, p2_p1_u2796, p2_p1_u2795, p2_p1_u2794, p2_p1_u2793, p2_p1_u2792, p2_p1_u2791, p2_p1_u2790, p2_p1_u2789, p2_p1_u2788, p2_p1_u2787, p2_p1_u2786, p2_p1_u2785, p2_p1_u2784, p2_p1_u2783, p2_p1_u2782, p2_p1_u2781, p2_p1_u2780, p2_p1_u2779, p2_p1_u2778, p2_p1_u2777, p2_p1_u2776, p2_p1_u2775, p2_p1_u2774, p2_p1_u2773, p2_p1_u2772, p2_p1_u2771, p2_p1_u2770, p2_p1_u2769, p2_p1_u2768, p2_p1_u2767, p2_p1_u2766, p2_p1_u2765, p2_p1_u2764, p2_p1_u2763, p2_p1_u2762, p2_p1_u2761, p2_p1_u2760, p2_p1_u2759, p2_p1_u2758, p2_p1_u2757, p2_p1_u2756, p2_p1_u2755, p2_p1_u2754, p2_p1_u2753, p2_p1_u2752, p2_p1_u2751, p2_p1_u2750, p2_p1_u2749, p2_p1_u2748, p2_p1_u2747, p2_p1_u2746, p2_p1_u2745, p2_p1_u2744, p2_p1_u2743, p2_p1_u2742, p2_p1_u2741, p2_p1_u2740, p2_p1_u2739, p2_p1_u2738, p2_p1_u2737, p2_p1_u2736, p2_p1_u2735, p2_p1_u2734, p2_p1_u2733, p2_p1_u2732, p2_p1_u2731, p2_p1_u2730, p2_p1_u2729, p2_p1_u2728, p2_p1_u2727, p2_p1_u2726, p2_p1_u2725, p2_p1_u2724, p2_p1_u2723, p2_p1_u2722, p2_p1_u2721, p2_p1_u2720, p2_p1_u2719, p2_p1_u2718, p2_p1_u2717, p2_p1_u2716, p2_p1_u2715, p2_p1_u2714, p2_p1_u2713, p2_p1_u2712, p2_p1_u2711, p2_p1_u2710, p2_p1_u2709, p2_p1_u2708, p2_p1_u2707, p2_p1_u2706, p2_p1_u2705, p2_p1_u2704, p2_p1_u2703, p2_p1_u2702, p2_p1_u2701, p2_p1_u2700, p2_p1_u2699, p2_p1_u2698, p2_p1_u2697, p2_p1_u2696, p2_p1_u2695, p2_p1_u2694, p2_p1_u2693, p2_p1_u2692, p2_p1_u2691, p2_p1_u2690, p2_p1_u2689, p2_p1_u2688, p2_p1_u2687, p2_p1_u2686, p2_p1_u2685, p2_p1_u2684, p2_p1_u2683, p2_p1_u2682, p2_p1_u2681, p2_p1_u2680, p2_p1_u2679, p2_p1_u2678, p2_p1_u2677, p2_p1_u2676, p2_p1_u2675, p2_p1_u2674, p2_p1_u2673, p2_p1_u2672, p2_p1_u2671, p2_p1_u2670, p2_p1_u2669, p2_p1_u2668, p2_p1_u2667, p2_p1_u2666, p2_p1_u2665, p2_p1_u2664, p2_p1_u2663, p2_p1_u2662, p2_p1_u2661, p2_p1_u2660, p2_p1_u2659, p2_p1_u2658, p2_p1_u2657, p2_p1_u2656, p2_p1_u2655, p2_p1_u3306, p2_p1_u2654, p2_p1_u3307, p2_p1_u3308, p2_p1_u2653, p2_p1_u3309, p2_p1_u2652, p2_p1_u3310, p2_p1_u2651, p2_p1_u3311, p2_p1_u2650, p2_p1_u2649, p2_p1_u3312, p2_p1_u3313);
	if(i == vec_length)begin
		$finish;
	end
end

integer fh_w;
initial begin
	fh_w = $fopen(`out_file, "w");
end
 
initial begin
	//$fsdbDumpfile("SET.fsdb");
	//$fsdbDumpvars;
	//$fsdbDumpMDA;
	$dumpfile("test_result.vcd");
    $dumpvars;

end
endmodule
