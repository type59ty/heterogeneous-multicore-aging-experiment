// b20
// 522 inputs  (32 PIs + 490 PPIs)
// 512 outputs (22 POs + 490 PPOs)
// 19682 gates (16614 gates + 3068 inverters + 0 buffers )
// ( 2036 AND + 480 OR + 13973 NAND + 125 NOR )
// Time: Wed Mar 25 17:47:24 2009
// All copyrigh from NCKU EE TestLAB, Taiwan. [2008.12. WCL]

module b20_ras ( P1_U3355 , P1_U3354 , P1_U3353 , P1_U3352 , P1_U3351 , P1_U3350 ,
             P1_U3349 , P1_U3348 , P1_U3347 , P1_U3346 , P1_U3345 , P1_U3344 ,
             P1_U3343 , P1_U3342 , P1_U3341 , P1_U3340 , P1_U3339 , P1_U3338 ,
             P1_U3337 , P1_U3336 , P1_U3335 , P1_U3334 , P1_U3333 , P1_U3332 ,
             P1_U3331 , P1_U3330 , P1_U3329 , P1_U3328 , P1_U3327 , P1_U3326 ,
             P1_U3325 , P1_U3324 , P1_U3439 , P1_U3440 , P1_U3323 , P1_U3322 ,
             P1_U3321 , P1_U3320 , P1_U3319 , P1_U3318 , P1_U3317 , P1_U3316 ,
             P1_U3315 , P1_U3314 , P1_U3313 , P1_U3312 , P1_U3311 , P1_U3310 ,
             P1_U3309 , P1_U3308 , P1_U3307 , P1_U3306 , P1_U3305 , P1_U3304 ,
             P1_U3303 , P1_U3302 , P1_U3301 , P1_U3300 , P1_U3299 , P1_U3298 ,
             P1_U3297 , P1_U3296 , P1_U3295 , P1_U3294 , P1_U3453 , P1_U3456 ,
             P1_U3459 , P1_U3462 , P1_U3465 , P1_U3468 , P1_U3471 , P1_U3474 ,
             P1_U3477 , P1_U3480 , P1_U3483 , P1_U3486 , P1_U3489 , P1_U3492 ,
             P1_U3495 , P1_U3498 , P1_U3501 , P1_U3504 , P1_U3507 , P1_U3509 ,
             P1_U3510 , P1_U3511 , P1_U3512 , P1_U3513 , P1_U3514 , P1_U3515 ,
             P1_U3516 , P1_U3517 , P1_U3518 , P1_U3519 , P1_U3520 , P1_U3521 ,
             P1_U3522 , P1_U3523 , P1_U3524 , P1_U3525 , P1_U3526 , P1_U3527 ,
             P1_U3528 , P1_U3529 , P1_U3530 , P1_U3531 , P1_U3532 , P1_U3533 ,
             P1_U3534 , P1_U3535 , P1_U3536 , P1_U3537 , P1_U3538 , P1_U3539 ,
             P1_U3540 , P1_U3541 , P1_U3542 , P1_U3543 , P1_U3544 , P1_U3545 ,
             P1_U3546 , P1_U3547 , P1_U3548 , P1_U3549 , P1_U3550 , P1_U3551 ,
             P1_U3552 , P1_U3553 , P1_U3293 , P1_U3292 , P1_U3291 , P1_U3290 ,
             P1_U3289 , P1_U3288 , P1_U3287 , P1_U3286 , P1_U3285 , P1_U3284 ,
             P1_U3283 , P1_U3282 , P1_U3281 , P1_U3280 , P1_U3279 , P1_U3278 ,
             P1_U3277 , P1_U3276 , P1_U3275 , P1_U3274 , P1_U3273 , P1_U3272 ,
             P1_U3271 , P1_U3270 , P1_U3269 , P1_U3268 , P1_U3267 , P1_U3266 ,
             P1_U3265 , P1_U3356 , P1_U3264 , P1_U3263 , P1_U3262 , P1_U3261 ,
             P1_U3260 , P1_U3259 , P1_U3258 , P1_U3257 , P1_U3256 , P1_U3255 ,
             P1_U3254 , P1_U3253 , P1_U3252 , P1_U3251 , P1_U3250 , P1_U3249 ,
             P1_U3248 , P1_U3247 , P1_U3246 , P1_U3245 , P1_U3244 , P1_U3243 ,
             P1_U3554 , P1_U3555 , P1_U3556 , P1_U3557 , P1_U3558 , P1_U3559 ,
             P1_U3560 , P1_U3561 , P1_U3562 , P1_U3563 , P1_U3564 , P1_U3565 ,
             P1_U3566 , P1_U3567 , P1_U3568 , P1_U3569 , P1_U3570 , P1_U3571 ,
             P1_U3572 , P1_U3573 , P1_U3574 , P1_U3575 , P1_U3576 , P1_U3577 ,
             P1_U3578 , P1_U3579 , P1_U3580 , P1_U3581 , P1_U3582 , P1_U3583 ,
             P1_U3584 , P1_U3585 , P1_U3242 , P1_U3241 , P1_U3240 , P1_U3239 ,
             P1_U3238 , P1_U3237 , P1_U3236 , P1_U3235 , P1_U3234 , P1_U3233 ,
             P1_U3232 , P1_U3231 , P1_U3230 , P1_U3229 , P1_U3228 , P1_U3227 ,
             P1_U3226 , P1_U3225 , P1_U3224 , P1_U3223 , P1_U3222 , P1_U3221 ,
             P1_U3220 , P1_U3219 , P1_U3218 , P1_U3217 , P1_U3216 , P1_U3215 ,
             P1_U3214 , P1_U3213 , P1_U3086 , P1_U3085 , P1_U3973 , P2_U3295 ,
             P2_U3294 , P2_U3293 , P2_U3292 , P2_U3291 , P2_U3290 , P2_U3289 ,
             P2_U3288 , P2_U3287 , P2_U3286 , P2_U3285 , P2_U3284 , P2_U3283 ,
             P2_U3282 , P2_U3281 , P2_U3280 , P2_U3279 , P2_U3278 , P2_U3277 ,
             P2_U3276 , P2_U3275 , P2_U3274 , P2_U3273 , P2_U3272 , P2_U3271 ,
             P2_U3270 , P2_U3269 , P2_U3268 , P2_U3267 , P2_U3266 , P2_U3265 ,
             P2_U3264 , P2_U3376 , P2_U3377 , P2_U3263 , P2_U3262 , P2_U3261 ,
             P2_U3260 , P2_U3259 , P2_U3258 , P2_U3257 , P2_U3256 , P2_U3255 ,
             P2_U3254 , P2_U3253 , P2_U3252 , P2_U3251 , P2_U3250 , P2_U3249 ,
             P2_U3248 , P2_U3247 , P2_U3246 , P2_U3245 , P2_U3244 , P2_U3243 ,
             P2_U3242 , P2_U3241 , P2_U3240 , P2_U3239 , P2_U3238 , P2_U3237 ,
             P2_U3236 , P2_U3235 , P2_U3234 , P2_U3390 , P2_U3393 , P2_U3396 ,
             P2_U3399 , P2_U3402 , P2_U3405 , P2_U3408 , P2_U3411 , P2_U3414 ,
             P2_U3417 , P2_U3420 , P2_U3423 , P2_U3426 , P2_U3429 , P2_U3432 ,
             P2_U3435 , P2_U3438 , P2_U3441 , P2_U3444 , P2_U3446 , P2_U3447 ,
             P2_U3448 , P2_U3449 , P2_U3450 , P2_U3451 , P2_U3452 , P2_U3453 ,
             P2_U3454 , P2_U3455 , P2_U3456 , P2_U3457 , P2_U3458 , P2_U3459 ,
             P2_U3460 , P2_U3461 , P2_U3462 , P2_U3463 , P2_U3464 , P2_U3465 ,
             P2_U3466 , P2_U3467 , P2_U3468 , P2_U3469 , P2_U3470 , P2_U3471 ,
             P2_U3472 , P2_U3473 , P2_U3474 , P2_U3475 , P2_U3476 , P2_U3477 ,
             P2_U3478 , P2_U3479 , P2_U3480 , P2_U3481 , P2_U3482 , P2_U3483 ,
             P2_U3484 , P2_U3485 , P2_U3486 , P2_U3487 , P2_U3488 , P2_U3489 ,
             P2_U3490 , P2_U3233 , P2_U3232 , P2_U3231 , P2_U3230 , P2_U3229 ,
             P2_U3228 , P2_U3227 , P2_U3226 , P2_U3225 , P2_U3224 , P2_U3223 ,
             P2_U3222 , P2_U3221 , P2_U3220 , P2_U3219 , P2_U3218 , P2_U3217 ,
             P2_U3216 , P2_U3215 , P2_U3214 , P2_U3213 , P2_U3212 , P2_U3211 ,
             P2_U3210 , P2_U3209 , P2_U3208 , P2_U3207 , P2_U3206 , P2_U3205 ,
             P2_U3204 , P2_U3203 , P2_U3202 , P2_U3201 , P2_U3200 , P2_U3199 ,
             P2_U3198 , P2_U3197 , P2_U3196 , P2_U3195 , P2_U3194 , P2_U3193 ,
             P2_U3192 , P2_U3191 , P2_U3190 , P2_U3189 , P2_U3188 , P2_U3187 ,
             P2_U3186 , P2_U3185 , P2_U3184 , P2_U3183 , P2_U3182 , P2_U3491 ,
             P2_U3492 , P2_U3493 , P2_U3494 , P2_U3495 , P2_U3496 , P2_U3497 ,
             P2_U3498 , P2_U3499 , P2_U3500 , P2_U3501 , P2_U3502 , P2_U3503 ,
             P2_U3504 , P2_U3505 , P2_U3506 , P2_U3507 , P2_U3508 , P2_U3509 ,
             P2_U3510 , P2_U3511 , P2_U3512 , P2_U3513 , P2_U3514 , P2_U3515 ,
             P2_U3516 , P2_U3517 , P2_U3518 , P2_U3519 , P2_U3520 , P2_U3521 ,
             P2_U3522 , P2_U3296 , P2_U3181 , P2_U3180 , P2_U3179 , P2_U3178 ,
             P2_U3177 , P2_U3176 , P2_U3175 , P2_U3174 , P2_U3173 , P2_U3172 ,
             P2_U3171 , P2_U3170 , P2_U3169 , P2_U3168 , P2_U3167 , P2_U3166 ,
             P2_U3165 , P2_U3164 , P2_U3163 , P2_U3162 , P2_U3161 , P2_U3160 ,
             P2_U3159 , P2_U3158 , P2_U3157 , P2_U3156 , P2_U3155 , P2_U3154 ,
             P2_U3153 , P2_U3151 , P2_U3150 , P2_U3893 , ADD_1068_U4 , ADD_1068_U55 ,
             ADD_1068_U56 , ADD_1068_U57 , ADD_1068_U58 , ADD_1068_U59 , ADD_1068_U60 , ADD_1068_U61 ,
             ADD_1068_U62 , ADD_1068_U63 , ADD_1068_U47 , ADD_1068_U48 , ADD_1068_U49 , ADD_1068_U50 ,
             ADD_1068_U51 , ADD_1068_U52 , ADD_1068_U53 , ADD_1068_U54 , ADD_1068_U5 , ADD_1068_U46 ,
             U126 , U123 ,
             P1_IR_REG_0_ , P1_IR_REG_1_ , P1_IR_REG_2_ , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ ,
             P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_10_ , P1_IR_REG_11_ ,
             P1_IR_REG_12_ , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_ ,
             P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_20_ , P1_IR_REG_21_ , P1_IR_REG_22_ , P1_IR_REG_23_ ,
             P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ , P1_IR_REG_27_ , P1_IR_REG_28_ , P1_IR_REG_29_ ,
             P1_IR_REG_30_ , P1_IR_REG_31_ , P1_D_REG_0_ , P1_D_REG_1_ , P1_D_REG_2_ , P1_D_REG_3_ ,
             P1_D_REG_4_ , P1_D_REG_5_ , P1_D_REG_6_ , P1_D_REG_7_ , P1_D_REG_8_ , P1_D_REG_9_ ,
             P1_D_REG_10_ , P1_D_REG_11_ , P1_D_REG_12_ , P1_D_REG_13_ , P1_D_REG_14_ , P1_D_REG_15_ ,
             P1_D_REG_16_ , P1_D_REG_17_ , P1_D_REG_18_ , P1_D_REG_19_ , P1_D_REG_20_ , P1_D_REG_21_ ,
             P1_D_REG_22_ , P1_D_REG_23_ , P1_D_REG_24_ , P1_D_REG_25_ , P1_D_REG_26_ , P1_D_REG_27_ ,
             P1_D_REG_28_ , P1_D_REG_29_ , P1_D_REG_30_ , P1_D_REG_31_ , P1_REG0_REG_0_ , P1_REG0_REG_1_ ,
             P1_REG0_REG_2_ , P1_REG0_REG_3_ , P1_REG0_REG_4_ , P1_REG0_REG_5_ , P1_REG0_REG_6_ , P1_REG0_REG_7_ ,
             P1_REG0_REG_8_ , P1_REG0_REG_9_ , P1_REG0_REG_10_ , P1_REG0_REG_11_ , P1_REG0_REG_12_ , P1_REG0_REG_13_ ,
             P1_REG0_REG_14_ , P1_REG0_REG_15_ , P1_REG0_REG_16_ , P1_REG0_REG_17_ , P1_REG0_REG_18_ , P1_REG0_REG_19_ ,
             P1_REG0_REG_20_ , P1_REG0_REG_21_ , P1_REG0_REG_22_ , P1_REG0_REG_23_ , P1_REG0_REG_24_ , P1_REG0_REG_25_ ,
             P1_REG0_REG_26_ , P1_REG0_REG_27_ , P1_REG0_REG_28_ , P1_REG0_REG_29_ , P1_REG0_REG_30_ , P1_REG0_REG_31_ ,
             P1_REG1_REG_0_ , P1_REG1_REG_1_ , P1_REG1_REG_2_ , P1_REG1_REG_3_ , P1_REG1_REG_4_ , P1_REG1_REG_5_ ,
             P1_REG1_REG_6_ , P1_REG1_REG_7_ , P1_REG1_REG_8_ , P1_REG1_REG_9_ , P1_REG1_REG_10_ , P1_REG1_REG_11_ ,
             P1_REG1_REG_12_ , P1_REG1_REG_13_ , P1_REG1_REG_14_ , P1_REG1_REG_15_ , P1_REG1_REG_16_ , P1_REG1_REG_17_ ,
             P1_REG1_REG_18_ , P1_REG1_REG_19_ , P1_REG1_REG_20_ , P1_REG1_REG_21_ , P1_REG1_REG_22_ , P1_REG1_REG_23_ ,
             P1_REG1_REG_24_ , P1_REG1_REG_25_ , P1_REG1_REG_26_ , P1_REG1_REG_27_ , P1_REG1_REG_28_ , P1_REG1_REG_29_ ,
             P1_REG1_REG_30_ , P1_REG1_REG_31_ , P1_REG2_REG_0_ , P1_REG2_REG_1_ , P1_REG2_REG_2_ , P1_REG2_REG_3_ ,
             P1_REG2_REG_4_ , P1_REG2_REG_5_ , P1_REG2_REG_6_ , P1_REG2_REG_7_ , P1_REG2_REG_8_ , P1_REG2_REG_9_ ,
             P1_REG2_REG_10_ , P1_REG2_REG_11_ , P1_REG2_REG_12_ , P1_REG2_REG_13_ , P1_REG2_REG_14_ , P1_REG2_REG_15_ ,
             P1_REG2_REG_16_ , P1_REG2_REG_17_ , P1_REG2_REG_18_ , P1_REG2_REG_19_ , P1_REG2_REG_20_ , P1_REG2_REG_21_ ,
             P1_REG2_REG_22_ , P1_REG2_REG_23_ , P1_REG2_REG_24_ , P1_REG2_REG_25_ , P1_REG2_REG_26_ , P1_REG2_REG_27_ ,
             P1_REG2_REG_28_ , P1_REG2_REG_29_ , P1_REG2_REG_30_ , P1_REG2_REG_31_ , P1_ADDR_REG_19_ , P1_ADDR_REG_18_ ,
             P1_ADDR_REG_17_ , P1_ADDR_REG_16_ , P1_ADDR_REG_15_ , P1_ADDR_REG_14_ , P1_ADDR_REG_13_ , P1_ADDR_REG_12_ ,
             P1_ADDR_REG_11_ , P1_ADDR_REG_10_ , P1_ADDR_REG_9_ , P1_ADDR_REG_8_ , P1_ADDR_REG_7_ , P1_ADDR_REG_6_ ,
             P1_ADDR_REG_5_ , P1_ADDR_REG_4_ , P1_ADDR_REG_3_ , P1_ADDR_REG_2_ , P1_ADDR_REG_1_ , P1_ADDR_REG_0_ ,
             P1_DATAO_REG_0_ , P1_DATAO_REG_1_ , P1_DATAO_REG_2_ , P1_DATAO_REG_3_ , P1_DATAO_REG_4_ , P1_DATAO_REG_5_ ,
             P1_DATAO_REG_6_ , P1_DATAO_REG_7_ , P1_DATAO_REG_8_ , P1_DATAO_REG_9_ , P1_DATAO_REG_10_ , P1_DATAO_REG_11_ ,
             P1_DATAO_REG_12_ , P1_DATAO_REG_13_ , P1_DATAO_REG_14_ , P1_DATAO_REG_15_ , P1_DATAO_REG_16_ , P1_DATAO_REG_17_ ,
             P1_DATAO_REG_18_ , P1_DATAO_REG_19_ , P1_DATAO_REG_20_ , P1_DATAO_REG_21_ , P1_DATAO_REG_22_ , P1_DATAO_REG_23_ ,
             P1_DATAO_REG_24_ , P1_DATAO_REG_25_ , P1_DATAO_REG_26_ , P1_DATAO_REG_27_ , P1_DATAO_REG_28_ , P1_DATAO_REG_29_ ,
             P1_DATAO_REG_30_ , P1_DATAO_REG_31_ , P1_B_REG , P1_REG3_REG_15_ , P1_REG3_REG_26_ , P1_REG3_REG_6_ ,
             P1_REG3_REG_18_ , P1_REG3_REG_2_ , P1_REG3_REG_11_ , P1_REG3_REG_22_ , P1_REG3_REG_13_ , P1_REG3_REG_20_ ,
             P1_REG3_REG_0_ , P1_REG3_REG_9_ , P1_REG3_REG_4_ , P1_REG3_REG_24_ , P1_REG3_REG_17_ , P1_REG3_REG_5_ ,
             P1_REG3_REG_16_ , P1_REG3_REG_25_ , P1_REG3_REG_12_ , P1_REG3_REG_21_ , P1_REG3_REG_1_ , P1_REG3_REG_8_ ,
             P1_REG3_REG_28_ , P1_REG3_REG_19_ , P1_REG3_REG_3_ , P1_REG3_REG_10_ , P1_REG3_REG_23_ , P1_REG3_REG_14_ ,
             P1_REG3_REG_27_ , P1_REG3_REG_7_ , P1_STATE_REG , P1_RD_REG , P1_WR_REG , P2_IR_REG_0_ ,
             P2_IR_REG_1_ , P2_IR_REG_2_ , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ , P2_IR_REG_6_ ,
             P2_IR_REG_7_ , P2_IR_REG_8_ , P2_IR_REG_9_ , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_ ,
             P2_IR_REG_13_ , P2_IR_REG_14_ , P2_IR_REG_15_ , P2_IR_REG_16_ , P2_IR_REG_17_ , P2_IR_REG_18_ ,
             P2_IR_REG_19_ , P2_IR_REG_20_ , P2_IR_REG_21_ , P2_IR_REG_22_ , P2_IR_REG_23_ , P2_IR_REG_24_ ,
             P2_IR_REG_25_ , P2_IR_REG_26_ , P2_IR_REG_27_ , P2_IR_REG_28_ , P2_IR_REG_29_ , P2_IR_REG_30_ ,
             P2_IR_REG_31_ , P2_D_REG_0_ , P2_D_REG_1_ , P2_D_REG_2_ , P2_D_REG_3_ , P2_D_REG_4_ ,
             P2_D_REG_5_ , P2_D_REG_6_ , P2_D_REG_7_ , P2_D_REG_8_ , P2_D_REG_9_ , P2_D_REG_10_ ,
             P2_D_REG_11_ , P2_D_REG_12_ , P2_D_REG_13_ , P2_D_REG_14_ , P2_D_REG_15_ , P2_D_REG_16_ ,
             P2_D_REG_17_ , P2_D_REG_18_ , P2_D_REG_19_ , P2_D_REG_20_ , P2_D_REG_21_ , P2_D_REG_22_ ,
             P2_D_REG_23_ , P2_D_REG_24_ , P2_D_REG_25_ , P2_D_REG_26_ , P2_D_REG_27_ , P2_D_REG_28_ ,
             P2_D_REG_29_ , P2_D_REG_30_ , P2_D_REG_31_ , P2_REG0_REG_0_ , P2_REG0_REG_1_ , P2_REG0_REG_2_ ,
             P2_REG0_REG_3_ , P2_REG0_REG_4_ , P2_REG0_REG_5_ , P2_REG0_REG_6_ , P2_REG0_REG_7_ , P2_REG0_REG_8_ ,
             P2_REG0_REG_9_ , P2_REG0_REG_10_ , P2_REG0_REG_11_ , P2_REG0_REG_12_ , P2_REG0_REG_13_ , P2_REG0_REG_14_ ,
             P2_REG0_REG_15_ , P2_REG0_REG_16_ , P2_REG0_REG_17_ , P2_REG0_REG_18_ , P2_REG0_REG_19_ , P2_REG0_REG_20_ ,
             P2_REG0_REG_21_ , P2_REG0_REG_22_ , P2_REG0_REG_23_ , P2_REG0_REG_24_ , P2_REG0_REG_25_ , P2_REG0_REG_26_ ,
             P2_REG0_REG_27_ , P2_REG0_REG_28_ , P2_REG0_REG_29_ , P2_REG0_REG_30_ , P2_REG0_REG_31_ , P2_REG1_REG_0_ ,
             P2_REG1_REG_1_ , P2_REG1_REG_2_ , P2_REG1_REG_3_ , P2_REG1_REG_4_ , P2_REG1_REG_5_ , P2_REG1_REG_6_ ,
             P2_REG1_REG_7_ , P2_REG1_REG_8_ , P2_REG1_REG_9_ , P2_REG1_REG_10_ , P2_REG1_REG_11_ , P2_REG1_REG_12_ ,
             P2_REG1_REG_13_ , P2_REG1_REG_14_ , P2_REG1_REG_15_ , P2_REG1_REG_16_ , P2_REG1_REG_17_ , P2_REG1_REG_18_ ,
             P2_REG1_REG_19_ , P2_REG1_REG_20_ , P2_REG1_REG_21_ , P2_REG1_REG_22_ , P2_REG1_REG_23_ , P2_REG1_REG_24_ ,
             P2_REG1_REG_25_ , P2_REG1_REG_26_ , P2_REG1_REG_27_ , P2_REG1_REG_28_ , P2_REG1_REG_29_ , P2_REG1_REG_30_ ,
             P2_REG1_REG_31_ , P2_REG2_REG_0_ , P2_REG2_REG_1_ , P2_REG2_REG_2_ , P2_REG2_REG_3_ , P2_REG2_REG_4_ ,
             P2_REG2_REG_5_ , P2_REG2_REG_6_ , P2_REG2_REG_7_ , P2_REG2_REG_8_ , P2_REG2_REG_9_ , P2_REG2_REG_10_ ,
             P2_REG2_REG_11_ , P2_REG2_REG_12_ , P2_REG2_REG_13_ , P2_REG2_REG_14_ , P2_REG2_REG_15_ , P2_REG2_REG_16_ ,
             P2_REG2_REG_17_ , P2_REG2_REG_18_ , P2_REG2_REG_19_ , P2_REG2_REG_20_ , P2_REG2_REG_21_ , P2_REG2_REG_22_ ,
             P2_REG2_REG_23_ , P2_REG2_REG_24_ , P2_REG2_REG_25_ , P2_REG2_REG_26_ , P2_REG2_REG_27_ , P2_REG2_REG_28_ ,
             P2_REG2_REG_29_ , P2_REG2_REG_30_ , P2_REG2_REG_31_ , P2_ADDR_REG_19_ , P2_ADDR_REG_18_ , P2_ADDR_REG_17_ ,
             P2_ADDR_REG_16_ , P2_ADDR_REG_15_ , P2_ADDR_REG_14_ , P2_ADDR_REG_13_ , P2_ADDR_REG_12_ , P2_ADDR_REG_11_ ,
             P2_ADDR_REG_10_ , P2_ADDR_REG_9_ , P2_ADDR_REG_8_ , P2_ADDR_REG_7_ , P2_ADDR_REG_6_ , P2_ADDR_REG_5_ ,
             P2_ADDR_REG_4_ , P2_ADDR_REG_3_ , P2_ADDR_REG_2_ , P2_ADDR_REG_1_ , P2_ADDR_REG_0_ , P2_DATAO_REG_0_ ,
             P2_DATAO_REG_1_ , P2_DATAO_REG_2_ , P2_DATAO_REG_3_ , P2_DATAO_REG_4_ , P2_DATAO_REG_5_ , P2_DATAO_REG_6_ ,
             P2_DATAO_REG_7_ , P2_DATAO_REG_8_ , P2_DATAO_REG_9_ , P2_DATAO_REG_10_ , P2_DATAO_REG_11_ , P2_DATAO_REG_12_ ,
             P2_DATAO_REG_13_ , P2_DATAO_REG_14_ , P2_DATAO_REG_15_ , P2_DATAO_REG_16_ , P2_DATAO_REG_17_ , P2_DATAO_REG_18_ ,
             P2_DATAO_REG_19_ , P2_DATAO_REG_20_ , P2_DATAO_REG_21_ , P2_DATAO_REG_22_ , P2_DATAO_REG_23_ , P2_DATAO_REG_24_ ,
             P2_DATAO_REG_25_ , P2_DATAO_REG_26_ , P2_DATAO_REG_27_ , P2_DATAO_REG_28_ , P2_DATAO_REG_29_ , P2_DATAO_REG_30_ ,
             P2_DATAO_REG_31_ , P2_B_REG , P2_REG3_REG_15_ , P2_REG3_REG_26_ , P2_REG3_REG_6_ , P2_REG3_REG_18_ ,
             P2_REG3_REG_2_ , P2_REG3_REG_11_ , P2_REG3_REG_22_ , P2_REG3_REG_13_ , P2_REG3_REG_20_ , P2_REG3_REG_0_ ,
             P2_REG3_REG_9_ , P2_REG3_REG_4_ , P2_REG3_REG_24_ , P2_REG3_REG_17_ , P2_REG3_REG_5_ , P2_REG3_REG_16_ ,
             P2_REG3_REG_25_ , P2_REG3_REG_12_ , P2_REG3_REG_21_ , P2_REG3_REG_1_ , P2_REG3_REG_8_ , P2_REG3_REG_28_ ,
             P2_REG3_REG_19_ , P2_REG3_REG_3_ , P2_REG3_REG_10_ , P2_REG3_REG_23_ , P2_REG3_REG_14_ , P2_REG3_REG_27_ ,
             P2_REG3_REG_7_ , P2_STATE_REG , P2_RD_REG , P2_WR_REG , SI_31_ , SI_30_ ,
             SI_29_ , SI_28_ , SI_27_ , SI_26_ , SI_25_ , SI_24_ ,
             SI_23_ , SI_22_ , SI_21_ , SI_20_ , SI_19_ , SI_18_ ,
             SI_17_ , SI_16_ , SI_15_ , SI_14_ , SI_13_ , SI_12_ ,
             SI_11_ , SI_10_ , SI_9_ , SI_8_ , SI_7_ , SI_6_ ,
             SI_5_ , SI_4_ , SI_3_ , SI_2_ , SI_1_ , SI_0_ );

output ADD_1068_U4 , ADD_1068_U55 , ADD_1068_U56 , ADD_1068_U57 , ADD_1068_U58 , ADD_1068_U59;
output ADD_1068_U60 , ADD_1068_U61 , ADD_1068_U62 , ADD_1068_U63 , ADD_1068_U47 , ADD_1068_U48;
output ADD_1068_U49 , ADD_1068_U50 , ADD_1068_U51 , ADD_1068_U52 , ADD_1068_U53 , ADD_1068_U54;
output ADD_1068_U5 , ADD_1068_U46 , U126 , U123;
output P1_U3355 , P1_U3354 , P1_U3353 , P1_U3352 , P1_U3351 , P1_U3350 , P1_U3349;
output P1_U3348 , P1_U3347 , P1_U3346 , P1_U3345 , P1_U3344 , P1_U3343 , P1_U3342;
output P1_U3341 , P1_U3340 , P1_U3339 , P1_U3338 , P1_U3337 , P1_U3336 , P1_U3335;
output P1_U3334 , P1_U3333 , P1_U3332 , P1_U3331 , P1_U3330 , P1_U3329 , P1_U3328;
output P1_U3327 , P1_U3326 , P1_U3325 , P1_U3324 , P1_U3439 , P1_U3440 , P1_U3323;
output P1_U3322 , P1_U3321 , P1_U3320 , P1_U3319 , P1_U3318 , P1_U3317 , P1_U3316;
output P1_U3315 , P1_U3314 , P1_U3313 , P1_U3312 , P1_U3311 , P1_U3310 , P1_U3309;
output P1_U3308 , P1_U3307 , P1_U3306 , P1_U3305 , P1_U3304 , P1_U3303 , P1_U3302;
output P1_U3301 , P1_U3300 , P1_U3299 , P1_U3298 , P1_U3297 , P1_U3296 , P1_U3295;
output P1_U3294 , P1_U3453 , P1_U3456 , P1_U3459 , P1_U3462 , P1_U3465 , P1_U3468;
output P1_U3471 , P1_U3474 , P1_U3477 , P1_U3480 , P1_U3483 , P1_U3486 , P1_U3489;
output P1_U3492 , P1_U3495 , P1_U3498 , P1_U3501 , P1_U3504 , P1_U3507 , P1_U3509;
output P1_U3510 , P1_U3511 , P1_U3512 , P1_U3513 , P1_U3514 , P1_U3515 , P1_U3516;
output P1_U3517 , P1_U3518 , P1_U3519 , P1_U3520 , P1_U3521 , P1_U3522 , P1_U3523;
output P1_U3524 , P1_U3525 , P1_U3526 , P1_U3527 , P1_U3528 , P1_U3529 , P1_U3530;
output P1_U3531 , P1_U3532 , P1_U3533 , P1_U3534 , P1_U3535 , P1_U3536 , P1_U3537;
output P1_U3538 , P1_U3539 , P1_U3540 , P1_U3541 , P1_U3542 , P1_U3543 , P1_U3544;
output P1_U3545 , P1_U3546 , P1_U3547 , P1_U3548 , P1_U3549 , P1_U3550 , P1_U3551;
output P1_U3552 , P1_U3553 , P1_U3293 , P1_U3292 , P1_U3291 , P1_U3290 , P1_U3289;
output P1_U3288 , P1_U3287 , P1_U3286 , P1_U3285 , P1_U3284 , P1_U3283 , P1_U3282;
output P1_U3281 , P1_U3280 , P1_U3279 , P1_U3278 , P1_U3277 , P1_U3276 , P1_U3275;
output P1_U3274 , P1_U3273 , P1_U3272 , P1_U3271 , P1_U3270 , P1_U3269 , P1_U3268;
output P1_U3267 , P1_U3266 , P1_U3265 , P1_U3356 , P1_U3264 , P1_U3263 , P1_U3262;
output P1_U3261 , P1_U3260 , P1_U3259 , P1_U3258 , P1_U3257 , P1_U3256 , P1_U3255;
output P1_U3254 , P1_U3253 , P1_U3252 , P1_U3251 , P1_U3250 , P1_U3249 , P1_U3248;
output P1_U3247 , P1_U3246 , P1_U3245 , P1_U3244 , P1_U3243 , P1_U3554 , P1_U3555;
output P1_U3556 , P1_U3557 , P1_U3558 , P1_U3559 , P1_U3560 , P1_U3561 , P1_U3562;
output P1_U3563 , P1_U3564 , P1_U3565 , P1_U3566 , P1_U3567 , P1_U3568 , P1_U3569;
output P1_U3570 , P1_U3571 , P1_U3572 , P1_U3573 , P1_U3574 , P1_U3575 , P1_U3576;
output P1_U3577 , P1_U3578 , P1_U3579 , P1_U3580 , P1_U3581 , P1_U3582 , P1_U3583;
output P1_U3584 , P1_U3585 , P1_U3242 , P1_U3241 , P1_U3240 , P1_U3239 , P1_U3238;
output P1_U3237 , P1_U3236 , P1_U3235 , P1_U3234 , P1_U3233 , P1_U3232 , P1_U3231;
output P1_U3230 , P1_U3229 , P1_U3228 , P1_U3227 , P1_U3226 , P1_U3225 , P1_U3224;
output P1_U3223 , P1_U3222 , P1_U3221 , P1_U3220 , P1_U3219 , P1_U3218 , P1_U3217;
output P1_U3216 , P1_U3215 , P1_U3214 , P1_U3213 , P1_U3086 , P1_U3085 , P1_U3973;
output P2_U3295 , P2_U3294 , P2_U3293 , P2_U3292 , P2_U3291 , P2_U3290 , P2_U3289;
output P2_U3288 , P2_U3287 , P2_U3286 , P2_U3285 , P2_U3284 , P2_U3283 , P2_U3282;
output P2_U3281 , P2_U3280 , P2_U3279 , P2_U3278 , P2_U3277 , P2_U3276 , P2_U3275;
output P2_U3274 , P2_U3273 , P2_U3272 , P2_U3271 , P2_U3270 , P2_U3269 , P2_U3268;
output P2_U3267 , P2_U3266 , P2_U3265 , P2_U3264 , P2_U3376 , P2_U3377 , P2_U3263;
output P2_U3262 , P2_U3261 , P2_U3260 , P2_U3259 , P2_U3258 , P2_U3257 , P2_U3256;
output P2_U3255 , P2_U3254 , P2_U3253 , P2_U3252 , P2_U3251 , P2_U3250 , P2_U3249;
output P2_U3248 , P2_U3247 , P2_U3246 , P2_U3245 , P2_U3244 , P2_U3243 , P2_U3242;
output P2_U3241 , P2_U3240 , P2_U3239 , P2_U3238 , P2_U3237 , P2_U3236 , P2_U3235;
output P2_U3234 , P2_U3390 , P2_U3393 , P2_U3396 , P2_U3399 , P2_U3402 , P2_U3405;
output P2_U3408 , P2_U3411 , P2_U3414 , P2_U3417 , P2_U3420 , P2_U3423 , P2_U3426;
output P2_U3429 , P2_U3432 , P2_U3435 , P2_U3438 , P2_U3441 , P2_U3444 , P2_U3446;
output P2_U3447 , P2_U3448 , P2_U3449 , P2_U3450 , P2_U3451 , P2_U3452 , P2_U3453;
output P2_U3454 , P2_U3455 , P2_U3456 , P2_U3457 , P2_U3458 , P2_U3459 , P2_U3460;
output P2_U3461 , P2_U3462 , P2_U3463 , P2_U3464 , P2_U3465 , P2_U3466 , P2_U3467;
output P2_U3468 , P2_U3469 , P2_U3470 , P2_U3471 , P2_U3472 , P2_U3473 , P2_U3474;
output P2_U3475 , P2_U3476 , P2_U3477 , P2_U3478 , P2_U3479 , P2_U3480 , P2_U3481;
output P2_U3482 , P2_U3483 , P2_U3484 , P2_U3485 , P2_U3486 , P2_U3487 , P2_U3488;
output P2_U3489 , P2_U3490 , P2_U3233 , P2_U3232 , P2_U3231 , P2_U3230 , P2_U3229;
output P2_U3228 , P2_U3227 , P2_U3226 , P2_U3225 , P2_U3224 , P2_U3223 , P2_U3222;
output P2_U3221 , P2_U3220 , P2_U3219 , P2_U3218 , P2_U3217 , P2_U3216 , P2_U3215;
output P2_U3214 , P2_U3213 , P2_U3212 , P2_U3211 , P2_U3210 , P2_U3209 , P2_U3208;
output P2_U3207 , P2_U3206 , P2_U3205 , P2_U3204 , P2_U3203 , P2_U3202 , P2_U3201;
output P2_U3200 , P2_U3199 , P2_U3198 , P2_U3197 , P2_U3196 , P2_U3195 , P2_U3194;
output P2_U3193 , P2_U3192 , P2_U3191 , P2_U3190 , P2_U3189 , P2_U3188 , P2_U3187;
output P2_U3186 , P2_U3185 , P2_U3184 , P2_U3183 , P2_U3182 , P2_U3491 , P2_U3492;
output P2_U3493 , P2_U3494 , P2_U3495 , P2_U3496 , P2_U3497 , P2_U3498 , P2_U3499;
output P2_U3500 , P2_U3501 , P2_U3502 , P2_U3503 , P2_U3504 , P2_U3505 , P2_U3506;
output P2_U3507 , P2_U3508 , P2_U3509 , P2_U3510 , P2_U3511 , P2_U3512 , P2_U3513;
output P2_U3514 , P2_U3515 , P2_U3516 , P2_U3517 , P2_U3518 , P2_U3519 , P2_U3520;
output P2_U3521 , P2_U3522 , P2_U3296 , P2_U3181 , P2_U3180 , P2_U3179 , P2_U3178;
output P2_U3177 , P2_U3176 , P2_U3175 , P2_U3174 , P2_U3173 , P2_U3172 , P2_U3171;
output P2_U3170 , P2_U3169 , P2_U3168 , P2_U3167 , P2_U3166 , P2_U3165 , P2_U3164;
output P2_U3163 , P2_U3162 , P2_U3161 , P2_U3160 , P2_U3159 , P2_U3158 , P2_U3157;
output P2_U3156 , P2_U3155 , P2_U3154 , P2_U3153 , P2_U3151 , P2_U3150 , P2_U3893;

input SI_31_ , SI_30_ , SI_29_ , SI_28_ , SI_27_ , SI_26_;
input SI_25_ , SI_24_ , SI_23_ , SI_22_ , SI_21_ , SI_20_;
input SI_19_ , SI_18_ , SI_17_ , SI_16_ , SI_15_ , SI_14_;
input SI_13_ , SI_12_ , SI_11_ , SI_10_ , SI_9_ , SI_8_;
input SI_7_ , SI_6_ , SI_5_ , SI_4_ , SI_3_ , SI_2_;
input SI_1_ , SI_0_;
input P1_IR_REG_0_ , P1_IR_REG_1_ , P1_IR_REG_2_ , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_;
input P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_10_ , P1_IR_REG_11_;
input P1_IR_REG_12_ , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_;
input P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_20_ , P1_IR_REG_21_ , P1_IR_REG_22_ , P1_IR_REG_23_;
input P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ , P1_IR_REG_27_ , P1_IR_REG_28_ , P1_IR_REG_29_;
input P1_IR_REG_30_ , P1_IR_REG_31_ , P1_D_REG_0_ , P1_D_REG_1_ , P1_D_REG_2_ , P1_D_REG_3_;
input P1_D_REG_4_ , P1_D_REG_5_ , P1_D_REG_6_ , P1_D_REG_7_ , P1_D_REG_8_ , P1_D_REG_9_;
input P1_D_REG_10_ , P1_D_REG_11_ , P1_D_REG_12_ , P1_D_REG_13_ , P1_D_REG_14_ , P1_D_REG_15_;
input P1_D_REG_16_ , P1_D_REG_17_ , P1_D_REG_18_ , P1_D_REG_19_ , P1_D_REG_20_ , P1_D_REG_21_;
input P1_D_REG_22_ , P1_D_REG_23_ , P1_D_REG_24_ , P1_D_REG_25_ , P1_D_REG_26_ , P1_D_REG_27_;
input P1_D_REG_28_ , P1_D_REG_29_ , P1_D_REG_30_ , P1_D_REG_31_ , P1_REG0_REG_0_ , P1_REG0_REG_1_;
input P1_REG0_REG_2_ , P1_REG0_REG_3_ , P1_REG0_REG_4_ , P1_REG0_REG_5_ , P1_REG0_REG_6_ , P1_REG0_REG_7_;
input P1_REG0_REG_8_ , P1_REG0_REG_9_ , P1_REG0_REG_10_ , P1_REG0_REG_11_ , P1_REG0_REG_12_ , P1_REG0_REG_13_;
input P1_REG0_REG_14_ , P1_REG0_REG_15_ , P1_REG0_REG_16_ , P1_REG0_REG_17_ , P1_REG0_REG_18_ , P1_REG0_REG_19_;
input P1_REG0_REG_20_ , P1_REG0_REG_21_ , P1_REG0_REG_22_ , P1_REG0_REG_23_ , P1_REG0_REG_24_ , P1_REG0_REG_25_;
input P1_REG0_REG_26_ , P1_REG0_REG_27_ , P1_REG0_REG_28_ , P1_REG0_REG_29_ , P1_REG0_REG_30_ , P1_REG0_REG_31_;
input P1_REG1_REG_0_ , P1_REG1_REG_1_ , P1_REG1_REG_2_ , P1_REG1_REG_3_ , P1_REG1_REG_4_ , P1_REG1_REG_5_;
input P1_REG1_REG_6_ , P1_REG1_REG_7_ , P1_REG1_REG_8_ , P1_REG1_REG_9_ , P1_REG1_REG_10_ , P1_REG1_REG_11_;
input P1_REG1_REG_12_ , P1_REG1_REG_13_ , P1_REG1_REG_14_ , P1_REG1_REG_15_ , P1_REG1_REG_16_ , P1_REG1_REG_17_;
input P1_REG1_REG_18_ , P1_REG1_REG_19_ , P1_REG1_REG_20_ , P1_REG1_REG_21_ , P1_REG1_REG_22_ , P1_REG1_REG_23_;
input P1_REG1_REG_24_ , P1_REG1_REG_25_ , P1_REG1_REG_26_ , P1_REG1_REG_27_ , P1_REG1_REG_28_ , P1_REG1_REG_29_;
input P1_REG1_REG_30_ , P1_REG1_REG_31_ , P1_REG2_REG_0_ , P1_REG2_REG_1_ , P1_REG2_REG_2_ , P1_REG2_REG_3_;
input P1_REG2_REG_4_ , P1_REG2_REG_5_ , P1_REG2_REG_6_ , P1_REG2_REG_7_ , P1_REG2_REG_8_ , P1_REG2_REG_9_;
input P1_REG2_REG_10_ , P1_REG2_REG_11_ , P1_REG2_REG_12_ , P1_REG2_REG_13_ , P1_REG2_REG_14_ , P1_REG2_REG_15_;
input P1_REG2_REG_16_ , P1_REG2_REG_17_ , P1_REG2_REG_18_ , P1_REG2_REG_19_ , P1_REG2_REG_20_ , P1_REG2_REG_21_;
input P1_REG2_REG_22_ , P1_REG2_REG_23_ , P1_REG2_REG_24_ , P1_REG2_REG_25_ , P1_REG2_REG_26_ , P1_REG2_REG_27_;
input P1_REG2_REG_28_ , P1_REG2_REG_29_ , P1_REG2_REG_30_ , P1_REG2_REG_31_ , P1_ADDR_REG_19_ , P1_ADDR_REG_18_;
input P1_ADDR_REG_17_ , P1_ADDR_REG_16_ , P1_ADDR_REG_15_ , P1_ADDR_REG_14_ , P1_ADDR_REG_13_ , P1_ADDR_REG_12_;
input P1_ADDR_REG_11_ , P1_ADDR_REG_10_ , P1_ADDR_REG_9_ , P1_ADDR_REG_8_ , P1_ADDR_REG_7_ , P1_ADDR_REG_6_;
input P1_ADDR_REG_5_ , P1_ADDR_REG_4_ , P1_ADDR_REG_3_ , P1_ADDR_REG_2_ , P1_ADDR_REG_1_ , P1_ADDR_REG_0_;
input P1_DATAO_REG_0_ , P1_DATAO_REG_1_ , P1_DATAO_REG_2_ , P1_DATAO_REG_3_ , P1_DATAO_REG_4_ , P1_DATAO_REG_5_;
input P1_DATAO_REG_6_ , P1_DATAO_REG_7_ , P1_DATAO_REG_8_ , P1_DATAO_REG_9_ , P1_DATAO_REG_10_ , P1_DATAO_REG_11_;
input P1_DATAO_REG_12_ , P1_DATAO_REG_13_ , P1_DATAO_REG_14_ , P1_DATAO_REG_15_ , P1_DATAO_REG_16_ , P1_DATAO_REG_17_;
input P1_DATAO_REG_18_ , P1_DATAO_REG_19_ , P1_DATAO_REG_20_ , P1_DATAO_REG_21_ , P1_DATAO_REG_22_ , P1_DATAO_REG_23_;
input P1_DATAO_REG_24_ , P1_DATAO_REG_25_ , P1_DATAO_REG_26_ , P1_DATAO_REG_27_ , P1_DATAO_REG_28_ , P1_DATAO_REG_29_;
input P1_DATAO_REG_30_ , P1_DATAO_REG_31_ , P1_B_REG , P1_REG3_REG_15_ , P1_REG3_REG_26_ , P1_REG3_REG_6_;
input P1_REG3_REG_18_ , P1_REG3_REG_2_ , P1_REG3_REG_11_ , P1_REG3_REG_22_ , P1_REG3_REG_13_ , P1_REG3_REG_20_;
input P1_REG3_REG_0_ , P1_REG3_REG_9_ , P1_REG3_REG_4_ , P1_REG3_REG_24_ , P1_REG3_REG_17_ , P1_REG3_REG_5_;
input P1_REG3_REG_16_ , P1_REG3_REG_25_ , P1_REG3_REG_12_ , P1_REG3_REG_21_ , P1_REG3_REG_1_ , P1_REG3_REG_8_;
input P1_REG3_REG_28_ , P1_REG3_REG_19_ , P1_REG3_REG_3_ , P1_REG3_REG_10_ , P1_REG3_REG_23_ , P1_REG3_REG_14_;
input P1_REG3_REG_27_ , P1_REG3_REG_7_ , P1_STATE_REG , P1_RD_REG , P1_WR_REG , P2_IR_REG_0_;
input P2_IR_REG_1_ , P2_IR_REG_2_ , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ , P2_IR_REG_6_;
input P2_IR_REG_7_ , P2_IR_REG_8_ , P2_IR_REG_9_ , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_;
input P2_IR_REG_13_ , P2_IR_REG_14_ , P2_IR_REG_15_ , P2_IR_REG_16_ , P2_IR_REG_17_ , P2_IR_REG_18_;
input P2_IR_REG_19_ , P2_IR_REG_20_ , P2_IR_REG_21_ , P2_IR_REG_22_ , P2_IR_REG_23_ , P2_IR_REG_24_;
input P2_IR_REG_25_ , P2_IR_REG_26_ , P2_IR_REG_27_ , P2_IR_REG_28_ , P2_IR_REG_29_ , P2_IR_REG_30_;
input P2_IR_REG_31_ , P2_D_REG_0_ , P2_D_REG_1_ , P2_D_REG_2_ , P2_D_REG_3_ , P2_D_REG_4_;
input P2_D_REG_5_ , P2_D_REG_6_ , P2_D_REG_7_ , P2_D_REG_8_ , P2_D_REG_9_ , P2_D_REG_10_;
input P2_D_REG_11_ , P2_D_REG_12_ , P2_D_REG_13_ , P2_D_REG_14_ , P2_D_REG_15_ , P2_D_REG_16_;
input P2_D_REG_17_ , P2_D_REG_18_ , P2_D_REG_19_ , P2_D_REG_20_ , P2_D_REG_21_ , P2_D_REG_22_;
input P2_D_REG_23_ , P2_D_REG_24_ , P2_D_REG_25_ , P2_D_REG_26_ , P2_D_REG_27_ , P2_D_REG_28_;
input P2_D_REG_29_ , P2_D_REG_30_ , P2_D_REG_31_ , P2_REG0_REG_0_ , P2_REG0_REG_1_ , P2_REG0_REG_2_;
input P2_REG0_REG_3_ , P2_REG0_REG_4_ , P2_REG0_REG_5_ , P2_REG0_REG_6_ , P2_REG0_REG_7_ , P2_REG0_REG_8_;
input P2_REG0_REG_9_ , P2_REG0_REG_10_ , P2_REG0_REG_11_ , P2_REG0_REG_12_ , P2_REG0_REG_13_ , P2_REG0_REG_14_;
input P2_REG0_REG_15_ , P2_REG0_REG_16_ , P2_REG0_REG_17_ , P2_REG0_REG_18_ , P2_REG0_REG_19_ , P2_REG0_REG_20_;
input P2_REG0_REG_21_ , P2_REG0_REG_22_ , P2_REG0_REG_23_ , P2_REG0_REG_24_ , P2_REG0_REG_25_ , P2_REG0_REG_26_;
input P2_REG0_REG_27_ , P2_REG0_REG_28_ , P2_REG0_REG_29_ , P2_REG0_REG_30_ , P2_REG0_REG_31_ , P2_REG1_REG_0_;
input P2_REG1_REG_1_ , P2_REG1_REG_2_ , P2_REG1_REG_3_ , P2_REG1_REG_4_ , P2_REG1_REG_5_ , P2_REG1_REG_6_;
input P2_REG1_REG_7_ , P2_REG1_REG_8_ , P2_REG1_REG_9_ , P2_REG1_REG_10_ , P2_REG1_REG_11_ , P2_REG1_REG_12_;
input P2_REG1_REG_13_ , P2_REG1_REG_14_ , P2_REG1_REG_15_ , P2_REG1_REG_16_ , P2_REG1_REG_17_ , P2_REG1_REG_18_;
input P2_REG1_REG_19_ , P2_REG1_REG_20_ , P2_REG1_REG_21_ , P2_REG1_REG_22_ , P2_REG1_REG_23_ , P2_REG1_REG_24_;
input P2_REG1_REG_25_ , P2_REG1_REG_26_ , P2_REG1_REG_27_ , P2_REG1_REG_28_ , P2_REG1_REG_29_ , P2_REG1_REG_30_;
input P2_REG1_REG_31_ , P2_REG2_REG_0_ , P2_REG2_REG_1_ , P2_REG2_REG_2_ , P2_REG2_REG_3_ , P2_REG2_REG_4_;
input P2_REG2_REG_5_ , P2_REG2_REG_6_ , P2_REG2_REG_7_ , P2_REG2_REG_8_ , P2_REG2_REG_9_ , P2_REG2_REG_10_;
input P2_REG2_REG_11_ , P2_REG2_REG_12_ , P2_REG2_REG_13_ , P2_REG2_REG_14_ , P2_REG2_REG_15_ , P2_REG2_REG_16_;
input P2_REG2_REG_17_ , P2_REG2_REG_18_ , P2_REG2_REG_19_ , P2_REG2_REG_20_ , P2_REG2_REG_21_ , P2_REG2_REG_22_;
input P2_REG2_REG_23_ , P2_REG2_REG_24_ , P2_REG2_REG_25_ , P2_REG2_REG_26_ , P2_REG2_REG_27_ , P2_REG2_REG_28_;
input P2_REG2_REG_29_ , P2_REG2_REG_30_ , P2_REG2_REG_31_ , P2_ADDR_REG_19_ , P2_ADDR_REG_18_ , P2_ADDR_REG_17_;
input P2_ADDR_REG_16_ , P2_ADDR_REG_15_ , P2_ADDR_REG_14_ , P2_ADDR_REG_13_ , P2_ADDR_REG_12_ , P2_ADDR_REG_11_;
input P2_ADDR_REG_10_ , P2_ADDR_REG_9_ , P2_ADDR_REG_8_ , P2_ADDR_REG_7_ , P2_ADDR_REG_6_ , P2_ADDR_REG_5_;
input P2_ADDR_REG_4_ , P2_ADDR_REG_3_ , P2_ADDR_REG_2_ , P2_ADDR_REG_1_ , P2_ADDR_REG_0_ , P2_DATAO_REG_0_;
input P2_DATAO_REG_1_ , P2_DATAO_REG_2_ , P2_DATAO_REG_3_ , P2_DATAO_REG_4_ , P2_DATAO_REG_5_ , P2_DATAO_REG_6_;
input P2_DATAO_REG_7_ , P2_DATAO_REG_8_ , P2_DATAO_REG_9_ , P2_DATAO_REG_10_ , P2_DATAO_REG_11_ , P2_DATAO_REG_12_;
input P2_DATAO_REG_13_ , P2_DATAO_REG_14_ , P2_DATAO_REG_15_ , P2_DATAO_REG_16_ , P2_DATAO_REG_17_ , P2_DATAO_REG_18_;
input P2_DATAO_REG_19_ , P2_DATAO_REG_20_ , P2_DATAO_REG_21_ , P2_DATAO_REG_22_ , P2_DATAO_REG_23_ , P2_DATAO_REG_24_;
input P2_DATAO_REG_25_ , P2_DATAO_REG_26_ , P2_DATAO_REG_27_ , P2_DATAO_REG_28_ , P2_DATAO_REG_29_ , P2_DATAO_REG_30_;
input P2_DATAO_REG_31_ , P2_B_REG , P2_REG3_REG_15_ , P2_REG3_REG_26_ , P2_REG3_REG_6_ , P2_REG3_REG_18_;
input P2_REG3_REG_2_ , P2_REG3_REG_11_ , P2_REG3_REG_22_ , P2_REG3_REG_13_ , P2_REG3_REG_20_ , P2_REG3_REG_0_;
input P2_REG3_REG_9_ , P2_REG3_REG_4_ , P2_REG3_REG_24_ , P2_REG3_REG_17_ , P2_REG3_REG_5_ , P2_REG3_REG_16_;
input P2_REG3_REG_25_ , P2_REG3_REG_12_ , P2_REG3_REG_21_ , P2_REG3_REG_1_ , P2_REG3_REG_8_ , P2_REG3_REG_28_;
input P2_REG3_REG_19_ , P2_REG3_REG_3_ , P2_REG3_REG_10_ , P2_REG3_REG_23_ , P2_REG3_REG_14_ , P2_REG3_REG_27_;
input P2_REG3_REG_7_ , P2_STATE_REG , P2_RD_REG , P2_WR_REG;

wire P2_R1161_U504 , P2_R1161_U503 , P2_R1161_U502 , U25 , U26 , U27 , U28 , U29 , U30 , U31;
wire U32 , U33 , U34 , U35 , U36 , U37 , U38 , U39 , U40 , U41;
wire U42 , U43 , U44 , U45 , U46 , U47 , U48 , U49 , U50 , U51;
wire U52 , U53 , U54 , U55 , U56 , U57 , U58 , U59 , U60 , U61;
wire U62 , U63 , U64 , U65 , U66 , U67 , U68 , U69 , U70 , U71;
wire U72 , U73 , U74 , U75 , U76 , U77 , U78 , U79 , U80 , U81;
wire U82 , U83 , U84 , U85 , U86 , U87 , U88 , U89 , U90 , U91;
wire U92 , U93 , U94 , U95 , U96 , U97 , U98 , U99 , U100 , U101;
wire U102 , U103 , U104 , U105 , U106 , U107 , U108 , U109 , U110 , U111;
wire U112 , U113 , U114 , U115 , U116 , U117 , U118 , U119 , U120 , U121;
wire U122 , U124 , U125 , U127 , U128 , U129 , U130 , U131 , U132 , U133;
wire U134 , U135 , U136 , U137 , U138 , U139 , U140 , U141 , U142 , U143;
wire U144 , U145 , U146 , U147 , U148 , U149 , U150 , U151 , U152 , U153;
wire U154 , U155 , U156 , U157 , U158 , U159 , U160 , U161 , U162 , U163;
wire U164 , U165 , U166 , U167 , U168 , U169 , U170 , U171 , U172 , U173;
wire U174 , U175 , U176 , U177 , U178 , U179 , U180 , U181 , U182 , U183;
wire U184 , U185 , U186 , U187 , U188 , U189 , U190 , U191 , U192 , U193;
wire U194 , U195 , U196 , U197 , U198 , U199 , U200 , U201 , U202 , U203;
wire U204 , U205 , U206 , U207 , U208 , U209 , U210 , U211 , U212 , U213;
wire U214 , U215 , U216 , U217 , U218 , U219 , U220 , U221 , U222 , U223;
wire U224 , U225 , U226 , U227 , U228 , U229 , U230 , U231 , U232 , U233;
wire U234 , U235 , U236 , U237 , U238 , U239 , U240 , U241 , U242 , U243;
wire U244 , U245 , U246 , U247 , U248 , U249 , U250 , U251 , U252 , U253;
wire U254 , U255 , U256 , U257 , U258 , U259 , U260 , U261 , U262 , U263;
wire U264 , U265 , U266 , U267 , U268 , U269 , U270 , U271 , U272 , U273;
wire U274 , U275 , U276 , U277 , U278 , U279 , U280 , U281 , U282 , U283;
wire U284 , U285 , U286 , U287 , U288 , U289 , U290 , U291 , U292 , U293;
wire U294 , U295 , U296 , U297 , U298 , U299 , U300 , U301 , U302 , U303;
wire U304 , U305 , U306 , U307 , U308 , U309 , U310 , U311 , U312 , U313;
wire U314 , U315 , U316 , U317 , U318 , U319 , U320 , U321 , U322 , U323;
wire U324 , U325 , U326 , P2_R1161_U501 , P2_R1161_U500 , P2_R1161_U499 , P2_R1161_U498 , P2_R1161_U497 , P2_R1161_U496 , P2_R1161_U495;
wire P2_R1161_U494 , P2_R1161_U493 , P2_R1161_U492 , P2_R1161_U491 , P2_R1161_U490 , P1_U3014 , P1_U3015 , P1_U3016 , P1_U3017 , P1_U3018;
wire P1_U3019 , P1_U3020 , P1_U3021 , P1_U3022 , P1_U3023 , P1_U3024 , P1_U3025 , P1_U3026 , P1_U3027 , P1_U3028;
wire P1_U3029 , P1_U3030 , P1_U3031 , P1_U3032 , P1_U3033 , P1_U3034 , P1_U3035 , P1_U3036 , P1_U3037 , P1_U3038;
wire P1_U3039 , P1_U3040 , P1_U3041 , P1_U3042 , P1_U3043 , P1_U3044 , P1_U3045 , P1_U3046 , P1_U3047 , P1_U3048;
wire P1_U3049 , P1_U3050 , P1_U3051 , P1_U3052 , P1_U3053 , P1_U3054 , P1_U3055 , P1_U3056 , P1_U3057 , P1_U3058;
wire P1_U3059 , P1_U3060 , P1_U3061 , P1_U3062 , P1_U3063 , P1_U3064 , P1_U3065 , P1_U3066 , P1_U3067 , P1_U3068;
wire P1_U3069 , P1_U3070 , P1_U3071 , P1_U3072 , P1_U3073 , P1_U3074 , P1_U3075 , P1_U3076 , P1_U3077 , P1_U3078;
wire P1_U3079 , P1_U3080 , P1_U3081 , P1_U3082 , P1_U3083 , P1_U3084 , P1_U3087 , P1_U3088 , P1_U3089 , P1_U3090;
wire P1_U3091 , P1_U3092 , P1_U3093 , P1_U3094 , P1_U3095 , P1_U3096 , P1_U3097 , P1_U3098 , P1_U3099 , P1_U3100;
wire P1_U3101 , P1_U3102 , P1_U3103 , P1_U3104 , P1_U3105 , P1_U3106 , P1_U3107 , P1_U3108 , P1_U3109 , P1_U3110;
wire P1_U3111 , P1_U3112 , P1_U3113 , P1_U3114 , P1_U3115 , P1_U3116 , P1_U3117 , P1_U3118 , P1_U3119 , P1_U3120;
wire P1_U3121 , P1_U3122 , P1_U3123 , P1_U3124 , P1_U3125 , P1_U3126 , P1_U3127 , P1_U3128 , P1_U3129 , P1_U3130;
wire P1_U3131 , P1_U3132 , P1_U3133 , P1_U3134 , P1_U3135 , P1_U3136 , P1_U3137 , P1_U3138 , P1_U3139 , P1_U3140;
wire P1_U3141 , P1_U3142 , P1_U3143 , P1_U3144 , P1_U3145 , P1_U3146 , P1_U3147 , P1_U3148 , P1_U3149 , P1_U3150;
wire P1_U3151 , P1_U3152 , P1_U3153 , P1_U3154 , P1_U3155 , P1_U3156 , P1_U3157 , P1_U3158 , P1_U3159 , P1_U3160;
wire P1_U3161 , P1_U3162 , P1_U3163 , P1_U3164 , P1_U3165 , P1_U3166 , P1_U3167 , P1_U3168 , P1_U3169 , P1_U3170;
wire P1_U3171 , P1_U3172 , P1_U3173 , P1_U3174 , P1_U3175 , P1_U3176 , P1_U3177 , P1_U3178 , P1_U3179 , P1_U3180;
wire P1_U3181 , P1_U3182 , P1_U3183 , P1_U3184 , P1_U3185 , P1_U3186 , P1_U3187 , P1_U3188 , P1_U3189 , P1_U3190;
wire P1_U3191 , P1_U3192 , P1_U3193 , P1_U3194 , P1_U3195 , P1_U3196 , P1_U3197 , P1_U3198 , P1_U3199 , P1_U3200;
wire P1_U3201 , P1_U3202 , P1_U3203 , P1_U3204 , P1_U3205 , P1_U3206 , P1_U3207 , P1_U3208 , P1_U3209 , P1_U3210;
wire P1_U3211 , P1_U3212 , P1_U3357 , P1_U3358 , P1_U3359 , P1_U3360 , P1_U3361 , P1_U3362 , P1_U3363 , P1_U3364;
wire P1_U3365 , P1_U3366 , P1_U3367 , P1_U3368 , P1_U3369 , P1_U3370 , P1_U3371 , P1_U3372 , P1_U3373 , P1_U3374;
wire P1_U3375 , P1_U3376 , P1_U3377 , P1_U3378 , P1_U3379 , P1_U3380 , P1_U3381 , P1_U3382 , P1_U3383 , P1_U3384;
wire P1_U3385 , P1_U3386 , P1_U3387 , P1_U3388 , P1_U3389 , P1_U3390 , P1_U3391 , P1_U3392 , P1_U3393 , P1_U3394;
wire P1_U3395 , P1_U3396 , P1_U3397 , P1_U3398 , P1_U3399 , P1_U3400 , P1_U3401 , P1_U3402 , P1_U3403 , P1_U3404;
wire P1_U3405 , P1_U3406 , P1_U3407 , P1_U3408 , P1_U3409 , P1_U3410 , P1_U3411 , P1_U3412 , P1_U3413 , P1_U3414;
wire P1_U3415 , P1_U3416 , P1_U3417 , P1_U3418 , P1_U3419 , P1_U3420 , P1_U3421 , P1_U3422 , P1_U3423 , P1_U3424;
wire P1_U3425 , P1_U3426 , P1_U3427 , P1_U3428 , P1_U3429 , P1_U3430 , P1_U3431 , P1_U3432 , P1_U3433 , P1_U3434;
wire P1_U3435 , P1_U3436 , P1_U3437 , P1_U3438 , P1_U3441 , P1_U3442 , P1_U3443 , P1_U3444 , P1_U3445 , P1_U3446;
wire P1_U3447 , P1_U3448 , P1_U3449 , P1_U3450 , P1_U3451 , P1_U3452 , P1_U3454 , P1_U3455 , P1_U3457 , P1_U3458;
wire P1_U3460 , P1_U3461 , P1_U3463 , P1_U3464 , P1_U3466 , P1_U3467 , P1_U3469 , P1_U3470 , P1_U3472 , P1_U3473;
wire P1_U3475 , P1_U3476 , P1_U3478 , P1_U3479 , P1_U3481 , P1_U3482 , P1_U3484 , P1_U3485 , P1_U3487 , P1_U3488;
wire P1_U3490 , P1_U3491 , P1_U3493 , P1_U3494 , P1_U3496 , P1_U3497 , P1_U3499 , P1_U3500 , P1_U3502 , P1_U3503;
wire P1_U3505 , P1_U3506 , P1_U3508 , P1_U3586 , P1_U3587 , P1_U3588 , P1_U3589 , P1_U3590 , P1_U3591 , P1_U3592;
wire P1_U3593 , P1_U3594 , P1_U3595 , P1_U3596 , P1_U3597 , P1_U3598 , P1_U3599 , P1_U3600 , P1_U3601 , P1_U3602;
wire P1_U3603 , P1_U3604 , P1_U3605 , P1_U3606 , P1_U3607 , P1_U3608 , P1_U3609 , P1_U3610 , P1_U3611 , P1_U3612;
wire P1_U3613 , P1_U3614 , P1_U3615 , P1_U3616 , P1_U3617 , P1_U3618 , P1_U3619 , P1_U3620 , P1_U3621 , P1_U3622;
wire P1_U3623 , P1_U3624 , P1_U3625 , P1_U3626 , P1_U3627 , P1_U3628 , P1_U3629 , P1_U3630 , P1_U3631 , P1_U3632;
wire P1_U3633 , P1_U3634 , P1_U3635 , P1_U3636 , P1_U3637 , P1_U3638 , P1_U3639 , P1_U3640 , P1_U3641 , P1_U3642;
wire P1_U3643 , P1_U3644 , P1_U3645 , P1_U3646 , P1_U3647 , P1_U3648 , P1_U3649 , P1_U3650 , P1_U3651 , P1_U3652;
wire P1_U3653 , P1_U3654 , P1_U3655 , P1_U3656 , P1_U3657 , P1_U3658 , P1_U3659 , P1_U3660 , P1_U3661 , P1_U3662;
wire P1_U3663 , P1_U3664 , P1_U3665 , P1_U3666 , P1_U3667 , P1_U3668 , P1_U3669 , P1_U3670 , P1_U3671 , P1_U3672;
wire P1_U3673 , P1_U3674 , P1_U3675 , P1_U3676 , P1_U3677 , P1_U3678 , P1_U3679 , P1_U3680 , P1_U3681 , P1_U3682;
wire P1_U3683 , P1_U3684 , P1_U3685 , P1_U3686 , P1_U3687 , P1_U3688 , P1_U3689 , P1_U3690 , P1_U3691 , P1_U3692;
wire P1_U3693 , P1_U3694 , P1_U3695 , P1_U3696 , P1_U3697 , P1_U3698 , P1_U3699 , P1_U3700 , P1_U3701 , P1_U3702;
wire P1_U3703 , P1_U3704 , P1_U3705 , P1_U3706 , P1_U3707 , P1_U3708 , P1_U3709 , P1_U3710 , P1_U3711 , P1_U3712;
wire P1_U3713 , P1_U3714 , P1_U3715 , P1_U3716 , P1_U3717 , P1_U3718 , P1_U3719 , P1_U3720 , P1_U3721 , P1_U3722;
wire P1_U3723 , P1_U3724 , P1_U3725 , P1_U3726 , P1_U3727 , P1_U3728 , P1_U3729 , P1_U3730 , P1_U3731 , P1_U3732;
wire P1_U3733 , P1_U3734 , P1_U3735 , P1_U3736 , P1_U3737 , P1_U3738 , P1_U3739 , P1_U3740 , P1_U3741 , P1_U3742;
wire P1_U3743 , P1_U3744 , P1_U3745 , P1_U3746 , P1_U3747 , P1_U3748 , P1_U3749 , P1_U3750 , P1_U3751 , P1_U3752;
wire P1_U3753 , P1_U3754 , P1_U3755 , P1_U3756 , P1_U3757 , P1_U3758 , P1_U3759 , P1_U3760 , P1_U3761 , P1_U3762;
wire P1_U3763 , P1_U3764 , P1_U3765 , P1_U3766 , P1_U3767 , P1_U3768 , P1_U3769 , P1_U3770 , P1_U3771 , P1_U3772;
wire P1_U3773 , P1_U3774 , P1_U3775 , P1_U3776 , P1_U3777 , P1_U3778 , P1_U3779 , P1_U3780 , P1_U3781 , P1_U3782;
wire P1_U3783 , P1_U3784 , P1_U3785 , P1_U3786 , P1_U3787 , P1_U3788 , P1_U3789 , P1_U3790 , P1_U3791 , P1_U3792;
wire P1_U3793 , P1_U3794 , P1_U3795 , P1_U3796 , P1_U3797 , P1_U3798 , P1_U3799 , P1_U3800 , P1_U3801 , P1_U3802;
wire P1_U3803 , P1_U3804 , P1_U3805 , P1_U3806 , P1_U3807 , P1_U3808 , P1_U3809 , P1_U3810 , P1_U3811 , P1_U3812;
wire P1_U3813 , P1_U3814 , P1_U3815 , P1_U3816 , P1_U3817 , P1_U3818 , P1_U3819 , P1_U3820 , P1_U3821 , P1_U3822;
wire P1_U3823 , P1_U3824 , P1_U3825 , P1_U3826 , P1_U3827 , P1_U3828 , P1_U3829 , P1_U3830 , P1_U3831 , P1_U3832;
wire P1_U3833 , P1_U3834 , P1_U3835 , P1_U3836 , P1_U3837 , P1_U3838 , P1_U3839 , P1_U3840 , P1_U3841 , P1_U3842;
wire P1_U3843 , P1_U3844 , P1_U3845 , P1_U3846 , P1_U3847 , P1_U3848 , P1_U3849 , P1_U3850 , P1_U3851 , P1_U3852;
wire P1_U3853 , P1_U3854 , P1_U3855 , P1_U3856 , P1_U3857 , P1_U3858 , P1_U3859 , P1_U3860 , P1_U3861 , P1_U3862;
wire P1_U3863 , P1_U3864 , P1_U3865 , P1_U3866 , P1_U3867 , P1_U3868 , P1_U3869 , P1_U3870 , P1_U3871 , P1_U3872;
wire P1_U3873 , P1_U3874 , P1_U3875 , P1_U3876 , P1_U3877 , P1_U3878 , P1_U3879 , P1_U3880 , P1_U3881 , P1_U3882;
wire P1_U3883 , P1_U3884 , P1_U3885 , P1_U3886 , P1_U3887 , P1_U3888 , P1_U3889 , P1_U3890 , P1_U3891 , P1_U3892;
wire P1_U3893 , P1_U3894 , P1_U3895 , P1_U3896 , P1_U3897 , P1_U3898 , P1_U3899 , P1_U3900 , P1_U3901 , P1_U3902;
wire P1_U3903 , P1_U3904 , P1_U3905 , P1_U3906 , P1_U3907 , P1_U3908 , P1_U3909 , P1_U3910 , P1_U3911 , P1_U3912;
wire P1_U3913 , P1_U3914 , P1_U3915 , P1_U3916 , P1_U3917 , P1_U3918 , P1_U3919 , P1_U3920 , P1_U3921 , P1_U3922;
wire P1_U3923 , P1_U3924 , P1_U3925 , P1_U3926 , P1_U3927 , P1_U3928 , P1_U3929 , P1_U3930 , P1_U3931 , P1_U3932;
wire P1_U3933 , P1_U3934 , P1_U3935 , P1_U3936 , P1_U3937 , P1_U3938 , P1_U3939 , P1_U3940 , P1_U3941 , P1_U3942;
wire P1_U3943 , P1_U3944 , P1_U3945 , P1_U3946 , P1_U3947 , P1_U3948 , P1_U3949 , P1_U3950 , P1_U3951 , P1_U3952;
wire P1_U3953 , P1_U3954 , P1_U3955 , P1_U3956 , P1_U3957 , P1_U3958 , P1_U3959 , P1_U3960 , P1_U3961 , P1_U3962;
wire P1_U3963 , P1_U3964 , P1_U3965 , P1_U3966 , P1_U3967 , P1_U3968 , P1_U3969 , P1_U3970 , P1_U3971 , P1_U3972;
wire P1_U3974 , P1_U3975 , P1_U3976 , P1_U3977 , P1_U3978 , P1_U3979 , P1_U3980 , P1_U3981 , P1_U3982 , P1_U3983;
wire P1_U3984 , P1_U3985 , P1_U3986 , P1_U3987 , P1_U3988 , P1_U3989 , P1_U3990 , P1_U3991 , P1_U3992 , P1_U3993;
wire P1_U3994 , P1_U3995 , P1_U3996 , P1_U3997 , P1_U3998 , P1_U3999 , P1_U4000 , P1_U4001 , P1_U4002 , P1_U4003;
wire P1_U4004 , P1_U4005 , P1_U4006 , P1_U4007 , P1_U4008 , P1_U4009 , P1_U4010 , P1_U4011 , P1_U4012 , P1_U4013;
wire P1_U4014 , P1_U4015 , P1_U4016 , P1_U4017 , P1_U4018 , P1_U4019 , P1_U4020 , P1_U4021 , P1_U4022 , P1_U4023;
wire P1_U4024 , P1_U4025 , P1_U4026 , P1_U4027 , P1_U4028 , P1_U4029 , P1_U4030 , P1_U4031 , P1_U4032 , P1_U4033;
wire P1_U4034 , P1_U4035 , P1_U4036 , P1_U4037 , P1_U4038 , P1_U4039 , P1_U4040 , P1_U4041 , P1_U4042 , P1_U4043;
wire P1_U4044 , P1_U4045 , P1_U4046 , P1_U4047 , P1_U4048 , P1_U4049 , P1_U4050 , P1_U4051 , P1_U4052 , P1_U4053;
wire P1_U4054 , P1_U4055 , P1_U4056 , P1_U4057 , P1_U4058 , P1_U4059 , P1_U4060 , P1_U4061 , P1_U4062 , P1_U4063;
wire P1_U4064 , P1_U4065 , P1_U4066 , P1_U4067 , P1_U4068 , P1_U4069 , P1_U4070 , P1_U4071 , P1_U4072 , P1_U4073;
wire P1_U4074 , P1_U4075 , P1_U4076 , P1_U4077 , P1_U4078 , P1_U4079 , P1_U4080 , P1_U4081 , P1_U4082 , P1_U4083;
wire P1_U4084 , P1_U4085 , P1_U4086 , P1_U4087 , P1_U4088 , P1_U4089 , P1_U4090 , P1_U4091 , P1_U4092 , P1_U4093;
wire P1_U4094 , P1_U4095 , P1_U4096 , P1_U4097 , P1_U4098 , P1_U4099 , P1_U4100 , P1_U4101 , P1_U4102 , P1_U4103;
wire P1_U4104 , P1_U4105 , P1_U4106 , P1_U4107 , P1_U4108 , P1_U4109 , P1_U4110 , P1_U4111 , P1_U4112 , P1_U4113;
wire P1_U4114 , P1_U4115 , P1_U4116 , P1_U4117 , P1_U4118 , P1_U4119 , P1_U4120 , P1_U4121 , P1_U4122 , P1_U4123;
wire P1_U4124 , P1_U4125 , P1_U4126 , P1_U4127 , P1_U4128 , P1_U4129 , P1_U4130 , P1_U4131 , P1_U4132 , P1_U4133;
wire P1_U4134 , P1_U4135 , P1_U4136 , P1_U4137 , P1_U4138 , P1_U4139 , P1_U4140 , P1_U4141 , P1_U4142 , P1_U4143;
wire P1_U4144 , P1_U4145 , P1_U4146 , P1_U4147 , P1_U4148 , P1_U4149 , P1_U4150 , P1_U4151 , P1_U4152 , P1_U4153;
wire P1_U4154 , P1_U4155 , P1_U4156 , P1_U4157 , P1_U4158 , P1_U4159 , P1_U4160 , P1_U4161 , P1_U4162 , P1_U4163;
wire P1_U4164 , P1_U4165 , P1_U4166 , P1_U4167 , P1_U4168 , P1_U4169 , P1_U4170 , P1_U4171 , P1_U4172 , P1_U4173;
wire P1_U4174 , P1_U4175 , P1_U4176 , P1_U4177 , P1_U4178 , P1_U4179 , P1_U4180 , P1_U4181 , P1_U4182 , P1_U4183;
wire P1_U4184 , P1_U4185 , P1_U4186 , P1_U4187 , P1_U4188 , P1_U4189 , P1_U4190 , P1_U4191 , P1_U4192 , P1_U4193;
wire P1_U4194 , P1_U4195 , P1_U4196 , P1_U4197 , P1_U4198 , P1_U4199 , P1_U4200 , P1_U4201 , P1_U4202 , P1_U4203;
wire P1_U4204 , P1_U4205 , P1_U4206 , P1_U4207 , P1_U4208 , P1_U4209 , P1_U4210 , P1_U4211 , P1_U4212 , P1_U4213;
wire P1_U4214 , P1_U4215 , P1_U4216 , P1_U4217 , P1_U4218 , P1_U4219 , P1_U4220 , P1_U4221 , P1_U4222 , P1_U4223;
wire P1_U4224 , P1_U4225 , P1_U4226 , P1_U4227 , P1_U4228 , P1_U4229 , P1_U4230 , P1_U4231 , P1_U4232 , P1_U4233;
wire P1_U4234 , P1_U4235 , P1_U4236 , P1_U4237 , P1_U4238 , P1_U4239 , P1_U4240 , P1_U4241 , P1_U4242 , P1_U4243;
wire P1_U4244 , P1_U4245 , P1_U4246 , P1_U4247 , P1_U4248 , P1_U4249 , P1_U4250 , P1_U4251 , P1_U4252 , P1_U4253;
wire P1_U4254 , P1_U4255 , P1_U4256 , P1_U4257 , P1_U4258 , P1_U4259 , P1_U4260 , P1_U4261 , P1_U4262 , P1_U4263;
wire P1_U4264 , P1_U4265 , P1_U4266 , P1_U4267 , P1_U4268 , P1_U4269 , P1_U4270 , P1_U4271 , P1_U4272 , P1_U4273;
wire P1_U4274 , P1_U4275 , P1_U4276 , P1_U4277 , P1_U4278 , P1_U4279 , P1_U4280 , P1_U4281 , P1_U4282 , P1_U4283;
wire P1_U4284 , P1_U4285 , P1_U4286 , P1_U4287 , P1_U4288 , P1_U4289 , P1_U4290 , P1_U4291 , P1_U4292 , P1_U4293;
wire P1_U4294 , P1_U4295 , P1_U4296 , P1_U4297 , P1_U4298 , P1_U4299 , P1_U4300 , P1_U4301 , P1_U4302 , P1_U4303;
wire P1_U4304 , P1_U4305 , P1_U4306 , P1_U4307 , P1_U4308 , P1_U4309 , P1_U4310 , P1_U4311 , P1_U4312 , P1_U4313;
wire P1_U4314 , P1_U4315 , P1_U4316 , P1_U4317 , P1_U4318 , P1_U4319 , P1_U4320 , P1_U4321 , P1_U4322 , P1_U4323;
wire P1_U4324 , P1_U4325 , P1_U4326 , P1_U4327 , P1_U4328 , P1_U4329 , P1_U4330 , P1_U4331 , P1_U4332 , P1_U4333;
wire P1_U4334 , P1_U4335 , P1_U4336 , P1_U4337 , P1_U4338 , P1_U4339 , P1_U4340 , P1_U4341 , P1_U4342 , P1_U4343;
wire P1_U4344 , P1_U4345 , P1_U4346 , P1_U4347 , P1_U4348 , P1_U4349 , P1_U4350 , P1_U4351 , P1_U4352 , P1_U4353;
wire P1_U4354 , P1_U4355 , P1_U4356 , P1_U4357 , P1_U4358 , P1_U4359 , P1_U4360 , P1_U4361 , P1_U4362 , P1_U4363;
wire P1_U4364 , P1_U4365 , P1_U4366 , P1_U4367 , P1_U4368 , P1_U4369 , P1_U4370 , P1_U4371 , P1_U4372 , P1_U4373;
wire P1_U4374 , P1_U4375 , P1_U4376 , P1_U4377 , P1_U4378 , P1_U4379 , P1_U4380 , P1_U4381 , P1_U4382 , P1_U4383;
wire P1_U4384 , P1_U4385 , P1_U4386 , P1_U4387 , P1_U4388 , P1_U4389 , P1_U4390 , P1_U4391 , P1_U4392 , P1_U4393;
wire P1_U4394 , P1_U4395 , P1_U4396 , P1_U4397 , P1_U4398 , P1_U4399 , P1_U4400 , P1_U4401 , P1_U4402 , P1_U4403;
wire P1_U4404 , P1_U4405 , P1_U4406 , P1_U4407 , P1_U4408 , P1_U4409 , P1_U4410 , P1_U4411 , P1_U4412 , P1_U4413;
wire P1_U4414 , P1_U4415 , P1_U4416 , P1_U4417 , P1_U4418 , P1_U4419 , P1_U4420 , P1_U4421 , P1_U4422 , P1_U4423;
wire P1_U4424 , P1_U4425 , P1_U4426 , P1_U4427 , P1_U4428 , P1_U4429 , P1_U4430 , P1_U4431 , P1_U4432 , P1_U4433;
wire P1_U4434 , P1_U4435 , P1_U4436 , P1_U4437 , P1_U4438 , P1_U4439 , P1_U4440 , P1_U4441 , P1_U4442 , P1_U4443;
wire P1_U4444 , P1_U4445 , P1_U4446 , P1_U4447 , P1_U4448 , P1_U4449 , P1_U4450 , P1_U4451 , P1_U4452 , P1_U4453;
wire P1_U4454 , P1_U4455 , P1_U4456 , P1_U4457 , P1_U4458 , P1_U4459 , P1_U4460 , P1_U4461 , P1_U4462 , P1_U4463;
wire P1_U4464 , P1_U4465 , P1_U4466 , P1_U4467 , P1_U4468 , P1_U4469 , P1_U4470 , P1_U4471 , P1_U4472 , P1_U4473;
wire P1_U4474 , P1_U4475 , P1_U4476 , P1_U4477 , P1_U4478 , P1_U4479 , P1_U4480 , P1_U4481 , P1_U4482 , P1_U4483;
wire P1_U4484 , P1_U4485 , P1_U4486 , P1_U4487 , P1_U4488 , P1_U4489 , P1_U4490 , P1_U4491 , P1_U4492 , P1_U4493;
wire P1_U4494 , P1_U4495 , P1_U4496 , P1_U4497 , P1_U4498 , P1_U4499 , P1_U4500 , P1_U4501 , P1_U4502 , P1_U4503;
wire P1_U4504 , P1_U4505 , P1_U4506 , P1_U4507 , P1_U4508 , P1_U4509 , P1_U4510 , P1_U4511 , P1_U4512 , P1_U4513;
wire P1_U4514 , P1_U4515 , P1_U4516 , P1_U4517 , P1_U4518 , P1_U4519 , P1_U4520 , P1_U4521 , P1_U4522 , P1_U4523;
wire P1_U4524 , P1_U4525 , P1_U4526 , P1_U4527 , P1_U4528 , P1_U4529 , P1_U4530 , P1_U4531 , P1_U4532 , P1_U4533;
wire P1_U4534 , P1_U4535 , P1_U4536 , P1_U4537 , P1_U4538 , P1_U4539 , P1_U4540 , P1_U4541 , P1_U4542 , P1_U4543;
wire P1_U4544 , P1_U4545 , P1_U4546 , P1_U4547 , P1_U4548 , P1_U4549 , P1_U4550 , P1_U4551 , P1_U4552 , P1_U4553;
wire P1_U4554 , P1_U4555 , P1_U4556 , P1_U4557 , P1_U4558 , P1_U4559 , P1_U4560 , P1_U4561 , P1_U4562 , P1_U4563;
wire P1_U4564 , P1_U4565 , P1_U4566 , P1_U4567 , P1_U4568 , P1_U4569 , P1_U4570 , P1_U4571 , P1_U4572 , P1_U4573;
wire P1_U4574 , P1_U4575 , P1_U4576 , P1_U4577 , P1_U4578 , P1_U4579 , P1_U4580 , P1_U4581 , P1_U4582 , P1_U4583;
wire P1_U4584 , P1_U4585 , P1_U4586 , P1_U4587 , P1_U4588 , P1_U4589 , P1_U4590 , P1_U4591 , P1_U4592 , P1_U4593;
wire P1_U4594 , P1_U4595 , P1_U4596 , P1_U4597 , P1_U4598 , P1_U4599 , P1_U4600 , P1_U4601 , P1_U4602 , P1_U4603;
wire P1_U4604 , P1_U4605 , P1_U4606 , P1_U4607 , P1_U4608 , P1_U4609 , P1_U4610 , P1_U4611 , P1_U4612 , P1_U4613;
wire P1_U4614 , P1_U4615 , P1_U4616 , P1_U4617 , P1_U4618 , P1_U4619 , P1_U4620 , P1_U4621 , P1_U4622 , P1_U4623;
wire P1_U4624 , P1_U4625 , P1_U4626 , P1_U4627 , P1_U4628 , P1_U4629 , P1_U4630 , P1_U4631 , P1_U4632 , P1_U4633;
wire P1_U4634 , P1_U4635 , P1_U4636 , P1_U4637 , P1_U4638 , P1_U4639 , P1_U4640 , P1_U4641 , P1_U4642 , P1_U4643;
wire P1_U4644 , P1_U4645 , P1_U4646 , P1_U4647 , P1_U4648 , P1_U4649 , P1_U4650 , P1_U4651 , P1_U4652 , P1_U4653;
wire P1_U4654 , P1_U4655 , P1_U4656 , P1_U4657 , P1_U4658 , P1_U4659 , P1_U4660 , P1_U4661 , P1_U4662 , P1_U4663;
wire P1_U4664 , P1_U4665 , P1_U4666 , P1_U4667 , P1_U4668 , P1_U4669 , P1_U4670 , P1_U4671 , P1_U4672 , P1_U4673;
wire P1_U4674 , P1_U4675 , P1_U4676 , P1_U4677 , P1_U4678 , P1_U4679 , P1_U4680 , P1_U4681 , P1_U4682 , P1_U4683;
wire P1_U4684 , P1_U4685 , P1_U4686 , P1_U4687 , P1_U4688 , P1_U4689 , P1_U4690 , P1_U4691 , P1_U4692 , P1_U4693;
wire P1_U4694 , P1_U4695 , P1_U4696 , P1_U4697 , P1_U4698 , P1_U4699 , P1_U4700 , P1_U4701 , P1_U4702 , P1_U4703;
wire P1_U4704 , P1_U4705 , P1_U4706 , P1_U4707 , P1_U4708 , P1_U4709 , P1_U4710 , P1_U4711 , P1_U4712 , P1_U4713;
wire P1_U4714 , P1_U4715 , P1_U4716 , P1_U4717 , P1_U4718 , P1_U4719 , P1_U4720 , P1_U4721 , P1_U4722 , P1_U4723;
wire P1_U4724 , P1_U4725 , P1_U4726 , P1_U4727 , P1_U4728 , P1_U4729 , P1_U4730 , P1_U4731 , P1_U4732 , P1_U4733;
wire P1_U4734 , P1_U4735 , P1_U4736 , P1_U4737 , P1_U4738 , P1_U4739 , P1_U4740 , P1_U4741 , P1_U4742 , P1_U4743;
wire P1_U4744 , P1_U4745 , P1_U4746 , P1_U4747 , P1_U4748 , P1_U4749 , P1_U4750 , P1_U4751 , P1_U4752 , P1_U4753;
wire P1_U4754 , P1_U4755 , P1_U4756 , P1_U4757 , P1_U4758 , P1_U4759 , P1_U4760 , P1_U4761 , P1_U4762 , P1_U4763;
wire P1_U4764 , P1_U4765 , P1_U4766 , P1_U4767 , P1_U4768 , P1_U4769 , P1_U4770 , P1_U4771 , P1_U4772 , P1_U4773;
wire P1_U4774 , P1_U4775 , P1_U4776 , P1_U4777 , P1_U4778 , P1_U4779 , P1_U4780 , P1_U4781 , P1_U4782 , P1_U4783;
wire P1_U4784 , P1_U4785 , P1_U4786 , P1_U4787 , P1_U4788 , P1_U4789 , P1_U4790 , P1_U4791 , P1_U4792 , P1_U4793;
wire P1_U4794 , P1_U4795 , P1_U4796 , P1_U4797 , P1_U4798 , P1_U4799 , P1_U4800 , P1_U4801 , P1_U4802 , P1_U4803;
wire P1_U4804 , P1_U4805 , P1_U4806 , P1_U4807 , P1_U4808 , P1_U4809 , P1_U4810 , P1_U4811 , P1_U4812 , P1_U4813;
wire P1_U4814 , P1_U4815 , P1_U4816 , P1_U4817 , P1_U4818 , P1_U4819 , P1_U4820 , P1_U4821 , P1_U4822 , P1_U4823;
wire P1_U4824 , P1_U4825 , P1_U4826 , P1_U4827 , P1_U4828 , P1_U4829 , P1_U4830 , P1_U4831 , P1_U4832 , P1_U4833;
wire P1_U4834 , P1_U4835 , P1_U4836 , P1_U4837 , P1_U4838 , P1_U4839 , P1_U4840 , P1_U4841 , P1_U4842 , P1_U4843;
wire P1_U4844 , P1_U4845 , P1_U4846 , P1_U4847 , P1_U4848 , P1_U4849 , P1_U4850 , P1_U4851 , P1_U4852 , P1_U4853;
wire P1_U4854 , P1_U4855 , P1_U4856 , P1_U4857 , P1_U4858 , P1_U4859 , P1_U4860 , P1_U4861 , P1_U4862 , P1_U4863;
wire P1_U4864 , P1_U4865 , P1_U4866 , P1_U4867 , P1_U4868 , P1_U4869 , P1_U4870 , P1_U4871 , P1_U4872 , P1_U4873;
wire P1_U4874 , P1_U4875 , P1_U4876 , P1_U4877 , P1_U4878 , P1_U4879 , P1_U4880 , P1_U4881 , P1_U4882 , P1_U4883;
wire P1_U4884 , P1_U4885 , P1_U4886 , P1_U4887 , P1_U4888 , P1_U4889 , P1_U4890 , P1_U4891 , P1_U4892 , P1_U4893;
wire P1_U4894 , P1_U4895 , P1_U4896 , P1_U4897 , P1_U4898 , P1_U4899 , P1_U4900 , P1_U4901 , P1_U4902 , P1_U4903;
wire P1_U4904 , P1_U4905 , P1_U4906 , P1_U4907 , P1_U4908 , P1_U4909 , P1_U4910 , P1_U4911 , P1_U4912 , P1_U4913;
wire P1_U4914 , P1_U4915 , P1_U4916 , P1_U4917 , P1_U4918 , P1_U4919 , P1_U4920 , P1_U4921 , P1_U4922 , P1_U4923;
wire P1_U4924 , P1_U4925 , P1_U4926 , P1_U4927 , P1_U4928 , P1_U4929 , P1_U4930 , P1_U4931 , P1_U4932 , P1_U4933;
wire P1_U4934 , P1_U4935 , P1_U4936 , P1_U4937 , P1_U4938 , P1_U4939 , P1_U4940 , P1_U4941 , P1_U4942 , P1_U4943;
wire P1_U4944 , P1_U4945 , P1_U4946 , P1_U4947 , P1_U4948 , P1_U4949 , P1_U4950 , P1_U4951 , P1_U4952 , P1_U4953;
wire P1_U4954 , P1_U4955 , P1_U4956 , P1_U4957 , P1_U4958 , P1_U4959 , P1_U4960 , P1_U4961 , P1_U4962 , P1_U4963;
wire P1_U4964 , P1_U4965 , P1_U4966 , P1_U4967 , P1_U4968 , P1_U4969 , P1_U4970 , P1_U4971 , P1_U4972 , P1_U4973;
wire P1_U4974 , P1_U4975 , P1_U4976 , P1_U4977 , P1_U4978 , P1_U4979 , P1_U4980 , P1_U4981 , P1_U4982 , P1_U4983;
wire P1_U4984 , P1_U4985 , P1_U4986 , P1_U4987 , P1_U4988 , P1_U4989 , P1_U4990 , P1_U4991 , P1_U4992 , P1_U4993;
wire P1_U4994 , P1_U4995 , P1_U4996 , P1_U4997 , P1_U4998 , P1_U4999 , P1_U5000 , P1_U5001 , P1_U5002 , P1_U5003;
wire P1_U5004 , P1_U5005 , P1_U5006 , P1_U5007 , P1_U5008 , P1_U5009 , P1_U5010 , P1_U5011 , P1_U5012 , P1_U5013;
wire P1_U5014 , P1_U5015 , P1_U5016 , P1_U5017 , P1_U5018 , P1_U5019 , P1_U5020 , P1_U5021 , P1_U5022 , P1_U5023;
wire P1_U5024 , P1_U5025 , P1_U5026 , P1_U5027 , P1_U5028 , P1_U5029 , P1_U5030 , P1_U5031 , P1_U5032 , P1_U5033;
wire P1_U5034 , P1_U5035 , P1_U5036 , P1_U5037 , P1_U5038 , P1_U5039 , P1_U5040 , P1_U5041 , P1_U5042 , P1_U5043;
wire P1_U5044 , P1_U5045 , P1_U5046 , P1_U5047 , P1_U5048 , P1_U5049 , P1_U5050 , P1_U5051 , P1_U5052 , P1_U5053;
wire P1_U5054 , P1_U5055 , P1_U5056 , P1_U5057 , P1_U5058 , P1_U5059 , P1_U5060 , P1_U5061 , P1_U5062 , P1_U5063;
wire P1_U5064 , P1_U5065 , P1_U5066 , P1_U5067 , P1_U5068 , P1_U5069 , P1_U5070 , P1_U5071 , P1_U5072 , P1_U5073;
wire P1_U5074 , P1_U5075 , P1_U5076 , P1_U5077 , P1_U5078 , P1_U5079 , P1_U5080 , P1_U5081 , P1_U5082 , P1_U5083;
wire P1_U5084 , P1_U5085 , P1_U5086 , P1_U5087 , P1_U5088 , P1_U5089 , P1_U5090 , P1_U5091 , P1_U5092 , P1_U5093;
wire P1_U5094 , P1_U5095 , P1_U5096 , P1_U5097 , P1_U5098 , P1_U5099 , P1_U5100 , P1_U5101 , P1_U5102 , P1_U5103;
wire P1_U5104 , P1_U5105 , P1_U5106 , P1_U5107 , P1_U5108 , P1_U5109 , P1_U5110 , P1_U5111 , P1_U5112 , P1_U5113;
wire P1_U5114 , P1_U5115 , P1_U5116 , P1_U5117 , P1_U5118 , P1_U5119 , P1_U5120 , P1_U5121 , P1_U5122 , P1_U5123;
wire P1_U5124 , P1_U5125 , P1_U5126 , P1_U5127 , P1_U5128 , P1_U5129 , P1_U5130 , P1_U5131 , P1_U5132 , P1_U5133;
wire P1_U5134 , P1_U5135 , P1_U5136 , P1_U5137 , P1_U5138 , P1_U5139 , P1_U5140 , P1_U5141 , P1_U5142 , P1_U5143;
wire P1_U5144 , P1_U5145 , P1_U5146 , P1_U5147 , P1_U5148 , P1_U5149 , P1_U5150 , P1_U5151 , P1_U5152 , P1_U5153;
wire P1_U5154 , P1_U5155 , P1_U5156 , P1_U5157 , P1_U5158 , P1_U5159 , P1_U5160 , P1_U5161 , P1_U5162 , P1_U5163;
wire P1_U5164 , P1_U5165 , P1_U5166 , P1_U5167 , P1_U5168 , P1_U5169 , P1_U5170 , P1_U5171 , P1_U5172 , P1_U5173;
wire P1_U5174 , P1_U5175 , P1_U5176 , P1_U5177 , P1_U5178 , P1_U5179 , P1_U5180 , P1_U5181 , P1_U5182 , P1_U5183;
wire P1_U5184 , P1_U5185 , P1_U5186 , P1_U5187 , P1_U5188 , P1_U5189 , P1_U5190 , P1_U5191 , P1_U5192 , P1_U5193;
wire P1_U5194 , P1_U5195 , P1_U5196 , P1_U5197 , P1_U5198 , P1_U5199 , P1_U5200 , P1_U5201 , P1_U5202 , P1_U5203;
wire P1_U5204 , P1_U5205 , P1_U5206 , P1_U5207 , P1_U5208 , P1_U5209 , P1_U5210 , P1_U5211 , P1_U5212 , P1_U5213;
wire P1_U5214 , P1_U5215 , P1_U5216 , P1_U5217 , P1_U5218 , P1_U5219 , P1_U5220 , P1_U5221 , P1_U5222 , P1_U5223;
wire P1_U5224 , P1_U5225 , P1_U5226 , P1_U5227 , P1_U5228 , P1_U5229 , P1_U5230 , P1_U5231 , P1_U5232 , P1_U5233;
wire P1_U5234 , P1_U5235 , P1_U5236 , P1_U5237 , P1_U5238 , P1_U5239 , P1_U5240 , P1_U5241 , P1_U5242 , P1_U5243;
wire P1_U5244 , P1_U5245 , P1_U5246 , P1_U5247 , P1_U5248 , P1_U5249 , P1_U5250 , P1_U5251 , P1_U5252 , P1_U5253;
wire P1_U5254 , P1_U5255 , P1_U5256 , P1_U5257 , P1_U5258 , P1_U5259 , P1_U5260 , P1_U5261 , P1_U5262 , P1_U5263;
wire P1_U5264 , P1_U5265 , P1_U5266 , P1_U5267 , P1_U5268 , P1_U5269 , P1_U5270 , P1_U5271 , P1_U5272 , P1_U5273;
wire P1_U5274 , P1_U5275 , P1_U5276 , P1_U5277 , P1_U5278 , P1_U5279 , P1_U5280 , P1_U5281 , P1_U5282 , P1_U5283;
wire P1_U5284 , P1_U5285 , P1_U5286 , P1_U5287 , P1_U5288 , P1_U5289 , P1_U5290 , P1_U5291 , P1_U5292 , P1_U5293;
wire P1_U5294 , P1_U5295 , P1_U5296 , P1_U5297 , P1_U5298 , P1_U5299 , P1_U5300 , P1_U5301 , P1_U5302 , P1_U5303;
wire P1_U5304 , P1_U5305 , P1_U5306 , P1_U5307 , P1_U5308 , P1_U5309 , P1_U5310 , P1_U5311 , P1_U5312 , P1_U5313;
wire P1_U5314 , P1_U5315 , P1_U5316 , P1_U5317 , P1_U5318 , P1_U5319 , P1_U5320 , P1_U5321 , P1_U5322 , P1_U5323;
wire P1_U5324 , P1_U5325 , P1_U5326 , P1_U5327 , P1_U5328 , P1_U5329 , P1_U5330 , P1_U5331 , P1_U5332 , P1_U5333;
wire P1_U5334 , P1_U5335 , P1_U5336 , P1_U5337 , P1_U5338 , P1_U5339 , P1_U5340 , P1_U5341 , P1_U5342 , P1_U5343;
wire P1_U5344 , P1_U5345 , P1_U5346 , P1_U5347 , P1_U5348 , P1_U5349 , P1_U5350 , P1_U5351 , P1_U5352 , P1_U5353;
wire P1_U5354 , P1_U5355 , P1_U5356 , P1_U5357 , P1_U5358 , P1_U5359 , P1_U5360 , P1_U5361 , P1_U5362 , P1_U5363;
wire P1_U5364 , P1_U5365 , P1_U5366 , P1_U5367 , P1_U5368 , P1_U5369 , P1_U5370 , P1_U5371 , P1_U5372 , P1_U5373;
wire P1_U5374 , P1_U5375 , P1_U5376 , P1_U5377 , P1_U5378 , P1_U5379 , P1_U5380 , P1_U5381 , P1_U5382 , P1_U5383;
wire P1_U5384 , P1_U5385 , P1_U5386 , P1_U5387 , P1_U5388 , P1_U5389 , P1_U5390 , P1_U5391 , P1_U5392 , P1_U5393;
wire P1_U5394 , P1_U5395 , P1_U5396 , P1_U5397 , P1_U5398 , P1_U5399 , P1_U5400 , P1_U5401 , P1_U5402 , P1_U5403;
wire P1_U5404 , P1_U5405 , P1_U5406 , P1_U5407 , P1_U5408 , P1_U5409 , P1_U5410 , P1_U5411 , P1_U5412 , P1_U5413;
wire P1_U5414 , P1_U5415 , P1_U5416 , P1_U5417 , P1_U5418 , P1_U5419 , P1_U5420 , P1_U5421 , P1_U5422 , P1_U5423;
wire P1_U5424 , P1_U5425 , P1_U5426 , P1_U5427 , P1_U5428 , P1_U5429 , P1_U5430 , P1_U5431 , P1_U5432 , P1_U5433;
wire P1_U5434 , P1_U5435 , P1_U5436 , P1_U5437 , P1_U5438 , P1_U5439 , P1_U5440 , P1_U5441 , P1_U5442 , P1_U5443;
wire P1_U5444 , P1_U5445 , P1_U5446 , P1_U5447 , P1_U5448 , P1_U5449 , P1_U5450 , P1_U5451 , P1_U5452 , P1_U5453;
wire P1_U5454 , P1_U5455 , P1_U5456 , P1_U5457 , P1_U5458 , P1_U5459 , P1_U5460 , P1_U5461 , P1_U5462 , P1_U5463;
wire P1_U5464 , P1_U5465 , P1_U5466 , P1_U5467 , P1_U5468 , P1_U5469 , P1_U5470 , P1_U5471 , P1_U5472 , P1_U5473;
wire P1_U5474 , P1_U5475 , P1_U5476 , P1_U5477 , P1_U5478 , P1_U5479 , P1_U5480 , P1_U5481 , P1_U5482 , P1_U5483;
wire P1_U5484 , P1_U5485 , P1_U5486 , P1_U5487 , P1_U5488 , P1_U5489 , P1_U5490 , P1_U5491 , P1_U5492 , P1_U5493;
wire P1_U5494 , P1_U5495 , P1_U5496 , P1_U5497 , P1_U5498 , P1_U5499 , P1_U5500 , P1_U5501 , P1_U5502 , P1_U5503;
wire P1_U5504 , P1_U5505 , P1_U5506 , P1_U5507 , P1_U5508 , P1_U5509 , P1_U5510 , P1_U5511 , P1_U5512 , P1_U5513;
wire P1_U5514 , P1_U5515 , P1_U5516 , P1_U5517 , P1_U5518 , P1_U5519 , P1_U5520 , P1_U5521 , P1_U5522 , P1_U5523;
wire P1_U5524 , P1_U5525 , P1_U5526 , P1_U5527 , P1_U5528 , P1_U5529 , P1_U5530 , P1_U5531 , P1_U5532 , P1_U5533;
wire P1_U5534 , P1_U5535 , P1_U5536 , P1_U5537 , P1_U5538 , P1_U5539 , P1_U5540 , P1_U5541 , P1_U5542 , P1_U5543;
wire P1_U5544 , P1_U5545 , P1_U5546 , P1_U5547 , P1_U5548 , P1_U5549 , P1_U5550 , P1_U5551 , P1_U5552 , P1_U5553;
wire P1_U5554 , P1_U5555 , P1_U5556 , P1_U5557 , P1_U5558 , P1_U5559 , P1_U5560 , P1_U5561 , P1_U5562 , P1_U5563;
wire P1_U5564 , P1_U5565 , P1_U5566 , P1_U5567 , P1_U5568 , P1_U5569 , P1_U5570 , P1_U5571 , P1_U5572 , P1_U5573;
wire P1_U5574 , P1_U5575 , P1_U5576 , P1_U5577 , P1_U5578 , P1_U5579 , P1_U5580 , P1_U5581 , P1_U5582 , P1_U5583;
wire P1_U5584 , P1_U5585 , P1_U5586 , P1_U5587 , P1_U5588 , P1_U5589 , P1_U5590 , P1_U5591 , P1_U5592 , P1_U5593;
wire P1_U5594 , P1_U5595 , P1_U5596 , P1_U5597 , P1_U5598 , P1_U5599 , P1_U5600 , P1_U5601 , P1_U5602 , P1_U5603;
wire P1_U5604 , P1_U5605 , P1_U5606 , P1_U5607 , P1_U5608 , P1_U5609 , P1_U5610 , P1_U5611 , P1_U5612 , P1_U5613;
wire P1_U5614 , P1_U5615 , P1_U5616 , P1_U5617 , P1_U5618 , P1_U5619 , P1_U5620 , P1_U5621 , P1_U5622 , P1_U5623;
wire P1_U5624 , P1_U5625 , P1_U5626 , P1_U5627 , P1_U5628 , P1_U5629 , P1_U5630 , P1_U5631 , P1_U5632 , P1_U5633;
wire P1_U5634 , P1_U5635 , P1_U5636 , P1_U5637 , P1_U5638 , P1_U5639 , P1_U5640 , P1_U5641 , P1_U5642 , P1_U5643;
wire P1_U5644 , P1_U5645 , P1_U5646 , P1_U5647 , P1_U5648 , P1_U5649 , P1_U5650 , P1_U5651 , P1_U5652 , P1_U5653;
wire P1_U5654 , P1_U5655 , P1_U5656 , P1_U5657 , P1_U5658 , P1_U5659 , P1_U5660 , P1_U5661 , P1_U5662 , P1_U5663;
wire P1_U5664 , P1_U5665 , P1_U5666 , P1_U5667 , P1_U5668 , P1_U5669 , P1_U5670 , P1_U5671 , P1_U5672 , P1_U5673;
wire P1_U5674 , P1_U5675 , P1_U5676 , P1_U5677 , P1_U5678 , P1_U5679 , P1_U5680 , P1_U5681 , P1_U5682 , P1_U5683;
wire P1_U5684 , P1_U5685 , P1_U5686 , P1_U5687 , P1_U5688 , P1_U5689 , P1_U5690 , P1_U5691 , P1_U5692 , P1_U5693;
wire P1_U5694 , P1_U5695 , P1_U5696 , P1_U5697 , P1_U5698 , P1_U5699 , P1_U5700 , P1_U5701 , P1_U5702 , P1_U5703;
wire P1_U5704 , P1_U5705 , P1_U5706 , P1_U5707 , P1_U5708 , P1_U5709 , P1_U5710 , P1_U5711 , P1_U5712 , P1_U5713;
wire P1_U5714 , P1_U5715 , P1_U5716 , P1_U5717 , P1_U5718 , P1_U5719 , P1_U5720 , P1_U5721 , P1_U5722 , P1_U5723;
wire P1_U5724 , P1_U5725 , P1_U5726 , P1_U5727 , P1_U5728 , P1_U5729 , P1_U5730 , P1_U5731 , P1_U5732 , P1_U5733;
wire P1_U5734 , P1_U5735 , P1_U5736 , P1_U5737 , P1_U5738 , P1_U5739 , P1_U5740 , P1_U5741 , P1_U5742 , P1_U5743;
wire P1_U5744 , P1_U5745 , P1_U5746 , P1_U5747 , P1_U5748 , P1_U5749 , P1_U5750 , P1_U5751 , P1_U5752 , P1_U5753;
wire P1_U5754 , P1_U5755 , P1_U5756 , P1_U5757 , P1_U5758 , P1_U5759 , P1_U5760 , P1_U5761 , P1_U5762 , P1_U5763;
wire P1_U5764 , P1_U5765 , P1_U5766 , P1_U5767 , P1_U5768 , P1_U5769 , P1_U5770 , P1_U5771 , P1_U5772 , P1_U5773;
wire P1_U5774 , P1_U5775 , P1_U5776 , P1_U5777 , P1_U5778 , P1_U5779 , P1_U5780 , P1_U5781 , P1_U5782 , P1_U5783;
wire P1_U5784 , P1_U5785 , P1_U5786 , P1_U5787 , P1_U5788 , P1_U5789 , P1_U5790 , P1_U5791 , P1_U5792 , P1_U5793;
wire P1_U5794 , P1_U5795 , P1_U5796 , P1_U5797 , P1_U5798 , P1_U5799 , P1_U5800 , P1_U5801 , P1_U5802 , P1_U5803;
wire P1_U5804 , P1_U5805 , P1_U5806 , P1_U5807 , P1_U5808 , P1_U5809 , P1_U5810 , P1_U5811 , P1_U5812 , P1_U5813;
wire P1_U5814 , P1_U5815 , P1_U5816 , P1_U5817 , P1_U5818 , P1_U5819 , P1_U5820 , P1_U5821 , P1_U5822 , P1_U5823;
wire P1_U5824 , P1_U5825 , P1_U5826 , P1_U5827 , P1_U5828 , P1_U5829 , P1_U5830 , P1_U5831 , P1_U5832 , P1_U5833;
wire P1_U5834 , P1_U5835 , P1_U5836 , P1_U5837 , P1_U5838 , P1_U5839 , P1_U5840 , P1_U5841 , P1_U5842 , P1_U5843;
wire P1_U5844 , P1_U5845 , P1_U5846 , P1_U5847 , P1_U5848 , P1_U5849 , P1_U5850 , P1_U5851 , P1_U5852 , P1_U5853;
wire P1_U5854 , P1_U5855 , P1_U5856 , P1_U5857 , P1_U5858 , P1_U5859 , P1_U5860 , P1_U5861 , P1_U5862 , P1_U5863;
wire P1_U5864 , P1_U5865 , P1_U5866 , P1_U5867 , P1_U5868 , P1_U5869 , P1_U5870 , P1_U5871 , P1_U5872 , P1_U5873;
wire P1_U5874 , P1_U5875 , P1_U5876 , P1_U5877 , P1_U5878 , P1_U5879 , P1_U5880 , P1_U5881 , P1_U5882 , P1_U5883;
wire P1_U5884 , P1_U5885 , P1_U5886 , P1_U5887 , P1_U5888 , P1_U5889 , P1_U5890 , P1_U5891 , P1_U5892 , P1_U5893;
wire P1_U5894 , P1_U5895 , P1_U5896 , P1_U5897 , P1_U5898 , P1_U5899 , P1_U5900 , P1_U5901 , P1_U5902 , P1_U5903;
wire P1_U5904 , P1_U5905 , P1_U5906 , P1_U5907 , P1_U5908 , P1_U5909 , P1_U5910 , P1_U5911 , P1_U5912 , P1_U5913;
wire P1_U5914 , P1_U5915 , P1_U5916 , P1_U5917 , P1_U5918 , P1_U5919 , P1_U5920 , P1_U5921 , P1_U5922 , P1_U5923;
wire P1_U5924 , P1_U5925 , P1_U5926 , P1_U5927 , P1_U5928 , P1_U5929 , P1_U5930 , P1_U5931 , P1_U5932 , P1_U5933;
wire P1_U5934 , P1_U5935 , P1_U5936 , P1_U5937 , P1_U5938 , P1_U5939 , P1_U5940 , P1_U5941 , P1_U5942 , P1_U5943;
wire P1_U5944 , P1_U5945 , P1_U5946 , P1_U5947 , P1_U5948 , P1_U5949 , P1_U5950 , P1_U5951 , P1_U5952 , P1_U5953;
wire P1_U5954 , P1_U5955 , P1_U5956 , P1_U5957 , P1_U5958 , P1_U5959 , P1_U5960 , P1_U5961 , P1_U5962 , P1_U5963;
wire P1_U5964 , P1_U5965 , P1_U5966 , P1_U5967 , P1_U5968 , P1_U5969 , P1_U5970 , P1_U5971 , P1_U5972 , P1_U5973;
wire P1_U5974 , P1_U5975 , P1_U5976 , P1_U5977 , P1_U5978 , P1_U5979 , P1_U5980 , P1_U5981 , P1_U5982 , P1_U5983;
wire P1_U5984 , P1_U5985 , P1_U5986 , P1_U5987 , P1_U5988 , P1_U5989 , P1_U5990 , P1_U5991 , P1_U5992 , P1_U5993;
wire P1_U5994 , P1_U5995 , P1_U5996 , P1_U5997 , P1_U5998 , P1_U5999 , P1_U6000 , P1_U6001 , P1_U6002 , P1_U6003;
wire P1_U6004 , P1_U6005 , P1_U6006 , P1_U6007 , P1_U6008 , P1_U6009 , P1_U6010 , P1_U6011 , P1_U6012 , P1_U6013;
wire P1_U6014 , P1_U6015 , P1_U6016 , P1_U6017 , P1_U6018 , P1_U6019 , P1_U6020 , P1_U6021 , P1_U6022 , P1_U6023;
wire P1_U6024 , P1_U6025 , P1_U6026 , P1_U6027 , P1_U6028 , P1_U6029 , P1_U6030 , P1_U6031 , P1_U6032 , P1_U6033;
wire P1_U6034 , P1_U6035 , P1_U6036 , P1_U6037 , P1_U6038 , P1_U6039 , P1_U6040 , P1_U6041 , P1_U6042 , P1_U6043;
wire P1_U6044 , P1_U6045 , P1_U6046 , P1_U6047 , P1_U6048 , P1_U6049 , P1_U6050 , P1_U6051 , P1_U6052 , P1_U6053;
wire P1_U6054 , P1_U6055 , P1_U6056 , P1_U6057 , P1_U6058 , P1_U6059 , P1_U6060 , P1_U6061 , P1_U6062 , P1_U6063;
wire P1_U6064 , P1_U6065 , P1_U6066 , P1_U6067 , P1_U6068 , P1_U6069 , P1_U6070 , P1_U6071 , P1_U6072 , P1_U6073;
wire P1_U6074 , P1_U6075 , P1_U6076 , P1_U6077 , P1_U6078 , P1_U6079 , P1_U6080 , P1_U6081 , P1_U6082 , P1_U6083;
wire P1_U6084 , P1_U6085 , P1_U6086 , P1_U6087 , P1_U6088 , P1_U6089 , P1_U6090 , P1_U6091 , P1_U6092 , P1_U6093;
wire P1_U6094 , P1_U6095 , P1_U6096 , P1_U6097 , P1_U6098 , P1_U6099 , P1_U6100 , P1_U6101 , P1_U6102 , P1_U6103;
wire P1_U6104 , P1_U6105 , P1_U6106 , P1_U6107 , P1_U6108 , P1_U6109 , P1_U6110 , P1_U6111 , P1_U6112 , P1_U6113;
wire P1_U6114 , P1_U6115 , P1_U6116 , P1_U6117 , P1_U6118 , P1_U6119 , P1_U6120 , P1_U6121 , P1_U6122 , P1_U6123;
wire P1_U6124 , P1_U6125 , P1_U6126 , P1_U6127 , P1_U6128 , P1_U6129 , P1_U6130 , P1_U6131 , P1_U6132 , P1_U6133;
wire P1_U6134 , P1_U6135 , P1_U6136 , P1_U6137 , P1_U6138 , P1_U6139 , P1_U6140 , P1_U6141 , P1_U6142 , P1_U6143;
wire P1_U6144 , P1_U6145 , P1_U6146 , P1_U6147 , P1_U6148 , P1_U6149 , P1_U6150 , P1_U6151 , P1_U6152 , P1_U6153;
wire P1_U6154 , P1_U6155 , P1_U6156 , P1_U6157 , P1_U6158 , P1_U6159 , P1_U6160 , P1_U6161 , P1_U6162 , P1_U6163;
wire P1_U6164 , P1_U6165 , P1_U6166 , P1_U6167 , P1_U6168 , P1_U6169 , P1_U6170 , P1_U6171 , P1_U6172 , P1_U6173;
wire P1_U6174 , P1_U6175 , P1_U6176 , P1_U6177 , P1_U6178 , P1_U6179 , P1_U6180 , P1_U6181 , P1_U6182 , P1_U6183;
wire P1_U6184 , P1_U6185 , P1_U6186 , P1_U6187 , P1_U6188 , P1_U6189 , P1_U6190 , P1_U6191 , P1_U6192 , P1_U6193;
wire P1_U6194 , P1_U6195 , P1_U6196 , P1_U6197 , P1_U6198 , P1_U6199 , P1_U6200 , P1_U6201 , P1_U6202 , P1_U6203;
wire P1_U6204 , P1_U6205 , P1_U6206 , P1_U6207 , P1_U6208 , P1_U6209 , P1_U6210 , P1_U6211 , P1_U6212 , P1_U6213;
wire P1_U6214 , P1_U6215 , P1_U6216 , P1_U6217 , P1_U6218 , P1_U6219 , P1_U6220 , P1_U6221 , P1_U6222 , P1_U6223;
wire P1_U6224 , P1_U6225 , P1_U6226 , P1_U6227 , P1_U6228 , P1_U6229 , P1_U6230 , P1_U6231 , P1_U6232 , P1_U6233;
wire P1_U6234 , P1_U6235 , P1_U6236 , P2_R1161_U489 , P2_R1161_U488 , P2_R1161_U487 , P2_R1161_U486 , P2_R1161_U485 , P2_R1161_U484 , P2_R1161_U483;
wire P2_R1161_U482 , P2_R1161_U481 , P2_R1161_U480 , P2_R1161_U479 , P2_R1161_U478 , P2_R1161_U477 , P2_R1161_U476 , P2_R1161_U475 , P2_R1161_U474 , P2_R1161_U473;
wire P2_R1161_U472 , P2_R1161_U471 , P2_R1161_U470 , P2_R1161_U469 , P2_R1161_U468 , P2_R1161_U467 , P2_R1161_U466 , P2_U3013 , P2_U3014 , P2_U3015;
wire P2_U3016 , P2_U3017 , P2_U3018 , P2_U3019 , P2_U3020 , P2_U3021 , P2_U3022 , P2_U3023 , P2_U3024 , P2_U3025;
wire P2_U3026 , P2_U3027 , P2_U3028 , P2_U3029 , P2_U3030 , P2_U3031 , P2_U3032 , P2_U3033 , P2_U3034 , P2_U3035;
wire P2_U3036 , P2_U3037 , P2_U3038 , P2_U3039 , P2_U3040 , P2_U3041 , P2_U3042 , P2_U3043 , P2_U3044 , P2_U3045;
wire P2_U3046 , P2_U3047 , P2_U3048 , P2_U3049 , P2_U3050 , P2_U3051 , P2_U3052 , P2_U3053 , P2_U3054 , P2_U3055;
wire P2_U3056 , P2_U3057 , P2_U3058 , P2_U3059 , P2_U3060 , P2_U3061 , P2_U3062 , P2_U3063 , P2_U3064 , P2_U3065;
wire P2_U3066 , P2_U3067 , P2_U3068 , P2_U3069 , P2_U3070 , P2_U3071 , P2_U3072 , P2_U3073 , P2_U3074 , P2_U3075;
wire P2_U3076 , P2_U3077 , P2_U3078 , P2_U3079 , P2_U3080 , P2_U3081 , P2_U3082 , P2_U3083 , P2_U3084 , P2_U3085;
wire P2_U3086 , P2_U3087 , P2_U3088 , P2_U3089 , P2_U3090 , P2_U3091 , P2_U3092 , P2_U3093 , P2_U3094 , P2_U3095;
wire P2_U3096 , P2_U3097 , P2_U3098 , P2_U3099 , P2_U3100 , P2_U3101 , P2_U3102 , P2_U3103 , P2_U3104 , P2_U3105;
wire P2_U3106 , P2_U3107 , P2_U3108 , P2_U3109 , P2_U3110 , P2_U3111 , P2_U3112 , P2_U3113 , P2_U3114 , P2_U3115;
wire P2_U3116 , P2_U3117 , P2_U3118 , P2_U3119 , P2_U3120 , P2_U3121 , P2_U3122 , P2_U3123 , P2_U3124 , P2_U3125;
wire P2_U3126 , P2_U3127 , P2_U3128 , P2_U3129 , P2_U3130 , P2_U3131 , P2_U3132 , P2_U3133 , P2_U3134 , P2_U3135;
wire P2_U3136 , P2_U3137 , P2_U3138 , P2_U3139 , P2_U3140 , P2_U3141 , P2_U3142 , P2_U3143 , P2_U3144 , P2_U3145;
wire P2_U3146 , P2_U3147 , P2_U3148 , P2_U3149 , P2_U3152 , P2_U3297 , P2_U3298 , P2_U3299 , P2_U3300 , P2_U3301;
wire P2_U3302 , P2_U3303 , P2_U3304 , P2_U3305 , P2_U3306 , P2_U3307 , P2_U3308 , P2_U3309 , P2_U3310 , P2_U3311;
wire P2_U3312 , P2_U3313 , P2_U3314 , P2_U3315 , P2_U3316 , P2_U3317 , P2_U3318 , P2_U3319 , P2_U3320 , P2_U3321;
wire P2_U3322 , P2_U3323 , P2_U3324 , P2_U3325 , P2_U3326 , P2_U3327 , P2_U3328 , P2_U3329 , P2_U3330 , P2_U3331;
wire P2_U3332 , P2_U3333 , P2_U3334 , P2_U3335 , P2_U3336 , P2_U3337 , P2_U3338 , P2_U3339 , P2_U3340 , P2_U3341;
wire P2_U3342 , P2_U3343 , P2_U3344 , P2_U3345 , P2_U3346 , P2_U3347 , P2_U3348 , P2_U3349 , P2_U3350 , P2_U3351;
wire P2_U3352 , P2_U3353 , P2_U3354 , P2_U3355 , P2_U3356 , P2_U3357 , P2_U3358 , P2_U3359 , P2_U3360 , P2_U3361;
wire P2_U3362 , P2_U3363 , P2_U3364 , P2_U3365 , P2_U3366 , P2_U3367 , P2_U3368 , P2_U3369 , P2_U3370 , P2_U3371;
wire P2_U3372 , P2_U3373 , P2_U3374 , P2_U3375 , P2_U3378 , P2_U3379 , P2_U3380 , P2_U3381 , P2_U3382 , P2_U3383;
wire P2_U3384 , P2_U3385 , P2_U3386 , P2_U3387 , P2_U3388 , P2_U3389 , P2_U3391 , P2_U3392 , P2_U3394 , P2_U3395;
wire P2_U3397 , P2_U3398 , P2_U3400 , P2_U3401 , P2_U3403 , P2_U3404 , P2_U3406 , P2_U3407 , P2_U3409 , P2_U3410;
wire P2_U3412 , P2_U3413 , P2_U3415 , P2_U3416 , P2_U3418 , P2_U3419 , P2_U3421 , P2_U3422 , P2_U3424 , P2_U3425;
wire P2_U3427 , P2_U3428 , P2_U3430 , P2_U3431 , P2_U3433 , P2_U3434 , P2_U3436 , P2_U3437 , P2_U3439 , P2_U3440;
wire P2_U3442 , P2_U3443 , P2_U3445 , P2_U3523 , P2_U3524 , P2_U3525 , P2_U3526 , P2_U3527 , P2_U3528 , P2_U3529;
wire P2_U3530 , P2_U3531 , P2_U3532 , P2_U3533 , P2_U3534 , P2_U3535 , P2_U3536 , P2_U3537 , P2_U3538 , P2_U3539;
wire P2_U3540 , P2_U3541 , P2_U3542 , P2_U3543 , P2_U3544 , P2_U3545 , P2_U3546 , P2_U3547 , P2_U3548 , P2_U3549;
wire P2_U3550 , P2_U3551 , P2_U3552 , P2_U3553 , P2_U3554 , P2_U3555 , P2_U3556 , P2_U3557 , P2_U3558 , P2_U3559;
wire P2_U3560 , P2_U3561 , P2_U3562 , P2_U3563 , P2_U3564 , P2_U3565 , P2_U3566 , P2_U3567 , P2_U3568 , P2_U3569;
wire P2_U3570 , P2_U3571 , P2_U3572 , P2_U3573 , P2_U3574 , P2_U3575 , P2_U3576 , P2_U3577 , P2_U3578 , P2_U3579;
wire P2_U3580 , P2_U3581 , P2_U3582 , P2_U3583 , P2_U3584 , P2_U3585 , P2_U3586 , P2_U3587 , P2_U3588 , P2_U3589;
wire P2_U3590 , P2_U3591 , P2_U3592 , P2_U3593 , P2_U3594 , P2_U3595 , P2_U3596 , P2_U3597 , P2_U3598 , P2_U3599;
wire P2_U3600 , P2_U3601 , P2_U3602 , P2_U3603 , P2_U3604 , P2_U3605 , P2_U3606 , P2_U3607 , P2_U3608 , P2_U3609;
wire P2_U3610 , P2_U3611 , P2_U3612 , P2_U3613 , P2_U3614 , P2_U3615 , P2_U3616 , P2_U3617 , P2_U3618 , P2_U3619;
wire P2_U3620 , P2_U3621 , P2_U3622 , P2_U3623 , P2_U3624 , P2_U3625 , P2_U3626 , P2_U3627 , P2_U3628 , P2_U3629;
wire P2_U3630 , P2_U3631 , P2_U3632 , P2_U3633 , P2_U3634 , P2_U3635 , P2_U3636 , P2_U3637 , P2_U3638 , P2_U3639;
wire P2_U3640 , P2_U3641 , P2_U3642 , P2_U3643 , P2_U3644 , P2_U3645 , P2_U3646 , P2_U3647 , P2_U3648 , P2_U3649;
wire P2_U3650 , P2_U3651 , P2_U3652 , P2_U3653 , P2_U3654 , P2_U3655 , P2_U3656 , P2_U3657 , P2_U3658 , P2_U3659;
wire P2_U3660 , P2_U3661 , P2_U3662 , P2_U3663 , P2_U3664 , P2_U3665 , P2_U3666 , P2_U3667 , P2_U3668 , P2_U3669;
wire P2_U3670 , P2_U3671 , P2_U3672 , P2_U3673 , P2_U3674 , P2_U3675 , P2_U3676 , P2_U3677 , P2_U3678 , P2_U3679;
wire P2_U3680 , P2_U3681 , P2_U3682 , P2_U3683 , P2_U3684 , P2_U3685 , P2_U3686 , P2_U3687 , P2_U3688 , P2_U3689;
wire P2_U3690 , P2_U3691 , P2_U3692 , P2_U3693 , P2_U3694 , P2_U3695 , P2_U3696 , P2_U3697 , P2_U3698 , P2_U3699;
wire P2_U3700 , P2_U3701 , P2_U3702 , P2_U3703 , P2_U3704 , P2_U3705 , P2_U3706 , P2_U3707 , P2_U3708 , P2_U3709;
wire P2_U3710 , P2_U3711 , P2_U3712 , P2_U3713 , P2_U3714 , P2_U3715 , P2_U3716 , P2_U3717 , P2_U3718 , P2_U3719;
wire P2_U3720 , P2_U3721 , P2_U3722 , P2_U3723 , P2_U3724 , P2_U3725 , P2_U3726 , P2_U3727 , P2_U3728 , P2_U3729;
wire P2_U3730 , P2_U3731 , P2_U3732 , P2_U3733 , P2_U3734 , P2_U3735 , P2_U3736 , P2_U3737 , P2_U3738 , P2_U3739;
wire P2_U3740 , P2_U3741 , P2_U3742 , P2_U3743 , P2_U3744 , P2_U3745 , P2_U3746 , P2_U3747 , P2_U3748 , P2_U3749;
wire P2_U3750 , P2_U3751 , P2_U3752 , P2_U3753 , P2_U3754 , P2_U3755 , P2_U3756 , P2_U3757 , P2_U3758 , P2_U3759;
wire P2_U3760 , P2_U3761 , P2_U3762 , P2_U3763 , P2_U3764 , P2_U3765 , P2_U3766 , P2_U3767 , P2_U3768 , P2_U3769;
wire P2_U3770 , P2_U3771 , P2_U3772 , P2_U3773 , P2_U3774 , P2_U3775 , P2_U3776 , P2_U3777 , P2_U3778 , P2_U3779;
wire P2_U3780 , P2_U3781 , P2_U3782 , P2_U3783 , P2_U3784 , P2_U3785 , P2_U3786 , P2_U3787 , P2_U3788 , P2_U3789;
wire P2_U3790 , P2_U3791 , P2_U3792 , P2_U3793 , P2_U3794 , P2_U3795 , P2_U3796 , P2_U3797 , P2_U3798 , P2_U3799;
wire P2_U3800 , P2_U3801 , P2_U3802 , P2_U3803 , P2_U3804 , P2_U3805 , P2_U3806 , P2_U3807 , P2_U3808 , P2_U3809;
wire P2_U3810 , P2_U3811 , P2_U3812 , P2_U3813 , P2_U3814 , P2_U3815 , P2_U3816 , P2_U3817 , P2_U3818 , P2_U3819;
wire P2_U3820 , P2_U3821 , P2_U3822 , P2_U3823 , P2_U3824 , P2_U3825 , P2_U3826 , P2_U3827 , P2_U3828 , P2_U3829;
wire P2_U3830 , P2_U3831 , P2_U3832 , P2_U3833 , P2_U3834 , P2_U3835 , P2_U3836 , P2_U3837 , P2_U3838 , P2_U3839;
wire P2_U3840 , P2_U3841 , P2_U3842 , P2_U3843 , P2_U3844 , P2_U3845 , P2_U3846 , P2_U3847 , P2_U3848 , P2_U3849;
wire P2_U3850 , P2_U3851 , P2_U3852 , P2_U3853 , P2_U3854 , P2_U3855 , P2_U3856 , P2_U3857 , P2_U3858 , P2_U3859;
wire P2_U3860 , P2_U3861 , P2_U3862 , P2_U3863 , P2_U3864 , P2_U3865 , P2_U3866 , P2_U3867 , P2_U3868 , P2_U3869;
wire P2_U3870 , P2_U3871 , P2_U3872 , P2_U3873 , P2_U3874 , P2_U3875 , P2_U3876 , P2_U3877 , P2_U3878 , P2_U3879;
wire P2_U3880 , P2_U3881 , P2_U3882 , P2_U3883 , P2_U3884 , P2_U3885 , P2_U3886 , P2_U3887 , P2_U3888 , P2_U3889;
wire P2_U3890 , P2_U3891 , P2_U3892 , P2_U3894 , P2_U3895 , P2_U3896 , P2_U3897 , P2_U3898 , P2_U3899 , P2_U3900;
wire P2_U3901 , P2_U3902 , P2_U3903 , P2_U3904 , P2_U3905 , P2_U3906 , P2_U3907 , P2_U3908 , P2_U3909 , P2_U3910;
wire P2_U3911 , P2_U3912 , P2_U3913 , P2_U3914 , P2_U3915 , P2_U3916 , P2_U3917 , P2_U3918 , P2_U3919 , P2_U3920;
wire P2_U3921 , P2_U3922 , P2_U3923 , P2_U3924 , P2_U3925 , P2_U3926 , P2_U3927 , P2_U3928 , P2_U3929 , P2_U3930;
wire P2_U3931 , P2_U3932 , P2_U3933 , P2_U3934 , P2_U3935 , P2_U3936 , P2_U3937 , P2_U3938 , P2_U3939 , P2_U3940;
wire P2_U3941 , P2_U3942 , P2_U3943 , P2_U3944 , P2_U3945 , P2_U3946 , P2_U3947 , P2_U3948 , P2_U3949 , P2_U3950;
wire P2_U3951 , P2_U3952 , P2_U3953 , P2_U3954 , P2_U3955 , P2_U3956 , P2_U3957 , P2_U3958 , P2_U3959 , P2_U3960;
wire P2_U3961 , P2_U3962 , P2_U3963 , P2_U3964 , P2_U3965 , P2_U3966 , P2_U3967 , P2_U3968 , P2_U3969 , P2_U3970;
wire P2_U3971 , P2_U3972 , P2_U3973 , P2_U3974 , P2_U3975 , P2_U3976 , P2_U3977 , P2_U3978 , P2_U3979 , P2_U3980;
wire P2_U3981 , P2_U3982 , P2_U3983 , P2_U3984 , P2_U3985 , P2_U3986 , P2_U3987 , P2_U3988 , P2_U3989 , P2_U3990;
wire P2_U3991 , P2_U3992 , P2_U3993 , P2_U3994 , P2_U3995 , P2_U3996 , P2_U3997 , P2_U3998 , P2_U3999 , P2_U4000;
wire P2_U4001 , P2_U4002 , P2_U4003 , P2_U4004 , P2_U4005 , P2_U4006 , P2_U4007 , P2_U4008 , P2_U4009 , P2_U4010;
wire P2_U4011 , P2_U4012 , P2_U4013 , P2_U4014 , P2_U4015 , P2_U4016 , P2_U4017 , P2_U4018 , P2_U4019 , P2_U4020;
wire P2_U4021 , P2_U4022 , P2_U4023 , P2_U4024 , P2_U4025 , P2_U4026 , P2_U4027 , P2_U4028 , P2_U4029 , P2_U4030;
wire P2_U4031 , P2_U4032 , P2_U4033 , P2_U4034 , P2_U4035 , P2_U4036 , P2_U4037 , P2_U4038 , P2_U4039 , P2_U4040;
wire P2_U4041 , P2_U4042 , P2_U4043 , P2_U4044 , P2_U4045 , P2_U4046 , P2_U4047 , P2_U4048 , P2_U4049 , P2_U4050;
wire P2_U4051 , P2_U4052 , P2_U4053 , P2_U4054 , P2_U4055 , P2_U4056 , P2_U4057 , P2_U4058 , P2_U4059 , P2_U4060;
wire P2_U4061 , P2_U4062 , P2_U4063 , P2_U4064 , P2_U4065 , P2_U4066 , P2_U4067 , P2_U4068 , P2_U4069 , P2_U4070;
wire P2_U4071 , P2_U4072 , P2_U4073 , P2_U4074 , P2_U4075 , P2_U4076 , P2_U4077 , P2_U4078 , P2_U4079 , P2_U4080;
wire P2_U4081 , P2_U4082 , P2_U4083 , P2_U4084 , P2_U4085 , P2_U4086 , P2_U4087 , P2_U4088 , P2_U4089 , P2_U4090;
wire P2_U4091 , P2_U4092 , P2_U4093 , P2_U4094 , P2_U4095 , P2_U4096 , P2_U4097 , P2_U4098 , P2_U4099 , P2_U4100;
wire P2_U4101 , P2_U4102 , P2_U4103 , P2_U4104 , P2_U4105 , P2_U4106 , P2_U4107 , P2_U4108 , P2_U4109 , P2_U4110;
wire P2_U4111 , P2_U4112 , P2_U4113 , P2_U4114 , P2_U4115 , P2_U4116 , P2_U4117 , P2_U4118 , P2_U4119 , P2_U4120;
wire P2_U4121 , P2_U4122 , P2_U4123 , P2_U4124 , P2_U4125 , P2_U4126 , P2_U4127 , P2_U4128 , P2_U4129 , P2_U4130;
wire P2_U4131 , P2_U4132 , P2_U4133 , P2_U4134 , P2_U4135 , P2_U4136 , P2_U4137 , P2_U4138 , P2_U4139 , P2_U4140;
wire P2_U4141 , P2_U4142 , P2_U4143 , P2_U4144 , P2_U4145 , P2_U4146 , P2_U4147 , P2_U4148 , P2_U4149 , P2_U4150;
wire P2_U4151 , P2_U4152 , P2_U4153 , P2_U4154 , P2_U4155 , P2_U4156 , P2_U4157 , P2_U4158 , P2_U4159 , P2_U4160;
wire P2_U4161 , P2_U4162 , P2_U4163 , P2_U4164 , P2_U4165 , P2_U4166 , P2_U4167 , P2_U4168 , P2_U4169 , P2_U4170;
wire P2_U4171 , P2_U4172 , P2_U4173 , P2_U4174 , P2_U4175 , P2_U4176 , P2_U4177 , P2_U4178 , P2_U4179 , P2_U4180;
wire P2_U4181 , P2_U4182 , P2_U4183 , P2_U4184 , P2_U4185 , P2_U4186 , P2_U4187 , P2_U4188 , P2_U4189 , P2_U4190;
wire P2_U4191 , P2_U4192 , P2_U4193 , P2_U4194 , P2_U4195 , P2_U4196 , P2_U4197 , P2_U4198 , P2_U4199 , P2_U4200;
wire P2_U4201 , P2_U4202 , P2_U4203 , P2_U4204 , P2_U4205 , P2_U4206 , P2_U4207 , P2_U4208 , P2_U4209 , P2_U4210;
wire P2_U4211 , P2_U4212 , P2_U4213 , P2_U4214 , P2_U4215 , P2_U4216 , P2_U4217 , P2_U4218 , P2_U4219 , P2_U4220;
wire P2_U4221 , P2_U4222 , P2_U4223 , P2_U4224 , P2_U4225 , P2_U4226 , P2_U4227 , P2_U4228 , P2_U4229 , P2_U4230;
wire P2_U4231 , P2_U4232 , P2_U4233 , P2_U4234 , P2_U4235 , P2_U4236 , P2_U4237 , P2_U4238 , P2_U4239 , P2_U4240;
wire P2_U4241 , P2_U4242 , P2_U4243 , P2_U4244 , P2_U4245 , P2_U4246 , P2_U4247 , P2_U4248 , P2_U4249 , P2_U4250;
wire P2_U4251 , P2_U4252 , P2_U4253 , P2_U4254 , P2_U4255 , P2_U4256 , P2_U4257 , P2_U4258 , P2_U4259 , P2_U4260;
wire P2_U4261 , P2_U4262 , P2_U4263 , P2_U4264 , P2_U4265 , P2_U4266 , P2_U4267 , P2_U4268 , P2_U4269 , P2_U4270;
wire P2_U4271 , P2_U4272 , P2_U4273 , P2_U4274 , P2_U4275 , P2_U4276 , P2_U4277 , P2_U4278 , P2_U4279 , P2_U4280;
wire P2_U4281 , P2_U4282 , P2_U4283 , P2_U4284 , P2_U4285 , P2_U4286 , P2_U4287 , P2_U4288 , P2_U4289 , P2_U4290;
wire P2_U4291 , P2_U4292 , P2_U4293 , P2_U4294 , P2_U4295 , P2_U4296 , P2_U4297 , P2_U4298 , P2_U4299 , P2_U4300;
wire P2_U4301 , P2_U4302 , P2_U4303 , P2_U4304 , P2_U4305 , P2_U4306 , P2_U4307 , P2_U4308 , P2_U4309 , P2_U4310;
wire P2_U4311 , P2_U4312 , P2_U4313 , P2_U4314 , P2_U4315 , P2_U4316 , P2_U4317 , P2_U4318 , P2_U4319 , P2_U4320;
wire P2_U4321 , P2_U4322 , P2_U4323 , P2_U4324 , P2_U4325 , P2_U4326 , P2_U4327 , P2_U4328 , P2_U4329 , P2_U4330;
wire P2_U4331 , P2_U4332 , P2_U4333 , P2_U4334 , P2_U4335 , P2_U4336 , P2_U4337 , P2_U4338 , P2_U4339 , P2_U4340;
wire P2_U4341 , P2_U4342 , P2_U4343 , P2_U4344 , P2_U4345 , P2_U4346 , P2_U4347 , P2_U4348 , P2_U4349 , P2_U4350;
wire P2_U4351 , P2_U4352 , P2_U4353 , P2_U4354 , P2_U4355 , P2_U4356 , P2_U4357 , P2_U4358 , P2_U4359 , P2_U4360;
wire P2_U4361 , P2_U4362 , P2_U4363 , P2_U4364 , P2_U4365 , P2_U4366 , P2_U4367 , P2_U4368 , P2_U4369 , P2_U4370;
wire P2_U4371 , P2_U4372 , P2_U4373 , P2_U4374 , P2_U4375 , P2_U4376 , P2_U4377 , P2_U4378 , P2_U4379 , P2_U4380;
wire P2_U4381 , P2_U4382 , P2_U4383 , P2_U4384 , P2_U4385 , P2_U4386 , P2_U4387 , P2_U4388 , P2_U4389 , P2_U4390;
wire P2_U4391 , P2_U4392 , P2_U4393 , P2_U4394 , P2_U4395 , P2_U4396 , P2_U4397 , P2_U4398 , P2_U4399 , P2_U4400;
wire P2_U4401 , P2_U4402 , P2_U4403 , P2_U4404 , P2_U4405 , P2_U4406 , P2_U4407 , P2_U4408 , P2_U4409 , P2_U4410;
wire P2_U4411 , P2_U4412 , P2_U4413 , P2_U4414 , P2_U4415 , P2_U4416 , P2_U4417 , P2_U4418 , P2_U4419 , P2_U4420;
wire P2_U4421 , P2_U4422 , P2_U4423 , P2_U4424 , P2_U4425 , P2_U4426 , P2_U4427 , P2_U4428 , P2_U4429 , P2_U4430;
wire P2_U4431 , P2_U4432 , P2_U4433 , P2_U4434 , P2_U4435 , P2_U4436 , P2_U4437 , P2_U4438 , P2_U4439 , P2_U4440;
wire P2_U4441 , P2_U4442 , P2_U4443 , P2_U4444 , P2_U4445 , P2_U4446 , P2_U4447 , P2_U4448 , P2_U4449 , P2_U4450;
wire P2_U4451 , P2_U4452 , P2_U4453 , P2_U4454 , P2_U4455 , P2_U4456 , P2_U4457 , P2_U4458 , P2_U4459 , P2_U4460;
wire P2_U4461 , P2_U4462 , P2_U4463 , P2_U4464 , P2_U4465 , P2_U4466 , P2_U4467 , P2_U4468 , P2_U4469 , P2_U4470;
wire P2_U4471 , P2_U4472 , P2_U4473 , P2_U4474 , P2_U4475 , P2_U4476 , P2_U4477 , P2_U4478 , P2_U4479 , P2_U4480;
wire P2_U4481 , P2_U4482 , P2_U4483 , P2_U4484 , P2_U4485 , P2_U4486 , P2_U4487 , P2_U4488 , P2_U4489 , P2_U4490;
wire P2_U4491 , P2_U4492 , P2_U4493 , P2_U4494 , P2_U4495 , P2_U4496 , P2_U4497 , P2_U4498 , P2_U4499 , P2_U4500;
wire P2_U4501 , P2_U4502 , P2_U4503 , P2_U4504 , P2_U4505 , P2_U4506 , P2_U4507 , P2_U4508 , P2_U4509 , P2_U4510;
wire P2_U4511 , P2_U4512 , P2_U4513 , P2_U4514 , P2_U4515 , P2_U4516 , P2_U4517 , P2_U4518 , P2_U4519 , P2_U4520;
wire P2_U4521 , P2_U4522 , P2_U4523 , P2_U4524 , P2_U4525 , P2_U4526 , P2_U4527 , P2_U4528 , P2_U4529 , P2_U4530;
wire P2_U4531 , P2_U4532 , P2_U4533 , P2_U4534 , P2_U4535 , P2_U4536 , P2_U4537 , P2_U4538 , P2_U4539 , P2_U4540;
wire P2_U4541 , P2_U4542 , P2_U4543 , P2_U4544 , P2_U4545 , P2_U4546 , P2_U4547 , P2_U4548 , P2_U4549 , P2_U4550;
wire P2_U4551 , P2_U4552 , P2_U4553 , P2_U4554 , P2_U4555 , P2_U4556 , P2_U4557 , P2_U4558 , P2_U4559 , P2_U4560;
wire P2_U4561 , P2_U4562 , P2_U4563 , P2_U4564 , P2_U4565 , P2_U4566 , P2_U4567 , P2_U4568 , P2_U4569 , P2_U4570;
wire P2_U4571 , P2_U4572 , P2_U4573 , P2_U4574 , P2_U4575 , P2_U4576 , P2_U4577 , P2_U4578 , P2_U4579 , P2_U4580;
wire P2_U4581 , P2_U4582 , P2_U4583 , P2_U4584 , P2_U4585 , P2_U4586 , P2_U4587 , P2_U4588 , P2_U4589 , P2_U4590;
wire P2_U4591 , P2_U4592 , P2_U4593 , P2_U4594 , P2_U4595 , P2_U4596 , P2_U4597 , P2_U4598 , P2_U4599 , P2_U4600;
wire P2_U4601 , P2_U4602 , P2_U4603 , P2_U4604 , P2_U4605 , P2_U4606 , P2_U4607 , P2_U4608 , P2_U4609 , P2_U4610;
wire P2_U4611 , P2_U4612 , P2_U4613 , P2_U4614 , P2_U4615 , P2_U4616 , P2_U4617 , P2_U4618 , P2_U4619 , P2_U4620;
wire P2_U4621 , P2_U4622 , P2_U4623 , P2_U4624 , P2_U4625 , P2_U4626 , P2_U4627 , P2_U4628 , P2_U4629 , P2_U4630;
wire P2_U4631 , P2_U4632 , P2_U4633 , P2_U4634 , P2_U4635 , P2_U4636 , P2_U4637 , P2_U4638 , P2_U4639 , P2_U4640;
wire P2_U4641 , P2_U4642 , P2_U4643 , P2_U4644 , P2_U4645 , P2_U4646 , P2_U4647 , P2_U4648 , P2_U4649 , P2_U4650;
wire P2_U4651 , P2_U4652 , P2_U4653 , P2_U4654 , P2_U4655 , P2_U4656 , P2_U4657 , P2_U4658 , P2_U4659 , P2_U4660;
wire P2_U4661 , P2_U4662 , P2_U4663 , P2_U4664 , P2_U4665 , P2_U4666 , P2_U4667 , P2_U4668 , P2_U4669 , P2_U4670;
wire P2_U4671 , P2_U4672 , P2_U4673 , P2_U4674 , P2_U4675 , P2_U4676 , P2_U4677 , P2_U4678 , P2_U4679 , P2_U4680;
wire P2_U4681 , P2_U4682 , P2_U4683 , P2_U4684 , P2_U4685 , P2_U4686 , P2_U4687 , P2_U4688 , P2_U4689 , P2_U4690;
wire P2_U4691 , P2_U4692 , P2_U4693 , P2_U4694 , P2_U4695 , P2_U4696 , P2_U4697 , P2_U4698 , P2_U4699 , P2_U4700;
wire P2_U4701 , P2_U4702 , P2_U4703 , P2_U4704 , P2_U4705 , P2_U4706 , P2_U4707 , P2_U4708 , P2_U4709 , P2_U4710;
wire P2_U4711 , P2_U4712 , P2_U4713 , P2_U4714 , P2_U4715 , P2_U4716 , P2_U4717 , P2_U4718 , P2_U4719 , P2_U4720;
wire P2_U4721 , P2_U4722 , P2_U4723 , P2_U4724 , P2_U4725 , P2_U4726 , P2_U4727 , P2_U4728 , P2_U4729 , P2_U4730;
wire P2_U4731 , P2_U4732 , P2_U4733 , P2_U4734 , P2_U4735 , P2_U4736 , P2_U4737 , P2_U4738 , P2_U4739 , P2_U4740;
wire P2_U4741 , P2_U4742 , P2_U4743 , P2_U4744 , P2_U4745 , P2_U4746 , P2_U4747 , P2_U4748 , P2_U4749 , P2_U4750;
wire P2_U4751 , P2_U4752 , P2_U4753 , P2_U4754 , P2_U4755 , P2_U4756 , P2_U4757 , P2_U4758 , P2_U4759 , P2_U4760;
wire P2_U4761 , P2_U4762 , P2_U4763 , P2_U4764 , P2_U4765 , P2_U4766 , P2_U4767 , P2_U4768 , P2_U4769 , P2_U4770;
wire P2_U4771 , P2_U4772 , P2_U4773 , P2_U4774 , P2_U4775 , P2_U4776 , P2_U4777 , P2_U4778 , P2_U4779 , P2_U4780;
wire P2_U4781 , P2_U4782 , P2_U4783 , P2_U4784 , P2_U4785 , P2_U4786 , P2_U4787 , P2_U4788 , P2_U4789 , P2_U4790;
wire P2_U4791 , P2_U4792 , P2_U4793 , P2_U4794 , P2_U4795 , P2_U4796 , P2_U4797 , P2_U4798 , P2_U4799 , P2_U4800;
wire P2_U4801 , P2_U4802 , P2_U4803 , P2_U4804 , P2_U4805 , P2_U4806 , P2_U4807 , P2_U4808 , P2_U4809 , P2_U4810;
wire P2_U4811 , P2_U4812 , P2_U4813 , P2_U4814 , P2_U4815 , P2_U4816 , P2_U4817 , P2_U4818 , P2_U4819 , P2_U4820;
wire P2_U4821 , P2_U4822 , P2_U4823 , P2_U4824 , P2_U4825 , P2_U4826 , P2_U4827 , P2_U4828 , P2_U4829 , P2_U4830;
wire P2_U4831 , P2_U4832 , P2_U4833 , P2_U4834 , P2_U4835 , P2_U4836 , P2_U4837 , P2_U4838 , P2_U4839 , P2_U4840;
wire P2_U4841 , P2_U4842 , P2_U4843 , P2_U4844 , P2_U4845 , P2_U4846 , P2_U4847 , P2_U4848 , P2_U4849 , P2_U4850;
wire P2_U4851 , P2_U4852 , P2_U4853 , P2_U4854 , P2_U4855 , P2_U4856 , P2_U4857 , P2_U4858 , P2_U4859 , P2_U4860;
wire P2_U4861 , P2_U4862 , P2_U4863 , P2_U4864 , P2_U4865 , P2_U4866 , P2_U4867 , P2_U4868 , P2_U4869 , P2_U4870;
wire P2_U4871 , P2_U4872 , P2_U4873 , P2_U4874 , P2_U4875 , P2_U4876 , P2_U4877 , P2_U4878 , P2_U4879 , P2_U4880;
wire P2_U4881 , P2_U4882 , P2_U4883 , P2_U4884 , P2_U4885 , P2_U4886 , P2_U4887 , P2_U4888 , P2_U4889 , P2_U4890;
wire P2_U4891 , P2_U4892 , P2_U4893 , P2_U4894 , P2_U4895 , P2_U4896 , P2_U4897 , P2_U4898 , P2_U4899 , P2_U4900;
wire P2_U4901 , P2_U4902 , P2_U4903 , P2_U4904 , P2_U4905 , P2_U4906 , P2_U4907 , P2_U4908 , P2_U4909 , P2_U4910;
wire P2_U4911 , P2_U4912 , P2_U4913 , P2_U4914 , P2_U4915 , P2_U4916 , P2_U4917 , P2_U4918 , P2_U4919 , P2_U4920;
wire P2_U4921 , P2_U4922 , P2_U4923 , P2_U4924 , P2_U4925 , P2_U4926 , P2_U4927 , P2_U4928 , P2_U4929 , P2_U4930;
wire P2_U4931 , P2_U4932 , P2_U4933 , P2_U4934 , P2_U4935 , P2_U4936 , P2_U4937 , P2_U4938 , P2_U4939 , P2_U4940;
wire P2_U4941 , P2_U4942 , P2_U4943 , P2_U4944 , P2_U4945 , P2_U4946 , P2_U4947 , P2_U4948 , P2_U4949 , P2_U4950;
wire P2_U4951 , P2_U4952 , P2_U4953 , P2_U4954 , P2_U4955 , P2_U4956 , P2_U4957 , P2_U4958 , P2_U4959 , P2_U4960;
wire P2_U4961 , P2_U4962 , P2_U4963 , P2_U4964 , P2_U4965 , P2_U4966 , P2_U4967 , P2_U4968 , P2_U4969 , P2_U4970;
wire P2_U4971 , P2_U4972 , P2_U4973 , P2_U4974 , P2_U4975 , P2_U4976 , P2_U4977 , P2_U4978 , P2_U4979 , P2_U4980;
wire P2_U4981 , P2_U4982 , P2_U4983 , P2_U4984 , P2_U4985 , P2_U4986 , P2_U4987 , P2_U4988 , P2_U4989 , P2_U4990;
wire P2_U4991 , P2_U4992 , P2_U4993 , P2_U4994 , P2_U4995 , P2_U4996 , P2_U4997 , P2_U4998 , P2_U4999 , P2_U5000;
wire P2_U5001 , P2_U5002 , P2_U5003 , P2_U5004 , P2_U5005 , P2_U5006 , P2_U5007 , P2_U5008 , P2_U5009 , P2_U5010;
wire P2_U5011 , P2_U5012 , P2_U5013 , P2_U5014 , P2_U5015 , P2_U5016 , P2_U5017 , P2_U5018 , P2_U5019 , P2_U5020;
wire P2_U5021 , P2_U5022 , P2_U5023 , P2_U5024 , P2_U5025 , P2_U5026 , P2_U5027 , P2_U5028 , P2_U5029 , P2_U5030;
wire P2_U5031 , P2_U5032 , P2_U5033 , P2_U5034 , P2_U5035 , P2_U5036 , P2_U5037 , P2_U5038 , P2_U5039 , P2_U5040;
wire P2_U5041 , P2_U5042 , P2_U5043 , P2_U5044 , P2_U5045 , P2_U5046 , P2_U5047 , P2_U5048 , P2_U5049 , P2_U5050;
wire P2_U5051 , P2_U5052 , P2_U5053 , P2_U5054 , P2_U5055 , P2_U5056 , P2_U5057 , P2_U5058 , P2_U5059 , P2_U5060;
wire P2_U5061 , P2_U5062 , P2_U5063 , P2_U5064 , P2_U5065 , P2_U5066 , P2_U5067 , P2_U5068 , P2_U5069 , P2_U5070;
wire P2_U5071 , P2_U5072 , P2_U5073 , P2_U5074 , P2_U5075 , P2_U5076 , P2_U5077 , P2_U5078 , P2_U5079 , P2_U5080;
wire P2_U5081 , P2_U5082 , P2_U5083 , P2_U5084 , P2_U5085 , P2_U5086 , P2_U5087 , P2_U5088 , P2_U5089 , P2_U5090;
wire P2_U5091 , P2_U5092 , P2_U5093 , P2_U5094 , P2_U5095 , P2_U5096 , P2_U5097 , P2_U5098 , P2_U5099 , P2_U5100;
wire P2_U5101 , P2_U5102 , P2_U5103 , P2_U5104 , P2_U5105 , P2_U5106 , P2_U5107 , P2_U5108 , P2_U5109 , P2_U5110;
wire P2_U5111 , P2_U5112 , P2_U5113 , P2_U5114 , P2_U5115 , P2_U5116 , P2_U5117 , P2_U5118 , P2_U5119 , P2_U5120;
wire P2_U5121 , P2_U5122 , P2_U5123 , P2_U5124 , P2_U5125 , P2_U5126 , P2_U5127 , P2_U5128 , P2_U5129 , P2_U5130;
wire P2_U5131 , P2_U5132 , P2_U5133 , P2_U5134 , P2_U5135 , P2_U5136 , P2_U5137 , P2_U5138 , P2_U5139 , P2_U5140;
wire P2_U5141 , P2_U5142 , P2_U5143 , P2_U5144 , P2_U5145 , P2_U5146 , P2_U5147 , P2_U5148 , P2_U5149 , P2_U5150;
wire P2_U5151 , P2_U5152 , P2_U5153 , P2_U5154 , P2_U5155 , P2_U5156 , P2_U5157 , P2_U5158 , P2_U5159 , P2_U5160;
wire P2_U5161 , P2_U5162 , P2_U5163 , P2_U5164 , P2_U5165 , P2_U5166 , P2_U5167 , P2_U5168 , P2_U5169 , P2_U5170;
wire P2_U5171 , P2_U5172 , P2_U5173 , P2_U5174 , P2_U5175 , P2_U5176 , P2_U5177 , P2_U5178 , P2_U5179 , P2_U5180;
wire P2_U5181 , P2_U5182 , P2_U5183 , P2_U5184 , P2_U5185 , P2_U5186 , P2_U5187 , P2_U5188 , P2_U5189 , P2_U5190;
wire P2_U5191 , P2_U5192 , P2_U5193 , P2_U5194 , P2_U5195 , P2_U5196 , P2_U5197 , P2_U5198 , P2_U5199 , P2_U5200;
wire P2_U5201 , P2_U5202 , P2_U5203 , P2_U5204 , P2_U5205 , P2_U5206 , P2_U5207 , P2_U5208 , P2_U5209 , P2_U5210;
wire P2_U5211 , P2_U5212 , P2_U5213 , P2_U5214 , P2_U5215 , P2_U5216 , P2_U5217 , P2_U5218 , P2_U5219 , P2_U5220;
wire P2_U5221 , P2_U5222 , P2_U5223 , P2_U5224 , P2_U5225 , P2_U5226 , P2_U5227 , P2_U5228 , P2_U5229 , P2_U5230;
wire P2_U5231 , P2_U5232 , P2_U5233 , P2_U5234 , P2_U5235 , P2_U5236 , P2_U5237 , P2_U5238 , P2_U5239 , P2_U5240;
wire P2_U5241 , P2_U5242 , P2_U5243 , P2_U5244 , P2_U5245 , P2_U5246 , P2_U5247 , P2_U5248 , P2_U5249 , P2_U5250;
wire P2_U5251 , P2_U5252 , P2_U5253 , P2_U5254 , P2_U5255 , P2_U5256 , P2_U5257 , P2_U5258 , P2_U5259 , P2_U5260;
wire P2_U5261 , P2_U5262 , P2_U5263 , P2_U5264 , P2_U5265 , P2_U5266 , P2_U5267 , P2_U5268 , P2_U5269 , P2_U5270;
wire P2_U5271 , P2_U5272 , P2_U5273 , P2_U5274 , P2_U5275 , P2_U5276 , P2_U5277 , P2_U5278 , P2_U5279 , P2_U5280;
wire P2_U5281 , P2_U5282 , P2_U5283 , P2_U5284 , P2_U5285 , P2_U5286 , P2_U5287 , P2_U5288 , P2_U5289 , P2_U5290;
wire P2_U5291 , P2_U5292 , P2_U5293 , P2_U5294 , P2_U5295 , P2_U5296 , P2_U5297 , P2_U5298 , P2_U5299 , P2_U5300;
wire P2_U5301 , P2_U5302 , P2_U5303 , P2_U5304 , P2_U5305 , P2_U5306 , P2_U5307 , P2_U5308 , P2_U5309 , P2_U5310;
wire P2_U5311 , P2_U5312 , P2_U5313 , P2_U5314 , P2_U5315 , P2_U5316 , P2_U5317 , P2_U5318 , P2_U5319 , P2_U5320;
wire P2_U5321 , P2_U5322 , P2_U5323 , P2_U5324 , P2_U5325 , P2_U5326 , P2_U5327 , P2_U5328 , P2_U5329 , P2_U5330;
wire P2_U5331 , P2_U5332 , P2_U5333 , P2_U5334 , P2_U5335 , P2_U5336 , P2_U5337 , P2_U5338 , P2_U5339 , P2_U5340;
wire P2_U5341 , P2_U5342 , P2_U5343 , P2_U5344 , P2_U5345 , P2_U5346 , P2_U5347 , P2_U5348 , P2_U5349 , P2_U5350;
wire P2_U5351 , P2_U5352 , P2_U5353 , P2_U5354 , P2_U5355 , P2_U5356 , P2_U5357 , P2_U5358 , P2_U5359 , P2_U5360;
wire P2_U5361 , P2_U5362 , P2_U5363 , P2_U5364 , P2_U5365 , P2_U5366 , P2_U5367 , P2_U5368 , P2_U5369 , P2_U5370;
wire P2_U5371 , P2_U5372 , P2_U5373 , P2_U5374 , P2_U5375 , P2_U5376 , P2_U5377 , P2_U5378 , P2_U5379 , P2_U5380;
wire P2_U5381 , P2_U5382 , P2_U5383 , P2_U5384 , P2_U5385 , P2_U5386 , P2_U5387 , P2_U5388 , P2_U5389 , P2_U5390;
wire P2_U5391 , P2_U5392 , P2_U5393 , P2_U5394 , P2_U5395 , P2_U5396 , P2_U5397 , P2_U5398 , P2_U5399 , P2_U5400;
wire P2_U5401 , P2_U5402 , P2_U5403 , P2_U5404 , P2_U5405 , P2_U5406 , P2_U5407 , P2_U5408 , P2_U5409 , P2_U5410;
wire P2_U5411 , P2_U5412 , P2_U5413 , P2_U5414 , P2_U5415 , P2_U5416 , P2_U5417 , P2_U5418 , P2_U5419 , P2_U5420;
wire P2_U5421 , P2_U5422 , P2_U5423 , P2_U5424 , P2_U5425 , P2_U5426 , P2_U5427 , P2_U5428 , P2_U5429 , P2_U5430;
wire P2_U5431 , P2_U5432 , P2_U5433 , P2_U5434 , P2_U5435 , P2_U5436 , P2_U5437 , P2_U5438 , P2_U5439 , P2_U5440;
wire P2_U5441 , P2_U5442 , P2_U5443 , P2_U5444 , P2_U5445 , P2_U5446 , P2_U5447 , P2_U5448 , P2_U5449 , P2_U5450;
wire P2_U5451 , P2_U5452 , P2_U5453 , P2_U5454 , P2_U5455 , P2_U5456 , P2_U5457 , P2_U5458 , P2_U5459 , P2_U5460;
wire P2_U5461 , P2_U5462 , P2_U5463 , P2_U5464 , P2_U5465 , P2_U5466 , P2_U5467 , P2_U5468 , P2_U5469 , P2_U5470;
wire P2_U5471 , P2_U5472 , P2_U5473 , P2_U5474 , P2_U5475 , P2_U5476 , P2_U5477 , P2_U5478 , P2_U5479 , P2_U5480;
wire P2_U5481 , P2_U5482 , P2_U5483 , P2_U5484 , P2_U5485 , P2_U5486 , P2_U5487 , P2_U5488 , P2_U5489 , P2_U5490;
wire P2_U5491 , P2_U5492 , P2_U5493 , P2_U5494 , P2_U5495 , P2_U5496 , P2_U5497 , P2_U5498 , P2_U5499 , P2_U5500;
wire P2_U5501 , P2_U5502 , P2_U5503 , P2_U5504 , P2_U5505 , P2_U5506 , P2_U5507 , P2_U5508 , P2_U5509 , P2_U5510;
wire P2_U5511 , P2_U5512 , P2_U5513 , P2_U5514 , P2_U5515 , P2_U5516 , P2_U5517 , P2_U5518 , P2_U5519 , P2_U5520;
wire P2_U5521 , P2_U5522 , P2_U5523 , P2_U5524 , P2_U5525 , P2_U5526 , P2_U5527 , P2_U5528 , P2_U5529 , P2_U5530;
wire P2_U5531 , P2_U5532 , P2_U5533 , P2_U5534 , P2_U5535 , P2_U5536 , P2_U5537 , P2_U5538 , P2_U5539 , P2_U5540;
wire P2_U5541 , P2_U5542 , P2_U5543 , P2_U5544 , P2_U5545 , P2_U5546 , P2_U5547 , P2_U5548 , P2_U5549 , P2_U5550;
wire P2_U5551 , P2_U5552 , P2_U5553 , P2_U5554 , P2_U5555 , P2_U5556 , P2_U5557 , P2_U5558 , P2_U5559 , P2_U5560;
wire P2_U5561 , P2_U5562 , P2_U5563 , P2_U5564 , P2_U5565 , P2_U5566 , P2_U5567 , P2_U5568 , P2_U5569 , P2_U5570;
wire P2_U5571 , P2_U5572 , P2_U5573 , P2_U5574 , P2_U5575 , P2_U5576 , P2_U5577 , P2_U5578 , P2_U5579 , P2_U5580;
wire P2_U5581 , P2_U5582 , P2_U5583 , P2_U5584 , P2_U5585 , P2_U5586 , P2_U5587 , P2_U5588 , P2_U5589 , P2_U5590;
wire P2_U5591 , P2_U5592 , P2_U5593 , P2_U5594 , P2_U5595 , P2_U5596 , P2_U5597 , P2_U5598 , P2_U5599 , P2_U5600;
wire P2_U5601 , P2_U5602 , P2_U5603 , P2_U5604 , P2_U5605 , P2_U5606 , P2_U5607 , P2_U5608 , P2_U5609 , P2_U5610;
wire P2_U5611 , P2_U5612 , P2_U5613 , P2_U5614 , P2_U5615 , P2_U5616 , P2_U5617 , P2_U5618 , P2_U5619 , P2_U5620;
wire P2_U5621 , P2_U5622 , P2_U5623 , P2_U5624 , P2_U5625 , P2_U5626 , P2_U5627 , P2_U5628 , P2_U5629 , P2_U5630;
wire P2_U5631 , P2_U5632 , P2_U5633 , P2_U5634 , P2_U5635 , P2_U5636 , P2_U5637 , P2_U5638 , P2_U5639 , P2_U5640;
wire P2_U5641 , P2_U5642 , P2_U5643 , P2_U5644 , P2_U5645 , P2_U5646 , P2_U5647 , P2_U5648 , P2_U5649 , P2_U5650;
wire P2_U5651 , P2_U5652 , P2_U5653 , P2_U5654 , P2_U5655 , P2_U5656 , P2_U5657 , P2_U5658 , P2_U5659 , P2_U5660;
wire P2_U5661 , P2_U5662 , P2_U5663 , P2_U5664 , P2_U5665 , P2_U5666 , P2_U5667 , P2_U5668 , P2_U5669 , P2_U5670;
wire P2_U5671 , P2_U5672 , P2_U5673 , P2_U5674 , P2_U5675 , P2_U5676 , P2_U5677 , P2_U5678 , P2_U5679 , P2_U5680;
wire P2_U5681 , P2_U5682 , P2_U5683 , P2_U5684 , P2_U5685 , P2_U5686 , P2_U5687 , P2_U5688 , P2_U5689 , P2_U5690;
wire P2_U5691 , P2_U5692 , P2_U5693 , P2_U5694 , P2_U5695 , P2_U5696 , P2_U5697 , P2_U5698 , P2_U5699 , P2_U5700;
wire P2_U5701 , P2_U5702 , P2_U5703 , P2_U5704 , P2_U5705 , P2_U5706 , P2_U5707 , P2_U5708 , P2_U5709 , P2_U5710;
wire P2_U5711 , P2_U5712 , P2_U5713 , P2_U5714 , P2_U5715 , P2_U5716 , P2_U5717 , P2_U5718 , P2_U5719 , P2_U5720;
wire P2_U5721 , P2_U5722 , P2_U5723 , P2_U5724 , P2_U5725 , P2_U5726 , P2_U5727 , P2_U5728 , P2_U5729 , P2_U5730;
wire P2_U5731 , P2_U5732 , P2_U5733 , P2_U5734 , P2_U5735 , P2_U5736 , P2_U5737 , P2_U5738 , P2_U5739 , P2_U5740;
wire P2_U5741 , P2_U5742 , P2_U5743 , P2_U5744 , P2_U5745 , P2_U5746 , P2_U5747 , P2_U5748 , P2_U5749 , P2_U5750;
wire P2_U5751 , P2_U5752 , P2_U5753 , P2_U5754 , P2_U5755 , P2_U5756 , P2_U5757 , P2_U5758 , P2_U5759 , P2_U5760;
wire P2_U5761 , P2_U5762 , P2_U5763 , P2_U5764 , P2_U5765 , P2_U5766 , P2_U5767 , P2_U5768 , P2_U5769 , P2_U5770;
wire P2_U5771 , P2_U5772 , P2_U5773 , P2_U5774 , P2_U5775 , P2_U5776 , P2_U5777 , P2_U5778 , P2_U5779 , P2_U5780;
wire P2_U5781 , P2_U5782 , P2_U5783 , P2_U5784 , P2_U5785 , P2_U5786 , P2_U5787 , P2_U5788 , P2_U5789 , P2_U5790;
wire P2_U5791 , P2_U5792 , P2_U5793 , P2_U5794 , P2_U5795 , P2_U5796 , P2_U5797 , P2_U5798 , P2_U5799 , P2_U5800;
wire P2_U5801 , P2_U5802 , P2_U5803 , P2_U5804 , P2_U5805 , P2_U5806 , P2_U5807 , P2_U5808 , P2_U5809 , P2_U5810;
wire P2_U5811 , P2_U5812 , P2_U5813 , P2_U5814 , P2_U5815 , P2_U5816 , P2_U5817 , P2_U5818 , P2_U5819 , P2_U5820;
wire P2_U5821 , P2_U5822 , P2_U5823 , P2_U5824 , P2_U5825 , P2_U5826 , P2_U5827 , P2_U5828 , P2_U5829 , P2_U5830;
wire P2_U5831 , P2_U5832 , P2_U5833 , P2_U5834 , P2_U5835 , P2_U5836 , P2_U5837 , P2_U5838 , P2_U5839 , P2_U5840;
wire P2_U5841 , P2_U5842 , P2_U5843 , P2_U5844 , P2_U5845 , P2_U5846 , P2_U5847 , P2_U5848 , P2_U5849 , P2_U5850;
wire P2_U5851 , P2_U5852 , P2_U5853 , P2_U5854 , P2_U5855 , P2_U5856 , P2_U5857 , P2_U5858 , P2_U5859 , P2_U5860;
wire P2_U5861 , P2_U5862 , P2_U5863 , P2_U5864 , P2_U5865 , P2_U5866 , P2_U5867 , P2_U5868 , P2_U5869 , P2_U5870;
wire P2_U5871 , P2_U5872 , P2_U5873 , P2_U5874 , P2_U5875 , P2_U5876 , P2_U5877 , P2_U5878 , P2_U5879 , P2_U5880;
wire P2_U5881 , P2_U5882 , P2_U5883 , P2_U5884 , P2_U5885 , P2_U5886 , P2_U5887 , P2_U5888 , P2_U5889 , P2_U5890;
wire P2_U5891 , P2_U5892 , P2_U5893 , P2_U5894 , P2_U5895 , P2_U5896 , P2_U5897 , P2_U5898 , P2_U5899 , P2_U5900;
wire P2_U5901 , P2_U5902 , P2_U5903 , P2_U5904 , P2_U5905 , P2_U5906 , P2_U5907 , P2_U5908 , P2_U5909 , P2_U5910;
wire P2_U5911 , P2_U5912 , P2_U5913 , P2_U5914 , P2_U5915 , P2_U5916 , P2_U5917 , P2_U5918 , P2_U5919 , P2_U5920;
wire P2_U5921 , P2_U5922 , P2_U5923 , P2_U5924 , P2_U5925 , P2_U5926 , P2_U5927 , P2_U5928 , P2_U5929 , P2_U5930;
wire P2_U5931 , P2_U5932 , P2_U5933 , P2_U5934 , P2_U5935 , P2_U5936 , P2_U5937 , P2_U5938 , P2_U5939 , P2_U5940;
wire P2_U5941 , P2_U5942 , P2_U5943 , P2_U5944 , P2_U5945 , P2_U5946 , P2_U5947 , P2_U5948 , P2_U5949 , P2_U5950;
wire P2_U5951 , P2_U5952 , P2_U5953 , P2_U5954 , P2_U5955 , P2_U5956 , P2_U5957 , P2_U5958 , P2_U5959 , P2_U5960;
wire P2_U5961 , P2_U5962 , P2_U5963 , P2_U5964 , P2_U5965 , P2_U5966 , P2_U5967 , P2_U5968 , P2_U5969 , P2_U5970;
wire P2_U5971 , P2_U5972 , P2_U5973 , P2_U5974 , P2_U5975 , P2_U5976 , P2_U5977 , P2_U5978 , P2_U5979 , P2_U5980;
wire P2_U5981 , P2_U5982 , P2_U5983 , P2_U5984 , P2_U5985 , P2_U5986 , P2_U5987 , P2_U5988 , P2_U5989 , P2_U5990;
wire P2_U5991 , P2_U5992 , P2_U5993 , P2_U5994 , P2_U5995 , P2_U5996 , P2_U5997 , P2_U5998 , P2_U5999 , P2_U6000;
wire P2_U6001 , P2_U6002 , P2_U6003 , P2_U6004 , P2_U6005 , P2_U6006 , P2_U6007 , P2_U6008 , P2_U6009 , P2_U6010;
wire P2_U6011 , P2_U6012 , P2_U6013 , P2_U6014 , P2_U6015 , P2_U6016 , P2_U6017 , P2_U6018 , P2_U6019 , P2_U6020;
wire P2_U6021 , P2_U6022 , P2_U6023 , P2_U6024 , P2_U6025 , P2_U6026 , P2_U6027 , P2_U6028 , P2_U6029 , P2_U6030;
wire P2_U6031 , P2_U6032 , P2_U6033 , P2_U6034 , P2_U6035 , P2_U6036 , P2_U6037 , P2_U6038 , P2_U6039 , P2_U6040;
wire P2_U6041 , P2_U6042 , P2_U6043 , P2_U6044 , P2_R1161_U465 , P2_R1161_U464 , P2_R1161_U463 , P2_R1161_U462 , P2_R1161_U461 , P2_R1161_U460;
wire P2_R1161_U459 , P2_R1161_U458 , P2_R1161_U457 , P2_R1161_U456 , P2_R1161_U455 , P2_R1161_U454 , P2_R1161_U453 , P2_R1161_U452 , P2_R1161_U451 , P2_R1161_U450;
wire P2_R1161_U449 , P2_R1161_U448 , P2_R1161_U447 , LT_1075_U6 , ADD_1068_U6 , ADD_1068_U7 , ADD_1068_U8 , ADD_1068_U9 , ADD_1068_U10 , ADD_1068_U11;
wire ADD_1068_U12 , ADD_1068_U13 , ADD_1068_U14 , ADD_1068_U15 , ADD_1068_U16 , ADD_1068_U17 , ADD_1068_U18 , ADD_1068_U19 , ADD_1068_U20 , ADD_1068_U21;
wire ADD_1068_U22 , ADD_1068_U23 , ADD_1068_U24 , ADD_1068_U25 , ADD_1068_U26 , ADD_1068_U27 , ADD_1068_U28 , ADD_1068_U29 , ADD_1068_U30 , ADD_1068_U31;
wire ADD_1068_U32 , ADD_1068_U33 , ADD_1068_U34 , ADD_1068_U35 , ADD_1068_U36 , ADD_1068_U37 , ADD_1068_U38 , ADD_1068_U39 , ADD_1068_U40 , ADD_1068_U41;
wire ADD_1068_U42 , ADD_1068_U43 , ADD_1068_U44 , ADD_1068_U45 , ADD_1068_U64 , ADD_1068_U65 , ADD_1068_U66 , ADD_1068_U67 , ADD_1068_U68 , ADD_1068_U69;
wire ADD_1068_U70 , ADD_1068_U71 , ADD_1068_U72 , ADD_1068_U73 , ADD_1068_U74 , ADD_1068_U75 , ADD_1068_U76 , ADD_1068_U77 , ADD_1068_U78 , ADD_1068_U79;
wire ADD_1068_U80 , ADD_1068_U81 , ADD_1068_U82 , ADD_1068_U83 , ADD_1068_U84 , ADD_1068_U85 , ADD_1068_U86 , ADD_1068_U87 , ADD_1068_U88 , ADD_1068_U89;
wire ADD_1068_U90 , ADD_1068_U91 , ADD_1068_U92 , ADD_1068_U93 , ADD_1068_U94 , ADD_1068_U95 , ADD_1068_U96 , ADD_1068_U97 , ADD_1068_U98 , ADD_1068_U99;
wire ADD_1068_U100 , ADD_1068_U101 , ADD_1068_U102 , ADD_1068_U103 , ADD_1068_U104 , ADD_1068_U105 , ADD_1068_U106 , ADD_1068_U107 , ADD_1068_U108 , ADD_1068_U109;
wire ADD_1068_U110 , ADD_1068_U111 , ADD_1068_U112 , ADD_1068_U113 , ADD_1068_U114 , ADD_1068_U115 , ADD_1068_U116 , ADD_1068_U117 , ADD_1068_U118 , ADD_1068_U119;
wire ADD_1068_U120 , ADD_1068_U121 , ADD_1068_U122 , ADD_1068_U123 , ADD_1068_U124 , ADD_1068_U125 , ADD_1068_U126 , ADD_1068_U127 , ADD_1068_U128 , ADD_1068_U129;
wire ADD_1068_U130 , ADD_1068_U131 , ADD_1068_U132 , ADD_1068_U133 , ADD_1068_U134 , ADD_1068_U135 , ADD_1068_U136 , ADD_1068_U137 , ADD_1068_U138 , ADD_1068_U139;
wire ADD_1068_U140 , ADD_1068_U141 , ADD_1068_U142 , ADD_1068_U143 , ADD_1068_U144 , ADD_1068_U145 , ADD_1068_U146 , ADD_1068_U147 , ADD_1068_U148 , ADD_1068_U149;
wire ADD_1068_U150 , ADD_1068_U151 , ADD_1068_U152 , ADD_1068_U153 , ADD_1068_U154 , ADD_1068_U155 , ADD_1068_U156 , ADD_1068_U157 , ADD_1068_U158 , ADD_1068_U159;
wire ADD_1068_U160 , ADD_1068_U161 , ADD_1068_U162 , ADD_1068_U163 , ADD_1068_U164 , ADD_1068_U165 , ADD_1068_U166 , ADD_1068_U167 , ADD_1068_U168 , ADD_1068_U169;
wire ADD_1068_U170 , ADD_1068_U171 , ADD_1068_U172 , ADD_1068_U173 , ADD_1068_U174 , ADD_1068_U175 , ADD_1068_U176 , ADD_1068_U177 , ADD_1068_U178 , ADD_1068_U179;
wire ADD_1068_U180 , ADD_1068_U181 , ADD_1068_U182 , ADD_1068_U183 , ADD_1068_U184 , ADD_1068_U185 , ADD_1068_U186 , ADD_1068_U187 , ADD_1068_U188 , ADD_1068_U189;
wire ADD_1068_U190 , ADD_1068_U191 , ADD_1068_U192 , ADD_1068_U193 , ADD_1068_U194 , ADD_1068_U195 , ADD_1068_U196 , ADD_1068_U197 , ADD_1068_U198 , ADD_1068_U199;
wire ADD_1068_U200 , ADD_1068_U201 , ADD_1068_U202 , ADD_1068_U203 , ADD_1068_U204 , ADD_1068_U205 , ADD_1068_U206 , ADD_1068_U207 , ADD_1068_U208 , ADD_1068_U209;
wire ADD_1068_U210 , ADD_1068_U211 , ADD_1068_U212 , ADD_1068_U213 , ADD_1068_U214 , ADD_1068_U215 , ADD_1068_U216 , ADD_1068_U217 , ADD_1068_U218 , ADD_1068_U219;
wire ADD_1068_U220 , ADD_1068_U221 , ADD_1068_U222 , ADD_1068_U223 , ADD_1068_U224 , ADD_1068_U225 , ADD_1068_U226 , ADD_1068_U227 , ADD_1068_U228 , ADD_1068_U229;
wire ADD_1068_U230 , ADD_1068_U231 , ADD_1068_U232 , ADD_1068_U233 , ADD_1068_U234 , ADD_1068_U235 , ADD_1068_U236 , ADD_1068_U237 , ADD_1068_U238 , ADD_1068_U239;
wire ADD_1068_U240 , ADD_1068_U241 , ADD_1068_U242 , ADD_1068_U243 , ADD_1068_U244 , ADD_1068_U245 , ADD_1068_U246 , ADD_1068_U247 , ADD_1068_U248 , ADD_1068_U249;
wire ADD_1068_U250 , ADD_1068_U251 , ADD_1068_U252 , ADD_1068_U253 , ADD_1068_U254 , ADD_1068_U255 , ADD_1068_U256 , ADD_1068_U257 , ADD_1068_U258 , ADD_1068_U259;
wire ADD_1068_U260 , ADD_1068_U261 , ADD_1068_U262 , ADD_1068_U263 , ADD_1068_U264 , ADD_1068_U265 , ADD_1068_U266 , ADD_1068_U267 , ADD_1068_U268 , ADD_1068_U269;
wire ADD_1068_U270 , ADD_1068_U271 , ADD_1068_U272 , ADD_1068_U273 , ADD_1068_U274 , ADD_1068_U275 , ADD_1068_U276 , ADD_1068_U277 , ADD_1068_U278 , ADD_1068_U279;
wire ADD_1068_U280 , ADD_1068_U281 , ADD_1068_U282 , ADD_1068_U283 , ADD_1068_U284 , ADD_1068_U285 , ADD_1068_U286 , ADD_1068_U287 , ADD_1068_U288 , ADD_1068_U289;
wire ADD_1068_U290 , ADD_1068_U291 , R140_U4 , R140_U5 , R140_U6 , R140_U7 , R140_U8 , R140_U9 , R140_U10 , R140_U11;
wire R140_U12 , R140_U13 , R140_U14 , R140_U15 , R140_U16 , R140_U17 , R140_U18 , R140_U19 , R140_U20 , R140_U21;
wire R140_U22 , R140_U23 , R140_U24 , R140_U25 , R140_U26 , R140_U27 , R140_U28 , R140_U29 , R140_U30 , R140_U31;
wire R140_U32 , R140_U33 , R140_U34 , R140_U35 , R140_U36 , R140_U37 , R140_U38 , R140_U39 , R140_U40 , R140_U41;
wire R140_U42 , R140_U43 , R140_U44 , R140_U45 , R140_U46 , R140_U47 , R140_U48 , R140_U49 , R140_U50 , R140_U51;
wire R140_U52 , R140_U53 , R140_U54 , R140_U55 , R140_U56 , R140_U57 , R140_U58 , R140_U59 , R140_U60 , R140_U61;
wire R140_U62 , R140_U63 , R140_U64 , R140_U65 , R140_U66 , R140_U67 , R140_U68 , R140_U69 , R140_U70 , R140_U71;
wire R140_U72 , R140_U73 , R140_U74 , R140_U75 , R140_U76 , R140_U77 , R140_U78 , R140_U79 , R140_U80 , R140_U81;
wire R140_U82 , R140_U83 , R140_U84 , R140_U85 , R140_U86 , R140_U87 , R140_U88 , R140_U89 , R140_U90 , R140_U91;
wire R140_U92 , R140_U93 , R140_U94 , R140_U95 , R140_U96 , R140_U97 , R140_U98 , R140_U99 , R140_U100 , R140_U101;
wire R140_U102 , R140_U103 , R140_U104 , R140_U105 , R140_U106 , R140_U107 , R140_U108 , R140_U109 , R140_U110 , R140_U111;
wire R140_U112 , R140_U113 , R140_U114 , R140_U115 , R140_U116 , R140_U117 , R140_U118 , R140_U119 , R140_U120 , R140_U121;
wire R140_U122 , R140_U123 , R140_U124 , R140_U125 , R140_U126 , R140_U127 , R140_U128 , R140_U129 , R140_U130 , R140_U131;
wire R140_U132 , R140_U133 , R140_U134 , R140_U135 , R140_U136 , R140_U137 , R140_U138 , R140_U139 , R140_U140 , R140_U141;
wire R140_U142 , R140_U143 , R140_U144 , R140_U145 , R140_U146 , R140_U147 , R140_U148 , R140_U149 , R140_U150 , R140_U151;
wire R140_U152 , R140_U153 , R140_U154 , R140_U155 , R140_U156 , R140_U157 , R140_U158 , R140_U159 , R140_U160 , R140_U161;
wire R140_U162 , R140_U163 , R140_U164 , R140_U165 , R140_U166 , R140_U167 , R140_U168 , R140_U169 , R140_U170 , R140_U171;
wire R140_U172 , R140_U173 , R140_U174 , R140_U175 , R140_U176 , R140_U177 , R140_U178 , R140_U179 , R140_U180 , R140_U181;
wire R140_U182 , R140_U183 , R140_U184 , R140_U185 , R140_U186 , R140_U187 , R140_U188 , R140_U189 , R140_U190 , R140_U191;
wire R140_U192 , R140_U193 , R140_U194 , R140_U195 , R140_U196 , R140_U197 , R140_U198 , R140_U199 , R140_U200 , R140_U201;
wire R140_U202 , R140_U203 , R140_U204 , R140_U205 , R140_U206 , R140_U207 , R140_U208 , R140_U209 , R140_U210 , R140_U211;
wire R140_U212 , R140_U213 , R140_U214 , R140_U215 , R140_U216 , R140_U217 , R140_U218 , R140_U219 , R140_U220 , R140_U221;
wire R140_U222 , R140_U223 , R140_U224 , R140_U225 , R140_U226 , R140_U227 , R140_U228 , R140_U229 , R140_U230 , R140_U231;
wire R140_U232 , R140_U233 , R140_U234 , R140_U235 , R140_U236 , R140_U237 , R140_U238 , R140_U239 , R140_U240 , R140_U241;
wire R140_U242 , R140_U243 , R140_U244 , R140_U245 , R140_U246 , R140_U247 , R140_U248 , R140_U249 , R140_U250 , R140_U251;
wire R140_U252 , R140_U253 , R140_U254 , R140_U255 , R140_U256 , R140_U257 , R140_U258 , R140_U259 , R140_U260 , R140_U261;
wire R140_U262 , R140_U263 , R140_U264 , R140_U265 , R140_U266 , R140_U267 , R140_U268 , R140_U269 , R140_U270 , R140_U271;
wire R140_U272 , R140_U273 , R140_U274 , R140_U275 , R140_U276 , R140_U277 , R140_U278 , R140_U279 , R140_U280 , R140_U281;
wire R140_U282 , R140_U283 , R140_U284 , R140_U285 , R140_U286 , R140_U287 , R140_U288 , R140_U289 , R140_U290 , R140_U291;
wire R140_U292 , R140_U293 , R140_U294 , R140_U295 , R140_U296 , R140_U297 , R140_U298 , R140_U299 , R140_U300 , R140_U301;
wire R140_U302 , R140_U303 , R140_U304 , R140_U305 , R140_U306 , R140_U307 , R140_U308 , R140_U309 , R140_U310 , R140_U311;
wire R140_U312 , R140_U313 , R140_U314 , R140_U315 , R140_U316 , R140_U317 , R140_U318 , R140_U319 , R140_U320 , R140_U321;
wire R140_U322 , R140_U323 , R140_U324 , R140_U325 , R140_U326 , R140_U327 , R140_U328 , R140_U329 , R140_U330 , R140_U331;
wire R140_U332 , R140_U333 , R140_U334 , R140_U335 , R140_U336 , R140_U337 , R140_U338 , R140_U339 , R140_U340 , R140_U341;
wire R140_U342 , R140_U343 , R140_U344 , R140_U345 , R140_U346 , R140_U347 , R140_U348 , R140_U349 , R140_U350 , R140_U351;
wire R140_U352 , R140_U353 , R140_U354 , R140_U355 , R140_U356 , R140_U357 , R140_U358 , R140_U359 , R140_U360 , R140_U361;
wire R140_U362 , R140_U363 , R140_U364 , R140_U365 , R140_U366 , R140_U367 , R140_U368 , R140_U369 , R140_U370 , R140_U371;
wire R140_U372 , R140_U373 , R140_U374 , R140_U375 , R140_U376 , R140_U377 , R140_U378 , R140_U379 , R140_U380 , R140_U381;
wire R140_U382 , R140_U383 , R140_U384 , R140_U385 , R140_U386 , R140_U387 , R140_U388 , R140_U389 , R140_U390 , R140_U391;
wire R140_U392 , R140_U393 , R140_U394 , R140_U395 , R140_U396 , R140_U397 , R140_U398 , R140_U399 , R140_U400 , R140_U401;
wire R140_U402 , R140_U403 , R140_U404 , R140_U405 , R140_U406 , R140_U407 , R140_U408 , R140_U409 , R140_U410 , R140_U411;
wire R140_U412 , R140_U413 , R140_U414 , R140_U415 , R140_U416 , R140_U417 , R140_U418 , R140_U419 , R140_U420 , R140_U421;
wire R140_U422 , R140_U423 , R140_U424 , R140_U425 , R140_U426 , R140_U427 , R140_U428 , R140_U429 , R140_U430 , R140_U431;
wire R140_U432 , R140_U433 , R140_U434 , R140_U435 , R140_U436 , R140_U437 , R140_U438 , R140_U439 , R140_U440 , R140_U441;
wire R140_U442 , R140_U443 , R140_U444 , R140_U445 , R140_U446 , R140_U447 , R140_U448 , R140_U449 , R140_U450 , R140_U451;
wire R140_U452 , R140_U453 , R140_U454 , R140_U455 , R140_U456 , R140_U457 , R140_U458 , R140_U459 , R140_U460 , R140_U461;
wire R140_U462 , R140_U463 , R140_U464 , R140_U465 , R140_U466 , R140_U467 , R140_U468 , R140_U469 , R140_U470 , R140_U471;
wire R140_U472 , R140_U473 , R140_U474 , R140_U475 , R140_U476 , R140_U477 , R140_U478 , R140_U479 , R140_U480 , R140_U481;
wire R140_U482 , R140_U483 , R140_U484 , R140_U485 , R140_U486 , R140_U487 , R140_U488 , R140_U489 , R140_U490 , R140_U491;
wire R140_U492 , R140_U493 , R140_U494 , R140_U495 , R140_U496 , R140_U497 , R140_U498 , R140_U499 , R140_U500 , R140_U501;
wire R140_U502 , R140_U503 , R140_U504 , R140_U505 , R140_U506 , R140_U507 , R140_U508 , R140_U509 , R140_U510 , R140_U511;
wire R140_U512 , R140_U513 , R140_U514 , R140_U515 , R140_U516 , R140_U517 , R140_U518 , R140_U519 , R140_U520 , R140_U521;
wire R140_U522 , R140_U523 , R140_U524 , R140_U525 , R140_U526 , R140_U527 , R140_U528 , R140_U529 , R140_U530 , R140_U531;
wire R140_U532 , R140_U533 , R140_U534 , R140_U535 , R140_U536 , R140_U537 , R140_U538 , R140_U539 , R140_U540 , R140_U541;
wire LT_1075_19_U6 , P1_ADD_95_U4 , P1_ADD_95_U5 , P1_ADD_95_U6 , P1_ADD_95_U7 , P1_ADD_95_U8 , P1_ADD_95_U9 , P1_ADD_95_U10 , P1_ADD_95_U11 , P1_ADD_95_U12;
wire P1_ADD_95_U13 , P1_ADD_95_U14 , P1_ADD_95_U15 , P1_ADD_95_U16 , P1_ADD_95_U17 , P1_ADD_95_U18 , P1_ADD_95_U19 , P1_ADD_95_U20 , P1_ADD_95_U21 , P1_ADD_95_U22;
wire P1_ADD_95_U23 , P1_ADD_95_U24 , P1_ADD_95_U25 , P1_ADD_95_U26 , P1_ADD_95_U27 , P1_ADD_95_U28 , P1_ADD_95_U29 , P1_ADD_95_U30 , P1_ADD_95_U31 , P1_ADD_95_U32;
wire P1_ADD_95_U33 , P1_ADD_95_U34 , P1_ADD_95_U35 , P1_ADD_95_U36 , P1_ADD_95_U37 , P1_ADD_95_U38 , P1_ADD_95_U39 , P1_ADD_95_U40 , P1_ADD_95_U41 , P1_ADD_95_U42;
wire P1_ADD_95_U43 , P1_ADD_95_U44 , P1_ADD_95_U45 , P1_ADD_95_U46 , P1_ADD_95_U47 , P1_ADD_95_U48 , P1_ADD_95_U49 , P1_ADD_95_U50 , P1_ADD_95_U51 , P1_ADD_95_U52;
wire P1_ADD_95_U53 , P1_ADD_95_U54 , P1_ADD_95_U55 , P1_ADD_95_U56 , P1_ADD_95_U57 , P1_ADD_95_U58 , P1_ADD_95_U59 , P1_ADD_95_U60 , P1_ADD_95_U61 , P1_ADD_95_U62;
wire P1_ADD_95_U63 , P1_ADD_95_U64 , P1_ADD_95_U65 , P1_ADD_95_U66 , P1_ADD_95_U67 , P1_ADD_95_U68 , P1_ADD_95_U69 , P1_ADD_95_U70 , P1_ADD_95_U71 , P1_ADD_95_U72;
wire P1_ADD_95_U73 , P1_ADD_95_U74 , P1_ADD_95_U75 , P1_ADD_95_U76 , P1_ADD_95_U77 , P1_ADD_95_U78 , P1_ADD_95_U79 , P1_ADD_95_U80 , P1_ADD_95_U81 , P1_ADD_95_U82;
wire P1_ADD_95_U83 , P1_ADD_95_U84 , P1_ADD_95_U85 , P1_ADD_95_U86 , P1_ADD_95_U87 , P1_ADD_95_U88 , P1_ADD_95_U89 , P1_ADD_95_U90 , P1_ADD_95_U91 , P1_ADD_95_U92;
wire P1_ADD_95_U93 , P1_ADD_95_U94 , P1_ADD_95_U95 , P1_ADD_95_U96 , P1_ADD_95_U97 , P1_ADD_95_U98 , P1_ADD_95_U99 , P1_ADD_95_U100 , P1_ADD_95_U101 , P1_ADD_95_U102;
wire P1_ADD_95_U103 , P1_ADD_95_U104 , P1_ADD_95_U105 , P1_ADD_95_U106 , P1_ADD_95_U107 , P1_ADD_95_U108 , P1_ADD_95_U109 , P1_ADD_95_U110 , P1_ADD_95_U111 , P1_ADD_95_U112;
wire P1_ADD_95_U113 , P1_ADD_95_U114 , P1_ADD_95_U115 , P1_ADD_95_U116 , P1_ADD_95_U117 , P1_ADD_95_U118 , P1_ADD_95_U119 , P1_ADD_95_U120 , P1_ADD_95_U121 , P1_ADD_95_U122;
wire P1_ADD_95_U123 , P1_ADD_95_U124 , P1_ADD_95_U125 , P1_ADD_95_U126 , P1_ADD_95_U127 , P1_ADD_95_U128 , P1_ADD_95_U129 , P1_ADD_95_U130 , P1_ADD_95_U131 , P1_ADD_95_U132;
wire P1_ADD_95_U133 , P1_ADD_95_U134 , P1_ADD_95_U135 , P1_ADD_95_U136 , P1_ADD_95_U137 , P1_ADD_95_U138 , P1_ADD_95_U139 , P1_ADD_95_U140 , P1_ADD_95_U141 , P1_ADD_95_U142;
wire P1_ADD_95_U143 , P1_ADD_95_U144 , P1_ADD_95_U145 , P1_ADD_95_U146 , P1_ADD_95_U147 , P1_ADD_95_U148 , P1_ADD_95_U149 , P1_ADD_95_U150 , P1_ADD_95_U151 , P1_ADD_95_U152;
wire P1_ADD_95_U153 , P1_R1105_U4 , P1_R1105_U5 , P1_R1105_U6 , P1_R1105_U7 , P1_R1105_U8 , P1_R1105_U9 , P1_R1105_U10 , P1_R1105_U11 , P1_R1105_U12;
wire P1_R1105_U13 , P1_R1105_U14 , P1_R1105_U15 , P1_R1105_U16 , P1_R1105_U17 , P1_R1105_U18 , P1_R1105_U19 , P1_R1105_U20 , P1_R1105_U21 , P1_R1105_U22;
wire P1_R1105_U23 , P1_R1105_U24 , P1_R1105_U25 , P1_R1105_U26 , P1_R1105_U27 , P1_R1105_U28 , P1_R1105_U29 , P1_R1105_U30 , P1_R1105_U31 , P1_R1105_U32;
wire P1_R1105_U33 , P1_R1105_U34 , P1_R1105_U35 , P1_R1105_U36 , P1_R1105_U37 , P1_R1105_U38 , P1_R1105_U39 , P1_R1105_U40 , P1_R1105_U41 , P1_R1105_U42;
wire P1_R1105_U43 , P1_R1105_U44 , P1_R1105_U45 , P1_R1105_U46 , P1_R1105_U47 , P1_R1105_U48 , P1_R1105_U49 , P1_R1105_U50 , P1_R1105_U51 , P1_R1105_U52;
wire P1_R1105_U53 , P1_R1105_U54 , P1_R1105_U55 , P1_R1105_U56 , P1_R1105_U57 , P1_R1105_U58 , P1_R1105_U59 , P1_R1105_U60 , P1_R1105_U61 , P1_R1105_U62;
wire P1_R1105_U63 , P1_R1105_U64 , P1_R1105_U65 , P1_R1105_U66 , P1_R1105_U67 , P1_R1105_U68 , P1_R1105_U69 , P1_R1105_U70 , P1_R1105_U71 , P1_R1105_U72;
wire P1_R1105_U73 , P1_R1105_U74 , P1_R1105_U75 , P1_R1105_U76 , P1_R1105_U77 , P1_R1105_U78 , P1_R1105_U79 , P1_R1105_U80 , P1_R1105_U81 , P1_R1105_U82;
wire P1_R1105_U83 , P1_R1105_U84 , P1_R1105_U85 , P1_R1105_U86 , P1_R1105_U87 , P1_R1105_U88 , P1_R1105_U89 , P1_R1105_U90 , P1_R1105_U91 , P1_R1105_U92;
wire P1_R1105_U93 , P1_R1105_U94 , P1_R1105_U95 , P1_R1105_U96 , P1_R1105_U97 , P1_R1105_U98 , P1_R1105_U99 , P1_R1105_U100 , P1_R1105_U101 , P1_R1105_U102;
wire P1_R1105_U103 , P1_R1105_U104 , P1_R1105_U105 , P1_R1105_U106 , P1_R1105_U107 , P1_R1105_U108 , P1_R1105_U109 , P1_R1105_U110 , P1_R1105_U111 , P1_R1105_U112;
wire P1_R1105_U113 , P1_R1105_U114 , P1_R1105_U115 , P1_R1105_U116 , P1_R1105_U117 , P1_R1105_U118 , P1_R1105_U119 , P1_R1105_U120 , P1_R1105_U121 , P1_R1105_U122;
wire P1_R1105_U123 , P1_R1105_U124 , P1_R1105_U125 , P1_R1105_U126 , P1_R1105_U127 , P1_R1105_U128 , P1_R1105_U129 , P1_R1105_U130 , P1_R1105_U131 , P1_R1105_U132;
wire P1_R1105_U133 , P1_R1105_U134 , P1_R1105_U135 , P1_R1105_U136 , P1_R1105_U137 , P1_R1105_U138 , P1_R1105_U139 , P1_R1105_U140 , P1_R1105_U141 , P1_R1105_U142;
wire P1_R1105_U143 , P1_R1105_U144 , P1_R1105_U145 , P1_R1105_U146 , P1_R1105_U147 , P1_R1105_U148 , P1_R1105_U149 , P1_R1105_U150 , P1_R1105_U151 , P1_R1105_U152;
wire P1_R1105_U153 , P1_R1105_U154 , P1_R1105_U155 , P1_R1105_U156 , P1_R1105_U157 , P1_R1105_U158 , P1_R1105_U159 , P1_R1105_U160 , P1_R1105_U161 , P1_R1105_U162;
wire P1_R1105_U163 , P1_R1105_U164 , P1_R1105_U165 , P1_R1105_U166 , P1_R1105_U167 , P1_R1105_U168 , P1_R1105_U169 , P1_R1105_U170 , P1_R1105_U171 , P1_R1105_U172;
wire P1_R1105_U173 , P1_R1105_U174 , P1_R1105_U175 , P1_R1105_U176 , P1_R1105_U177 , P1_R1105_U178 , P1_R1105_U179 , P1_R1105_U180 , P1_R1105_U181 , P1_R1105_U182;
wire P1_R1105_U183 , P1_R1105_U184 , P1_R1105_U185 , P1_R1105_U186 , P1_R1105_U187 , P1_R1105_U188 , P1_R1105_U189 , P1_R1105_U190 , P1_R1105_U191 , P1_R1105_U192;
wire P1_R1105_U193 , P1_R1105_U194 , P1_R1105_U195 , P1_R1105_U196 , P1_R1105_U197 , P1_R1105_U198 , P1_R1105_U199 , P1_R1105_U200 , P1_R1105_U201 , P1_R1105_U202;
wire P1_R1105_U203 , P1_R1105_U204 , P1_R1105_U205 , P1_R1105_U206 , P1_R1105_U207 , P1_R1105_U208 , P1_R1105_U209 , P1_R1105_U210 , P1_R1105_U211 , P1_R1105_U212;
wire P1_R1105_U213 , P1_R1105_U214 , P1_R1105_U215 , P1_R1105_U216 , P1_R1105_U217 , P1_R1105_U218 , P1_R1105_U219 , P1_R1105_U220 , P1_R1105_U221 , P1_R1105_U222;
wire P1_R1105_U223 , P1_R1105_U224 , P1_R1105_U225 , P1_R1105_U226 , P1_R1105_U227 , P1_R1105_U228 , P1_R1105_U229 , P1_R1105_U230 , P1_R1105_U231 , P1_R1105_U232;
wire P1_R1105_U233 , P1_R1105_U234 , P1_R1105_U235 , P1_R1105_U236 , P1_R1105_U237 , P1_R1105_U238 , P1_R1105_U239 , P1_R1105_U240 , P1_R1105_U241 , P1_R1105_U242;
wire P1_R1105_U243 , P1_R1105_U244 , P1_R1105_U245 , P1_R1105_U246 , P1_R1105_U247 , P1_R1105_U248 , P1_R1105_U249 , P1_R1105_U250 , P1_R1105_U251 , P1_R1105_U252;
wire P1_R1105_U253 , P1_R1105_U254 , P1_R1105_U255 , P1_R1105_U256 , P1_R1105_U257 , P1_R1105_U258 , P1_R1105_U259 , P1_R1105_U260 , P1_R1105_U261 , P1_R1105_U262;
wire P1_R1105_U263 , P1_R1105_U264 , P1_R1105_U265 , P1_R1105_U266 , P1_R1105_U267 , P1_R1105_U268 , P1_R1105_U269 , P1_R1105_U270 , P1_R1105_U271 , P1_R1105_U272;
wire P1_R1105_U273 , P1_R1105_U274 , P1_R1105_U275 , P1_R1105_U276 , P1_R1105_U277 , P1_R1105_U278 , P1_R1105_U279 , P1_R1105_U280 , P1_R1105_U281 , P1_R1105_U282;
wire P1_R1105_U283 , P1_R1105_U284 , P1_R1105_U285 , P1_R1105_U286 , P1_R1105_U287 , P1_R1105_U288 , P1_R1105_U289 , P1_R1105_U290 , P1_R1105_U291 , P1_R1105_U292;
wire P1_R1105_U293 , P1_R1105_U294 , P1_R1105_U295 , P1_R1105_U296 , P1_R1105_U297 , P1_R1105_U298 , P1_R1105_U299 , P1_R1105_U300 , P1_R1105_U301 , P1_R1105_U302;
wire P1_R1105_U303 , P1_R1105_U304 , P1_R1105_U305 , P1_R1105_U306 , P1_R1105_U307 , P1_R1105_U308 , P1_SUB_84_U6 , P1_SUB_84_U7 , P1_SUB_84_U8 , P1_SUB_84_U9;
wire P1_SUB_84_U10 , P1_SUB_84_U11 , P1_SUB_84_U12 , P1_SUB_84_U13 , P1_SUB_84_U14 , P1_SUB_84_U15 , P1_SUB_84_U16 , P1_SUB_84_U17 , P1_SUB_84_U18 , P1_SUB_84_U19;
wire P1_SUB_84_U20 , P1_SUB_84_U21 , P1_SUB_84_U22 , P1_SUB_84_U23 , P1_SUB_84_U24 , P1_SUB_84_U25 , P1_SUB_84_U26 , P1_SUB_84_U27 , P1_SUB_84_U28 , P1_SUB_84_U29;
wire P1_SUB_84_U30 , P1_SUB_84_U31 , P1_SUB_84_U32 , P1_SUB_84_U33 , P1_SUB_84_U34 , P1_SUB_84_U35 , P1_SUB_84_U36 , P1_SUB_84_U37 , P1_SUB_84_U38 , P1_SUB_84_U39;
wire P1_SUB_84_U40 , P1_SUB_84_U41 , P1_SUB_84_U42 , P1_SUB_84_U43 , P1_SUB_84_U44 , P1_SUB_84_U45 , P1_SUB_84_U46 , P1_SUB_84_U47 , P1_SUB_84_U48 , P1_SUB_84_U49;
wire P1_SUB_84_U50 , P1_SUB_84_U51 , P1_SUB_84_U52 , P1_SUB_84_U53 , P1_SUB_84_U54 , P1_SUB_84_U55 , P1_SUB_84_U56 , P1_SUB_84_U57 , P1_SUB_84_U58 , P1_SUB_84_U59;
wire P1_SUB_84_U60 , P1_SUB_84_U61 , P1_SUB_84_U62 , P1_SUB_84_U63 , P1_SUB_84_U64 , P1_SUB_84_U65 , P1_SUB_84_U66 , P1_SUB_84_U67 , P1_SUB_84_U68 , P1_SUB_84_U69;
wire P1_SUB_84_U70 , P1_SUB_84_U71 , P1_SUB_84_U72 , P1_SUB_84_U73 , P1_SUB_84_U74 , P1_SUB_84_U75 , P1_SUB_84_U76 , P1_SUB_84_U77 , P1_SUB_84_U78 , P1_SUB_84_U79;
wire P1_SUB_84_U80 , P1_SUB_84_U81 , P1_SUB_84_U82 , P1_SUB_84_U83 , P1_SUB_84_U84 , P1_SUB_84_U85 , P1_SUB_84_U86 , P1_SUB_84_U87 , P1_SUB_84_U88 , P1_SUB_84_U89;
wire P1_SUB_84_U90 , P1_SUB_84_U91 , P1_SUB_84_U92 , P1_SUB_84_U93 , P1_SUB_84_U94 , P1_SUB_84_U95 , P1_SUB_84_U96 , P1_SUB_84_U97 , P1_SUB_84_U98 , P1_SUB_84_U99;
wire P1_SUB_84_U100 , P1_SUB_84_U101 , P1_SUB_84_U102 , P1_SUB_84_U103 , P1_SUB_84_U104 , P1_SUB_84_U105 , P1_SUB_84_U106 , P1_SUB_84_U107 , P1_SUB_84_U108 , P1_SUB_84_U109;
wire P1_SUB_84_U110 , P1_SUB_84_U111 , P1_SUB_84_U112 , P1_SUB_84_U113 , P1_SUB_84_U114 , P1_SUB_84_U115 , P1_SUB_84_U116 , P1_SUB_84_U117 , P1_SUB_84_U118 , P1_SUB_84_U119;
wire P1_SUB_84_U120 , P1_SUB_84_U121 , P1_SUB_84_U122 , P1_SUB_84_U123 , P1_SUB_84_U124 , P1_SUB_84_U125 , P1_SUB_84_U126 , P1_SUB_84_U127 , P1_SUB_84_U128 , P1_SUB_84_U129;
wire P1_SUB_84_U130 , P1_SUB_84_U131 , P1_SUB_84_U132 , P1_SUB_84_U133 , P1_SUB_84_U134 , P1_SUB_84_U135 , P1_SUB_84_U136 , P1_SUB_84_U137 , P1_SUB_84_U138 , P1_SUB_84_U139;
wire P1_SUB_84_U140 , P1_SUB_84_U141 , P1_SUB_84_U142 , P1_SUB_84_U143 , P1_SUB_84_U144 , P1_SUB_84_U145 , P1_SUB_84_U146 , P1_SUB_84_U147 , P1_SUB_84_U148 , P1_SUB_84_U149;
wire P1_SUB_84_U150 , P1_SUB_84_U151 , P1_SUB_84_U152 , P1_SUB_84_U153 , P1_SUB_84_U154 , P1_SUB_84_U155 , P1_SUB_84_U156 , P1_SUB_84_U157 , P1_SUB_84_U158 , P1_SUB_84_U159;
wire P1_SUB_84_U160 , P1_SUB_84_U161 , P1_SUB_84_U162 , P1_SUB_84_U163 , P1_SUB_84_U164 , P1_SUB_84_U165 , P1_SUB_84_U166 , P1_SUB_84_U167 , P1_SUB_84_U168 , P1_SUB_84_U169;
wire P1_SUB_84_U170 , P1_SUB_84_U171 , P1_SUB_84_U172 , P1_SUB_84_U173 , P1_SUB_84_U174 , P1_SUB_84_U175 , P1_SUB_84_U176 , P1_SUB_84_U177 , P1_SUB_84_U178 , P1_SUB_84_U179;
wire P1_SUB_84_U180 , P1_SUB_84_U181 , P1_SUB_84_U182 , P1_SUB_84_U183 , P1_SUB_84_U184 , P1_SUB_84_U185 , P1_SUB_84_U186 , P1_SUB_84_U187 , P1_SUB_84_U188 , P1_SUB_84_U189;
wire P1_SUB_84_U190 , P1_SUB_84_U191 , P1_SUB_84_U192 , P1_SUB_84_U193 , P1_SUB_84_U194 , P1_SUB_84_U195 , P1_SUB_84_U196 , P1_SUB_84_U197 , P1_SUB_84_U198 , P1_SUB_84_U199;
wire P1_SUB_84_U200 , P1_SUB_84_U201 , P1_SUB_84_U202 , P1_SUB_84_U203 , P1_SUB_84_U204 , P1_SUB_84_U205 , P1_SUB_84_U206 , P1_SUB_84_U207 , P1_SUB_84_U208 , P1_SUB_84_U209;
wire P1_SUB_84_U210 , P1_SUB_84_U211 , P1_SUB_84_U212 , P1_SUB_84_U213 , P1_SUB_84_U214 , P1_SUB_84_U215 , P1_SUB_84_U216 , P1_SUB_84_U217 , P1_SUB_84_U218 , P1_SUB_84_U219;
wire P1_SUB_84_U220 , P1_SUB_84_U221 , P1_SUB_84_U222 , P1_SUB_84_U223 , P1_SUB_84_U224 , P1_SUB_84_U225 , P1_SUB_84_U226 , P1_SUB_84_U227 , P1_SUB_84_U228 , P1_SUB_84_U229;
wire P1_SUB_84_U230 , P1_SUB_84_U231 , P1_SUB_84_U232 , P1_SUB_84_U233 , P1_SUB_84_U234 , P1_SUB_84_U235 , P1_SUB_84_U236 , P1_SUB_84_U237 , P1_SUB_84_U238 , P1_SUB_84_U239;
wire P1_SUB_84_U240 , P1_SUB_84_U241 , P1_SUB_84_U242 , P1_SUB_84_U243 , P1_SUB_84_U244 , P1_SUB_84_U245 , P1_SUB_84_U246 , P1_SUB_84_U247 , P1_SUB_84_U248 , P1_SUB_84_U249;
wire P1_SUB_84_U250 , P1_SUB_84_U251 , P1_R1309_U6 , P1_R1309_U7 , P1_R1309_U8 , P1_R1309_U9 , P1_R1309_U10 , P1_R1282_U6 , P1_R1282_U7 , P1_R1282_U8;
wire P1_R1282_U9 , P1_R1282_U10 , P1_R1282_U11 , P1_R1282_U12 , P1_R1282_U13 , P1_R1282_U14 , P1_R1282_U15 , P1_R1282_U16 , P1_R1282_U17 , P1_R1282_U18;
wire P1_R1282_U19 , P1_R1282_U20 , P1_R1282_U21 , P1_R1282_U22 , P1_R1282_U23 , P1_R1282_U24 , P1_R1282_U25 , P1_R1282_U26 , P1_R1282_U27 , P1_R1282_U28;
wire P1_R1282_U29 , P1_R1282_U30 , P1_R1282_U31 , P1_R1282_U32 , P1_R1282_U33 , P1_R1282_U34 , P1_R1282_U35 , P1_R1282_U36 , P1_R1282_U37 , P1_R1282_U38;
wire P1_R1282_U39 , P1_R1282_U40 , P1_R1282_U41 , P1_R1282_U42 , P1_R1282_U43 , P1_R1282_U44 , P1_R1282_U45 , P1_R1282_U46 , P1_R1282_U47 , P1_R1282_U48;
wire P1_R1282_U49 , P1_R1282_U50 , P1_R1282_U51 , P1_R1282_U52 , P1_R1282_U53 , P1_R1282_U54 , P1_R1282_U55 , P1_R1282_U56 , P1_R1282_U57 , P1_R1282_U58;
wire P1_R1282_U59 , P1_R1282_U60 , P1_R1282_U61 , P1_R1282_U62 , P1_R1282_U63 , P1_R1282_U64 , P1_R1282_U65 , P1_R1282_U66 , P1_R1282_U67 , P1_R1282_U68;
wire P1_R1282_U69 , P1_R1282_U70 , P1_R1282_U71 , P1_R1282_U72 , P1_R1282_U73 , P1_R1282_U74 , P1_R1282_U75 , P1_R1282_U76 , P1_R1282_U77 , P1_R1282_U78;
wire P1_R1282_U79 , P1_R1282_U80 , P1_R1282_U81 , P1_R1282_U82 , P1_R1282_U83 , P1_R1282_U84 , P1_R1282_U85 , P1_R1282_U86 , P1_R1282_U87 , P1_R1282_U88;
wire P1_R1282_U89 , P1_R1282_U90 , P1_R1282_U91 , P1_R1282_U92 , P1_R1282_U93 , P1_R1282_U94 , P1_R1282_U95 , P1_R1282_U96 , P1_R1282_U97 , P1_R1282_U98;
wire P1_R1282_U99 , P1_R1282_U100 , P1_R1282_U101 , P1_R1282_U102 , P1_R1282_U103 , P1_R1282_U104 , P1_R1282_U105 , P1_R1282_U106 , P1_R1282_U107 , P1_R1282_U108;
wire P1_R1282_U109 , P1_R1282_U110 , P1_R1282_U111 , P1_R1282_U112 , P1_R1282_U113 , P1_R1282_U114 , P1_R1282_U115 , P1_R1282_U116 , P1_R1282_U117 , P1_R1282_U118;
wire P1_R1282_U119 , P1_R1282_U120 , P1_R1282_U121 , P1_R1282_U122 , P1_R1282_U123 , P1_R1282_U124 , P1_R1282_U125 , P1_R1282_U126 , P1_R1282_U127 , P1_R1282_U128;
wire P1_R1282_U129 , P1_R1282_U130 , P1_R1282_U131 , P1_R1282_U132 , P1_R1282_U133 , P1_R1282_U134 , P1_R1282_U135 , P1_R1282_U136 , P1_R1282_U137 , P1_R1282_U138;
wire P1_R1282_U139 , P1_R1282_U140 , P1_R1282_U141 , P1_R1282_U142 , P1_R1282_U143 , P1_R1282_U144 , P1_R1282_U145 , P1_R1282_U146 , P1_R1282_U147 , P1_R1282_U148;
wire P1_R1282_U149 , P1_R1282_U150 , P1_R1282_U151 , P1_R1282_U152 , P1_R1282_U153 , P1_R1282_U154 , P1_R1282_U155 , P1_R1282_U156 , P1_R1282_U157 , P1_R1282_U158;
wire P1_R1282_U159 , P1_R1240_U4 , P1_R1240_U5 , P1_R1240_U6 , P1_R1240_U7 , P1_R1240_U8 , P1_R1240_U9 , P1_R1240_U10 , P1_R1240_U11 , P1_R1240_U12;
wire P1_R1240_U13 , P1_R1240_U14 , P1_R1240_U15 , P1_R1240_U16 , P1_R1240_U17 , P1_R1240_U18 , P1_R1240_U19 , P1_R1240_U20 , P1_R1240_U21 , P1_R1240_U22;
wire P1_R1240_U23 , P1_R1240_U24 , P1_R1240_U25 , P1_R1240_U26 , P1_R1240_U27 , P1_R1240_U28 , P1_R1240_U29 , P1_R1240_U30 , P1_R1240_U31 , P1_R1240_U32;
wire P1_R1240_U33 , P1_R1240_U34 , P1_R1240_U35 , P1_R1240_U36 , P1_R1240_U37 , P1_R1240_U38 , P1_R1240_U39 , P1_R1240_U40 , P1_R1240_U41 , P1_R1240_U42;
wire P1_R1240_U43 , P1_R1240_U44 , P1_R1240_U45 , P1_R1240_U46 , P1_R1240_U47 , P1_R1240_U48 , P1_R1240_U49 , P1_R1240_U50 , P1_R1240_U51 , P1_R1240_U52;
wire P1_R1240_U53 , P1_R1240_U54 , P1_R1240_U55 , P1_R1240_U56 , P1_R1240_U57 , P1_R1240_U58 , P1_R1240_U59 , P1_R1240_U60 , P1_R1240_U61 , P1_R1240_U62;
wire P1_R1240_U63 , P1_R1240_U64 , P1_R1240_U65 , P1_R1240_U66 , P1_R1240_U67 , P1_R1240_U68 , P1_R1240_U69 , P1_R1240_U70 , P1_R1240_U71 , P1_R1240_U72;
wire P1_R1240_U73 , P1_R1240_U74 , P1_R1240_U75 , P1_R1240_U76 , P1_R1240_U77 , P1_R1240_U78 , P1_R1240_U79 , P1_R1240_U80 , P1_R1240_U81 , P1_R1240_U82;
wire P1_R1240_U83 , P1_R1240_U84 , P1_R1240_U85 , P1_R1240_U86 , P1_R1240_U87 , P1_R1240_U88 , P1_R1240_U89 , P1_R1240_U90 , P1_R1240_U91 , P1_R1240_U92;
wire P1_R1240_U93 , P1_R1240_U94 , P1_R1240_U95 , P1_R1240_U96 , P1_R1240_U97 , P1_R1240_U98 , P1_R1240_U99 , P1_R1240_U100 , P1_R1240_U101 , P1_R1240_U102;
wire P1_R1240_U103 , P1_R1240_U104 , P1_R1240_U105 , P1_R1240_U106 , P1_R1240_U107 , P1_R1240_U108 , P1_R1240_U109 , P1_R1240_U110 , P1_R1240_U111 , P1_R1240_U112;
wire P1_R1240_U113 , P1_R1240_U114 , P1_R1240_U115 , P1_R1240_U116 , P1_R1240_U117 , P1_R1240_U118 , P1_R1240_U119 , P1_R1240_U120 , P1_R1240_U121 , P1_R1240_U122;
wire P1_R1240_U123 , P1_R1240_U124 , P1_R1240_U125 , P1_R1240_U126 , P1_R1240_U127 , P1_R1240_U128 , P1_R1240_U129 , P1_R1240_U130 , P1_R1240_U131 , P1_R1240_U132;
wire P1_R1240_U133 , P1_R1240_U134 , P1_R1240_U135 , P1_R1240_U136 , P1_R1240_U137 , P1_R1240_U138 , P1_R1240_U139 , P1_R1240_U140 , P1_R1240_U141 , P1_R1240_U142;
wire P1_R1240_U143 , P1_R1240_U144 , P1_R1240_U145 , P1_R1240_U146 , P1_R1240_U147 , P1_R1240_U148 , P1_R1240_U149 , P1_R1240_U150 , P1_R1240_U151 , P1_R1240_U152;
wire P1_R1240_U153 , P1_R1240_U154 , P1_R1240_U155 , P1_R1240_U156 , P1_R1240_U157 , P1_R1240_U158 , P1_R1240_U159 , P1_R1240_U160 , P1_R1240_U161 , P1_R1240_U162;
wire P1_R1240_U163 , P1_R1240_U164 , P1_R1240_U165 , P1_R1240_U166 , P1_R1240_U167 , P1_R1240_U168 , P1_R1240_U169 , P1_R1240_U170 , P1_R1240_U171 , P1_R1240_U172;
wire P1_R1240_U173 , P1_R1240_U174 , P1_R1240_U175 , P1_R1240_U176 , P1_R1240_U177 , P1_R1240_U178 , P1_R1240_U179 , P1_R1240_U180 , P1_R1240_U181 , P1_R1240_U182;
wire P1_R1240_U183 , P1_R1240_U184 , P1_R1240_U185 , P1_R1240_U186 , P1_R1240_U187 , P1_R1240_U188 , P1_R1240_U189 , P1_R1240_U190 , P1_R1240_U191 , P1_R1240_U192;
wire P1_R1240_U193 , P1_R1240_U194 , P1_R1240_U195 , P1_R1240_U196 , P1_R1240_U197 , P1_R1240_U198 , P1_R1240_U199 , P1_R1240_U200 , P1_R1240_U201 , P1_R1240_U202;
wire P1_R1240_U203 , P1_R1240_U204 , P1_R1240_U205 , P1_R1240_U206 , P1_R1240_U207 , P1_R1240_U208 , P1_R1240_U209 , P1_R1240_U210 , P1_R1240_U211 , P1_R1240_U212;
wire P1_R1240_U213 , P1_R1240_U214 , P1_R1240_U215 , P1_R1240_U216 , P1_R1240_U217 , P1_R1240_U218 , P1_R1240_U219 , P1_R1240_U220 , P1_R1240_U221 , P1_R1240_U222;
wire P1_R1240_U223 , P1_R1240_U224 , P1_R1240_U225 , P1_R1240_U226 , P1_R1240_U227 , P1_R1240_U228 , P1_R1240_U229 , P1_R1240_U230 , P1_R1240_U231 , P1_R1240_U232;
wire P1_R1240_U233 , P1_R1240_U234 , P1_R1240_U235 , P1_R1240_U236 , P1_R1240_U237 , P1_R1240_U238 , P1_R1240_U239 , P1_R1240_U240 , P1_R1240_U241 , P1_R1240_U242;
wire P1_R1240_U243 , P1_R1240_U244 , P1_R1240_U245 , P1_R1240_U246 , P1_R1240_U247 , P1_R1240_U248 , P1_R1240_U249 , P1_R1240_U250 , P1_R1240_U251 , P1_R1240_U252;
wire P1_R1240_U253 , P1_R1240_U254 , P1_R1240_U255 , P1_R1240_U256 , P1_R1240_U257 , P1_R1240_U258 , P1_R1240_U259 , P1_R1240_U260 , P1_R1240_U261 , P1_R1240_U262;
wire P1_R1240_U263 , P1_R1240_U264 , P1_R1240_U265 , P1_R1240_U266 , P1_R1240_U267 , P1_R1240_U268 , P1_R1240_U269 , P1_R1240_U270 , P1_R1240_U271 , P1_R1240_U272;
wire P1_R1240_U273 , P1_R1240_U274 , P1_R1240_U275 , P1_R1240_U276 , P1_R1240_U277 , P1_R1240_U278 , P1_R1240_U279 , P1_R1240_U280 , P1_R1240_U281 , P1_R1240_U282;
wire P1_R1240_U283 , P1_R1240_U284 , P1_R1240_U285 , P1_R1240_U286 , P1_R1240_U287 , P1_R1240_U288 , P1_R1240_U289 , P1_R1240_U290 , P1_R1240_U291 , P1_R1240_U292;
wire P1_R1240_U293 , P1_R1240_U294 , P1_R1240_U295 , P1_R1240_U296 , P1_R1240_U297 , P1_R1240_U298 , P1_R1240_U299 , P1_R1240_U300 , P1_R1240_U301 , P1_R1240_U302;
wire P1_R1240_U303 , P1_R1240_U304 , P1_R1240_U305 , P1_R1240_U306 , P1_R1240_U307 , P1_R1240_U308 , P1_R1240_U309 , P1_R1240_U310 , P1_R1240_U311 , P1_R1240_U312;
wire P1_R1240_U313 , P1_R1240_U314 , P1_R1240_U315 , P1_R1240_U316 , P1_R1240_U317 , P1_R1240_U318 , P1_R1240_U319 , P1_R1240_U320 , P1_R1240_U321 , P1_R1240_U322;
wire P1_R1240_U323 , P1_R1240_U324 , P1_R1240_U325 , P1_R1240_U326 , P1_R1240_U327 , P1_R1240_U328 , P1_R1240_U329 , P1_R1240_U330 , P1_R1240_U331 , P1_R1240_U332;
wire P1_R1240_U333 , P1_R1240_U334 , P1_R1240_U335 , P1_R1240_U336 , P1_R1240_U337 , P1_R1240_U338 , P1_R1240_U339 , P1_R1240_U340 , P1_R1240_U341 , P1_R1240_U342;
wire P1_R1240_U343 , P1_R1240_U344 , P1_R1240_U345 , P1_R1240_U346 , P1_R1240_U347 , P1_R1240_U348 , P1_R1240_U349 , P1_R1240_U350 , P1_R1240_U351 , P1_R1240_U352;
wire P1_R1240_U353 , P1_R1240_U354 , P1_R1240_U355 , P1_R1240_U356 , P1_R1240_U357 , P1_R1240_U358 , P1_R1240_U359 , P1_R1240_U360 , P1_R1240_U361 , P1_R1240_U362;
wire P1_R1240_U363 , P1_R1240_U364 , P1_R1240_U365 , P1_R1240_U366 , P1_R1240_U367 , P1_R1240_U368 , P1_R1240_U369 , P1_R1240_U370 , P1_R1240_U371 , P1_R1240_U372;
wire P1_R1240_U373 , P1_R1240_U374 , P1_R1240_U375 , P1_R1240_U376 , P1_R1240_U377 , P1_R1240_U378 , P1_R1240_U379 , P1_R1240_U380 , P1_R1240_U381 , P1_R1240_U382;
wire P1_R1240_U383 , P1_R1240_U384 , P1_R1240_U385 , P1_R1240_U386 , P1_R1240_U387 , P1_R1240_U388 , P1_R1240_U389 , P1_R1240_U390 , P1_R1240_U391 , P1_R1240_U392;
wire P1_R1240_U393 , P1_R1240_U394 , P1_R1240_U395 , P1_R1240_U396 , P1_R1240_U397 , P1_R1240_U398 , P1_R1240_U399 , P1_R1240_U400 , P1_R1240_U401 , P1_R1240_U402;
wire P1_R1240_U403 , P1_R1240_U404 , P1_R1240_U405 , P1_R1240_U406 , P1_R1240_U407 , P1_R1240_U408 , P1_R1240_U409 , P1_R1240_U410 , P1_R1240_U411 , P1_R1240_U412;
wire P1_R1240_U413 , P1_R1240_U414 , P1_R1240_U415 , P1_R1240_U416 , P1_R1240_U417 , P1_R1240_U418 , P1_R1240_U419 , P1_R1240_U420 , P1_R1240_U421 , P1_R1240_U422;
wire P1_R1240_U423 , P1_R1240_U424 , P1_R1240_U425 , P1_R1240_U426 , P1_R1240_U427 , P1_R1240_U428 , P1_R1240_U429 , P1_R1240_U430 , P1_R1240_U431 , P1_R1240_U432;
wire P1_R1240_U433 , P1_R1240_U434 , P1_R1240_U435 , P1_R1240_U436 , P1_R1240_U437 , P1_R1240_U438 , P1_R1240_U439 , P1_R1240_U440 , P1_R1240_U441 , P1_R1240_U442;
wire P1_R1240_U443 , P1_R1240_U444 , P1_R1240_U445 , P1_R1240_U446 , P1_R1240_U447 , P1_R1240_U448 , P1_R1240_U449 , P1_R1240_U450 , P1_R1240_U451 , P1_R1240_U452;
wire P1_R1240_U453 , P1_R1240_U454 , P1_R1240_U455 , P1_R1240_U456 , P1_R1240_U457 , P1_R1240_U458 , P1_R1240_U459 , P1_R1240_U460 , P1_R1240_U461 , P1_R1240_U462;
wire P1_R1240_U463 , P1_R1240_U464 , P1_R1240_U465 , P1_R1240_U466 , P1_R1240_U467 , P1_R1240_U468 , P1_R1240_U469 , P1_R1240_U470 , P1_R1240_U471 , P1_R1240_U472;
wire P1_R1240_U473 , P1_R1240_U474 , P1_R1240_U475 , P1_R1240_U476 , P1_R1240_U477 , P1_R1240_U478 , P1_R1240_U479 , P1_R1240_U480 , P1_R1240_U481 , P1_R1240_U482;
wire P1_R1240_U483 , P1_R1240_U484 , P1_R1240_U485 , P1_R1240_U486 , P1_R1240_U487 , P1_R1240_U488 , P1_R1240_U489 , P1_R1240_U490 , P1_R1240_U491 , P1_R1240_U492;
wire P1_R1240_U493 , P1_R1240_U494 , P1_R1240_U495 , P1_R1240_U496 , P1_R1240_U497 , P1_R1240_U498 , P1_R1240_U499 , P1_R1240_U500 , P1_R1240_U501 , P1_R1240_U502;
wire P1_R1240_U503 , P1_R1162_U4 , P1_R1162_U5 , P1_R1162_U6 , P1_R1162_U7 , P1_R1162_U8 , P1_R1162_U9 , P1_R1162_U10 , P1_R1162_U11 , P1_R1162_U12;
wire P1_R1162_U13 , P1_R1162_U14 , P1_R1162_U15 , P1_R1162_U16 , P1_R1162_U17 , P1_R1162_U18 , P1_R1162_U19 , P1_R1162_U20 , P1_R1162_U21 , P1_R1162_U22;
wire P1_R1162_U23 , P1_R1162_U24 , P1_R1162_U25 , P1_R1162_U26 , P1_R1162_U27 , P1_R1162_U28 , P1_R1162_U29 , P1_R1162_U30 , P1_R1162_U31 , P1_R1162_U32;
wire P1_R1162_U33 , P1_R1162_U34 , P1_R1162_U35 , P1_R1162_U36 , P1_R1162_U37 , P1_R1162_U38 , P1_R1162_U39 , P1_R1162_U40 , P1_R1162_U41 , P1_R1162_U42;
wire P1_R1162_U43 , P1_R1162_U44 , P1_R1162_U45 , P1_R1162_U46 , P1_R1162_U47 , P1_R1162_U48 , P1_R1162_U49 , P1_R1162_U50 , P1_R1162_U51 , P1_R1162_U52;
wire P1_R1162_U53 , P1_R1162_U54 , P1_R1162_U55 , P1_R1162_U56 , P1_R1162_U57 , P1_R1162_U58 , P1_R1162_U59 , P1_R1162_U60 , P1_R1162_U61 , P1_R1162_U62;
wire P1_R1162_U63 , P1_R1162_U64 , P1_R1162_U65 , P1_R1162_U66 , P1_R1162_U67 , P1_R1162_U68 , P1_R1162_U69 , P1_R1162_U70 , P1_R1162_U71 , P1_R1162_U72;
wire P1_R1162_U73 , P1_R1162_U74 , P1_R1162_U75 , P1_R1162_U76 , P1_R1162_U77 , P1_R1162_U78 , P1_R1162_U79 , P1_R1162_U80 , P1_R1162_U81 , P1_R1162_U82;
wire P1_R1162_U83 , P1_R1162_U84 , P1_R1162_U85 , P1_R1162_U86 , P1_R1162_U87 , P1_R1162_U88 , P1_R1162_U89 , P1_R1162_U90 , P1_R1162_U91 , P1_R1162_U92;
wire P1_R1162_U93 , P1_R1162_U94 , P1_R1162_U95 , P1_R1162_U96 , P1_R1162_U97 , P1_R1162_U98 , P1_R1162_U99 , P1_R1162_U100 , P1_R1162_U101 , P1_R1162_U102;
wire P1_R1162_U103 , P1_R1162_U104 , P1_R1162_U105 , P1_R1162_U106 , P1_R1162_U107 , P1_R1162_U108 , P1_R1162_U109 , P1_R1162_U110 , P1_R1162_U111 , P1_R1162_U112;
wire P1_R1162_U113 , P1_R1162_U114 , P1_R1162_U115 , P1_R1162_U116 , P1_R1162_U117 , P1_R1162_U118 , P1_R1162_U119 , P1_R1162_U120 , P1_R1162_U121 , P1_R1162_U122;
wire P1_R1162_U123 , P1_R1162_U124 , P1_R1162_U125 , P1_R1162_U126 , P1_R1162_U127 , P1_R1162_U128 , P1_R1162_U129 , P1_R1162_U130 , P1_R1162_U131 , P1_R1162_U132;
wire P1_R1162_U133 , P1_R1162_U134 , P1_R1162_U135 , P1_R1162_U136 , P1_R1162_U137 , P1_R1162_U138 , P1_R1162_U139 , P1_R1162_U140 , P1_R1162_U141 , P1_R1162_U142;
wire P1_R1162_U143 , P1_R1162_U144 , P1_R1162_U145 , P1_R1162_U146 , P1_R1162_U147 , P1_R1162_U148 , P1_R1162_U149 , P1_R1162_U150 , P1_R1162_U151 , P1_R1162_U152;
wire P1_R1162_U153 , P1_R1162_U154 , P1_R1162_U155 , P1_R1162_U156 , P1_R1162_U157 , P1_R1162_U158 , P1_R1162_U159 , P1_R1162_U160 , P1_R1162_U161 , P1_R1162_U162;
wire P1_R1162_U163 , P1_R1162_U164 , P1_R1162_U165 , P1_R1162_U166 , P1_R1162_U167 , P1_R1162_U168 , P1_R1162_U169 , P1_R1162_U170 , P1_R1162_U171 , P1_R1162_U172;
wire P1_R1162_U173 , P1_R1162_U174 , P1_R1162_U175 , P1_R1162_U176 , P1_R1162_U177 , P1_R1162_U178 , P1_R1162_U179 , P1_R1162_U180 , P1_R1162_U181 , P1_R1162_U182;
wire P1_R1162_U183 , P1_R1162_U184 , P1_R1162_U185 , P1_R1162_U186 , P1_R1162_U187 , P1_R1162_U188 , P1_R1162_U189 , P1_R1162_U190 , P1_R1162_U191 , P1_R1162_U192;
wire P1_R1162_U193 , P1_R1162_U194 , P1_R1162_U195 , P1_R1162_U196 , P1_R1162_U197 , P1_R1162_U198 , P1_R1162_U199 , P1_R1162_U200 , P1_R1162_U201 , P1_R1162_U202;
wire P1_R1162_U203 , P1_R1162_U204 , P1_R1162_U205 , P1_R1162_U206 , P1_R1162_U207 , P1_R1162_U208 , P1_R1162_U209 , P1_R1162_U210 , P1_R1162_U211 , P1_R1162_U212;
wire P1_R1162_U213 , P1_R1162_U214 , P1_R1162_U215 , P1_R1162_U216 , P1_R1162_U217 , P1_R1162_U218 , P1_R1162_U219 , P1_R1162_U220 , P1_R1162_U221 , P1_R1162_U222;
wire P1_R1162_U223 , P1_R1162_U224 , P1_R1162_U225 , P1_R1162_U226 , P1_R1162_U227 , P1_R1162_U228 , P1_R1162_U229 , P1_R1162_U230 , P1_R1162_U231 , P1_R1162_U232;
wire P1_R1162_U233 , P1_R1162_U234 , P1_R1162_U235 , P1_R1162_U236 , P1_R1162_U237 , P1_R1162_U238 , P1_R1162_U239 , P1_R1162_U240 , P1_R1162_U241 , P1_R1162_U242;
wire P1_R1162_U243 , P1_R1162_U244 , P1_R1162_U245 , P1_R1162_U246 , P1_R1162_U247 , P1_R1162_U248 , P1_R1162_U249 , P1_R1162_U250 , P1_R1162_U251 , P1_R1162_U252;
wire P1_R1162_U253 , P1_R1162_U254 , P1_R1162_U255 , P1_R1162_U256 , P1_R1162_U257 , P1_R1162_U258 , P1_R1162_U259 , P1_R1162_U260 , P1_R1162_U261 , P1_R1162_U262;
wire P1_R1162_U263 , P1_R1162_U264 , P1_R1162_U265 , P1_R1162_U266 , P1_R1162_U267 , P1_R1162_U268 , P1_R1162_U269 , P1_R1162_U270 , P1_R1162_U271 , P1_R1162_U272;
wire P1_R1162_U273 , P1_R1162_U274 , P1_R1162_U275 , P1_R1162_U276 , P1_R1162_U277 , P1_R1162_U278 , P1_R1162_U279 , P1_R1162_U280 , P1_R1162_U281 , P1_R1162_U282;
wire P1_R1162_U283 , P1_R1162_U284 , P1_R1162_U285 , P1_R1162_U286 , P1_R1162_U287 , P1_R1162_U288 , P1_R1162_U289 , P1_R1162_U290 , P1_R1162_U291 , P1_R1162_U292;
wire P1_R1162_U293 , P1_R1162_U294 , P1_R1162_U295 , P1_R1162_U296 , P1_R1162_U297 , P1_R1162_U298 , P1_R1162_U299 , P1_R1162_U300 , P1_R1162_U301 , P1_R1162_U302;
wire P1_R1162_U303 , P1_R1162_U304 , P1_R1162_U305 , P1_R1162_U306 , P1_R1162_U307 , P1_R1162_U308 , P1_R1117_U6 , P1_R1117_U7 , P1_R1117_U8 , P1_R1117_U9;
wire P1_R1117_U10 , P1_R1117_U11 , P1_R1117_U12 , P1_R1117_U13 , P1_R1117_U14 , P1_R1117_U15 , P1_R1117_U16 , P1_R1117_U17 , P1_R1117_U18 , P1_R1117_U19;
wire P1_R1117_U20 , P1_R1117_U21 , P1_R1117_U22 , P1_R1117_U23 , P1_R1117_U24 , P1_R1117_U25 , P1_R1117_U26 , P1_R1117_U27 , P1_R1117_U28 , P1_R1117_U29;
wire P1_R1117_U30 , P1_R1117_U31 , P1_R1117_U32 , P1_R1117_U33 , P1_R1117_U34 , P1_R1117_U35 , P1_R1117_U36 , P1_R1117_U37 , P1_R1117_U38 , P1_R1117_U39;
wire P1_R1117_U40 , P1_R1117_U41 , P1_R1117_U42 , P1_R1117_U43 , P1_R1117_U44 , P1_R1117_U45 , P1_R1117_U46 , P1_R1117_U47 , P1_R1117_U48 , P1_R1117_U49;
wire P1_R1117_U50 , P1_R1117_U51 , P1_R1117_U52 , P1_R1117_U53 , P1_R1117_U54 , P1_R1117_U55 , P1_R1117_U56 , P1_R1117_U57 , P1_R1117_U58 , P1_R1117_U59;
wire P1_R1117_U60 , P1_R1117_U61 , P1_R1117_U62 , P1_R1117_U63 , P1_R1117_U64 , P1_R1117_U65 , P1_R1117_U66 , P1_R1117_U67 , P1_R1117_U68 , P1_R1117_U69;
wire P1_R1117_U70 , P1_R1117_U71 , P1_R1117_U72 , P1_R1117_U73 , P1_R1117_U74 , P1_R1117_U75 , P1_R1117_U76 , P1_R1117_U77 , P1_R1117_U78 , P1_R1117_U79;
wire P1_R1117_U80 , P1_R1117_U81 , P1_R1117_U82 , P1_R1117_U83 , P1_R1117_U84 , P1_R1117_U85 , P1_R1117_U86 , P1_R1117_U87 , P1_R1117_U88 , P1_R1117_U89;
wire P1_R1117_U90 , P1_R1117_U91 , P1_R1117_U92 , P1_R1117_U93 , P1_R1117_U94 , P1_R1117_U95 , P1_R1117_U96 , P1_R1117_U97 , P1_R1117_U98 , P1_R1117_U99;
wire P1_R1117_U100 , P1_R1117_U101 , P1_R1117_U102 , P1_R1117_U103 , P1_R1117_U104 , P1_R1117_U105 , P1_R1117_U106 , P1_R1117_U107 , P1_R1117_U108 , P1_R1117_U109;
wire P1_R1117_U110 , P1_R1117_U111 , P1_R1117_U112 , P1_R1117_U113 , P1_R1117_U114 , P1_R1117_U115 , P1_R1117_U116 , P1_R1117_U117 , P1_R1117_U118 , P1_R1117_U119;
wire P1_R1117_U120 , P1_R1117_U121 , P1_R1117_U122 , P1_R1117_U123 , P1_R1117_U124 , P1_R1117_U125 , P1_R1117_U126 , P1_R1117_U127 , P1_R1117_U128 , P1_R1117_U129;
wire P1_R1117_U130 , P1_R1117_U131 , P1_R1117_U132 , P1_R1117_U133 , P1_R1117_U134 , P1_R1117_U135 , P1_R1117_U136 , P1_R1117_U137 , P1_R1117_U138 , P1_R1117_U139;
wire P1_R1117_U140 , P1_R1117_U141 , P1_R1117_U142 , P1_R1117_U143 , P1_R1117_U144 , P1_R1117_U145 , P1_R1117_U146 , P1_R1117_U147 , P1_R1117_U148 , P1_R1117_U149;
wire P1_R1117_U150 , P1_R1117_U151 , P1_R1117_U152 , P1_R1117_U153 , P1_R1117_U154 , P1_R1117_U155 , P1_R1117_U156 , P1_R1117_U157 , P1_R1117_U158 , P1_R1117_U159;
wire P1_R1117_U160 , P1_R1117_U161 , P1_R1117_U162 , P1_R1117_U163 , P1_R1117_U164 , P1_R1117_U165 , P1_R1117_U166 , P1_R1117_U167 , P1_R1117_U168 , P1_R1117_U169;
wire P1_R1117_U170 , P1_R1117_U171 , P1_R1117_U172 , P1_R1117_U173 , P1_R1117_U174 , P1_R1117_U175 , P1_R1117_U176 , P1_R1117_U177 , P1_R1117_U178 , P1_R1117_U179;
wire P1_R1117_U180 , P1_R1117_U181 , P1_R1117_U182 , P1_R1117_U183 , P1_R1117_U184 , P1_R1117_U185 , P1_R1117_U186 , P1_R1117_U187 , P1_R1117_U188 , P1_R1117_U189;
wire P1_R1117_U190 , P1_R1117_U191 , P1_R1117_U192 , P1_R1117_U193 , P1_R1117_U194 , P1_R1117_U195 , P1_R1117_U196 , P1_R1117_U197 , P1_R1117_U198 , P1_R1117_U199;
wire P1_R1117_U200 , P1_R1117_U201 , P1_R1117_U202 , P1_R1117_U203 , P1_R1117_U204 , P1_R1117_U205 , P1_R1117_U206 , P1_R1117_U207 , P1_R1117_U208 , P1_R1117_U209;
wire P1_R1117_U210 , P1_R1117_U211 , P1_R1117_U212 , P1_R1117_U213 , P1_R1117_U214 , P1_R1117_U215 , P1_R1117_U216 , P1_R1117_U217 , P1_R1117_U218 , P1_R1117_U219;
wire P1_R1117_U220 , P1_R1117_U221 , P1_R1117_U222 , P1_R1117_U223 , P1_R1117_U224 , P1_R1117_U225 , P1_R1117_U226 , P1_R1117_U227 , P1_R1117_U228 , P1_R1117_U229;
wire P1_R1117_U230 , P1_R1117_U231 , P1_R1117_U232 , P1_R1117_U233 , P1_R1117_U234 , P1_R1117_U235 , P1_R1117_U236 , P1_R1117_U237 , P1_R1117_U238 , P1_R1117_U239;
wire P1_R1117_U240 , P1_R1117_U241 , P1_R1117_U242 , P1_R1117_U243 , P1_R1117_U244 , P1_R1117_U245 , P1_R1117_U246 , P1_R1117_U247 , P1_R1117_U248 , P1_R1117_U249;
wire P1_R1117_U250 , P1_R1117_U251 , P1_R1117_U252 , P1_R1117_U253 , P1_R1117_U254 , P1_R1117_U255 , P1_R1117_U256 , P1_R1117_U257 , P1_R1117_U258 , P1_R1117_U259;
wire P1_R1117_U260 , P1_R1117_U261 , P1_R1117_U262 , P1_R1117_U263 , P1_R1117_U264 , P1_R1117_U265 , P1_R1117_U266 , P1_R1117_U267 , P1_R1117_U268 , P1_R1117_U269;
wire P1_R1117_U270 , P1_R1117_U271 , P1_R1117_U272 , P1_R1117_U273 , P1_R1117_U274 , P1_R1117_U275 , P1_R1117_U276 , P1_R1117_U277 , P1_R1117_U278 , P1_R1117_U279;
wire P1_R1117_U280 , P1_R1117_U281 , P1_R1117_U282 , P1_R1117_U283 , P1_R1117_U284 , P1_R1117_U285 , P1_R1117_U286 , P1_R1117_U287 , P1_R1117_U288 , P1_R1117_U289;
wire P1_R1117_U290 , P1_R1117_U291 , P1_R1117_U292 , P1_R1117_U293 , P1_R1117_U294 , P1_R1117_U295 , P1_R1117_U296 , P1_R1117_U297 , P1_R1117_U298 , P1_R1117_U299;
wire P1_R1117_U300 , P1_R1117_U301 , P1_R1117_U302 , P1_R1117_U303 , P1_R1117_U304 , P1_R1117_U305 , P1_R1117_U306 , P1_R1117_U307 , P1_R1117_U308 , P1_R1117_U309;
wire P1_R1117_U310 , P1_R1117_U311 , P1_R1117_U312 , P1_R1117_U313 , P1_R1117_U314 , P1_R1117_U315 , P1_R1117_U316 , P1_R1117_U317 , P1_R1117_U318 , P1_R1117_U319;
wire P1_R1117_U320 , P1_R1117_U321 , P1_R1117_U322 , P1_R1117_U323 , P1_R1117_U324 , P1_R1117_U325 , P1_R1117_U326 , P1_R1117_U327 , P1_R1117_U328 , P1_R1117_U329;
wire P1_R1117_U330 , P1_R1117_U331 , P1_R1117_U332 , P1_R1117_U333 , P1_R1117_U334 , P1_R1117_U335 , P1_R1117_U336 , P1_R1117_U337 , P1_R1117_U338 , P1_R1117_U339;
wire P1_R1117_U340 , P1_R1117_U341 , P1_R1117_U342 , P1_R1117_U343 , P1_R1117_U344 , P1_R1117_U345 , P1_R1117_U346 , P1_R1117_U347 , P1_R1117_U348 , P1_R1117_U349;
wire P1_R1117_U350 , P1_R1117_U351 , P1_R1117_U352 , P1_R1117_U353 , P1_R1117_U354 , P1_R1117_U355 , P1_R1117_U356 , P1_R1117_U357 , P1_R1117_U358 , P1_R1117_U359;
wire P1_R1117_U360 , P1_R1117_U361 , P1_R1117_U362 , P1_R1117_U363 , P1_R1117_U364 , P1_R1117_U365 , P1_R1117_U366 , P1_R1117_U367 , P1_R1117_U368 , P1_R1117_U369;
wire P1_R1117_U370 , P1_R1117_U371 , P1_R1117_U372 , P1_R1117_U373 , P1_R1117_U374 , P1_R1117_U375 , P1_R1117_U376 , P1_R1117_U377 , P1_R1117_U378 , P1_R1117_U379;
wire P1_R1117_U380 , P1_R1117_U381 , P1_R1117_U382 , P1_R1117_U383 , P1_R1117_U384 , P1_R1117_U385 , P1_R1117_U386 , P1_R1117_U387 , P1_R1117_U388 , P1_R1117_U389;
wire P1_R1117_U390 , P1_R1117_U391 , P1_R1117_U392 , P1_R1117_U393 , P1_R1117_U394 , P1_R1117_U395 , P1_R1117_U396 , P1_R1117_U397 , P1_R1117_U398 , P1_R1117_U399;
wire P1_R1117_U400 , P1_R1117_U401 , P1_R1117_U402 , P1_R1117_U403 , P1_R1117_U404 , P1_R1117_U405 , P1_R1117_U406 , P1_R1117_U407 , P1_R1117_U408 , P1_R1117_U409;
wire P1_R1117_U410 , P1_R1117_U411 , P1_R1117_U412 , P1_R1117_U413 , P1_R1117_U414 , P1_R1117_U415 , P1_R1117_U416 , P1_R1117_U417 , P1_R1117_U418 , P1_R1117_U419;
wire P1_R1117_U420 , P1_R1117_U421 , P1_R1117_U422 , P1_R1117_U423 , P1_R1117_U424 , P1_R1117_U425 , P1_R1117_U426 , P1_R1117_U427 , P1_R1117_U428 , P1_R1117_U429;
wire P1_R1117_U430 , P1_R1117_U431 , P1_R1117_U432 , P1_R1117_U433 , P1_R1117_U434 , P1_R1117_U435 , P1_R1117_U436 , P1_R1117_U437 , P1_R1117_U438 , P1_R1117_U439;
wire P1_R1117_U440 , P1_R1117_U441 , P1_R1117_U442 , P1_R1117_U443 , P1_R1117_U444 , P1_R1117_U445 , P1_R1117_U446 , P1_R1117_U447 , P1_R1117_U448 , P1_R1117_U449;
wire P1_R1117_U450 , P1_R1117_U451 , P1_R1117_U452 , P1_R1117_U453 , P1_R1117_U454 , P1_R1117_U455 , P1_R1117_U456 , P1_R1117_U457 , P1_R1117_U458 , P1_R1117_U459;
wire P1_R1117_U460 , P1_R1117_U461 , P1_R1117_U462 , P1_R1117_U463 , P1_R1117_U464 , P1_R1117_U465 , P1_R1117_U466 , P1_R1117_U467 , P1_R1117_U468 , P1_R1117_U469;
wire P1_R1117_U470 , P1_R1117_U471 , P1_R1117_U472 , P1_R1117_U473 , P1_R1375_U6 , P1_R1375_U7 , P1_R1375_U8 , P1_R1375_U9 , P1_R1375_U10 , P1_R1375_U11;
wire P1_R1375_U12 , P1_R1375_U13 , P1_R1375_U14 , P1_R1375_U15 , P1_R1375_U16 , P1_R1375_U17 , P1_R1375_U18 , P1_R1375_U19 , P1_R1375_U20 , P1_R1375_U21;
wire P1_R1375_U22 , P1_R1375_U23 , P1_R1375_U24 , P1_R1375_U25 , P1_R1375_U26 , P1_R1375_U27 , P1_R1375_U28 , P1_R1375_U29 , P1_R1375_U30 , P1_R1375_U31;
wire P1_R1375_U32 , P1_R1375_U33 , P1_R1375_U34 , P1_R1375_U35 , P1_R1375_U36 , P1_R1375_U37 , P1_R1375_U38 , P1_R1375_U39 , P1_R1375_U40 , P1_R1375_U41;
wire P1_R1375_U42 , P1_R1375_U43 , P1_R1375_U44 , P1_R1375_U45 , P1_R1375_U46 , P1_R1375_U47 , P1_R1375_U48 , P1_R1375_U49 , P1_R1375_U50 , P1_R1375_U51;
wire P1_R1375_U52 , P1_R1375_U53 , P1_R1375_U54 , P1_R1375_U55 , P1_R1375_U56 , P1_R1375_U57 , P1_R1375_U58 , P1_R1375_U59 , P1_R1375_U60 , P1_R1375_U61;
wire P1_R1375_U62 , P1_R1375_U63 , P1_R1375_U64 , P1_R1375_U65 , P1_R1375_U66 , P1_R1375_U67 , P1_R1375_U68 , P1_R1375_U69 , P1_R1375_U70 , P1_R1375_U71;
wire P1_R1375_U72 , P1_R1375_U73 , P1_R1375_U74 , P1_R1375_U75 , P1_R1375_U76 , P1_R1375_U77 , P1_R1375_U78 , P1_R1375_U79 , P1_R1375_U80 , P1_R1375_U81;
wire P1_R1375_U82 , P1_R1375_U83 , P1_R1375_U84 , P1_R1375_U85 , P1_R1375_U86 , P1_R1375_U87 , P1_R1375_U88 , P1_R1375_U89 , P1_R1375_U90 , P1_R1375_U91;
wire P1_R1375_U92 , P1_R1375_U93 , P1_R1375_U94 , P1_R1375_U95 , P1_R1375_U96 , P1_R1375_U97 , P1_R1375_U98 , P1_R1375_U99 , P1_R1375_U100 , P1_R1375_U101;
wire P1_R1375_U102 , P1_R1375_U103 , P1_R1375_U104 , P1_R1375_U105 , P1_R1375_U106 , P1_R1375_U107 , P1_R1375_U108 , P1_R1375_U109 , P1_R1375_U110 , P1_R1375_U111;
wire P1_R1375_U112 , P1_R1375_U113 , P1_R1375_U114 , P1_R1375_U115 , P1_R1375_U116 , P1_R1375_U117 , P1_R1375_U118 , P1_R1375_U119 , P1_R1375_U120 , P1_R1375_U121;
wire P1_R1375_U122 , P1_R1375_U123 , P1_R1375_U124 , P1_R1375_U125 , P1_R1375_U126 , P1_R1375_U127 , P1_R1375_U128 , P1_R1375_U129 , P1_R1375_U130 , P1_R1375_U131;
wire P1_R1375_U132 , P1_R1375_U133 , P1_R1375_U134 , P1_R1375_U135 , P1_R1375_U136 , P1_R1375_U137 , P1_R1375_U138 , P1_R1375_U139 , P1_R1375_U140 , P1_R1375_U141;
wire P1_R1375_U142 , P1_R1375_U143 , P1_R1375_U144 , P1_R1375_U145 , P1_R1375_U146 , P1_R1375_U147 , P1_R1375_U148 , P1_R1375_U149 , P1_R1375_U150 , P1_R1375_U151;
wire P1_R1375_U152 , P1_R1375_U153 , P1_R1375_U154 , P1_R1375_U155 , P1_R1375_U156 , P1_R1375_U157 , P1_R1375_U158 , P1_R1375_U159 , P1_R1375_U160 , P1_R1375_U161;
wire P1_R1375_U162 , P1_R1375_U163 , P1_R1375_U164 , P1_R1375_U165 , P1_R1375_U166 , P1_R1375_U167 , P1_R1375_U168 , P1_R1375_U169 , P1_R1375_U170 , P1_R1375_U171;
wire P1_R1375_U172 , P1_R1375_U173 , P1_R1375_U174 , P1_R1375_U175 , P1_R1375_U176 , P1_R1375_U177 , P1_R1375_U178 , P1_R1375_U179 , P1_R1375_U180 , P1_R1375_U181;
wire P1_R1375_U182 , P1_R1375_U183 , P1_R1375_U184 , P1_R1375_U185 , P1_R1375_U186 , P1_R1375_U187 , P1_R1375_U188 , P1_R1375_U189 , P1_R1375_U190 , P1_R1375_U191;
wire P1_R1375_U192 , P1_R1375_U193 , P1_R1375_U194 , P1_R1375_U195 , P1_R1375_U196 , P1_R1375_U197 , P1_R1375_U198 , P1_R1375_U199 , P1_R1375_U200 , P1_R1375_U201;
wire P1_R1375_U202 , P1_R1375_U203 , P1_R1375_U204 , P1_R1375_U205 , P1_R1375_U206 , P1_R1375_U207 , P1_R1352_U6 , P1_R1352_U7 , P1_R1207_U6 , P1_R1207_U7;
wire P1_R1207_U8 , P1_R1207_U9 , P1_R1207_U10 , P1_R1207_U11 , P1_R1207_U12 , P1_R1207_U13 , P1_R1207_U14 , P1_R1207_U15 , P1_R1207_U16 , P1_R1207_U17;
wire P1_R1207_U18 , P1_R1207_U19 , P1_R1207_U20 , P1_R1207_U21 , P1_R1207_U22 , P1_R1207_U23 , P1_R1207_U24 , P1_R1207_U25 , P1_R1207_U26 , P1_R1207_U27;
wire P1_R1207_U28 , P1_R1207_U29 , P1_R1207_U30 , P1_R1207_U31 , P1_R1207_U32 , P1_R1207_U33 , P1_R1207_U34 , P1_R1207_U35 , P1_R1207_U36 , P1_R1207_U37;
wire P1_R1207_U38 , P1_R1207_U39 , P1_R1207_U40 , P1_R1207_U41 , P1_R1207_U42 , P1_R1207_U43 , P1_R1207_U44 , P1_R1207_U45 , P1_R1207_U46 , P1_R1207_U47;
wire P1_R1207_U48 , P1_R1207_U49 , P1_R1207_U50 , P1_R1207_U51 , P1_R1207_U52 , P1_R1207_U53 , P1_R1207_U54 , P1_R1207_U55 , P1_R1207_U56 , P1_R1207_U57;
wire P1_R1207_U58 , P1_R1207_U59 , P1_R1207_U60 , P1_R1207_U61 , P1_R1207_U62 , P1_R1207_U63 , P1_R1207_U64 , P1_R1207_U65 , P1_R1207_U66 , P1_R1207_U67;
wire P1_R1207_U68 , P1_R1207_U69 , P1_R1207_U70 , P1_R1207_U71 , P1_R1207_U72 , P1_R1207_U73 , P1_R1207_U74 , P1_R1207_U75 , P1_R1207_U76 , P1_R1207_U77;
wire P1_R1207_U78 , P1_R1207_U79 , P1_R1207_U80 , P1_R1207_U81 , P1_R1207_U82 , P1_R1207_U83 , P1_R1207_U84 , P1_R1207_U85 , P1_R1207_U86 , P1_R1207_U87;
wire P1_R1207_U88 , P1_R1207_U89 , P1_R1207_U90 , P1_R1207_U91 , P1_R1207_U92 , P1_R1207_U93 , P1_R1207_U94 , P1_R1207_U95 , P1_R1207_U96 , P1_R1207_U97;
wire P1_R1207_U98 , P1_R1207_U99 , P1_R1207_U100 , P1_R1207_U101 , P1_R1207_U102 , P1_R1207_U103 , P1_R1207_U104 , P1_R1207_U105 , P1_R1207_U106 , P1_R1207_U107;
wire P1_R1207_U108 , P1_R1207_U109 , P1_R1207_U110 , P1_R1207_U111 , P1_R1207_U112 , P1_R1207_U113 , P1_R1207_U114 , P1_R1207_U115 , P1_R1207_U116 , P1_R1207_U117;
wire P1_R1207_U118 , P1_R1207_U119 , P1_R1207_U120 , P1_R1207_U121 , P1_R1207_U122 , P1_R1207_U123 , P1_R1207_U124 , P1_R1207_U125 , P1_R1207_U126 , P1_R1207_U127;
wire P1_R1207_U128 , P1_R1207_U129 , P1_R1207_U130 , P1_R1207_U131 , P1_R1207_U132 , P1_R1207_U133 , P1_R1207_U134 , P1_R1207_U135 , P1_R1207_U136 , P1_R1207_U137;
wire P1_R1207_U138 , P1_R1207_U139 , P1_R1207_U140 , P1_R1207_U141 , P1_R1207_U142 , P1_R1207_U143 , P1_R1207_U144 , P1_R1207_U145 , P1_R1207_U146 , P1_R1207_U147;
wire P1_R1207_U148 , P1_R1207_U149 , P1_R1207_U150 , P1_R1207_U151 , P1_R1207_U152 , P1_R1207_U153 , P1_R1207_U154 , P1_R1207_U155 , P1_R1207_U156 , P1_R1207_U157;
wire P1_R1207_U158 , P1_R1207_U159 , P1_R1207_U160 , P1_R1207_U161 , P1_R1207_U162 , P1_R1207_U163 , P1_R1207_U164 , P1_R1207_U165 , P1_R1207_U166 , P1_R1207_U167;
wire P1_R1207_U168 , P1_R1207_U169 , P1_R1207_U170 , P1_R1207_U171 , P1_R1207_U172 , P1_R1207_U173 , P1_R1207_U174 , P1_R1207_U175 , P1_R1207_U176 , P1_R1207_U177;
wire P1_R1207_U178 , P1_R1207_U179 , P1_R1207_U180 , P1_R1207_U181 , P1_R1207_U182 , P1_R1207_U183 , P1_R1207_U184 , P1_R1207_U185 , P1_R1207_U186 , P1_R1207_U187;
wire P1_R1207_U188 , P1_R1207_U189 , P1_R1207_U190 , P1_R1207_U191 , P1_R1207_U192 , P1_R1207_U193 , P1_R1207_U194 , P1_R1207_U195 , P1_R1207_U196 , P1_R1207_U197;
wire P1_R1207_U198 , P1_R1207_U199 , P1_R1207_U200 , P1_R1207_U201 , P1_R1207_U202 , P1_R1207_U203 , P1_R1207_U204 , P1_R1207_U205 , P1_R1207_U206 , P1_R1207_U207;
wire P1_R1207_U208 , P1_R1207_U209 , P1_R1207_U210 , P1_R1207_U211 , P1_R1207_U212 , P1_R1207_U213 , P1_R1207_U214 , P1_R1207_U215 , P1_R1207_U216 , P1_R1207_U217;
wire P1_R1207_U218 , P1_R1207_U219 , P1_R1207_U220 , P1_R1207_U221 , P1_R1207_U222 , P1_R1207_U223 , P1_R1207_U224 , P1_R1207_U225 , P1_R1207_U226 , P1_R1207_U227;
wire P1_R1207_U228 , P1_R1207_U229 , P1_R1207_U230 , P1_R1207_U231 , P1_R1207_U232 , P1_R1207_U233 , P1_R1207_U234 , P1_R1207_U235 , P1_R1207_U236 , P1_R1207_U237;
wire P1_R1207_U238 , P1_R1207_U239 , P1_R1207_U240 , P1_R1207_U241 , P1_R1207_U242 , P1_R1207_U243 , P1_R1207_U244 , P1_R1207_U245 , P1_R1207_U246 , P1_R1207_U247;
wire P1_R1207_U248 , P1_R1207_U249 , P1_R1207_U250 , P1_R1207_U251 , P1_R1207_U252 , P1_R1207_U253 , P1_R1207_U254 , P1_R1207_U255 , P1_R1207_U256 , P1_R1207_U257;
wire P1_R1207_U258 , P1_R1207_U259 , P1_R1207_U260 , P1_R1207_U261 , P1_R1207_U262 , P1_R1207_U263 , P1_R1207_U264 , P1_R1207_U265 , P1_R1207_U266 , P1_R1207_U267;
wire P1_R1207_U268 , P1_R1207_U269 , P1_R1207_U270 , P1_R1207_U271 , P1_R1207_U272 , P1_R1207_U273 , P1_R1207_U274 , P1_R1207_U275 , P1_R1207_U276 , P1_R1207_U277;
wire P1_R1207_U278 , P1_R1207_U279 , P1_R1207_U280 , P1_R1207_U281 , P1_R1207_U282 , P1_R1207_U283 , P1_R1207_U284 , P1_R1207_U285 , P1_R1207_U286 , P1_R1207_U287;
wire P1_R1207_U288 , P1_R1207_U289 , P1_R1207_U290 , P1_R1207_U291 , P1_R1207_U292 , P1_R1207_U293 , P1_R1207_U294 , P1_R1207_U295 , P1_R1207_U296 , P1_R1207_U297;
wire P1_R1207_U298 , P1_R1207_U299 , P1_R1207_U300 , P1_R1207_U301 , P1_R1207_U302 , P1_R1207_U303 , P1_R1207_U304 , P1_R1207_U305 , P1_R1207_U306 , P1_R1207_U307;
wire P1_R1207_U308 , P1_R1207_U309 , P1_R1207_U310 , P1_R1207_U311 , P1_R1207_U312 , P1_R1207_U313 , P1_R1207_U314 , P1_R1207_U315 , P1_R1207_U316 , P1_R1207_U317;
wire P1_R1207_U318 , P1_R1207_U319 , P1_R1207_U320 , P1_R1207_U321 , P1_R1207_U322 , P1_R1207_U323 , P1_R1207_U324 , P1_R1207_U325 , P1_R1207_U326 , P1_R1207_U327;
wire P1_R1207_U328 , P1_R1207_U329 , P1_R1207_U330 , P1_R1207_U331 , P1_R1207_U332 , P1_R1207_U333 , P1_R1207_U334 , P1_R1207_U335 , P1_R1207_U336 , P1_R1207_U337;
wire P1_R1207_U338 , P1_R1207_U339 , P1_R1207_U340 , P1_R1207_U341 , P1_R1207_U342 , P1_R1207_U343 , P1_R1207_U344 , P1_R1207_U345 , P1_R1207_U346 , P1_R1207_U347;
wire P1_R1207_U348 , P1_R1207_U349 , P1_R1207_U350 , P1_R1207_U351 , P1_R1207_U352 , P1_R1207_U353 , P1_R1207_U354 , P1_R1207_U355 , P1_R1207_U356 , P1_R1207_U357;
wire P1_R1207_U358 , P1_R1207_U359 , P1_R1207_U360 , P1_R1207_U361 , P1_R1207_U362 , P1_R1207_U363 , P1_R1207_U364 , P1_R1207_U365 , P1_R1207_U366 , P1_R1207_U367;
wire P1_R1207_U368 , P1_R1207_U369 , P1_R1207_U370 , P1_R1207_U371 , P1_R1207_U372 , P1_R1207_U373 , P1_R1207_U374 , P1_R1207_U375 , P1_R1207_U376 , P1_R1207_U377;
wire P1_R1207_U378 , P1_R1207_U379 , P1_R1207_U380 , P1_R1207_U381 , P1_R1207_U382 , P1_R1207_U383 , P1_R1207_U384 , P1_R1207_U385 , P1_R1207_U386 , P1_R1207_U387;
wire P1_R1207_U388 , P1_R1207_U389 , P1_R1207_U390 , P1_R1207_U391 , P1_R1207_U392 , P1_R1207_U393 , P1_R1207_U394 , P1_R1207_U395 , P1_R1207_U396 , P1_R1207_U397;
wire P1_R1207_U398 , P1_R1207_U399 , P1_R1207_U400 , P1_R1207_U401 , P1_R1207_U402 , P1_R1207_U403 , P1_R1207_U404 , P1_R1207_U405 , P1_R1207_U406 , P1_R1207_U407;
wire P1_R1207_U408 , P1_R1207_U409 , P1_R1207_U410 , P1_R1207_U411 , P1_R1207_U412 , P1_R1207_U413 , P1_R1207_U414 , P1_R1207_U415 , P1_R1207_U416 , P1_R1207_U417;
wire P1_R1207_U418 , P1_R1207_U419 , P1_R1207_U420 , P1_R1207_U421 , P1_R1207_U422 , P1_R1207_U423 , P1_R1207_U424 , P1_R1207_U425 , P1_R1207_U426 , P1_R1207_U427;
wire P1_R1207_U428 , P1_R1207_U429 , P1_R1207_U430 , P1_R1207_U431 , P1_R1207_U432 , P1_R1207_U433 , P1_R1207_U434 , P1_R1207_U435 , P1_R1207_U436 , P1_R1207_U437;
wire P1_R1207_U438 , P1_R1207_U439 , P1_R1207_U440 , P1_R1207_U441 , P1_R1207_U442 , P1_R1207_U443 , P1_R1207_U444 , P1_R1207_U445 , P1_R1207_U446 , P1_R1207_U447;
wire P1_R1207_U448 , P1_R1207_U449 , P1_R1207_U450 , P1_R1207_U451 , P1_R1207_U452 , P1_R1207_U453 , P1_R1207_U454 , P1_R1207_U455 , P1_R1207_U456 , P1_R1207_U457;
wire P1_R1207_U458 , P1_R1207_U459 , P1_R1207_U460 , P1_R1207_U461 , P1_R1207_U462 , P1_R1207_U463 , P1_R1207_U464 , P1_R1207_U465 , P1_R1207_U466 , P1_R1207_U467;
wire P1_R1207_U468 , P1_R1207_U469 , P1_R1207_U470 , P1_R1207_U471 , P1_R1207_U472 , P1_R1207_U473 , P1_R1165_U4 , P1_R1165_U5 , P1_R1165_U6 , P1_R1165_U7;
wire P1_R1165_U8 , P1_R1165_U9 , P1_R1165_U10 , P1_R1165_U11 , P1_R1165_U12 , P1_R1165_U13 , P1_R1165_U14 , P1_R1165_U15 , P1_R1165_U16 , P1_R1165_U17;
wire P1_R1165_U18 , P1_R1165_U19 , P1_R1165_U20 , P1_R1165_U21 , P1_R1165_U22 , P1_R1165_U23 , P1_R1165_U24 , P1_R1165_U25 , P1_R1165_U26 , P1_R1165_U27;
wire P1_R1165_U28 , P1_R1165_U29 , P1_R1165_U30 , P1_R1165_U31 , P1_R1165_U32 , P1_R1165_U33 , P1_R1165_U34 , P1_R1165_U35 , P1_R1165_U36 , P1_R1165_U37;
wire P1_R1165_U38 , P1_R1165_U39 , P1_R1165_U40 , P1_R1165_U41 , P1_R1165_U42 , P1_R1165_U43 , P1_R1165_U44 , P1_R1165_U45 , P1_R1165_U46 , P1_R1165_U47;
wire P1_R1165_U48 , P1_R1165_U49 , P1_R1165_U50 , P1_R1165_U51 , P1_R1165_U52 , P1_R1165_U53 , P1_R1165_U54 , P1_R1165_U55 , P1_R1165_U56 , P1_R1165_U57;
wire P1_R1165_U58 , P1_R1165_U59 , P1_R1165_U60 , P1_R1165_U61 , P1_R1165_U62 , P1_R1165_U63 , P1_R1165_U64 , P1_R1165_U65 , P1_R1165_U66 , P1_R1165_U67;
wire P1_R1165_U68 , P1_R1165_U69 , P1_R1165_U70 , P1_R1165_U71 , P1_R1165_U72 , P1_R1165_U73 , P1_R1165_U74 , P1_R1165_U75 , P1_R1165_U76 , P1_R1165_U77;
wire P1_R1165_U78 , P1_R1165_U79 , P1_R1165_U80 , P1_R1165_U81 , P1_R1165_U82 , P1_R1165_U83 , P1_R1165_U84 , P1_R1165_U85 , P1_R1165_U86 , P1_R1165_U87;
wire P1_R1165_U88 , P1_R1165_U89 , P1_R1165_U90 , P1_R1165_U91 , P1_R1165_U92 , P1_R1165_U93 , P1_R1165_U94 , P1_R1165_U95 , P1_R1165_U96 , P1_R1165_U97;
wire P1_R1165_U98 , P1_R1165_U99 , P1_R1165_U100 , P1_R1165_U101 , P1_R1165_U102 , P1_R1165_U103 , P1_R1165_U104 , P1_R1165_U105 , P1_R1165_U106 , P1_R1165_U107;
wire P1_R1165_U108 , P1_R1165_U109 , P1_R1165_U110 , P1_R1165_U111 , P1_R1165_U112 , P1_R1165_U113 , P1_R1165_U114 , P1_R1165_U115 , P1_R1165_U116 , P1_R1165_U117;
wire P1_R1165_U118 , P1_R1165_U119 , P1_R1165_U120 , P1_R1165_U121 , P1_R1165_U122 , P1_R1165_U123 , P1_R1165_U124 , P1_R1165_U125 , P1_R1165_U126 , P1_R1165_U127;
wire P1_R1165_U128 , P1_R1165_U129 , P1_R1165_U130 , P1_R1165_U131 , P1_R1165_U132 , P1_R1165_U133 , P1_R1165_U134 , P1_R1165_U135 , P1_R1165_U136 , P1_R1165_U137;
wire P1_R1165_U138 , P1_R1165_U139 , P1_R1165_U140 , P1_R1165_U141 , P1_R1165_U142 , P1_R1165_U143 , P1_R1165_U144 , P1_R1165_U145 , P1_R1165_U146 , P1_R1165_U147;
wire P1_R1165_U148 , P1_R1165_U149 , P1_R1165_U150 , P1_R1165_U151 , P1_R1165_U152 , P1_R1165_U153 , P1_R1165_U154 , P1_R1165_U155 , P1_R1165_U156 , P1_R1165_U157;
wire P1_R1165_U158 , P1_R1165_U159 , P1_R1165_U160 , P1_R1165_U161 , P1_R1165_U162 , P1_R1165_U163 , P1_R1165_U164 , P1_R1165_U165 , P1_R1165_U166 , P1_R1165_U167;
wire P1_R1165_U168 , P1_R1165_U169 , P1_R1165_U170 , P1_R1165_U171 , P1_R1165_U172 , P1_R1165_U173 , P1_R1165_U174 , P1_R1165_U175 , P1_R1165_U176 , P1_R1165_U177;
wire P1_R1165_U178 , P1_R1165_U179 , P1_R1165_U180 , P1_R1165_U181 , P1_R1165_U182 , P1_R1165_U183 , P1_R1165_U184 , P1_R1165_U185 , P1_R1165_U186 , P1_R1165_U187;
wire P1_R1165_U188 , P1_R1165_U189 , P1_R1165_U190 , P1_R1165_U191 , P1_R1165_U192 , P1_R1165_U193 , P1_R1165_U194 , P1_R1165_U195 , P1_R1165_U196 , P1_R1165_U197;
wire P1_R1165_U198 , P1_R1165_U199 , P1_R1165_U200 , P1_R1165_U201 , P1_R1165_U202 , P1_R1165_U203 , P1_R1165_U204 , P1_R1165_U205 , P1_R1165_U206 , P1_R1165_U207;
wire P1_R1165_U208 , P1_R1165_U209 , P1_R1165_U210 , P1_R1165_U211 , P1_R1165_U212 , P1_R1165_U213 , P1_R1165_U214 , P1_R1165_U215 , P1_R1165_U216 , P1_R1165_U217;
wire P1_R1165_U218 , P1_R1165_U219 , P1_R1165_U220 , P1_R1165_U221 , P1_R1165_U222 , P1_R1165_U223 , P1_R1165_U224 , P1_R1165_U225 , P1_R1165_U226 , P1_R1165_U227;
wire P1_R1165_U228 , P1_R1165_U229 , P1_R1165_U230 , P1_R1165_U231 , P1_R1165_U232 , P1_R1165_U233 , P1_R1165_U234 , P1_R1165_U235 , P1_R1165_U236 , P1_R1165_U237;
wire P1_R1165_U238 , P1_R1165_U239 , P1_R1165_U240 , P1_R1165_U241 , P1_R1165_U242 , P1_R1165_U243 , P1_R1165_U244 , P1_R1165_U245 , P1_R1165_U246 , P1_R1165_U247;
wire P1_R1165_U248 , P1_R1165_U249 , P1_R1165_U250 , P1_R1165_U251 , P1_R1165_U252 , P1_R1165_U253 , P1_R1165_U254 , P1_R1165_U255 , P1_R1165_U256 , P1_R1165_U257;
wire P1_R1165_U258 , P1_R1165_U259 , P1_R1165_U260 , P1_R1165_U261 , P1_R1165_U262 , P1_R1165_U263 , P1_R1165_U264 , P1_R1165_U265 , P1_R1165_U266 , P1_R1165_U267;
wire P1_R1165_U268 , P1_R1165_U269 , P1_R1165_U270 , P1_R1165_U271 , P1_R1165_U272 , P1_R1165_U273 , P1_R1165_U274 , P1_R1165_U275 , P1_R1165_U276 , P1_R1165_U277;
wire P1_R1165_U278 , P1_R1165_U279 , P1_R1165_U280 , P1_R1165_U281 , P1_R1165_U282 , P1_R1165_U283 , P1_R1165_U284 , P1_R1165_U285 , P1_R1165_U286 , P1_R1165_U287;
wire P1_R1165_U288 , P1_R1165_U289 , P1_R1165_U290 , P1_R1165_U291 , P1_R1165_U292 , P1_R1165_U293 , P1_R1165_U294 , P1_R1165_U295 , P1_R1165_U296 , P1_R1165_U297;
wire P1_R1165_U298 , P1_R1165_U299 , P1_R1165_U300 , P1_R1165_U301 , P1_R1165_U302 , P1_R1165_U303 , P1_R1165_U304 , P1_R1165_U305 , P1_R1165_U306 , P1_R1165_U307;
wire P1_R1165_U308 , P1_R1165_U309 , P1_R1165_U310 , P1_R1165_U311 , P1_R1165_U312 , P1_R1165_U313 , P1_R1165_U314 , P1_R1165_U315 , P1_R1165_U316 , P1_R1165_U317;
wire P1_R1165_U318 , P1_R1165_U319 , P1_R1165_U320 , P1_R1165_U321 , P1_R1165_U322 , P1_R1165_U323 , P1_R1165_U324 , P1_R1165_U325 , P1_R1165_U326 , P1_R1165_U327;
wire P1_R1165_U328 , P1_R1165_U329 , P1_R1165_U330 , P1_R1165_U331 , P1_R1165_U332 , P1_R1165_U333 , P1_R1165_U334 , P1_R1165_U335 , P1_R1165_U336 , P1_R1165_U337;
wire P1_R1165_U338 , P1_R1165_U339 , P1_R1165_U340 , P1_R1165_U341 , P1_R1165_U342 , P1_R1165_U343 , P1_R1165_U344 , P1_R1165_U345 , P1_R1165_U346 , P1_R1165_U347;
wire P1_R1165_U348 , P1_R1165_U349 , P1_R1165_U350 , P1_R1165_U351 , P1_R1165_U352 , P1_R1165_U353 , P1_R1165_U354 , P1_R1165_U355 , P1_R1165_U356 , P1_R1165_U357;
wire P1_R1165_U358 , P1_R1165_U359 , P1_R1165_U360 , P1_R1165_U361 , P1_R1165_U362 , P1_R1165_U363 , P1_R1165_U364 , P1_R1165_U365 , P1_R1165_U366 , P1_R1165_U367;
wire P1_R1165_U368 , P1_R1165_U369 , P1_R1165_U370 , P1_R1165_U371 , P1_R1165_U372 , P1_R1165_U373 , P1_R1165_U374 , P1_R1165_U375 , P1_R1165_U376 , P1_R1165_U377;
wire P1_R1165_U378 , P1_R1165_U379 , P1_R1165_U380 , P1_R1165_U381 , P1_R1165_U382 , P1_R1165_U383 , P1_R1165_U384 , P1_R1165_U385 , P1_R1165_U386 , P1_R1165_U387;
wire P1_R1165_U388 , P1_R1165_U389 , P1_R1165_U390 , P1_R1165_U391 , P1_R1165_U392 , P1_R1165_U393 , P1_R1165_U394 , P1_R1165_U395 , P1_R1165_U396 , P1_R1165_U397;
wire P1_R1165_U398 , P1_R1165_U399 , P1_R1165_U400 , P1_R1165_U401 , P1_R1165_U402 , P1_R1165_U403 , P1_R1165_U404 , P1_R1165_U405 , P1_R1165_U406 , P1_R1165_U407;
wire P1_R1165_U408 , P1_R1165_U409 , P1_R1165_U410 , P1_R1165_U411 , P1_R1165_U412 , P1_R1165_U413 , P1_R1165_U414 , P1_R1165_U415 , P1_R1165_U416 , P1_R1165_U417;
wire P1_R1165_U418 , P1_R1165_U419 , P1_R1165_U420 , P1_R1165_U421 , P1_R1165_U422 , P1_R1165_U423 , P1_R1165_U424 , P1_R1165_U425 , P1_R1165_U426 , P1_R1165_U427;
wire P1_R1165_U428 , P1_R1165_U429 , P1_R1165_U430 , P1_R1165_U431 , P1_R1165_U432 , P1_R1165_U433 , P1_R1165_U434 , P1_R1165_U435 , P1_R1165_U436 , P1_R1165_U437;
wire P1_R1165_U438 , P1_R1165_U439 , P1_R1165_U440 , P1_R1165_U441 , P1_R1165_U442 , P1_R1165_U443 , P1_R1165_U444 , P1_R1165_U445 , P1_R1165_U446 , P1_R1165_U447;
wire P1_R1165_U448 , P1_R1165_U449 , P1_R1165_U450 , P1_R1165_U451 , P1_R1165_U452 , P1_R1165_U453 , P1_R1165_U454 , P1_R1165_U455 , P1_R1165_U456 , P1_R1165_U457;
wire P1_R1165_U458 , P1_R1165_U459 , P1_R1165_U460 , P1_R1165_U461 , P1_R1165_U462 , P1_R1165_U463 , P1_R1165_U464 , P1_R1165_U465 , P1_R1165_U466 , P1_R1165_U467;
wire P1_R1165_U468 , P1_R1165_U469 , P1_R1165_U470 , P1_R1165_U471 , P1_R1165_U472 , P1_R1165_U473 , P1_R1165_U474 , P1_R1165_U475 , P1_R1165_U476 , P1_R1165_U477;
wire P1_R1165_U478 , P1_R1165_U479 , P1_R1165_U480 , P1_R1165_U481 , P1_R1165_U482 , P1_R1165_U483 , P1_R1165_U484 , P1_R1165_U485 , P1_R1165_U486 , P1_R1165_U487;
wire P1_R1165_U488 , P1_R1165_U489 , P1_R1165_U490 , P1_R1165_U491 , P1_R1165_U492 , P1_R1165_U493 , P1_R1165_U494 , P1_R1165_U495 , P1_R1165_U496 , P1_R1165_U497;
wire P1_R1165_U498 , P1_R1165_U499 , P1_R1165_U500 , P1_R1165_U501 , P1_R1165_U502 , P1_R1165_U503 , P1_R1165_U504 , P1_R1165_U505 , P1_R1165_U506 , P1_R1165_U507;
wire P1_R1165_U508 , P1_R1165_U509 , P1_R1165_U510 , P1_R1165_U511 , P1_R1165_U512 , P1_R1165_U513 , P1_R1165_U514 , P1_R1165_U515 , P1_R1165_U516 , P1_R1165_U517;
wire P1_R1165_U518 , P1_R1165_U519 , P1_R1165_U520 , P1_R1165_U521 , P1_R1165_U522 , P1_R1165_U523 , P1_R1165_U524 , P1_R1165_U525 , P1_R1165_U526 , P1_R1165_U527;
wire P1_R1165_U528 , P1_R1165_U529 , P1_R1165_U530 , P1_R1165_U531 , P1_R1165_U532 , P1_R1165_U533 , P1_R1165_U534 , P1_R1165_U535 , P1_R1165_U536 , P1_R1165_U537;
wire P1_R1165_U538 , P1_R1165_U539 , P1_R1165_U540 , P1_R1165_U541 , P1_R1165_U542 , P1_R1165_U543 , P1_R1165_U544 , P1_R1165_U545 , P1_R1165_U546 , P1_R1165_U547;
wire P1_R1165_U548 , P1_R1165_U549 , P1_R1165_U550 , P1_R1165_U551 , P1_R1165_U552 , P1_R1165_U553 , P1_R1165_U554 , P1_R1165_U555 , P1_R1165_U556 , P1_R1165_U557;
wire P1_R1165_U558 , P1_R1165_U559 , P1_R1165_U560 , P1_R1165_U561 , P1_R1165_U562 , P1_R1165_U563 , P1_R1165_U564 , P1_R1165_U565 , P1_R1165_U566 , P1_R1165_U567;
wire P1_R1165_U568 , P1_R1165_U569 , P1_R1165_U570 , P1_R1165_U571 , P1_R1165_U572 , P1_R1165_U573 , P1_R1165_U574 , P1_R1165_U575 , P1_R1165_U576 , P1_R1165_U577;
wire P1_R1165_U578 , P1_R1165_U579 , P1_R1165_U580 , P1_R1165_U581 , P1_R1165_U582 , P1_R1165_U583 , P1_R1165_U584 , P1_R1165_U585 , P1_R1165_U586 , P1_R1165_U587;
wire P1_R1165_U588 , P1_R1165_U589 , P1_R1165_U590 , P1_R1165_U591 , P1_R1165_U592 , P1_R1165_U593 , P1_R1165_U594 , P1_R1165_U595 , P1_R1165_U596 , P1_R1165_U597;
wire P1_R1165_U598 , P1_R1165_U599 , P1_R1165_U600 , P1_R1165_U601 , P1_R1165_U602 , P1_R1150_U6 , P1_R1150_U7 , P1_R1150_U8 , P1_R1150_U9 , P1_R1150_U10;
wire P1_R1150_U11 , P1_R1150_U12 , P1_R1150_U13 , P1_R1150_U14 , P1_R1150_U15 , P1_R1150_U16 , P1_R1150_U17 , P1_R1150_U18 , P1_R1150_U19 , P1_R1150_U20;
wire P1_R1150_U21 , P1_R1150_U22 , P1_R1150_U23 , P1_R1150_U24 , P1_R1150_U25 , P1_R1150_U26 , P1_R1150_U27 , P1_R1150_U28 , P1_R1150_U29 , P1_R1150_U30;
wire P1_R1150_U31 , P1_R1150_U32 , P1_R1150_U33 , P1_R1150_U34 , P1_R1150_U35 , P1_R1150_U36 , P1_R1150_U37 , P1_R1150_U38 , P1_R1150_U39 , P1_R1150_U40;
wire P1_R1150_U41 , P1_R1150_U42 , P1_R1150_U43 , P1_R1150_U44 , P1_R1150_U45 , P1_R1150_U46 , P1_R1150_U47 , P1_R1150_U48 , P1_R1150_U49 , P1_R1150_U50;
wire P1_R1150_U51 , P1_R1150_U52 , P1_R1150_U53 , P1_R1150_U54 , P1_R1150_U55 , P1_R1150_U56 , P1_R1150_U57 , P1_R1150_U58 , P1_R1150_U59 , P1_R1150_U60;
wire P1_R1150_U61 , P1_R1150_U62 , P1_R1150_U63 , P1_R1150_U64 , P1_R1150_U65 , P1_R1150_U66 , P1_R1150_U67 , P1_R1150_U68 , P1_R1150_U69 , P1_R1150_U70;
wire P1_R1150_U71 , P1_R1150_U72 , P1_R1150_U73 , P1_R1150_U74 , P1_R1150_U75 , P1_R1150_U76 , P1_R1150_U77 , P1_R1150_U78 , P1_R1150_U79 , P1_R1150_U80;
wire P1_R1150_U81 , P1_R1150_U82 , P1_R1150_U83 , P1_R1150_U84 , P1_R1150_U85 , P1_R1150_U86 , P1_R1150_U87 , P1_R1150_U88 , P1_R1150_U89 , P1_R1150_U90;
wire P1_R1150_U91 , P1_R1150_U92 , P1_R1150_U93 , P1_R1150_U94 , P1_R1150_U95 , P1_R1150_U96 , P1_R1150_U97 , P1_R1150_U98 , P1_R1150_U99 , P1_R1150_U100;
wire P1_R1150_U101 , P1_R1150_U102 , P1_R1150_U103 , P1_R1150_U104 , P1_R1150_U105 , P1_R1150_U106 , P1_R1150_U107 , P1_R1150_U108 , P1_R1150_U109 , P1_R1150_U110;
wire P1_R1150_U111 , P1_R1150_U112 , P1_R1150_U113 , P1_R1150_U114 , P1_R1150_U115 , P1_R1150_U116 , P1_R1150_U117 , P1_R1150_U118 , P1_R1150_U119 , P1_R1150_U120;
wire P1_R1150_U121 , P1_R1150_U122 , P1_R1150_U123 , P1_R1150_U124 , P1_R1150_U125 , P1_R1150_U126 , P1_R1150_U127 , P1_R1150_U128 , P1_R1150_U129 , P1_R1150_U130;
wire P1_R1150_U131 , P1_R1150_U132 , P1_R1150_U133 , P1_R1150_U134 , P1_R1150_U135 , P1_R1150_U136 , P1_R1150_U137 , P1_R1150_U138 , P1_R1150_U139 , P1_R1150_U140;
wire P1_R1150_U141 , P1_R1150_U142 , P1_R1150_U143 , P1_R1150_U144 , P1_R1150_U145 , P1_R1150_U146 , P1_R1150_U147 , P1_R1150_U148 , P1_R1150_U149 , P1_R1150_U150;
wire P1_R1150_U151 , P1_R1150_U152 , P1_R1150_U153 , P1_R1150_U154 , P1_R1150_U155 , P1_R1150_U156 , P1_R1150_U157 , P1_R1150_U158 , P1_R1150_U159 , P1_R1150_U160;
wire P1_R1150_U161 , P1_R1150_U162 , P1_R1150_U163 , P1_R1150_U164 , P1_R1150_U165 , P1_R1150_U166 , P1_R1150_U167 , P1_R1150_U168 , P1_R1150_U169 , P1_R1150_U170;
wire P1_R1150_U171 , P1_R1150_U172 , P1_R1150_U173 , P1_R1150_U174 , P1_R1150_U175 , P1_R1150_U176 , P1_R1150_U177 , P1_R1150_U178 , P1_R1150_U179 , P1_R1150_U180;
wire P1_R1150_U181 , P1_R1150_U182 , P1_R1150_U183 , P1_R1150_U184 , P1_R1150_U185 , P1_R1150_U186 , P1_R1150_U187 , P1_R1150_U188 , P1_R1150_U189 , P1_R1150_U190;
wire P1_R1150_U191 , P1_R1150_U192 , P1_R1150_U193 , P1_R1150_U194 , P1_R1150_U195 , P1_R1150_U196 , P1_R1150_U197 , P1_R1150_U198 , P1_R1150_U199 , P1_R1150_U200;
wire P1_R1150_U201 , P1_R1150_U202 , P1_R1150_U203 , P1_R1150_U204 , P1_R1150_U205 , P1_R1150_U206 , P1_R1150_U207 , P1_R1150_U208 , P1_R1150_U209 , P1_R1150_U210;
wire P1_R1150_U211 , P1_R1150_U212 , P1_R1150_U213 , P1_R1150_U214 , P1_R1150_U215 , P1_R1150_U216 , P1_R1150_U217 , P1_R1150_U218 , P1_R1150_U219 , P1_R1150_U220;
wire P1_R1150_U221 , P1_R1150_U222 , P1_R1150_U223 , P1_R1150_U224 , P1_R1150_U225 , P1_R1150_U226 , P1_R1150_U227 , P1_R1150_U228 , P1_R1150_U229 , P1_R1150_U230;
wire P1_R1150_U231 , P1_R1150_U232 , P1_R1150_U233 , P1_R1150_U234 , P1_R1150_U235 , P1_R1150_U236 , P1_R1150_U237 , P1_R1150_U238 , P1_R1150_U239 , P1_R1150_U240;
wire P1_R1150_U241 , P1_R1150_U242 , P1_R1150_U243 , P1_R1150_U244 , P1_R1150_U245 , P1_R1150_U246 , P1_R1150_U247 , P1_R1150_U248 , P1_R1150_U249 , P1_R1150_U250;
wire P1_R1150_U251 , P1_R1150_U252 , P1_R1150_U253 , P1_R1150_U254 , P1_R1150_U255 , P1_R1150_U256 , P1_R1150_U257 , P1_R1150_U258 , P1_R1150_U259 , P1_R1150_U260;
wire P1_R1150_U261 , P1_R1150_U262 , P1_R1150_U263 , P1_R1150_U264 , P1_R1150_U265 , P1_R1150_U266 , P1_R1150_U267 , P1_R1150_U268 , P1_R1150_U269 , P1_R1150_U270;
wire P1_R1150_U271 , P1_R1150_U272 , P1_R1150_U273 , P1_R1150_U274 , P1_R1150_U275 , P1_R1150_U276 , P1_R1150_U277 , P1_R1150_U278 , P1_R1150_U279 , P1_R1150_U280;
wire P1_R1150_U281 , P1_R1150_U282 , P1_R1150_U283 , P1_R1150_U284 , P1_R1150_U285 , P1_R1150_U286 , P1_R1150_U287 , P1_R1150_U288 , P1_R1150_U289 , P1_R1150_U290;
wire P1_R1150_U291 , P1_R1150_U292 , P1_R1150_U293 , P1_R1150_U294 , P1_R1150_U295 , P1_R1150_U296 , P1_R1150_U297 , P1_R1150_U298 , P1_R1150_U299 , P1_R1150_U300;
wire P1_R1150_U301 , P1_R1150_U302 , P1_R1150_U303 , P1_R1150_U304 , P1_R1150_U305 , P1_R1150_U306 , P1_R1150_U307 , P1_R1150_U308 , P1_R1150_U309 , P1_R1150_U310;
wire P1_R1150_U311 , P1_R1150_U312 , P1_R1150_U313 , P1_R1150_U314 , P1_R1150_U315 , P1_R1150_U316 , P1_R1150_U317 , P1_R1150_U318 , P1_R1150_U319 , P1_R1150_U320;
wire P1_R1150_U321 , P1_R1150_U322 , P1_R1150_U323 , P1_R1150_U324 , P1_R1150_U325 , P1_R1150_U326 , P1_R1150_U327 , P1_R1150_U328 , P1_R1150_U329 , P1_R1150_U330;
wire P1_R1150_U331 , P1_R1150_U332 , P1_R1150_U333 , P1_R1150_U334 , P1_R1150_U335 , P1_R1150_U336 , P1_R1150_U337 , P1_R1150_U338 , P1_R1150_U339 , P1_R1150_U340;
wire P1_R1150_U341 , P1_R1150_U342 , P1_R1150_U343 , P1_R1150_U344 , P1_R1150_U345 , P1_R1150_U346 , P1_R1150_U347 , P1_R1150_U348 , P1_R1150_U349 , P1_R1150_U350;
wire P1_R1150_U351 , P1_R1150_U352 , P1_R1150_U353 , P1_R1150_U354 , P1_R1150_U355 , P1_R1150_U356 , P1_R1150_U357 , P1_R1150_U358 , P1_R1150_U359 , P1_R1150_U360;
wire P1_R1150_U361 , P1_R1150_U362 , P1_R1150_U363 , P1_R1150_U364 , P1_R1150_U365 , P1_R1150_U366 , P1_R1150_U367 , P1_R1150_U368 , P1_R1150_U369 , P1_R1150_U370;
wire P1_R1150_U371 , P1_R1150_U372 , P1_R1150_U373 , P1_R1150_U374 , P1_R1150_U375 , P1_R1150_U376 , P1_R1150_U377 , P1_R1150_U378 , P1_R1150_U379 , P1_R1150_U380;
wire P1_R1150_U381 , P1_R1150_U382 , P1_R1150_U383 , P1_R1150_U384 , P1_R1150_U385 , P1_R1150_U386 , P1_R1150_U387 , P1_R1150_U388 , P1_R1150_U389 , P1_R1150_U390;
wire P1_R1150_U391 , P1_R1150_U392 , P1_R1150_U393 , P1_R1150_U394 , P1_R1150_U395 , P1_R1150_U396 , P1_R1150_U397 , P1_R1150_U398 , P1_R1150_U399 , P1_R1150_U400;
wire P1_R1150_U401 , P1_R1150_U402 , P1_R1150_U403 , P1_R1150_U404 , P1_R1150_U405 , P1_R1150_U406 , P1_R1150_U407 , P1_R1150_U408 , P1_R1150_U409 , P1_R1150_U410;
wire P1_R1150_U411 , P1_R1150_U412 , P1_R1150_U413 , P1_R1150_U414 , P1_R1150_U415 , P1_R1150_U416 , P1_R1150_U417 , P1_R1150_U418 , P1_R1150_U419 , P1_R1150_U420;
wire P1_R1150_U421 , P1_R1150_U422 , P1_R1150_U423 , P1_R1150_U424 , P1_R1150_U425 , P1_R1150_U426 , P1_R1150_U427 , P1_R1150_U428 , P1_R1150_U429 , P1_R1150_U430;
wire P1_R1150_U431 , P1_R1150_U432 , P1_R1150_U433 , P1_R1150_U434 , P1_R1150_U435 , P1_R1150_U436 , P1_R1150_U437 , P1_R1150_U438 , P1_R1150_U439 , P1_R1150_U440;
wire P1_R1150_U441 , P1_R1150_U442 , P1_R1150_U443 , P1_R1150_U444 , P1_R1150_U445 , P1_R1150_U446 , P1_R1150_U447 , P1_R1150_U448 , P1_R1150_U449 , P1_R1150_U450;
wire P1_R1150_U451 , P1_R1150_U452 , P1_R1150_U453 , P1_R1150_U454 , P1_R1150_U455 , P1_R1150_U456 , P1_R1150_U457 , P1_R1150_U458 , P1_R1150_U459 , P1_R1150_U460;
wire P1_R1150_U461 , P1_R1150_U462 , P1_R1150_U463 , P1_R1150_U464 , P1_R1150_U465 , P1_R1150_U466 , P1_R1150_U467 , P1_R1150_U468 , P1_R1150_U469 , P1_R1150_U470;
wire P1_R1150_U471 , P1_R1150_U472 , P1_R1150_U473 , P1_R1192_U6 , P1_R1192_U7 , P1_R1192_U8 , P1_R1192_U9 , P1_R1192_U10 , P1_R1192_U11 , P1_R1192_U12;
wire P1_R1192_U13 , P1_R1192_U14 , P1_R1192_U15 , P1_R1192_U16 , P1_R1192_U17 , P1_R1192_U18 , P1_R1192_U19 , P1_R1192_U20 , P1_R1192_U21 , P1_R1192_U22;
wire P1_R1192_U23 , P1_R1192_U24 , P1_R1192_U25 , P1_R1192_U26 , P1_R1192_U27 , P1_R1192_U28 , P1_R1192_U29 , P1_R1192_U30 , P1_R1192_U31 , P1_R1192_U32;
wire P1_R1192_U33 , P1_R1192_U34 , P1_R1192_U35 , P1_R1192_U36 , P1_R1192_U37 , P1_R1192_U38 , P1_R1192_U39 , P1_R1192_U40 , P1_R1192_U41 , P1_R1192_U42;
wire P1_R1192_U43 , P1_R1192_U44 , P1_R1192_U45 , P1_R1192_U46 , P1_R1192_U47 , P1_R1192_U48 , P1_R1192_U49 , P1_R1192_U50 , P1_R1192_U51 , P1_R1192_U52;
wire P1_R1192_U53 , P1_R1192_U54 , P1_R1192_U55 , P1_R1192_U56 , P1_R1192_U57 , P1_R1192_U58 , P1_R1192_U59 , P1_R1192_U60 , P1_R1192_U61 , P1_R1192_U62;
wire P1_R1192_U63 , P1_R1192_U64 , P1_R1192_U65 , P1_R1192_U66 , P1_R1192_U67 , P1_R1192_U68 , P1_R1192_U69 , P1_R1192_U70 , P1_R1192_U71 , P1_R1192_U72;
wire P1_R1192_U73 , P1_R1192_U74 , P1_R1192_U75 , P1_R1192_U76 , P1_R1192_U77 , P1_R1192_U78 , P1_R1192_U79 , P1_R1192_U80 , P1_R1192_U81 , P1_R1192_U82;
wire P1_R1192_U83 , P1_R1192_U84 , P1_R1192_U85 , P1_R1192_U86 , P1_R1192_U87 , P1_R1192_U88 , P1_R1192_U89 , P1_R1192_U90 , P1_R1192_U91 , P1_R1192_U92;
wire P1_R1192_U93 , P1_R1192_U94 , P1_R1192_U95 , P1_R1192_U96 , P1_R1192_U97 , P1_R1192_U98 , P1_R1192_U99 , P1_R1192_U100 , P1_R1192_U101 , P1_R1192_U102;
wire P1_R1192_U103 , P1_R1192_U104 , P1_R1192_U105 , P1_R1192_U106 , P1_R1192_U107 , P1_R1192_U108 , P1_R1192_U109 , P1_R1192_U110 , P1_R1192_U111 , P1_R1192_U112;
wire P1_R1192_U113 , P1_R1192_U114 , P1_R1192_U115 , P1_R1192_U116 , P1_R1192_U117 , P1_R1192_U118 , P1_R1192_U119 , P1_R1192_U120 , P1_R1192_U121 , P1_R1192_U122;
wire P1_R1192_U123 , P1_R1192_U124 , P1_R1192_U125 , P1_R1192_U126 , P1_R1192_U127 , P1_R1192_U128 , P1_R1192_U129 , P1_R1192_U130 , P1_R1192_U131 , P1_R1192_U132;
wire P1_R1192_U133 , P1_R1192_U134 , P1_R1192_U135 , P1_R1192_U136 , P1_R1192_U137 , P1_R1192_U138 , P1_R1192_U139 , P1_R1192_U140 , P1_R1192_U141 , P1_R1192_U142;
wire P1_R1192_U143 , P1_R1192_U144 , P1_R1192_U145 , P1_R1192_U146 , P1_R1192_U147 , P1_R1192_U148 , P1_R1192_U149 , P1_R1192_U150 , P1_R1192_U151 , P1_R1192_U152;
wire P1_R1192_U153 , P1_R1192_U154 , P1_R1192_U155 , P1_R1192_U156 , P1_R1192_U157 , P1_R1192_U158 , P1_R1192_U159 , P1_R1192_U160 , P1_R1192_U161 , P1_R1192_U162;
wire P1_R1192_U163 , P1_R1192_U164 , P1_R1192_U165 , P1_R1192_U166 , P1_R1192_U167 , P1_R1192_U168 , P1_R1192_U169 , P1_R1192_U170 , P1_R1192_U171 , P1_R1192_U172;
wire P1_R1192_U173 , P1_R1192_U174 , P1_R1192_U175 , P1_R1192_U176 , P1_R1192_U177 , P1_R1192_U178 , P1_R1192_U179 , P1_R1192_U180 , P1_R1192_U181 , P1_R1192_U182;
wire P1_R1192_U183 , P1_R1192_U184 , P1_R1192_U185 , P1_R1192_U186 , P1_R1192_U187 , P1_R1192_U188 , P1_R1192_U189 , P1_R1192_U190 , P1_R1192_U191 , P1_R1192_U192;
wire P1_R1192_U193 , P1_R1192_U194 , P1_R1192_U195 , P1_R1192_U196 , P1_R1192_U197 , P1_R1192_U198 , P1_R1192_U199 , P1_R1192_U200 , P1_R1192_U201 , P1_R1192_U202;
wire P1_R1192_U203 , P1_R1192_U204 , P1_R1192_U205 , P1_R1192_U206 , P1_R1192_U207 , P1_R1192_U208 , P1_R1192_U209 , P1_R1192_U210 , P1_R1192_U211 , P1_R1192_U212;
wire P1_R1192_U213 , P1_R1192_U214 , P1_R1192_U215 , P1_R1192_U216 , P1_R1192_U217 , P1_R1192_U218 , P1_R1192_U219 , P1_R1192_U220 , P1_R1192_U221 , P1_R1192_U222;
wire P1_R1192_U223 , P1_R1192_U224 , P1_R1192_U225 , P1_R1192_U226 , P1_R1192_U227 , P1_R1192_U228 , P1_R1192_U229 , P1_R1192_U230 , P1_R1192_U231 , P1_R1192_U232;
wire P1_R1192_U233 , P1_R1192_U234 , P1_R1192_U235 , P1_R1192_U236 , P1_R1192_U237 , P1_R1192_U238 , P1_R1192_U239 , P1_R1192_U240 , P1_R1192_U241 , P1_R1192_U242;
wire P1_R1192_U243 , P1_R1192_U244 , P1_R1192_U245 , P1_R1192_U246 , P1_R1192_U247 , P1_R1192_U248 , P1_R1192_U249 , P1_R1192_U250 , P1_R1192_U251 , P1_R1192_U252;
wire P1_R1192_U253 , P1_R1192_U254 , P1_R1192_U255 , P1_R1192_U256 , P1_R1192_U257 , P1_R1192_U258 , P1_R1192_U259 , P1_R1192_U260 , P1_R1192_U261 , P1_R1192_U262;
wire P1_R1192_U263 , P1_R1192_U264 , P1_R1192_U265 , P1_R1192_U266 , P1_R1192_U267 , P1_R1192_U268 , P1_R1192_U269 , P1_R1192_U270 , P1_R1192_U271 , P1_R1192_U272;
wire P1_R1192_U273 , P1_R1192_U274 , P1_R1192_U275 , P1_R1192_U276 , P1_R1192_U277 , P1_R1192_U278 , P1_R1192_U279 , P1_R1192_U280 , P1_R1192_U281 , P1_R1192_U282;
wire P1_R1192_U283 , P1_R1192_U284 , P1_R1192_U285 , P1_R1192_U286 , P1_R1192_U287 , P1_R1192_U288 , P1_R1192_U289 , P1_R1192_U290 , P1_R1192_U291 , P1_R1192_U292;
wire P1_R1192_U293 , P1_R1192_U294 , P1_R1192_U295 , P1_R1192_U296 , P1_R1192_U297 , P1_R1192_U298 , P1_R1192_U299 , P1_R1192_U300 , P1_R1192_U301 , P1_R1192_U302;
wire P1_R1192_U303 , P1_R1192_U304 , P1_R1192_U305 , P1_R1192_U306 , P1_R1192_U307 , P1_R1192_U308 , P1_R1192_U309 , P1_R1192_U310 , P1_R1192_U311 , P1_R1192_U312;
wire P1_R1192_U313 , P1_R1192_U314 , P1_R1192_U315 , P1_R1192_U316 , P1_R1192_U317 , P1_R1192_U318 , P1_R1192_U319 , P1_R1192_U320 , P1_R1192_U321 , P1_R1192_U322;
wire P1_R1192_U323 , P1_R1192_U324 , P1_R1192_U325 , P1_R1192_U326 , P1_R1192_U327 , P1_R1192_U328 , P1_R1192_U329 , P1_R1192_U330 , P1_R1192_U331 , P1_R1192_U332;
wire P1_R1192_U333 , P1_R1192_U334 , P1_R1192_U335 , P1_R1192_U336 , P1_R1192_U337 , P1_R1192_U338 , P1_R1192_U339 , P1_R1192_U340 , P1_R1192_U341 , P1_R1192_U342;
wire P1_R1192_U343 , P1_R1192_U344 , P1_R1192_U345 , P1_R1192_U346 , P1_R1192_U347 , P1_R1192_U348 , P1_R1192_U349 , P1_R1192_U350 , P1_R1192_U351 , P1_R1192_U352;
wire P1_R1192_U353 , P1_R1192_U354 , P1_R1192_U355 , P1_R1192_U356 , P1_R1192_U357 , P1_R1192_U358 , P1_R1192_U359 , P1_R1192_U360 , P1_R1192_U361 , P1_R1192_U362;
wire P1_R1192_U363 , P1_R1192_U364 , P1_R1192_U365 , P1_R1192_U366 , P1_R1192_U367 , P1_R1192_U368 , P1_R1192_U369 , P1_R1192_U370 , P1_R1192_U371 , P1_R1192_U372;
wire P1_R1192_U373 , P1_R1192_U374 , P1_R1192_U375 , P1_R1192_U376 , P1_R1192_U377 , P1_R1192_U378 , P1_R1192_U379 , P1_R1192_U380 , P1_R1192_U381 , P1_R1192_U382;
wire P1_R1192_U383 , P1_R1192_U384 , P1_R1192_U385 , P1_R1192_U386 , P1_R1192_U387 , P1_R1192_U388 , P1_R1192_U389 , P1_R1192_U390 , P1_R1192_U391 , P1_R1192_U392;
wire P1_R1192_U393 , P1_R1192_U394 , P1_R1192_U395 , P1_R1192_U396 , P1_R1192_U397 , P1_R1192_U398 , P1_R1192_U399 , P1_R1192_U400 , P1_R1192_U401 , P1_R1192_U402;
wire P1_R1192_U403 , P1_R1192_U404 , P1_R1192_U405 , P1_R1192_U406 , P1_R1192_U407 , P1_R1192_U408 , P1_R1192_U409 , P1_R1192_U410 , P1_R1192_U411 , P1_R1192_U412;
wire P1_R1192_U413 , P1_R1192_U414 , P1_R1192_U415 , P1_R1192_U416 , P1_R1192_U417 , P1_R1192_U418 , P1_R1192_U419 , P1_R1192_U420 , P1_R1192_U421 , P1_R1192_U422;
wire P1_R1192_U423 , P1_R1192_U424 , P1_R1192_U425 , P1_R1192_U426 , P1_R1192_U427 , P1_R1192_U428 , P1_R1192_U429 , P1_R1192_U430 , P1_R1192_U431 , P1_R1192_U432;
wire P1_R1192_U433 , P1_R1192_U434 , P1_R1192_U435 , P1_R1192_U436 , P1_R1192_U437 , P1_R1192_U438 , P1_R1192_U439 , P1_R1192_U440 , P1_R1192_U441 , P1_R1192_U442;
wire P1_R1192_U443 , P1_R1192_U444 , P1_R1192_U445 , P1_R1192_U446 , P1_R1192_U447 , P1_R1192_U448 , P1_R1192_U449 , P1_R1192_U450 , P1_R1192_U451 , P1_R1192_U452;
wire P1_R1192_U453 , P1_R1192_U454 , P1_R1192_U455 , P1_R1192_U456 , P1_R1192_U457 , P1_R1192_U458 , P1_R1192_U459 , P1_R1192_U460 , P1_R1192_U461 , P1_R1192_U462;
wire P1_R1192_U463 , P1_R1192_U464 , P1_R1192_U465 , P1_R1192_U466 , P1_R1192_U467 , P1_R1192_U468 , P1_R1192_U469 , P1_R1192_U470 , P1_R1192_U471 , P1_R1192_U472;
wire P1_R1192_U473 , P1_LT_197_U6 , P1_LT_197_U7 , P1_LT_197_U8 , P1_LT_197_U9 , P1_LT_197_U10 , P1_LT_197_U11 , P1_LT_197_U12 , P1_LT_197_U13 , P1_LT_197_U14;
wire P1_LT_197_U15 , P1_LT_197_U16 , P1_LT_197_U17 , P1_LT_197_U18 , P1_LT_197_U19 , P1_LT_197_U20 , P1_LT_197_U21 , P1_LT_197_U22 , P1_LT_197_U23 , P1_LT_197_U24;
wire P1_LT_197_U25 , P1_LT_197_U26 , P1_LT_197_U27 , P1_LT_197_U28 , P1_LT_197_U29 , P1_LT_197_U30 , P1_LT_197_U31 , P1_LT_197_U32 , P1_LT_197_U33 , P1_LT_197_U34;
wire P1_LT_197_U35 , P1_LT_197_U36 , P1_LT_197_U37 , P1_LT_197_U38 , P1_LT_197_U39 , P1_LT_197_U40 , P1_LT_197_U41 , P1_LT_197_U42 , P1_LT_197_U43 , P1_LT_197_U44;
wire P1_LT_197_U45 , P1_LT_197_U46 , P1_LT_197_U47 , P1_LT_197_U48 , P1_LT_197_U49 , P1_LT_197_U50 , P1_LT_197_U51 , P1_LT_197_U52 , P1_LT_197_U53 , P1_LT_197_U54;
wire P1_LT_197_U55 , P1_LT_197_U56 , P1_LT_197_U57 , P1_LT_197_U58 , P1_LT_197_U59 , P1_LT_197_U60 , P1_LT_197_U61 , P1_LT_197_U62 , P1_LT_197_U63 , P1_LT_197_U64;
wire P1_LT_197_U65 , P1_LT_197_U66 , P1_LT_197_U67 , P1_LT_197_U68 , P1_LT_197_U69 , P1_LT_197_U70 , P1_LT_197_U71 , P1_LT_197_U72 , P1_LT_197_U73 , P1_LT_197_U74;
wire P1_LT_197_U75 , P1_LT_197_U76 , P1_LT_197_U77 , P1_LT_197_U78 , P1_LT_197_U79 , P1_LT_197_U80 , P1_LT_197_U81 , P1_LT_197_U82 , P1_LT_197_U83 , P1_LT_197_U84;
wire P1_LT_197_U85 , P1_LT_197_U86 , P1_LT_197_U87 , P1_LT_197_U88 , P1_LT_197_U89 , P1_LT_197_U90 , P1_LT_197_U91 , P1_LT_197_U92 , P1_LT_197_U93 , P1_LT_197_U94;
wire P1_LT_197_U95 , P1_LT_197_U96 , P1_LT_197_U97 , P1_LT_197_U98 , P1_LT_197_U99 , P1_LT_197_U100 , P1_LT_197_U101 , P1_LT_197_U102 , P1_LT_197_U103 , P1_LT_197_U104;
wire P1_LT_197_U105 , P1_LT_197_U106 , P1_LT_197_U107 , P1_LT_197_U108 , P1_LT_197_U109 , P1_LT_197_U110 , P1_LT_197_U111 , P1_LT_197_U112 , P1_LT_197_U113 , P1_LT_197_U114;
wire P1_LT_197_U115 , P1_LT_197_U116 , P1_LT_197_U117 , P1_LT_197_U118 , P1_LT_197_U119 , P1_LT_197_U120 , P1_LT_197_U121 , P1_LT_197_U122 , P1_LT_197_U123 , P1_LT_197_U124;
wire P1_LT_197_U125 , P1_LT_197_U126 , P1_LT_197_U127 , P1_LT_197_U128 , P1_LT_197_U129 , P1_LT_197_U130 , P1_LT_197_U131 , P1_LT_197_U132 , P1_LT_197_U133 , P1_LT_197_U134;
wire P1_LT_197_U135 , P1_LT_197_U136 , P1_LT_197_U137 , P1_LT_197_U138 , P1_LT_197_U139 , P1_LT_197_U140 , P1_LT_197_U141 , P1_LT_197_U142 , P1_LT_197_U143 , P1_LT_197_U144;
wire P1_LT_197_U145 , P1_LT_197_U146 , P1_LT_197_U147 , P1_LT_197_U148 , P1_LT_197_U149 , P1_LT_197_U150 , P1_LT_197_U151 , P1_LT_197_U152 , P1_LT_197_U153 , P1_LT_197_U154;
wire P1_LT_197_U155 , P1_LT_197_U156 , P1_LT_197_U157 , P1_LT_197_U158 , P1_LT_197_U159 , P1_LT_197_U160 , P1_LT_197_U161 , P1_LT_197_U162 , P1_LT_197_U163 , P1_LT_197_U164;
wire P1_LT_197_U165 , P1_LT_197_U166 , P1_LT_197_U167 , P1_LT_197_U168 , P1_LT_197_U169 , P1_LT_197_U170 , P1_LT_197_U171 , P1_LT_197_U172 , P1_LT_197_U173 , P1_LT_197_U174;
wire P1_LT_197_U175 , P1_LT_197_U176 , P1_LT_197_U177 , P1_LT_197_U178 , P1_LT_197_U179 , P1_LT_197_U180 , P1_LT_197_U181 , P1_LT_197_U182 , P1_LT_197_U183 , P1_LT_197_U184;
wire P1_LT_197_U185 , P1_LT_197_U186 , P1_LT_197_U187 , P1_LT_197_U188 , P1_LT_197_U189 , P1_LT_197_U190 , P1_LT_197_U191 , P1_LT_197_U192 , P1_LT_197_U193 , P1_LT_197_U194;
wire P1_LT_197_U195 , P1_LT_197_U196 , P1_LT_197_U197 , P1_LT_197_U198 , P1_LT_197_U199 , P1_LT_197_U200 , P1_R1360_U6 , P1_R1360_U7 , P1_R1360_U8 , P1_R1360_U9;
wire P1_R1360_U10 , P1_R1360_U11 , P1_R1360_U12 , P1_R1360_U13 , P1_R1360_U14 , P1_R1360_U15 , P1_R1360_U16 , P1_R1360_U17 , P1_R1360_U18 , P1_R1360_U19;
wire P1_R1360_U20 , P1_R1360_U21 , P1_R1360_U22 , P1_R1360_U23 , P1_R1360_U24 , P1_R1360_U25 , P1_R1360_U26 , P1_R1360_U27 , P1_R1360_U28 , P1_R1360_U29;
wire P1_R1360_U30 , P1_R1360_U31 , P1_R1360_U32 , P1_R1360_U33 , P1_R1360_U34 , P1_R1360_U35 , P1_R1360_U36 , P1_R1360_U37 , P1_R1360_U38 , P1_R1360_U39;
wire P1_R1360_U40 , P1_R1360_U41 , P1_R1360_U42 , P1_R1360_U43 , P1_R1360_U44 , P1_R1360_U45 , P1_R1360_U46 , P1_R1360_U47 , P1_R1360_U48 , P1_R1360_U49;
wire P1_R1360_U50 , P1_R1360_U51 , P1_R1360_U52 , P1_R1360_U53 , P1_R1360_U54 , P1_R1360_U55 , P1_R1360_U56 , P1_R1360_U57 , P1_R1360_U58 , P1_R1360_U59;
wire P1_R1360_U60 , P1_R1360_U61 , P1_R1360_U62 , P1_R1360_U63 , P1_R1360_U64 , P1_R1360_U65 , P1_R1360_U66 , P1_R1360_U67 , P1_R1360_U68 , P1_R1360_U69;
wire P1_R1360_U70 , P1_R1360_U71 , P1_R1360_U72 , P1_R1360_U73 , P1_R1360_U74 , P1_R1360_U75 , P1_R1360_U76 , P1_R1360_U77 , P1_R1360_U78 , P1_R1360_U79;
wire P1_R1360_U80 , P1_R1360_U81 , P1_R1360_U82 , P1_R1360_U83 , P1_R1360_U84 , P1_R1360_U85 , P1_R1360_U86 , P1_R1360_U87 , P1_R1360_U88 , P1_R1360_U89;
wire P1_R1360_U90 , P1_R1360_U91 , P1_R1360_U92 , P1_R1360_U93 , P1_R1360_U94 , P1_R1360_U95 , P1_R1360_U96 , P1_R1360_U97 , P1_R1360_U98 , P1_R1360_U99;
wire P1_R1360_U100 , P1_R1360_U101 , P1_R1360_U102 , P1_R1360_U103 , P1_R1360_U104 , P1_R1360_U105 , P1_R1360_U106 , P1_R1360_U107 , P1_R1360_U108 , P1_R1360_U109;
wire P1_R1360_U110 , P1_R1360_U111 , P1_R1360_U112 , P1_R1360_U113 , P1_R1360_U114 , P1_R1360_U115 , P1_R1360_U116 , P1_R1360_U117 , P1_R1360_U118 , P1_R1360_U119;
wire P1_R1360_U120 , P1_R1360_U121 , P1_R1360_U122 , P1_R1360_U123 , P1_R1360_U124 , P1_R1360_U125 , P1_R1360_U126 , P1_R1360_U127 , P1_R1360_U128 , P1_R1360_U129;
wire P1_R1360_U130 , P1_R1360_U131 , P1_R1360_U132 , P1_R1360_U133 , P1_R1360_U134 , P1_R1360_U135 , P1_R1360_U136 , P1_R1360_U137 , P1_R1360_U138 , P1_R1360_U139;
wire P1_R1360_U140 , P1_R1360_U141 , P1_R1360_U142 , P1_R1360_U143 , P1_R1360_U144 , P1_R1360_U145 , P1_R1360_U146 , P1_R1360_U147 , P1_R1360_U148 , P1_R1360_U149;
wire P1_R1360_U150 , P1_R1360_U151 , P1_R1360_U152 , P1_R1360_U153 , P1_R1360_U154 , P1_R1360_U155 , P1_R1360_U156 , P1_R1360_U157 , P1_R1360_U158 , P1_R1360_U159;
wire P1_R1360_U160 , P1_R1360_U161 , P1_R1360_U162 , P1_R1360_U163 , P1_R1360_U164 , P1_R1360_U165 , P1_R1360_U166 , P1_R1360_U167 , P1_R1360_U168 , P1_R1360_U169;
wire P1_R1360_U170 , P1_R1360_U171 , P1_R1360_U172 , P1_R1360_U173 , P1_R1360_U174 , P1_R1360_U175 , P1_R1360_U176 , P1_R1360_U177 , P1_R1360_U178 , P1_R1360_U179;
wire P1_R1360_U180 , P1_R1360_U181 , P1_R1360_U182 , P1_R1360_U183 , P1_R1360_U184 , P1_R1360_U185 , P1_R1360_U186 , P1_R1360_U187 , P1_R1360_U188 , P1_R1360_U189;
wire P1_R1360_U190 , P1_R1360_U191 , P1_R1360_U192 , P1_R1360_U193 , P1_R1360_U194 , P1_R1360_U195 , P1_R1360_U196 , P1_R1360_U197 , P1_R1360_U198 , P1_R1360_U199;
wire P1_R1360_U200 , P1_R1360_U201 , P1_R1360_U202 , P1_R1360_U203 , P1_R1360_U204 , P1_R1360_U205 , P1_R1171_U4 , P1_R1171_U5 , P1_R1171_U6 , P1_R1171_U7;
wire P1_R1171_U8 , P1_R1171_U9 , P1_R1171_U10 , P1_R1171_U11 , P1_R1171_U12 , P1_R1171_U13 , P1_R1171_U14 , P1_R1171_U15 , P1_R1171_U16 , P1_R1171_U17;
wire P1_R1171_U18 , P1_R1171_U19 , P1_R1171_U20 , P1_R1171_U21 , P1_R1171_U22 , P1_R1171_U23 , P1_R1171_U24 , P1_R1171_U25 , P1_R1171_U26 , P1_R1171_U27;
wire P1_R1171_U28 , P1_R1171_U29 , P1_R1171_U30 , P1_R1171_U31 , P1_R1171_U32 , P1_R1171_U33 , P1_R1171_U34 , P1_R1171_U35 , P1_R1171_U36 , P1_R1171_U37;
wire P1_R1171_U38 , P1_R1171_U39 , P1_R1171_U40 , P1_R1171_U41 , P1_R1171_U42 , P1_R1171_U43 , P1_R1171_U44 , P1_R1171_U45 , P1_R1171_U46 , P1_R1171_U47;
wire P1_R1171_U48 , P1_R1171_U49 , P1_R1171_U50 , P1_R1171_U51 , P1_R1171_U52 , P1_R1171_U53 , P1_R1171_U54 , P1_R1171_U55 , P1_R1171_U56 , P1_R1171_U57;
wire P1_R1171_U58 , P1_R1171_U59 , P1_R1171_U60 , P1_R1171_U61 , P1_R1171_U62 , P1_R1171_U63 , P1_R1171_U64 , P1_R1171_U65 , P1_R1171_U66 , P1_R1171_U67;
wire P1_R1171_U68 , P1_R1171_U69 , P1_R1171_U70 , P1_R1171_U71 , P1_R1171_U72 , P1_R1171_U73 , P1_R1171_U74 , P1_R1171_U75 , P1_R1171_U76 , P1_R1171_U77;
wire P1_R1171_U78 , P1_R1171_U79 , P1_R1171_U80 , P1_R1171_U81 , P1_R1171_U82 , P1_R1171_U83 , P1_R1171_U84 , P1_R1171_U85 , P1_R1171_U86 , P1_R1171_U87;
wire P1_R1171_U88 , P1_R1171_U89 , P1_R1171_U90 , P1_R1171_U91 , P1_R1171_U92 , P1_R1171_U93 , P1_R1171_U94 , P1_R1171_U95 , P1_R1171_U96 , P1_R1171_U97;
wire P1_R1171_U98 , P1_R1171_U99 , P1_R1171_U100 , P1_R1171_U101 , P1_R1171_U102 , P1_R1171_U103 , P1_R1171_U104 , P1_R1171_U105 , P1_R1171_U106 , P1_R1171_U107;
wire P1_R1171_U108 , P1_R1171_U109 , P1_R1171_U110 , P1_R1171_U111 , P1_R1171_U112 , P1_R1171_U113 , P1_R1171_U114 , P1_R1171_U115 , P1_R1171_U116 , P1_R1171_U117;
wire P1_R1171_U118 , P1_R1171_U119 , P1_R1171_U120 , P1_R1171_U121 , P1_R1171_U122 , P1_R1171_U123 , P1_R1171_U124 , P1_R1171_U125 , P1_R1171_U126 , P1_R1171_U127;
wire P1_R1171_U128 , P1_R1171_U129 , P1_R1171_U130 , P1_R1171_U131 , P1_R1171_U132 , P1_R1171_U133 , P1_R1171_U134 , P1_R1171_U135 , P1_R1171_U136 , P1_R1171_U137;
wire P1_R1171_U138 , P1_R1171_U139 , P1_R1171_U140 , P1_R1171_U141 , P1_R1171_U142 , P1_R1171_U143 , P1_R1171_U144 , P1_R1171_U145 , P1_R1171_U146 , P1_R1171_U147;
wire P1_R1171_U148 , P1_R1171_U149 , P1_R1171_U150 , P1_R1171_U151 , P1_R1171_U152 , P1_R1171_U153 , P1_R1171_U154 , P1_R1171_U155 , P1_R1171_U156 , P1_R1171_U157;
wire P1_R1171_U158 , P1_R1171_U159 , P1_R1171_U160 , P1_R1171_U161 , P1_R1171_U162 , P1_R1171_U163 , P1_R1171_U164 , P1_R1171_U165 , P1_R1171_U166 , P1_R1171_U167;
wire P1_R1171_U168 , P1_R1171_U169 , P1_R1171_U170 , P1_R1171_U171 , P1_R1171_U172 , P1_R1171_U173 , P1_R1171_U174 , P1_R1171_U175 , P1_R1171_U176 , P1_R1171_U177;
wire P1_R1171_U178 , P1_R1171_U179 , P1_R1171_U180 , P1_R1171_U181 , P1_R1171_U182 , P1_R1171_U183 , P1_R1171_U184 , P1_R1171_U185 , P1_R1171_U186 , P1_R1171_U187;
wire P1_R1171_U188 , P1_R1171_U189 , P1_R1171_U190 , P1_R1171_U191 , P1_R1171_U192 , P1_R1171_U193 , P1_R1171_U194 , P1_R1171_U195 , P1_R1171_U196 , P1_R1171_U197;
wire P1_R1171_U198 , P1_R1171_U199 , P1_R1171_U200 , P1_R1171_U201 , P1_R1171_U202 , P1_R1171_U203 , P1_R1171_U204 , P1_R1171_U205 , P1_R1171_U206 , P1_R1171_U207;
wire P1_R1171_U208 , P1_R1171_U209 , P1_R1171_U210 , P1_R1171_U211 , P1_R1171_U212 , P1_R1171_U213 , P1_R1171_U214 , P1_R1171_U215 , P1_R1171_U216 , P1_R1171_U217;
wire P1_R1171_U218 , P1_R1171_U219 , P1_R1171_U220 , P1_R1171_U221 , P1_R1171_U222 , P1_R1171_U223 , P1_R1171_U224 , P1_R1171_U225 , P1_R1171_U226 , P1_R1171_U227;
wire P1_R1171_U228 , P1_R1171_U229 , P1_R1171_U230 , P1_R1171_U231 , P1_R1171_U232 , P1_R1171_U233 , P1_R1171_U234 , P1_R1171_U235 , P1_R1171_U236 , P1_R1171_U237;
wire P1_R1171_U238 , P1_R1171_U239 , P1_R1171_U240 , P1_R1171_U241 , P1_R1171_U242 , P1_R1171_U243 , P1_R1171_U244 , P1_R1171_U245 , P1_R1171_U246 , P1_R1171_U247;
wire P1_R1171_U248 , P1_R1171_U249 , P1_R1171_U250 , P1_R1171_U251 , P1_R1171_U252 , P1_R1171_U253 , P1_R1171_U254 , P1_R1171_U255 , P1_R1171_U256 , P1_R1171_U257;
wire P1_R1171_U258 , P1_R1171_U259 , P1_R1171_U260 , P1_R1171_U261 , P1_R1171_U262 , P1_R1171_U263 , P1_R1171_U264 , P1_R1171_U265 , P1_R1171_U266 , P1_R1171_U267;
wire P1_R1171_U268 , P1_R1171_U269 , P1_R1171_U270 , P1_R1171_U271 , P1_R1171_U272 , P1_R1171_U273 , P1_R1171_U274 , P1_R1171_U275 , P1_R1171_U276 , P1_R1171_U277;
wire P1_R1171_U278 , P1_R1171_U279 , P1_R1171_U280 , P1_R1171_U281 , P1_R1171_U282 , P1_R1171_U283 , P1_R1171_U284 , P1_R1171_U285 , P1_R1171_U286 , P1_R1171_U287;
wire P1_R1171_U288 , P1_R1171_U289 , P1_R1171_U290 , P1_R1171_U291 , P1_R1171_U292 , P1_R1171_U293 , P1_R1171_U294 , P1_R1171_U295 , P1_R1171_U296 , P1_R1171_U297;
wire P1_R1171_U298 , P1_R1171_U299 , P1_R1171_U300 , P1_R1171_U301 , P1_R1171_U302 , P1_R1171_U303 , P1_R1171_U304 , P1_R1171_U305 , P1_R1171_U306 , P1_R1171_U307;
wire P1_R1171_U308 , P1_R1171_U309 , P1_R1171_U310 , P1_R1171_U311 , P1_R1171_U312 , P1_R1171_U313 , P1_R1171_U314 , P1_R1171_U315 , P1_R1171_U316 , P1_R1171_U317;
wire P1_R1171_U318 , P1_R1171_U319 , P1_R1171_U320 , P1_R1171_U321 , P1_R1171_U322 , P1_R1171_U323 , P1_R1171_U324 , P1_R1171_U325 , P1_R1171_U326 , P1_R1171_U327;
wire P1_R1171_U328 , P1_R1171_U329 , P1_R1171_U330 , P1_R1171_U331 , P1_R1171_U332 , P1_R1171_U333 , P1_R1171_U334 , P1_R1171_U335 , P1_R1171_U336 , P1_R1171_U337;
wire P1_R1171_U338 , P1_R1171_U339 , P1_R1171_U340 , P1_R1171_U341 , P1_R1171_U342 , P1_R1171_U343 , P1_R1171_U344 , P1_R1171_U345 , P1_R1171_U346 , P1_R1171_U347;
wire P1_R1171_U348 , P1_R1171_U349 , P1_R1171_U350 , P1_R1171_U351 , P1_R1171_U352 , P1_R1171_U353 , P1_R1171_U354 , P1_R1171_U355 , P1_R1171_U356 , P1_R1171_U357;
wire P1_R1171_U358 , P1_R1171_U359 , P1_R1171_U360 , P1_R1171_U361 , P1_R1171_U362 , P1_R1171_U363 , P1_R1171_U364 , P1_R1171_U365 , P1_R1171_U366 , P1_R1171_U367;
wire P1_R1171_U368 , P1_R1171_U369 , P1_R1171_U370 , P1_R1171_U371 , P1_R1171_U372 , P1_R1171_U373 , P1_R1171_U374 , P1_R1171_U375 , P1_R1171_U376 , P1_R1171_U377;
wire P1_R1171_U378 , P1_R1171_U379 , P1_R1171_U380 , P1_R1171_U381 , P1_R1171_U382 , P1_R1171_U383 , P1_R1171_U384 , P1_R1171_U385 , P1_R1171_U386 , P1_R1171_U387;
wire P1_R1171_U388 , P1_R1171_U389 , P1_R1171_U390 , P1_R1171_U391 , P1_R1171_U392 , P1_R1171_U393 , P1_R1171_U394 , P1_R1171_U395 , P1_R1171_U396 , P1_R1171_U397;
wire P1_R1171_U398 , P1_R1171_U399 , P1_R1171_U400 , P1_R1171_U401 , P1_R1171_U402 , P1_R1171_U403 , P1_R1171_U404 , P1_R1171_U405 , P1_R1171_U406 , P1_R1171_U407;
wire P1_R1171_U408 , P1_R1171_U409 , P1_R1171_U410 , P1_R1171_U411 , P1_R1171_U412 , P1_R1171_U413 , P1_R1171_U414 , P1_R1171_U415 , P1_R1171_U416 , P1_R1171_U417;
wire P1_R1171_U418 , P1_R1171_U419 , P1_R1171_U420 , P1_R1171_U421 , P1_R1171_U422 , P1_R1171_U423 , P1_R1171_U424 , P1_R1171_U425 , P1_R1171_U426 , P1_R1171_U427;
wire P1_R1171_U428 , P1_R1171_U429 , P1_R1171_U430 , P1_R1171_U431 , P1_R1171_U432 , P1_R1171_U433 , P1_R1171_U434 , P1_R1171_U435 , P1_R1171_U436 , P1_R1171_U437;
wire P1_R1171_U438 , P1_R1171_U439 , P1_R1171_U440 , P1_R1171_U441 , P1_R1171_U442 , P1_R1171_U443 , P1_R1171_U444 , P1_R1171_U445 , P1_R1171_U446 , P1_R1171_U447;
wire P1_R1171_U448 , P1_R1171_U449 , P1_R1171_U450 , P1_R1171_U451 , P1_R1171_U452 , P1_R1171_U453 , P1_R1171_U454 , P1_R1171_U455 , P1_R1171_U456 , P1_R1171_U457;
wire P1_R1171_U458 , P1_R1171_U459 , P1_R1171_U460 , P1_R1171_U461 , P1_R1171_U462 , P1_R1171_U463 , P1_R1171_U464 , P1_R1171_U465 , P1_R1171_U466 , P1_R1171_U467;
wire P1_R1171_U468 , P1_R1171_U469 , P1_R1171_U470 , P1_R1171_U471 , P1_R1171_U472 , P1_R1171_U473 , P1_R1171_U474 , P1_R1171_U475 , P1_R1171_U476 , P1_R1171_U477;
wire P1_R1171_U478 , P1_R1171_U479 , P1_R1171_U480 , P1_R1171_U481 , P1_R1171_U482 , P1_R1171_U483 , P1_R1171_U484 , P1_R1171_U485 , P1_R1171_U486 , P1_R1171_U487;
wire P1_R1171_U488 , P1_R1171_U489 , P1_R1171_U490 , P1_R1171_U491 , P1_R1171_U492 , P1_R1171_U493 , P1_R1171_U494 , P1_R1171_U495 , P1_R1171_U496 , P1_R1171_U497;
wire P1_R1171_U498 , P1_R1171_U499 , P1_R1171_U500 , P1_R1171_U501 , P1_R1171_U502 , P1_R1171_U503 , P1_R1138_U4 , P1_R1138_U5 , P1_R1138_U6 , P1_R1138_U7;
wire P1_R1138_U8 , P1_R1138_U9 , P1_R1138_U10 , P1_R1138_U11 , P1_R1138_U12 , P1_R1138_U13 , P1_R1138_U14 , P1_R1138_U15 , P1_R1138_U16 , P1_R1138_U17;
wire P1_R1138_U18 , P1_R1138_U19 , P1_R1138_U20 , P1_R1138_U21 , P1_R1138_U22 , P1_R1138_U23 , P1_R1138_U24 , P1_R1138_U25 , P1_R1138_U26 , P1_R1138_U27;
wire P1_R1138_U28 , P1_R1138_U29 , P1_R1138_U30 , P1_R1138_U31 , P1_R1138_U32 , P1_R1138_U33 , P1_R1138_U34 , P1_R1138_U35 , P1_R1138_U36 , P1_R1138_U37;
wire P1_R1138_U38 , P1_R1138_U39 , P1_R1138_U40 , P1_R1138_U41 , P1_R1138_U42 , P1_R1138_U43 , P1_R1138_U44 , P1_R1138_U45 , P1_R1138_U46 , P1_R1138_U47;
wire P1_R1138_U48 , P1_R1138_U49 , P1_R1138_U50 , P1_R1138_U51 , P1_R1138_U52 , P1_R1138_U53 , P1_R1138_U54 , P1_R1138_U55 , P1_R1138_U56 , P1_R1138_U57;
wire P1_R1138_U58 , P1_R1138_U59 , P1_R1138_U60 , P1_R1138_U61 , P1_R1138_U62 , P1_R1138_U63 , P1_R1138_U64 , P1_R1138_U65 , P1_R1138_U66 , P1_R1138_U67;
wire P1_R1138_U68 , P1_R1138_U69 , P1_R1138_U70 , P1_R1138_U71 , P1_R1138_U72 , P1_R1138_U73 , P1_R1138_U74 , P1_R1138_U75 , P1_R1138_U76 , P1_R1138_U77;
wire P1_R1138_U78 , P1_R1138_U79 , P1_R1138_U80 , P1_R1138_U81 , P1_R1138_U82 , P1_R1138_U83 , P1_R1138_U84 , P1_R1138_U85 , P1_R1138_U86 , P1_R1138_U87;
wire P1_R1138_U88 , P1_R1138_U89 , P1_R1138_U90 , P1_R1138_U91 , P1_R1138_U92 , P1_R1138_U93 , P1_R1138_U94 , P1_R1138_U95 , P1_R1138_U96 , P1_R1138_U97;
wire P1_R1138_U98 , P1_R1138_U99 , P1_R1138_U100 , P1_R1138_U101 , P1_R1138_U102 , P1_R1138_U103 , P1_R1138_U104 , P1_R1138_U105 , P1_R1138_U106 , P1_R1138_U107;
wire P1_R1138_U108 , P1_R1138_U109 , P1_R1138_U110 , P1_R1138_U111 , P1_R1138_U112 , P1_R1138_U113 , P1_R1138_U114 , P1_R1138_U115 , P1_R1138_U116 , P1_R1138_U117;
wire P1_R1138_U118 , P1_R1138_U119 , P1_R1138_U120 , P1_R1138_U121 , P1_R1138_U122 , P1_R1138_U123 , P1_R1138_U124 , P1_R1138_U125 , P1_R1138_U126 , P1_R1138_U127;
wire P1_R1138_U128 , P1_R1138_U129 , P1_R1138_U130 , P1_R1138_U131 , P1_R1138_U132 , P1_R1138_U133 , P1_R1138_U134 , P1_R1138_U135 , P1_R1138_U136 , P1_R1138_U137;
wire P1_R1138_U138 , P1_R1138_U139 , P1_R1138_U140 , P1_R1138_U141 , P1_R1138_U142 , P1_R1138_U143 , P1_R1138_U144 , P1_R1138_U145 , P1_R1138_U146 , P1_R1138_U147;
wire P1_R1138_U148 , P1_R1138_U149 , P1_R1138_U150 , P1_R1138_U151 , P1_R1138_U152 , P1_R1138_U153 , P1_R1138_U154 , P1_R1138_U155 , P1_R1138_U156 , P1_R1138_U157;
wire P1_R1138_U158 , P1_R1138_U159 , P1_R1138_U160 , P1_R1138_U161 , P1_R1138_U162 , P1_R1138_U163 , P1_R1138_U164 , P1_R1138_U165 , P1_R1138_U166 , P1_R1138_U167;
wire P1_R1138_U168 , P1_R1138_U169 , P1_R1138_U170 , P1_R1138_U171 , P1_R1138_U172 , P1_R1138_U173 , P1_R1138_U174 , P1_R1138_U175 , P1_R1138_U176 , P1_R1138_U177;
wire P1_R1138_U178 , P1_R1138_U179 , P1_R1138_U180 , P1_R1138_U181 , P1_R1138_U182 , P1_R1138_U183 , P1_R1138_U184 , P1_R1138_U185 , P1_R1138_U186 , P1_R1138_U187;
wire P1_R1138_U188 , P1_R1138_U189 , P1_R1138_U190 , P1_R1138_U191 , P1_R1138_U192 , P1_R1138_U193 , P1_R1138_U194 , P1_R1138_U195 , P1_R1138_U196 , P1_R1138_U197;
wire P1_R1138_U198 , P1_R1138_U199 , P1_R1138_U200 , P1_R1138_U201 , P1_R1138_U202 , P1_R1138_U203 , P1_R1138_U204 , P1_R1138_U205 , P1_R1138_U206 , P1_R1138_U207;
wire P1_R1138_U208 , P1_R1138_U209 , P1_R1138_U210 , P1_R1138_U211 , P1_R1138_U212 , P1_R1138_U213 , P1_R1138_U214 , P1_R1138_U215 , P1_R1138_U216 , P1_R1138_U217;
wire P1_R1138_U218 , P1_R1138_U219 , P1_R1138_U220 , P1_R1138_U221 , P1_R1138_U222 , P1_R1138_U223 , P1_R1138_U224 , P1_R1138_U225 , P1_R1138_U226 , P1_R1138_U227;
wire P1_R1138_U228 , P1_R1138_U229 , P1_R1138_U230 , P1_R1138_U231 , P1_R1138_U232 , P1_R1138_U233 , P1_R1138_U234 , P1_R1138_U235 , P1_R1138_U236 , P1_R1138_U237;
wire P1_R1138_U238 , P1_R1138_U239 , P1_R1138_U240 , P1_R1138_U241 , P1_R1138_U242 , P1_R1138_U243 , P1_R1138_U244 , P1_R1138_U245 , P1_R1138_U246 , P1_R1138_U247;
wire P1_R1138_U248 , P1_R1138_U249 , P1_R1138_U250 , P1_R1138_U251 , P1_R1138_U252 , P1_R1138_U253 , P1_R1138_U254 , P1_R1138_U255 , P1_R1138_U256 , P1_R1138_U257;
wire P1_R1138_U258 , P1_R1138_U259 , P1_R1138_U260 , P1_R1138_U261 , P1_R1138_U262 , P1_R1138_U263 , P1_R1138_U264 , P1_R1138_U265 , P1_R1138_U266 , P1_R1138_U267;
wire P1_R1138_U268 , P1_R1138_U269 , P1_R1138_U270 , P1_R1138_U271 , P1_R1138_U272 , P1_R1138_U273 , P1_R1138_U274 , P1_R1138_U275 , P1_R1138_U276 , P1_R1138_U277;
wire P1_R1138_U278 , P1_R1138_U279 , P1_R1138_U280 , P1_R1138_U281 , P1_R1138_U282 , P1_R1138_U283 , P1_R1138_U284 , P1_R1138_U285 , P1_R1138_U286 , P1_R1138_U287;
wire P1_R1138_U288 , P1_R1138_U289 , P1_R1138_U290 , P1_R1138_U291 , P1_R1138_U292 , P1_R1138_U293 , P1_R1138_U294 , P1_R1138_U295 , P1_R1138_U296 , P1_R1138_U297;
wire P1_R1138_U298 , P1_R1138_U299 , P1_R1138_U300 , P1_R1138_U301 , P1_R1138_U302 , P1_R1138_U303 , P1_R1138_U304 , P1_R1138_U305 , P1_R1138_U306 , P1_R1138_U307;
wire P1_R1138_U308 , P1_R1138_U309 , P1_R1138_U310 , P1_R1138_U311 , P1_R1138_U312 , P1_R1138_U313 , P1_R1138_U314 , P1_R1138_U315 , P1_R1138_U316 , P1_R1138_U317;
wire P1_R1138_U318 , P1_R1138_U319 , P1_R1138_U320 , P1_R1138_U321 , P1_R1138_U322 , P1_R1138_U323 , P1_R1138_U324 , P1_R1138_U325 , P1_R1138_U326 , P1_R1138_U327;
wire P1_R1138_U328 , P1_R1138_U329 , P1_R1138_U330 , P1_R1138_U331 , P1_R1138_U332 , P1_R1138_U333 , P1_R1138_U334 , P1_R1138_U335 , P1_R1138_U336 , P1_R1138_U337;
wire P1_R1138_U338 , P1_R1138_U339 , P1_R1138_U340 , P1_R1138_U341 , P1_R1138_U342 , P1_R1138_U343 , P1_R1138_U344 , P1_R1138_U345 , P1_R1138_U346 , P1_R1138_U347;
wire P1_R1138_U348 , P1_R1138_U349 , P1_R1138_U350 , P1_R1138_U351 , P1_R1138_U352 , P1_R1138_U353 , P1_R1138_U354 , P1_R1138_U355 , P1_R1138_U356 , P1_R1138_U357;
wire P1_R1138_U358 , P1_R1138_U359 , P1_R1138_U360 , P1_R1138_U361 , P1_R1138_U362 , P1_R1138_U363 , P1_R1138_U364 , P1_R1138_U365 , P1_R1138_U366 , P1_R1138_U367;
wire P1_R1138_U368 , P1_R1138_U369 , P1_R1138_U370 , P1_R1138_U371 , P1_R1138_U372 , P1_R1138_U373 , P1_R1138_U374 , P1_R1138_U375 , P1_R1138_U376 , P1_R1138_U377;
wire P1_R1138_U378 , P1_R1138_U379 , P1_R1138_U380 , P1_R1138_U381 , P1_R1138_U382 , P1_R1138_U383 , P1_R1138_U384 , P1_R1138_U385 , P1_R1138_U386 , P1_R1138_U387;
wire P1_R1138_U388 , P1_R1138_U389 , P1_R1138_U390 , P1_R1138_U391 , P1_R1138_U392 , P1_R1138_U393 , P1_R1138_U394 , P1_R1138_U395 , P1_R1138_U396 , P1_R1138_U397;
wire P1_R1138_U398 , P1_R1138_U399 , P1_R1138_U400 , P1_R1138_U401 , P1_R1138_U402 , P1_R1138_U403 , P1_R1138_U404 , P1_R1138_U405 , P1_R1138_U406 , P1_R1138_U407;
wire P1_R1138_U408 , P1_R1138_U409 , P1_R1138_U410 , P1_R1138_U411 , P1_R1138_U412 , P1_R1138_U413 , P1_R1138_U414 , P1_R1138_U415 , P1_R1138_U416 , P1_R1138_U417;
wire P1_R1138_U418 , P1_R1138_U419 , P1_R1138_U420 , P1_R1138_U421 , P1_R1138_U422 , P1_R1138_U423 , P1_R1138_U424 , P1_R1138_U425 , P1_R1138_U426 , P1_R1138_U427;
wire P1_R1138_U428 , P1_R1138_U429 , P1_R1138_U430 , P1_R1138_U431 , P1_R1138_U432 , P1_R1138_U433 , P1_R1138_U434 , P1_R1138_U435 , P1_R1138_U436 , P1_R1138_U437;
wire P1_R1138_U438 , P1_R1138_U439 , P1_R1138_U440 , P1_R1138_U441 , P1_R1138_U442 , P1_R1138_U443 , P1_R1138_U444 , P1_R1138_U445 , P1_R1138_U446 , P1_R1138_U447;
wire P1_R1138_U448 , P1_R1138_U449 , P1_R1138_U450 , P1_R1138_U451 , P1_R1138_U452 , P1_R1138_U453 , P1_R1138_U454 , P1_R1138_U455 , P1_R1138_U456 , P1_R1138_U457;
wire P1_R1138_U458 , P1_R1138_U459 , P1_R1138_U460 , P1_R1138_U461 , P1_R1138_U462 , P1_R1138_U463 , P1_R1138_U464 , P1_R1138_U465 , P1_R1138_U466 , P1_R1138_U467;
wire P1_R1138_U468 , P1_R1138_U469 , P1_R1138_U470 , P1_R1138_U471 , P1_R1138_U472 , P1_R1138_U473 , P1_R1138_U474 , P1_R1138_U475 , P1_R1138_U476 , P1_R1138_U477;
wire P1_R1138_U478 , P1_R1138_U479 , P1_R1138_U480 , P1_R1138_U481 , P1_R1138_U482 , P1_R1138_U483 , P1_R1138_U484 , P1_R1138_U485 , P1_R1138_U486 , P1_R1138_U487;
wire P1_R1138_U488 , P1_R1138_U489 , P1_R1138_U490 , P1_R1138_U491 , P1_R1138_U492 , P1_R1138_U493 , P1_R1138_U494 , P1_R1138_U495 , P1_R1138_U496 , P1_R1138_U497;
wire P1_R1138_U498 , P1_R1138_U499 , P1_R1138_U500 , P1_R1138_U501 , P1_R1138_U502 , P1_R1138_U503 , P1_R1222_U4 , P1_R1222_U5 , P1_R1222_U6 , P1_R1222_U7;
wire P1_R1222_U8 , P1_R1222_U9 , P1_R1222_U10 , P1_R1222_U11 , P1_R1222_U12 , P1_R1222_U13 , P1_R1222_U14 , P1_R1222_U15 , P1_R1222_U16 , P1_R1222_U17;
wire P1_R1222_U18 , P1_R1222_U19 , P1_R1222_U20 , P1_R1222_U21 , P1_R1222_U22 , P1_R1222_U23 , P1_R1222_U24 , P1_R1222_U25 , P1_R1222_U26 , P1_R1222_U27;
wire P1_R1222_U28 , P1_R1222_U29 , P1_R1222_U30 , P1_R1222_U31 , P1_R1222_U32 , P1_R1222_U33 , P1_R1222_U34 , P1_R1222_U35 , P1_R1222_U36 , P1_R1222_U37;
wire P1_R1222_U38 , P1_R1222_U39 , P1_R1222_U40 , P1_R1222_U41 , P1_R1222_U42 , P1_R1222_U43 , P1_R1222_U44 , P1_R1222_U45 , P1_R1222_U46 , P1_R1222_U47;
wire P1_R1222_U48 , P1_R1222_U49 , P1_R1222_U50 , P1_R1222_U51 , P1_R1222_U52 , P1_R1222_U53 , P1_R1222_U54 , P1_R1222_U55 , P1_R1222_U56 , P1_R1222_U57;
wire P1_R1222_U58 , P1_R1222_U59 , P1_R1222_U60 , P1_R1222_U61 , P1_R1222_U62 , P1_R1222_U63 , P1_R1222_U64 , P1_R1222_U65 , P1_R1222_U66 , P1_R1222_U67;
wire P1_R1222_U68 , P1_R1222_U69 , P1_R1222_U70 , P1_R1222_U71 , P1_R1222_U72 , P1_R1222_U73 , P1_R1222_U74 , P1_R1222_U75 , P1_R1222_U76 , P1_R1222_U77;
wire P1_R1222_U78 , P1_R1222_U79 , P1_R1222_U80 , P1_R1222_U81 , P1_R1222_U82 , P1_R1222_U83 , P1_R1222_U84 , P1_R1222_U85 , P1_R1222_U86 , P1_R1222_U87;
wire P1_R1222_U88 , P1_R1222_U89 , P1_R1222_U90 , P1_R1222_U91 , P1_R1222_U92 , P1_R1222_U93 , P1_R1222_U94 , P1_R1222_U95 , P1_R1222_U96 , P1_R1222_U97;
wire P1_R1222_U98 , P1_R1222_U99 , P1_R1222_U100 , P1_R1222_U101 , P1_R1222_U102 , P1_R1222_U103 , P1_R1222_U104 , P1_R1222_U105 , P1_R1222_U106 , P1_R1222_U107;
wire P1_R1222_U108 , P1_R1222_U109 , P1_R1222_U110 , P1_R1222_U111 , P1_R1222_U112 , P1_R1222_U113 , P1_R1222_U114 , P1_R1222_U115 , P1_R1222_U116 , P1_R1222_U117;
wire P1_R1222_U118 , P1_R1222_U119 , P1_R1222_U120 , P1_R1222_U121 , P1_R1222_U122 , P1_R1222_U123 , P1_R1222_U124 , P1_R1222_U125 , P1_R1222_U126 , P1_R1222_U127;
wire P1_R1222_U128 , P1_R1222_U129 , P1_R1222_U130 , P1_R1222_U131 , P1_R1222_U132 , P1_R1222_U133 , P1_R1222_U134 , P1_R1222_U135 , P1_R1222_U136 , P1_R1222_U137;
wire P1_R1222_U138 , P1_R1222_U139 , P1_R1222_U140 , P1_R1222_U141 , P1_R1222_U142 , P1_R1222_U143 , P1_R1222_U144 , P1_R1222_U145 , P1_R1222_U146 , P1_R1222_U147;
wire P1_R1222_U148 , P1_R1222_U149 , P1_R1222_U150 , P1_R1222_U151 , P1_R1222_U152 , P1_R1222_U153 , P1_R1222_U154 , P1_R1222_U155 , P1_R1222_U156 , P1_R1222_U157;
wire P1_R1222_U158 , P1_R1222_U159 , P1_R1222_U160 , P1_R1222_U161 , P1_R1222_U162 , P1_R1222_U163 , P1_R1222_U164 , P1_R1222_U165 , P1_R1222_U166 , P1_R1222_U167;
wire P1_R1222_U168 , P1_R1222_U169 , P1_R1222_U170 , P1_R1222_U171 , P1_R1222_U172 , P1_R1222_U173 , P1_R1222_U174 , P1_R1222_U175 , P1_R1222_U176 , P1_R1222_U177;
wire P1_R1222_U178 , P1_R1222_U179 , P1_R1222_U180 , P1_R1222_U181 , P1_R1222_U182 , P1_R1222_U183 , P1_R1222_U184 , P1_R1222_U185 , P1_R1222_U186 , P1_R1222_U187;
wire P1_R1222_U188 , P1_R1222_U189 , P1_R1222_U190 , P1_R1222_U191 , P1_R1222_U192 , P1_R1222_U193 , P1_R1222_U194 , P1_R1222_U195 , P1_R1222_U196 , P1_R1222_U197;
wire P1_R1222_U198 , P1_R1222_U199 , P1_R1222_U200 , P1_R1222_U201 , P1_R1222_U202 , P1_R1222_U203 , P1_R1222_U204 , P1_R1222_U205 , P1_R1222_U206 , P1_R1222_U207;
wire P1_R1222_U208 , P1_R1222_U209 , P1_R1222_U210 , P1_R1222_U211 , P1_R1222_U212 , P1_R1222_U213 , P1_R1222_U214 , P1_R1222_U215 , P1_R1222_U216 , P1_R1222_U217;
wire P1_R1222_U218 , P1_R1222_U219 , P1_R1222_U220 , P1_R1222_U221 , P1_R1222_U222 , P1_R1222_U223 , P1_R1222_U224 , P1_R1222_U225 , P1_R1222_U226 , P1_R1222_U227;
wire P1_R1222_U228 , P1_R1222_U229 , P1_R1222_U230 , P1_R1222_U231 , P1_R1222_U232 , P1_R1222_U233 , P1_R1222_U234 , P1_R1222_U235 , P1_R1222_U236 , P1_R1222_U237;
wire P1_R1222_U238 , P1_R1222_U239 , P1_R1222_U240 , P1_R1222_U241 , P1_R1222_U242 , P1_R1222_U243 , P1_R1222_U244 , P1_R1222_U245 , P1_R1222_U246 , P1_R1222_U247;
wire P1_R1222_U248 , P1_R1222_U249 , P1_R1222_U250 , P1_R1222_U251 , P1_R1222_U252 , P1_R1222_U253 , P1_R1222_U254 , P1_R1222_U255 , P1_R1222_U256 , P1_R1222_U257;
wire P1_R1222_U258 , P1_R1222_U259 , P1_R1222_U260 , P1_R1222_U261 , P1_R1222_U262 , P1_R1222_U263 , P1_R1222_U264 , P1_R1222_U265 , P1_R1222_U266 , P1_R1222_U267;
wire P1_R1222_U268 , P1_R1222_U269 , P1_R1222_U270 , P1_R1222_U271 , P1_R1222_U272 , P1_R1222_U273 , P1_R1222_U274 , P1_R1222_U275 , P1_R1222_U276 , P1_R1222_U277;
wire P1_R1222_U278 , P1_R1222_U279 , P1_R1222_U280 , P1_R1222_U281 , P1_R1222_U282 , P1_R1222_U283 , P1_R1222_U284 , P1_R1222_U285 , P1_R1222_U286 , P1_R1222_U287;
wire P1_R1222_U288 , P1_R1222_U289 , P1_R1222_U290 , P1_R1222_U291 , P1_R1222_U292 , P1_R1222_U293 , P1_R1222_U294 , P1_R1222_U295 , P1_R1222_U296 , P1_R1222_U297;
wire P1_R1222_U298 , P1_R1222_U299 , P1_R1222_U300 , P1_R1222_U301 , P1_R1222_U302 , P1_R1222_U303 , P1_R1222_U304 , P1_R1222_U305 , P1_R1222_U306 , P1_R1222_U307;
wire P1_R1222_U308 , P1_R1222_U309 , P1_R1222_U310 , P1_R1222_U311 , P1_R1222_U312 , P1_R1222_U313 , P1_R1222_U314 , P1_R1222_U315 , P1_R1222_U316 , P1_R1222_U317;
wire P1_R1222_U318 , P1_R1222_U319 , P1_R1222_U320 , P1_R1222_U321 , P1_R1222_U322 , P1_R1222_U323 , P1_R1222_U324 , P1_R1222_U325 , P1_R1222_U326 , P1_R1222_U327;
wire P1_R1222_U328 , P1_R1222_U329 , P1_R1222_U330 , P1_R1222_U331 , P1_R1222_U332 , P1_R1222_U333 , P1_R1222_U334 , P1_R1222_U335 , P1_R1222_U336 , P1_R1222_U337;
wire P1_R1222_U338 , P1_R1222_U339 , P1_R1222_U340 , P1_R1222_U341 , P1_R1222_U342 , P1_R1222_U343 , P1_R1222_U344 , P1_R1222_U345 , P1_R1222_U346 , P1_R1222_U347;
wire P1_R1222_U348 , P1_R1222_U349 , P1_R1222_U350 , P1_R1222_U351 , P1_R1222_U352 , P1_R1222_U353 , P1_R1222_U354 , P1_R1222_U355 , P1_R1222_U356 , P1_R1222_U357;
wire P1_R1222_U358 , P1_R1222_U359 , P1_R1222_U360 , P1_R1222_U361 , P1_R1222_U362 , P1_R1222_U363 , P1_R1222_U364 , P1_R1222_U365 , P1_R1222_U366 , P1_R1222_U367;
wire P1_R1222_U368 , P1_R1222_U369 , P1_R1222_U370 , P1_R1222_U371 , P1_R1222_U372 , P1_R1222_U373 , P1_R1222_U374 , P1_R1222_U375 , P1_R1222_U376 , P1_R1222_U377;
wire P1_R1222_U378 , P1_R1222_U379 , P1_R1222_U380 , P1_R1222_U381 , P1_R1222_U382 , P1_R1222_U383 , P1_R1222_U384 , P1_R1222_U385 , P1_R1222_U386 , P1_R1222_U387;
wire P1_R1222_U388 , P1_R1222_U389 , P1_R1222_U390 , P1_R1222_U391 , P1_R1222_U392 , P1_R1222_U393 , P1_R1222_U394 , P1_R1222_U395 , P1_R1222_U396 , P1_R1222_U397;
wire P1_R1222_U398 , P1_R1222_U399 , P1_R1222_U400 , P1_R1222_U401 , P1_R1222_U402 , P1_R1222_U403 , P1_R1222_U404 , P1_R1222_U405 , P1_R1222_U406 , P1_R1222_U407;
wire P1_R1222_U408 , P1_R1222_U409 , P1_R1222_U410 , P1_R1222_U411 , P1_R1222_U412 , P1_R1222_U413 , P1_R1222_U414 , P1_R1222_U415 , P1_R1222_U416 , P1_R1222_U417;
wire P1_R1222_U418 , P1_R1222_U419 , P1_R1222_U420 , P1_R1222_U421 , P1_R1222_U422 , P1_R1222_U423 , P1_R1222_U424 , P1_R1222_U425 , P1_R1222_U426 , P1_R1222_U427;
wire P1_R1222_U428 , P1_R1222_U429 , P1_R1222_U430 , P1_R1222_U431 , P1_R1222_U432 , P1_R1222_U433 , P1_R1222_U434 , P1_R1222_U435 , P1_R1222_U436 , P1_R1222_U437;
wire P1_R1222_U438 , P1_R1222_U439 , P1_R1222_U440 , P1_R1222_U441 , P1_R1222_U442 , P1_R1222_U443 , P1_R1222_U444 , P1_R1222_U445 , P1_R1222_U446 , P1_R1222_U447;
wire P1_R1222_U448 , P1_R1222_U449 , P1_R1222_U450 , P1_R1222_U451 , P1_R1222_U452 , P1_R1222_U453 , P1_R1222_U454 , P1_R1222_U455 , P1_R1222_U456 , P1_R1222_U457;
wire P1_R1222_U458 , P1_R1222_U459 , P1_R1222_U460 , P1_R1222_U461 , P1_R1222_U462 , P1_R1222_U463 , P1_R1222_U464 , P1_R1222_U465 , P1_R1222_U466 , P1_R1222_U467;
wire P1_R1222_U468 , P1_R1222_U469 , P1_R1222_U470 , P1_R1222_U471 , P1_R1222_U472 , P1_R1222_U473 , P1_R1222_U474 , P1_R1222_U475 , P1_R1222_U476 , P1_R1222_U477;
wire P1_R1222_U478 , P1_R1222_U479 , P1_R1222_U480 , P1_R1222_U481 , P1_R1222_U482 , P1_R1222_U483 , P1_R1222_U484 , P1_R1222_U485 , P1_R1222_U486 , P1_R1222_U487;
wire P1_R1222_U488 , P1_R1222_U489 , P1_R1222_U490 , P1_R1222_U491 , P1_R1222_U492 , P1_R1222_U493 , P1_R1222_U494 , P1_R1222_U495 , P1_R1222_U496 , P1_R1222_U497;
wire P1_R1222_U498 , P1_R1222_U499 , P1_R1222_U500 , P1_R1222_U501 , P1_R1222_U502 , P1_R1222_U503 , P2_SUB_594_U6 , P2_SUB_594_U7 , P2_SUB_594_U8 , P2_SUB_594_U9;
wire P2_SUB_594_U10 , P2_SUB_594_U11 , P2_SUB_594_U12 , P2_SUB_594_U13 , P2_SUB_594_U14 , P2_SUB_594_U15 , P2_SUB_594_U16 , P2_SUB_594_U17 , P2_SUB_594_U18 , P2_SUB_594_U19;
wire P2_SUB_594_U20 , P2_SUB_594_U21 , P2_SUB_594_U22 , P2_SUB_594_U23 , P2_SUB_594_U24 , P2_SUB_594_U25 , P2_SUB_594_U26 , P2_SUB_594_U27 , P2_SUB_594_U28 , P2_SUB_594_U29;
wire P2_SUB_594_U30 , P2_SUB_594_U31 , P2_SUB_594_U32 , P2_SUB_594_U33 , P2_SUB_594_U34 , P2_SUB_594_U35 , P2_SUB_594_U36 , P2_SUB_594_U37 , P2_SUB_594_U38 , P2_SUB_594_U39;
wire P2_SUB_594_U40 , P2_SUB_594_U41 , P2_SUB_594_U42 , P2_SUB_594_U43 , P2_SUB_594_U44 , P2_SUB_594_U45 , P2_SUB_594_U46 , P2_SUB_594_U47 , P2_SUB_594_U48 , P2_SUB_594_U49;
wire P2_SUB_594_U50 , P2_SUB_594_U51 , P2_SUB_594_U52 , P2_SUB_594_U53 , P2_SUB_594_U54 , P2_SUB_594_U55 , P2_SUB_594_U56 , P2_SUB_594_U57 , P2_SUB_594_U58 , P2_SUB_594_U59;
wire P2_SUB_594_U60 , P2_SUB_594_U61 , P2_SUB_594_U62 , P2_SUB_594_U63 , P2_SUB_594_U64 , P2_SUB_594_U65 , P2_SUB_594_U66 , P2_SUB_594_U67 , P2_SUB_594_U68 , P2_SUB_594_U69;
wire P2_SUB_594_U70 , P2_SUB_594_U71 , P2_SUB_594_U72 , P2_SUB_594_U73 , P2_SUB_594_U74 , P2_SUB_594_U75 , P2_SUB_594_U76 , P2_SUB_594_U77 , P2_SUB_594_U78 , P2_SUB_594_U79;
wire P2_SUB_594_U80 , P2_SUB_594_U81 , P2_SUB_594_U82 , P2_SUB_594_U83 , P2_SUB_594_U84 , P2_SUB_594_U85 , P2_SUB_594_U86 , P2_SUB_594_U87 , P2_SUB_594_U88 , P2_SUB_594_U89;
wire P2_SUB_594_U90 , P2_SUB_594_U91 , P2_SUB_594_U92 , P2_SUB_594_U93 , P2_SUB_594_U94 , P2_SUB_594_U95 , P2_SUB_594_U96 , P2_SUB_594_U97 , P2_SUB_594_U98 , P2_SUB_594_U99;
wire P2_SUB_594_U100 , P2_SUB_594_U101 , P2_SUB_594_U102 , P2_SUB_594_U103 , P2_SUB_594_U104 , P2_SUB_594_U105 , P2_SUB_594_U106 , P2_SUB_594_U107 , P2_SUB_594_U108 , P2_SUB_594_U109;
wire P2_SUB_594_U110 , P2_SUB_594_U111 , P2_SUB_594_U112 , P2_SUB_594_U113 , P2_SUB_594_U114 , P2_SUB_594_U115 , P2_SUB_594_U116 , P2_SUB_594_U117 , P2_SUB_594_U118 , P2_SUB_594_U119;
wire P2_SUB_594_U120 , P2_SUB_594_U121 , P2_SUB_594_U122 , P2_SUB_594_U123 , P2_SUB_594_U124 , P2_SUB_594_U125 , P2_SUB_594_U126 , P2_SUB_594_U127 , P2_SUB_594_U128 , P2_SUB_594_U129;
wire P2_SUB_594_U130 , P2_SUB_594_U131 , P2_SUB_594_U132 , P2_SUB_594_U133 , P2_SUB_594_U134 , P2_SUB_594_U135 , P2_SUB_594_U136 , P2_SUB_594_U137 , P2_SUB_594_U138 , P2_SUB_594_U139;
wire P2_SUB_594_U140 , P2_SUB_594_U141 , P2_SUB_594_U142 , P2_SUB_594_U143 , P2_SUB_594_U144 , P2_SUB_594_U145 , P2_SUB_594_U146 , P2_SUB_594_U147 , P2_SUB_594_U148 , P2_SUB_594_U149;
wire P2_SUB_594_U150 , P2_SUB_594_U151 , P2_SUB_594_U152 , P2_SUB_594_U153 , P2_SUB_594_U154 , P2_SUB_594_U155 , P2_SUB_594_U156 , P2_SUB_594_U157 , P2_SUB_594_U158 , P2_R693_U6;
wire P2_R693_U7 , P2_R693_U8 , P2_R693_U9 , P2_R693_U10 , P2_R693_U11 , P2_R693_U12 , P2_R693_U13 , P2_R693_U14 , P2_R693_U15 , P2_R693_U16;
wire P2_R693_U17 , P2_R693_U18 , P2_R693_U19 , P2_R693_U20 , P2_R693_U21 , P2_R693_U22 , P2_R693_U23 , P2_R693_U24 , P2_R693_U25 , P2_R693_U26;
wire P2_R693_U27 , P2_R693_U28 , P2_R693_U29 , P2_R693_U30 , P2_R693_U31 , P2_R693_U32 , P2_R693_U33 , P2_R693_U34 , P2_R693_U35 , P2_R693_U36;
wire P2_R693_U37 , P2_R693_U38 , P2_R693_U39 , P2_R693_U40 , P2_R693_U41 , P2_R693_U42 , P2_R693_U43 , P2_R693_U44 , P2_R693_U45 , P2_R693_U46;
wire P2_R693_U47 , P2_R693_U48 , P2_R693_U49 , P2_R693_U50 , P2_R693_U51 , P2_R693_U52 , P2_R693_U53 , P2_R693_U54 , P2_R693_U55 , P2_R693_U56;
wire P2_R693_U57 , P2_R693_U58 , P2_R693_U59 , P2_R693_U60 , P2_R693_U61 , P2_R693_U62 , P2_R693_U63 , P2_R693_U64 , P2_R693_U65 , P2_R693_U66;
wire P2_R693_U67 , P2_R693_U68 , P2_R693_U69 , P2_R693_U70 , P2_R693_U71 , P2_R693_U72 , P2_R693_U73 , P2_R693_U74 , P2_R693_U75 , P2_R693_U76;
wire P2_R693_U77 , P2_R693_U78 , P2_R693_U79 , P2_R693_U80 , P2_R693_U81 , P2_R693_U82 , P2_R693_U83 , P2_R693_U84 , P2_R693_U85 , P2_R693_U86;
wire P2_R693_U87 , P2_R693_U88 , P2_R693_U89 , P2_R693_U90 , P2_R693_U91 , P2_R693_U92 , P2_R693_U93 , P2_R693_U94 , P2_R693_U95 , P2_R693_U96;
wire P2_R693_U97 , P2_R693_U98 , P2_R693_U99 , P2_R693_U100 , P2_R693_U101 , P2_R693_U102 , P2_R693_U103 , P2_R693_U104 , P2_R693_U105 , P2_R693_U106;
wire P2_R693_U107 , P2_R693_U108 , P2_R693_U109 , P2_R693_U110 , P2_R693_U111 , P2_R693_U112 , P2_R693_U113 , P2_R693_U114 , P2_R693_U115 , P2_R693_U116;
wire P2_R693_U117 , P2_R693_U118 , P2_R693_U119 , P2_R693_U120 , P2_R693_U121 , P2_R693_U122 , P2_R693_U123 , P2_R693_U124 , P2_R693_U125 , P2_R693_U126;
wire P2_R693_U127 , P2_R693_U128 , P2_R693_U129 , P2_R693_U130 , P2_R693_U131 , P2_R693_U132 , P2_R693_U133 , P2_R693_U134 , P2_R693_U135 , P2_R693_U136;
wire P2_R693_U137 , P2_R693_U138 , P2_R693_U139 , P2_R693_U140 , P2_R693_U141 , P2_R693_U142 , P2_R693_U143 , P2_R693_U144 , P2_R693_U145 , P2_R693_U146;
wire P2_R693_U147 , P2_R693_U148 , P2_R693_U149 , P2_R693_U150 , P2_R693_U151 , P2_R693_U152 , P2_R693_U153 , P2_R693_U154 , P2_R693_U155 , P2_R693_U156;
wire P2_R693_U157 , P2_R693_U158 , P2_R693_U159 , P2_R693_U160 , P2_R693_U161 , P2_R693_U162 , P2_R693_U163 , P2_R693_U164 , P2_R693_U165 , P2_R693_U166;
wire P2_R693_U167 , P2_R693_U168 , P2_R693_U169 , P2_R693_U170 , P2_R693_U171 , P2_R693_U172 , P2_R693_U173 , P2_R693_U174 , P2_R693_U175 , P2_R693_U176;
wire P2_R693_U177 , P2_R693_U178 , P2_R693_U179 , P2_R693_U180 , P2_R693_U181 , P2_R693_U182 , P2_R693_U183 , P2_R693_U184 , P2_R693_U185 , P2_R693_U186;
wire P2_R693_U187 , P2_R693_U188 , P2_R693_U189 , P2_R693_U190 , P2_R693_U191 , P2_R693_U192 , P2_R693_U193 , P2_SUB_605_U6 , P2_SUB_605_U7 , P2_SUB_605_U8;
wire P2_SUB_605_U9 , P2_SUB_605_U10 , P2_SUB_605_U11 , P2_SUB_605_U12 , P2_SUB_605_U13 , P2_SUB_605_U14 , P2_SUB_605_U15 , P2_SUB_605_U16 , P2_SUB_605_U17 , P2_SUB_605_U18;
wire P2_SUB_605_U19 , P2_SUB_605_U20 , P2_SUB_605_U21 , P2_SUB_605_U22 , P2_SUB_605_U23 , P2_SUB_605_U24 , P2_SUB_605_U25 , P2_SUB_605_U26 , P2_SUB_605_U27 , P2_SUB_605_U28;
wire P2_SUB_605_U29 , P2_SUB_605_U30 , P2_SUB_605_U31 , P2_SUB_605_U32 , P2_SUB_605_U33 , P2_SUB_605_U34 , P2_SUB_605_U35 , P2_SUB_605_U36 , P2_SUB_605_U37 , P2_SUB_605_U38;
wire P2_SUB_605_U39 , P2_SUB_605_U40 , P2_SUB_605_U41 , P2_SUB_605_U42 , P2_SUB_605_U43 , P2_SUB_605_U44 , P2_SUB_605_U45 , P2_SUB_605_U46 , P2_SUB_605_U47 , P2_SUB_605_U48;
wire P2_SUB_605_U49 , P2_SUB_605_U50 , P2_SUB_605_U51 , P2_SUB_605_U52 , P2_SUB_605_U53 , P2_SUB_605_U54 , P2_SUB_605_U55 , P2_SUB_605_U56 , P2_SUB_605_U57 , P2_SUB_605_U58;
wire P2_SUB_605_U59 , P2_SUB_605_U60 , P2_SUB_605_U61 , P2_SUB_605_U62 , P2_SUB_605_U63 , P2_SUB_605_U64 , P2_SUB_605_U65 , P2_SUB_605_U66 , P2_SUB_605_U67 , P2_SUB_605_U68;
wire P2_SUB_605_U69 , P2_SUB_605_U70 , P2_SUB_605_U71 , P2_SUB_605_U72 , P2_SUB_605_U73 , P2_SUB_605_U74 , P2_SUB_605_U75 , P2_SUB_605_U76 , P2_SUB_605_U77 , P2_SUB_605_U78;
wire P2_SUB_605_U79 , P2_SUB_605_U80 , P2_SUB_605_U81 , P2_SUB_605_U82 , P2_SUB_605_U83 , P2_SUB_605_U84 , P2_SUB_605_U85 , P2_SUB_605_U86 , P2_SUB_605_U87 , P2_SUB_605_U88;
wire P2_SUB_605_U89 , P2_SUB_605_U90 , P2_SUB_605_U91 , P2_SUB_605_U92 , P2_SUB_605_U93 , P2_SUB_605_U94 , P2_SUB_605_U95 , P2_SUB_605_U96 , P2_SUB_605_U97 , P2_SUB_605_U98;
wire P2_SUB_605_U99 , P2_SUB_605_U100 , P2_SUB_605_U101 , P2_SUB_605_U102 , P2_SUB_605_U103 , P2_SUB_605_U104 , P2_SUB_605_U105 , P2_SUB_605_U106 , P2_SUB_605_U107 , P2_SUB_605_U108;
wire P2_SUB_605_U109 , P2_SUB_605_U110 , P2_SUB_605_U111 , P2_SUB_605_U112 , P2_SUB_605_U113 , P2_R1095_U6 , P2_R1095_U7 , P2_R1095_U8 , P2_R1095_U9 , P2_R1095_U10;
wire P2_R1095_U11 , P2_R1095_U12 , P2_R1095_U13 , P2_R1095_U14 , P2_R1095_U15 , P2_R1095_U16 , P2_R1095_U17 , P2_R1095_U18 , P2_R1095_U19 , P2_R1095_U20;
wire P2_R1095_U21 , P2_R1095_U22 , P2_R1095_U23 , P2_R1095_U24 , P2_R1095_U25 , P2_R1095_U26 , P2_R1095_U27 , P2_R1095_U28 , P2_R1095_U29 , P2_R1095_U30;
wire P2_R1095_U31 , P2_R1095_U32 , P2_R1095_U33 , P2_R1095_U34 , P2_R1095_U35 , P2_R1095_U36 , P2_R1095_U37 , P2_R1095_U38 , P2_R1095_U39 , P2_R1095_U40;
wire P2_R1095_U41 , P2_R1095_U42 , P2_R1095_U43 , P2_R1095_U44 , P2_R1095_U45 , P2_R1095_U46 , P2_R1095_U47 , P2_R1095_U48 , P2_R1095_U49 , P2_R1095_U50;
wire P2_R1095_U51 , P2_R1095_U52 , P2_R1095_U53 , P2_R1095_U54 , P2_R1095_U55 , P2_R1095_U56 , P2_R1095_U57 , P2_R1095_U58 , P2_R1095_U59 , P2_R1095_U60;
wire P2_R1095_U61 , P2_R1095_U62 , P2_R1095_U63 , P2_R1095_U64 , P2_R1095_U65 , P2_R1095_U66 , P2_R1095_U67 , P2_R1095_U68 , P2_R1095_U69 , P2_R1095_U70;
wire P2_R1095_U71 , P2_R1095_U72 , P2_R1095_U73 , P2_R1095_U74 , P2_R1095_U75 , P2_R1095_U76 , P2_R1095_U77 , P2_R1095_U78 , P2_R1095_U79 , P2_R1095_U80;
wire P2_R1095_U81 , P2_R1095_U82 , P2_R1095_U83 , P2_R1095_U84 , P2_R1095_U85 , P2_R1095_U86 , P2_R1095_U87 , P2_R1095_U88 , P2_R1095_U89 , P2_R1095_U90;
wire P2_R1095_U91 , P2_R1095_U92 , P2_R1095_U93 , P2_R1095_U94 , P2_R1095_U95 , P2_R1095_U96 , P2_R1095_U97 , P2_R1095_U98 , P2_R1095_U99 , P2_R1095_U100;
wire P2_R1095_U101 , P2_R1095_U102 , P2_R1095_U103 , P2_R1095_U104 , P2_R1095_U105 , P2_R1095_U106 , P2_R1095_U107 , P2_R1095_U108 , P2_R1095_U109 , P2_R1095_U110;
wire P2_R1095_U111 , P2_R1095_U112 , P2_R1095_U113 , P2_R1095_U114 , P2_R1095_U115 , P2_R1095_U116 , P2_R1095_U117 , P2_R1095_U118 , P2_R1095_U119 , P2_R1095_U120;
wire P2_R1095_U121 , P2_R1095_U122 , P2_R1095_U123 , P2_R1095_U124 , P2_R1095_U125 , P2_R1095_U126 , P2_R1095_U127 , P2_R1095_U128 , P2_R1095_U129 , P2_R1095_U130;
wire P2_R1095_U131 , P2_R1095_U132 , P2_R1095_U133 , P2_R1095_U134 , P2_R1095_U135 , P2_R1095_U136 , P2_R1095_U137 , P2_R1095_U138 , P2_R1095_U139 , P2_R1095_U140;
wire P2_R1095_U141 , P2_R1095_U142 , P2_R1095_U143 , P2_R1095_U144 , P2_R1095_U145 , P2_R1095_U146 , P2_R1095_U147 , P2_R1095_U148 , P2_R1095_U149 , P2_R1095_U150;
wire P2_R1095_U151 , P2_R1095_U152 , P2_R1095_U153 , P2_R1095_U154 , P2_R1095_U155 , P2_R1095_U156 , P2_R1095_U157 , P2_R1095_U158 , P2_R1095_U159 , P2_R1095_U160;
wire P2_R1095_U161 , P2_R1095_U162 , P2_R1095_U163 , P2_R1095_U164 , P2_R1095_U165 , P2_R1095_U166 , P2_R1095_U167 , P2_R1095_U168 , P2_R1095_U169 , P2_R1095_U170;
wire P2_R1095_U171 , P2_R1095_U172 , P2_R1095_U173 , P2_R1095_U174 , P2_R1095_U175 , P2_R1095_U176 , P2_R1095_U177 , P2_R1095_U178 , P2_R1095_U179 , P2_R1095_U180;
wire P2_R1095_U181 , P2_R1095_U182 , P2_R1095_U183 , P2_R1095_U184 , P2_R1095_U185 , P2_R1095_U186 , P2_R1095_U187 , P2_R1095_U188 , P2_R1095_U189 , P2_R1095_U190;
wire P2_R1095_U191 , P2_R1095_U192 , P2_R1095_U193 , P2_R1095_U194 , P2_R1095_U195 , P2_R1095_U196 , P2_R1095_U197 , P2_R1095_U198 , P2_R1095_U199 , P2_R1095_U200;
wire P2_R1095_U201 , P2_R1095_U202 , P2_R1095_U203 , P2_R1095_U204 , P2_R1095_U205 , P2_R1095_U206 , P2_R1095_U207 , P2_R1095_U208 , P2_R1095_U209 , P2_R1095_U210;
wire P2_R1095_U211 , P2_R1095_U212 , P2_R1095_U213 , P2_R1095_U214 , P2_R1095_U215 , P2_R1095_U216 , P2_R1095_U217 , P2_R1095_U218 , P2_R1095_U219 , P2_R1095_U220;
wire P2_R1095_U221 , P2_R1095_U222 , P2_R1095_U223 , P2_R1095_U224 , P2_R1095_U225 , P2_R1095_U226 , P2_R1095_U227 , P2_R1095_U228 , P2_R1095_U229 , P2_R1095_U230;
wire P2_R1095_U231 , P2_R1095_U232 , P2_R1095_U233 , P2_R1095_U234 , P2_R1095_U235 , P2_R1095_U236 , P2_R1095_U237 , P2_R1095_U238 , P2_R1095_U239 , P2_R1095_U240;
wire P2_R1095_U241 , P2_R1095_U242 , P2_R1095_U243 , P2_R1095_U244 , P2_R1095_U245 , P2_R1095_U246 , P2_R1095_U247 , P2_R1095_U248 , P2_R1095_U249 , P2_R1095_U250;
wire P2_R1095_U251 , P2_R1095_U252 , P2_R1095_U253 , P2_R1095_U254 , P2_R1095_U255 , P2_R1095_U256 , P2_R1095_U257 , P2_R1095_U258 , P2_R1095_U259 , P2_R1095_U260;
wire P2_R1095_U261 , P2_R1095_U262 , P2_R1095_U263 , P2_R1095_U264 , P2_R1095_U265 , P2_R1095_U266 , P2_R1095_U267 , P2_R1095_U268 , P2_R1095_U269 , P2_R1095_U270;
wire P2_R1095_U271 , P2_R1095_U272 , P2_R1095_U273 , P2_R1095_U274 , P2_R1095_U275 , P2_R1095_U276 , P2_R1095_U277 , P2_R1095_U278 , P2_R1095_U279 , P2_R1095_U280;
wire P2_R1095_U281 , P2_R1095_U282 , P2_R1095_U283 , P2_R1095_U284 , P2_R1095_U285 , P2_R1095_U286 , P2_R1095_U287 , P2_R1095_U288 , P2_R1095_U289 , P2_R1095_U290;
wire P2_R1095_U291 , P2_R1095_U292 , P2_R1095_U293 , P2_R1095_U294 , P2_R1095_U295 , P2_R1095_U296 , P2_R1095_U297 , P2_R1095_U298 , P2_R1095_U299 , P2_R1095_U300;
wire P2_R1095_U301 , P2_R1095_U302 , P2_R1095_U303 , P2_R1095_U304 , P2_R1095_U305 , P2_R1095_U306 , P2_R1095_U307 , P2_R1095_U308 , P2_R1095_U309 , P2_R1095_U310;
wire P2_R1095_U311 , P2_R1095_U312 , P2_R1095_U313 , P2_R1095_U314 , P2_R1095_U315 , P2_R1095_U316 , P2_R1095_U317 , P2_R1095_U318 , P2_R1095_U319 , P2_R1095_U320;
wire P2_R1095_U321 , P2_R1095_U322 , P2_R1095_U323 , P2_R1095_U324 , P2_R1095_U325 , P2_R1095_U326 , P2_R1095_U327 , P2_R1095_U328 , P2_R1095_U329 , P2_R1095_U330;
wire P2_R1095_U331 , P2_R1095_U332 , P2_R1095_U333 , P2_R1095_U334 , P2_R1095_U335 , P2_R1095_U336 , P2_R1095_U337 , P2_R1095_U338 , P2_R1095_U339 , P2_R1095_U340;
wire P2_R1095_U341 , P2_R1095_U342 , P2_R1095_U343 , P2_R1095_U344 , P2_R1095_U345 , P2_R1095_U346 , P2_R1095_U347 , P2_R1095_U348 , P2_R1095_U349 , P2_R1095_U350;
wire P2_R1095_U351 , P2_R1095_U352 , P2_R1095_U353 , P2_R1095_U354 , P2_R1095_U355 , P2_R1095_U356 , P2_R1095_U357 , P2_R1095_U358 , P2_R1095_U359 , P2_R1095_U360;
wire P2_R1095_U361 , P2_R1095_U362 , P2_R1095_U363 , P2_R1095_U364 , P2_R1095_U365 , P2_R1095_U366 , P2_R1095_U367 , P2_R1095_U368 , P2_R1095_U369 , P2_R1095_U370;
wire P2_R1095_U371 , P2_R1095_U372 , P2_R1095_U373 , P2_R1095_U374 , P2_R1095_U375 , P2_R1095_U376 , P2_R1095_U377 , P2_R1095_U378 , P2_R1095_U379 , P2_R1095_U380;
wire P2_R1095_U381 , P2_R1095_U382 , P2_R1095_U383 , P2_R1095_U384 , P2_R1095_U385 , P2_R1095_U386 , P2_R1095_U387 , P2_R1095_U388 , P2_R1095_U389 , P2_R1095_U390;
wire P2_R1095_U391 , P2_R1095_U392 , P2_R1095_U393 , P2_R1095_U394 , P2_R1095_U395 , P2_R1095_U396 , P2_R1095_U397 , P2_R1095_U398 , P2_R1095_U399 , P2_R1095_U400;
wire P2_R1095_U401 , P2_R1095_U402 , P2_R1095_U403 , P2_R1095_U404 , P2_R1095_U405 , P2_R1095_U406 , P2_R1095_U407 , P2_R1095_U408 , P2_R1095_U409 , P2_R1095_U410;
wire P2_R1095_U411 , P2_R1095_U412 , P2_R1095_U413 , P2_R1095_U414 , P2_R1095_U415 , P2_R1095_U416 , P2_R1095_U417 , P2_R1095_U418 , P2_R1095_U419 , P2_R1095_U420;
wire P2_R1095_U421 , P2_R1095_U422 , P2_R1095_U423 , P2_R1095_U424 , P2_R1095_U425 , P2_R1095_U426 , P2_R1095_U427 , P2_R1095_U428 , P2_R1095_U429 , P2_R1095_U430;
wire P2_R1095_U431 , P2_R1095_U432 , P2_R1095_U433 , P2_R1095_U434 , P2_R1095_U435 , P2_R1095_U436 , P2_R1095_U437 , P2_R1095_U438 , P2_R1095_U439 , P2_R1095_U440;
wire P2_R1095_U441 , P2_R1095_U442 , P2_R1095_U443 , P2_R1095_U444 , P2_R1095_U445 , P2_R1095_U446 , P2_R1095_U447 , P2_R1095_U448 , P2_R1095_U449 , P2_R1095_U450;
wire P2_R1095_U451 , P2_R1095_U452 , P2_R1095_U453 , P2_R1095_U454 , P2_R1095_U455 , P2_R1095_U456 , P2_R1095_U457 , P2_R1095_U458 , P2_R1095_U459 , P2_R1095_U460;
wire P2_R1095_U461 , P2_R1095_U462 , P2_R1095_U463 , P2_R1095_U464 , P2_R1095_U465 , P2_R1095_U466 , P2_R1095_U467 , P2_R1095_U468 , P2_R1095_U469 , P2_R1095_U470;
wire P2_R1095_U471 , P2_R1095_U472 , P2_R1095_U473 , P2_R1095_U474 , P2_R1095_U475 , P2_R1095_U476 , P2_R1095_U477 , P2_R1095_U478 , P2_R1095_U479 , P2_R1095_U480;
wire P2_R1095_U481 , P2_R1095_U482 , P2_R1095_U483 , P2_R1095_U484 , P2_R1095_U485 , P2_R1095_U486 , P2_R1095_U487 , P2_R1095_U488 , P2_R1095_U489 , P2_R1212_U6;
wire P2_R1212_U7 , P2_R1212_U8 , P2_R1212_U9 , P2_R1212_U10 , P2_R1212_U11 , P2_R1212_U12 , P2_R1212_U13 , P2_R1212_U14 , P2_R1212_U15 , P2_R1212_U16;
wire P2_R1212_U17 , P2_R1212_U18 , P2_R1212_U19 , P2_R1212_U20 , P2_R1212_U21 , P2_R1212_U22 , P2_R1212_U23 , P2_R1212_U24 , P2_R1212_U25 , P2_R1212_U26;
wire P2_R1212_U27 , P2_R1212_U28 , P2_R1212_U29 , P2_R1212_U30 , P2_R1212_U31 , P2_R1212_U32 , P2_R1212_U33 , P2_R1212_U34 , P2_R1212_U35 , P2_R1212_U36;
wire P2_R1212_U37 , P2_R1212_U38 , P2_R1212_U39 , P2_R1212_U40 , P2_R1212_U41 , P2_R1212_U42 , P2_R1212_U43 , P2_R1212_U44 , P2_R1212_U45 , P2_R1212_U46;
wire P2_R1212_U47 , P2_R1212_U48 , P2_R1212_U49 , P2_R1212_U50 , P2_R1212_U51 , P2_R1212_U52 , P2_R1212_U53 , P2_R1212_U54 , P2_R1212_U55 , P2_R1212_U56;
wire P2_R1212_U57 , P2_R1212_U58 , P2_R1212_U59 , P2_R1212_U60 , P2_R1212_U61 , P2_R1212_U62 , P2_R1212_U63 , P2_R1212_U64 , P2_R1212_U65 , P2_R1212_U66;
wire P2_R1212_U67 , P2_R1212_U68 , P2_R1212_U69 , P2_R1212_U70 , P2_R1212_U71 , P2_R1212_U72 , P2_R1212_U73 , P2_R1212_U74 , P2_R1212_U75 , P2_R1212_U76;
wire P2_R1212_U77 , P2_R1212_U78 , P2_R1212_U79 , P2_R1212_U80 , P2_R1212_U81 , P2_R1212_U82 , P2_R1212_U83 , P2_R1212_U84 , P2_R1212_U85 , P2_R1212_U86;
wire P2_R1212_U87 , P2_R1212_U88 , P2_R1212_U89 , P2_R1212_U90 , P2_R1212_U91 , P2_R1212_U92 , P2_R1212_U93 , P2_R1212_U94 , P2_R1212_U95 , P2_R1212_U96;
wire P2_R1212_U97 , P2_R1212_U98 , P2_R1212_U99 , P2_R1212_U100 , P2_R1212_U101 , P2_R1212_U102 , P2_R1212_U103 , P2_R1212_U104 , P2_R1212_U105 , P2_R1212_U106;
wire P2_R1212_U107 , P2_R1212_U108 , P2_R1212_U109 , P2_R1212_U110 , P2_R1212_U111 , P2_R1212_U112 , P2_R1212_U113 , P2_R1212_U114 , P2_R1212_U115 , P2_R1212_U116;
wire P2_R1212_U117 , P2_R1212_U118 , P2_R1212_U119 , P2_R1212_U120 , P2_R1212_U121 , P2_R1212_U122 , P2_R1212_U123 , P2_R1212_U124 , P2_R1212_U125 , P2_R1212_U126;
wire P2_R1212_U127 , P2_R1212_U128 , P2_R1212_U129 , P2_R1212_U130 , P2_R1212_U131 , P2_R1212_U132 , P2_R1212_U133 , P2_R1212_U134 , P2_R1212_U135 , P2_R1212_U136;
wire P2_R1212_U137 , P2_R1212_U138 , P2_R1212_U139 , P2_R1212_U140 , P2_R1212_U141 , P2_R1212_U142 , P2_R1212_U143 , P2_R1212_U144 , P2_R1212_U145 , P2_R1212_U146;
wire P2_R1212_U147 , P2_R1212_U148 , P2_R1212_U149 , P2_R1212_U150 , P2_R1212_U151 , P2_R1212_U152 , P2_R1212_U153 , P2_R1212_U154 , P2_R1212_U155 , P2_R1212_U156;
wire P2_R1212_U157 , P2_R1212_U158 , P2_R1212_U159 , P2_R1212_U160 , P2_R1212_U161 , P2_R1212_U162 , P2_R1212_U163 , P2_R1212_U164 , P2_R1212_U165 , P2_R1212_U166;
wire P2_R1212_U167 , P2_R1212_U168 , P2_R1212_U169 , P2_R1212_U170 , P2_R1212_U171 , P2_R1212_U172 , P2_R1212_U173 , P2_R1212_U174 , P2_R1212_U175 , P2_R1212_U176;
wire P2_R1212_U177 , P2_R1212_U178 , P2_R1212_U179 , P2_R1212_U180 , P2_R1212_U181 , P2_R1212_U182 , P2_R1212_U183 , P2_R1212_U184 , P2_R1212_U185 , P2_R1212_U186;
wire P2_R1212_U187 , P2_R1212_U188 , P2_R1212_U189 , P2_R1212_U190 , P2_R1212_U191 , P2_R1212_U192 , P2_R1212_U193 , P2_R1212_U194 , P2_R1212_U195 , P2_R1212_U196;
wire P2_R1212_U197 , P2_R1212_U198 , P2_R1212_U199 , P2_R1212_U200 , P2_R1212_U201 , P2_R1212_U202 , P2_R1212_U203 , P2_R1212_U204 , P2_R1212_U205 , P2_R1212_U206;
wire P2_R1212_U207 , P2_R1212_U208 , P2_R1212_U209 , P2_R1212_U210 , P2_R1212_U211 , P2_R1212_U212 , P2_R1212_U213 , P2_R1212_U214 , P2_R1212_U215 , P2_R1212_U216;
wire P2_R1212_U217 , P2_R1212_U218 , P2_R1212_U219 , P2_R1212_U220 , P2_R1212_U221 , P2_R1212_U222 , P2_R1212_U223 , P2_R1212_U224 , P2_R1212_U225 , P2_R1212_U226;
wire P2_R1212_U227 , P2_R1212_U228 , P2_R1212_U229 , P2_R1212_U230 , P2_R1212_U231 , P2_R1212_U232 , P2_R1212_U233 , P2_R1212_U234 , P2_R1212_U235 , P2_R1212_U236;
wire P2_R1212_U237 , P2_R1212_U238 , P2_R1212_U239 , P2_R1212_U240 , P2_R1212_U241 , P2_R1212_U242 , P2_R1212_U243 , P2_R1212_U244 , P2_R1212_U245 , P2_R1212_U246;
wire P2_R1212_U247 , P2_R1212_U248 , P2_R1212_U249 , P2_R1212_U250 , P2_R1212_U251 , P2_R1212_U252 , P2_R1212_U253 , P2_R1212_U254 , P2_R1212_U255 , P2_R1212_U256;
wire P2_R1212_U257 , P2_R1212_U258 , P2_R1212_U259 , P2_R1212_U260 , P2_R1212_U261 , P2_R1212_U262 , P2_R1212_U263 , P2_R1212_U264 , P2_R1212_U265 , P2_R1212_U266;
wire P2_R1212_U267 , P2_R1212_U268 , P2_R1212_U269 , P2_R1212_U270 , P2_R1212_U271 , P2_R1212_U272 , P2_R1212_U273 , P2_R1212_U274 , P2_R1212_U275 , P2_R1212_U276;
wire P2_R1209_U6 , P2_R1209_U7 , P2_R1209_U8 , P2_R1209_U9 , P2_R1209_U10 , P2_R1209_U11 , P2_R1209_U12 , P2_R1209_U13 , P2_R1209_U14 , P2_R1209_U15;
wire P2_R1209_U16 , P2_R1209_U17 , P2_R1209_U18 , P2_R1209_U19 , P2_R1209_U20 , P2_R1209_U21 , P2_R1209_U22 , P2_R1209_U23 , P2_R1209_U24 , P2_R1209_U25;
wire P2_R1209_U26 , P2_R1209_U27 , P2_R1209_U28 , P2_R1209_U29 , P2_R1209_U30 , P2_R1209_U31 , P2_R1209_U32 , P2_R1209_U33 , P2_R1209_U34 , P2_R1209_U35;
wire P2_R1209_U36 , P2_R1209_U37 , P2_R1209_U38 , P2_R1209_U39 , P2_R1209_U40 , P2_R1209_U41 , P2_R1209_U42 , P2_R1209_U43 , P2_R1209_U44 , P2_R1209_U45;
wire P2_R1209_U46 , P2_R1209_U47 , P2_R1209_U48 , P2_R1209_U49 , P2_R1209_U50 , P2_R1209_U51 , P2_R1209_U52 , P2_R1209_U53 , P2_R1209_U54 , P2_R1209_U55;
wire P2_R1209_U56 , P2_R1209_U57 , P2_R1209_U58 , P2_R1209_U59 , P2_R1209_U60 , P2_R1209_U61 , P2_R1209_U62 , P2_R1209_U63 , P2_R1209_U64 , P2_R1209_U65;
wire P2_R1209_U66 , P2_R1209_U67 , P2_R1209_U68 , P2_R1209_U69 , P2_R1209_U70 , P2_R1209_U71 , P2_R1209_U72 , P2_R1209_U73 , P2_R1209_U74 , P2_R1209_U75;
wire P2_R1209_U76 , P2_R1209_U77 , P2_R1209_U78 , P2_R1209_U79 , P2_R1209_U80 , P2_R1209_U81 , P2_R1209_U82 , P2_R1209_U83 , P2_R1209_U84 , P2_R1209_U85;
wire P2_R1209_U86 , P2_R1209_U87 , P2_R1209_U88 , P2_R1209_U89 , P2_R1209_U90 , P2_R1209_U91 , P2_R1209_U92 , P2_R1209_U93 , P2_R1209_U94 , P2_R1209_U95;
wire P2_R1209_U96 , P2_R1209_U97 , P2_R1209_U98 , P2_R1209_U99 , P2_R1209_U100 , P2_R1209_U101 , P2_R1209_U102 , P2_R1209_U103 , P2_R1209_U104 , P2_R1209_U105;
wire P2_R1209_U106 , P2_R1209_U107 , P2_R1209_U108 , P2_R1209_U109 , P2_R1209_U110 , P2_R1209_U111 , P2_R1209_U112 , P2_R1209_U113 , P2_R1209_U114 , P2_R1209_U115;
wire P2_R1209_U116 , P2_R1209_U117 , P2_R1209_U118 , P2_R1209_U119 , P2_R1209_U120 , P2_R1209_U121 , P2_R1209_U122 , P2_R1209_U123 , P2_R1209_U124 , P2_R1209_U125;
wire P2_R1209_U126 , P2_R1209_U127 , P2_R1209_U128 , P2_R1209_U129 , P2_R1209_U130 , P2_R1209_U131 , P2_R1209_U132 , P2_R1209_U133 , P2_R1209_U134 , P2_R1209_U135;
wire P2_R1209_U136 , P2_R1209_U137 , P2_R1209_U138 , P2_R1209_U139 , P2_R1209_U140 , P2_R1209_U141 , P2_R1209_U142 , P2_R1209_U143 , P2_R1209_U144 , P2_R1209_U145;
wire P2_R1209_U146 , P2_R1209_U147 , P2_R1209_U148 , P2_R1209_U149 , P2_R1209_U150 , P2_R1209_U151 , P2_R1209_U152 , P2_R1209_U153 , P2_R1209_U154 , P2_R1209_U155;
wire P2_R1209_U156 , P2_R1209_U157 , P2_R1209_U158 , P2_R1209_U159 , P2_R1209_U160 , P2_R1209_U161 , P2_R1209_U162 , P2_R1209_U163 , P2_R1209_U164 , P2_R1209_U165;
wire P2_R1209_U166 , P2_R1209_U167 , P2_R1209_U168 , P2_R1209_U169 , P2_R1209_U170 , P2_R1209_U171 , P2_R1209_U172 , P2_R1209_U173 , P2_R1209_U174 , P2_R1209_U175;
wire P2_R1209_U176 , P2_R1209_U177 , P2_R1209_U178 , P2_R1209_U179 , P2_R1209_U180 , P2_R1209_U181 , P2_R1209_U182 , P2_R1209_U183 , P2_R1209_U184 , P2_R1209_U185;
wire P2_R1209_U186 , P2_R1209_U187 , P2_R1209_U188 , P2_R1209_U189 , P2_R1209_U190 , P2_R1209_U191 , P2_R1209_U192 , P2_R1209_U193 , P2_R1209_U194 , P2_R1209_U195;
wire P2_R1209_U196 , P2_R1209_U197 , P2_R1209_U198 , P2_R1209_U199 , P2_R1209_U200 , P2_R1209_U201 , P2_R1209_U202 , P2_R1209_U203 , P2_R1209_U204 , P2_R1209_U205;
wire P2_R1209_U206 , P2_R1209_U207 , P2_R1209_U208 , P2_R1209_U209 , P2_R1209_U210 , P2_R1209_U211 , P2_R1209_U212 , P2_R1209_U213 , P2_R1209_U214 , P2_R1209_U215;
wire P2_R1209_U216 , P2_R1209_U217 , P2_R1209_U218 , P2_R1209_U219 , P2_R1209_U220 , P2_R1209_U221 , P2_R1209_U222 , P2_R1209_U223 , P2_R1209_U224 , P2_R1209_U225;
wire P2_R1209_U226 , P2_R1209_U227 , P2_R1209_U228 , P2_R1209_U229 , P2_R1209_U230 , P2_R1209_U231 , P2_R1209_U232 , P2_R1209_U233 , P2_R1209_U234 , P2_R1209_U235;
wire P2_R1209_U236 , P2_R1209_U237 , P2_R1209_U238 , P2_R1209_U239 , P2_R1209_U240 , P2_R1209_U241 , P2_R1209_U242 , P2_R1209_U243 , P2_R1209_U244 , P2_R1209_U245;
wire P2_R1209_U246 , P2_R1209_U247 , P2_R1209_U248 , P2_R1209_U249 , P2_R1209_U250 , P2_R1209_U251 , P2_R1209_U252 , P2_R1209_U253 , P2_R1209_U254 , P2_R1209_U255;
wire P2_R1209_U256 , P2_R1209_U257 , P2_R1209_U258 , P2_R1209_U259 , P2_R1209_U260 , P2_R1209_U261 , P2_R1209_U262 , P2_R1209_U263 , P2_R1209_U264 , P2_R1209_U265;
wire P2_R1209_U266 , P2_R1209_U267 , P2_R1209_U268 , P2_R1209_U269 , P2_R1209_U270 , P2_R1209_U271 , P2_R1209_U272 , P2_R1209_U273 , P2_R1209_U274 , P2_R1209_U275;
wire P2_R1209_U276 , P2_R1300_U6 , P2_R1300_U7 , P2_R1300_U8 , P2_R1300_U9 , P2_R1300_U10 , P2_R1200_U6 , P2_R1200_U7 , P2_R1200_U8 , P2_R1200_U9;
wire P2_R1200_U10 , P2_R1200_U11 , P2_R1200_U12 , P2_R1200_U13 , P2_R1200_U14 , P2_R1200_U15 , P2_R1200_U16 , P2_R1200_U17 , P2_R1200_U18 , P2_R1200_U19;
wire P2_R1200_U20 , P2_R1200_U21 , P2_R1200_U22 , P2_R1200_U23 , P2_R1200_U24 , P2_R1200_U25 , P2_R1200_U26 , P2_R1200_U27 , P2_R1200_U28 , P2_R1200_U29;
wire P2_R1200_U30 , P2_R1200_U31 , P2_R1200_U32 , P2_R1200_U33 , P2_R1200_U34 , P2_R1200_U35 , P2_R1200_U36 , P2_R1200_U37 , P2_R1200_U38 , P2_R1200_U39;
wire P2_R1200_U40 , P2_R1200_U41 , P2_R1200_U42 , P2_R1200_U43 , P2_R1200_U44 , P2_R1200_U45 , P2_R1200_U46 , P2_R1200_U47 , P2_R1200_U48 , P2_R1200_U49;
wire P2_R1200_U50 , P2_R1200_U51 , P2_R1200_U52 , P2_R1200_U53 , P2_R1200_U54 , P2_R1200_U55 , P2_R1200_U56 , P2_R1200_U57 , P2_R1200_U58 , P2_R1200_U59;
wire P2_R1200_U60 , P2_R1200_U61 , P2_R1200_U62 , P2_R1200_U63 , P2_R1200_U64 , P2_R1200_U65 , P2_R1200_U66 , P2_R1200_U67 , P2_R1200_U68 , P2_R1200_U69;
wire P2_R1200_U70 , P2_R1200_U71 , P2_R1200_U72 , P2_R1200_U73 , P2_R1200_U74 , P2_R1200_U75 , P2_R1200_U76 , P2_R1200_U77 , P2_R1200_U78 , P2_R1200_U79;
wire P2_R1200_U80 , P2_R1200_U81 , P2_R1200_U82 , P2_R1200_U83 , P2_R1200_U84 , P2_R1200_U85 , P2_R1200_U86 , P2_R1200_U87 , P2_R1200_U88 , P2_R1200_U89;
wire P2_R1200_U90 , P2_R1200_U91 , P2_R1200_U92 , P2_R1200_U93 , P2_R1200_U94 , P2_R1200_U95 , P2_R1200_U96 , P2_R1200_U97 , P2_R1200_U98 , P2_R1200_U99;
wire P2_R1200_U100 , P2_R1200_U101 , P2_R1200_U102 , P2_R1200_U103 , P2_R1200_U104 , P2_R1200_U105 , P2_R1200_U106 , P2_R1200_U107 , P2_R1200_U108 , P2_R1200_U109;
wire P2_R1200_U110 , P2_R1200_U111 , P2_R1200_U112 , P2_R1200_U113 , P2_R1200_U114 , P2_R1200_U115 , P2_R1200_U116 , P2_R1200_U117 , P2_R1200_U118 , P2_R1200_U119;
wire P2_R1200_U120 , P2_R1200_U121 , P2_R1200_U122 , P2_R1200_U123 , P2_R1200_U124 , P2_R1200_U125 , P2_R1200_U126 , P2_R1200_U127 , P2_R1200_U128 , P2_R1200_U129;
wire P2_R1200_U130 , P2_R1200_U131 , P2_R1200_U132 , P2_R1200_U133 , P2_R1200_U134 , P2_R1200_U135 , P2_R1200_U136 , P2_R1200_U137 , P2_R1200_U138 , P2_R1200_U139;
wire P2_R1200_U140 , P2_R1200_U141 , P2_R1200_U142 , P2_R1200_U143 , P2_R1200_U144 , P2_R1200_U145 , P2_R1200_U146 , P2_R1200_U147 , P2_R1200_U148 , P2_R1200_U149;
wire P2_R1200_U150 , P2_R1200_U151 , P2_R1200_U152 , P2_R1200_U153 , P2_R1200_U154 , P2_R1200_U155 , P2_R1200_U156 , P2_R1200_U157 , P2_R1200_U158 , P2_R1200_U159;
wire P2_R1200_U160 , P2_R1200_U161 , P2_R1200_U162 , P2_R1200_U163 , P2_R1200_U164 , P2_R1200_U165 , P2_R1200_U166 , P2_R1200_U167 , P2_R1200_U168 , P2_R1200_U169;
wire P2_R1200_U170 , P2_R1200_U171 , P2_R1200_U172 , P2_R1200_U173 , P2_R1200_U174 , P2_R1200_U175 , P2_R1200_U176 , P2_R1200_U177 , P2_R1200_U178 , P2_R1200_U179;
wire P2_R1200_U180 , P2_R1200_U181 , P2_R1200_U182 , P2_R1200_U183 , P2_R1200_U184 , P2_R1200_U185 , P2_R1200_U186 , P2_R1200_U187 , P2_R1200_U188 , P2_R1200_U189;
wire P2_R1200_U190 , P2_R1200_U191 , P2_R1200_U192 , P2_R1200_U193 , P2_R1200_U194 , P2_R1200_U195 , P2_R1200_U196 , P2_R1200_U197 , P2_R1200_U198 , P2_R1200_U199;
wire P2_R1200_U200 , P2_R1200_U201 , P2_R1200_U202 , P2_R1200_U203 , P2_R1200_U204 , P2_R1200_U205 , P2_R1200_U206 , P2_R1200_U207 , P2_R1200_U208 , P2_R1200_U209;
wire P2_R1200_U210 , P2_R1200_U211 , P2_R1200_U212 , P2_R1200_U213 , P2_R1200_U214 , P2_R1200_U215 , P2_R1200_U216 , P2_R1200_U217 , P2_R1200_U218 , P2_R1200_U219;
wire P2_R1200_U220 , P2_R1200_U221 , P2_R1200_U222 , P2_R1200_U223 , P2_R1200_U224 , P2_R1200_U225 , P2_R1200_U226 , P2_R1200_U227 , P2_R1200_U228 , P2_R1200_U229;
wire P2_R1200_U230 , P2_R1200_U231 , P2_R1200_U232 , P2_R1200_U233 , P2_R1200_U234 , P2_R1200_U235 , P2_R1200_U236 , P2_R1200_U237 , P2_R1200_U238 , P2_R1200_U239;
wire P2_R1200_U240 , P2_R1200_U241 , P2_R1200_U242 , P2_R1200_U243 , P2_R1200_U244 , P2_R1200_U245 , P2_R1200_U246 , P2_R1200_U247 , P2_R1200_U248 , P2_R1200_U249;
wire P2_R1200_U250 , P2_R1200_U251 , P2_R1200_U252 , P2_R1200_U253 , P2_R1200_U254 , P2_R1200_U255 , P2_R1200_U256 , P2_R1200_U257 , P2_R1200_U258 , P2_R1200_U259;
wire P2_R1200_U260 , P2_R1200_U261 , P2_R1200_U262 , P2_R1200_U263 , P2_R1200_U264 , P2_R1200_U265 , P2_R1200_U266 , P2_R1200_U267 , P2_R1200_U268 , P2_R1200_U269;
wire P2_R1200_U270 , P2_R1200_U271 , P2_R1200_U272 , P2_R1200_U273 , P2_R1200_U274 , P2_R1200_U275 , P2_R1200_U276 , P2_R1200_U277 , P2_R1200_U278 , P2_R1200_U279;
wire P2_R1200_U280 , P2_R1200_U281 , P2_R1200_U282 , P2_R1200_U283 , P2_R1200_U284 , P2_R1200_U285 , P2_R1200_U286 , P2_R1200_U287 , P2_R1200_U288 , P2_R1200_U289;
wire P2_R1200_U290 , P2_R1200_U291 , P2_R1200_U292 , P2_R1200_U293 , P2_R1200_U294 , P2_R1200_U295 , P2_R1200_U296 , P2_R1200_U297 , P2_R1200_U298 , P2_R1200_U299;
wire P2_R1200_U300 , P2_R1200_U301 , P2_R1200_U302 , P2_R1200_U303 , P2_R1200_U304 , P2_R1200_U305 , P2_R1200_U306 , P2_R1200_U307 , P2_R1200_U308 , P2_R1200_U309;
wire P2_R1200_U310 , P2_R1200_U311 , P2_R1200_U312 , P2_R1200_U313 , P2_R1200_U314 , P2_R1200_U315 , P2_R1200_U316 , P2_R1200_U317 , P2_R1200_U318 , P2_R1200_U319;
wire P2_R1200_U320 , P2_R1200_U321 , P2_R1200_U322 , P2_R1200_U323 , P2_R1200_U324 , P2_R1200_U325 , P2_R1200_U326 , P2_R1200_U327 , P2_R1200_U328 , P2_R1200_U329;
wire P2_R1200_U330 , P2_R1200_U331 , P2_R1200_U332 , P2_R1200_U333 , P2_R1200_U334 , P2_R1200_U335 , P2_R1200_U336 , P2_R1200_U337 , P2_R1200_U338 , P2_R1200_U339;
wire P2_R1200_U340 , P2_R1200_U341 , P2_R1200_U342 , P2_R1200_U343 , P2_R1200_U344 , P2_R1200_U345 , P2_R1200_U346 , P2_R1200_U347 , P2_R1200_U348 , P2_R1200_U349;
wire P2_R1200_U350 , P2_R1200_U351 , P2_R1200_U352 , P2_R1200_U353 , P2_R1200_U354 , P2_R1200_U355 , P2_R1200_U356 , P2_R1200_U357 , P2_R1200_U358 , P2_R1200_U359;
wire P2_R1200_U360 , P2_R1200_U361 , P2_R1200_U362 , P2_R1200_U363 , P2_R1200_U364 , P2_R1200_U365 , P2_R1200_U366 , P2_R1200_U367 , P2_R1200_U368 , P2_R1200_U369;
wire P2_R1200_U370 , P2_R1200_U371 , P2_R1200_U372 , P2_R1200_U373 , P2_R1200_U374 , P2_R1200_U375 , P2_R1200_U376 , P2_R1200_U377 , P2_R1200_U378 , P2_R1200_U379;
wire P2_R1200_U380 , P2_R1200_U381 , P2_R1200_U382 , P2_R1200_U383 , P2_R1200_U384 , P2_R1200_U385 , P2_R1200_U386 , P2_R1200_U387 , P2_R1200_U388 , P2_R1200_U389;
wire P2_R1200_U390 , P2_R1200_U391 , P2_R1200_U392 , P2_R1200_U393 , P2_R1200_U394 , P2_R1200_U395 , P2_R1200_U396 , P2_R1200_U397 , P2_R1200_U398 , P2_R1200_U399;
wire P2_R1200_U400 , P2_R1200_U401 , P2_R1200_U402 , P2_R1200_U403 , P2_R1200_U404 , P2_R1200_U405 , P2_R1200_U406 , P2_R1200_U407 , P2_R1200_U408 , P2_R1200_U409;
wire P2_R1200_U410 , P2_R1200_U411 , P2_R1200_U412 , P2_R1200_U413 , P2_R1200_U414 , P2_R1200_U415 , P2_R1200_U416 , P2_R1200_U417 , P2_R1200_U418 , P2_R1200_U419;
wire P2_R1200_U420 , P2_R1200_U421 , P2_R1200_U422 , P2_R1200_U423 , P2_R1200_U424 , P2_R1200_U425 , P2_R1200_U426 , P2_R1200_U427 , P2_R1200_U428 , P2_R1200_U429;
wire P2_R1200_U430 , P2_R1200_U431 , P2_R1200_U432 , P2_R1200_U433 , P2_R1200_U434 , P2_R1200_U435 , P2_R1200_U436 , P2_R1200_U437 , P2_R1200_U438 , P2_R1200_U439;
wire P2_R1200_U440 , P2_R1200_U441 , P2_R1200_U442 , P2_R1200_U443 , P2_R1200_U444 , P2_R1200_U445 , P2_R1200_U446 , P2_R1200_U447 , P2_R1200_U448 , P2_R1200_U449;
wire P2_R1200_U450 , P2_R1200_U451 , P2_R1200_U452 , P2_R1200_U453 , P2_R1200_U454 , P2_R1200_U455 , P2_R1200_U456 , P2_R1200_U457 , P2_R1200_U458 , P2_R1200_U459;
wire P2_R1200_U460 , P2_R1200_U461 , P2_R1200_U462 , P2_R1200_U463 , P2_R1200_U464 , P2_R1200_U465 , P2_R1200_U466 , P2_R1200_U467 , P2_R1200_U468 , P2_R1200_U469;
wire P2_R1200_U470 , P2_R1200_U471 , P2_R1200_U472 , P2_R1200_U473 , P2_R1200_U474 , P2_R1200_U475 , P2_R1200_U476 , P2_R1200_U477 , P2_R1200_U478 , P2_R1200_U479;
wire P2_R1200_U480 , P2_R1200_U481 , P2_R1200_U482 , P2_R1200_U483 , P2_R1200_U484 , P2_R1200_U485 , P2_R1200_U486 , P2_R1200_U487 , P2_R1200_U488 , P2_R1200_U489;
wire P2_R1179_U6 , P2_R1179_U7 , P2_R1179_U8 , P2_R1179_U9 , P2_R1179_U10 , P2_R1179_U11 , P2_R1179_U12 , P2_R1179_U13 , P2_R1179_U14 , P2_R1179_U15;
wire P2_R1179_U16 , P2_R1179_U17 , P2_R1179_U18 , P2_R1179_U19 , P2_R1179_U20 , P2_R1179_U21 , P2_R1179_U22 , P2_R1179_U23 , P2_R1179_U24 , P2_R1179_U25;
wire P2_R1179_U26 , P2_R1179_U27 , P2_R1179_U28 , P2_R1179_U29 , P2_R1179_U30 , P2_R1179_U31 , P2_R1179_U32 , P2_R1179_U33 , P2_R1179_U34 , P2_R1179_U35;
wire P2_R1179_U36 , P2_R1179_U37 , P2_R1179_U38 , P2_R1179_U39 , P2_R1179_U40 , P2_R1179_U41 , P2_R1179_U42 , P2_R1179_U43 , P2_R1179_U44 , P2_R1179_U45;
wire P2_R1179_U46 , P2_R1179_U47 , P2_R1179_U48 , P2_R1179_U49 , P2_R1179_U50 , P2_R1179_U51 , P2_R1179_U52 , P2_R1179_U53 , P2_R1179_U54 , P2_R1179_U55;
wire P2_R1179_U56 , P2_R1179_U57 , P2_R1179_U58 , P2_R1179_U59 , P2_R1179_U60 , P2_R1179_U61 , P2_R1179_U62 , P2_R1179_U63 , P2_R1179_U64 , P2_R1179_U65;
wire P2_R1179_U66 , P2_R1179_U67 , P2_R1179_U68 , P2_R1179_U69 , P2_R1179_U70 , P2_R1179_U71 , P2_R1179_U72 , P2_R1179_U73 , P2_R1179_U74 , P2_R1179_U75;
wire P2_R1179_U76 , P2_R1179_U77 , P2_R1179_U78 , P2_R1179_U79 , P2_R1179_U80 , P2_R1179_U81 , P2_R1179_U82 , P2_R1179_U83 , P2_R1179_U84 , P2_R1179_U85;
wire P2_R1179_U86 , P2_R1179_U87 , P2_R1179_U88 , P2_R1179_U89 , P2_R1179_U90 , P2_R1179_U91 , P2_R1179_U92 , P2_R1179_U93 , P2_R1179_U94 , P2_R1179_U95;
wire P2_R1179_U96 , P2_R1179_U97 , P2_R1179_U98 , P2_R1179_U99 , P2_R1179_U100 , P2_R1179_U101 , P2_R1179_U102 , P2_R1179_U103 , P2_R1179_U104 , P2_R1179_U105;
wire P2_R1179_U106 , P2_R1179_U107 , P2_R1179_U108 , P2_R1179_U109 , P2_R1179_U110 , P2_R1179_U111 , P2_R1179_U112 , P2_R1179_U113 , P2_R1179_U114 , P2_R1179_U115;
wire P2_R1179_U116 , P2_R1179_U117 , P2_R1179_U118 , P2_R1179_U119 , P2_R1179_U120 , P2_R1179_U121 , P2_R1179_U122 , P2_R1179_U123 , P2_R1179_U124 , P2_R1179_U125;
wire P2_R1179_U126 , P2_R1179_U127 , P2_R1179_U128 , P2_R1179_U129 , P2_R1179_U130 , P2_R1179_U131 , P2_R1179_U132 , P2_R1179_U133 , P2_R1179_U134 , P2_R1179_U135;
wire P2_R1179_U136 , P2_R1179_U137 , P2_R1179_U138 , P2_R1179_U139 , P2_R1179_U140 , P2_R1179_U141 , P2_R1179_U142 , P2_R1179_U143 , P2_R1179_U144 , P2_R1179_U145;
wire P2_R1179_U146 , P2_R1179_U147 , P2_R1179_U148 , P2_R1179_U149 , P2_R1179_U150 , P2_R1179_U151 , P2_R1179_U152 , P2_R1179_U153 , P2_R1179_U154 , P2_R1179_U155;
wire P2_R1179_U156 , P2_R1179_U157 , P2_R1179_U158 , P2_R1179_U159 , P2_R1179_U160 , P2_R1179_U161 , P2_R1179_U162 , P2_R1179_U163 , P2_R1179_U164 , P2_R1179_U165;
wire P2_R1179_U166 , P2_R1179_U167 , P2_R1179_U168 , P2_R1179_U169 , P2_R1179_U170 , P2_R1179_U171 , P2_R1179_U172 , P2_R1179_U173 , P2_R1179_U174 , P2_R1179_U175;
wire P2_R1179_U176 , P2_R1179_U177 , P2_R1179_U178 , P2_R1179_U179 , P2_R1179_U180 , P2_R1179_U181 , P2_R1179_U182 , P2_R1179_U183 , P2_R1179_U184 , P2_R1179_U185;
wire P2_R1179_U186 , P2_R1179_U187 , P2_R1179_U188 , P2_R1179_U189 , P2_R1179_U190 , P2_R1179_U191 , P2_R1179_U192 , P2_R1179_U193 , P2_R1179_U194 , P2_R1179_U195;
wire P2_R1179_U196 , P2_R1179_U197 , P2_R1179_U198 , P2_R1179_U199 , P2_R1179_U200 , P2_R1179_U201 , P2_R1179_U202 , P2_R1179_U203 , P2_R1179_U204 , P2_R1179_U205;
wire P2_R1179_U206 , P2_R1179_U207 , P2_R1179_U208 , P2_R1179_U209 , P2_R1179_U210 , P2_R1179_U211 , P2_R1179_U212 , P2_R1179_U213 , P2_R1179_U214 , P2_R1179_U215;
wire P2_R1179_U216 , P2_R1179_U217 , P2_R1179_U218 , P2_R1179_U219 , P2_R1179_U220 , P2_R1179_U221 , P2_R1179_U222 , P2_R1179_U223 , P2_R1179_U224 , P2_R1179_U225;
wire P2_R1179_U226 , P2_R1179_U227 , P2_R1179_U228 , P2_R1179_U229 , P2_R1179_U230 , P2_R1179_U231 , P2_R1179_U232 , P2_R1179_U233 , P2_R1179_U234 , P2_R1179_U235;
wire P2_R1179_U236 , P2_R1179_U237 , P2_R1179_U238 , P2_R1179_U239 , P2_R1179_U240 , P2_R1179_U241 , P2_R1179_U242 , P2_R1179_U243 , P2_R1179_U244 , P2_R1179_U245;
wire P2_R1179_U246 , P2_R1179_U247 , P2_R1179_U248 , P2_R1179_U249 , P2_R1179_U250 , P2_R1179_U251 , P2_R1179_U252 , P2_R1179_U253 , P2_R1179_U254 , P2_R1179_U255;
wire P2_R1179_U256 , P2_R1179_U257 , P2_R1179_U258 , P2_R1179_U259 , P2_R1179_U260 , P2_R1179_U261 , P2_R1179_U262 , P2_R1179_U263 , P2_R1179_U264 , P2_R1179_U265;
wire P2_R1179_U266 , P2_R1179_U267 , P2_R1179_U268 , P2_R1179_U269 , P2_R1179_U270 , P2_R1179_U271 , P2_R1179_U272 , P2_R1179_U273 , P2_R1179_U274 , P2_R1179_U275;
wire P2_R1179_U276 , P2_R1179_U277 , P2_R1179_U278 , P2_R1179_U279 , P2_R1179_U280 , P2_R1179_U281 , P2_R1179_U282 , P2_R1179_U283 , P2_R1179_U284 , P2_R1179_U285;
wire P2_R1179_U286 , P2_R1179_U287 , P2_R1179_U288 , P2_R1179_U289 , P2_R1179_U290 , P2_R1179_U291 , P2_R1179_U292 , P2_R1179_U293 , P2_R1179_U294 , P2_R1179_U295;
wire P2_R1179_U296 , P2_R1179_U297 , P2_R1179_U298 , P2_R1179_U299 , P2_R1179_U300 , P2_R1179_U301 , P2_R1179_U302 , P2_R1179_U303 , P2_R1179_U304 , P2_R1179_U305;
wire P2_R1179_U306 , P2_R1179_U307 , P2_R1179_U308 , P2_R1179_U309 , P2_R1179_U310 , P2_R1179_U311 , P2_R1179_U312 , P2_R1179_U313 , P2_R1179_U314 , P2_R1179_U315;
wire P2_R1179_U316 , P2_R1179_U317 , P2_R1179_U318 , P2_R1179_U319 , P2_R1179_U320 , P2_R1179_U321 , P2_R1179_U322 , P2_R1179_U323 , P2_R1179_U324 , P2_R1179_U325;
wire P2_R1179_U326 , P2_R1179_U327 , P2_R1179_U328 , P2_R1179_U329 , P2_R1179_U330 , P2_R1179_U331 , P2_R1179_U332 , P2_R1179_U333 , P2_R1179_U334 , P2_R1179_U335;
wire P2_R1179_U336 , P2_R1179_U337 , P2_R1179_U338 , P2_R1179_U339 , P2_R1179_U340 , P2_R1179_U341 , P2_R1179_U342 , P2_R1179_U343 , P2_R1179_U344 , P2_R1179_U345;
wire P2_R1179_U346 , P2_R1179_U347 , P2_R1179_U348 , P2_R1179_U349 , P2_R1179_U350 , P2_R1179_U351 , P2_R1179_U352 , P2_R1179_U353 , P2_R1179_U354 , P2_R1179_U355;
wire P2_R1179_U356 , P2_R1179_U357 , P2_R1179_U358 , P2_R1179_U359 , P2_R1179_U360 , P2_R1179_U361 , P2_R1179_U362 , P2_R1179_U363 , P2_R1179_U364 , P2_R1179_U365;
wire P2_R1179_U366 , P2_R1179_U367 , P2_R1179_U368 , P2_R1179_U369 , P2_R1179_U370 , P2_R1179_U371 , P2_R1179_U372 , P2_R1179_U373 , P2_R1179_U374 , P2_R1179_U375;
wire P2_R1179_U376 , P2_R1179_U377 , P2_R1179_U378 , P2_R1179_U379 , P2_R1179_U380 , P2_R1179_U381 , P2_R1179_U382 , P2_R1179_U383 , P2_R1179_U384 , P2_R1179_U385;
wire P2_R1179_U386 , P2_R1179_U387 , P2_R1179_U388 , P2_R1179_U389 , P2_R1179_U390 , P2_R1179_U391 , P2_R1179_U392 , P2_R1179_U393 , P2_R1179_U394 , P2_R1179_U395;
wire P2_R1179_U396 , P2_R1179_U397 , P2_R1179_U398 , P2_R1179_U399 , P2_R1179_U400 , P2_R1179_U401 , P2_R1179_U402 , P2_R1179_U403 , P2_R1179_U404 , P2_R1179_U405;
wire P2_R1179_U406 , P2_R1179_U407 , P2_R1179_U408 , P2_R1179_U409 , P2_R1179_U410 , P2_R1179_U411 , P2_R1179_U412 , P2_R1179_U413 , P2_R1179_U414 , P2_R1179_U415;
wire P2_R1179_U416 , P2_R1179_U417 , P2_R1179_U418 , P2_R1179_U419 , P2_R1179_U420 , P2_R1179_U421 , P2_R1179_U422 , P2_R1179_U423 , P2_R1179_U424 , P2_R1179_U425;
wire P2_R1179_U426 , P2_R1179_U427 , P2_R1179_U428 , P2_R1179_U429 , P2_R1179_U430 , P2_R1179_U431 , P2_R1179_U432 , P2_R1179_U433 , P2_R1179_U434 , P2_R1179_U435;
wire P2_R1179_U436 , P2_R1179_U437 , P2_R1179_U438 , P2_R1179_U439 , P2_R1179_U440 , P2_R1179_U441 , P2_R1179_U442 , P2_R1179_U443 , P2_R1179_U444 , P2_R1179_U445;
wire P2_R1179_U446 , P2_R1179_U447 , P2_R1179_U448 , P2_R1179_U449 , P2_R1179_U450 , P2_R1179_U451 , P2_R1179_U452 , P2_R1179_U453 , P2_R1179_U454 , P2_R1179_U455;
wire P2_R1179_U456 , P2_R1179_U457 , P2_R1179_U458 , P2_R1179_U459 , P2_R1179_U460 , P2_R1179_U461 , P2_R1179_U462 , P2_R1179_U463 , P2_R1179_U464 , P2_R1179_U465;
wire P2_R1179_U466 , P2_R1179_U467 , P2_R1179_U468 , P2_R1179_U469 , P2_R1179_U470 , P2_R1179_U471 , P2_R1179_U472 , P2_R1179_U473 , P2_R1179_U474 , P2_R1179_U475;
wire P2_R1179_U476 , P2_R1179_U477 , P2_R1179_U478 , P2_R1179_U479 , P2_R1179_U480 , P2_R1179_U481 , P2_R1179_U482 , P2_R1179_U483 , P2_R1179_U484 , P2_R1179_U485;
wire P2_R1179_U486 , P2_R1179_U487 , P2_R1179_U488 , P2_R1179_U489 , P2_R1269_U6 , P2_R1269_U7 , P2_R1269_U8 , P2_R1269_U9 , P2_R1269_U10 , P2_R1269_U11;
wire P2_R1269_U12 , P2_R1269_U13 , P2_R1269_U14 , P2_R1269_U15 , P2_R1269_U16 , P2_R1269_U17 , P2_R1269_U18 , P2_R1269_U19 , P2_R1269_U20 , P2_R1269_U21;
wire P2_R1269_U22 , P2_R1269_U23 , P2_R1269_U24 , P2_R1269_U25 , P2_R1269_U26 , P2_R1269_U27 , P2_R1269_U28 , P2_R1269_U29 , P2_R1269_U30 , P2_R1269_U31;
wire P2_R1269_U32 , P2_R1269_U33 , P2_R1269_U34 , P2_R1269_U35 , P2_R1269_U36 , P2_R1269_U37 , P2_R1269_U38 , P2_R1269_U39 , P2_R1269_U40 , P2_R1269_U41;
wire P2_R1269_U42 , P2_R1269_U43 , P2_R1269_U44 , P2_R1269_U45 , P2_R1269_U46 , P2_R1269_U47 , P2_R1269_U48 , P2_R1269_U49 , P2_R1269_U50 , P2_R1269_U51;
wire P2_R1269_U52 , P2_R1269_U53 , P2_R1269_U54 , P2_R1269_U55 , P2_R1269_U56 , P2_R1269_U57 , P2_R1269_U58 , P2_R1269_U59 , P2_R1269_U60 , P2_R1269_U61;
wire P2_R1269_U62 , P2_R1269_U63 , P2_R1269_U64 , P2_R1269_U65 , P2_R1269_U66 , P2_R1269_U67 , P2_R1269_U68 , P2_R1269_U69 , P2_R1269_U70 , P2_R1269_U71;
wire P2_R1269_U72 , P2_R1269_U73 , P2_R1269_U74 , P2_R1269_U75 , P2_R1269_U76 , P2_R1269_U77 , P2_R1269_U78 , P2_R1269_U79 , P2_R1269_U80 , P2_R1269_U81;
wire P2_R1269_U82 , P2_R1269_U83 , P2_R1269_U84 , P2_R1269_U85 , P2_R1269_U86 , P2_R1269_U87 , P2_R1269_U88 , P2_R1269_U89 , P2_R1269_U90 , P2_R1269_U91;
wire P2_R1269_U92 , P2_R1269_U93 , P2_R1269_U94 , P2_R1269_U95 , P2_R1269_U96 , P2_R1269_U97 , P2_R1269_U98 , P2_R1269_U99 , P2_R1269_U100 , P2_R1269_U101;
wire P2_R1269_U102 , P2_R1269_U103 , P2_R1269_U104 , P2_R1269_U105 , P2_R1269_U106 , P2_R1269_U107 , P2_R1269_U108 , P2_R1269_U109 , P2_R1269_U110 , P2_R1269_U111;
wire P2_R1269_U112 , P2_R1269_U113 , P2_R1269_U114 , P2_R1269_U115 , P2_R1269_U116 , P2_R1269_U117 , P2_R1269_U118 , P2_R1269_U119 , P2_R1269_U120 , P2_R1269_U121;
wire P2_R1269_U122 , P2_R1269_U123 , P2_R1269_U124 , P2_R1269_U125 , P2_R1269_U126 , P2_R1269_U127 , P2_R1269_U128 , P2_R1269_U129 , P2_R1269_U130 , P2_R1269_U131;
wire P2_R1269_U132 , P2_R1269_U133 , P2_R1269_U134 , P2_R1269_U135 , P2_R1269_U136 , P2_R1269_U137 , P2_R1269_U138 , P2_R1269_U139 , P2_R1269_U140 , P2_R1269_U141;
wire P2_R1269_U142 , P2_R1269_U143 , P2_R1269_U144 , P2_R1269_U145 , P2_R1269_U146 , P2_R1269_U147 , P2_R1269_U148 , P2_R1269_U149 , P2_R1269_U150 , P2_R1269_U151;
wire P2_R1269_U152 , P2_R1269_U153 , P2_R1269_U154 , P2_R1269_U155 , P2_R1269_U156 , P2_R1269_U157 , P2_R1269_U158 , P2_R1269_U159 , P2_R1269_U160 , P2_R1269_U161;
wire P2_R1269_U162 , P2_R1269_U163 , P2_R1269_U164 , P2_R1269_U165 , P2_R1269_U166 , P2_R1269_U167 , P2_R1269_U168 , P2_R1269_U169 , P2_R1269_U170 , P2_R1269_U171;
wire P2_R1269_U172 , P2_R1269_U173 , P2_R1269_U174 , P2_R1269_U175 , P2_R1269_U176 , P2_R1269_U177 , P2_R1269_U178 , P2_R1269_U179 , P2_R1269_U180 , P2_R1269_U181;
wire P2_R1269_U182 , P2_R1269_U183 , P2_R1269_U184 , P2_R1269_U185 , P2_R1269_U186 , P2_R1269_U187 , P2_R1269_U188 , P2_R1269_U189 , P2_R1269_U190 , P2_R1269_U191;
wire P2_R1269_U192 , P2_R1269_U193 , P2_R1269_U194 , P2_R1269_U195 , P2_R1269_U196 , P2_R1269_U197 , P2_R1269_U198 , P2_R1269_U199 , P2_R1269_U200 , P2_R1269_U201;
wire P2_R1269_U202 , P2_R1269_U203 , P2_R1269_U204 , P2_R1269_U205 , P2_R1269_U206 , P2_R1269_U207 , P2_R1269_U208 , P2_R1269_U209 , P2_R1110_U4 , P2_R1110_U5;
wire P2_R1110_U6 , P2_R1110_U7 , P2_R1110_U8 , P2_R1110_U9 , P2_R1110_U10 , P2_R1110_U11 , P2_R1110_U12 , P2_R1110_U13 , P2_R1110_U14 , P2_R1110_U15;
wire P2_R1110_U16 , P2_R1110_U17 , P2_R1110_U18 , P2_R1110_U19 , P2_R1110_U20 , P2_R1110_U21 , P2_R1110_U22 , P2_R1110_U23 , P2_R1110_U24 , P2_R1110_U25;
wire P2_R1110_U26 , P2_R1110_U27 , P2_R1110_U28 , P2_R1110_U29 , P2_R1110_U30 , P2_R1110_U31 , P2_R1110_U32 , P2_R1110_U33 , P2_R1110_U34 , P2_R1110_U35;
wire P2_R1110_U36 , P2_R1110_U37 , P2_R1110_U38 , P2_R1110_U39 , P2_R1110_U40 , P2_R1110_U41 , P2_R1110_U42 , P2_R1110_U43 , P2_R1110_U44 , P2_R1110_U45;
wire P2_R1110_U46 , P2_R1110_U47 , P2_R1110_U48 , P2_R1110_U49 , P2_R1110_U50 , P2_R1110_U51 , P2_R1110_U52 , P2_R1110_U53 , P2_R1110_U54 , P2_R1110_U55;
wire P2_R1110_U56 , P2_R1110_U57 , P2_R1110_U58 , P2_R1110_U59 , P2_R1110_U60 , P2_R1110_U61 , P2_R1110_U62 , P2_R1110_U63 , P2_R1110_U64 , P2_R1110_U65;
wire P2_R1110_U66 , P2_R1110_U67 , P2_R1110_U68 , P2_R1110_U69 , P2_R1110_U70 , P2_R1110_U71 , P2_R1110_U72 , P2_R1110_U73 , P2_R1110_U74 , P2_R1110_U75;
wire P2_R1110_U76 , P2_R1110_U77 , P2_R1110_U78 , P2_R1110_U79 , P2_R1110_U80 , P2_R1110_U81 , P2_R1110_U82 , P2_R1110_U83 , P2_R1110_U84 , P2_R1110_U85;
wire P2_R1110_U86 , P2_R1110_U87 , P2_R1110_U88 , P2_R1110_U89 , P2_R1110_U90 , P2_R1110_U91 , P2_R1110_U92 , P2_R1110_U93 , P2_R1110_U94 , P2_R1110_U95;
wire P2_R1110_U96 , P2_R1110_U97 , P2_R1110_U98 , P2_R1110_U99 , P2_R1110_U100 , P2_R1110_U101 , P2_R1110_U102 , P2_R1110_U103 , P2_R1110_U104 , P2_R1110_U105;
wire P2_R1110_U106 , P2_R1110_U107 , P2_R1110_U108 , P2_R1110_U109 , P2_R1110_U110 , P2_R1110_U111 , P2_R1110_U112 , P2_R1110_U113 , P2_R1110_U114 , P2_R1110_U115;
wire P2_R1110_U116 , P2_R1110_U117 , P2_R1110_U118 , P2_R1110_U119 , P2_R1110_U120 , P2_R1110_U121 , P2_R1110_U122 , P2_R1110_U123 , P2_R1110_U124 , P2_R1110_U125;
wire P2_R1110_U126 , P2_R1110_U127 , P2_R1110_U128 , P2_R1110_U129 , P2_R1110_U130 , P2_R1110_U131 , P2_R1110_U132 , P2_R1110_U133 , P2_R1110_U134 , P2_R1110_U135;
wire P2_R1110_U136 , P2_R1110_U137 , P2_R1110_U138 , P2_R1110_U139 , P2_R1110_U140 , P2_R1110_U141 , P2_R1110_U142 , P2_R1110_U143 , P2_R1110_U144 , P2_R1110_U145;
wire P2_R1110_U146 , P2_R1110_U147 , P2_R1110_U148 , P2_R1110_U149 , P2_R1110_U150 , P2_R1110_U151 , P2_R1110_U152 , P2_R1110_U153 , P2_R1110_U154 , P2_R1110_U155;
wire P2_R1110_U156 , P2_R1110_U157 , P2_R1110_U158 , P2_R1110_U159 , P2_R1110_U160 , P2_R1110_U161 , P2_R1110_U162 , P2_R1110_U163 , P2_R1110_U164 , P2_R1110_U165;
wire P2_R1110_U166 , P2_R1110_U167 , P2_R1110_U168 , P2_R1110_U169 , P2_R1110_U170 , P2_R1110_U171 , P2_R1110_U172 , P2_R1110_U173 , P2_R1110_U174 , P2_R1110_U175;
wire P2_R1110_U176 , P2_R1110_U177 , P2_R1110_U178 , P2_R1110_U179 , P2_R1110_U180 , P2_R1110_U181 , P2_R1110_U182 , P2_R1110_U183 , P2_R1110_U184 , P2_R1110_U185;
wire P2_R1110_U186 , P2_R1110_U187 , P2_R1110_U188 , P2_R1110_U189 , P2_R1110_U190 , P2_R1110_U191 , P2_R1110_U192 , P2_R1110_U193 , P2_R1110_U194 , P2_R1110_U195;
wire P2_R1110_U196 , P2_R1110_U197 , P2_R1110_U198 , P2_R1110_U199 , P2_R1110_U200 , P2_R1110_U201 , P2_R1110_U202 , P2_R1110_U203 , P2_R1110_U204 , P2_R1110_U205;
wire P2_R1110_U206 , P2_R1110_U207 , P2_R1110_U208 , P2_R1110_U209 , P2_R1110_U210 , P2_R1110_U211 , P2_R1110_U212 , P2_R1110_U213 , P2_R1110_U214 , P2_R1110_U215;
wire P2_R1110_U216 , P2_R1110_U217 , P2_R1110_U218 , P2_R1110_U219 , P2_R1110_U220 , P2_R1110_U221 , P2_R1110_U222 , P2_R1110_U223 , P2_R1110_U224 , P2_R1110_U225;
wire P2_R1110_U226 , P2_R1110_U227 , P2_R1110_U228 , P2_R1110_U229 , P2_R1110_U230 , P2_R1110_U231 , P2_R1110_U232 , P2_R1110_U233 , P2_R1110_U234 , P2_R1110_U235;
wire P2_R1110_U236 , P2_R1110_U237 , P2_R1110_U238 , P2_R1110_U239 , P2_R1110_U240 , P2_R1110_U241 , P2_R1110_U242 , P2_R1110_U243 , P2_R1110_U244 , P2_R1110_U245;
wire P2_R1110_U246 , P2_R1110_U247 , P2_R1110_U248 , P2_R1110_U249 , P2_R1110_U250 , P2_R1110_U251 , P2_R1110_U252 , P2_R1110_U253 , P2_R1110_U254 , P2_R1110_U255;
wire P2_R1110_U256 , P2_R1110_U257 , P2_R1110_U258 , P2_R1110_U259 , P2_R1110_U260 , P2_R1110_U261 , P2_R1110_U262 , P2_R1110_U263 , P2_R1110_U264 , P2_R1110_U265;
wire P2_R1110_U266 , P2_R1110_U267 , P2_R1110_U268 , P2_R1110_U269 , P2_R1110_U270 , P2_R1110_U271 , P2_R1110_U272 , P2_R1110_U273 , P2_R1110_U274 , P2_R1110_U275;
wire P2_R1110_U276 , P2_R1110_U277 , P2_R1110_U278 , P2_R1110_U279 , P2_R1110_U280 , P2_R1110_U281 , P2_R1110_U282 , P2_R1110_U283 , P2_R1110_U284 , P2_R1110_U285;
wire P2_R1110_U286 , P2_R1110_U287 , P2_R1110_U288 , P2_R1110_U289 , P2_R1110_U290 , P2_R1110_U291 , P2_R1110_U292 , P2_R1110_U293 , P2_R1110_U294 , P2_R1110_U295;
wire P2_R1110_U296 , P2_R1110_U297 , P2_R1110_U298 , P2_R1110_U299 , P2_R1110_U300 , P2_R1110_U301 , P2_R1110_U302 , P2_R1110_U303 , P2_R1110_U304 , P2_R1110_U305;
wire P2_R1110_U306 , P2_R1110_U307 , P2_R1110_U308 , P2_R1110_U309 , P2_R1110_U310 , P2_R1110_U311 , P2_R1110_U312 , P2_R1110_U313 , P2_R1110_U314 , P2_R1110_U315;
wire P2_R1110_U316 , P2_R1110_U317 , P2_R1110_U318 , P2_R1110_U319 , P2_R1110_U320 , P2_R1110_U321 , P2_R1110_U322 , P2_R1110_U323 , P2_R1110_U324 , P2_R1110_U325;
wire P2_R1110_U326 , P2_R1110_U327 , P2_R1110_U328 , P2_R1110_U329 , P2_R1110_U330 , P2_R1110_U331 , P2_R1110_U332 , P2_R1110_U333 , P2_R1110_U334 , P2_R1110_U335;
wire P2_R1110_U336 , P2_R1110_U337 , P2_R1110_U338 , P2_R1110_U339 , P2_R1110_U340 , P2_R1110_U341 , P2_R1110_U342 , P2_R1110_U343 , P2_R1110_U344 , P2_R1110_U345;
wire P2_R1110_U346 , P2_R1110_U347 , P2_R1110_U348 , P2_R1110_U349 , P2_R1110_U350 , P2_R1110_U351 , P2_R1110_U352 , P2_R1110_U353 , P2_R1110_U354 , P2_R1110_U355;
wire P2_R1110_U356 , P2_R1110_U357 , P2_R1110_U358 , P2_R1110_U359 , P2_R1110_U360 , P2_R1110_U361 , P2_R1110_U362 , P2_R1110_U363 , P2_R1110_U364 , P2_R1110_U365;
wire P2_R1110_U366 , P2_R1110_U367 , P2_R1110_U368 , P2_R1110_U369 , P2_R1110_U370 , P2_R1110_U371 , P2_R1110_U372 , P2_R1110_U373 , P2_R1110_U374 , P2_R1110_U375;
wire P2_R1110_U376 , P2_R1110_U377 , P2_R1110_U378 , P2_R1110_U379 , P2_R1110_U380 , P2_R1110_U381 , P2_R1110_U382 , P2_R1110_U383 , P2_R1110_U384 , P2_R1110_U385;
wire P2_R1110_U386 , P2_R1110_U387 , P2_R1110_U388 , P2_R1110_U389 , P2_R1110_U390 , P2_R1110_U391 , P2_R1110_U392 , P2_R1110_U393 , P2_R1110_U394 , P2_R1110_U395;
wire P2_R1110_U396 , P2_R1110_U397 , P2_R1110_U398 , P2_R1110_U399 , P2_R1110_U400 , P2_R1110_U401 , P2_R1110_U402 , P2_R1110_U403 , P2_R1110_U404 , P2_R1110_U405;
wire P2_R1110_U406 , P2_R1110_U407 , P2_R1110_U408 , P2_R1110_U409 , P2_R1110_U410 , P2_R1110_U411 , P2_R1110_U412 , P2_R1110_U413 , P2_R1110_U414 , P2_R1110_U415;
wire P2_R1110_U416 , P2_R1110_U417 , P2_R1110_U418 , P2_R1110_U419 , P2_R1110_U420 , P2_R1110_U421 , P2_R1110_U422 , P2_R1110_U423 , P2_R1110_U424 , P2_R1110_U425;
wire P2_R1110_U426 , P2_R1110_U427 , P2_R1110_U428 , P2_R1110_U429 , P2_R1110_U430 , P2_R1110_U431 , P2_R1110_U432 , P2_R1110_U433 , P2_R1110_U434 , P2_R1110_U435;
wire P2_R1110_U436 , P2_R1110_U437 , P2_R1110_U438 , P2_R1110_U439 , P2_R1110_U440 , P2_R1110_U441 , P2_R1110_U442 , P2_R1110_U443 , P2_R1110_U444 , P2_R1110_U445;
wire P2_R1110_U446 , P2_R1110_U447 , P2_R1110_U448 , P2_R1110_U449 , P2_R1110_U450 , P2_R1110_U451 , P2_R1110_U452 , P2_R1110_U453 , P2_R1110_U454 , P2_R1110_U455;
wire P2_R1110_U456 , P2_R1110_U457 , P2_R1110_U458 , P2_R1110_U459 , P2_R1110_U460 , P2_R1110_U461 , P2_R1110_U462 , P2_R1110_U463 , P2_R1110_U464 , P2_R1110_U465;
wire P2_R1110_U466 , P2_R1110_U467 , P2_R1110_U468 , P2_R1110_U469 , P2_R1110_U470 , P2_R1110_U471 , P2_R1110_U472 , P2_R1110_U473 , P2_R1110_U474 , P2_R1110_U475;
wire P2_R1110_U476 , P2_R1110_U477 , P2_R1110_U478 , P2_R1110_U479 , P2_R1110_U480 , P2_R1110_U481 , P2_R1110_U482 , P2_R1110_U483 , P2_R1110_U484 , P2_R1110_U485;
wire P2_R1110_U486 , P2_R1110_U487 , P2_R1110_U488 , P2_R1110_U489 , P2_R1110_U490 , P2_R1110_U491 , P2_R1110_U492 , P2_R1110_U493 , P2_R1110_U494 , P2_R1110_U495;
wire P2_R1110_U496 , P2_R1110_U497 , P2_R1110_U498 , P2_R1110_U499 , P2_R1110_U500 , P2_R1110_U501 , P2_R1110_U502 , P2_R1110_U503 , P2_R1110_U504 , P2_R1297_U6;
wire P2_R1297_U7 , P2_R1077_U4 , P2_R1077_U5 , P2_R1077_U6 , P2_R1077_U7 , P2_R1077_U8 , P2_R1077_U9 , P2_R1077_U10 , P2_R1077_U11 , P2_R1077_U12;
wire P2_R1077_U13 , P2_R1077_U14 , P2_R1077_U15 , P2_R1077_U16 , P2_R1077_U17 , P2_R1077_U18 , P2_R1077_U19 , P2_R1077_U20 , P2_R1077_U21 , P2_R1077_U22;
wire P2_R1077_U23 , P2_R1077_U24 , P2_R1077_U25 , P2_R1077_U26 , P2_R1077_U27 , P2_R1077_U28 , P2_R1077_U29 , P2_R1077_U30 , P2_R1077_U31 , P2_R1077_U32;
wire P2_R1077_U33 , P2_R1077_U34 , P2_R1077_U35 , P2_R1077_U36 , P2_R1077_U37 , P2_R1077_U38 , P2_R1077_U39 , P2_R1077_U40 , P2_R1077_U41 , P2_R1077_U42;
wire P2_R1077_U43 , P2_R1077_U44 , P2_R1077_U45 , P2_R1077_U46 , P2_R1077_U47 , P2_R1077_U48 , P2_R1077_U49 , P2_R1077_U50 , P2_R1077_U51 , P2_R1077_U52;
wire P2_R1077_U53 , P2_R1077_U54 , P2_R1077_U55 , P2_R1077_U56 , P2_R1077_U57 , P2_R1077_U58 , P2_R1077_U59 , P2_R1077_U60 , P2_R1077_U61 , P2_R1077_U62;
wire P2_R1077_U63 , P2_R1077_U64 , P2_R1077_U65 , P2_R1077_U66 , P2_R1077_U67 , P2_R1077_U68 , P2_R1077_U69 , P2_R1077_U70 , P2_R1077_U71 , P2_R1077_U72;
wire P2_R1077_U73 , P2_R1077_U74 , P2_R1077_U75 , P2_R1077_U76 , P2_R1077_U77 , P2_R1077_U78 , P2_R1077_U79 , P2_R1077_U80 , P2_R1077_U81 , P2_R1077_U82;
wire P2_R1077_U83 , P2_R1077_U84 , P2_R1077_U85 , P2_R1077_U86 , P2_R1077_U87 , P2_R1077_U88 , P2_R1077_U89 , P2_R1077_U90 , P2_R1077_U91 , P2_R1077_U92;
wire P2_R1077_U93 , P2_R1077_U94 , P2_R1077_U95 , P2_R1077_U96 , P2_R1077_U97 , P2_R1077_U98 , P2_R1077_U99 , P2_R1077_U100 , P2_R1077_U101 , P2_R1077_U102;
wire P2_R1077_U103 , P2_R1077_U104 , P2_R1077_U105 , P2_R1077_U106 , P2_R1077_U107 , P2_R1077_U108 , P2_R1077_U109 , P2_R1077_U110 , P2_R1077_U111 , P2_R1077_U112;
wire P2_R1077_U113 , P2_R1077_U114 , P2_R1077_U115 , P2_R1077_U116 , P2_R1077_U117 , P2_R1077_U118 , P2_R1077_U119 , P2_R1077_U120 , P2_R1077_U121 , P2_R1077_U122;
wire P2_R1077_U123 , P2_R1077_U124 , P2_R1077_U125 , P2_R1077_U126 , P2_R1077_U127 , P2_R1077_U128 , P2_R1077_U129 , P2_R1077_U130 , P2_R1077_U131 , P2_R1077_U132;
wire P2_R1077_U133 , P2_R1077_U134 , P2_R1077_U135 , P2_R1077_U136 , P2_R1077_U137 , P2_R1077_U138 , P2_R1077_U139 , P2_R1077_U140 , P2_R1077_U141 , P2_R1077_U142;
wire P2_R1077_U143 , P2_R1077_U144 , P2_R1077_U145 , P2_R1077_U146 , P2_R1077_U147 , P2_R1077_U148 , P2_R1077_U149 , P2_R1077_U150 , P2_R1077_U151 , P2_R1077_U152;
wire P2_R1077_U153 , P2_R1077_U154 , P2_R1077_U155 , P2_R1077_U156 , P2_R1077_U157 , P2_R1077_U158 , P2_R1077_U159 , P2_R1077_U160 , P2_R1077_U161 , P2_R1077_U162;
wire P2_R1077_U163 , P2_R1077_U164 , P2_R1077_U165 , P2_R1077_U166 , P2_R1077_U167 , P2_R1077_U168 , P2_R1077_U169 , P2_R1077_U170 , P2_R1077_U171 , P2_R1077_U172;
wire P2_R1077_U173 , P2_R1077_U174 , P2_R1077_U175 , P2_R1077_U176 , P2_R1077_U177 , P2_R1077_U178 , P2_R1077_U179 , P2_R1077_U180 , P2_R1077_U181 , P2_R1077_U182;
wire P2_R1077_U183 , P2_R1077_U184 , P2_R1077_U185 , P2_R1077_U186 , P2_R1077_U187 , P2_R1077_U188 , P2_R1077_U189 , P2_R1077_U190 , P2_R1077_U191 , P2_R1077_U192;
wire P2_R1077_U193 , P2_R1077_U194 , P2_R1077_U195 , P2_R1077_U196 , P2_R1077_U197 , P2_R1077_U198 , P2_R1077_U199 , P2_R1077_U200 , P2_R1077_U201 , P2_R1077_U202;
wire P2_R1077_U203 , P2_R1077_U204 , P2_R1077_U205 , P2_R1077_U206 , P2_R1077_U207 , P2_R1077_U208 , P2_R1077_U209 , P2_R1077_U210 , P2_R1077_U211 , P2_R1077_U212;
wire P2_R1077_U213 , P2_R1077_U214 , P2_R1077_U215 , P2_R1077_U216 , P2_R1077_U217 , P2_R1077_U218 , P2_R1077_U219 , P2_R1077_U220 , P2_R1077_U221 , P2_R1077_U222;
wire P2_R1077_U223 , P2_R1077_U224 , P2_R1077_U225 , P2_R1077_U226 , P2_R1077_U227 , P2_R1077_U228 , P2_R1077_U229 , P2_R1077_U230 , P2_R1077_U231 , P2_R1077_U232;
wire P2_R1077_U233 , P2_R1077_U234 , P2_R1077_U235 , P2_R1077_U236 , P2_R1077_U237 , P2_R1077_U238 , P2_R1077_U239 , P2_R1077_U240 , P2_R1077_U241 , P2_R1077_U242;
wire P2_R1077_U243 , P2_R1077_U244 , P2_R1077_U245 , P2_R1077_U246 , P2_R1077_U247 , P2_R1077_U248 , P2_R1077_U249 , P2_R1077_U250 , P2_R1077_U251 , P2_R1077_U252;
wire P2_R1077_U253 , P2_R1077_U254 , P2_R1077_U255 , P2_R1077_U256 , P2_R1077_U257 , P2_R1077_U258 , P2_R1077_U259 , P2_R1077_U260 , P2_R1077_U261 , P2_R1077_U262;
wire P2_R1077_U263 , P2_R1077_U264 , P2_R1077_U265 , P2_R1077_U266 , P2_R1077_U267 , P2_R1077_U268 , P2_R1077_U269 , P2_R1077_U270 , P2_R1077_U271 , P2_R1077_U272;
wire P2_R1077_U273 , P2_R1077_U274 , P2_R1077_U275 , P2_R1077_U276 , P2_R1077_U277 , P2_R1077_U278 , P2_R1077_U279 , P2_R1077_U280 , P2_R1077_U281 , P2_R1077_U282;
wire P2_R1077_U283 , P2_R1077_U284 , P2_R1077_U285 , P2_R1077_U286 , P2_R1077_U287 , P2_R1077_U288 , P2_R1077_U289 , P2_R1077_U290 , P2_R1077_U291 , P2_R1077_U292;
wire P2_R1077_U293 , P2_R1077_U294 , P2_R1077_U295 , P2_R1077_U296 , P2_R1077_U297 , P2_R1077_U298 , P2_R1077_U299 , P2_R1077_U300 , P2_R1077_U301 , P2_R1077_U302;
wire P2_R1077_U303 , P2_R1077_U304 , P2_R1077_U305 , P2_R1077_U306 , P2_R1077_U307 , P2_R1077_U308 , P2_R1077_U309 , P2_R1077_U310 , P2_R1077_U311 , P2_R1077_U312;
wire P2_R1077_U313 , P2_R1077_U314 , P2_R1077_U315 , P2_R1077_U316 , P2_R1077_U317 , P2_R1077_U318 , P2_R1077_U319 , P2_R1077_U320 , P2_R1077_U321 , P2_R1077_U322;
wire P2_R1077_U323 , P2_R1077_U324 , P2_R1077_U325 , P2_R1077_U326 , P2_R1077_U327 , P2_R1077_U328 , P2_R1077_U329 , P2_R1077_U330 , P2_R1077_U331 , P2_R1077_U332;
wire P2_R1077_U333 , P2_R1077_U334 , P2_R1077_U335 , P2_R1077_U336 , P2_R1077_U337 , P2_R1077_U338 , P2_R1077_U339 , P2_R1077_U340 , P2_R1077_U341 , P2_R1077_U342;
wire P2_R1077_U343 , P2_R1077_U344 , P2_R1077_U345 , P2_R1077_U346 , P2_R1077_U347 , P2_R1077_U348 , P2_R1077_U349 , P2_R1077_U350 , P2_R1077_U351 , P2_R1077_U352;
wire P2_R1077_U353 , P2_R1077_U354 , P2_R1077_U355 , P2_R1077_U356 , P2_R1077_U357 , P2_R1077_U358 , P2_R1077_U359 , P2_R1077_U360 , P2_R1077_U361 , P2_R1077_U362;
wire P2_R1077_U363 , P2_R1077_U364 , P2_R1077_U365 , P2_R1077_U366 , P2_R1077_U367 , P2_R1077_U368 , P2_R1077_U369 , P2_R1077_U370 , P2_R1077_U371 , P2_R1077_U372;
wire P2_R1077_U373 , P2_R1077_U374 , P2_R1077_U375 , P2_R1077_U376 , P2_R1077_U377 , P2_R1077_U378 , P2_R1077_U379 , P2_R1077_U380 , P2_R1077_U381 , P2_R1077_U382;
wire P2_R1077_U383 , P2_R1077_U384 , P2_R1077_U385 , P2_R1077_U386 , P2_R1077_U387 , P2_R1077_U388 , P2_R1077_U389 , P2_R1077_U390 , P2_R1077_U391 , P2_R1077_U392;
wire P2_R1077_U393 , P2_R1077_U394 , P2_R1077_U395 , P2_R1077_U396 , P2_R1077_U397 , P2_R1077_U398 , P2_R1077_U399 , P2_R1077_U400 , P2_R1077_U401 , P2_R1077_U402;
wire P2_R1077_U403 , P2_R1077_U404 , P2_R1077_U405 , P2_R1077_U406 , P2_R1077_U407 , P2_R1077_U408 , P2_R1077_U409 , P2_R1077_U410 , P2_R1077_U411 , P2_R1077_U412;
wire P2_R1077_U413 , P2_R1077_U414 , P2_R1077_U415 , P2_R1077_U416 , P2_R1077_U417 , P2_R1077_U418 , P2_R1077_U419 , P2_R1077_U420 , P2_R1077_U421 , P2_R1077_U422;
wire P2_R1077_U423 , P2_R1077_U424 , P2_R1077_U425 , P2_R1077_U426 , P2_R1077_U427 , P2_R1077_U428 , P2_R1077_U429 , P2_R1077_U430 , P2_R1077_U431 , P2_R1077_U432;
wire P2_R1077_U433 , P2_R1077_U434 , P2_R1077_U435 , P2_R1077_U436 , P2_R1077_U437 , P2_R1077_U438 , P2_R1077_U439 , P2_R1077_U440 , P2_R1077_U441 , P2_R1077_U442;
wire P2_R1077_U443 , P2_R1077_U444 , P2_R1077_U445 , P2_R1077_U446 , P2_R1077_U447 , P2_R1077_U448 , P2_R1077_U449 , P2_R1077_U450 , P2_R1077_U451 , P2_R1077_U452;
wire P2_R1077_U453 , P2_R1077_U454 , P2_R1077_U455 , P2_R1077_U456 , P2_R1077_U457 , P2_R1077_U458 , P2_R1077_U459 , P2_R1077_U460 , P2_R1077_U461 , P2_R1077_U462;
wire P2_R1077_U463 , P2_R1077_U464 , P2_R1077_U465 , P2_R1077_U466 , P2_R1077_U467 , P2_R1077_U468 , P2_R1077_U469 , P2_R1077_U470 , P2_R1077_U471 , P2_R1077_U472;
wire P2_R1077_U473 , P2_R1077_U474 , P2_R1077_U475 , P2_R1077_U476 , P2_R1077_U477 , P2_R1077_U478 , P2_R1077_U479 , P2_R1077_U480 , P2_R1077_U481 , P2_R1077_U482;
wire P2_R1077_U483 , P2_R1077_U484 , P2_R1077_U485 , P2_R1077_U486 , P2_R1077_U487 , P2_R1077_U488 , P2_R1077_U489 , P2_R1077_U490 , P2_R1077_U491 , P2_R1077_U492;
wire P2_R1077_U493 , P2_R1077_U494 , P2_R1077_U495 , P2_R1077_U496 , P2_R1077_U497 , P2_R1077_U498 , P2_R1077_U499 , P2_R1077_U500 , P2_R1077_U501 , P2_R1077_U502;
wire P2_R1077_U503 , P2_R1077_U504 , P2_R1143_U4 , P2_R1143_U5 , P2_R1143_U6 , P2_R1143_U7 , P2_R1143_U8 , P2_R1143_U9 , P2_R1143_U10 , P2_R1143_U11;
wire P2_R1143_U12 , P2_R1143_U13 , P2_R1143_U14 , P2_R1143_U15 , P2_R1143_U16 , P2_R1143_U17 , P2_R1143_U18 , P2_R1143_U19 , P2_R1143_U20 , P2_R1143_U21;
wire P2_R1143_U22 , P2_R1143_U23 , P2_R1143_U24 , P2_R1143_U25 , P2_R1143_U26 , P2_R1143_U27 , P2_R1143_U28 , P2_R1143_U29 , P2_R1143_U30 , P2_R1143_U31;
wire P2_R1143_U32 , P2_R1143_U33 , P2_R1143_U34 , P2_R1143_U35 , P2_R1143_U36 , P2_R1143_U37 , P2_R1143_U38 , P2_R1143_U39 , P2_R1143_U40 , P2_R1143_U41;
wire P2_R1143_U42 , P2_R1143_U43 , P2_R1143_U44 , P2_R1143_U45 , P2_R1143_U46 , P2_R1143_U47 , P2_R1143_U48 , P2_R1143_U49 , P2_R1143_U50 , P2_R1143_U51;
wire P2_R1143_U52 , P2_R1143_U53 , P2_R1143_U54 , P2_R1143_U55 , P2_R1143_U56 , P2_R1143_U57 , P2_R1143_U58 , P2_R1143_U59 , P2_R1143_U60 , P2_R1143_U61;
wire P2_R1143_U62 , P2_R1143_U63 , P2_R1143_U64 , P2_R1143_U65 , P2_R1143_U66 , P2_R1143_U67 , P2_R1143_U68 , P2_R1143_U69 , P2_R1143_U70 , P2_R1143_U71;
wire P2_R1143_U72 , P2_R1143_U73 , P2_R1143_U74 , P2_R1143_U75 , P2_R1143_U76 , P2_R1143_U77 , P2_R1143_U78 , P2_R1143_U79 , P2_R1143_U80 , P2_R1143_U81;
wire P2_R1143_U82 , P2_R1143_U83 , P2_R1143_U84 , P2_R1143_U85 , P2_R1143_U86 , P2_R1143_U87 , P2_R1143_U88 , P2_R1143_U89 , P2_R1143_U90 , P2_R1143_U91;
wire P2_R1143_U92 , P2_R1143_U93 , P2_R1143_U94 , P2_R1143_U95 , P2_R1143_U96 , P2_R1143_U97 , P2_R1143_U98 , P2_R1143_U99 , P2_R1143_U100 , P2_R1143_U101;
wire P2_R1143_U102 , P2_R1143_U103 , P2_R1143_U104 , P2_R1143_U105 , P2_R1143_U106 , P2_R1143_U107 , P2_R1143_U108 , P2_R1143_U109 , P2_R1143_U110 , P2_R1143_U111;
wire P2_R1143_U112 , P2_R1143_U113 , P2_R1143_U114 , P2_R1143_U115 , P2_R1143_U116 , P2_R1143_U117 , P2_R1143_U118 , P2_R1143_U119 , P2_R1143_U120 , P2_R1143_U121;
wire P2_R1143_U122 , P2_R1143_U123 , P2_R1143_U124 , P2_R1143_U125 , P2_R1143_U126 , P2_R1143_U127 , P2_R1143_U128 , P2_R1143_U129 , P2_R1143_U130 , P2_R1143_U131;
wire P2_R1143_U132 , P2_R1143_U133 , P2_R1143_U134 , P2_R1143_U135 , P2_R1143_U136 , P2_R1143_U137 , P2_R1143_U138 , P2_R1143_U139 , P2_R1143_U140 , P2_R1143_U141;
wire P2_R1143_U142 , P2_R1143_U143 , P2_R1143_U144 , P2_R1143_U145 , P2_R1143_U146 , P2_R1143_U147 , P2_R1143_U148 , P2_R1143_U149 , P2_R1143_U150 , P2_R1143_U151;
wire P2_R1143_U152 , P2_R1143_U153 , P2_R1143_U154 , P2_R1143_U155 , P2_R1143_U156 , P2_R1143_U157 , P2_R1143_U158 , P2_R1143_U159 , P2_R1143_U160 , P2_R1143_U161;
wire P2_R1143_U162 , P2_R1143_U163 , P2_R1143_U164 , P2_R1143_U165 , P2_R1143_U166 , P2_R1143_U167 , P2_R1143_U168 , P2_R1143_U169 , P2_R1143_U170 , P2_R1143_U171;
wire P2_R1143_U172 , P2_R1143_U173 , P2_R1143_U174 , P2_R1143_U175 , P2_R1143_U176 , P2_R1143_U177 , P2_R1143_U178 , P2_R1143_U179 , P2_R1143_U180 , P2_R1143_U181;
wire P2_R1143_U182 , P2_R1143_U183 , P2_R1143_U184 , P2_R1143_U185 , P2_R1143_U186 , P2_R1143_U187 , P2_R1143_U188 , P2_R1143_U189 , P2_R1143_U190 , P2_R1143_U191;
wire P2_R1143_U192 , P2_R1143_U193 , P2_R1143_U194 , P2_R1143_U195 , P2_R1143_U196 , P2_R1143_U197 , P2_R1143_U198 , P2_R1143_U199 , P2_R1143_U200 , P2_R1143_U201;
wire P2_R1143_U202 , P2_R1143_U203 , P2_R1143_U204 , P2_R1143_U205 , P2_R1143_U206 , P2_R1143_U207 , P2_R1143_U208 , P2_R1143_U209 , P2_R1143_U210 , P2_R1143_U211;
wire P2_R1143_U212 , P2_R1143_U213 , P2_R1143_U214 , P2_R1143_U215 , P2_R1143_U216 , P2_R1143_U217 , P2_R1143_U218 , P2_R1143_U219 , P2_R1143_U220 , P2_R1143_U221;
wire P2_R1143_U222 , P2_R1143_U223 , P2_R1143_U224 , P2_R1143_U225 , P2_R1143_U226 , P2_R1143_U227 , P2_R1143_U228 , P2_R1143_U229 , P2_R1143_U230 , P2_R1143_U231;
wire P2_R1143_U232 , P2_R1143_U233 , P2_R1143_U234 , P2_R1143_U235 , P2_R1143_U236 , P2_R1143_U237 , P2_R1143_U238 , P2_R1143_U239 , P2_R1143_U240 , P2_R1143_U241;
wire P2_R1143_U242 , P2_R1143_U243 , P2_R1143_U244 , P2_R1143_U245 , P2_R1143_U246 , P2_R1143_U247 , P2_R1143_U248 , P2_R1143_U249 , P2_R1143_U250 , P2_R1143_U251;
wire P2_R1143_U252 , P2_R1143_U253 , P2_R1143_U254 , P2_R1143_U255 , P2_R1143_U256 , P2_R1143_U257 , P2_R1143_U258 , P2_R1143_U259 , P2_R1143_U260 , P2_R1143_U261;
wire P2_R1143_U262 , P2_R1143_U263 , P2_R1143_U264 , P2_R1143_U265 , P2_R1143_U266 , P2_R1143_U267 , P2_R1143_U268 , P2_R1143_U269 , P2_R1143_U270 , P2_R1143_U271;
wire P2_R1143_U272 , P2_R1143_U273 , P2_R1143_U274 , P2_R1143_U275 , P2_R1143_U276 , P2_R1143_U277 , P2_R1143_U278 , P2_R1143_U279 , P2_R1143_U280 , P2_R1143_U281;
wire P2_R1143_U282 , P2_R1143_U283 , P2_R1143_U284 , P2_R1143_U285 , P2_R1143_U286 , P2_R1143_U287 , P2_R1143_U288 , P2_R1143_U289 , P2_R1143_U290 , P2_R1143_U291;
wire P2_R1143_U292 , P2_R1143_U293 , P2_R1143_U294 , P2_R1143_U295 , P2_R1143_U296 , P2_R1143_U297 , P2_R1143_U298 , P2_R1143_U299 , P2_R1143_U300 , P2_R1143_U301;
wire P2_R1143_U302 , P2_R1143_U303 , P2_R1143_U304 , P2_R1143_U305 , P2_R1143_U306 , P2_R1143_U307 , P2_R1143_U308 , P2_R1143_U309 , P2_R1143_U310 , P2_R1143_U311;
wire P2_R1143_U312 , P2_R1143_U313 , P2_R1143_U314 , P2_R1143_U315 , P2_R1143_U316 , P2_R1143_U317 , P2_R1143_U318 , P2_R1143_U319 , P2_R1143_U320 , P2_R1143_U321;
wire P2_R1143_U322 , P2_R1143_U323 , P2_R1143_U324 , P2_R1143_U325 , P2_R1143_U326 , P2_R1143_U327 , P2_R1143_U328 , P2_R1143_U329 , P2_R1143_U330 , P2_R1143_U331;
wire P2_R1143_U332 , P2_R1143_U333 , P2_R1143_U334 , P2_R1143_U335 , P2_R1143_U336 , P2_R1143_U337 , P2_R1143_U338 , P2_R1143_U339 , P2_R1143_U340 , P2_R1143_U341;
wire P2_R1143_U342 , P2_R1143_U343 , P2_R1143_U344 , P2_R1143_U345 , P2_R1143_U346 , P2_R1143_U347 , P2_R1143_U348 , P2_R1143_U349 , P2_R1143_U350 , P2_R1143_U351;
wire P2_R1143_U352 , P2_R1143_U353 , P2_R1143_U354 , P2_R1143_U355 , P2_R1143_U356 , P2_R1143_U357 , P2_R1143_U358 , P2_R1143_U359 , P2_R1143_U360 , P2_R1143_U361;
wire P2_R1143_U362 , P2_R1143_U363 , P2_R1143_U364 , P2_R1143_U365 , P2_R1143_U366 , P2_R1143_U367 , P2_R1143_U368 , P2_R1143_U369 , P2_R1143_U370 , P2_R1143_U371;
wire P2_R1143_U372 , P2_R1143_U373 , P2_R1143_U374 , P2_R1143_U375 , P2_R1143_U376 , P2_R1143_U377 , P2_R1143_U378 , P2_R1143_U379 , P2_R1143_U380 , P2_R1143_U381;
wire P2_R1143_U382 , P2_R1143_U383 , P2_R1143_U384 , P2_R1143_U385 , P2_R1143_U386 , P2_R1143_U387 , P2_R1143_U388 , P2_R1143_U389 , P2_R1143_U390 , P2_R1143_U391;
wire P2_R1143_U392 , P2_R1143_U393 , P2_R1143_U394 , P2_R1143_U395 , P2_R1143_U396 , P2_R1143_U397 , P2_R1143_U398 , P2_R1143_U399 , P2_R1143_U400 , P2_R1143_U401;
wire P2_R1143_U402 , P2_R1143_U403 , P2_R1143_U404 , P2_R1143_U405 , P2_R1143_U406 , P2_R1143_U407 , P2_R1143_U408 , P2_R1143_U409 , P2_R1143_U410 , P2_R1143_U411;
wire P2_R1143_U412 , P2_R1143_U413 , P2_R1143_U414 , P2_R1143_U415 , P2_R1143_U416 , P2_R1143_U417 , P2_R1143_U418 , P2_R1143_U419 , P2_R1143_U420 , P2_R1143_U421;
wire P2_R1143_U422 , P2_R1143_U423 , P2_R1143_U424 , P2_R1143_U425 , P2_R1143_U426 , P2_R1143_U427 , P2_R1143_U428 , P2_R1143_U429 , P2_R1143_U430 , P2_R1143_U431;
wire P2_R1143_U432 , P2_R1143_U433 , P2_R1143_U434 , P2_R1143_U435 , P2_R1143_U436 , P2_R1143_U437 , P2_R1143_U438 , P2_R1143_U439 , P2_R1143_U440 , P2_R1143_U441;
wire P2_R1143_U442 , P2_R1143_U443 , P2_R1143_U444 , P2_R1143_U445 , P2_R1143_U446 , P2_R1143_U447 , P2_R1143_U448 , P2_R1143_U449 , P2_R1143_U450 , P2_R1143_U451;
wire P2_R1143_U452 , P2_R1143_U453 , P2_R1143_U454 , P2_R1143_U455 , P2_R1143_U456 , P2_R1143_U457 , P2_R1143_U458 , P2_R1143_U459 , P2_R1143_U460 , P2_R1143_U461;
wire P2_R1143_U462 , P2_R1143_U463 , P2_R1143_U464 , P2_R1143_U465 , P2_R1143_U466 , P2_R1143_U467 , P2_R1143_U468 , P2_R1143_U469 , P2_R1143_U470 , P2_R1143_U471;
wire P2_R1143_U472 , P2_R1143_U473 , P2_R1143_U474 , P2_R1143_U475 , P2_R1143_U476 , P2_R1143_U477 , P2_R1143_U478 , P2_R1143_U479 , P2_R1143_U480 , P2_R1143_U481;
wire P2_R1143_U482 , P2_R1143_U483 , P2_R1143_U484 , P2_R1143_U485 , P2_R1143_U486 , P2_R1143_U487 , P2_R1143_U488 , P2_R1143_U489 , P2_R1143_U490 , P2_R1143_U491;
wire P2_R1143_U492 , P2_R1143_U493 , P2_R1143_U494 , P2_R1143_U495 , P2_R1143_U496 , P2_R1143_U497 , P2_R1143_U498 , P2_R1143_U499 , P2_R1143_U500 , P2_R1143_U501;
wire P2_R1143_U502 , P2_R1143_U503 , P2_R1143_U504 , P2_R1158_U4 , P2_R1158_U5 , P2_R1158_U6 , P2_R1158_U7 , P2_R1158_U8 , P2_R1158_U9 , P2_R1158_U10;
wire P2_R1158_U11 , P2_R1158_U12 , P2_R1158_U13 , P2_R1158_U14 , P2_R1158_U15 , P2_R1158_U16 , P2_R1158_U17 , P2_R1158_U18 , P2_R1158_U19 , P2_R1158_U20;
wire P2_R1158_U21 , P2_R1158_U22 , P2_R1158_U23 , P2_R1158_U24 , P2_R1158_U25 , P2_R1158_U26 , P2_R1158_U27 , P2_R1158_U28 , P2_R1158_U29 , P2_R1158_U30;
wire P2_R1158_U31 , P2_R1158_U32 , P2_R1158_U33 , P2_R1158_U34 , P2_R1158_U35 , P2_R1158_U36 , P2_R1158_U37 , P2_R1158_U38 , P2_R1158_U39 , P2_R1158_U40;
wire P2_R1158_U41 , P2_R1158_U42 , P2_R1158_U43 , P2_R1158_U44 , P2_R1158_U45 , P2_R1158_U46 , P2_R1158_U47 , P2_R1158_U48 , P2_R1158_U49 , P2_R1158_U50;
wire P2_R1158_U51 , P2_R1158_U52 , P2_R1158_U53 , P2_R1158_U54 , P2_R1158_U55 , P2_R1158_U56 , P2_R1158_U57 , P2_R1158_U58 , P2_R1158_U59 , P2_R1158_U60;
wire P2_R1158_U61 , P2_R1158_U62 , P2_R1158_U63 , P2_R1158_U64 , P2_R1158_U65 , P2_R1158_U66 , P2_R1158_U67 , P2_R1158_U68 , P2_R1158_U69 , P2_R1158_U70;
wire P2_R1158_U71 , P2_R1158_U72 , P2_R1158_U73 , P2_R1158_U74 , P2_R1158_U75 , P2_R1158_U76 , P2_R1158_U77 , P2_R1158_U78 , P2_R1158_U79 , P2_R1158_U80;
wire P2_R1158_U81 , P2_R1158_U82 , P2_R1158_U83 , P2_R1158_U84 , P2_R1158_U85 , P2_R1158_U86 , P2_R1158_U87 , P2_R1158_U88 , P2_R1158_U89 , P2_R1158_U90;
wire P2_R1158_U91 , P2_R1158_U92 , P2_R1158_U93 , P2_R1158_U94 , P2_R1158_U95 , P2_R1158_U96 , P2_R1158_U97 , P2_R1158_U98 , P2_R1158_U99 , P2_R1158_U100;
wire P2_R1158_U101 , P2_R1158_U102 , P2_R1158_U103 , P2_R1158_U104 , P2_R1158_U105 , P2_R1158_U106 , P2_R1158_U107 , P2_R1158_U108 , P2_R1158_U109 , P2_R1158_U110;
wire P2_R1158_U111 , P2_R1158_U112 , P2_R1158_U113 , P2_R1158_U114 , P2_R1158_U115 , P2_R1158_U116 , P2_R1158_U117 , P2_R1158_U118 , P2_R1158_U119 , P2_R1158_U120;
wire P2_R1158_U121 , P2_R1158_U122 , P2_R1158_U123 , P2_R1158_U124 , P2_R1158_U125 , P2_R1158_U126 , P2_R1158_U127 , P2_R1158_U128 , P2_R1158_U129 , P2_R1158_U130;
wire P2_R1158_U131 , P2_R1158_U132 , P2_R1158_U133 , P2_R1158_U134 , P2_R1158_U135 , P2_R1158_U136 , P2_R1158_U137 , P2_R1158_U138 , P2_R1158_U139 , P2_R1158_U140;
wire P2_R1158_U141 , P2_R1158_U142 , P2_R1158_U143 , P2_R1158_U144 , P2_R1158_U145 , P2_R1158_U146 , P2_R1158_U147 , P2_R1158_U148 , P2_R1158_U149 , P2_R1158_U150;
wire P2_R1158_U151 , P2_R1158_U152 , P2_R1158_U153 , P2_R1158_U154 , P2_R1158_U155 , P2_R1158_U156 , P2_R1158_U157 , P2_R1158_U158 , P2_R1158_U159 , P2_R1158_U160;
wire P2_R1158_U161 , P2_R1158_U162 , P2_R1158_U163 , P2_R1158_U164 , P2_R1158_U165 , P2_R1158_U166 , P2_R1158_U167 , P2_R1158_U168 , P2_R1158_U169 , P2_R1158_U170;
wire P2_R1158_U171 , P2_R1158_U172 , P2_R1158_U173 , P2_R1158_U174 , P2_R1158_U175 , P2_R1158_U176 , P2_R1158_U177 , P2_R1158_U178 , P2_R1158_U179 , P2_R1158_U180;
wire P2_R1158_U181 , P2_R1158_U182 , P2_R1158_U183 , P2_R1158_U184 , P2_R1158_U185 , P2_R1158_U186 , P2_R1158_U187 , P2_R1158_U188 , P2_R1158_U189 , P2_R1158_U190;
wire P2_R1158_U191 , P2_R1158_U192 , P2_R1158_U193 , P2_R1158_U194 , P2_R1158_U195 , P2_R1158_U196 , P2_R1158_U197 , P2_R1158_U198 , P2_R1158_U199 , P2_R1158_U200;
wire P2_R1158_U201 , P2_R1158_U202 , P2_R1158_U203 , P2_R1158_U204 , P2_R1158_U205 , P2_R1158_U206 , P2_R1158_U207 , P2_R1158_U208 , P2_R1158_U209 , P2_R1158_U210;
wire P2_R1158_U211 , P2_R1158_U212 , P2_R1158_U213 , P2_R1158_U214 , P2_R1158_U215 , P2_R1158_U216 , P2_R1158_U217 , P2_R1158_U218 , P2_R1158_U219 , P2_R1158_U220;
wire P2_R1158_U221 , P2_R1158_U222 , P2_R1158_U223 , P2_R1158_U224 , P2_R1158_U225 , P2_R1158_U226 , P2_R1158_U227 , P2_R1158_U228 , P2_R1158_U229 , P2_R1158_U230;
wire P2_R1158_U231 , P2_R1158_U232 , P2_R1158_U233 , P2_R1158_U234 , P2_R1158_U235 , P2_R1158_U236 , P2_R1158_U237 , P2_R1158_U238 , P2_R1158_U239 , P2_R1158_U240;
wire P2_R1158_U241 , P2_R1158_U242 , P2_R1158_U243 , P2_R1158_U244 , P2_R1158_U245 , P2_R1158_U246 , P2_R1158_U247 , P2_R1158_U248 , P2_R1158_U249 , P2_R1158_U250;
wire P2_R1158_U251 , P2_R1158_U252 , P2_R1158_U253 , P2_R1158_U254 , P2_R1158_U255 , P2_R1158_U256 , P2_R1158_U257 , P2_R1158_U258 , P2_R1158_U259 , P2_R1158_U260;
wire P2_R1158_U261 , P2_R1158_U262 , P2_R1158_U263 , P2_R1158_U264 , P2_R1158_U265 , P2_R1158_U266 , P2_R1158_U267 , P2_R1158_U268 , P2_R1158_U269 , P2_R1158_U270;
wire P2_R1158_U271 , P2_R1158_U272 , P2_R1158_U273 , P2_R1158_U274 , P2_R1158_U275 , P2_R1158_U276 , P2_R1158_U277 , P2_R1158_U278 , P2_R1158_U279 , P2_R1158_U280;
wire P2_R1158_U281 , P2_R1158_U282 , P2_R1158_U283 , P2_R1158_U284 , P2_R1158_U285 , P2_R1158_U286 , P2_R1158_U287 , P2_R1158_U288 , P2_R1158_U289 , P2_R1158_U290;
wire P2_R1158_U291 , P2_R1158_U292 , P2_R1158_U293 , P2_R1158_U294 , P2_R1158_U295 , P2_R1158_U296 , P2_R1158_U297 , P2_R1158_U298 , P2_R1158_U299 , P2_R1158_U300;
wire P2_R1158_U301 , P2_R1158_U302 , P2_R1158_U303 , P2_R1158_U304 , P2_R1158_U305 , P2_R1158_U306 , P2_R1158_U307 , P2_R1158_U308 , P2_R1158_U309 , P2_R1158_U310;
wire P2_R1158_U311 , P2_R1158_U312 , P2_R1158_U313 , P2_R1158_U314 , P2_R1158_U315 , P2_R1158_U316 , P2_R1158_U317 , P2_R1158_U318 , P2_R1158_U319 , P2_R1158_U320;
wire P2_R1158_U321 , P2_R1158_U322 , P2_R1158_U323 , P2_R1158_U324 , P2_R1158_U325 , P2_R1158_U326 , P2_R1158_U327 , P2_R1158_U328 , P2_R1158_U329 , P2_R1158_U330;
wire P2_R1158_U331 , P2_R1158_U332 , P2_R1158_U333 , P2_R1158_U334 , P2_R1158_U335 , P2_R1158_U336 , P2_R1158_U337 , P2_R1158_U338 , P2_R1158_U339 , P2_R1158_U340;
wire P2_R1158_U341 , P2_R1158_U342 , P2_R1158_U343 , P2_R1158_U344 , P2_R1158_U345 , P2_R1158_U346 , P2_R1158_U347 , P2_R1158_U348 , P2_R1158_U349 , P2_R1158_U350;
wire P2_R1158_U351 , P2_R1158_U352 , P2_R1158_U353 , P2_R1158_U354 , P2_R1158_U355 , P2_R1158_U356 , P2_R1158_U357 , P2_R1158_U358 , P2_R1158_U359 , P2_R1158_U360;
wire P2_R1158_U361 , P2_R1158_U362 , P2_R1158_U363 , P2_R1158_U364 , P2_R1158_U365 , P2_R1158_U366 , P2_R1158_U367 , P2_R1158_U368 , P2_R1158_U369 , P2_R1158_U370;
wire P2_R1158_U371 , P2_R1158_U372 , P2_R1158_U373 , P2_R1158_U374 , P2_R1158_U375 , P2_R1158_U376 , P2_R1158_U377 , P2_R1158_U378 , P2_R1158_U379 , P2_R1158_U380;
wire P2_R1158_U381 , P2_R1158_U382 , P2_R1158_U383 , P2_R1158_U384 , P2_R1158_U385 , P2_R1158_U386 , P2_R1158_U387 , P2_R1158_U388 , P2_R1158_U389 , P2_R1158_U390;
wire P2_R1158_U391 , P2_R1158_U392 , P2_R1158_U393 , P2_R1158_U394 , P2_R1158_U395 , P2_R1158_U396 , P2_R1158_U397 , P2_R1158_U398 , P2_R1158_U399 , P2_R1158_U400;
wire P2_R1158_U401 , P2_R1158_U402 , P2_R1158_U403 , P2_R1158_U404 , P2_R1158_U405 , P2_R1158_U406 , P2_R1158_U407 , P2_R1158_U408 , P2_R1158_U409 , P2_R1158_U410;
wire P2_R1158_U411 , P2_R1158_U412 , P2_R1158_U413 , P2_R1158_U414 , P2_R1158_U415 , P2_R1158_U416 , P2_R1158_U417 , P2_R1158_U418 , P2_R1158_U419 , P2_R1158_U420;
wire P2_R1158_U421 , P2_R1158_U422 , P2_R1158_U423 , P2_R1158_U424 , P2_R1158_U425 , P2_R1158_U426 , P2_R1158_U427 , P2_R1158_U428 , P2_R1158_U429 , P2_R1158_U430;
wire P2_R1158_U431 , P2_R1158_U432 , P2_R1158_U433 , P2_R1158_U434 , P2_R1158_U435 , P2_R1158_U436 , P2_R1158_U437 , P2_R1158_U438 , P2_R1158_U439 , P2_R1158_U440;
wire P2_R1158_U441 , P2_R1158_U442 , P2_R1158_U443 , P2_R1158_U444 , P2_R1158_U445 , P2_R1158_U446 , P2_R1158_U447 , P2_R1158_U448 , P2_R1158_U449 , P2_R1158_U450;
wire P2_R1158_U451 , P2_R1158_U452 , P2_R1158_U453 , P2_R1158_U454 , P2_R1158_U455 , P2_R1158_U456 , P2_R1158_U457 , P2_R1158_U458 , P2_R1158_U459 , P2_R1158_U460;
wire P2_R1158_U461 , P2_R1158_U462 , P2_R1158_U463 , P2_R1158_U464 , P2_R1158_U465 , P2_R1158_U466 , P2_R1158_U467 , P2_R1158_U468 , P2_R1158_U469 , P2_R1158_U470;
wire P2_R1158_U471 , P2_R1158_U472 , P2_R1158_U473 , P2_R1158_U474 , P2_R1158_U475 , P2_R1158_U476 , P2_R1158_U477 , P2_R1158_U478 , P2_R1158_U479 , P2_R1158_U480;
wire P2_R1158_U481 , P2_R1158_U482 , P2_R1158_U483 , P2_R1158_U484 , P2_R1158_U485 , P2_R1158_U486 , P2_R1158_U487 , P2_R1158_U488 , P2_R1158_U489 , P2_R1158_U490;
wire P2_R1158_U491 , P2_R1158_U492 , P2_R1158_U493 , P2_R1158_U494 , P2_R1158_U495 , P2_R1158_U496 , P2_R1158_U497 , P2_R1158_U498 , P2_R1158_U499 , P2_R1158_U500;
wire P2_R1158_U501 , P2_R1158_U502 , P2_R1158_U503 , P2_R1158_U504 , P2_R1158_U505 , P2_R1158_U506 , P2_R1158_U507 , P2_R1158_U508 , P2_R1158_U509 , P2_R1158_U510;
wire P2_R1158_U511 , P2_R1158_U512 , P2_R1158_U513 , P2_R1158_U514 , P2_R1158_U515 , P2_R1158_U516 , P2_R1158_U517 , P2_R1158_U518 , P2_R1158_U519 , P2_R1158_U520;
wire P2_R1158_U521 , P2_R1158_U522 , P2_R1158_U523 , P2_R1158_U524 , P2_R1158_U525 , P2_R1158_U526 , P2_R1158_U527 , P2_R1158_U528 , P2_R1158_U529 , P2_R1158_U530;
wire P2_R1158_U531 , P2_R1158_U532 , P2_R1158_U533 , P2_R1158_U534 , P2_R1158_U535 , P2_R1158_U536 , P2_R1158_U537 , P2_R1158_U538 , P2_R1158_U539 , P2_R1158_U540;
wire P2_R1158_U541 , P2_R1158_U542 , P2_R1158_U543 , P2_R1158_U544 , P2_R1158_U545 , P2_R1158_U546 , P2_R1158_U547 , P2_R1158_U548 , P2_R1158_U549 , P2_R1158_U550;
wire P2_R1158_U551 , P2_R1158_U552 , P2_R1158_U553 , P2_R1158_U554 , P2_R1158_U555 , P2_R1158_U556 , P2_R1158_U557 , P2_R1158_U558 , P2_R1158_U559 , P2_R1158_U560;
wire P2_R1158_U561 , P2_R1158_U562 , P2_R1158_U563 , P2_R1158_U564 , P2_R1158_U565 , P2_R1158_U566 , P2_R1158_U567 , P2_R1158_U568 , P2_R1158_U569 , P2_R1158_U570;
wire P2_R1158_U571 , P2_R1158_U572 , P2_R1158_U573 , P2_R1158_U574 , P2_R1158_U575 , P2_R1158_U576 , P2_R1158_U577 , P2_R1158_U578 , P2_R1158_U579 , P2_R1158_U580;
wire P2_R1158_U581 , P2_R1158_U582 , P2_R1158_U583 , P2_R1158_U584 , P2_R1158_U585 , P2_R1158_U586 , P2_R1158_U587 , P2_R1158_U588 , P2_R1158_U589 , P2_R1158_U590;
wire P2_R1158_U591 , P2_R1158_U592 , P2_R1158_U593 , P2_R1158_U594 , P2_R1158_U595 , P2_R1158_U596 , P2_R1158_U597 , P2_R1158_U598 , P2_R1158_U599 , P2_R1158_U600;
wire P2_R1158_U601 , P2_R1158_U602 , P2_R1158_U603 , P2_R1158_U604 , P2_R1158_U605 , P2_R1158_U606 , P2_R1158_U607 , P2_R1158_U608 , P2_R1158_U609 , P2_R1158_U610;
wire P2_R1158_U611 , P2_R1158_U612 , P2_R1158_U613 , P2_R1158_U614 , P2_R1158_U615 , P2_R1158_U616 , P2_R1158_U617 , P2_R1158_U618 , P2_R1158_U619 , P2_R1158_U620;
wire P2_R1158_U621 , P2_R1158_U622 , P2_R1158_U623 , P2_R1158_U624 , P2_R1158_U625 , P2_R1158_U626 , P2_R1158_U627 , P2_R1158_U628 , P2_R1158_U629 , P2_R1158_U630;
wire P2_R1158_U631 , P2_R1158_U632 , P2_R1158_U633 , P2_R1158_U634 , P2_R1131_U6 , P2_R1131_U7 , P2_R1131_U8 , P2_R1131_U9 , P2_R1131_U10 , P2_R1131_U11;
wire P2_R1131_U12 , P2_R1131_U13 , P2_R1131_U14 , P2_R1131_U15 , P2_R1131_U16 , P2_R1131_U17 , P2_R1131_U18 , P2_R1131_U19 , P2_R1131_U20 , P2_R1131_U21;
wire P2_R1131_U22 , P2_R1131_U23 , P2_R1131_U24 , P2_R1131_U25 , P2_R1131_U26 , P2_R1131_U27 , P2_R1131_U28 , P2_R1131_U29 , P2_R1131_U30 , P2_R1131_U31;
wire P2_R1131_U32 , P2_R1131_U33 , P2_R1131_U34 , P2_R1131_U35 , P2_R1131_U36 , P2_R1131_U37 , P2_R1131_U38 , P2_R1131_U39 , P2_R1131_U40 , P2_R1131_U41;
wire P2_R1131_U42 , P2_R1131_U43 , P2_R1131_U44 , P2_R1131_U45 , P2_R1131_U46 , P2_R1131_U47 , P2_R1131_U48 , P2_R1131_U49 , P2_R1131_U50 , P2_R1131_U51;
wire P2_R1131_U52 , P2_R1131_U53 , P2_R1131_U54 , P2_R1131_U55 , P2_R1131_U56 , P2_R1131_U57 , P2_R1131_U58 , P2_R1131_U59 , P2_R1131_U60 , P2_R1131_U61;
wire P2_R1131_U62 , P2_R1131_U63 , P2_R1131_U64 , P2_R1131_U65 , P2_R1131_U66 , P2_R1131_U67 , P2_R1131_U68 , P2_R1131_U69 , P2_R1131_U70 , P2_R1131_U71;
wire P2_R1131_U72 , P2_R1131_U73 , P2_R1131_U74 , P2_R1131_U75 , P2_R1131_U76 , P2_R1131_U77 , P2_R1131_U78 , P2_R1131_U79 , P2_R1131_U80 , P2_R1131_U81;
wire P2_R1131_U82 , P2_R1131_U83 , P2_R1131_U84 , P2_R1131_U85 , P2_R1131_U86 , P2_R1131_U87 , P2_R1131_U88 , P2_R1131_U89 , P2_R1131_U90 , P2_R1131_U91;
wire P2_R1131_U92 , P2_R1131_U93 , P2_R1131_U94 , P2_R1131_U95 , P2_R1131_U96 , P2_R1131_U97 , P2_R1131_U98 , P2_R1131_U99 , P2_R1131_U100 , P2_R1131_U101;
wire P2_R1131_U102 , P2_R1131_U103 , P2_R1131_U104 , P2_R1131_U105 , P2_R1131_U106 , P2_R1131_U107 , P2_R1131_U108 , P2_R1131_U109 , P2_R1131_U110 , P2_R1131_U111;
wire P2_R1131_U112 , P2_R1131_U113 , P2_R1131_U114 , P2_R1131_U115 , P2_R1131_U116 , P2_R1131_U117 , P2_R1131_U118 , P2_R1131_U119 , P2_R1131_U120 , P2_R1131_U121;
wire P2_R1131_U122 , P2_R1131_U123 , P2_R1131_U124 , P2_R1131_U125 , P2_R1131_U126 , P2_R1131_U127 , P2_R1131_U128 , P2_R1131_U129 , P2_R1131_U130 , P2_R1131_U131;
wire P2_R1131_U132 , P2_R1131_U133 , P2_R1131_U134 , P2_R1131_U135 , P2_R1131_U136 , P2_R1131_U137 , P2_R1131_U138 , P2_R1131_U139 , P2_R1131_U140 , P2_R1131_U141;
wire P2_R1131_U142 , P2_R1131_U143 , P2_R1131_U144 , P2_R1131_U145 , P2_R1131_U146 , P2_R1131_U147 , P2_R1131_U148 , P2_R1131_U149 , P2_R1131_U150 , P2_R1131_U151;
wire P2_R1131_U152 , P2_R1131_U153 , P2_R1131_U154 , P2_R1131_U155 , P2_R1131_U156 , P2_R1131_U157 , P2_R1131_U158 , P2_R1131_U159 , P2_R1131_U160 , P2_R1131_U161;
wire P2_R1131_U162 , P2_R1131_U163 , P2_R1131_U164 , P2_R1131_U165 , P2_R1131_U166 , P2_R1131_U167 , P2_R1131_U168 , P2_R1131_U169 , P2_R1131_U170 , P2_R1131_U171;
wire P2_R1131_U172 , P2_R1131_U173 , P2_R1131_U174 , P2_R1131_U175 , P2_R1131_U176 , P2_R1131_U177 , P2_R1131_U178 , P2_R1131_U179 , P2_R1131_U180 , P2_R1131_U181;
wire P2_R1131_U182 , P2_R1131_U183 , P2_R1131_U184 , P2_R1131_U185 , P2_R1131_U186 , P2_R1131_U187 , P2_R1131_U188 , P2_R1131_U189 , P2_R1131_U190 , P2_R1131_U191;
wire P2_R1131_U192 , P2_R1131_U193 , P2_R1131_U194 , P2_R1131_U195 , P2_R1131_U196 , P2_R1131_U197 , P2_R1131_U198 , P2_R1131_U199 , P2_R1131_U200 , P2_R1131_U201;
wire P2_R1131_U202 , P2_R1131_U203 , P2_R1131_U204 , P2_R1131_U205 , P2_R1131_U206 , P2_R1131_U207 , P2_R1131_U208 , P2_R1131_U209 , P2_R1131_U210 , P2_R1131_U211;
wire P2_R1131_U212 , P2_R1131_U213 , P2_R1131_U214 , P2_R1131_U215 , P2_R1131_U216 , P2_R1131_U217 , P2_R1131_U218 , P2_R1131_U219 , P2_R1131_U220 , P2_R1131_U221;
wire P2_R1131_U222 , P2_R1131_U223 , P2_R1131_U224 , P2_R1131_U225 , P2_R1131_U226 , P2_R1131_U227 , P2_R1131_U228 , P2_R1131_U229 , P2_R1131_U230 , P2_R1131_U231;
wire P2_R1131_U232 , P2_R1131_U233 , P2_R1131_U234 , P2_R1131_U235 , P2_R1131_U236 , P2_R1131_U237 , P2_R1131_U238 , P2_R1131_U239 , P2_R1131_U240 , P2_R1131_U241;
wire P2_R1131_U242 , P2_R1131_U243 , P2_R1131_U244 , P2_R1131_U245 , P2_R1131_U246 , P2_R1131_U247 , P2_R1131_U248 , P2_R1131_U249 , P2_R1131_U250 , P2_R1131_U251;
wire P2_R1131_U252 , P2_R1131_U253 , P2_R1131_U254 , P2_R1131_U255 , P2_R1131_U256 , P2_R1131_U257 , P2_R1131_U258 , P2_R1131_U259 , P2_R1131_U260 , P2_R1131_U261;
wire P2_R1131_U262 , P2_R1131_U263 , P2_R1131_U264 , P2_R1131_U265 , P2_R1131_U266 , P2_R1131_U267 , P2_R1131_U268 , P2_R1131_U269 , P2_R1131_U270 , P2_R1131_U271;
wire P2_R1131_U272 , P2_R1131_U273 , P2_R1131_U274 , P2_R1131_U275 , P2_R1131_U276 , P2_R1131_U277 , P2_R1131_U278 , P2_R1131_U279 , P2_R1131_U280 , P2_R1131_U281;
wire P2_R1131_U282 , P2_R1131_U283 , P2_R1131_U284 , P2_R1131_U285 , P2_R1131_U286 , P2_R1131_U287 , P2_R1131_U288 , P2_R1131_U289 , P2_R1131_U290 , P2_R1131_U291;
wire P2_R1131_U292 , P2_R1131_U293 , P2_R1131_U294 , P2_R1131_U295 , P2_R1131_U296 , P2_R1131_U297 , P2_R1131_U298 , P2_R1131_U299 , P2_R1131_U300 , P2_R1131_U301;
wire P2_R1131_U302 , P2_R1131_U303 , P2_R1131_U304 , P2_R1131_U305 , P2_R1131_U306 , P2_R1131_U307 , P2_R1131_U308 , P2_R1131_U309 , P2_R1131_U310 , P2_R1131_U311;
wire P2_R1131_U312 , P2_R1131_U313 , P2_R1131_U314 , P2_R1131_U315 , P2_R1131_U316 , P2_R1131_U317 , P2_R1131_U318 , P2_R1131_U319 , P2_R1131_U320 , P2_R1131_U321;
wire P2_R1131_U322 , P2_R1131_U323 , P2_R1131_U324 , P2_R1131_U325 , P2_R1131_U326 , P2_R1131_U327 , P2_R1131_U328 , P2_R1131_U329 , P2_R1131_U330 , P2_R1131_U331;
wire P2_R1131_U332 , P2_R1131_U333 , P2_R1131_U334 , P2_R1131_U335 , P2_R1131_U336 , P2_R1131_U337 , P2_R1131_U338 , P2_R1131_U339 , P2_R1131_U340 , P2_R1131_U341;
wire P2_R1131_U342 , P2_R1131_U343 , P2_R1131_U344 , P2_R1131_U345 , P2_R1131_U346 , P2_R1131_U347 , P2_R1131_U348 , P2_R1131_U349 , P2_R1131_U350 , P2_R1131_U351;
wire P2_R1131_U352 , P2_R1131_U353 , P2_R1131_U354 , P2_R1131_U355 , P2_R1131_U356 , P2_R1131_U357 , P2_R1131_U358 , P2_R1131_U359 , P2_R1131_U360 , P2_R1131_U361;
wire P2_R1131_U362 , P2_R1131_U363 , P2_R1131_U364 , P2_R1131_U365 , P2_R1131_U366 , P2_R1131_U367 , P2_R1131_U368 , P2_R1131_U369 , P2_R1131_U370 , P2_R1131_U371;
wire P2_R1131_U372 , P2_R1131_U373 , P2_R1131_U374 , P2_R1131_U375 , P2_R1131_U376 , P2_R1131_U377 , P2_R1131_U378 , P2_R1131_U379 , P2_R1131_U380 , P2_R1131_U381;
wire P2_R1131_U382 , P2_R1131_U383 , P2_R1131_U384 , P2_R1131_U385 , P2_R1131_U386 , P2_R1131_U387 , P2_R1131_U388 , P2_R1131_U389 , P2_R1131_U390 , P2_R1131_U391;
wire P2_R1131_U392 , P2_R1131_U393 , P2_R1131_U394 , P2_R1131_U395 , P2_R1131_U396 , P2_R1131_U397 , P2_R1131_U398 , P2_R1131_U399 , P2_R1131_U400 , P2_R1131_U401;
wire P2_R1131_U402 , P2_R1131_U403 , P2_R1131_U404 , P2_R1131_U405 , P2_R1131_U406 , P2_R1131_U407 , P2_R1131_U408 , P2_R1131_U409 , P2_R1131_U410 , P2_R1131_U411;
wire P2_R1131_U412 , P2_R1131_U413 , P2_R1131_U414 , P2_R1131_U415 , P2_R1131_U416 , P2_R1131_U417 , P2_R1131_U418 , P2_R1131_U419 , P2_R1131_U420 , P2_R1131_U421;
wire P2_R1131_U422 , P2_R1131_U423 , P2_R1131_U424 , P2_R1131_U425 , P2_R1131_U426 , P2_R1131_U427 , P2_R1131_U428 , P2_R1131_U429 , P2_R1131_U430 , P2_R1131_U431;
wire P2_R1131_U432 , P2_R1131_U433 , P2_R1131_U434 , P2_R1131_U435 , P2_R1131_U436 , P2_R1131_U437 , P2_R1131_U438 , P2_R1131_U439 , P2_R1131_U440 , P2_R1131_U441;
wire P2_R1131_U442 , P2_R1131_U443 , P2_R1131_U444 , P2_R1131_U445 , P2_R1131_U446 , P2_R1131_U447 , P2_R1131_U448 , P2_R1131_U449 , P2_R1131_U450 , P2_R1131_U451;
wire P2_R1131_U452 , P2_R1131_U453 , P2_R1131_U454 , P2_R1131_U455 , P2_R1131_U456 , P2_R1131_U457 , P2_R1131_U458 , P2_R1131_U459 , P2_R1131_U460 , P2_R1131_U461;
wire P2_R1131_U462 , P2_R1131_U463 , P2_R1131_U464 , P2_R1131_U465 , P2_R1131_U466 , P2_R1131_U467 , P2_R1131_U468 , P2_R1131_U469 , P2_R1131_U470 , P2_R1131_U471;
wire P2_R1131_U472 , P2_R1131_U473 , P2_R1131_U474 , P2_R1131_U475 , P2_R1131_U476 , P2_R1131_U477 , P2_R1131_U478 , P2_R1131_U479 , P2_R1131_U480 , P2_R1131_U481;
wire P2_R1131_U482 , P2_R1131_U483 , P2_R1131_U484 , P2_R1131_U485 , P2_R1131_U486 , P2_R1131_U487 , P2_R1131_U488 , P2_R1131_U489 , P2_R1054_U6 , P2_R1054_U7;
wire P2_R1054_U8 , P2_R1054_U9 , P2_R1054_U10 , P2_R1054_U11 , P2_R1054_U12 , P2_R1054_U13 , P2_R1054_U14 , P2_R1054_U15 , P2_R1054_U16 , P2_R1054_U17;
wire P2_R1054_U18 , P2_R1054_U19 , P2_R1054_U20 , P2_R1054_U21 , P2_R1054_U22 , P2_R1054_U23 , P2_R1054_U24 , P2_R1054_U25 , P2_R1054_U26 , P2_R1054_U27;
wire P2_R1054_U28 , P2_R1054_U29 , P2_R1054_U30 , P2_R1054_U31 , P2_R1054_U32 , P2_R1054_U33 , P2_R1054_U34 , P2_R1054_U35 , P2_R1054_U36 , P2_R1054_U37;
wire P2_R1054_U38 , P2_R1054_U39 , P2_R1054_U40 , P2_R1054_U41 , P2_R1054_U42 , P2_R1054_U43 , P2_R1054_U44 , P2_R1054_U45 , P2_R1054_U46 , P2_R1054_U47;
wire P2_R1054_U48 , P2_R1054_U49 , P2_R1054_U50 , P2_R1054_U51 , P2_R1054_U52 , P2_R1054_U53 , P2_R1054_U54 , P2_R1054_U55 , P2_R1054_U56 , P2_R1054_U57;
wire P2_R1054_U58 , P2_R1054_U59 , P2_R1054_U60 , P2_R1054_U61 , P2_R1054_U62 , P2_R1054_U63 , P2_R1054_U64 , P2_R1054_U65 , P2_R1054_U66 , P2_R1054_U67;
wire P2_R1054_U68 , P2_R1054_U69 , P2_R1054_U70 , P2_R1054_U71 , P2_R1054_U72 , P2_R1054_U73 , P2_R1054_U74 , P2_R1054_U75 , P2_R1054_U76 , P2_R1054_U77;
wire P2_R1054_U78 , P2_R1054_U79 , P2_R1054_U80 , P2_R1054_U81 , P2_R1054_U82 , P2_R1054_U83 , P2_R1054_U84 , P2_R1054_U85 , P2_R1054_U86 , P2_R1054_U87;
wire P2_R1054_U88 , P2_R1054_U89 , P2_R1054_U90 , P2_R1054_U91 , P2_R1054_U92 , P2_R1054_U93 , P2_R1054_U94 , P2_R1054_U95 , P2_R1054_U96 , P2_R1054_U97;
wire P2_R1054_U98 , P2_R1054_U99 , P2_R1054_U100 , P2_R1054_U101 , P2_R1054_U102 , P2_R1054_U103 , P2_R1054_U104 , P2_R1054_U105 , P2_R1054_U106 , P2_R1054_U107;
wire P2_R1054_U108 , P2_R1054_U109 , P2_R1054_U110 , P2_R1054_U111 , P2_R1054_U112 , P2_R1054_U113 , P2_R1054_U114 , P2_R1054_U115 , P2_R1054_U116 , P2_R1054_U117;
wire P2_R1054_U118 , P2_R1054_U119 , P2_R1054_U120 , P2_R1054_U121 , P2_R1054_U122 , P2_R1054_U123 , P2_R1054_U124 , P2_R1054_U125 , P2_R1054_U126 , P2_R1054_U127;
wire P2_R1054_U128 , P2_R1054_U129 , P2_R1054_U130 , P2_R1054_U131 , P2_R1054_U132 , P2_R1054_U133 , P2_R1054_U134 , P2_R1054_U135 , P2_R1054_U136 , P2_R1054_U137;
wire P2_R1054_U138 , P2_R1054_U139 , P2_R1054_U140 , P2_R1054_U141 , P2_R1054_U142 , P2_R1054_U143 , P2_R1054_U144 , P2_R1054_U145 , P2_R1054_U146 , P2_R1054_U147;
wire P2_R1054_U148 , P2_R1054_U149 , P2_R1054_U150 , P2_R1054_U151 , P2_R1054_U152 , P2_R1054_U153 , P2_R1054_U154 , P2_R1054_U155 , P2_R1054_U156 , P2_R1054_U157;
wire P2_R1054_U158 , P2_R1054_U159 , P2_R1054_U160 , P2_R1054_U161 , P2_R1054_U162 , P2_R1054_U163 , P2_R1054_U164 , P2_R1054_U165 , P2_R1054_U166 , P2_R1054_U167;
wire P2_R1054_U168 , P2_R1054_U169 , P2_R1054_U170 , P2_R1054_U171 , P2_R1054_U172 , P2_R1054_U173 , P2_R1054_U174 , P2_R1054_U175 , P2_R1054_U176 , P2_R1054_U177;
wire P2_R1054_U178 , P2_R1054_U179 , P2_R1054_U180 , P2_R1054_U181 , P2_R1054_U182 , P2_R1054_U183 , P2_R1054_U184 , P2_R1054_U185 , P2_R1054_U186 , P2_R1054_U187;
wire P2_R1054_U188 , P2_R1054_U189 , P2_R1054_U190 , P2_R1054_U191 , P2_R1054_U192 , P2_R1054_U193 , P2_R1054_U194 , P2_R1054_U195 , P2_R1054_U196 , P2_R1054_U197;
wire P2_R1054_U198 , P2_R1054_U199 , P2_R1054_U200 , P2_R1054_U201 , P2_R1054_U202 , P2_R1054_U203 , P2_R1054_U204 , P2_R1054_U205 , P2_R1054_U206 , P2_R1054_U207;
wire P2_R1054_U208 , P2_R1054_U209 , P2_R1054_U210 , P2_R1054_U211 , P2_R1054_U212 , P2_R1054_U213 , P2_R1054_U214 , P2_R1054_U215 , P2_R1054_U216 , P2_R1054_U217;
wire P2_R1054_U218 , P2_R1054_U219 , P2_R1054_U220 , P2_R1054_U221 , P2_R1054_U222 , P2_R1054_U223 , P2_R1054_U224 , P2_R1054_U225 , P2_R1054_U226 , P2_R1054_U227;
wire P2_R1054_U228 , P2_R1054_U229 , P2_R1054_U230 , P2_R1054_U231 , P2_R1054_U232 , P2_R1054_U233 , P2_R1054_U234 , P2_R1054_U235 , P2_R1054_U236 , P2_R1054_U237;
wire P2_R1054_U238 , P2_R1054_U239 , P2_R1054_U240 , P2_R1054_U241 , P2_R1054_U242 , P2_R1054_U243 , P2_R1054_U244 , P2_R1054_U245 , P2_R1054_U246 , P2_R1054_U247;
wire P2_R1054_U248 , P2_R1054_U249 , P2_R1054_U250 , P2_R1054_U251 , P2_R1054_U252 , P2_R1054_U253 , P2_R1054_U254 , P2_R1054_U255 , P2_R1054_U256 , P2_R1054_U257;
wire P2_R1054_U258 , P2_R1054_U259 , P2_R1054_U260 , P2_R1054_U261 , P2_R1054_U262 , P2_R1054_U263 , P2_R1054_U264 , P2_R1054_U265 , P2_R1054_U266 , P2_R1054_U267;
wire P2_R1054_U268 , P2_R1054_U269 , P2_R1054_U270 , P2_R1054_U271 , P2_R1054_U272 , P2_R1054_U273 , P2_R1054_U274 , P2_R1054_U275 , P2_R1054_U276 , P2_R1054_U277;
wire P2_R1054_U278 , P2_R1054_U279 , P2_R1054_U280 , P2_R1054_U281 , P2_R1054_U282 , P2_R1054_U283 , P2_R1054_U284 , P2_R1054_U285 , P2_R1054_U286 , P2_R1054_U287;
wire P2_R1054_U288 , P2_R1054_U289 , P2_R1054_U290 , P2_R1054_U291 , P2_R1054_U292 , P2_R1054_U293 , P2_R1054_U294 , P2_R1161_U4 , P2_R1161_U5 , P2_R1161_U6;
wire P2_R1161_U7 , P2_R1161_U8 , P2_R1161_U9 , P2_R1161_U10 , P2_R1161_U11 , P2_R1161_U12 , P2_R1161_U13 , P2_R1161_U14 , P2_R1161_U15 , P2_R1161_U16;
wire P2_R1161_U17 , P2_R1161_U18 , P2_R1161_U19 , P2_R1161_U20 , P2_R1161_U21 , P2_R1161_U22 , P2_R1161_U23 , P2_R1161_U24 , P2_R1161_U25 , P2_R1161_U26;
wire P2_R1161_U27 , P2_R1161_U28 , P2_R1161_U29 , P2_R1161_U30 , P2_R1161_U31 , P2_R1161_U32 , P2_R1161_U33 , P2_R1161_U34 , P2_R1161_U35 , P2_R1161_U36;
wire P2_R1161_U37 , P2_R1161_U38 , P2_R1161_U39 , P2_R1161_U40 , P2_R1161_U41 , P2_R1161_U42 , P2_R1161_U43 , P2_R1161_U44 , P2_R1161_U45 , P2_R1161_U46;
wire P2_R1161_U47 , P2_R1161_U48 , P2_R1161_U49 , P2_R1161_U50 , P2_R1161_U51 , P2_R1161_U52 , P2_R1161_U53 , P2_R1161_U54 , P2_R1161_U55 , P2_R1161_U56;
wire P2_R1161_U57 , P2_R1161_U58 , P2_R1161_U59 , P2_R1161_U60 , P2_R1161_U61 , P2_R1161_U62 , P2_R1161_U63 , P2_R1161_U64 , P2_R1161_U65 , P2_R1161_U66;
wire P2_R1161_U67 , P2_R1161_U68 , P2_R1161_U69 , P2_R1161_U70 , P2_R1161_U71 , P2_R1161_U72 , P2_R1161_U73 , P2_R1161_U74 , P2_R1161_U75 , P2_R1161_U76;
wire P2_R1161_U77 , P2_R1161_U78 , P2_R1161_U79 , P2_R1161_U80 , P2_R1161_U81 , P2_R1161_U82 , P2_R1161_U83 , P2_R1161_U84 , P2_R1161_U85 , P2_R1161_U86;
wire P2_R1161_U87 , P2_R1161_U88 , P2_R1161_U89 , P2_R1161_U90 , P2_R1161_U91 , P2_R1161_U92 , P2_R1161_U93 , P2_R1161_U94 , P2_R1161_U95 , P2_R1161_U96;
wire P2_R1161_U97 , P2_R1161_U98 , P2_R1161_U99 , P2_R1161_U100 , P2_R1161_U101 , P2_R1161_U102 , P2_R1161_U103 , P2_R1161_U104 , P2_R1161_U105 , P2_R1161_U106;
wire P2_R1161_U107 , P2_R1161_U108 , P2_R1161_U109 , P2_R1161_U110 , P2_R1161_U111 , P2_R1161_U112 , P2_R1161_U113 , P2_R1161_U114 , P2_R1161_U115 , P2_R1161_U116;
wire P2_R1161_U117 , P2_R1161_U118 , P2_R1161_U119 , P2_R1161_U120 , P2_R1161_U121 , P2_R1161_U122 , P2_R1161_U123 , P2_R1161_U124 , P2_R1161_U125 , P2_R1161_U126;
wire P2_R1161_U127 , P2_R1161_U128 , P2_R1161_U129 , P2_R1161_U130 , P2_R1161_U131 , P2_R1161_U132 , P2_R1161_U133 , P2_R1161_U134 , P2_R1161_U135 , P2_R1161_U136;
wire P2_R1161_U137 , P2_R1161_U138 , P2_R1161_U139 , P2_R1161_U140 , P2_R1161_U141 , P2_R1161_U142 , P2_R1161_U143 , P2_R1161_U144 , P2_R1161_U145 , P2_R1161_U146;
wire P2_R1161_U147 , P2_R1161_U148 , P2_R1161_U149 , P2_R1161_U150 , P2_R1161_U151 , P2_R1161_U152 , P2_R1161_U153 , P2_R1161_U154 , P2_R1161_U155 , P2_R1161_U156;
wire P2_R1161_U157 , P2_R1161_U158 , P2_R1161_U159 , P2_R1161_U160 , P2_R1161_U161 , P2_R1161_U162 , P2_R1161_U163 , P2_R1161_U164 , P2_R1161_U165 , P2_R1161_U166;
wire P2_R1161_U167 , P2_R1161_U168 , P2_R1161_U169 , P2_R1161_U170 , P2_R1161_U171 , P2_R1161_U172 , P2_R1161_U173 , P2_R1161_U174 , P2_R1161_U175 , P2_R1161_U176;
wire P2_R1161_U177 , P2_R1161_U178 , P2_R1161_U179 , P2_R1161_U180 , P2_R1161_U181 , P2_R1161_U182 , P2_R1161_U183 , P2_R1161_U184 , P2_R1161_U185 , P2_R1161_U186;
wire P2_R1161_U187 , P2_R1161_U188 , P2_R1161_U189 , P2_R1161_U190 , P2_R1161_U191 , P2_R1161_U192 , P2_R1161_U193 , P2_R1161_U194 , P2_R1161_U195 , P2_R1161_U196;
wire P2_R1161_U197 , P2_R1161_U198 , P2_R1161_U199 , P2_R1161_U200 , P2_R1161_U201 , P2_R1161_U202 , P2_R1161_U203 , P2_R1161_U204 , P2_R1161_U205 , P2_R1161_U206;
wire P2_R1161_U207 , P2_R1161_U208 , P2_R1161_U209 , P2_R1161_U210 , P2_R1161_U211 , P2_R1161_U212 , P2_R1161_U213 , P2_R1161_U214 , P2_R1161_U215 , P2_R1161_U216;
wire P2_R1161_U217 , P2_R1161_U218 , P2_R1161_U219 , P2_R1161_U220 , P2_R1161_U221 , P2_R1161_U222 , P2_R1161_U223 , P2_R1161_U224 , P2_R1161_U225 , P2_R1161_U226;
wire P2_R1161_U227 , P2_R1161_U228 , P2_R1161_U229 , P2_R1161_U230 , P2_R1161_U231 , P2_R1161_U232 , P2_R1161_U233 , P2_R1161_U234 , P2_R1161_U235 , P2_R1161_U236;
wire P2_R1161_U237 , P2_R1161_U238 , P2_R1161_U239 , P2_R1161_U240 , P2_R1161_U241 , P2_R1161_U242 , P2_R1161_U243 , P2_R1161_U244 , P2_R1161_U245 , P2_R1161_U246;
wire P2_R1161_U247 , P2_R1161_U248 , P2_R1161_U249 , P2_R1161_U250 , P2_R1161_U251 , P2_R1161_U252 , P2_R1161_U253 , P2_R1161_U254 , P2_R1161_U255 , P2_R1161_U256;
wire P2_R1161_U257 , P2_R1161_U258 , P2_R1161_U259 , P2_R1161_U260 , P2_R1161_U261 , P2_R1161_U262 , P2_R1161_U263 , P2_R1161_U264 , P2_R1161_U265 , P2_R1161_U266;
wire P2_R1161_U267 , P2_R1161_U268 , P2_R1161_U269 , P2_R1161_U270 , P2_R1161_U271 , P2_R1161_U272 , P2_R1161_U273 , P2_R1161_U274 , P2_R1161_U275 , P2_R1161_U276;
wire P2_R1161_U277 , P2_R1161_U278 , P2_R1161_U279 , P2_R1161_U280 , P2_R1161_U281 , P2_R1161_U282 , P2_R1161_U283 , P2_R1161_U284 , P2_R1161_U285 , P2_R1161_U286;
wire P2_R1161_U287 , P2_R1161_U288 , P2_R1161_U289 , P2_R1161_U290 , P2_R1161_U291 , P2_R1161_U292 , P2_R1161_U293 , P2_R1161_U294 , P2_R1161_U295 , P2_R1161_U296;
wire P2_R1161_U297 , P2_R1161_U298 , P2_R1161_U299 , P2_R1161_U300 , P2_R1161_U301 , P2_R1161_U302 , P2_R1161_U303 , P2_R1161_U304 , P2_R1161_U305 , P2_R1161_U306;
wire P2_R1161_U307 , P2_R1161_U308 , P2_R1161_U309 , P2_R1161_U310 , P2_R1161_U311 , P2_R1161_U312 , P2_R1161_U313 , P2_R1161_U314 , P2_R1161_U315 , P2_R1161_U316;
wire P2_R1161_U317 , P2_R1161_U318 , P2_R1161_U319 , P2_R1161_U320 , P2_R1161_U321 , P2_R1161_U322 , P2_R1161_U323 , P2_R1161_U324 , P2_R1161_U325 , P2_R1161_U326;
wire P2_R1161_U327 , P2_R1161_U328 , P2_R1161_U329 , P2_R1161_U330 , P2_R1161_U331 , P2_R1161_U332 , P2_R1161_U333 , P2_R1161_U334 , P2_R1161_U335 , P2_R1161_U336;
wire P2_R1161_U337 , P2_R1161_U338 , P2_R1161_U339 , P2_R1161_U340 , P2_R1161_U341 , P2_R1161_U342 , P2_R1161_U343 , P2_R1161_U344 , P2_R1161_U345 , P2_R1161_U346;
wire P2_R1161_U347 , P2_R1161_U348 , P2_R1161_U349 , P2_R1161_U350 , P2_R1161_U351 , P2_R1161_U352 , P2_R1161_U353 , P2_R1161_U354 , P2_R1161_U355 , P2_R1161_U356;
wire P2_R1161_U357 , P2_R1161_U358 , P2_R1161_U359 , P2_R1161_U360 , P2_R1161_U361 , P2_R1161_U362 , P2_R1161_U363 , P2_R1161_U364 , P2_R1161_U365 , P2_R1161_U366;
wire P2_R1161_U367 , P2_R1161_U368 , P2_R1161_U369 , P2_R1161_U370 , P2_R1161_U371 , P2_R1161_U372 , P2_R1161_U373 , P2_R1161_U374 , P2_R1161_U375 , P2_R1161_U376;
wire P2_R1161_U377 , P2_R1161_U378 , P2_R1161_U379 , P2_R1161_U380 , P2_R1161_U381 , P2_R1161_U382 , P2_R1161_U383 , P2_R1161_U384 , P2_R1161_U385 , P2_R1161_U386;
wire P2_R1161_U387 , P2_R1161_U388 , P2_R1161_U389 , P2_R1161_U390 , P2_R1161_U391 , P2_R1161_U392 , P2_R1161_U393 , P2_R1161_U394 , P2_R1161_U395 , P2_R1161_U396;
wire P2_R1161_U397 , P2_R1161_U398 , P2_R1161_U399 , P2_R1161_U400 , P2_R1161_U401 , P2_R1161_U402 , P2_R1161_U403 , P2_R1161_U404 , P2_R1161_U405 , P2_R1161_U406;
wire P2_R1161_U407 , P2_R1161_U408 , P2_R1161_U409 , P2_R1161_U410 , P2_R1161_U411 , P2_R1161_U412 , P2_R1161_U413 , P2_R1161_U414 , P2_R1161_U415 , P2_R1161_U416;
wire P2_R1161_U417 , P2_R1161_U418 , P2_R1161_U419 , P2_R1161_U420 , P2_R1161_U421 , P2_R1161_U422 , P2_R1161_U423 , P2_R1161_U424 , P2_R1161_U425 , P2_R1161_U426;
wire P2_R1161_U427 , P2_R1161_U428 , P2_R1161_U429 , P2_R1161_U430 , P2_R1161_U431 , P2_R1161_U432 , P2_R1161_U433 , P2_R1161_U434 , P2_R1161_U435 , P2_R1161_U436;
wire P2_R1161_U437 , P2_R1161_U438 , P2_R1161_U439 , P2_R1161_U440 , P2_R1161_U441 , P2_R1161_U442 , P2_R1161_U443 , P2_R1161_U444 , P2_R1161_U445 , P2_R1161_U446;


nand NAND2_1 ( P2_R1161_U504 , P2_U3387 , P2_R1161_U30 );
nand NAND2_2 ( P2_R1161_U503 , P2_U3076 , P2_R1161_U29 );
nand NAND2_3 ( P2_R1161_U502 , P2_U3419 , P2_R1161_U64 );
nand NAND2_4 ( U25 , U136 , U135 );
nand NAND2_5 ( U26 , U138 , U137 );
nand NAND2_6 ( U27 , U140 , U139 );
nand NAND2_7 ( U28 , U142 , U141 );
nand NAND2_8 ( U29 , U144 , U143 );
nand NAND2_9 ( U30 , U146 , U145 );
nand NAND2_10 ( U31 , U148 , U147 );
nand NAND2_11 ( U32 , U150 , U149 );
nand NAND2_12 ( U33 , U152 , U151 );
nand NAND2_13 ( U34 , U154 , U153 );
nand NAND2_14 ( U35 , U156 , U155 );
nand NAND2_15 ( U36 , U158 , U157 );
nand NAND2_16 ( U37 , U160 , U159 );
nand NAND2_17 ( U38 , U162 , U161 );
nand NAND2_18 ( U39 , U164 , U163 );
nand NAND2_19 ( U40 , U166 , U165 );
nand NAND2_20 ( U41 , U168 , U167 );
nand NAND2_21 ( U42 , U170 , U169 );
nand NAND2_22 ( U43 , U172 , U171 );
nand NAND2_23 ( U44 , U174 , U173 );
nand NAND2_24 ( U45 , U176 , U175 );
nand NAND2_25 ( U46 , U178 , U177 );
nand NAND2_26 ( U47 , U180 , U179 );
nand NAND2_27 ( U48 , U182 , U181 );
nand NAND2_28 ( U49 , U184 , U183 );
nand NAND2_29 ( U50 , U186 , U185 );
nand NAND2_30 ( U51 , U188 , U187 );
nand NAND2_31 ( U52 , U190 , U189 );
nand NAND2_32 ( U53 , U192 , U191 );
nand NAND2_33 ( U54 , U194 , U193 );
nand NAND2_34 ( U55 , U196 , U195 );
nand NAND2_35 ( U56 , U198 , U197 );
nand NAND2_36 ( U57 , U200 , U199 );
nand NAND2_37 ( U58 , U202 , U201 );
nand NAND2_38 ( U59 , U204 , U203 );
nand NAND2_39 ( U60 , U206 , U205 );
nand NAND2_40 ( U61 , U208 , U207 );
nand NAND2_41 ( U62 , U210 , U209 );
nand NAND2_42 ( U63 , U212 , U211 );
nand NAND2_43 ( U64 , U214 , U213 );
nand NAND2_44 ( U65 , U216 , U215 );
nand NAND2_45 ( U66 , U218 , U217 );
nand NAND2_46 ( U67 , U220 , U219 );
nand NAND2_47 ( U68 , U222 , U221 );
nand NAND2_48 ( U69 , U224 , U223 );
nand NAND2_49 ( U70 , U226 , U225 );
nand NAND2_50 ( U71 , U228 , U227 );
nand NAND2_51 ( U72 , U230 , U229 );
nand NAND2_52 ( U73 , U232 , U231 );
nand NAND2_53 ( U74 , U234 , U233 );
nand NAND2_54 ( U75 , U236 , U235 );
nand NAND2_55 ( U76 , U238 , U237 );
nand NAND2_56 ( U77 , U240 , U239 );
nand NAND2_57 ( U78 , U242 , U241 );
nand NAND2_58 ( U79 , U244 , U243 );
nand NAND2_59 ( U80 , U246 , U245 );
nand NAND2_60 ( U81 , U248 , U247 );
nand NAND2_61 ( U82 , U250 , U249 );
nand NAND2_62 ( U83 , U252 , U251 );
nand NAND2_63 ( U84 , U254 , U253 );
nand NAND2_64 ( U85 , U256 , U255 );
nand NAND2_65 ( U86 , U258 , U257 );
nand NAND2_66 ( U87 , U260 , U259 );
nand NAND2_67 ( U88 , U262 , U261 );
nand NAND2_68 ( U89 , U264 , U263 );
nand NAND2_69 ( U90 , U266 , U265 );
nand NAND2_70 ( U91 , U268 , U267 );
nand NAND2_71 ( U92 , U270 , U269 );
nand NAND2_72 ( U93 , U272 , U271 );
nand NAND2_73 ( U94 , U274 , U273 );
nand NAND2_74 ( U95 , U276 , U275 );
nand NAND2_75 ( U96 , U278 , U277 );
nand NAND2_76 ( U97 , U280 , U279 );
nand NAND2_77 ( U98 , U282 , U281 );
nand NAND2_78 ( U99 , U284 , U283 );
nand NAND2_79 ( U100 , U286 , U285 );
nand NAND2_80 ( U101 , U288 , U287 );
nand NAND2_81 ( U102 , U290 , U289 );
nand NAND2_82 ( U103 , U292 , U291 );
nand NAND2_83 ( U104 , U294 , U293 );
nand NAND2_84 ( U105 , U296 , U295 );
nand NAND2_85 ( U106 , U298 , U297 );
nand NAND2_86 ( U107 , U300 , U299 );
nand NAND2_87 ( U108 , U302 , U301 );
nand NAND2_88 ( U109 , U304 , U303 );
nand NAND2_89 ( U110 , U306 , U305 );
nand NAND2_90 ( U111 , U308 , U307 );
nand NAND2_91 ( U112 , U310 , U309 );
nand NAND2_92 ( U113 , U312 , U311 );
nand NAND2_93 ( U114 , U314 , U313 );
nand NAND2_94 ( U115 , U316 , U315 );
nand NAND2_95 ( U116 , U318 , U317 );
nand NAND2_96 ( U117 , U320 , U319 );
nand NAND2_97 ( U118 , U322 , U321 );
nand NAND2_98 ( U119 , U324 , U323 );
nand NAND2_99 ( U120 , U326 , U325 );
not NOT1_100 ( U121 , P2_WR_REG );
not NOT1_101 ( U122 , P1_WR_REG );
and AND2_102 ( U123 , U132 , U131 );
not NOT1_103 ( U124 , P2_RD_REG );
not NOT1_104 ( U125 , P1_RD_REG );
and AND2_105 ( U126 , U134 , U133 );
nand NAND2_106 ( U127 , U129 , U128 );
nand NAND3_107 ( U128 , LT_1075_U6 , U125 , LT_1075_19_U6 );
nand NAND3_108 ( U129 , P1_ADDR_REG_19_ , U124 , P2_ADDR_REG_19_ );
not NOT1_109 ( U130 , U127 );
nand NAND2_110 ( U131 , P2_WR_REG , U122 );
nand NAND2_111 ( U132 , P1_WR_REG , U121 );
nand NAND2_112 ( U133 , P2_RD_REG , U125 );
nand NAND2_113 ( U134 , P1_RD_REG , U124 );
nand NAND2_114 ( U135 , P1_DATAO_REG_9_ , U127 );
nand NAND2_115 ( U136 , R140_U84 , U130 );
nand NAND2_116 ( U137 , P1_DATAO_REG_8_ , U127 );
nand NAND2_117 ( U138 , R140_U85 , U130 );
nand NAND2_118 ( U139 , P1_DATAO_REG_7_ , U127 );
nand NAND2_119 ( U140 , R140_U86 , U130 );
nand NAND2_120 ( U141 , P1_DATAO_REG_6_ , U127 );
nand NAND2_121 ( U142 , R140_U87 , U130 );
nand NAND2_122 ( U143 , P1_DATAO_REG_5_ , U127 );
nand NAND2_123 ( U144 , R140_U88 , U130 );
nand NAND2_124 ( U145 , P1_DATAO_REG_4_ , U127 );
nand NAND2_125 ( U146 , R140_U89 , U130 );
nand NAND2_126 ( U147 , P1_DATAO_REG_3_ , U127 );
nand NAND2_127 ( U148 , R140_U90 , U130 );
nand NAND2_128 ( U149 , P1_DATAO_REG_31_ , U127 );
nand NAND2_129 ( U150 , R140_U11 , U130 );
nand NAND2_130 ( U151 , P1_DATAO_REG_30_ , U127 );
nand NAND2_131 ( U152 , R140_U91 , U130 );
nand NAND2_132 ( U153 , P1_DATAO_REG_2_ , U127 );
nand NAND2_133 ( U154 , R140_U92 , U130 );
nand NAND2_134 ( U155 , P1_DATAO_REG_29_ , U127 );
nand NAND2_135 ( U156 , R140_U93 , U130 );
nand NAND2_136 ( U157 , P1_DATAO_REG_28_ , U127 );
nand NAND2_137 ( U158 , R140_U94 , U130 );
nand NAND2_138 ( U159 , P1_DATAO_REG_27_ , U127 );
nand NAND2_139 ( U160 , R140_U95 , U130 );
nand NAND2_140 ( U161 , P1_DATAO_REG_26_ , U127 );
nand NAND2_141 ( U162 , R140_U96 , U130 );
nand NAND2_142 ( U163 , P1_DATAO_REG_25_ , U127 );
nand NAND2_143 ( U164 , R140_U97 , U130 );
nand NAND2_144 ( U165 , P1_DATAO_REG_24_ , U127 );
nand NAND2_145 ( U166 , R140_U98 , U130 );
nand NAND2_146 ( U167 , P1_DATAO_REG_23_ , U127 );
nand NAND2_147 ( U168 , R140_U99 , U130 );
nand NAND2_148 ( U169 , P1_DATAO_REG_22_ , U127 );
nand NAND2_149 ( U170 , R140_U100 , U130 );
nand NAND2_150 ( U171 , P1_DATAO_REG_21_ , U127 );
nand NAND2_151 ( U172 , R140_U101 , U130 );
nand NAND2_152 ( U173 , P1_DATAO_REG_20_ , U127 );
nand NAND2_153 ( U174 , R140_U102 , U130 );
nand NAND2_154 ( U175 , P1_DATAO_REG_1_ , U127 );
nand NAND2_155 ( U176 , R140_U10 , U130 );
nand NAND2_156 ( U177 , P1_DATAO_REG_19_ , U127 );
nand NAND2_157 ( U178 , R140_U103 , U130 );
nand NAND2_158 ( U179 , P1_DATAO_REG_18_ , U127 );
nand NAND2_159 ( U180 , R140_U104 , U130 );
nand NAND2_160 ( U181 , P1_DATAO_REG_17_ , U127 );
nand NAND2_161 ( U182 , R140_U105 , U130 );
nand NAND2_162 ( U183 , P1_DATAO_REG_16_ , U127 );
nand NAND2_163 ( U184 , R140_U106 , U130 );
nand NAND2_164 ( U185 , P1_DATAO_REG_15_ , U127 );
nand NAND2_165 ( U186 , R140_U107 , U130 );
nand NAND2_166 ( U187 , P1_DATAO_REG_14_ , U127 );
nand NAND2_167 ( U188 , R140_U108 , U130 );
nand NAND2_168 ( U189 , P1_DATAO_REG_13_ , U127 );
nand NAND2_169 ( U190 , R140_U109 , U130 );
nand NAND2_170 ( U191 , P1_DATAO_REG_12_ , U127 );
nand NAND2_171 ( U192 , R140_U110 , U130 );
nand NAND2_172 ( U193 , P1_DATAO_REG_11_ , U127 );
nand NAND2_173 ( U194 , R140_U111 , U130 );
nand NAND2_174 ( U195 , P1_DATAO_REG_10_ , U127 );
nand NAND2_175 ( U196 , R140_U112 , U130 );
nand NAND2_176 ( U197 , P1_DATAO_REG_0_ , U127 );
nand NAND2_177 ( U198 , R140_U83 , U130 );
nand NAND2_178 ( U199 , R140_U84 , U127 );
nand NAND2_179 ( U200 , P2_DATAO_REG_9_ , U130 );
nand NAND2_180 ( U201 , R140_U85 , U127 );
nand NAND2_181 ( U202 , P2_DATAO_REG_8_ , U130 );
nand NAND2_182 ( U203 , R140_U86 , U127 );
nand NAND2_183 ( U204 , P2_DATAO_REG_7_ , U130 );
nand NAND2_184 ( U205 , R140_U87 , U127 );
nand NAND2_185 ( U206 , P2_DATAO_REG_6_ , U130 );
nand NAND2_186 ( U207 , R140_U88 , U127 );
nand NAND2_187 ( U208 , P2_DATAO_REG_5_ , U130 );
nand NAND2_188 ( U209 , R140_U89 , U127 );
nand NAND2_189 ( U210 , P2_DATAO_REG_4_ , U130 );
nand NAND2_190 ( U211 , R140_U90 , U127 );
nand NAND2_191 ( U212 , P2_DATAO_REG_3_ , U130 );
nand NAND2_192 ( U213 , R140_U11 , U127 );
nand NAND2_193 ( U214 , P2_DATAO_REG_31_ , U130 );
nand NAND2_194 ( U215 , R140_U91 , U127 );
nand NAND2_195 ( U216 , P2_DATAO_REG_30_ , U130 );
nand NAND2_196 ( U217 , R140_U92 , U127 );
nand NAND2_197 ( U218 , P2_DATAO_REG_2_ , U130 );
nand NAND2_198 ( U219 , R140_U93 , U127 );
nand NAND2_199 ( U220 , P2_DATAO_REG_29_ , U130 );
nand NAND2_200 ( U221 , R140_U94 , U127 );
nand NAND2_201 ( U222 , P2_DATAO_REG_28_ , U130 );
nand NAND2_202 ( U223 , R140_U95 , U127 );
nand NAND2_203 ( U224 , P2_DATAO_REG_27_ , U130 );
nand NAND2_204 ( U225 , R140_U96 , U127 );
nand NAND2_205 ( U226 , P2_DATAO_REG_26_ , U130 );
nand NAND2_206 ( U227 , R140_U97 , U127 );
nand NAND2_207 ( U228 , P2_DATAO_REG_25_ , U130 );
nand NAND2_208 ( U229 , R140_U98 , U127 );
nand NAND2_209 ( U230 , P2_DATAO_REG_24_ , U130 );
nand NAND2_210 ( U231 , R140_U99 , U127 );
nand NAND2_211 ( U232 , P2_DATAO_REG_23_ , U130 );
nand NAND2_212 ( U233 , R140_U100 , U127 );
nand NAND2_213 ( U234 , P2_DATAO_REG_22_ , U130 );
nand NAND2_214 ( U235 , R140_U101 , U127 );
nand NAND2_215 ( U236 , P2_DATAO_REG_21_ , U130 );
nand NAND2_216 ( U237 , R140_U102 , U127 );
nand NAND2_217 ( U238 , P2_DATAO_REG_20_ , U130 );
nand NAND2_218 ( U239 , R140_U10 , U127 );
nand NAND2_219 ( U240 , P2_DATAO_REG_1_ , U130 );
nand NAND2_220 ( U241 , R140_U103 , U127 );
nand NAND2_221 ( U242 , P2_DATAO_REG_19_ , U130 );
nand NAND2_222 ( U243 , R140_U104 , U127 );
nand NAND2_223 ( U244 , P2_DATAO_REG_18_ , U130 );
nand NAND2_224 ( U245 , R140_U105 , U127 );
nand NAND2_225 ( U246 , P2_DATAO_REG_17_ , U130 );
nand NAND2_226 ( U247 , R140_U106 , U127 );
nand NAND2_227 ( U248 , P2_DATAO_REG_16_ , U130 );
nand NAND2_228 ( U249 , R140_U107 , U127 );
nand NAND2_229 ( U250 , P2_DATAO_REG_15_ , U130 );
nand NAND2_230 ( U251 , R140_U108 , U127 );
nand NAND2_231 ( U252 , P2_DATAO_REG_14_ , U130 );
nand NAND2_232 ( U253 , R140_U109 , U127 );
nand NAND2_233 ( U254 , P2_DATAO_REG_13_ , U130 );
nand NAND2_234 ( U255 , R140_U110 , U127 );
nand NAND2_235 ( U256 , P2_DATAO_REG_12_ , U130 );
nand NAND2_236 ( U257 , R140_U111 , U127 );
nand NAND2_237 ( U258 , P2_DATAO_REG_11_ , U130 );
nand NAND2_238 ( U259 , R140_U112 , U127 );
nand NAND2_239 ( U260 , P2_DATAO_REG_10_ , U130 );
nand NAND2_240 ( U261 , R140_U83 , U127 );
nand NAND2_241 ( U262 , P2_DATAO_REG_0_ , U130 );
nand NAND2_242 ( U263 , P2_DATAO_REG_9_ , U127 );
nand NAND2_243 ( U264 , U130 , P1_DATAO_REG_9_ );
nand NAND2_244 ( U265 , P2_DATAO_REG_8_ , U127 );
nand NAND2_245 ( U266 , P1_DATAO_REG_8_ , U130 );
nand NAND2_246 ( U267 , P2_DATAO_REG_7_ , U127 );
nand NAND2_247 ( U268 , P1_DATAO_REG_7_ , U130 );
nand NAND2_248 ( U269 , P2_DATAO_REG_6_ , U127 );
nand NAND2_249 ( U270 , P1_DATAO_REG_6_ , U130 );
nand NAND2_250 ( U271 , P2_DATAO_REG_5_ , U127 );
nand NAND2_251 ( U272 , P1_DATAO_REG_5_ , U130 );
nand NAND2_252 ( U273 , P2_DATAO_REG_4_ , U127 );
nand NAND2_253 ( U274 , P1_DATAO_REG_4_ , U130 );
nand NAND2_254 ( U275 , P2_DATAO_REG_31_ , U127 );
nand NAND2_255 ( U276 , P1_DATAO_REG_31_ , U130 );
nand NAND2_256 ( U277 , P2_DATAO_REG_30_ , U127 );
nand NAND2_257 ( U278 , P1_DATAO_REG_30_ , U130 );
nand NAND2_258 ( U279 , P2_DATAO_REG_3_ , U127 );
nand NAND2_259 ( U280 , P1_DATAO_REG_3_ , U130 );
nand NAND2_260 ( U281 , P2_DATAO_REG_29_ , U127 );
nand NAND2_261 ( U282 , P1_DATAO_REG_29_ , U130 );
nand NAND2_262 ( U283 , P2_DATAO_REG_28_ , U127 );
nand NAND2_263 ( U284 , P1_DATAO_REG_28_ , U130 );
nand NAND2_264 ( U285 , P2_DATAO_REG_27_ , U127 );
nand NAND2_265 ( U286 , P1_DATAO_REG_27_ , U130 );
nand NAND2_266 ( U287 , P2_DATAO_REG_26_ , U127 );
nand NAND2_267 ( U288 , P1_DATAO_REG_26_ , U130 );
nand NAND2_268 ( U289 , P2_DATAO_REG_25_ , U127 );
nand NAND2_269 ( U290 , P1_DATAO_REG_25_ , U130 );
nand NAND2_270 ( U291 , P2_DATAO_REG_24_ , U127 );
nand NAND2_271 ( U292 , P1_DATAO_REG_24_ , U130 );
nand NAND2_272 ( U293 , P2_DATAO_REG_23_ , U127 );
nand NAND2_273 ( U294 , P1_DATAO_REG_23_ , U130 );
nand NAND2_274 ( U295 , P2_DATAO_REG_22_ , U127 );
nand NAND2_275 ( U296 , P1_DATAO_REG_22_ , U130 );
nand NAND2_276 ( U297 , P2_DATAO_REG_21_ , U127 );
nand NAND2_277 ( U298 , P1_DATAO_REG_21_ , U130 );
nand NAND2_278 ( U299 , P2_DATAO_REG_20_ , U127 );
nand NAND2_279 ( U300 , P1_DATAO_REG_20_ , U130 );
nand NAND2_280 ( U301 , P2_DATAO_REG_2_ , U127 );
nand NAND2_281 ( U302 , P1_DATAO_REG_2_ , U130 );
nand NAND2_282 ( U303 , P2_DATAO_REG_19_ , U127 );
nand NAND2_283 ( U304 , P1_DATAO_REG_19_ , U130 );
nand NAND2_284 ( U305 , P2_DATAO_REG_18_ , U127 );
nand NAND2_285 ( U306 , P1_DATAO_REG_18_ , U130 );
nand NAND2_286 ( U307 , P2_DATAO_REG_17_ , U127 );
nand NAND2_287 ( U308 , P1_DATAO_REG_17_ , U130 );
nand NAND2_288 ( U309 , P2_DATAO_REG_16_ , U127 );
nand NAND2_289 ( U310 , P1_DATAO_REG_16_ , U130 );
nand NAND2_290 ( U311 , P2_DATAO_REG_15_ , U127 );
nand NAND2_291 ( U312 , P1_DATAO_REG_15_ , U130 );
nand NAND2_292 ( U313 , P2_DATAO_REG_14_ , U127 );
nand NAND2_293 ( U314 , P1_DATAO_REG_14_ , U130 );
nand NAND2_294 ( U315 , P2_DATAO_REG_13_ , U127 );
nand NAND2_295 ( U316 , P1_DATAO_REG_13_ , U130 );
nand NAND2_296 ( U317 , P2_DATAO_REG_12_ , U127 );
nand NAND2_297 ( U318 , P1_DATAO_REG_12_ , U130 );
nand NAND2_298 ( U319 , P2_DATAO_REG_11_ , U127 );
nand NAND2_299 ( U320 , P1_DATAO_REG_11_ , U130 );
nand NAND2_300 ( U321 , P2_DATAO_REG_10_ , U127 );
nand NAND2_301 ( U322 , P1_DATAO_REG_10_ , U130 );
nand NAND2_302 ( U323 , P2_DATAO_REG_1_ , U127 );
nand NAND2_303 ( U324 , P1_DATAO_REG_1_ , U130 );
nand NAND2_304 ( U325 , P2_DATAO_REG_0_ , U127 );
nand NAND2_305 ( U326 , P1_DATAO_REG_0_ , U130 );
nand NAND2_306 ( P2_R1161_U501 , P2_U3061 , P2_R1161_U63 );
nand NAND2_307 ( P2_R1161_U500 , P2_R1161_U244 , P2_R1161_U498 );
nand NAND2_308 ( P2_R1161_U499 , P2_R1161_U363 , P2_R1161_U167 );
nand NAND2_309 ( P2_R1161_U498 , P2_R1161_U497 , P2_R1161_U496 );
nand NAND2_310 ( P2_R1161_U497 , P2_U3422 , P2_R1161_U67 );
nand NAND2_311 ( P2_R1161_U496 , P2_U3062 , P2_R1161_U66 );
nand NAND2_312 ( P2_R1161_U495 , P2_R1161_U493 , P2_R1161_U338 );
nand NAND2_313 ( P2_R1161_U494 , P2_R1161_U362 , P2_R1161_U93 );
nand NAND2_314 ( P2_R1161_U493 , P2_R1161_U492 , P2_R1161_U491 );
nand NAND2_315 ( P2_R1161_U492 , P2_U3425 , P2_R1161_U70 );
nand NAND2_316 ( P2_R1161_U491 , P2_U3071 , P2_R1161_U69 );
nand NAND2_317 ( P2_R1161_U490 , P2_U3428 , P2_R1161_U62 );
and AND2_318 ( P1_U3014 , P1_U3956 , P1_U3443 );
and AND2_319 ( P1_U3015 , P1_U3449 , P1_U3446 );
and AND2_320 ( P1_U3016 , P1_U3630 , P1_U3625 );
and AND2_321 ( P1_U3017 , P1_U3444 , P1_U3445 );
and AND2_322 ( P1_U3018 , P1_U5711 , P1_U3444 );
and AND2_323 ( P1_U3019 , P1_U5708 , P1_U3445 );
and AND2_324 ( P1_U3020 , P1_U5708 , P1_U5711 );
and AND2_325 ( P1_U3021 , P1_U5368 , P1_U3421 );
and AND2_326 ( P1_U3022 , P1_U3046 , P1_STATE_REG );
and AND2_327 ( P1_U3023 , P1_U3049 , P1_U5690 );
and AND2_328 ( P1_U3024 , P1_U3807 , P1_U3423 );
and AND2_329 ( P1_U3025 , P1_U3987 , P1_U5699 );
and AND2_330 ( P1_U3026 , P1_U3953 , P1_U5690 );
and AND2_331 ( P1_U3027 , P1_U3871 , P1_U3972 );
and AND2_332 ( P1_U3028 , P1_U3357 , P1_STATE_REG );
and AND2_333 ( P1_U3029 , P1_U3964 , P1_U3989 );
and AND2_334 ( P1_U3030 , P1_U3989 , P1_U3422 );
and AND2_335 ( P1_U3031 , P1_U3957 , P1_U3989 );
and AND2_336 ( P1_U3032 , P1_U3965 , P1_U3989 );
and AND2_337 ( P1_U3033 , P1_U3987 , P1_U3446 );
and AND2_338 ( P1_U3034 , P1_U3972 , P1_U5699 );
and AND2_339 ( P1_U3035 , P1_U3989 , P1_U3025 );
and AND2_340 ( P1_U3036 , P1_U3972 , P1_U3446 );
and AND2_341 ( P1_U3037 , P1_U5702 , P1_U4880 );
and AND2_342 ( P1_U3038 , P1_U3024 , P1_U5702 );
and AND2_343 ( P1_U3039 , P1_U5699 , P1_U4880 );
and AND2_344 ( P1_U3040 , P1_U3024 , P1_U5699 );
and AND2_345 ( P1_U3041 , P1_U3015 , P1_U4880 );
and AND2_346 ( P1_U3042 , P1_U3024 , P1_U3015 );
and AND2_347 ( P1_U3043 , P1_U3022 , P1_U3423 );
and AND2_348 ( P1_U3044 , P1_U5113 , P1_STATE_REG );
and AND2_349 ( P1_U3045 , P1_U3022 , P1_U5115 );
and AND2_350 ( P1_U3046 , P1_U5677 , P1_U3421 );
and AND2_351 ( P1_U3047 , P1_U3631 , P1_U3016 );
and AND2_352 ( P1_U3048 , P1_U5690 , P1_U3442 );
and AND2_353 ( P1_U3049 , P1_U5684 , P1_U5693 );
and AND2_354 ( P1_U3050 , P1_U3435 , P1_U3437 );
and AND4_355 ( P1_U3051 , P1_U4706 , P1_U4703 , P1_U4700 , P1_U4699 );
and AND2_356 ( P1_U3052 , P1_U6070 , P1_U6069 );
nand NAND4_357 ( P1_U3053 , P1_U4637 , P1_U4638 , P1_U4636 , P1_U4639 );
nand NAND4_358 ( P1_U3054 , P1_U4656 , P1_U4657 , P1_U4655 , P1_U4658 );
nand NAND4_359 ( P1_U3055 , P1_U4677 , P1_U4676 , P1_U4675 , P1_U4674 );
nand NAND3_360 ( P1_U3056 , P1_U4714 , P1_U4715 , P1_U4713 );
nand NAND4_361 ( P1_U3057 , P1_U4618 , P1_U4619 , P1_U4617 , P1_U4620 );
nand NAND4_362 ( P1_U3058 , P1_U4599 , P1_U4600 , P1_U4598 , P1_U4601 );
nand NAND3_363 ( P1_U3059 , P1_U4694 , P1_U4695 , P1_U4693 );
nand NAND4_364 ( P1_U3060 , P1_U4202 , P1_U4201 , P1_U4200 , P1_U4199 );
nand NAND4_365 ( P1_U3061 , P1_U4542 , P1_U4543 , P1_U4541 , P1_U4544 );
nand NAND4_366 ( P1_U3062 , P1_U4314 , P1_U4315 , P1_U4313 , P1_U4316 );
nand NAND4_367 ( P1_U3063 , P1_U4333 , P1_U4334 , P1_U4332 , P1_U4335 );
nand NAND4_368 ( P1_U3064 , P1_U4183 , P1_U4182 , P1_U4181 , P1_U4180 );
nand NAND4_369 ( P1_U3065 , P1_U4580 , P1_U4581 , P1_U4579 , P1_U4582 );
nand NAND4_370 ( P1_U3066 , P1_U4561 , P1_U4562 , P1_U4560 , P1_U4563 );
nand NAND4_371 ( P1_U3067 , P1_U4221 , P1_U4220 , P1_U4219 , P1_U4218 );
nand NAND4_372 ( P1_U3068 , P1_U4159 , P1_U4158 , P1_U4157 , P1_U4156 );
nand NAND4_373 ( P1_U3069 , P1_U4447 , P1_U4448 , P1_U4446 , P1_U4449 );
nand NAND4_374 ( P1_U3070 , P1_U4259 , P1_U4258 , P1_U4257 , P1_U4256 );
nand NAND4_375 ( P1_U3071 , P1_U4240 , P1_U4239 , P1_U4238 , P1_U4237 );
nand NAND4_376 ( P1_U3072 , P1_U4352 , P1_U4353 , P1_U4351 , P1_U4354 );
nand NAND4_377 ( P1_U3073 , P1_U4428 , P1_U4429 , P1_U4427 , P1_U4430 );
nand NAND4_378 ( P1_U3074 , P1_U4409 , P1_U4410 , P1_U4408 , P1_U4411 );
nand NAND4_379 ( P1_U3075 , P1_U4523 , P1_U4524 , P1_U4522 , P1_U4525 );
nand NAND4_380 ( P1_U3076 , P1_U4504 , P1_U4505 , P1_U4503 , P1_U4506 );
nand NAND4_381 ( P1_U3077 , P1_U4164 , P1_U4163 , P1_U4162 , P1_U4161 );
nand NAND4_382 ( P1_U3078 , P1_U4140 , P1_U4139 , P1_U4138 , P1_U4137 );
nand NAND4_383 ( P1_U3079 , P1_U4390 , P1_U4391 , P1_U4389 , P1_U4392 );
nand NAND4_384 ( P1_U3080 , P1_U4371 , P1_U4372 , P1_U4370 , P1_U4373 );
nand NAND4_385 ( P1_U3081 , P1_U4485 , P1_U4486 , P1_U4484 , P1_U4487 );
nand NAND4_386 ( P1_U3082 , P1_U4466 , P1_U4467 , P1_U4465 , P1_U4468 );
nand NAND4_387 ( P1_U3083 , P1_U4295 , P1_U4296 , P1_U4294 , P1_U4297 );
nand NAND4_388 ( P1_U3084 , P1_U4278 , P1_U4277 , P1_U4276 , P1_U4275 );
nand NAND2_389 ( P1_U3085 , P1_U4887 , P1_STATE_REG );
not NOT1_390 ( P1_U3086 , P1_STATE_REG );
nand NAND2_391 ( P1_U3087 , P1_U5576 , P1_U5575 );
nand NAND2_392 ( P1_U3088 , P1_U5578 , P1_U5577 );
nand NAND3_393 ( P1_U3089 , P1_U5583 , P1_U5584 , P1_U5582 );
nand NAND2_394 ( P1_U3090 , P1_U3895 , P1_U5586 );
nand NAND2_395 ( P1_U3091 , P1_U3896 , P1_U5589 );
nand NAND2_396 ( P1_U3092 , P1_U3897 , P1_U5592 );
nand NAND2_397 ( P1_U3093 , P1_U3898 , P1_U5595 );
nand NAND2_398 ( P1_U3094 , P1_U3899 , P1_U5598 );
nand NAND2_399 ( P1_U3095 , P1_U3900 , P1_U5601 );
nand NAND2_400 ( P1_U3096 , P1_U3901 , P1_U5604 );
nand NAND2_401 ( P1_U3097 , P1_U3902 , P1_U5607 );
nand NAND2_402 ( P1_U3098 , P1_U3903 , P1_U5610 );
nand NAND2_403 ( P1_U3099 , P1_U3904 , P1_U5616 );
nand NAND2_404 ( P1_U3100 , P1_U3905 , P1_U5619 );
nand NAND2_405 ( P1_U3101 , P1_U3906 , P1_U5622 );
nand NAND2_406 ( P1_U3102 , P1_U3907 , P1_U5625 );
nand NAND2_407 ( P1_U3103 , P1_U3908 , P1_U5628 );
nand NAND2_408 ( P1_U3104 , P1_U3909 , P1_U5631 );
nand NAND3_409 ( P1_U3105 , P1_U5634 , P1_U5635 , P1_U5633 );
nand NAND3_410 ( P1_U3106 , P1_U5637 , P1_U5638 , P1_U5636 );
nand NAND3_411 ( P1_U3107 , P1_U5640 , P1_U5641 , P1_U5639 );
nand NAND3_412 ( P1_U3108 , P1_U5643 , P1_U5644 , P1_U5642 );
nand NAND3_413 ( P1_U3109 , P1_U5558 , P1_U5559 , P1_U5557 );
nand NAND3_414 ( P1_U3110 , P1_U5561 , P1_U5562 , P1_U5560 );
nand NAND3_415 ( P1_U3111 , P1_U5564 , P1_U5565 , P1_U5563 );
nand NAND3_416 ( P1_U3112 , P1_U5567 , P1_U5568 , P1_U5566 );
nand NAND3_417 ( P1_U3113 , P1_U5570 , P1_U5571 , P1_U5569 );
nand NAND3_418 ( P1_U3114 , P1_U5573 , P1_U5574 , P1_U5572 );
nand NAND3_419 ( P1_U3115 , P1_U5580 , P1_U5581 , P1_U5579 );
nand NAND3_420 ( P1_U3116 , P1_U5613 , P1_U5614 , P1_U5612 );
nand NAND3_421 ( P1_U3117 , P1_U5646 , P1_U5647 , P1_U5645 );
nand NAND2_422 ( P1_U3118 , P1_U5649 , P1_U5648 );
nand NAND2_423 ( P1_U3119 , P1_U5506 , P1_U5505 );
nand NAND2_424 ( P1_U3120 , P1_U5508 , P1_U5507 );
nand NAND3_425 ( P1_U3121 , P1_U3438 , P1_U5511 , P1_U5512 );
nand NAND2_426 ( P1_U3122 , P1_U3879 , P1_U5513 );
nand NAND2_427 ( P1_U3123 , P1_U3880 , P1_U5515 );
nand NAND2_428 ( P1_U3124 , P1_U3881 , P1_U5517 );
nand NAND2_429 ( P1_U3125 , P1_U3882 , P1_U5519 );
nand NAND2_430 ( P1_U3126 , P1_U3883 , P1_U5521 );
nand NAND2_431 ( P1_U3127 , P1_U3884 , P1_U5523 );
nand NAND2_432 ( P1_U3128 , P1_U3885 , P1_U5525 );
nand NAND2_433 ( P1_U3129 , P1_U3886 , P1_U5527 );
nand NAND2_434 ( P1_U3130 , P1_U3887 , P1_U5529 );
nand NAND2_435 ( P1_U3131 , P1_U3888 , P1_U5534 );
nand NAND2_436 ( P1_U3132 , P1_U3889 , P1_U5536 );
nand NAND2_437 ( P1_U3133 , P1_U3890 , P1_U5538 );
nand NAND2_438 ( P1_U3134 , P1_U3891 , P1_U5540 );
nand NAND2_439 ( P1_U3135 , P1_U3892 , P1_U5542 );
nand NAND2_440 ( P1_U3136 , P1_U3893 , P1_U5544 );
nand NAND3_441 ( P1_U3137 , P1_U5546 , P1_U3438 , P1_U5545 );
nand NAND3_442 ( P1_U3138 , P1_U5548 , P1_U3438 , P1_U5547 );
nand NAND3_443 ( P1_U3139 , P1_U5550 , P1_U3438 , P1_U5549 );
nand NAND3_444 ( P1_U3140 , P1_U5552 , P1_U3438 , P1_U5551 );
nand NAND3_445 ( P1_U3141 , P1_U5494 , P1_U3438 , P1_U5493 );
nand NAND3_446 ( P1_U3142 , P1_U5496 , P1_U3438 , P1_U5495 );
nand NAND3_447 ( P1_U3143 , P1_U5498 , P1_U3438 , P1_U5497 );
nand NAND3_448 ( P1_U3144 , P1_U5500 , P1_U3438 , P1_U5499 );
nand NAND3_449 ( P1_U3145 , P1_U5502 , P1_U3438 , P1_U5501 );
nand NAND3_450 ( P1_U3146 , P1_U5504 , P1_U3438 , P1_U5503 );
nand NAND3_451 ( P1_U3147 , P1_U5510 , P1_U3438 , P1_U5509 );
nand NAND3_452 ( P1_U3148 , P1_U5532 , P1_U3438 , P1_U5531 );
nand NAND3_453 ( P1_U3149 , P1_U5554 , P1_U3438 , P1_U5553 );
nand NAND2_454 ( P1_U3150 , P1_U3894 , P1_U5556 );
nand NAND2_455 ( P1_U3151 , P1_U3953 , P1_U3438 );
nand NAND2_456 ( P1_U3152 , P1_U5677 , P1_U3372 );
nand NAND2_457 ( P1_U3153 , P1_U5448 , P1_U5447 );
nand NAND2_458 ( P1_U3154 , P1_U5450 , P1_U5449 );
nand NAND2_459 ( P1_U3155 , P1_U5452 , P1_U5451 );
nand NAND2_460 ( P1_U3156 , P1_U5454 , P1_U5453 );
nand NAND2_461 ( P1_U3157 , P1_U5456 , P1_U5455 );
nand NAND2_462 ( P1_U3158 , P1_U5458 , P1_U5457 );
nand NAND2_463 ( P1_U3159 , P1_U5460 , P1_U5459 );
nand NAND2_464 ( P1_U3160 , P1_U5462 , P1_U5461 );
nand NAND2_465 ( P1_U3161 , P1_U5464 , P1_U5463 );
nand NAND2_466 ( P1_U3162 , P1_U5468 , P1_U5467 );
nand NAND2_467 ( P1_U3163 , P1_U5470 , P1_U5469 );
nand NAND2_468 ( P1_U3164 , P1_U5472 , P1_U5471 );
nand NAND2_469 ( P1_U3165 , P1_U5474 , P1_U5473 );
nand NAND2_470 ( P1_U3166 , P1_U5476 , P1_U5475 );
nand NAND2_471 ( P1_U3167 , P1_U5478 , P1_U5477 );
nand NAND2_472 ( P1_U3168 , P1_U5480 , P1_U5479 );
nand NAND2_473 ( P1_U3169 , P1_U5482 , P1_U5481 );
nand NAND2_474 ( P1_U3170 , P1_U5484 , P1_U5483 );
nand NAND2_475 ( P1_U3171 , P1_U5486 , P1_U5485 );
nand NAND2_476 ( P1_U3172 , P1_U5434 , P1_U5433 );
nand NAND2_477 ( P1_U3173 , P1_U5436 , P1_U5435 );
nand NAND2_478 ( P1_U3174 , P1_U5438 , P1_U5437 );
nand NAND2_479 ( P1_U3175 , P1_U5440 , P1_U5439 );
nand NAND2_480 ( P1_U3176 , P1_U5442 , P1_U5441 );
nand NAND2_481 ( P1_U3177 , P1_U5444 , P1_U5443 );
nand NAND2_482 ( P1_U3178 , P1_U5446 , P1_U5445 );
nand NAND2_483 ( P1_U3179 , P1_U5466 , P1_U5465 );
nand NAND2_484 ( P1_U3180 , P1_U5488 , P1_U5487 );
nand NAND3_485 ( P1_U3181 , P1_U5490 , P1_U5491 , P1_U5489 );
nand NAND2_486 ( P1_U3182 , P1_U5389 , P1_U5388 );
nand NAND2_487 ( P1_U3183 , P1_U5391 , P1_U5390 );
nand NAND2_488 ( P1_U3184 , P1_U5393 , P1_U5392 );
nand NAND2_489 ( P1_U3185 , P1_U5395 , P1_U5394 );
nand NAND2_490 ( P1_U3186 , P1_U5397 , P1_U5396 );
nand NAND2_491 ( P1_U3187 , P1_U5399 , P1_U5398 );
nand NAND2_492 ( P1_U3188 , P1_U5401 , P1_U5400 );
nand NAND2_493 ( P1_U3189 , P1_U5403 , P1_U5402 );
nand NAND2_494 ( P1_U3190 , P1_U5405 , P1_U5404 );
nand NAND2_495 ( P1_U3191 , P1_U5409 , P1_U5408 );
nand NAND2_496 ( P1_U3192 , P1_U5411 , P1_U5410 );
nand NAND2_497 ( P1_U3193 , P1_U5413 , P1_U5412 );
nand NAND2_498 ( P1_U3194 , P1_U5415 , P1_U5414 );
nand NAND2_499 ( P1_U3195 , P1_U5417 , P1_U5416 );
nand NAND2_500 ( P1_U3196 , P1_U5419 , P1_U5418 );
nand NAND2_501 ( P1_U3197 , P1_U5421 , P1_U5420 );
nand NAND2_502 ( P1_U3198 , P1_U5423 , P1_U5422 );
nand NAND2_503 ( P1_U3199 , P1_U5425 , P1_U5424 );
nand NAND2_504 ( P1_U3200 , P1_U5427 , P1_U5426 );
nand NAND2_505 ( P1_U3201 , P1_U5375 , P1_U5374 );
nand NAND2_506 ( P1_U3202 , P1_U5377 , P1_U5376 );
nand NAND2_507 ( P1_U3203 , P1_U5379 , P1_U5378 );
nand NAND2_508 ( P1_U3204 , P1_U5381 , P1_U5380 );
nand NAND2_509 ( P1_U3205 , P1_U5383 , P1_U5382 );
nand NAND2_510 ( P1_U3206 , P1_U5385 , P1_U5384 );
nand NAND2_511 ( P1_U3207 , P1_U5387 , P1_U5386 );
nand NAND2_512 ( P1_U3208 , P1_U5407 , P1_U5406 );
nand NAND2_513 ( P1_U3209 , P1_U5429 , P1_U5428 );
nand NAND2_514 ( P1_U3210 , P1_U3878 , P1_U5430 );
and AND2_515 ( P1_U3211 , P1_U5367 , P1_U3421 );
nand NAND3_516 ( P1_U3212 , P1_U6236 , P1_U6235 , P1_U5365 );
nand NAND5_517 ( P1_U3213 , P1_U5359 , P1_U5358 , P1_U5362 , P1_U5360 , P1_U5361 );
nand NAND5_518 ( P1_U3214 , P1_U5350 , P1_U5349 , P1_U5353 , P1_U5351 , P1_U5352 );
nand NAND5_519 ( P1_U3215 , P1_U5341 , P1_U5340 , P1_U5344 , P1_U5342 , P1_U5343 );
nand NAND5_520 ( P1_U3216 , P1_U5332 , P1_U5331 , P1_U5335 , P1_U5333 , P1_U5334 );
nand NAND5_521 ( P1_U3217 , P1_U5323 , P1_U5322 , P1_U5326 , P1_U5324 , P1_U5325 );
nand NAND5_522 ( P1_U3218 , P1_U5314 , P1_U5313 , P1_U5317 , P1_U5315 , P1_U5316 );
nand NAND5_523 ( P1_U3219 , P1_U5305 , P1_U5304 , P1_U5308 , P1_U5306 , P1_U5307 );
nand NAND5_524 ( P1_U3220 , P1_U5296 , P1_U5295 , P1_U5299 , P1_U5297 , P1_U5298 );
nand NAND5_525 ( P1_U3221 , P1_U5287 , P1_U5286 , P1_U5290 , P1_U5288 , P1_U5289 );
nand NAND4_526 ( P1_U3222 , P1_U5278 , P1_U5277 , P1_U3876 , P1_U5279 );
nand NAND5_527 ( P1_U3223 , P1_U5269 , P1_U5268 , P1_U5272 , P1_U5270 , P1_U5271 );
nand NAND5_528 ( P1_U3224 , P1_U5260 , P1_U5259 , P1_U5263 , P1_U5261 , P1_U5262 );
nand NAND5_529 ( P1_U3225 , P1_U5251 , P1_U5250 , P1_U5254 , P1_U5252 , P1_U5253 );
nand NAND5_530 ( P1_U3226 , P1_U5242 , P1_U5241 , P1_U5245 , P1_U5243 , P1_U5244 );
nand NAND5_531 ( P1_U3227 , P1_U5233 , P1_U5232 , P1_U5236 , P1_U5234 , P1_U5235 );
nand NAND5_532 ( P1_U3228 , P1_U5224 , P1_U5223 , P1_U5227 , P1_U5225 , P1_U5226 );
nand NAND5_533 ( P1_U3229 , P1_U5215 , P1_U5214 , P1_U5218 , P1_U5216 , P1_U5217 );
nand NAND5_534 ( P1_U3230 , P1_U5206 , P1_U5205 , P1_U5209 , P1_U5207 , P1_U5208 );
nand NAND5_535 ( P1_U3231 , P1_U5197 , P1_U5196 , P1_U5200 , P1_U5198 , P1_U5199 );
nand NAND3_536 ( P1_U3232 , P1_U3875 , P1_U5189 , P1_U3874 );
nand NAND5_537 ( P1_U3233 , P1_U5180 , P1_U5179 , P1_U5183 , P1_U5181 , P1_U5182 );
nand NAND5_538 ( P1_U3234 , P1_U5171 , P1_U5170 , P1_U5174 , P1_U5172 , P1_U5173 );
nand NAND5_539 ( P1_U3235 , P1_U5162 , P1_U5161 , P1_U5165 , P1_U5163 , P1_U5164 );
nand NAND5_540 ( P1_U3236 , P1_U5153 , P1_U5152 , P1_U5156 , P1_U5154 , P1_U5155 );
nand NAND4_541 ( P1_U3237 , P1_U5144 , P1_U5143 , P1_U5145 , P1_U3872 );
nand NAND5_542 ( P1_U3238 , P1_U5135 , P1_U5134 , P1_U5138 , P1_U5136 , P1_U5137 );
nand NAND5_543 ( P1_U3239 , P1_U5126 , P1_U5125 , P1_U5129 , P1_U5127 , P1_U5128 );
nand NAND5_544 ( P1_U3240 , P1_U5117 , P1_U5116 , P1_U5120 , P1_U5118 , P1_U5119 );
nand NAND5_545 ( P1_U3241 , P1_U5104 , P1_U5103 , P1_U5107 , P1_U5105 , P1_U5106 );
and AND2_546 ( P1_U3242 , P1_U3866 , P1_U5650 );
nand NAND2_547 ( P1_U3243 , P1_U3849 , P1_U3848 );
nand NAND2_548 ( P1_U3244 , P1_U3847 , P1_U3846 );
nand NAND2_549 ( P1_U3245 , P1_U3845 , P1_U3844 );
nand NAND2_550 ( P1_U3246 , P1_U3842 , P1_U3841 );
nand NAND2_551 ( P1_U3247 , P1_U3840 , P1_U3839 );
nand NAND2_552 ( P1_U3248 , P1_U3837 , P1_U3836 );
nand NAND2_553 ( P1_U3249 , P1_U3835 , P1_U3834 );
nand NAND3_554 ( P1_U3250 , P1_U3832 , P1_U3833 , P1_U5010 );
nand NAND3_555 ( P1_U3251 , P1_U3830 , P1_U3831 , P1_U5000 );
nand NAND3_556 ( P1_U3252 , P1_U3828 , P1_U3829 , P1_U4990 );
nand NAND3_557 ( P1_U3253 , P1_U3826 , P1_U3827 , P1_U4980 );
nand NAND3_558 ( P1_U3254 , P1_U3824 , P1_U3825 , P1_U4970 );
nand NAND3_559 ( P1_U3255 , P1_U3822 , P1_U3823 , P1_U4960 );
nand NAND3_560 ( P1_U3256 , P1_U3820 , P1_U3821 , P1_U4950 );
nand NAND3_561 ( P1_U3257 , P1_U3818 , P1_U3819 , P1_U4940 );
nand NAND3_562 ( P1_U3258 , P1_U3816 , P1_U3817 , P1_U4930 );
nand NAND3_563 ( P1_U3259 , P1_U3814 , P1_U3815 , P1_U4920 );
nand NAND3_564 ( P1_U3260 , P1_U3812 , P1_U3813 , P1_U4910 );
nand NAND3_565 ( P1_U3261 , P1_U3810 , P1_U3811 , P1_U4900 );
nand NAND3_566 ( P1_U3262 , P1_U3808 , P1_U3809 , P1_U4890 );
nand NAND3_567 ( P1_U3263 , P1_U3947 , P1_U4878 , P1_U4879 );
nand NAND3_568 ( P1_U3264 , P1_U3946 , P1_U4876 , P1_U4877 );
nand NAND4_569 ( P1_U3265 , P1_U3799 , P1_U3800 , P1_U4869 , P1_U3943 );
nand NAND4_570 ( P1_U3266 , P1_U3797 , P1_U3798 , P1_U4864 , P1_U3942 );
nand NAND4_571 ( P1_U3267 , P1_U3795 , P1_U3796 , P1_U4859 , P1_U3941 );
nand NAND4_572 ( P1_U3268 , P1_U3793 , P1_U3794 , P1_U4854 , P1_U3940 );
nand NAND4_573 ( P1_U3269 , P1_U3791 , P1_U3792 , P1_U4849 , P1_U3939 );
nand NAND3_574 ( P1_U3270 , P1_U3790 , P1_U3789 , P1_U3938 );
nand NAND3_575 ( P1_U3271 , P1_U3788 , P1_U3787 , P1_U3937 );
nand NAND2_576 ( P1_U3272 , P1_U3786 , P1_U3936 );
nand NAND3_577 ( P1_U3273 , P1_U3785 , P1_U3784 , P1_U3935 );
nand NAND2_578 ( P1_U3274 , P1_U3783 , P1_U3934 );
nand NAND2_579 ( P1_U3275 , P1_U3782 , P1_U3933 );
nand NAND2_580 ( P1_U3276 , P1_U3781 , P1_U3932 );
nand NAND2_581 ( P1_U3277 , P1_U3780 , P1_U3931 );
nand NAND2_582 ( P1_U3278 , P1_U3779 , P1_U3930 );
nand NAND2_583 ( P1_U3279 , P1_U3778 , P1_U3929 );
nand NAND3_584 ( P1_U3280 , P1_U3777 , P1_U3776 , P1_U3928 );
nand NAND3_585 ( P1_U3281 , P1_U3775 , P1_U3774 , P1_U3927 );
nand NAND3_586 ( P1_U3282 , P1_U3773 , P1_U3772 , P1_U3926 );
nand NAND4_587 ( P1_U3283 , P1_U3770 , P1_U3771 , P1_U4779 , P1_U3925 );
nand NAND4_588 ( P1_U3284 , P1_U3768 , P1_U3769 , P1_U4774 , P1_U3924 );
nand NAND4_589 ( P1_U3285 , P1_U3766 , P1_U3767 , P1_U4769 , P1_U3923 );
nand NAND4_590 ( P1_U3286 , P1_U3764 , P1_U3765 , P1_U4764 , P1_U3922 );
nand NAND4_591 ( P1_U3287 , P1_U3762 , P1_U3763 , P1_U4759 , P1_U3921 );
nand NAND4_592 ( P1_U3288 , P1_U3760 , P1_U3761 , P1_U4754 , P1_U3920 );
nand NAND4_593 ( P1_U3289 , P1_U3758 , P1_U3759 , P1_U4749 , P1_U3919 );
nand NAND3_594 ( P1_U3290 , P1_U3757 , P1_U3756 , P1_U3918 );
nand NAND2_595 ( P1_U3291 , P1_U3755 , P1_U3754 );
nand NAND2_596 ( P1_U3292 , P1_U3753 , P1_U3752 );
nand NAND2_597 ( P1_U3293 , P1_U3751 , P1_U3750 );
and AND2_598 ( P1_U3294 , P1_D_REG_31_ , P1_U3911 );
and AND2_599 ( P1_U3295 , P1_D_REG_30_ , P1_U3911 );
and AND2_600 ( P1_U3296 , P1_D_REG_29_ , P1_U3911 );
and AND2_601 ( P1_U3297 , P1_D_REG_28_ , P1_U3911 );
and AND2_602 ( P1_U3298 , P1_D_REG_27_ , P1_U3911 );
and AND2_603 ( P1_U3299 , P1_D_REG_26_ , P1_U3911 );
and AND2_604 ( P1_U3300 , P1_D_REG_25_ , P1_U3911 );
and AND2_605 ( P1_U3301 , P1_D_REG_24_ , P1_U3911 );
and AND2_606 ( P1_U3302 , P1_D_REG_23_ , P1_U3911 );
and AND2_607 ( P1_U3303 , P1_D_REG_22_ , P1_U3911 );
and AND2_608 ( P1_U3304 , P1_D_REG_21_ , P1_U3911 );
and AND2_609 ( P1_U3305 , P1_D_REG_20_ , P1_U3911 );
and AND2_610 ( P1_U3306 , P1_D_REG_19_ , P1_U3911 );
and AND2_611 ( P1_U3307 , P1_D_REG_18_ , P1_U3911 );
and AND2_612 ( P1_U3308 , P1_D_REG_17_ , P1_U3911 );
and AND2_613 ( P1_U3309 , P1_D_REG_16_ , P1_U3911 );
and AND2_614 ( P1_U3310 , P1_D_REG_15_ , P1_U3911 );
and AND2_615 ( P1_U3311 , P1_D_REG_14_ , P1_U3911 );
and AND2_616 ( P1_U3312 , P1_D_REG_13_ , P1_U3911 );
and AND2_617 ( P1_U3313 , P1_D_REG_12_ , P1_U3911 );
and AND2_618 ( P1_U3314 , P1_D_REG_11_ , P1_U3911 );
and AND2_619 ( P1_U3315 , P1_D_REG_10_ , P1_U3911 );
and AND2_620 ( P1_U3316 , P1_D_REG_9_ , P1_U3911 );
and AND2_621 ( P1_U3317 , P1_D_REG_8_ , P1_U3911 );
and AND2_622 ( P1_U3318 , P1_D_REG_7_ , P1_U3911 );
and AND2_623 ( P1_U3319 , P1_D_REG_6_ , P1_U3911 );
and AND2_624 ( P1_U3320 , P1_D_REG_5_ , P1_U3911 );
and AND2_625 ( P1_U3321 , P1_D_REG_4_ , P1_U3911 );
and AND2_626 ( P1_U3322 , P1_D_REG_3_ , P1_U3911 );
and AND2_627 ( P1_U3323 , P1_D_REG_2_ , P1_U3911 );
nand NAND3_628 ( P1_U3324 , P1_U4099 , P1_U4100 , P1_U4098 );
nand NAND3_629 ( P1_U3325 , P1_U4096 , P1_U4097 , P1_U4095 );
nand NAND3_630 ( P1_U3326 , P1_U4093 , P1_U4094 , P1_U4092 );
nand NAND3_631 ( P1_U3327 , P1_U4090 , P1_U4091 , P1_U4089 );
nand NAND3_632 ( P1_U3328 , P1_U4087 , P1_U4088 , P1_U4086 );
nand NAND3_633 ( P1_U3329 , P1_U4084 , P1_U4085 , P1_U4083 );
nand NAND3_634 ( P1_U3330 , P1_U4081 , P1_U4082 , P1_U4080 );
nand NAND3_635 ( P1_U3331 , P1_U4078 , P1_U4079 , P1_U4077 );
nand NAND3_636 ( P1_U3332 , P1_U4075 , P1_U4076 , P1_U4074 );
nand NAND3_637 ( P1_U3333 , P1_U4072 , P1_U4073 , P1_U4071 );
nand NAND3_638 ( P1_U3334 , P1_U4069 , P1_U4070 , P1_U4068 );
nand NAND3_639 ( P1_U3335 , P1_U4066 , P1_U4067 , P1_U4065 );
nand NAND3_640 ( P1_U3336 , P1_U4063 , P1_U4064 , P1_U4062 );
nand NAND3_641 ( P1_U3337 , P1_U4060 , P1_U4061 , P1_U4059 );
nand NAND3_642 ( P1_U3338 , P1_U4057 , P1_U4058 , P1_U4056 );
nand NAND3_643 ( P1_U3339 , P1_U4054 , P1_U4055 , P1_U4053 );
nand NAND3_644 ( P1_U3340 , P1_U4051 , P1_U4052 , P1_U4050 );
nand NAND3_645 ( P1_U3341 , P1_U4048 , P1_U4049 , P1_U4047 );
nand NAND3_646 ( P1_U3342 , P1_U4045 , P1_U4046 , P1_U4044 );
nand NAND3_647 ( P1_U3343 , P1_U4042 , P1_U4043 , P1_U4041 );
nand NAND3_648 ( P1_U3344 , P1_U4039 , P1_U4040 , P1_U4038 );
nand NAND3_649 ( P1_U3345 , P1_U4036 , P1_U4037 , P1_U4035 );
nand NAND3_650 ( P1_U3346 , P1_U4033 , P1_U4034 , P1_U4032 );
nand NAND3_651 ( P1_U3347 , P1_U4030 , P1_U4031 , P1_U4029 );
nand NAND3_652 ( P1_U3348 , P1_U4027 , P1_U4028 , P1_U4026 );
nand NAND3_653 ( P1_U3349 , P1_U4024 , P1_U4025 , P1_U4023 );
nand NAND3_654 ( P1_U3350 , P1_U4021 , P1_U4022 , P1_U4020 );
nand NAND3_655 ( P1_U3351 , P1_U4018 , P1_U4019 , P1_U4017 );
nand NAND3_656 ( P1_U3352 , P1_U4015 , P1_U4016 , P1_U4014 );
nand NAND3_657 ( P1_U3353 , P1_U4012 , P1_U4013 , P1_U4011 );
nand NAND3_658 ( P1_U3354 , P1_U4009 , P1_U4010 , P1_U4008 );
nand NAND3_659 ( P1_U3355 , P1_U4006 , P1_U4007 , P1_U4005 );
nand NAND5_660 ( P1_U3356 , P1_U4874 , P1_U4872 , P1_U4875 , P1_U4873 , P1_U3944 );
nand NAND2_661 ( P1_U3357 , P1_STATE_REG , P1_U3910 );
nand NAND2_662 ( P1_U3358 , P1_U3437 , P1_U5669 );
not NOT1_663 ( P1_U3359 , P1_B_REG );
nand NAND3_664 ( P1_U3360 , P1_U5674 , P1_U5673 , P1_U3437 );
nand NAND2_665 ( P1_U3361 , P1_U3048 , P1_U3443 );
nand NAND3_666 ( P1_U3362 , P1_U3441 , P1_U3442 , P1_U3443 );
nand NAND2_667 ( P1_U3363 , P1_U3441 , P1_U5687 );
nand NAND2_668 ( P1_U3364 , P1_U4001 , P1_U3443 );
nand NAND3_669 ( P1_U3365 , P1_U3441 , P1_U3442 , P1_U3447 );
nand NAND2_670 ( P1_U3366 , P1_U4001 , P1_U3447 );
nand NAND2_671 ( P1_U3367 , P1_U5690 , P1_U5687 );
nand NAND2_672 ( P1_U3368 , P1_U4002 , P1_U3443 );
nand NAND2_673 ( P1_U3369 , P1_U3960 , P1_U5693 );
nand NAND2_674 ( P1_U3370 , P1_U4002 , P1_U3447 );
nand NAND2_675 ( P1_U3371 , P1_U3956 , P1_U5684 );
nand NAND2_676 ( P1_U3372 , P1_U5684 , P1_U3442 );
nand NAND2_677 ( P1_U3373 , P1_U3443 , P1_U3447 );
nand NAND5_678 ( P1_U3374 , P1_U4148 , P1_U4147 , P1_U4149 , P1_U3619 , P1_U3618 );
not NOT1_679 ( P1_U3375 , P1_REG2_REG_0_ );
nand NAND4_680 ( P1_U3376 , P1_U4167 , P1_U4166 , P1_U3633 , P1_U3635 );
nand NAND4_681 ( P1_U3377 , P1_U4186 , P1_U4185 , P1_U3637 , P1_U3639 );
nand NAND5_682 ( P1_U3378 , P1_U4205 , P1_U4204 , P1_U4206 , P1_U4207 , P1_U3642 );
nand NAND5_683 ( P1_U3379 , P1_U4224 , P1_U4223 , P1_U4225 , P1_U4226 , P1_U3645 );
nand NAND4_684 ( P1_U3380 , P1_U4243 , P1_U4242 , P1_U3647 , P1_U3649 );
nand NAND4_685 ( P1_U3381 , P1_U4262 , P1_U4261 , P1_U3651 , P1_U3653 );
nand NAND4_686 ( P1_U3382 , P1_U4281 , P1_U4280 , P1_U3655 , P1_U3657 );
nand NAND4_687 ( P1_U3383 , P1_U4300 , P1_U4299 , P1_U3659 , P1_U3661 );
nand NAND4_688 ( P1_U3384 , P1_U4319 , P1_U4318 , P1_U3663 , P1_U3665 );
nand NAND4_689 ( P1_U3385 , P1_U4338 , P1_U4337 , P1_U3667 , P1_U3669 );
nand NAND4_690 ( P1_U3386 , P1_U4357 , P1_U4356 , P1_U3671 , P1_U3673 );
nand NAND4_691 ( P1_U3387 , P1_U4376 , P1_U4375 , P1_U3675 , P1_U3677 );
nand NAND4_692 ( P1_U3388 , P1_U4395 , P1_U4394 , P1_U3679 , P1_U3681 );
nand NAND4_693 ( P1_U3389 , P1_U4414 , P1_U4413 , P1_U3683 , P1_U3685 );
nand NAND4_694 ( P1_U3390 , P1_U4433 , P1_U4432 , P1_U3687 , P1_U3689 );
nand NAND4_695 ( P1_U3391 , P1_U4452 , P1_U4451 , P1_U3691 , P1_U3693 );
nand NAND4_696 ( P1_U3392 , P1_U4471 , P1_U4470 , P1_U3695 , P1_U3697 );
nand NAND4_697 ( P1_U3393 , P1_U4490 , P1_U4489 , P1_U3699 , P1_U3701 );
nand NAND4_698 ( P1_U3394 , P1_U4509 , P1_U4508 , P1_U3703 , P1_U3705 );
nand NAND2_699 ( P1_U3395 , U76 , P1_U3912 );
nand NAND4_700 ( P1_U3396 , P1_U4528 , P1_U4527 , P1_U3707 , P1_U3709 );
nand NAND2_701 ( P1_U3397 , U75 , P1_U3912 );
nand NAND4_702 ( P1_U3398 , P1_U4547 , P1_U4546 , P1_U3711 , P1_U3713 );
nand NAND2_703 ( P1_U3399 , U74 , P1_U3912 );
nand NAND4_704 ( P1_U3400 , P1_U4566 , P1_U4565 , P1_U3715 , P1_U3717 );
nand NAND2_705 ( P1_U3401 , U73 , P1_U3912 );
nand NAND4_706 ( P1_U3402 , P1_U4585 , P1_U4584 , P1_U3719 , P1_U3721 );
nand NAND2_707 ( P1_U3403 , U72 , P1_U3912 );
nand NAND4_708 ( P1_U3404 , P1_U4604 , P1_U4603 , P1_U3723 , P1_U3725 );
nand NAND2_709 ( P1_U3405 , U71 , P1_U3912 );
nand NAND4_710 ( P1_U3406 , P1_U4623 , P1_U4622 , P1_U3727 , P1_U3729 );
nand NAND2_711 ( P1_U3407 , U70 , P1_U3912 );
nand NAND4_712 ( P1_U3408 , P1_U4642 , P1_U4641 , P1_U3731 , P1_U3733 );
nand NAND2_713 ( P1_U3409 , U69 , P1_U3912 );
nand NAND4_714 ( P1_U3410 , P1_U4661 , P1_U4660 , P1_U3735 , P1_U3737 );
nand NAND2_715 ( P1_U3411 , U68 , P1_U3912 );
nand NAND4_716 ( P1_U3412 , P1_U4680 , P1_U4679 , P1_U3739 , P1_U3741 );
nand NAND2_717 ( P1_U3413 , U67 , P1_U3912 );
nand NAND2_718 ( P1_U3414 , U65 , P1_U3912 );
nand NAND2_719 ( P1_U3415 , U64 , P1_U3912 );
nand NAND2_720 ( P1_U3416 , P1_U3953 , P1_U5693 );
nand NAND2_721 ( P1_U3417 , P1_U3022 , P1_U4724 );
nand NAND2_722 ( P1_U3418 , P1_U3988 , P1_U5690 );
nand NAND2_723 ( P1_U3419 , P1_U3048 , P1_U3447 );
nand NAND2_724 ( P1_U3420 , P1_U3023 , P1_U5687 );
nand NAND2_725 ( P1_U3421 , P1_U3050 , P1_U3436 );
nand NAND2_726 ( P1_U3422 , P1_U3966 , P1_U4725 );
nand NAND2_727 ( P1_U3423 , P1_U3424 , P1_U4888 );
nand NAND2_728 ( P1_U3424 , P1_U4102 , P1_U5677 );
nand NAND2_729 ( P1_U3425 , P1_U3999 , P1_STATE_REG );
nand NAND2_730 ( P1_U3426 , P1_U3438 , P1_U5687 );
nand NAND2_731 ( P1_U3427 , P1_U3014 , P1_U3015 );
nand NAND2_732 ( P1_U3428 , P1_U3443 , P1_U3438 );
nand NAND2_733 ( P1_U3429 , P1_U3022 , P1_U3422 );
nand NAND2_734 ( P1_U3430 , P1_U3867 , P1_U3016 );
nand NAND2_735 ( P1_U3431 , P1_U3014 , P1_U3022 );
nand NAND2_736 ( P1_U3432 , P1_U3870 , P1_U5101 );
nand NAND2_737 ( P1_U3433 , P1_U3442 , P1_U5693 );
nand NAND2_738 ( P1_U3434 , P1_U5371 , P1_U5370 );
nand NAND2_739 ( P1_U3435 , P1_U5665 , P1_U5664 );
nand NAND2_740 ( P1_U3436 , P1_U5668 , P1_U5667 );
nand NAND2_741 ( P1_U3437 , P1_U5671 , P1_U5670 );
nand NAND2_742 ( P1_U3438 , P1_U5676 , P1_U5675 );
nand NAND2_743 ( P1_U3439 , P1_U5679 , P1_U5678 );
nand NAND2_744 ( P1_U3440 , P1_U5681 , P1_U5680 );
nand NAND2_745 ( P1_U3441 , P1_U5689 , P1_U5688 );
nand NAND2_746 ( P1_U3442 , P1_U5686 , P1_U5685 );
nand NAND2_747 ( P1_U3443 , P1_U5683 , P1_U5682 );
nand NAND2_748 ( P1_U3444 , P1_U5707 , P1_U5706 );
nand NAND2_749 ( P1_U3445 , P1_U5710 , P1_U5709 );
nand NAND2_750 ( P1_U3446 , P1_U5698 , P1_U5697 );
nand NAND2_751 ( P1_U3447 , P1_U5692 , P1_U5691 );
nand NAND2_752 ( P1_U3448 , P1_U5695 , P1_U5694 );
nand NAND2_753 ( P1_U3449 , P1_U5701 , P1_U5700 );
nand NAND2_754 ( P1_U3450 , P1_U5704 , P1_U5703 );
nand NAND2_755 ( P1_U3451 , P1_U5718 , P1_U5717 );
nand NAND2_756 ( P1_U3452 , P1_U5715 , P1_U5714 );
nand NAND2_757 ( P1_U3453 , P1_U5721 , P1_U5720 );
nand NAND2_758 ( P1_U3454 , P1_U5723 , P1_U5722 );
nand NAND2_759 ( P1_U3455 , P1_U5725 , P1_U5724 );
nand NAND2_760 ( P1_U3456 , P1_U5728 , P1_U5727 );
nand NAND2_761 ( P1_U3457 , P1_U5730 , P1_U5729 );
nand NAND2_762 ( P1_U3458 , P1_U5732 , P1_U5731 );
nand NAND2_763 ( P1_U3459 , P1_U5735 , P1_U5734 );
nand NAND2_764 ( P1_U3460 , P1_U5737 , P1_U5736 );
nand NAND2_765 ( P1_U3461 , P1_U5739 , P1_U5738 );
nand NAND2_766 ( P1_U3462 , P1_U5742 , P1_U5741 );
nand NAND2_767 ( P1_U3463 , P1_U5744 , P1_U5743 );
nand NAND2_768 ( P1_U3464 , P1_U5746 , P1_U5745 );
nand NAND2_769 ( P1_U3465 , P1_U5749 , P1_U5748 );
nand NAND2_770 ( P1_U3466 , P1_U5751 , P1_U5750 );
nand NAND2_771 ( P1_U3467 , P1_U5753 , P1_U5752 );
nand NAND2_772 ( P1_U3468 , P1_U5756 , P1_U5755 );
nand NAND2_773 ( P1_U3469 , P1_U5758 , P1_U5757 );
nand NAND2_774 ( P1_U3470 , P1_U5760 , P1_U5759 );
nand NAND2_775 ( P1_U3471 , P1_U5763 , P1_U5762 );
nand NAND2_776 ( P1_U3472 , P1_U5765 , P1_U5764 );
nand NAND2_777 ( P1_U3473 , P1_U5767 , P1_U5766 );
nand NAND2_778 ( P1_U3474 , P1_U5770 , P1_U5769 );
nand NAND2_779 ( P1_U3475 , P1_U5772 , P1_U5771 );
nand NAND2_780 ( P1_U3476 , P1_U5774 , P1_U5773 );
nand NAND2_781 ( P1_U3477 , P1_U5777 , P1_U5776 );
nand NAND2_782 ( P1_U3478 , P1_U5779 , P1_U5778 );
nand NAND2_783 ( P1_U3479 , P1_U5781 , P1_U5780 );
nand NAND2_784 ( P1_U3480 , P1_U5784 , P1_U5783 );
nand NAND2_785 ( P1_U3481 , P1_U5786 , P1_U5785 );
nand NAND2_786 ( P1_U3482 , P1_U5788 , P1_U5787 );
nand NAND2_787 ( P1_U3483 , P1_U5791 , P1_U5790 );
nand NAND2_788 ( P1_U3484 , P1_U5793 , P1_U5792 );
nand NAND2_789 ( P1_U3485 , P1_U5795 , P1_U5794 );
nand NAND2_790 ( P1_U3486 , P1_U5798 , P1_U5797 );
nand NAND2_791 ( P1_U3487 , P1_U5800 , P1_U5799 );
nand NAND2_792 ( P1_U3488 , P1_U5802 , P1_U5801 );
nand NAND2_793 ( P1_U3489 , P1_U5805 , P1_U5804 );
nand NAND2_794 ( P1_U3490 , P1_U5807 , P1_U5806 );
nand NAND2_795 ( P1_U3491 , P1_U5809 , P1_U5808 );
nand NAND2_796 ( P1_U3492 , P1_U5812 , P1_U5811 );
nand NAND2_797 ( P1_U3493 , P1_U5814 , P1_U5813 );
nand NAND2_798 ( P1_U3494 , P1_U5816 , P1_U5815 );
nand NAND2_799 ( P1_U3495 , P1_U5819 , P1_U5818 );
nand NAND2_800 ( P1_U3496 , P1_U5821 , P1_U5820 );
nand NAND2_801 ( P1_U3497 , P1_U5823 , P1_U5822 );
nand NAND2_802 ( P1_U3498 , P1_U5826 , P1_U5825 );
nand NAND2_803 ( P1_U3499 , P1_U5828 , P1_U5827 );
nand NAND2_804 ( P1_U3500 , P1_U5830 , P1_U5829 );
nand NAND2_805 ( P1_U3501 , P1_U5833 , P1_U5832 );
nand NAND2_806 ( P1_U3502 , P1_U5835 , P1_U5834 );
nand NAND2_807 ( P1_U3503 , P1_U5837 , P1_U5836 );
nand NAND2_808 ( P1_U3504 , P1_U5840 , P1_U5839 );
nand NAND2_809 ( P1_U3505 , P1_U5842 , P1_U5841 );
nand NAND2_810 ( P1_U3506 , P1_U5844 , P1_U5843 );
nand NAND2_811 ( P1_U3507 , P1_U5847 , P1_U5846 );
nand NAND2_812 ( P1_U3508 , P1_U5849 , P1_U5848 );
nand NAND2_813 ( P1_U3509 , P1_U5852 , P1_U5851 );
nand NAND2_814 ( P1_U3510 , P1_U5854 , P1_U5853 );
nand NAND2_815 ( P1_U3511 , P1_U5856 , P1_U5855 );
nand NAND2_816 ( P1_U3512 , P1_U5858 , P1_U5857 );
nand NAND2_817 ( P1_U3513 , P1_U5860 , P1_U5859 );
nand NAND2_818 ( P1_U3514 , P1_U5862 , P1_U5861 );
nand NAND2_819 ( P1_U3515 , P1_U5864 , P1_U5863 );
nand NAND2_820 ( P1_U3516 , P1_U5866 , P1_U5865 );
nand NAND2_821 ( P1_U3517 , P1_U5868 , P1_U5867 );
nand NAND2_822 ( P1_U3518 , P1_U5870 , P1_U5869 );
nand NAND2_823 ( P1_U3519 , P1_U5872 , P1_U5871 );
nand NAND2_824 ( P1_U3520 , P1_U5874 , P1_U5873 );
nand NAND2_825 ( P1_U3521 , P1_U5876 , P1_U5875 );
nand NAND2_826 ( P1_U3522 , P1_U5878 , P1_U5877 );
nand NAND2_827 ( P1_U3523 , P1_U5880 , P1_U5879 );
nand NAND2_828 ( P1_U3524 , P1_U5882 , P1_U5881 );
nand NAND2_829 ( P1_U3525 , P1_U5884 , P1_U5883 );
nand NAND2_830 ( P1_U3526 , P1_U5886 , P1_U5885 );
nand NAND2_831 ( P1_U3527 , P1_U5888 , P1_U5887 );
nand NAND2_832 ( P1_U3528 , P1_U5890 , P1_U5889 );
nand NAND2_833 ( P1_U3529 , P1_U5892 , P1_U5891 );
nand NAND2_834 ( P1_U3530 , P1_U5894 , P1_U5893 );
nand NAND2_835 ( P1_U3531 , P1_U5896 , P1_U5895 );
nand NAND2_836 ( P1_U3532 , P1_U5898 , P1_U5897 );
nand NAND2_837 ( P1_U3533 , P1_U5900 , P1_U5899 );
nand NAND2_838 ( P1_U3534 , P1_U5902 , P1_U5901 );
nand NAND2_839 ( P1_U3535 , P1_U5904 , P1_U5903 );
nand NAND2_840 ( P1_U3536 , P1_U5906 , P1_U5905 );
nand NAND2_841 ( P1_U3537 , P1_U5908 , P1_U5907 );
nand NAND2_842 ( P1_U3538 , P1_U5910 , P1_U5909 );
nand NAND2_843 ( P1_U3539 , P1_U5912 , P1_U5911 );
nand NAND2_844 ( P1_U3540 , P1_U5914 , P1_U5913 );
nand NAND2_845 ( P1_U3541 , P1_U5916 , P1_U5915 );
nand NAND2_846 ( P1_U3542 , P1_U5918 , P1_U5917 );
nand NAND2_847 ( P1_U3543 , P1_U5920 , P1_U5919 );
nand NAND2_848 ( P1_U3544 , P1_U5922 , P1_U5921 );
nand NAND2_849 ( P1_U3545 , P1_U5924 , P1_U5923 );
nand NAND2_850 ( P1_U3546 , P1_U5926 , P1_U5925 );
nand NAND2_851 ( P1_U3547 , P1_U5928 , P1_U5927 );
nand NAND2_852 ( P1_U3548 , P1_U5930 , P1_U5929 );
nand NAND2_853 ( P1_U3549 , P1_U5932 , P1_U5931 );
nand NAND2_854 ( P1_U3550 , P1_U5934 , P1_U5933 );
nand NAND2_855 ( P1_U3551 , P1_U5936 , P1_U5935 );
nand NAND2_856 ( P1_U3552 , P1_U5938 , P1_U5937 );
nand NAND2_857 ( P1_U3553 , P1_U5940 , P1_U5939 );
nand NAND2_858 ( P1_U3554 , P1_U6006 , P1_U6005 );
nand NAND2_859 ( P1_U3555 , P1_U6008 , P1_U6007 );
nand NAND2_860 ( P1_U3556 , P1_U6010 , P1_U6009 );
nand NAND2_861 ( P1_U3557 , P1_U6012 , P1_U6011 );
nand NAND2_862 ( P1_U3558 , P1_U6014 , P1_U6013 );
nand NAND2_863 ( P1_U3559 , P1_U6016 , P1_U6015 );
nand NAND2_864 ( P1_U3560 , P1_U6018 , P1_U6017 );
nand NAND2_865 ( P1_U3561 , P1_U6020 , P1_U6019 );
nand NAND2_866 ( P1_U3562 , P1_U6022 , P1_U6021 );
nand NAND2_867 ( P1_U3563 , P1_U6024 , P1_U6023 );
nand NAND2_868 ( P1_U3564 , P1_U6026 , P1_U6025 );
nand NAND2_869 ( P1_U3565 , P1_U6028 , P1_U6027 );
nand NAND2_870 ( P1_U3566 , P1_U6030 , P1_U6029 );
nand NAND2_871 ( P1_U3567 , P1_U6032 , P1_U6031 );
nand NAND2_872 ( P1_U3568 , P1_U6034 , P1_U6033 );
nand NAND2_873 ( P1_U3569 , P1_U6036 , P1_U6035 );
nand NAND2_874 ( P1_U3570 , P1_U6038 , P1_U6037 );
nand NAND2_875 ( P1_U3571 , P1_U6040 , P1_U6039 );
nand NAND2_876 ( P1_U3572 , P1_U6042 , P1_U6041 );
nand NAND2_877 ( P1_U3573 , P1_U6044 , P1_U6043 );
nand NAND2_878 ( P1_U3574 , P1_U6046 , P1_U6045 );
nand NAND2_879 ( P1_U3575 , P1_U6048 , P1_U6047 );
nand NAND2_880 ( P1_U3576 , P1_U6050 , P1_U6049 );
nand NAND2_881 ( P1_U3577 , P1_U6052 , P1_U6051 );
nand NAND2_882 ( P1_U3578 , P1_U6054 , P1_U6053 );
nand NAND2_883 ( P1_U3579 , P1_U6056 , P1_U6055 );
nand NAND2_884 ( P1_U3580 , P1_U6058 , P1_U6057 );
nand NAND2_885 ( P1_U3581 , P1_U6060 , P1_U6059 );
nand NAND2_886 ( P1_U3582 , P1_U6062 , P1_U6061 );
nand NAND2_887 ( P1_U3583 , P1_U6064 , P1_U6063 );
nand NAND2_888 ( P1_U3584 , P1_U6066 , P1_U6065 );
nand NAND2_889 ( P1_U3585 , P1_U6068 , P1_U6067 );
nand NAND2_890 ( P1_U3586 , P1_U6172 , P1_U6171 );
nand NAND2_891 ( P1_U3587 , P1_U6174 , P1_U6173 );
nand NAND2_892 ( P1_U3588 , P1_U6176 , P1_U6175 );
nand NAND2_893 ( P1_U3589 , P1_U6178 , P1_U6177 );
nand NAND2_894 ( P1_U3590 , P1_U6180 , P1_U6179 );
nand NAND2_895 ( P1_U3591 , P1_U6182 , P1_U6181 );
nand NAND2_896 ( P1_U3592 , P1_U6184 , P1_U6183 );
nand NAND2_897 ( P1_U3593 , P1_U6186 , P1_U6185 );
nand NAND2_898 ( P1_U3594 , P1_U6188 , P1_U6187 );
nand NAND2_899 ( P1_U3595 , P1_U6190 , P1_U6189 );
nand NAND2_900 ( P1_U3596 , P1_U6192 , P1_U6191 );
nand NAND2_901 ( P1_U3597 , P1_U6194 , P1_U6193 );
nand NAND2_902 ( P1_U3598 , P1_U6196 , P1_U6195 );
nand NAND2_903 ( P1_U3599 , P1_U6198 , P1_U6197 );
nand NAND2_904 ( P1_U3600 , P1_U6200 , P1_U6199 );
nand NAND2_905 ( P1_U3601 , P1_U6202 , P1_U6201 );
nand NAND2_906 ( P1_U3602 , P1_U6204 , P1_U6203 );
nand NAND2_907 ( P1_U3603 , P1_U6206 , P1_U6205 );
nand NAND2_908 ( P1_U3604 , P1_U6208 , P1_U6207 );
nand NAND2_909 ( P1_U3605 , P1_U6210 , P1_U6209 );
nand NAND2_910 ( P1_U3606 , P1_U6212 , P1_U6211 );
nand NAND2_911 ( P1_U3607 , P1_U6214 , P1_U6213 );
nand NAND2_912 ( P1_U3608 , P1_U6216 , P1_U6215 );
nand NAND2_913 ( P1_U3609 , P1_U6218 , P1_U6217 );
nand NAND2_914 ( P1_U3610 , P1_U6220 , P1_U6219 );
nand NAND2_915 ( P1_U3611 , P1_U6222 , P1_U6221 );
nand NAND2_916 ( P1_U3612 , P1_U6224 , P1_U6223 );
nand NAND2_917 ( P1_U3613 , P1_U6226 , P1_U6225 );
nand NAND2_918 ( P1_U3614 , P1_U6228 , P1_U6227 );
nand NAND2_919 ( P1_U3615 , P1_U6230 , P1_U6229 );
nand NAND2_920 ( P1_U3616 , P1_U6232 , P1_U6231 );
nand NAND2_921 ( P1_U3617 , P1_U6234 , P1_U6233 );
and AND2_922 ( P1_U3618 , P1_U4144 , P1_U4143 );
and AND2_923 ( P1_U3619 , P1_U4146 , P1_U4145 );
and AND4_924 ( P1_U3620 , P1_U4152 , P1_U4153 , P1_U4154 , P1_U4151 );
and AND4_925 ( P1_U3621 , P1_U4108 , P1_U4107 , P1_U4106 , P1_U4105 );
and AND4_926 ( P1_U3622 , P1_U4112 , P1_U4111 , P1_U4110 , P1_U4109 );
and AND4_927 ( P1_U3623 , P1_U4116 , P1_U4115 , P1_U4114 , P1_U4113 );
and AND3_928 ( P1_U3624 , P1_U4118 , P1_U4117 , P1_U4119 );
and AND4_929 ( P1_U3625 , P1_U3624 , P1_U3623 , P1_U3622 , P1_U3621 );
and AND4_930 ( P1_U3626 , P1_U4123 , P1_U4122 , P1_U4121 , P1_U4120 );
and AND4_931 ( P1_U3627 , P1_U4127 , P1_U4126 , P1_U4125 , P1_U4124 );
and AND4_932 ( P1_U3628 , P1_U4131 , P1_U4130 , P1_U4129 , P1_U4128 );
and AND3_933 ( P1_U3629 , P1_U4133 , P1_U4132 , P1_U4134 );
and AND4_934 ( P1_U3630 , P1_U3629 , P1_U3628 , P1_U3627 , P1_U3626 );
and AND2_935 ( P1_U3631 , P1_U5716 , P1_U4136 );
and AND2_936 ( P1_U3632 , P1_U5719 , P1_U3022 );
and AND2_937 ( P1_U3633 , P1_U4169 , P1_U4168 );
and AND2_938 ( P1_U3634 , P1_U4171 , P1_U4170 );
and AND3_939 ( P1_U3635 , P1_U4173 , P1_U4172 , P1_U3634 );
and AND4_940 ( P1_U3636 , P1_U4176 , P1_U4177 , P1_U4178 , P1_U4175 );
and AND2_941 ( P1_U3637 , P1_U4188 , P1_U4187 );
and AND2_942 ( P1_U3638 , P1_U4190 , P1_U4189 );
and AND3_943 ( P1_U3639 , P1_U4192 , P1_U4191 , P1_U3638 );
and AND4_944 ( P1_U3640 , P1_U4195 , P1_U4196 , P1_U4197 , P1_U4194 );
and AND2_945 ( P1_U3641 , P1_U4209 , P1_U4208 );
and AND3_946 ( P1_U3642 , P1_U4211 , P1_U4210 , P1_U3641 );
and AND4_947 ( P1_U3643 , P1_U4214 , P1_U4215 , P1_U4216 , P1_U4213 );
and AND2_948 ( P1_U3644 , P1_U4228 , P1_U4227 );
and AND3_949 ( P1_U3645 , P1_U4230 , P1_U4229 , P1_U3644 );
and AND4_950 ( P1_U3646 , P1_U4233 , P1_U4234 , P1_U4235 , P1_U4232 );
and AND2_951 ( P1_U3647 , P1_U4245 , P1_U4244 );
and AND2_952 ( P1_U3648 , P1_U4247 , P1_U4246 );
and AND3_953 ( P1_U3649 , P1_U4249 , P1_U4248 , P1_U3648 );
and AND4_954 ( P1_U3650 , P1_U4252 , P1_U4253 , P1_U4254 , P1_U4251 );
and AND2_955 ( P1_U3651 , P1_U4264 , P1_U4263 );
and AND2_956 ( P1_U3652 , P1_U4266 , P1_U4265 );
and AND3_957 ( P1_U3653 , P1_U4268 , P1_U4267 , P1_U3652 );
and AND4_958 ( P1_U3654 , P1_U4271 , P1_U4272 , P1_U4273 , P1_U4270 );
and AND2_959 ( P1_U3655 , P1_U4283 , P1_U4282 );
and AND2_960 ( P1_U3656 , P1_U4285 , P1_U4284 );
and AND3_961 ( P1_U3657 , P1_U4287 , P1_U4286 , P1_U3656 );
and AND4_962 ( P1_U3658 , P1_U4290 , P1_U4291 , P1_U4292 , P1_U4289 );
and AND2_963 ( P1_U3659 , P1_U4302 , P1_U4301 );
and AND2_964 ( P1_U3660 , P1_U4304 , P1_U4303 );
and AND3_965 ( P1_U3661 , P1_U4306 , P1_U4305 , P1_U3660 );
and AND4_966 ( P1_U3662 , P1_U4309 , P1_U4310 , P1_U4311 , P1_U4308 );
and AND2_967 ( P1_U3663 , P1_U4321 , P1_U4320 );
and AND2_968 ( P1_U3664 , P1_U4323 , P1_U4322 );
and AND3_969 ( P1_U3665 , P1_U4325 , P1_U4324 , P1_U3664 );
and AND4_970 ( P1_U3666 , P1_U4328 , P1_U4329 , P1_U4330 , P1_U4327 );
and AND2_971 ( P1_U3667 , P1_U4340 , P1_U4339 );
and AND2_972 ( P1_U3668 , P1_U4342 , P1_U4341 );
and AND3_973 ( P1_U3669 , P1_U4344 , P1_U4343 , P1_U3668 );
and AND4_974 ( P1_U3670 , P1_U4347 , P1_U4348 , P1_U4349 , P1_U4346 );
and AND2_975 ( P1_U3671 , P1_U4359 , P1_U4358 );
and AND2_976 ( P1_U3672 , P1_U4361 , P1_U4360 );
and AND3_977 ( P1_U3673 , P1_U4363 , P1_U4362 , P1_U3672 );
and AND4_978 ( P1_U3674 , P1_U4368 , P1_U4365 , P1_U4366 , P1_U4367 );
and AND2_979 ( P1_U3675 , P1_U4378 , P1_U4377 );
and AND2_980 ( P1_U3676 , P1_U4380 , P1_U4379 );
and AND3_981 ( P1_U3677 , P1_U4382 , P1_U4381 , P1_U3676 );
and AND4_982 ( P1_U3678 , P1_U4387 , P1_U4384 , P1_U4385 , P1_U4386 );
and AND2_983 ( P1_U3679 , P1_U4397 , P1_U4396 );
and AND2_984 ( P1_U3680 , P1_U4399 , P1_U4398 );
and AND3_985 ( P1_U3681 , P1_U4401 , P1_U4400 , P1_U3680 );
and AND4_986 ( P1_U3682 , P1_U4406 , P1_U4405 , P1_U4404 , P1_U4403 );
and AND2_987 ( P1_U3683 , P1_U4416 , P1_U4415 );
and AND2_988 ( P1_U3684 , P1_U4418 , P1_U4417 );
and AND3_989 ( P1_U3685 , P1_U4420 , P1_U4419 , P1_U3684 );
and AND4_990 ( P1_U3686 , P1_U4423 , P1_U4422 , P1_U4425 , P1_U4424 );
and AND2_991 ( P1_U3687 , P1_U4435 , P1_U4434 );
and AND2_992 ( P1_U3688 , P1_U4437 , P1_U4436 );
and AND3_993 ( P1_U3689 , P1_U4439 , P1_U4438 , P1_U3688 );
and AND4_994 ( P1_U3690 , P1_U4442 , P1_U4441 , P1_U4444 , P1_U4443 );
and AND2_995 ( P1_U3691 , P1_U4454 , P1_U4453 );
and AND2_996 ( P1_U3692 , P1_U4456 , P1_U4455 );
and AND3_997 ( P1_U3693 , P1_U4458 , P1_U4457 , P1_U3692 );
and AND4_998 ( P1_U3694 , P1_U4461 , P1_U4460 , P1_U4463 , P1_U4462 );
and AND2_999 ( P1_U3695 , P1_U4473 , P1_U4472 );
and AND2_1000 ( P1_U3696 , P1_U4475 , P1_U4474 );
and AND3_1001 ( P1_U3697 , P1_U4477 , P1_U4476 , P1_U3696 );
and AND4_1002 ( P1_U3698 , P1_U4480 , P1_U4479 , P1_U4482 , P1_U4481 );
and AND2_1003 ( P1_U3699 , P1_U4492 , P1_U4491 );
and AND2_1004 ( P1_U3700 , P1_U4494 , P1_U4493 );
and AND3_1005 ( P1_U3701 , P1_U4496 , P1_U4495 , P1_U3700 );
and AND4_1006 ( P1_U3702 , P1_U4499 , P1_U4498 , P1_U4501 , P1_U4500 );
and AND2_1007 ( P1_U3703 , P1_U4511 , P1_U4510 );
and AND2_1008 ( P1_U3704 , P1_U4513 , P1_U4512 );
and AND3_1009 ( P1_U3705 , P1_U4515 , P1_U4514 , P1_U3704 );
and AND4_1010 ( P1_U3706 , P1_U4518 , P1_U4517 , P1_U4520 , P1_U4519 );
and AND2_1011 ( P1_U3707 , P1_U4530 , P1_U4529 );
and AND2_1012 ( P1_U3708 , P1_U4532 , P1_U4531 );
and AND3_1013 ( P1_U3709 , P1_U4534 , P1_U4533 , P1_U3708 );
and AND4_1014 ( P1_U3710 , P1_U4539 , P1_U4538 , P1_U4537 , P1_U4536 );
and AND2_1015 ( P1_U3711 , P1_U4549 , P1_U4548 );
and AND2_1016 ( P1_U3712 , P1_U4551 , P1_U4550 );
and AND3_1017 ( P1_U3713 , P1_U4553 , P1_U4552 , P1_U3712 );
and AND4_1018 ( P1_U3714 , P1_U4556 , P1_U4555 , P1_U4558 , P1_U4557 );
and AND2_1019 ( P1_U3715 , P1_U4568 , P1_U4567 );
and AND2_1020 ( P1_U3716 , P1_U4570 , P1_U4569 );
and AND3_1021 ( P1_U3717 , P1_U4572 , P1_U4571 , P1_U3716 );
and AND4_1022 ( P1_U3718 , P1_U4577 , P1_U4576 , P1_U4575 , P1_U4574 );
and AND2_1023 ( P1_U3719 , P1_U4587 , P1_U4586 );
and AND2_1024 ( P1_U3720 , P1_U4589 , P1_U4588 );
and AND3_1025 ( P1_U3721 , P1_U4591 , P1_U4590 , P1_U3720 );
and AND4_1026 ( P1_U3722 , P1_U4596 , P1_U4593 , P1_U4594 , P1_U4595 );
and AND2_1027 ( P1_U3723 , P1_U4606 , P1_U4605 );
and AND2_1028 ( P1_U3724 , P1_U4608 , P1_U4607 );
and AND3_1029 ( P1_U3725 , P1_U4610 , P1_U4609 , P1_U3724 );
and AND4_1030 ( P1_U3726 , P1_U4613 , P1_U4614 , P1_U4615 , P1_U4612 );
and AND2_1031 ( P1_U3727 , P1_U4625 , P1_U4624 );
and AND2_1032 ( P1_U3728 , P1_U4627 , P1_U4626 );
and AND3_1033 ( P1_U3729 , P1_U4629 , P1_U4628 , P1_U3728 );
and AND4_1034 ( P1_U3730 , P1_U4632 , P1_U4633 , P1_U4634 , P1_U4631 );
and AND2_1035 ( P1_U3731 , P1_U4644 , P1_U4643 );
and AND2_1036 ( P1_U3732 , P1_U4646 , P1_U4645 );
and AND3_1037 ( P1_U3733 , P1_U4648 , P1_U4647 , P1_U3732 );
and AND4_1038 ( P1_U3734 , P1_U4651 , P1_U4652 , P1_U4653 , P1_U4650 );
and AND2_1039 ( P1_U3735 , P1_U4663 , P1_U4662 );
and AND2_1040 ( P1_U3736 , P1_U4665 , P1_U4664 );
and AND3_1041 ( P1_U3737 , P1_U4667 , P1_U4666 , P1_U3736 );
and AND4_1042 ( P1_U3738 , P1_U4670 , P1_U4671 , P1_U4672 , P1_U4669 );
and AND2_1043 ( P1_U3739 , P1_U4682 , P1_U4681 );
and AND2_1044 ( P1_U3740 , P1_U4684 , P1_U4683 );
and AND3_1045 ( P1_U3741 , P1_U4686 , P1_U4685 , P1_U3740 );
and AND4_1046 ( P1_U3742 , P1_U4689 , P1_U4690 , P1_U4691 , P1_U4688 );
and AND2_1047 ( P1_U3743 , P1_U4698 , P1_U3987 );
and AND3_1048 ( P1_U3744 , P1_U4702 , P1_U4701 , P1_U4704 );
and AND2_1049 ( P1_U3745 , P1_U4707 , P1_U4705 );
and AND3_1050 ( P1_U3746 , P1_U4710 , P1_U4711 , P1_U4709 );
and AND2_1051 ( P1_U3747 , P1_U3987 , P1_U4698 );
and AND2_1052 ( P1_U3748 , P1_U3022 , P1_U3451 );
and AND3_1053 ( P1_U3749 , P1_U5719 , P1_U3969 , P1_U3452 );
and AND3_1054 ( P1_U3750 , P1_U4728 , P1_U4727 , P1_U4729 );
and AND3_1055 ( P1_U3751 , P1_U4731 , P1_U4730 , P1_U3915 );
and AND3_1056 ( P1_U3752 , P1_U4733 , P1_U4732 , P1_U4734 );
and AND3_1057 ( P1_U3753 , P1_U4736 , P1_U4735 , P1_U3916 );
and AND3_1058 ( P1_U3754 , P1_U4738 , P1_U4737 , P1_U4739 );
and AND3_1059 ( P1_U3755 , P1_U4741 , P1_U4740 , P1_U3917 );
and AND3_1060 ( P1_U3756 , P1_U4743 , P1_U4742 , P1_U4744 );
and AND2_1061 ( P1_U3757 , P1_U4746 , P1_U4745 );
and AND2_1062 ( P1_U3758 , P1_U4748 , P1_U4747 );
and AND2_1063 ( P1_U3759 , P1_U4751 , P1_U4750 );
and AND2_1064 ( P1_U3760 , P1_U4753 , P1_U4752 );
and AND2_1065 ( P1_U3761 , P1_U4756 , P1_U4755 );
and AND2_1066 ( P1_U3762 , P1_U4758 , P1_U4757 );
and AND2_1067 ( P1_U3763 , P1_U4761 , P1_U4760 );
and AND2_1068 ( P1_U3764 , P1_U4763 , P1_U4762 );
and AND2_1069 ( P1_U3765 , P1_U4766 , P1_U4765 );
and AND2_1070 ( P1_U3766 , P1_U4768 , P1_U4767 );
and AND2_1071 ( P1_U3767 , P1_U4771 , P1_U4770 );
and AND2_1072 ( P1_U3768 , P1_U4773 , P1_U4772 );
and AND2_1073 ( P1_U3769 , P1_U4776 , P1_U4775 );
and AND2_1074 ( P1_U3770 , P1_U4778 , P1_U4777 );
and AND2_1075 ( P1_U3771 , P1_U4781 , P1_U4780 );
and AND3_1076 ( P1_U3772 , P1_U4783 , P1_U4782 , P1_U4784 );
and AND2_1077 ( P1_U3773 , P1_U4786 , P1_U4785 );
and AND3_1078 ( P1_U3774 , P1_U4788 , P1_U4787 , P1_U4789 );
and AND2_1079 ( P1_U3775 , P1_U4791 , P1_U4790 );
and AND3_1080 ( P1_U3776 , P1_U4793 , P1_U4792 , P1_U4794 );
and AND2_1081 ( P1_U3777 , P1_U4796 , P1_U4795 );
and AND5_1082 ( P1_U3778 , P1_U4798 , P1_U4797 , P1_U4799 , P1_U4800 , P1_U4801 );
and AND5_1083 ( P1_U3779 , P1_U4803 , P1_U4802 , P1_U4804 , P1_U4805 , P1_U4806 );
and AND5_1084 ( P1_U3780 , P1_U4808 , P1_U4807 , P1_U4809 , P1_U4810 , P1_U4811 );
and AND5_1085 ( P1_U3781 , P1_U4813 , P1_U4812 , P1_U4814 , P1_U4815 , P1_U4816 );
and AND5_1086 ( P1_U3782 , P1_U4818 , P1_U4817 , P1_U4819 , P1_U4820 , P1_U4821 );
and AND5_1087 ( P1_U3783 , P1_U4823 , P1_U4822 , P1_U4824 , P1_U4825 , P1_U4826 );
and AND3_1088 ( P1_U3784 , P1_U4828 , P1_U4827 , P1_U4829 );
and AND2_1089 ( P1_U3785 , P1_U4831 , P1_U4830 );
and AND5_1090 ( P1_U3786 , P1_U4833 , P1_U4832 , P1_U4834 , P1_U4835 , P1_U4836 );
and AND3_1091 ( P1_U3787 , P1_U4838 , P1_U4837 , P1_U4839 );
and AND2_1092 ( P1_U3788 , P1_U4841 , P1_U4840 );
and AND3_1093 ( P1_U3789 , P1_U4843 , P1_U4842 , P1_U4844 );
and AND2_1094 ( P1_U3790 , P1_U4846 , P1_U4845 );
and AND2_1095 ( P1_U3791 , P1_U4848 , P1_U4847 );
and AND2_1096 ( P1_U3792 , P1_U4851 , P1_U4850 );
and AND2_1097 ( P1_U3793 , P1_U4853 , P1_U4852 );
and AND2_1098 ( P1_U3794 , P1_U4856 , P1_U4855 );
and AND2_1099 ( P1_U3795 , P1_U4858 , P1_U4857 );
and AND2_1100 ( P1_U3796 , P1_U4861 , P1_U4860 );
and AND2_1101 ( P1_U3797 , P1_U4863 , P1_U4862 );
and AND2_1102 ( P1_U3798 , P1_U4866 , P1_U4865 );
and AND2_1103 ( P1_U3799 , P1_U4868 , P1_U4867 );
and AND2_1104 ( P1_U3800 , P1_U4871 , P1_U4870 );
and AND3_1105 ( P1_U3801 , P1_U5657 , P1_U4707 , P1_U5658 );
and AND2_1106 ( P1_U3802 , P1_U5660 , P1_U5659 );
and AND3_1107 ( P1_U3803 , P1_U3419 , P1_U3370 , P1_U3366 );
and AND3_1108 ( P1_U3804 , P1_U3368 , P1_U3365 , P1_U3361 );
and AND2_1109 ( P1_U3805 , P1_U3362 , P1_U3364 );
and AND2_1110 ( P1_U3806 , P1_U3805 , P1_U3420 );
and AND2_1111 ( P1_U3807 , P1_U3438 , P1_STATE_REG );
and AND2_1112 ( P1_U3808 , P1_U4891 , P1_U4892 );
and AND3_1113 ( P1_U3809 , P1_U4895 , P1_U4893 , P1_U4894 );
and AND2_1114 ( P1_U3810 , P1_U4901 , P1_U4902 );
and AND3_1115 ( P1_U3811 , P1_U4905 , P1_U4903 , P1_U4904 );
and AND2_1116 ( P1_U3812 , P1_U4911 , P1_U4912 );
and AND3_1117 ( P1_U3813 , P1_U4915 , P1_U4913 , P1_U4914 );
and AND2_1118 ( P1_U3814 , P1_U4921 , P1_U4922 );
and AND3_1119 ( P1_U3815 , P1_U4925 , P1_U4923 , P1_U4924 );
and AND2_1120 ( P1_U3816 , P1_U4931 , P1_U4932 );
and AND3_1121 ( P1_U3817 , P1_U4935 , P1_U4933 , P1_U4934 );
and AND2_1122 ( P1_U3818 , P1_U4941 , P1_U4942 );
and AND3_1123 ( P1_U3819 , P1_U4945 , P1_U4943 , P1_U4944 );
and AND2_1124 ( P1_U3820 , P1_U4951 , P1_U4952 );
and AND3_1125 ( P1_U3821 , P1_U4955 , P1_U4953 , P1_U4954 );
and AND2_1126 ( P1_U3822 , P1_U4961 , P1_U4962 );
and AND3_1127 ( P1_U3823 , P1_U4965 , P1_U4963 , P1_U4964 );
and AND2_1128 ( P1_U3824 , P1_U4971 , P1_U4972 );
and AND3_1129 ( P1_U3825 , P1_U4975 , P1_U4973 , P1_U4974 );
and AND2_1130 ( P1_U3826 , P1_U4981 , P1_U4982 );
and AND3_1131 ( P1_U3827 , P1_U4985 , P1_U4983 , P1_U4984 );
and AND2_1132 ( P1_U3828 , P1_U4991 , P1_U4992 );
and AND3_1133 ( P1_U3829 , P1_U4995 , P1_U4993 , P1_U4994 );
and AND2_1134 ( P1_U3830 , P1_U5001 , P1_U5002 );
and AND3_1135 ( P1_U3831 , P1_U5005 , P1_U5003 , P1_U5004 );
and AND2_1136 ( P1_U3832 , P1_U5011 , P1_U5012 );
and AND3_1137 ( P1_U3833 , P1_U5014 , P1_U5013 , P1_U5015 );
and AND3_1138 ( P1_U3834 , P1_U5021 , P1_U5022 , P1_U5020 );
and AND3_1139 ( P1_U3835 , P1_U5024 , P1_U5023 , P1_U5025 );
and AND3_1140 ( P1_U3836 , P1_U5031 , P1_U5032 , P1_U5030 );
and AND3_1141 ( P1_U3837 , P1_U5034 , P1_U5033 , P1_U5035 );
and AND2_1142 ( P1_U3838 , P1_U5040 , P1_U3998 );
and AND3_1143 ( P1_U3839 , P1_U5042 , P1_U5041 , P1_U3838 );
and AND3_1144 ( P1_U3840 , P1_U5044 , P1_U5043 , P1_U5045 );
and AND3_1145 ( P1_U3841 , P1_U5051 , P1_U5052 , P1_U5050 );
and AND3_1146 ( P1_U3842 , P1_U5054 , P1_U5053 , P1_U5055 );
and AND2_1147 ( P1_U3843 , P1_U5060 , P1_U3998 );
and AND3_1148 ( P1_U3844 , P1_U5062 , P1_U5061 , P1_U3843 );
and AND3_1149 ( P1_U3845 , P1_U5064 , P1_U5063 , P1_U5065 );
and AND3_1150 ( P1_U3846 , P1_U5071 , P1_U5072 , P1_U5070 );
and AND3_1151 ( P1_U3847 , P1_U5074 , P1_U5073 , P1_U5075 );
and AND3_1152 ( P1_U3848 , P1_U5081 , P1_U5082 , P1_U5080 );
and AND3_1153 ( P1_U3849 , P1_U5084 , P1_U5083 , P1_U5085 );
and AND2_1154 ( P1_U3850 , P1_STATE_REG , P1_U3428 );
and AND2_1155 ( P1_U3851 , P1_U3850 , P1_U3424 );
and AND3_1156 ( P1_U3852 , P1_U6114 , P1_U6111 , P1_U6117 );
and AND3_1157 ( P1_U3853 , P1_U3854 , P1_U3852 , P1_U6129 );
and AND3_1158 ( P1_U3854 , P1_U6126 , P1_U6123 , P1_U6120 );
and AND3_1159 ( P1_U3855 , P1_U6138 , P1_U6135 , P1_U6141 );
and AND3_1160 ( P1_U3856 , P1_U6147 , P1_U6144 , P1_U6150 );
and AND3_1161 ( P1_U3857 , P1_U3856 , P1_U3855 , P1_U6132 );
and AND5_1162 ( P1_U3858 , P1_U3863 , P1_U3862 , P1_U6081 , P1_U6078 , P1_U6075 );
and AND5_1163 ( P1_U3859 , P1_U6165 , P1_U6162 , P1_U6159 , P1_U6156 , P1_U6168 );
and AND5_1164 ( P1_U3860 , P1_U3857 , P1_U3853 , P1_U6108 , P1_U6153 , P1_U3859 );
and AND2_1165 ( P1_U3861 , P1_U6102 , P1_U3858 );
and AND4_1166 ( P1_U3862 , P1_U6093 , P1_U6090 , P1_U6087 , P1_U6084 );
and AND2_1167 ( P1_U3863 , P1_U6099 , P1_U6096 );
and AND3_1168 ( P1_U3864 , P1_U5090 , P1_U5091 , P1_U5087 );
and AND2_1169 ( P1_U3865 , P1_U3052 , P1_U5690 );
and AND2_1170 ( P1_U3866 , P1_U5651 , P1_U5652 );
and AND2_1171 ( P1_U3867 , P1_U3451 , P1_U3452 );
and AND3_1172 ( P1_U3868 , P1_U3371 , P1_U3369 , P1_U3420 );
and AND2_1173 ( P1_U3869 , P1_U5677 , P1_U3969 );
and AND2_1174 ( P1_U3870 , P1_U3424 , P1_U3869 );
and AND2_1175 ( P1_U3871 , P1_U3022 , P1_U5100 );
and AND2_1176 ( P1_U3872 , P1_U5147 , P1_U5146 );
and AND2_1177 ( P1_U3873 , P1_U3994 , P1_U3078 );
and AND2_1178 ( P1_U3874 , P1_U5188 , P1_U5187 );
and AND2_1179 ( P1_U3875 , P1_U5191 , P1_U5190 );
and AND2_1180 ( P1_U3876 , P1_U5281 , P1_U5280 );
and AND2_1181 ( P1_U3877 , P1_U3433 , P1_U5366 );
and AND2_1182 ( P1_U3878 , P1_U5431 , P1_U5432 );
and AND2_1183 ( P1_U3879 , P1_U5514 , P1_U3438 );
and AND2_1184 ( P1_U3880 , P1_U5516 , P1_U3438 );
and AND2_1185 ( P1_U3881 , P1_U5518 , P1_U3438 );
and AND2_1186 ( P1_U3882 , P1_U5520 , P1_U3438 );
and AND2_1187 ( P1_U3883 , P1_U5522 , P1_U3438 );
and AND2_1188 ( P1_U3884 , P1_U5524 , P1_U3438 );
and AND2_1189 ( P1_U3885 , P1_U5526 , P1_U3438 );
and AND2_1190 ( P1_U3886 , P1_U5528 , P1_U3438 );
and AND2_1191 ( P1_U3887 , P1_U5530 , P1_U3438 );
and AND2_1192 ( P1_U3888 , P1_U3438 , P1_U5533 );
and AND2_1193 ( P1_U3889 , P1_U3438 , P1_U5535 );
and AND2_1194 ( P1_U3890 , P1_U3438 , P1_U5537 );
and AND2_1195 ( P1_U3891 , P1_U3438 , P1_U5539 );
and AND2_1196 ( P1_U3892 , P1_U3438 , P1_U5541 );
and AND2_1197 ( P1_U3893 , P1_U3438 , P1_U5543 );
and AND2_1198 ( P1_U3894 , P1_U3438 , P1_U5555 );
and AND2_1199 ( P1_U3895 , P1_U5587 , P1_U5585 );
and AND2_1200 ( P1_U3896 , P1_U5590 , P1_U5588 );
and AND2_1201 ( P1_U3897 , P1_U5593 , P1_U5591 );
and AND2_1202 ( P1_U3898 , P1_U5596 , P1_U5594 );
and AND2_1203 ( P1_U3899 , P1_U5599 , P1_U5597 );
and AND2_1204 ( P1_U3900 , P1_U5602 , P1_U5600 );
and AND2_1205 ( P1_U3901 , P1_U5605 , P1_U5603 );
and AND2_1206 ( P1_U3902 , P1_U5608 , P1_U5606 );
and AND2_1207 ( P1_U3903 , P1_U5611 , P1_U5609 );
and AND2_1208 ( P1_U3904 , P1_U5617 , P1_U5615 );
and AND2_1209 ( P1_U3905 , P1_U5620 , P1_U5618 );
and AND2_1210 ( P1_U3906 , P1_U5623 , P1_U5621 );
and AND2_1211 ( P1_U3907 , P1_U5626 , P1_U5624 );
and AND2_1212 ( P1_U3908 , P1_U5629 , P1_U5627 );
and AND2_1213 ( P1_U3909 , P1_U5632 , P1_U5630 );
not NOT1_1214 ( P1_U3910 , P1_IR_REG_31_ );
nand NAND2_1215 ( P1_U3911 , P1_U3022 , P1_U3360 );
nand NAND2_1216 ( P1_U3912 , P1_U5702 , P1_U5699 );
nand NAND2_1217 ( P1_U3913 , P1_U3632 , P1_U3047 );
nand NAND2_1218 ( P1_U3914 , P1_U3748 , P1_U3047 );
and AND2_1219 ( P1_U3915 , P1_U5942 , P1_U5941 );
and AND2_1220 ( P1_U3916 , P1_U5944 , P1_U5943 );
and AND2_1221 ( P1_U3917 , P1_U5946 , P1_U5945 );
and AND2_1222 ( P1_U3918 , P1_U5948 , P1_U5947 );
and AND2_1223 ( P1_U3919 , P1_U5950 , P1_U5949 );
and AND2_1224 ( P1_U3920 , P1_U5952 , P1_U5951 );
and AND2_1225 ( P1_U3921 , P1_U5954 , P1_U5953 );
and AND2_1226 ( P1_U3922 , P1_U5956 , P1_U5955 );
and AND2_1227 ( P1_U3923 , P1_U5958 , P1_U5957 );
and AND2_1228 ( P1_U3924 , P1_U5960 , P1_U5959 );
and AND2_1229 ( P1_U3925 , P1_U5962 , P1_U5961 );
and AND2_1230 ( P1_U3926 , P1_U5964 , P1_U5963 );
and AND2_1231 ( P1_U3927 , P1_U5966 , P1_U5965 );
and AND2_1232 ( P1_U3928 , P1_U5968 , P1_U5967 );
and AND2_1233 ( P1_U3929 , P1_U5970 , P1_U5969 );
and AND2_1234 ( P1_U3930 , P1_U5972 , P1_U5971 );
and AND2_1235 ( P1_U3931 , P1_U5974 , P1_U5973 );
and AND2_1236 ( P1_U3932 , P1_U5976 , P1_U5975 );
and AND2_1237 ( P1_U3933 , P1_U5978 , P1_U5977 );
and AND2_1238 ( P1_U3934 , P1_U5980 , P1_U5979 );
and AND2_1239 ( P1_U3935 , P1_U5982 , P1_U5981 );
and AND2_1240 ( P1_U3936 , P1_U5984 , P1_U5983 );
and AND2_1241 ( P1_U3937 , P1_U5986 , P1_U5985 );
and AND2_1242 ( P1_U3938 , P1_U5988 , P1_U5987 );
and AND2_1243 ( P1_U3939 , P1_U5990 , P1_U5989 );
and AND2_1244 ( P1_U3940 , P1_U5992 , P1_U5991 );
and AND2_1245 ( P1_U3941 , P1_U5994 , P1_U5993 );
and AND2_1246 ( P1_U3942 , P1_U5996 , P1_U5995 );
and AND2_1247 ( P1_U3943 , P1_U5998 , P1_U5997 );
and AND2_1248 ( P1_U3944 , P1_U6000 , P1_U5999 );
nand NAND2_1249 ( P1_U3945 , P1_U3747 , P1_U3056 );
and AND2_1250 ( P1_U3946 , P1_U6002 , P1_U6001 );
and AND2_1251 ( P1_U3947 , P1_U6004 , P1_U6003 );
not NOT1_1252 ( P1_U3948 , P1_R1375_U14 );
not NOT1_1253 ( P1_U3949 , P1_R1360_U14 );
and AND2_1254 ( P1_U3950 , P1_U6072 , P1_U6071 );
nand NAND3_1255 ( P1_U3951 , P1_U3860 , P1_U6105 , P1_U3861 );
not NOT1_1256 ( P1_U3952 , P1_R1352_U6 );
not NOT1_1257 ( P1_U3953 , P1_U3372 );
not NOT1_1258 ( P1_U3954 , P1_U3426 );
not NOT1_1259 ( P1_U3955 , P1_U3428 );
not NOT1_1260 ( P1_U3956 , P1_U3370 );
not NOT1_1261 ( P1_U3957 , P1_U3419 );
not NOT1_1262 ( P1_U3958 , P1_U3366 );
not NOT1_1263 ( P1_U3959 , P1_U3365 );
not NOT1_1264 ( P1_U3960 , P1_U3368 );
not NOT1_1265 ( P1_U3961 , P1_U3361 );
not NOT1_1266 ( P1_U3962 , P1_U3364 );
not NOT1_1267 ( P1_U3963 , P1_U3362 );
not NOT1_1268 ( P1_U3964 , P1_U3420 );
not NOT1_1269 ( P1_U3965 , P1_U3418 );
nand NAND2_1270 ( P1_U3966 , P1_U3049 , P1_U4001 );
not NOT1_1271 ( P1_U3967 , P1_U3371 );
not NOT1_1272 ( P1_U3968 , P1_U3369 );
nand NAND2_1273 ( P1_U3969 , P1_U3987 , P1_U3367 );
nand NAND2_1274 ( P1_U3970 , P1_U3049 , P1_U3421 );
not NOT1_1275 ( P1_U3971 , P1_U3912 );
not NOT1_1276 ( P1_U3972 , P1_U3430 );
not NOT1_1277 ( P1_U3973 , P1_U3425 );
not NOT1_1278 ( P1_U3974 , P1_U3411 );
not NOT1_1279 ( P1_U3975 , P1_U3409 );
not NOT1_1280 ( P1_U3976 , P1_U3407 );
not NOT1_1281 ( P1_U3977 , P1_U3405 );
not NOT1_1282 ( P1_U3978 , P1_U3403 );
not NOT1_1283 ( P1_U3979 , P1_U3401 );
not NOT1_1284 ( P1_U3980 , P1_U3399 );
not NOT1_1285 ( P1_U3981 , P1_U3397 );
not NOT1_1286 ( P1_U3982 , P1_U3395 );
not NOT1_1287 ( P1_U3983 , P1_U3415 );
not NOT1_1288 ( P1_U3984 , P1_U3414 );
not NOT1_1289 ( P1_U3985 , P1_U3413 );
not NOT1_1290 ( P1_U3986 , P1_U3427 );
not NOT1_1291 ( P1_U3987 , P1_U3373 );
not NOT1_1292 ( P1_U3988 , P1_U3416 );
not NOT1_1293 ( P1_U3989 , P1_U3417 );
not NOT1_1294 ( P1_U3990 , P1_U3914 );
not NOT1_1295 ( P1_U3991 , P1_U3913 );
not NOT1_1296 ( P1_U3992 , P1_U3911 );
not NOT1_1297 ( P1_U3993 , P1_U3945 );
not NOT1_1298 ( P1_U3994 , P1_U3431 );
nand NAND2_1299 ( P1_U3995 , P1_U3432 , P1_STATE_REG );
nand NAND2_1300 ( P1_U3996 , P1_U3965 , P1_U3022 );
not NOT1_1301 ( P1_U3997 , P1_U3429 );
nand NAND2_1302 ( P1_U3998 , P1_U3973 , P1_U3212 );
not NOT1_1303 ( P1_U3999 , P1_U3424 );
not NOT1_1304 ( P1_U4000 , P1_U3433 );
not NOT1_1305 ( P1_U4001 , P1_U3363 );
not NOT1_1306 ( P1_U4002 , P1_U3367 );
not NOT1_1307 ( P1_U4003 , P1_U3358 );
not NOT1_1308 ( P1_U4004 , P1_U3357 );
nand NAND2_1309 ( P1_U4005 , U88 , P1_U3086 );
nand NAND2_1310 ( P1_U4006 , P1_IR_REG_0_ , P1_U3028 );
nand NAND2_1311 ( P1_U4007 , P1_IR_REG_0_ , P1_U4004 );
nand NAND2_1312 ( P1_U4008 , U77 , P1_U3086 );
nand NAND2_1313 ( P1_U4009 , P1_SUB_84_U40 , P1_U3028 );
nand NAND2_1314 ( P1_U4010 , P1_IR_REG_1_ , P1_U4004 );
nand NAND2_1315 ( P1_U4011 , U66 , P1_U3086 );
nand NAND2_1316 ( P1_U4012 , P1_SUB_84_U21 , P1_U3028 );
nand NAND2_1317 ( P1_U4013 , P1_IR_REG_2_ , P1_U4004 );
nand NAND2_1318 ( P1_U4014 , U63 , P1_U3086 );
nand NAND2_1319 ( P1_U4015 , P1_SUB_84_U22 , P1_U3028 );
nand NAND2_1320 ( P1_U4016 , P1_IR_REG_3_ , P1_U4004 );
nand NAND2_1321 ( P1_U4017 , U62 , P1_U3086 );
nand NAND2_1322 ( P1_U4018 , P1_SUB_84_U23 , P1_U3028 );
nand NAND2_1323 ( P1_U4019 , P1_IR_REG_4_ , P1_U4004 );
nand NAND2_1324 ( P1_U4020 , U61 , P1_U3086 );
nand NAND2_1325 ( P1_U4021 , P1_SUB_84_U162 , P1_U3028 );
nand NAND2_1326 ( P1_U4022 , P1_IR_REG_5_ , P1_U4004 );
nand NAND2_1327 ( P1_U4023 , U60 , P1_U3086 );
nand NAND2_1328 ( P1_U4024 , P1_SUB_84_U24 , P1_U3028 );
nand NAND2_1329 ( P1_U4025 , P1_IR_REG_6_ , P1_U4004 );
nand NAND2_1330 ( P1_U4026 , U59 , P1_U3086 );
nand NAND2_1331 ( P1_U4027 , P1_SUB_84_U25 , P1_U3028 );
nand NAND2_1332 ( P1_U4028 , P1_IR_REG_7_ , P1_U4004 );
nand NAND2_1333 ( P1_U4029 , U58 , P1_U3086 );
nand NAND2_1334 ( P1_U4030 , P1_SUB_84_U26 , P1_U3028 );
nand NAND2_1335 ( P1_U4031 , P1_IR_REG_8_ , P1_U4004 );
nand NAND2_1336 ( P1_U4032 , U57 , P1_U3086 );
nand NAND2_1337 ( P1_U4033 , P1_SUB_84_U160 , P1_U3028 );
nand NAND2_1338 ( P1_U4034 , P1_IR_REG_9_ , P1_U4004 );
nand NAND2_1339 ( P1_U4035 , U87 , P1_U3086 );
nand NAND2_1340 ( P1_U4036 , P1_SUB_84_U6 , P1_U3028 );
nand NAND2_1341 ( P1_U4037 , P1_IR_REG_10_ , P1_U4004 );
nand NAND2_1342 ( P1_U4038 , U86 , P1_U3086 );
nand NAND2_1343 ( P1_U4039 , P1_SUB_84_U7 , P1_U3028 );
nand NAND2_1344 ( P1_U4040 , P1_IR_REG_11_ , P1_U4004 );
nand NAND2_1345 ( P1_U4041 , U85 , P1_U3086 );
nand NAND2_1346 ( P1_U4042 , P1_SUB_84_U8 , P1_U3028 );
nand NAND2_1347 ( P1_U4043 , P1_IR_REG_12_ , P1_U4004 );
nand NAND2_1348 ( P1_U4044 , U84 , P1_U3086 );
nand NAND2_1349 ( P1_U4045 , P1_SUB_84_U179 , P1_U3028 );
nand NAND2_1350 ( P1_U4046 , P1_IR_REG_13_ , P1_U4004 );
nand NAND2_1351 ( P1_U4047 , U83 , P1_U3086 );
nand NAND2_1352 ( P1_U4048 , P1_SUB_84_U9 , P1_U3028 );
nand NAND2_1353 ( P1_U4049 , P1_IR_REG_14_ , P1_U4004 );
nand NAND2_1354 ( P1_U4050 , U82 , P1_U3086 );
nand NAND2_1355 ( P1_U4051 , P1_SUB_84_U10 , P1_U3028 );
nand NAND2_1356 ( P1_U4052 , P1_IR_REG_15_ , P1_U4004 );
nand NAND2_1357 ( P1_U4053 , U81 , P1_U3086 );
nand NAND2_1358 ( P1_U4054 , P1_SUB_84_U11 , P1_U3028 );
nand NAND2_1359 ( P1_U4055 , P1_IR_REG_16_ , P1_U4004 );
nand NAND2_1360 ( P1_U4056 , U80 , P1_U3086 );
nand NAND2_1361 ( P1_U4057 , P1_SUB_84_U177 , P1_U3028 );
nand NAND2_1362 ( P1_U4058 , P1_IR_REG_17_ , P1_U4004 );
nand NAND2_1363 ( P1_U4059 , U79 , P1_U3086 );
nand NAND2_1364 ( P1_U4060 , P1_SUB_84_U12 , P1_U3028 );
nand NAND2_1365 ( P1_U4061 , P1_IR_REG_18_ , P1_U4004 );
nand NAND2_1366 ( P1_U4062 , U78 , P1_U3086 );
nand NAND2_1367 ( P1_U4063 , P1_SUB_84_U13 , P1_U3028 );
nand NAND2_1368 ( P1_U4064 , P1_IR_REG_19_ , P1_U4004 );
nand NAND2_1369 ( P1_U4065 , U76 , P1_U3086 );
nand NAND2_1370 ( P1_U4066 , P1_SUB_84_U14 , P1_U3028 );
nand NAND2_1371 ( P1_U4067 , P1_IR_REG_20_ , P1_U4004 );
nand NAND2_1372 ( P1_U4068 , U75 , P1_U3086 );
nand NAND2_1373 ( P1_U4069 , P1_SUB_84_U173 , P1_U3028 );
nand NAND2_1374 ( P1_U4070 , P1_IR_REG_21_ , P1_U4004 );
nand NAND2_1375 ( P1_U4071 , U74 , P1_U3086 );
nand NAND2_1376 ( P1_U4072 , P1_SUB_84_U15 , P1_U3028 );
nand NAND2_1377 ( P1_U4073 , P1_IR_REG_22_ , P1_U4004 );
nand NAND2_1378 ( P1_U4074 , U73 , P1_U3086 );
nand NAND2_1379 ( P1_U4075 , P1_SUB_84_U16 , P1_U3028 );
nand NAND2_1380 ( P1_U4076 , P1_IR_REG_23_ , P1_U4004 );
nand NAND2_1381 ( P1_U4077 , U72 , P1_U3086 );
nand NAND2_1382 ( P1_U4078 , P1_SUB_84_U17 , P1_U3028 );
nand NAND2_1383 ( P1_U4079 , P1_IR_REG_24_ , P1_U4004 );
nand NAND2_1384 ( P1_U4080 , U71 , P1_U3086 );
nand NAND2_1385 ( P1_U4081 , P1_SUB_84_U170 , P1_U3028 );
nand NAND2_1386 ( P1_U4082 , P1_IR_REG_25_ , P1_U4004 );
nand NAND2_1387 ( P1_U4083 , U70 , P1_U3086 );
nand NAND2_1388 ( P1_U4084 , P1_SUB_84_U18 , P1_U3028 );
nand NAND2_1389 ( P1_U4085 , P1_IR_REG_26_ , P1_U4004 );
nand NAND2_1390 ( P1_U4086 , U69 , P1_U3086 );
nand NAND2_1391 ( P1_U4087 , P1_SUB_84_U42 , P1_U3028 );
nand NAND2_1392 ( P1_U4088 , P1_IR_REG_27_ , P1_U4004 );
nand NAND2_1393 ( P1_U4089 , U68 , P1_U3086 );
nand NAND2_1394 ( P1_U4090 , P1_SUB_84_U19 , P1_U3028 );
nand NAND2_1395 ( P1_U4091 , P1_IR_REG_28_ , P1_U4004 );
nand NAND2_1396 ( P1_U4092 , U67 , P1_U3086 );
nand NAND2_1397 ( P1_U4093 , P1_SUB_84_U20 , P1_U3028 );
nand NAND2_1398 ( P1_U4094 , P1_IR_REG_29_ , P1_U4004 );
nand NAND2_1399 ( P1_U4095 , U65 , P1_U3086 );
nand NAND2_1400 ( P1_U4096 , P1_SUB_84_U165 , P1_U3028 );
nand NAND2_1401 ( P1_U4097 , P1_IR_REG_30_ , P1_U4004 );
nand NAND2_1402 ( P1_U4098 , U64 , P1_U3086 );
nand NAND2_1403 ( P1_U4099 , P1_SUB_84_U41 , P1_U3028 );
nand NAND2_1404 ( P1_U4100 , P1_IR_REG_31_ , P1_U4004 );
not NOT1_1405 ( P1_U4101 , P1_U3360 );
not NOT1_1406 ( P1_U4102 , P1_U3421 );
nand NAND2_1407 ( P1_U4103 , P1_U3358 , P1_U5666 );
nand NAND2_1408 ( P1_U4104 , P1_U3358 , P1_U5669 );
nand NAND2_1409 ( P1_U4105 , P1_U4101 , P1_D_REG_10_ );
nand NAND2_1410 ( P1_U4106 , P1_U4101 , P1_D_REG_11_ );
nand NAND2_1411 ( P1_U4107 , P1_U4101 , P1_D_REG_12_ );
nand NAND2_1412 ( P1_U4108 , P1_U4101 , P1_D_REG_13_ );
nand NAND2_1413 ( P1_U4109 , P1_U4101 , P1_D_REG_14_ );
nand NAND2_1414 ( P1_U4110 , P1_U4101 , P1_D_REG_15_ );
nand NAND2_1415 ( P1_U4111 , P1_U4101 , P1_D_REG_16_ );
nand NAND2_1416 ( P1_U4112 , P1_U4101 , P1_D_REG_17_ );
nand NAND2_1417 ( P1_U4113 , P1_U4101 , P1_D_REG_18_ );
nand NAND2_1418 ( P1_U4114 , P1_U4101 , P1_D_REG_19_ );
nand NAND2_1419 ( P1_U4115 , P1_U4101 , P1_D_REG_20_ );
nand NAND2_1420 ( P1_U4116 , P1_U4101 , P1_D_REG_21_ );
nand NAND2_1421 ( P1_U4117 , P1_U4101 , P1_D_REG_22_ );
nand NAND2_1422 ( P1_U4118 , P1_U4101 , P1_D_REG_23_ );
nand NAND2_1423 ( P1_U4119 , P1_U4101 , P1_D_REG_24_ );
nand NAND2_1424 ( P1_U4120 , P1_U4101 , P1_D_REG_25_ );
nand NAND2_1425 ( P1_U4121 , P1_U4101 , P1_D_REG_26_ );
nand NAND2_1426 ( P1_U4122 , P1_U4101 , P1_D_REG_27_ );
nand NAND2_1427 ( P1_U4123 , P1_U4101 , P1_D_REG_28_ );
nand NAND2_1428 ( P1_U4124 , P1_U4101 , P1_D_REG_29_ );
nand NAND2_1429 ( P1_U4125 , P1_U4101 , P1_D_REG_2_ );
nand NAND2_1430 ( P1_U4126 , P1_U4101 , P1_D_REG_30_ );
nand NAND2_1431 ( P1_U4127 , P1_U4101 , P1_D_REG_31_ );
nand NAND2_1432 ( P1_U4128 , P1_U4101 , P1_D_REG_3_ );
nand NAND2_1433 ( P1_U4129 , P1_U4101 , P1_D_REG_4_ );
nand NAND2_1434 ( P1_U4130 , P1_U4101 , P1_D_REG_5_ );
nand NAND2_1435 ( P1_U4131 , P1_U4101 , P1_D_REG_6_ );
nand NAND2_1436 ( P1_U4132 , P1_U4101 , P1_D_REG_7_ );
nand NAND2_1437 ( P1_U4133 , P1_U4101 , P1_D_REG_8_ );
nand NAND2_1438 ( P1_U4134 , P1_U4101 , P1_D_REG_9_ );
nand NAND2_1439 ( P1_U4135 , P1_U5690 , P1_U5693 );
nand NAND3_1440 ( P1_U4136 , P1_U5713 , P1_U5712 , P1_U3367 );
nand NAND2_1441 ( P1_U4137 , P1_U3018 , P1_REG2_REG_1_ );
nand NAND2_1442 ( P1_U4138 , P1_U3019 , P1_REG1_REG_1_ );
nand NAND2_1443 ( P1_U4139 , P1_U3020 , P1_REG0_REG_1_ );
nand NAND2_1444 ( P1_U4140 , P1_REG3_REG_1_ , P1_U3017 );
not NOT1_1445 ( P1_U4141 , P1_U3078 );
nand NAND2_1446 ( P1_U4142 , P1_U3966 , P1_U3416 );
nand NAND2_1447 ( P1_U4143 , P1_U3961 , P1_R1150_U18 );
nand NAND2_1448 ( P1_U4144 , P1_U3963 , P1_R1117_U18 );
nand NAND2_1449 ( P1_U4145 , P1_U3962 , P1_R1138_U96 );
nand NAND2_1450 ( P1_U4146 , P1_U3959 , P1_R1192_U18 );
nand NAND2_1451 ( P1_U4147 , P1_U3958 , P1_R1207_U18 );
nand NAND2_1452 ( P1_U4148 , P1_U3968 , P1_R1171_U96 );
nand NAND2_1453 ( P1_U4149 , P1_U3967 , P1_R1240_U96 );
not NOT1_1454 ( P1_U4150 , P1_U3374 );
nand NAND2_1455 ( P1_U4151 , P1_R1222_U96 , P1_U3026 );
nand NAND2_1456 ( P1_U4152 , P1_U3025 , P1_U3078 );
nand NAND2_1457 ( P1_U4153 , P1_U3450 , P1_U3023 );
nand NAND2_1458 ( P1_U4154 , P1_U3450 , P1_U4142 );
nand NAND2_1459 ( P1_U4155 , P1_U3620 , P1_U4150 );
nand NAND2_1460 ( P1_U4156 , P1_REG2_REG_2_ , P1_U3018 );
nand NAND2_1461 ( P1_U4157 , P1_REG1_REG_2_ , P1_U3019 );
nand NAND2_1462 ( P1_U4158 , P1_REG0_REG_2_ , P1_U3020 );
nand NAND2_1463 ( P1_U4159 , P1_REG3_REG_2_ , P1_U3017 );
not NOT1_1464 ( P1_U4160 , P1_U3068 );
nand NAND2_1465 ( P1_U4161 , P1_REG0_REG_0_ , P1_U3020 );
nand NAND2_1466 ( P1_U4162 , P1_REG1_REG_0_ , P1_U3019 );
nand NAND2_1467 ( P1_U4163 , P1_REG2_REG_0_ , P1_U3018 );
nand NAND2_1468 ( P1_U4164 , P1_REG3_REG_0_ , P1_U3017 );
not NOT1_1469 ( P1_U4165 , P1_U3077 );
nand NAND2_1470 ( P1_U4166 , P1_U3033 , P1_U3077 );
nand NAND2_1471 ( P1_U4167 , P1_R1150_U96 , P1_U3961 );
nand NAND2_1472 ( P1_U4168 , P1_R1117_U96 , P1_U3963 );
nand NAND2_1473 ( P1_U4169 , P1_R1138_U95 , P1_U3962 );
nand NAND2_1474 ( P1_U4170 , P1_R1192_U96 , P1_U3959 );
nand NAND2_1475 ( P1_U4171 , P1_R1207_U96 , P1_U3958 );
nand NAND2_1476 ( P1_U4172 , P1_R1171_U95 , P1_U3968 );
nand NAND2_1477 ( P1_U4173 , P1_R1240_U95 , P1_U3967 );
not NOT1_1478 ( P1_U4174 , P1_U3376 );
nand NAND2_1479 ( P1_U4175 , P1_R1222_U95 , P1_U3026 );
nand NAND2_1480 ( P1_U4176 , P1_U3025 , P1_U3068 );
nand NAND2_1481 ( P1_U4177 , P1_R1282_U57 , P1_U3023 );
nand NAND2_1482 ( P1_U4178 , P1_U3455 , P1_U4142 );
nand NAND2_1483 ( P1_U4179 , P1_U3636 , P1_U4174 );
nand NAND2_1484 ( P1_U4180 , P1_REG2_REG_3_ , P1_U3018 );
nand NAND2_1485 ( P1_U4181 , P1_REG1_REG_3_ , P1_U3019 );
nand NAND2_1486 ( P1_U4182 , P1_REG0_REG_3_ , P1_U3020 );
nand NAND2_1487 ( P1_U4183 , P1_ADD_95_U4 , P1_U3017 );
not NOT1_1488 ( P1_U4184 , P1_U3064 );
nand NAND2_1489 ( P1_U4185 , P1_U3033 , P1_U3078 );
nand NAND2_1490 ( P1_U4186 , P1_R1150_U106 , P1_U3961 );
nand NAND2_1491 ( P1_U4187 , P1_R1117_U106 , P1_U3963 );
nand NAND2_1492 ( P1_U4188 , P1_R1138_U17 , P1_U3962 );
nand NAND2_1493 ( P1_U4189 , P1_R1192_U106 , P1_U3959 );
nand NAND2_1494 ( P1_U4190 , P1_R1207_U106 , P1_U3958 );
nand NAND2_1495 ( P1_U4191 , P1_R1171_U17 , P1_U3968 );
nand NAND2_1496 ( P1_U4192 , P1_R1240_U17 , P1_U3967 );
not NOT1_1497 ( P1_U4193 , P1_U3377 );
nand NAND2_1498 ( P1_U4194 , P1_R1222_U17 , P1_U3026 );
nand NAND2_1499 ( P1_U4195 , P1_U3025 , P1_U3064 );
nand NAND2_1500 ( P1_U4196 , P1_R1282_U18 , P1_U3023 );
nand NAND2_1501 ( P1_U4197 , P1_U3458 , P1_U4142 );
nand NAND2_1502 ( P1_U4198 , P1_U3640 , P1_U4193 );
nand NAND2_1503 ( P1_U4199 , P1_REG2_REG_4_ , P1_U3018 );
nand NAND2_1504 ( P1_U4200 , P1_REG1_REG_4_ , P1_U3019 );
nand NAND2_1505 ( P1_U4201 , P1_REG0_REG_4_ , P1_U3020 );
nand NAND2_1506 ( P1_U4202 , P1_ADD_95_U59 , P1_U3017 );
not NOT1_1507 ( P1_U4203 , P1_U3060 );
nand NAND2_1508 ( P1_U4204 , P1_U3033 , P1_U3068 );
nand NAND2_1509 ( P1_U4205 , P1_R1150_U15 , P1_U3961 );
nand NAND2_1510 ( P1_U4206 , P1_R1117_U15 , P1_U3963 );
nand NAND2_1511 ( P1_U4207 , P1_R1138_U101 , P1_U3962 );
nand NAND2_1512 ( P1_U4208 , P1_R1192_U15 , P1_U3959 );
nand NAND2_1513 ( P1_U4209 , P1_R1207_U15 , P1_U3958 );
nand NAND2_1514 ( P1_U4210 , P1_R1171_U101 , P1_U3968 );
nand NAND2_1515 ( P1_U4211 , P1_R1240_U101 , P1_U3967 );
not NOT1_1516 ( P1_U4212 , P1_U3378 );
nand NAND2_1517 ( P1_U4213 , P1_R1222_U101 , P1_U3026 );
nand NAND2_1518 ( P1_U4214 , P1_U3025 , P1_U3060 );
nand NAND2_1519 ( P1_U4215 , P1_R1282_U20 , P1_U3023 );
nand NAND2_1520 ( P1_U4216 , P1_U3461 , P1_U4142 );
nand NAND2_1521 ( P1_U4217 , P1_U3643 , P1_U4212 );
nand NAND2_1522 ( P1_U4218 , P1_REG2_REG_5_ , P1_U3018 );
nand NAND2_1523 ( P1_U4219 , P1_REG1_REG_5_ , P1_U3019 );
nand NAND2_1524 ( P1_U4220 , P1_REG0_REG_5_ , P1_U3020 );
nand NAND2_1525 ( P1_U4221 , P1_ADD_95_U58 , P1_U3017 );
not NOT1_1526 ( P1_U4222 , P1_U3067 );
nand NAND2_1527 ( P1_U4223 , P1_U3033 , P1_U3064 );
nand NAND2_1528 ( P1_U4224 , P1_R1150_U105 , P1_U3961 );
nand NAND2_1529 ( P1_U4225 , P1_R1117_U105 , P1_U3963 );
nand NAND2_1530 ( P1_U4226 , P1_R1138_U100 , P1_U3962 );
nand NAND2_1531 ( P1_U4227 , P1_R1192_U105 , P1_U3959 );
nand NAND2_1532 ( P1_U4228 , P1_R1207_U105 , P1_U3958 );
nand NAND2_1533 ( P1_U4229 , P1_R1171_U100 , P1_U3968 );
nand NAND2_1534 ( P1_U4230 , P1_R1240_U100 , P1_U3967 );
not NOT1_1535 ( P1_U4231 , P1_U3379 );
nand NAND2_1536 ( P1_U4232 , P1_R1222_U100 , P1_U3026 );
nand NAND2_1537 ( P1_U4233 , P1_U3025 , P1_U3067 );
nand NAND2_1538 ( P1_U4234 , P1_R1282_U21 , P1_U3023 );
nand NAND2_1539 ( P1_U4235 , P1_U3464 , P1_U4142 );
nand NAND2_1540 ( P1_U4236 , P1_U3646 , P1_U4231 );
nand NAND2_1541 ( P1_U4237 , P1_REG2_REG_6_ , P1_U3018 );
nand NAND2_1542 ( P1_U4238 , P1_REG1_REG_6_ , P1_U3019 );
nand NAND2_1543 ( P1_U4239 , P1_REG0_REG_6_ , P1_U3020 );
nand NAND2_1544 ( P1_U4240 , P1_ADD_95_U57 , P1_U3017 );
not NOT1_1545 ( P1_U4241 , P1_U3071 );
nand NAND2_1546 ( P1_U4242 , P1_U3033 , P1_U3060 );
nand NAND2_1547 ( P1_U4243 , P1_R1150_U104 , P1_U3961 );
nand NAND2_1548 ( P1_U4244 , P1_R1117_U104 , P1_U3963 );
nand NAND2_1549 ( P1_U4245 , P1_R1138_U18 , P1_U3962 );
nand NAND2_1550 ( P1_U4246 , P1_R1192_U104 , P1_U3959 );
nand NAND2_1551 ( P1_U4247 , P1_R1207_U104 , P1_U3958 );
nand NAND2_1552 ( P1_U4248 , P1_R1171_U18 , P1_U3968 );
nand NAND2_1553 ( P1_U4249 , P1_R1240_U18 , P1_U3967 );
not NOT1_1554 ( P1_U4250 , P1_U3380 );
nand NAND2_1555 ( P1_U4251 , P1_R1222_U18 , P1_U3026 );
nand NAND2_1556 ( P1_U4252 , P1_U3025 , P1_U3071 );
nand NAND2_1557 ( P1_U4253 , P1_R1282_U65 , P1_U3023 );
nand NAND2_1558 ( P1_U4254 , P1_U3467 , P1_U4142 );
nand NAND2_1559 ( P1_U4255 , P1_U3650 , P1_U4250 );
nand NAND2_1560 ( P1_U4256 , P1_REG2_REG_7_ , P1_U3018 );
nand NAND2_1561 ( P1_U4257 , P1_REG1_REG_7_ , P1_U3019 );
nand NAND2_1562 ( P1_U4258 , P1_REG0_REG_7_ , P1_U3020 );
nand NAND2_1563 ( P1_U4259 , P1_ADD_95_U56 , P1_U3017 );
not NOT1_1564 ( P1_U4260 , P1_U3070 );
nand NAND2_1565 ( P1_U4261 , P1_U3033 , P1_U3067 );
nand NAND2_1566 ( P1_U4262 , P1_R1150_U16 , P1_U3961 );
nand NAND2_1567 ( P1_U4263 , P1_R1117_U16 , P1_U3963 );
nand NAND2_1568 ( P1_U4264 , P1_R1138_U99 , P1_U3962 );
nand NAND2_1569 ( P1_U4265 , P1_R1192_U16 , P1_U3959 );
nand NAND2_1570 ( P1_U4266 , P1_R1207_U16 , P1_U3958 );
nand NAND2_1571 ( P1_U4267 , P1_R1171_U99 , P1_U3968 );
nand NAND2_1572 ( P1_U4268 , P1_R1240_U99 , P1_U3967 );
not NOT1_1573 ( P1_U4269 , P1_U3381 );
nand NAND2_1574 ( P1_U4270 , P1_R1222_U99 , P1_U3026 );
nand NAND2_1575 ( P1_U4271 , P1_U3025 , P1_U3070 );
nand NAND2_1576 ( P1_U4272 , P1_R1282_U22 , P1_U3023 );
nand NAND2_1577 ( P1_U4273 , P1_U3470 , P1_U4142 );
nand NAND2_1578 ( P1_U4274 , P1_U3654 , P1_U4269 );
nand NAND2_1579 ( P1_U4275 , P1_REG2_REG_8_ , P1_U3018 );
nand NAND2_1580 ( P1_U4276 , P1_REG1_REG_8_ , P1_U3019 );
nand NAND2_1581 ( P1_U4277 , P1_REG0_REG_8_ , P1_U3020 );
nand NAND2_1582 ( P1_U4278 , P1_ADD_95_U55 , P1_U3017 );
not NOT1_1583 ( P1_U4279 , P1_U3084 );
nand NAND2_1584 ( P1_U4280 , P1_U3033 , P1_U3071 );
nand NAND2_1585 ( P1_U4281 , P1_R1150_U103 , P1_U3961 );
nand NAND2_1586 ( P1_U4282 , P1_R1117_U103 , P1_U3963 );
nand NAND2_1587 ( P1_U4283 , P1_R1138_U19 , P1_U3962 );
nand NAND2_1588 ( P1_U4284 , P1_R1192_U103 , P1_U3959 );
nand NAND2_1589 ( P1_U4285 , P1_R1207_U103 , P1_U3958 );
nand NAND2_1590 ( P1_U4286 , P1_R1171_U19 , P1_U3968 );
nand NAND2_1591 ( P1_U4287 , P1_R1240_U19 , P1_U3967 );
not NOT1_1592 ( P1_U4288 , P1_U3382 );
nand NAND2_1593 ( P1_U4289 , P1_R1222_U19 , P1_U3026 );
nand NAND2_1594 ( P1_U4290 , P1_U3025 , P1_U3084 );
nand NAND2_1595 ( P1_U4291 , P1_R1282_U23 , P1_U3023 );
nand NAND2_1596 ( P1_U4292 , P1_U3473 , P1_U4142 );
nand NAND2_1597 ( P1_U4293 , P1_U3658 , P1_U4288 );
nand NAND2_1598 ( P1_U4294 , P1_REG2_REG_9_ , P1_U3018 );
nand NAND2_1599 ( P1_U4295 , P1_REG1_REG_9_ , P1_U3019 );
nand NAND2_1600 ( P1_U4296 , P1_REG0_REG_9_ , P1_U3020 );
nand NAND2_1601 ( P1_U4297 , P1_ADD_95_U54 , P1_U3017 );
not NOT1_1602 ( P1_U4298 , P1_U3083 );
nand NAND2_1603 ( P1_U4299 , P1_U3033 , P1_U3070 );
nand NAND2_1604 ( P1_U4300 , P1_R1150_U17 , P1_U3961 );
nand NAND2_1605 ( P1_U4301 , P1_R1117_U17 , P1_U3963 );
nand NAND2_1606 ( P1_U4302 , P1_R1138_U98 , P1_U3962 );
nand NAND2_1607 ( P1_U4303 , P1_R1192_U17 , P1_U3959 );
nand NAND2_1608 ( P1_U4304 , P1_R1207_U17 , P1_U3958 );
nand NAND2_1609 ( P1_U4305 , P1_R1171_U98 , P1_U3968 );
nand NAND2_1610 ( P1_U4306 , P1_R1240_U98 , P1_U3967 );
not NOT1_1611 ( P1_U4307 , P1_U3383 );
nand NAND2_1612 ( P1_U4308 , P1_R1222_U98 , P1_U3026 );
nand NAND2_1613 ( P1_U4309 , P1_U3025 , P1_U3083 );
nand NAND2_1614 ( P1_U4310 , P1_R1282_U24 , P1_U3023 );
nand NAND2_1615 ( P1_U4311 , P1_U3476 , P1_U4142 );
nand NAND2_1616 ( P1_U4312 , P1_U3662 , P1_U4307 );
nand NAND2_1617 ( P1_U4313 , P1_REG2_REG_10_ , P1_U3018 );
nand NAND2_1618 ( P1_U4314 , P1_REG1_REG_10_ , P1_U3019 );
nand NAND2_1619 ( P1_U4315 , P1_REG0_REG_10_ , P1_U3020 );
nand NAND2_1620 ( P1_U4316 , P1_ADD_95_U78 , P1_U3017 );
not NOT1_1621 ( P1_U4317 , P1_U3062 );
nand NAND2_1622 ( P1_U4318 , P1_U3033 , P1_U3084 );
nand NAND2_1623 ( P1_U4319 , P1_R1150_U102 , P1_U3961 );
nand NAND2_1624 ( P1_U4320 , P1_R1117_U102 , P1_U3963 );
nand NAND2_1625 ( P1_U4321 , P1_R1138_U97 , P1_U3962 );
nand NAND2_1626 ( P1_U4322 , P1_R1192_U102 , P1_U3959 );
nand NAND2_1627 ( P1_U4323 , P1_R1207_U102 , P1_U3958 );
nand NAND2_1628 ( P1_U4324 , P1_R1171_U97 , P1_U3968 );
nand NAND2_1629 ( P1_U4325 , P1_R1240_U97 , P1_U3967 );
not NOT1_1630 ( P1_U4326 , P1_U3384 );
nand NAND2_1631 ( P1_U4327 , P1_R1222_U97 , P1_U3026 );
nand NAND2_1632 ( P1_U4328 , P1_U3025 , P1_U3062 );
nand NAND2_1633 ( P1_U4329 , P1_R1282_U63 , P1_U3023 );
nand NAND2_1634 ( P1_U4330 , P1_U3479 , P1_U4142 );
nand NAND2_1635 ( P1_U4331 , P1_U3666 , P1_U4326 );
nand NAND2_1636 ( P1_U4332 , P1_REG2_REG_11_ , P1_U3018 );
nand NAND2_1637 ( P1_U4333 , P1_REG1_REG_11_ , P1_U3019 );
nand NAND2_1638 ( P1_U4334 , P1_REG0_REG_11_ , P1_U3020 );
nand NAND2_1639 ( P1_U4335 , P1_ADD_95_U77 , P1_U3017 );
not NOT1_1640 ( P1_U4336 , P1_U3063 );
nand NAND2_1641 ( P1_U4337 , P1_U3033 , P1_U3083 );
nand NAND2_1642 ( P1_U4338 , P1_R1150_U112 , P1_U3961 );
nand NAND2_1643 ( P1_U4339 , P1_R1117_U112 , P1_U3963 );
nand NAND2_1644 ( P1_U4340 , P1_R1138_U11 , P1_U3962 );
nand NAND2_1645 ( P1_U4341 , P1_R1192_U112 , P1_U3959 );
nand NAND2_1646 ( P1_U4342 , P1_R1207_U112 , P1_U3958 );
nand NAND2_1647 ( P1_U4343 , P1_R1171_U11 , P1_U3968 );
nand NAND2_1648 ( P1_U4344 , P1_R1240_U11 , P1_U3967 );
not NOT1_1649 ( P1_U4345 , P1_U3385 );
nand NAND2_1650 ( P1_U4346 , P1_R1222_U11 , P1_U3026 );
nand NAND2_1651 ( P1_U4347 , P1_U3025 , P1_U3063 );
nand NAND2_1652 ( P1_U4348 , P1_R1282_U6 , P1_U3023 );
nand NAND2_1653 ( P1_U4349 , P1_U3482 , P1_U4142 );
nand NAND2_1654 ( P1_U4350 , P1_U3670 , P1_U4345 );
nand NAND2_1655 ( P1_U4351 , P1_REG2_REG_12_ , P1_U3018 );
nand NAND2_1656 ( P1_U4352 , P1_REG1_REG_12_ , P1_U3019 );
nand NAND2_1657 ( P1_U4353 , P1_REG0_REG_12_ , P1_U3020 );
nand NAND2_1658 ( P1_U4354 , P1_ADD_95_U76 , P1_U3017 );
not NOT1_1659 ( P1_U4355 , P1_U3072 );
nand NAND2_1660 ( P1_U4356 , P1_U3033 , P1_U3062 );
nand NAND2_1661 ( P1_U4357 , P1_R1150_U10 , P1_U3961 );
nand NAND2_1662 ( P1_U4358 , P1_R1117_U10 , P1_U3963 );
nand NAND2_1663 ( P1_U4359 , P1_R1138_U115 , P1_U3962 );
nand NAND2_1664 ( P1_U4360 , P1_R1192_U10 , P1_U3959 );
nand NAND2_1665 ( P1_U4361 , P1_R1207_U10 , P1_U3958 );
nand NAND2_1666 ( P1_U4362 , P1_R1171_U115 , P1_U3968 );
nand NAND2_1667 ( P1_U4363 , P1_R1240_U115 , P1_U3967 );
not NOT1_1668 ( P1_U4364 , P1_U3386 );
nand NAND2_1669 ( P1_U4365 , P1_R1222_U115 , P1_U3026 );
nand NAND2_1670 ( P1_U4366 , P1_U3025 , P1_U3072 );
nand NAND2_1671 ( P1_U4367 , P1_R1282_U7 , P1_U3023 );
nand NAND2_1672 ( P1_U4368 , P1_U3485 , P1_U4142 );
nand NAND2_1673 ( P1_U4369 , P1_U3674 , P1_U4364 );
nand NAND2_1674 ( P1_U4370 , P1_REG2_REG_13_ , P1_U3018 );
nand NAND2_1675 ( P1_U4371 , P1_REG1_REG_13_ , P1_U3019 );
nand NAND2_1676 ( P1_U4372 , P1_REG0_REG_13_ , P1_U3020 );
nand NAND2_1677 ( P1_U4373 , P1_ADD_95_U75 , P1_U3017 );
not NOT1_1678 ( P1_U4374 , P1_U3080 );
nand NAND2_1679 ( P1_U4375 , P1_U3033 , P1_U3063 );
nand NAND2_1680 ( P1_U4376 , P1_R1150_U101 , P1_U3961 );
nand NAND2_1681 ( P1_U4377 , P1_R1117_U101 , P1_U3963 );
nand NAND2_1682 ( P1_U4378 , P1_R1138_U114 , P1_U3962 );
nand NAND2_1683 ( P1_U4379 , P1_R1192_U101 , P1_U3959 );
nand NAND2_1684 ( P1_U4380 , P1_R1207_U101 , P1_U3958 );
nand NAND2_1685 ( P1_U4381 , P1_R1171_U114 , P1_U3968 );
nand NAND2_1686 ( P1_U4382 , P1_R1240_U114 , P1_U3967 );
not NOT1_1687 ( P1_U4383 , P1_U3387 );
nand NAND2_1688 ( P1_U4384 , P1_R1222_U114 , P1_U3026 );
nand NAND2_1689 ( P1_U4385 , P1_U3025 , P1_U3080 );
nand NAND2_1690 ( P1_U4386 , P1_R1282_U8 , P1_U3023 );
nand NAND2_1691 ( P1_U4387 , P1_U3488 , P1_U4142 );
nand NAND2_1692 ( P1_U4388 , P1_U3678 , P1_U4383 );
nand NAND2_1693 ( P1_U4389 , P1_REG2_REG_14_ , P1_U3018 );
nand NAND2_1694 ( P1_U4390 , P1_REG1_REG_14_ , P1_U3019 );
nand NAND2_1695 ( P1_U4391 , P1_REG0_REG_14_ , P1_U3020 );
nand NAND2_1696 ( P1_U4392 , P1_ADD_95_U74 , P1_U3017 );
not NOT1_1697 ( P1_U4393 , P1_U3079 );
nand NAND2_1698 ( P1_U4394 , P1_U3033 , P1_U3072 );
nand NAND2_1699 ( P1_U4395 , P1_R1150_U100 , P1_U3961 );
nand NAND2_1700 ( P1_U4396 , P1_R1117_U100 , P1_U3963 );
nand NAND2_1701 ( P1_U4397 , P1_R1138_U12 , P1_U3962 );
nand NAND2_1702 ( P1_U4398 , P1_R1192_U100 , P1_U3959 );
nand NAND2_1703 ( P1_U4399 , P1_R1207_U100 , P1_U3958 );
nand NAND2_1704 ( P1_U4400 , P1_R1171_U12 , P1_U3968 );
nand NAND2_1705 ( P1_U4401 , P1_R1240_U12 , P1_U3967 );
not NOT1_1706 ( P1_U4402 , P1_U3388 );
nand NAND2_1707 ( P1_U4403 , P1_R1222_U12 , P1_U3026 );
nand NAND2_1708 ( P1_U4404 , P1_U3025 , P1_U3079 );
nand NAND2_1709 ( P1_U4405 , P1_R1282_U86 , P1_U3023 );
nand NAND2_1710 ( P1_U4406 , P1_U3491 , P1_U4142 );
nand NAND2_1711 ( P1_U4407 , P1_U3682 , P1_U4402 );
nand NAND2_1712 ( P1_U4408 , P1_REG2_REG_15_ , P1_U3018 );
nand NAND2_1713 ( P1_U4409 , P1_REG1_REG_15_ , P1_U3019 );
nand NAND2_1714 ( P1_U4410 , P1_REG0_REG_15_ , P1_U3020 );
nand NAND2_1715 ( P1_U4411 , P1_ADD_95_U73 , P1_U3017 );
not NOT1_1716 ( P1_U4412 , P1_U3074 );
nand NAND2_1717 ( P1_U4413 , P1_U3033 , P1_U3080 );
nand NAND2_1718 ( P1_U4414 , P1_R1150_U111 , P1_U3961 );
nand NAND2_1719 ( P1_U4415 , P1_R1117_U111 , P1_U3963 );
nand NAND2_1720 ( P1_U4416 , P1_R1138_U113 , P1_U3962 );
nand NAND2_1721 ( P1_U4417 , P1_R1192_U111 , P1_U3959 );
nand NAND2_1722 ( P1_U4418 , P1_R1207_U111 , P1_U3958 );
nand NAND2_1723 ( P1_U4419 , P1_R1171_U113 , P1_U3968 );
nand NAND2_1724 ( P1_U4420 , P1_R1240_U113 , P1_U3967 );
not NOT1_1725 ( P1_U4421 , P1_U3389 );
nand NAND2_1726 ( P1_U4422 , P1_R1222_U113 , P1_U3026 );
nand NAND2_1727 ( P1_U4423 , P1_U3025 , P1_U3074 );
nand NAND2_1728 ( P1_U4424 , P1_R1282_U9 , P1_U3023 );
nand NAND2_1729 ( P1_U4425 , P1_U3494 , P1_U4142 );
nand NAND2_1730 ( P1_U4426 , P1_U3686 , P1_U4421 );
nand NAND2_1731 ( P1_U4427 , P1_REG2_REG_16_ , P1_U3018 );
nand NAND2_1732 ( P1_U4428 , P1_REG1_REG_16_ , P1_U3019 );
nand NAND2_1733 ( P1_U4429 , P1_REG0_REG_16_ , P1_U3020 );
nand NAND2_1734 ( P1_U4430 , P1_ADD_95_U72 , P1_U3017 );
not NOT1_1735 ( P1_U4431 , P1_U3073 );
nand NAND2_1736 ( P1_U4432 , P1_U3033 , P1_U3079 );
nand NAND2_1737 ( P1_U4433 , P1_R1150_U110 , P1_U3961 );
nand NAND2_1738 ( P1_U4434 , P1_R1117_U110 , P1_U3963 );
nand NAND2_1739 ( P1_U4435 , P1_R1138_U112 , P1_U3962 );
nand NAND2_1740 ( P1_U4436 , P1_R1192_U110 , P1_U3959 );
nand NAND2_1741 ( P1_U4437 , P1_R1207_U110 , P1_U3958 );
nand NAND2_1742 ( P1_U4438 , P1_R1171_U112 , P1_U3968 );
nand NAND2_1743 ( P1_U4439 , P1_R1240_U112 , P1_U3967 );
not NOT1_1744 ( P1_U4440 , P1_U3390 );
nand NAND2_1745 ( P1_U4441 , P1_R1222_U112 , P1_U3026 );
nand NAND2_1746 ( P1_U4442 , P1_U3025 , P1_U3073 );
nand NAND2_1747 ( P1_U4443 , P1_R1282_U10 , P1_U3023 );
nand NAND2_1748 ( P1_U4444 , P1_U3497 , P1_U4142 );
nand NAND2_1749 ( P1_U4445 , P1_U3690 , P1_U4440 );
nand NAND2_1750 ( P1_U4446 , P1_REG2_REG_17_ , P1_U3018 );
nand NAND2_1751 ( P1_U4447 , P1_REG1_REG_17_ , P1_U3019 );
nand NAND2_1752 ( P1_U4448 , P1_REG0_REG_17_ , P1_U3020 );
nand NAND2_1753 ( P1_U4449 , P1_ADD_95_U71 , P1_U3017 );
not NOT1_1754 ( P1_U4450 , P1_U3069 );
nand NAND2_1755 ( P1_U4451 , P1_U3033 , P1_U3074 );
nand NAND2_1756 ( P1_U4452 , P1_R1150_U11 , P1_U3961 );
nand NAND2_1757 ( P1_U4453 , P1_R1117_U11 , P1_U3963 );
nand NAND2_1758 ( P1_U4454 , P1_R1138_U111 , P1_U3962 );
nand NAND2_1759 ( P1_U4455 , P1_R1192_U11 , P1_U3959 );
nand NAND2_1760 ( P1_U4456 , P1_R1207_U11 , P1_U3958 );
nand NAND2_1761 ( P1_U4457 , P1_R1171_U111 , P1_U3968 );
nand NAND2_1762 ( P1_U4458 , P1_R1240_U111 , P1_U3967 );
not NOT1_1763 ( P1_U4459 , P1_U3391 );
nand NAND2_1764 ( P1_U4460 , P1_R1222_U111 , P1_U3026 );
nand NAND2_1765 ( P1_U4461 , P1_U3025 , P1_U3069 );
nand NAND2_1766 ( P1_U4462 , P1_R1282_U11 , P1_U3023 );
nand NAND2_1767 ( P1_U4463 , P1_U3500 , P1_U4142 );
nand NAND2_1768 ( P1_U4464 , P1_U3694 , P1_U4459 );
nand NAND2_1769 ( P1_U4465 , P1_REG2_REG_18_ , P1_U3018 );
nand NAND2_1770 ( P1_U4466 , P1_REG1_REG_18_ , P1_U3019 );
nand NAND2_1771 ( P1_U4467 , P1_REG0_REG_18_ , P1_U3020 );
nand NAND2_1772 ( P1_U4468 , P1_ADD_95_U70 , P1_U3017 );
not NOT1_1773 ( P1_U4469 , P1_U3082 );
nand NAND2_1774 ( P1_U4470 , P1_U3033 , P1_U3073 );
nand NAND2_1775 ( P1_U4471 , P1_R1150_U99 , P1_U3961 );
nand NAND2_1776 ( P1_U4472 , P1_R1117_U99 , P1_U3963 );
nand NAND2_1777 ( P1_U4473 , P1_R1138_U13 , P1_U3962 );
nand NAND2_1778 ( P1_U4474 , P1_R1192_U99 , P1_U3959 );
nand NAND2_1779 ( P1_U4475 , P1_R1207_U99 , P1_U3958 );
nand NAND2_1780 ( P1_U4476 , P1_R1171_U13 , P1_U3968 );
nand NAND2_1781 ( P1_U4477 , P1_R1240_U13 , P1_U3967 );
not NOT1_1782 ( P1_U4478 , P1_U3392 );
nand NAND2_1783 ( P1_U4479 , P1_R1222_U13 , P1_U3026 );
nand NAND2_1784 ( P1_U4480 , P1_U3025 , P1_U3082 );
nand NAND2_1785 ( P1_U4481 , P1_R1282_U84 , P1_U3023 );
nand NAND2_1786 ( P1_U4482 , P1_U3503 , P1_U4142 );
nand NAND2_1787 ( P1_U4483 , P1_U3698 , P1_U4478 );
nand NAND2_1788 ( P1_U4484 , P1_REG2_REG_19_ , P1_U3018 );
nand NAND2_1789 ( P1_U4485 , P1_REG1_REG_19_ , P1_U3019 );
nand NAND2_1790 ( P1_U4486 , P1_REG0_REG_19_ , P1_U3020 );
nand NAND2_1791 ( P1_U4487 , P1_ADD_95_U69 , P1_U3017 );
not NOT1_1792 ( P1_U4488 , P1_U3081 );
nand NAND2_1793 ( P1_U4489 , P1_U3033 , P1_U3069 );
nand NAND2_1794 ( P1_U4490 , P1_R1150_U98 , P1_U3961 );
nand NAND2_1795 ( P1_U4491 , P1_R1117_U98 , P1_U3963 );
nand NAND2_1796 ( P1_U4492 , P1_R1138_U110 , P1_U3962 );
nand NAND2_1797 ( P1_U4493 , P1_R1192_U98 , P1_U3959 );
nand NAND2_1798 ( P1_U4494 , P1_R1207_U98 , P1_U3958 );
nand NAND2_1799 ( P1_U4495 , P1_R1171_U110 , P1_U3968 );
nand NAND2_1800 ( P1_U4496 , P1_R1240_U110 , P1_U3967 );
not NOT1_1801 ( P1_U4497 , P1_U3393 );
nand NAND2_1802 ( P1_U4498 , P1_R1222_U110 , P1_U3026 );
nand NAND2_1803 ( P1_U4499 , P1_U3025 , P1_U3081 );
nand NAND2_1804 ( P1_U4500 , P1_R1282_U12 , P1_U3023 );
nand NAND2_1805 ( P1_U4501 , P1_U3506 , P1_U4142 );
nand NAND2_1806 ( P1_U4502 , P1_U3702 , P1_U4497 );
nand NAND2_1807 ( P1_U4503 , P1_REG2_REG_20_ , P1_U3018 );
nand NAND2_1808 ( P1_U4504 , P1_REG1_REG_20_ , P1_U3019 );
nand NAND2_1809 ( P1_U4505 , P1_REG0_REG_20_ , P1_U3020 );
nand NAND2_1810 ( P1_U4506 , P1_ADD_95_U68 , P1_U3017 );
not NOT1_1811 ( P1_U4507 , P1_U3076 );
nand NAND2_1812 ( P1_U4508 , P1_U3033 , P1_U3082 );
nand NAND2_1813 ( P1_U4509 , P1_R1150_U97 , P1_U3961 );
nand NAND2_1814 ( P1_U4510 , P1_R1117_U97 , P1_U3963 );
nand NAND2_1815 ( P1_U4511 , P1_R1138_U109 , P1_U3962 );
nand NAND2_1816 ( P1_U4512 , P1_R1192_U97 , P1_U3959 );
nand NAND2_1817 ( P1_U4513 , P1_R1207_U97 , P1_U3958 );
nand NAND2_1818 ( P1_U4514 , P1_R1171_U109 , P1_U3968 );
nand NAND2_1819 ( P1_U4515 , P1_R1240_U109 , P1_U3967 );
not NOT1_1820 ( P1_U4516 , P1_U3394 );
nand NAND2_1821 ( P1_U4517 , P1_R1222_U109 , P1_U3026 );
nand NAND2_1822 ( P1_U4518 , P1_U3025 , P1_U3076 );
nand NAND2_1823 ( P1_U4519 , P1_R1282_U82 , P1_U3023 );
nand NAND2_1824 ( P1_U4520 , P1_U3508 , P1_U4142 );
nand NAND2_1825 ( P1_U4521 , P1_U3706 , P1_U4516 );
nand NAND2_1826 ( P1_U4522 , P1_REG2_REG_21_ , P1_U3018 );
nand NAND2_1827 ( P1_U4523 , P1_REG1_REG_21_ , P1_U3019 );
nand NAND2_1828 ( P1_U4524 , P1_REG0_REG_21_ , P1_U3020 );
nand NAND2_1829 ( P1_U4525 , P1_ADD_95_U67 , P1_U3017 );
not NOT1_1830 ( P1_U4526 , P1_U3075 );
nand NAND2_1831 ( P1_U4527 , P1_U3033 , P1_U3081 );
nand NAND2_1832 ( P1_U4528 , P1_R1150_U95 , P1_U3961 );
nand NAND2_1833 ( P1_U4529 , P1_R1117_U95 , P1_U3963 );
nand NAND2_1834 ( P1_U4530 , P1_R1138_U14 , P1_U3962 );
nand NAND2_1835 ( P1_U4531 , P1_R1192_U95 , P1_U3959 );
nand NAND2_1836 ( P1_U4532 , P1_R1207_U95 , P1_U3958 );
nand NAND2_1837 ( P1_U4533 , P1_R1171_U14 , P1_U3968 );
nand NAND2_1838 ( P1_U4534 , P1_R1240_U14 , P1_U3967 );
not NOT1_1839 ( P1_U4535 , P1_U3396 );
nand NAND2_1840 ( P1_U4536 , P1_R1222_U14 , P1_U3026 );
nand NAND2_1841 ( P1_U4537 , P1_U3025 , P1_U3075 );
nand NAND2_1842 ( P1_U4538 , P1_R1282_U13 , P1_U3023 );
nand NAND2_1843 ( P1_U4539 , P1_U3982 , P1_U4142 );
nand NAND2_1844 ( P1_U4540 , P1_U3710 , P1_U4535 );
nand NAND2_1845 ( P1_U4541 , P1_REG2_REG_22_ , P1_U3018 );
nand NAND2_1846 ( P1_U4542 , P1_REG1_REG_22_ , P1_U3019 );
nand NAND2_1847 ( P1_U4543 , P1_REG0_REG_22_ , P1_U3020 );
nand NAND2_1848 ( P1_U4544 , P1_ADD_95_U66 , P1_U3017 );
not NOT1_1849 ( P1_U4545 , P1_U3061 );
nand NAND2_1850 ( P1_U4546 , P1_U3033 , P1_U3076 );
nand NAND2_1851 ( P1_U4547 , P1_R1150_U109 , P1_U3961 );
nand NAND2_1852 ( P1_U4548 , P1_R1117_U109 , P1_U3963 );
nand NAND2_1853 ( P1_U4549 , P1_R1138_U15 , P1_U3962 );
nand NAND2_1854 ( P1_U4550 , P1_R1192_U109 , P1_U3959 );
nand NAND2_1855 ( P1_U4551 , P1_R1207_U109 , P1_U3958 );
nand NAND2_1856 ( P1_U4552 , P1_R1171_U15 , P1_U3968 );
nand NAND2_1857 ( P1_U4553 , P1_R1240_U15 , P1_U3967 );
not NOT1_1858 ( P1_U4554 , P1_U3398 );
nand NAND2_1859 ( P1_U4555 , P1_R1222_U15 , P1_U3026 );
nand NAND2_1860 ( P1_U4556 , P1_U3025 , P1_U3061 );
nand NAND2_1861 ( P1_U4557 , P1_R1282_U78 , P1_U3023 );
nand NAND2_1862 ( P1_U4558 , P1_U3981 , P1_U4142 );
nand NAND2_1863 ( P1_U4559 , P1_U3714 , P1_U4554 );
nand NAND2_1864 ( P1_U4560 , P1_REG2_REG_23_ , P1_U3018 );
nand NAND2_1865 ( P1_U4561 , P1_REG1_REG_23_ , P1_U3019 );
nand NAND2_1866 ( P1_U4562 , P1_REG0_REG_23_ , P1_U3020 );
nand NAND2_1867 ( P1_U4563 , P1_ADD_95_U65 , P1_U3017 );
not NOT1_1868 ( P1_U4564 , P1_U3066 );
nand NAND2_1869 ( P1_U4565 , P1_U3033 , P1_U3075 );
nand NAND2_1870 ( P1_U4566 , P1_R1150_U108 , P1_U3961 );
nand NAND2_1871 ( P1_U4567 , P1_R1117_U108 , P1_U3963 );
nand NAND2_1872 ( P1_U4568 , P1_R1138_U108 , P1_U3962 );
nand NAND2_1873 ( P1_U4569 , P1_R1192_U108 , P1_U3959 );
nand NAND2_1874 ( P1_U4570 , P1_R1207_U108 , P1_U3958 );
nand NAND2_1875 ( P1_U4571 , P1_R1171_U108 , P1_U3968 );
nand NAND2_1876 ( P1_U4572 , P1_R1240_U108 , P1_U3967 );
not NOT1_1877 ( P1_U4573 , P1_U3400 );
nand NAND2_1878 ( P1_U4574 , P1_R1222_U108 , P1_U3026 );
nand NAND2_1879 ( P1_U4575 , P1_U3025 , P1_U3066 );
nand NAND2_1880 ( P1_U4576 , P1_R1282_U14 , P1_U3023 );
nand NAND2_1881 ( P1_U4577 , P1_U3980 , P1_U4142 );
nand NAND2_1882 ( P1_U4578 , P1_U3718 , P1_U4573 );
nand NAND2_1883 ( P1_U4579 , P1_REG2_REG_24_ , P1_U3018 );
nand NAND2_1884 ( P1_U4580 , P1_REG1_REG_24_ , P1_U3019 );
nand NAND2_1885 ( P1_U4581 , P1_REG0_REG_24_ , P1_U3020 );
nand NAND2_1886 ( P1_U4582 , P1_ADD_95_U64 , P1_U3017 );
not NOT1_1887 ( P1_U4583 , P1_U3065 );
nand NAND2_1888 ( P1_U4584 , P1_U3033 , P1_U3061 );
nand NAND2_1889 ( P1_U4585 , P1_R1150_U12 , P1_U3961 );
nand NAND2_1890 ( P1_U4586 , P1_R1117_U12 , P1_U3963 );
nand NAND2_1891 ( P1_U4587 , P1_R1138_U107 , P1_U3962 );
nand NAND2_1892 ( P1_U4588 , P1_R1192_U12 , P1_U3959 );
nand NAND2_1893 ( P1_U4589 , P1_R1207_U12 , P1_U3958 );
nand NAND2_1894 ( P1_U4590 , P1_R1171_U107 , P1_U3968 );
nand NAND2_1895 ( P1_U4591 , P1_R1240_U107 , P1_U3967 );
not NOT1_1896 ( P1_U4592 , P1_U3402 );
nand NAND2_1897 ( P1_U4593 , P1_R1222_U107 , P1_U3026 );
nand NAND2_1898 ( P1_U4594 , P1_U3025 , P1_U3065 );
nand NAND2_1899 ( P1_U4595 , P1_R1282_U76 , P1_U3023 );
nand NAND2_1900 ( P1_U4596 , P1_U3979 , P1_U4142 );
nand NAND2_1901 ( P1_U4597 , P1_U3722 , P1_U4592 );
nand NAND2_1902 ( P1_U4598 , P1_REG2_REG_25_ , P1_U3018 );
nand NAND2_1903 ( P1_U4599 , P1_REG1_REG_25_ , P1_U3019 );
nand NAND2_1904 ( P1_U4600 , P1_REG0_REG_25_ , P1_U3020 );
nand NAND2_1905 ( P1_U4601 , P1_ADD_95_U63 , P1_U3017 );
not NOT1_1906 ( P1_U4602 , P1_U3058 );
nand NAND2_1907 ( P1_U4603 , P1_U3033 , P1_U3066 );
nand NAND2_1908 ( P1_U4604 , P1_R1150_U94 , P1_U3961 );
nand NAND2_1909 ( P1_U4605 , P1_R1117_U94 , P1_U3963 );
nand NAND2_1910 ( P1_U4606 , P1_R1138_U106 , P1_U3962 );
nand NAND2_1911 ( P1_U4607 , P1_R1192_U94 , P1_U3959 );
nand NAND2_1912 ( P1_U4608 , P1_R1207_U94 , P1_U3958 );
nand NAND2_1913 ( P1_U4609 , P1_R1171_U106 , P1_U3968 );
nand NAND2_1914 ( P1_U4610 , P1_R1240_U106 , P1_U3967 );
not NOT1_1915 ( P1_U4611 , P1_U3404 );
nand NAND2_1916 ( P1_U4612 , P1_R1222_U106 , P1_U3026 );
nand NAND2_1917 ( P1_U4613 , P1_U3025 , P1_U3058 );
nand NAND2_1918 ( P1_U4614 , P1_R1282_U15 , P1_U3023 );
nand NAND2_1919 ( P1_U4615 , P1_U3978 , P1_U4142 );
nand NAND2_1920 ( P1_U4616 , P1_U3726 , P1_U4611 );
nand NAND2_1921 ( P1_U4617 , P1_REG2_REG_26_ , P1_U3018 );
nand NAND2_1922 ( P1_U4618 , P1_REG1_REG_26_ , P1_U3019 );
nand NAND2_1923 ( P1_U4619 , P1_REG0_REG_26_ , P1_U3020 );
nand NAND2_1924 ( P1_U4620 , P1_ADD_95_U62 , P1_U3017 );
not NOT1_1925 ( P1_U4621 , P1_U3057 );
nand NAND2_1926 ( P1_U4622 , P1_U3033 , P1_U3065 );
nand NAND2_1927 ( P1_U4623 , P1_R1150_U93 , P1_U3961 );
nand NAND2_1928 ( P1_U4624 , P1_R1117_U93 , P1_U3963 );
nand NAND2_1929 ( P1_U4625 , P1_R1138_U105 , P1_U3962 );
nand NAND2_1930 ( P1_U4626 , P1_R1192_U93 , P1_U3959 );
nand NAND2_1931 ( P1_U4627 , P1_R1207_U93 , P1_U3958 );
nand NAND2_1932 ( P1_U4628 , P1_R1171_U105 , P1_U3968 );
nand NAND2_1933 ( P1_U4629 , P1_R1240_U105 , P1_U3967 );
not NOT1_1934 ( P1_U4630 , P1_U3406 );
nand NAND2_1935 ( P1_U4631 , P1_R1222_U105 , P1_U3026 );
nand NAND2_1936 ( P1_U4632 , P1_U3025 , P1_U3057 );
nand NAND2_1937 ( P1_U4633 , P1_R1282_U74 , P1_U3023 );
nand NAND2_1938 ( P1_U4634 , P1_U3977 , P1_U4142 );
nand NAND2_1939 ( P1_U4635 , P1_U3730 , P1_U4630 );
nand NAND2_1940 ( P1_U4636 , P1_REG2_REG_27_ , P1_U3018 );
nand NAND2_1941 ( P1_U4637 , P1_REG1_REG_27_ , P1_U3019 );
nand NAND2_1942 ( P1_U4638 , P1_REG0_REG_27_ , P1_U3020 );
nand NAND2_1943 ( P1_U4639 , P1_ADD_95_U61 , P1_U3017 );
not NOT1_1944 ( P1_U4640 , P1_U3053 );
nand NAND2_1945 ( P1_U4641 , P1_U3033 , P1_U3058 );
nand NAND2_1946 ( P1_U4642 , P1_R1150_U107 , P1_U3961 );
nand NAND2_1947 ( P1_U4643 , P1_R1117_U107 , P1_U3963 );
nand NAND2_1948 ( P1_U4644 , P1_R1138_U16 , P1_U3962 );
nand NAND2_1949 ( P1_U4645 , P1_R1192_U107 , P1_U3959 );
nand NAND2_1950 ( P1_U4646 , P1_R1207_U107 , P1_U3958 );
nand NAND2_1951 ( P1_U4647 , P1_R1171_U16 , P1_U3968 );
nand NAND2_1952 ( P1_U4648 , P1_R1240_U16 , P1_U3967 );
not NOT1_1953 ( P1_U4649 , P1_U3408 );
nand NAND2_1954 ( P1_U4650 , P1_R1222_U16 , P1_U3026 );
nand NAND2_1955 ( P1_U4651 , P1_U3025 , P1_U3053 );
nand NAND2_1956 ( P1_U4652 , P1_R1282_U16 , P1_U3023 );
nand NAND2_1957 ( P1_U4653 , P1_U3976 , P1_U4142 );
nand NAND2_1958 ( P1_U4654 , P1_U3734 , P1_U4649 );
nand NAND2_1959 ( P1_U4655 , P1_REG2_REG_28_ , P1_U3018 );
nand NAND2_1960 ( P1_U4656 , P1_REG1_REG_28_ , P1_U3019 );
nand NAND2_1961 ( P1_U4657 , P1_REG0_REG_28_ , P1_U3020 );
nand NAND2_1962 ( P1_U4658 , P1_ADD_95_U60 , P1_U3017 );
not NOT1_1963 ( P1_U4659 , P1_U3054 );
nand NAND2_1964 ( P1_U4660 , P1_U3033 , P1_U3057 );
nand NAND2_1965 ( P1_U4661 , P1_R1150_U13 , P1_U3961 );
nand NAND2_1966 ( P1_U4662 , P1_R1117_U13 , P1_U3963 );
nand NAND2_1967 ( P1_U4663 , P1_R1138_U104 , P1_U3962 );
nand NAND2_1968 ( P1_U4664 , P1_R1192_U13 , P1_U3959 );
nand NAND2_1969 ( P1_U4665 , P1_R1207_U13 , P1_U3958 );
nand NAND2_1970 ( P1_U4666 , P1_R1171_U104 , P1_U3968 );
nand NAND2_1971 ( P1_U4667 , P1_R1240_U104 , P1_U3967 );
not NOT1_1972 ( P1_U4668 , P1_U3410 );
nand NAND2_1973 ( P1_U4669 , P1_R1222_U104 , P1_U3026 );
nand NAND2_1974 ( P1_U4670 , P1_U3025 , P1_U3054 );
nand NAND2_1975 ( P1_U4671 , P1_R1282_U72 , P1_U3023 );
nand NAND2_1976 ( P1_U4672 , P1_U3975 , P1_U4142 );
nand NAND2_1977 ( P1_U4673 , P1_U3738 , P1_U4668 );
nand NAND2_1978 ( P1_U4674 , P1_ADD_95_U5 , P1_U3017 );
nand NAND2_1979 ( P1_U4675 , P1_REG2_REG_29_ , P1_U3018 );
nand NAND2_1980 ( P1_U4676 , P1_REG1_REG_29_ , P1_U3019 );
nand NAND2_1981 ( P1_U4677 , P1_REG0_REG_29_ , P1_U3020 );
not NOT1_1982 ( P1_U4678 , P1_U3055 );
nand NAND2_1983 ( P1_U4679 , P1_U3033 , P1_U3053 );
nand NAND2_1984 ( P1_U4680 , P1_R1150_U92 , P1_U3961 );
nand NAND2_1985 ( P1_U4681 , P1_R1117_U92 , P1_U3963 );
nand NAND2_1986 ( P1_U4682 , P1_R1138_U103 , P1_U3962 );
nand NAND2_1987 ( P1_U4683 , P1_R1192_U92 , P1_U3959 );
nand NAND2_1988 ( P1_U4684 , P1_R1207_U92 , P1_U3958 );
nand NAND2_1989 ( P1_U4685 , P1_R1171_U103 , P1_U3968 );
nand NAND2_1990 ( P1_U4686 , P1_R1240_U103 , P1_U3967 );
not NOT1_1991 ( P1_U4687 , P1_U3412 );
nand NAND2_1992 ( P1_U4688 , P1_R1222_U103 , P1_U3026 );
nand NAND2_1993 ( P1_U4689 , P1_U3025 , P1_U3055 );
nand NAND2_1994 ( P1_U4690 , P1_R1282_U17 , P1_U3023 );
nand NAND2_1995 ( P1_U4691 , P1_U3974 , P1_U4142 );
nand NAND2_1996 ( P1_U4692 , P1_U3742 , P1_U4687 );
nand NAND2_1997 ( P1_U4693 , P1_REG2_REG_30_ , P1_U3018 );
nand NAND2_1998 ( P1_U4694 , P1_REG1_REG_30_ , P1_U3019 );
nand NAND2_1999 ( P1_U4695 , P1_REG0_REG_30_ , P1_U3020 );
not NOT1_2000 ( P1_U4696 , P1_U3059 );
nand NAND2_2001 ( P1_U4697 , P1_U5699 , P1_U3359 );
nand NAND2_2002 ( P1_U4698 , P1_U3912 , P1_U4697 );
nand NAND2_2003 ( P1_U4699 , P1_U3743 , P1_U3059 );
nand NAND2_2004 ( P1_U4700 , P1_U3033 , P1_U3054 );
nand NAND2_2005 ( P1_U4701 , P1_R1150_U14 , P1_U3961 );
nand NAND2_2006 ( P1_U4702 , P1_R1117_U14 , P1_U3963 );
nand NAND2_2007 ( P1_U4703 , P1_R1138_U102 , P1_U3962 );
nand NAND2_2008 ( P1_U4704 , P1_R1192_U14 , P1_U3959 );
nand NAND2_2009 ( P1_U4705 , P1_R1207_U14 , P1_U3958 );
nand NAND2_2010 ( P1_U4706 , P1_R1171_U102 , P1_U3968 );
nand NAND2_2011 ( P1_U4707 , P1_R1240_U102 , P1_U3967 );
nand NAND3_2012 ( P1_U4708 , P1_U3802 , P1_U3051 , P1_U3801 );
nand NAND2_2013 ( P1_U4709 , P1_R1222_U102 , P1_U3026 );
nand NAND2_2014 ( P1_U4710 , P1_R1282_U70 , P1_U3023 );
nand NAND2_2015 ( P1_U4711 , P1_U3985 , P1_U4142 );
nand NAND4_2016 ( P1_U4712 , P1_U3746 , P1_U3051 , P1_U3745 , P1_U3744 );
nand NAND2_2017 ( P1_U4713 , P1_REG2_REG_31_ , P1_U3018 );
nand NAND2_2018 ( P1_U4714 , P1_REG1_REG_31_ , P1_U3019 );
nand NAND2_2019 ( P1_U4715 , P1_REG0_REG_31_ , P1_U3020 );
not NOT1_2020 ( P1_U4716 , P1_U3056 );
nand NAND2_2021 ( P1_U4717 , P1_R1282_U19 , P1_U3023 );
nand NAND2_2022 ( P1_U4718 , P1_U3984 , P1_U4142 );
nand NAND3_2023 ( P1_U4719 , P1_U4718 , P1_U3945 , P1_U4717 );
nand NAND2_2024 ( P1_U4720 , P1_R1282_U68 , P1_U3023 );
nand NAND2_2025 ( P1_U4721 , P1_U3983 , P1_U4142 );
nand NAND3_2026 ( P1_U4722 , P1_U4721 , P1_U3945 , P1_U4720 );
nand NAND2_2027 ( P1_U4723 , P1_U3749 , P1_U3016 );
nand NAND2_2028 ( P1_U4724 , P1_U3418 , P1_U4723 );
nand NAND2_2029 ( P1_U4725 , P1_U3988 , P1_U3441 );
not NOT1_2030 ( P1_U4726 , P1_U3422 );
nand NAND2_2031 ( P1_U4727 , P1_U3035 , P1_U3078 );
nand NAND2_2032 ( P1_U4728 , P1_U3032 , P1_REG3_REG_0_ );
nand NAND2_2033 ( P1_U4729 , P1_U3031 , P1_R1222_U96 );
nand NAND2_2034 ( P1_U4730 , P1_U3030 , P1_U3450 );
nand NAND2_2035 ( P1_U4731 , P1_U3029 , P1_U3450 );
nand NAND2_2036 ( P1_U4732 , P1_U3035 , P1_U3068 );
nand NAND2_2037 ( P1_U4733 , P1_U3032 , P1_REG3_REG_1_ );
nand NAND2_2038 ( P1_U4734 , P1_U3031 , P1_R1222_U95 );
nand NAND2_2039 ( P1_U4735 , P1_U3030 , P1_U3455 );
nand NAND2_2040 ( P1_U4736 , P1_U3029 , P1_R1282_U57 );
nand NAND2_2041 ( P1_U4737 , P1_U3035 , P1_U3064 );
nand NAND2_2042 ( P1_U4738 , P1_U3032 , P1_REG3_REG_2_ );
nand NAND2_2043 ( P1_U4739 , P1_U3031 , P1_R1222_U17 );
nand NAND2_2044 ( P1_U4740 , P1_U3030 , P1_U3458 );
nand NAND2_2045 ( P1_U4741 , P1_U3029 , P1_R1282_U18 );
nand NAND2_2046 ( P1_U4742 , P1_U3035 , P1_U3060 );
nand NAND2_2047 ( P1_U4743 , P1_U3032 , P1_ADD_95_U4 );
nand NAND2_2048 ( P1_U4744 , P1_U3031 , P1_R1222_U101 );
nand NAND2_2049 ( P1_U4745 , P1_U3030 , P1_U3461 );
nand NAND2_2050 ( P1_U4746 , P1_U3029 , P1_R1282_U20 );
nand NAND2_2051 ( P1_U4747 , P1_U3035 , P1_U3067 );
nand NAND2_2052 ( P1_U4748 , P1_U3032 , P1_ADD_95_U59 );
nand NAND2_2053 ( P1_U4749 , P1_U3031 , P1_R1222_U100 );
nand NAND2_2054 ( P1_U4750 , P1_U3030 , P1_U3464 );
nand NAND2_2055 ( P1_U4751 , P1_U3029 , P1_R1282_U21 );
nand NAND2_2056 ( P1_U4752 , P1_U3035 , P1_U3071 );
nand NAND2_2057 ( P1_U4753 , P1_U3032 , P1_ADD_95_U58 );
nand NAND2_2058 ( P1_U4754 , P1_U3031 , P1_R1222_U18 );
nand NAND2_2059 ( P1_U4755 , P1_U3030 , P1_U3467 );
nand NAND2_2060 ( P1_U4756 , P1_U3029 , P1_R1282_U65 );
nand NAND2_2061 ( P1_U4757 , P1_U3035 , P1_U3070 );
nand NAND2_2062 ( P1_U4758 , P1_U3032 , P1_ADD_95_U57 );
nand NAND2_2063 ( P1_U4759 , P1_U3031 , P1_R1222_U99 );
nand NAND2_2064 ( P1_U4760 , P1_U3030 , P1_U3470 );
nand NAND2_2065 ( P1_U4761 , P1_U3029 , P1_R1282_U22 );
nand NAND2_2066 ( P1_U4762 , P1_U3035 , P1_U3084 );
nand NAND2_2067 ( P1_U4763 , P1_U3032 , P1_ADD_95_U56 );
nand NAND2_2068 ( P1_U4764 , P1_U3031 , P1_R1222_U19 );
nand NAND2_2069 ( P1_U4765 , P1_U3030 , P1_U3473 );
nand NAND2_2070 ( P1_U4766 , P1_U3029 , P1_R1282_U23 );
nand NAND2_2071 ( P1_U4767 , P1_U3035 , P1_U3083 );
nand NAND2_2072 ( P1_U4768 , P1_U3032 , P1_ADD_95_U55 );
nand NAND2_2073 ( P1_U4769 , P1_U3031 , P1_R1222_U98 );
nand NAND2_2074 ( P1_U4770 , P1_U3030 , P1_U3476 );
nand NAND2_2075 ( P1_U4771 , P1_U3029 , P1_R1282_U24 );
nand NAND2_2076 ( P1_U4772 , P1_U3035 , P1_U3062 );
nand NAND2_2077 ( P1_U4773 , P1_U3032 , P1_ADD_95_U54 );
nand NAND2_2078 ( P1_U4774 , P1_U3031 , P1_R1222_U97 );
nand NAND2_2079 ( P1_U4775 , P1_U3030 , P1_U3479 );
nand NAND2_2080 ( P1_U4776 , P1_U3029 , P1_R1282_U63 );
nand NAND2_2081 ( P1_U4777 , P1_U3035 , P1_U3063 );
nand NAND2_2082 ( P1_U4778 , P1_U3032 , P1_ADD_95_U78 );
nand NAND2_2083 ( P1_U4779 , P1_U3031 , P1_R1222_U11 );
nand NAND2_2084 ( P1_U4780 , P1_U3030 , P1_U3482 );
nand NAND2_2085 ( P1_U4781 , P1_U3029 , P1_R1282_U6 );
nand NAND2_2086 ( P1_U4782 , P1_U3035 , P1_U3072 );
nand NAND2_2087 ( P1_U4783 , P1_U3032 , P1_ADD_95_U77 );
nand NAND2_2088 ( P1_U4784 , P1_U3031 , P1_R1222_U115 );
nand NAND2_2089 ( P1_U4785 , P1_U3030 , P1_U3485 );
nand NAND2_2090 ( P1_U4786 , P1_U3029 , P1_R1282_U7 );
nand NAND2_2091 ( P1_U4787 , P1_U3035 , P1_U3080 );
nand NAND2_2092 ( P1_U4788 , P1_U3032 , P1_ADD_95_U76 );
nand NAND2_2093 ( P1_U4789 , P1_U3031 , P1_R1222_U114 );
nand NAND2_2094 ( P1_U4790 , P1_U3030 , P1_U3488 );
nand NAND2_2095 ( P1_U4791 , P1_U3029 , P1_R1282_U8 );
nand NAND2_2096 ( P1_U4792 , P1_U3035 , P1_U3079 );
nand NAND2_2097 ( P1_U4793 , P1_U3032 , P1_ADD_95_U75 );
nand NAND2_2098 ( P1_U4794 , P1_U3031 , P1_R1222_U12 );
nand NAND2_2099 ( P1_U4795 , P1_U3030 , P1_U3491 );
nand NAND2_2100 ( P1_U4796 , P1_U3029 , P1_R1282_U86 );
nand NAND2_2101 ( P1_U4797 , P1_U3035 , P1_U3074 );
nand NAND2_2102 ( P1_U4798 , P1_U3032 , P1_ADD_95_U74 );
nand NAND2_2103 ( P1_U4799 , P1_U3031 , P1_R1222_U113 );
nand NAND2_2104 ( P1_U4800 , P1_U3030 , P1_U3494 );
nand NAND2_2105 ( P1_U4801 , P1_U3029 , P1_R1282_U9 );
nand NAND2_2106 ( P1_U4802 , P1_U3035 , P1_U3073 );
nand NAND2_2107 ( P1_U4803 , P1_U3032 , P1_ADD_95_U73 );
nand NAND2_2108 ( P1_U4804 , P1_U3031 , P1_R1222_U112 );
nand NAND2_2109 ( P1_U4805 , P1_U3030 , P1_U3497 );
nand NAND2_2110 ( P1_U4806 , P1_U3029 , P1_R1282_U10 );
nand NAND2_2111 ( P1_U4807 , P1_U3035 , P1_U3069 );
nand NAND2_2112 ( P1_U4808 , P1_U3032 , P1_ADD_95_U72 );
nand NAND2_2113 ( P1_U4809 , P1_U3031 , P1_R1222_U111 );
nand NAND2_2114 ( P1_U4810 , P1_U3030 , P1_U3500 );
nand NAND2_2115 ( P1_U4811 , P1_U3029 , P1_R1282_U11 );
nand NAND2_2116 ( P1_U4812 , P1_U3035 , P1_U3082 );
nand NAND2_2117 ( P1_U4813 , P1_U3032 , P1_ADD_95_U71 );
nand NAND2_2118 ( P1_U4814 , P1_U3031 , P1_R1222_U13 );
nand NAND2_2119 ( P1_U4815 , P1_U3030 , P1_U3503 );
nand NAND2_2120 ( P1_U4816 , P1_U3029 , P1_R1282_U84 );
nand NAND2_2121 ( P1_U4817 , P1_U3035 , P1_U3081 );
nand NAND2_2122 ( P1_U4818 , P1_U3032 , P1_ADD_95_U70 );
nand NAND2_2123 ( P1_U4819 , P1_U3031 , P1_R1222_U110 );
nand NAND2_2124 ( P1_U4820 , P1_U3030 , P1_U3506 );
nand NAND2_2125 ( P1_U4821 , P1_U3029 , P1_R1282_U12 );
nand NAND2_2126 ( P1_U4822 , P1_U3035 , P1_U3076 );
nand NAND2_2127 ( P1_U4823 , P1_U3032 , P1_ADD_95_U69 );
nand NAND2_2128 ( P1_U4824 , P1_U3031 , P1_R1222_U109 );
nand NAND2_2129 ( P1_U4825 , P1_U3030 , P1_U3508 );
nand NAND2_2130 ( P1_U4826 , P1_U3029 , P1_R1282_U82 );
nand NAND2_2131 ( P1_U4827 , P1_U3035 , P1_U3075 );
nand NAND2_2132 ( P1_U4828 , P1_U3032 , P1_ADD_95_U68 );
nand NAND2_2133 ( P1_U4829 , P1_U3031 , P1_R1222_U14 );
nand NAND2_2134 ( P1_U4830 , P1_U3030 , P1_U3982 );
nand NAND2_2135 ( P1_U4831 , P1_U3029 , P1_R1282_U13 );
nand NAND2_2136 ( P1_U4832 , P1_U3035 , P1_U3061 );
nand NAND2_2137 ( P1_U4833 , P1_U3032 , P1_ADD_95_U67 );
nand NAND2_2138 ( P1_U4834 , P1_U3031 , P1_R1222_U15 );
nand NAND2_2139 ( P1_U4835 , P1_U3030 , P1_U3981 );
nand NAND2_2140 ( P1_U4836 , P1_U3029 , P1_R1282_U78 );
nand NAND2_2141 ( P1_U4837 , P1_U3035 , P1_U3066 );
nand NAND2_2142 ( P1_U4838 , P1_U3032 , P1_ADD_95_U66 );
nand NAND2_2143 ( P1_U4839 , P1_U3031 , P1_R1222_U108 );
nand NAND2_2144 ( P1_U4840 , P1_U3030 , P1_U3980 );
nand NAND2_2145 ( P1_U4841 , P1_U3029 , P1_R1282_U14 );
nand NAND2_2146 ( P1_U4842 , P1_U3035 , P1_U3065 );
nand NAND2_2147 ( P1_U4843 , P1_U3032 , P1_ADD_95_U65 );
nand NAND2_2148 ( P1_U4844 , P1_U3031 , P1_R1222_U107 );
nand NAND2_2149 ( P1_U4845 , P1_U3030 , P1_U3979 );
nand NAND2_2150 ( P1_U4846 , P1_U3029 , P1_R1282_U76 );
nand NAND2_2151 ( P1_U4847 , P1_U3035 , P1_U3058 );
nand NAND2_2152 ( P1_U4848 , P1_U3032 , P1_ADD_95_U64 );
nand NAND2_2153 ( P1_U4849 , P1_U3031 , P1_R1222_U106 );
nand NAND2_2154 ( P1_U4850 , P1_U3030 , P1_U3978 );
nand NAND2_2155 ( P1_U4851 , P1_U3029 , P1_R1282_U15 );
nand NAND2_2156 ( P1_U4852 , P1_U3035 , P1_U3057 );
nand NAND2_2157 ( P1_U4853 , P1_U3032 , P1_ADD_95_U63 );
nand NAND2_2158 ( P1_U4854 , P1_U3031 , P1_R1222_U105 );
nand NAND2_2159 ( P1_U4855 , P1_U3030 , P1_U3977 );
nand NAND2_2160 ( P1_U4856 , P1_U3029 , P1_R1282_U74 );
nand NAND2_2161 ( P1_U4857 , P1_U3035 , P1_U3053 );
nand NAND2_2162 ( P1_U4858 , P1_U3032 , P1_ADD_95_U62 );
nand NAND2_2163 ( P1_U4859 , P1_U3031 , P1_R1222_U16 );
nand NAND2_2164 ( P1_U4860 , P1_U3030 , P1_U3976 );
nand NAND2_2165 ( P1_U4861 , P1_U3029 , P1_R1282_U16 );
nand NAND2_2166 ( P1_U4862 , P1_U3035 , P1_U3054 );
nand NAND2_2167 ( P1_U4863 , P1_U3032 , P1_ADD_95_U61 );
nand NAND2_2168 ( P1_U4864 , P1_U3031 , P1_R1222_U104 );
nand NAND2_2169 ( P1_U4865 , P1_U3030 , P1_U3975 );
nand NAND2_2170 ( P1_U4866 , P1_U3029 , P1_R1282_U72 );
nand NAND2_2171 ( P1_U4867 , P1_U3035 , P1_U3055 );
nand NAND2_2172 ( P1_U4868 , P1_U3032 , P1_ADD_95_U60 );
nand NAND2_2173 ( P1_U4869 , P1_U3031 , P1_R1222_U103 );
nand NAND2_2174 ( P1_U4870 , P1_U3030 , P1_U3974 );
nand NAND2_2175 ( P1_U4871 , P1_U3029 , P1_R1282_U17 );
nand NAND2_2176 ( P1_U4872 , P1_U3032 , P1_ADD_95_U5 );
nand NAND2_2177 ( P1_U4873 , P1_U3031 , P1_R1222_U102 );
nand NAND2_2178 ( P1_U4874 , P1_U3030 , P1_U3985 );
nand NAND2_2179 ( P1_U4875 , P1_U3029 , P1_R1282_U70 );
nand NAND2_2180 ( P1_U4876 , P1_U3030 , P1_U3984 );
nand NAND2_2181 ( P1_U4877 , P1_U3029 , P1_R1282_U19 );
nand NAND2_2182 ( P1_U4878 , P1_U3030 , P1_U3983 );
nand NAND2_2183 ( P1_U4879 , P1_U3029 , P1_R1282_U68 );
nand NAND5_2184 ( P1_U4880 , P1_U3804 , P1_U3803 , P1_U3806 , P1_U4726 , P1_U3418 );
nand NAND2_2185 ( P1_U4881 , P1_R1105_U13 , P1_U3041 );
nand NAND2_2186 ( P1_U4882 , P1_U3039 , P1_U3442 );
nand NAND2_2187 ( P1_U4883 , P1_R1162_U13 , P1_U3037 );
nand NAND3_2188 ( P1_U4884 , P1_U4882 , P1_U4881 , P1_U4883 );
nand NAND2_2189 ( P1_U4885 , P1_U3046 , P1_U3373 );
nand NAND2_2190 ( P1_U4886 , P1_U5677 , P1_U4885 );
nand NAND2_2191 ( P1_U4887 , P1_U4886 , P1_U3912 );
not NOT1_2192 ( P1_U4888 , P1_U3085 );
not NOT1_2193 ( P1_U4889 , P1_U3423 );
nand NAND2_2194 ( P1_U4890 , P1_U3043 , P1_U4884 );
nand NAND2_2195 ( P1_U4891 , P1_U3042 , P1_R1105_U13 );
nand NAND2_2196 ( P1_U4892 , P1_REG3_REG_19_ , P1_U3086 );
nand NAND2_2197 ( P1_U4893 , P1_U3040 , P1_U3442 );
nand NAND2_2198 ( P1_U4894 , P1_U3038 , P1_R1162_U13 );
nand NAND2_2199 ( P1_U4895 , P1_ADDR_REG_19_ , P1_U4889 );
nand NAND2_2200 ( P1_U4896 , P1_R1105_U75 , P1_U3041 );
nand NAND2_2201 ( P1_U4897 , P1_U3039 , P1_U3505 );
nand NAND2_2202 ( P1_U4898 , P1_R1162_U75 , P1_U3037 );
nand NAND3_2203 ( P1_U4899 , P1_U4897 , P1_U4896 , P1_U4898 );
nand NAND2_2204 ( P1_U4900 , P1_U3043 , P1_U4899 );
nand NAND2_2205 ( P1_U4901 , P1_R1105_U75 , P1_U3042 );
nand NAND2_2206 ( P1_U4902 , P1_REG3_REG_18_ , P1_U3086 );
nand NAND2_2207 ( P1_U4903 , P1_U3040 , P1_U3505 );
nand NAND2_2208 ( P1_U4904 , P1_R1162_U75 , P1_U3038 );
nand NAND2_2209 ( P1_U4905 , P1_ADDR_REG_18_ , P1_U4889 );
nand NAND2_2210 ( P1_U4906 , P1_R1105_U12 , P1_U3041 );
nand NAND2_2211 ( P1_U4907 , P1_U3039 , P1_U3502 );
nand NAND2_2212 ( P1_U4908 , P1_R1162_U12 , P1_U3037 );
nand NAND3_2213 ( P1_U4909 , P1_U4907 , P1_U4906 , P1_U4908 );
nand NAND2_2214 ( P1_U4910 , P1_U3043 , P1_U4909 );
nand NAND2_2215 ( P1_U4911 , P1_R1105_U12 , P1_U3042 );
nand NAND2_2216 ( P1_U4912 , P1_REG3_REG_17_ , P1_U3086 );
nand NAND2_2217 ( P1_U4913 , P1_U3040 , P1_U3502 );
nand NAND2_2218 ( P1_U4914 , P1_R1162_U12 , P1_U3038 );
nand NAND2_2219 ( P1_U4915 , P1_ADDR_REG_17_ , P1_U4889 );
nand NAND2_2220 ( P1_U4916 , P1_R1105_U76 , P1_U3041 );
nand NAND2_2221 ( P1_U4917 , P1_U3039 , P1_U3499 );
nand NAND2_2222 ( P1_U4918 , P1_R1162_U76 , P1_U3037 );
nand NAND3_2223 ( P1_U4919 , P1_U4917 , P1_U4916 , P1_U4918 );
nand NAND2_2224 ( P1_U4920 , P1_U3043 , P1_U4919 );
nand NAND2_2225 ( P1_U4921 , P1_R1105_U76 , P1_U3042 );
nand NAND2_2226 ( P1_U4922 , P1_REG3_REG_16_ , P1_U3086 );
nand NAND2_2227 ( P1_U4923 , P1_U3040 , P1_U3499 );
nand NAND2_2228 ( P1_U4924 , P1_R1162_U76 , P1_U3038 );
nand NAND2_2229 ( P1_U4925 , P1_ADDR_REG_16_ , P1_U4889 );
nand NAND2_2230 ( P1_U4926 , P1_R1105_U77 , P1_U3041 );
nand NAND2_2231 ( P1_U4927 , P1_U3039 , P1_U3496 );
nand NAND2_2232 ( P1_U4928 , P1_R1162_U77 , P1_U3037 );
nand NAND3_2233 ( P1_U4929 , P1_U4927 , P1_U4926 , P1_U4928 );
nand NAND2_2234 ( P1_U4930 , P1_U3043 , P1_U4929 );
nand NAND2_2235 ( P1_U4931 , P1_R1105_U77 , P1_U3042 );
nand NAND2_2236 ( P1_U4932 , P1_REG3_REG_15_ , P1_U3086 );
nand NAND2_2237 ( P1_U4933 , P1_U3040 , P1_U3496 );
nand NAND2_2238 ( P1_U4934 , P1_R1162_U77 , P1_U3038 );
nand NAND2_2239 ( P1_U4935 , P1_ADDR_REG_15_ , P1_U4889 );
nand NAND2_2240 ( P1_U4936 , P1_R1105_U78 , P1_U3041 );
nand NAND2_2241 ( P1_U4937 , P1_U3039 , P1_U3493 );
nand NAND2_2242 ( P1_U4938 , P1_R1162_U78 , P1_U3037 );
nand NAND3_2243 ( P1_U4939 , P1_U4937 , P1_U4936 , P1_U4938 );
nand NAND2_2244 ( P1_U4940 , P1_U3043 , P1_U4939 );
nand NAND2_2245 ( P1_U4941 , P1_R1105_U78 , P1_U3042 );
nand NAND2_2246 ( P1_U4942 , P1_REG3_REG_14_ , P1_U3086 );
nand NAND2_2247 ( P1_U4943 , P1_U3040 , P1_U3493 );
nand NAND2_2248 ( P1_U4944 , P1_R1162_U78 , P1_U3038 );
nand NAND2_2249 ( P1_U4945 , P1_ADDR_REG_14_ , P1_U4889 );
nand NAND2_2250 ( P1_U4946 , P1_R1105_U11 , P1_U3041 );
nand NAND2_2251 ( P1_U4947 , P1_U3039 , P1_U3490 );
nand NAND2_2252 ( P1_U4948 , P1_R1162_U11 , P1_U3037 );
nand NAND3_2253 ( P1_U4949 , P1_U4947 , P1_U4946 , P1_U4948 );
nand NAND2_2254 ( P1_U4950 , P1_U3043 , P1_U4949 );
nand NAND2_2255 ( P1_U4951 , P1_R1105_U11 , P1_U3042 );
nand NAND2_2256 ( P1_U4952 , P1_REG3_REG_13_ , P1_U3086 );
nand NAND2_2257 ( P1_U4953 , P1_U3040 , P1_U3490 );
nand NAND2_2258 ( P1_U4954 , P1_R1162_U11 , P1_U3038 );
nand NAND2_2259 ( P1_U4955 , P1_ADDR_REG_13_ , P1_U4889 );
nand NAND2_2260 ( P1_U4956 , P1_R1105_U79 , P1_U3041 );
nand NAND2_2261 ( P1_U4957 , P1_U3039 , P1_U3487 );
nand NAND2_2262 ( P1_U4958 , P1_R1162_U79 , P1_U3037 );
nand NAND3_2263 ( P1_U4959 , P1_U4957 , P1_U4956 , P1_U4958 );
nand NAND2_2264 ( P1_U4960 , P1_U3043 , P1_U4959 );
nand NAND2_2265 ( P1_U4961 , P1_R1105_U79 , P1_U3042 );
nand NAND2_2266 ( P1_U4962 , P1_REG3_REG_12_ , P1_U3086 );
nand NAND2_2267 ( P1_U4963 , P1_U3040 , P1_U3487 );
nand NAND2_2268 ( P1_U4964 , P1_R1162_U79 , P1_U3038 );
nand NAND2_2269 ( P1_U4965 , P1_ADDR_REG_12_ , P1_U4889 );
nand NAND2_2270 ( P1_U4966 , P1_R1105_U80 , P1_U3041 );
nand NAND2_2271 ( P1_U4967 , P1_U3039 , P1_U3484 );
nand NAND2_2272 ( P1_U4968 , P1_R1162_U80 , P1_U3037 );
nand NAND3_2273 ( P1_U4969 , P1_U4967 , P1_U4966 , P1_U4968 );
nand NAND2_2274 ( P1_U4970 , P1_U3043 , P1_U4969 );
nand NAND2_2275 ( P1_U4971 , P1_R1105_U80 , P1_U3042 );
nand NAND2_2276 ( P1_U4972 , P1_REG3_REG_11_ , P1_U3086 );
nand NAND2_2277 ( P1_U4973 , P1_U3040 , P1_U3484 );
nand NAND2_2278 ( P1_U4974 , P1_R1162_U80 , P1_U3038 );
nand NAND2_2279 ( P1_U4975 , P1_ADDR_REG_11_ , P1_U4889 );
nand NAND2_2280 ( P1_U4976 , P1_R1105_U10 , P1_U3041 );
nand NAND2_2281 ( P1_U4977 , P1_U3039 , P1_U3481 );
nand NAND2_2282 ( P1_U4978 , P1_R1162_U10 , P1_U3037 );
nand NAND3_2283 ( P1_U4979 , P1_U4977 , P1_U4976 , P1_U4978 );
nand NAND2_2284 ( P1_U4980 , P1_U3043 , P1_U4979 );
nand NAND2_2285 ( P1_U4981 , P1_R1105_U10 , P1_U3042 );
nand NAND2_2286 ( P1_U4982 , P1_REG3_REG_10_ , P1_U3086 );
nand NAND2_2287 ( P1_U4983 , P1_U3040 , P1_U3481 );
nand NAND2_2288 ( P1_U4984 , P1_R1162_U10 , P1_U3038 );
nand NAND2_2289 ( P1_U4985 , P1_ADDR_REG_10_ , P1_U4889 );
nand NAND2_2290 ( P1_U4986 , P1_R1105_U70 , P1_U3041 );
nand NAND2_2291 ( P1_U4987 , P1_U3039 , P1_U3478 );
nand NAND2_2292 ( P1_U4988 , P1_R1162_U70 , P1_U3037 );
nand NAND3_2293 ( P1_U4989 , P1_U4987 , P1_U4986 , P1_U4988 );
nand NAND2_2294 ( P1_U4990 , P1_U3043 , P1_U4989 );
nand NAND2_2295 ( P1_U4991 , P1_R1105_U70 , P1_U3042 );
nand NAND2_2296 ( P1_U4992 , P1_REG3_REG_9_ , P1_U3086 );
nand NAND2_2297 ( P1_U4993 , P1_U3040 , P1_U3478 );
nand NAND2_2298 ( P1_U4994 , P1_R1162_U70 , P1_U3038 );
nand NAND2_2299 ( P1_U4995 , P1_ADDR_REG_9_ , P1_U4889 );
nand NAND2_2300 ( P1_U4996 , P1_R1105_U71 , P1_U3041 );
nand NAND2_2301 ( P1_U4997 , P1_U3039 , P1_U3475 );
nand NAND2_2302 ( P1_U4998 , P1_R1162_U71 , P1_U3037 );
nand NAND3_2303 ( P1_U4999 , P1_U4997 , P1_U4996 , P1_U4998 );
nand NAND2_2304 ( P1_U5000 , P1_U3043 , P1_U4999 );
nand NAND2_2305 ( P1_U5001 , P1_R1105_U71 , P1_U3042 );
nand NAND2_2306 ( P1_U5002 , P1_REG3_REG_8_ , P1_U3086 );
nand NAND2_2307 ( P1_U5003 , P1_U3040 , P1_U3475 );
nand NAND2_2308 ( P1_U5004 , P1_R1162_U71 , P1_U3038 );
nand NAND2_2309 ( P1_U5005 , P1_ADDR_REG_8_ , P1_U4889 );
nand NAND2_2310 ( P1_U5006 , P1_R1105_U16 , P1_U3041 );
nand NAND2_2311 ( P1_U5007 , P1_U3039 , P1_U3472 );
nand NAND2_2312 ( P1_U5008 , P1_R1162_U16 , P1_U3037 );
nand NAND3_2313 ( P1_U5009 , P1_U5007 , P1_U5006 , P1_U5008 );
nand NAND2_2314 ( P1_U5010 , P1_U3043 , P1_U5009 );
nand NAND2_2315 ( P1_U5011 , P1_R1105_U16 , P1_U3042 );
nand NAND2_2316 ( P1_U5012 , P1_REG3_REG_7_ , P1_U3086 );
nand NAND2_2317 ( P1_U5013 , P1_U3040 , P1_U3472 );
nand NAND2_2318 ( P1_U5014 , P1_R1162_U16 , P1_U3038 );
nand NAND2_2319 ( P1_U5015 , P1_ADDR_REG_7_ , P1_U4889 );
nand NAND2_2320 ( P1_U5016 , P1_R1105_U72 , P1_U3041 );
nand NAND2_2321 ( P1_U5017 , P1_U3039 , P1_U3469 );
nand NAND2_2322 ( P1_U5018 , P1_R1162_U72 , P1_U3037 );
nand NAND3_2323 ( P1_U5019 , P1_U5017 , P1_U5016 , P1_U5018 );
nand NAND2_2324 ( P1_U5020 , P1_U3043 , P1_U5019 );
nand NAND2_2325 ( P1_U5021 , P1_R1105_U72 , P1_U3042 );
nand NAND2_2326 ( P1_U5022 , P1_REG3_REG_6_ , P1_U3086 );
nand NAND2_2327 ( P1_U5023 , P1_U3040 , P1_U3469 );
nand NAND2_2328 ( P1_U5024 , P1_R1162_U72 , P1_U3038 );
nand NAND2_2329 ( P1_U5025 , P1_ADDR_REG_6_ , P1_U4889 );
nand NAND2_2330 ( P1_U5026 , P1_R1105_U15 , P1_U3041 );
nand NAND2_2331 ( P1_U5027 , P1_U3039 , P1_U3466 );
nand NAND2_2332 ( P1_U5028 , P1_R1162_U15 , P1_U3037 );
nand NAND3_2333 ( P1_U5029 , P1_U5027 , P1_U5026 , P1_U5028 );
nand NAND2_2334 ( P1_U5030 , P1_U3043 , P1_U5029 );
nand NAND2_2335 ( P1_U5031 , P1_R1105_U15 , P1_U3042 );
nand NAND2_2336 ( P1_U5032 , P1_REG3_REG_5_ , P1_U3086 );
nand NAND2_2337 ( P1_U5033 , P1_U3040 , P1_U3466 );
nand NAND2_2338 ( P1_U5034 , P1_R1162_U15 , P1_U3038 );
nand NAND2_2339 ( P1_U5035 , P1_ADDR_REG_5_ , P1_U4889 );
nand NAND2_2340 ( P1_U5036 , P1_R1105_U73 , P1_U3041 );
nand NAND2_2341 ( P1_U5037 , P1_U3039 , P1_U3463 );
nand NAND2_2342 ( P1_U5038 , P1_R1162_U73 , P1_U3037 );
nand NAND3_2343 ( P1_U5039 , P1_U5037 , P1_U5036 , P1_U5038 );
nand NAND2_2344 ( P1_U5040 , P1_U3043 , P1_U5039 );
nand NAND2_2345 ( P1_U5041 , P1_R1105_U73 , P1_U3042 );
nand NAND2_2346 ( P1_U5042 , P1_REG3_REG_4_ , P1_U3086 );
nand NAND2_2347 ( P1_U5043 , P1_U3040 , P1_U3463 );
nand NAND2_2348 ( P1_U5044 , P1_R1162_U73 , P1_U3038 );
nand NAND2_2349 ( P1_U5045 , P1_ADDR_REG_4_ , P1_U4889 );
nand NAND2_2350 ( P1_U5046 , P1_R1105_U74 , P1_U3041 );
nand NAND2_2351 ( P1_U5047 , P1_U3039 , P1_U3460 );
nand NAND2_2352 ( P1_U5048 , P1_R1162_U74 , P1_U3037 );
nand NAND3_2353 ( P1_U5049 , P1_U5047 , P1_U5046 , P1_U5048 );
nand NAND2_2354 ( P1_U5050 , P1_U3043 , P1_U5049 );
nand NAND2_2355 ( P1_U5051 , P1_R1105_U74 , P1_U3042 );
nand NAND2_2356 ( P1_U5052 , P1_REG3_REG_3_ , P1_U3086 );
nand NAND2_2357 ( P1_U5053 , P1_U3040 , P1_U3460 );
nand NAND2_2358 ( P1_U5054 , P1_R1162_U74 , P1_U3038 );
nand NAND2_2359 ( P1_U5055 , P1_ADDR_REG_3_ , P1_U4889 );
nand NAND2_2360 ( P1_U5056 , P1_R1105_U14 , P1_U3041 );
nand NAND2_2361 ( P1_U5057 , P1_U3039 , P1_U3457 );
nand NAND2_2362 ( P1_U5058 , P1_R1162_U14 , P1_U3037 );
nand NAND3_2363 ( P1_U5059 , P1_U5057 , P1_U5056 , P1_U5058 );
nand NAND2_2364 ( P1_U5060 , P1_U3043 , P1_U5059 );
nand NAND2_2365 ( P1_U5061 , P1_R1105_U14 , P1_U3042 );
nand NAND2_2366 ( P1_U5062 , P1_REG3_REG_2_ , P1_U3086 );
nand NAND2_2367 ( P1_U5063 , P1_U3040 , P1_U3457 );
nand NAND2_2368 ( P1_U5064 , P1_R1162_U14 , P1_U3038 );
nand NAND2_2369 ( P1_U5065 , P1_ADDR_REG_2_ , P1_U4889 );
nand NAND2_2370 ( P1_U5066 , P1_R1105_U68 , P1_U3041 );
nand NAND2_2371 ( P1_U5067 , P1_U3039 , P1_U3454 );
nand NAND2_2372 ( P1_U5068 , P1_R1162_U68 , P1_U3037 );
nand NAND3_2373 ( P1_U5069 , P1_U5067 , P1_U5066 , P1_U5068 );
nand NAND2_2374 ( P1_U5070 , P1_U3043 , P1_U5069 );
nand NAND2_2375 ( P1_U5071 , P1_R1105_U68 , P1_U3042 );
nand NAND2_2376 ( P1_U5072 , P1_REG3_REG_1_ , P1_U3086 );
nand NAND2_2377 ( P1_U5073 , P1_U3040 , P1_U3454 );
nand NAND2_2378 ( P1_U5074 , P1_R1162_U68 , P1_U3038 );
nand NAND2_2379 ( P1_U5075 , P1_ADDR_REG_1_ , P1_U4889 );
nand NAND2_2380 ( P1_U5076 , P1_R1105_U69 , P1_U3041 );
nand NAND2_2381 ( P1_U5077 , P1_U3039 , P1_U3448 );
nand NAND2_2382 ( P1_U5078 , P1_R1162_U69 , P1_U3037 );
nand NAND3_2383 ( P1_U5079 , P1_U5077 , P1_U5076 , P1_U5078 );
nand NAND2_2384 ( P1_U5080 , P1_U3043 , P1_U5079 );
nand NAND2_2385 ( P1_U5081 , P1_R1105_U69 , P1_U3042 );
nand NAND2_2386 ( P1_U5082 , P1_REG3_REG_0_ , P1_U3086 );
nand NAND2_2387 ( P1_U5083 , P1_U3040 , P1_U3448 );
nand NAND2_2388 ( P1_U5084 , P1_R1162_U69 , P1_U3038 );
nand NAND2_2389 ( P1_U5085 , P1_ADDR_REG_0_ , P1_U4889 );
not NOT1_2390 ( P1_U5086 , P1_U3951 );
nand NAND3_2391 ( P1_U5087 , P1_U3954 , P1_U3987 , P1_LT_197_U13 );
nand NAND2_2392 ( P1_U5088 , P1_U5677 , P1_U3427 );
nand NAND2_2393 ( P1_U5089 , P1_U3851 , P1_U5088 );
nand NAND3_2394 ( P1_U5090 , P1_U3022 , P1_U3986 , P1_U3949 );
nand NAND2_2395 ( P1_U5091 , P1_B_REG , P1_U5089 );
nand NAND2_2396 ( P1_U5092 , P1_U3036 , P1_U3079 );
nand NAND2_2397 ( P1_U5093 , P1_U3034 , P1_U3073 );
nand NAND2_2398 ( P1_U5094 , P1_ADD_95_U73 , P1_U3430 );
nand NAND3_2399 ( P1_U5095 , P1_U5094 , P1_U5092 , P1_U5093 );
nand NAND3_2400 ( P1_U5096 , P1_U3364 , P1_U3361 , P1_U3362 );
nand NAND3_2401 ( P1_U5097 , P1_U3366 , P1_U3419 , P1_U3365 );
nand NAND2_2402 ( P1_U5098 , P1_U5684 , P1_U5097 );
nand NAND2_2403 ( P1_U5099 , P1_U5693 , P1_U5096 );
nand NAND3_2404 ( P1_U5100 , P1_U5099 , P1_U5098 , P1_U3868 );
nand NAND2_2405 ( P1_U5101 , P1_U5100 , P1_U3430 );
not NOT1_2406 ( P1_U5102 , P1_U3432 );
nand NAND2_2407 ( P1_U5103 , P1_U3497 , P1_U5656 );
nand NAND2_2408 ( P1_U5104 , P1_ADD_95_U73 , P1_U5655 );
nand NAND2_2409 ( P1_U5105 , P1_U3994 , P1_U5095 );
nand NAND2_2410 ( P1_U5106 , P1_R1165_U104 , P1_U3027 );
nand NAND2_2411 ( P1_U5107 , P1_REG3_REG_15_ , P1_U3086 );
nand NAND2_2412 ( P1_U5108 , P1_U3036 , P1_U3058 );
nand NAND2_2413 ( P1_U5109 , P1_U3034 , P1_U3053 );
nand NAND2_2414 ( P1_U5110 , P1_ADD_95_U62 , P1_U3430 );
nand NAND3_2415 ( P1_U5111 , P1_U5110 , P1_U5108 , P1_U5109 );
nand NAND2_2416 ( P1_U5112 , P1_U3422 , P1_U3430 );
nand NAND2_2417 ( P1_U5113 , P1_U5102 , P1_U5112 );
nand NAND2_2418 ( P1_U5114 , P1_U3972 , P1_U3422 );
nand NAND2_2419 ( P1_U5115 , P1_U3418 , P1_U5114 );
nand NAND2_2420 ( P1_U5116 , P1_U3045 , P1_U3976 );
nand NAND2_2421 ( P1_U5117 , P1_U3044 , P1_ADD_95_U62 );
nand NAND2_2422 ( P1_U5118 , P1_U3994 , P1_U5111 );
nand NAND2_2423 ( P1_U5119 , P1_R1165_U13 , P1_U3027 );
nand NAND2_2424 ( P1_U5120 , P1_REG3_REG_26_ , P1_U3086 );
nand NAND2_2425 ( P1_U5121 , P1_U3036 , P1_U3067 );
nand NAND2_2426 ( P1_U5122 , P1_U3034 , P1_U3070 );
nand NAND2_2427 ( P1_U5123 , P1_ADD_95_U57 , P1_U3430 );
nand NAND3_2428 ( P1_U5124 , P1_U5122 , P1_U5121 , P1_U5123 );
nand NAND2_2429 ( P1_U5125 , P1_U3470 , P1_U5656 );
nand NAND2_2430 ( P1_U5126 , P1_ADD_95_U57 , P1_U5655 );
nand NAND2_2431 ( P1_U5127 , P1_U3994 , P1_U5124 );
nand NAND2_2432 ( P1_U5128 , P1_R1165_U89 , P1_U3027 );
nand NAND2_2433 ( P1_U5129 , P1_REG3_REG_6_ , P1_U3086 );
nand NAND2_2434 ( P1_U5130 , P1_U3036 , P1_U3069 );
nand NAND2_2435 ( P1_U5131 , P1_U3034 , P1_U3081 );
nand NAND2_2436 ( P1_U5132 , P1_ADD_95_U70 , P1_U3430 );
nand NAND3_2437 ( P1_U5133 , P1_U5132 , P1_U5130 , P1_U5131 );
nand NAND2_2438 ( P1_U5134 , P1_U3506 , P1_U5656 );
nand NAND2_2439 ( P1_U5135 , P1_ADD_95_U70 , P1_U5655 );
nand NAND2_2440 ( P1_U5136 , P1_U3994 , P1_U5133 );
nand NAND2_2441 ( P1_U5137 , P1_R1165_U102 , P1_U3027 );
nand NAND2_2442 ( P1_U5138 , P1_REG3_REG_18_ , P1_U3086 );
nand NAND2_2443 ( P1_U5139 , P1_U3036 , P1_U3078 );
nand NAND2_2444 ( P1_U5140 , P1_U3034 , P1_U3064 );
nand NAND2_2445 ( P1_U5141 , P1_REG3_REG_2_ , P1_U3430 );
nand NAND3_2446 ( P1_U5142 , P1_U5140 , P1_U5139 , P1_U5141 );
nand NAND2_2447 ( P1_U5143 , P1_U3458 , P1_U5656 );
nand NAND2_2448 ( P1_U5144 , P1_REG3_REG_2_ , P1_U5655 );
nand NAND2_2449 ( P1_U5145 , P1_U3994 , P1_U5142 );
nand NAND2_2450 ( P1_U5146 , P1_R1165_U92 , P1_U3027 );
nand NAND2_2451 ( P1_U5147 , P1_REG3_REG_2_ , P1_U3086 );
nand NAND2_2452 ( P1_U5148 , P1_U3036 , P1_U3062 );
nand NAND2_2453 ( P1_U5149 , P1_U3034 , P1_U3072 );
nand NAND2_2454 ( P1_U5150 , P1_ADD_95_U77 , P1_U3430 );
nand NAND3_2455 ( P1_U5151 , P1_U5149 , P1_U5148 , P1_U5150 );
nand NAND2_2456 ( P1_U5152 , P1_U3485 , P1_U5656 );
nand NAND2_2457 ( P1_U5153 , P1_ADD_95_U77 , P1_U5655 );
nand NAND2_2458 ( P1_U5154 , P1_U3994 , P1_U5151 );
nand NAND2_2459 ( P1_U5155 , P1_R1165_U107 , P1_U3027 );
nand NAND2_2460 ( P1_U5156 , P1_REG3_REG_11_ , P1_U3086 );
nand NAND2_2461 ( P1_U5157 , P1_U3036 , P1_U3075 );
nand NAND2_2462 ( P1_U5158 , P1_U3034 , P1_U3066 );
nand NAND2_2463 ( P1_U5159 , P1_ADD_95_U66 , P1_U3430 );
nand NAND3_2464 ( P1_U5160 , P1_U5159 , P1_U5157 , P1_U5158 );
nand NAND2_2465 ( P1_U5161 , P1_U3045 , P1_U3980 );
nand NAND2_2466 ( P1_U5162 , P1_U3044 , P1_ADD_95_U66 );
nand NAND2_2467 ( P1_U5163 , P1_U3994 , P1_U5160 );
nand NAND2_2468 ( P1_U5164 , P1_R1165_U98 , P1_U3027 );
nand NAND2_2469 ( P1_U5165 , P1_REG3_REG_22_ , P1_U3086 );
nand NAND2_2470 ( P1_U5166 , P1_U3036 , P1_U3072 );
nand NAND2_2471 ( P1_U5167 , P1_U3034 , P1_U3079 );
nand NAND2_2472 ( P1_U5168 , P1_ADD_95_U75 , P1_U3430 );
nand NAND3_2473 ( P1_U5169 , P1_U5168 , P1_U5166 , P1_U5167 );
nand NAND2_2474 ( P1_U5170 , P1_U3491 , P1_U5656 );
nand NAND2_2475 ( P1_U5171 , P1_ADD_95_U75 , P1_U5655 );
nand NAND2_2476 ( P1_U5172 , P1_U3994 , P1_U5169 );
nand NAND2_2477 ( P1_U5173 , P1_R1165_U10 , P1_U3027 );
nand NAND2_2478 ( P1_U5174 , P1_REG3_REG_13_ , P1_U3086 );
nand NAND2_2479 ( P1_U5175 , P1_U3036 , P1_U3081 );
nand NAND2_2480 ( P1_U5176 , P1_U3034 , P1_U3075 );
nand NAND2_2481 ( P1_U5177 , P1_ADD_95_U68 , P1_U3430 );
nand NAND3_2482 ( P1_U5178 , P1_U5177 , P1_U5175 , P1_U5176 );
nand NAND2_2483 ( P1_U5179 , P1_U3045 , P1_U3982 );
nand NAND2_2484 ( P1_U5180 , P1_U3044 , P1_ADD_95_U68 );
nand NAND2_2485 ( P1_U5181 , P1_U3994 , P1_U5178 );
nand NAND2_2486 ( P1_U5182 , P1_R1165_U99 , P1_U3027 );
nand NAND2_2487 ( P1_U5183 , P1_REG3_REG_20_ , P1_U3086 );
nand NAND2_2488 ( P1_U5184 , P1_U3431 , P1_U3429 );
nand NAND2_2489 ( P1_U5185 , P1_U5184 , P1_U3430 );
nand NAND2_2490 ( P1_U5186 , P1_U3995 , P1_U5185 );
nand NAND2_2491 ( P1_U5187 , P1_U3873 , P1_U3034 );
nand NAND2_2492 ( P1_U5188 , P1_U3450 , P1_U5656 );
nand NAND2_2493 ( P1_U5189 , P1_REG3_REG_0_ , P1_U5186 );
nand NAND2_2494 ( P1_U5190 , P1_R1165_U86 , P1_U3027 );
nand NAND2_2495 ( P1_U5191 , P1_REG3_REG_0_ , P1_U3086 );
nand NAND2_2496 ( P1_U5192 , P1_U3036 , P1_U3084 );
nand NAND2_2497 ( P1_U5193 , P1_U3034 , P1_U3062 );
nand NAND2_2498 ( P1_U5194 , P1_ADD_95_U54 , P1_U3430 );
nand NAND3_2499 ( P1_U5195 , P1_U5193 , P1_U5192 , P1_U5194 );
nand NAND2_2500 ( P1_U5196 , P1_U3479 , P1_U5656 );
nand NAND2_2501 ( P1_U5197 , P1_ADD_95_U54 , P1_U5655 );
nand NAND2_2502 ( P1_U5198 , P1_U3994 , P1_U5195 );
nand NAND2_2503 ( P1_U5199 , P1_R1165_U87 , P1_U3027 );
nand NAND2_2504 ( P1_U5200 , P1_REG3_REG_9_ , P1_U3086 );
nand NAND2_2505 ( P1_U5201 , P1_U3036 , P1_U3064 );
nand NAND2_2506 ( P1_U5202 , P1_U3034 , P1_U3067 );
nand NAND2_2507 ( P1_U5203 , P1_ADD_95_U59 , P1_U3430 );
nand NAND3_2508 ( P1_U5204 , P1_U5202 , P1_U5201 , P1_U5203 );
nand NAND2_2509 ( P1_U5205 , P1_U3464 , P1_U5656 );
nand NAND2_2510 ( P1_U5206 , P1_ADD_95_U59 , P1_U5655 );
nand NAND2_2511 ( P1_U5207 , P1_U3994 , P1_U5204 );
nand NAND2_2512 ( P1_U5208 , P1_R1165_U91 , P1_U3027 );
nand NAND2_2513 ( P1_U5209 , P1_REG3_REG_4_ , P1_U3086 );
nand NAND2_2514 ( P1_U5210 , P1_U3036 , P1_U3066 );
nand NAND2_2515 ( P1_U5211 , P1_U3034 , P1_U3058 );
nand NAND2_2516 ( P1_U5212 , P1_ADD_95_U64 , P1_U3430 );
nand NAND3_2517 ( P1_U5213 , P1_U5212 , P1_U5210 , P1_U5211 );
nand NAND2_2518 ( P1_U5214 , P1_U3045 , P1_U3978 );
nand NAND2_2519 ( P1_U5215 , P1_U3044 , P1_ADD_95_U64 );
nand NAND2_2520 ( P1_U5216 , P1_U3994 , P1_U5213 );
nand NAND2_2521 ( P1_U5217 , P1_R1165_U96 , P1_U3027 );
nand NAND2_2522 ( P1_U5218 , P1_REG3_REG_24_ , P1_U3086 );
nand NAND2_2523 ( P1_U5219 , P1_U3036 , P1_U3073 );
nand NAND2_2524 ( P1_U5220 , P1_U3034 , P1_U3082 );
nand NAND2_2525 ( P1_U5221 , P1_ADD_95_U71 , P1_U3430 );
nand NAND3_2526 ( P1_U5222 , P1_U5221 , P1_U5219 , P1_U5220 );
nand NAND2_2527 ( P1_U5223 , P1_U3503 , P1_U5656 );
nand NAND2_2528 ( P1_U5224 , P1_ADD_95_U71 , P1_U5655 );
nand NAND2_2529 ( P1_U5225 , P1_U3994 , P1_U5222 );
nand NAND2_2530 ( P1_U5226 , P1_R1165_U11 , P1_U3027 );
nand NAND2_2531 ( P1_U5227 , P1_REG3_REG_17_ , P1_U3086 );
nand NAND2_2532 ( P1_U5228 , P1_U3036 , P1_U3060 );
nand NAND2_2533 ( P1_U5229 , P1_U3034 , P1_U3071 );
nand NAND2_2534 ( P1_U5230 , P1_ADD_95_U58 , P1_U3430 );
nand NAND3_2535 ( P1_U5231 , P1_U5229 , P1_U5228 , P1_U5230 );
nand NAND2_2536 ( P1_U5232 , P1_U3467 , P1_U5656 );
nand NAND2_2537 ( P1_U5233 , P1_ADD_95_U58 , P1_U5655 );
nand NAND2_2538 ( P1_U5234 , P1_U3994 , P1_U5231 );
nand NAND2_2539 ( P1_U5235 , P1_R1165_U90 , P1_U3027 );
nand NAND2_2540 ( P1_U5236 , P1_REG3_REG_5_ , P1_U3086 );
nand NAND2_2541 ( P1_U5237 , P1_U3036 , P1_U3074 );
nand NAND2_2542 ( P1_U5238 , P1_U3034 , P1_U3069 );
nand NAND2_2543 ( P1_U5239 , P1_ADD_95_U72 , P1_U3430 );
nand NAND3_2544 ( P1_U5240 , P1_U5239 , P1_U5237 , P1_U5238 );
nand NAND2_2545 ( P1_U5241 , P1_U3500 , P1_U5656 );
nand NAND2_2546 ( P1_U5242 , P1_ADD_95_U72 , P1_U5655 );
nand NAND2_2547 ( P1_U5243 , P1_U3994 , P1_U5240 );
nand NAND2_2548 ( P1_U5244 , P1_R1165_U103 , P1_U3027 );
nand NAND2_2549 ( P1_U5245 , P1_REG3_REG_16_ , P1_U3086 );
nand NAND2_2550 ( P1_U5246 , P1_U3036 , P1_U3065 );
nand NAND2_2551 ( P1_U5247 , P1_U3034 , P1_U3057 );
nand NAND2_2552 ( P1_U5248 , P1_ADD_95_U63 , P1_U3430 );
nand NAND3_2553 ( P1_U5249 , P1_U5248 , P1_U5246 , P1_U5247 );
nand NAND2_2554 ( P1_U5250 , P1_U3045 , P1_U3977 );
nand NAND2_2555 ( P1_U5251 , P1_U3044 , P1_ADD_95_U63 );
nand NAND2_2556 ( P1_U5252 , P1_U3994 , P1_U5249 );
nand NAND2_2557 ( P1_U5253 , P1_R1165_U95 , P1_U3027 );
nand NAND2_2558 ( P1_U5254 , P1_REG3_REG_25_ , P1_U3086 );
nand NAND2_2559 ( P1_U5255 , P1_U3036 , P1_U3063 );
nand NAND2_2560 ( P1_U5256 , P1_U3034 , P1_U3080 );
nand NAND2_2561 ( P1_U5257 , P1_ADD_95_U76 , P1_U3430 );
nand NAND3_2562 ( P1_U5258 , P1_U5257 , P1_U5255 , P1_U5256 );
nand NAND2_2563 ( P1_U5259 , P1_U3488 , P1_U5656 );
nand NAND2_2564 ( P1_U5260 , P1_ADD_95_U76 , P1_U5655 );
nand NAND2_2565 ( P1_U5261 , P1_U3994 , P1_U5258 );
nand NAND2_2566 ( P1_U5262 , P1_R1165_U106 , P1_U3027 );
nand NAND2_2567 ( P1_U5263 , P1_REG3_REG_12_ , P1_U3086 );
nand NAND2_2568 ( P1_U5264 , P1_U3036 , P1_U3076 );
nand NAND2_2569 ( P1_U5265 , P1_U3034 , P1_U3061 );
nand NAND2_2570 ( P1_U5266 , P1_ADD_95_U67 , P1_U3430 );
nand NAND3_2571 ( P1_U5267 , P1_U5266 , P1_U5264 , P1_U5265 );
nand NAND2_2572 ( P1_U5268 , P1_U3045 , P1_U3981 );
nand NAND2_2573 ( P1_U5269 , P1_U3044 , P1_ADD_95_U67 );
nand NAND2_2574 ( P1_U5270 , P1_U3994 , P1_U5267 );
nand NAND2_2575 ( P1_U5271 , P1_R1165_U12 , P1_U3027 );
nand NAND2_2576 ( P1_U5272 , P1_REG3_REG_21_ , P1_U3086 );
nand NAND2_2577 ( P1_U5273 , P1_U3036 , P1_U3077 );
nand NAND2_2578 ( P1_U5274 , P1_U3034 , P1_U3068 );
nand NAND2_2579 ( P1_U5275 , P1_REG3_REG_1_ , P1_U3430 );
nand NAND3_2580 ( P1_U5276 , P1_U5274 , P1_U5273 , P1_U5275 );
nand NAND2_2581 ( P1_U5277 , P1_U3455 , P1_U5656 );
nand NAND2_2582 ( P1_U5278 , P1_REG3_REG_1_ , P1_U5655 );
nand NAND2_2583 ( P1_U5279 , P1_U3994 , P1_U5276 );
nand NAND2_2584 ( P1_U5280 , P1_R1165_U100 , P1_U3027 );
nand NAND2_2585 ( P1_U5281 , P1_REG3_REG_1_ , P1_U3086 );
nand NAND2_2586 ( P1_U5282 , P1_U3036 , P1_U3070 );
nand NAND2_2587 ( P1_U5283 , P1_U3034 , P1_U3083 );
nand NAND2_2588 ( P1_U5284 , P1_ADD_95_U55 , P1_U3430 );
nand NAND3_2589 ( P1_U5285 , P1_U5283 , P1_U5282 , P1_U5284 );
nand NAND2_2590 ( P1_U5286 , P1_U3476 , P1_U5656 );
nand NAND2_2591 ( P1_U5287 , P1_ADD_95_U55 , P1_U5655 );
nand NAND2_2592 ( P1_U5288 , P1_U3994 , P1_U5285 );
nand NAND2_2593 ( P1_U5289 , P1_R1165_U88 , P1_U3027 );
nand NAND2_2594 ( P1_U5290 , P1_REG3_REG_8_ , P1_U3086 );
nand NAND2_2595 ( P1_U5291 , P1_U3036 , P1_U3053 );
nand NAND2_2596 ( P1_U5292 , P1_U3034 , P1_U3055 );
nand NAND2_2597 ( P1_U5293 , P1_ADD_95_U60 , P1_U3430 );
nand NAND3_2598 ( P1_U5294 , P1_U5292 , P1_U5291 , P1_U5293 );
nand NAND2_2599 ( P1_U5295 , P1_U3045 , P1_U3974 );
nand NAND2_2600 ( P1_U5296 , P1_U3044 , P1_ADD_95_U60 );
nand NAND2_2601 ( P1_U5297 , P1_U3994 , P1_U5294 );
nand NAND2_2602 ( P1_U5298 , P1_R1165_U93 , P1_U3027 );
nand NAND2_2603 ( P1_U5299 , P1_REG3_REG_28_ , P1_U3086 );
nand NAND2_2604 ( P1_U5300 , P1_U3036 , P1_U3082 );
nand NAND2_2605 ( P1_U5301 , P1_U3034 , P1_U3076 );
nand NAND2_2606 ( P1_U5302 , P1_ADD_95_U69 , P1_U3430 );
nand NAND3_2607 ( P1_U5303 , P1_U5302 , P1_U5300 , P1_U5301 );
nand NAND2_2608 ( P1_U5304 , P1_U3508 , P1_U5656 );
nand NAND2_2609 ( P1_U5305 , P1_ADD_95_U69 , P1_U5655 );
nand NAND2_2610 ( P1_U5306 , P1_U3994 , P1_U5303 );
nand NAND2_2611 ( P1_U5307 , P1_R1165_U101 , P1_U3027 );
nand NAND2_2612 ( P1_U5308 , P1_REG3_REG_19_ , P1_U3086 );
nand NAND2_2613 ( P1_U5309 , P1_U3036 , P1_U3068 );
nand NAND2_2614 ( P1_U5310 , P1_U3034 , P1_U3060 );
nand NAND2_2615 ( P1_U5311 , P1_ADD_95_U4 , P1_U3430 );
nand NAND3_2616 ( P1_U5312 , P1_U5310 , P1_U5309 , P1_U5311 );
nand NAND2_2617 ( P1_U5313 , P1_U3461 , P1_U5656 );
nand NAND2_2618 ( P1_U5314 , P1_ADD_95_U4 , P1_U5655 );
nand NAND2_2619 ( P1_U5315 , P1_U3994 , P1_U5312 );
nand NAND2_2620 ( P1_U5316 , P1_R1165_U14 , P1_U3027 );
nand NAND2_2621 ( P1_U5317 , P1_REG3_REG_3_ , P1_U3086 );
nand NAND2_2622 ( P1_U5318 , P1_U3036 , P1_U3083 );
nand NAND2_2623 ( P1_U5319 , P1_U3034 , P1_U3063 );
nand NAND2_2624 ( P1_U5320 , P1_ADD_95_U78 , P1_U3430 );
nand NAND3_2625 ( P1_U5321 , P1_U5319 , P1_U5318 , P1_U5320 );
nand NAND2_2626 ( P1_U5322 , P1_U3482 , P1_U5656 );
nand NAND2_2627 ( P1_U5323 , P1_ADD_95_U78 , P1_U5655 );
nand NAND2_2628 ( P1_U5324 , P1_U3994 , P1_U5321 );
nand NAND2_2629 ( P1_U5325 , P1_R1165_U108 , P1_U3027 );
nand NAND2_2630 ( P1_U5326 , P1_REG3_REG_10_ , P1_U3086 );
nand NAND2_2631 ( P1_U5327 , P1_U3036 , P1_U3061 );
nand NAND2_2632 ( P1_U5328 , P1_U3034 , P1_U3065 );
nand NAND2_2633 ( P1_U5329 , P1_ADD_95_U65 , P1_U3430 );
nand NAND3_2634 ( P1_U5330 , P1_U5329 , P1_U5327 , P1_U5328 );
nand NAND2_2635 ( P1_U5331 , P1_U3045 , P1_U3979 );
nand NAND2_2636 ( P1_U5332 , P1_U3044 , P1_ADD_95_U65 );
nand NAND2_2637 ( P1_U5333 , P1_U3994 , P1_U5330 );
nand NAND2_2638 ( P1_U5334 , P1_R1165_U97 , P1_U3027 );
nand NAND2_2639 ( P1_U5335 , P1_REG3_REG_23_ , P1_U3086 );
nand NAND2_2640 ( P1_U5336 , P1_U3036 , P1_U3080 );
nand NAND2_2641 ( P1_U5337 , P1_U3034 , P1_U3074 );
nand NAND2_2642 ( P1_U5338 , P1_ADD_95_U74 , P1_U3430 );
nand NAND3_2643 ( P1_U5339 , P1_U5338 , P1_U5336 , P1_U5337 );
nand NAND2_2644 ( P1_U5340 , P1_U3494 , P1_U5656 );
nand NAND2_2645 ( P1_U5341 , P1_ADD_95_U74 , P1_U5655 );
nand NAND2_2646 ( P1_U5342 , P1_U3994 , P1_U5339 );
nand NAND2_2647 ( P1_U5343 , P1_R1165_U105 , P1_U3027 );
nand NAND2_2648 ( P1_U5344 , P1_REG3_REG_14_ , P1_U3086 );
nand NAND2_2649 ( P1_U5345 , P1_U3036 , P1_U3057 );
nand NAND2_2650 ( P1_U5346 , P1_U3034 , P1_U3054 );
nand NAND2_2651 ( P1_U5347 , P1_ADD_95_U61 , P1_U3430 );
nand NAND3_2652 ( P1_U5348 , P1_U5347 , P1_U5345 , P1_U5346 );
nand NAND2_2653 ( P1_U5349 , P1_U3045 , P1_U3975 );
nand NAND2_2654 ( P1_U5350 , P1_U3044 , P1_ADD_95_U61 );
nand NAND2_2655 ( P1_U5351 , P1_U3994 , P1_U5348 );
nand NAND2_2656 ( P1_U5352 , P1_R1165_U94 , P1_U3027 );
nand NAND2_2657 ( P1_U5353 , P1_REG3_REG_27_ , P1_U3086 );
nand NAND2_2658 ( P1_U5354 , P1_U3036 , P1_U3071 );
nand NAND2_2659 ( P1_U5355 , P1_U3034 , P1_U3084 );
nand NAND2_2660 ( P1_U5356 , P1_ADD_95_U56 , P1_U3430 );
nand NAND3_2661 ( P1_U5357 , P1_U5355 , P1_U5354 , P1_U5356 );
nand NAND2_2662 ( P1_U5358 , P1_U3473 , P1_U5656 );
nand NAND2_2663 ( P1_U5359 , P1_ADD_95_U56 , P1_U5655 );
nand NAND2_2664 ( P1_U5360 , P1_U3994 , P1_U5357 );
nand NAND2_2665 ( P1_U5361 , P1_R1165_U15 , P1_U3027 );
nand NAND2_2666 ( P1_U5362 , P1_REG3_REG_7_ , P1_U3086 );
nand NAND2_2667 ( P1_U5363 , P1_U3449 , P1_U3375 );
nand NAND2_2668 ( P1_U5364 , P1_U3446 , P1_U5363 );
nand NAND3_2669 ( P1_U5365 , P1_U5702 , P1_U3446 , P1_R1165_U86 );
nand NAND2_2670 ( P1_U5366 , P1_U3447 , P1_U3441 );
nand NAND2_2671 ( P1_U5367 , P1_U3877 , P1_U3970 );
nand NAND2_2672 ( P1_U5368 , P1_U3370 , P1_U3419 );
nand NAND3_2673 ( P1_U5369 , P1_U3368 , P1_U3363 , P1_U3365 );
nand NAND2_2674 ( P1_U5370 , P1_U4000 , P1_U3421 );
nand NAND2_2675 ( P1_U5371 , P1_U5369 , P1_U3421 );
not NOT1_2676 ( P1_U5372 , P1_U3434 );
nand NAND2_2677 ( P1_U5373 , P1_U5372 , P1_U3970 );
nand NAND2_2678 ( P1_U5374 , P1_U3479 , P1_U5373 );
nand NAND2_2679 ( P1_U5375 , P1_U3021 , P1_U3083 );
nand NAND2_2680 ( P1_U5376 , P1_U3476 , P1_U5373 );
nand NAND2_2681 ( P1_U5377 , P1_U3021 , P1_U3084 );
nand NAND2_2682 ( P1_U5378 , P1_U3473 , P1_U5373 );
nand NAND2_2683 ( P1_U5379 , P1_U3021 , P1_U3070 );
nand NAND2_2684 ( P1_U5380 , P1_U3470 , P1_U5373 );
nand NAND2_2685 ( P1_U5381 , P1_U3021 , P1_U3071 );
nand NAND2_2686 ( P1_U5382 , P1_U3467 , P1_U5373 );
nand NAND2_2687 ( P1_U5383 , P1_U3021 , P1_U3067 );
nand NAND2_2688 ( P1_U5384 , P1_U3464 , P1_U5373 );
nand NAND2_2689 ( P1_U5385 , P1_U3021 , P1_U3060 );
nand NAND2_2690 ( P1_U5386 , P1_U3461 , P1_U5373 );
nand NAND2_2691 ( P1_U5387 , P1_U3021 , P1_U3064 );
nand NAND2_2692 ( P1_U5388 , P1_U3974 , P1_U5373 );
nand NAND2_2693 ( P1_U5389 , P1_U3021 , P1_U3054 );
nand NAND2_2694 ( P1_U5390 , P1_U3975 , P1_U5373 );
nand NAND2_2695 ( P1_U5391 , P1_U3021 , P1_U3053 );
nand NAND2_2696 ( P1_U5392 , P1_U3976 , P1_U5373 );
nand NAND2_2697 ( P1_U5393 , P1_U3021 , P1_U3057 );
nand NAND2_2698 ( P1_U5394 , P1_U3977 , P1_U5373 );
nand NAND2_2699 ( P1_U5395 , P1_U3021 , P1_U3058 );
nand NAND2_2700 ( P1_U5396 , P1_U3978 , P1_U5373 );
nand NAND2_2701 ( P1_U5397 , P1_U3021 , P1_U3065 );
nand NAND2_2702 ( P1_U5398 , P1_U3979 , P1_U5373 );
nand NAND2_2703 ( P1_U5399 , P1_U3021 , P1_U3066 );
nand NAND2_2704 ( P1_U5400 , P1_U3980 , P1_U5373 );
nand NAND2_2705 ( P1_U5401 , P1_U3021 , P1_U3061 );
nand NAND2_2706 ( P1_U5402 , P1_U3981 , P1_U5373 );
nand NAND2_2707 ( P1_U5403 , P1_U3021 , P1_U3075 );
nand NAND2_2708 ( P1_U5404 , P1_U3982 , P1_U5373 );
nand NAND2_2709 ( P1_U5405 , P1_U3021 , P1_U3076 );
nand NAND2_2710 ( P1_U5406 , P1_U3458 , P1_U5373 );
nand NAND2_2711 ( P1_U5407 , P1_U3021 , P1_U3068 );
nand NAND2_2712 ( P1_U5408 , P1_U3508 , P1_U5373 );
nand NAND2_2713 ( P1_U5409 , P1_U3021 , P1_U3081 );
nand NAND2_2714 ( P1_U5410 , P1_U3506 , P1_U5373 );
nand NAND2_2715 ( P1_U5411 , P1_U3021 , P1_U3082 );
nand NAND2_2716 ( P1_U5412 , P1_U3503 , P1_U5373 );
nand NAND2_2717 ( P1_U5413 , P1_U3021 , P1_U3069 );
nand NAND2_2718 ( P1_U5414 , P1_U3500 , P1_U5373 );
nand NAND2_2719 ( P1_U5415 , P1_U3021 , P1_U3073 );
nand NAND2_2720 ( P1_U5416 , P1_U3497 , P1_U5373 );
nand NAND2_2721 ( P1_U5417 , P1_U3021 , P1_U3074 );
nand NAND2_2722 ( P1_U5418 , P1_U3494 , P1_U5373 );
nand NAND2_2723 ( P1_U5419 , P1_U3021 , P1_U3079 );
nand NAND2_2724 ( P1_U5420 , P1_U3491 , P1_U5373 );
nand NAND2_2725 ( P1_U5421 , P1_U3021 , P1_U3080 );
nand NAND2_2726 ( P1_U5422 , P1_U3488 , P1_U5373 );
nand NAND2_2727 ( P1_U5423 , P1_U3021 , P1_U3072 );
nand NAND2_2728 ( P1_U5424 , P1_U3485 , P1_U5373 );
nand NAND2_2729 ( P1_U5425 , P1_U3021 , P1_U3063 );
nand NAND2_2730 ( P1_U5426 , P1_U3482 , P1_U5373 );
nand NAND2_2731 ( P1_U5427 , P1_U3021 , P1_U3062 );
nand NAND2_2732 ( P1_U5428 , P1_U3455 , P1_U5373 );
nand NAND2_2733 ( P1_U5429 , P1_U3021 , P1_U3078 );
nand NAND2_2734 ( P1_U5430 , P1_U3450 , P1_U5373 );
nand NAND2_2735 ( P1_U5431 , P1_U3021 , P1_U3077 );
nand NAND2_2736 ( P1_U5432 , P1_U4102 , P1_REG1_REG_0_ );
nand NAND2_2737 ( P1_U5433 , P1_U3021 , P1_U3479 );
nand NAND2_2738 ( P1_U5434 , P1_U3434 , P1_U3083 );
nand NAND2_2739 ( P1_U5435 , P1_U3021 , P1_U3476 );
nand NAND2_2740 ( P1_U5436 , P1_U3434 , P1_U3084 );
nand NAND2_2741 ( P1_U5437 , P1_U3021 , P1_U3473 );
nand NAND2_2742 ( P1_U5438 , P1_U3434 , P1_U3070 );
nand NAND2_2743 ( P1_U5439 , P1_U3021 , P1_U3470 );
nand NAND2_2744 ( P1_U5440 , P1_U3434 , P1_U3071 );
nand NAND2_2745 ( P1_U5441 , P1_U3021 , P1_U3467 );
nand NAND2_2746 ( P1_U5442 , P1_U3434 , P1_U3067 );
nand NAND2_2747 ( P1_U5443 , P1_U3021 , P1_U3464 );
nand NAND2_2748 ( P1_U5444 , P1_U3434 , P1_U3060 );
nand NAND2_2749 ( P1_U5445 , P1_U3021 , P1_U3461 );
nand NAND2_2750 ( P1_U5446 , P1_U3434 , P1_U3064 );
nand NAND2_2751 ( P1_U5447 , P1_U3021 , P1_U3974 );
nand NAND2_2752 ( P1_U5448 , P1_U3434 , P1_U3054 );
nand NAND2_2753 ( P1_U5449 , P1_U3021 , P1_U3975 );
nand NAND2_2754 ( P1_U5450 , P1_U3434 , P1_U3053 );
nand NAND2_2755 ( P1_U5451 , P1_U3021 , P1_U3976 );
nand NAND2_2756 ( P1_U5452 , P1_U3434 , P1_U3057 );
nand NAND2_2757 ( P1_U5453 , P1_U3021 , P1_U3977 );
nand NAND2_2758 ( P1_U5454 , P1_U3434 , P1_U3058 );
nand NAND2_2759 ( P1_U5455 , P1_U3021 , P1_U3978 );
nand NAND2_2760 ( P1_U5456 , P1_U3434 , P1_U3065 );
nand NAND2_2761 ( P1_U5457 , P1_U3021 , P1_U3979 );
nand NAND2_2762 ( P1_U5458 , P1_U3434 , P1_U3066 );
nand NAND2_2763 ( P1_U5459 , P1_U3021 , P1_U3980 );
nand NAND2_2764 ( P1_U5460 , P1_U3434 , P1_U3061 );
nand NAND2_2765 ( P1_U5461 , P1_U3021 , P1_U3981 );
nand NAND2_2766 ( P1_U5462 , P1_U3434 , P1_U3075 );
nand NAND2_2767 ( P1_U5463 , P1_U3021 , P1_U3982 );
nand NAND2_2768 ( P1_U5464 , P1_U3434 , P1_U3076 );
nand NAND2_2769 ( P1_U5465 , P1_U3021 , P1_U3458 );
nand NAND2_2770 ( P1_U5466 , P1_U3434 , P1_U3068 );
nand NAND2_2771 ( P1_U5467 , P1_U3021 , P1_U3508 );
nand NAND2_2772 ( P1_U5468 , P1_U3434 , P1_U3081 );
nand NAND2_2773 ( P1_U5469 , P1_U3021 , P1_U3506 );
nand NAND2_2774 ( P1_U5470 , P1_U3434 , P1_U3082 );
nand NAND2_2775 ( P1_U5471 , P1_U3021 , P1_U3503 );
nand NAND2_2776 ( P1_U5472 , P1_U3434 , P1_U3069 );
nand NAND2_2777 ( P1_U5473 , P1_U3021 , P1_U3500 );
nand NAND2_2778 ( P1_U5474 , P1_U3434 , P1_U3073 );
nand NAND2_2779 ( P1_U5475 , P1_U3021 , P1_U3497 );
nand NAND2_2780 ( P1_U5476 , P1_U3434 , P1_U3074 );
nand NAND2_2781 ( P1_U5477 , P1_U3021 , P1_U3494 );
nand NAND2_2782 ( P1_U5478 , P1_U3434 , P1_U3079 );
nand NAND2_2783 ( P1_U5479 , P1_U3021 , P1_U3491 );
nand NAND2_2784 ( P1_U5480 , P1_U3434 , P1_U3080 );
nand NAND2_2785 ( P1_U5481 , P1_U3021 , P1_U3488 );
nand NAND2_2786 ( P1_U5482 , P1_U3434 , P1_U3072 );
nand NAND2_2787 ( P1_U5483 , P1_U3021 , P1_U3485 );
nand NAND2_2788 ( P1_U5484 , P1_U3434 , P1_U3063 );
nand NAND2_2789 ( P1_U5485 , P1_U3021 , P1_U3482 );
nand NAND2_2790 ( P1_U5486 , P1_U3434 , P1_U3062 );
nand NAND2_2791 ( P1_U5487 , P1_U3021 , P1_U3455 );
nand NAND2_2792 ( P1_U5488 , P1_U3434 , P1_U3078 );
nand NAND2_2793 ( P1_U5489 , P1_U3021 , P1_U3450 );
nand NAND2_2794 ( P1_U5490 , P1_U3434 , P1_U3077 );
nand NAND2_2795 ( P1_U5491 , P1_U4102 , P1_U3448 );
nand NAND2_2796 ( P1_U5492 , P1_U3426 , P1_U3428 );
nand NAND2_2797 ( P1_U5493 , P1_U3953 , P1_U3479 );
nand NAND2_2798 ( P1_U5494 , P1_U3586 , P1_U5492 );
nand NAND2_2799 ( P1_U5495 , P1_U3953 , P1_U3476 );
nand NAND2_2800 ( P1_U5496 , P1_U3587 , P1_U5492 );
nand NAND2_2801 ( P1_U5497 , P1_U3953 , P1_U3473 );
nand NAND2_2802 ( P1_U5498 , P1_U3588 , P1_U5492 );
nand NAND2_2803 ( P1_U5499 , P1_U3953 , P1_U3470 );
nand NAND2_2804 ( P1_U5500 , P1_U3589 , P1_U5492 );
nand NAND2_2805 ( P1_U5501 , P1_U3953 , P1_U3467 );
nand NAND2_2806 ( P1_U5502 , P1_U3590 , P1_U5492 );
nand NAND2_2807 ( P1_U5503 , P1_U3953 , P1_U3464 );
nand NAND2_2808 ( P1_U5504 , P1_U3591 , P1_U5492 );
nand NAND2_2809 ( P1_U5505 , P1_U3593 , P1_U5492 );
nand NAND2_2810 ( P1_U5506 , P1_U3983 , P1_U3953 );
nand NAND2_2811 ( P1_U5507 , P1_U3594 , P1_U5492 );
nand NAND2_2812 ( P1_U5508 , P1_U3984 , P1_U3953 );
nand NAND2_2813 ( P1_U5509 , P1_U3953 , P1_U3461 );
nand NAND2_2814 ( P1_U5510 , P1_U3592 , P1_U5492 );
nand NAND2_2815 ( P1_U5511 , P1_U3596 , P1_U5492 );
nand NAND2_2816 ( P1_U5512 , P1_U3985 , P1_U3953 );
nand NAND2_2817 ( P1_U5513 , P1_U3597 , P1_U5492 );
nand NAND2_2818 ( P1_U5514 , P1_U3974 , P1_U3953 );
nand NAND2_2819 ( P1_U5515 , P1_U3598 , P1_U5492 );
nand NAND2_2820 ( P1_U5516 , P1_U3975 , P1_U3953 );
nand NAND2_2821 ( P1_U5517 , P1_U3599 , P1_U5492 );
nand NAND2_2822 ( P1_U5518 , P1_U3976 , P1_U3953 );
nand NAND2_2823 ( P1_U5519 , P1_U3600 , P1_U5492 );
nand NAND2_2824 ( P1_U5520 , P1_U3977 , P1_U3953 );
nand NAND2_2825 ( P1_U5521 , P1_U3601 , P1_U5492 );
nand NAND2_2826 ( P1_U5522 , P1_U3978 , P1_U3953 );
nand NAND2_2827 ( P1_U5523 , P1_U3602 , P1_U5492 );
nand NAND2_2828 ( P1_U5524 , P1_U3979 , P1_U3953 );
nand NAND2_2829 ( P1_U5525 , P1_U3603 , P1_U5492 );
nand NAND2_2830 ( P1_U5526 , P1_U3980 , P1_U3953 );
nand NAND2_2831 ( P1_U5527 , P1_U3604 , P1_U5492 );
nand NAND2_2832 ( P1_U5528 , P1_U3981 , P1_U3953 );
nand NAND2_2833 ( P1_U5529 , P1_U3605 , P1_U5492 );
nand NAND2_2834 ( P1_U5530 , P1_U3982 , P1_U3953 );
nand NAND2_2835 ( P1_U5531 , P1_U3953 , P1_U3458 );
nand NAND2_2836 ( P1_U5532 , P1_U3595 , P1_U5492 );
nand NAND2_2837 ( P1_U5533 , P1_U3953 , P1_U3508 );
nand NAND2_2838 ( P1_U5534 , P1_U3607 , P1_U5492 );
nand NAND2_2839 ( P1_U5535 , P1_U3953 , P1_U3506 );
nand NAND2_2840 ( P1_U5536 , P1_U3608 , P1_U5492 );
nand NAND2_2841 ( P1_U5537 , P1_U3953 , P1_U3503 );
nand NAND2_2842 ( P1_U5538 , P1_U3609 , P1_U5492 );
nand NAND2_2843 ( P1_U5539 , P1_U3953 , P1_U3500 );
nand NAND2_2844 ( P1_U5540 , P1_U3610 , P1_U5492 );
nand NAND2_2845 ( P1_U5541 , P1_U3953 , P1_U3497 );
nand NAND2_2846 ( P1_U5542 , P1_U3611 , P1_U5492 );
nand NAND2_2847 ( P1_U5543 , P1_U3953 , P1_U3494 );
nand NAND2_2848 ( P1_U5544 , P1_U3612 , P1_U5492 );
nand NAND2_2849 ( P1_U5545 , P1_U3953 , P1_U3491 );
nand NAND2_2850 ( P1_U5546 , P1_U3613 , P1_U5492 );
nand NAND2_2851 ( P1_U5547 , P1_U3953 , P1_U3488 );
nand NAND2_2852 ( P1_U5548 , P1_U3614 , P1_U5492 );
nand NAND2_2853 ( P1_U5549 , P1_U3953 , P1_U3485 );
nand NAND2_2854 ( P1_U5550 , P1_U3615 , P1_U5492 );
nand NAND2_2855 ( P1_U5551 , P1_U3953 , P1_U3482 );
nand NAND2_2856 ( P1_U5552 , P1_U3616 , P1_U5492 );
nand NAND2_2857 ( P1_U5553 , P1_U3953 , P1_U3455 );
nand NAND2_2858 ( P1_U5554 , P1_U3606 , P1_U5492 );
nand NAND2_2859 ( P1_U5555 , P1_U3953 , P1_U3450 );
nand NAND2_2860 ( P1_U5556 , P1_U3617 , P1_U5492 );
nand NAND2_2861 ( P1_U5557 , P1_U3479 , P1_U5492 );
nand NAND2_2862 ( P1_U5558 , P1_U3953 , P1_U3586 );
nand NAND2_2863 ( P1_U5559 , P1_U5677 , P1_U3084 );
nand NAND2_2864 ( P1_U5560 , P1_U3476 , P1_U5492 );
nand NAND2_2865 ( P1_U5561 , P1_U3953 , P1_U3587 );
nand NAND2_2866 ( P1_U5562 , P1_U5677 , P1_U3070 );
nand NAND2_2867 ( P1_U5563 , P1_U3473 , P1_U5492 );
nand NAND2_2868 ( P1_U5564 , P1_U3953 , P1_U3588 );
nand NAND2_2869 ( P1_U5565 , P1_U5677 , P1_U3071 );
nand NAND2_2870 ( P1_U5566 , P1_U3470 , P1_U5492 );
nand NAND2_2871 ( P1_U5567 , P1_U3953 , P1_U3589 );
nand NAND2_2872 ( P1_U5568 , P1_U5677 , P1_U3067 );
nand NAND2_2873 ( P1_U5569 , P1_U3467 , P1_U5492 );
nand NAND2_2874 ( P1_U5570 , P1_U3953 , P1_U3590 );
nand NAND2_2875 ( P1_U5571 , P1_U5677 , P1_U3060 );
nand NAND2_2876 ( P1_U5572 , P1_U3464 , P1_U5492 );
nand NAND2_2877 ( P1_U5573 , P1_U3953 , P1_U3591 );
nand NAND2_2878 ( P1_U5574 , P1_U5677 , P1_U3064 );
nand NAND2_2879 ( P1_U5575 , P1_U3983 , P1_U5492 );
nand NAND2_2880 ( P1_U5576 , P1_U3953 , P1_U3593 );
nand NAND2_2881 ( P1_U5577 , P1_U3984 , P1_U5492 );
nand NAND2_2882 ( P1_U5578 , P1_U3953 , P1_U3594 );
nand NAND2_2883 ( P1_U5579 , P1_U3461 , P1_U5492 );
nand NAND2_2884 ( P1_U5580 , P1_U3953 , P1_U3592 );
nand NAND2_2885 ( P1_U5581 , P1_U5677 , P1_U3068 );
nand NAND2_2886 ( P1_U5582 , P1_U3985 , P1_U5492 );
nand NAND2_2887 ( P1_U5583 , P1_U3953 , P1_U3596 );
nand NAND2_2888 ( P1_U5584 , P1_U5677 , P1_U3054 );
nand NAND2_2889 ( P1_U5585 , P1_U3974 , P1_U5492 );
nand NAND2_2890 ( P1_U5586 , P1_U3953 , P1_U3597 );
nand NAND2_2891 ( P1_U5587 , P1_U5677 , P1_U3053 );
nand NAND2_2892 ( P1_U5588 , P1_U3975 , P1_U5492 );
nand NAND2_2893 ( P1_U5589 , P1_U3953 , P1_U3598 );
nand NAND2_2894 ( P1_U5590 , P1_U5677 , P1_U3057 );
nand NAND2_2895 ( P1_U5591 , P1_U3976 , P1_U5492 );
nand NAND2_2896 ( P1_U5592 , P1_U3953 , P1_U3599 );
nand NAND2_2897 ( P1_U5593 , P1_U5677 , P1_U3058 );
nand NAND2_2898 ( P1_U5594 , P1_U3977 , P1_U5492 );
nand NAND2_2899 ( P1_U5595 , P1_U3953 , P1_U3600 );
nand NAND2_2900 ( P1_U5596 , P1_U5677 , P1_U3065 );
nand NAND2_2901 ( P1_U5597 , P1_U3978 , P1_U5492 );
nand NAND2_2902 ( P1_U5598 , P1_U3953 , P1_U3601 );
nand NAND2_2903 ( P1_U5599 , P1_U5677 , P1_U3066 );
nand NAND2_2904 ( P1_U5600 , P1_U3979 , P1_U5492 );
nand NAND2_2905 ( P1_U5601 , P1_U3953 , P1_U3602 );
nand NAND2_2906 ( P1_U5602 , P1_U5677 , P1_U3061 );
nand NAND2_2907 ( P1_U5603 , P1_U3980 , P1_U5492 );
nand NAND2_2908 ( P1_U5604 , P1_U3953 , P1_U3603 );
nand NAND2_2909 ( P1_U5605 , P1_U5677 , P1_U3075 );
nand NAND2_2910 ( P1_U5606 , P1_U3981 , P1_U5492 );
nand NAND2_2911 ( P1_U5607 , P1_U3953 , P1_U3604 );
nand NAND2_2912 ( P1_U5608 , P1_U5677 , P1_U3076 );
nand NAND2_2913 ( P1_U5609 , P1_U3982 , P1_U5492 );
nand NAND2_2914 ( P1_U5610 , P1_U3953 , P1_U3605 );
nand NAND2_2915 ( P1_U5611 , P1_U5677 , P1_U3081 );
nand NAND2_2916 ( P1_U5612 , P1_U3458 , P1_U5492 );
nand NAND2_2917 ( P1_U5613 , P1_U3953 , P1_U3595 );
nand NAND2_2918 ( P1_U5614 , P1_U5677 , P1_U3078 );
nand NAND2_2919 ( P1_U5615 , P1_U3508 , P1_U5492 );
nand NAND2_2920 ( P1_U5616 , P1_U3953 , P1_U3607 );
nand NAND2_2921 ( P1_U5617 , P1_U5677 , P1_U3082 );
nand NAND2_2922 ( P1_U5618 , P1_U3506 , P1_U5492 );
nand NAND2_2923 ( P1_U5619 , P1_U3953 , P1_U3608 );
nand NAND2_2924 ( P1_U5620 , P1_U5677 , P1_U3069 );
nand NAND2_2925 ( P1_U5621 , P1_U3503 , P1_U5492 );
nand NAND2_2926 ( P1_U5622 , P1_U3953 , P1_U3609 );
nand NAND2_2927 ( P1_U5623 , P1_U5677 , P1_U3073 );
nand NAND2_2928 ( P1_U5624 , P1_U3500 , P1_U5492 );
nand NAND2_2929 ( P1_U5625 , P1_U3953 , P1_U3610 );
nand NAND2_2930 ( P1_U5626 , P1_U5677 , P1_U3074 );
nand NAND2_2931 ( P1_U5627 , P1_U3497 , P1_U5492 );
nand NAND2_2932 ( P1_U5628 , P1_U3953 , P1_U3611 );
nand NAND2_2933 ( P1_U5629 , P1_U5677 , P1_U3079 );
nand NAND2_2934 ( P1_U5630 , P1_U3494 , P1_U5492 );
nand NAND2_2935 ( P1_U5631 , P1_U3953 , P1_U3612 );
nand NAND2_2936 ( P1_U5632 , P1_U5677 , P1_U3080 );
nand NAND2_2937 ( P1_U5633 , P1_U3491 , P1_U5492 );
nand NAND2_2938 ( P1_U5634 , P1_U3953 , P1_U3613 );
nand NAND2_2939 ( P1_U5635 , P1_U5677 , P1_U3072 );
nand NAND2_2940 ( P1_U5636 , P1_U3488 , P1_U5492 );
nand NAND2_2941 ( P1_U5637 , P1_U3953 , P1_U3614 );
nand NAND2_2942 ( P1_U5638 , P1_U5677 , P1_U3063 );
nand NAND2_2943 ( P1_U5639 , P1_U3485 , P1_U5492 );
nand NAND2_2944 ( P1_U5640 , P1_U3953 , P1_U3615 );
nand NAND2_2945 ( P1_U5641 , P1_U5677 , P1_U3062 );
nand NAND2_2946 ( P1_U5642 , P1_U3482 , P1_U5492 );
nand NAND2_2947 ( P1_U5643 , P1_U3953 , P1_U3616 );
nand NAND2_2948 ( P1_U5644 , P1_U5677 , P1_U3083 );
nand NAND2_2949 ( P1_U5645 , P1_U3455 , P1_U5492 );
nand NAND2_2950 ( P1_U5646 , P1_U3953 , P1_U3606 );
nand NAND2_2951 ( P1_U5647 , P1_U5677 , P1_U3077 );
nand NAND2_2952 ( P1_U5648 , P1_U3450 , P1_U5492 );
nand NAND2_2953 ( P1_U5649 , P1_U3953 , P1_U3617 );
nand NAND4_2954 ( P1_U5650 , P1_U5662 , P1_U3950 , P1_U3052 , P1_U3864 );
nand NAND2_2955 ( P1_U5651 , P1_U3086 , P1_U5091 );
nand NAND3_2956 ( P1_U5652 , P1_U5091 , P1_U5090 , P1_U3865 );
nand NAND2_2957 ( P1_U5653 , P1_U3997 , P1_U3430 );
nand NAND2_2958 ( P1_U5654 , P1_U3972 , P1_U3997 );
nand NAND2_2959 ( P1_U5655 , P1_U5653 , P1_U3995 );
nand NAND2_2960 ( P1_U5656 , P1_U5654 , P1_U3996 );
nand NAND2_2961 ( P1_U5657 , P1_R1207_U14 , P1_U3958 );
nand NAND2_2962 ( P1_U5658 , P1_R1192_U14 , P1_U3959 );
nand NAND2_2963 ( P1_U5659 , P1_R1150_U14 , P1_U3961 );
nand NAND2_2964 ( P1_U5660 , P1_R1117_U14 , P1_U3963 );
nand NAND2_2965 ( P1_U5661 , P1_U5666 , P1_U5672 );
nand NAND3_2966 ( P1_U5662 , P1_U6170 , P1_U6169 , P1_U5693 );
nand NAND2_2967 ( P1_U5663 , P1_U3442 , P1_U3438 );
nand NAND2_2968 ( P1_U5664 , P1_IR_REG_24_ , P1_U3910 );
nand NAND2_2969 ( P1_U5665 , P1_IR_REG_31_ , P1_SUB_84_U17 );
not NOT1_2970 ( P1_U5666 , P1_U3435 );
nand NAND2_2971 ( P1_U5667 , P1_IR_REG_25_ , P1_U3910 );
nand NAND2_2972 ( P1_U5668 , P1_IR_REG_31_ , P1_SUB_84_U170 );
not NOT1_2973 ( P1_U5669 , P1_U3436 );
nand NAND2_2974 ( P1_U5670 , P1_IR_REG_26_ , P1_U3910 );
nand NAND2_2975 ( P1_U5671 , P1_IR_REG_31_ , P1_SUB_84_U18 );
not NOT1_2976 ( P1_U5672 , P1_U3437 );
nand NAND2_2977 ( P1_U5673 , P1_U3050 , P1_U3359 );
nand NAND3_2978 ( P1_U5674 , P1_U4003 , P1_U5666 , P1_B_REG );
nand NAND2_2979 ( P1_U5675 , P1_IR_REG_23_ , P1_U3910 );
nand NAND2_2980 ( P1_U5676 , P1_IR_REG_31_ , P1_SUB_84_U16 );
not NOT1_2981 ( P1_U5677 , P1_U3438 );
nand NAND2_2982 ( P1_U5678 , P1_D_REG_0_ , P1_U3911 );
nand NAND2_2983 ( P1_U5679 , P1_U3992 , P1_U4103 );
nand NAND2_2984 ( P1_U5680 , P1_D_REG_1_ , P1_U3911 );
nand NAND2_2985 ( P1_U5681 , P1_U3992 , P1_U4104 );
nand NAND2_2986 ( P1_U5682 , P1_IR_REG_22_ , P1_U3910 );
nand NAND2_2987 ( P1_U5683 , P1_IR_REG_31_ , P1_SUB_84_U15 );
not NOT1_2988 ( P1_U5684 , P1_U3443 );
nand NAND2_2989 ( P1_U5685 , P1_IR_REG_19_ , P1_U3910 );
nand NAND2_2990 ( P1_U5686 , P1_IR_REG_31_ , P1_SUB_84_U13 );
not NOT1_2991 ( P1_U5687 , P1_U3442 );
nand NAND2_2992 ( P1_U5688 , P1_IR_REG_20_ , P1_U3910 );
nand NAND2_2993 ( P1_U5689 , P1_IR_REG_31_ , P1_SUB_84_U14 );
not NOT1_2994 ( P1_U5690 , P1_U3441 );
nand NAND2_2995 ( P1_U5691 , P1_IR_REG_21_ , P1_U3910 );
nand NAND2_2996 ( P1_U5692 , P1_IR_REG_31_ , P1_SUB_84_U173 );
not NOT1_2997 ( P1_U5693 , P1_U3447 );
nand NAND2_2998 ( P1_U5694 , P1_IR_REG_0_ , P1_U3910 );
nand NAND2_2999 ( P1_U5695 , P1_IR_REG_31_ , P1_IR_REG_0_ );
not NOT1_3000 ( P1_U5696 , P1_U3448 );
nand NAND2_3001 ( P1_U5697 , P1_IR_REG_28_ , P1_U3910 );
nand NAND2_3002 ( P1_U5698 , P1_IR_REG_31_ , P1_SUB_84_U19 );
not NOT1_3003 ( P1_U5699 , P1_U3446 );
nand NAND2_3004 ( P1_U5700 , P1_IR_REG_27_ , P1_U3910 );
nand NAND2_3005 ( P1_U5701 , P1_IR_REG_31_ , P1_SUB_84_U42 );
not NOT1_3006 ( P1_U5702 , P1_U3449 );
nand NAND2_3007 ( P1_U5703 , U88 , P1_U3912 );
nand NAND2_3008 ( P1_U5704 , P1_U3971 , P1_U3448 );
not NOT1_3009 ( P1_U5705 , P1_U3450 );
nand NAND2_3010 ( P1_U5706 , P1_IR_REG_30_ , P1_U3910 );
nand NAND2_3011 ( P1_U5707 , P1_IR_REG_31_ , P1_SUB_84_U165 );
not NOT1_3012 ( P1_U5708 , P1_U3444 );
nand NAND2_3013 ( P1_U5709 , P1_IR_REG_29_ , P1_U3910 );
nand NAND2_3014 ( P1_U5710 , P1_IR_REG_31_ , P1_SUB_84_U20 );
not NOT1_3015 ( P1_U5711 , P1_U3445 );
nand NAND2_3016 ( P1_U5712 , P1_U3443 , P1_U5693 );
nand NAND2_3017 ( P1_U5713 , P1_U5684 , P1_U4135 );
nand NAND2_3018 ( P1_U5714 , P1_D_REG_1_ , P1_U4101 );
nand NAND2_3019 ( P1_U5715 , P1_U4104 , P1_U3360 );
not NOT1_3020 ( P1_U5716 , P1_U3452 );
nand NAND2_3021 ( P1_U5717 , P1_U5661 , P1_U3360 );
nand NAND2_3022 ( P1_U5718 , P1_D_REG_0_ , P1_U4101 );
not NOT1_3023 ( P1_U5719 , P1_U3451 );
nand NAND2_3024 ( P1_U5720 , P1_REG0_REG_0_ , P1_U3913 );
nand NAND2_3025 ( P1_U5721 , P1_U3991 , P1_U4155 );
nand NAND2_3026 ( P1_U5722 , P1_IR_REG_1_ , P1_U3910 );
nand NAND2_3027 ( P1_U5723 , P1_IR_REG_31_ , P1_SUB_84_U40 );
nand NAND2_3028 ( P1_U5724 , U77 , P1_U3912 );
nand NAND2_3029 ( P1_U5725 , P1_U3454 , P1_U3971 );
not NOT1_3030 ( P1_U5726 , P1_U3455 );
nand NAND2_3031 ( P1_U5727 , P1_REG0_REG_1_ , P1_U3913 );
nand NAND2_3032 ( P1_U5728 , P1_U3991 , P1_U4179 );
nand NAND2_3033 ( P1_U5729 , P1_IR_REG_2_ , P1_U3910 );
nand NAND2_3034 ( P1_U5730 , P1_IR_REG_31_ , P1_SUB_84_U21 );
nand NAND2_3035 ( P1_U5731 , U66 , P1_U3912 );
nand NAND2_3036 ( P1_U5732 , P1_U3457 , P1_U3971 );
not NOT1_3037 ( P1_U5733 , P1_U3458 );
nand NAND2_3038 ( P1_U5734 , P1_REG0_REG_2_ , P1_U3913 );
nand NAND2_3039 ( P1_U5735 , P1_U3991 , P1_U4198 );
nand NAND2_3040 ( P1_U5736 , P1_IR_REG_3_ , P1_U3910 );
nand NAND2_3041 ( P1_U5737 , P1_IR_REG_31_ , P1_SUB_84_U22 );
nand NAND2_3042 ( P1_U5738 , U63 , P1_U3912 );
nand NAND2_3043 ( P1_U5739 , P1_U3460 , P1_U3971 );
not NOT1_3044 ( P1_U5740 , P1_U3461 );
nand NAND2_3045 ( P1_U5741 , P1_REG0_REG_3_ , P1_U3913 );
nand NAND2_3046 ( P1_U5742 , P1_U3991 , P1_U4217 );
nand NAND2_3047 ( P1_U5743 , P1_IR_REG_4_ , P1_U3910 );
nand NAND2_3048 ( P1_U5744 , P1_IR_REG_31_ , P1_SUB_84_U23 );
nand NAND2_3049 ( P1_U5745 , U62 , P1_U3912 );
nand NAND2_3050 ( P1_U5746 , P1_U3463 , P1_U3971 );
not NOT1_3051 ( P1_U5747 , P1_U3464 );
nand NAND2_3052 ( P1_U5748 , P1_REG0_REG_4_ , P1_U3913 );
nand NAND2_3053 ( P1_U5749 , P1_U3991 , P1_U4236 );
nand NAND2_3054 ( P1_U5750 , P1_IR_REG_5_ , P1_U3910 );
nand NAND2_3055 ( P1_U5751 , P1_IR_REG_31_ , P1_SUB_84_U162 );
nand NAND2_3056 ( P1_U5752 , U61 , P1_U3912 );
nand NAND2_3057 ( P1_U5753 , P1_U3466 , P1_U3971 );
not NOT1_3058 ( P1_U5754 , P1_U3467 );
nand NAND2_3059 ( P1_U5755 , P1_REG0_REG_5_ , P1_U3913 );
nand NAND2_3060 ( P1_U5756 , P1_U3991 , P1_U4255 );
nand NAND2_3061 ( P1_U5757 , P1_IR_REG_6_ , P1_U3910 );
nand NAND2_3062 ( P1_U5758 , P1_IR_REG_31_ , P1_SUB_84_U24 );
nand NAND2_3063 ( P1_U5759 , U60 , P1_U3912 );
nand NAND2_3064 ( P1_U5760 , P1_U3469 , P1_U3971 );
not NOT1_3065 ( P1_U5761 , P1_U3470 );
nand NAND2_3066 ( P1_U5762 , P1_REG0_REG_6_ , P1_U3913 );
nand NAND2_3067 ( P1_U5763 , P1_U3991 , P1_U4274 );
nand NAND2_3068 ( P1_U5764 , P1_IR_REG_7_ , P1_U3910 );
nand NAND2_3069 ( P1_U5765 , P1_IR_REG_31_ , P1_SUB_84_U25 );
nand NAND2_3070 ( P1_U5766 , U59 , P1_U3912 );
nand NAND2_3071 ( P1_U5767 , P1_U3472 , P1_U3971 );
not NOT1_3072 ( P1_U5768 , P1_U3473 );
nand NAND2_3073 ( P1_U5769 , P1_REG0_REG_7_ , P1_U3913 );
nand NAND2_3074 ( P1_U5770 , P1_U3991 , P1_U4293 );
nand NAND2_3075 ( P1_U5771 , P1_IR_REG_8_ , P1_U3910 );
nand NAND2_3076 ( P1_U5772 , P1_IR_REG_31_ , P1_SUB_84_U26 );
nand NAND2_3077 ( P1_U5773 , U58 , P1_U3912 );
nand NAND2_3078 ( P1_U5774 , P1_U3475 , P1_U3971 );
not NOT1_3079 ( P1_U5775 , P1_U3476 );
nand NAND2_3080 ( P1_U5776 , P1_REG0_REG_8_ , P1_U3913 );
nand NAND2_3081 ( P1_U5777 , P1_U3991 , P1_U4312 );
nand NAND2_3082 ( P1_U5778 , P1_IR_REG_9_ , P1_U3910 );
nand NAND2_3083 ( P1_U5779 , P1_IR_REG_31_ , P1_SUB_84_U160 );
nand NAND2_3084 ( P1_U5780 , U57 , P1_U3912 );
nand NAND2_3085 ( P1_U5781 , P1_U3478 , P1_U3971 );
not NOT1_3086 ( P1_U5782 , P1_U3479 );
nand NAND2_3087 ( P1_U5783 , P1_REG0_REG_9_ , P1_U3913 );
nand NAND2_3088 ( P1_U5784 , P1_U3991 , P1_U4331 );
nand NAND2_3089 ( P1_U5785 , P1_IR_REG_10_ , P1_U3910 );
nand NAND2_3090 ( P1_U5786 , P1_IR_REG_31_ , P1_SUB_84_U6 );
nand NAND2_3091 ( P1_U5787 , U87 , P1_U3912 );
nand NAND2_3092 ( P1_U5788 , P1_U3481 , P1_U3971 );
not NOT1_3093 ( P1_U5789 , P1_U3482 );
nand NAND2_3094 ( P1_U5790 , P1_REG0_REG_10_ , P1_U3913 );
nand NAND2_3095 ( P1_U5791 , P1_U3991 , P1_U4350 );
nand NAND2_3096 ( P1_U5792 , P1_IR_REG_11_ , P1_U3910 );
nand NAND2_3097 ( P1_U5793 , P1_IR_REG_31_ , P1_SUB_84_U7 );
nand NAND2_3098 ( P1_U5794 , U86 , P1_U3912 );
nand NAND2_3099 ( P1_U5795 , P1_U3484 , P1_U3971 );
not NOT1_3100 ( P1_U5796 , P1_U3485 );
nand NAND2_3101 ( P1_U5797 , P1_REG0_REG_11_ , P1_U3913 );
nand NAND2_3102 ( P1_U5798 , P1_U3991 , P1_U4369 );
nand NAND2_3103 ( P1_U5799 , P1_IR_REG_12_ , P1_U3910 );
nand NAND2_3104 ( P1_U5800 , P1_IR_REG_31_ , P1_SUB_84_U8 );
nand NAND2_3105 ( P1_U5801 , U85 , P1_U3912 );
nand NAND2_3106 ( P1_U5802 , P1_U3487 , P1_U3971 );
not NOT1_3107 ( P1_U5803 , P1_U3488 );
nand NAND2_3108 ( P1_U5804 , P1_REG0_REG_12_ , P1_U3913 );
nand NAND2_3109 ( P1_U5805 , P1_U3991 , P1_U4388 );
nand NAND2_3110 ( P1_U5806 , P1_IR_REG_13_ , P1_U3910 );
nand NAND2_3111 ( P1_U5807 , P1_IR_REG_31_ , P1_SUB_84_U179 );
nand NAND2_3112 ( P1_U5808 , U84 , P1_U3912 );
nand NAND2_3113 ( P1_U5809 , P1_U3490 , P1_U3971 );
not NOT1_3114 ( P1_U5810 , P1_U3491 );
nand NAND2_3115 ( P1_U5811 , P1_REG0_REG_13_ , P1_U3913 );
nand NAND2_3116 ( P1_U5812 , P1_U3991 , P1_U4407 );
nand NAND2_3117 ( P1_U5813 , P1_IR_REG_14_ , P1_U3910 );
nand NAND2_3118 ( P1_U5814 , P1_IR_REG_31_ , P1_SUB_84_U9 );
nand NAND2_3119 ( P1_U5815 , U83 , P1_U3912 );
nand NAND2_3120 ( P1_U5816 , P1_U3493 , P1_U3971 );
not NOT1_3121 ( P1_U5817 , P1_U3494 );
nand NAND2_3122 ( P1_U5818 , P1_REG0_REG_14_ , P1_U3913 );
nand NAND2_3123 ( P1_U5819 , P1_U3991 , P1_U4426 );
nand NAND2_3124 ( P1_U5820 , P1_IR_REG_15_ , P1_U3910 );
nand NAND2_3125 ( P1_U5821 , P1_IR_REG_31_ , P1_SUB_84_U10 );
nand NAND2_3126 ( P1_U5822 , U82 , P1_U3912 );
nand NAND2_3127 ( P1_U5823 , P1_U3496 , P1_U3971 );
not NOT1_3128 ( P1_U5824 , P1_U3497 );
nand NAND2_3129 ( P1_U5825 , P1_REG0_REG_15_ , P1_U3913 );
nand NAND2_3130 ( P1_U5826 , P1_U3991 , P1_U4445 );
nand NAND2_3131 ( P1_U5827 , P1_IR_REG_16_ , P1_U3910 );
nand NAND2_3132 ( P1_U5828 , P1_IR_REG_31_ , P1_SUB_84_U11 );
nand NAND2_3133 ( P1_U5829 , U81 , P1_U3912 );
nand NAND2_3134 ( P1_U5830 , P1_U3499 , P1_U3971 );
not NOT1_3135 ( P1_U5831 , P1_U3500 );
nand NAND2_3136 ( P1_U5832 , P1_REG0_REG_16_ , P1_U3913 );
nand NAND2_3137 ( P1_U5833 , P1_U3991 , P1_U4464 );
nand NAND2_3138 ( P1_U5834 , P1_IR_REG_17_ , P1_U3910 );
nand NAND2_3139 ( P1_U5835 , P1_IR_REG_31_ , P1_SUB_84_U177 );
nand NAND2_3140 ( P1_U5836 , U80 , P1_U3912 );
nand NAND2_3141 ( P1_U5837 , P1_U3502 , P1_U3971 );
not NOT1_3142 ( P1_U5838 , P1_U3503 );
nand NAND2_3143 ( P1_U5839 , P1_REG0_REG_17_ , P1_U3913 );
nand NAND2_3144 ( P1_U5840 , P1_U3991 , P1_U4483 );
nand NAND2_3145 ( P1_U5841 , P1_IR_REG_18_ , P1_U3910 );
nand NAND2_3146 ( P1_U5842 , P1_IR_REG_31_ , P1_SUB_84_U12 );
nand NAND2_3147 ( P1_U5843 , U79 , P1_U3912 );
nand NAND2_3148 ( P1_U5844 , P1_U3505 , P1_U3971 );
not NOT1_3149 ( P1_U5845 , P1_U3506 );
nand NAND2_3150 ( P1_U5846 , P1_REG0_REG_18_ , P1_U3913 );
nand NAND2_3151 ( P1_U5847 , P1_U3991 , P1_U4502 );
nand NAND2_3152 ( P1_U5848 , U78 , P1_U3912 );
nand NAND2_3153 ( P1_U5849 , P1_U3971 , P1_U3442 );
not NOT1_3154 ( P1_U5850 , P1_U3508 );
nand NAND2_3155 ( P1_U5851 , P1_REG0_REG_19_ , P1_U3913 );
nand NAND2_3156 ( P1_U5852 , P1_U3991 , P1_U4521 );
nand NAND2_3157 ( P1_U5853 , P1_REG0_REG_20_ , P1_U3913 );
nand NAND2_3158 ( P1_U5854 , P1_U3991 , P1_U4540 );
nand NAND2_3159 ( P1_U5855 , P1_REG0_REG_21_ , P1_U3913 );
nand NAND2_3160 ( P1_U5856 , P1_U3991 , P1_U4559 );
nand NAND2_3161 ( P1_U5857 , P1_REG0_REG_22_ , P1_U3913 );
nand NAND2_3162 ( P1_U5858 , P1_U3991 , P1_U4578 );
nand NAND2_3163 ( P1_U5859 , P1_REG0_REG_23_ , P1_U3913 );
nand NAND2_3164 ( P1_U5860 , P1_U3991 , P1_U4597 );
nand NAND2_3165 ( P1_U5861 , P1_REG0_REG_24_ , P1_U3913 );
nand NAND2_3166 ( P1_U5862 , P1_U3991 , P1_U4616 );
nand NAND2_3167 ( P1_U5863 , P1_REG0_REG_25_ , P1_U3913 );
nand NAND2_3168 ( P1_U5864 , P1_U3991 , P1_U4635 );
nand NAND2_3169 ( P1_U5865 , P1_REG0_REG_26_ , P1_U3913 );
nand NAND2_3170 ( P1_U5866 , P1_U3991 , P1_U4654 );
nand NAND2_3171 ( P1_U5867 , P1_REG0_REG_27_ , P1_U3913 );
nand NAND2_3172 ( P1_U5868 , P1_U3991 , P1_U4673 );
nand NAND2_3173 ( P1_U5869 , P1_REG0_REG_28_ , P1_U3913 );
nand NAND2_3174 ( P1_U5870 , P1_U3991 , P1_U4692 );
nand NAND2_3175 ( P1_U5871 , P1_REG0_REG_29_ , P1_U3913 );
nand NAND2_3176 ( P1_U5872 , P1_U3991 , P1_U4712 );
nand NAND2_3177 ( P1_U5873 , P1_REG0_REG_30_ , P1_U3913 );
nand NAND2_3178 ( P1_U5874 , P1_U3991 , P1_U4719 );
nand NAND2_3179 ( P1_U5875 , P1_REG0_REG_31_ , P1_U3913 );
nand NAND2_3180 ( P1_U5876 , P1_U3991 , P1_U4722 );
nand NAND2_3181 ( P1_U5877 , P1_REG1_REG_0_ , P1_U3914 );
nand NAND2_3182 ( P1_U5878 , P1_U3990 , P1_U4155 );
nand NAND2_3183 ( P1_U5879 , P1_REG1_REG_1_ , P1_U3914 );
nand NAND2_3184 ( P1_U5880 , P1_U3990 , P1_U4179 );
nand NAND2_3185 ( P1_U5881 , P1_REG1_REG_2_ , P1_U3914 );
nand NAND2_3186 ( P1_U5882 , P1_U3990 , P1_U4198 );
nand NAND2_3187 ( P1_U5883 , P1_REG1_REG_3_ , P1_U3914 );
nand NAND2_3188 ( P1_U5884 , P1_U3990 , P1_U4217 );
nand NAND2_3189 ( P1_U5885 , P1_REG1_REG_4_ , P1_U3914 );
nand NAND2_3190 ( P1_U5886 , P1_U3990 , P1_U4236 );
nand NAND2_3191 ( P1_U5887 , P1_REG1_REG_5_ , P1_U3914 );
nand NAND2_3192 ( P1_U5888 , P1_U3990 , P1_U4255 );
nand NAND2_3193 ( P1_U5889 , P1_REG1_REG_6_ , P1_U3914 );
nand NAND2_3194 ( P1_U5890 , P1_U3990 , P1_U4274 );
nand NAND2_3195 ( P1_U5891 , P1_REG1_REG_7_ , P1_U3914 );
nand NAND2_3196 ( P1_U5892 , P1_U3990 , P1_U4293 );
nand NAND2_3197 ( P1_U5893 , P1_REG1_REG_8_ , P1_U3914 );
nand NAND2_3198 ( P1_U5894 , P1_U3990 , P1_U4312 );
nand NAND2_3199 ( P1_U5895 , P1_REG1_REG_9_ , P1_U3914 );
nand NAND2_3200 ( P1_U5896 , P1_U3990 , P1_U4331 );
nand NAND2_3201 ( P1_U5897 , P1_REG1_REG_10_ , P1_U3914 );
nand NAND2_3202 ( P1_U5898 , P1_U3990 , P1_U4350 );
nand NAND2_3203 ( P1_U5899 , P1_REG1_REG_11_ , P1_U3914 );
nand NAND2_3204 ( P1_U5900 , P1_U3990 , P1_U4369 );
nand NAND2_3205 ( P1_U5901 , P1_REG1_REG_12_ , P1_U3914 );
nand NAND2_3206 ( P1_U5902 , P1_U3990 , P1_U4388 );
nand NAND2_3207 ( P1_U5903 , P1_REG1_REG_13_ , P1_U3914 );
nand NAND2_3208 ( P1_U5904 , P1_U3990 , P1_U4407 );
nand NAND2_3209 ( P1_U5905 , P1_REG1_REG_14_ , P1_U3914 );
nand NAND2_3210 ( P1_U5906 , P1_U3990 , P1_U4426 );
nand NAND2_3211 ( P1_U5907 , P1_REG1_REG_15_ , P1_U3914 );
nand NAND2_3212 ( P1_U5908 , P1_U3990 , P1_U4445 );
nand NAND2_3213 ( P1_U5909 , P1_REG1_REG_16_ , P1_U3914 );
nand NAND2_3214 ( P1_U5910 , P1_U3990 , P1_U4464 );
nand NAND2_3215 ( P1_U5911 , P1_REG1_REG_17_ , P1_U3914 );
nand NAND2_3216 ( P1_U5912 , P1_U3990 , P1_U4483 );
nand NAND2_3217 ( P1_U5913 , P1_REG1_REG_18_ , P1_U3914 );
nand NAND2_3218 ( P1_U5914 , P1_U3990 , P1_U4502 );
nand NAND2_3219 ( P1_U5915 , P1_REG1_REG_19_ , P1_U3914 );
nand NAND2_3220 ( P1_U5916 , P1_U3990 , P1_U4521 );
nand NAND2_3221 ( P1_U5917 , P1_REG1_REG_20_ , P1_U3914 );
nand NAND2_3222 ( P1_U5918 , P1_U3990 , P1_U4540 );
nand NAND2_3223 ( P1_U5919 , P1_REG1_REG_21_ , P1_U3914 );
nand NAND2_3224 ( P1_U5920 , P1_U3990 , P1_U4559 );
nand NAND2_3225 ( P1_U5921 , P1_REG1_REG_22_ , P1_U3914 );
nand NAND2_3226 ( P1_U5922 , P1_U3990 , P1_U4578 );
nand NAND2_3227 ( P1_U5923 , P1_REG1_REG_23_ , P1_U3914 );
nand NAND2_3228 ( P1_U5924 , P1_U3990 , P1_U4597 );
nand NAND2_3229 ( P1_U5925 , P1_REG1_REG_24_ , P1_U3914 );
nand NAND2_3230 ( P1_U5926 , P1_U3990 , P1_U4616 );
nand NAND2_3231 ( P1_U5927 , P1_REG1_REG_25_ , P1_U3914 );
nand NAND2_3232 ( P1_U5928 , P1_U3990 , P1_U4635 );
nand NAND2_3233 ( P1_U5929 , P1_REG1_REG_26_ , P1_U3914 );
nand NAND2_3234 ( P1_U5930 , P1_U3990 , P1_U4654 );
nand NAND2_3235 ( P1_U5931 , P1_REG1_REG_27_ , P1_U3914 );
nand NAND2_3236 ( P1_U5932 , P1_U3990 , P1_U4673 );
nand NAND2_3237 ( P1_U5933 , P1_REG1_REG_28_ , P1_U3914 );
nand NAND2_3238 ( P1_U5934 , P1_U3990 , P1_U4692 );
nand NAND2_3239 ( P1_U5935 , P1_REG1_REG_29_ , P1_U3914 );
nand NAND2_3240 ( P1_U5936 , P1_U3990 , P1_U4712 );
nand NAND2_3241 ( P1_U5937 , P1_REG1_REG_30_ , P1_U3914 );
nand NAND2_3242 ( P1_U5938 , P1_U3990 , P1_U4719 );
nand NAND2_3243 ( P1_U5939 , P1_REG1_REG_31_ , P1_U3914 );
nand NAND2_3244 ( P1_U5940 , P1_U3990 , P1_U4722 );
nand NAND2_3245 ( P1_U5941 , P1_REG2_REG_0_ , P1_U3417 );
nand NAND2_3246 ( P1_U5942 , P1_U3989 , P1_U3374 );
nand NAND2_3247 ( P1_U5943 , P1_REG2_REG_1_ , P1_U3417 );
nand NAND2_3248 ( P1_U5944 , P1_U3989 , P1_U3376 );
nand NAND2_3249 ( P1_U5945 , P1_REG2_REG_2_ , P1_U3417 );
nand NAND2_3250 ( P1_U5946 , P1_U3989 , P1_U3377 );
nand NAND2_3251 ( P1_U5947 , P1_REG2_REG_3_ , P1_U3417 );
nand NAND2_3252 ( P1_U5948 , P1_U3989 , P1_U3378 );
nand NAND2_3253 ( P1_U5949 , P1_REG2_REG_4_ , P1_U3417 );
nand NAND2_3254 ( P1_U5950 , P1_U3989 , P1_U3379 );
nand NAND2_3255 ( P1_U5951 , P1_REG2_REG_5_ , P1_U3417 );
nand NAND2_3256 ( P1_U5952 , P1_U3989 , P1_U3380 );
nand NAND2_3257 ( P1_U5953 , P1_REG2_REG_6_ , P1_U3417 );
nand NAND2_3258 ( P1_U5954 , P1_U3989 , P1_U3381 );
nand NAND2_3259 ( P1_U5955 , P1_REG2_REG_7_ , P1_U3417 );
nand NAND2_3260 ( P1_U5956 , P1_U3989 , P1_U3382 );
nand NAND2_3261 ( P1_U5957 , P1_REG2_REG_8_ , P1_U3417 );
nand NAND2_3262 ( P1_U5958 , P1_U3989 , P1_U3383 );
nand NAND2_3263 ( P1_U5959 , P1_REG2_REG_9_ , P1_U3417 );
nand NAND2_3264 ( P1_U5960 , P1_U3989 , P1_U3384 );
nand NAND2_3265 ( P1_U5961 , P1_REG2_REG_10_ , P1_U3417 );
nand NAND2_3266 ( P1_U5962 , P1_U3989 , P1_U3385 );
nand NAND2_3267 ( P1_U5963 , P1_REG2_REG_11_ , P1_U3417 );
nand NAND2_3268 ( P1_U5964 , P1_U3989 , P1_U3386 );
nand NAND2_3269 ( P1_U5965 , P1_REG2_REG_12_ , P1_U3417 );
nand NAND2_3270 ( P1_U5966 , P1_U3989 , P1_U3387 );
nand NAND2_3271 ( P1_U5967 , P1_REG2_REG_13_ , P1_U3417 );
nand NAND2_3272 ( P1_U5968 , P1_U3989 , P1_U3388 );
nand NAND2_3273 ( P1_U5969 , P1_REG2_REG_14_ , P1_U3417 );
nand NAND2_3274 ( P1_U5970 , P1_U3989 , P1_U3389 );
nand NAND2_3275 ( P1_U5971 , P1_REG2_REG_15_ , P1_U3417 );
nand NAND2_3276 ( P1_U5972 , P1_U3989 , P1_U3390 );
nand NAND2_3277 ( P1_U5973 , P1_REG2_REG_16_ , P1_U3417 );
nand NAND2_3278 ( P1_U5974 , P1_U3989 , P1_U3391 );
nand NAND2_3279 ( P1_U5975 , P1_REG2_REG_17_ , P1_U3417 );
nand NAND2_3280 ( P1_U5976 , P1_U3989 , P1_U3392 );
nand NAND2_3281 ( P1_U5977 , P1_REG2_REG_18_ , P1_U3417 );
nand NAND2_3282 ( P1_U5978 , P1_U3989 , P1_U3393 );
nand NAND2_3283 ( P1_U5979 , P1_REG2_REG_19_ , P1_U3417 );
nand NAND2_3284 ( P1_U5980 , P1_U3989 , P1_U3394 );
nand NAND2_3285 ( P1_U5981 , P1_REG2_REG_20_ , P1_U3417 );
nand NAND2_3286 ( P1_U5982 , P1_U3989 , P1_U3396 );
nand NAND2_3287 ( P1_U5983 , P1_REG2_REG_21_ , P1_U3417 );
nand NAND2_3288 ( P1_U5984 , P1_U3989 , P1_U3398 );
nand NAND2_3289 ( P1_U5985 , P1_REG2_REG_22_ , P1_U3417 );
nand NAND2_3290 ( P1_U5986 , P1_U3989 , P1_U3400 );
nand NAND2_3291 ( P1_U5987 , P1_REG2_REG_23_ , P1_U3417 );
nand NAND2_3292 ( P1_U5988 , P1_U3989 , P1_U3402 );
nand NAND2_3293 ( P1_U5989 , P1_REG2_REG_24_ , P1_U3417 );
nand NAND2_3294 ( P1_U5990 , P1_U3989 , P1_U3404 );
nand NAND2_3295 ( P1_U5991 , P1_REG2_REG_25_ , P1_U3417 );
nand NAND2_3296 ( P1_U5992 , P1_U3989 , P1_U3406 );
nand NAND2_3297 ( P1_U5993 , P1_REG2_REG_26_ , P1_U3417 );
nand NAND2_3298 ( P1_U5994 , P1_U3989 , P1_U3408 );
nand NAND2_3299 ( P1_U5995 , P1_REG2_REG_27_ , P1_U3417 );
nand NAND2_3300 ( P1_U5996 , P1_U3989 , P1_U3410 );
nand NAND2_3301 ( P1_U5997 , P1_REG2_REG_28_ , P1_U3417 );
nand NAND2_3302 ( P1_U5998 , P1_U3989 , P1_U3412 );
nand NAND2_3303 ( P1_U5999 , P1_REG2_REG_29_ , P1_U3417 );
nand NAND2_3304 ( P1_U6000 , P1_U3989 , P1_U4708 );
nand NAND2_3305 ( P1_U6001 , P1_REG2_REG_30_ , P1_U3417 );
nand NAND2_3306 ( P1_U6002 , P1_U3993 , P1_U3989 );
nand NAND2_3307 ( P1_U6003 , P1_REG2_REG_31_ , P1_U3417 );
nand NAND2_3308 ( P1_U6004 , P1_U3993 , P1_U3989 );
nand NAND2_3309 ( P1_U6005 , P1_DATAO_REG_0_ , P1_U3425 );
nand NAND2_3310 ( P1_U6006 , P1_U3973 , P1_U3077 );
nand NAND2_3311 ( P1_U6007 , P1_DATAO_REG_1_ , P1_U3425 );
nand NAND2_3312 ( P1_U6008 , P1_U3973 , P1_U3078 );
nand NAND2_3313 ( P1_U6009 , P1_DATAO_REG_2_ , P1_U3425 );
nand NAND2_3314 ( P1_U6010 , P1_U3973 , P1_U3068 );
nand NAND2_3315 ( P1_U6011 , P1_DATAO_REG_3_ , P1_U3425 );
nand NAND2_3316 ( P1_U6012 , P1_U3973 , P1_U3064 );
nand NAND2_3317 ( P1_U6013 , P1_DATAO_REG_4_ , P1_U3425 );
nand NAND2_3318 ( P1_U6014 , P1_U3973 , P1_U3060 );
nand NAND2_3319 ( P1_U6015 , P1_DATAO_REG_5_ , P1_U3425 );
nand NAND2_3320 ( P1_U6016 , P1_U3973 , P1_U3067 );
nand NAND2_3321 ( P1_U6017 , P1_DATAO_REG_6_ , P1_U3425 );
nand NAND2_3322 ( P1_U6018 , P1_U3973 , P1_U3071 );
nand NAND2_3323 ( P1_U6019 , P1_DATAO_REG_7_ , P1_U3425 );
nand NAND2_3324 ( P1_U6020 , P1_U3973 , P1_U3070 );
nand NAND2_3325 ( P1_U6021 , P1_DATAO_REG_8_ , P1_U3425 );
nand NAND2_3326 ( P1_U6022 , P1_U3973 , P1_U3084 );
nand NAND2_3327 ( P1_U6023 , P1_DATAO_REG_9_ , P1_U3425 );
nand NAND2_3328 ( P1_U6024 , P1_U3973 , P1_U3083 );
nand NAND2_3329 ( P1_U6025 , P1_DATAO_REG_10_ , P1_U3425 );
nand NAND2_3330 ( P1_U6026 , P1_U3973 , P1_U3062 );
nand NAND2_3331 ( P1_U6027 , P1_DATAO_REG_11_ , P1_U3425 );
nand NAND2_3332 ( P1_U6028 , P1_U3973 , P1_U3063 );
nand NAND2_3333 ( P1_U6029 , P1_DATAO_REG_12_ , P1_U3425 );
nand NAND2_3334 ( P1_U6030 , P1_U3973 , P1_U3072 );
nand NAND2_3335 ( P1_U6031 , P1_DATAO_REG_13_ , P1_U3425 );
nand NAND2_3336 ( P1_U6032 , P1_U3973 , P1_U3080 );
nand NAND2_3337 ( P1_U6033 , P1_DATAO_REG_14_ , P1_U3425 );
nand NAND2_3338 ( P1_U6034 , P1_U3973 , P1_U3079 );
nand NAND2_3339 ( P1_U6035 , P1_DATAO_REG_15_ , P1_U3425 );
nand NAND2_3340 ( P1_U6036 , P1_U3973 , P1_U3074 );
nand NAND2_3341 ( P1_U6037 , P1_DATAO_REG_16_ , P1_U3425 );
nand NAND2_3342 ( P1_U6038 , P1_U3973 , P1_U3073 );
nand NAND2_3343 ( P1_U6039 , P1_DATAO_REG_17_ , P1_U3425 );
nand NAND2_3344 ( P1_U6040 , P1_U3973 , P1_U3069 );
nand NAND2_3345 ( P1_U6041 , P1_DATAO_REG_18_ , P1_U3425 );
nand NAND2_3346 ( P1_U6042 , P1_U3973 , P1_U3082 );
nand NAND2_3347 ( P1_U6043 , P1_DATAO_REG_19_ , P1_U3425 );
nand NAND2_3348 ( P1_U6044 , P1_U3973 , P1_U3081 );
nand NAND2_3349 ( P1_U6045 , P1_DATAO_REG_20_ , P1_U3425 );
nand NAND2_3350 ( P1_U6046 , P1_U3973 , P1_U3076 );
nand NAND2_3351 ( P1_U6047 , P1_DATAO_REG_21_ , P1_U3425 );
nand NAND2_3352 ( P1_U6048 , P1_U3973 , P1_U3075 );
nand NAND2_3353 ( P1_U6049 , P1_DATAO_REG_22_ , P1_U3425 );
nand NAND2_3354 ( P1_U6050 , P1_U3973 , P1_U3061 );
nand NAND2_3355 ( P1_U6051 , P1_DATAO_REG_23_ , P1_U3425 );
nand NAND2_3356 ( P1_U6052 , P1_U3973 , P1_U3066 );
nand NAND2_3357 ( P1_U6053 , P1_DATAO_REG_24_ , P1_U3425 );
nand NAND2_3358 ( P1_U6054 , P1_U3973 , P1_U3065 );
nand NAND2_3359 ( P1_U6055 , P1_DATAO_REG_25_ , P1_U3425 );
nand NAND2_3360 ( P1_U6056 , P1_U3973 , P1_U3058 );
nand NAND2_3361 ( P1_U6057 , P1_DATAO_REG_26_ , P1_U3425 );
nand NAND2_3362 ( P1_U6058 , P1_U3973 , P1_U3057 );
nand NAND2_3363 ( P1_U6059 , P1_DATAO_REG_27_ , P1_U3425 );
nand NAND2_3364 ( P1_U6060 , P1_U3973 , P1_U3053 );
nand NAND2_3365 ( P1_U6061 , P1_DATAO_REG_28_ , P1_U3425 );
nand NAND2_3366 ( P1_U6062 , P1_U3973 , P1_U3054 );
nand NAND2_3367 ( P1_U6063 , P1_DATAO_REG_29_ , P1_U3425 );
nand NAND2_3368 ( P1_U6064 , P1_U3973 , P1_U3055 );
nand NAND2_3369 ( P1_U6065 , P1_DATAO_REG_30_ , P1_U3425 );
nand NAND2_3370 ( P1_U6066 , P1_U3973 , P1_U3059 );
nand NAND2_3371 ( P1_U6067 , P1_DATAO_REG_31_ , P1_U3425 );
nand NAND2_3372 ( P1_U6068 , P1_U3973 , P1_U3056 );
nand NAND3_3373 ( P1_U6069 , P1_U3048 , P1_U3438 , P1_U3948 );
nand NAND3_3374 ( P1_U6070 , P1_U3954 , P1_U5690 , P1_R1375_U14 );
nand NAND4_3375 ( P1_U6071 , P1_U5684 , P1_U3447 , P1_U3438 , P1_U3949 );
nand NAND3_3376 ( P1_U6072 , P1_U3955 , P1_U3959 , P1_R1360_U14 );
nand NAND2_3377 ( P1_U6073 , P1_U3985 , P1_U3055 );
nand NAND2_3378 ( P1_U6074 , P1_U3413 , P1_U4678 );
nand NAND2_3379 ( P1_U6075 , P1_U6074 , P1_U6073 );
nand NAND2_3380 ( P1_U6076 , P1_U3974 , P1_U3054 );
nand NAND2_3381 ( P1_U6077 , P1_U3411 , P1_U4659 );
nand NAND2_3382 ( P1_U6078 , P1_U6077 , P1_U6076 );
nand NAND2_3383 ( P1_U6079 , P1_U3975 , P1_U3053 );
nand NAND2_3384 ( P1_U6080 , P1_U3409 , P1_U4640 );
nand NAND2_3385 ( P1_U6081 , P1_U6080 , P1_U6079 );
nand NAND2_3386 ( P1_U6082 , P1_U3978 , P1_U3065 );
nand NAND2_3387 ( P1_U6083 , P1_U3403 , P1_U4583 );
nand NAND2_3388 ( P1_U6084 , P1_U6083 , P1_U6082 );
nand NAND2_3389 ( P1_U6085 , P1_U3979 , P1_U3066 );
nand NAND2_3390 ( P1_U6086 , P1_U3401 , P1_U4564 );
nand NAND2_3391 ( P1_U6087 , P1_U6086 , P1_U6085 );
nand NAND2_3392 ( P1_U6088 , P1_U3981 , P1_U3075 );
nand NAND2_3393 ( P1_U6089 , P1_U3397 , P1_U4526 );
nand NAND2_3394 ( P1_U6090 , P1_U6089 , P1_U6088 );
nand NAND2_3395 ( P1_U6091 , P1_U3980 , P1_U3061 );
nand NAND2_3396 ( P1_U6092 , P1_U3399 , P1_U4545 );
nand NAND2_3397 ( P1_U6093 , P1_U6092 , P1_U6091 );
nand NAND2_3398 ( P1_U6094 , P1_U3977 , P1_U3058 );
nand NAND2_3399 ( P1_U6095 , P1_U3405 , P1_U4602 );
nand NAND2_3400 ( P1_U6096 , P1_U6095 , P1_U6094 );
nand NAND2_3401 ( P1_U6097 , P1_U3976 , P1_U3057 );
nand NAND2_3402 ( P1_U6098 , P1_U3407 , P1_U4621 );
nand NAND2_3403 ( P1_U6099 , P1_U6098 , P1_U6097 );
nand NAND2_3404 ( P1_U6100 , P1_U3984 , P1_U3059 );
nand NAND2_3405 ( P1_U6101 , P1_U3414 , P1_U4696 );
nand NAND2_3406 ( P1_U6102 , P1_U6101 , P1_U6100 );
nand NAND2_3407 ( P1_U6103 , P1_U3983 , P1_U3056 );
nand NAND2_3408 ( P1_U6104 , P1_U3415 , P1_U4716 );
nand NAND2_3409 ( P1_U6105 , P1_U6104 , P1_U6103 );
nand NAND2_3410 ( P1_U6106 , P1_U5838 , P1_U4450 );
nand NAND2_3411 ( P1_U6107 , P1_U3503 , P1_U3069 );
nand NAND2_3412 ( P1_U6108 , P1_U6107 , P1_U6106 );
nand NAND2_3413 ( P1_U6109 , P1_U5775 , P1_U4279 );
nand NAND2_3414 ( P1_U6110 , P1_U3476 , P1_U3084 );
nand NAND2_3415 ( P1_U6111 , P1_U6110 , P1_U6109 );
nand NAND2_3416 ( P1_U6112 , P1_U5782 , P1_U4298 );
nand NAND2_3417 ( P1_U6113 , P1_U3479 , P1_U3083 );
nand NAND2_3418 ( P1_U6114 , P1_U6113 , P1_U6112 );
nand NAND2_3419 ( P1_U6115 , P1_U5810 , P1_U4374 );
nand NAND2_3420 ( P1_U6116 , P1_U3491 , P1_U3080 );
nand NAND2_3421 ( P1_U6117 , P1_U6116 , P1_U6115 );
nand NAND2_3422 ( P1_U6118 , P1_U5817 , P1_U4393 );
nand NAND2_3423 ( P1_U6119 , P1_U3494 , P1_U3079 );
nand NAND2_3424 ( P1_U6120 , P1_U6119 , P1_U6118 );
nand NAND2_3425 ( P1_U6121 , P1_U5705 , P1_U4165 );
nand NAND2_3426 ( P1_U6122 , P1_U3450 , P1_U3077 );
nand NAND2_3427 ( P1_U6123 , P1_U6122 , P1_U6121 );
nand NAND2_3428 ( P1_U6124 , P1_U5726 , P1_U4141 );
nand NAND2_3429 ( P1_U6125 , P1_U3455 , P1_U3078 );
nand NAND2_3430 ( P1_U6126 , P1_U6125 , P1_U6124 );
nand NAND2_3431 ( P1_U6127 , P1_U5824 , P1_U4412 );
nand NAND2_3432 ( P1_U6128 , P1_U3497 , P1_U3074 );
nand NAND2_3433 ( P1_U6129 , P1_U6128 , P1_U6127 );
nand NAND2_3434 ( P1_U6130 , P1_U5831 , P1_U4431 );
nand NAND2_3435 ( P1_U6131 , P1_U3500 , P1_U3073 );
nand NAND2_3436 ( P1_U6132 , P1_U6131 , P1_U6130 );
nand NAND2_3437 ( P1_U6133 , P1_U5761 , P1_U4241 );
nand NAND2_3438 ( P1_U6134 , P1_U3470 , P1_U3071 );
nand NAND2_3439 ( P1_U6135 , P1_U6134 , P1_U6133 );
nand NAND2_3440 ( P1_U6136 , P1_U5768 , P1_U4260 );
nand NAND2_3441 ( P1_U6137 , P1_U3473 , P1_U3070 );
nand NAND2_3442 ( P1_U6138 , P1_U6137 , P1_U6136 );
nand NAND2_3443 ( P1_U6139 , P1_U5803 , P1_U4355 );
nand NAND2_3444 ( P1_U6140 , P1_U3488 , P1_U3072 );
nand NAND2_3445 ( P1_U6141 , P1_U6140 , P1_U6139 );
nand NAND2_3446 ( P1_U6142 , P1_U5733 , P1_U4160 );
nand NAND2_3447 ( P1_U6143 , P1_U3458 , P1_U3068 );
nand NAND2_3448 ( P1_U6144 , P1_U6143 , P1_U6142 );
nand NAND2_3449 ( P1_U6145 , P1_U5740 , P1_U4184 );
nand NAND2_3450 ( P1_U6146 , P1_U3461 , P1_U3064 );
nand NAND2_3451 ( P1_U6147 , P1_U6146 , P1_U6145 );
nand NAND2_3452 ( P1_U6148 , P1_U5754 , P1_U4222 );
nand NAND2_3453 ( P1_U6149 , P1_U3467 , P1_U3067 );
nand NAND2_3454 ( P1_U6150 , P1_U6149 , P1_U6148 );
nand NAND2_3455 ( P1_U6151 , P1_U5845 , P1_U4469 );
nand NAND2_3456 ( P1_U6152 , P1_U3506 , P1_U3082 );
nand NAND2_3457 ( P1_U6153 , P1_U6152 , P1_U6151 );
nand NAND2_3458 ( P1_U6154 , P1_U5850 , P1_U4488 );
nand NAND2_3459 ( P1_U6155 , P1_U3508 , P1_U3081 );
nand NAND2_3460 ( P1_U6156 , P1_U6155 , P1_U6154 );
nand NAND2_3461 ( P1_U6157 , P1_U5747 , P1_U4203 );
nand NAND2_3462 ( P1_U6158 , P1_U3464 , P1_U3060 );
nand NAND2_3463 ( P1_U6159 , P1_U6158 , P1_U6157 );
nand NAND2_3464 ( P1_U6160 , P1_U5796 , P1_U4336 );
nand NAND2_3465 ( P1_U6161 , P1_U3485 , P1_U3063 );
nand NAND2_3466 ( P1_U6162 , P1_U6161 , P1_U6160 );
nand NAND2_3467 ( P1_U6163 , P1_U5789 , P1_U4317 );
nand NAND2_3468 ( P1_U6164 , P1_U3482 , P1_U3062 );
nand NAND2_3469 ( P1_U6165 , P1_U6164 , P1_U6163 );
nand NAND2_3470 ( P1_U6166 , P1_U3982 , P1_U3076 );
nand NAND2_3471 ( P1_U6167 , P1_U3395 , P1_U4507 );
nand NAND2_3472 ( P1_U6168 , P1_U6167 , P1_U6166 );
nand NAND2_3473 ( P1_U6169 , P1_U5663 , P1_U3951 );
nand NAND2_3474 ( P1_U6170 , P1_U5086 , P1_U3426 );
nand NAND2_3475 ( P1_U6171 , P1_U3083 , P1_R1352_U6 );
nand NAND2_3476 ( P1_U6172 , P1_U3083 , P1_U3952 );
nand NAND2_3477 ( P1_U6173 , P1_U3084 , P1_R1352_U6 );
nand NAND2_3478 ( P1_U6174 , P1_U3084 , P1_U3952 );
nand NAND2_3479 ( P1_U6175 , P1_U3070 , P1_R1352_U6 );
nand NAND2_3480 ( P1_U6176 , P1_U3070 , P1_U3952 );
nand NAND2_3481 ( P1_U6177 , P1_U3071 , P1_R1352_U6 );
nand NAND2_3482 ( P1_U6178 , P1_U3071 , P1_U3952 );
nand NAND2_3483 ( P1_U6179 , P1_U3067 , P1_R1352_U6 );
nand NAND2_3484 ( P1_U6180 , P1_U3067 , P1_U3952 );
nand NAND2_3485 ( P1_U6181 , P1_U3060 , P1_R1352_U6 );
nand NAND2_3486 ( P1_U6182 , P1_U3060 , P1_U3952 );
nand NAND2_3487 ( P1_U6183 , P1_U3064 , P1_R1352_U6 );
nand NAND2_3488 ( P1_U6184 , P1_U3064 , P1_U3952 );
nand NAND2_3489 ( P1_U6185 , P1_R1309_U8 , P1_R1352_U6 );
nand NAND2_3490 ( P1_U6186 , P1_U3056 , P1_U3952 );
nand NAND2_3491 ( P1_U6187 , P1_R1309_U6 , P1_R1352_U6 );
nand NAND2_3492 ( P1_U6188 , P1_U3059 , P1_U3952 );
nand NAND2_3493 ( P1_U6189 , P1_U3068 , P1_R1352_U6 );
nand NAND2_3494 ( P1_U6190 , P1_U3068 , P1_U3952 );
nand NAND2_3495 ( P1_U6191 , P1_U3055 , P1_R1352_U6 );
nand NAND2_3496 ( P1_U6192 , P1_U3055 , P1_U3952 );
nand NAND2_3497 ( P1_U6193 , P1_U3054 , P1_R1352_U6 );
nand NAND2_3498 ( P1_U6194 , P1_U3054 , P1_U3952 );
nand NAND2_3499 ( P1_U6195 , P1_U3053 , P1_R1352_U6 );
nand NAND2_3500 ( P1_U6196 , P1_U3053 , P1_U3952 );
nand NAND2_3501 ( P1_U6197 , P1_U3057 , P1_R1352_U6 );
nand NAND2_3502 ( P1_U6198 , P1_U3057 , P1_U3952 );
nand NAND2_3503 ( P1_U6199 , P1_U3058 , P1_R1352_U6 );
nand NAND2_3504 ( P1_U6200 , P1_U3058 , P1_U3952 );
nand NAND2_3505 ( P1_U6201 , P1_U3065 , P1_R1352_U6 );
nand NAND2_3506 ( P1_U6202 , P1_U3065 , P1_U3952 );
nand NAND2_3507 ( P1_U6203 , P1_U3066 , P1_R1352_U6 );
nand NAND2_3508 ( P1_U6204 , P1_U3066 , P1_U3952 );
nand NAND2_3509 ( P1_U6205 , P1_U3061 , P1_R1352_U6 );
nand NAND2_3510 ( P1_U6206 , P1_U3061 , P1_U3952 );
nand NAND2_3511 ( P1_U6207 , P1_U3075 , P1_R1352_U6 );
nand NAND2_3512 ( P1_U6208 , P1_U3075 , P1_U3952 );
nand NAND2_3513 ( P1_U6209 , P1_U3076 , P1_R1352_U6 );
nand NAND2_3514 ( P1_U6210 , P1_U3076 , P1_U3952 );
nand NAND2_3515 ( P1_U6211 , P1_U3078 , P1_R1352_U6 );
nand NAND2_3516 ( P1_U6212 , P1_U3078 , P1_U3952 );
nand NAND2_3517 ( P1_U6213 , P1_U3081 , P1_R1352_U6 );
nand NAND2_3518 ( P1_U6214 , P1_U3081 , P1_U3952 );
nand NAND2_3519 ( P1_U6215 , P1_U3082 , P1_R1352_U6 );
nand NAND2_3520 ( P1_U6216 , P1_U3082 , P1_U3952 );
nand NAND2_3521 ( P1_U6217 , P1_U3069 , P1_R1352_U6 );
nand NAND2_3522 ( P1_U6218 , P1_U3069 , P1_U3952 );
nand NAND2_3523 ( P1_U6219 , P1_U3073 , P1_R1352_U6 );
nand NAND2_3524 ( P1_U6220 , P1_U3073 , P1_U3952 );
nand NAND2_3525 ( P1_U6221 , P1_U3074 , P1_R1352_U6 );
nand NAND2_3526 ( P1_U6222 , P1_U3074 , P1_U3952 );
nand NAND2_3527 ( P1_U6223 , P1_U3079 , P1_R1352_U6 );
nand NAND2_3528 ( P1_U6224 , P1_U3079 , P1_U3952 );
nand NAND2_3529 ( P1_U6225 , P1_U3080 , P1_R1352_U6 );
nand NAND2_3530 ( P1_U6226 , P1_U3080 , P1_U3952 );
nand NAND2_3531 ( P1_U6227 , P1_U3072 , P1_R1352_U6 );
nand NAND2_3532 ( P1_U6228 , P1_U3072 , P1_U3952 );
nand NAND2_3533 ( P1_U6229 , P1_U3063 , P1_R1352_U6 );
nand NAND2_3534 ( P1_U6230 , P1_U3063 , P1_U3952 );
nand NAND2_3535 ( P1_U6231 , P1_U3062 , P1_R1352_U6 );
nand NAND2_3536 ( P1_U6232 , P1_U3062 , P1_U3952 );
nand NAND2_3537 ( P1_U6233 , P1_U3077 , P1_R1352_U6 );
nand NAND2_3538 ( P1_U6234 , P1_U3077 , P1_U3952 );
nand NAND2_3539 ( P1_U6235 , P1_U3448 , P1_U5364 );
nand NAND3_3540 ( P1_U6236 , P1_U3015 , P1_REG2_REG_0_ , P1_U5696 );
nand NAND2_3541 ( P2_R1161_U489 , P2_U3079 , P2_R1161_U61 );
nand NAND2_3542 ( P2_R1161_U488 , P2_R1161_U254 , P2_R1161_U486 );
nand NAND2_3543 ( P2_R1161_U487 , P2_R1161_U165 , P2_R1161_U166 );
nand NAND2_3544 ( P2_R1161_U486 , P2_R1161_U485 , P2_R1161_U484 );
nand NAND2_3545 ( P2_R1161_U485 , P2_U3431 , P2_R1161_U72 );
nand NAND2_3546 ( P2_R1161_U484 , P2_U3078 , P2_R1161_U71 );
nand NAND2_3547 ( P2_R1161_U483 , P2_U3431 , P2_R1161_U72 );
nand NAND2_3548 ( P2_R1161_U482 , P2_U3078 , P2_R1161_U71 );
nand NAND2_3549 ( P2_R1161_U481 , P2_R1161_U258 , P2_R1161_U479 );
nand NAND2_3550 ( P2_R1161_U480 , P2_R1161_U163 , P2_R1161_U164 );
nand NAND2_3551 ( P2_R1161_U479 , P2_R1161_U478 , P2_R1161_U477 );
nand NAND2_3552 ( P2_R1161_U478 , P2_U3434 , P2_R1161_U74 );
nand NAND2_3553 ( P2_R1161_U477 , P2_U3073 , P2_R1161_U73 );
nand NAND2_3554 ( P2_R1161_U476 , P2_U3434 , P2_R1161_U74 );
nand NAND2_3555 ( P2_R1161_U475 , P2_U3073 , P2_R1161_U73 );
nand NAND2_3556 ( P2_R1161_U474 , P2_R1161_U472 , P2_R1161_U262 );
nand NAND2_3557 ( P2_R1161_U473 , P2_R1161_U361 , P2_R1161_U92 );
nand NAND2_3558 ( P2_R1161_U472 , P2_R1161_U471 , P2_R1161_U470 );
nand NAND2_3559 ( P2_R1161_U471 , P2_U3437 , P2_R1161_U57 );
nand NAND2_3560 ( P2_R1161_U470 , P2_U3072 , P2_R1161_U56 );
nand NAND2_3561 ( P2_R1161_U469 , P2_U3440 , P2_R1161_U58 );
nand NAND2_3562 ( P2_R1161_U468 , P2_U3068 , P2_R1161_U60 );
nand NAND2_3563 ( P2_R1161_U467 , P2_R1161_U270 , P2_R1161_U465 );
nand NAND2_3564 ( P2_R1161_U466 , P2_R1161_U360 , P2_R1161_U162 );
and AND2_3565 ( P2_U3013 , P2_U3380 , P2_U5446 );
and AND2_3566 ( P2_U3014 , P2_U3380 , P2_U3379 );
and AND2_3567 ( P2_U3015 , P2_U5449 , P2_U3379 );
and AND2_3568 ( P2_U3016 , P2_U5449 , P2_U5446 );
and AND2_3569 ( P2_U3017 , P2_U3870 , P2_U5443 );
and AND2_3570 ( P2_U3018 , P2_U3587 , P2_U3582 );
and AND2_3571 ( P2_U3019 , P2_U3381 , P2_U3382 );
and AND2_3572 ( P2_U3020 , P2_U5458 , P2_U3381 );
and AND2_3573 ( P2_U3021 , P2_U5455 , P2_U3382 );
and AND2_3574 ( P2_U3022 , P2_U5458 , P2_U5455 );
and AND2_3575 ( P2_U3023 , P2_U3046 , P2_STATE_REG );
and AND2_3576 ( P2_U3024 , P2_U3701 , P2_U3366 );
and AND2_3577 ( P2_U3025 , P2_U3907 , P2_U4069 );
and AND2_3578 ( P2_U3026 , P2_U3015 , P2_U5443 );
and AND2_3579 ( P2_U3027 , P2_U3297 , P2_STATE_REG );
and AND2_3580 ( P2_U3028 , P2_U3882 , P2_U3908 );
and AND2_3581 ( P2_U3029 , P2_U3908 , P2_U3365 );
and AND2_3582 ( P2_U3030 , P2_U3698 , P2_U3908 );
and AND2_3583 ( P2_U3031 , P2_U3886 , P2_U3023 );
and AND2_3584 ( P2_U3032 , P2_U3891 , P2_U4069 );
and AND2_3585 ( P2_U3033 , P2_U3907 , P2_U4085 );
and AND2_3586 ( P2_U3034 , P2_U3908 , P2_U3025 );
and AND2_3587 ( P2_U3035 , P2_U3023 , P2_U4985 );
and AND2_3588 ( P2_U3036 , P2_U3891 , P2_U4085 );
and AND2_3589 ( P2_U3037 , P2_U5464 , P2_U4750 );
and AND2_3590 ( P2_U3038 , P2_U3024 , P2_U5464 );
and AND2_3591 ( P2_U3039 , P2_U5461 , P2_U4750 );
and AND2_3592 ( P2_U3040 , P2_U3888 , P2_U4750 );
and AND2_3593 ( P2_U3041 , P2_U3024 , P2_U3888 );
and AND2_3594 ( P2_U3042 , P2_U3023 , P2_U3366 );
and AND2_3595 ( P2_U3043 , P2_U3023 , P2_U3365 );
and AND2_3596 ( P2_U3044 , P2_U5000 , P2_STATE_REG );
and AND2_3597 ( P2_U3045 , P2_U3023 , P2_U5002 );
and AND2_3598 ( P2_U3046 , P2_U5436 , P2_U3362 );
and AND2_3599 ( P2_U3047 , P2_U3697 , P2_U3018 );
and AND2_3600 ( P2_U3048 , P2_U3696 , P2_U3018 );
and AND2_3601 ( P2_U3049 , P2_U4745 , P2_U4744 );
and AND2_3602 ( P2_U3050 , P2_U4755 , P2_STATE_REG );
and AND2_3603 ( P2_U3051 , P2_U3893 , P2_U4757 );
nand NAND4_3604 ( P2_U3052 , P2_U4534 , P2_U4533 , P2_U4532 , P2_U4531 );
nand NAND4_3605 ( P2_U3053 , P2_U4552 , P2_U4551 , P2_U4550 , P2_U4549 );
nand NAND4_3606 ( P2_U3054 , P2_U4570 , P2_U4569 , P2_U4568 , P2_U4567 );
nand NAND4_3607 ( P2_U3055 , P2_U4608 , P2_U4607 , P2_U4606 , P2_U4605 );
nand NAND4_3608 ( P2_U3056 , P2_U4516 , P2_U4515 , P2_U4514 , P2_U4513 );
nand NAND4_3609 ( P2_U3057 , P2_U4498 , P2_U4497 , P2_U4496 , P2_U4495 );
nand NAND4_3610 ( P2_U3058 , P2_U4588 , P2_U4587 , P2_U4586 , P2_U4585 );
nand NAND4_3611 ( P2_U3059 , P2_U4120 , P2_U4119 , P2_U4118 , P2_U4117 );
nand NAND4_3612 ( P2_U3060 , P2_U4444 , P2_U4443 , P2_U4442 , P2_U4441 );
nand NAND4_3613 ( P2_U3061 , P2_U4228 , P2_U4227 , P2_U4226 , P2_U4225 );
nand NAND4_3614 ( P2_U3062 , P2_U4246 , P2_U4245 , P2_U4244 , P2_U4243 );
nand NAND4_3615 ( P2_U3063 , P2_U4102 , P2_U4101 , P2_U4100 , P2_U4099 );
nand NAND4_3616 ( P2_U3064 , P2_U4480 , P2_U4479 , P2_U4478 , P2_U4477 );
nand NAND4_3617 ( P2_U3065 , P2_U4462 , P2_U4461 , P2_U4460 , P2_U4459 );
nand NAND4_3618 ( P2_U3066 , P2_U4138 , P2_U4137 , P2_U4136 , P2_U4135 );
nand NAND4_3619 ( P2_U3067 , P2_U4077 , P2_U4076 , P2_U4075 , P2_U4074 );
nand NAND4_3620 ( P2_U3068 , P2_U4354 , P2_U4353 , P2_U4352 , P2_U4351 );
nand NAND4_3621 ( P2_U3069 , P2_U4174 , P2_U4173 , P2_U4172 , P2_U4171 );
nand NAND4_3622 ( P2_U3070 , P2_U4156 , P2_U4155 , P2_U4154 , P2_U4153 );
nand NAND4_3623 ( P2_U3071 , P2_U4264 , P2_U4263 , P2_U4262 , P2_U4261 );
nand NAND4_3624 ( P2_U3072 , P2_U4336 , P2_U4335 , P2_U4334 , P2_U4333 );
nand NAND4_3625 ( P2_U3073 , P2_U4318 , P2_U4317 , P2_U4316 , P2_U4315 );
nand NAND4_3626 ( P2_U3074 , P2_U4426 , P2_U4425 , P2_U4424 , P2_U4423 );
nand NAND4_3627 ( P2_U3075 , P2_U4408 , P2_U4407 , P2_U4406 , P2_U4405 );
nand NAND4_3628 ( P2_U3076 , P2_U4082 , P2_U4081 , P2_U4080 , P2_U4079 );
nand NAND4_3629 ( P2_U3077 , P2_U4058 , P2_U4057 , P2_U4056 , P2_U4055 );
nand NAND4_3630 ( P2_U3078 , P2_U4300 , P2_U4299 , P2_U4298 , P2_U4297 );
nand NAND4_3631 ( P2_U3079 , P2_U4282 , P2_U4281 , P2_U4280 , P2_U4279 );
nand NAND4_3632 ( P2_U3080 , P2_U4390 , P2_U4389 , P2_U4388 , P2_U4387 );
nand NAND4_3633 ( P2_U3081 , P2_U4372 , P2_U4371 , P2_U4370 , P2_U4369 );
nand NAND4_3634 ( P2_U3082 , P2_U4210 , P2_U4209 , P2_U4208 , P2_U4207 );
nand NAND4_3635 ( P2_U3083 , P2_U4192 , P2_U4191 , P2_U4190 , P2_U4189 );
nand NAND2_3636 ( P2_U3084 , P2_U5337 , P2_U5336 );
nand NAND2_3637 ( P2_U3085 , P2_U5339 , P2_U5338 );
nand NAND3_3638 ( P2_U3086 , P2_U5345 , P2_U5343 , P2_U5344 );
nand NAND3_3639 ( P2_U3087 , P2_U5348 , P2_U5346 , P2_U5347 );
nand NAND3_3640 ( P2_U3088 , P2_U5351 , P2_U5349 , P2_U5350 );
nand NAND3_3641 ( P2_U3089 , P2_U5354 , P2_U5352 , P2_U5353 );
nand NAND3_3642 ( P2_U3090 , P2_U5357 , P2_U5355 , P2_U5356 );
nand NAND3_3643 ( P2_U3091 , P2_U5360 , P2_U5358 , P2_U5359 );
nand NAND3_3644 ( P2_U3092 , P2_U5363 , P2_U5361 , P2_U5362 );
nand NAND3_3645 ( P2_U3093 , P2_U5366 , P2_U5364 , P2_U5365 );
nand NAND3_3646 ( P2_U3094 , P2_U5369 , P2_U5367 , P2_U5368 );
nand NAND3_3647 ( P2_U3095 , P2_U5372 , P2_U5370 , P2_U5371 );
nand NAND3_3648 ( P2_U3096 , P2_U5377 , P2_U5378 , P2_U5376 );
nand NAND3_3649 ( P2_U3097 , P2_U5380 , P2_U5381 , P2_U5379 );
nand NAND3_3650 ( P2_U3098 , P2_U5383 , P2_U5384 , P2_U5382 );
nand NAND3_3651 ( P2_U3099 , P2_U5386 , P2_U5387 , P2_U5385 );
nand NAND3_3652 ( P2_U3100 , P2_U5389 , P2_U5390 , P2_U5388 );
nand NAND3_3653 ( P2_U3101 , P2_U5392 , P2_U5393 , P2_U5391 );
nand NAND3_3654 ( P2_U3102 , P2_U5395 , P2_U5396 , P2_U5394 );
nand NAND3_3655 ( P2_U3103 , P2_U5398 , P2_U5399 , P2_U5397 );
nand NAND3_3656 ( P2_U3104 , P2_U5401 , P2_U5402 , P2_U5400 );
nand NAND3_3657 ( P2_U3105 , P2_U5404 , P2_U5405 , P2_U5403 );
nand NAND3_3658 ( P2_U3106 , P2_U5319 , P2_U5320 , P2_U5318 );
nand NAND3_3659 ( P2_U3107 , P2_U5322 , P2_U5323 , P2_U5321 );
nand NAND3_3660 ( P2_U3108 , P2_U5325 , P2_U5326 , P2_U5324 );
nand NAND3_3661 ( P2_U3109 , P2_U5328 , P2_U5329 , P2_U5327 );
nand NAND3_3662 ( P2_U3110 , P2_U5331 , P2_U5332 , P2_U5330 );
nand NAND3_3663 ( P2_U3111 , P2_U5334 , P2_U5333 , P2_U5335 );
nand NAND3_3664 ( P2_U3112 , P2_U5341 , P2_U5340 , P2_U5342 );
nand NAND3_3665 ( P2_U3113 , P2_U5374 , P2_U5373 , P2_U5375 );
nand NAND3_3666 ( P2_U3114 , P2_U5407 , P2_U5406 , P2_U5408 );
nand NAND2_3667 ( P2_U3115 , P2_U5410 , P2_U5409 );
nand NAND2_3668 ( P2_U3116 , P2_U5267 , P2_U5266 );
nand NAND2_3669 ( P2_U3117 , P2_U5269 , P2_U5268 );
nand NAND3_3670 ( P2_U3118 , P2_U5273 , P2_U3375 , P2_U5272 );
nand NAND3_3671 ( P2_U3119 , P2_U5275 , P2_U3375 , P2_U5274 );
nand NAND3_3672 ( P2_U3120 , P2_U5277 , P2_U3375 , P2_U5276 );
nand NAND3_3673 ( P2_U3121 , P2_U5279 , P2_U3375 , P2_U5278 );
nand NAND3_3674 ( P2_U3122 , P2_U5281 , P2_U3375 , P2_U5280 );
nand NAND3_3675 ( P2_U3123 , P2_U5283 , P2_U3375 , P2_U5282 );
nand NAND3_3676 ( P2_U3124 , P2_U5285 , P2_U3375 , P2_U5284 );
nand NAND3_3677 ( P2_U3125 , P2_U5287 , P2_U3375 , P2_U5286 );
nand NAND3_3678 ( P2_U3126 , P2_U5289 , P2_U3375 , P2_U5288 );
nand NAND3_3679 ( P2_U3127 , P2_U5291 , P2_U3375 , P2_U5290 );
nand NAND3_3680 ( P2_U3128 , P2_U5295 , P2_U3375 , P2_U5294 );
nand NAND3_3681 ( P2_U3129 , P2_U5297 , P2_U3375 , P2_U5296 );
nand NAND3_3682 ( P2_U3130 , P2_U5299 , P2_U3375 , P2_U5298 );
nand NAND3_3683 ( P2_U3131 , P2_U5301 , P2_U3375 , P2_U5300 );
nand NAND3_3684 ( P2_U3132 , P2_U5303 , P2_U3375 , P2_U5302 );
nand NAND3_3685 ( P2_U3133 , P2_U5305 , P2_U3375 , P2_U5304 );
nand NAND3_3686 ( P2_U3134 , P2_U5307 , P2_U3375 , P2_U5306 );
nand NAND3_3687 ( P2_U3135 , P2_U5309 , P2_U3375 , P2_U5308 );
nand NAND3_3688 ( P2_U3136 , P2_U5311 , P2_U3375 , P2_U5310 );
nand NAND3_3689 ( P2_U3137 , P2_U5313 , P2_U3375 , P2_U5312 );
nand NAND3_3690 ( P2_U3138 , P2_U5255 , P2_U3375 , P2_U5254 );
nand NAND3_3691 ( P2_U3139 , P2_U5257 , P2_U3375 , P2_U5256 );
nand NAND3_3692 ( P2_U3140 , P2_U5259 , P2_U3375 , P2_U5258 );
nand NAND3_3693 ( P2_U3141 , P2_U5261 , P2_U3375 , P2_U5260 );
nand NAND3_3694 ( P2_U3142 , P2_U5263 , P2_U3375 , P2_U5262 );
nand NAND2_3695 ( P2_U3143 , P2_U3822 , P2_U5265 );
nand NAND2_3696 ( P2_U3144 , P2_U3823 , P2_U5271 );
nand NAND2_3697 ( P2_U3145 , P2_U3824 , P2_U5293 );
nand NAND2_3698 ( P2_U3146 , P2_U3825 , P2_U5315 );
nand NAND2_3699 ( P2_U3147 , P2_U3826 , P2_U5317 );
nand NAND3_3700 ( P2_U3148 , P2_U3385 , P2_U5449 , P2_U3375 );
nand NAND2_3701 ( P2_U3149 , P2_U3818 , P2_U3013 );
nand NAND2_3702 ( P2_U3150 , P2_U3817 , P2_U5249 );
not NOT1_3703 ( P2_U3151 , P2_STATE_REG );
nand NAND3_3704 ( P2_U3152 , P2_U5940 , P2_U5939 , P2_U3359 );
nand NAND4_3705 ( P2_U3153 , P2_U5245 , P2_U5244 , P2_U3816 , P2_U5246 );
nand NAND4_3706 ( P2_U3154 , P2_U5236 , P2_U3815 , P2_U5235 , P2_U5237 );
nand NAND4_3707 ( P2_U3155 , P2_U5227 , P2_U5226 , P2_U3814 , P2_U5228 );
nand NAND4_3708 ( P2_U3156 , P2_U5218 , P2_U3813 , P2_U5217 , P2_U5219 );
nand NAND4_3709 ( P2_U3157 , P2_U5209 , P2_U5208 , P2_U3812 , P2_U5210 );
nand NAND3_3710 ( P2_U3158 , P2_U3810 , P2_U5200 , P2_U3811 );
nand NAND4_3711 ( P2_U3159 , P2_U5191 , P2_U3809 , P2_U5190 , P2_U5192 );
nand NAND4_3712 ( P2_U3160 , P2_U5182 , P2_U3808 , P2_U5181 , P2_U5183 );
nand NAND4_3713 ( P2_U3161 , P2_U5173 , P2_U5172 , P2_U3807 , P2_U5174 );
nand NAND3_3714 ( P2_U3162 , P2_U3805 , P2_U5164 , P2_U3806 );
nand NAND4_3715 ( P2_U3163 , P2_U5155 , P2_U3804 , P2_U5154 , P2_U5156 );
nand NAND4_3716 ( P2_U3164 , P2_U5146 , P2_U5145 , P2_U3803 , P2_U5147 );
nand NAND4_3717 ( P2_U3165 , P2_U5137 , P2_U3802 , P2_U5136 , P2_U5138 );
nand NAND4_3718 ( P2_U3166 , P2_U5128 , P2_U5127 , P2_U3801 , P2_U5129 );
nand NAND4_3719 ( P2_U3167 , P2_U5119 , P2_U5118 , P2_U3800 , P2_U5120 );
nand NAND4_3720 ( P2_U3168 , P2_U5110 , P2_U5109 , P2_U3799 , P2_U5111 );
nand NAND4_3721 ( P2_U3169 , P2_U5101 , P2_U3798 , P2_U5100 , P2_U5102 );
nand NAND3_3722 ( P2_U3170 , P2_U3796 , P2_U5092 , P2_U3797 );
nand NAND4_3723 ( P2_U3171 , P2_U5083 , P2_U5082 , P2_U3795 , P2_U5084 );
nand NAND2_3724 ( P2_U3172 , P2_U5075 , P2_U3794 );
nand NAND4_3725 ( P2_U3173 , P2_U5067 , P2_U3791 , P2_U5066 , P2_U5068 );
nand NAND4_3726 ( P2_U3174 , P2_U5058 , P2_U5057 , P2_U3790 , P2_U5059 );
nand NAND4_3727 ( P2_U3175 , P2_U5049 , P2_U3789 , P2_U5048 , P2_U5050 );
nand NAND4_3728 ( P2_U3176 , P2_U5040 , P2_U5039 , P2_U3788 , P2_U5041 );
nand NAND3_3729 ( P2_U3177 , P2_U3786 , P2_U5031 , P2_U3787 );
nand NAND4_3730 ( P2_U3178 , P2_U5022 , P2_U5021 , P2_U3785 , P2_U5023 );
nand NAND4_3731 ( P2_U3179 , P2_U5013 , P2_U5012 , P2_U3784 , P2_U5014 );
nand NAND4_3732 ( P2_U3180 , P2_U5004 , P2_U3783 , P2_U5003 , P2_U5005 );
nand NAND4_3733 ( P2_U3181 , P2_U4991 , P2_U4990 , P2_U3782 , P2_U4992 );
nand NAND2_3734 ( P2_U3182 , P2_U4969 , P2_U3761 );
nand NAND2_3735 ( P2_U3183 , P2_U4958 , P2_U3758 );
nand NAND2_3736 ( P2_U3184 , P2_U4947 , P2_U3755 );
nand NAND3_3737 ( P2_U3185 , P2_U4937 , P2_U4936 , P2_U3752 );
nand NAND3_3738 ( P2_U3186 , P2_U4926 , P2_U4925 , P2_U3749 );
nand NAND4_3739 ( P2_U3187 , P2_U4914 , P2_U3746 , P2_U3748 , P2_U4912 );
nand NAND3_3740 ( P2_U3188 , P2_U4903 , P2_U3743 , P2_U4901 );
nand NAND3_3741 ( P2_U3189 , P2_U3741 , P2_U4892 , P2_U3740 );
nand NAND3_3742 ( P2_U3190 , P2_U3738 , P2_U4881 , P2_U3737 );
nand NAND2_3743 ( P2_U3191 , P2_U4870 , P2_U3734 );
nand NAND2_3744 ( P2_U3192 , P2_U4859 , P2_U3731 );
nand NAND2_3745 ( P2_U3193 , P2_U4848 , P2_U3728 );
nand NAND2_3746 ( P2_U3194 , P2_U4837 , P2_U3725 );
nand NAND2_3747 ( P2_U3195 , P2_U4826 , P2_U3722 );
nand NAND2_3748 ( P2_U3196 , P2_U4815 , P2_U3719 );
nand NAND2_3749 ( P2_U3197 , P2_U4804 , P2_U3716 );
nand NAND2_3750 ( P2_U3198 , P2_U4793 , P2_U3713 );
nand NAND2_3751 ( P2_U3199 , P2_U4782 , P2_U3710 );
nand NAND2_3752 ( P2_U3200 , P2_U4771 , P2_U3707 );
nand NAND2_3753 ( P2_U3201 , P2_U4760 , P2_U3704 );
nand NAND3_3754 ( P2_U3202 , P2_U4749 , P2_U3049 , P2_U4748 );
nand NAND3_3755 ( P2_U3203 , P2_U4747 , P2_U3049 , P2_U4746 );
nand NAND4_3756 ( P2_U3204 , P2_U4742 , P2_U4743 , P2_U4741 , P2_U3862 );
nand NAND5_3757 ( P2_U3205 , P2_U4739 , P2_U4737 , P2_U4740 , P2_U4738 , P2_U3861 );
nand NAND5_3758 ( P2_U3206 , P2_U4735 , P2_U4733 , P2_U4736 , P2_U4734 , P2_U3860 );
nand NAND5_3759 ( P2_U3207 , P2_U4731 , P2_U4729 , P2_U4732 , P2_U4730 , P2_U3859 );
nand NAND5_3760 ( P2_U3208 , P2_U4727 , P2_U4725 , P2_U4728 , P2_U4726 , P2_U3858 );
nand NAND5_3761 ( P2_U3209 , P2_U4723 , P2_U4721 , P2_U4724 , P2_U4722 , P2_U3857 );
nand NAND5_3762 ( P2_U3210 , P2_U4719 , P2_U4717 , P2_U4720 , P2_U4718 , P2_U3856 );
nand NAND5_3763 ( P2_U3211 , P2_U4715 , P2_U4713 , P2_U4716 , P2_U4714 , P2_U3855 );
nand NAND5_3764 ( P2_U3212 , P2_U4711 , P2_U4709 , P2_U4712 , P2_U4710 , P2_U3854 );
nand NAND5_3765 ( P2_U3213 , P2_U4707 , P2_U4705 , P2_U4708 , P2_U4706 , P2_U3853 );
nand NAND5_3766 ( P2_U3214 , P2_U4703 , P2_U4701 , P2_U4704 , P2_U4702 , P2_U3852 );
nand NAND5_3767 ( P2_U3215 , P2_U4699 , P2_U4697 , P2_U4700 , P2_U4698 , P2_U3851 );
nand NAND5_3768 ( P2_U3216 , P2_U4695 , P2_U4693 , P2_U4696 , P2_U4694 , P2_U3850 );
nand NAND5_3769 ( P2_U3217 , P2_U4691 , P2_U4689 , P2_U4692 , P2_U4690 , P2_U3849 );
nand NAND5_3770 ( P2_U3218 , P2_U4687 , P2_U4685 , P2_U4688 , P2_U4686 , P2_U3848 );
nand NAND5_3771 ( P2_U3219 , P2_U4683 , P2_U4681 , P2_U4684 , P2_U4682 , P2_U3847 );
nand NAND5_3772 ( P2_U3220 , P2_U4679 , P2_U4677 , P2_U4680 , P2_U4678 , P2_U3846 );
nand NAND5_3773 ( P2_U3221 , P2_U4675 , P2_U4673 , P2_U4676 , P2_U4674 , P2_U3845 );
nand NAND5_3774 ( P2_U3222 , P2_U4671 , P2_U4669 , P2_U4672 , P2_U4670 , P2_U3844 );
nand NAND5_3775 ( P2_U3223 , P2_U4667 , P2_U4665 , P2_U4668 , P2_U4666 , P2_U3843 );
nand NAND5_3776 ( P2_U3224 , P2_U4663 , P2_U4661 , P2_U4664 , P2_U4662 , P2_U3842 );
nand NAND5_3777 ( P2_U3225 , P2_U4660 , P2_U4659 , P2_U4658 , P2_U4657 , P2_U3841 );
nand NAND5_3778 ( P2_U3226 , P2_U4656 , P2_U4655 , P2_U4654 , P2_U4653 , P2_U3840 );
nand NAND5_3779 ( P2_U3227 , P2_U4650 , P2_U4649 , P2_U4651 , P2_U3839 , P2_U4652 );
nand NAND5_3780 ( P2_U3228 , P2_U4646 , P2_U4645 , P2_U4647 , P2_U3838 , P2_U4648 );
nand NAND5_3781 ( P2_U3229 , P2_U4642 , P2_U4641 , P2_U4643 , P2_U3837 , P2_U4644 );
nand NAND5_3782 ( P2_U3230 , P2_U4638 , P2_U4637 , P2_U4639 , P2_U3836 , P2_U4640 );
nand NAND5_3783 ( P2_U3231 , P2_U4634 , P2_U4633 , P2_U4635 , P2_U3835 , P2_U4636 );
nand NAND5_3784 ( P2_U3232 , P2_U4630 , P2_U4629 , P2_U4631 , P2_U3834 , P2_U4632 );
nand NAND5_3785 ( P2_U3233 , P2_U4626 , P2_U4625 , P2_U4627 , P2_U3833 , P2_U4628 );
and AND2_3786 ( P2_U3234 , P2_D_REG_31_ , P2_U3828 );
and AND2_3787 ( P2_U3235 , P2_D_REG_30_ , P2_U3828 );
and AND2_3788 ( P2_U3236 , P2_D_REG_29_ , P2_U3828 );
and AND2_3789 ( P2_U3237 , P2_D_REG_28_ , P2_U3828 );
and AND2_3790 ( P2_U3238 , P2_D_REG_27_ , P2_U3828 );
and AND2_3791 ( P2_U3239 , P2_D_REG_26_ , P2_U3828 );
and AND2_3792 ( P2_U3240 , P2_D_REG_25_ , P2_U3828 );
and AND2_3793 ( P2_U3241 , P2_D_REG_24_ , P2_U3828 );
and AND2_3794 ( P2_U3242 , P2_D_REG_23_ , P2_U3828 );
and AND2_3795 ( P2_U3243 , P2_D_REG_22_ , P2_U3828 );
and AND2_3796 ( P2_U3244 , P2_D_REG_21_ , P2_U3828 );
and AND2_3797 ( P2_U3245 , P2_D_REG_20_ , P2_U3828 );
and AND2_3798 ( P2_U3246 , P2_D_REG_19_ , P2_U3828 );
and AND2_3799 ( P2_U3247 , P2_D_REG_18_ , P2_U3828 );
and AND2_3800 ( P2_U3248 , P2_D_REG_17_ , P2_U3828 );
and AND2_3801 ( P2_U3249 , P2_D_REG_16_ , P2_U3828 );
and AND2_3802 ( P2_U3250 , P2_D_REG_15_ , P2_U3828 );
and AND2_3803 ( P2_U3251 , P2_D_REG_14_ , P2_U3828 );
and AND2_3804 ( P2_U3252 , P2_D_REG_13_ , P2_U3828 );
and AND2_3805 ( P2_U3253 , P2_D_REG_12_ , P2_U3828 );
and AND2_3806 ( P2_U3254 , P2_D_REG_11_ , P2_U3828 );
and AND2_3807 ( P2_U3255 , P2_D_REG_10_ , P2_U3828 );
and AND2_3808 ( P2_U3256 , P2_D_REG_9_ , P2_U3828 );
and AND2_3809 ( P2_U3257 , P2_D_REG_8_ , P2_U3828 );
and AND2_3810 ( P2_U3258 , P2_D_REG_7_ , P2_U3828 );
and AND2_3811 ( P2_U3259 , P2_D_REG_6_ , P2_U3828 );
and AND2_3812 ( P2_U3260 , P2_D_REG_5_ , P2_U3828 );
and AND2_3813 ( P2_U3261 , P2_D_REG_4_ , P2_U3828 );
and AND2_3814 ( P2_U3262 , P2_D_REG_3_ , P2_U3828 );
and AND2_3815 ( P2_U3263 , P2_D_REG_2_ , P2_U3828 );
nand NAND3_3816 ( P2_U3264 , P2_U4012 , P2_U4013 , P2_U4011 );
nand NAND3_3817 ( P2_U3265 , P2_U4009 , P2_U4010 , P2_U4008 );
nand NAND3_3818 ( P2_U3266 , P2_U4006 , P2_U4007 , P2_U4005 );
nand NAND3_3819 ( P2_U3267 , P2_U4003 , P2_U4004 , P2_U4002 );
nand NAND3_3820 ( P2_U3268 , P2_U4000 , P2_U4001 , P2_U3999 );
nand NAND3_3821 ( P2_U3269 , P2_U3997 , P2_U3998 , P2_U3996 );
nand NAND3_3822 ( P2_U3270 , P2_U3994 , P2_U3995 , P2_U3993 );
nand NAND3_3823 ( P2_U3271 , P2_U3991 , P2_U3992 , P2_U3990 );
nand NAND3_3824 ( P2_U3272 , P2_U3988 , P2_U3989 , P2_U3987 );
nand NAND3_3825 ( P2_U3273 , P2_U3985 , P2_U3986 , P2_U3984 );
nand NAND3_3826 ( P2_U3274 , P2_U3982 , P2_U3983 , P2_U3981 );
nand NAND3_3827 ( P2_U3275 , P2_U3979 , P2_U3980 , P2_U3978 );
nand NAND3_3828 ( P2_U3276 , P2_U3976 , P2_U3977 , P2_U3975 );
nand NAND3_3829 ( P2_U3277 , P2_U3973 , P2_U3974 , P2_U3972 );
nand NAND3_3830 ( P2_U3278 , P2_U3970 , P2_U3971 , P2_U3969 );
nand NAND3_3831 ( P2_U3279 , P2_U3967 , P2_U3968 , P2_U3966 );
nand NAND3_3832 ( P2_U3280 , P2_U3964 , P2_U3965 , P2_U3963 );
nand NAND3_3833 ( P2_U3281 , P2_U3961 , P2_U3962 , P2_U3960 );
nand NAND3_3834 ( P2_U3282 , P2_U3958 , P2_U3959 , P2_U3957 );
nand NAND3_3835 ( P2_U3283 , P2_U3955 , P2_U3956 , P2_U3954 );
nand NAND3_3836 ( P2_U3284 , P2_U3952 , P2_U3953 , P2_U3951 );
nand NAND3_3837 ( P2_U3285 , P2_U3949 , P2_U3950 , P2_U3948 );
nand NAND3_3838 ( P2_U3286 , P2_U3946 , P2_U3947 , P2_U3945 );
nand NAND3_3839 ( P2_U3287 , P2_U3943 , P2_U3944 , P2_U3942 );
nand NAND3_3840 ( P2_U3288 , P2_U3940 , P2_U3941 , P2_U3939 );
nand NAND3_3841 ( P2_U3289 , P2_U3937 , P2_U3938 , P2_U3936 );
nand NAND3_3842 ( P2_U3290 , P2_U3934 , P2_U3935 , P2_U3933 );
nand NAND3_3843 ( P2_U3291 , P2_U3931 , P2_U3932 , P2_U3930 );
nand NAND3_3844 ( P2_U3292 , P2_U3928 , P2_U3929 , P2_U3927 );
nand NAND3_3845 ( P2_U3293 , P2_U3925 , P2_U3926 , P2_U3924 );
nand NAND3_3846 ( P2_U3294 , P2_U3922 , P2_U3923 , P2_U3921 );
nand NAND3_3847 ( P2_U3295 , P2_U3919 , P2_U3920 , P2_U3918 );
and AND2_3848 ( P2_U3296 , P2_U3780 , P2_U5417 );
nand NAND2_3849 ( P2_U3297 , P2_STATE_REG , P2_U3827 );
not NOT1_3850 ( P2_U3298 , P2_B_REG );
nand NAND2_3851 ( P2_U3299 , P2_U3374 , P2_U5427 );
nand NAND2_3852 ( P2_U3300 , P2_U3374 , P2_U4014 );
nand NAND2_3853 ( P2_U3301 , P2_U3013 , P2_U5443 );
nand NAND2_3854 ( P2_U3302 , P2_U3014 , P2_U5452 );
nand NAND2_3855 ( P2_U3303 , P2_U3588 , P2_U3018 );
nand NAND2_3856 ( P2_U3304 , P2_U3589 , P2_U3018 );
nand NAND2_3857 ( P2_U3305 , P2_U3014 , P2_U5443 );
nand NAND2_3858 ( P2_U3306 , P2_U3014 , P2_U3378 );
nand NAND2_3859 ( P2_U3307 , P2_U3013 , P2_U3378 );
nand NAND3_3860 ( P2_U3308 , P2_U3385 , P2_U3379 , P2_U3378 );
nand NAND3_3861 ( P2_U3309 , P2_U5446 , P2_U3385 , P2_U3378 );
nand NAND2_3862 ( P2_U3310 , P2_U5452 , P2_U3013 );
nand NAND2_3863 ( P2_U3311 , P2_U3874 , P2_U5443 );
nand NAND2_3864 ( P2_U3312 , P2_U3016 , P2_U3385 );
nand NAND2_3865 ( P2_U3313 , P2_U3385 , P2_U3380 );
nand NAND5_3866 ( P2_U3314 , P2_U4066 , P2_U4065 , P2_U4067 , P2_U3576 , P2_U3575 );
nand NAND4_3867 ( P2_U3315 , P2_U4087 , P2_U4086 , P2_U3590 , P2_U3592 );
nand NAND4_3868 ( P2_U3316 , P2_U4105 , P2_U4104 , P2_U3594 , P2_U3596 );
nand NAND4_3869 ( P2_U3317 , P2_U4123 , P2_U4122 , P2_U3598 , P2_U3600 );
nand NAND4_3870 ( P2_U3318 , P2_U4141 , P2_U4140 , P2_U3602 , P2_U3604 );
nand NAND4_3871 ( P2_U3319 , P2_U4159 , P2_U4158 , P2_U3606 , P2_U3608 );
nand NAND4_3872 ( P2_U3320 , P2_U4177 , P2_U4176 , P2_U3610 , P2_U3612 );
nand NAND4_3873 ( P2_U3321 , P2_U4195 , P2_U4194 , P2_U3614 , P2_U3616 );
nand NAND5_3874 ( P2_U3322 , P2_U4213 , P2_U4212 , P2_U4214 , P2_U4215 , P2_U3619 );
nand NAND5_3875 ( P2_U3323 , P2_U4231 , P2_U4230 , P2_U4232 , P2_U4233 , P2_U3622 );
nand NAND5_3876 ( P2_U3324 , P2_U4249 , P2_U4248 , P2_U4250 , P2_U4251 , P2_U3625 );
nand NAND5_3877 ( P2_U3325 , P2_U4267 , P2_U4266 , P2_U4268 , P2_U4269 , P2_U3628 );
nand NAND4_3878 ( P2_U3326 , P2_U4285 , P2_U4284 , P2_U3630 , P2_U3632 );
nand NAND4_3879 ( P2_U3327 , P2_U4303 , P2_U4302 , P2_U3634 , P2_U3636 );
nand NAND5_3880 ( P2_U3328 , P2_U4321 , P2_U4320 , P2_U4322 , P2_U4323 , P2_U3639 );
nand NAND5_3881 ( P2_U3329 , P2_U4339 , P2_U4338 , P2_U4340 , P2_U4341 , P2_U3642 );
nand NAND5_3882 ( P2_U3330 , P2_U4357 , P2_U4356 , P2_U4358 , P2_U4359 , P2_U3645 );
nand NAND4_3883 ( P2_U3331 , P2_U4375 , P2_U4374 , P2_U3647 , P2_U3649 );
nand NAND4_3884 ( P2_U3332 , P2_U4393 , P2_U4392 , P2_U3651 , P2_U3653 );
nand NAND4_3885 ( P2_U3333 , P2_U4411 , P2_U4410 , P2_U3655 , P2_U3657 );
nand NAND2_3886 ( P2_U3334 , U44 , P2_U3829 );
nand NAND4_3887 ( P2_U3335 , P2_U4429 , P2_U4428 , P2_U3659 , P2_U3661 );
nand NAND2_3888 ( P2_U3336 , U43 , P2_U3829 );
nand NAND5_3889 ( P2_U3337 , P2_U4447 , P2_U4446 , P2_U4448 , P2_U4449 , P2_U3664 );
nand NAND2_3890 ( P2_U3338 , U42 , P2_U3829 );
nand NAND5_3891 ( P2_U3339 , P2_U4465 , P2_U4464 , P2_U4466 , P2_U4467 , P2_U3667 );
nand NAND2_3892 ( P2_U3340 , U41 , P2_U3829 );
nand NAND5_3893 ( P2_U3341 , P2_U4483 , P2_U4482 , P2_U4484 , P2_U4485 , P2_U3670 );
nand NAND2_3894 ( P2_U3342 , U40 , P2_U3829 );
nand NAND4_3895 ( P2_U3343 , P2_U4501 , P2_U4500 , P2_U3672 , P2_U3674 );
nand NAND2_3896 ( P2_U3344 , U39 , P2_U3829 );
nand NAND4_3897 ( P2_U3345 , P2_U4519 , P2_U4518 , P2_U3676 , P2_U3678 );
nand NAND2_3898 ( P2_U3346 , U38 , P2_U3829 );
nand NAND4_3899 ( P2_U3347 , P2_U4537 , P2_U4536 , P2_U3680 , P2_U3682 );
nand NAND2_3900 ( P2_U3348 , U37 , P2_U3829 );
nand NAND4_3901 ( P2_U3349 , P2_U4555 , P2_U4554 , P2_U3684 , P2_U3686 );
nand NAND2_3902 ( P2_U3350 , U36 , P2_U3829 );
nand NAND4_3903 ( P2_U3351 , P2_U4573 , P2_U4572 , P2_U3688 , P2_U3690 );
nand NAND2_3904 ( P2_U3352 , P2_U3383 , P2_U3384 );
nand NAND2_3905 ( P2_U3353 , U35 , P2_U3829 );
nand NAND2_3906 ( P2_U3354 , P2_U3694 , P2_U3692 );
nand NAND2_3907 ( P2_U3355 , U33 , P2_U3829 );
nand NAND2_3908 ( P2_U3356 , U32 , P2_U3829 );
nand NAND2_3909 ( P2_U3357 , P2_U3015 , P2_U5452 );
nand NAND2_3910 ( P2_U3358 , P2_U3023 , P2_U4623 );
nand NAND2_3911 ( P2_U3359 , P2_U5443 , P2_U3385 );
nand NAND2_3912 ( P2_U3360 , P2_U3875 , P2_U5443 );
nand NAND3_3913 ( P2_U3361 , P2_U3907 , P2_U4591 , P2_U3055 );
nand NAND3_3914 ( P2_U3362 , P2_U3373 , P2_U3374 , P2_U3372 );
nand NAND2_3915 ( P2_U3363 , P2_U3699 , P2_U3906 );
nand NAND2_3916 ( P2_U3364 , P2_U3313 , P2_U3829 );
nand NAND2_3917 ( P2_U3365 , P2_U3873 , P2_U5419 );
nand NAND2_3918 ( P2_U3366 , P2_U3700 , P2_U3050 );
nand NAND2_3919 ( P2_U3367 , P2_U3878 , P2_U3385 );
nand NAND2_3920 ( P2_U3368 , P2_U3764 , P2_U3886 );
nand NAND2_3921 ( P2_U3369 , P2_U3872 , P2_U3378 );
nand NAND3_3922 ( P2_U3370 , P2_U4988 , P2_U4987 , P2_U3781 );
nand NAND2_3923 ( P2_U3371 , P2_U5413 , P2_U3913 );
nand NAND2_3924 ( P2_U3372 , P2_U5423 , P2_U5422 );
nand NAND2_3925 ( P2_U3373 , P2_U5426 , P2_U5425 );
nand NAND2_3926 ( P2_U3374 , P2_U5429 , P2_U5428 );
nand NAND2_3927 ( P2_U3375 , P2_U5435 , P2_U5434 );
nand NAND2_3928 ( P2_U3376 , P2_U5438 , P2_U5437 );
nand NAND2_3929 ( P2_U3377 , P2_U5440 , P2_U5439 );
nand NAND2_3930 ( P2_U3378 , P2_U5442 , P2_U5441 );
nand NAND2_3931 ( P2_U3379 , P2_U5445 , P2_U5444 );
nand NAND2_3932 ( P2_U3380 , P2_U5448 , P2_U5447 );
nand NAND2_3933 ( P2_U3381 , P2_U5454 , P2_U5453 );
nand NAND2_3934 ( P2_U3382 , P2_U5457 , P2_U5456 );
nand NAND2_3935 ( P2_U3383 , P2_U5460 , P2_U5459 );
nand NAND2_3936 ( P2_U3384 , P2_U5463 , P2_U5462 );
nand NAND2_3937 ( P2_U3385 , P2_U5451 , P2_U5450 );
nand NAND2_3938 ( P2_U3386 , P2_U5466 , P2_U5465 );
nand NAND2_3939 ( P2_U3387 , P2_U5468 , P2_U5467 );
nand NAND2_3940 ( P2_U3388 , P2_U5471 , P2_U5470 );
nand NAND2_3941 ( P2_U3389 , P2_U5474 , P2_U5473 );
nand NAND2_3942 ( P2_U3390 , P2_U5480 , P2_U5479 );
nand NAND2_3943 ( P2_U3391 , P2_U5482 , P2_U5481 );
nand NAND2_3944 ( P2_U3392 , P2_U5484 , P2_U5483 );
nand NAND2_3945 ( P2_U3393 , P2_U5487 , P2_U5486 );
nand NAND2_3946 ( P2_U3394 , P2_U5489 , P2_U5488 );
nand NAND2_3947 ( P2_U3395 , P2_U5491 , P2_U5490 );
nand NAND2_3948 ( P2_U3396 , P2_U5494 , P2_U5493 );
nand NAND2_3949 ( P2_U3397 , P2_U5496 , P2_U5495 );
nand NAND2_3950 ( P2_U3398 , P2_U5498 , P2_U5497 );
nand NAND2_3951 ( P2_U3399 , P2_U5501 , P2_U5500 );
nand NAND2_3952 ( P2_U3400 , P2_U5503 , P2_U5502 );
nand NAND2_3953 ( P2_U3401 , P2_U5505 , P2_U5504 );
nand NAND2_3954 ( P2_U3402 , P2_U5508 , P2_U5507 );
nand NAND2_3955 ( P2_U3403 , P2_U5510 , P2_U5509 );
nand NAND2_3956 ( P2_U3404 , P2_U5512 , P2_U5511 );
nand NAND2_3957 ( P2_U3405 , P2_U5515 , P2_U5514 );
nand NAND2_3958 ( P2_U3406 , P2_U5517 , P2_U5516 );
nand NAND2_3959 ( P2_U3407 , P2_U5519 , P2_U5518 );
nand NAND2_3960 ( P2_U3408 , P2_U5522 , P2_U5521 );
nand NAND2_3961 ( P2_U3409 , P2_U5524 , P2_U5523 );
nand NAND2_3962 ( P2_U3410 , P2_U5526 , P2_U5525 );
nand NAND2_3963 ( P2_U3411 , P2_U5529 , P2_U5528 );
nand NAND2_3964 ( P2_U3412 , P2_U5531 , P2_U5530 );
nand NAND2_3965 ( P2_U3413 , P2_U5533 , P2_U5532 );
nand NAND2_3966 ( P2_U3414 , P2_U5536 , P2_U5535 );
nand NAND2_3967 ( P2_U3415 , P2_U5538 , P2_U5537 );
nand NAND2_3968 ( P2_U3416 , P2_U5540 , P2_U5539 );
nand NAND2_3969 ( P2_U3417 , P2_U5543 , P2_U5542 );
nand NAND2_3970 ( P2_U3418 , P2_U5545 , P2_U5544 );
nand NAND2_3971 ( P2_U3419 , P2_U5547 , P2_U5546 );
nand NAND2_3972 ( P2_U3420 , P2_U5550 , P2_U5549 );
nand NAND2_3973 ( P2_U3421 , P2_U5552 , P2_U5551 );
nand NAND2_3974 ( P2_U3422 , P2_U5554 , P2_U5553 );
nand NAND2_3975 ( P2_U3423 , P2_U5557 , P2_U5556 );
nand NAND2_3976 ( P2_U3424 , P2_U5559 , P2_U5558 );
nand NAND2_3977 ( P2_U3425 , P2_U5561 , P2_U5560 );
nand NAND2_3978 ( P2_U3426 , P2_U5564 , P2_U5563 );
nand NAND2_3979 ( P2_U3427 , P2_U5566 , P2_U5565 );
nand NAND2_3980 ( P2_U3428 , P2_U5568 , P2_U5567 );
nand NAND2_3981 ( P2_U3429 , P2_U5571 , P2_U5570 );
nand NAND2_3982 ( P2_U3430 , P2_U5573 , P2_U5572 );
nand NAND2_3983 ( P2_U3431 , P2_U5575 , P2_U5574 );
nand NAND2_3984 ( P2_U3432 , P2_U5578 , P2_U5577 );
nand NAND2_3985 ( P2_U3433 , P2_U5580 , P2_U5579 );
nand NAND2_3986 ( P2_U3434 , P2_U5582 , P2_U5581 );
nand NAND2_3987 ( P2_U3435 , P2_U5585 , P2_U5584 );
nand NAND2_3988 ( P2_U3436 , P2_U5587 , P2_U5586 );
nand NAND2_3989 ( P2_U3437 , P2_U5589 , P2_U5588 );
nand NAND2_3990 ( P2_U3438 , P2_U5592 , P2_U5591 );
nand NAND2_3991 ( P2_U3439 , P2_U5594 , P2_U5593 );
nand NAND2_3992 ( P2_U3440 , P2_U5596 , P2_U5595 );
nand NAND2_3993 ( P2_U3441 , P2_U5599 , P2_U5598 );
nand NAND2_3994 ( P2_U3442 , P2_U5601 , P2_U5600 );
nand NAND2_3995 ( P2_U3443 , P2_U5603 , P2_U5602 );
nand NAND2_3996 ( P2_U3444 , P2_U5606 , P2_U5605 );
nand NAND2_3997 ( P2_U3445 , P2_U5608 , P2_U5607 );
nand NAND2_3998 ( P2_U3446 , P2_U5611 , P2_U5610 );
nand NAND2_3999 ( P2_U3447 , P2_U5613 , P2_U5612 );
nand NAND2_4000 ( P2_U3448 , P2_U5615 , P2_U5614 );
nand NAND2_4001 ( P2_U3449 , P2_U5617 , P2_U5616 );
nand NAND2_4002 ( P2_U3450 , P2_U5619 , P2_U5618 );
nand NAND2_4003 ( P2_U3451 , P2_U5621 , P2_U5620 );
nand NAND2_4004 ( P2_U3452 , P2_U5623 , P2_U5622 );
nand NAND2_4005 ( P2_U3453 , P2_U5625 , P2_U5624 );
nand NAND2_4006 ( P2_U3454 , P2_U5627 , P2_U5626 );
nand NAND2_4007 ( P2_U3455 , P2_U5629 , P2_U5628 );
nand NAND2_4008 ( P2_U3456 , P2_U5631 , P2_U5630 );
nand NAND2_4009 ( P2_U3457 , P2_U5633 , P2_U5632 );
nand NAND2_4010 ( P2_U3458 , P2_U5635 , P2_U5634 );
nand NAND2_4011 ( P2_U3459 , P2_U5639 , P2_U5638 );
nand NAND2_4012 ( P2_U3460 , P2_U5641 , P2_U5640 );
nand NAND2_4013 ( P2_U3461 , P2_U5643 , P2_U5642 );
nand NAND2_4014 ( P2_U3462 , P2_U5645 , P2_U5644 );
nand NAND2_4015 ( P2_U3463 , P2_U5647 , P2_U5646 );
nand NAND2_4016 ( P2_U3464 , P2_U5649 , P2_U5648 );
nand NAND2_4017 ( P2_U3465 , P2_U5651 , P2_U5650 );
nand NAND2_4018 ( P2_U3466 , P2_U5653 , P2_U5652 );
nand NAND2_4019 ( P2_U3467 , P2_U5655 , P2_U5654 );
nand NAND2_4020 ( P2_U3468 , P2_U5657 , P2_U5656 );
nand NAND2_4021 ( P2_U3469 , P2_U5659 , P2_U5658 );
nand NAND2_4022 ( P2_U3470 , P2_U5661 , P2_U5660 );
nand NAND2_4023 ( P2_U3471 , P2_U5663 , P2_U5662 );
nand NAND2_4024 ( P2_U3472 , P2_U5665 , P2_U5664 );
nand NAND2_4025 ( P2_U3473 , P2_U5667 , P2_U5666 );
nand NAND2_4026 ( P2_U3474 , P2_U5669 , P2_U5668 );
nand NAND2_4027 ( P2_U3475 , P2_U5671 , P2_U5670 );
nand NAND2_4028 ( P2_U3476 , P2_U5673 , P2_U5672 );
nand NAND2_4029 ( P2_U3477 , P2_U5675 , P2_U5674 );
nand NAND2_4030 ( P2_U3478 , P2_U5677 , P2_U5676 );
nand NAND2_4031 ( P2_U3479 , P2_U5679 , P2_U5678 );
nand NAND2_4032 ( P2_U3480 , P2_U5681 , P2_U5680 );
nand NAND2_4033 ( P2_U3481 , P2_U5683 , P2_U5682 );
nand NAND2_4034 ( P2_U3482 , P2_U5685 , P2_U5684 );
nand NAND2_4035 ( P2_U3483 , P2_U5687 , P2_U5686 );
nand NAND2_4036 ( P2_U3484 , P2_U5689 , P2_U5688 );
nand NAND2_4037 ( P2_U3485 , P2_U5691 , P2_U5690 );
nand NAND2_4038 ( P2_U3486 , P2_U5693 , P2_U5692 );
nand NAND2_4039 ( P2_U3487 , P2_U5695 , P2_U5694 );
nand NAND2_4040 ( P2_U3488 , P2_U5697 , P2_U5696 );
nand NAND2_4041 ( P2_U3489 , P2_U5699 , P2_U5698 );
nand NAND2_4042 ( P2_U3490 , P2_U5701 , P2_U5700 );
nand NAND2_4043 ( P2_U3491 , P2_U5766 , P2_U5765 );
nand NAND2_4044 ( P2_U3492 , P2_U5768 , P2_U5767 );
nand NAND2_4045 ( P2_U3493 , P2_U5770 , P2_U5769 );
nand NAND2_4046 ( P2_U3494 , P2_U5772 , P2_U5771 );
nand NAND2_4047 ( P2_U3495 , P2_U5774 , P2_U5773 );
nand NAND2_4048 ( P2_U3496 , P2_U5776 , P2_U5775 );
nand NAND2_4049 ( P2_U3497 , P2_U5778 , P2_U5777 );
nand NAND2_4050 ( P2_U3498 , P2_U5780 , P2_U5779 );
nand NAND2_4051 ( P2_U3499 , P2_U5782 , P2_U5781 );
nand NAND2_4052 ( P2_U3500 , P2_U5784 , P2_U5783 );
nand NAND2_4053 ( P2_U3501 , P2_U5786 , P2_U5785 );
nand NAND2_4054 ( P2_U3502 , P2_U5788 , P2_U5787 );
nand NAND2_4055 ( P2_U3503 , P2_U5790 , P2_U5789 );
nand NAND2_4056 ( P2_U3504 , P2_U5792 , P2_U5791 );
nand NAND2_4057 ( P2_U3505 , P2_U5794 , P2_U5793 );
nand NAND2_4058 ( P2_U3506 , P2_U5796 , P2_U5795 );
nand NAND2_4059 ( P2_U3507 , P2_U5798 , P2_U5797 );
nand NAND2_4060 ( P2_U3508 , P2_U5800 , P2_U5799 );
nand NAND2_4061 ( P2_U3509 , P2_U5802 , P2_U5801 );
nand NAND2_4062 ( P2_U3510 , P2_U5804 , P2_U5803 );
nand NAND2_4063 ( P2_U3511 , P2_U5806 , P2_U5805 );
nand NAND2_4064 ( P2_U3512 , P2_U5808 , P2_U5807 );
nand NAND2_4065 ( P2_U3513 , P2_U5810 , P2_U5809 );
nand NAND2_4066 ( P2_U3514 , P2_U5812 , P2_U5811 );
nand NAND2_4067 ( P2_U3515 , P2_U5814 , P2_U5813 );
nand NAND2_4068 ( P2_U3516 , P2_U5816 , P2_U5815 );
nand NAND2_4069 ( P2_U3517 , P2_U5818 , P2_U5817 );
nand NAND2_4070 ( P2_U3518 , P2_U5820 , P2_U5819 );
nand NAND2_4071 ( P2_U3519 , P2_U5822 , P2_U5821 );
nand NAND2_4072 ( P2_U3520 , P2_U5824 , P2_U5823 );
nand NAND2_4073 ( P2_U3521 , P2_U5826 , P2_U5825 );
nand NAND2_4074 ( P2_U3522 , P2_U5828 , P2_U5827 );
nand NAND2_4075 ( P2_U3523 , P2_U5942 , P2_U5941 );
nand NAND2_4076 ( P2_U3524 , P2_U5944 , P2_U5943 );
nand NAND2_4077 ( P2_U3525 , P2_U5946 , P2_U5945 );
nand NAND2_4078 ( P2_U3526 , P2_U5948 , P2_U5947 );
nand NAND2_4079 ( P2_U3527 , P2_U5950 , P2_U5949 );
nand NAND2_4080 ( P2_U3528 , P2_U5952 , P2_U5951 );
nand NAND2_4081 ( P2_U3529 , P2_U5954 , P2_U5953 );
nand NAND2_4082 ( P2_U3530 , P2_U5956 , P2_U5955 );
nand NAND2_4083 ( P2_U3531 , P2_U5958 , P2_U5957 );
nand NAND2_4084 ( P2_U3532 , P2_U5960 , P2_U5959 );
nand NAND2_4085 ( P2_U3533 , P2_U5962 , P2_U5961 );
nand NAND2_4086 ( P2_U3534 , P2_U5964 , P2_U5963 );
nand NAND2_4087 ( P2_U3535 , P2_U5966 , P2_U5965 );
nand NAND2_4088 ( P2_U3536 , P2_U5968 , P2_U5967 );
nand NAND2_4089 ( P2_U3537 , P2_U5970 , P2_U5969 );
nand NAND2_4090 ( P2_U3538 , P2_U5972 , P2_U5971 );
nand NAND2_4091 ( P2_U3539 , P2_U5974 , P2_U5973 );
nand NAND2_4092 ( P2_U3540 , P2_U5976 , P2_U5975 );
nand NAND2_4093 ( P2_U3541 , P2_U5978 , P2_U5977 );
nand NAND2_4094 ( P2_U3542 , P2_U5980 , P2_U5979 );
nand NAND2_4095 ( P2_U3543 , P2_U5982 , P2_U5981 );
nand NAND2_4096 ( P2_U3544 , P2_U5984 , P2_U5983 );
nand NAND2_4097 ( P2_U3545 , P2_U5986 , P2_U5985 );
nand NAND2_4098 ( P2_U3546 , P2_U5988 , P2_U5987 );
nand NAND2_4099 ( P2_U3547 , P2_U5990 , P2_U5989 );
nand NAND2_4100 ( P2_U3548 , P2_U5992 , P2_U5991 );
nand NAND2_4101 ( P2_U3549 , P2_U5994 , P2_U5993 );
nand NAND2_4102 ( P2_U3550 , P2_U5996 , P2_U5995 );
nand NAND2_4103 ( P2_U3551 , P2_U5998 , P2_U5997 );
nand NAND2_4104 ( P2_U3552 , P2_U6000 , P2_U5999 );
nand NAND2_4105 ( P2_U3553 , P2_U6002 , P2_U6001 );
nand NAND2_4106 ( P2_U3554 , P2_U6004 , P2_U6003 );
nand NAND2_4107 ( P2_U3555 , P2_U6006 , P2_U6005 );
nand NAND2_4108 ( P2_U3556 , P2_U6008 , P2_U6007 );
nand NAND2_4109 ( P2_U3557 , P2_U6010 , P2_U6009 );
nand NAND2_4110 ( P2_U3558 , P2_U6012 , P2_U6011 );
nand NAND2_4111 ( P2_U3559 , P2_U6014 , P2_U6013 );
nand NAND2_4112 ( P2_U3560 , P2_U6016 , P2_U6015 );
nand NAND2_4113 ( P2_U3561 , P2_U6018 , P2_U6017 );
nand NAND2_4114 ( P2_U3562 , P2_U6020 , P2_U6019 );
nand NAND2_4115 ( P2_U3563 , P2_U6022 , P2_U6021 );
nand NAND2_4116 ( P2_U3564 , P2_U6024 , P2_U6023 );
nand NAND2_4117 ( P2_U3565 , P2_U6026 , P2_U6025 );
nand NAND2_4118 ( P2_U3566 , P2_U6028 , P2_U6027 );
nand NAND2_4119 ( P2_U3567 , P2_U6030 , P2_U6029 );
nand NAND2_4120 ( P2_U3568 , P2_U6032 , P2_U6031 );
nand NAND2_4121 ( P2_U3569 , P2_U6034 , P2_U6033 );
nand NAND2_4122 ( P2_U3570 , P2_U6036 , P2_U6035 );
nand NAND2_4123 ( P2_U3571 , P2_U6038 , P2_U6037 );
nand NAND2_4124 ( P2_U3572 , P2_U6040 , P2_U6039 );
nand NAND2_4125 ( P2_U3573 , P2_U6042 , P2_U6041 );
nand NAND2_4126 ( P2_U3574 , P2_U6044 , P2_U6043 );
and AND2_4127 ( P2_U3575 , P2_U4062 , P2_U4061 );
and AND2_4128 ( P2_U3576 , P2_U4064 , P2_U4063 );
and AND3_4129 ( P2_U3577 , P2_U4072 , P2_U4070 , P2_U4071 );
and AND4_4130 ( P2_U3578 , P2_U4021 , P2_U4020 , P2_U4019 , P2_U4018 );
and AND4_4131 ( P2_U3579 , P2_U4025 , P2_U4024 , P2_U4023 , P2_U4022 );
and AND4_4132 ( P2_U3580 , P2_U4029 , P2_U4028 , P2_U4027 , P2_U4026 );
and AND3_4133 ( P2_U3581 , P2_U4031 , P2_U4030 , P2_U4032 );
and AND4_4134 ( P2_U3582 , P2_U3581 , P2_U3580 , P2_U3579 , P2_U3578 );
and AND4_4135 ( P2_U3583 , P2_U4036 , P2_U4035 , P2_U4034 , P2_U4033 );
and AND4_4136 ( P2_U3584 , P2_U4040 , P2_U4039 , P2_U4038 , P2_U4037 );
and AND4_4137 ( P2_U3585 , P2_U4044 , P2_U4043 , P2_U4042 , P2_U4041 );
and AND3_4138 ( P2_U3586 , P2_U4046 , P2_U4045 , P2_U4047 );
and AND4_4139 ( P2_U3587 , P2_U3586 , P2_U3585 , P2_U3584 , P2_U3583 );
and AND2_4140 ( P2_U3588 , P2_U3389 , P2_U3388 );
and AND2_4141 ( P2_U3589 , P2_U5475 , P2_U5472 );
and AND2_4142 ( P2_U3590 , P2_U4089 , P2_U4088 );
and AND2_4143 ( P2_U3591 , P2_U4091 , P2_U4090 );
and AND3_4144 ( P2_U3592 , P2_U4093 , P2_U4092 , P2_U3591 );
and AND3_4145 ( P2_U3593 , P2_U4096 , P2_U4097 , P2_U4095 );
and AND2_4146 ( P2_U3594 , P2_U4107 , P2_U4106 );
and AND2_4147 ( P2_U3595 , P2_U4109 , P2_U4108 );
and AND3_4148 ( P2_U3596 , P2_U4111 , P2_U4110 , P2_U3595 );
and AND3_4149 ( P2_U3597 , P2_U4114 , P2_U4115 , P2_U4113 );
and AND2_4150 ( P2_U3598 , P2_U4125 , P2_U4124 );
and AND2_4151 ( P2_U3599 , P2_U4127 , P2_U4126 );
and AND3_4152 ( P2_U3600 , P2_U4129 , P2_U4128 , P2_U3599 );
and AND3_4153 ( P2_U3601 , P2_U4132 , P2_U4133 , P2_U4131 );
and AND2_4154 ( P2_U3602 , P2_U4143 , P2_U4142 );
and AND2_4155 ( P2_U3603 , P2_U4145 , P2_U4144 );
and AND3_4156 ( P2_U3604 , P2_U4147 , P2_U4146 , P2_U3603 );
and AND3_4157 ( P2_U3605 , P2_U4150 , P2_U4151 , P2_U4149 );
and AND2_4158 ( P2_U3606 , P2_U4161 , P2_U4160 );
and AND2_4159 ( P2_U3607 , P2_U4163 , P2_U4162 );
and AND3_4160 ( P2_U3608 , P2_U4165 , P2_U4164 , P2_U3607 );
and AND3_4161 ( P2_U3609 , P2_U4168 , P2_U4169 , P2_U4167 );
and AND2_4162 ( P2_U3610 , P2_U4179 , P2_U4178 );
and AND2_4163 ( P2_U3611 , P2_U4181 , P2_U4180 );
and AND3_4164 ( P2_U3612 , P2_U4183 , P2_U4182 , P2_U3611 );
and AND3_4165 ( P2_U3613 , P2_U4186 , P2_U4187 , P2_U4185 );
and AND2_4166 ( P2_U3614 , P2_U4197 , P2_U4196 );
and AND2_4167 ( P2_U3615 , P2_U4199 , P2_U4198 );
and AND3_4168 ( P2_U3616 , P2_U4201 , P2_U4200 , P2_U3615 );
and AND3_4169 ( P2_U3617 , P2_U4204 , P2_U4205 , P2_U4203 );
and AND2_4170 ( P2_U3618 , P2_U4217 , P2_U4216 );
and AND3_4171 ( P2_U3619 , P2_U4219 , P2_U4218 , P2_U3618 );
and AND3_4172 ( P2_U3620 , P2_U4222 , P2_U4223 , P2_U4221 );
and AND2_4173 ( P2_U3621 , P2_U4235 , P2_U4234 );
and AND3_4174 ( P2_U3622 , P2_U4237 , P2_U4236 , P2_U3621 );
and AND3_4175 ( P2_U3623 , P2_U4240 , P2_U4241 , P2_U4239 );
and AND2_4176 ( P2_U3624 , P2_U4253 , P2_U4252 );
and AND3_4177 ( P2_U3625 , P2_U4255 , P2_U4254 , P2_U3624 );
and AND3_4178 ( P2_U3626 , P2_U4258 , P2_U4259 , P2_U4257 );
and AND2_4179 ( P2_U3627 , P2_U4271 , P2_U4270 );
and AND3_4180 ( P2_U3628 , P2_U4273 , P2_U4272 , P2_U3627 );
and AND3_4181 ( P2_U3629 , P2_U4276 , P2_U4277 , P2_U4275 );
and AND2_4182 ( P2_U3630 , P2_U4287 , P2_U4286 );
and AND2_4183 ( P2_U3631 , P2_U4289 , P2_U4288 );
and AND3_4184 ( P2_U3632 , P2_U4291 , P2_U4290 , P2_U3631 );
and AND3_4185 ( P2_U3633 , P2_U4294 , P2_U4295 , P2_U4293 );
and AND2_4186 ( P2_U3634 , P2_U4305 , P2_U4304 );
and AND2_4187 ( P2_U3635 , P2_U4307 , P2_U4306 );
and AND3_4188 ( P2_U3636 , P2_U4309 , P2_U4308 , P2_U3635 );
and AND3_4189 ( P2_U3637 , P2_U4312 , P2_U4313 , P2_U4311 );
and AND2_4190 ( P2_U3638 , P2_U4325 , P2_U4324 );
and AND3_4191 ( P2_U3639 , P2_U4327 , P2_U4326 , P2_U3638 );
and AND3_4192 ( P2_U3640 , P2_U4330 , P2_U4331 , P2_U4329 );
and AND2_4193 ( P2_U3641 , P2_U4343 , P2_U4342 );
and AND3_4194 ( P2_U3642 , P2_U4345 , P2_U4344 , P2_U3641 );
and AND3_4195 ( P2_U3643 , P2_U4348 , P2_U4349 , P2_U4347 );
and AND2_4196 ( P2_U3644 , P2_U4361 , P2_U4360 );
and AND3_4197 ( P2_U3645 , P2_U4363 , P2_U4362 , P2_U3644 );
and AND3_4198 ( P2_U3646 , P2_U4366 , P2_U4367 , P2_U4365 );
and AND2_4199 ( P2_U3647 , P2_U4377 , P2_U4376 );
and AND2_4200 ( P2_U3648 , P2_U4379 , P2_U4378 );
and AND3_4201 ( P2_U3649 , P2_U4381 , P2_U4380 , P2_U3648 );
and AND3_4202 ( P2_U3650 , P2_U4384 , P2_U4385 , P2_U4383 );
and AND2_4203 ( P2_U3651 , P2_U4395 , P2_U4394 );
and AND2_4204 ( P2_U3652 , P2_U4397 , P2_U4396 );
and AND3_4205 ( P2_U3653 , P2_U4399 , P2_U4398 , P2_U3652 );
and AND3_4206 ( P2_U3654 , P2_U4402 , P2_U4403 , P2_U4401 );
and AND2_4207 ( P2_U3655 , P2_U4413 , P2_U4412 );
and AND2_4208 ( P2_U3656 , P2_U4415 , P2_U4414 );
and AND3_4209 ( P2_U3657 , P2_U4417 , P2_U4416 , P2_U3656 );
and AND3_4210 ( P2_U3658 , P2_U4420 , P2_U4421 , P2_U4419 );
and AND2_4211 ( P2_U3659 , P2_U4431 , P2_U4430 );
and AND2_4212 ( P2_U3660 , P2_U4433 , P2_U4432 );
and AND3_4213 ( P2_U3661 , P2_U4435 , P2_U4434 , P2_U3660 );
and AND3_4214 ( P2_U3662 , P2_U4438 , P2_U4439 , P2_U4437 );
and AND2_4215 ( P2_U3663 , P2_U4451 , P2_U4450 );
and AND3_4216 ( P2_U3664 , P2_U4453 , P2_U4452 , P2_U3663 );
and AND3_4217 ( P2_U3665 , P2_U4456 , P2_U4457 , P2_U4455 );
and AND2_4218 ( P2_U3666 , P2_U4469 , P2_U4468 );
and AND3_4219 ( P2_U3667 , P2_U4471 , P2_U4470 , P2_U3666 );
and AND3_4220 ( P2_U3668 , P2_U4474 , P2_U4475 , P2_U4473 );
and AND2_4221 ( P2_U3669 , P2_U4487 , P2_U4486 );
and AND3_4222 ( P2_U3670 , P2_U4489 , P2_U4488 , P2_U3669 );
and AND3_4223 ( P2_U3671 , P2_U4492 , P2_U4493 , P2_U4491 );
and AND2_4224 ( P2_U3672 , P2_U4503 , P2_U4502 );
and AND2_4225 ( P2_U3673 , P2_U4505 , P2_U4504 );
and AND3_4226 ( P2_U3674 , P2_U4507 , P2_U4506 , P2_U3673 );
and AND3_4227 ( P2_U3675 , P2_U4510 , P2_U4511 , P2_U4509 );
and AND2_4228 ( P2_U3676 , P2_U4521 , P2_U4520 );
and AND2_4229 ( P2_U3677 , P2_U4523 , P2_U4522 );
and AND3_4230 ( P2_U3678 , P2_U4525 , P2_U4524 , P2_U3677 );
and AND3_4231 ( P2_U3679 , P2_U4528 , P2_U4529 , P2_U4527 );
and AND2_4232 ( P2_U3680 , P2_U4539 , P2_U4538 );
and AND2_4233 ( P2_U3681 , P2_U4541 , P2_U4540 );
and AND3_4234 ( P2_U3682 , P2_U4543 , P2_U4542 , P2_U3681 );
and AND3_4235 ( P2_U3683 , P2_U4546 , P2_U4547 , P2_U4545 );
and AND2_4236 ( P2_U3684 , P2_U4557 , P2_U4556 );
and AND2_4237 ( P2_U3685 , P2_U4559 , P2_U4558 );
and AND3_4238 ( P2_U3686 , P2_U4561 , P2_U4560 , P2_U3685 );
and AND3_4239 ( P2_U3687 , P2_U4564 , P2_U4565 , P2_U4563 );
and AND2_4240 ( P2_U3688 , P2_U4575 , P2_U4574 );
and AND2_4241 ( P2_U3689 , P2_U4577 , P2_U4576 );
and AND3_4242 ( P2_U3690 , P2_U4579 , P2_U4578 , P2_U3689 );
and AND3_4243 ( P2_U3691 , P2_U4582 , P2_U4583 , P2_U4581 );
and AND5_4244 ( P2_U3692 , P2_U4593 , P2_U4592 , P2_U4594 , P2_U4595 , P2_U4596 );
and AND2_4245 ( P2_U3693 , P2_U4598 , P2_U4597 );
and AND3_4246 ( P2_U3694 , P2_U4600 , P2_U4599 , P2_U3693 );
and AND2_4247 ( P2_U3695 , P2_U4603 , P2_U4602 );
and AND2_4248 ( P2_U3696 , P2_U5472 , P2_U3389 );
and AND2_4249 ( P2_U3697 , P2_U5475 , P2_U3388 );
and AND2_4250 ( P2_U3698 , P2_U3916 , P2_U3379 );
and AND2_4251 ( P2_U3699 , P2_U5436 , P2_STATE_REG );
and AND2_4252 ( P2_U3700 , P2_U5420 , P2_U3364 );
and AND2_4253 ( P2_U3701 , P2_U3375 , P2_STATE_REG );
and AND5_4254 ( P2_U3702 , P2_U3301 , P2_U3308 , P2_U3305 , P2_U3306 , P2_U3307 );
and AND2_4255 ( P2_U3703 , P2_U3309 , P2_U3360 );
and AND4_4256 ( P2_U3704 , P2_U4759 , P2_U4758 , P2_U4761 , P2_U3706 );
and AND2_4257 ( P2_U3705 , P2_U4764 , P2_U4762 );
and AND2_4258 ( P2_U3706 , P2_U3705 , P2_U4763 );
and AND4_4259 ( P2_U3707 , P2_U4770 , P2_U4769 , P2_U4772 , P2_U3709 );
and AND2_4260 ( P2_U3708 , P2_U4775 , P2_U4773 );
and AND2_4261 ( P2_U3709 , P2_U3708 , P2_U4774 );
and AND4_4262 ( P2_U3710 , P2_U4781 , P2_U4780 , P2_U4783 , P2_U3712 );
and AND2_4263 ( P2_U3711 , P2_U4786 , P2_U4784 );
and AND2_4264 ( P2_U3712 , P2_U3711 , P2_U4785 );
and AND4_4265 ( P2_U3713 , P2_U4792 , P2_U4791 , P2_U4794 , P2_U3715 );
and AND2_4266 ( P2_U3714 , P2_U4797 , P2_U4795 );
and AND2_4267 ( P2_U3715 , P2_U3714 , P2_U4796 );
and AND4_4268 ( P2_U3716 , P2_U4803 , P2_U4802 , P2_U4805 , P2_U3718 );
and AND2_4269 ( P2_U3717 , P2_U4808 , P2_U4806 );
and AND2_4270 ( P2_U3718 , P2_U3717 , P2_U4807 );
and AND4_4271 ( P2_U3719 , P2_U4814 , P2_U4813 , P2_U4816 , P2_U3721 );
and AND2_4272 ( P2_U3720 , P2_U4819 , P2_U4817 );
and AND2_4273 ( P2_U3721 , P2_U3720 , P2_U4818 );
and AND4_4274 ( P2_U3722 , P2_U4825 , P2_U4824 , P2_U4827 , P2_U3724 );
and AND2_4275 ( P2_U3723 , P2_U4830 , P2_U4828 );
and AND2_4276 ( P2_U3724 , P2_U3723 , P2_U4829 );
and AND4_4277 ( P2_U3725 , P2_U4836 , P2_U4835 , P2_U4838 , P2_U3727 );
and AND2_4278 ( P2_U3726 , P2_U4841 , P2_U4839 );
and AND2_4279 ( P2_U3727 , P2_U3726 , P2_U4840 );
and AND4_4280 ( P2_U3728 , P2_U4847 , P2_U4849 , P2_U4846 , P2_U3730 );
and AND2_4281 ( P2_U3729 , P2_U4852 , P2_U4850 );
and AND2_4282 ( P2_U3730 , P2_U3729 , P2_U4851 );
and AND4_4283 ( P2_U3731 , P2_U4858 , P2_U4860 , P2_U4857 , P2_U3733 );
and AND2_4284 ( P2_U3732 , P2_U4863 , P2_U4861 );
and AND2_4285 ( P2_U3733 , P2_U3732 , P2_U4862 );
and AND4_4286 ( P2_U3734 , P2_U4869 , P2_U4871 , P2_U4868 , P2_U3736 );
and AND2_4287 ( P2_U3735 , P2_U4874 , P2_U4872 );
and AND2_4288 ( P2_U3736 , P2_U3735 , P2_U4873 );
and AND2_4289 ( P2_U3737 , P2_U4880 , P2_U4879 );
and AND3_4290 ( P2_U3738 , P2_U3739 , P2_U4884 , P2_U4882 );
and AND2_4291 ( P2_U3739 , P2_U4885 , P2_U4883 );
and AND2_4292 ( P2_U3740 , P2_U4891 , P2_U4890 );
and AND3_4293 ( P2_U3741 , P2_U3742 , P2_U4895 , P2_U4893 );
and AND2_4294 ( P2_U3742 , P2_U4896 , P2_U4894 );
and AND3_4295 ( P2_U3743 , P2_U4904 , P2_U4902 , P2_U3745 );
and AND2_4296 ( P2_U3744 , P2_U4907 , P2_U4905 );
and AND2_4297 ( P2_U3745 , P2_U3744 , P2_U4906 );
and AND2_4298 ( P2_U3746 , P2_U4915 , P2_U4913 );
and AND2_4299 ( P2_U3747 , P2_U4918 , P2_U4916 );
and AND2_4300 ( P2_U3748 , P2_U3747 , P2_U4917 );
and AND3_4301 ( P2_U3749 , P2_U4924 , P2_U3751 , P2_U4923 );
and AND2_4302 ( P2_U3750 , P2_U4929 , P2_U4927 );
and AND2_4303 ( P2_U3751 , P2_U3750 , P2_U4928 );
and AND3_4304 ( P2_U3752 , P2_U4935 , P2_U3754 , P2_U4934 );
and AND2_4305 ( P2_U3753 , P2_U4940 , P2_U4938 );
and AND2_4306 ( P2_U3754 , P2_U3753 , P2_U4939 );
and AND4_4307 ( P2_U3755 , P2_U4946 , P2_U4948 , P2_U4945 , P2_U3757 );
and AND2_4308 ( P2_U3756 , P2_U4951 , P2_U4949 );
and AND2_4309 ( P2_U3757 , P2_U3756 , P2_U4950 );
and AND4_4310 ( P2_U3758 , P2_U4957 , P2_U4956 , P2_U4959 , P2_U3760 );
and AND2_4311 ( P2_U3759 , P2_U4962 , P2_U4960 );
and AND2_4312 ( P2_U3760 , P2_U3759 , P2_U4961 );
and AND4_4313 ( P2_U3761 , P2_U4968 , P2_U4967 , P2_U4970 , P2_U3763 );
and AND2_4314 ( P2_U3762 , P2_U4973 , P2_U4971 );
and AND2_4315 ( P2_U3763 , P2_U3762 , P2_U4972 );
and AND2_4316 ( P2_U3764 , P2_U5464 , P2_U3383 );
nand NAND2_4317 ( P2_U3765 , P2_U5830 , P2_U5829 );
and AND2_4318 ( P2_U3766 , P2_U5911 , P2_U5908 );
and AND4_4319 ( P2_U3767 , P2_U3769 , P2_U3768 , P2_U3766 , P2_U5893 );
and AND2_4320 ( P2_U3768 , P2_U5899 , P2_U5896 );
and AND2_4321 ( P2_U3769 , P2_U5905 , P2_U5902 );
and AND3_4322 ( P2_U3770 , P2_U5878 , P2_U5875 , P2_U5872 );
and AND4_4323 ( P2_U3771 , P2_U5887 , P2_U5884 , P2_U5881 , P2_U5890 );
and AND3_4324 ( P2_U3772 , P2_U3771 , P2_U3770 , P2_U5869 );
and AND4_4325 ( P2_U3773 , P2_U5863 , P2_U5860 , P2_U5857 , P2_U5854 );
and AND2_4326 ( P2_U3774 , P2_U5851 , P2_U5848 );
and AND4_4327 ( P2_U3775 , P2_U5926 , P2_U5923 , P2_U5920 , P2_U5917 );
and AND3_4328 ( P2_U3776 , P2_U5839 , P2_U5836 , P2_U5842 );
and AND5_4329 ( P2_U3777 , P2_U3773 , P2_U3774 , P2_U5866 , P2_U5845 , P2_U3776 );
and AND5_4330 ( P2_U3778 , P2_U3767 , P2_U3772 , P2_U5914 , P2_U3775 , P2_U5929 );
and AND3_4331 ( P2_U3779 , P2_U4977 , P2_U3866 , P2_U4976 );
and AND2_4332 ( P2_U3780 , P2_U5412 , P2_U5411 );
and AND4_4333 ( P2_U3781 , P2_U5436 , P2_U3362 , P2_U4986 , P2_U3876 );
and AND2_4334 ( P2_U3782 , P2_U4994 , P2_U4993 );
and AND2_4335 ( P2_U3783 , P2_U5007 , P2_U5006 );
and AND2_4336 ( P2_U3784 , P2_U5016 , P2_U5015 );
and AND2_4337 ( P2_U3785 , P2_U5025 , P2_U5024 );
and AND2_4338 ( P2_U3786 , P2_U5032 , P2_U5030 );
and AND2_4339 ( P2_U3787 , P2_U5034 , P2_U5033 );
and AND2_4340 ( P2_U3788 , P2_U5043 , P2_U5042 );
and AND2_4341 ( P2_U3789 , P2_U5052 , P2_U5051 );
and AND2_4342 ( P2_U3790 , P2_U5061 , P2_U5060 );
and AND2_4343 ( P2_U3791 , P2_U5070 , P2_U5069 );
and AND2_4344 ( P2_U3792 , P2_U3031 , P2_U3077 );
and AND2_4345 ( P2_U3793 , P2_U5074 , P2_U5073 );
and AND3_4346 ( P2_U3794 , P2_U5077 , P2_U5076 , P2_U3793 );
and AND2_4347 ( P2_U3795 , P2_U5086 , P2_U5085 );
and AND2_4348 ( P2_U3796 , P2_U5093 , P2_U5091 );
and AND2_4349 ( P2_U3797 , P2_U5095 , P2_U5094 );
and AND2_4350 ( P2_U3798 , P2_U5104 , P2_U5103 );
and AND2_4351 ( P2_U3799 , P2_U5113 , P2_U5112 );
and AND2_4352 ( P2_U3800 , P2_U5122 , P2_U5121 );
and AND2_4353 ( P2_U3801 , P2_U5131 , P2_U5130 );
and AND2_4354 ( P2_U3802 , P2_U5140 , P2_U5139 );
and AND2_4355 ( P2_U3803 , P2_U5149 , P2_U5148 );
and AND2_4356 ( P2_U3804 , P2_U5158 , P2_U5157 );
and AND2_4357 ( P2_U3805 , P2_U5165 , P2_U5163 );
and AND2_4358 ( P2_U3806 , P2_U5167 , P2_U5166 );
and AND2_4359 ( P2_U3807 , P2_U5176 , P2_U5175 );
and AND2_4360 ( P2_U3808 , P2_U5185 , P2_U5184 );
and AND2_4361 ( P2_U3809 , P2_U5194 , P2_U5193 );
and AND2_4362 ( P2_U3810 , P2_U5201 , P2_U5199 );
and AND2_4363 ( P2_U3811 , P2_U5203 , P2_U5202 );
and AND2_4364 ( P2_U3812 , P2_U5212 , P2_U5211 );
and AND2_4365 ( P2_U3813 , P2_U5221 , P2_U5220 );
and AND2_4366 ( P2_U3814 , P2_U5230 , P2_U5229 );
and AND2_4367 ( P2_U3815 , P2_U5239 , P2_U5238 );
and AND2_4368 ( P2_U3816 , P2_U5248 , P2_U5247 );
and AND2_4369 ( P2_U3817 , P2_U5250 , P2_STATE_REG );
and AND2_4370 ( P2_U3818 , P2_U5436 , P2_U3385 );
and AND2_4371 ( P2_U3819 , P2_U3385 , P2_U3375 );
and AND3_4372 ( P2_U3820 , P2_U3871 , P2_U3312 , P2_U3302 );
and AND3_4373 ( P2_U3821 , P2_U3357 , P2_U3873 , P2_U3310 );
and AND2_4374 ( P2_U3822 , P2_U3375 , P2_U5264 );
and AND2_4375 ( P2_U3823 , P2_U3375 , P2_U5270 );
and AND2_4376 ( P2_U3824 , P2_U3375 , P2_U5292 );
and AND2_4377 ( P2_U3825 , P2_U3375 , P2_U5314 );
and AND2_4378 ( P2_U3826 , P2_U3375 , P2_U5316 );
not NOT1_4379 ( P2_U3827 , P2_IR_REG_31_ );
nand NAND2_4380 ( P2_U3828 , P2_U3023 , P2_U3300 );
nand NAND2_4381 ( P2_U3829 , P2_U5464 , P2_U5461 );
nand NAND2_4382 ( P2_U3830 , P2_U5452 , P2_U5443 );
nand NAND2_4383 ( P2_U3831 , P2_U3023 , P2_U4054 );
nand NAND2_4384 ( P2_U3832 , P2_U3023 , P2_U4618 );
and AND2_4385 ( P2_U3833 , P2_U5703 , P2_U5702 );
and AND2_4386 ( P2_U3834 , P2_U5705 , P2_U5704 );
and AND2_4387 ( P2_U3835 , P2_U5707 , P2_U5706 );
and AND2_4388 ( P2_U3836 , P2_U5709 , P2_U5708 );
and AND2_4389 ( P2_U3837 , P2_U5711 , P2_U5710 );
and AND2_4390 ( P2_U3838 , P2_U5713 , P2_U5712 );
and AND2_4391 ( P2_U3839 , P2_U5715 , P2_U5714 );
and AND2_4392 ( P2_U3840 , P2_U5717 , P2_U5716 );
and AND2_4393 ( P2_U3841 , P2_U5719 , P2_U5718 );
and AND2_4394 ( P2_U3842 , P2_U5721 , P2_U5720 );
and AND2_4395 ( P2_U3843 , P2_U5723 , P2_U5722 );
and AND2_4396 ( P2_U3844 , P2_U5725 , P2_U5724 );
and AND2_4397 ( P2_U3845 , P2_U5727 , P2_U5726 );
and AND2_4398 ( P2_U3846 , P2_U5729 , P2_U5728 );
and AND2_4399 ( P2_U3847 , P2_U5731 , P2_U5730 );
and AND2_4400 ( P2_U3848 , P2_U5733 , P2_U5732 );
and AND2_4401 ( P2_U3849 , P2_U5735 , P2_U5734 );
and AND2_4402 ( P2_U3850 , P2_U5737 , P2_U5736 );
and AND2_4403 ( P2_U3851 , P2_U5739 , P2_U5738 );
and AND2_4404 ( P2_U3852 , P2_U5741 , P2_U5740 );
and AND2_4405 ( P2_U3853 , P2_U5743 , P2_U5742 );
and AND2_4406 ( P2_U3854 , P2_U5745 , P2_U5744 );
and AND2_4407 ( P2_U3855 , P2_U5747 , P2_U5746 );
and AND2_4408 ( P2_U3856 , P2_U5749 , P2_U5748 );
and AND2_4409 ( P2_U3857 , P2_U5751 , P2_U5750 );
and AND2_4410 ( P2_U3858 , P2_U5753 , P2_U5752 );
and AND2_4411 ( P2_U3859 , P2_U5755 , P2_U5754 );
and AND2_4412 ( P2_U3860 , P2_U5757 , P2_U5756 );
and AND2_4413 ( P2_U3861 , P2_U5759 , P2_U5758 );
and AND2_4414 ( P2_U3862 , P2_U5761 , P2_U5760 );
not NOT1_4415 ( P2_U3863 , P2_R1269_U22 );
nand NAND2_4416 ( P2_U3864 , P2_U3778 , P2_U3777 );
not NOT1_4417 ( P2_U3865 , P2_R693_U14 );
and AND2_4418 ( P2_U3866 , P2_U5936 , P2_U5935 );
not NOT1_4419 ( P2_U3867 , P2_R1297_U6 );
not NOT1_4420 ( P2_U3868 , P2_U3356 );
not NOT1_4421 ( P2_U3869 , P2_U3355 );
not NOT1_4422 ( P2_U3870 , P2_U3312 );
nand NAND2_4423 ( P2_U3871 , P2_U3015 , P2_U3385 );
not NOT1_4424 ( P2_U3872 , P2_U3302 );
nand NAND2_4425 ( P2_U3873 , P2_U3016 , P2_U5452 );
not NOT1_4426 ( P2_U3874 , P2_U3310 );
not NOT1_4427 ( P2_U3875 , P2_U3357 );
nand NAND2_4428 ( P2_U3876 , P2_U3014 , P2_U3385 );
not NOT1_4429 ( P2_U3877 , P2_U3308 );
not NOT1_4430 ( P2_U3878 , P2_U3301 );
not NOT1_4431 ( P2_U3879 , P2_U3305 );
not NOT1_4432 ( P2_U3880 , P2_U3307 );
not NOT1_4433 ( P2_U3881 , P2_U3306 );
not NOT1_4434 ( P2_U3882 , P2_U3360 );
not NOT1_4435 ( P2_U3883 , P2_U3311 );
nand NAND2_4436 ( P2_U3884 , P2_U3874 , P2_U3378 );
not NOT1_4437 ( P2_U3885 , P2_U3369 );
not NOT1_4438 ( P2_U3886 , P2_U3367 );
not NOT1_4439 ( P2_U3887 , P2_U3309 );
not NOT1_4440 ( P2_U3888 , P2_U3352 );
not NOT1_4441 ( P2_U3889 , P2_U3829 );
not NOT1_4442 ( P2_U3890 , P2_U3303 );
not NOT1_4443 ( P2_U3891 , P2_U3304 );
nand NAND2_4444 ( P2_U3892 , P2_U5461 , P2_U3384 );
not NOT1_4445 ( P2_U3893 , P2_U3363 );
not NOT1_4446 ( P2_U3894 , P2_U3364 );
not NOT1_4447 ( P2_U3895 , P2_U3350 );
not NOT1_4448 ( P2_U3896 , P2_U3348 );
not NOT1_4449 ( P2_U3897 , P2_U3346 );
not NOT1_4450 ( P2_U3898 , P2_U3344 );
not NOT1_4451 ( P2_U3899 , P2_U3342 );
not NOT1_4452 ( P2_U3900 , P2_U3340 );
not NOT1_4453 ( P2_U3901 , P2_U3338 );
not NOT1_4454 ( P2_U3902 , P2_U3336 );
not NOT1_4455 ( P2_U3903 , P2_U3334 );
not NOT1_4456 ( P2_U3904 , P2_U3353 );
not NOT1_4457 ( P2_U3905 , P2_U3368 );
not NOT1_4458 ( P2_U3906 , P2_U3362 );
not NOT1_4459 ( P2_U3907 , P2_U3313 );
not NOT1_4460 ( P2_U3908 , P2_U3358 );
not NOT1_4461 ( P2_U3909 , P2_U3832 );
not NOT1_4462 ( P2_U3910 , P2_U3831 );
not NOT1_4463 ( P2_U3911 , P2_U3828 );
not NOT1_4464 ( P2_U3912 , P2_U3361 );
nand NAND2_4465 ( P2_U3913 , P2_U3370 , P2_STATE_REG );
nand NAND2_4466 ( P2_U3914 , P2_U3882 , P2_U3023 );
not NOT1_4467 ( P2_U3915 , P2_U3299 );
not NOT1_4468 ( P2_U3916 , P2_U3359 );
not NOT1_4469 ( P2_U3917 , P2_U3297 );
nand NAND2_4470 ( P2_U3918 , U56 , P2_U3151 );
nand NAND2_4471 ( P2_U3919 , P2_IR_REG_0_ , P2_U3027 );
nand NAND2_4472 ( P2_U3920 , P2_IR_REG_0_ , P2_U3917 );
nand NAND2_4473 ( P2_U3921 , U45 , P2_U3151 );
nand NAND2_4474 ( P2_U3922 , P2_SUB_594_U53 , P2_U3027 );
nand NAND2_4475 ( P2_U3923 , P2_IR_REG_1_ , P2_U3917 );
nand NAND2_4476 ( P2_U3924 , U34 , P2_U3151 );
nand NAND2_4477 ( P2_U3925 , P2_SUB_594_U23 , P2_U3027 );
nand NAND2_4478 ( P2_U3926 , P2_IR_REG_2_ , P2_U3917 );
nand NAND2_4479 ( P2_U3927 , U31 , P2_U3151 );
nand NAND2_4480 ( P2_U3928 , P2_SUB_594_U24 , P2_U3027 );
nand NAND2_4481 ( P2_U3929 , P2_IR_REG_3_ , P2_U3917 );
nand NAND2_4482 ( P2_U3930 , U30 , P2_U3151 );
nand NAND2_4483 ( P2_U3931 , P2_SUB_594_U25 , P2_U3027 );
nand NAND2_4484 ( P2_U3932 , P2_IR_REG_4_ , P2_U3917 );
nand NAND2_4485 ( P2_U3933 , U29 , P2_U3151 );
nand NAND2_4486 ( P2_U3934 , P2_SUB_594_U72 , P2_U3027 );
nand NAND2_4487 ( P2_U3935 , P2_IR_REG_5_ , P2_U3917 );
nand NAND2_4488 ( P2_U3936 , U28 , P2_U3151 );
nand NAND2_4489 ( P2_U3937 , P2_SUB_594_U26 , P2_U3027 );
nand NAND2_4490 ( P2_U3938 , P2_IR_REG_6_ , P2_U3917 );
nand NAND2_4491 ( P2_U3939 , U27 , P2_U3151 );
nand NAND2_4492 ( P2_U3940 , P2_SUB_594_U27 , P2_U3027 );
nand NAND2_4493 ( P2_U3941 , P2_IR_REG_7_ , P2_U3917 );
nand NAND2_4494 ( P2_U3942 , U26 , P2_U3151 );
nand NAND2_4495 ( P2_U3943 , P2_SUB_594_U28 , P2_U3027 );
nand NAND2_4496 ( P2_U3944 , P2_IR_REG_8_ , P2_U3917 );
nand NAND2_4497 ( P2_U3945 , U25 , P2_U3151 );
nand NAND2_4498 ( P2_U3946 , P2_SUB_594_U70 , P2_U3027 );
nand NAND2_4499 ( P2_U3947 , P2_IR_REG_9_ , P2_U3917 );
nand NAND2_4500 ( P2_U3948 , U55 , P2_U3151 );
nand NAND2_4501 ( P2_U3949 , P2_SUB_594_U8 , P2_U3027 );
nand NAND2_4502 ( P2_U3950 , P2_IR_REG_10_ , P2_U3917 );
nand NAND2_4503 ( P2_U3951 , U54 , P2_U3151 );
nand NAND2_4504 ( P2_U3952 , P2_SUB_594_U9 , P2_U3027 );
nand NAND2_4505 ( P2_U3953 , P2_IR_REG_11_ , P2_U3917 );
nand NAND2_4506 ( P2_U3954 , U53 , P2_U3151 );
nand NAND2_4507 ( P2_U3955 , P2_SUB_594_U10 , P2_U3027 );
nand NAND2_4508 ( P2_U3956 , P2_IR_REG_12_ , P2_U3917 );
nand NAND2_4509 ( P2_U3957 , U52 , P2_U3151 );
nand NAND2_4510 ( P2_U3958 , P2_SUB_594_U87 , P2_U3027 );
nand NAND2_4511 ( P2_U3959 , P2_IR_REG_13_ , P2_U3917 );
nand NAND2_4512 ( P2_U3960 , U51 , P2_U3151 );
nand NAND2_4513 ( P2_U3961 , P2_SUB_594_U11 , P2_U3027 );
nand NAND2_4514 ( P2_U3962 , P2_IR_REG_14_ , P2_U3917 );
nand NAND2_4515 ( P2_U3963 , U50 , P2_U3151 );
nand NAND2_4516 ( P2_U3964 , P2_SUB_594_U12 , P2_U3027 );
nand NAND2_4517 ( P2_U3965 , P2_IR_REG_15_ , P2_U3917 );
nand NAND2_4518 ( P2_U3966 , U49 , P2_U3151 );
nand NAND2_4519 ( P2_U3967 , P2_SUB_594_U13 , P2_U3027 );
nand NAND2_4520 ( P2_U3968 , P2_IR_REG_16_ , P2_U3917 );
nand NAND2_4521 ( P2_U3969 , U48 , P2_U3151 );
nand NAND2_4522 ( P2_U3970 , P2_SUB_594_U85 , P2_U3027 );
nand NAND2_4523 ( P2_U3971 , P2_IR_REG_17_ , P2_U3917 );
nand NAND2_4524 ( P2_U3972 , U47 , P2_U3151 );
nand NAND2_4525 ( P2_U3973 , P2_SUB_594_U14 , P2_U3027 );
nand NAND2_4526 ( P2_U3974 , P2_IR_REG_18_ , P2_U3917 );
nand NAND2_4527 ( P2_U3975 , U46 , P2_U3151 );
nand NAND2_4528 ( P2_U3976 , P2_SUB_594_U15 , P2_U3027 );
nand NAND2_4529 ( P2_U3977 , P2_IR_REG_19_ , P2_U3917 );
nand NAND2_4530 ( P2_U3978 , U44 , P2_U3151 );
nand NAND2_4531 ( P2_U3979 , P2_SUB_594_U16 , P2_U3027 );
nand NAND2_4532 ( P2_U3980 , P2_IR_REG_20_ , P2_U3917 );
nand NAND2_4533 ( P2_U3981 , U43 , P2_U3151 );
nand NAND2_4534 ( P2_U3982 , P2_SUB_594_U81 , P2_U3027 );
nand NAND2_4535 ( P2_U3983 , P2_IR_REG_21_ , P2_U3917 );
nand NAND2_4536 ( P2_U3984 , U42 , P2_U3151 );
nand NAND2_4537 ( P2_U3985 , P2_SUB_594_U17 , P2_U3027 );
nand NAND2_4538 ( P2_U3986 , P2_IR_REG_22_ , P2_U3917 );
nand NAND2_4539 ( P2_U3987 , U41 , P2_U3151 );
nand NAND2_4540 ( P2_U3988 , P2_SUB_594_U18 , P2_U3027 );
nand NAND2_4541 ( P2_U3989 , P2_IR_REG_23_ , P2_U3917 );
nand NAND2_4542 ( P2_U3990 , U40 , P2_U3151 );
nand NAND2_4543 ( P2_U3991 , P2_SUB_594_U19 , P2_U3027 );
nand NAND2_4544 ( P2_U3992 , P2_IR_REG_24_ , P2_U3917 );
nand NAND2_4545 ( P2_U3993 , U39 , P2_U3151 );
nand NAND2_4546 ( P2_U3994 , P2_SUB_594_U79 , P2_U3027 );
nand NAND2_4547 ( P2_U3995 , P2_IR_REG_25_ , P2_U3917 );
nand NAND2_4548 ( P2_U3996 , U38 , P2_U3151 );
nand NAND2_4549 ( P2_U3997 , P2_SUB_594_U20 , P2_U3027 );
nand NAND2_4550 ( P2_U3998 , P2_IR_REG_26_ , P2_U3917 );
nand NAND2_4551 ( P2_U3999 , U37 , P2_U3151 );
nand NAND2_4552 ( P2_U4000 , P2_SUB_594_U77 , P2_U3027 );
nand NAND2_4553 ( P2_U4001 , P2_IR_REG_27_ , P2_U3917 );
nand NAND2_4554 ( P2_U4002 , U36 , P2_U3151 );
nand NAND2_4555 ( P2_U4003 , P2_SUB_594_U21 , P2_U3027 );
nand NAND2_4556 ( P2_U4004 , P2_IR_REG_28_ , P2_U3917 );
nand NAND2_4557 ( P2_U4005 , U35 , P2_U3151 );
nand NAND2_4558 ( P2_U4006 , P2_SUB_594_U22 , P2_U3027 );
nand NAND2_4559 ( P2_U4007 , P2_IR_REG_29_ , P2_U3917 );
nand NAND2_4560 ( P2_U4008 , U33 , P2_U3151 );
nand NAND2_4561 ( P2_U4009 , P2_SUB_594_U75 , P2_U3027 );
nand NAND2_4562 ( P2_U4010 , P2_IR_REG_30_ , P2_U3917 );
nand NAND2_4563 ( P2_U4011 , U32 , P2_U3151 );
nand NAND2_4564 ( P2_U4012 , P2_SUB_594_U54 , P2_U3027 );
nand NAND2_4565 ( P2_U4013 , P2_IR_REG_31_ , P2_U3917 );
nand NAND2_4566 ( P2_U4014 , P2_U3915 , P2_U5433 );
not NOT1_4567 ( P2_U4015 , P2_U3300 );
nand NAND2_4568 ( P2_U4016 , P2_U3299 , P2_U5424 );
nand NAND2_4569 ( P2_U4017 , P2_U3299 , P2_U5427 );
nand NAND2_4570 ( P2_U4018 , P2_U4015 , P2_D_REG_10_ );
nand NAND2_4571 ( P2_U4019 , P2_U4015 , P2_D_REG_11_ );
nand NAND2_4572 ( P2_U4020 , P2_U4015 , P2_D_REG_12_ );
nand NAND2_4573 ( P2_U4021 , P2_U4015 , P2_D_REG_13_ );
nand NAND2_4574 ( P2_U4022 , P2_U4015 , P2_D_REG_14_ );
nand NAND2_4575 ( P2_U4023 , P2_U4015 , P2_D_REG_15_ );
nand NAND2_4576 ( P2_U4024 , P2_U4015 , P2_D_REG_16_ );
nand NAND2_4577 ( P2_U4025 , P2_U4015 , P2_D_REG_17_ );
nand NAND2_4578 ( P2_U4026 , P2_U4015 , P2_D_REG_18_ );
nand NAND2_4579 ( P2_U4027 , P2_U4015 , P2_D_REG_19_ );
nand NAND2_4580 ( P2_U4028 , P2_U4015 , P2_D_REG_20_ );
nand NAND2_4581 ( P2_U4029 , P2_U4015 , P2_D_REG_21_ );
nand NAND2_4582 ( P2_U4030 , P2_U4015 , P2_D_REG_22_ );
nand NAND2_4583 ( P2_U4031 , P2_U4015 , P2_D_REG_23_ );
nand NAND2_4584 ( P2_U4032 , P2_U4015 , P2_D_REG_24_ );
nand NAND2_4585 ( P2_U4033 , P2_U4015 , P2_D_REG_25_ );
nand NAND2_4586 ( P2_U4034 , P2_U4015 , P2_D_REG_26_ );
nand NAND2_4587 ( P2_U4035 , P2_U4015 , P2_D_REG_27_ );
nand NAND2_4588 ( P2_U4036 , P2_U4015 , P2_D_REG_28_ );
nand NAND2_4589 ( P2_U4037 , P2_U4015 , P2_D_REG_29_ );
nand NAND2_4590 ( P2_U4038 , P2_U4015 , P2_D_REG_2_ );
nand NAND2_4591 ( P2_U4039 , P2_U4015 , P2_D_REG_30_ );
nand NAND2_4592 ( P2_U4040 , P2_U4015 , P2_D_REG_31_ );
nand NAND2_4593 ( P2_U4041 , P2_U4015 , P2_D_REG_3_ );
nand NAND2_4594 ( P2_U4042 , P2_U4015 , P2_D_REG_4_ );
nand NAND2_4595 ( P2_U4043 , P2_U4015 , P2_D_REG_5_ );
nand NAND2_4596 ( P2_U4044 , P2_U4015 , P2_D_REG_6_ );
nand NAND2_4597 ( P2_U4045 , P2_U4015 , P2_D_REG_7_ );
nand NAND2_4598 ( P2_U4046 , P2_U4015 , P2_D_REG_8_ );
nand NAND2_4599 ( P2_U4047 , P2_U4015 , P2_D_REG_9_ );
not NOT1_4600 ( P2_U4048 , P2_U3830 );
nand NAND2_4601 ( P2_U4049 , P2_U5452 , P2_U5446 );
nand NAND2_4602 ( P2_U4050 , P2_U5478 , P2_U4049 );
nand NAND2_4603 ( P2_U4051 , P2_U3369 , P2_U3367 );
nand NAND2_4604 ( P2_U4052 , P2_U3890 , P2_U4051 );
nand NAND2_4605 ( P2_U4053 , P2_U3891 , P2_U4050 );
nand NAND2_4606 ( P2_U4054 , P2_U4053 , P2_U4052 );
nand NAND2_4607 ( P2_U4055 , P2_U3022 , P2_REG0_REG_1_ );
nand NAND2_4608 ( P2_U4056 , P2_REG1_REG_1_ , P2_U3021 );
nand NAND2_4609 ( P2_U4057 , P2_REG2_REG_1_ , P2_U3020 );
nand NAND2_4610 ( P2_U4058 , P2_REG3_REG_1_ , P2_U3019 );
not NOT1_4611 ( P2_U4059 , P2_U3077 );
nand NAND2_4612 ( P2_U4060 , P2_U3873 , P2_U3357 );
nand NAND2_4613 ( P2_U4061 , P2_U3879 , P2_R1110_U95 );
nand NAND2_4614 ( P2_U4062 , P2_U3881 , P2_R1077_U95 );
nand NAND2_4615 ( P2_U4063 , P2_U3880 , P2_R1095_U25 );
nand NAND2_4616 ( P2_U4064 , P2_U3877 , P2_R1143_U95 );
nand NAND2_4617 ( P2_U4065 , P2_U3887 , P2_R1161_U95 );
nand NAND2_4618 ( P2_U4066 , P2_U3883 , P2_R1131_U25 );
nand NAND2_4619 ( P2_U4067 , P2_U3017 , P2_R1200_U25 );
not NOT1_4620 ( P2_U4068 , P2_U3314 );
nand NAND2_4621 ( P2_U4069 , P2_U3352 , P2_U3829 );
nand NAND2_4622 ( P2_U4070 , P2_R1179_U25 , P2_U3026 );
nand NAND2_4623 ( P2_U4071 , P2_U3025 , P2_U3077 );
nand NAND2_4624 ( P2_U4072 , P2_U3387 , P2_U4060 );
nand NAND2_4625 ( P2_U4073 , P2_U3577 , P2_U4068 );
nand NAND2_4626 ( P2_U4074 , P2_REG0_REG_2_ , P2_U3022 );
nand NAND2_4627 ( P2_U4075 , P2_REG1_REG_2_ , P2_U3021 );
nand NAND2_4628 ( P2_U4076 , P2_REG2_REG_2_ , P2_U3020 );
nand NAND2_4629 ( P2_U4077 , P2_REG3_REG_2_ , P2_U3019 );
not NOT1_4630 ( P2_U4078 , P2_U3067 );
nand NAND2_4631 ( P2_U4079 , P2_REG0_REG_0_ , P2_U3022 );
nand NAND2_4632 ( P2_U4080 , P2_REG1_REG_0_ , P2_U3021 );
nand NAND2_4633 ( P2_U4081 , P2_REG2_REG_0_ , P2_U3020 );
nand NAND2_4634 ( P2_U4082 , P2_REG3_REG_0_ , P2_U3019 );
not NOT1_4635 ( P2_U4083 , P2_U3076 );
nand NAND2_4636 ( P2_U4084 , P2_U5464 , P2_U3383 );
nand NAND2_4637 ( P2_U4085 , P2_U3892 , P2_U4084 );
nand NAND2_4638 ( P2_U4086 , P2_U3033 , P2_U3076 );
nand NAND2_4639 ( P2_U4087 , P2_R1110_U94 , P2_U3879 );
nand NAND2_4640 ( P2_U4088 , P2_R1077_U94 , P2_U3881 );
nand NAND2_4641 ( P2_U4089 , P2_R1095_U102 , P2_U3880 );
nand NAND2_4642 ( P2_U4090 , P2_R1143_U94 , P2_U3877 );
nand NAND2_4643 ( P2_U4091 , P2_R1161_U94 , P2_U3887 );
nand NAND2_4644 ( P2_U4092 , P2_R1131_U102 , P2_U3883 );
nand NAND2_4645 ( P2_U4093 , P2_R1200_U102 , P2_U3017 );
not NOT1_4646 ( P2_U4094 , P2_U3315 );
nand NAND2_4647 ( P2_U4095 , P2_R1179_U102 , P2_U3026 );
nand NAND2_4648 ( P2_U4096 , P2_U3025 , P2_U3067 );
nand NAND2_4649 ( P2_U4097 , P2_U3392 , P2_U4060 );
nand NAND2_4650 ( P2_U4098 , P2_U3593 , P2_U4094 );
nand NAND2_4651 ( P2_U4099 , P2_REG0_REG_3_ , P2_U3022 );
nand NAND2_4652 ( P2_U4100 , P2_REG1_REG_3_ , P2_U3021 );
nand NAND2_4653 ( P2_U4101 , P2_REG2_REG_3_ , P2_U3020 );
nand NAND2_4654 ( P2_U4102 , P2_SUB_605_U26 , P2_U3019 );
not NOT1_4655 ( P2_U4103 , P2_U3063 );
nand NAND2_4656 ( P2_U4104 , P2_U3033 , P2_U3077 );
nand NAND2_4657 ( P2_U4105 , P2_R1110_U16 , P2_U3879 );
nand NAND2_4658 ( P2_U4106 , P2_R1077_U16 , P2_U3881 );
nand NAND2_4659 ( P2_U4107 , P2_R1095_U112 , P2_U3880 );
nand NAND2_4660 ( P2_U4108 , P2_R1143_U16 , P2_U3877 );
nand NAND2_4661 ( P2_U4109 , P2_R1161_U16 , P2_U3887 );
nand NAND2_4662 ( P2_U4110 , P2_R1131_U112 , P2_U3883 );
nand NAND2_4663 ( P2_U4111 , P2_R1200_U112 , P2_U3017 );
not NOT1_4664 ( P2_U4112 , P2_U3316 );
nand NAND2_4665 ( P2_U4113 , P2_R1179_U112 , P2_U3026 );
nand NAND2_4666 ( P2_U4114 , P2_U3025 , P2_U3063 );
nand NAND2_4667 ( P2_U4115 , P2_U3395 , P2_U4060 );
nand NAND2_4668 ( P2_U4116 , P2_U3597 , P2_U4112 );
nand NAND2_4669 ( P2_U4117 , P2_REG0_REG_4_ , P2_U3022 );
nand NAND2_4670 ( P2_U4118 , P2_REG1_REG_4_ , P2_U3021 );
nand NAND2_4671 ( P2_U4119 , P2_REG2_REG_4_ , P2_U3020 );
nand NAND2_4672 ( P2_U4120 , P2_SUB_605_U30 , P2_U3019 );
not NOT1_4673 ( P2_U4121 , P2_U3059 );
nand NAND2_4674 ( P2_U4122 , P2_U3033 , P2_U3067 );
nand NAND2_4675 ( P2_U4123 , P2_R1110_U100 , P2_U3879 );
nand NAND2_4676 ( P2_U4124 , P2_R1077_U100 , P2_U3881 );
nand NAND2_4677 ( P2_U4125 , P2_R1095_U22 , P2_U3880 );
nand NAND2_4678 ( P2_U4126 , P2_R1143_U100 , P2_U3877 );
nand NAND2_4679 ( P2_U4127 , P2_R1161_U100 , P2_U3887 );
nand NAND2_4680 ( P2_U4128 , P2_R1131_U22 , P2_U3883 );
nand NAND2_4681 ( P2_U4129 , P2_R1200_U22 , P2_U3017 );
not NOT1_4682 ( P2_U4130 , P2_U3317 );
nand NAND2_4683 ( P2_U4131 , P2_R1179_U22 , P2_U3026 );
nand NAND2_4684 ( P2_U4132 , P2_U3025 , P2_U3059 );
nand NAND2_4685 ( P2_U4133 , P2_U3398 , P2_U4060 );
nand NAND2_4686 ( P2_U4134 , P2_U3601 , P2_U4130 );
nand NAND2_4687 ( P2_U4135 , P2_REG0_REG_5_ , P2_U3022 );
nand NAND2_4688 ( P2_U4136 , P2_REG1_REG_5_ , P2_U3021 );
nand NAND2_4689 ( P2_U4137 , P2_REG2_REG_5_ , P2_U3020 );
nand NAND2_4690 ( P2_U4138 , P2_SUB_605_U22 , P2_U3019 );
not NOT1_4691 ( P2_U4139 , P2_U3066 );
nand NAND2_4692 ( P2_U4140 , P2_U3033 , P2_U3063 );
nand NAND2_4693 ( P2_U4141 , P2_R1110_U99 , P2_U3879 );
nand NAND2_4694 ( P2_U4142 , P2_R1077_U99 , P2_U3881 );
nand NAND2_4695 ( P2_U4143 , P2_R1095_U111 , P2_U3880 );
nand NAND2_4696 ( P2_U4144 , P2_R1143_U99 , P2_U3877 );
nand NAND2_4697 ( P2_U4145 , P2_R1161_U99 , P2_U3887 );
nand NAND2_4698 ( P2_U4146 , P2_R1131_U111 , P2_U3883 );
nand NAND2_4699 ( P2_U4147 , P2_R1200_U111 , P2_U3017 );
not NOT1_4700 ( P2_U4148 , P2_U3318 );
nand NAND2_4701 ( P2_U4149 , P2_R1179_U111 , P2_U3026 );
nand NAND2_4702 ( P2_U4150 , P2_U3025 , P2_U3066 );
nand NAND2_4703 ( P2_U4151 , P2_U3401 , P2_U4060 );
nand NAND2_4704 ( P2_U4152 , P2_U3605 , P2_U4148 );
nand NAND2_4705 ( P2_U4153 , P2_REG0_REG_6_ , P2_U3022 );
nand NAND2_4706 ( P2_U4154 , P2_REG1_REG_6_ , P2_U3021 );
nand NAND2_4707 ( P2_U4155 , P2_REG2_REG_6_ , P2_U3020 );
nand NAND2_4708 ( P2_U4156 , P2_SUB_605_U8 , P2_U3019 );
not NOT1_4709 ( P2_U4157 , P2_U3070 );
nand NAND2_4710 ( P2_U4158 , P2_U3033 , P2_U3059 );
nand NAND2_4711 ( P2_U4159 , P2_R1110_U17 , P2_U3879 );
nand NAND2_4712 ( P2_U4160 , P2_R1077_U17 , P2_U3881 );
nand NAND2_4713 ( P2_U4161 , P2_R1095_U110 , P2_U3880 );
nand NAND2_4714 ( P2_U4162 , P2_R1143_U17 , P2_U3877 );
nand NAND2_4715 ( P2_U4163 , P2_R1161_U17 , P2_U3887 );
nand NAND2_4716 ( P2_U4164 , P2_R1131_U110 , P2_U3883 );
nand NAND2_4717 ( P2_U4165 , P2_R1200_U110 , P2_U3017 );
not NOT1_4718 ( P2_U4166 , P2_U3319 );
nand NAND2_4719 ( P2_U4167 , P2_R1179_U110 , P2_U3026 );
nand NAND2_4720 ( P2_U4168 , P2_U3025 , P2_U3070 );
nand NAND2_4721 ( P2_U4169 , P2_U3404 , P2_U4060 );
nand NAND2_4722 ( P2_U4170 , P2_U3609 , P2_U4166 );
nand NAND2_4723 ( P2_U4171 , P2_REG0_REG_7_ , P2_U3022 );
nand NAND2_4724 ( P2_U4172 , P2_REG1_REG_7_ , P2_U3021 );
nand NAND2_4725 ( P2_U4173 , P2_REG2_REG_7_ , P2_U3020 );
nand NAND2_4726 ( P2_U4174 , P2_SUB_605_U18 , P2_U3019 );
not NOT1_4727 ( P2_U4175 , P2_U3069 );
nand NAND2_4728 ( P2_U4176 , P2_U3033 , P2_U3066 );
nand NAND2_4729 ( P2_U4177 , P2_R1110_U98 , P2_U3879 );
nand NAND2_4730 ( P2_U4178 , P2_R1077_U98 , P2_U3881 );
nand NAND2_4731 ( P2_U4179 , P2_R1095_U23 , P2_U3880 );
nand NAND2_4732 ( P2_U4180 , P2_R1143_U98 , P2_U3877 );
nand NAND2_4733 ( P2_U4181 , P2_R1161_U98 , P2_U3887 );
nand NAND2_4734 ( P2_U4182 , P2_R1131_U23 , P2_U3883 );
nand NAND2_4735 ( P2_U4183 , P2_R1200_U23 , P2_U3017 );
not NOT1_4736 ( P2_U4184 , P2_U3320 );
nand NAND2_4737 ( P2_U4185 , P2_R1179_U23 , P2_U3026 );
nand NAND2_4738 ( P2_U4186 , P2_U3025 , P2_U3069 );
nand NAND2_4739 ( P2_U4187 , P2_U3407 , P2_U4060 );
nand NAND2_4740 ( P2_U4188 , P2_U3613 , P2_U4184 );
nand NAND2_4741 ( P2_U4189 , P2_REG0_REG_8_ , P2_U3022 );
nand NAND2_4742 ( P2_U4190 , P2_REG1_REG_8_ , P2_U3021 );
nand NAND2_4743 ( P2_U4191 , P2_REG2_REG_8_ , P2_U3020 );
nand NAND2_4744 ( P2_U4192 , P2_SUB_605_U12 , P2_U3019 );
not NOT1_4745 ( P2_U4193 , P2_U3083 );
nand NAND2_4746 ( P2_U4194 , P2_U3033 , P2_U3070 );
nand NAND2_4747 ( P2_U4195 , P2_R1110_U18 , P2_U3879 );
nand NAND2_4748 ( P2_U4196 , P2_R1077_U18 , P2_U3881 );
nand NAND2_4749 ( P2_U4197 , P2_R1095_U109 , P2_U3880 );
nand NAND2_4750 ( P2_U4198 , P2_R1143_U18 , P2_U3877 );
nand NAND2_4751 ( P2_U4199 , P2_R1161_U18 , P2_U3887 );
nand NAND2_4752 ( P2_U4200 , P2_R1131_U109 , P2_U3883 );
nand NAND2_4753 ( P2_U4201 , P2_R1200_U109 , P2_U3017 );
not NOT1_4754 ( P2_U4202 , P2_U3321 );
nand NAND2_4755 ( P2_U4203 , P2_R1179_U109 , P2_U3026 );
nand NAND2_4756 ( P2_U4204 , P2_U3025 , P2_U3083 );
nand NAND2_4757 ( P2_U4205 , P2_U3410 , P2_U4060 );
nand NAND2_4758 ( P2_U4206 , P2_U3617 , P2_U4202 );
nand NAND2_4759 ( P2_U4207 , P2_REG0_REG_9_ , P2_U3022 );
nand NAND2_4760 ( P2_U4208 , P2_REG1_REG_9_ , P2_U3021 );
nand NAND2_4761 ( P2_U4209 , P2_REG2_REG_9_ , P2_U3020 );
nand NAND2_4762 ( P2_U4210 , P2_SUB_605_U14 , P2_U3019 );
not NOT1_4763 ( P2_U4211 , P2_U3082 );
nand NAND2_4764 ( P2_U4212 , P2_U3033 , P2_U3069 );
nand NAND2_4765 ( P2_U4213 , P2_R1110_U97 , P2_U3879 );
nand NAND2_4766 ( P2_U4214 , P2_R1077_U97 , P2_U3881 );
nand NAND2_4767 ( P2_U4215 , P2_R1095_U24 , P2_U3880 );
nand NAND2_4768 ( P2_U4216 , P2_R1143_U97 , P2_U3877 );
nand NAND2_4769 ( P2_U4217 , P2_R1161_U97 , P2_U3887 );
nand NAND2_4770 ( P2_U4218 , P2_R1131_U24 , P2_U3883 );
nand NAND2_4771 ( P2_U4219 , P2_R1200_U24 , P2_U3017 );
not NOT1_4772 ( P2_U4220 , P2_U3322 );
nand NAND2_4773 ( P2_U4221 , P2_R1179_U24 , P2_U3026 );
nand NAND2_4774 ( P2_U4222 , P2_U3025 , P2_U3082 );
nand NAND2_4775 ( P2_U4223 , P2_U3413 , P2_U4060 );
nand NAND2_4776 ( P2_U4224 , P2_U3620 , P2_U4220 );
nand NAND2_4777 ( P2_U4225 , P2_REG0_REG_10_ , P2_U3022 );
nand NAND2_4778 ( P2_U4226 , P2_REG1_REG_10_ , P2_U3021 );
nand NAND2_4779 ( P2_U4227 , P2_REG2_REG_10_ , P2_U3020 );
nand NAND2_4780 ( P2_U4228 , P2_SUB_605_U13 , P2_U3019 );
not NOT1_4781 ( P2_U4229 , P2_U3061 );
nand NAND2_4782 ( P2_U4230 , P2_U3033 , P2_U3083 );
nand NAND2_4783 ( P2_U4231 , P2_R1110_U96 , P2_U3879 );
nand NAND2_4784 ( P2_U4232 , P2_R1077_U96 , P2_U3881 );
nand NAND2_4785 ( P2_U4233 , P2_R1095_U108 , P2_U3880 );
nand NAND2_4786 ( P2_U4234 , P2_R1143_U96 , P2_U3877 );
nand NAND2_4787 ( P2_U4235 , P2_R1161_U96 , P2_U3887 );
nand NAND2_4788 ( P2_U4236 , P2_R1131_U108 , P2_U3883 );
nand NAND2_4789 ( P2_U4237 , P2_R1200_U108 , P2_U3017 );
not NOT1_4790 ( P2_U4238 , P2_U3323 );
nand NAND2_4791 ( P2_U4239 , P2_R1179_U108 , P2_U3026 );
nand NAND2_4792 ( P2_U4240 , P2_U3025 , P2_U3061 );
nand NAND2_4793 ( P2_U4241 , P2_U3416 , P2_U4060 );
nand NAND2_4794 ( P2_U4242 , P2_U3623 , P2_U4238 );
nand NAND2_4795 ( P2_U4243 , P2_REG0_REG_11_ , P2_U3022 );
nand NAND2_4796 ( P2_U4244 , P2_REG1_REG_11_ , P2_U3021 );
nand NAND2_4797 ( P2_U4245 , P2_REG2_REG_11_ , P2_U3020 );
nand NAND2_4798 ( P2_U4246 , P2_SUB_605_U9 , P2_U3019 );
not NOT1_4799 ( P2_U4247 , P2_U3062 );
nand NAND2_4800 ( P2_U4248 , P2_U3033 , P2_U3082 );
nand NAND2_4801 ( P2_U4249 , P2_R1110_U10 , P2_U3879 );
nand NAND2_4802 ( P2_U4250 , P2_R1077_U10 , P2_U3881 );
nand NAND2_4803 ( P2_U4251 , P2_R1095_U118 , P2_U3880 );
nand NAND2_4804 ( P2_U4252 , P2_R1143_U10 , P2_U3877 );
nand NAND2_4805 ( P2_U4253 , P2_R1161_U10 , P2_U3887 );
nand NAND2_4806 ( P2_U4254 , P2_R1131_U118 , P2_U3883 );
nand NAND2_4807 ( P2_U4255 , P2_R1200_U118 , P2_U3017 );
not NOT1_4808 ( P2_U4256 , P2_U3324 );
nand NAND2_4809 ( P2_U4257 , P2_R1179_U118 , P2_U3026 );
nand NAND2_4810 ( P2_U4258 , P2_U3025 , P2_U3062 );
nand NAND2_4811 ( P2_U4259 , P2_U3419 , P2_U4060 );
nand NAND2_4812 ( P2_U4260 , P2_U3626 , P2_U4256 );
nand NAND2_4813 ( P2_U4261 , P2_REG0_REG_12_ , P2_U3022 );
nand NAND2_4814 ( P2_U4262 , P2_REG1_REG_12_ , P2_U3021 );
nand NAND2_4815 ( P2_U4263 , P2_REG2_REG_12_ , P2_U3020 );
nand NAND2_4816 ( P2_U4264 , P2_SUB_605_U24 , P2_U3019 );
not NOT1_4817 ( P2_U4265 , P2_U3071 );
nand NAND2_4818 ( P2_U4266 , P2_U3033 , P2_U3061 );
nand NAND2_4819 ( P2_U4267 , P2_R1110_U114 , P2_U3879 );
nand NAND2_4820 ( P2_U4268 , P2_R1077_U114 , P2_U3881 );
nand NAND2_4821 ( P2_U4269 , P2_R1095_U17 , P2_U3880 );
nand NAND2_4822 ( P2_U4270 , P2_R1143_U114 , P2_U3877 );
nand NAND2_4823 ( P2_U4271 , P2_R1161_U114 , P2_U3887 );
nand NAND2_4824 ( P2_U4272 , P2_R1131_U17 , P2_U3883 );
nand NAND2_4825 ( P2_U4273 , P2_R1200_U17 , P2_U3017 );
not NOT1_4826 ( P2_U4274 , P2_U3325 );
nand NAND2_4827 ( P2_U4275 , P2_R1179_U17 , P2_U3026 );
nand NAND2_4828 ( P2_U4276 , P2_U3025 , P2_U3071 );
nand NAND2_4829 ( P2_U4277 , P2_U3422 , P2_U4060 );
nand NAND2_4830 ( P2_U4278 , P2_U3629 , P2_U4274 );
nand NAND2_4831 ( P2_U4279 , P2_REG0_REG_13_ , P2_U3022 );
nand NAND2_4832 ( P2_U4280 , P2_REG1_REG_13_ , P2_U3021 );
nand NAND2_4833 ( P2_U4281 , P2_REG2_REG_13_ , P2_U3020 );
nand NAND2_4834 ( P2_U4282 , P2_SUB_605_U25 , P2_U3019 );
not NOT1_4835 ( P2_U4283 , P2_U3079 );
nand NAND2_4836 ( P2_U4284 , P2_U3033 , P2_U3062 );
nand NAND2_4837 ( P2_U4285 , P2_R1110_U113 , P2_U3879 );
nand NAND2_4838 ( P2_U4286 , P2_R1077_U113 , P2_U3881 );
nand NAND2_4839 ( P2_U4287 , P2_R1095_U107 , P2_U3880 );
nand NAND2_4840 ( P2_U4288 , P2_R1143_U113 , P2_U3877 );
nand NAND2_4841 ( P2_U4289 , P2_R1161_U113 , P2_U3887 );
nand NAND2_4842 ( P2_U4290 , P2_R1131_U107 , P2_U3883 );
nand NAND2_4843 ( P2_U4291 , P2_R1200_U107 , P2_U3017 );
not NOT1_4844 ( P2_U4292 , P2_U3326 );
nand NAND2_4845 ( P2_U4293 , P2_R1179_U107 , P2_U3026 );
nand NAND2_4846 ( P2_U4294 , P2_U3025 , P2_U3079 );
nand NAND2_4847 ( P2_U4295 , P2_U3425 , P2_U4060 );
nand NAND2_4848 ( P2_U4296 , P2_U3633 , P2_U4292 );
nand NAND2_4849 ( P2_U4297 , P2_REG0_REG_14_ , P2_U3022 );
nand NAND2_4850 ( P2_U4298 , P2_REG1_REG_14_ , P2_U3021 );
nand NAND2_4851 ( P2_U4299 , P2_REG2_REG_14_ , P2_U3020 );
nand NAND2_4852 ( P2_U4300 , P2_SUB_605_U31 , P2_U3019 );
not NOT1_4853 ( P2_U4301 , P2_U3078 );
nand NAND2_4854 ( P2_U4302 , P2_U3033 , P2_U3071 );
nand NAND2_4855 ( P2_U4303 , P2_R1110_U11 , P2_U3879 );
nand NAND2_4856 ( P2_U4304 , P2_R1077_U11 , P2_U3881 );
nand NAND2_4857 ( P2_U4305 , P2_R1095_U106 , P2_U3880 );
nand NAND2_4858 ( P2_U4306 , P2_R1143_U11 , P2_U3877 );
nand NAND2_4859 ( P2_U4307 , P2_R1161_U11 , P2_U3887 );
nand NAND2_4860 ( P2_U4308 , P2_R1131_U106 , P2_U3883 );
nand NAND2_4861 ( P2_U4309 , P2_R1200_U106 , P2_U3017 );
not NOT1_4862 ( P2_U4310 , P2_U3327 );
nand NAND2_4863 ( P2_U4311 , P2_R1179_U106 , P2_U3026 );
nand NAND2_4864 ( P2_U4312 , P2_U3025 , P2_U3078 );
nand NAND2_4865 ( P2_U4313 , P2_U3428 , P2_U4060 );
nand NAND2_4866 ( P2_U4314 , P2_U3637 , P2_U4310 );
nand NAND2_4867 ( P2_U4315 , P2_REG0_REG_15_ , P2_U3022 );
nand NAND2_4868 ( P2_U4316 , P2_REG1_REG_15_ , P2_U3021 );
nand NAND2_4869 ( P2_U4317 , P2_REG2_REG_15_ , P2_U3020 );
nand NAND2_4870 ( P2_U4318 , P2_SUB_605_U21 , P2_U3019 );
not NOT1_4871 ( P2_U4319 , P2_U3073 );
nand NAND2_4872 ( P2_U4320 , P2_U3033 , P2_U3079 );
nand NAND2_4873 ( P2_U4321 , P2_R1110_U112 , P2_U3879 );
nand NAND2_4874 ( P2_U4322 , P2_R1077_U112 , P2_U3881 );
nand NAND2_4875 ( P2_U4323 , P2_R1095_U117 , P2_U3880 );
nand NAND2_4876 ( P2_U4324 , P2_R1143_U112 , P2_U3877 );
nand NAND2_4877 ( P2_U4325 , P2_R1161_U112 , P2_U3887 );
nand NAND2_4878 ( P2_U4326 , P2_R1131_U117 , P2_U3883 );
nand NAND2_4879 ( P2_U4327 , P2_R1200_U117 , P2_U3017 );
not NOT1_4880 ( P2_U4328 , P2_U3328 );
nand NAND2_4881 ( P2_U4329 , P2_R1179_U117 , P2_U3026 );
nand NAND2_4882 ( P2_U4330 , P2_U3025 , P2_U3073 );
nand NAND2_4883 ( P2_U4331 , P2_U3431 , P2_U4060 );
nand NAND2_4884 ( P2_U4332 , P2_U3640 , P2_U4328 );
nand NAND2_4885 ( P2_U4333 , P2_REG0_REG_16_ , P2_U3022 );
nand NAND2_4886 ( P2_U4334 , P2_REG1_REG_16_ , P2_U3021 );
nand NAND2_4887 ( P2_U4335 , P2_REG2_REG_16_ , P2_U3020 );
nand NAND2_4888 ( P2_U4336 , P2_SUB_605_U7 , P2_U3019 );
not NOT1_4889 ( P2_U4337 , P2_U3072 );
nand NAND2_4890 ( P2_U4338 , P2_U3033 , P2_U3078 );
nand NAND2_4891 ( P2_U4339 , P2_R1110_U111 , P2_U3879 );
nand NAND2_4892 ( P2_U4340 , P2_R1077_U111 , P2_U3881 );
nand NAND2_4893 ( P2_U4341 , P2_R1095_U116 , P2_U3880 );
nand NAND2_4894 ( P2_U4342 , P2_R1143_U111 , P2_U3877 );
nand NAND2_4895 ( P2_U4343 , P2_R1161_U111 , P2_U3887 );
nand NAND2_4896 ( P2_U4344 , P2_R1131_U116 , P2_U3883 );
nand NAND2_4897 ( P2_U4345 , P2_R1200_U116 , P2_U3017 );
not NOT1_4898 ( P2_U4346 , P2_U3329 );
nand NAND2_4899 ( P2_U4347 , P2_R1179_U116 , P2_U3026 );
nand NAND2_4900 ( P2_U4348 , P2_U3025 , P2_U3072 );
nand NAND2_4901 ( P2_U4349 , P2_U3434 , P2_U4060 );
nand NAND2_4902 ( P2_U4350 , P2_U3643 , P2_U4346 );
nand NAND2_4903 ( P2_U4351 , P2_REG0_REG_17_ , P2_U3022 );
nand NAND2_4904 ( P2_U4352 , P2_REG1_REG_17_ , P2_U3021 );
nand NAND2_4905 ( P2_U4353 , P2_REG2_REG_17_ , P2_U3020 );
nand NAND2_4906 ( P2_U4354 , P2_SUB_605_U19 , P2_U3019 );
not NOT1_4907 ( P2_U4355 , P2_U3068 );
nand NAND2_4908 ( P2_U4356 , P2_U3033 , P2_U3073 );
nand NAND2_4909 ( P2_U4357 , P2_R1110_U110 , P2_U3879 );
nand NAND2_4910 ( P2_U4358 , P2_R1077_U110 , P2_U3881 );
nand NAND2_4911 ( P2_U4359 , P2_R1095_U18 , P2_U3880 );
nand NAND2_4912 ( P2_U4360 , P2_R1143_U110 , P2_U3877 );
nand NAND2_4913 ( P2_U4361 , P2_R1161_U110 , P2_U3887 );
nand NAND2_4914 ( P2_U4362 , P2_R1131_U18 , P2_U3883 );
nand NAND2_4915 ( P2_U4363 , P2_R1200_U18 , P2_U3017 );
not NOT1_4916 ( P2_U4364 , P2_U3330 );
nand NAND2_4917 ( P2_U4365 , P2_R1179_U18 , P2_U3026 );
nand NAND2_4918 ( P2_U4366 , P2_U3025 , P2_U3068 );
nand NAND2_4919 ( P2_U4367 , P2_U3437 , P2_U4060 );
nand NAND2_4920 ( P2_U4368 , P2_U3646 , P2_U4364 );
nand NAND2_4921 ( P2_U4369 , P2_REG0_REG_18_ , P2_U3022 );
nand NAND2_4922 ( P2_U4370 , P2_REG1_REG_18_ , P2_U3021 );
nand NAND2_4923 ( P2_U4371 , P2_REG2_REG_18_ , P2_U3020 );
nand NAND2_4924 ( P2_U4372 , P2_SUB_605_U11 , P2_U3019 );
not NOT1_4925 ( P2_U4373 , P2_U3081 );
nand NAND2_4926 ( P2_U4374 , P2_U3033 , P2_U3072 );
nand NAND2_4927 ( P2_U4375 , P2_R1110_U12 , P2_U3879 );
nand NAND2_4928 ( P2_U4376 , P2_R1077_U12 , P2_U3881 );
nand NAND2_4929 ( P2_U4377 , P2_R1095_U105 , P2_U3880 );
nand NAND2_4930 ( P2_U4378 , P2_R1143_U12 , P2_U3877 );
nand NAND2_4931 ( P2_U4379 , P2_R1161_U12 , P2_U3887 );
nand NAND2_4932 ( P2_U4380 , P2_R1131_U105 , P2_U3883 );
nand NAND2_4933 ( P2_U4381 , P2_R1200_U105 , P2_U3017 );
not NOT1_4934 ( P2_U4382 , P2_U3331 );
nand NAND2_4935 ( P2_U4383 , P2_R1179_U105 , P2_U3026 );
nand NAND2_4936 ( P2_U4384 , P2_U3025 , P2_U3081 );
nand NAND2_4937 ( P2_U4385 , P2_U3440 , P2_U4060 );
nand NAND2_4938 ( P2_U4386 , P2_U3650 , P2_U4382 );
nand NAND2_4939 ( P2_U4387 , P2_REG0_REG_19_ , P2_U3022 );
nand NAND2_4940 ( P2_U4388 , P2_REG1_REG_19_ , P2_U3021 );
nand NAND2_4941 ( P2_U4389 , P2_REG2_REG_19_ , P2_U3020 );
nand NAND2_4942 ( P2_U4390 , P2_SUB_605_U15 , P2_U3019 );
not NOT1_4943 ( P2_U4391 , P2_U3080 );
nand NAND2_4944 ( P2_U4392 , P2_U3033 , P2_U3068 );
nand NAND2_4945 ( P2_U4393 , P2_R1110_U109 , P2_U3879 );
nand NAND2_4946 ( P2_U4394 , P2_R1077_U109 , P2_U3881 );
nand NAND2_4947 ( P2_U4395 , P2_R1095_U104 , P2_U3880 );
nand NAND2_4948 ( P2_U4396 , P2_R1143_U109 , P2_U3877 );
nand NAND2_4949 ( P2_U4397 , P2_R1161_U109 , P2_U3887 );
nand NAND2_4950 ( P2_U4398 , P2_R1131_U104 , P2_U3883 );
nand NAND2_4951 ( P2_U4399 , P2_R1200_U104 , P2_U3017 );
not NOT1_4952 ( P2_U4400 , P2_U3332 );
nand NAND2_4953 ( P2_U4401 , P2_R1179_U104 , P2_U3026 );
nand NAND2_4954 ( P2_U4402 , P2_U3025 , P2_U3080 );
nand NAND2_4955 ( P2_U4403 , P2_U3443 , P2_U4060 );
nand NAND2_4956 ( P2_U4404 , P2_U3654 , P2_U4400 );
nand NAND2_4957 ( P2_U4405 , P2_REG2_REG_20_ , P2_U3020 );
nand NAND2_4958 ( P2_U4406 , P2_REG1_REG_20_ , P2_U3021 );
nand NAND2_4959 ( P2_U4407 , P2_REG0_REG_20_ , P2_U3022 );
nand NAND2_4960 ( P2_U4408 , P2_SUB_605_U20 , P2_U3019 );
not NOT1_4961 ( P2_U4409 , P2_U3075 );
nand NAND2_4962 ( P2_U4410 , P2_U3033 , P2_U3081 );
nand NAND2_4963 ( P2_U4411 , P2_R1110_U108 , P2_U3879 );
nand NAND2_4964 ( P2_U4412 , P2_R1077_U108 , P2_U3881 );
nand NAND2_4965 ( P2_U4413 , P2_R1095_U103 , P2_U3880 );
nand NAND2_4966 ( P2_U4414 , P2_R1143_U108 , P2_U3877 );
nand NAND2_4967 ( P2_U4415 , P2_R1161_U108 , P2_U3887 );
nand NAND2_4968 ( P2_U4416 , P2_R1131_U103 , P2_U3883 );
nand NAND2_4969 ( P2_U4417 , P2_R1200_U103 , P2_U3017 );
not NOT1_4970 ( P2_U4418 , P2_U3333 );
nand NAND2_4971 ( P2_U4419 , P2_R1179_U103 , P2_U3026 );
nand NAND2_4972 ( P2_U4420 , P2_U3025 , P2_U3075 );
nand NAND2_4973 ( P2_U4421 , P2_U3445 , P2_U4060 );
nand NAND2_4974 ( P2_U4422 , P2_U3658 , P2_U4418 );
nand NAND2_4975 ( P2_U4423 , P2_REG2_REG_21_ , P2_U3020 );
nand NAND2_4976 ( P2_U4424 , P2_REG1_REG_21_ , P2_U3021 );
nand NAND2_4977 ( P2_U4425 , P2_REG0_REG_21_ , P2_U3022 );
nand NAND2_4978 ( P2_U4426 , P2_SUB_605_U28 , P2_U3019 );
not NOT1_4979 ( P2_U4427 , P2_U3074 );
nand NAND2_4980 ( P2_U4428 , P2_U3033 , P2_U3080 );
nand NAND2_4981 ( P2_U4429 , P2_R1110_U13 , P2_U3879 );
nand NAND2_4982 ( P2_U4430 , P2_R1077_U13 , P2_U3881 );
nand NAND2_4983 ( P2_U4431 , P2_R1095_U101 , P2_U3880 );
nand NAND2_4984 ( P2_U4432 , P2_R1143_U13 , P2_U3877 );
nand NAND2_4985 ( P2_U4433 , P2_R1161_U13 , P2_U3887 );
nand NAND2_4986 ( P2_U4434 , P2_R1131_U101 , P2_U3883 );
nand NAND2_4987 ( P2_U4435 , P2_R1200_U101 , P2_U3017 );
not NOT1_4988 ( P2_U4436 , P2_U3335 );
nand NAND2_4989 ( P2_U4437 , P2_R1179_U101 , P2_U3026 );
nand NAND2_4990 ( P2_U4438 , P2_U3025 , P2_U3074 );
nand NAND2_4991 ( P2_U4439 , P2_U3903 , P2_U4060 );
nand NAND2_4992 ( P2_U4440 , P2_U3662 , P2_U4436 );
nand NAND2_4993 ( P2_U4441 , P2_REG2_REG_22_ , P2_U3020 );
nand NAND2_4994 ( P2_U4442 , P2_REG1_REG_22_ , P2_U3021 );
nand NAND2_4995 ( P2_U4443 , P2_REG0_REG_22_ , P2_U3022 );
nand NAND2_4996 ( P2_U4444 , P2_SUB_605_U17 , P2_U3019 );
not NOT1_4997 ( P2_U4445 , P2_U3060 );
nand NAND2_4998 ( P2_U4446 , P2_U3033 , P2_U3075 );
nand NAND2_4999 ( P2_U4447 , P2_R1110_U14 , P2_U3879 );
nand NAND2_5000 ( P2_U4448 , P2_R1077_U14 , P2_U3881 );
nand NAND2_5001 ( P2_U4449 , P2_R1095_U115 , P2_U3880 );
nand NAND2_5002 ( P2_U4450 , P2_R1143_U14 , P2_U3877 );
nand NAND2_5003 ( P2_U4451 , P2_R1161_U14 , P2_U3887 );
nand NAND2_5004 ( P2_U4452 , P2_R1131_U115 , P2_U3883 );
nand NAND2_5005 ( P2_U4453 , P2_R1200_U115 , P2_U3017 );
not NOT1_5006 ( P2_U4454 , P2_U3337 );
nand NAND2_5007 ( P2_U4455 , P2_R1179_U115 , P2_U3026 );
nand NAND2_5008 ( P2_U4456 , P2_U3025 , P2_U3060 );
nand NAND2_5009 ( P2_U4457 , P2_U3902 , P2_U4060 );
nand NAND2_5010 ( P2_U4458 , P2_U3665 , P2_U4454 );
nand NAND2_5011 ( P2_U4459 , P2_REG2_REG_23_ , P2_U3020 );
nand NAND2_5012 ( P2_U4460 , P2_REG1_REG_23_ , P2_U3021 );
nand NAND2_5013 ( P2_U4461 , P2_REG0_REG_23_ , P2_U3022 );
nand NAND2_5014 ( P2_U4462 , P2_SUB_605_U6 , P2_U3019 );
not NOT1_5015 ( P2_U4463 , P2_U3065 );
nand NAND2_5016 ( P2_U4464 , P2_U3033 , P2_U3074 );
nand NAND2_5017 ( P2_U4465 , P2_R1110_U107 , P2_U3879 );
nand NAND2_5018 ( P2_U4466 , P2_R1077_U107 , P2_U3881 );
nand NAND2_5019 ( P2_U4467 , P2_R1095_U114 , P2_U3880 );
nand NAND2_5020 ( P2_U4468 , P2_R1143_U107 , P2_U3877 );
nand NAND2_5021 ( P2_U4469 , P2_R1161_U107 , P2_U3887 );
nand NAND2_5022 ( P2_U4470 , P2_R1131_U114 , P2_U3883 );
nand NAND2_5023 ( P2_U4471 , P2_R1200_U114 , P2_U3017 );
not NOT1_5024 ( P2_U4472 , P2_U3339 );
nand NAND2_5025 ( P2_U4473 , P2_R1179_U114 , P2_U3026 );
nand NAND2_5026 ( P2_U4474 , P2_U3025 , P2_U3065 );
nand NAND2_5027 ( P2_U4475 , P2_U3901 , P2_U4060 );
nand NAND2_5028 ( P2_U4476 , P2_U3668 , P2_U4472 );
nand NAND2_5029 ( P2_U4477 , P2_REG2_REG_24_ , P2_U3020 );
nand NAND2_5030 ( P2_U4478 , P2_REG1_REG_24_ , P2_U3021 );
nand NAND2_5031 ( P2_U4479 , P2_REG0_REG_24_ , P2_U3022 );
nand NAND2_5032 ( P2_U4480 , P2_SUB_605_U10 , P2_U3019 );
not NOT1_5033 ( P2_U4481 , P2_U3064 );
nand NAND2_5034 ( P2_U4482 , P2_U3033 , P2_U3060 );
nand NAND2_5035 ( P2_U4483 , P2_R1110_U106 , P2_U3879 );
nand NAND2_5036 ( P2_U4484 , P2_R1077_U106 , P2_U3881 );
nand NAND2_5037 ( P2_U4485 , P2_R1095_U19 , P2_U3880 );
nand NAND2_5038 ( P2_U4486 , P2_R1143_U106 , P2_U3877 );
nand NAND2_5039 ( P2_U4487 , P2_R1161_U106 , P2_U3887 );
nand NAND2_5040 ( P2_U4488 , P2_R1131_U19 , P2_U3883 );
nand NAND2_5041 ( P2_U4489 , P2_R1200_U19 , P2_U3017 );
not NOT1_5042 ( P2_U4490 , P2_U3341 );
nand NAND2_5043 ( P2_U4491 , P2_R1179_U19 , P2_U3026 );
nand NAND2_5044 ( P2_U4492 , P2_U3025 , P2_U3064 );
nand NAND2_5045 ( P2_U4493 , P2_U3900 , P2_U4060 );
nand NAND2_5046 ( P2_U4494 , P2_U3671 , P2_U4490 );
nand NAND2_5047 ( P2_U4495 , P2_REG2_REG_25_ , P2_U3020 );
nand NAND2_5048 ( P2_U4496 , P2_REG1_REG_25_ , P2_U3021 );
nand NAND2_5049 ( P2_U4497 , P2_REG0_REG_25_ , P2_U3022 );
nand NAND2_5050 ( P2_U4498 , P2_SUB_605_U16 , P2_U3019 );
not NOT1_5051 ( P2_U4499 , P2_U3057 );
nand NAND2_5052 ( P2_U4500 , P2_U3033 , P2_U3065 );
nand NAND2_5053 ( P2_U4501 , P2_R1110_U105 , P2_U3879 );
nand NAND2_5054 ( P2_U4502 , P2_R1077_U105 , P2_U3881 );
nand NAND2_5055 ( P2_U4503 , P2_R1095_U100 , P2_U3880 );
nand NAND2_5056 ( P2_U4504 , P2_R1143_U105 , P2_U3877 );
nand NAND2_5057 ( P2_U4505 , P2_R1161_U105 , P2_U3887 );
nand NAND2_5058 ( P2_U4506 , P2_R1131_U100 , P2_U3883 );
nand NAND2_5059 ( P2_U4507 , P2_R1200_U100 , P2_U3017 );
not NOT1_5060 ( P2_U4508 , P2_U3343 );
nand NAND2_5061 ( P2_U4509 , P2_R1179_U100 , P2_U3026 );
nand NAND2_5062 ( P2_U4510 , P2_U3025 , P2_U3057 );
nand NAND2_5063 ( P2_U4511 , P2_U3899 , P2_U4060 );
nand NAND2_5064 ( P2_U4512 , P2_U3675 , P2_U4508 );
nand NAND2_5065 ( P2_U4513 , P2_REG2_REG_26_ , P2_U3020 );
nand NAND2_5066 ( P2_U4514 , P2_REG1_REG_26_ , P2_U3021 );
nand NAND2_5067 ( P2_U4515 , P2_REG0_REG_26_ , P2_U3022 );
nand NAND2_5068 ( P2_U4516 , P2_SUB_605_U27 , P2_U3019 );
not NOT1_5069 ( P2_U4517 , P2_U3056 );
nand NAND2_5070 ( P2_U4518 , P2_U3033 , P2_U3064 );
nand NAND2_5071 ( P2_U4519 , P2_R1110_U104 , P2_U3879 );
nand NAND2_5072 ( P2_U4520 , P2_R1077_U104 , P2_U3881 );
nand NAND2_5073 ( P2_U4521 , P2_R1095_U99 , P2_U3880 );
nand NAND2_5074 ( P2_U4522 , P2_R1143_U104 , P2_U3877 );
nand NAND2_5075 ( P2_U4523 , P2_R1161_U104 , P2_U3887 );
nand NAND2_5076 ( P2_U4524 , P2_R1131_U99 , P2_U3883 );
nand NAND2_5077 ( P2_U4525 , P2_R1200_U99 , P2_U3017 );
not NOT1_5078 ( P2_U4526 , P2_U3345 );
nand NAND2_5079 ( P2_U4527 , P2_R1179_U99 , P2_U3026 );
nand NAND2_5080 ( P2_U4528 , P2_U3025 , P2_U3056 );
nand NAND2_5081 ( P2_U4529 , P2_U3898 , P2_U4060 );
nand NAND2_5082 ( P2_U4530 , P2_U3679 , P2_U4526 );
nand NAND2_5083 ( P2_U4531 , P2_REG2_REG_27_ , P2_U3020 );
nand NAND2_5084 ( P2_U4532 , P2_REG1_REG_27_ , P2_U3021 );
nand NAND2_5085 ( P2_U4533 , P2_REG0_REG_27_ , P2_U3022 );
nand NAND2_5086 ( P2_U4534 , P2_SUB_605_U23 , P2_U3019 );
not NOT1_5087 ( P2_U4535 , P2_U3052 );
nand NAND2_5088 ( P2_U4536 , P2_U3033 , P2_U3057 );
nand NAND2_5089 ( P2_U4537 , P2_R1110_U15 , P2_U3879 );
nand NAND2_5090 ( P2_U4538 , P2_R1077_U15 , P2_U3881 );
nand NAND2_5091 ( P2_U4539 , P2_R1095_U113 , P2_U3880 );
nand NAND2_5092 ( P2_U4540 , P2_R1143_U15 , P2_U3877 );
nand NAND2_5093 ( P2_U4541 , P2_R1161_U15 , P2_U3887 );
nand NAND2_5094 ( P2_U4542 , P2_R1131_U113 , P2_U3883 );
nand NAND2_5095 ( P2_U4543 , P2_R1200_U113 , P2_U3017 );
not NOT1_5096 ( P2_U4544 , P2_U3347 );
nand NAND2_5097 ( P2_U4545 , P2_R1179_U113 , P2_U3026 );
nand NAND2_5098 ( P2_U4546 , P2_U3025 , P2_U3052 );
nand NAND2_5099 ( P2_U4547 , P2_U3897 , P2_U4060 );
nand NAND2_5100 ( P2_U4548 , P2_U3683 , P2_U4544 );
nand NAND2_5101 ( P2_U4549 , P2_REG2_REG_28_ , P2_U3020 );
nand NAND2_5102 ( P2_U4550 , P2_REG1_REG_28_ , P2_U3021 );
nand NAND2_5103 ( P2_U4551 , P2_REG0_REG_28_ , P2_U3022 );
nand NAND2_5104 ( P2_U4552 , P2_SUB_605_U29 , P2_U3019 );
not NOT1_5105 ( P2_U4553 , P2_U3053 );
nand NAND2_5106 ( P2_U4554 , P2_U3033 , P2_U3056 );
nand NAND2_5107 ( P2_U4555 , P2_R1110_U103 , P2_U3879 );
nand NAND2_5108 ( P2_U4556 , P2_R1077_U103 , P2_U3881 );
nand NAND2_5109 ( P2_U4557 , P2_R1095_U20 , P2_U3880 );
nand NAND2_5110 ( P2_U4558 , P2_R1143_U103 , P2_U3877 );
nand NAND2_5111 ( P2_U4559 , P2_R1161_U103 , P2_U3887 );
nand NAND2_5112 ( P2_U4560 , P2_R1131_U20 , P2_U3883 );
nand NAND2_5113 ( P2_U4561 , P2_R1200_U20 , P2_U3017 );
not NOT1_5114 ( P2_U4562 , P2_U3349 );
nand NAND2_5115 ( P2_U4563 , P2_R1179_U20 , P2_U3026 );
nand NAND2_5116 ( P2_U4564 , P2_U3025 , P2_U3053 );
nand NAND2_5117 ( P2_U4565 , P2_U3896 , P2_U4060 );
nand NAND2_5118 ( P2_U4566 , P2_U3687 , P2_U4562 );
nand NAND2_5119 ( P2_U4567 , P2_SUB_605_U94 , P2_U3019 );
nand NAND2_5120 ( P2_U4568 , P2_REG2_REG_29_ , P2_U3020 );
nand NAND2_5121 ( P2_U4569 , P2_REG1_REG_29_ , P2_U3021 );
nand NAND2_5122 ( P2_U4570 , P2_REG0_REG_29_ , P2_U3022 );
not NOT1_5123 ( P2_U4571 , P2_U3054 );
nand NAND2_5124 ( P2_U4572 , P2_U3033 , P2_U3052 );
nand NAND2_5125 ( P2_U4573 , P2_R1110_U102 , P2_U3879 );
nand NAND2_5126 ( P2_U4574 , P2_R1077_U102 , P2_U3881 );
nand NAND2_5127 ( P2_U4575 , P2_R1095_U98 , P2_U3880 );
nand NAND2_5128 ( P2_U4576 , P2_R1143_U102 , P2_U3877 );
nand NAND2_5129 ( P2_U4577 , P2_R1161_U102 , P2_U3887 );
nand NAND2_5130 ( P2_U4578 , P2_R1131_U98 , P2_U3883 );
nand NAND2_5131 ( P2_U4579 , P2_R1200_U98 , P2_U3017 );
not NOT1_5132 ( P2_U4580 , P2_U3351 );
nand NAND2_5133 ( P2_U4581 , P2_R1179_U98 , P2_U3026 );
nand NAND2_5134 ( P2_U4582 , P2_U3025 , P2_U3054 );
nand NAND2_5135 ( P2_U4583 , P2_U3895 , P2_U4060 );
nand NAND2_5136 ( P2_U4584 , P2_U3691 , P2_U4580 );
nand NAND2_5137 ( P2_U4585 , P2_REG2_REG_30_ , P2_U3020 );
nand NAND2_5138 ( P2_U4586 , P2_REG1_REG_30_ , P2_U3021 );
nand NAND2_5139 ( P2_U4587 , P2_REG0_REG_30_ , P2_U3022 );
nand NAND2_5140 ( P2_U4588 , P2_SUB_605_U94 , P2_U3019 );
not NOT1_5141 ( P2_U4589 , P2_U3058 );
nand NAND2_5142 ( P2_U4590 , P2_U3888 , P2_U3298 );
nand NAND2_5143 ( P2_U4591 , P2_U3829 , P2_U4590 );
nand NAND3_5144 ( P2_U4592 , P2_U4591 , P2_U3907 , P2_U3058 );
nand NAND2_5145 ( P2_U4593 , P2_U3033 , P2_U3053 );
nand NAND2_5146 ( P2_U4594 , P2_R1110_U101 , P2_U3879 );
nand NAND2_5147 ( P2_U4595 , P2_R1077_U101 , P2_U3881 );
nand NAND2_5148 ( P2_U4596 , P2_R1095_U21 , P2_U3880 );
nand NAND2_5149 ( P2_U4597 , P2_R1143_U101 , P2_U3877 );
nand NAND2_5150 ( P2_U4598 , P2_R1161_U101 , P2_U3887 );
nand NAND2_5151 ( P2_U4599 , P2_R1131_U21 , P2_U3883 );
nand NAND2_5152 ( P2_U4600 , P2_R1200_U21 , P2_U3017 );
not NOT1_5153 ( P2_U4601 , P2_U3354 );
nand NAND2_5154 ( P2_U4602 , P2_R1179_U21 , P2_U3026 );
nand NAND2_5155 ( P2_U4603 , P2_U3904 , P2_U4060 );
nand NAND2_5156 ( P2_U4604 , P2_U3695 , P2_U4601 );
nand NAND2_5157 ( P2_U4605 , P2_SUB_605_U94 , P2_U3019 );
nand NAND2_5158 ( P2_U4606 , P2_REG2_REG_31_ , P2_U3020 );
nand NAND2_5159 ( P2_U4607 , P2_REG1_REG_31_ , P2_U3021 );
nand NAND2_5160 ( P2_U4608 , P2_REG0_REG_31_ , P2_U3022 );
not NOT1_5161 ( P2_U4609 , P2_U3055 );
nand NAND2_5162 ( P2_U4610 , P2_U3869 , P2_U4060 );
nand NAND2_5163 ( P2_U4611 , P2_U3361 , P2_U4610 );
nand NAND2_5164 ( P2_U4612 , P2_U3868 , P2_U4060 );
nand NAND2_5165 ( P2_U4613 , P2_U3361 , P2_U4612 );
nand NAND3_5166 ( P2_U4614 , P2_U5637 , P2_U5636 , P2_U3302 );
nand NAND2_5167 ( P2_U4615 , P2_U3884 , P2_U3367 );
nand NAND2_5168 ( P2_U4616 , P2_U3048 , P2_U4615 );
nand NAND2_5169 ( P2_U4617 , P2_U3047 , P2_U4614 );
nand NAND2_5170 ( P2_U4618 , P2_U4617 , P2_U4616 );
nand NAND2_5171 ( P2_U4619 , P2_U5452 , P2_U3379 );
nand NAND3_5172 ( P2_U4620 , P2_U4619 , P2_U3380 , P2_U3830 );
nand NAND2_5173 ( P2_U4621 , P2_U3048 , P2_U4620 );
nand NAND2_5174 ( P2_U4622 , P2_U3047 , P2_U4615 );
nand NAND3_5175 ( P2_U4623 , P2_U4621 , P2_U3360 , P2_U4622 );
not NOT1_5176 ( P2_U4624 , P2_U3365 );
nand NAND2_5177 ( P2_U4625 , P2_U3034 , P2_U3077 );
nand NAND2_5178 ( P2_U4626 , P2_U3030 , P2_R1179_U25 );
nand NAND2_5179 ( P2_U4627 , P2_U3029 , P2_U3387 );
nand NAND2_5180 ( P2_U4628 , P2_U3028 , P2_REG3_REG_0_ );
nand NAND2_5181 ( P2_U4629 , P2_U3034 , P2_U3067 );
nand NAND2_5182 ( P2_U4630 , P2_U3030 , P2_R1179_U102 );
nand NAND2_5183 ( P2_U4631 , P2_U3029 , P2_U3392 );
nand NAND2_5184 ( P2_U4632 , P2_U3028 , P2_REG3_REG_1_ );
nand NAND2_5185 ( P2_U4633 , P2_U3034 , P2_U3063 );
nand NAND2_5186 ( P2_U4634 , P2_U3030 , P2_R1179_U112 );
nand NAND2_5187 ( P2_U4635 , P2_U3029 , P2_U3395 );
nand NAND2_5188 ( P2_U4636 , P2_U3028 , P2_REG3_REG_2_ );
nand NAND2_5189 ( P2_U4637 , P2_U3034 , P2_U3059 );
nand NAND2_5190 ( P2_U4638 , P2_U3030 , P2_R1179_U22 );
nand NAND2_5191 ( P2_U4639 , P2_U3029 , P2_U3398 );
nand NAND2_5192 ( P2_U4640 , P2_U3028 , P2_SUB_605_U26 );
nand NAND2_5193 ( P2_U4641 , P2_U3034 , P2_U3066 );
nand NAND2_5194 ( P2_U4642 , P2_U3030 , P2_R1179_U111 );
nand NAND2_5195 ( P2_U4643 , P2_U3029 , P2_U3401 );
nand NAND2_5196 ( P2_U4644 , P2_U3028 , P2_SUB_605_U30 );
nand NAND2_5197 ( P2_U4645 , P2_U3034 , P2_U3070 );
nand NAND2_5198 ( P2_U4646 , P2_U3030 , P2_R1179_U110 );
nand NAND2_5199 ( P2_U4647 , P2_U3029 , P2_U3404 );
nand NAND2_5200 ( P2_U4648 , P2_U3028 , P2_SUB_605_U22 );
nand NAND2_5201 ( P2_U4649 , P2_U3034 , P2_U3069 );
nand NAND2_5202 ( P2_U4650 , P2_U3030 , P2_R1179_U23 );
nand NAND2_5203 ( P2_U4651 , P2_U3029 , P2_U3407 );
nand NAND2_5204 ( P2_U4652 , P2_U3028 , P2_SUB_605_U8 );
nand NAND2_5205 ( P2_U4653 , P2_U3034 , P2_U3083 );
nand NAND2_5206 ( P2_U4654 , P2_U3030 , P2_R1179_U109 );
nand NAND2_5207 ( P2_U4655 , P2_U3029 , P2_U3410 );
nand NAND2_5208 ( P2_U4656 , P2_U3028 , P2_SUB_605_U18 );
nand NAND2_5209 ( P2_U4657 , P2_U3034 , P2_U3082 );
nand NAND2_5210 ( P2_U4658 , P2_U3030 , P2_R1179_U24 );
nand NAND2_5211 ( P2_U4659 , P2_U3029 , P2_U3413 );
nand NAND2_5212 ( P2_U4660 , P2_U3028 , P2_SUB_605_U12 );
nand NAND2_5213 ( P2_U4661 , P2_U3034 , P2_U3061 );
nand NAND2_5214 ( P2_U4662 , P2_U3030 , P2_R1179_U108 );
nand NAND2_5215 ( P2_U4663 , P2_U3029 , P2_U3416 );
nand NAND2_5216 ( P2_U4664 , P2_U3028 , P2_SUB_605_U14 );
nand NAND2_5217 ( P2_U4665 , P2_U3034 , P2_U3062 );
nand NAND2_5218 ( P2_U4666 , P2_U3030 , P2_R1179_U118 );
nand NAND2_5219 ( P2_U4667 , P2_U3029 , P2_U3419 );
nand NAND2_5220 ( P2_U4668 , P2_U3028 , P2_SUB_605_U13 );
nand NAND2_5221 ( P2_U4669 , P2_U3034 , P2_U3071 );
nand NAND2_5222 ( P2_U4670 , P2_U3030 , P2_R1179_U17 );
nand NAND2_5223 ( P2_U4671 , P2_U3029 , P2_U3422 );
nand NAND2_5224 ( P2_U4672 , P2_U3028 , P2_SUB_605_U9 );
nand NAND2_5225 ( P2_U4673 , P2_U3034 , P2_U3079 );
nand NAND2_5226 ( P2_U4674 , P2_U3030 , P2_R1179_U107 );
nand NAND2_5227 ( P2_U4675 , P2_U3029 , P2_U3425 );
nand NAND2_5228 ( P2_U4676 , P2_U3028 , P2_SUB_605_U24 );
nand NAND2_5229 ( P2_U4677 , P2_U3034 , P2_U3078 );
nand NAND2_5230 ( P2_U4678 , P2_U3030 , P2_R1179_U106 );
nand NAND2_5231 ( P2_U4679 , P2_U3029 , P2_U3428 );
nand NAND2_5232 ( P2_U4680 , P2_U3028 , P2_SUB_605_U25 );
nand NAND2_5233 ( P2_U4681 , P2_U3034 , P2_U3073 );
nand NAND2_5234 ( P2_U4682 , P2_U3030 , P2_R1179_U117 );
nand NAND2_5235 ( P2_U4683 , P2_U3029 , P2_U3431 );
nand NAND2_5236 ( P2_U4684 , P2_U3028 , P2_SUB_605_U31 );
nand NAND2_5237 ( P2_U4685 , P2_U3034 , P2_U3072 );
nand NAND2_5238 ( P2_U4686 , P2_U3030 , P2_R1179_U116 );
nand NAND2_5239 ( P2_U4687 , P2_U3029 , P2_U3434 );
nand NAND2_5240 ( P2_U4688 , P2_U3028 , P2_SUB_605_U21 );
nand NAND2_5241 ( P2_U4689 , P2_U3034 , P2_U3068 );
nand NAND2_5242 ( P2_U4690 , P2_U3030 , P2_R1179_U18 );
nand NAND2_5243 ( P2_U4691 , P2_U3029 , P2_U3437 );
nand NAND2_5244 ( P2_U4692 , P2_U3028 , P2_SUB_605_U7 );
nand NAND2_5245 ( P2_U4693 , P2_U3034 , P2_U3081 );
nand NAND2_5246 ( P2_U4694 , P2_U3030 , P2_R1179_U105 );
nand NAND2_5247 ( P2_U4695 , P2_U3029 , P2_U3440 );
nand NAND2_5248 ( P2_U4696 , P2_U3028 , P2_SUB_605_U19 );
nand NAND2_5249 ( P2_U4697 , P2_U3034 , P2_U3080 );
nand NAND2_5250 ( P2_U4698 , P2_U3030 , P2_R1179_U104 );
nand NAND2_5251 ( P2_U4699 , P2_U3029 , P2_U3443 );
nand NAND2_5252 ( P2_U4700 , P2_U3028 , P2_SUB_605_U11 );
nand NAND2_5253 ( P2_U4701 , P2_U3034 , P2_U3075 );
nand NAND2_5254 ( P2_U4702 , P2_U3030 , P2_R1179_U103 );
nand NAND2_5255 ( P2_U4703 , P2_U3029 , P2_U3445 );
nand NAND2_5256 ( P2_U4704 , P2_U3028 , P2_SUB_605_U15 );
nand NAND2_5257 ( P2_U4705 , P2_U3034 , P2_U3074 );
nand NAND2_5258 ( P2_U4706 , P2_U3030 , P2_R1179_U101 );
nand NAND2_5259 ( P2_U4707 , P2_U3029 , P2_U3903 );
nand NAND2_5260 ( P2_U4708 , P2_U3028 , P2_SUB_605_U20 );
nand NAND2_5261 ( P2_U4709 , P2_U3034 , P2_U3060 );
nand NAND2_5262 ( P2_U4710 , P2_U3030 , P2_R1179_U115 );
nand NAND2_5263 ( P2_U4711 , P2_U3029 , P2_U3902 );
nand NAND2_5264 ( P2_U4712 , P2_U3028 , P2_SUB_605_U28 );
nand NAND2_5265 ( P2_U4713 , P2_U3034 , P2_U3065 );
nand NAND2_5266 ( P2_U4714 , P2_U3030 , P2_R1179_U114 );
nand NAND2_5267 ( P2_U4715 , P2_U3029 , P2_U3901 );
nand NAND2_5268 ( P2_U4716 , P2_U3028 , P2_SUB_605_U17 );
nand NAND2_5269 ( P2_U4717 , P2_U3034 , P2_U3064 );
nand NAND2_5270 ( P2_U4718 , P2_U3030 , P2_R1179_U19 );
nand NAND2_5271 ( P2_U4719 , P2_U3029 , P2_U3900 );
nand NAND2_5272 ( P2_U4720 , P2_U3028 , P2_SUB_605_U6 );
nand NAND2_5273 ( P2_U4721 , P2_U3034 , P2_U3057 );
nand NAND2_5274 ( P2_U4722 , P2_U3030 , P2_R1179_U100 );
nand NAND2_5275 ( P2_U4723 , P2_U3029 , P2_U3899 );
nand NAND2_5276 ( P2_U4724 , P2_U3028 , P2_SUB_605_U10 );
nand NAND2_5277 ( P2_U4725 , P2_U3034 , P2_U3056 );
nand NAND2_5278 ( P2_U4726 , P2_U3030 , P2_R1179_U99 );
nand NAND2_5279 ( P2_U4727 , P2_U3029 , P2_U3898 );
nand NAND2_5280 ( P2_U4728 , P2_U3028 , P2_SUB_605_U16 );
nand NAND2_5281 ( P2_U4729 , P2_U3034 , P2_U3052 );
nand NAND2_5282 ( P2_U4730 , P2_U3030 , P2_R1179_U113 );
nand NAND2_5283 ( P2_U4731 , P2_U3029 , P2_U3897 );
nand NAND2_5284 ( P2_U4732 , P2_U3028 , P2_SUB_605_U27 );
nand NAND2_5285 ( P2_U4733 , P2_U3034 , P2_U3053 );
nand NAND2_5286 ( P2_U4734 , P2_U3030 , P2_R1179_U20 );
nand NAND2_5287 ( P2_U4735 , P2_U3029 , P2_U3896 );
nand NAND2_5288 ( P2_U4736 , P2_U3028 , P2_SUB_605_U23 );
nand NAND2_5289 ( P2_U4737 , P2_U3034 , P2_U3054 );
nand NAND2_5290 ( P2_U4738 , P2_U3030 , P2_R1179_U98 );
nand NAND2_5291 ( P2_U4739 , P2_U3029 , P2_U3895 );
nand NAND2_5292 ( P2_U4740 , P2_U3028 , P2_SUB_605_U29 );
nand NAND2_5293 ( P2_U4741 , P2_U3030 , P2_R1179_U21 );
nand NAND2_5294 ( P2_U4742 , P2_U3029 , P2_U3904 );
nand NAND2_5295 ( P2_U4743 , P2_U3028 , P2_SUB_605_U94 );
nand NAND2_5296 ( P2_U4744 , P2_U3028 , P2_SUB_605_U94 );
nand NAND2_5297 ( P2_U4745 , P2_U3912 , P2_U3908 );
nand NAND2_5298 ( P2_U4746 , P2_U3029 , P2_U3869 );
nand NAND2_5299 ( P2_U4747 , P2_REG2_REG_30_ , P2_U3358 );
nand NAND2_5300 ( P2_U4748 , P2_U3029 , P2_U3868 );
nand NAND2_5301 ( P2_U4749 , P2_REG2_REG_31_ , P2_U3358 );
nand NAND4_5302 ( P2_U4750 , P2_U4624 , P2_U3359 , P2_U3703 , P2_U3702 );
nand NAND2_5303 ( P2_U4751 , P2_R1212_U6 , P2_U3040 );
nand NAND2_5304 ( P2_U4752 , P2_U3039 , P2_U3379 );
nand NAND2_5305 ( P2_U4753 , P2_R1209_U6 , P2_U3037 );
nand NAND3_5306 ( P2_U4754 , P2_U4752 , P2_U4751 , P2_U4753 );
nand NAND2_5307 ( P2_U4755 , P2_U3906 , P2_U5436 );
not NOT1_5308 ( P2_U4756 , P2_U3366 );
nand NAND2_5309 ( P2_U4757 , P2_U3829 , P2_U3892 );
nand NAND2_5310 ( P2_U4758 , P2_R1054_U67 , P2_U3051 );
nand NAND2_5311 ( P2_U4759 , P2_U5764 , P2_U3379 );
nand NAND2_5312 ( P2_U4760 , P2_U3042 , P2_U4754 );
nand NAND2_5313 ( P2_U4761 , P2_U3041 , P2_R1212_U6 );
nand NAND2_5314 ( P2_U4762 , P2_REG3_REG_19_ , P2_U3151 );
nand NAND2_5315 ( P2_U4763 , P2_U3038 , P2_R1209_U6 );
nand NAND2_5316 ( P2_U4764 , P2_ADDR_REG_19_ , P2_U4756 );
nand NAND2_5317 ( P2_U4765 , P2_R1212_U58 , P2_U3040 );
nand NAND2_5318 ( P2_U4766 , P2_U3039 , P2_U3442 );
nand NAND2_5319 ( P2_U4767 , P2_R1209_U58 , P2_U3037 );
nand NAND3_5320 ( P2_U4768 , P2_U4766 , P2_U4765 , P2_U4767 );
nand NAND2_5321 ( P2_U4769 , P2_R1054_U68 , P2_U3051 );
nand NAND2_5322 ( P2_U4770 , P2_U5764 , P2_U3442 );
nand NAND2_5323 ( P2_U4771 , P2_U3042 , P2_U4768 );
nand NAND2_5324 ( P2_U4772 , P2_R1212_U58 , P2_U3041 );
nand NAND2_5325 ( P2_U4773 , P2_REG3_REG_18_ , P2_U3151 );
nand NAND2_5326 ( P2_U4774 , P2_R1209_U58 , P2_U3038 );
nand NAND2_5327 ( P2_U4775 , P2_ADDR_REG_18_ , P2_U4756 );
nand NAND2_5328 ( P2_U4776 , P2_R1212_U59 , P2_U3040 );
nand NAND2_5329 ( P2_U4777 , P2_U3039 , P2_U3439 );
nand NAND2_5330 ( P2_U4778 , P2_R1209_U59 , P2_U3037 );
nand NAND3_5331 ( P2_U4779 , P2_U4777 , P2_U4776 , P2_U4778 );
nand NAND2_5332 ( P2_U4780 , P2_R1054_U69 , P2_U3051 );
nand NAND2_5333 ( P2_U4781 , P2_U5764 , P2_U3439 );
nand NAND2_5334 ( P2_U4782 , P2_U3042 , P2_U4779 );
nand NAND2_5335 ( P2_U4783 , P2_R1212_U59 , P2_U3041 );
nand NAND2_5336 ( P2_U4784 , P2_REG3_REG_17_ , P2_U3151 );
nand NAND2_5337 ( P2_U4785 , P2_R1209_U59 , P2_U3038 );
nand NAND2_5338 ( P2_U4786 , P2_ADDR_REG_17_ , P2_U4756 );
nand NAND2_5339 ( P2_U4787 , P2_R1212_U60 , P2_U3040 );
nand NAND2_5340 ( P2_U4788 , P2_U3039 , P2_U3436 );
nand NAND2_5341 ( P2_U4789 , P2_R1209_U60 , P2_U3037 );
nand NAND3_5342 ( P2_U4790 , P2_U4788 , P2_U4787 , P2_U4789 );
nand NAND2_5343 ( P2_U4791 , P2_R1054_U13 , P2_U3051 );
nand NAND2_5344 ( P2_U4792 , P2_U5764 , P2_U3436 );
nand NAND2_5345 ( P2_U4793 , P2_U3042 , P2_U4790 );
nand NAND2_5346 ( P2_U4794 , P2_R1212_U60 , P2_U3041 );
nand NAND2_5347 ( P2_U4795 , P2_REG3_REG_16_ , P2_U3151 );
nand NAND2_5348 ( P2_U4796 , P2_R1209_U60 , P2_U3038 );
nand NAND2_5349 ( P2_U4797 , P2_ADDR_REG_16_ , P2_U4756 );
nand NAND2_5350 ( P2_U4798 , P2_R1212_U61 , P2_U3040 );
nand NAND2_5351 ( P2_U4799 , P2_U3039 , P2_U3433 );
nand NAND2_5352 ( P2_U4800 , P2_R1209_U61 , P2_U3037 );
nand NAND3_5353 ( P2_U4801 , P2_U4799 , P2_U4798 , P2_U4800 );
nand NAND2_5354 ( P2_U4802 , P2_R1054_U77 , P2_U3051 );
nand NAND2_5355 ( P2_U4803 , P2_U5764 , P2_U3433 );
nand NAND2_5356 ( P2_U4804 , P2_U3042 , P2_U4801 );
nand NAND2_5357 ( P2_U4805 , P2_R1212_U61 , P2_U3041 );
nand NAND2_5358 ( P2_U4806 , P2_REG3_REG_15_ , P2_U3151 );
nand NAND2_5359 ( P2_U4807 , P2_R1209_U61 , P2_U3038 );
nand NAND2_5360 ( P2_U4808 , P2_ADDR_REG_15_ , P2_U4756 );
nand NAND2_5361 ( P2_U4809 , P2_R1212_U62 , P2_U3040 );
nand NAND2_5362 ( P2_U4810 , P2_U3039 , P2_U3430 );
nand NAND2_5363 ( P2_U4811 , P2_R1209_U62 , P2_U3037 );
nand NAND3_5364 ( P2_U4812 , P2_U4810 , P2_U4809 , P2_U4811 );
nand NAND2_5365 ( P2_U4813 , P2_R1054_U78 , P2_U3051 );
nand NAND2_5366 ( P2_U4814 , P2_U5764 , P2_U3430 );
nand NAND2_5367 ( P2_U4815 , P2_U3042 , P2_U4812 );
nand NAND2_5368 ( P2_U4816 , P2_R1212_U62 , P2_U3041 );
nand NAND2_5369 ( P2_U4817 , P2_REG3_REG_14_ , P2_U3151 );
nand NAND2_5370 ( P2_U4818 , P2_R1209_U62 , P2_U3038 );
nand NAND2_5371 ( P2_U4819 , P2_ADDR_REG_14_ , P2_U4756 );
nand NAND2_5372 ( P2_U4820 , P2_R1212_U63 , P2_U3040 );
nand NAND2_5373 ( P2_U4821 , P2_U3039 , P2_U3427 );
nand NAND2_5374 ( P2_U4822 , P2_R1209_U63 , P2_U3037 );
nand NAND3_5375 ( P2_U4823 , P2_U4821 , P2_U4820 , P2_U4822 );
nand NAND2_5376 ( P2_U4824 , P2_R1054_U70 , P2_U3051 );
nand NAND2_5377 ( P2_U4825 , P2_U5764 , P2_U3427 );
nand NAND2_5378 ( P2_U4826 , P2_U3042 , P2_U4823 );
nand NAND2_5379 ( P2_U4827 , P2_R1212_U63 , P2_U3041 );
nand NAND2_5380 ( P2_U4828 , P2_REG3_REG_13_ , P2_U3151 );
nand NAND2_5381 ( P2_U4829 , P2_R1209_U63 , P2_U3038 );
nand NAND2_5382 ( P2_U4830 , P2_ADDR_REG_13_ , P2_U4756 );
nand NAND2_5383 ( P2_U4831 , P2_R1212_U64 , P2_U3040 );
nand NAND2_5384 ( P2_U4832 , P2_U3039 , P2_U3424 );
nand NAND2_5385 ( P2_U4833 , P2_R1209_U64 , P2_U3037 );
nand NAND3_5386 ( P2_U4834 , P2_U4832 , P2_U4831 , P2_U4833 );
nand NAND2_5387 ( P2_U4835 , P2_R1054_U71 , P2_U3051 );
nand NAND2_5388 ( P2_U4836 , P2_U5764 , P2_U3424 );
nand NAND2_5389 ( P2_U4837 , P2_U3042 , P2_U4834 );
nand NAND2_5390 ( P2_U4838 , P2_R1212_U64 , P2_U3041 );
nand NAND2_5391 ( P2_U4839 , P2_REG3_REG_12_ , P2_U3151 );
nand NAND2_5392 ( P2_U4840 , P2_R1209_U64 , P2_U3038 );
nand NAND2_5393 ( P2_U4841 , P2_ADDR_REG_12_ , P2_U4756 );
nand NAND2_5394 ( P2_U4842 , P2_R1212_U65 , P2_U3040 );
nand NAND2_5395 ( P2_U4843 , P2_U3039 , P2_U3421 );
nand NAND2_5396 ( P2_U4844 , P2_R1209_U65 , P2_U3037 );
nand NAND3_5397 ( P2_U4845 , P2_U4843 , P2_U4842 , P2_U4844 );
nand NAND2_5398 ( P2_U4846 , P2_R1054_U12 , P2_U3051 );
nand NAND2_5399 ( P2_U4847 , P2_U5764 , P2_U3421 );
nand NAND2_5400 ( P2_U4848 , P2_U3042 , P2_U4845 );
nand NAND2_5401 ( P2_U4849 , P2_R1212_U65 , P2_U3041 );
nand NAND2_5402 ( P2_U4850 , P2_REG3_REG_11_ , P2_U3151 );
nand NAND2_5403 ( P2_U4851 , P2_R1209_U65 , P2_U3038 );
nand NAND2_5404 ( P2_U4852 , P2_ADDR_REG_11_ , P2_U4756 );
nand NAND2_5405 ( P2_U4853 , P2_R1212_U66 , P2_U3040 );
nand NAND2_5406 ( P2_U4854 , P2_U3039 , P2_U3418 );
nand NAND2_5407 ( P2_U4855 , P2_R1209_U66 , P2_U3037 );
nand NAND3_5408 ( P2_U4856 , P2_U4854 , P2_U4853 , P2_U4855 );
nand NAND2_5409 ( P2_U4857 , P2_R1054_U79 , P2_U3051 );
nand NAND2_5410 ( P2_U4858 , P2_U5764 , P2_U3418 );
nand NAND2_5411 ( P2_U4859 , P2_U3042 , P2_U4856 );
nand NAND2_5412 ( P2_U4860 , P2_R1212_U66 , P2_U3041 );
nand NAND2_5413 ( P2_U4861 , P2_REG3_REG_10_ , P2_U3151 );
nand NAND2_5414 ( P2_U4862 , P2_R1209_U66 , P2_U3038 );
nand NAND2_5415 ( P2_U4863 , P2_ADDR_REG_10_ , P2_U4756 );
nand NAND2_5416 ( P2_U4864 , P2_R1212_U49 , P2_U3040 );
nand NAND2_5417 ( P2_U4865 , P2_U3039 , P2_U3415 );
nand NAND2_5418 ( P2_U4866 , P2_R1209_U49 , P2_U3037 );
nand NAND3_5419 ( P2_U4867 , P2_U4865 , P2_U4864 , P2_U4866 );
nand NAND2_5420 ( P2_U4868 , P2_R1054_U72 , P2_U3051 );
nand NAND2_5421 ( P2_U4869 , P2_U5764 , P2_U3415 );
nand NAND2_5422 ( P2_U4870 , P2_U3042 , P2_U4867 );
nand NAND2_5423 ( P2_U4871 , P2_R1212_U49 , P2_U3041 );
nand NAND2_5424 ( P2_U4872 , P2_REG3_REG_9_ , P2_U3151 );
nand NAND2_5425 ( P2_U4873 , P2_R1209_U49 , P2_U3038 );
nand NAND2_5426 ( P2_U4874 , P2_ADDR_REG_9_ , P2_U4756 );
nand NAND2_5427 ( P2_U4875 , P2_R1212_U50 , P2_U3040 );
nand NAND2_5428 ( P2_U4876 , P2_U3039 , P2_U3412 );
nand NAND2_5429 ( P2_U4877 , P2_R1209_U50 , P2_U3037 );
nand NAND3_5430 ( P2_U4878 , P2_U4876 , P2_U4875 , P2_U4877 );
nand NAND2_5431 ( P2_U4879 , P2_R1054_U16 , P2_U3051 );
nand NAND2_5432 ( P2_U4880 , P2_U5764 , P2_U3412 );
nand NAND2_5433 ( P2_U4881 , P2_U3042 , P2_U4878 );
nand NAND2_5434 ( P2_U4882 , P2_R1212_U50 , P2_U3041 );
nand NAND2_5435 ( P2_U4883 , P2_REG3_REG_8_ , P2_U3151 );
nand NAND2_5436 ( P2_U4884 , P2_R1209_U50 , P2_U3038 );
nand NAND2_5437 ( P2_U4885 , P2_ADDR_REG_8_ , P2_U4756 );
nand NAND2_5438 ( P2_U4886 , P2_R1212_U51 , P2_U3040 );
nand NAND2_5439 ( P2_U4887 , P2_U3039 , P2_U3409 );
nand NAND2_5440 ( P2_U4888 , P2_R1209_U51 , P2_U3037 );
nand NAND3_5441 ( P2_U4889 , P2_U4887 , P2_U4886 , P2_U4888 );
nand NAND2_5442 ( P2_U4890 , P2_R1054_U73 , P2_U3051 );
nand NAND2_5443 ( P2_U4891 , P2_U5764 , P2_U3409 );
nand NAND2_5444 ( P2_U4892 , P2_U3042 , P2_U4889 );
nand NAND2_5445 ( P2_U4893 , P2_R1212_U51 , P2_U3041 );
nand NAND2_5446 ( P2_U4894 , P2_REG3_REG_7_ , P2_U3151 );
nand NAND2_5447 ( P2_U4895 , P2_R1209_U51 , P2_U3038 );
nand NAND2_5448 ( P2_U4896 , P2_ADDR_REG_7_ , P2_U4756 );
nand NAND2_5449 ( P2_U4897 , P2_R1212_U52 , P2_U3040 );
nand NAND2_5450 ( P2_U4898 , P2_U3039 , P2_U3406 );
nand NAND2_5451 ( P2_U4899 , P2_R1209_U52 , P2_U3037 );
nand NAND3_5452 ( P2_U4900 , P2_U4898 , P2_U4897 , P2_U4899 );
nand NAND2_5453 ( P2_U4901 , P2_R1054_U15 , P2_U3051 );
nand NAND2_5454 ( P2_U4902 , P2_U5764 , P2_U3406 );
nand NAND2_5455 ( P2_U4903 , P2_U3042 , P2_U4900 );
nand NAND2_5456 ( P2_U4904 , P2_R1212_U52 , P2_U3041 );
nand NAND2_5457 ( P2_U4905 , P2_REG3_REG_6_ , P2_U3151 );
nand NAND2_5458 ( P2_U4906 , P2_R1209_U52 , P2_U3038 );
nand NAND2_5459 ( P2_U4907 , P2_ADDR_REG_6_ , P2_U4756 );
nand NAND2_5460 ( P2_U4908 , P2_R1212_U53 , P2_U3040 );
nand NAND2_5461 ( P2_U4909 , P2_U3039 , P2_U3403 );
nand NAND2_5462 ( P2_U4910 , P2_R1209_U53 , P2_U3037 );
nand NAND3_5463 ( P2_U4911 , P2_U4909 , P2_U4908 , P2_U4910 );
nand NAND2_5464 ( P2_U4912 , P2_R1054_U74 , P2_U3051 );
nand NAND2_5465 ( P2_U4913 , P2_U5764 , P2_U3403 );
nand NAND2_5466 ( P2_U4914 , P2_U3042 , P2_U4911 );
nand NAND2_5467 ( P2_U4915 , P2_R1212_U53 , P2_U3041 );
nand NAND2_5468 ( P2_U4916 , P2_REG3_REG_5_ , P2_U3151 );
nand NAND2_5469 ( P2_U4917 , P2_R1209_U53 , P2_U3038 );
nand NAND2_5470 ( P2_U4918 , P2_ADDR_REG_5_ , P2_U4756 );
nand NAND2_5471 ( P2_U4919 , P2_R1212_U54 , P2_U3040 );
nand NAND2_5472 ( P2_U4920 , P2_U3039 , P2_U3400 );
nand NAND2_5473 ( P2_U4921 , P2_R1209_U54 , P2_U3037 );
nand NAND3_5474 ( P2_U4922 , P2_U4920 , P2_U4919 , P2_U4921 );
nand NAND2_5475 ( P2_U4923 , P2_R1054_U75 , P2_U3051 );
nand NAND2_5476 ( P2_U4924 , P2_U5764 , P2_U3400 );
nand NAND2_5477 ( P2_U4925 , P2_U3042 , P2_U4922 );
nand NAND2_5478 ( P2_U4926 , P2_R1212_U54 , P2_U3041 );
nand NAND2_5479 ( P2_U4927 , P2_REG3_REG_4_ , P2_U3151 );
nand NAND2_5480 ( P2_U4928 , P2_R1209_U54 , P2_U3038 );
nand NAND2_5481 ( P2_U4929 , P2_ADDR_REG_4_ , P2_U4756 );
nand NAND2_5482 ( P2_U4930 , P2_R1212_U55 , P2_U3040 );
nand NAND2_5483 ( P2_U4931 , P2_U3039 , P2_U3397 );
nand NAND2_5484 ( P2_U4932 , P2_R1209_U55 , P2_U3037 );
nand NAND3_5485 ( P2_U4933 , P2_U4931 , P2_U4930 , P2_U4932 );
nand NAND2_5486 ( P2_U4934 , P2_R1054_U14 , P2_U3051 );
nand NAND2_5487 ( P2_U4935 , P2_U5764 , P2_U3397 );
nand NAND2_5488 ( P2_U4936 , P2_U3042 , P2_U4933 );
nand NAND2_5489 ( P2_U4937 , P2_R1212_U55 , P2_U3041 );
nand NAND2_5490 ( P2_U4938 , P2_REG3_REG_3_ , P2_U3151 );
nand NAND2_5491 ( P2_U4939 , P2_R1209_U55 , P2_U3038 );
nand NAND2_5492 ( P2_U4940 , P2_ADDR_REG_3_ , P2_U4756 );
nand NAND2_5493 ( P2_U4941 , P2_R1212_U56 , P2_U3040 );
nand NAND2_5494 ( P2_U4942 , P2_U3039 , P2_U3394 );
nand NAND2_5495 ( P2_U4943 , P2_R1209_U56 , P2_U3037 );
nand NAND3_5496 ( P2_U4944 , P2_U4942 , P2_U4941 , P2_U4943 );
nand NAND2_5497 ( P2_U4945 , P2_R1054_U76 , P2_U3051 );
nand NAND2_5498 ( P2_U4946 , P2_U5764 , P2_U3394 );
nand NAND2_5499 ( P2_U4947 , P2_U3042 , P2_U4944 );
nand NAND2_5500 ( P2_U4948 , P2_R1212_U56 , P2_U3041 );
nand NAND2_5501 ( P2_U4949 , P2_REG3_REG_2_ , P2_U3151 );
nand NAND2_5502 ( P2_U4950 , P2_R1209_U56 , P2_U3038 );
nand NAND2_5503 ( P2_U4951 , P2_ADDR_REG_2_ , P2_U4756 );
nand NAND2_5504 ( P2_U4952 , P2_R1212_U57 , P2_U3040 );
nand NAND2_5505 ( P2_U4953 , P2_U3039 , P2_U3391 );
nand NAND2_5506 ( P2_U4954 , P2_R1209_U57 , P2_U3037 );
nand NAND3_5507 ( P2_U4955 , P2_U4953 , P2_U4952 , P2_U4954 );
nand NAND2_5508 ( P2_U4956 , P2_R1054_U66 , P2_U3051 );
nand NAND2_5509 ( P2_U4957 , P2_U5764 , P2_U3391 );
nand NAND2_5510 ( P2_U4958 , P2_U3042 , P2_U4955 );
nand NAND2_5511 ( P2_U4959 , P2_R1212_U57 , P2_U3041 );
nand NAND2_5512 ( P2_U4960 , P2_REG3_REG_1_ , P2_U3151 );
nand NAND2_5513 ( P2_U4961 , P2_R1209_U57 , P2_U3038 );
nand NAND2_5514 ( P2_U4962 , P2_ADDR_REG_1_ , P2_U4756 );
nand NAND2_5515 ( P2_U4963 , P2_R1212_U7 , P2_U3040 );
nand NAND2_5516 ( P2_U4964 , P2_U3039 , P2_U3386 );
nand NAND2_5517 ( P2_U4965 , P2_R1209_U7 , P2_U3037 );
nand NAND3_5518 ( P2_U4966 , P2_U4964 , P2_U4963 , P2_U4965 );
nand NAND2_5519 ( P2_U4967 , P2_R1054_U17 , P2_U3051 );
nand NAND2_5520 ( P2_U4968 , P2_U5764 , P2_U3386 );
nand NAND2_5521 ( P2_U4969 , P2_U3042 , P2_U4966 );
nand NAND2_5522 ( P2_U4970 , P2_R1212_U7 , P2_U3041 );
nand NAND2_5523 ( P2_U4971 , P2_REG3_REG_0_ , P2_U3151 );
nand NAND2_5524 ( P2_U4972 , P2_R1209_U7 , P2_U3038 );
nand NAND2_5525 ( P2_U4973 , P2_ADDR_REG_0_ , P2_U4756 );
not NOT1_5526 ( P2_U4974 , P2_U3864 );
nand NAND3_5527 ( P2_U4975 , P2_U5938 , P2_U5937 , P2_U3050 );
nand NAND3_5528 ( P2_U4976 , P2_U3023 , P2_U3905 , P2_U3863 );
nand NAND2_5529 ( P2_U4977 , P2_B_REG , P2_U4975 );
nand NAND2_5530 ( P2_U4978 , P2_U3036 , P2_U3078 );
nand NAND2_5531 ( P2_U4979 , P2_U3032 , P2_U3072 );
nand NAND2_5532 ( P2_U4980 , P2_SUB_605_U21 , P2_U3304 );
nand NAND3_5533 ( P2_U4981 , P2_U4979 , P2_U4978 , P2_U4980 );
nand NAND5_5534 ( P2_U4982 , P2_U3311 , P2_U3871 , P2_U3884 , P2_U5421 , P2_U3312 );
nand NAND2_5535 ( P2_U4983 , P2_U3890 , P2_U4982 );
nand NAND2_5536 ( P2_U4984 , P2_U3885 , P2_U3891 );
nand NAND2_5537 ( P2_U4985 , P2_U4984 , P2_U4983 );
nand NAND2_5538 ( P2_U4986 , P2_U3907 , P2_U3378 );
nand NAND2_5539 ( P2_U4987 , P2_U3885 , P2_U3304 );
nand NAND2_5540 ( P2_U4988 , P2_U4982 , P2_U3303 );
not NOT1_5541 ( P2_U4989 , P2_U3370 );
nand NAND2_5542 ( P2_U4990 , P2_U3434 , P2_U5416 );
nand NAND2_5543 ( P2_U4991 , P2_SUB_605_U21 , P2_U3371 );
nand NAND2_5544 ( P2_U4992 , P2_R1158_U114 , P2_U3035 );
nand NAND2_5545 ( P2_U4993 , P2_U3031 , P2_U4981 );
nand NAND2_5546 ( P2_U4994 , P2_REG3_REG_15_ , P2_U3151 );
nand NAND2_5547 ( P2_U4995 , P2_U3036 , P2_U3057 );
nand NAND2_5548 ( P2_U4996 , P2_U3032 , P2_U3052 );
nand NAND2_5549 ( P2_U4997 , P2_SUB_605_U27 , P2_U3304 );
nand NAND3_5550 ( P2_U4998 , P2_U4996 , P2_U4995 , P2_U4997 );
nand NAND2_5551 ( P2_U4999 , P2_U3365 , P2_U3303 );
nand NAND2_5552 ( P2_U5000 , P2_U4989 , P2_U4999 );
nand NAND2_5553 ( P2_U5001 , P2_U3890 , P2_U3365 );
nand NAND2_5554 ( P2_U5002 , P2_U3360 , P2_U5001 );
nand NAND2_5555 ( P2_U5003 , P2_U3045 , P2_U3897 );
nand NAND2_5556 ( P2_U5004 , P2_U3044 , P2_SUB_605_U27 );
nand NAND2_5557 ( P2_U5005 , P2_R1158_U17 , P2_U3035 );
nand NAND2_5558 ( P2_U5006 , P2_U3031 , P2_U4998 );
nand NAND2_5559 ( P2_U5007 , P2_REG3_REG_26_ , P2_U3151 );
nand NAND2_5560 ( P2_U5008 , P2_U3036 , P2_U3066 );
nand NAND2_5561 ( P2_U5009 , P2_U3032 , P2_U3069 );
nand NAND2_5562 ( P2_U5010 , P2_SUB_605_U8 , P2_U3304 );
nand NAND3_5563 ( P2_U5011 , P2_U5009 , P2_U5008 , P2_U5010 );
nand NAND2_5564 ( P2_U5012 , P2_U3407 , P2_U5416 );
nand NAND2_5565 ( P2_U5013 , P2_SUB_605_U8 , P2_U3371 );
nand NAND2_5566 ( P2_U5014 , P2_R1158_U99 , P2_U3035 );
nand NAND2_5567 ( P2_U5015 , P2_U3031 , P2_U5011 );
nand NAND2_5568 ( P2_U5016 , P2_REG3_REG_6_ , P2_U3151 );
nand NAND2_5569 ( P2_U5017 , P2_U3036 , P2_U3068 );
nand NAND2_5570 ( P2_U5018 , P2_U3032 , P2_U3080 );
nand NAND2_5571 ( P2_U5019 , P2_SUB_605_U11 , P2_U3304 );
nand NAND3_5572 ( P2_U5020 , P2_U5018 , P2_U5017 , P2_U5019 );
nand NAND2_5573 ( P2_U5021 , P2_U3443 , P2_U5416 );
nand NAND2_5574 ( P2_U5022 , P2_SUB_605_U11 , P2_U3371 );
nand NAND2_5575 ( P2_U5023 , P2_R1158_U112 , P2_U3035 );
nand NAND2_5576 ( P2_U5024 , P2_U3031 , P2_U5020 );
nand NAND2_5577 ( P2_U5025 , P2_REG3_REG_18_ , P2_U3151 );
nand NAND2_5578 ( P2_U5026 , P2_U3036 , P2_U3077 );
nand NAND2_5579 ( P2_U5027 , P2_U3032 , P2_U3063 );
nand NAND2_5580 ( P2_U5028 , P2_REG3_REG_2_ , P2_U3304 );
nand NAND3_5581 ( P2_U5029 , P2_U5027 , P2_U5026 , P2_U5028 );
nand NAND2_5582 ( P2_U5030 , P2_U3395 , P2_U5416 );
nand NAND2_5583 ( P2_U5031 , P2_REG3_REG_2_ , P2_U3371 );
nand NAND2_5584 ( P2_U5032 , P2_R1158_U102 , P2_U3035 );
nand NAND2_5585 ( P2_U5033 , P2_U3031 , P2_U5029 );
nand NAND2_5586 ( P2_U5034 , P2_REG3_REG_2_ , P2_U3151 );
nand NAND2_5587 ( P2_U5035 , P2_U3036 , P2_U3061 );
nand NAND2_5588 ( P2_U5036 , P2_U3032 , P2_U3071 );
nand NAND2_5589 ( P2_U5037 , P2_SUB_605_U9 , P2_U3304 );
nand NAND3_5590 ( P2_U5038 , P2_U5036 , P2_U5035 , P2_U5037 );
nand NAND2_5591 ( P2_U5039 , P2_U3422 , P2_U5416 );
nand NAND2_5592 ( P2_U5040 , P2_SUB_605_U9 , P2_U3371 );
nand NAND2_5593 ( P2_U5041 , P2_R1158_U117 , P2_U3035 );
nand NAND2_5594 ( P2_U5042 , P2_U3031 , P2_U5038 );
nand NAND2_5595 ( P2_U5043 , P2_REG3_REG_11_ , P2_U3151 );
nand NAND2_5596 ( P2_U5044 , P2_U3036 , P2_U3074 );
nand NAND2_5597 ( P2_U5045 , P2_U3032 , P2_U3065 );
nand NAND2_5598 ( P2_U5046 , P2_SUB_605_U17 , P2_U3304 );
nand NAND3_5599 ( P2_U5047 , P2_U5045 , P2_U5044 , P2_U5046 );
nand NAND2_5600 ( P2_U5048 , P2_U3045 , P2_U3901 );
nand NAND2_5601 ( P2_U5049 , P2_U3044 , P2_SUB_605_U17 );
nand NAND2_5602 ( P2_U5050 , P2_R1158_U108 , P2_U3035 );
nand NAND2_5603 ( P2_U5051 , P2_U3031 , P2_U5047 );
nand NAND2_5604 ( P2_U5052 , P2_REG3_REG_22_ , P2_U3151 );
nand NAND2_5605 ( P2_U5053 , P2_U3036 , P2_U3071 );
nand NAND2_5606 ( P2_U5054 , P2_U3032 , P2_U3078 );
nand NAND2_5607 ( P2_U5055 , P2_SUB_605_U25 , P2_U3304 );
nand NAND3_5608 ( P2_U5056 , P2_U5054 , P2_U5053 , P2_U5055 );
nand NAND2_5609 ( P2_U5057 , P2_U3428 , P2_U5416 );
nand NAND2_5610 ( P2_U5058 , P2_SUB_605_U25 , P2_U3371 );
nand NAND2_5611 ( P2_U5059 , P2_R1158_U14 , P2_U3035 );
nand NAND2_5612 ( P2_U5060 , P2_U3031 , P2_U5056 );
nand NAND2_5613 ( P2_U5061 , P2_REG3_REG_13_ , P2_U3151 );
nand NAND2_5614 ( P2_U5062 , P2_U3036 , P2_U3080 );
nand NAND2_5615 ( P2_U5063 , P2_U3032 , P2_U3074 );
nand NAND2_5616 ( P2_U5064 , P2_SUB_605_U20 , P2_U3304 );
nand NAND3_5617 ( P2_U5065 , P2_U5063 , P2_U5062 , P2_U5064 );
nand NAND2_5618 ( P2_U5066 , P2_U3045 , P2_U3903 );
nand NAND2_5619 ( P2_U5067 , P2_U3044 , P2_SUB_605_U20 );
nand NAND2_5620 ( P2_U5068 , P2_R1158_U109 , P2_U3035 );
nand NAND2_5621 ( P2_U5069 , P2_U3031 , P2_U5065 );
nand NAND2_5622 ( P2_U5070 , P2_REG3_REG_20_ , P2_U3151 );
nand NAND2_5623 ( P2_U5071 , P2_U3031 , P2_U3304 );
nand NAND2_5624 ( P2_U5072 , P2_U5415 , P2_U5071 );
nand NAND2_5625 ( P2_U5073 , P2_U3792 , P2_U3032 );
nand NAND2_5626 ( P2_U5074 , P2_U3387 , P2_U5416 );
nand NAND2_5627 ( P2_U5075 , P2_REG3_REG_0_ , P2_U5072 );
nand NAND2_5628 ( P2_U5076 , P2_R1158_U96 , P2_U3035 );
nand NAND2_5629 ( P2_U5077 , P2_REG3_REG_0_ , P2_U3151 );
nand NAND2_5630 ( P2_U5078 , P2_U3036 , P2_U3083 );
nand NAND2_5631 ( P2_U5079 , P2_U3032 , P2_U3061 );
nand NAND2_5632 ( P2_U5080 , P2_SUB_605_U14 , P2_U3304 );
nand NAND3_5633 ( P2_U5081 , P2_U5079 , P2_U5078 , P2_U5080 );
nand NAND2_5634 ( P2_U5082 , P2_U3416 , P2_U5416 );
nand NAND2_5635 ( P2_U5083 , P2_SUB_605_U14 , P2_U3371 );
nand NAND2_5636 ( P2_U5084 , P2_R1158_U97 , P2_U3035 );
nand NAND2_5637 ( P2_U5085 , P2_U3031 , P2_U5081 );
nand NAND2_5638 ( P2_U5086 , P2_REG3_REG_9_ , P2_U3151 );
nand NAND2_5639 ( P2_U5087 , P2_U3036 , P2_U3063 );
nand NAND2_5640 ( P2_U5088 , P2_U3032 , P2_U3066 );
nand NAND2_5641 ( P2_U5089 , P2_SUB_605_U30 , P2_U3304 );
nand NAND3_5642 ( P2_U5090 , P2_U5088 , P2_U5087 , P2_U5089 );
nand NAND2_5643 ( P2_U5091 , P2_U3401 , P2_U5416 );
nand NAND2_5644 ( P2_U5092 , P2_SUB_605_U30 , P2_U3371 );
nand NAND2_5645 ( P2_U5093 , P2_R1158_U101 , P2_U3035 );
nand NAND2_5646 ( P2_U5094 , P2_U3031 , P2_U5090 );
nand NAND2_5647 ( P2_U5095 , P2_REG3_REG_4_ , P2_U3151 );
nand NAND2_5648 ( P2_U5096 , P2_U3036 , P2_U3065 );
nand NAND2_5649 ( P2_U5097 , P2_U3032 , P2_U3057 );
nand NAND2_5650 ( P2_U5098 , P2_SUB_605_U10 , P2_U3304 );
nand NAND3_5651 ( P2_U5099 , P2_U5097 , P2_U5096 , P2_U5098 );
nand NAND2_5652 ( P2_U5100 , P2_U3045 , P2_U3899 );
nand NAND2_5653 ( P2_U5101 , P2_U3044 , P2_SUB_605_U10 );
nand NAND2_5654 ( P2_U5102 , P2_R1158_U106 , P2_U3035 );
nand NAND2_5655 ( P2_U5103 , P2_U3031 , P2_U5099 );
nand NAND2_5656 ( P2_U5104 , P2_REG3_REG_24_ , P2_U3151 );
nand NAND2_5657 ( P2_U5105 , P2_U3036 , P2_U3072 );
nand NAND2_5658 ( P2_U5106 , P2_U3032 , P2_U3081 );
nand NAND2_5659 ( P2_U5107 , P2_SUB_605_U19 , P2_U3304 );
nand NAND3_5660 ( P2_U5108 , P2_U5106 , P2_U5105 , P2_U5107 );
nand NAND2_5661 ( P2_U5109 , P2_U3440 , P2_U5416 );
nand NAND2_5662 ( P2_U5110 , P2_SUB_605_U19 , P2_U3371 );
nand NAND2_5663 ( P2_U5111 , P2_R1158_U15 , P2_U3035 );
nand NAND2_5664 ( P2_U5112 , P2_U3031 , P2_U5108 );
nand NAND2_5665 ( P2_U5113 , P2_REG3_REG_17_ , P2_U3151 );
nand NAND2_5666 ( P2_U5114 , P2_U3036 , P2_U3059 );
nand NAND2_5667 ( P2_U5115 , P2_U3032 , P2_U3070 );
nand NAND2_5668 ( P2_U5116 , P2_SUB_605_U22 , P2_U3304 );
nand NAND3_5669 ( P2_U5117 , P2_U5115 , P2_U5114 , P2_U5116 );
nand NAND2_5670 ( P2_U5118 , P2_U3404 , P2_U5416 );
nand NAND2_5671 ( P2_U5119 , P2_SUB_605_U22 , P2_U3371 );
nand NAND2_5672 ( P2_U5120 , P2_R1158_U100 , P2_U3035 );
nand NAND2_5673 ( P2_U5121 , P2_U3031 , P2_U5117 );
nand NAND2_5674 ( P2_U5122 , P2_REG3_REG_5_ , P2_U3151 );
nand NAND2_5675 ( P2_U5123 , P2_U3036 , P2_U3073 );
nand NAND2_5676 ( P2_U5124 , P2_U3032 , P2_U3068 );
nand NAND2_5677 ( P2_U5125 , P2_SUB_605_U7 , P2_U3304 );
nand NAND3_5678 ( P2_U5126 , P2_U5124 , P2_U5123 , P2_U5125 );
nand NAND2_5679 ( P2_U5127 , P2_U3437 , P2_U5416 );
nand NAND2_5680 ( P2_U5128 , P2_SUB_605_U7 , P2_U3371 );
nand NAND2_5681 ( P2_U5129 , P2_R1158_U113 , P2_U3035 );
nand NAND2_5682 ( P2_U5130 , P2_U3031 , P2_U5126 );
nand NAND2_5683 ( P2_U5131 , P2_REG3_REG_16_ , P2_U3151 );
nand NAND2_5684 ( P2_U5132 , P2_U3036 , P2_U3064 );
nand NAND2_5685 ( P2_U5133 , P2_U3032 , P2_U3056 );
nand NAND2_5686 ( P2_U5134 , P2_SUB_605_U16 , P2_U3304 );
nand NAND3_5687 ( P2_U5135 , P2_U5133 , P2_U5132 , P2_U5134 );
nand NAND2_5688 ( P2_U5136 , P2_U3045 , P2_U3898 );
nand NAND2_5689 ( P2_U5137 , P2_U3044 , P2_SUB_605_U16 );
nand NAND2_5690 ( P2_U5138 , P2_R1158_U105 , P2_U3035 );
nand NAND2_5691 ( P2_U5139 , P2_U3031 , P2_U5135 );
nand NAND2_5692 ( P2_U5140 , P2_REG3_REG_25_ , P2_U3151 );
nand NAND2_5693 ( P2_U5141 , P2_U3036 , P2_U3062 );
nand NAND2_5694 ( P2_U5142 , P2_U3032 , P2_U3079 );
nand NAND2_5695 ( P2_U5143 , P2_SUB_605_U24 , P2_U3304 );
nand NAND3_5696 ( P2_U5144 , P2_U5142 , P2_U5141 , P2_U5143 );
nand NAND2_5697 ( P2_U5145 , P2_U3425 , P2_U5416 );
nand NAND2_5698 ( P2_U5146 , P2_SUB_605_U24 , P2_U3371 );
nand NAND2_5699 ( P2_U5147 , P2_R1158_U116 , P2_U3035 );
nand NAND2_5700 ( P2_U5148 , P2_U3031 , P2_U5144 );
nand NAND2_5701 ( P2_U5149 , P2_REG3_REG_12_ , P2_U3151 );
nand NAND2_5702 ( P2_U5150 , P2_U3036 , P2_U3075 );
nand NAND2_5703 ( P2_U5151 , P2_U3032 , P2_U3060 );
nand NAND2_5704 ( P2_U5152 , P2_SUB_605_U28 , P2_U3304 );
nand NAND3_5705 ( P2_U5153 , P2_U5151 , P2_U5150 , P2_U5152 );
nand NAND2_5706 ( P2_U5154 , P2_U3045 , P2_U3902 );
nand NAND2_5707 ( P2_U5155 , P2_U3044 , P2_SUB_605_U28 );
nand NAND2_5708 ( P2_U5156 , P2_R1158_U16 , P2_U3035 );
nand NAND2_5709 ( P2_U5157 , P2_U3031 , P2_U5153 );
nand NAND2_5710 ( P2_U5158 , P2_REG3_REG_21_ , P2_U3151 );
nand NAND2_5711 ( P2_U5159 , P2_U3036 , P2_U3076 );
nand NAND2_5712 ( P2_U5160 , P2_U3032 , P2_U3067 );
nand NAND2_5713 ( P2_U5161 , P2_REG3_REG_1_ , P2_U3304 );
nand NAND3_5714 ( P2_U5162 , P2_U5160 , P2_U5159 , P2_U5161 );
nand NAND2_5715 ( P2_U5163 , P2_U3392 , P2_U5416 );
nand NAND2_5716 ( P2_U5164 , P2_REG3_REG_1_ , P2_U3371 );
nand NAND2_5717 ( P2_U5165 , P2_R1158_U110 , P2_U3035 );
nand NAND2_5718 ( P2_U5166 , P2_U3031 , P2_U5162 );
nand NAND2_5719 ( P2_U5167 , P2_REG3_REG_1_ , P2_U3151 );
nand NAND2_5720 ( P2_U5168 , P2_U3036 , P2_U3069 );
nand NAND2_5721 ( P2_U5169 , P2_U3032 , P2_U3082 );
nand NAND2_5722 ( P2_U5170 , P2_SUB_605_U12 , P2_U3304 );
nand NAND3_5723 ( P2_U5171 , P2_U5169 , P2_U5168 , P2_U5170 );
nand NAND2_5724 ( P2_U5172 , P2_U3413 , P2_U5416 );
nand NAND2_5725 ( P2_U5173 , P2_SUB_605_U12 , P2_U3371 );
nand NAND2_5726 ( P2_U5174 , P2_R1158_U98 , P2_U3035 );
nand NAND2_5727 ( P2_U5175 , P2_U3031 , P2_U5171 );
nand NAND2_5728 ( P2_U5176 , P2_REG3_REG_8_ , P2_U3151 );
nand NAND2_5729 ( P2_U5177 , P2_U3036 , P2_U3052 );
nand NAND2_5730 ( P2_U5178 , P2_U3032 , P2_U3054 );
nand NAND2_5731 ( P2_U5179 , P2_SUB_605_U29 , P2_U3304 );
nand NAND3_5732 ( P2_U5180 , P2_U5178 , P2_U5177 , P2_U5179 );
nand NAND2_5733 ( P2_U5181 , P2_U3045 , P2_U3895 );
nand NAND2_5734 ( P2_U5182 , P2_U3044 , P2_SUB_605_U29 );
nand NAND2_5735 ( P2_U5183 , P2_R1158_U103 , P2_U3035 );
nand NAND2_5736 ( P2_U5184 , P2_U3031 , P2_U5180 );
nand NAND2_5737 ( P2_U5185 , P2_REG3_REG_28_ , P2_U3151 );
nand NAND2_5738 ( P2_U5186 , P2_U3036 , P2_U3081 );
nand NAND2_5739 ( P2_U5187 , P2_U3032 , P2_U3075 );
nand NAND2_5740 ( P2_U5188 , P2_SUB_605_U15 , P2_U3304 );
nand NAND3_5741 ( P2_U5189 , P2_U5187 , P2_U5186 , P2_U5188 );
nand NAND2_5742 ( P2_U5190 , P2_U3445 , P2_U5416 );
nand NAND2_5743 ( P2_U5191 , P2_SUB_605_U15 , P2_U3371 );
nand NAND2_5744 ( P2_U5192 , P2_R1158_U111 , P2_U3035 );
nand NAND2_5745 ( P2_U5193 , P2_U3031 , P2_U5189 );
nand NAND2_5746 ( P2_U5194 , P2_REG3_REG_19_ , P2_U3151 );
nand NAND2_5747 ( P2_U5195 , P2_U3036 , P2_U3067 );
nand NAND2_5748 ( P2_U5196 , P2_U3032 , P2_U3059 );
nand NAND2_5749 ( P2_U5197 , P2_SUB_605_U26 , P2_U3304 );
nand NAND3_5750 ( P2_U5198 , P2_U5196 , P2_U5195 , P2_U5197 );
nand NAND2_5751 ( P2_U5199 , P2_U3398 , P2_U5416 );
nand NAND2_5752 ( P2_U5200 , P2_SUB_605_U26 , P2_U3371 );
nand NAND2_5753 ( P2_U5201 , P2_R1158_U18 , P2_U3035 );
nand NAND2_5754 ( P2_U5202 , P2_U3031 , P2_U5198 );
nand NAND2_5755 ( P2_U5203 , P2_REG3_REG_3_ , P2_U3151 );
nand NAND2_5756 ( P2_U5204 , P2_U3036 , P2_U3082 );
nand NAND2_5757 ( P2_U5205 , P2_U3032 , P2_U3062 );
nand NAND2_5758 ( P2_U5206 , P2_SUB_605_U13 , P2_U3304 );
nand NAND3_5759 ( P2_U5207 , P2_U5205 , P2_U5204 , P2_U5206 );
nand NAND2_5760 ( P2_U5208 , P2_U3419 , P2_U5416 );
nand NAND2_5761 ( P2_U5209 , P2_SUB_605_U13 , P2_U3371 );
nand NAND2_5762 ( P2_U5210 , P2_R1158_U118 , P2_U3035 );
nand NAND2_5763 ( P2_U5211 , P2_U3031 , P2_U5207 );
nand NAND2_5764 ( P2_U5212 , P2_REG3_REG_10_ , P2_U3151 );
nand NAND2_5765 ( P2_U5213 , P2_U3036 , P2_U3060 );
nand NAND2_5766 ( P2_U5214 , P2_U3032 , P2_U3064 );
nand NAND2_5767 ( P2_U5215 , P2_SUB_605_U6 , P2_U3304 );
nand NAND3_5768 ( P2_U5216 , P2_U5214 , P2_U5213 , P2_U5215 );
nand NAND2_5769 ( P2_U5217 , P2_U3045 , P2_U3900 );
nand NAND2_5770 ( P2_U5218 , P2_U3044 , P2_SUB_605_U6 );
nand NAND2_5771 ( P2_U5219 , P2_R1158_U107 , P2_U3035 );
nand NAND2_5772 ( P2_U5220 , P2_U3031 , P2_U5216 );
nand NAND2_5773 ( P2_U5221 , P2_REG3_REG_23_ , P2_U3151 );
nand NAND2_5774 ( P2_U5222 , P2_U3036 , P2_U3079 );
nand NAND2_5775 ( P2_U5223 , P2_U3032 , P2_U3073 );
nand NAND2_5776 ( P2_U5224 , P2_SUB_605_U31 , P2_U3304 );
nand NAND3_5777 ( P2_U5225 , P2_U5223 , P2_U5222 , P2_U5224 );
nand NAND2_5778 ( P2_U5226 , P2_U3431 , P2_U5416 );
nand NAND2_5779 ( P2_U5227 , P2_SUB_605_U31 , P2_U3371 );
nand NAND2_5780 ( P2_U5228 , P2_R1158_U115 , P2_U3035 );
nand NAND2_5781 ( P2_U5229 , P2_U3031 , P2_U5225 );
nand NAND2_5782 ( P2_U5230 , P2_REG3_REG_14_ , P2_U3151 );
nand NAND2_5783 ( P2_U5231 , P2_U3036 , P2_U3056 );
nand NAND2_5784 ( P2_U5232 , P2_U3032 , P2_U3053 );
nand NAND2_5785 ( P2_U5233 , P2_SUB_605_U23 , P2_U3304 );
nand NAND3_5786 ( P2_U5234 , P2_U5232 , P2_U5231 , P2_U5233 );
nand NAND2_5787 ( P2_U5235 , P2_U3045 , P2_U3896 );
nand NAND2_5788 ( P2_U5236 , P2_U3044 , P2_SUB_605_U23 );
nand NAND2_5789 ( P2_U5237 , P2_R1158_U104 , P2_U3035 );
nand NAND2_5790 ( P2_U5238 , P2_U3031 , P2_U5234 );
nand NAND2_5791 ( P2_U5239 , P2_REG3_REG_27_ , P2_U3151 );
nand NAND2_5792 ( P2_U5240 , P2_U3036 , P2_U3070 );
nand NAND2_5793 ( P2_U5241 , P2_U3032 , P2_U3083 );
nand NAND2_5794 ( P2_U5242 , P2_SUB_605_U18 , P2_U3304 );
nand NAND3_5795 ( P2_U5243 , P2_U5241 , P2_U5240 , P2_U5242 );
nand NAND2_5796 ( P2_U5244 , P2_U3410 , P2_U5416 );
nand NAND2_5797 ( P2_U5245 , P2_SUB_605_U18 , P2_U3371 );
nand NAND2_5798 ( P2_U5246 , P2_R1158_U19 , P2_U3035 );
nand NAND2_5799 ( P2_U5247 , P2_U3031 , P2_U5243 );
nand NAND2_5800 ( P2_U5248 , P2_REG3_REG_7_ , P2_U3151 );
nand NAND2_5801 ( P2_U5249 , P2_U3894 , P2_U3046 );
nand NAND2_5802 ( P2_U5250 , P2_U3375 , P2_U3829 );
nand NAND2_5803 ( P2_U5251 , P2_U3821 , P2_U3820 );
nand NAND2_5804 ( P2_U5252 , P2_U3819 , P2_U3013 );
nand NAND2_5805 ( P2_U5253 , P2_U3876 , P2_U5252 );
nand NAND2_5806 ( P2_U5254 , P2_U3416 , P2_U5253 );
nand NAND2_5807 ( P2_U5255 , P2_U5251 , P2_U3082 );
nand NAND2_5808 ( P2_U5256 , P2_U3413 , P2_U5253 );
nand NAND2_5809 ( P2_U5257 , P2_U5251 , P2_U3083 );
nand NAND2_5810 ( P2_U5258 , P2_U3410 , P2_U5253 );
nand NAND2_5811 ( P2_U5259 , P2_U5251 , P2_U3069 );
nand NAND2_5812 ( P2_U5260 , P2_U3407 , P2_U5253 );
nand NAND2_5813 ( P2_U5261 , P2_U5251 , P2_U3070 );
nand NAND2_5814 ( P2_U5262 , P2_U3404 , P2_U5253 );
nand NAND2_5815 ( P2_U5263 , P2_U5251 , P2_U3066 );
nand NAND2_5816 ( P2_U5264 , P2_U3401 , P2_U5253 );
nand NAND2_5817 ( P2_U5265 , P2_U5251 , P2_U3059 );
nand NAND2_5818 ( P2_U5266 , P2_U3868 , P2_U5253 );
nand NAND2_5819 ( P2_U5267 , P2_U5251 , P2_U3055 );
nand NAND2_5820 ( P2_U5268 , P2_U3869 , P2_U5253 );
nand NAND2_5821 ( P2_U5269 , P2_U5251 , P2_U3058 );
nand NAND2_5822 ( P2_U5270 , P2_U3398 , P2_U5253 );
nand NAND2_5823 ( P2_U5271 , P2_U5251 , P2_U3063 );
nand NAND2_5824 ( P2_U5272 , P2_U3904 , P2_U5253 );
nand NAND2_5825 ( P2_U5273 , P2_U5251 , P2_U3054 );
nand NAND2_5826 ( P2_U5274 , P2_U3895 , P2_U5253 );
nand NAND2_5827 ( P2_U5275 , P2_U5251 , P2_U3053 );
nand NAND2_5828 ( P2_U5276 , P2_U3896 , P2_U5253 );
nand NAND2_5829 ( P2_U5277 , P2_U5251 , P2_U3052 );
nand NAND2_5830 ( P2_U5278 , P2_U3897 , P2_U5253 );
nand NAND2_5831 ( P2_U5279 , P2_U5251 , P2_U3056 );
nand NAND2_5832 ( P2_U5280 , P2_U3898 , P2_U5253 );
nand NAND2_5833 ( P2_U5281 , P2_U5251 , P2_U3057 );
nand NAND2_5834 ( P2_U5282 , P2_U3899 , P2_U5253 );
nand NAND2_5835 ( P2_U5283 , P2_U5251 , P2_U3064 );
nand NAND2_5836 ( P2_U5284 , P2_U3900 , P2_U5253 );
nand NAND2_5837 ( P2_U5285 , P2_U5251 , P2_U3065 );
nand NAND2_5838 ( P2_U5286 , P2_U3901 , P2_U5253 );
nand NAND2_5839 ( P2_U5287 , P2_U5251 , P2_U3060 );
nand NAND2_5840 ( P2_U5288 , P2_U3902 , P2_U5253 );
nand NAND2_5841 ( P2_U5289 , P2_U5251 , P2_U3074 );
nand NAND2_5842 ( P2_U5290 , P2_U3903 , P2_U5253 );
nand NAND2_5843 ( P2_U5291 , P2_U5251 , P2_U3075 );
nand NAND2_5844 ( P2_U5292 , P2_U3395 , P2_U5253 );
nand NAND2_5845 ( P2_U5293 , P2_U5251 , P2_U3067 );
nand NAND2_5846 ( P2_U5294 , P2_U3445 , P2_U5253 );
nand NAND2_5847 ( P2_U5295 , P2_U5251 , P2_U3080 );
nand NAND2_5848 ( P2_U5296 , P2_U3443 , P2_U5253 );
nand NAND2_5849 ( P2_U5297 , P2_U5251 , P2_U3081 );
nand NAND2_5850 ( P2_U5298 , P2_U3440 , P2_U5253 );
nand NAND2_5851 ( P2_U5299 , P2_U5251 , P2_U3068 );
nand NAND2_5852 ( P2_U5300 , P2_U3437 , P2_U5253 );
nand NAND2_5853 ( P2_U5301 , P2_U5251 , P2_U3072 );
nand NAND2_5854 ( P2_U5302 , P2_U3434 , P2_U5253 );
nand NAND2_5855 ( P2_U5303 , P2_U5251 , P2_U3073 );
nand NAND2_5856 ( P2_U5304 , P2_U3431 , P2_U5253 );
nand NAND2_5857 ( P2_U5305 , P2_U5251 , P2_U3078 );
nand NAND2_5858 ( P2_U5306 , P2_U3428 , P2_U5253 );
nand NAND2_5859 ( P2_U5307 , P2_U5251 , P2_U3079 );
nand NAND2_5860 ( P2_U5308 , P2_U3425 , P2_U5253 );
nand NAND2_5861 ( P2_U5309 , P2_U5251 , P2_U3071 );
nand NAND2_5862 ( P2_U5310 , P2_U3422 , P2_U5253 );
nand NAND2_5863 ( P2_U5311 , P2_U5251 , P2_U3062 );
nand NAND2_5864 ( P2_U5312 , P2_U3419 , P2_U5253 );
nand NAND2_5865 ( P2_U5313 , P2_U5251 , P2_U3061 );
nand NAND2_5866 ( P2_U5314 , P2_U3392 , P2_U5253 );
nand NAND2_5867 ( P2_U5315 , P2_U5251 , P2_U3077 );
nand NAND2_5868 ( P2_U5316 , P2_U3387 , P2_U5253 );
nand NAND2_5869 ( P2_U5317 , P2_U5251 , P2_U3076 );
nand NAND2_5870 ( P2_U5318 , P2_U3416 , P2_U5251 );
nand NAND2_5871 ( P2_U5319 , P2_U5253 , P2_U3082 );
nand NAND2_5872 ( P2_U5320 , P2_U5436 , P2_U3083 );
nand NAND2_5873 ( P2_U5321 , P2_U3413 , P2_U5251 );
nand NAND2_5874 ( P2_U5322 , P2_U5253 , P2_U3083 );
nand NAND2_5875 ( P2_U5323 , P2_U5436 , P2_U3069 );
nand NAND2_5876 ( P2_U5324 , P2_U3410 , P2_U5251 );
nand NAND2_5877 ( P2_U5325 , P2_U5253 , P2_U3069 );
nand NAND2_5878 ( P2_U5326 , P2_U5436 , P2_U3070 );
nand NAND2_5879 ( P2_U5327 , P2_U3407 , P2_U5251 );
nand NAND2_5880 ( P2_U5328 , P2_U5253 , P2_U3070 );
nand NAND2_5881 ( P2_U5329 , P2_U5436 , P2_U3066 );
nand NAND2_5882 ( P2_U5330 , P2_U3404 , P2_U5251 );
nand NAND2_5883 ( P2_U5331 , P2_U5253 , P2_U3066 );
nand NAND2_5884 ( P2_U5332 , P2_U5436 , P2_U3059 );
nand NAND2_5885 ( P2_U5333 , P2_U3401 , P2_U5251 );
nand NAND2_5886 ( P2_U5334 , P2_U5253 , P2_U3059 );
nand NAND2_5887 ( P2_U5335 , P2_U5436 , P2_U3063 );
nand NAND2_5888 ( P2_U5336 , P2_U5253 , P2_U3055 );
nand NAND2_5889 ( P2_U5337 , P2_U3868 , P2_U5251 );
nand NAND2_5890 ( P2_U5338 , P2_U5253 , P2_U3058 );
nand NAND2_5891 ( P2_U5339 , P2_U3869 , P2_U5251 );
nand NAND2_5892 ( P2_U5340 , P2_U3398 , P2_U5251 );
nand NAND2_5893 ( P2_U5341 , P2_U5253 , P2_U3063 );
nand NAND2_5894 ( P2_U5342 , P2_U5436 , P2_U3067 );
nand NAND2_5895 ( P2_U5343 , P2_U5253 , P2_U3054 );
nand NAND2_5896 ( P2_U5344 , P2_U3904 , P2_U5251 );
nand NAND2_5897 ( P2_U5345 , P2_U5436 , P2_U3053 );
nand NAND2_5898 ( P2_U5346 , P2_U5253 , P2_U3053 );
nand NAND2_5899 ( P2_U5347 , P2_U3895 , P2_U5251 );
nand NAND2_5900 ( P2_U5348 , P2_U5436 , P2_U3052 );
nand NAND2_5901 ( P2_U5349 , P2_U5253 , P2_U3052 );
nand NAND2_5902 ( P2_U5350 , P2_U3896 , P2_U5251 );
nand NAND2_5903 ( P2_U5351 , P2_U5436 , P2_U3056 );
nand NAND2_5904 ( P2_U5352 , P2_U5253 , P2_U3056 );
nand NAND2_5905 ( P2_U5353 , P2_U3897 , P2_U5251 );
nand NAND2_5906 ( P2_U5354 , P2_U5436 , P2_U3057 );
nand NAND2_5907 ( P2_U5355 , P2_U5253 , P2_U3057 );
nand NAND2_5908 ( P2_U5356 , P2_U3898 , P2_U5251 );
nand NAND2_5909 ( P2_U5357 , P2_U5436 , P2_U3064 );
nand NAND2_5910 ( P2_U5358 , P2_U5253 , P2_U3064 );
nand NAND2_5911 ( P2_U5359 , P2_U3899 , P2_U5251 );
nand NAND2_5912 ( P2_U5360 , P2_U5436 , P2_U3065 );
nand NAND2_5913 ( P2_U5361 , P2_U5253 , P2_U3065 );
nand NAND2_5914 ( P2_U5362 , P2_U3900 , P2_U5251 );
nand NAND2_5915 ( P2_U5363 , P2_U5436 , P2_U3060 );
nand NAND2_5916 ( P2_U5364 , P2_U5253 , P2_U3060 );
nand NAND2_5917 ( P2_U5365 , P2_U3901 , P2_U5251 );
nand NAND2_5918 ( P2_U5366 , P2_U5436 , P2_U3074 );
nand NAND2_5919 ( P2_U5367 , P2_U5253 , P2_U3074 );
nand NAND2_5920 ( P2_U5368 , P2_U3902 , P2_U5251 );
nand NAND2_5921 ( P2_U5369 , P2_U5436 , P2_U3075 );
nand NAND2_5922 ( P2_U5370 , P2_U5253 , P2_U3075 );
nand NAND2_5923 ( P2_U5371 , P2_U3903 , P2_U5251 );
nand NAND2_5924 ( P2_U5372 , P2_U5436 , P2_U3080 );
nand NAND2_5925 ( P2_U5373 , P2_U3395 , P2_U5251 );
nand NAND2_5926 ( P2_U5374 , P2_U5253 , P2_U3067 );
nand NAND2_5927 ( P2_U5375 , P2_U5436 , P2_U3077 );
nand NAND2_5928 ( P2_U5376 , P2_U3445 , P2_U5251 );
nand NAND2_5929 ( P2_U5377 , P2_U5253 , P2_U3080 );
nand NAND2_5930 ( P2_U5378 , P2_U5436 , P2_U3081 );
nand NAND2_5931 ( P2_U5379 , P2_U3443 , P2_U5251 );
nand NAND2_5932 ( P2_U5380 , P2_U5253 , P2_U3081 );
nand NAND2_5933 ( P2_U5381 , P2_U5436 , P2_U3068 );
nand NAND2_5934 ( P2_U5382 , P2_U3440 , P2_U5251 );
nand NAND2_5935 ( P2_U5383 , P2_U5253 , P2_U3068 );
nand NAND2_5936 ( P2_U5384 , P2_U5436 , P2_U3072 );
nand NAND2_5937 ( P2_U5385 , P2_U3437 , P2_U5251 );
nand NAND2_5938 ( P2_U5386 , P2_U5253 , P2_U3072 );
nand NAND2_5939 ( P2_U5387 , P2_U5436 , P2_U3073 );
nand NAND2_5940 ( P2_U5388 , P2_U3434 , P2_U5251 );
nand NAND2_5941 ( P2_U5389 , P2_U5253 , P2_U3073 );
nand NAND2_5942 ( P2_U5390 , P2_U5436 , P2_U3078 );
nand NAND2_5943 ( P2_U5391 , P2_U3431 , P2_U5251 );
nand NAND2_5944 ( P2_U5392 , P2_U5253 , P2_U3078 );
nand NAND2_5945 ( P2_U5393 , P2_U5436 , P2_U3079 );
nand NAND2_5946 ( P2_U5394 , P2_U3428 , P2_U5251 );
nand NAND2_5947 ( P2_U5395 , P2_U5253 , P2_U3079 );
nand NAND2_5948 ( P2_U5396 , P2_U5436 , P2_U3071 );
nand NAND2_5949 ( P2_U5397 , P2_U3425 , P2_U5251 );
nand NAND2_5950 ( P2_U5398 , P2_U5253 , P2_U3071 );
nand NAND2_5951 ( P2_U5399 , P2_U5436 , P2_U3062 );
nand NAND2_5952 ( P2_U5400 , P2_U3422 , P2_U5251 );
nand NAND2_5953 ( P2_U5401 , P2_U5253 , P2_U3062 );
nand NAND2_5954 ( P2_U5402 , P2_U5436 , P2_U3061 );
nand NAND2_5955 ( P2_U5403 , P2_U3419 , P2_U5251 );
nand NAND2_5956 ( P2_U5404 , P2_U5253 , P2_U3061 );
nand NAND2_5957 ( P2_U5405 , P2_U5436 , P2_U3082 );
nand NAND2_5958 ( P2_U5406 , P2_U3392 , P2_U5251 );
nand NAND2_5959 ( P2_U5407 , P2_U5253 , P2_U3077 );
nand NAND2_5960 ( P2_U5408 , P2_U5436 , P2_U3076 );
nand NAND2_5961 ( P2_U5409 , P2_U3387 , P2_U5251 );
nand NAND2_5962 ( P2_U5410 , P2_U5253 , P2_U3076 );
nand NAND2_5963 ( P2_U5411 , P2_U4977 , P2_U3151 );
nand NAND3_5964 ( P2_U5412 , P2_U4977 , P2_U5436 , P2_U4976 );
nand NAND2_5965 ( P2_U5413 , P2_U3043 , P2_U3303 );
nand NAND2_5966 ( P2_U5414 , P2_U3043 , P2_U3890 );
not NOT1_5967 ( P2_U5415 , P2_U3371 );
nand NAND2_5968 ( P2_U5416 , P2_U5414 , P2_U3914 );
nand NAND3_5969 ( P2_U5417 , P2_U5934 , P2_U5933 , P2_U3779 );
nand NAND2_5970 ( P2_U5418 , P2_U5430 , P2_U5424 );
nand NAND2_5971 ( P2_U5419 , P2_U3875 , P2_U3378 );
nand NAND2_5972 ( P2_U5420 , P2_U3375 , P2_U3829 );
nand NAND2_5973 ( P2_U5421 , P2_U3872 , P2_U5443 );
nand NAND2_5974 ( P2_U5422 , P2_IR_REG_24_ , P2_U3827 );
nand NAND2_5975 ( P2_U5423 , P2_IR_REG_31_ , P2_SUB_594_U19 );
not NOT1_5976 ( P2_U5424 , P2_U3372 );
nand NAND2_5977 ( P2_U5425 , P2_IR_REG_25_ , P2_U3827 );
nand NAND2_5978 ( P2_U5426 , P2_IR_REG_31_ , P2_SUB_594_U79 );
not NOT1_5979 ( P2_U5427 , P2_U3373 );
nand NAND2_5980 ( P2_U5428 , P2_IR_REG_26_ , P2_U3827 );
nand NAND2_5981 ( P2_U5429 , P2_IR_REG_31_ , P2_SUB_594_U20 );
not NOT1_5982 ( P2_U5430 , P2_U3374 );
nand NAND2_5983 ( P2_U5431 , P2_U5424 , P2_B_REG );
nand NAND2_5984 ( P2_U5432 , P2_U3372 , P2_U3298 );
nand NAND2_5985 ( P2_U5433 , P2_U5432 , P2_U5431 );
nand NAND2_5986 ( P2_U5434 , P2_IR_REG_23_ , P2_U3827 );
nand NAND2_5987 ( P2_U5435 , P2_IR_REG_31_ , P2_SUB_594_U18 );
not NOT1_5988 ( P2_U5436 , P2_U3375 );
nand NAND2_5989 ( P2_U5437 , P2_D_REG_0_ , P2_U3828 );
nand NAND2_5990 ( P2_U5438 , P2_U3911 , P2_U4016 );
nand NAND2_5991 ( P2_U5439 , P2_D_REG_1_ , P2_U3828 );
nand NAND2_5992 ( P2_U5440 , P2_U3911 , P2_U4017 );
nand NAND2_5993 ( P2_U5441 , P2_IR_REG_20_ , P2_U3827 );
nand NAND2_5994 ( P2_U5442 , P2_IR_REG_31_ , P2_SUB_594_U16 );
not NOT1_5995 ( P2_U5443 , P2_U3378 );
nand NAND2_5996 ( P2_U5444 , P2_IR_REG_19_ , P2_U3827 );
nand NAND2_5997 ( P2_U5445 , P2_IR_REG_31_ , P2_SUB_594_U15 );
not NOT1_5998 ( P2_U5446 , P2_U3379 );
nand NAND2_5999 ( P2_U5447 , P2_IR_REG_22_ , P2_U3827 );
nand NAND2_6000 ( P2_U5448 , P2_IR_REG_31_ , P2_SUB_594_U17 );
not NOT1_6001 ( P2_U5449 , P2_U3380 );
nand NAND2_6002 ( P2_U5450 , P2_IR_REG_21_ , P2_U3827 );
nand NAND2_6003 ( P2_U5451 , P2_IR_REG_31_ , P2_SUB_594_U81 );
not NOT1_6004 ( P2_U5452 , P2_U3385 );
nand NAND2_6005 ( P2_U5453 , P2_IR_REG_30_ , P2_U3827 );
nand NAND2_6006 ( P2_U5454 , P2_IR_REG_31_ , P2_SUB_594_U75 );
not NOT1_6007 ( P2_U5455 , P2_U3381 );
nand NAND2_6008 ( P2_U5456 , P2_IR_REG_29_ , P2_U3827 );
nand NAND2_6009 ( P2_U5457 , P2_IR_REG_31_ , P2_SUB_594_U22 );
not NOT1_6010 ( P2_U5458 , P2_U3382 );
nand NAND2_6011 ( P2_U5459 , P2_IR_REG_28_ , P2_U3827 );
nand NAND2_6012 ( P2_U5460 , P2_IR_REG_31_ , P2_SUB_594_U21 );
not NOT1_6013 ( P2_U5461 , P2_U3383 );
nand NAND2_6014 ( P2_U5462 , P2_IR_REG_27_ , P2_U3827 );
nand NAND2_6015 ( P2_U5463 , P2_IR_REG_31_ , P2_SUB_594_U77 );
not NOT1_6016 ( P2_U5464 , P2_U3384 );
nand NAND2_6017 ( P2_U5465 , P2_IR_REG_0_ , P2_U3827 );
nand NAND2_6018 ( P2_U5466 , P2_IR_REG_31_ , P2_IR_REG_0_ );
nand NAND2_6019 ( P2_U5467 , U56 , P2_U3829 );
nand NAND2_6020 ( P2_U5468 , P2_U3889 , P2_U3386 );
not NOT1_6021 ( P2_U5469 , P2_U3387 );
nand NAND2_6022 ( P2_U5470 , P2_U5418 , P2_U3300 );
nand NAND2_6023 ( P2_U5471 , P2_D_REG_0_ , P2_U4015 );
not NOT1_6024 ( P2_U5472 , P2_U3388 );
nand NAND2_6025 ( P2_U5473 , P2_D_REG_1_ , P2_U4015 );
nand NAND2_6026 ( P2_U5474 , P2_U4017 , P2_U3300 );
not NOT1_6027 ( P2_U5475 , P2_U3389 );
nand NAND2_6028 ( P2_U5476 , P2_U4048 , P2_U5449 );
nand NAND2_6029 ( P2_U5477 , P2_U3380 , P2_U3830 );
nand NAND2_6030 ( P2_U5478 , P2_U5477 , P2_U5476 );
nand NAND2_6031 ( P2_U5479 , P2_REG0_REG_0_ , P2_U3831 );
nand NAND2_6032 ( P2_U5480 , P2_U3910 , P2_U4073 );
nand NAND2_6033 ( P2_U5481 , P2_IR_REG_1_ , P2_U3827 );
nand NAND2_6034 ( P2_U5482 , P2_IR_REG_31_ , P2_SUB_594_U53 );
nand NAND2_6035 ( P2_U5483 , U45 , P2_U3829 );
nand NAND2_6036 ( P2_U5484 , P2_U3391 , P2_U3889 );
not NOT1_6037 ( P2_U5485 , P2_U3392 );
nand NAND2_6038 ( P2_U5486 , P2_REG0_REG_1_ , P2_U3831 );
nand NAND2_6039 ( P2_U5487 , P2_U3910 , P2_U4098 );
nand NAND2_6040 ( P2_U5488 , P2_IR_REG_2_ , P2_U3827 );
nand NAND2_6041 ( P2_U5489 , P2_IR_REG_31_ , P2_SUB_594_U23 );
nand NAND2_6042 ( P2_U5490 , U34 , P2_U3829 );
nand NAND2_6043 ( P2_U5491 , P2_U3394 , P2_U3889 );
not NOT1_6044 ( P2_U5492 , P2_U3395 );
nand NAND2_6045 ( P2_U5493 , P2_REG0_REG_2_ , P2_U3831 );
nand NAND2_6046 ( P2_U5494 , P2_U3910 , P2_U4116 );
nand NAND2_6047 ( P2_U5495 , P2_IR_REG_3_ , P2_U3827 );
nand NAND2_6048 ( P2_U5496 , P2_IR_REG_31_ , P2_SUB_594_U24 );
nand NAND2_6049 ( P2_U5497 , U31 , P2_U3829 );
nand NAND2_6050 ( P2_U5498 , P2_U3397 , P2_U3889 );
not NOT1_6051 ( P2_U5499 , P2_U3398 );
nand NAND2_6052 ( P2_U5500 , P2_REG0_REG_3_ , P2_U3831 );
nand NAND2_6053 ( P2_U5501 , P2_U3910 , P2_U4134 );
nand NAND2_6054 ( P2_U5502 , P2_IR_REG_4_ , P2_U3827 );
nand NAND2_6055 ( P2_U5503 , P2_IR_REG_31_ , P2_SUB_594_U25 );
nand NAND2_6056 ( P2_U5504 , U30 , P2_U3829 );
nand NAND2_6057 ( P2_U5505 , P2_U3400 , P2_U3889 );
not NOT1_6058 ( P2_U5506 , P2_U3401 );
nand NAND2_6059 ( P2_U5507 , P2_REG0_REG_4_ , P2_U3831 );
nand NAND2_6060 ( P2_U5508 , P2_U3910 , P2_U4152 );
nand NAND2_6061 ( P2_U5509 , P2_IR_REG_5_ , P2_U3827 );
nand NAND2_6062 ( P2_U5510 , P2_IR_REG_31_ , P2_SUB_594_U72 );
nand NAND2_6063 ( P2_U5511 , U29 , P2_U3829 );
nand NAND2_6064 ( P2_U5512 , P2_U3403 , P2_U3889 );
not NOT1_6065 ( P2_U5513 , P2_U3404 );
nand NAND2_6066 ( P2_U5514 , P2_REG0_REG_5_ , P2_U3831 );
nand NAND2_6067 ( P2_U5515 , P2_U3910 , P2_U4170 );
nand NAND2_6068 ( P2_U5516 , P2_IR_REG_6_ , P2_U3827 );
nand NAND2_6069 ( P2_U5517 , P2_IR_REG_31_ , P2_SUB_594_U26 );
nand NAND2_6070 ( P2_U5518 , U28 , P2_U3829 );
nand NAND2_6071 ( P2_U5519 , P2_U3406 , P2_U3889 );
not NOT1_6072 ( P2_U5520 , P2_U3407 );
nand NAND2_6073 ( P2_U5521 , P2_REG0_REG_6_ , P2_U3831 );
nand NAND2_6074 ( P2_U5522 , P2_U3910 , P2_U4188 );
nand NAND2_6075 ( P2_U5523 , P2_IR_REG_7_ , P2_U3827 );
nand NAND2_6076 ( P2_U5524 , P2_IR_REG_31_ , P2_SUB_594_U27 );
nand NAND2_6077 ( P2_U5525 , U27 , P2_U3829 );
nand NAND2_6078 ( P2_U5526 , P2_U3409 , P2_U3889 );
not NOT1_6079 ( P2_U5527 , P2_U3410 );
nand NAND2_6080 ( P2_U5528 , P2_REG0_REG_7_ , P2_U3831 );
nand NAND2_6081 ( P2_U5529 , P2_U3910 , P2_U4206 );
nand NAND2_6082 ( P2_U5530 , P2_IR_REG_8_ , P2_U3827 );
nand NAND2_6083 ( P2_U5531 , P2_IR_REG_31_ , P2_SUB_594_U28 );
nand NAND2_6084 ( P2_U5532 , U26 , P2_U3829 );
nand NAND2_6085 ( P2_U5533 , P2_U3412 , P2_U3889 );
not NOT1_6086 ( P2_U5534 , P2_U3413 );
nand NAND2_6087 ( P2_U5535 , P2_REG0_REG_8_ , P2_U3831 );
nand NAND2_6088 ( P2_U5536 , P2_U3910 , P2_U4224 );
nand NAND2_6089 ( P2_U5537 , P2_IR_REG_9_ , P2_U3827 );
nand NAND2_6090 ( P2_U5538 , P2_IR_REG_31_ , P2_SUB_594_U70 );
nand NAND2_6091 ( P2_U5539 , U25 , P2_U3829 );
nand NAND2_6092 ( P2_U5540 , P2_U3415 , P2_U3889 );
not NOT1_6093 ( P2_U5541 , P2_U3416 );
nand NAND2_6094 ( P2_U5542 , P2_REG0_REG_9_ , P2_U3831 );
nand NAND2_6095 ( P2_U5543 , P2_U3910 , P2_U4242 );
nand NAND2_6096 ( P2_U5544 , P2_IR_REG_10_ , P2_U3827 );
nand NAND2_6097 ( P2_U5545 , P2_IR_REG_31_ , P2_SUB_594_U8 );
nand NAND2_6098 ( P2_U5546 , U55 , P2_U3829 );
nand NAND2_6099 ( P2_U5547 , P2_U3418 , P2_U3889 );
not NOT1_6100 ( P2_U5548 , P2_U3419 );
nand NAND2_6101 ( P2_U5549 , P2_REG0_REG_10_ , P2_U3831 );
nand NAND2_6102 ( P2_U5550 , P2_U3910 , P2_U4260 );
nand NAND2_6103 ( P2_U5551 , P2_IR_REG_11_ , P2_U3827 );
nand NAND2_6104 ( P2_U5552 , P2_IR_REG_31_ , P2_SUB_594_U9 );
nand NAND2_6105 ( P2_U5553 , U54 , P2_U3829 );
nand NAND2_6106 ( P2_U5554 , P2_U3421 , P2_U3889 );
not NOT1_6107 ( P2_U5555 , P2_U3422 );
nand NAND2_6108 ( P2_U5556 , P2_REG0_REG_11_ , P2_U3831 );
nand NAND2_6109 ( P2_U5557 , P2_U3910 , P2_U4278 );
nand NAND2_6110 ( P2_U5558 , P2_IR_REG_12_ , P2_U3827 );
nand NAND2_6111 ( P2_U5559 , P2_IR_REG_31_ , P2_SUB_594_U10 );
nand NAND2_6112 ( P2_U5560 , U53 , P2_U3829 );
nand NAND2_6113 ( P2_U5561 , P2_U3424 , P2_U3889 );
not NOT1_6114 ( P2_U5562 , P2_U3425 );
nand NAND2_6115 ( P2_U5563 , P2_REG0_REG_12_ , P2_U3831 );
nand NAND2_6116 ( P2_U5564 , P2_U3910 , P2_U4296 );
nand NAND2_6117 ( P2_U5565 , P2_IR_REG_13_ , P2_U3827 );
nand NAND2_6118 ( P2_U5566 , P2_IR_REG_31_ , P2_SUB_594_U87 );
nand NAND2_6119 ( P2_U5567 , U52 , P2_U3829 );
nand NAND2_6120 ( P2_U5568 , P2_U3427 , P2_U3889 );
not NOT1_6121 ( P2_U5569 , P2_U3428 );
nand NAND2_6122 ( P2_U5570 , P2_REG0_REG_13_ , P2_U3831 );
nand NAND2_6123 ( P2_U5571 , P2_U3910 , P2_U4314 );
nand NAND2_6124 ( P2_U5572 , P2_IR_REG_14_ , P2_U3827 );
nand NAND2_6125 ( P2_U5573 , P2_IR_REG_31_ , P2_SUB_594_U11 );
nand NAND2_6126 ( P2_U5574 , U51 , P2_U3829 );
nand NAND2_6127 ( P2_U5575 , P2_U3430 , P2_U3889 );
not NOT1_6128 ( P2_U5576 , P2_U3431 );
nand NAND2_6129 ( P2_U5577 , P2_REG0_REG_14_ , P2_U3831 );
nand NAND2_6130 ( P2_U5578 , P2_U3910 , P2_U4332 );
nand NAND2_6131 ( P2_U5579 , P2_IR_REG_15_ , P2_U3827 );
nand NAND2_6132 ( P2_U5580 , P2_IR_REG_31_ , P2_SUB_594_U12 );
nand NAND2_6133 ( P2_U5581 , U50 , P2_U3829 );
nand NAND2_6134 ( P2_U5582 , P2_U3433 , P2_U3889 );
not NOT1_6135 ( P2_U5583 , P2_U3434 );
nand NAND2_6136 ( P2_U5584 , P2_REG0_REG_15_ , P2_U3831 );
nand NAND2_6137 ( P2_U5585 , P2_U3910 , P2_U4350 );
nand NAND2_6138 ( P2_U5586 , P2_IR_REG_16_ , P2_U3827 );
nand NAND2_6139 ( P2_U5587 , P2_IR_REG_31_ , P2_SUB_594_U13 );
nand NAND2_6140 ( P2_U5588 , U49 , P2_U3829 );
nand NAND2_6141 ( P2_U5589 , P2_U3436 , P2_U3889 );
not NOT1_6142 ( P2_U5590 , P2_U3437 );
nand NAND2_6143 ( P2_U5591 , P2_REG0_REG_16_ , P2_U3831 );
nand NAND2_6144 ( P2_U5592 , P2_U3910 , P2_U4368 );
nand NAND2_6145 ( P2_U5593 , P2_IR_REG_17_ , P2_U3827 );
nand NAND2_6146 ( P2_U5594 , P2_IR_REG_31_ , P2_SUB_594_U85 );
nand NAND2_6147 ( P2_U5595 , U48 , P2_U3829 );
nand NAND2_6148 ( P2_U5596 , P2_U3439 , P2_U3889 );
not NOT1_6149 ( P2_U5597 , P2_U3440 );
nand NAND2_6150 ( P2_U5598 , P2_REG0_REG_17_ , P2_U3831 );
nand NAND2_6151 ( P2_U5599 , P2_U3910 , P2_U4386 );
nand NAND2_6152 ( P2_U5600 , P2_IR_REG_18_ , P2_U3827 );
nand NAND2_6153 ( P2_U5601 , P2_IR_REG_31_ , P2_SUB_594_U14 );
nand NAND2_6154 ( P2_U5602 , U47 , P2_U3829 );
nand NAND2_6155 ( P2_U5603 , P2_U3442 , P2_U3889 );
not NOT1_6156 ( P2_U5604 , P2_U3443 );
nand NAND2_6157 ( P2_U5605 , P2_REG0_REG_18_ , P2_U3831 );
nand NAND2_6158 ( P2_U5606 , P2_U3910 , P2_U4404 );
nand NAND2_6159 ( P2_U5607 , U46 , P2_U3829 );
nand NAND2_6160 ( P2_U5608 , P2_U3889 , P2_U3379 );
not NOT1_6161 ( P2_U5609 , P2_U3445 );
nand NAND2_6162 ( P2_U5610 , P2_REG0_REG_19_ , P2_U3831 );
nand NAND2_6163 ( P2_U5611 , P2_U3910 , P2_U4422 );
nand NAND2_6164 ( P2_U5612 , P2_REG0_REG_20_ , P2_U3831 );
nand NAND2_6165 ( P2_U5613 , P2_U3910 , P2_U4440 );
nand NAND2_6166 ( P2_U5614 , P2_REG0_REG_21_ , P2_U3831 );
nand NAND2_6167 ( P2_U5615 , P2_U3910 , P2_U4458 );
nand NAND2_6168 ( P2_U5616 , P2_REG0_REG_22_ , P2_U3831 );
nand NAND2_6169 ( P2_U5617 , P2_U3910 , P2_U4476 );
nand NAND2_6170 ( P2_U5618 , P2_REG0_REG_23_ , P2_U3831 );
nand NAND2_6171 ( P2_U5619 , P2_U3910 , P2_U4494 );
nand NAND2_6172 ( P2_U5620 , P2_REG0_REG_24_ , P2_U3831 );
nand NAND2_6173 ( P2_U5621 , P2_U3910 , P2_U4512 );
nand NAND2_6174 ( P2_U5622 , P2_REG0_REG_25_ , P2_U3831 );
nand NAND2_6175 ( P2_U5623 , P2_U3910 , P2_U4530 );
nand NAND2_6176 ( P2_U5624 , P2_REG0_REG_26_ , P2_U3831 );
nand NAND2_6177 ( P2_U5625 , P2_U3910 , P2_U4548 );
nand NAND2_6178 ( P2_U5626 , P2_REG0_REG_27_ , P2_U3831 );
nand NAND2_6179 ( P2_U5627 , P2_U3910 , P2_U4566 );
nand NAND2_6180 ( P2_U5628 , P2_REG0_REG_28_ , P2_U3831 );
nand NAND2_6181 ( P2_U5629 , P2_U3910 , P2_U4584 );
nand NAND2_6182 ( P2_U5630 , P2_REG0_REG_29_ , P2_U3831 );
nand NAND2_6183 ( P2_U5631 , P2_U3910 , P2_U4604 );
nand NAND2_6184 ( P2_U5632 , P2_REG0_REG_30_ , P2_U3831 );
nand NAND2_6185 ( P2_U5633 , P2_U3910 , P2_U4611 );
nand NAND2_6186 ( P2_U5634 , P2_REG0_REG_31_ , P2_U3831 );
nand NAND2_6187 ( P2_U5635 , P2_U3910 , P2_U4613 );
nand NAND2_6188 ( P2_U5636 , P2_U5449 , P2_U3830 );
nand NAND2_6189 ( P2_U5637 , P2_U4048 , P2_U5446 );
nand NAND2_6190 ( P2_U5638 , P2_REG1_REG_0_ , P2_U3832 );
nand NAND2_6191 ( P2_U5639 , P2_U3909 , P2_U4073 );
nand NAND2_6192 ( P2_U5640 , P2_REG1_REG_1_ , P2_U3832 );
nand NAND2_6193 ( P2_U5641 , P2_U3909 , P2_U4098 );
nand NAND2_6194 ( P2_U5642 , P2_REG1_REG_2_ , P2_U3832 );
nand NAND2_6195 ( P2_U5643 , P2_U3909 , P2_U4116 );
nand NAND2_6196 ( P2_U5644 , P2_REG1_REG_3_ , P2_U3832 );
nand NAND2_6197 ( P2_U5645 , P2_U3909 , P2_U4134 );
nand NAND2_6198 ( P2_U5646 , P2_REG1_REG_4_ , P2_U3832 );
nand NAND2_6199 ( P2_U5647 , P2_U3909 , P2_U4152 );
nand NAND2_6200 ( P2_U5648 , P2_REG1_REG_5_ , P2_U3832 );
nand NAND2_6201 ( P2_U5649 , P2_U3909 , P2_U4170 );
nand NAND2_6202 ( P2_U5650 , P2_REG1_REG_6_ , P2_U3832 );
nand NAND2_6203 ( P2_U5651 , P2_U3909 , P2_U4188 );
nand NAND2_6204 ( P2_U5652 , P2_REG1_REG_7_ , P2_U3832 );
nand NAND2_6205 ( P2_U5653 , P2_U3909 , P2_U4206 );
nand NAND2_6206 ( P2_U5654 , P2_REG1_REG_8_ , P2_U3832 );
nand NAND2_6207 ( P2_U5655 , P2_U3909 , P2_U4224 );
nand NAND2_6208 ( P2_U5656 , P2_REG1_REG_9_ , P2_U3832 );
nand NAND2_6209 ( P2_U5657 , P2_U3909 , P2_U4242 );
nand NAND2_6210 ( P2_U5658 , P2_REG1_REG_10_ , P2_U3832 );
nand NAND2_6211 ( P2_U5659 , P2_U3909 , P2_U4260 );
nand NAND2_6212 ( P2_U5660 , P2_REG1_REG_11_ , P2_U3832 );
nand NAND2_6213 ( P2_U5661 , P2_U3909 , P2_U4278 );
nand NAND2_6214 ( P2_U5662 , P2_REG1_REG_12_ , P2_U3832 );
nand NAND2_6215 ( P2_U5663 , P2_U3909 , P2_U4296 );
nand NAND2_6216 ( P2_U5664 , P2_REG1_REG_13_ , P2_U3832 );
nand NAND2_6217 ( P2_U5665 , P2_U3909 , P2_U4314 );
nand NAND2_6218 ( P2_U5666 , P2_REG1_REG_14_ , P2_U3832 );
nand NAND2_6219 ( P2_U5667 , P2_U3909 , P2_U4332 );
nand NAND2_6220 ( P2_U5668 , P2_REG1_REG_15_ , P2_U3832 );
nand NAND2_6221 ( P2_U5669 , P2_U3909 , P2_U4350 );
nand NAND2_6222 ( P2_U5670 , P2_REG1_REG_16_ , P2_U3832 );
nand NAND2_6223 ( P2_U5671 , P2_U3909 , P2_U4368 );
nand NAND2_6224 ( P2_U5672 , P2_REG1_REG_17_ , P2_U3832 );
nand NAND2_6225 ( P2_U5673 , P2_U3909 , P2_U4386 );
nand NAND2_6226 ( P2_U5674 , P2_REG1_REG_18_ , P2_U3832 );
nand NAND2_6227 ( P2_U5675 , P2_U3909 , P2_U4404 );
nand NAND2_6228 ( P2_U5676 , P2_REG1_REG_19_ , P2_U3832 );
nand NAND2_6229 ( P2_U5677 , P2_U3909 , P2_U4422 );
nand NAND2_6230 ( P2_U5678 , P2_REG1_REG_20_ , P2_U3832 );
nand NAND2_6231 ( P2_U5679 , P2_U3909 , P2_U4440 );
nand NAND2_6232 ( P2_U5680 , P2_REG1_REG_21_ , P2_U3832 );
nand NAND2_6233 ( P2_U5681 , P2_U3909 , P2_U4458 );
nand NAND2_6234 ( P2_U5682 , P2_REG1_REG_22_ , P2_U3832 );
nand NAND2_6235 ( P2_U5683 , P2_U3909 , P2_U4476 );
nand NAND2_6236 ( P2_U5684 , P2_REG1_REG_23_ , P2_U3832 );
nand NAND2_6237 ( P2_U5685 , P2_U3909 , P2_U4494 );
nand NAND2_6238 ( P2_U5686 , P2_REG1_REG_24_ , P2_U3832 );
nand NAND2_6239 ( P2_U5687 , P2_U3909 , P2_U4512 );
nand NAND2_6240 ( P2_U5688 , P2_REG1_REG_25_ , P2_U3832 );
nand NAND2_6241 ( P2_U5689 , P2_U3909 , P2_U4530 );
nand NAND2_6242 ( P2_U5690 , P2_REG1_REG_26_ , P2_U3832 );
nand NAND2_6243 ( P2_U5691 , P2_U3909 , P2_U4548 );
nand NAND2_6244 ( P2_U5692 , P2_REG1_REG_27_ , P2_U3832 );
nand NAND2_6245 ( P2_U5693 , P2_U3909 , P2_U4566 );
nand NAND2_6246 ( P2_U5694 , P2_REG1_REG_28_ , P2_U3832 );
nand NAND2_6247 ( P2_U5695 , P2_U3909 , P2_U4584 );
nand NAND2_6248 ( P2_U5696 , P2_REG1_REG_29_ , P2_U3832 );
nand NAND2_6249 ( P2_U5697 , P2_U3909 , P2_U4604 );
nand NAND2_6250 ( P2_U5698 , P2_REG1_REG_30_ , P2_U3832 );
nand NAND2_6251 ( P2_U5699 , P2_U3909 , P2_U4611 );
nand NAND2_6252 ( P2_U5700 , P2_REG1_REG_31_ , P2_U3832 );
nand NAND2_6253 ( P2_U5701 , P2_U3909 , P2_U4613 );
nand NAND2_6254 ( P2_U5702 , P2_REG2_REG_0_ , P2_U3358 );
nand NAND2_6255 ( P2_U5703 , P2_U3908 , P2_U3314 );
nand NAND2_6256 ( P2_U5704 , P2_REG2_REG_1_ , P2_U3358 );
nand NAND2_6257 ( P2_U5705 , P2_U3908 , P2_U3315 );
nand NAND2_6258 ( P2_U5706 , P2_REG2_REG_2_ , P2_U3358 );
nand NAND2_6259 ( P2_U5707 , P2_U3908 , P2_U3316 );
nand NAND2_6260 ( P2_U5708 , P2_REG2_REG_3_ , P2_U3358 );
nand NAND2_6261 ( P2_U5709 , P2_U3908 , P2_U3317 );
nand NAND2_6262 ( P2_U5710 , P2_REG2_REG_4_ , P2_U3358 );
nand NAND2_6263 ( P2_U5711 , P2_U3908 , P2_U3318 );
nand NAND2_6264 ( P2_U5712 , P2_REG2_REG_5_ , P2_U3358 );
nand NAND2_6265 ( P2_U5713 , P2_U3908 , P2_U3319 );
nand NAND2_6266 ( P2_U5714 , P2_REG2_REG_6_ , P2_U3358 );
nand NAND2_6267 ( P2_U5715 , P2_U3908 , P2_U3320 );
nand NAND2_6268 ( P2_U5716 , P2_REG2_REG_7_ , P2_U3358 );
nand NAND2_6269 ( P2_U5717 , P2_U3908 , P2_U3321 );
nand NAND2_6270 ( P2_U5718 , P2_REG2_REG_8_ , P2_U3358 );
nand NAND2_6271 ( P2_U5719 , P2_U3908 , P2_U3322 );
nand NAND2_6272 ( P2_U5720 , P2_REG2_REG_9_ , P2_U3358 );
nand NAND2_6273 ( P2_U5721 , P2_U3908 , P2_U3323 );
nand NAND2_6274 ( P2_U5722 , P2_REG2_REG_10_ , P2_U3358 );
nand NAND2_6275 ( P2_U5723 , P2_U3908 , P2_U3324 );
nand NAND2_6276 ( P2_U5724 , P2_REG2_REG_11_ , P2_U3358 );
nand NAND2_6277 ( P2_U5725 , P2_U3908 , P2_U3325 );
nand NAND2_6278 ( P2_U5726 , P2_REG2_REG_12_ , P2_U3358 );
nand NAND2_6279 ( P2_U5727 , P2_U3908 , P2_U3326 );
nand NAND2_6280 ( P2_U5728 , P2_REG2_REG_13_ , P2_U3358 );
nand NAND2_6281 ( P2_U5729 , P2_U3908 , P2_U3327 );
nand NAND2_6282 ( P2_U5730 , P2_REG2_REG_14_ , P2_U3358 );
nand NAND2_6283 ( P2_U5731 , P2_U3908 , P2_U3328 );
nand NAND2_6284 ( P2_U5732 , P2_REG2_REG_15_ , P2_U3358 );
nand NAND2_6285 ( P2_U5733 , P2_U3908 , P2_U3329 );
nand NAND2_6286 ( P2_U5734 , P2_REG2_REG_16_ , P2_U3358 );
nand NAND2_6287 ( P2_U5735 , P2_U3908 , P2_U3330 );
nand NAND2_6288 ( P2_U5736 , P2_REG2_REG_17_ , P2_U3358 );
nand NAND2_6289 ( P2_U5737 , P2_U3908 , P2_U3331 );
nand NAND2_6290 ( P2_U5738 , P2_REG2_REG_18_ , P2_U3358 );
nand NAND2_6291 ( P2_U5739 , P2_U3908 , P2_U3332 );
nand NAND2_6292 ( P2_U5740 , P2_REG2_REG_19_ , P2_U3358 );
nand NAND2_6293 ( P2_U5741 , P2_U3908 , P2_U3333 );
nand NAND2_6294 ( P2_U5742 , P2_REG2_REG_20_ , P2_U3358 );
nand NAND2_6295 ( P2_U5743 , P2_U3908 , P2_U3335 );
nand NAND2_6296 ( P2_U5744 , P2_REG2_REG_21_ , P2_U3358 );
nand NAND2_6297 ( P2_U5745 , P2_U3908 , P2_U3337 );
nand NAND2_6298 ( P2_U5746 , P2_REG2_REG_22_ , P2_U3358 );
nand NAND2_6299 ( P2_U5747 , P2_U3908 , P2_U3339 );
nand NAND2_6300 ( P2_U5748 , P2_REG2_REG_23_ , P2_U3358 );
nand NAND2_6301 ( P2_U5749 , P2_U3908 , P2_U3341 );
nand NAND2_6302 ( P2_U5750 , P2_REG2_REG_24_ , P2_U3358 );
nand NAND2_6303 ( P2_U5751 , P2_U3908 , P2_U3343 );
nand NAND2_6304 ( P2_U5752 , P2_REG2_REG_25_ , P2_U3358 );
nand NAND2_6305 ( P2_U5753 , P2_U3908 , P2_U3345 );
nand NAND2_6306 ( P2_U5754 , P2_REG2_REG_26_ , P2_U3358 );
nand NAND2_6307 ( P2_U5755 , P2_U3908 , P2_U3347 );
nand NAND2_6308 ( P2_U5756 , P2_REG2_REG_27_ , P2_U3358 );
nand NAND2_6309 ( P2_U5757 , P2_U3908 , P2_U3349 );
nand NAND2_6310 ( P2_U5758 , P2_REG2_REG_28_ , P2_U3358 );
nand NAND2_6311 ( P2_U5759 , P2_U3908 , P2_U3351 );
nand NAND2_6312 ( P2_U5760 , P2_REG2_REG_29_ , P2_U3358 );
nand NAND2_6313 ( P2_U5761 , P2_U3908 , P2_U3354 );
nand NAND2_6314 ( P2_U5762 , P2_U5461 , P2_U3024 );
nand NAND2_6315 ( P2_U5763 , P2_U3383 , P2_U3893 );
nand NAND2_6316 ( P2_U5764 , P2_U5763 , P2_U5762 );
nand NAND2_6317 ( P2_U5765 , P2_DATAO_REG_0_ , P2_U3363 );
nand NAND2_6318 ( P2_U5766 , P2_U3893 , P2_U3076 );
nand NAND2_6319 ( P2_U5767 , P2_DATAO_REG_1_ , P2_U3363 );
nand NAND2_6320 ( P2_U5768 , P2_U3893 , P2_U3077 );
nand NAND2_6321 ( P2_U5769 , P2_DATAO_REG_2_ , P2_U3363 );
nand NAND2_6322 ( P2_U5770 , P2_U3893 , P2_U3067 );
nand NAND2_6323 ( P2_U5771 , P2_DATAO_REG_3_ , P2_U3363 );
nand NAND2_6324 ( P2_U5772 , P2_U3893 , P2_U3063 );
nand NAND2_6325 ( P2_U5773 , P2_DATAO_REG_4_ , P2_U3363 );
nand NAND2_6326 ( P2_U5774 , P2_U3893 , P2_U3059 );
nand NAND2_6327 ( P2_U5775 , P2_DATAO_REG_5_ , P2_U3363 );
nand NAND2_6328 ( P2_U5776 , P2_U3893 , P2_U3066 );
nand NAND2_6329 ( P2_U5777 , P2_DATAO_REG_6_ , P2_U3363 );
nand NAND2_6330 ( P2_U5778 , P2_U3893 , P2_U3070 );
nand NAND2_6331 ( P2_U5779 , P2_DATAO_REG_7_ , P2_U3363 );
nand NAND2_6332 ( P2_U5780 , P2_U3893 , P2_U3069 );
nand NAND2_6333 ( P2_U5781 , P2_DATAO_REG_8_ , P2_U3363 );
nand NAND2_6334 ( P2_U5782 , P2_U3893 , P2_U3083 );
nand NAND2_6335 ( P2_U5783 , P2_DATAO_REG_9_ , P2_U3363 );
nand NAND2_6336 ( P2_U5784 , P2_U3893 , P2_U3082 );
nand NAND2_6337 ( P2_U5785 , P2_DATAO_REG_10_ , P2_U3363 );
nand NAND2_6338 ( P2_U5786 , P2_U3893 , P2_U3061 );
nand NAND2_6339 ( P2_U5787 , P2_DATAO_REG_11_ , P2_U3363 );
nand NAND2_6340 ( P2_U5788 , P2_U3893 , P2_U3062 );
nand NAND2_6341 ( P2_U5789 , P2_DATAO_REG_12_ , P2_U3363 );
nand NAND2_6342 ( P2_U5790 , P2_U3893 , P2_U3071 );
nand NAND2_6343 ( P2_U5791 , P2_DATAO_REG_13_ , P2_U3363 );
nand NAND2_6344 ( P2_U5792 , P2_U3893 , P2_U3079 );
nand NAND2_6345 ( P2_U5793 , P2_DATAO_REG_14_ , P2_U3363 );
nand NAND2_6346 ( P2_U5794 , P2_U3893 , P2_U3078 );
nand NAND2_6347 ( P2_U5795 , P2_DATAO_REG_15_ , P2_U3363 );
nand NAND2_6348 ( P2_U5796 , P2_U3893 , P2_U3073 );
nand NAND2_6349 ( P2_U5797 , P2_DATAO_REG_16_ , P2_U3363 );
nand NAND2_6350 ( P2_U5798 , P2_U3893 , P2_U3072 );
nand NAND2_6351 ( P2_U5799 , P2_DATAO_REG_17_ , P2_U3363 );
nand NAND2_6352 ( P2_U5800 , P2_U3893 , P2_U3068 );
nand NAND2_6353 ( P2_U5801 , P2_DATAO_REG_18_ , P2_U3363 );
nand NAND2_6354 ( P2_U5802 , P2_U3893 , P2_U3081 );
nand NAND2_6355 ( P2_U5803 , P2_DATAO_REG_19_ , P2_U3363 );
nand NAND2_6356 ( P2_U5804 , P2_U3893 , P2_U3080 );
nand NAND2_6357 ( P2_U5805 , P2_DATAO_REG_20_ , P2_U3363 );
nand NAND2_6358 ( P2_U5806 , P2_U3893 , P2_U3075 );
nand NAND2_6359 ( P2_U5807 , P2_DATAO_REG_21_ , P2_U3363 );
nand NAND2_6360 ( P2_U5808 , P2_U3893 , P2_U3074 );
nand NAND2_6361 ( P2_U5809 , P2_DATAO_REG_22_ , P2_U3363 );
nand NAND2_6362 ( P2_U5810 , P2_U3893 , P2_U3060 );
nand NAND2_6363 ( P2_U5811 , P2_DATAO_REG_23_ , P2_U3363 );
nand NAND2_6364 ( P2_U5812 , P2_U3893 , P2_U3065 );
nand NAND2_6365 ( P2_U5813 , P2_DATAO_REG_24_ , P2_U3363 );
nand NAND2_6366 ( P2_U5814 , P2_U3893 , P2_U3064 );
nand NAND2_6367 ( P2_U5815 , P2_DATAO_REG_25_ , P2_U3363 );
nand NAND2_6368 ( P2_U5816 , P2_U3893 , P2_U3057 );
nand NAND2_6369 ( P2_U5817 , P2_DATAO_REG_26_ , P2_U3363 );
nand NAND2_6370 ( P2_U5818 , P2_U3893 , P2_U3056 );
nand NAND2_6371 ( P2_U5819 , P2_DATAO_REG_27_ , P2_U3363 );
nand NAND2_6372 ( P2_U5820 , P2_U3893 , P2_U3052 );
nand NAND2_6373 ( P2_U5821 , P2_DATAO_REG_28_ , P2_U3363 );
nand NAND2_6374 ( P2_U5822 , P2_U3893 , P2_U3053 );
nand NAND2_6375 ( P2_U5823 , P2_DATAO_REG_29_ , P2_U3363 );
nand NAND2_6376 ( P2_U5824 , P2_U3893 , P2_U3054 );
nand NAND2_6377 ( P2_U5825 , P2_DATAO_REG_30_ , P2_U3363 );
nand NAND2_6378 ( P2_U5826 , P2_U3893 , P2_U3058 );
nand NAND2_6379 ( P2_U5827 , P2_DATAO_REG_31_ , P2_U3363 );
nand NAND2_6380 ( P2_U5828 , P2_U3893 , P2_U3055 );
nand NAND2_6381 ( P2_U5829 , P2_U3379 , P2_U3313 );
nand NAND2_6382 ( P2_U5830 , P2_U5446 , P2_U3907 );
not NOT1_6383 ( P2_U5831 , P2_U3765 );
nand NAND2_6384 ( P2_U5832 , P2_R1269_U22 , P2_U5831 );
nand NAND2_6385 ( P2_U5833 , P2_U3765 , P2_U3863 );
nand NAND2_6386 ( P2_U5834 , P2_U3896 , P2_U3052 );
nand NAND2_6387 ( P2_U5835 , P2_U3348 , P2_U4535 );
nand NAND2_6388 ( P2_U5836 , P2_U5835 , P2_U5834 );
nand NAND2_6389 ( P2_U5837 , P2_U3895 , P2_U3053 );
nand NAND2_6390 ( P2_U5838 , P2_U3350 , P2_U4553 );
nand NAND2_6391 ( P2_U5839 , P2_U5838 , P2_U5837 );
nand NAND2_6392 ( P2_U5840 , P2_U3868 , P2_U3055 );
nand NAND2_6393 ( P2_U5841 , P2_U3356 , P2_U4609 );
nand NAND2_6394 ( P2_U5842 , P2_U5841 , P2_U5840 );
nand NAND2_6395 ( P2_U5843 , P2_U3904 , P2_U3054 );
nand NAND2_6396 ( P2_U5844 , P2_U3353 , P2_U4571 );
nand NAND2_6397 ( P2_U5845 , P2_U5844 , P2_U5843 );
nand NAND2_6398 ( P2_U5846 , P2_U3902 , P2_U3074 );
nand NAND2_6399 ( P2_U5847 , P2_U3336 , P2_U4427 );
nand NAND2_6400 ( P2_U5848 , P2_U5847 , P2_U5846 );
nand NAND2_6401 ( P2_U5849 , P2_U3903 , P2_U3075 );
nand NAND2_6402 ( P2_U5850 , P2_U3334 , P2_U4409 );
nand NAND2_6403 ( P2_U5851 , P2_U5850 , P2_U5849 );
nand NAND2_6404 ( P2_U5852 , P2_U5499 , P2_U4103 );
nand NAND2_6405 ( P2_U5853 , P2_U3398 , P2_U3063 );
nand NAND2_6406 ( P2_U5854 , P2_U5853 , P2_U5852 );
nand NAND2_6407 ( P2_U5855 , P2_U5555 , P2_U4247 );
nand NAND2_6408 ( P2_U5856 , P2_U3422 , P2_U3062 );
nand NAND2_6409 ( P2_U5857 , P2_U5856 , P2_U5855 );
nand NAND2_6410 ( P2_U5858 , P2_U5548 , P2_U4229 );
nand NAND2_6411 ( P2_U5859 , P2_U3419 , P2_U3061 );
nand NAND2_6412 ( P2_U5860 , P2_U5859 , P2_U5858 );
nand NAND2_6413 ( P2_U5861 , P2_U5506 , P2_U4121 );
nand NAND2_6414 ( P2_U5862 , P2_U3401 , P2_U3059 );
nand NAND2_6415 ( P2_U5863 , P2_U5862 , P2_U5861 );
nand NAND2_6416 ( P2_U5864 , P2_U3901 , P2_U3060 );
nand NAND2_6417 ( P2_U5865 , P2_U3338 , P2_U4445 );
nand NAND2_6418 ( P2_U5866 , P2_U5865 , P2_U5864 );
nand NAND2_6419 ( P2_U5867 , P2_U5597 , P2_U4355 );
nand NAND2_6420 ( P2_U5868 , P2_U3440 , P2_U3068 );
nand NAND2_6421 ( P2_U5869 , P2_U5868 , P2_U5867 );
nand NAND2_6422 ( P2_U5870 , P2_U5583 , P2_U4319 );
nand NAND2_6423 ( P2_U5871 , P2_U3434 , P2_U3073 );
nand NAND2_6424 ( P2_U5872 , P2_U5871 , P2_U5870 );
nand NAND2_6425 ( P2_U5873 , P2_U5562 , P2_U4265 );
nand NAND2_6426 ( P2_U5874 , P2_U3425 , P2_U3071 );
nand NAND2_6427 ( P2_U5875 , P2_U5874 , P2_U5873 );
nand NAND2_6428 ( P2_U5876 , P2_U5520 , P2_U4157 );
nand NAND2_6429 ( P2_U5877 , P2_U3407 , P2_U3070 );
nand NAND2_6430 ( P2_U5878 , P2_U5877 , P2_U5876 );
nand NAND2_6431 ( P2_U5879 , P2_U5527 , P2_U4175 );
nand NAND2_6432 ( P2_U5880 , P2_U3410 , P2_U3069 );
nand NAND2_6433 ( P2_U5881 , P2_U5880 , P2_U5879 );
nand NAND2_6434 ( P2_U5882 , P2_U5492 , P2_U4078 );
nand NAND2_6435 ( P2_U5883 , P2_U3395 , P2_U3067 );
nand NAND2_6436 ( P2_U5884 , P2_U5883 , P2_U5882 );
nand NAND2_6437 ( P2_U5885 , P2_U5513 , P2_U4139 );
nand NAND2_6438 ( P2_U5886 , P2_U3404 , P2_U3066 );
nand NAND2_6439 ( P2_U5887 , P2_U5886 , P2_U5885 );
nand NAND2_6440 ( P2_U5888 , P2_U5590 , P2_U4337 );
nand NAND2_6441 ( P2_U5889 , P2_U3437 , P2_U3072 );
nand NAND2_6442 ( P2_U5890 , P2_U5889 , P2_U5888 );
nand NAND2_6443 ( P2_U5891 , P2_U5604 , P2_U4373 );
nand NAND2_6444 ( P2_U5892 , P2_U3443 , P2_U3081 );
nand NAND2_6445 ( P2_U5893 , P2_U5892 , P2_U5891 );
nand NAND2_6446 ( P2_U5894 , P2_U5569 , P2_U4283 );
nand NAND2_6447 ( P2_U5895 , P2_U3428 , P2_U3079 );
nand NAND2_6448 ( P2_U5896 , P2_U5895 , P2_U5894 );
nand NAND2_6449 ( P2_U5897 , P2_U5576 , P2_U4301 );
nand NAND2_6450 ( P2_U5898 , P2_U3431 , P2_U3078 );
nand NAND2_6451 ( P2_U5899 , P2_U5898 , P2_U5897 );
nand NAND2_6452 ( P2_U5900 , P2_U5485 , P2_U4059 );
nand NAND2_6453 ( P2_U5901 , P2_U3392 , P2_U3077 );
nand NAND2_6454 ( P2_U5902 , P2_U5901 , P2_U5900 );
nand NAND2_6455 ( P2_U5903 , P2_U5469 , P2_U4083 );
nand NAND2_6456 ( P2_U5904 , P2_U3387 , P2_U3076 );
nand NAND2_6457 ( P2_U5905 , P2_U5904 , P2_U5903 );
nand NAND2_6458 ( P2_U5906 , P2_U5534 , P2_U4193 );
nand NAND2_6459 ( P2_U5907 , P2_U3413 , P2_U3083 );
nand NAND2_6460 ( P2_U5908 , P2_U5907 , P2_U5906 );
nand NAND2_6461 ( P2_U5909 , P2_U5541 , P2_U4211 );
nand NAND2_6462 ( P2_U5910 , P2_U3416 , P2_U3082 );
nand NAND2_6463 ( P2_U5911 , P2_U5910 , P2_U5909 );
nand NAND2_6464 ( P2_U5912 , P2_U5609 , P2_U4391 );
nand NAND2_6465 ( P2_U5913 , P2_U3445 , P2_U3080 );
nand NAND2_6466 ( P2_U5914 , P2_U5913 , P2_U5912 );
nand NAND2_6467 ( P2_U5915 , P2_U3897 , P2_U3056 );
nand NAND2_6468 ( P2_U5916 , P2_U3346 , P2_U4517 );
nand NAND2_6469 ( P2_U5917 , P2_U5916 , P2_U5915 );
nand NAND2_6470 ( P2_U5918 , P2_U3898 , P2_U3057 );
nand NAND2_6471 ( P2_U5919 , P2_U3344 , P2_U4499 );
nand NAND2_6472 ( P2_U5920 , P2_U5919 , P2_U5918 );
nand NAND2_6473 ( P2_U5921 , P2_U3900 , P2_U3065 );
nand NAND2_6474 ( P2_U5922 , P2_U3340 , P2_U4463 );
nand NAND2_6475 ( P2_U5923 , P2_U5922 , P2_U5921 );
nand NAND2_6476 ( P2_U5924 , P2_U3899 , P2_U3064 );
nand NAND2_6477 ( P2_U5925 , P2_U3342 , P2_U4481 );
nand NAND2_6478 ( P2_U5926 , P2_U5925 , P2_U5924 );
nand NAND2_6479 ( P2_U5927 , P2_U3869 , P2_U3058 );
nand NAND2_6480 ( P2_U5928 , P2_U3355 , P2_U4589 );
nand NAND2_6481 ( P2_U5929 , P2_U5928 , P2_U5927 );
nand NAND2_6482 ( P2_U5930 , P2_U4974 , P2_U5446 );
nand NAND2_6483 ( P2_U5931 , P2_U3379 , P2_U3864 );
nand NAND2_6484 ( P2_U5932 , P2_U5931 , P2_U5930 );
nand NAND3_6485 ( P2_U5933 , P2_U5833 , P2_U5832 , P2_U5443 );
nand NAND3_6486 ( P2_U5934 , P2_U5452 , P2_U5932 , P2_U3378 );
nand NAND2_6487 ( P2_U5935 , P2_U3877 , P2_U3865 );
nand NAND2_6488 ( P2_U5936 , P2_R693_U14 , P2_U3887 );
nand NAND2_6489 ( P2_U5937 , P2_U5436 , P2_U3368 );
nand NAND2_6490 ( P2_U5938 , P2_U3380 , P2_U3375 );
nand NAND2_6491 ( P2_U5939 , P2_U5446 , P2_U5443 );
nand NAND3_6492 ( P2_U5940 , P2_U3388 , P2_U5452 , P2_U3378 );
nand NAND2_6493 ( P2_U5941 , P2_U3082 , P2_R1297_U6 );
nand NAND2_6494 ( P2_U5942 , P2_U3082 , P2_U3867 );
nand NAND2_6495 ( P2_U5943 , P2_U3083 , P2_R1297_U6 );
nand NAND2_6496 ( P2_U5944 , P2_U3083 , P2_U3867 );
nand NAND2_6497 ( P2_U5945 , P2_U3069 , P2_R1297_U6 );
nand NAND2_6498 ( P2_U5946 , P2_U3069 , P2_U3867 );
nand NAND2_6499 ( P2_U5947 , P2_U3070 , P2_R1297_U6 );
nand NAND2_6500 ( P2_U5948 , P2_U3070 , P2_U3867 );
nand NAND2_6501 ( P2_U5949 , P2_U3066 , P2_R1297_U6 );
nand NAND2_6502 ( P2_U5950 , P2_U3066 , P2_U3867 );
nand NAND2_6503 ( P2_U5951 , P2_U3059 , P2_R1297_U6 );
nand NAND2_6504 ( P2_U5952 , P2_U3059 , P2_U3867 );
nand NAND2_6505 ( P2_U5953 , P2_R1300_U8 , P2_R1297_U6 );
nand NAND2_6506 ( P2_U5954 , P2_U3055 , P2_U3867 );
nand NAND2_6507 ( P2_U5955 , P2_R1300_U6 , P2_R1297_U6 );
nand NAND2_6508 ( P2_U5956 , P2_U3058 , P2_U3867 );
nand NAND2_6509 ( P2_U5957 , P2_U3063 , P2_R1297_U6 );
nand NAND2_6510 ( P2_U5958 , P2_U3063 , P2_U3867 );
nand NAND2_6511 ( P2_U5959 , P2_U3054 , P2_R1297_U6 );
nand NAND2_6512 ( P2_U5960 , P2_U3054 , P2_U3867 );
nand NAND2_6513 ( P2_U5961 , P2_U3053 , P2_R1297_U6 );
nand NAND2_6514 ( P2_U5962 , P2_U3053 , P2_U3867 );
nand NAND2_6515 ( P2_U5963 , P2_U3052 , P2_R1297_U6 );
nand NAND2_6516 ( P2_U5964 , P2_U3052 , P2_U3867 );
nand NAND2_6517 ( P2_U5965 , P2_U3056 , P2_R1297_U6 );
nand NAND2_6518 ( P2_U5966 , P2_U3056 , P2_U3867 );
nand NAND2_6519 ( P2_U5967 , P2_U3057 , P2_R1297_U6 );
nand NAND2_6520 ( P2_U5968 , P2_U3057 , P2_U3867 );
nand NAND2_6521 ( P2_U5969 , P2_U3064 , P2_R1297_U6 );
nand NAND2_6522 ( P2_U5970 , P2_U3064 , P2_U3867 );
nand NAND2_6523 ( P2_U5971 , P2_U3065 , P2_R1297_U6 );
nand NAND2_6524 ( P2_U5972 , P2_U3065 , P2_U3867 );
nand NAND2_6525 ( P2_U5973 , P2_U3060 , P2_R1297_U6 );
nand NAND2_6526 ( P2_U5974 , P2_U3060 , P2_U3867 );
nand NAND2_6527 ( P2_U5975 , P2_U3074 , P2_R1297_U6 );
nand NAND2_6528 ( P2_U5976 , P2_U3074 , P2_U3867 );
nand NAND2_6529 ( P2_U5977 , P2_U3075 , P2_R1297_U6 );
nand NAND2_6530 ( P2_U5978 , P2_U3075 , P2_U3867 );
nand NAND2_6531 ( P2_U5979 , P2_U3067 , P2_R1297_U6 );
nand NAND2_6532 ( P2_U5980 , P2_U3067 , P2_U3867 );
nand NAND2_6533 ( P2_U5981 , P2_U3080 , P2_R1297_U6 );
nand NAND2_6534 ( P2_U5982 , P2_U3080 , P2_U3867 );
nand NAND2_6535 ( P2_U5983 , P2_U3081 , P2_R1297_U6 );
nand NAND2_6536 ( P2_U5984 , P2_U3081 , P2_U3867 );
nand NAND2_6537 ( P2_U5985 , P2_U3068 , P2_R1297_U6 );
nand NAND2_6538 ( P2_U5986 , P2_U3068 , P2_U3867 );
nand NAND2_6539 ( P2_U5987 , P2_U3072 , P2_R1297_U6 );
nand NAND2_6540 ( P2_U5988 , P2_U3072 , P2_U3867 );
nand NAND2_6541 ( P2_U5989 , P2_U3073 , P2_R1297_U6 );
nand NAND2_6542 ( P2_U5990 , P2_U3073 , P2_U3867 );
nand NAND2_6543 ( P2_U5991 , P2_U3078 , P2_R1297_U6 );
nand NAND2_6544 ( P2_U5992 , P2_U3078 , P2_U3867 );
nand NAND2_6545 ( P2_U5993 , P2_U3079 , P2_R1297_U6 );
nand NAND2_6546 ( P2_U5994 , P2_U3079 , P2_U3867 );
nand NAND2_6547 ( P2_U5995 , P2_U3071 , P2_R1297_U6 );
nand NAND2_6548 ( P2_U5996 , P2_U3071 , P2_U3867 );
nand NAND2_6549 ( P2_U5997 , P2_U3062 , P2_R1297_U6 );
nand NAND2_6550 ( P2_U5998 , P2_U3062 , P2_U3867 );
nand NAND2_6551 ( P2_U5999 , P2_U3061 , P2_R1297_U6 );
nand NAND2_6552 ( P2_U6000 , P2_U3061 , P2_U3867 );
nand NAND2_6553 ( P2_U6001 , P2_U3077 , P2_R1297_U6 );
nand NAND2_6554 ( P2_U6002 , P2_U3077 , P2_U3867 );
nand NAND2_6555 ( P2_U6003 , P2_U3076 , P2_R1297_U6 );
nand NAND2_6556 ( P2_U6004 , P2_U3076 , P2_U3867 );
nand NAND2_6557 ( P2_U6005 , P2_U5464 , P2_REG1_REG_9_ );
nand NAND2_6558 ( P2_U6006 , P2_U3384 , P2_REG2_REG_9_ );
nand NAND2_6559 ( P2_U6007 , P2_U5464 , P2_REG1_REG_8_ );
nand NAND2_6560 ( P2_U6008 , P2_U3384 , P2_REG2_REG_8_ );
nand NAND2_6561 ( P2_U6009 , P2_U5464 , P2_REG1_REG_7_ );
nand NAND2_6562 ( P2_U6010 , P2_U3384 , P2_REG2_REG_7_ );
nand NAND2_6563 ( P2_U6011 , P2_U5464 , P2_REG1_REG_6_ );
nand NAND2_6564 ( P2_U6012 , P2_U3384 , P2_REG2_REG_6_ );
nand NAND2_6565 ( P2_U6013 , P2_U5464 , P2_REG1_REG_5_ );
nand NAND2_6566 ( P2_U6014 , P2_U3384 , P2_REG2_REG_5_ );
nand NAND2_6567 ( P2_U6015 , P2_U5464 , P2_REG1_REG_4_ );
nand NAND2_6568 ( P2_U6016 , P2_U3384 , P2_REG2_REG_4_ );
nand NAND2_6569 ( P2_U6017 , P2_U5464 , P2_REG1_REG_3_ );
nand NAND2_6570 ( P2_U6018 , P2_U3384 , P2_REG2_REG_3_ );
nand NAND2_6571 ( P2_U6019 , P2_U5464 , P2_REG1_REG_2_ );
nand NAND2_6572 ( P2_U6020 , P2_U3384 , P2_REG2_REG_2_ );
nand NAND2_6573 ( P2_U6021 , P2_U5464 , P2_REG1_REG_19_ );
nand NAND2_6574 ( P2_U6022 , P2_U3384 , P2_REG2_REG_19_ );
nand NAND2_6575 ( P2_U6023 , P2_U5464 , P2_REG1_REG_18_ );
nand NAND2_6576 ( P2_U6024 , P2_U3384 , P2_REG2_REG_18_ );
nand NAND2_6577 ( P2_U6025 , P2_U5464 , P2_REG1_REG_17_ );
nand NAND2_6578 ( P2_U6026 , P2_U3384 , P2_REG2_REG_17_ );
nand NAND2_6579 ( P2_U6027 , P2_U5464 , P2_REG1_REG_16_ );
nand NAND2_6580 ( P2_U6028 , P2_U3384 , P2_REG2_REG_16_ );
nand NAND2_6581 ( P2_U6029 , P2_U5464 , P2_REG1_REG_15_ );
nand NAND2_6582 ( P2_U6030 , P2_U3384 , P2_REG2_REG_15_ );
nand NAND2_6583 ( P2_U6031 , P2_U5464 , P2_REG1_REG_14_ );
nand NAND2_6584 ( P2_U6032 , P2_U3384 , P2_REG2_REG_14_ );
nand NAND2_6585 ( P2_U6033 , P2_U5464 , P2_REG1_REG_13_ );
nand NAND2_6586 ( P2_U6034 , P2_U3384 , P2_REG2_REG_13_ );
nand NAND2_6587 ( P2_U6035 , P2_U5464 , P2_REG1_REG_12_ );
nand NAND2_6588 ( P2_U6036 , P2_U3384 , P2_REG2_REG_12_ );
nand NAND2_6589 ( P2_U6037 , P2_U5464 , P2_REG1_REG_11_ );
nand NAND2_6590 ( P2_U6038 , P2_U3384 , P2_REG2_REG_11_ );
nand NAND2_6591 ( P2_U6039 , P2_U5464 , P2_REG1_REG_10_ );
nand NAND2_6592 ( P2_U6040 , P2_U3384 , P2_REG2_REG_10_ );
nand NAND2_6593 ( P2_U6041 , P2_U5464 , P2_REG1_REG_1_ );
nand NAND2_6594 ( P2_U6042 , P2_U3384 , P2_REG2_REG_1_ );
nand NAND2_6595 ( P2_U6043 , P2_U5464 , P2_REG1_REG_0_ );
nand NAND2_6596 ( P2_U6044 , P2_U3384 , P2_REG2_REG_0_ );
nand NAND2_6597 ( P2_R1161_U465 , P2_R1161_U464 , P2_R1161_U463 );
nand NAND2_6598 ( P2_R1161_U464 , P2_U3443 , P2_R1161_U76 );
nand NAND2_6599 ( P2_R1161_U463 , P2_U3081 , P2_R1161_U75 );
nand NAND2_6600 ( P2_R1161_U462 , P2_R1161_U460 , P2_R1161_U316 );
nand NAND2_6601 ( P2_R1161_U461 , P2_R1161_U359 , P2_R1161_U91 );
nand NAND2_6602 ( P2_R1161_U460 , P2_R1161_U459 , P2_R1161_U458 );
nand NAND2_6603 ( P2_R1161_U459 , P2_U3445 , P2_R1161_U79 );
nand NAND2_6604 ( P2_R1161_U458 , P2_U3080 , P2_R1161_U78 );
nand NAND2_6605 ( P2_R1161_U457 , P2_R1161_U328 , P2_R1161_U31 );
nand NAND2_6606 ( P2_R1161_U456 , P2_R1161_U182 , P2_R1161_U161 );
nand NAND2_6607 ( P2_R1161_U455 , P2_U3903 , P2_R1161_U90 );
nand NAND2_6608 ( P2_R1161_U454 , P2_U3075 , P2_R1161_U81 );
nand NAND2_6609 ( P2_R1161_U453 , P2_R1161_U452 , P2_R1161_U451 );
nand NAND2_6610 ( P2_R1161_U452 , P2_U3902 , P2_R1161_U55 );
nand NAND2_6611 ( P2_R1161_U451 , P2_U3074 , P2_R1161_U54 );
nand NAND2_6612 ( P2_R1161_U450 , P2_U3902 , P2_R1161_U55 );
nand NAND2_6613 ( P2_R1161_U449 , P2_U3074 , P2_R1161_U54 );
nand NAND2_6614 ( P2_R1161_U448 , P2_R1161_U286 , P2_R1161_U446 );
nand NAND2_6615 ( P2_R1161_U447 , P2_R1161_U158 , P2_R1161_U159 );
not NOT1_6616 ( LT_1075_U6 , P1_ADDR_REG_19_ );
and AND2_6617 ( ADD_1068_U4 , ADD_1068_U159 , ADD_1068_U155 );
nand NAND3_6618 ( ADD_1068_U5 , ADD_1068_U221 , ADD_1068_U220 , ADD_1068_U160 );
not NOT1_6619 ( ADD_1068_U6 , P1_ADDR_REG_0_ );
not NOT1_6620 ( ADD_1068_U7 , P2_ADDR_REG_0_ );
not NOT1_6621 ( ADD_1068_U8 , P2_ADDR_REG_1_ );
nand NAND2_6622 ( ADD_1068_U9 , P2_ADDR_REG_0_ , P1_ADDR_REG_0_ );
not NOT1_6623 ( ADD_1068_U10 , P1_ADDR_REG_1_ );
not NOT1_6624 ( ADD_1068_U11 , P1_ADDR_REG_2_ );
not NOT1_6625 ( ADD_1068_U12 , P2_ADDR_REG_2_ );
not NOT1_6626 ( ADD_1068_U13 , P1_ADDR_REG_3_ );
not NOT1_6627 ( ADD_1068_U14 , P2_ADDR_REG_3_ );
not NOT1_6628 ( ADD_1068_U15 , P1_ADDR_REG_4_ );
not NOT1_6629 ( ADD_1068_U16 , P2_ADDR_REG_4_ );
not NOT1_6630 ( ADD_1068_U17 , P1_ADDR_REG_5_ );
not NOT1_6631 ( ADD_1068_U18 , P2_ADDR_REG_5_ );
not NOT1_6632 ( ADD_1068_U19 , P1_ADDR_REG_6_ );
not NOT1_6633 ( ADD_1068_U20 , P2_ADDR_REG_6_ );
not NOT1_6634 ( ADD_1068_U21 , P1_ADDR_REG_7_ );
not NOT1_6635 ( ADD_1068_U22 , P2_ADDR_REG_7_ );
not NOT1_6636 ( ADD_1068_U23 , P1_ADDR_REG_8_ );
not NOT1_6637 ( ADD_1068_U24 , P2_ADDR_REG_8_ );
not NOT1_6638 ( ADD_1068_U25 , P2_ADDR_REG_9_ );
not NOT1_6639 ( ADD_1068_U26 , P1_ADDR_REG_9_ );
not NOT1_6640 ( ADD_1068_U27 , P1_ADDR_REG_10_ );
not NOT1_6641 ( ADD_1068_U28 , P2_ADDR_REG_10_ );
not NOT1_6642 ( ADD_1068_U29 , P1_ADDR_REG_11_ );
not NOT1_6643 ( ADD_1068_U30 , P2_ADDR_REG_11_ );
not NOT1_6644 ( ADD_1068_U31 , P1_ADDR_REG_12_ );
not NOT1_6645 ( ADD_1068_U32 , P2_ADDR_REG_12_ );
not NOT1_6646 ( ADD_1068_U33 , P1_ADDR_REG_13_ );
not NOT1_6647 ( ADD_1068_U34 , P2_ADDR_REG_13_ );
not NOT1_6648 ( ADD_1068_U35 , P1_ADDR_REG_14_ );
not NOT1_6649 ( ADD_1068_U36 , P2_ADDR_REG_14_ );
not NOT1_6650 ( ADD_1068_U37 , P1_ADDR_REG_15_ );
not NOT1_6651 ( ADD_1068_U38 , P2_ADDR_REG_15_ );
not NOT1_6652 ( ADD_1068_U39 , P1_ADDR_REG_16_ );
not NOT1_6653 ( ADD_1068_U40 , P2_ADDR_REG_16_ );
not NOT1_6654 ( ADD_1068_U41 , P1_ADDR_REG_17_ );
not NOT1_6655 ( ADD_1068_U42 , P2_ADDR_REG_17_ );
not NOT1_6656 ( ADD_1068_U43 , P1_ADDR_REG_18_ );
not NOT1_6657 ( ADD_1068_U44 , P2_ADDR_REG_18_ );
nand NAND2_6658 ( ADD_1068_U45 , ADD_1068_U150 , ADD_1068_U149 );
nand NAND2_6659 ( ADD_1068_U46 , ADD_1068_U291 , ADD_1068_U290 );
nand NAND2_6660 ( ADD_1068_U47 , ADD_1068_U167 , ADD_1068_U166 );
nand NAND2_6661 ( ADD_1068_U48 , ADD_1068_U174 , ADD_1068_U173 );
nand NAND2_6662 ( ADD_1068_U49 , ADD_1068_U181 , ADD_1068_U180 );
nand NAND2_6663 ( ADD_1068_U50 , ADD_1068_U188 , ADD_1068_U187 );
nand NAND2_6664 ( ADD_1068_U51 , ADD_1068_U195 , ADD_1068_U194 );
nand NAND2_6665 ( ADD_1068_U52 , ADD_1068_U202 , ADD_1068_U201 );
nand NAND2_6666 ( ADD_1068_U53 , ADD_1068_U209 , ADD_1068_U208 );
nand NAND2_6667 ( ADD_1068_U54 , ADD_1068_U216 , ADD_1068_U215 );
nand NAND2_6668 ( ADD_1068_U55 , ADD_1068_U233 , ADD_1068_U232 );
nand NAND2_6669 ( ADD_1068_U56 , ADD_1068_U240 , ADD_1068_U239 );
nand NAND2_6670 ( ADD_1068_U57 , ADD_1068_U247 , ADD_1068_U246 );
nand NAND2_6671 ( ADD_1068_U58 , ADD_1068_U254 , ADD_1068_U253 );
nand NAND2_6672 ( ADD_1068_U59 , ADD_1068_U261 , ADD_1068_U260 );
nand NAND2_6673 ( ADD_1068_U60 , ADD_1068_U268 , ADD_1068_U267 );
nand NAND2_6674 ( ADD_1068_U61 , ADD_1068_U275 , ADD_1068_U274 );
nand NAND2_6675 ( ADD_1068_U62 , ADD_1068_U282 , ADD_1068_U281 );
nand NAND2_6676 ( ADD_1068_U63 , ADD_1068_U289 , ADD_1068_U288 );
nand NAND2_6677 ( ADD_1068_U64 , ADD_1068_U114 , ADD_1068_U113 );
nand NAND2_6678 ( ADD_1068_U65 , ADD_1068_U110 , ADD_1068_U109 );
nand NAND2_6679 ( ADD_1068_U66 , ADD_1068_U106 , ADD_1068_U105 );
nand NAND2_6680 ( ADD_1068_U67 , ADD_1068_U102 , ADD_1068_U101 );
nand NAND2_6681 ( ADD_1068_U68 , ADD_1068_U98 , ADD_1068_U97 );
nand NAND2_6682 ( ADD_1068_U69 , ADD_1068_U94 , ADD_1068_U93 );
nand NAND2_6683 ( ADD_1068_U70 , ADD_1068_U90 , ADD_1068_U89 );
nand NAND2_6684 ( ADD_1068_U71 , ADD_1068_U72 , ADD_1068_U86 );
nand NAND2_6685 ( ADD_1068_U72 , P1_ADDR_REG_1_ , ADD_1068_U84 );
not NOT1_6686 ( ADD_1068_U73 , P2_ADDR_REG_19_ );
not NOT1_6687 ( ADD_1068_U74 , P1_ADDR_REG_19_ );
nand NAND2_6688 ( ADD_1068_U75 , ADD_1068_U146 , ADD_1068_U145 );
nand NAND2_6689 ( ADD_1068_U76 , ADD_1068_U142 , ADD_1068_U141 );
nand NAND2_6690 ( ADD_1068_U77 , ADD_1068_U138 , ADD_1068_U137 );
nand NAND2_6691 ( ADD_1068_U78 , ADD_1068_U134 , ADD_1068_U133 );
nand NAND2_6692 ( ADD_1068_U79 , ADD_1068_U130 , ADD_1068_U129 );
nand NAND2_6693 ( ADD_1068_U80 , ADD_1068_U126 , ADD_1068_U125 );
nand NAND2_6694 ( ADD_1068_U81 , ADD_1068_U122 , ADD_1068_U121 );
nand NAND2_6695 ( ADD_1068_U82 , ADD_1068_U118 , ADD_1068_U117 );
not NOT1_6696 ( ADD_1068_U83 , ADD_1068_U72 );
not NOT1_6697 ( ADD_1068_U84 , ADD_1068_U9 );
nand NAND2_6698 ( ADD_1068_U85 , ADD_1068_U10 , ADD_1068_U9 );
nand NAND2_6699 ( ADD_1068_U86 , P2_ADDR_REG_1_ , ADD_1068_U85 );
not NOT1_6700 ( ADD_1068_U87 , ADD_1068_U71 );
or OR2_6701 ( ADD_1068_U88 , P1_ADDR_REG_2_ , P2_ADDR_REG_2_ );
nand NAND2_6702 ( ADD_1068_U89 , ADD_1068_U88 , ADD_1068_U71 );
nand NAND2_6703 ( ADD_1068_U90 , P2_ADDR_REG_2_ , P1_ADDR_REG_2_ );
not NOT1_6704 ( ADD_1068_U91 , ADD_1068_U70 );
or OR2_6705 ( ADD_1068_U92 , P1_ADDR_REG_3_ , P2_ADDR_REG_3_ );
nand NAND2_6706 ( ADD_1068_U93 , ADD_1068_U92 , ADD_1068_U70 );
nand NAND2_6707 ( ADD_1068_U94 , P2_ADDR_REG_3_ , P1_ADDR_REG_3_ );
not NOT1_6708 ( ADD_1068_U95 , ADD_1068_U69 );
or OR2_6709 ( ADD_1068_U96 , P1_ADDR_REG_4_ , P2_ADDR_REG_4_ );
nand NAND2_6710 ( ADD_1068_U97 , ADD_1068_U96 , ADD_1068_U69 );
nand NAND2_6711 ( ADD_1068_U98 , P2_ADDR_REG_4_ , P1_ADDR_REG_4_ );
not NOT1_6712 ( ADD_1068_U99 , ADD_1068_U68 );
or OR2_6713 ( ADD_1068_U100 , P1_ADDR_REG_5_ , P2_ADDR_REG_5_ );
nand NAND2_6714 ( ADD_1068_U101 , ADD_1068_U100 , ADD_1068_U68 );
nand NAND2_6715 ( ADD_1068_U102 , P2_ADDR_REG_5_ , P1_ADDR_REG_5_ );
not NOT1_6716 ( ADD_1068_U103 , ADD_1068_U67 );
or OR2_6717 ( ADD_1068_U104 , P1_ADDR_REG_6_ , P2_ADDR_REG_6_ );
nand NAND2_6718 ( ADD_1068_U105 , ADD_1068_U104 , ADD_1068_U67 );
nand NAND2_6719 ( ADD_1068_U106 , P2_ADDR_REG_6_ , P1_ADDR_REG_6_ );
not NOT1_6720 ( ADD_1068_U107 , ADD_1068_U66 );
or OR2_6721 ( ADD_1068_U108 , P1_ADDR_REG_7_ , P2_ADDR_REG_7_ );
nand NAND2_6722 ( ADD_1068_U109 , ADD_1068_U108 , ADD_1068_U66 );
nand NAND2_6723 ( ADD_1068_U110 , P2_ADDR_REG_7_ , P1_ADDR_REG_7_ );
not NOT1_6724 ( ADD_1068_U111 , ADD_1068_U65 );
or OR2_6725 ( ADD_1068_U112 , P1_ADDR_REG_8_ , P2_ADDR_REG_8_ );
nand NAND2_6726 ( ADD_1068_U113 , ADD_1068_U112 , ADD_1068_U65 );
nand NAND2_6727 ( ADD_1068_U114 , P2_ADDR_REG_8_ , P1_ADDR_REG_8_ );
not NOT1_6728 ( ADD_1068_U115 , ADD_1068_U64 );
or OR2_6729 ( ADD_1068_U116 , P1_ADDR_REG_9_ , P2_ADDR_REG_9_ );
nand NAND2_6730 ( ADD_1068_U117 , ADD_1068_U116 , ADD_1068_U64 );
nand NAND2_6731 ( ADD_1068_U118 , P1_ADDR_REG_9_ , P2_ADDR_REG_9_ );
not NOT1_6732 ( ADD_1068_U119 , ADD_1068_U82 );
or OR2_6733 ( ADD_1068_U120 , P1_ADDR_REG_10_ , P2_ADDR_REG_10_ );
nand NAND2_6734 ( ADD_1068_U121 , ADD_1068_U120 , ADD_1068_U82 );
nand NAND2_6735 ( ADD_1068_U122 , P2_ADDR_REG_10_ , P1_ADDR_REG_10_ );
not NOT1_6736 ( ADD_1068_U123 , ADD_1068_U81 );
or OR2_6737 ( ADD_1068_U124 , P1_ADDR_REG_11_ , P2_ADDR_REG_11_ );
nand NAND2_6738 ( ADD_1068_U125 , ADD_1068_U124 , ADD_1068_U81 );
nand NAND2_6739 ( ADD_1068_U126 , P2_ADDR_REG_11_ , P1_ADDR_REG_11_ );
not NOT1_6740 ( ADD_1068_U127 , ADD_1068_U80 );
or OR2_6741 ( ADD_1068_U128 , P1_ADDR_REG_12_ , P2_ADDR_REG_12_ );
nand NAND2_6742 ( ADD_1068_U129 , ADD_1068_U128 , ADD_1068_U80 );
nand NAND2_6743 ( ADD_1068_U130 , P2_ADDR_REG_12_ , P1_ADDR_REG_12_ );
not NOT1_6744 ( ADD_1068_U131 , ADD_1068_U79 );
or OR2_6745 ( ADD_1068_U132 , P1_ADDR_REG_13_ , P2_ADDR_REG_13_ );
nand NAND2_6746 ( ADD_1068_U133 , ADD_1068_U132 , ADD_1068_U79 );
nand NAND2_6747 ( ADD_1068_U134 , P2_ADDR_REG_13_ , P1_ADDR_REG_13_ );
not NOT1_6748 ( ADD_1068_U135 , ADD_1068_U78 );
or OR2_6749 ( ADD_1068_U136 , P1_ADDR_REG_14_ , P2_ADDR_REG_14_ );
nand NAND2_6750 ( ADD_1068_U137 , ADD_1068_U136 , ADD_1068_U78 );
nand NAND2_6751 ( ADD_1068_U138 , P2_ADDR_REG_14_ , P1_ADDR_REG_14_ );
not NOT1_6752 ( ADD_1068_U139 , ADD_1068_U77 );
or OR2_6753 ( ADD_1068_U140 , P1_ADDR_REG_15_ , P2_ADDR_REG_15_ );
nand NAND2_6754 ( ADD_1068_U141 , ADD_1068_U140 , ADD_1068_U77 );
nand NAND2_6755 ( ADD_1068_U142 , P2_ADDR_REG_15_ , P1_ADDR_REG_15_ );
not NOT1_6756 ( ADD_1068_U143 , ADD_1068_U76 );
or OR2_6757 ( ADD_1068_U144 , P1_ADDR_REG_16_ , P2_ADDR_REG_16_ );
nand NAND2_6758 ( ADD_1068_U145 , ADD_1068_U144 , ADD_1068_U76 );
nand NAND2_6759 ( ADD_1068_U146 , P2_ADDR_REG_16_ , P1_ADDR_REG_16_ );
not NOT1_6760 ( ADD_1068_U147 , ADD_1068_U75 );
or OR2_6761 ( ADD_1068_U148 , P1_ADDR_REG_17_ , P2_ADDR_REG_17_ );
nand NAND2_6762 ( ADD_1068_U149 , ADD_1068_U148 , ADD_1068_U75 );
nand NAND2_6763 ( ADD_1068_U150 , P2_ADDR_REG_17_ , P1_ADDR_REG_17_ );
not NOT1_6764 ( ADD_1068_U151 , ADD_1068_U45 );
or OR2_6765 ( ADD_1068_U152 , P1_ADDR_REG_18_ , P2_ADDR_REG_18_ );
nand NAND2_6766 ( ADD_1068_U153 , ADD_1068_U152 , ADD_1068_U45 );
nand NAND2_6767 ( ADD_1068_U154 , P2_ADDR_REG_18_ , P1_ADDR_REG_18_ );
nand NAND4_6768 ( ADD_1068_U155 , ADD_1068_U223 , ADD_1068_U222 , ADD_1068_U154 , ADD_1068_U153 );
nand NAND2_6769 ( ADD_1068_U156 , P2_ADDR_REG_18_ , P1_ADDR_REG_18_ );
nand NAND2_6770 ( ADD_1068_U157 , ADD_1068_U151 , ADD_1068_U156 );
or OR2_6771 ( ADD_1068_U158 , P2_ADDR_REG_18_ , P1_ADDR_REG_18_ );
nand NAND3_6772 ( ADD_1068_U159 , ADD_1068_U158 , ADD_1068_U226 , ADD_1068_U157 );
nand NAND2_6773 ( ADD_1068_U160 , ADD_1068_U219 , ADD_1068_U10 );
nand NAND2_6774 ( ADD_1068_U161 , P2_ADDR_REG_9_ , ADD_1068_U26 );
nand NAND2_6775 ( ADD_1068_U162 , P1_ADDR_REG_9_ , ADD_1068_U25 );
nand NAND2_6776 ( ADD_1068_U163 , P2_ADDR_REG_9_ , ADD_1068_U26 );
nand NAND2_6777 ( ADD_1068_U164 , P1_ADDR_REG_9_ , ADD_1068_U25 );
nand NAND2_6778 ( ADD_1068_U165 , ADD_1068_U164 , ADD_1068_U163 );
nand NAND3_6779 ( ADD_1068_U166 , ADD_1068_U162 , ADD_1068_U161 , ADD_1068_U64 );
nand NAND2_6780 ( ADD_1068_U167 , ADD_1068_U115 , ADD_1068_U165 );
nand NAND2_6781 ( ADD_1068_U168 , P2_ADDR_REG_8_ , ADD_1068_U23 );
nand NAND2_6782 ( ADD_1068_U169 , P1_ADDR_REG_8_ , ADD_1068_U24 );
nand NAND2_6783 ( ADD_1068_U170 , P2_ADDR_REG_8_ , ADD_1068_U23 );
nand NAND2_6784 ( ADD_1068_U171 , P1_ADDR_REG_8_ , ADD_1068_U24 );
nand NAND2_6785 ( ADD_1068_U172 , ADD_1068_U171 , ADD_1068_U170 );
nand NAND3_6786 ( ADD_1068_U173 , ADD_1068_U169 , ADD_1068_U168 , ADD_1068_U65 );
nand NAND2_6787 ( ADD_1068_U174 , ADD_1068_U111 , ADD_1068_U172 );
nand NAND2_6788 ( ADD_1068_U175 , P2_ADDR_REG_7_ , ADD_1068_U21 );
nand NAND2_6789 ( ADD_1068_U176 , P1_ADDR_REG_7_ , ADD_1068_U22 );
nand NAND2_6790 ( ADD_1068_U177 , P2_ADDR_REG_7_ , ADD_1068_U21 );
nand NAND2_6791 ( ADD_1068_U178 , P1_ADDR_REG_7_ , ADD_1068_U22 );
nand NAND2_6792 ( ADD_1068_U179 , ADD_1068_U178 , ADD_1068_U177 );
nand NAND3_6793 ( ADD_1068_U180 , ADD_1068_U176 , ADD_1068_U175 , ADD_1068_U66 );
nand NAND2_6794 ( ADD_1068_U181 , ADD_1068_U107 , ADD_1068_U179 );
nand NAND2_6795 ( ADD_1068_U182 , P2_ADDR_REG_6_ , ADD_1068_U19 );
nand NAND2_6796 ( ADD_1068_U183 , P1_ADDR_REG_6_ , ADD_1068_U20 );
nand NAND2_6797 ( ADD_1068_U184 , P2_ADDR_REG_6_ , ADD_1068_U19 );
nand NAND2_6798 ( ADD_1068_U185 , P1_ADDR_REG_6_ , ADD_1068_U20 );
nand NAND2_6799 ( ADD_1068_U186 , ADD_1068_U185 , ADD_1068_U184 );
nand NAND3_6800 ( ADD_1068_U187 , ADD_1068_U183 , ADD_1068_U182 , ADD_1068_U67 );
nand NAND2_6801 ( ADD_1068_U188 , ADD_1068_U103 , ADD_1068_U186 );
nand NAND2_6802 ( ADD_1068_U189 , P2_ADDR_REG_5_ , ADD_1068_U17 );
nand NAND2_6803 ( ADD_1068_U190 , P1_ADDR_REG_5_ , ADD_1068_U18 );
nand NAND2_6804 ( ADD_1068_U191 , P2_ADDR_REG_5_ , ADD_1068_U17 );
nand NAND2_6805 ( ADD_1068_U192 , P1_ADDR_REG_5_ , ADD_1068_U18 );
nand NAND2_6806 ( ADD_1068_U193 , ADD_1068_U192 , ADD_1068_U191 );
nand NAND3_6807 ( ADD_1068_U194 , ADD_1068_U190 , ADD_1068_U189 , ADD_1068_U68 );
nand NAND2_6808 ( ADD_1068_U195 , ADD_1068_U99 , ADD_1068_U193 );
nand NAND2_6809 ( ADD_1068_U196 , P2_ADDR_REG_4_ , ADD_1068_U15 );
nand NAND2_6810 ( ADD_1068_U197 , P1_ADDR_REG_4_ , ADD_1068_U16 );
nand NAND2_6811 ( ADD_1068_U198 , P2_ADDR_REG_4_ , ADD_1068_U15 );
nand NAND2_6812 ( ADD_1068_U199 , P1_ADDR_REG_4_ , ADD_1068_U16 );
nand NAND2_6813 ( ADD_1068_U200 , ADD_1068_U199 , ADD_1068_U198 );
nand NAND3_6814 ( ADD_1068_U201 , ADD_1068_U197 , ADD_1068_U196 , ADD_1068_U69 );
nand NAND2_6815 ( ADD_1068_U202 , ADD_1068_U95 , ADD_1068_U200 );
nand NAND2_6816 ( ADD_1068_U203 , P2_ADDR_REG_3_ , ADD_1068_U13 );
nand NAND2_6817 ( ADD_1068_U204 , P1_ADDR_REG_3_ , ADD_1068_U14 );
nand NAND2_6818 ( ADD_1068_U205 , P2_ADDR_REG_3_ , ADD_1068_U13 );
nand NAND2_6819 ( ADD_1068_U206 , P1_ADDR_REG_3_ , ADD_1068_U14 );
nand NAND2_6820 ( ADD_1068_U207 , ADD_1068_U206 , ADD_1068_U205 );
nand NAND3_6821 ( ADD_1068_U208 , ADD_1068_U204 , ADD_1068_U203 , ADD_1068_U70 );
nand NAND2_6822 ( ADD_1068_U209 , ADD_1068_U91 , ADD_1068_U207 );
nand NAND2_6823 ( ADD_1068_U210 , P2_ADDR_REG_2_ , ADD_1068_U11 );
nand NAND2_6824 ( ADD_1068_U211 , P1_ADDR_REG_2_ , ADD_1068_U12 );
nand NAND2_6825 ( ADD_1068_U212 , P2_ADDR_REG_2_ , ADD_1068_U11 );
nand NAND2_6826 ( ADD_1068_U213 , P1_ADDR_REG_2_ , ADD_1068_U12 );
nand NAND2_6827 ( ADD_1068_U214 , ADD_1068_U213 , ADD_1068_U212 );
nand NAND3_6828 ( ADD_1068_U215 , ADD_1068_U211 , ADD_1068_U210 , ADD_1068_U71 );
nand NAND2_6829 ( ADD_1068_U216 , ADD_1068_U87 , ADD_1068_U214 );
nand NAND2_6830 ( ADD_1068_U217 , P2_ADDR_REG_1_ , ADD_1068_U9 );
nand NAND2_6831 ( ADD_1068_U218 , ADD_1068_U84 , ADD_1068_U8 );
nand NAND2_6832 ( ADD_1068_U219 , ADD_1068_U218 , ADD_1068_U217 );
nand NAND3_6833 ( ADD_1068_U220 , P1_ADDR_REG_1_ , ADD_1068_U9 , ADD_1068_U8 );
nand NAND2_6834 ( ADD_1068_U221 , ADD_1068_U83 , P2_ADDR_REG_1_ );
nand NAND2_6835 ( ADD_1068_U222 , P2_ADDR_REG_19_ , ADD_1068_U74 );
nand NAND2_6836 ( ADD_1068_U223 , P1_ADDR_REG_19_ , ADD_1068_U73 );
nand NAND2_6837 ( ADD_1068_U224 , P2_ADDR_REG_19_ , ADD_1068_U74 );
nand NAND2_6838 ( ADD_1068_U225 , P1_ADDR_REG_19_ , ADD_1068_U73 );
nand NAND2_6839 ( ADD_1068_U226 , ADD_1068_U225 , ADD_1068_U224 );
nand NAND2_6840 ( ADD_1068_U227 , P2_ADDR_REG_18_ , ADD_1068_U43 );
nand NAND2_6841 ( ADD_1068_U228 , P1_ADDR_REG_18_ , ADD_1068_U44 );
nand NAND2_6842 ( ADD_1068_U229 , P2_ADDR_REG_18_ , ADD_1068_U43 );
nand NAND2_6843 ( ADD_1068_U230 , P1_ADDR_REG_18_ , ADD_1068_U44 );
nand NAND2_6844 ( ADD_1068_U231 , ADD_1068_U230 , ADD_1068_U229 );
nand NAND3_6845 ( ADD_1068_U232 , ADD_1068_U228 , ADD_1068_U227 , ADD_1068_U45 );
nand NAND2_6846 ( ADD_1068_U233 , ADD_1068_U231 , ADD_1068_U151 );
nand NAND2_6847 ( ADD_1068_U234 , P2_ADDR_REG_17_ , ADD_1068_U41 );
nand NAND2_6848 ( ADD_1068_U235 , P1_ADDR_REG_17_ , ADD_1068_U42 );
nand NAND2_6849 ( ADD_1068_U236 , P2_ADDR_REG_17_ , ADD_1068_U41 );
nand NAND2_6850 ( ADD_1068_U237 , P1_ADDR_REG_17_ , ADD_1068_U42 );
nand NAND2_6851 ( ADD_1068_U238 , ADD_1068_U237 , ADD_1068_U236 );
nand NAND3_6852 ( ADD_1068_U239 , ADD_1068_U235 , ADD_1068_U234 , ADD_1068_U75 );
nand NAND2_6853 ( ADD_1068_U240 , ADD_1068_U147 , ADD_1068_U238 );
nand NAND2_6854 ( ADD_1068_U241 , P2_ADDR_REG_16_ , ADD_1068_U39 );
nand NAND2_6855 ( ADD_1068_U242 , P1_ADDR_REG_16_ , ADD_1068_U40 );
nand NAND2_6856 ( ADD_1068_U243 , P2_ADDR_REG_16_ , ADD_1068_U39 );
nand NAND2_6857 ( ADD_1068_U244 , P1_ADDR_REG_16_ , ADD_1068_U40 );
nand NAND2_6858 ( ADD_1068_U245 , ADD_1068_U244 , ADD_1068_U243 );
nand NAND3_6859 ( ADD_1068_U246 , ADD_1068_U242 , ADD_1068_U241 , ADD_1068_U76 );
nand NAND2_6860 ( ADD_1068_U247 , ADD_1068_U143 , ADD_1068_U245 );
nand NAND2_6861 ( ADD_1068_U248 , P2_ADDR_REG_15_ , ADD_1068_U37 );
nand NAND2_6862 ( ADD_1068_U249 , P1_ADDR_REG_15_ , ADD_1068_U38 );
nand NAND2_6863 ( ADD_1068_U250 , P2_ADDR_REG_15_ , ADD_1068_U37 );
nand NAND2_6864 ( ADD_1068_U251 , P1_ADDR_REG_15_ , ADD_1068_U38 );
nand NAND2_6865 ( ADD_1068_U252 , ADD_1068_U251 , ADD_1068_U250 );
nand NAND3_6866 ( ADD_1068_U253 , ADD_1068_U249 , ADD_1068_U248 , ADD_1068_U77 );
nand NAND2_6867 ( ADD_1068_U254 , ADD_1068_U139 , ADD_1068_U252 );
nand NAND2_6868 ( ADD_1068_U255 , P2_ADDR_REG_14_ , ADD_1068_U35 );
nand NAND2_6869 ( ADD_1068_U256 , P1_ADDR_REG_14_ , ADD_1068_U36 );
nand NAND2_6870 ( ADD_1068_U257 , P2_ADDR_REG_14_ , ADD_1068_U35 );
nand NAND2_6871 ( ADD_1068_U258 , P1_ADDR_REG_14_ , ADD_1068_U36 );
nand NAND2_6872 ( ADD_1068_U259 , ADD_1068_U258 , ADD_1068_U257 );
nand NAND3_6873 ( ADD_1068_U260 , ADD_1068_U256 , ADD_1068_U255 , ADD_1068_U78 );
nand NAND2_6874 ( ADD_1068_U261 , ADD_1068_U135 , ADD_1068_U259 );
nand NAND2_6875 ( ADD_1068_U262 , P2_ADDR_REG_13_ , ADD_1068_U33 );
nand NAND2_6876 ( ADD_1068_U263 , P1_ADDR_REG_13_ , ADD_1068_U34 );
nand NAND2_6877 ( ADD_1068_U264 , P2_ADDR_REG_13_ , ADD_1068_U33 );
nand NAND2_6878 ( ADD_1068_U265 , P1_ADDR_REG_13_ , ADD_1068_U34 );
nand NAND2_6879 ( ADD_1068_U266 , ADD_1068_U265 , ADD_1068_U264 );
nand NAND3_6880 ( ADD_1068_U267 , ADD_1068_U263 , ADD_1068_U262 , ADD_1068_U79 );
nand NAND2_6881 ( ADD_1068_U268 , ADD_1068_U131 , ADD_1068_U266 );
nand NAND2_6882 ( ADD_1068_U269 , P2_ADDR_REG_12_ , ADD_1068_U31 );
nand NAND2_6883 ( ADD_1068_U270 , P1_ADDR_REG_12_ , ADD_1068_U32 );
nand NAND2_6884 ( ADD_1068_U271 , P2_ADDR_REG_12_ , ADD_1068_U31 );
nand NAND2_6885 ( ADD_1068_U272 , P1_ADDR_REG_12_ , ADD_1068_U32 );
nand NAND2_6886 ( ADD_1068_U273 , ADD_1068_U272 , ADD_1068_U271 );
nand NAND3_6887 ( ADD_1068_U274 , ADD_1068_U270 , ADD_1068_U269 , ADD_1068_U80 );
nand NAND2_6888 ( ADD_1068_U275 , ADD_1068_U127 , ADD_1068_U273 );
nand NAND2_6889 ( ADD_1068_U276 , P2_ADDR_REG_11_ , ADD_1068_U29 );
nand NAND2_6890 ( ADD_1068_U277 , P1_ADDR_REG_11_ , ADD_1068_U30 );
nand NAND2_6891 ( ADD_1068_U278 , P2_ADDR_REG_11_ , ADD_1068_U29 );
nand NAND2_6892 ( ADD_1068_U279 , P1_ADDR_REG_11_ , ADD_1068_U30 );
nand NAND2_6893 ( ADD_1068_U280 , ADD_1068_U279 , ADD_1068_U278 );
nand NAND3_6894 ( ADD_1068_U281 , ADD_1068_U277 , ADD_1068_U276 , ADD_1068_U81 );
nand NAND2_6895 ( ADD_1068_U282 , ADD_1068_U123 , ADD_1068_U280 );
nand NAND2_6896 ( ADD_1068_U283 , P2_ADDR_REG_10_ , ADD_1068_U27 );
nand NAND2_6897 ( ADD_1068_U284 , P1_ADDR_REG_10_ , ADD_1068_U28 );
nand NAND2_6898 ( ADD_1068_U285 , P2_ADDR_REG_10_ , ADD_1068_U27 );
nand NAND2_6899 ( ADD_1068_U286 , P1_ADDR_REG_10_ , ADD_1068_U28 );
nand NAND2_6900 ( ADD_1068_U287 , ADD_1068_U286 , ADD_1068_U285 );
nand NAND3_6901 ( ADD_1068_U288 , ADD_1068_U284 , ADD_1068_U283 , ADD_1068_U82 );
nand NAND2_6902 ( ADD_1068_U289 , ADD_1068_U119 , ADD_1068_U287 );
nand NAND2_6903 ( ADD_1068_U290 , P2_ADDR_REG_0_ , ADD_1068_U6 );
nand NAND2_6904 ( ADD_1068_U291 , P1_ADDR_REG_0_ , ADD_1068_U7 );
and AND2_6905 ( R140_U4 , R140_U197 , R140_U195 );
and AND2_6906 ( R140_U5 , R140_U203 , R140_U201 );
and AND2_6907 ( R140_U6 , R140_U5 , R140_U205 );
and AND2_6908 ( R140_U7 , R140_U213 , R140_U209 );
and AND2_6909 ( R140_U8 , R140_U7 , R140_U216 );
and AND2_6910 ( R140_U9 , R140_U378 , R140_U377 );
nand NAND3_6911 ( R140_U10 , R140_U469 , R140_U468 , R140_U324 );
and AND2_6912 ( R140_U11 , R140_U124 , R140_U323 );
not NOT1_6913 ( R140_U12 , SI_8_ );
not NOT1_6914 ( R140_U13 , U90 );
not NOT1_6915 ( R140_U14 , SI_7_ );
not NOT1_6916 ( R140_U15 , U91 );
nand NAND2_6917 ( R140_U16 , U91 , SI_7_ );
not NOT1_6918 ( R140_U17 , SI_6_ );
not NOT1_6919 ( R140_U18 , U92 );
not NOT1_6920 ( R140_U19 , SI_5_ );
not NOT1_6921 ( R140_U20 , U93 );
not NOT1_6922 ( R140_U21 , SI_4_ );
not NOT1_6923 ( R140_U22 , U94 );
nand NAND2_6924 ( R140_U23 , U94 , SI_4_ );
not NOT1_6925 ( R140_U24 , SI_3_ );
not NOT1_6926 ( R140_U25 , U97 );
not NOT1_6927 ( R140_U26 , SI_2_ );
not NOT1_6928 ( R140_U27 , U108 );
nand NAND2_6929 ( R140_U28 , U108 , SI_2_ );
not NOT1_6930 ( R140_U29 , SI_1_ );
not NOT1_6931 ( R140_U30 , SI_0_ );
not NOT1_6932 ( R140_U31 , U120 );
not NOT1_6933 ( R140_U32 , U119 );
not NOT1_6934 ( R140_U33 , U89 );
not NOT1_6935 ( R140_U34 , SI_9_ );
nand NAND2_6936 ( R140_U35 , R140_U288 , R140_U198 );
not NOT1_6937 ( R140_U36 , SI_14_ );
not NOT1_6938 ( R140_U37 , U114 );
not NOT1_6939 ( R140_U38 , SI_10_ );
not NOT1_6940 ( R140_U39 , U118 );
not NOT1_6941 ( R140_U40 , SI_13_ );
not NOT1_6942 ( R140_U41 , U115 );
not NOT1_6943 ( R140_U42 , SI_12_ );
not NOT1_6944 ( R140_U43 , U116 );
not NOT1_6945 ( R140_U44 , SI_11_ );
not NOT1_6946 ( R140_U45 , U117 );
nand NAND2_6947 ( R140_U46 , U117 , SI_11_ );
not NOT1_6948 ( R140_U47 , SI_15_ );
not NOT1_6949 ( R140_U48 , U113 );
not NOT1_6950 ( R140_U49 , SI_16_ );
not NOT1_6951 ( R140_U50 , U112 );
not NOT1_6952 ( R140_U51 , SI_17_ );
not NOT1_6953 ( R140_U52 , U111 );
not NOT1_6954 ( R140_U53 , SI_18_ );
not NOT1_6955 ( R140_U54 , U110 );
not NOT1_6956 ( R140_U55 , SI_19_ );
not NOT1_6957 ( R140_U56 , U109 );
not NOT1_6958 ( R140_U57 , SI_20_ );
not NOT1_6959 ( R140_U58 , U107 );
not NOT1_6960 ( R140_U59 , SI_21_ );
not NOT1_6961 ( R140_U60 , U106 );
not NOT1_6962 ( R140_U61 , SI_22_ );
not NOT1_6963 ( R140_U62 , U105 );
not NOT1_6964 ( R140_U63 , SI_23_ );
not NOT1_6965 ( R140_U64 , U104 );
not NOT1_6966 ( R140_U65 , SI_24_ );
not NOT1_6967 ( R140_U66 , U103 );
not NOT1_6968 ( R140_U67 , SI_25_ );
not NOT1_6969 ( R140_U68 , U102 );
not NOT1_6970 ( R140_U69 , SI_26_ );
not NOT1_6971 ( R140_U70 , U101 );
not NOT1_6972 ( R140_U71 , SI_27_ );
not NOT1_6973 ( R140_U72 , U100 );
not NOT1_6974 ( R140_U73 , SI_28_ );
not NOT1_6975 ( R140_U74 , U99 );
not NOT1_6976 ( R140_U75 , SI_29_ );
not NOT1_6977 ( R140_U76 , U98 );
not NOT1_6978 ( R140_U77 , SI_30_ );
not NOT1_6979 ( R140_U78 , U96 );
nand NAND3_6980 ( R140_U79 , SI_0_ , SI_1_ , U120 );
nand NAND2_6981 ( R140_U80 , R140_U300 , R140_U217 );
nand NAND2_6982 ( R140_U81 , R140_U297 , R140_U214 );
nand NAND2_6983 ( R140_U82 , R140_U293 , R140_U206 );
nand NAND2_6984 ( R140_U83 , R140_U541 , R140_U540 );
nand NAND2_6985 ( R140_U84 , R140_U331 , R140_U330 );
nand NAND2_6986 ( R140_U85 , R140_U338 , R140_U337 );
nand NAND2_6987 ( R140_U86 , R140_U345 , R140_U344 );
nand NAND2_6988 ( R140_U87 , R140_U352 , R140_U351 );
nand NAND2_6989 ( R140_U88 , R140_U359 , R140_U358 );
nand NAND2_6990 ( R140_U89 , R140_U366 , R140_U365 );
nand NAND2_6991 ( R140_U90 , R140_U373 , R140_U372 );
nand NAND2_6992 ( R140_U91 , R140_U387 , R140_U386 );
nand NAND2_6993 ( R140_U92 , R140_U394 , R140_U393 );
nand NAND2_6994 ( R140_U93 , R140_U401 , R140_U400 );
nand NAND2_6995 ( R140_U94 , R140_U408 , R140_U407 );
nand NAND2_6996 ( R140_U95 , R140_U415 , R140_U414 );
nand NAND2_6997 ( R140_U96 , R140_U422 , R140_U421 );
nand NAND2_6998 ( R140_U97 , R140_U429 , R140_U428 );
nand NAND2_6999 ( R140_U98 , R140_U436 , R140_U435 );
nand NAND2_7000 ( R140_U99 , R140_U443 , R140_U442 );
nand NAND2_7001 ( R140_U100 , R140_U450 , R140_U449 );
nand NAND2_7002 ( R140_U101 , R140_U457 , R140_U456 );
nand NAND2_7003 ( R140_U102 , R140_U464 , R140_U463 );
nand NAND2_7004 ( R140_U103 , R140_U476 , R140_U475 );
nand NAND2_7005 ( R140_U104 , R140_U483 , R140_U482 );
nand NAND2_7006 ( R140_U105 , R140_U490 , R140_U489 );
nand NAND2_7007 ( R140_U106 , R140_U497 , R140_U496 );
nand NAND2_7008 ( R140_U107 , R140_U504 , R140_U503 );
nand NAND2_7009 ( R140_U108 , R140_U511 , R140_U510 );
nand NAND2_7010 ( R140_U109 , R140_U518 , R140_U517 );
nand NAND2_7011 ( R140_U110 , R140_U525 , R140_U524 );
nand NAND2_7012 ( R140_U111 , R140_U532 , R140_U531 );
nand NAND2_7013 ( R140_U112 , R140_U539 , R140_U538 );
and AND2_7014 ( R140_U113 , R140_U189 , R140_U193 );
and AND2_7015 ( R140_U114 , R140_U287 , R140_U194 );
and AND2_7016 ( R140_U115 , R140_U4 , R140_U199 );
and AND2_7017 ( R140_U116 , R140_U290 , R140_U200 );
and AND2_7018 ( R140_U117 , R140_U291 , R140_U204 );
and AND2_7019 ( R140_U118 , R140_U6 , R140_U207 );
and AND2_7020 ( R140_U119 , R140_U295 , R140_U208 );
and AND2_7021 ( R140_U120 , R140_U8 , R140_U219 );
and AND2_7022 ( R140_U121 , R140_U303 , R140_U220 );
and AND3_7023 ( R140_U122 , R140_U9 , R140_U282 , R140_U280 );
and AND2_7024 ( R140_U123 , R140_U283 , R140_U376 );
and AND2_7025 ( R140_U124 , R140_U141 , R140_U284 );
and AND2_7026 ( R140_U125 , R140_U326 , R140_U325 );
nand NAND2_7027 ( R140_U126 , R140_U117 , R140_U309 );
and AND2_7028 ( R140_U127 , R140_U333 , R140_U332 );
nand NAND2_7029 ( R140_U128 , R140_U307 , R140_U16 );
and AND2_7030 ( R140_U129 , R140_U340 , R140_U339 );
nand NAND2_7031 ( R140_U130 , R140_U116 , R140_U319 );
and AND2_7032 ( R140_U131 , R140_U347 , R140_U346 );
nand NAND2_7033 ( R140_U132 , R140_U289 , R140_U317 );
and AND2_7034 ( R140_U133 , R140_U354 , R140_U353 );
nand NAND2_7035 ( R140_U134 , R140_U315 , R140_U23 );
and AND2_7036 ( R140_U135 , R140_U361 , R140_U360 );
nand NAND2_7037 ( R140_U136 , R140_U114 , R140_U321 );
and AND2_7038 ( R140_U137 , R140_U368 , R140_U367 );
nand NAND2_7039 ( R140_U138 , R140_U28 , R140_U190 );
not NOT1_7040 ( R140_U139 , U95 );
not NOT1_7041 ( R140_U140 , SI_31_ );
and AND2_7042 ( R140_U141 , R140_U380 , R140_U379 );
and AND2_7043 ( R140_U142 , R140_U382 , R140_U381 );
nand NAND2_7044 ( R140_U143 , R140_U280 , R140_U279 );
nand NAND3_7045 ( R140_U144 , R140_U286 , R140_U79 , R140_U285 );
and AND2_7046 ( R140_U145 , R140_U396 , R140_U395 );
nand NAND2_7047 ( R140_U146 , R140_U276 , R140_U275 );
and AND2_7048 ( R140_U147 , R140_U403 , R140_U402 );
nand NAND2_7049 ( R140_U148 , R140_U272 , R140_U271 );
and AND2_7050 ( R140_U149 , R140_U410 , R140_U409 );
nand NAND2_7051 ( R140_U150 , R140_U268 , R140_U267 );
and AND2_7052 ( R140_U151 , R140_U417 , R140_U416 );
nand NAND2_7053 ( R140_U152 , R140_U264 , R140_U263 );
and AND2_7054 ( R140_U153 , R140_U424 , R140_U423 );
nand NAND2_7055 ( R140_U154 , R140_U260 , R140_U259 );
and AND2_7056 ( R140_U155 , R140_U431 , R140_U430 );
nand NAND2_7057 ( R140_U156 , R140_U256 , R140_U255 );
and AND2_7058 ( R140_U157 , R140_U438 , R140_U437 );
nand NAND2_7059 ( R140_U158 , R140_U252 , R140_U251 );
and AND2_7060 ( R140_U159 , R140_U445 , R140_U444 );
nand NAND2_7061 ( R140_U160 , R140_U248 , R140_U247 );
and AND2_7062 ( R140_U161 , R140_U452 , R140_U451 );
nand NAND2_7063 ( R140_U162 , R140_U244 , R140_U243 );
and AND2_7064 ( R140_U163 , R140_U459 , R140_U458 );
nand NAND2_7065 ( R140_U164 , R140_U240 , R140_U239 );
nand NAND2_7066 ( R140_U165 , U120 , SI_0_ );
and AND2_7067 ( R140_U166 , R140_U471 , R140_U470 );
nand NAND2_7068 ( R140_U167 , R140_U236 , R140_U235 );
and AND2_7069 ( R140_U168 , R140_U478 , R140_U477 );
nand NAND2_7070 ( R140_U169 , R140_U232 , R140_U231 );
and AND2_7071 ( R140_U170 , R140_U485 , R140_U484 );
nand NAND2_7072 ( R140_U171 , R140_U228 , R140_U227 );
and AND2_7073 ( R140_U172 , R140_U492 , R140_U491 );
nand NAND2_7074 ( R140_U173 , R140_U224 , R140_U223 );
and AND2_7075 ( R140_U174 , R140_U499 , R140_U498 );
nand NAND2_7076 ( R140_U175 , R140_U121 , R140_U302 );
and AND2_7077 ( R140_U176 , R140_U506 , R140_U505 );
nand NAND2_7078 ( R140_U177 , R140_U301 , R140_U299 );
and AND2_7079 ( R140_U178 , R140_U513 , R140_U512 );
nand NAND2_7080 ( R140_U179 , R140_U298 , R140_U296 );
and AND2_7081 ( R140_U180 , R140_U520 , R140_U519 );
nand NAND2_7082 ( R140_U181 , R140_U46 , R140_U210 );
and AND2_7083 ( R140_U182 , R140_U527 , R140_U526 );
nand NAND2_7084 ( R140_U183 , R140_U119 , R140_U313 );
and AND2_7085 ( R140_U184 , R140_U534 , R140_U533 );
nand NAND2_7086 ( R140_U185 , R140_U294 , R140_U311 );
not NOT1_7087 ( R140_U186 , R140_U79 );
not NOT1_7088 ( R140_U187 , R140_U165 );
not NOT1_7089 ( R140_U188 , R140_U144 );
or OR2_7090 ( R140_U189 , SI_2_ , U108 );
nand NAND2_7091 ( R140_U190 , R140_U304 , R140_U189 );
not NOT1_7092 ( R140_U191 , R140_U28 );
not NOT1_7093 ( R140_U192 , R140_U138 );
or OR2_7094 ( R140_U193 , SI_3_ , U97 );
nand NAND2_7095 ( R140_U194 , U97 , SI_3_ );
or OR2_7096 ( R140_U195 , SI_4_ , U94 );
not NOT1_7097 ( R140_U196 , R140_U23 );
or OR2_7098 ( R140_U197 , SI_5_ , U93 );
nand NAND2_7099 ( R140_U198 , U93 , SI_5_ );
or OR2_7100 ( R140_U199 , SI_6_ , U92 );
nand NAND2_7101 ( R140_U200 , U92 , SI_6_ );
or OR2_7102 ( R140_U201 , SI_7_ , U91 );
not NOT1_7103 ( R140_U202 , R140_U16 );
or OR2_7104 ( R140_U203 , SI_8_ , U90 );
nand NAND2_7105 ( R140_U204 , U90 , SI_8_ );
or OR2_7106 ( R140_U205 , SI_9_ , U89 );
nand NAND2_7107 ( R140_U206 , SI_9_ , U89 );
or OR2_7108 ( R140_U207 , SI_10_ , U118 );
nand NAND2_7109 ( R140_U208 , U118 , SI_10_ );
or OR2_7110 ( R140_U209 , SI_11_ , U117 );
nand NAND2_7111 ( R140_U210 , R140_U209 , R140_U183 );
not NOT1_7112 ( R140_U211 , R140_U46 );
not NOT1_7113 ( R140_U212 , R140_U181 );
or OR2_7114 ( R140_U213 , SI_12_ , U116 );
nand NAND2_7115 ( R140_U214 , U116 , SI_12_ );
not NOT1_7116 ( R140_U215 , R140_U179 );
or OR2_7117 ( R140_U216 , SI_13_ , U115 );
nand NAND2_7118 ( R140_U217 , U115 , SI_13_ );
not NOT1_7119 ( R140_U218 , R140_U177 );
or OR2_7120 ( R140_U219 , SI_14_ , U114 );
nand NAND2_7121 ( R140_U220 , U114 , SI_14_ );
not NOT1_7122 ( R140_U221 , R140_U175 );
or OR2_7123 ( R140_U222 , SI_15_ , U113 );
nand NAND2_7124 ( R140_U223 , R140_U222 , R140_U175 );
nand NAND2_7125 ( R140_U224 , U113 , SI_15_ );
not NOT1_7126 ( R140_U225 , R140_U173 );
or OR2_7127 ( R140_U226 , SI_16_ , U112 );
nand NAND2_7128 ( R140_U227 , R140_U226 , R140_U173 );
nand NAND2_7129 ( R140_U228 , U112 , SI_16_ );
not NOT1_7130 ( R140_U229 , R140_U171 );
or OR2_7131 ( R140_U230 , SI_17_ , U111 );
nand NAND2_7132 ( R140_U231 , R140_U230 , R140_U171 );
nand NAND2_7133 ( R140_U232 , U111 , SI_17_ );
not NOT1_7134 ( R140_U233 , R140_U169 );
or OR2_7135 ( R140_U234 , SI_18_ , U110 );
nand NAND2_7136 ( R140_U235 , R140_U234 , R140_U169 );
nand NAND2_7137 ( R140_U236 , U110 , SI_18_ );
not NOT1_7138 ( R140_U237 , R140_U167 );
or OR2_7139 ( R140_U238 , SI_19_ , U109 );
nand NAND2_7140 ( R140_U239 , R140_U238 , R140_U167 );
nand NAND2_7141 ( R140_U240 , U109 , SI_19_ );
not NOT1_7142 ( R140_U241 , R140_U164 );
or OR2_7143 ( R140_U242 , SI_20_ , U107 );
nand NAND2_7144 ( R140_U243 , R140_U242 , R140_U164 );
nand NAND2_7145 ( R140_U244 , U107 , SI_20_ );
not NOT1_7146 ( R140_U245 , R140_U162 );
or OR2_7147 ( R140_U246 , SI_21_ , U106 );
nand NAND2_7148 ( R140_U247 , R140_U246 , R140_U162 );
nand NAND2_7149 ( R140_U248 , U106 , SI_21_ );
not NOT1_7150 ( R140_U249 , R140_U160 );
or OR2_7151 ( R140_U250 , SI_22_ , U105 );
nand NAND2_7152 ( R140_U251 , R140_U250 , R140_U160 );
nand NAND2_7153 ( R140_U252 , U105 , SI_22_ );
not NOT1_7154 ( R140_U253 , R140_U158 );
or OR2_7155 ( R140_U254 , SI_23_ , U104 );
nand NAND2_7156 ( R140_U255 , R140_U254 , R140_U158 );
nand NAND2_7157 ( R140_U256 , U104 , SI_23_ );
not NOT1_7158 ( R140_U257 , R140_U156 );
or OR2_7159 ( R140_U258 , SI_24_ , U103 );
nand NAND2_7160 ( R140_U259 , R140_U258 , R140_U156 );
nand NAND2_7161 ( R140_U260 , U103 , SI_24_ );
not NOT1_7162 ( R140_U261 , R140_U154 );
or OR2_7163 ( R140_U262 , SI_25_ , U102 );
nand NAND2_7164 ( R140_U263 , R140_U262 , R140_U154 );
nand NAND2_7165 ( R140_U264 , U102 , SI_25_ );
not NOT1_7166 ( R140_U265 , R140_U152 );
or OR2_7167 ( R140_U266 , SI_26_ , U101 );
nand NAND2_7168 ( R140_U267 , R140_U266 , R140_U152 );
nand NAND2_7169 ( R140_U268 , U101 , SI_26_ );
not NOT1_7170 ( R140_U269 , R140_U150 );
or OR2_7171 ( R140_U270 , SI_27_ , U100 );
nand NAND2_7172 ( R140_U271 , R140_U270 , R140_U150 );
nand NAND2_7173 ( R140_U272 , U100 , SI_27_ );
not NOT1_7174 ( R140_U273 , R140_U148 );
or OR2_7175 ( R140_U274 , SI_28_ , U99 );
nand NAND2_7176 ( R140_U275 , R140_U274 , R140_U148 );
nand NAND2_7177 ( R140_U276 , U99 , SI_28_ );
not NOT1_7178 ( R140_U277 , R140_U146 );
or OR2_7179 ( R140_U278 , SI_29_ , U98 );
nand NAND2_7180 ( R140_U279 , R140_U278 , R140_U146 );
nand NAND2_7181 ( R140_U280 , U98 , SI_29_ );
not NOT1_7182 ( R140_U281 , R140_U143 );
nand NAND2_7183 ( R140_U282 , U96 , SI_30_ );
or OR2_7184 ( R140_U283 , U96 , SI_30_ );
nand NAND2_7185 ( R140_U284 , R140_U279 , R140_U122 );
nand NAND3_7186 ( R140_U285 , U120 , SI_0_ , U119 );
nand NAND2_7187 ( R140_U286 , U119 , SI_1_ );
nand NAND2_7188 ( R140_U287 , R140_U191 , R140_U193 );
nand NAND2_7189 ( R140_U288 , R140_U196 , R140_U197 );
not NOT1_7190 ( R140_U289 , R140_U35 );
nand NAND2_7191 ( R140_U290 , R140_U35 , R140_U199 );
nand NAND2_7192 ( R140_U291 , R140_U202 , R140_U203 );
nand NAND2_7193 ( R140_U292 , R140_U291 , R140_U204 );
nand NAND2_7194 ( R140_U293 , R140_U292 , R140_U205 );
not NOT1_7195 ( R140_U294 , R140_U82 );
nand NAND2_7196 ( R140_U295 , R140_U82 , R140_U207 );
nand NAND2_7197 ( R140_U296 , R140_U7 , R140_U183 );
nand NAND2_7198 ( R140_U297 , R140_U211 , R140_U213 );
not NOT1_7199 ( R140_U298 , R140_U81 );
nand NAND2_7200 ( R140_U299 , R140_U8 , R140_U183 );
nand NAND2_7201 ( R140_U300 , R140_U81 , R140_U216 );
not NOT1_7202 ( R140_U301 , R140_U80 );
nand NAND2_7203 ( R140_U302 , R140_U120 , R140_U183 );
nand NAND2_7204 ( R140_U303 , R140_U80 , R140_U219 );
nand NAND3_7205 ( R140_U304 , R140_U306 , R140_U286 , R140_U305 );
nand NAND3_7206 ( R140_U305 , U120 , SI_0_ , U119 );
nand NAND3_7207 ( R140_U306 , SI_0_ , SI_1_ , U120 );
nand NAND2_7208 ( R140_U307 , R140_U201 , R140_U130 );
not NOT1_7209 ( R140_U308 , R140_U128 );
nand NAND2_7210 ( R140_U309 , R140_U5 , R140_U130 );
not NOT1_7211 ( R140_U310 , R140_U126 );
nand NAND2_7212 ( R140_U311 , R140_U6 , R140_U130 );
not NOT1_7213 ( R140_U312 , R140_U185 );
nand NAND2_7214 ( R140_U313 , R140_U118 , R140_U130 );
not NOT1_7215 ( R140_U314 , R140_U183 );
nand NAND2_7216 ( R140_U315 , R140_U195 , R140_U136 );
not NOT1_7217 ( R140_U316 , R140_U134 );
nand NAND2_7218 ( R140_U317 , R140_U4 , R140_U136 );
not NOT1_7219 ( R140_U318 , R140_U132 );
nand NAND2_7220 ( R140_U319 , R140_U115 , R140_U136 );
not NOT1_7221 ( R140_U320 , R140_U130 );
nand NAND2_7222 ( R140_U321 , R140_U113 , R140_U144 );
not NOT1_7223 ( R140_U322 , R140_U136 );
nand NAND2_7224 ( R140_U323 , R140_U123 , R140_U143 );
nand NAND2_7225 ( R140_U324 , R140_U186 , U119 );
nand NAND2_7226 ( R140_U325 , U89 , R140_U34 );
nand NAND2_7227 ( R140_U326 , SI_9_ , R140_U33 );
nand NAND2_7228 ( R140_U327 , U89 , R140_U34 );
nand NAND2_7229 ( R140_U328 , SI_9_ , R140_U33 );
nand NAND2_7230 ( R140_U329 , R140_U328 , R140_U327 );
nand NAND2_7231 ( R140_U330 , R140_U125 , R140_U126 );
nand NAND2_7232 ( R140_U331 , R140_U310 , R140_U329 );
nand NAND2_7233 ( R140_U332 , U90 , R140_U12 );
nand NAND2_7234 ( R140_U333 , SI_8_ , R140_U13 );
nand NAND2_7235 ( R140_U334 , U90 , R140_U12 );
nand NAND2_7236 ( R140_U335 , SI_8_ , R140_U13 );
nand NAND2_7237 ( R140_U336 , R140_U335 , R140_U334 );
nand NAND2_7238 ( R140_U337 , R140_U127 , R140_U128 );
nand NAND2_7239 ( R140_U338 , R140_U308 , R140_U336 );
nand NAND2_7240 ( R140_U339 , U91 , R140_U14 );
nand NAND2_7241 ( R140_U340 , SI_7_ , R140_U15 );
nand NAND2_7242 ( R140_U341 , U91 , R140_U14 );
nand NAND2_7243 ( R140_U342 , SI_7_ , R140_U15 );
nand NAND2_7244 ( R140_U343 , R140_U342 , R140_U341 );
nand NAND2_7245 ( R140_U344 , R140_U129 , R140_U130 );
nand NAND2_7246 ( R140_U345 , R140_U320 , R140_U343 );
nand NAND2_7247 ( R140_U346 , U92 , R140_U17 );
nand NAND2_7248 ( R140_U347 , SI_6_ , R140_U18 );
nand NAND2_7249 ( R140_U348 , U92 , R140_U17 );
nand NAND2_7250 ( R140_U349 , SI_6_ , R140_U18 );
nand NAND2_7251 ( R140_U350 , R140_U349 , R140_U348 );
nand NAND2_7252 ( R140_U351 , R140_U131 , R140_U132 );
nand NAND2_7253 ( R140_U352 , R140_U318 , R140_U350 );
nand NAND2_7254 ( R140_U353 , U93 , R140_U19 );
nand NAND2_7255 ( R140_U354 , SI_5_ , R140_U20 );
nand NAND2_7256 ( R140_U355 , U93 , R140_U19 );
nand NAND2_7257 ( R140_U356 , SI_5_ , R140_U20 );
nand NAND2_7258 ( R140_U357 , R140_U356 , R140_U355 );
nand NAND2_7259 ( R140_U358 , R140_U133 , R140_U134 );
nand NAND2_7260 ( R140_U359 , R140_U316 , R140_U357 );
nand NAND2_7261 ( R140_U360 , U94 , R140_U21 );
nand NAND2_7262 ( R140_U361 , SI_4_ , R140_U22 );
nand NAND2_7263 ( R140_U362 , U94 , R140_U21 );
nand NAND2_7264 ( R140_U363 , SI_4_ , R140_U22 );
nand NAND2_7265 ( R140_U364 , R140_U363 , R140_U362 );
nand NAND2_7266 ( R140_U365 , R140_U135 , R140_U136 );
nand NAND2_7267 ( R140_U366 , R140_U322 , R140_U364 );
nand NAND2_7268 ( R140_U367 , U97 , R140_U24 );
nand NAND2_7269 ( R140_U368 , SI_3_ , R140_U25 );
nand NAND2_7270 ( R140_U369 , U97 , R140_U24 );
nand NAND2_7271 ( R140_U370 , SI_3_ , R140_U25 );
nand NAND2_7272 ( R140_U371 , R140_U370 , R140_U369 );
nand NAND2_7273 ( R140_U372 , R140_U137 , R140_U138 );
nand NAND2_7274 ( R140_U373 , R140_U192 , R140_U371 );
nand NAND2_7275 ( R140_U374 , U95 , R140_U140 );
nand NAND2_7276 ( R140_U375 , SI_31_ , R140_U139 );
nand NAND2_7277 ( R140_U376 , R140_U375 , R140_U374 );
nand NAND2_7278 ( R140_U377 , U95 , R140_U140 );
nand NAND2_7279 ( R140_U378 , SI_31_ , R140_U139 );
nand NAND3_7280 ( R140_U379 , R140_U9 , R140_U77 , R140_U78 );
nand NAND3_7281 ( R140_U380 , SI_30_ , R140_U376 , U96 );
nand NAND2_7282 ( R140_U381 , U96 , R140_U77 );
nand NAND2_7283 ( R140_U382 , SI_30_ , R140_U78 );
nand NAND2_7284 ( R140_U383 , U96 , R140_U77 );
nand NAND2_7285 ( R140_U384 , SI_30_ , R140_U78 );
nand NAND2_7286 ( R140_U385 , R140_U384 , R140_U383 );
nand NAND2_7287 ( R140_U386 , R140_U142 , R140_U143 );
nand NAND2_7288 ( R140_U387 , R140_U281 , R140_U385 );
nand NAND2_7289 ( R140_U388 , U108 , R140_U26 );
nand NAND2_7290 ( R140_U389 , SI_2_ , R140_U27 );
nand NAND2_7291 ( R140_U390 , U108 , R140_U26 );
nand NAND2_7292 ( R140_U391 , SI_2_ , R140_U27 );
nand NAND2_7293 ( R140_U392 , R140_U391 , R140_U390 );
nand NAND3_7294 ( R140_U393 , R140_U389 , R140_U388 , R140_U144 );
nand NAND2_7295 ( R140_U394 , R140_U188 , R140_U392 );
nand NAND2_7296 ( R140_U395 , U98 , R140_U75 );
nand NAND2_7297 ( R140_U396 , SI_29_ , R140_U76 );
nand NAND2_7298 ( R140_U397 , U98 , R140_U75 );
nand NAND2_7299 ( R140_U398 , SI_29_ , R140_U76 );
nand NAND2_7300 ( R140_U399 , R140_U398 , R140_U397 );
nand NAND2_7301 ( R140_U400 , R140_U145 , R140_U146 );
nand NAND2_7302 ( R140_U401 , R140_U277 , R140_U399 );
nand NAND2_7303 ( R140_U402 , U99 , R140_U73 );
nand NAND2_7304 ( R140_U403 , SI_28_ , R140_U74 );
nand NAND2_7305 ( R140_U404 , U99 , R140_U73 );
nand NAND2_7306 ( R140_U405 , SI_28_ , R140_U74 );
nand NAND2_7307 ( R140_U406 , R140_U405 , R140_U404 );
nand NAND2_7308 ( R140_U407 , R140_U147 , R140_U148 );
nand NAND2_7309 ( R140_U408 , R140_U273 , R140_U406 );
nand NAND2_7310 ( R140_U409 , U100 , R140_U71 );
nand NAND2_7311 ( R140_U410 , SI_27_ , R140_U72 );
nand NAND2_7312 ( R140_U411 , U100 , R140_U71 );
nand NAND2_7313 ( R140_U412 , SI_27_ , R140_U72 );
nand NAND2_7314 ( R140_U413 , R140_U412 , R140_U411 );
nand NAND2_7315 ( R140_U414 , R140_U149 , R140_U150 );
nand NAND2_7316 ( R140_U415 , R140_U269 , R140_U413 );
nand NAND2_7317 ( R140_U416 , U101 , R140_U69 );
nand NAND2_7318 ( R140_U417 , SI_26_ , R140_U70 );
nand NAND2_7319 ( R140_U418 , U101 , R140_U69 );
nand NAND2_7320 ( R140_U419 , SI_26_ , R140_U70 );
nand NAND2_7321 ( R140_U420 , R140_U419 , R140_U418 );
nand NAND2_7322 ( R140_U421 , R140_U151 , R140_U152 );
nand NAND2_7323 ( R140_U422 , R140_U265 , R140_U420 );
nand NAND2_7324 ( R140_U423 , U102 , R140_U67 );
nand NAND2_7325 ( R140_U424 , SI_25_ , R140_U68 );
nand NAND2_7326 ( R140_U425 , U102 , R140_U67 );
nand NAND2_7327 ( R140_U426 , SI_25_ , R140_U68 );
nand NAND2_7328 ( R140_U427 , R140_U426 , R140_U425 );
nand NAND2_7329 ( R140_U428 , R140_U153 , R140_U154 );
nand NAND2_7330 ( R140_U429 , R140_U261 , R140_U427 );
nand NAND2_7331 ( R140_U430 , U103 , R140_U65 );
nand NAND2_7332 ( R140_U431 , SI_24_ , R140_U66 );
nand NAND2_7333 ( R140_U432 , U103 , R140_U65 );
nand NAND2_7334 ( R140_U433 , SI_24_ , R140_U66 );
nand NAND2_7335 ( R140_U434 , R140_U433 , R140_U432 );
nand NAND2_7336 ( R140_U435 , R140_U155 , R140_U156 );
nand NAND2_7337 ( R140_U436 , R140_U257 , R140_U434 );
nand NAND2_7338 ( R140_U437 , U104 , R140_U63 );
nand NAND2_7339 ( R140_U438 , SI_23_ , R140_U64 );
nand NAND2_7340 ( R140_U439 , U104 , R140_U63 );
nand NAND2_7341 ( R140_U440 , SI_23_ , R140_U64 );
nand NAND2_7342 ( R140_U441 , R140_U440 , R140_U439 );
nand NAND2_7343 ( R140_U442 , R140_U157 , R140_U158 );
nand NAND2_7344 ( R140_U443 , R140_U253 , R140_U441 );
nand NAND2_7345 ( R140_U444 , U105 , R140_U61 );
nand NAND2_7346 ( R140_U445 , SI_22_ , R140_U62 );
nand NAND2_7347 ( R140_U446 , U105 , R140_U61 );
nand NAND2_7348 ( R140_U447 , SI_22_ , R140_U62 );
nand NAND2_7349 ( R140_U448 , R140_U447 , R140_U446 );
nand NAND2_7350 ( R140_U449 , R140_U159 , R140_U160 );
nand NAND2_7351 ( R140_U450 , R140_U249 , R140_U448 );
nand NAND2_7352 ( R140_U451 , U106 , R140_U59 );
nand NAND2_7353 ( R140_U452 , SI_21_ , R140_U60 );
nand NAND2_7354 ( R140_U453 , U106 , R140_U59 );
nand NAND2_7355 ( R140_U454 , SI_21_ , R140_U60 );
nand NAND2_7356 ( R140_U455 , R140_U454 , R140_U453 );
nand NAND2_7357 ( R140_U456 , R140_U161 , R140_U162 );
nand NAND2_7358 ( R140_U457 , R140_U245 , R140_U455 );
nand NAND2_7359 ( R140_U458 , U107 , R140_U57 );
nand NAND2_7360 ( R140_U459 , SI_20_ , R140_U58 );
nand NAND2_7361 ( R140_U460 , U107 , R140_U57 );
nand NAND2_7362 ( R140_U461 , SI_20_ , R140_U58 );
nand NAND2_7363 ( R140_U462 , R140_U461 , R140_U460 );
nand NAND2_7364 ( R140_U463 , R140_U163 , R140_U164 );
nand NAND2_7365 ( R140_U464 , R140_U241 , R140_U462 );
nand NAND2_7366 ( R140_U465 , U119 , R140_U165 );
nand NAND2_7367 ( R140_U466 , R140_U187 , R140_U32 );
nand NAND2_7368 ( R140_U467 , R140_U466 , R140_U465 );
nand NAND3_7369 ( R140_U468 , R140_U165 , R140_U32 , SI_1_ );
nand NAND2_7370 ( R140_U469 , R140_U467 , R140_U29 );
nand NAND2_7371 ( R140_U470 , U109 , R140_U55 );
nand NAND2_7372 ( R140_U471 , SI_19_ , R140_U56 );
nand NAND2_7373 ( R140_U472 , U109 , R140_U55 );
nand NAND2_7374 ( R140_U473 , SI_19_ , R140_U56 );
nand NAND2_7375 ( R140_U474 , R140_U473 , R140_U472 );
nand NAND2_7376 ( R140_U475 , R140_U166 , R140_U167 );
nand NAND2_7377 ( R140_U476 , R140_U237 , R140_U474 );
nand NAND2_7378 ( R140_U477 , U110 , R140_U53 );
nand NAND2_7379 ( R140_U478 , SI_18_ , R140_U54 );
nand NAND2_7380 ( R140_U479 , U110 , R140_U53 );
nand NAND2_7381 ( R140_U480 , SI_18_ , R140_U54 );
nand NAND2_7382 ( R140_U481 , R140_U480 , R140_U479 );
nand NAND2_7383 ( R140_U482 , R140_U168 , R140_U169 );
nand NAND2_7384 ( R140_U483 , R140_U233 , R140_U481 );
nand NAND2_7385 ( R140_U484 , U111 , R140_U51 );
nand NAND2_7386 ( R140_U485 , SI_17_ , R140_U52 );
nand NAND2_7387 ( R140_U486 , U111 , R140_U51 );
nand NAND2_7388 ( R140_U487 , SI_17_ , R140_U52 );
nand NAND2_7389 ( R140_U488 , R140_U487 , R140_U486 );
nand NAND2_7390 ( R140_U489 , R140_U170 , R140_U171 );
nand NAND2_7391 ( R140_U490 , R140_U229 , R140_U488 );
nand NAND2_7392 ( R140_U491 , U112 , R140_U49 );
nand NAND2_7393 ( R140_U492 , SI_16_ , R140_U50 );
nand NAND2_7394 ( R140_U493 , U112 , R140_U49 );
nand NAND2_7395 ( R140_U494 , SI_16_ , R140_U50 );
nand NAND2_7396 ( R140_U495 , R140_U494 , R140_U493 );
nand NAND2_7397 ( R140_U496 , R140_U172 , R140_U173 );
nand NAND2_7398 ( R140_U497 , R140_U225 , R140_U495 );
nand NAND2_7399 ( R140_U498 , U113 , R140_U47 );
nand NAND2_7400 ( R140_U499 , SI_15_ , R140_U48 );
nand NAND2_7401 ( R140_U500 , U113 , R140_U47 );
nand NAND2_7402 ( R140_U501 , SI_15_ , R140_U48 );
nand NAND2_7403 ( R140_U502 , R140_U501 , R140_U500 );
nand NAND2_7404 ( R140_U503 , R140_U174 , R140_U175 );
nand NAND2_7405 ( R140_U504 , R140_U221 , R140_U502 );
nand NAND2_7406 ( R140_U505 , U114 , R140_U36 );
nand NAND2_7407 ( R140_U506 , SI_14_ , R140_U37 );
nand NAND2_7408 ( R140_U507 , U114 , R140_U36 );
nand NAND2_7409 ( R140_U508 , SI_14_ , R140_U37 );
nand NAND2_7410 ( R140_U509 , R140_U508 , R140_U507 );
nand NAND2_7411 ( R140_U510 , R140_U176 , R140_U177 );
nand NAND2_7412 ( R140_U511 , R140_U218 , R140_U509 );
nand NAND2_7413 ( R140_U512 , U115 , R140_U40 );
nand NAND2_7414 ( R140_U513 , SI_13_ , R140_U41 );
nand NAND2_7415 ( R140_U514 , U115 , R140_U40 );
nand NAND2_7416 ( R140_U515 , SI_13_ , R140_U41 );
nand NAND2_7417 ( R140_U516 , R140_U515 , R140_U514 );
nand NAND2_7418 ( R140_U517 , R140_U178 , R140_U179 );
nand NAND2_7419 ( R140_U518 , R140_U215 , R140_U516 );
nand NAND2_7420 ( R140_U519 , U116 , R140_U42 );
nand NAND2_7421 ( R140_U520 , SI_12_ , R140_U43 );
nand NAND2_7422 ( R140_U521 , U116 , R140_U42 );
nand NAND2_7423 ( R140_U522 , SI_12_ , R140_U43 );
nand NAND2_7424 ( R140_U523 , R140_U522 , R140_U521 );
nand NAND2_7425 ( R140_U524 , R140_U180 , R140_U181 );
nand NAND2_7426 ( R140_U525 , R140_U212 , R140_U523 );
nand NAND2_7427 ( R140_U526 , U117 , R140_U44 );
nand NAND2_7428 ( R140_U527 , SI_11_ , R140_U45 );
nand NAND2_7429 ( R140_U528 , U117 , R140_U44 );
nand NAND2_7430 ( R140_U529 , SI_11_ , R140_U45 );
nand NAND2_7431 ( R140_U530 , R140_U529 , R140_U528 );
nand NAND2_7432 ( R140_U531 , R140_U182 , R140_U183 );
nand NAND2_7433 ( R140_U532 , R140_U314 , R140_U530 );
nand NAND2_7434 ( R140_U533 , U118 , R140_U38 );
nand NAND2_7435 ( R140_U534 , SI_10_ , R140_U39 );
nand NAND2_7436 ( R140_U535 , U118 , R140_U38 );
nand NAND2_7437 ( R140_U536 , SI_10_ , R140_U39 );
nand NAND2_7438 ( R140_U537 , R140_U536 , R140_U535 );
nand NAND2_7439 ( R140_U538 , R140_U184 , R140_U185 );
nand NAND2_7440 ( R140_U539 , R140_U312 , R140_U537 );
nand NAND2_7441 ( R140_U540 , U120 , R140_U30 );
nand NAND2_7442 ( R140_U541 , SI_0_ , R140_U31 );
not NOT1_7443 ( LT_1075_19_U6 , P2_ADDR_REG_19_ );
not NOT1_7444 ( P1_ADD_95_U4 , P1_REG3_REG_3_ );
and AND3_7445 ( P1_ADD_95_U5 , P1_REG3_REG_28_ , P1_REG3_REG_27_ , P1_ADD_95_U102 );
not NOT1_7446 ( P1_ADD_95_U6 , P1_REG3_REG_4_ );
nand NAND2_7447 ( P1_ADD_95_U7 , P1_REG3_REG_4_ , P1_REG3_REG_3_ );
not NOT1_7448 ( P1_ADD_95_U8 , P1_REG3_REG_5_ );
nand NAND2_7449 ( P1_ADD_95_U9 , P1_REG3_REG_5_ , P1_ADD_95_U80 );
not NOT1_7450 ( P1_ADD_95_U10 , P1_REG3_REG_6_ );
nand NAND2_7451 ( P1_ADD_95_U11 , P1_REG3_REG_6_ , P1_ADD_95_U81 );
not NOT1_7452 ( P1_ADD_95_U12 , P1_REG3_REG_7_ );
nand NAND2_7453 ( P1_ADD_95_U13 , P1_REG3_REG_7_ , P1_ADD_95_U82 );
not NOT1_7454 ( P1_ADD_95_U14 , P1_REG3_REG_8_ );
not NOT1_7455 ( P1_ADD_95_U15 , P1_REG3_REG_9_ );
nand NAND2_7456 ( P1_ADD_95_U16 , P1_REG3_REG_8_ , P1_ADD_95_U83 );
nand NAND2_7457 ( P1_ADD_95_U17 , P1_ADD_95_U84 , P1_REG3_REG_9_ );
not NOT1_7458 ( P1_ADD_95_U18 , P1_REG3_REG_10_ );
nand NAND2_7459 ( P1_ADD_95_U19 , P1_REG3_REG_10_ , P1_ADD_95_U85 );
not NOT1_7460 ( P1_ADD_95_U20 , P1_REG3_REG_11_ );
nand NAND2_7461 ( P1_ADD_95_U21 , P1_REG3_REG_11_ , P1_ADD_95_U86 );
not NOT1_7462 ( P1_ADD_95_U22 , P1_REG3_REG_12_ );
nand NAND2_7463 ( P1_ADD_95_U23 , P1_REG3_REG_12_ , P1_ADD_95_U87 );
not NOT1_7464 ( P1_ADD_95_U24 , P1_REG3_REG_13_ );
nand NAND2_7465 ( P1_ADD_95_U25 , P1_REG3_REG_13_ , P1_ADD_95_U88 );
not NOT1_7466 ( P1_ADD_95_U26 , P1_REG3_REG_14_ );
nand NAND2_7467 ( P1_ADD_95_U27 , P1_REG3_REG_14_ , P1_ADD_95_U89 );
not NOT1_7468 ( P1_ADD_95_U28 , P1_REG3_REG_15_ );
nand NAND2_7469 ( P1_ADD_95_U29 , P1_REG3_REG_15_ , P1_ADD_95_U90 );
not NOT1_7470 ( P1_ADD_95_U30 , P1_REG3_REG_16_ );
nand NAND2_7471 ( P1_ADD_95_U31 , P1_REG3_REG_16_ , P1_ADD_95_U91 );
not NOT1_7472 ( P1_ADD_95_U32 , P1_REG3_REG_17_ );
nand NAND2_7473 ( P1_ADD_95_U33 , P1_REG3_REG_17_ , P1_ADD_95_U92 );
not NOT1_7474 ( P1_ADD_95_U34 , P1_REG3_REG_18_ );
nand NAND2_7475 ( P1_ADD_95_U35 , P1_REG3_REG_18_ , P1_ADD_95_U93 );
not NOT1_7476 ( P1_ADD_95_U36 , P1_REG3_REG_19_ );
nand NAND2_7477 ( P1_ADD_95_U37 , P1_REG3_REG_19_ , P1_ADD_95_U94 );
not NOT1_7478 ( P1_ADD_95_U38 , P1_REG3_REG_20_ );
nand NAND2_7479 ( P1_ADD_95_U39 , P1_REG3_REG_20_ , P1_ADD_95_U95 );
not NOT1_7480 ( P1_ADD_95_U40 , P1_REG3_REG_21_ );
nand NAND2_7481 ( P1_ADD_95_U41 , P1_REG3_REG_21_ , P1_ADD_95_U96 );
not NOT1_7482 ( P1_ADD_95_U42 , P1_REG3_REG_22_ );
nand NAND2_7483 ( P1_ADD_95_U43 , P1_REG3_REG_22_ , P1_ADD_95_U97 );
not NOT1_7484 ( P1_ADD_95_U44 , P1_REG3_REG_23_ );
nand NAND2_7485 ( P1_ADD_95_U45 , P1_REG3_REG_23_ , P1_ADD_95_U98 );
not NOT1_7486 ( P1_ADD_95_U46 , P1_REG3_REG_24_ );
nand NAND2_7487 ( P1_ADD_95_U47 , P1_REG3_REG_24_ , P1_ADD_95_U99 );
not NOT1_7488 ( P1_ADD_95_U48 , P1_REG3_REG_25_ );
nand NAND2_7489 ( P1_ADD_95_U49 , P1_REG3_REG_25_ , P1_ADD_95_U100 );
not NOT1_7490 ( P1_ADD_95_U50 , P1_REG3_REG_26_ );
nand NAND2_7491 ( P1_ADD_95_U51 , P1_REG3_REG_26_ , P1_ADD_95_U101 );
not NOT1_7492 ( P1_ADD_95_U52 , P1_REG3_REG_28_ );
not NOT1_7493 ( P1_ADD_95_U53 , P1_REG3_REG_27_ );
nand NAND2_7494 ( P1_ADD_95_U54 , P1_ADD_95_U105 , P1_ADD_95_U104 );
nand NAND2_7495 ( P1_ADD_95_U55 , P1_ADD_95_U107 , P1_ADD_95_U106 );
nand NAND2_7496 ( P1_ADD_95_U56 , P1_ADD_95_U109 , P1_ADD_95_U108 );
nand NAND2_7497 ( P1_ADD_95_U57 , P1_ADD_95_U111 , P1_ADD_95_U110 );
nand NAND2_7498 ( P1_ADD_95_U58 , P1_ADD_95_U113 , P1_ADD_95_U112 );
nand NAND2_7499 ( P1_ADD_95_U59 , P1_ADD_95_U115 , P1_ADD_95_U114 );
nand NAND2_7500 ( P1_ADD_95_U60 , P1_ADD_95_U117 , P1_ADD_95_U116 );
nand NAND2_7501 ( P1_ADD_95_U61 , P1_ADD_95_U119 , P1_ADD_95_U118 );
nand NAND2_7502 ( P1_ADD_95_U62 , P1_ADD_95_U121 , P1_ADD_95_U120 );
nand NAND2_7503 ( P1_ADD_95_U63 , P1_ADD_95_U123 , P1_ADD_95_U122 );
nand NAND2_7504 ( P1_ADD_95_U64 , P1_ADD_95_U125 , P1_ADD_95_U124 );
nand NAND2_7505 ( P1_ADD_95_U65 , P1_ADD_95_U127 , P1_ADD_95_U126 );
nand NAND2_7506 ( P1_ADD_95_U66 , P1_ADD_95_U129 , P1_ADD_95_U128 );
nand NAND2_7507 ( P1_ADD_95_U67 , P1_ADD_95_U131 , P1_ADD_95_U130 );
nand NAND2_7508 ( P1_ADD_95_U68 , P1_ADD_95_U133 , P1_ADD_95_U132 );
nand NAND2_7509 ( P1_ADD_95_U69 , P1_ADD_95_U135 , P1_ADD_95_U134 );
nand NAND2_7510 ( P1_ADD_95_U70 , P1_ADD_95_U137 , P1_ADD_95_U136 );
nand NAND2_7511 ( P1_ADD_95_U71 , P1_ADD_95_U139 , P1_ADD_95_U138 );
nand NAND2_7512 ( P1_ADD_95_U72 , P1_ADD_95_U141 , P1_ADD_95_U140 );
nand NAND2_7513 ( P1_ADD_95_U73 , P1_ADD_95_U143 , P1_ADD_95_U142 );
nand NAND2_7514 ( P1_ADD_95_U74 , P1_ADD_95_U145 , P1_ADD_95_U144 );
nand NAND2_7515 ( P1_ADD_95_U75 , P1_ADD_95_U147 , P1_ADD_95_U146 );
nand NAND2_7516 ( P1_ADD_95_U76 , P1_ADD_95_U149 , P1_ADD_95_U148 );
nand NAND2_7517 ( P1_ADD_95_U77 , P1_ADD_95_U151 , P1_ADD_95_U150 );
nand NAND2_7518 ( P1_ADD_95_U78 , P1_ADD_95_U153 , P1_ADD_95_U152 );
nand NAND2_7519 ( P1_ADD_95_U79 , P1_REG3_REG_27_ , P1_ADD_95_U102 );
not NOT1_7520 ( P1_ADD_95_U80 , P1_ADD_95_U7 );
not NOT1_7521 ( P1_ADD_95_U81 , P1_ADD_95_U9 );
not NOT1_7522 ( P1_ADD_95_U82 , P1_ADD_95_U11 );
not NOT1_7523 ( P1_ADD_95_U83 , P1_ADD_95_U13 );
not NOT1_7524 ( P1_ADD_95_U84 , P1_ADD_95_U16 );
not NOT1_7525 ( P1_ADD_95_U85 , P1_ADD_95_U17 );
not NOT1_7526 ( P1_ADD_95_U86 , P1_ADD_95_U19 );
not NOT1_7527 ( P1_ADD_95_U87 , P1_ADD_95_U21 );
not NOT1_7528 ( P1_ADD_95_U88 , P1_ADD_95_U23 );
not NOT1_7529 ( P1_ADD_95_U89 , P1_ADD_95_U25 );
not NOT1_7530 ( P1_ADD_95_U90 , P1_ADD_95_U27 );
not NOT1_7531 ( P1_ADD_95_U91 , P1_ADD_95_U29 );
not NOT1_7532 ( P1_ADD_95_U92 , P1_ADD_95_U31 );
not NOT1_7533 ( P1_ADD_95_U93 , P1_ADD_95_U33 );
not NOT1_7534 ( P1_ADD_95_U94 , P1_ADD_95_U35 );
not NOT1_7535 ( P1_ADD_95_U95 , P1_ADD_95_U37 );
not NOT1_7536 ( P1_ADD_95_U96 , P1_ADD_95_U39 );
not NOT1_7537 ( P1_ADD_95_U97 , P1_ADD_95_U41 );
not NOT1_7538 ( P1_ADD_95_U98 , P1_ADD_95_U43 );
not NOT1_7539 ( P1_ADD_95_U99 , P1_ADD_95_U45 );
not NOT1_7540 ( P1_ADD_95_U100 , P1_ADD_95_U47 );
not NOT1_7541 ( P1_ADD_95_U101 , P1_ADD_95_U49 );
not NOT1_7542 ( P1_ADD_95_U102 , P1_ADD_95_U51 );
not NOT1_7543 ( P1_ADD_95_U103 , P1_ADD_95_U79 );
nand NAND2_7544 ( P1_ADD_95_U104 , P1_REG3_REG_9_ , P1_ADD_95_U16 );
nand NAND2_7545 ( P1_ADD_95_U105 , P1_ADD_95_U84 , P1_ADD_95_U15 );
nand NAND2_7546 ( P1_ADD_95_U106 , P1_REG3_REG_8_ , P1_ADD_95_U13 );
nand NAND2_7547 ( P1_ADD_95_U107 , P1_ADD_95_U83 , P1_ADD_95_U14 );
nand NAND2_7548 ( P1_ADD_95_U108 , P1_REG3_REG_7_ , P1_ADD_95_U11 );
nand NAND2_7549 ( P1_ADD_95_U109 , P1_ADD_95_U82 , P1_ADD_95_U12 );
nand NAND2_7550 ( P1_ADD_95_U110 , P1_REG3_REG_6_ , P1_ADD_95_U9 );
nand NAND2_7551 ( P1_ADD_95_U111 , P1_ADD_95_U81 , P1_ADD_95_U10 );
nand NAND2_7552 ( P1_ADD_95_U112 , P1_REG3_REG_5_ , P1_ADD_95_U7 );
nand NAND2_7553 ( P1_ADD_95_U113 , P1_ADD_95_U80 , P1_ADD_95_U8 );
nand NAND2_7554 ( P1_ADD_95_U114 , P1_REG3_REG_4_ , P1_ADD_95_U4 );
nand NAND2_7555 ( P1_ADD_95_U115 , P1_REG3_REG_3_ , P1_ADD_95_U6 );
nand NAND2_7556 ( P1_ADD_95_U116 , P1_REG3_REG_28_ , P1_ADD_95_U79 );
nand NAND2_7557 ( P1_ADD_95_U117 , P1_ADD_95_U103 , P1_ADD_95_U52 );
nand NAND2_7558 ( P1_ADD_95_U118 , P1_REG3_REG_27_ , P1_ADD_95_U51 );
nand NAND2_7559 ( P1_ADD_95_U119 , P1_ADD_95_U102 , P1_ADD_95_U53 );
nand NAND2_7560 ( P1_ADD_95_U120 , P1_REG3_REG_26_ , P1_ADD_95_U49 );
nand NAND2_7561 ( P1_ADD_95_U121 , P1_ADD_95_U101 , P1_ADD_95_U50 );
nand NAND2_7562 ( P1_ADD_95_U122 , P1_REG3_REG_25_ , P1_ADD_95_U47 );
nand NAND2_7563 ( P1_ADD_95_U123 , P1_ADD_95_U100 , P1_ADD_95_U48 );
nand NAND2_7564 ( P1_ADD_95_U124 , P1_REG3_REG_24_ , P1_ADD_95_U45 );
nand NAND2_7565 ( P1_ADD_95_U125 , P1_ADD_95_U99 , P1_ADD_95_U46 );
nand NAND2_7566 ( P1_ADD_95_U126 , P1_REG3_REG_23_ , P1_ADD_95_U43 );
nand NAND2_7567 ( P1_ADD_95_U127 , P1_ADD_95_U98 , P1_ADD_95_U44 );
nand NAND2_7568 ( P1_ADD_95_U128 , P1_REG3_REG_22_ , P1_ADD_95_U41 );
nand NAND2_7569 ( P1_ADD_95_U129 , P1_ADD_95_U97 , P1_ADD_95_U42 );
nand NAND2_7570 ( P1_ADD_95_U130 , P1_REG3_REG_21_ , P1_ADD_95_U39 );
nand NAND2_7571 ( P1_ADD_95_U131 , P1_ADD_95_U96 , P1_ADD_95_U40 );
nand NAND2_7572 ( P1_ADD_95_U132 , P1_REG3_REG_20_ , P1_ADD_95_U37 );
nand NAND2_7573 ( P1_ADD_95_U133 , P1_ADD_95_U95 , P1_ADD_95_U38 );
nand NAND2_7574 ( P1_ADD_95_U134 , P1_REG3_REG_19_ , P1_ADD_95_U35 );
nand NAND2_7575 ( P1_ADD_95_U135 , P1_ADD_95_U94 , P1_ADD_95_U36 );
nand NAND2_7576 ( P1_ADD_95_U136 , P1_REG3_REG_18_ , P1_ADD_95_U33 );
nand NAND2_7577 ( P1_ADD_95_U137 , P1_ADD_95_U93 , P1_ADD_95_U34 );
nand NAND2_7578 ( P1_ADD_95_U138 , P1_REG3_REG_17_ , P1_ADD_95_U31 );
nand NAND2_7579 ( P1_ADD_95_U139 , P1_ADD_95_U92 , P1_ADD_95_U32 );
nand NAND2_7580 ( P1_ADD_95_U140 , P1_REG3_REG_16_ , P1_ADD_95_U29 );
nand NAND2_7581 ( P1_ADD_95_U141 , P1_ADD_95_U91 , P1_ADD_95_U30 );
nand NAND2_7582 ( P1_ADD_95_U142 , P1_REG3_REG_15_ , P1_ADD_95_U27 );
nand NAND2_7583 ( P1_ADD_95_U143 , P1_ADD_95_U90 , P1_ADD_95_U28 );
nand NAND2_7584 ( P1_ADD_95_U144 , P1_REG3_REG_14_ , P1_ADD_95_U25 );
nand NAND2_7585 ( P1_ADD_95_U145 , P1_ADD_95_U89 , P1_ADD_95_U26 );
nand NAND2_7586 ( P1_ADD_95_U146 , P1_REG3_REG_13_ , P1_ADD_95_U23 );
nand NAND2_7587 ( P1_ADD_95_U147 , P1_ADD_95_U88 , P1_ADD_95_U24 );
nand NAND2_7588 ( P1_ADD_95_U148 , P1_REG3_REG_12_ , P1_ADD_95_U21 );
nand NAND2_7589 ( P1_ADD_95_U149 , P1_ADD_95_U87 , P1_ADD_95_U22 );
nand NAND2_7590 ( P1_ADD_95_U150 , P1_REG3_REG_11_ , P1_ADD_95_U19 );
nand NAND2_7591 ( P1_ADD_95_U151 , P1_ADD_95_U86 , P1_ADD_95_U20 );
nand NAND2_7592 ( P1_ADD_95_U152 , P1_REG3_REG_10_ , P1_ADD_95_U17 );
nand NAND2_7593 ( P1_ADD_95_U153 , P1_ADD_95_U85 , P1_ADD_95_U18 );
and AND2_7594 ( P1_R1105_U4 , P1_R1105_U95 , P1_R1105_U94 );
and AND2_7595 ( P1_R1105_U5 , P1_R1105_U96 , P1_R1105_U97 );
and AND2_7596 ( P1_R1105_U6 , P1_R1105_U113 , P1_R1105_U112 );
and AND2_7597 ( P1_R1105_U7 , P1_R1105_U155 , P1_R1105_U154 );
and AND2_7598 ( P1_R1105_U8 , P1_R1105_U164 , P1_R1105_U163 );
and AND2_7599 ( P1_R1105_U9 , P1_R1105_U182 , P1_R1105_U181 );
and AND2_7600 ( P1_R1105_U10 , P1_R1105_U218 , P1_R1105_U215 );
and AND2_7601 ( P1_R1105_U11 , P1_R1105_U211 , P1_R1105_U208 );
and AND2_7602 ( P1_R1105_U12 , P1_R1105_U202 , P1_R1105_U199 );
and AND2_7603 ( P1_R1105_U13 , P1_R1105_U196 , P1_R1105_U192 );
and AND2_7604 ( P1_R1105_U14 , P1_R1105_U151 , P1_R1105_U148 );
and AND2_7605 ( P1_R1105_U15 , P1_R1105_U143 , P1_R1105_U140 );
and AND2_7606 ( P1_R1105_U16 , P1_R1105_U129 , P1_R1105_U126 );
not NOT1_7607 ( P1_R1105_U17 , P1_REG2_REG_6_ );
not NOT1_7608 ( P1_R1105_U18 , P1_U3469 );
not NOT1_7609 ( P1_R1105_U19 , P1_U3472 );
nand NAND2_7610 ( P1_R1105_U20 , P1_U3469 , P1_REG2_REG_6_ );
not NOT1_7611 ( P1_R1105_U21 , P1_REG2_REG_7_ );
not NOT1_7612 ( P1_R1105_U22 , P1_REG2_REG_4_ );
not NOT1_7613 ( P1_R1105_U23 , P1_U3463 );
not NOT1_7614 ( P1_R1105_U24 , P1_U3466 );
not NOT1_7615 ( P1_R1105_U25 , P1_REG2_REG_2_ );
not NOT1_7616 ( P1_R1105_U26 , P1_U3457 );
not NOT1_7617 ( P1_R1105_U27 , P1_REG2_REG_0_ );
not NOT1_7618 ( P1_R1105_U28 , P1_U3448 );
nand NAND2_7619 ( P1_R1105_U29 , P1_U3448 , P1_REG2_REG_0_ );
not NOT1_7620 ( P1_R1105_U30 , P1_REG2_REG_3_ );
not NOT1_7621 ( P1_R1105_U31 , P1_U3460 );
nand NAND2_7622 ( P1_R1105_U32 , P1_U3463 , P1_REG2_REG_4_ );
not NOT1_7623 ( P1_R1105_U33 , P1_REG2_REG_5_ );
not NOT1_7624 ( P1_R1105_U34 , P1_REG2_REG_8_ );
not NOT1_7625 ( P1_R1105_U35 , P1_U3475 );
not NOT1_7626 ( P1_R1105_U36 , P1_U3478 );
not NOT1_7627 ( P1_R1105_U37 , P1_REG2_REG_9_ );
nand NAND2_7628 ( P1_R1105_U38 , P1_R1105_U49 , P1_R1105_U121 );
nand NAND3_7629 ( P1_R1105_U39 , P1_R1105_U110 , P1_R1105_U108 , P1_R1105_U109 );
nand NAND2_7630 ( P1_R1105_U40 , P1_R1105_U98 , P1_R1105_U99 );
nand NAND2_7631 ( P1_R1105_U41 , P1_REG2_REG_1_ , P1_U3454 );
nand NAND3_7632 ( P1_R1105_U42 , P1_R1105_U136 , P1_R1105_U134 , P1_R1105_U135 );
nand NAND2_7633 ( P1_R1105_U43 , P1_R1105_U132 , P1_R1105_U131 );
not NOT1_7634 ( P1_R1105_U44 , P1_REG2_REG_16_ );
not NOT1_7635 ( P1_R1105_U45 , P1_U3499 );
not NOT1_7636 ( P1_R1105_U46 , P1_U3502 );
nand NAND2_7637 ( P1_R1105_U47 , P1_U3499 , P1_REG2_REG_16_ );
not NOT1_7638 ( P1_R1105_U48 , P1_REG2_REG_17_ );
nand NAND2_7639 ( P1_R1105_U49 , P1_U3475 , P1_REG2_REG_8_ );
not NOT1_7640 ( P1_R1105_U50 , P1_REG2_REG_10_ );
not NOT1_7641 ( P1_R1105_U51 , P1_U3481 );
not NOT1_7642 ( P1_R1105_U52 , P1_REG2_REG_12_ );
not NOT1_7643 ( P1_R1105_U53 , P1_U3487 );
not NOT1_7644 ( P1_R1105_U54 , P1_REG2_REG_11_ );
not NOT1_7645 ( P1_R1105_U55 , P1_U3484 );
nand NAND2_7646 ( P1_R1105_U56 , P1_U3484 , P1_REG2_REG_11_ );
not NOT1_7647 ( P1_R1105_U57 , P1_REG2_REG_13_ );
not NOT1_7648 ( P1_R1105_U58 , P1_U3490 );
not NOT1_7649 ( P1_R1105_U59 , P1_REG2_REG_14_ );
not NOT1_7650 ( P1_R1105_U60 , P1_U3493 );
not NOT1_7651 ( P1_R1105_U61 , P1_REG2_REG_15_ );
not NOT1_7652 ( P1_R1105_U62 , P1_U3496 );
not NOT1_7653 ( P1_R1105_U63 , P1_REG2_REG_18_ );
not NOT1_7654 ( P1_R1105_U64 , P1_U3505 );
nand NAND3_7655 ( P1_R1105_U65 , P1_R1105_U186 , P1_R1105_U185 , P1_R1105_U187 );
nand NAND2_7656 ( P1_R1105_U66 , P1_R1105_U179 , P1_R1105_U178 );
nand NAND2_7657 ( P1_R1105_U67 , P1_R1105_U56 , P1_R1105_U204 );
nand NAND2_7658 ( P1_R1105_U68 , P1_R1105_U259 , P1_R1105_U258 );
nand NAND2_7659 ( P1_R1105_U69 , P1_R1105_U308 , P1_R1105_U307 );
nand NAND2_7660 ( P1_R1105_U70 , P1_R1105_U231 , P1_R1105_U230 );
nand NAND2_7661 ( P1_R1105_U71 , P1_R1105_U236 , P1_R1105_U235 );
nand NAND2_7662 ( P1_R1105_U72 , P1_R1105_U243 , P1_R1105_U242 );
nand NAND2_7663 ( P1_R1105_U73 , P1_R1105_U250 , P1_R1105_U249 );
nand NAND2_7664 ( P1_R1105_U74 , P1_R1105_U255 , P1_R1105_U254 );
nand NAND2_7665 ( P1_R1105_U75 , P1_R1105_U271 , P1_R1105_U270 );
nand NAND2_7666 ( P1_R1105_U76 , P1_R1105_U278 , P1_R1105_U277 );
nand NAND2_7667 ( P1_R1105_U77 , P1_R1105_U285 , P1_R1105_U284 );
nand NAND2_7668 ( P1_R1105_U78 , P1_R1105_U292 , P1_R1105_U291 );
nand NAND2_7669 ( P1_R1105_U79 , P1_R1105_U299 , P1_R1105_U298 );
nand NAND2_7670 ( P1_R1105_U80 , P1_R1105_U304 , P1_R1105_U303 );
nand NAND3_7671 ( P1_R1105_U81 , P1_R1105_U117 , P1_R1105_U116 , P1_R1105_U118 );
nand NAND2_7672 ( P1_R1105_U82 , P1_R1105_U133 , P1_R1105_U145 );
nand NAND2_7673 ( P1_R1105_U83 , P1_R1105_U41 , P1_R1105_U152 );
not NOT1_7674 ( P1_R1105_U84 , P1_U3442 );
not NOT1_7675 ( P1_R1105_U85 , P1_REG2_REG_19_ );
nand NAND2_7676 ( P1_R1105_U86 , P1_R1105_U175 , P1_R1105_U174 );
nand NAND2_7677 ( P1_R1105_U87 , P1_R1105_U171 , P1_R1105_U170 );
nand NAND2_7678 ( P1_R1105_U88 , P1_R1105_U161 , P1_R1105_U160 );
not NOT1_7679 ( P1_R1105_U89 , P1_R1105_U32 );
nand NAND2_7680 ( P1_R1105_U90 , P1_REG2_REG_9_ , P1_U3478 );
nand NAND2_7681 ( P1_R1105_U91 , P1_U3487 , P1_REG2_REG_12_ );
not NOT1_7682 ( P1_R1105_U92 , P1_R1105_U56 );
not NOT1_7683 ( P1_R1105_U93 , P1_R1105_U49 );
or OR2_7684 ( P1_R1105_U94 , P1_U3466 , P1_REG2_REG_5_ );
or OR2_7685 ( P1_R1105_U95 , P1_U3463 , P1_REG2_REG_4_ );
or OR2_7686 ( P1_R1105_U96 , P1_REG2_REG_3_ , P1_U3460 );
or OR2_7687 ( P1_R1105_U97 , P1_REG2_REG_2_ , P1_U3457 );
not NOT1_7688 ( P1_R1105_U98 , P1_R1105_U29 );
or OR2_7689 ( P1_R1105_U99 , P1_REG2_REG_1_ , P1_U3454 );
not NOT1_7690 ( P1_R1105_U100 , P1_R1105_U40 );
not NOT1_7691 ( P1_R1105_U101 , P1_R1105_U41 );
nand NAND2_7692 ( P1_R1105_U102 , P1_R1105_U40 , P1_R1105_U41 );
nand NAND3_7693 ( P1_R1105_U103 , P1_REG2_REG_2_ , P1_U3457 , P1_R1105_U96 );
nand NAND2_7694 ( P1_R1105_U104 , P1_R1105_U5 , P1_R1105_U102 );
nand NAND2_7695 ( P1_R1105_U105 , P1_U3460 , P1_REG2_REG_3_ );
nand NAND3_7696 ( P1_R1105_U106 , P1_R1105_U105 , P1_R1105_U103 , P1_R1105_U104 );
nand NAND2_7697 ( P1_R1105_U107 , P1_R1105_U33 , P1_R1105_U32 );
nand NAND2_7698 ( P1_R1105_U108 , P1_U3466 , P1_R1105_U107 );
nand NAND2_7699 ( P1_R1105_U109 , P1_R1105_U4 , P1_R1105_U106 );
nand NAND2_7700 ( P1_R1105_U110 , P1_REG2_REG_5_ , P1_R1105_U89 );
not NOT1_7701 ( P1_R1105_U111 , P1_R1105_U39 );
or OR2_7702 ( P1_R1105_U112 , P1_U3472 , P1_REG2_REG_7_ );
or OR2_7703 ( P1_R1105_U113 , P1_U3469 , P1_REG2_REG_6_ );
not NOT1_7704 ( P1_R1105_U114 , P1_R1105_U20 );
nand NAND2_7705 ( P1_R1105_U115 , P1_R1105_U21 , P1_R1105_U20 );
nand NAND2_7706 ( P1_R1105_U116 , P1_U3472 , P1_R1105_U115 );
nand NAND2_7707 ( P1_R1105_U117 , P1_REG2_REG_7_ , P1_R1105_U114 );
nand NAND2_7708 ( P1_R1105_U118 , P1_R1105_U6 , P1_R1105_U39 );
not NOT1_7709 ( P1_R1105_U119 , P1_R1105_U81 );
or OR2_7710 ( P1_R1105_U120 , P1_REG2_REG_8_ , P1_U3475 );
nand NAND2_7711 ( P1_R1105_U121 , P1_R1105_U120 , P1_R1105_U81 );
not NOT1_7712 ( P1_R1105_U122 , P1_R1105_U38 );
or OR2_7713 ( P1_R1105_U123 , P1_U3478 , P1_REG2_REG_9_ );
or OR2_7714 ( P1_R1105_U124 , P1_REG2_REG_6_ , P1_U3469 );
nand NAND2_7715 ( P1_R1105_U125 , P1_R1105_U124 , P1_R1105_U39 );
nand NAND4_7716 ( P1_R1105_U126 , P1_R1105_U238 , P1_R1105_U237 , P1_R1105_U20 , P1_R1105_U125 );
nand NAND2_7717 ( P1_R1105_U127 , P1_R1105_U111 , P1_R1105_U20 );
nand NAND2_7718 ( P1_R1105_U128 , P1_REG2_REG_7_ , P1_U3472 );
nand NAND3_7719 ( P1_R1105_U129 , P1_R1105_U128 , P1_R1105_U6 , P1_R1105_U127 );
or OR2_7720 ( P1_R1105_U130 , P1_U3469 , P1_REG2_REG_6_ );
nand NAND2_7721 ( P1_R1105_U131 , P1_R1105_U101 , P1_R1105_U97 );
nand NAND2_7722 ( P1_R1105_U132 , P1_U3457 , P1_REG2_REG_2_ );
not NOT1_7723 ( P1_R1105_U133 , P1_R1105_U43 );
nand NAND2_7724 ( P1_R1105_U134 , P1_R1105_U100 , P1_R1105_U5 );
nand NAND2_7725 ( P1_R1105_U135 , P1_R1105_U43 , P1_R1105_U96 );
nand NAND2_7726 ( P1_R1105_U136 , P1_U3460 , P1_REG2_REG_3_ );
not NOT1_7727 ( P1_R1105_U137 , P1_R1105_U42 );
or OR2_7728 ( P1_R1105_U138 , P1_REG2_REG_4_ , P1_U3463 );
nand NAND2_7729 ( P1_R1105_U139 , P1_R1105_U138 , P1_R1105_U42 );
nand NAND4_7730 ( P1_R1105_U140 , P1_R1105_U245 , P1_R1105_U244 , P1_R1105_U32 , P1_R1105_U139 );
nand NAND2_7731 ( P1_R1105_U141 , P1_R1105_U137 , P1_R1105_U32 );
nand NAND2_7732 ( P1_R1105_U142 , P1_REG2_REG_5_ , P1_U3466 );
nand NAND3_7733 ( P1_R1105_U143 , P1_R1105_U142 , P1_R1105_U4 , P1_R1105_U141 );
or OR2_7734 ( P1_R1105_U144 , P1_U3463 , P1_REG2_REG_4_ );
nand NAND2_7735 ( P1_R1105_U145 , P1_R1105_U100 , P1_R1105_U97 );
not NOT1_7736 ( P1_R1105_U146 , P1_R1105_U82 );
nand NAND2_7737 ( P1_R1105_U147 , P1_U3460 , P1_REG2_REG_3_ );
nand NAND4_7738 ( P1_R1105_U148 , P1_R1105_U41 , P1_R1105_U40 , P1_R1105_U257 , P1_R1105_U256 );
nand NAND2_7739 ( P1_R1105_U149 , P1_R1105_U41 , P1_R1105_U40 );
nand NAND2_7740 ( P1_R1105_U150 , P1_U3457 , P1_REG2_REG_2_ );
nand NAND3_7741 ( P1_R1105_U151 , P1_R1105_U150 , P1_R1105_U97 , P1_R1105_U149 );
or OR2_7742 ( P1_R1105_U152 , P1_REG2_REG_1_ , P1_U3454 );
not NOT1_7743 ( P1_R1105_U153 , P1_R1105_U83 );
or OR2_7744 ( P1_R1105_U154 , P1_U3478 , P1_REG2_REG_9_ );
or OR2_7745 ( P1_R1105_U155 , P1_U3481 , P1_REG2_REG_10_ );
nand NAND2_7746 ( P1_R1105_U156 , P1_R1105_U93 , P1_R1105_U7 );
nand NAND2_7747 ( P1_R1105_U157 , P1_U3481 , P1_REG2_REG_10_ );
nand NAND3_7748 ( P1_R1105_U158 , P1_R1105_U157 , P1_R1105_U90 , P1_R1105_U156 );
or OR2_7749 ( P1_R1105_U159 , P1_REG2_REG_10_ , P1_U3481 );
nand NAND3_7750 ( P1_R1105_U160 , P1_R1105_U120 , P1_R1105_U7 , P1_R1105_U81 );
nand NAND2_7751 ( P1_R1105_U161 , P1_R1105_U159 , P1_R1105_U158 );
not NOT1_7752 ( P1_R1105_U162 , P1_R1105_U88 );
or OR2_7753 ( P1_R1105_U163 , P1_U3490 , P1_REG2_REG_13_ );
or OR2_7754 ( P1_R1105_U164 , P1_U3487 , P1_REG2_REG_12_ );
nand NAND2_7755 ( P1_R1105_U165 , P1_R1105_U92 , P1_R1105_U8 );
nand NAND2_7756 ( P1_R1105_U166 , P1_U3490 , P1_REG2_REG_13_ );
nand NAND3_7757 ( P1_R1105_U167 , P1_R1105_U166 , P1_R1105_U91 , P1_R1105_U165 );
or OR2_7758 ( P1_R1105_U168 , P1_REG2_REG_11_ , P1_U3484 );
or OR2_7759 ( P1_R1105_U169 , P1_REG2_REG_13_ , P1_U3490 );
nand NAND3_7760 ( P1_R1105_U170 , P1_R1105_U168 , P1_R1105_U8 , P1_R1105_U88 );
nand NAND2_7761 ( P1_R1105_U171 , P1_R1105_U169 , P1_R1105_U167 );
not NOT1_7762 ( P1_R1105_U172 , P1_R1105_U87 );
or OR2_7763 ( P1_R1105_U173 , P1_REG2_REG_14_ , P1_U3493 );
nand NAND2_7764 ( P1_R1105_U174 , P1_R1105_U173 , P1_R1105_U87 );
nand NAND2_7765 ( P1_R1105_U175 , P1_U3493 , P1_REG2_REG_14_ );
not NOT1_7766 ( P1_R1105_U176 , P1_R1105_U86 );
or OR2_7767 ( P1_R1105_U177 , P1_REG2_REG_15_ , P1_U3496 );
nand NAND2_7768 ( P1_R1105_U178 , P1_R1105_U177 , P1_R1105_U86 );
nand NAND2_7769 ( P1_R1105_U179 , P1_U3496 , P1_REG2_REG_15_ );
not NOT1_7770 ( P1_R1105_U180 , P1_R1105_U66 );
or OR2_7771 ( P1_R1105_U181 , P1_U3502 , P1_REG2_REG_17_ );
or OR2_7772 ( P1_R1105_U182 , P1_U3499 , P1_REG2_REG_16_ );
not NOT1_7773 ( P1_R1105_U183 , P1_R1105_U47 );
nand NAND2_7774 ( P1_R1105_U184 , P1_R1105_U48 , P1_R1105_U47 );
nand NAND2_7775 ( P1_R1105_U185 , P1_U3502 , P1_R1105_U184 );
nand NAND2_7776 ( P1_R1105_U186 , P1_REG2_REG_17_ , P1_R1105_U183 );
nand NAND2_7777 ( P1_R1105_U187 , P1_R1105_U9 , P1_R1105_U66 );
not NOT1_7778 ( P1_R1105_U188 , P1_R1105_U65 );
or OR2_7779 ( P1_R1105_U189 , P1_REG2_REG_18_ , P1_U3505 );
nand NAND2_7780 ( P1_R1105_U190 , P1_R1105_U189 , P1_R1105_U65 );
nand NAND2_7781 ( P1_R1105_U191 , P1_U3505 , P1_REG2_REG_18_ );
nand NAND4_7782 ( P1_R1105_U192 , P1_R1105_U261 , P1_R1105_U260 , P1_R1105_U191 , P1_R1105_U190 );
nand NAND2_7783 ( P1_R1105_U193 , P1_U3505 , P1_REG2_REG_18_ );
nand NAND2_7784 ( P1_R1105_U194 , P1_R1105_U188 , P1_R1105_U193 );
or OR2_7785 ( P1_R1105_U195 , P1_U3505 , P1_REG2_REG_18_ );
nand NAND3_7786 ( P1_R1105_U196 , P1_R1105_U195 , P1_R1105_U264 , P1_R1105_U194 );
or OR2_7787 ( P1_R1105_U197 , P1_REG2_REG_16_ , P1_U3499 );
nand NAND2_7788 ( P1_R1105_U198 , P1_R1105_U197 , P1_R1105_U66 );
nand NAND4_7789 ( P1_R1105_U199 , P1_R1105_U273 , P1_R1105_U272 , P1_R1105_U47 , P1_R1105_U198 );
nand NAND2_7790 ( P1_R1105_U200 , P1_R1105_U180 , P1_R1105_U47 );
nand NAND2_7791 ( P1_R1105_U201 , P1_REG2_REG_17_ , P1_U3502 );
nand NAND3_7792 ( P1_R1105_U202 , P1_R1105_U201 , P1_R1105_U9 , P1_R1105_U200 );
or OR2_7793 ( P1_R1105_U203 , P1_U3499 , P1_REG2_REG_16_ );
nand NAND2_7794 ( P1_R1105_U204 , P1_R1105_U168 , P1_R1105_U88 );
not NOT1_7795 ( P1_R1105_U205 , P1_R1105_U67 );
or OR2_7796 ( P1_R1105_U206 , P1_REG2_REG_12_ , P1_U3487 );
nand NAND2_7797 ( P1_R1105_U207 , P1_R1105_U206 , P1_R1105_U67 );
nand NAND4_7798 ( P1_R1105_U208 , P1_R1105_U294 , P1_R1105_U293 , P1_R1105_U91 , P1_R1105_U207 );
nand NAND2_7799 ( P1_R1105_U209 , P1_R1105_U205 , P1_R1105_U91 );
nand NAND2_7800 ( P1_R1105_U210 , P1_U3490 , P1_REG2_REG_13_ );
nand NAND3_7801 ( P1_R1105_U211 , P1_R1105_U210 , P1_R1105_U8 , P1_R1105_U209 );
or OR2_7802 ( P1_R1105_U212 , P1_U3487 , P1_REG2_REG_12_ );
or OR2_7803 ( P1_R1105_U213 , P1_REG2_REG_9_ , P1_U3478 );
nand NAND2_7804 ( P1_R1105_U214 , P1_R1105_U213 , P1_R1105_U38 );
nand NAND4_7805 ( P1_R1105_U215 , P1_R1105_U306 , P1_R1105_U305 , P1_R1105_U90 , P1_R1105_U214 );
nand NAND2_7806 ( P1_R1105_U216 , P1_R1105_U122 , P1_R1105_U90 );
nand NAND2_7807 ( P1_R1105_U217 , P1_U3481 , P1_REG2_REG_10_ );
nand NAND3_7808 ( P1_R1105_U218 , P1_R1105_U217 , P1_R1105_U7 , P1_R1105_U216 );
nand NAND2_7809 ( P1_R1105_U219 , P1_R1105_U123 , P1_R1105_U90 );
nand NAND2_7810 ( P1_R1105_U220 , P1_R1105_U120 , P1_R1105_U49 );
nand NAND2_7811 ( P1_R1105_U221 , P1_R1105_U130 , P1_R1105_U20 );
nand NAND2_7812 ( P1_R1105_U222 , P1_R1105_U144 , P1_R1105_U32 );
nand NAND2_7813 ( P1_R1105_U223 , P1_R1105_U147 , P1_R1105_U96 );
nand NAND2_7814 ( P1_R1105_U224 , P1_R1105_U203 , P1_R1105_U47 );
nand NAND2_7815 ( P1_R1105_U225 , P1_R1105_U212 , P1_R1105_U91 );
nand NAND2_7816 ( P1_R1105_U226 , P1_R1105_U168 , P1_R1105_U56 );
nand NAND2_7817 ( P1_R1105_U227 , P1_U3478 , P1_R1105_U37 );
nand NAND2_7818 ( P1_R1105_U228 , P1_REG2_REG_9_ , P1_R1105_U36 );
nand NAND2_7819 ( P1_R1105_U229 , P1_R1105_U228 , P1_R1105_U227 );
nand NAND2_7820 ( P1_R1105_U230 , P1_R1105_U219 , P1_R1105_U38 );
nand NAND2_7821 ( P1_R1105_U231 , P1_R1105_U229 , P1_R1105_U122 );
nand NAND2_7822 ( P1_R1105_U232 , P1_U3475 , P1_R1105_U34 );
nand NAND2_7823 ( P1_R1105_U233 , P1_REG2_REG_8_ , P1_R1105_U35 );
nand NAND2_7824 ( P1_R1105_U234 , P1_R1105_U233 , P1_R1105_U232 );
nand NAND2_7825 ( P1_R1105_U235 , P1_R1105_U220 , P1_R1105_U81 );
nand NAND2_7826 ( P1_R1105_U236 , P1_R1105_U119 , P1_R1105_U234 );
nand NAND2_7827 ( P1_R1105_U237 , P1_U3472 , P1_R1105_U21 );
nand NAND2_7828 ( P1_R1105_U238 , P1_REG2_REG_7_ , P1_R1105_U19 );
nand NAND2_7829 ( P1_R1105_U239 , P1_U3469 , P1_R1105_U17 );
nand NAND2_7830 ( P1_R1105_U240 , P1_REG2_REG_6_ , P1_R1105_U18 );
nand NAND2_7831 ( P1_R1105_U241 , P1_R1105_U240 , P1_R1105_U239 );
nand NAND2_7832 ( P1_R1105_U242 , P1_R1105_U221 , P1_R1105_U39 );
nand NAND2_7833 ( P1_R1105_U243 , P1_R1105_U241 , P1_R1105_U111 );
nand NAND2_7834 ( P1_R1105_U244 , P1_U3466 , P1_R1105_U33 );
nand NAND2_7835 ( P1_R1105_U245 , P1_REG2_REG_5_ , P1_R1105_U24 );
nand NAND2_7836 ( P1_R1105_U246 , P1_U3463 , P1_R1105_U22 );
nand NAND2_7837 ( P1_R1105_U247 , P1_REG2_REG_4_ , P1_R1105_U23 );
nand NAND2_7838 ( P1_R1105_U248 , P1_R1105_U247 , P1_R1105_U246 );
nand NAND2_7839 ( P1_R1105_U249 , P1_R1105_U222 , P1_R1105_U42 );
nand NAND2_7840 ( P1_R1105_U250 , P1_R1105_U248 , P1_R1105_U137 );
nand NAND2_7841 ( P1_R1105_U251 , P1_U3460 , P1_R1105_U30 );
nand NAND2_7842 ( P1_R1105_U252 , P1_REG2_REG_3_ , P1_R1105_U31 );
nand NAND2_7843 ( P1_R1105_U253 , P1_R1105_U252 , P1_R1105_U251 );
nand NAND2_7844 ( P1_R1105_U254 , P1_R1105_U223 , P1_R1105_U82 );
nand NAND2_7845 ( P1_R1105_U255 , P1_R1105_U146 , P1_R1105_U253 );
nand NAND2_7846 ( P1_R1105_U256 , P1_U3457 , P1_R1105_U25 );
nand NAND2_7847 ( P1_R1105_U257 , P1_REG2_REG_2_ , P1_R1105_U26 );
nand NAND2_7848 ( P1_R1105_U258 , P1_R1105_U98 , P1_R1105_U83 );
nand NAND2_7849 ( P1_R1105_U259 , P1_R1105_U153 , P1_R1105_U29 );
nand NAND2_7850 ( P1_R1105_U260 , P1_U3442 , P1_R1105_U85 );
nand NAND2_7851 ( P1_R1105_U261 , P1_REG2_REG_19_ , P1_R1105_U84 );
nand NAND2_7852 ( P1_R1105_U262 , P1_U3442 , P1_R1105_U85 );
nand NAND2_7853 ( P1_R1105_U263 , P1_REG2_REG_19_ , P1_R1105_U84 );
nand NAND2_7854 ( P1_R1105_U264 , P1_R1105_U263 , P1_R1105_U262 );
nand NAND2_7855 ( P1_R1105_U265 , P1_U3505 , P1_R1105_U63 );
nand NAND2_7856 ( P1_R1105_U266 , P1_REG2_REG_18_ , P1_R1105_U64 );
nand NAND2_7857 ( P1_R1105_U267 , P1_U3505 , P1_R1105_U63 );
nand NAND2_7858 ( P1_R1105_U268 , P1_REG2_REG_18_ , P1_R1105_U64 );
nand NAND2_7859 ( P1_R1105_U269 , P1_R1105_U268 , P1_R1105_U267 );
nand NAND3_7860 ( P1_R1105_U270 , P1_R1105_U266 , P1_R1105_U265 , P1_R1105_U65 );
nand NAND2_7861 ( P1_R1105_U271 , P1_R1105_U269 , P1_R1105_U188 );
nand NAND2_7862 ( P1_R1105_U272 , P1_U3502 , P1_R1105_U48 );
nand NAND2_7863 ( P1_R1105_U273 , P1_REG2_REG_17_ , P1_R1105_U46 );
nand NAND2_7864 ( P1_R1105_U274 , P1_U3499 , P1_R1105_U44 );
nand NAND2_7865 ( P1_R1105_U275 , P1_REG2_REG_16_ , P1_R1105_U45 );
nand NAND2_7866 ( P1_R1105_U276 , P1_R1105_U275 , P1_R1105_U274 );
nand NAND2_7867 ( P1_R1105_U277 , P1_R1105_U224 , P1_R1105_U66 );
nand NAND2_7868 ( P1_R1105_U278 , P1_R1105_U276 , P1_R1105_U180 );
nand NAND2_7869 ( P1_R1105_U279 , P1_U3496 , P1_R1105_U61 );
nand NAND2_7870 ( P1_R1105_U280 , P1_REG2_REG_15_ , P1_R1105_U62 );
nand NAND2_7871 ( P1_R1105_U281 , P1_U3496 , P1_R1105_U61 );
nand NAND2_7872 ( P1_R1105_U282 , P1_REG2_REG_15_ , P1_R1105_U62 );
nand NAND2_7873 ( P1_R1105_U283 , P1_R1105_U282 , P1_R1105_U281 );
nand NAND3_7874 ( P1_R1105_U284 , P1_R1105_U280 , P1_R1105_U279 , P1_R1105_U86 );
nand NAND2_7875 ( P1_R1105_U285 , P1_R1105_U176 , P1_R1105_U283 );
nand NAND2_7876 ( P1_R1105_U286 , P1_U3493 , P1_R1105_U59 );
nand NAND2_7877 ( P1_R1105_U287 , P1_REG2_REG_14_ , P1_R1105_U60 );
nand NAND2_7878 ( P1_R1105_U288 , P1_U3493 , P1_R1105_U59 );
nand NAND2_7879 ( P1_R1105_U289 , P1_REG2_REG_14_ , P1_R1105_U60 );
nand NAND2_7880 ( P1_R1105_U290 , P1_R1105_U289 , P1_R1105_U288 );
nand NAND3_7881 ( P1_R1105_U291 , P1_R1105_U287 , P1_R1105_U286 , P1_R1105_U87 );
nand NAND2_7882 ( P1_R1105_U292 , P1_R1105_U172 , P1_R1105_U290 );
nand NAND2_7883 ( P1_R1105_U293 , P1_U3490 , P1_R1105_U57 );
nand NAND2_7884 ( P1_R1105_U294 , P1_REG2_REG_13_ , P1_R1105_U58 );
nand NAND2_7885 ( P1_R1105_U295 , P1_U3487 , P1_R1105_U52 );
nand NAND2_7886 ( P1_R1105_U296 , P1_REG2_REG_12_ , P1_R1105_U53 );
nand NAND2_7887 ( P1_R1105_U297 , P1_R1105_U296 , P1_R1105_U295 );
nand NAND2_7888 ( P1_R1105_U298 , P1_R1105_U225 , P1_R1105_U67 );
nand NAND2_7889 ( P1_R1105_U299 , P1_R1105_U297 , P1_R1105_U205 );
nand NAND2_7890 ( P1_R1105_U300 , P1_U3484 , P1_R1105_U54 );
nand NAND2_7891 ( P1_R1105_U301 , P1_REG2_REG_11_ , P1_R1105_U55 );
nand NAND2_7892 ( P1_R1105_U302 , P1_R1105_U301 , P1_R1105_U300 );
nand NAND2_7893 ( P1_R1105_U303 , P1_R1105_U226 , P1_R1105_U88 );
nand NAND2_7894 ( P1_R1105_U304 , P1_R1105_U162 , P1_R1105_U302 );
nand NAND2_7895 ( P1_R1105_U305 , P1_U3481 , P1_R1105_U50 );
nand NAND2_7896 ( P1_R1105_U306 , P1_REG2_REG_10_ , P1_R1105_U51 );
nand NAND2_7897 ( P1_R1105_U307 , P1_U3448 , P1_R1105_U27 );
nand NAND2_7898 ( P1_R1105_U308 , P1_REG2_REG_0_ , P1_R1105_U28 );
and AND2_7899 ( P1_SUB_84_U6 , P1_SUB_84_U227 , P1_SUB_84_U38 );
and AND2_7900 ( P1_SUB_84_U7 , P1_SUB_84_U225 , P1_SUB_84_U192 );
and AND2_7901 ( P1_SUB_84_U8 , P1_SUB_84_U224 , P1_SUB_84_U35 );
and AND2_7902 ( P1_SUB_84_U9 , P1_SUB_84_U223 , P1_SUB_84_U36 );
and AND2_7903 ( P1_SUB_84_U10 , P1_SUB_84_U221 , P1_SUB_84_U195 );
and AND2_7904 ( P1_SUB_84_U11 , P1_SUB_84_U220 , P1_SUB_84_U34 );
and AND2_7905 ( P1_SUB_84_U12 , P1_SUB_84_U219 , P1_SUB_84_U197 );
and AND2_7906 ( P1_SUB_84_U13 , P1_SUB_84_U217 , P1_SUB_84_U198 );
and AND2_7907 ( P1_SUB_84_U14 , P1_SUB_84_U216 , P1_SUB_84_U172 );
and AND2_7908 ( P1_SUB_84_U15 , P1_SUB_84_U215 , P1_SUB_84_U200 );
and AND2_7909 ( P1_SUB_84_U16 , P1_SUB_84_U213 , P1_SUB_84_U201 );
and AND2_7910 ( P1_SUB_84_U17 , P1_SUB_84_U212 , P1_SUB_84_U169 );
and AND2_7911 ( P1_SUB_84_U18 , P1_SUB_84_U211 , P1_SUB_84_U167 );
and AND2_7912 ( P1_SUB_84_U19 , P1_SUB_84_U209 , P1_SUB_84_U204 );
and AND2_7913 ( P1_SUB_84_U20 , P1_SUB_84_U208 , P1_SUB_84_U33 );
and AND2_7914 ( P1_SUB_84_U21 , P1_SUB_84_U207 , P1_SUB_84_U27 );
and AND2_7915 ( P1_SUB_84_U22 , P1_SUB_84_U190 , P1_SUB_84_U180 );
and AND2_7916 ( P1_SUB_84_U23 , P1_SUB_84_U189 , P1_SUB_84_U29 );
and AND2_7917 ( P1_SUB_84_U24 , P1_SUB_84_U188 , P1_SUB_84_U30 );
and AND2_7918 ( P1_SUB_84_U25 , P1_SUB_84_U186 , P1_SUB_84_U183 );
and AND2_7919 ( P1_SUB_84_U26 , P1_SUB_84_U185 , P1_SUB_84_U28 );
or OR3_7920 ( P1_SUB_84_U27 , P1_IR_REG_1_ , P1_IR_REG_0_ , P1_IR_REG_2_ );
nand NAND3_7921 ( P1_SUB_84_U28 , P1_SUB_84_U44 , P1_SUB_84_U230 , P1_SUB_84_U43 );
nand NAND2_7922 ( P1_SUB_84_U29 , P1_SUB_84_U45 , P1_SUB_84_U230 );
nand NAND2_7923 ( P1_SUB_84_U30 , P1_SUB_84_U46 , P1_SUB_84_U181 );
not NOT1_7924 ( P1_SUB_84_U31 , P1_IR_REG_7_ );
not NOT1_7925 ( P1_SUB_84_U32 , P1_IR_REG_3_ );
nand NAND2_7926 ( P1_SUB_84_U33 , P1_SUB_84_U56 , P1_SUB_84_U51 );
nand NAND4_7927 ( P1_SUB_84_U34 , P1_SUB_84_U130 , P1_SUB_84_U129 , P1_SUB_84_U128 , P1_SUB_84_U127 );
nand NAND2_7928 ( P1_SUB_84_U35 , P1_SUB_84_U156 , P1_SUB_84_U184 );
nand NAND2_7929 ( P1_SUB_84_U36 , P1_SUB_84_U157 , P1_SUB_84_U193 );
not NOT1_7930 ( P1_SUB_84_U37 , P1_IR_REG_15_ );
nand NAND2_7931 ( P1_SUB_84_U38 , P1_SUB_84_U158 , P1_SUB_84_U184 );
not NOT1_7932 ( P1_SUB_84_U39 , P1_IR_REG_11_ );
nand NAND2_7933 ( P1_SUB_84_U40 , P1_SUB_84_U247 , P1_SUB_84_U246 );
nand NAND2_7934 ( P1_SUB_84_U41 , P1_SUB_84_U237 , P1_SUB_84_U236 );
nand NAND2_7935 ( P1_SUB_84_U42 , P1_SUB_84_U241 , P1_SUB_84_U240 );
nor nor_7936 ( P1_SUB_84_U43 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_7937 ( P1_SUB_84_U44 , P1_IR_REG_7_ , P1_IR_REG_8_ );
nor nor_7938 ( P1_SUB_84_U45 , P1_IR_REG_3_ , P1_IR_REG_4_ );
nor nor_7939 ( P1_SUB_84_U46 , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_7940 ( P1_SUB_84_U47 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_7941 ( P1_SUB_84_U48 , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_7942 ( P1_SUB_84_U49 , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_7943 ( P1_SUB_84_U50 , P1_IR_REG_22_ , P1_IR_REG_20_ , P1_IR_REG_21_ );
and AND4_7944 ( P1_SUB_84_U51 , P1_SUB_84_U50 , P1_SUB_84_U49 , P1_SUB_84_U48 , P1_SUB_84_U47 );
nor nor_7945 ( P1_SUB_84_U52 , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ );
nor nor_7946 ( P1_SUB_84_U53 , P1_IR_REG_27_ , P1_IR_REG_28_ , P1_IR_REG_29_ , P1_IR_REG_2_ );
nor nor_7947 ( P1_SUB_84_U54 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_7948 ( P1_SUB_84_U55 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_7949 ( P1_SUB_84_U56 , P1_SUB_84_U55 , P1_SUB_84_U54 , P1_SUB_84_U53 , P1_SUB_84_U52 );
nor nor_7950 ( P1_SUB_84_U57 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_7951 ( P1_SUB_84_U58 , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_7952 ( P1_SUB_84_U59 , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_7953 ( P1_SUB_84_U60 , P1_IR_REG_22_ , P1_IR_REG_20_ , P1_IR_REG_21_ );
and AND4_7954 ( P1_SUB_84_U61 , P1_SUB_84_U60 , P1_SUB_84_U59 , P1_SUB_84_U58 , P1_SUB_84_U57 );
nor nor_7955 ( P1_SUB_84_U62 , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ );
nor nor_7956 ( P1_SUB_84_U63 , P1_IR_REG_2_ , P1_IR_REG_27_ , P1_IR_REG_28_ );
nor nor_7957 ( P1_SUB_84_U64 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_7958 ( P1_SUB_84_U65 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_7959 ( P1_SUB_84_U66 , P1_SUB_84_U65 , P1_SUB_84_U64 , P1_SUB_84_U63 , P1_SUB_84_U62 );
nor nor_7960 ( P1_SUB_84_U67 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_7961 ( P1_SUB_84_U68 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_7962 ( P1_SUB_84_U69 , P1_IR_REG_17_ , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
nor nor_7963 ( P1_SUB_84_U70 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
and AND4_7964 ( P1_SUB_84_U71 , P1_SUB_84_U70 , P1_SUB_84_U69 , P1_SUB_84_U68 , P1_SUB_84_U67 );
nor nor_7965 ( P1_SUB_84_U72 , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ );
nor nor_7966 ( P1_SUB_84_U73 , P1_IR_REG_2_ , P1_IR_REG_26_ , P1_IR_REG_27_ );
nor nor_7967 ( P1_SUB_84_U74 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_7968 ( P1_SUB_84_U75 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_7969 ( P1_SUB_84_U76 , P1_SUB_84_U75 , P1_SUB_84_U74 , P1_SUB_84_U73 , P1_SUB_84_U72 );
nor nor_7970 ( P1_SUB_84_U77 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_7971 ( P1_SUB_84_U78 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_7972 ( P1_SUB_84_U79 , P1_IR_REG_17_ , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
nor nor_7973 ( P1_SUB_84_U80 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
and AND4_7974 ( P1_SUB_84_U81 , P1_SUB_84_U80 , P1_SUB_84_U79 , P1_SUB_84_U78 , P1_SUB_84_U77 );
nor nor_7975 ( P1_SUB_84_U82 , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ );
nor nor_7976 ( P1_SUB_84_U83 , P1_IR_REG_3_ , P1_IR_REG_26_ , P1_IR_REG_2_ );
nor nor_7977 ( P1_SUB_84_U84 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_7978 ( P1_SUB_84_U85 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_7979 ( P1_SUB_84_U86 , P1_SUB_84_U85 , P1_SUB_84_U84 , P1_SUB_84_U83 , P1_SUB_84_U82 );
nor nor_7980 ( P1_SUB_84_U87 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_7981 ( P1_SUB_84_U88 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_7982 ( P1_SUB_84_U89 , P1_IR_REG_17_ , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
nor nor_7983 ( P1_SUB_84_U90 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
and AND4_7984 ( P1_SUB_84_U91 , P1_SUB_84_U90 , P1_SUB_84_U89 , P1_SUB_84_U88 , P1_SUB_84_U87 );
nor nor_7985 ( P1_SUB_84_U92 , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ );
nor nor_7986 ( P1_SUB_84_U93 , P1_IR_REG_3_ , P1_IR_REG_26_ , P1_IR_REG_2_ );
nor nor_7987 ( P1_SUB_84_U94 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_7988 ( P1_SUB_84_U95 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_7989 ( P1_SUB_84_U96 , P1_SUB_84_U95 , P1_SUB_84_U94 , P1_SUB_84_U93 , P1_SUB_84_U92 );
nor nor_7990 ( P1_SUB_84_U97 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_7991 ( P1_SUB_84_U98 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_7992 ( P1_SUB_84_U99 , P1_IR_REG_19_ , P1_IR_REG_17_ , P1_IR_REG_18_ );
nor nor_7993 ( P1_SUB_84_U100 , P1_IR_REG_20_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
and AND4_7994 ( P1_SUB_84_U101 , P1_SUB_84_U100 , P1_SUB_84_U99 , P1_SUB_84_U98 , P1_SUB_84_U97 );
nor nor_7995 ( P1_SUB_84_U102 , P1_IR_REG_21_ , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ );
nor nor_7996 ( P1_SUB_84_U103 , P1_IR_REG_3_ , P1_IR_REG_25_ , P1_IR_REG_2_ );
nor nor_7997 ( P1_SUB_84_U104 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_7998 ( P1_SUB_84_U105 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_7999 ( P1_SUB_84_U106 , P1_SUB_84_U105 , P1_SUB_84_U104 , P1_SUB_84_U103 , P1_SUB_84_U102 );
nor nor_8000 ( P1_SUB_84_U107 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_8001 ( P1_SUB_84_U108 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_8002 ( P1_SUB_84_U109 , P1_IR_REG_19_ , P1_IR_REG_17_ , P1_IR_REG_18_ );
nor nor_8003 ( P1_SUB_84_U110 , P1_IR_REG_20_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
and AND4_8004 ( P1_SUB_84_U111 , P1_SUB_84_U110 , P1_SUB_84_U109 , P1_SUB_84_U108 , P1_SUB_84_U107 );
nor nor_8005 ( P1_SUB_84_U112 , P1_IR_REG_23_ , P1_IR_REG_21_ , P1_IR_REG_22_ );
nor nor_8006 ( P1_SUB_84_U113 , P1_IR_REG_3_ , P1_IR_REG_24_ , P1_IR_REG_2_ );
nor nor_8007 ( P1_SUB_84_U114 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_8008 ( P1_SUB_84_U115 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_8009 ( P1_SUB_84_U116 , P1_SUB_84_U115 , P1_SUB_84_U114 , P1_SUB_84_U113 , P1_SUB_84_U112 );
nor nor_8010 ( P1_SUB_84_U117 , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8011 ( P1_SUB_84_U118 , P1_IR_REG_15_ , P1_IR_REG_13_ , P1_IR_REG_14_ );
nor nor_8012 ( P1_SUB_84_U119 , P1_IR_REG_18_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_8013 ( P1_SUB_84_U120 , P1_IR_REG_0_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
and AND4_8014 ( P1_SUB_84_U121 , P1_SUB_84_U120 , P1_SUB_84_U119 , P1_SUB_84_U118 , P1_SUB_84_U117 );
nor nor_8015 ( P1_SUB_84_U122 , P1_IR_REG_22_ , P1_IR_REG_20_ , P1_IR_REG_21_ );
nor nor_8016 ( P1_SUB_84_U123 , P1_IR_REG_3_ , P1_IR_REG_23_ , P1_IR_REG_2_ );
nor nor_8017 ( P1_SUB_84_U124 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_8018 ( P1_SUB_84_U125 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_8019 ( P1_SUB_84_U126 , P1_SUB_84_U125 , P1_SUB_84_U124 , P1_SUB_84_U123 , P1_SUB_84_U122 );
nor nor_8020 ( P1_SUB_84_U127 , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8021 ( P1_SUB_84_U128 , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_8022 ( P1_SUB_84_U129 , P1_IR_REG_2_ , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_8023 ( P1_SUB_84_U130 , P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ );
nor nor_8024 ( P1_SUB_84_U131 , P1_IR_REG_17_ , P1_IR_REG_18_ );
nor nor_8025 ( P1_SUB_84_U132 , P1_IR_REG_19_ , P1_IR_REG_20_ );
nor nor_8026 ( P1_SUB_84_U133 , P1_IR_REG_21_ , P1_IR_REG_22_ );
and AND3_8027 ( P1_SUB_84_U134 , P1_SUB_84_U132 , P1_SUB_84_U131 , P1_SUB_84_U133 );
nor nor_8028 ( P1_SUB_84_U135 , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8029 ( P1_SUB_84_U136 , P1_IR_REG_15_ , P1_IR_REG_13_ , P1_IR_REG_14_ );
and AND2_8030 ( P1_SUB_84_U137 , P1_SUB_84_U136 , P1_SUB_84_U135 );
nor nor_8031 ( P1_SUB_84_U138 , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_18_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_8032 ( P1_SUB_84_U139 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
nor nor_8033 ( P1_SUB_84_U140 , P1_IR_REG_4_ , P1_IR_REG_2_ , P1_IR_REG_3_ );
and AND2_8034 ( P1_SUB_84_U141 , P1_SUB_84_U140 , P1_SUB_84_U139 );
nor nor_8035 ( P1_SUB_84_U142 , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8036 ( P1_SUB_84_U143 , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8037 ( P1_SUB_84_U144 , P1_IR_REG_15_ , P1_IR_REG_13_ , P1_IR_REG_14_ );
nor nor_8038 ( P1_SUB_84_U145 , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_18_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_8039 ( P1_SUB_84_U146 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_2_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
nor nor_8040 ( P1_SUB_84_U147 , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8041 ( P1_SUB_84_U148 , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8042 ( P1_SUB_84_U149 , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_17_ , P1_IR_REG_15_ , P1_IR_REG_16_ );
nor nor_8043 ( P1_SUB_84_U150 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_2_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_8044 ( P1_SUB_84_U151 , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_8045 ( P1_SUB_84_U152 , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_8046 ( P1_SUB_84_U153 , P1_IR_REG_18_ , P1_IR_REG_1_ , P1_IR_REG_17_ , P1_IR_REG_15_ , P1_IR_REG_16_ );
nor nor_8047 ( P1_SUB_84_U154 , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_3_ , P1_IR_REG_0_ , P1_IR_REG_2_ );
nor nor_8048 ( P1_SUB_84_U155 , P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ );
nor nor_8049 ( P1_SUB_84_U156 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_9_ );
nor nor_8050 ( P1_SUB_84_U157 , P1_IR_REG_13_ , P1_IR_REG_14_ );
nor nor_8051 ( P1_SUB_84_U158 , P1_IR_REG_10_ , P1_IR_REG_9_ );
not NOT1_8052 ( P1_SUB_84_U159 , P1_IR_REG_9_ );
and AND2_8053 ( P1_SUB_84_U160 , P1_SUB_84_U233 , P1_SUB_84_U232 );
not NOT1_8054 ( P1_SUB_84_U161 , P1_IR_REG_5_ );
and AND2_8055 ( P1_SUB_84_U162 , P1_SUB_84_U235 , P1_SUB_84_U234 );
not NOT1_8056 ( P1_SUB_84_U163 , P1_IR_REG_31_ );
not NOT1_8057 ( P1_SUB_84_U164 , P1_IR_REG_30_ );
and AND2_8058 ( P1_SUB_84_U165 , P1_SUB_84_U239 , P1_SUB_84_U238 );
not NOT1_8059 ( P1_SUB_84_U166 , P1_IR_REG_27_ );
nand NAND2_8060 ( P1_SUB_84_U167 , P1_SUB_84_U96 , P1_SUB_84_U91 );
not NOT1_8061 ( P1_SUB_84_U168 , P1_IR_REG_25_ );
nand NAND2_8062 ( P1_SUB_84_U169 , P1_SUB_84_U116 , P1_SUB_84_U111 );
and AND2_8063 ( P1_SUB_84_U170 , P1_SUB_84_U243 , P1_SUB_84_U242 );
not NOT1_8064 ( P1_SUB_84_U171 , P1_IR_REG_21_ );
nand NAND5_8065 ( P1_SUB_84_U172 , P1_SUB_84_U144 , P1_SUB_84_U143 , P1_SUB_84_U145 , P1_SUB_84_U147 , P1_SUB_84_U146 );
and AND2_8066 ( P1_SUB_84_U173 , P1_SUB_84_U245 , P1_SUB_84_U244 );
not NOT1_8067 ( P1_SUB_84_U174 , P1_IR_REG_1_ );
not NOT1_8068 ( P1_SUB_84_U175 , P1_IR_REG_0_ );
not NOT1_8069 ( P1_SUB_84_U176 , P1_IR_REG_17_ );
and AND2_8070 ( P1_SUB_84_U177 , P1_SUB_84_U249 , P1_SUB_84_U248 );
not NOT1_8071 ( P1_SUB_84_U178 , P1_IR_REG_13_ );
and AND2_8072 ( P1_SUB_84_U179 , P1_SUB_84_U251 , P1_SUB_84_U250 );
nand NAND2_8073 ( P1_SUB_84_U180 , P1_SUB_84_U230 , P1_SUB_84_U32 );
not NOT1_8074 ( P1_SUB_84_U181 , P1_SUB_84_U29 );
not NOT1_8075 ( P1_SUB_84_U182 , P1_SUB_84_U30 );
nand NAND2_8076 ( P1_SUB_84_U183 , P1_SUB_84_U182 , P1_SUB_84_U31 );
not NOT1_8077 ( P1_SUB_84_U184 , P1_SUB_84_U28 );
nand NAND2_8078 ( P1_SUB_84_U185 , P1_IR_REG_8_ , P1_SUB_84_U183 );
nand NAND2_8079 ( P1_SUB_84_U186 , P1_IR_REG_7_ , P1_SUB_84_U30 );
nand NAND2_8080 ( P1_SUB_84_U187 , P1_SUB_84_U181 , P1_SUB_84_U161 );
nand NAND2_8081 ( P1_SUB_84_U188 , P1_IR_REG_6_ , P1_SUB_84_U187 );
nand NAND2_8082 ( P1_SUB_84_U189 , P1_IR_REG_4_ , P1_SUB_84_U180 );
nand NAND2_8083 ( P1_SUB_84_U190 , P1_IR_REG_3_ , P1_SUB_84_U27 );
not NOT1_8084 ( P1_SUB_84_U191 , P1_SUB_84_U38 );
nand NAND2_8085 ( P1_SUB_84_U192 , P1_SUB_84_U191 , P1_SUB_84_U39 );
not NOT1_8086 ( P1_SUB_84_U193 , P1_SUB_84_U35 );
not NOT1_8087 ( P1_SUB_84_U194 , P1_SUB_84_U36 );
nand NAND2_8088 ( P1_SUB_84_U195 , P1_SUB_84_U194 , P1_SUB_84_U37 );
not NOT1_8089 ( P1_SUB_84_U196 , P1_SUB_84_U34 );
nand NAND4_8090 ( P1_SUB_84_U197 , P1_SUB_84_U155 , P1_SUB_84_U154 , P1_SUB_84_U153 , P1_SUB_84_U152 );
nand NAND4_8091 ( P1_SUB_84_U198 , P1_SUB_84_U151 , P1_SUB_84_U150 , P1_SUB_84_U149 , P1_SUB_84_U148 );
not NOT1_8092 ( P1_SUB_84_U199 , P1_SUB_84_U172 );
nand NAND2_8093 ( P1_SUB_84_U200 , P1_SUB_84_U134 , P1_SUB_84_U196 );
nand NAND2_8094 ( P1_SUB_84_U201 , P1_SUB_84_U126 , P1_SUB_84_U121 );
not NOT1_8095 ( P1_SUB_84_U202 , P1_SUB_84_U169 );
not NOT1_8096 ( P1_SUB_84_U203 , P1_SUB_84_U167 );
nand NAND2_8097 ( P1_SUB_84_U204 , P1_SUB_84_U66 , P1_SUB_84_U61 );
not NOT1_8098 ( P1_SUB_84_U205 , P1_SUB_84_U33 );
or OR2_8099 ( P1_SUB_84_U206 , P1_IR_REG_1_ , P1_IR_REG_0_ );
nand NAND2_8100 ( P1_SUB_84_U207 , P1_IR_REG_2_ , P1_SUB_84_U206 );
nand NAND2_8101 ( P1_SUB_84_U208 , P1_IR_REG_29_ , P1_SUB_84_U204 );
nand NAND2_8102 ( P1_SUB_84_U209 , P1_IR_REG_28_ , P1_SUB_84_U229 );
nand NAND2_8103 ( P1_SUB_84_U210 , P1_SUB_84_U106 , P1_SUB_84_U101 );
nand NAND2_8104 ( P1_SUB_84_U211 , P1_IR_REG_26_ , P1_SUB_84_U210 );
nand NAND2_8105 ( P1_SUB_84_U212 , P1_IR_REG_24_ , P1_SUB_84_U201 );
nand NAND2_8106 ( P1_SUB_84_U213 , P1_IR_REG_23_ , P1_SUB_84_U200 );
nand NAND4_8107 ( P1_SUB_84_U214 , P1_SUB_84_U142 , P1_SUB_84_U141 , P1_SUB_84_U138 , P1_SUB_84_U137 );
nand NAND2_8108 ( P1_SUB_84_U215 , P1_IR_REG_22_ , P1_SUB_84_U214 );
nand NAND2_8109 ( P1_SUB_84_U216 , P1_IR_REG_20_ , P1_SUB_84_U198 );
nand NAND2_8110 ( P1_SUB_84_U217 , P1_IR_REG_19_ , P1_SUB_84_U197 );
nand NAND2_8111 ( P1_SUB_84_U218 , P1_SUB_84_U196 , P1_SUB_84_U176 );
nand NAND2_8112 ( P1_SUB_84_U219 , P1_IR_REG_18_ , P1_SUB_84_U218 );
nand NAND2_8113 ( P1_SUB_84_U220 , P1_IR_REG_16_ , P1_SUB_84_U195 );
nand NAND2_8114 ( P1_SUB_84_U221 , P1_IR_REG_15_ , P1_SUB_84_U36 );
nand NAND2_8115 ( P1_SUB_84_U222 , P1_SUB_84_U193 , P1_SUB_84_U178 );
nand NAND2_8116 ( P1_SUB_84_U223 , P1_IR_REG_14_ , P1_SUB_84_U222 );
nand NAND2_8117 ( P1_SUB_84_U224 , P1_IR_REG_12_ , P1_SUB_84_U192 );
nand NAND2_8118 ( P1_SUB_84_U225 , P1_IR_REG_11_ , P1_SUB_84_U38 );
nand NAND2_8119 ( P1_SUB_84_U226 , P1_SUB_84_U184 , P1_SUB_84_U159 );
nand NAND2_8120 ( P1_SUB_84_U227 , P1_IR_REG_10_ , P1_SUB_84_U226 );
nand NAND2_8121 ( P1_SUB_84_U228 , P1_SUB_84_U205 , P1_SUB_84_U164 );
nand NAND2_8122 ( P1_SUB_84_U229 , P1_SUB_84_U76 , P1_SUB_84_U71 );
not NOT1_8123 ( P1_SUB_84_U230 , P1_SUB_84_U27 );
nand NAND2_8124 ( P1_SUB_84_U231 , P1_SUB_84_U86 , P1_SUB_84_U81 );
nand NAND2_8125 ( P1_SUB_84_U232 , P1_IR_REG_9_ , P1_SUB_84_U28 );
nand NAND2_8126 ( P1_SUB_84_U233 , P1_SUB_84_U184 , P1_SUB_84_U159 );
nand NAND2_8127 ( P1_SUB_84_U234 , P1_IR_REG_5_ , P1_SUB_84_U29 );
nand NAND2_8128 ( P1_SUB_84_U235 , P1_SUB_84_U181 , P1_SUB_84_U161 );
nand NAND2_8129 ( P1_SUB_84_U236 , P1_SUB_84_U228 , P1_SUB_84_U163 );
nand NAND3_8130 ( P1_SUB_84_U237 , P1_SUB_84_U205 , P1_SUB_84_U164 , P1_IR_REG_31_ );
nand NAND2_8131 ( P1_SUB_84_U238 , P1_IR_REG_30_ , P1_SUB_84_U33 );
nand NAND2_8132 ( P1_SUB_84_U239 , P1_SUB_84_U205 , P1_SUB_84_U164 );
nand NAND2_8133 ( P1_SUB_84_U240 , P1_SUB_84_U203 , P1_IR_REG_27_ );
nand NAND2_8134 ( P1_SUB_84_U241 , P1_SUB_84_U231 , P1_SUB_84_U166 );
nand NAND2_8135 ( P1_SUB_84_U242 , P1_IR_REG_25_ , P1_SUB_84_U169 );
nand NAND2_8136 ( P1_SUB_84_U243 , P1_SUB_84_U202 , P1_SUB_84_U168 );
nand NAND2_8137 ( P1_SUB_84_U244 , P1_IR_REG_21_ , P1_SUB_84_U172 );
nand NAND2_8138 ( P1_SUB_84_U245 , P1_SUB_84_U199 , P1_SUB_84_U171 );
nand NAND2_8139 ( P1_SUB_84_U246 , P1_IR_REG_1_ , P1_SUB_84_U175 );
nand NAND2_8140 ( P1_SUB_84_U247 , P1_IR_REG_0_ , P1_SUB_84_U174 );
nand NAND2_8141 ( P1_SUB_84_U248 , P1_IR_REG_17_ , P1_SUB_84_U34 );
nand NAND2_8142 ( P1_SUB_84_U249 , P1_SUB_84_U196 , P1_SUB_84_U176 );
nand NAND2_8143 ( P1_SUB_84_U250 , P1_IR_REG_13_ , P1_SUB_84_U35 );
nand NAND2_8144 ( P1_SUB_84_U251 , P1_SUB_84_U193 , P1_SUB_84_U178 );
not NOT1_8145 ( P1_R1309_U6 , P1_U3059 );
not NOT1_8146 ( P1_R1309_U7 , P1_U3056 );
and AND2_8147 ( P1_R1309_U8 , P1_R1309_U10 , P1_R1309_U9 );
nand NAND2_8148 ( P1_R1309_U9 , P1_U3056 , P1_R1309_U6 );
nand NAND2_8149 ( P1_R1309_U10 , P1_U3059 , P1_R1309_U7 );
and AND2_8150 ( P1_R1282_U6 , P1_R1282_U135 , P1_R1282_U35 );
and AND2_8151 ( P1_R1282_U7 , P1_R1282_U133 , P1_R1282_U36 );
and AND2_8152 ( P1_R1282_U8 , P1_R1282_U132 , P1_R1282_U37 );
and AND2_8153 ( P1_R1282_U9 , P1_R1282_U131 , P1_R1282_U38 );
and AND2_8154 ( P1_R1282_U10 , P1_R1282_U129 , P1_R1282_U39 );
and AND2_8155 ( P1_R1282_U11 , P1_R1282_U128 , P1_R1282_U40 );
and AND2_8156 ( P1_R1282_U12 , P1_R1282_U127 , P1_R1282_U41 );
and AND2_8157 ( P1_R1282_U13 , P1_R1282_U125 , P1_R1282_U42 );
and AND2_8158 ( P1_R1282_U14 , P1_R1282_U123 , P1_R1282_U43 );
and AND2_8159 ( P1_R1282_U15 , P1_R1282_U121 , P1_R1282_U44 );
and AND2_8160 ( P1_R1282_U16 , P1_R1282_U119 , P1_R1282_U45 );
and AND2_8161 ( P1_R1282_U17 , P1_R1282_U117 , P1_R1282_U46 );
and AND2_8162 ( P1_R1282_U18 , P1_R1282_U115 , P1_R1282_U25 );
and AND2_8163 ( P1_R1282_U19 , P1_R1282_U113 , P1_R1282_U67 );
and AND2_8164 ( P1_R1282_U20 , P1_R1282_U98 , P1_R1282_U26 );
and AND2_8165 ( P1_R1282_U21 , P1_R1282_U97 , P1_R1282_U27 );
and AND2_8166 ( P1_R1282_U22 , P1_R1282_U96 , P1_R1282_U28 );
and AND2_8167 ( P1_R1282_U23 , P1_R1282_U94 , P1_R1282_U29 );
and AND2_8168 ( P1_R1282_U24 , P1_R1282_U93 , P1_R1282_U30 );
or OR3_8169 ( P1_R1282_U25 , P1_U3458 , P1_U3450 , P1_U3455 );
nand NAND2_8170 ( P1_R1282_U26 , P1_R1282_U87 , P1_R1282_U34 );
nand NAND2_8171 ( P1_R1282_U27 , P1_R1282_U88 , P1_R1282_U33 );
nand NAND2_8172 ( P1_R1282_U28 , P1_R1282_U58 , P1_R1282_U89 );
nand NAND2_8173 ( P1_R1282_U29 , P1_R1282_U90 , P1_R1282_U32 );
nand NAND2_8174 ( P1_R1282_U30 , P1_R1282_U91 , P1_R1282_U31 );
not NOT1_8175 ( P1_R1282_U31 , P1_U3476 );
not NOT1_8176 ( P1_R1282_U32 , P1_U3473 );
not NOT1_8177 ( P1_R1282_U33 , P1_U3464 );
not NOT1_8178 ( P1_R1282_U34 , P1_U3461 );
nand NAND2_8179 ( P1_R1282_U35 , P1_R1282_U59 , P1_R1282_U92 );
nand NAND2_8180 ( P1_R1282_U36 , P1_R1282_U99 , P1_R1282_U56 );
nand NAND2_8181 ( P1_R1282_U37 , P1_R1282_U100 , P1_R1282_U55 );
nand NAND2_8182 ( P1_R1282_U38 , P1_R1282_U60 , P1_R1282_U101 );
nand NAND2_8183 ( P1_R1282_U39 , P1_R1282_U102 , P1_R1282_U54 );
nand NAND2_8184 ( P1_R1282_U40 , P1_R1282_U103 , P1_R1282_U53 );
nand NAND2_8185 ( P1_R1282_U41 , P1_R1282_U61 , P1_R1282_U104 );
nand NAND3_8186 ( P1_R1282_U42 , P1_R1282_U105 , P1_R1282_U81 , P1_R1282_U52 );
nand NAND3_8187 ( P1_R1282_U43 , P1_R1282_U106 , P1_R1282_U77 , P1_R1282_U51 );
nand NAND3_8188 ( P1_R1282_U44 , P1_R1282_U107 , P1_R1282_U75 , P1_R1282_U50 );
nand NAND3_8189 ( P1_R1282_U45 , P1_R1282_U108 , P1_R1282_U73 , P1_R1282_U49 );
nand NAND3_8190 ( P1_R1282_U46 , P1_R1282_U109 , P1_R1282_U71 , P1_R1282_U48 );
not NOT1_8191 ( P1_R1282_U47 , P1_U3984 );
not NOT1_8192 ( P1_R1282_U48 , P1_U3974 );
not NOT1_8193 ( P1_R1282_U49 , P1_U3976 );
not NOT1_8194 ( P1_R1282_U50 , P1_U3978 );
not NOT1_8195 ( P1_R1282_U51 , P1_U3980 );
not NOT1_8196 ( P1_R1282_U52 , P1_U3982 );
not NOT1_8197 ( P1_R1282_U53 , P1_U3500 );
not NOT1_8198 ( P1_R1282_U54 , P1_U3497 );
not NOT1_8199 ( P1_R1282_U55 , P1_U3488 );
not NOT1_8200 ( P1_R1282_U56 , P1_U3485 );
nand NAND2_8201 ( P1_R1282_U57 , P1_R1282_U153 , P1_R1282_U152 );
nor nor_8202 ( P1_R1282_U58 , P1_U3467 , P1_U3470 );
nor nor_8203 ( P1_R1282_U59 , P1_U3482 , P1_U3479 );
nor nor_8204 ( P1_R1282_U60 , P1_U3491 , P1_U3494 );
nor nor_8205 ( P1_R1282_U61 , P1_U3503 , P1_U3506 );
not NOT1_8206 ( P1_R1282_U62 , P1_U3479 );
and AND2_8207 ( P1_R1282_U63 , P1_R1282_U137 , P1_R1282_U136 );
not NOT1_8208 ( P1_R1282_U64 , P1_U3467 );
and AND2_8209 ( P1_R1282_U65 , P1_R1282_U139 , P1_R1282_U138 );
not NOT1_8210 ( P1_R1282_U66 , P1_U3983 );
nand NAND3_8211 ( P1_R1282_U67 , P1_R1282_U110 , P1_R1282_U69 , P1_R1282_U47 );
and AND2_8212 ( P1_R1282_U68 , P1_R1282_U141 , P1_R1282_U140 );
not NOT1_8213 ( P1_R1282_U69 , P1_U3985 );
and AND2_8214 ( P1_R1282_U70 , P1_R1282_U143 , P1_R1282_U142 );
not NOT1_8215 ( P1_R1282_U71 , P1_U3975 );
and AND2_8216 ( P1_R1282_U72 , P1_R1282_U145 , P1_R1282_U144 );
not NOT1_8217 ( P1_R1282_U73 , P1_U3977 );
and AND2_8218 ( P1_R1282_U74 , P1_R1282_U147 , P1_R1282_U146 );
not NOT1_8219 ( P1_R1282_U75 , P1_U3979 );
and AND2_8220 ( P1_R1282_U76 , P1_R1282_U149 , P1_R1282_U148 );
not NOT1_8221 ( P1_R1282_U77 , P1_U3981 );
and AND2_8222 ( P1_R1282_U78 , P1_R1282_U151 , P1_R1282_U150 );
not NOT1_8223 ( P1_R1282_U79 , P1_U3455 );
not NOT1_8224 ( P1_R1282_U80 , P1_U3450 );
not NOT1_8225 ( P1_R1282_U81 , P1_U3508 );
and AND2_8226 ( P1_R1282_U82 , P1_R1282_U155 , P1_R1282_U154 );
not NOT1_8227 ( P1_R1282_U83 , P1_U3503 );
and AND2_8228 ( P1_R1282_U84 , P1_R1282_U157 , P1_R1282_U156 );
not NOT1_8229 ( P1_R1282_U85 , P1_U3491 );
and AND2_8230 ( P1_R1282_U86 , P1_R1282_U159 , P1_R1282_U158 );
not NOT1_8231 ( P1_R1282_U87 , P1_R1282_U25 );
not NOT1_8232 ( P1_R1282_U88 , P1_R1282_U26 );
not NOT1_8233 ( P1_R1282_U89 , P1_R1282_U27 );
not NOT1_8234 ( P1_R1282_U90 , P1_R1282_U28 );
not NOT1_8235 ( P1_R1282_U91 , P1_R1282_U29 );
not NOT1_8236 ( P1_R1282_U92 , P1_R1282_U30 );
nand NAND2_8237 ( P1_R1282_U93 , P1_U3476 , P1_R1282_U29 );
nand NAND2_8238 ( P1_R1282_U94 , P1_U3473 , P1_R1282_U28 );
nand NAND2_8239 ( P1_R1282_U95 , P1_R1282_U89 , P1_R1282_U64 );
nand NAND2_8240 ( P1_R1282_U96 , P1_U3470 , P1_R1282_U95 );
nand NAND2_8241 ( P1_R1282_U97 , P1_U3464 , P1_R1282_U26 );
nand NAND2_8242 ( P1_R1282_U98 , P1_U3461 , P1_R1282_U25 );
not NOT1_8243 ( P1_R1282_U99 , P1_R1282_U35 );
not NOT1_8244 ( P1_R1282_U100 , P1_R1282_U36 );
not NOT1_8245 ( P1_R1282_U101 , P1_R1282_U37 );
not NOT1_8246 ( P1_R1282_U102 , P1_R1282_U38 );
not NOT1_8247 ( P1_R1282_U103 , P1_R1282_U39 );
not NOT1_8248 ( P1_R1282_U104 , P1_R1282_U40 );
not NOT1_8249 ( P1_R1282_U105 , P1_R1282_U41 );
not NOT1_8250 ( P1_R1282_U106 , P1_R1282_U42 );
not NOT1_8251 ( P1_R1282_U107 , P1_R1282_U43 );
not NOT1_8252 ( P1_R1282_U108 , P1_R1282_U44 );
not NOT1_8253 ( P1_R1282_U109 , P1_R1282_U45 );
not NOT1_8254 ( P1_R1282_U110 , P1_R1282_U46 );
not NOT1_8255 ( P1_R1282_U111 , P1_R1282_U67 );
nand NAND2_8256 ( P1_R1282_U112 , P1_R1282_U110 , P1_R1282_U69 );
nand NAND2_8257 ( P1_R1282_U113 , P1_U3984 , P1_R1282_U112 );
or OR2_8258 ( P1_R1282_U114 , P1_U3455 , P1_U3450 );
nand NAND2_8259 ( P1_R1282_U115 , P1_U3458 , P1_R1282_U114 );
nand NAND2_8260 ( P1_R1282_U116 , P1_R1282_U109 , P1_R1282_U71 );
nand NAND2_8261 ( P1_R1282_U117 , P1_U3974 , P1_R1282_U116 );
nand NAND2_8262 ( P1_R1282_U118 , P1_R1282_U108 , P1_R1282_U73 );
nand NAND2_8263 ( P1_R1282_U119 , P1_U3976 , P1_R1282_U118 );
nand NAND2_8264 ( P1_R1282_U120 , P1_R1282_U107 , P1_R1282_U75 );
nand NAND2_8265 ( P1_R1282_U121 , P1_U3978 , P1_R1282_U120 );
nand NAND2_8266 ( P1_R1282_U122 , P1_R1282_U106 , P1_R1282_U77 );
nand NAND2_8267 ( P1_R1282_U123 , P1_U3980 , P1_R1282_U122 );
nand NAND2_8268 ( P1_R1282_U124 , P1_R1282_U105 , P1_R1282_U81 );
nand NAND2_8269 ( P1_R1282_U125 , P1_U3982 , P1_R1282_U124 );
nand NAND2_8270 ( P1_R1282_U126 , P1_R1282_U104 , P1_R1282_U83 );
nand NAND2_8271 ( P1_R1282_U127 , P1_U3506 , P1_R1282_U126 );
nand NAND2_8272 ( P1_R1282_U128 , P1_U3500 , P1_R1282_U39 );
nand NAND2_8273 ( P1_R1282_U129 , P1_U3497 , P1_R1282_U38 );
nand NAND2_8274 ( P1_R1282_U130 , P1_R1282_U101 , P1_R1282_U85 );
nand NAND2_8275 ( P1_R1282_U131 , P1_U3494 , P1_R1282_U130 );
nand NAND2_8276 ( P1_R1282_U132 , P1_U3488 , P1_R1282_U36 );
nand NAND2_8277 ( P1_R1282_U133 , P1_U3485 , P1_R1282_U35 );
nand NAND2_8278 ( P1_R1282_U134 , P1_R1282_U92 , P1_R1282_U62 );
nand NAND2_8279 ( P1_R1282_U135 , P1_U3482 , P1_R1282_U134 );
nand NAND2_8280 ( P1_R1282_U136 , P1_U3479 , P1_R1282_U30 );
nand NAND2_8281 ( P1_R1282_U137 , P1_R1282_U92 , P1_R1282_U62 );
nand NAND2_8282 ( P1_R1282_U138 , P1_U3467 , P1_R1282_U27 );
nand NAND2_8283 ( P1_R1282_U139 , P1_R1282_U89 , P1_R1282_U64 );
nand NAND2_8284 ( P1_R1282_U140 , P1_U3983 , P1_R1282_U67 );
nand NAND2_8285 ( P1_R1282_U141 , P1_R1282_U111 , P1_R1282_U66 );
nand NAND2_8286 ( P1_R1282_U142 , P1_U3985 , P1_R1282_U46 );
nand NAND2_8287 ( P1_R1282_U143 , P1_R1282_U110 , P1_R1282_U69 );
nand NAND2_8288 ( P1_R1282_U144 , P1_U3975 , P1_R1282_U45 );
nand NAND2_8289 ( P1_R1282_U145 , P1_R1282_U109 , P1_R1282_U71 );
nand NAND2_8290 ( P1_R1282_U146 , P1_U3977 , P1_R1282_U44 );
nand NAND2_8291 ( P1_R1282_U147 , P1_R1282_U108 , P1_R1282_U73 );
nand NAND2_8292 ( P1_R1282_U148 , P1_U3979 , P1_R1282_U43 );
nand NAND2_8293 ( P1_R1282_U149 , P1_R1282_U107 , P1_R1282_U75 );
nand NAND2_8294 ( P1_R1282_U150 , P1_U3981 , P1_R1282_U42 );
nand NAND2_8295 ( P1_R1282_U151 , P1_R1282_U106 , P1_R1282_U77 );
nand NAND2_8296 ( P1_R1282_U152 , P1_U3455 , P1_R1282_U80 );
nand NAND2_8297 ( P1_R1282_U153 , P1_U3450 , P1_R1282_U79 );
nand NAND2_8298 ( P1_R1282_U154 , P1_U3508 , P1_R1282_U41 );
nand NAND2_8299 ( P1_R1282_U155 , P1_R1282_U105 , P1_R1282_U81 );
nand NAND2_8300 ( P1_R1282_U156 , P1_U3503 , P1_R1282_U40 );
nand NAND2_8301 ( P1_R1282_U157 , P1_R1282_U104 , P1_R1282_U83 );
nand NAND2_8302 ( P1_R1282_U158 , P1_U3491 , P1_R1282_U37 );
nand NAND2_8303 ( P1_R1282_U159 , P1_R1282_U101 , P1_R1282_U85 );
and AND2_8304 ( P1_R1240_U4 , P1_R1240_U178 , P1_R1240_U177 );
and AND2_8305 ( P1_R1240_U5 , P1_R1240_U179 , P1_R1240_U180 );
and AND2_8306 ( P1_R1240_U6 , P1_R1240_U196 , P1_R1240_U195 );
and AND2_8307 ( P1_R1240_U7 , P1_R1240_U236 , P1_R1240_U235 );
and AND2_8308 ( P1_R1240_U8 , P1_R1240_U245 , P1_R1240_U244 );
and AND2_8309 ( P1_R1240_U9 , P1_R1240_U263 , P1_R1240_U262 );
and AND2_8310 ( P1_R1240_U10 , P1_R1240_U271 , P1_R1240_U270 );
and AND2_8311 ( P1_R1240_U11 , P1_R1240_U350 , P1_R1240_U347 );
and AND2_8312 ( P1_R1240_U12 , P1_R1240_U343 , P1_R1240_U340 );
and AND2_8313 ( P1_R1240_U13 , P1_R1240_U334 , P1_R1240_U331 );
and AND2_8314 ( P1_R1240_U14 , P1_R1240_U325 , P1_R1240_U322 );
and AND2_8315 ( P1_R1240_U15 , P1_R1240_U319 , P1_R1240_U317 );
and AND2_8316 ( P1_R1240_U16 , P1_R1240_U312 , P1_R1240_U309 );
and AND2_8317 ( P1_R1240_U17 , P1_R1240_U234 , P1_R1240_U231 );
and AND2_8318 ( P1_R1240_U18 , P1_R1240_U226 , P1_R1240_U223 );
and AND2_8319 ( P1_R1240_U19 , P1_R1240_U212 , P1_R1240_U209 );
not NOT1_8320 ( P1_R1240_U20 , P1_U3470 );
not NOT1_8321 ( P1_R1240_U21 , P1_U3071 );
not NOT1_8322 ( P1_R1240_U22 , P1_U3070 );
nand NAND2_8323 ( P1_R1240_U23 , P1_U3071 , P1_U3470 );
not NOT1_8324 ( P1_R1240_U24 , P1_U3473 );
not NOT1_8325 ( P1_R1240_U25 , P1_U3464 );
not NOT1_8326 ( P1_R1240_U26 , P1_U3060 );
not NOT1_8327 ( P1_R1240_U27 , P1_U3067 );
not NOT1_8328 ( P1_R1240_U28 , P1_U3458 );
not NOT1_8329 ( P1_R1240_U29 , P1_U3068 );
not NOT1_8330 ( P1_R1240_U30 , P1_U3450 );
not NOT1_8331 ( P1_R1240_U31 , P1_U3077 );
nand NAND2_8332 ( P1_R1240_U32 , P1_U3077 , P1_U3450 );
not NOT1_8333 ( P1_R1240_U33 , P1_U3461 );
not NOT1_8334 ( P1_R1240_U34 , P1_U3064 );
nand NAND2_8335 ( P1_R1240_U35 , P1_U3060 , P1_U3464 );
not NOT1_8336 ( P1_R1240_U36 , P1_U3467 );
not NOT1_8337 ( P1_R1240_U37 , P1_U3476 );
not NOT1_8338 ( P1_R1240_U38 , P1_U3084 );
not NOT1_8339 ( P1_R1240_U39 , P1_U3083 );
not NOT1_8340 ( P1_R1240_U40 , P1_U3479 );
nand NAND2_8341 ( P1_R1240_U41 , P1_R1240_U62 , P1_R1240_U204 );
nand NAND2_8342 ( P1_R1240_U42 , P1_R1240_U118 , P1_R1240_U192 );
nand NAND2_8343 ( P1_R1240_U43 , P1_R1240_U181 , P1_R1240_U182 );
nand NAND2_8344 ( P1_R1240_U44 , P1_U3455 , P1_U3078 );
nand NAND2_8345 ( P1_R1240_U45 , P1_R1240_U122 , P1_R1240_U218 );
nand NAND2_8346 ( P1_R1240_U46 , P1_R1240_U215 , P1_R1240_U214 );
not NOT1_8347 ( P1_R1240_U47 , P1_U3975 );
not NOT1_8348 ( P1_R1240_U48 , P1_U3053 );
not NOT1_8349 ( P1_R1240_U49 , P1_U3057 );
not NOT1_8350 ( P1_R1240_U50 , P1_U3976 );
not NOT1_8351 ( P1_R1240_U51 , P1_U3977 );
not NOT1_8352 ( P1_R1240_U52 , P1_U3058 );
not NOT1_8353 ( P1_R1240_U53 , P1_U3978 );
not NOT1_8354 ( P1_R1240_U54 , P1_U3065 );
not NOT1_8355 ( P1_R1240_U55 , P1_U3981 );
not NOT1_8356 ( P1_R1240_U56 , P1_U3075 );
not NOT1_8357 ( P1_R1240_U57 , P1_U3500 );
not NOT1_8358 ( P1_R1240_U58 , P1_U3073 );
not NOT1_8359 ( P1_R1240_U59 , P1_U3069 );
nand NAND2_8360 ( P1_R1240_U60 , P1_U3073 , P1_U3500 );
not NOT1_8361 ( P1_R1240_U61 , P1_U3503 );
nand NAND2_8362 ( P1_R1240_U62 , P1_U3084 , P1_U3476 );
not NOT1_8363 ( P1_R1240_U63 , P1_U3482 );
not NOT1_8364 ( P1_R1240_U64 , P1_U3062 );
not NOT1_8365 ( P1_R1240_U65 , P1_U3488 );
not NOT1_8366 ( P1_R1240_U66 , P1_U3072 );
not NOT1_8367 ( P1_R1240_U67 , P1_U3485 );
not NOT1_8368 ( P1_R1240_U68 , P1_U3063 );
nand NAND2_8369 ( P1_R1240_U69 , P1_U3063 , P1_U3485 );
not NOT1_8370 ( P1_R1240_U70 , P1_U3491 );
not NOT1_8371 ( P1_R1240_U71 , P1_U3080 );
not NOT1_8372 ( P1_R1240_U72 , P1_U3494 );
not NOT1_8373 ( P1_R1240_U73 , P1_U3079 );
not NOT1_8374 ( P1_R1240_U74 , P1_U3497 );
not NOT1_8375 ( P1_R1240_U75 , P1_U3074 );
not NOT1_8376 ( P1_R1240_U76 , P1_U3506 );
not NOT1_8377 ( P1_R1240_U77 , P1_U3082 );
nand NAND2_8378 ( P1_R1240_U78 , P1_U3082 , P1_U3506 );
not NOT1_8379 ( P1_R1240_U79 , P1_U3508 );
not NOT1_8380 ( P1_R1240_U80 , P1_U3081 );
nand NAND2_8381 ( P1_R1240_U81 , P1_U3081 , P1_U3508 );
not NOT1_8382 ( P1_R1240_U82 , P1_U3982 );
not NOT1_8383 ( P1_R1240_U83 , P1_U3980 );
not NOT1_8384 ( P1_R1240_U84 , P1_U3061 );
not NOT1_8385 ( P1_R1240_U85 , P1_U3979 );
not NOT1_8386 ( P1_R1240_U86 , P1_U3066 );
nand NAND2_8387 ( P1_R1240_U87 , P1_U3976 , P1_U3057 );
not NOT1_8388 ( P1_R1240_U88 , P1_U3054 );
not NOT1_8389 ( P1_R1240_U89 , P1_U3974 );
nand NAND2_8390 ( P1_R1240_U90 , P1_R1240_U305 , P1_R1240_U175 );
not NOT1_8391 ( P1_R1240_U91 , P1_U3076 );
nand NAND2_8392 ( P1_R1240_U92 , P1_R1240_U78 , P1_R1240_U314 );
nand NAND2_8393 ( P1_R1240_U93 , P1_R1240_U260 , P1_R1240_U259 );
nand NAND2_8394 ( P1_R1240_U94 , P1_R1240_U69 , P1_R1240_U336 );
nand NAND2_8395 ( P1_R1240_U95 , P1_R1240_U456 , P1_R1240_U455 );
nand NAND2_8396 ( P1_R1240_U96 , P1_R1240_U503 , P1_R1240_U502 );
nand NAND2_8397 ( P1_R1240_U97 , P1_R1240_U374 , P1_R1240_U373 );
nand NAND2_8398 ( P1_R1240_U98 , P1_R1240_U379 , P1_R1240_U378 );
nand NAND2_8399 ( P1_R1240_U99 , P1_R1240_U386 , P1_R1240_U385 );
nand NAND2_8400 ( P1_R1240_U100 , P1_R1240_U393 , P1_R1240_U392 );
nand NAND2_8401 ( P1_R1240_U101 , P1_R1240_U398 , P1_R1240_U397 );
nand NAND2_8402 ( P1_R1240_U102 , P1_R1240_U407 , P1_R1240_U406 );
nand NAND2_8403 ( P1_R1240_U103 , P1_R1240_U414 , P1_R1240_U413 );
nand NAND2_8404 ( P1_R1240_U104 , P1_R1240_U421 , P1_R1240_U420 );
nand NAND2_8405 ( P1_R1240_U105 , P1_R1240_U428 , P1_R1240_U427 );
nand NAND2_8406 ( P1_R1240_U106 , P1_R1240_U433 , P1_R1240_U432 );
nand NAND2_8407 ( P1_R1240_U107 , P1_R1240_U440 , P1_R1240_U439 );
nand NAND2_8408 ( P1_R1240_U108 , P1_R1240_U447 , P1_R1240_U446 );
nand NAND2_8409 ( P1_R1240_U109 , P1_R1240_U461 , P1_R1240_U460 );
nand NAND2_8410 ( P1_R1240_U110 , P1_R1240_U466 , P1_R1240_U465 );
nand NAND2_8411 ( P1_R1240_U111 , P1_R1240_U473 , P1_R1240_U472 );
nand NAND2_8412 ( P1_R1240_U112 , P1_R1240_U480 , P1_R1240_U479 );
nand NAND2_8413 ( P1_R1240_U113 , P1_R1240_U487 , P1_R1240_U486 );
nand NAND2_8414 ( P1_R1240_U114 , P1_R1240_U494 , P1_R1240_U493 );
nand NAND2_8415 ( P1_R1240_U115 , P1_R1240_U499 , P1_R1240_U498 );
and AND2_8416 ( P1_R1240_U116 , P1_U3458 , P1_U3068 );
and AND2_8417 ( P1_R1240_U117 , P1_R1240_U188 , P1_R1240_U186 );
and AND2_8418 ( P1_R1240_U118 , P1_R1240_U193 , P1_R1240_U191 );
and AND2_8419 ( P1_R1240_U119 , P1_R1240_U200 , P1_R1240_U199 );
and AND3_8420 ( P1_R1240_U120 , P1_R1240_U381 , P1_R1240_U380 , P1_R1240_U23 );
and AND2_8421 ( P1_R1240_U121 , P1_R1240_U211 , P1_R1240_U6 );
and AND2_8422 ( P1_R1240_U122 , P1_R1240_U219 , P1_R1240_U217 );
and AND3_8423 ( P1_R1240_U123 , P1_R1240_U388 , P1_R1240_U387 , P1_R1240_U35 );
and AND2_8424 ( P1_R1240_U124 , P1_R1240_U225 , P1_R1240_U4 );
and AND2_8425 ( P1_R1240_U125 , P1_R1240_U233 , P1_R1240_U180 );
and AND2_8426 ( P1_R1240_U126 , P1_R1240_U203 , P1_R1240_U7 );
and AND2_8427 ( P1_R1240_U127 , P1_R1240_U238 , P1_R1240_U170 );
and AND2_8428 ( P1_R1240_U128 , P1_R1240_U249 , P1_R1240_U8 );
and AND2_8429 ( P1_R1240_U129 , P1_R1240_U247 , P1_R1240_U171 );
and AND2_8430 ( P1_R1240_U130 , P1_R1240_U267 , P1_R1240_U266 );
and AND2_8431 ( P1_R1240_U131 , P1_R1240_U10 , P1_R1240_U281 );
and AND2_8432 ( P1_R1240_U132 , P1_R1240_U284 , P1_R1240_U279 );
and AND2_8433 ( P1_R1240_U133 , P1_R1240_U300 , P1_R1240_U297 );
and AND2_8434 ( P1_R1240_U134 , P1_R1240_U367 , P1_R1240_U301 );
and AND2_8435 ( P1_R1240_U135 , P1_R1240_U159 , P1_R1240_U277 );
and AND3_8436 ( P1_R1240_U136 , P1_R1240_U454 , P1_R1240_U453 , P1_R1240_U81 );
and AND3_8437 ( P1_R1240_U137 , P1_R1240_U468 , P1_R1240_U467 , P1_R1240_U60 );
and AND2_8438 ( P1_R1240_U138 , P1_R1240_U333 , P1_R1240_U9 );
and AND3_8439 ( P1_R1240_U139 , P1_R1240_U489 , P1_R1240_U488 , P1_R1240_U171 );
and AND2_8440 ( P1_R1240_U140 , P1_R1240_U342 , P1_R1240_U8 );
and AND3_8441 ( P1_R1240_U141 , P1_R1240_U501 , P1_R1240_U500 , P1_R1240_U170 );
and AND2_8442 ( P1_R1240_U142 , P1_R1240_U349 , P1_R1240_U7 );
nand NAND2_8443 ( P1_R1240_U143 , P1_R1240_U119 , P1_R1240_U201 );
nand NAND2_8444 ( P1_R1240_U144 , P1_R1240_U216 , P1_R1240_U228 );
not NOT1_8445 ( P1_R1240_U145 , P1_U3055 );
not NOT1_8446 ( P1_R1240_U146 , P1_U3985 );
and AND2_8447 ( P1_R1240_U147 , P1_R1240_U402 , P1_R1240_U401 );
nand NAND3_8448 ( P1_R1240_U148 , P1_R1240_U303 , P1_R1240_U168 , P1_R1240_U363 );
and AND2_8449 ( P1_R1240_U149 , P1_R1240_U409 , P1_R1240_U408 );
nand NAND3_8450 ( P1_R1240_U150 , P1_R1240_U369 , P1_R1240_U368 , P1_R1240_U134 );
and AND2_8451 ( P1_R1240_U151 , P1_R1240_U416 , P1_R1240_U415 );
nand NAND3_8452 ( P1_R1240_U152 , P1_R1240_U364 , P1_R1240_U298 , P1_R1240_U87 );
and AND2_8453 ( P1_R1240_U153 , P1_R1240_U423 , P1_R1240_U422 );
nand NAND2_8454 ( P1_R1240_U154 , P1_R1240_U292 , P1_R1240_U291 );
and AND2_8455 ( P1_R1240_U155 , P1_R1240_U435 , P1_R1240_U434 );
nand NAND2_8456 ( P1_R1240_U156 , P1_R1240_U288 , P1_R1240_U287 );
and AND2_8457 ( P1_R1240_U157 , P1_R1240_U442 , P1_R1240_U441 );
nand NAND2_8458 ( P1_R1240_U158 , P1_R1240_U132 , P1_R1240_U283 );
and AND2_8459 ( P1_R1240_U159 , P1_R1240_U449 , P1_R1240_U448 );
nand NAND2_8460 ( P1_R1240_U160 , P1_R1240_U44 , P1_R1240_U326 );
nand NAND2_8461 ( P1_R1240_U161 , P1_R1240_U130 , P1_R1240_U268 );
and AND2_8462 ( P1_R1240_U162 , P1_R1240_U475 , P1_R1240_U474 );
nand NAND2_8463 ( P1_R1240_U163 , P1_R1240_U256 , P1_R1240_U255 );
and AND2_8464 ( P1_R1240_U164 , P1_R1240_U482 , P1_R1240_U481 );
nand NAND2_8465 ( P1_R1240_U165 , P1_R1240_U252 , P1_R1240_U251 );
nand NAND2_8466 ( P1_R1240_U166 , P1_R1240_U242 , P1_R1240_U241 );
nand NAND2_8467 ( P1_R1240_U167 , P1_R1240_U366 , P1_R1240_U365 );
nand NAND2_8468 ( P1_R1240_U168 , P1_U3054 , P1_R1240_U150 );
not NOT1_8469 ( P1_R1240_U169 , P1_R1240_U35 );
nand NAND2_8470 ( P1_R1240_U170 , P1_U3479 , P1_U3083 );
nand NAND2_8471 ( P1_R1240_U171 , P1_U3072 , P1_U3488 );
nand NAND2_8472 ( P1_R1240_U172 , P1_U3058 , P1_U3977 );
not NOT1_8473 ( P1_R1240_U173 , P1_R1240_U69 );
not NOT1_8474 ( P1_R1240_U174 , P1_R1240_U78 );
nand NAND2_8475 ( P1_R1240_U175 , P1_U3065 , P1_U3978 );
not NOT1_8476 ( P1_R1240_U176 , P1_R1240_U62 );
or OR2_8477 ( P1_R1240_U177 , P1_U3067 , P1_U3467 );
or OR2_8478 ( P1_R1240_U178 , P1_U3060 , P1_U3464 );
or OR2_8479 ( P1_R1240_U179 , P1_U3461 , P1_U3064 );
or OR2_8480 ( P1_R1240_U180 , P1_U3458 , P1_U3068 );
not NOT1_8481 ( P1_R1240_U181 , P1_R1240_U32 );
or OR2_8482 ( P1_R1240_U182 , P1_U3455 , P1_U3078 );
not NOT1_8483 ( P1_R1240_U183 , P1_R1240_U43 );
not NOT1_8484 ( P1_R1240_U184 , P1_R1240_U44 );
nand NAND2_8485 ( P1_R1240_U185 , P1_R1240_U43 , P1_R1240_U44 );
nand NAND2_8486 ( P1_R1240_U186 , P1_R1240_U116 , P1_R1240_U179 );
nand NAND2_8487 ( P1_R1240_U187 , P1_R1240_U5 , P1_R1240_U185 );
nand NAND2_8488 ( P1_R1240_U188 , P1_U3064 , P1_U3461 );
nand NAND2_8489 ( P1_R1240_U189 , P1_R1240_U117 , P1_R1240_U187 );
nand NAND2_8490 ( P1_R1240_U190 , P1_R1240_U36 , P1_R1240_U35 );
nand NAND2_8491 ( P1_R1240_U191 , P1_U3067 , P1_R1240_U190 );
nand NAND2_8492 ( P1_R1240_U192 , P1_R1240_U4 , P1_R1240_U189 );
nand NAND2_8493 ( P1_R1240_U193 , P1_U3467 , P1_R1240_U169 );
not NOT1_8494 ( P1_R1240_U194 , P1_R1240_U42 );
or OR2_8495 ( P1_R1240_U195 , P1_U3070 , P1_U3473 );
or OR2_8496 ( P1_R1240_U196 , P1_U3071 , P1_U3470 );
not NOT1_8497 ( P1_R1240_U197 , P1_R1240_U23 );
nand NAND2_8498 ( P1_R1240_U198 , P1_R1240_U24 , P1_R1240_U23 );
nand NAND2_8499 ( P1_R1240_U199 , P1_U3070 , P1_R1240_U198 );
nand NAND2_8500 ( P1_R1240_U200 , P1_U3473 , P1_R1240_U197 );
nand NAND2_8501 ( P1_R1240_U201 , P1_R1240_U6 , P1_R1240_U42 );
not NOT1_8502 ( P1_R1240_U202 , P1_R1240_U143 );
or OR2_8503 ( P1_R1240_U203 , P1_U3476 , P1_U3084 );
nand NAND2_8504 ( P1_R1240_U204 , P1_R1240_U203 , P1_R1240_U143 );
not NOT1_8505 ( P1_R1240_U205 , P1_R1240_U41 );
or OR2_8506 ( P1_R1240_U206 , P1_U3083 , P1_U3479 );
or OR2_8507 ( P1_R1240_U207 , P1_U3470 , P1_U3071 );
nand NAND2_8508 ( P1_R1240_U208 , P1_R1240_U207 , P1_R1240_U42 );
nand NAND2_8509 ( P1_R1240_U209 , P1_R1240_U120 , P1_R1240_U208 );
nand NAND2_8510 ( P1_R1240_U210 , P1_R1240_U194 , P1_R1240_U23 );
nand NAND2_8511 ( P1_R1240_U211 , P1_U3473 , P1_U3070 );
nand NAND2_8512 ( P1_R1240_U212 , P1_R1240_U121 , P1_R1240_U210 );
or OR2_8513 ( P1_R1240_U213 , P1_U3071 , P1_U3470 );
nand NAND2_8514 ( P1_R1240_U214 , P1_R1240_U184 , P1_R1240_U180 );
nand NAND2_8515 ( P1_R1240_U215 , P1_U3068 , P1_U3458 );
not NOT1_8516 ( P1_R1240_U216 , P1_R1240_U46 );
nand NAND2_8517 ( P1_R1240_U217 , P1_R1240_U183 , P1_R1240_U5 );
nand NAND2_8518 ( P1_R1240_U218 , P1_R1240_U46 , P1_R1240_U179 );
nand NAND2_8519 ( P1_R1240_U219 , P1_U3064 , P1_U3461 );
not NOT1_8520 ( P1_R1240_U220 , P1_R1240_U45 );
or OR2_8521 ( P1_R1240_U221 , P1_U3464 , P1_U3060 );
nand NAND2_8522 ( P1_R1240_U222 , P1_R1240_U221 , P1_R1240_U45 );
nand NAND2_8523 ( P1_R1240_U223 , P1_R1240_U123 , P1_R1240_U222 );
nand NAND2_8524 ( P1_R1240_U224 , P1_R1240_U220 , P1_R1240_U35 );
nand NAND2_8525 ( P1_R1240_U225 , P1_U3467 , P1_U3067 );
nand NAND2_8526 ( P1_R1240_U226 , P1_R1240_U124 , P1_R1240_U224 );
or OR2_8527 ( P1_R1240_U227 , P1_U3060 , P1_U3464 );
nand NAND2_8528 ( P1_R1240_U228 , P1_R1240_U183 , P1_R1240_U180 );
not NOT1_8529 ( P1_R1240_U229 , P1_R1240_U144 );
nand NAND2_8530 ( P1_R1240_U230 , P1_U3064 , P1_U3461 );
nand NAND4_8531 ( P1_R1240_U231 , P1_R1240_U400 , P1_R1240_U399 , P1_R1240_U44 , P1_R1240_U43 );
nand NAND2_8532 ( P1_R1240_U232 , P1_R1240_U44 , P1_R1240_U43 );
nand NAND2_8533 ( P1_R1240_U233 , P1_U3068 , P1_U3458 );
nand NAND2_8534 ( P1_R1240_U234 , P1_R1240_U125 , P1_R1240_U232 );
or OR2_8535 ( P1_R1240_U235 , P1_U3083 , P1_U3479 );
or OR2_8536 ( P1_R1240_U236 , P1_U3062 , P1_U3482 );
nand NAND2_8537 ( P1_R1240_U237 , P1_R1240_U176 , P1_R1240_U7 );
nand NAND2_8538 ( P1_R1240_U238 , P1_U3062 , P1_U3482 );
nand NAND2_8539 ( P1_R1240_U239 , P1_R1240_U127 , P1_R1240_U237 );
or OR2_8540 ( P1_R1240_U240 , P1_U3482 , P1_U3062 );
nand NAND2_8541 ( P1_R1240_U241 , P1_R1240_U126 , P1_R1240_U143 );
nand NAND2_8542 ( P1_R1240_U242 , P1_R1240_U240 , P1_R1240_U239 );
not NOT1_8543 ( P1_R1240_U243 , P1_R1240_U166 );
or OR2_8544 ( P1_R1240_U244 , P1_U3080 , P1_U3491 );
or OR2_8545 ( P1_R1240_U245 , P1_U3072 , P1_U3488 );
nand NAND2_8546 ( P1_R1240_U246 , P1_R1240_U173 , P1_R1240_U8 );
nand NAND2_8547 ( P1_R1240_U247 , P1_U3080 , P1_U3491 );
nand NAND2_8548 ( P1_R1240_U248 , P1_R1240_U129 , P1_R1240_U246 );
or OR2_8549 ( P1_R1240_U249 , P1_U3485 , P1_U3063 );
or OR2_8550 ( P1_R1240_U250 , P1_U3491 , P1_U3080 );
nand NAND2_8551 ( P1_R1240_U251 , P1_R1240_U128 , P1_R1240_U166 );
nand NAND2_8552 ( P1_R1240_U252 , P1_R1240_U250 , P1_R1240_U248 );
not NOT1_8553 ( P1_R1240_U253 , P1_R1240_U165 );
or OR2_8554 ( P1_R1240_U254 , P1_U3494 , P1_U3079 );
nand NAND2_8555 ( P1_R1240_U255 , P1_R1240_U254 , P1_R1240_U165 );
nand NAND2_8556 ( P1_R1240_U256 , P1_U3079 , P1_U3494 );
not NOT1_8557 ( P1_R1240_U257 , P1_R1240_U163 );
or OR2_8558 ( P1_R1240_U258 , P1_U3497 , P1_U3074 );
nand NAND2_8559 ( P1_R1240_U259 , P1_R1240_U258 , P1_R1240_U163 );
nand NAND2_8560 ( P1_R1240_U260 , P1_U3074 , P1_U3497 );
not NOT1_8561 ( P1_R1240_U261 , P1_R1240_U93 );
or OR2_8562 ( P1_R1240_U262 , P1_U3069 , P1_U3503 );
or OR2_8563 ( P1_R1240_U263 , P1_U3073 , P1_U3500 );
not NOT1_8564 ( P1_R1240_U264 , P1_R1240_U60 );
nand NAND2_8565 ( P1_R1240_U265 , P1_R1240_U61 , P1_R1240_U60 );
nand NAND2_8566 ( P1_R1240_U266 , P1_U3069 , P1_R1240_U265 );
nand NAND2_8567 ( P1_R1240_U267 , P1_U3503 , P1_R1240_U264 );
nand NAND2_8568 ( P1_R1240_U268 , P1_R1240_U9 , P1_R1240_U93 );
not NOT1_8569 ( P1_R1240_U269 , P1_R1240_U161 );
or OR2_8570 ( P1_R1240_U270 , P1_U3076 , P1_U3982 );
or OR2_8571 ( P1_R1240_U271 , P1_U3081 , P1_U3508 );
or OR2_8572 ( P1_R1240_U272 , P1_U3075 , P1_U3981 );
not NOT1_8573 ( P1_R1240_U273 , P1_R1240_U81 );
nand NAND2_8574 ( P1_R1240_U274 , P1_U3982 , P1_R1240_U273 );
nand NAND2_8575 ( P1_R1240_U275 , P1_R1240_U274 , P1_R1240_U91 );
nand NAND2_8576 ( P1_R1240_U276 , P1_R1240_U81 , P1_R1240_U82 );
nand NAND2_8577 ( P1_R1240_U277 , P1_R1240_U276 , P1_R1240_U275 );
nand NAND2_8578 ( P1_R1240_U278 , P1_R1240_U174 , P1_R1240_U10 );
nand NAND2_8579 ( P1_R1240_U279 , P1_U3075 , P1_U3981 );
nand NAND2_8580 ( P1_R1240_U280 , P1_R1240_U277 , P1_R1240_U278 );
or OR2_8581 ( P1_R1240_U281 , P1_U3506 , P1_U3082 );
or OR2_8582 ( P1_R1240_U282 , P1_U3981 , P1_U3075 );
nand NAND3_8583 ( P1_R1240_U283 , P1_R1240_U272 , P1_R1240_U161 , P1_R1240_U131 );
nand NAND2_8584 ( P1_R1240_U284 , P1_R1240_U282 , P1_R1240_U280 );
not NOT1_8585 ( P1_R1240_U285 , P1_R1240_U158 );
or OR2_8586 ( P1_R1240_U286 , P1_U3980 , P1_U3061 );
nand NAND2_8587 ( P1_R1240_U287 , P1_R1240_U286 , P1_R1240_U158 );
nand NAND2_8588 ( P1_R1240_U288 , P1_U3061 , P1_U3980 );
not NOT1_8589 ( P1_R1240_U289 , P1_R1240_U156 );
or OR2_8590 ( P1_R1240_U290 , P1_U3979 , P1_U3066 );
nand NAND2_8591 ( P1_R1240_U291 , P1_R1240_U290 , P1_R1240_U156 );
nand NAND2_8592 ( P1_R1240_U292 , P1_U3066 , P1_U3979 );
not NOT1_8593 ( P1_R1240_U293 , P1_R1240_U154 );
or OR2_8594 ( P1_R1240_U294 , P1_U3058 , P1_U3977 );
nand NAND2_8595 ( P1_R1240_U295 , P1_R1240_U175 , P1_R1240_U172 );
not NOT1_8596 ( P1_R1240_U296 , P1_R1240_U87 );
or OR2_8597 ( P1_R1240_U297 , P1_U3978 , P1_U3065 );
nand NAND3_8598 ( P1_R1240_U298 , P1_R1240_U154 , P1_R1240_U297 , P1_R1240_U167 );
not NOT1_8599 ( P1_R1240_U299 , P1_R1240_U152 );
or OR2_8600 ( P1_R1240_U300 , P1_U3975 , P1_U3053 );
nand NAND2_8601 ( P1_R1240_U301 , P1_U3053 , P1_U3975 );
not NOT1_8602 ( P1_R1240_U302 , P1_R1240_U150 );
nand NAND2_8603 ( P1_R1240_U303 , P1_U3974 , P1_R1240_U150 );
not NOT1_8604 ( P1_R1240_U304 , P1_R1240_U148 );
nand NAND2_8605 ( P1_R1240_U305 , P1_R1240_U297 , P1_R1240_U154 );
not NOT1_8606 ( P1_R1240_U306 , P1_R1240_U90 );
or OR2_8607 ( P1_R1240_U307 , P1_U3977 , P1_U3058 );
nand NAND2_8608 ( P1_R1240_U308 , P1_R1240_U307 , P1_R1240_U90 );
nand NAND3_8609 ( P1_R1240_U309 , P1_R1240_U308 , P1_R1240_U172 , P1_R1240_U153 );
nand NAND2_8610 ( P1_R1240_U310 , P1_R1240_U306 , P1_R1240_U172 );
nand NAND2_8611 ( P1_R1240_U311 , P1_U3976 , P1_U3057 );
nand NAND3_8612 ( P1_R1240_U312 , P1_R1240_U310 , P1_R1240_U311 , P1_R1240_U167 );
or OR2_8613 ( P1_R1240_U313 , P1_U3058 , P1_U3977 );
nand NAND2_8614 ( P1_R1240_U314 , P1_R1240_U281 , P1_R1240_U161 );
not NOT1_8615 ( P1_R1240_U315 , P1_R1240_U92 );
nand NAND2_8616 ( P1_R1240_U316 , P1_R1240_U10 , P1_R1240_U92 );
nand NAND2_8617 ( P1_R1240_U317 , P1_R1240_U135 , P1_R1240_U316 );
nand NAND2_8618 ( P1_R1240_U318 , P1_R1240_U316 , P1_R1240_U277 );
nand NAND2_8619 ( P1_R1240_U319 , P1_R1240_U452 , P1_R1240_U318 );
or OR2_8620 ( P1_R1240_U320 , P1_U3508 , P1_U3081 );
nand NAND2_8621 ( P1_R1240_U321 , P1_R1240_U320 , P1_R1240_U92 );
nand NAND2_8622 ( P1_R1240_U322 , P1_R1240_U136 , P1_R1240_U321 );
nand NAND2_8623 ( P1_R1240_U323 , P1_R1240_U315 , P1_R1240_U81 );
nand NAND2_8624 ( P1_R1240_U324 , P1_U3076 , P1_U3982 );
nand NAND3_8625 ( P1_R1240_U325 , P1_R1240_U324 , P1_R1240_U323 , P1_R1240_U10 );
or OR2_8626 ( P1_R1240_U326 , P1_U3455 , P1_U3078 );
not NOT1_8627 ( P1_R1240_U327 , P1_R1240_U160 );
or OR2_8628 ( P1_R1240_U328 , P1_U3081 , P1_U3508 );
or OR2_8629 ( P1_R1240_U329 , P1_U3500 , P1_U3073 );
nand NAND2_8630 ( P1_R1240_U330 , P1_R1240_U329 , P1_R1240_U93 );
nand NAND2_8631 ( P1_R1240_U331 , P1_R1240_U137 , P1_R1240_U330 );
nand NAND2_8632 ( P1_R1240_U332 , P1_R1240_U261 , P1_R1240_U60 );
nand NAND2_8633 ( P1_R1240_U333 , P1_U3503 , P1_U3069 );
nand NAND2_8634 ( P1_R1240_U334 , P1_R1240_U138 , P1_R1240_U332 );
or OR2_8635 ( P1_R1240_U335 , P1_U3073 , P1_U3500 );
nand NAND2_8636 ( P1_R1240_U336 , P1_R1240_U249 , P1_R1240_U166 );
not NOT1_8637 ( P1_R1240_U337 , P1_R1240_U94 );
or OR2_8638 ( P1_R1240_U338 , P1_U3488 , P1_U3072 );
nand NAND2_8639 ( P1_R1240_U339 , P1_R1240_U338 , P1_R1240_U94 );
nand NAND2_8640 ( P1_R1240_U340 , P1_R1240_U139 , P1_R1240_U339 );
nand NAND2_8641 ( P1_R1240_U341 , P1_R1240_U337 , P1_R1240_U171 );
nand NAND2_8642 ( P1_R1240_U342 , P1_U3080 , P1_U3491 );
nand NAND2_8643 ( P1_R1240_U343 , P1_R1240_U140 , P1_R1240_U341 );
or OR2_8644 ( P1_R1240_U344 , P1_U3072 , P1_U3488 );
or OR2_8645 ( P1_R1240_U345 , P1_U3479 , P1_U3083 );
nand NAND2_8646 ( P1_R1240_U346 , P1_R1240_U345 , P1_R1240_U41 );
nand NAND2_8647 ( P1_R1240_U347 , P1_R1240_U141 , P1_R1240_U346 );
nand NAND2_8648 ( P1_R1240_U348 , P1_R1240_U205 , P1_R1240_U170 );
nand NAND2_8649 ( P1_R1240_U349 , P1_U3062 , P1_U3482 );
nand NAND2_8650 ( P1_R1240_U350 , P1_R1240_U142 , P1_R1240_U348 );
nand NAND2_8651 ( P1_R1240_U351 , P1_R1240_U206 , P1_R1240_U170 );
nand NAND2_8652 ( P1_R1240_U352 , P1_R1240_U203 , P1_R1240_U62 );
nand NAND2_8653 ( P1_R1240_U353 , P1_R1240_U213 , P1_R1240_U23 );
nand NAND2_8654 ( P1_R1240_U354 , P1_R1240_U227 , P1_R1240_U35 );
nand NAND2_8655 ( P1_R1240_U355 , P1_R1240_U230 , P1_R1240_U179 );
nand NAND2_8656 ( P1_R1240_U356 , P1_R1240_U313 , P1_R1240_U172 );
nand NAND2_8657 ( P1_R1240_U357 , P1_R1240_U297 , P1_R1240_U175 );
nand NAND2_8658 ( P1_R1240_U358 , P1_R1240_U328 , P1_R1240_U81 );
nand NAND2_8659 ( P1_R1240_U359 , P1_R1240_U281 , P1_R1240_U78 );
nand NAND2_8660 ( P1_R1240_U360 , P1_R1240_U335 , P1_R1240_U60 );
nand NAND2_8661 ( P1_R1240_U361 , P1_R1240_U344 , P1_R1240_U171 );
nand NAND2_8662 ( P1_R1240_U362 , P1_R1240_U249 , P1_R1240_U69 );
nand NAND2_8663 ( P1_R1240_U363 , P1_U3974 , P1_U3054 );
nand NAND2_8664 ( P1_R1240_U364 , P1_R1240_U295 , P1_R1240_U167 );
nand NAND2_8665 ( P1_R1240_U365 , P1_U3057 , P1_R1240_U294 );
nand NAND2_8666 ( P1_R1240_U366 , P1_U3976 , P1_R1240_U294 );
nand NAND3_8667 ( P1_R1240_U367 , P1_R1240_U295 , P1_R1240_U167 , P1_R1240_U300 );
nand NAND3_8668 ( P1_R1240_U368 , P1_R1240_U154 , P1_R1240_U167 , P1_R1240_U133 );
nand NAND2_8669 ( P1_R1240_U369 , P1_R1240_U296 , P1_R1240_U300 );
nand NAND2_8670 ( P1_R1240_U370 , P1_U3083 , P1_R1240_U40 );
nand NAND2_8671 ( P1_R1240_U371 , P1_U3479 , P1_R1240_U39 );
nand NAND2_8672 ( P1_R1240_U372 , P1_R1240_U371 , P1_R1240_U370 );
nand NAND2_8673 ( P1_R1240_U373 , P1_R1240_U351 , P1_R1240_U41 );
nand NAND2_8674 ( P1_R1240_U374 , P1_R1240_U372 , P1_R1240_U205 );
nand NAND2_8675 ( P1_R1240_U375 , P1_U3084 , P1_R1240_U37 );
nand NAND2_8676 ( P1_R1240_U376 , P1_U3476 , P1_R1240_U38 );
nand NAND2_8677 ( P1_R1240_U377 , P1_R1240_U376 , P1_R1240_U375 );
nand NAND2_8678 ( P1_R1240_U378 , P1_R1240_U352 , P1_R1240_U143 );
nand NAND2_8679 ( P1_R1240_U379 , P1_R1240_U202 , P1_R1240_U377 );
nand NAND2_8680 ( P1_R1240_U380 , P1_U3070 , P1_R1240_U24 );
nand NAND2_8681 ( P1_R1240_U381 , P1_U3473 , P1_R1240_U22 );
nand NAND2_8682 ( P1_R1240_U382 , P1_U3071 , P1_R1240_U20 );
nand NAND2_8683 ( P1_R1240_U383 , P1_U3470 , P1_R1240_U21 );
nand NAND2_8684 ( P1_R1240_U384 , P1_R1240_U383 , P1_R1240_U382 );
nand NAND2_8685 ( P1_R1240_U385 , P1_R1240_U353 , P1_R1240_U42 );
nand NAND2_8686 ( P1_R1240_U386 , P1_R1240_U384 , P1_R1240_U194 );
nand NAND2_8687 ( P1_R1240_U387 , P1_U3067 , P1_R1240_U36 );
nand NAND2_8688 ( P1_R1240_U388 , P1_U3467 , P1_R1240_U27 );
nand NAND2_8689 ( P1_R1240_U389 , P1_U3060 , P1_R1240_U25 );
nand NAND2_8690 ( P1_R1240_U390 , P1_U3464 , P1_R1240_U26 );
nand NAND2_8691 ( P1_R1240_U391 , P1_R1240_U390 , P1_R1240_U389 );
nand NAND2_8692 ( P1_R1240_U392 , P1_R1240_U354 , P1_R1240_U45 );
nand NAND2_8693 ( P1_R1240_U393 , P1_R1240_U391 , P1_R1240_U220 );
nand NAND2_8694 ( P1_R1240_U394 , P1_U3064 , P1_R1240_U33 );
nand NAND2_8695 ( P1_R1240_U395 , P1_U3461 , P1_R1240_U34 );
nand NAND2_8696 ( P1_R1240_U396 , P1_R1240_U395 , P1_R1240_U394 );
nand NAND2_8697 ( P1_R1240_U397 , P1_R1240_U355 , P1_R1240_U144 );
nand NAND2_8698 ( P1_R1240_U398 , P1_R1240_U229 , P1_R1240_U396 );
nand NAND2_8699 ( P1_R1240_U399 , P1_U3068 , P1_R1240_U28 );
nand NAND2_8700 ( P1_R1240_U400 , P1_U3458 , P1_R1240_U29 );
nand NAND2_8701 ( P1_R1240_U401 , P1_U3055 , P1_R1240_U146 );
nand NAND2_8702 ( P1_R1240_U402 , P1_U3985 , P1_R1240_U145 );
nand NAND2_8703 ( P1_R1240_U403 , P1_U3055 , P1_R1240_U146 );
nand NAND2_8704 ( P1_R1240_U404 , P1_U3985 , P1_R1240_U145 );
nand NAND2_8705 ( P1_R1240_U405 , P1_R1240_U404 , P1_R1240_U403 );
nand NAND2_8706 ( P1_R1240_U406 , P1_R1240_U147 , P1_R1240_U148 );
nand NAND2_8707 ( P1_R1240_U407 , P1_R1240_U304 , P1_R1240_U405 );
nand NAND2_8708 ( P1_R1240_U408 , P1_U3054 , P1_R1240_U89 );
nand NAND2_8709 ( P1_R1240_U409 , P1_U3974 , P1_R1240_U88 );
nand NAND2_8710 ( P1_R1240_U410 , P1_U3054 , P1_R1240_U89 );
nand NAND2_8711 ( P1_R1240_U411 , P1_U3974 , P1_R1240_U88 );
nand NAND2_8712 ( P1_R1240_U412 , P1_R1240_U411 , P1_R1240_U410 );
nand NAND2_8713 ( P1_R1240_U413 , P1_R1240_U149 , P1_R1240_U150 );
nand NAND2_8714 ( P1_R1240_U414 , P1_R1240_U302 , P1_R1240_U412 );
nand NAND2_8715 ( P1_R1240_U415 , P1_U3053 , P1_R1240_U47 );
nand NAND2_8716 ( P1_R1240_U416 , P1_U3975 , P1_R1240_U48 );
nand NAND2_8717 ( P1_R1240_U417 , P1_U3053 , P1_R1240_U47 );
nand NAND2_8718 ( P1_R1240_U418 , P1_U3975 , P1_R1240_U48 );
nand NAND2_8719 ( P1_R1240_U419 , P1_R1240_U418 , P1_R1240_U417 );
nand NAND2_8720 ( P1_R1240_U420 , P1_R1240_U151 , P1_R1240_U152 );
nand NAND2_8721 ( P1_R1240_U421 , P1_R1240_U299 , P1_R1240_U419 );
nand NAND2_8722 ( P1_R1240_U422 , P1_U3057 , P1_R1240_U50 );
nand NAND2_8723 ( P1_R1240_U423 , P1_U3976 , P1_R1240_U49 );
nand NAND2_8724 ( P1_R1240_U424 , P1_U3058 , P1_R1240_U51 );
nand NAND2_8725 ( P1_R1240_U425 , P1_U3977 , P1_R1240_U52 );
nand NAND2_8726 ( P1_R1240_U426 , P1_R1240_U425 , P1_R1240_U424 );
nand NAND2_8727 ( P1_R1240_U427 , P1_R1240_U356 , P1_R1240_U90 );
nand NAND2_8728 ( P1_R1240_U428 , P1_R1240_U426 , P1_R1240_U306 );
nand NAND2_8729 ( P1_R1240_U429 , P1_U3065 , P1_R1240_U53 );
nand NAND2_8730 ( P1_R1240_U430 , P1_U3978 , P1_R1240_U54 );
nand NAND2_8731 ( P1_R1240_U431 , P1_R1240_U430 , P1_R1240_U429 );
nand NAND2_8732 ( P1_R1240_U432 , P1_R1240_U357 , P1_R1240_U154 );
nand NAND2_8733 ( P1_R1240_U433 , P1_R1240_U293 , P1_R1240_U431 );
nand NAND2_8734 ( P1_R1240_U434 , P1_U3066 , P1_R1240_U85 );
nand NAND2_8735 ( P1_R1240_U435 , P1_U3979 , P1_R1240_U86 );
nand NAND2_8736 ( P1_R1240_U436 , P1_U3066 , P1_R1240_U85 );
nand NAND2_8737 ( P1_R1240_U437 , P1_U3979 , P1_R1240_U86 );
nand NAND2_8738 ( P1_R1240_U438 , P1_R1240_U437 , P1_R1240_U436 );
nand NAND2_8739 ( P1_R1240_U439 , P1_R1240_U155 , P1_R1240_U156 );
nand NAND2_8740 ( P1_R1240_U440 , P1_R1240_U289 , P1_R1240_U438 );
nand NAND2_8741 ( P1_R1240_U441 , P1_U3061 , P1_R1240_U83 );
nand NAND2_8742 ( P1_R1240_U442 , P1_U3980 , P1_R1240_U84 );
nand NAND2_8743 ( P1_R1240_U443 , P1_U3061 , P1_R1240_U83 );
nand NAND2_8744 ( P1_R1240_U444 , P1_U3980 , P1_R1240_U84 );
nand NAND2_8745 ( P1_R1240_U445 , P1_R1240_U444 , P1_R1240_U443 );
nand NAND2_8746 ( P1_R1240_U446 , P1_R1240_U157 , P1_R1240_U158 );
nand NAND2_8747 ( P1_R1240_U447 , P1_R1240_U285 , P1_R1240_U445 );
nand NAND2_8748 ( P1_R1240_U448 , P1_U3075 , P1_R1240_U55 );
nand NAND2_8749 ( P1_R1240_U449 , P1_U3981 , P1_R1240_U56 );
nand NAND2_8750 ( P1_R1240_U450 , P1_U3075 , P1_R1240_U55 );
nand NAND2_8751 ( P1_R1240_U451 , P1_U3981 , P1_R1240_U56 );
nand NAND2_8752 ( P1_R1240_U452 , P1_R1240_U451 , P1_R1240_U450 );
nand NAND2_8753 ( P1_R1240_U453 , P1_U3076 , P1_R1240_U82 );
nand NAND2_8754 ( P1_R1240_U454 , P1_U3982 , P1_R1240_U91 );
nand NAND2_8755 ( P1_R1240_U455 , P1_R1240_U181 , P1_R1240_U160 );
nand NAND2_8756 ( P1_R1240_U456 , P1_R1240_U327 , P1_R1240_U32 );
nand NAND2_8757 ( P1_R1240_U457 , P1_U3081 , P1_R1240_U79 );
nand NAND2_8758 ( P1_R1240_U458 , P1_U3508 , P1_R1240_U80 );
nand NAND2_8759 ( P1_R1240_U459 , P1_R1240_U458 , P1_R1240_U457 );
nand NAND2_8760 ( P1_R1240_U460 , P1_R1240_U358 , P1_R1240_U92 );
nand NAND2_8761 ( P1_R1240_U461 , P1_R1240_U459 , P1_R1240_U315 );
nand NAND2_8762 ( P1_R1240_U462 , P1_U3082 , P1_R1240_U76 );
nand NAND2_8763 ( P1_R1240_U463 , P1_U3506 , P1_R1240_U77 );
nand NAND2_8764 ( P1_R1240_U464 , P1_R1240_U463 , P1_R1240_U462 );
nand NAND2_8765 ( P1_R1240_U465 , P1_R1240_U359 , P1_R1240_U161 );
nand NAND2_8766 ( P1_R1240_U466 , P1_R1240_U269 , P1_R1240_U464 );
nand NAND2_8767 ( P1_R1240_U467 , P1_U3069 , P1_R1240_U61 );
nand NAND2_8768 ( P1_R1240_U468 , P1_U3503 , P1_R1240_U59 );
nand NAND2_8769 ( P1_R1240_U469 , P1_U3073 , P1_R1240_U57 );
nand NAND2_8770 ( P1_R1240_U470 , P1_U3500 , P1_R1240_U58 );
nand NAND2_8771 ( P1_R1240_U471 , P1_R1240_U470 , P1_R1240_U469 );
nand NAND2_8772 ( P1_R1240_U472 , P1_R1240_U360 , P1_R1240_U93 );
nand NAND2_8773 ( P1_R1240_U473 , P1_R1240_U471 , P1_R1240_U261 );
nand NAND2_8774 ( P1_R1240_U474 , P1_U3074 , P1_R1240_U74 );
nand NAND2_8775 ( P1_R1240_U475 , P1_U3497 , P1_R1240_U75 );
nand NAND2_8776 ( P1_R1240_U476 , P1_U3074 , P1_R1240_U74 );
nand NAND2_8777 ( P1_R1240_U477 , P1_U3497 , P1_R1240_U75 );
nand NAND2_8778 ( P1_R1240_U478 , P1_R1240_U477 , P1_R1240_U476 );
nand NAND2_8779 ( P1_R1240_U479 , P1_R1240_U162 , P1_R1240_U163 );
nand NAND2_8780 ( P1_R1240_U480 , P1_R1240_U257 , P1_R1240_U478 );
nand NAND2_8781 ( P1_R1240_U481 , P1_U3079 , P1_R1240_U72 );
nand NAND2_8782 ( P1_R1240_U482 , P1_U3494 , P1_R1240_U73 );
nand NAND2_8783 ( P1_R1240_U483 , P1_U3079 , P1_R1240_U72 );
nand NAND2_8784 ( P1_R1240_U484 , P1_U3494 , P1_R1240_U73 );
nand NAND2_8785 ( P1_R1240_U485 , P1_R1240_U484 , P1_R1240_U483 );
nand NAND2_8786 ( P1_R1240_U486 , P1_R1240_U164 , P1_R1240_U165 );
nand NAND2_8787 ( P1_R1240_U487 , P1_R1240_U253 , P1_R1240_U485 );
nand NAND2_8788 ( P1_R1240_U488 , P1_U3080 , P1_R1240_U70 );
nand NAND2_8789 ( P1_R1240_U489 , P1_U3491 , P1_R1240_U71 );
nand NAND2_8790 ( P1_R1240_U490 , P1_U3072 , P1_R1240_U65 );
nand NAND2_8791 ( P1_R1240_U491 , P1_U3488 , P1_R1240_U66 );
nand NAND2_8792 ( P1_R1240_U492 , P1_R1240_U491 , P1_R1240_U490 );
nand NAND2_8793 ( P1_R1240_U493 , P1_R1240_U361 , P1_R1240_U94 );
nand NAND2_8794 ( P1_R1240_U494 , P1_R1240_U492 , P1_R1240_U337 );
nand NAND2_8795 ( P1_R1240_U495 , P1_U3063 , P1_R1240_U67 );
nand NAND2_8796 ( P1_R1240_U496 , P1_U3485 , P1_R1240_U68 );
nand NAND2_8797 ( P1_R1240_U497 , P1_R1240_U496 , P1_R1240_U495 );
nand NAND2_8798 ( P1_R1240_U498 , P1_R1240_U362 , P1_R1240_U166 );
nand NAND2_8799 ( P1_R1240_U499 , P1_R1240_U243 , P1_R1240_U497 );
nand NAND2_8800 ( P1_R1240_U500 , P1_U3062 , P1_R1240_U63 );
nand NAND2_8801 ( P1_R1240_U501 , P1_U3482 , P1_R1240_U64 );
nand NAND2_8802 ( P1_R1240_U502 , P1_U3077 , P1_R1240_U30 );
nand NAND2_8803 ( P1_R1240_U503 , P1_U3450 , P1_R1240_U31 );
and AND2_8804 ( P1_R1162_U4 , P1_R1162_U95 , P1_R1162_U94 );
and AND2_8805 ( P1_R1162_U5 , P1_R1162_U96 , P1_R1162_U97 );
and AND2_8806 ( P1_R1162_U6 , P1_R1162_U113 , P1_R1162_U112 );
and AND2_8807 ( P1_R1162_U7 , P1_R1162_U155 , P1_R1162_U154 );
and AND2_8808 ( P1_R1162_U8 , P1_R1162_U164 , P1_R1162_U163 );
and AND2_8809 ( P1_R1162_U9 , P1_R1162_U182 , P1_R1162_U181 );
and AND2_8810 ( P1_R1162_U10 , P1_R1162_U218 , P1_R1162_U215 );
and AND2_8811 ( P1_R1162_U11 , P1_R1162_U211 , P1_R1162_U208 );
and AND2_8812 ( P1_R1162_U12 , P1_R1162_U202 , P1_R1162_U199 );
and AND2_8813 ( P1_R1162_U13 , P1_R1162_U196 , P1_R1162_U192 );
and AND2_8814 ( P1_R1162_U14 , P1_R1162_U151 , P1_R1162_U148 );
and AND2_8815 ( P1_R1162_U15 , P1_R1162_U143 , P1_R1162_U140 );
and AND2_8816 ( P1_R1162_U16 , P1_R1162_U129 , P1_R1162_U126 );
not NOT1_8817 ( P1_R1162_U17 , P1_REG1_REG_6_ );
not NOT1_8818 ( P1_R1162_U18 , P1_U3469 );
not NOT1_8819 ( P1_R1162_U19 , P1_U3472 );
nand NAND2_8820 ( P1_R1162_U20 , P1_U3469 , P1_REG1_REG_6_ );
not NOT1_8821 ( P1_R1162_U21 , P1_REG1_REG_7_ );
not NOT1_8822 ( P1_R1162_U22 , P1_REG1_REG_4_ );
not NOT1_8823 ( P1_R1162_U23 , P1_U3463 );
not NOT1_8824 ( P1_R1162_U24 , P1_U3466 );
not NOT1_8825 ( P1_R1162_U25 , P1_REG1_REG_2_ );
not NOT1_8826 ( P1_R1162_U26 , P1_U3457 );
not NOT1_8827 ( P1_R1162_U27 , P1_REG1_REG_0_ );
not NOT1_8828 ( P1_R1162_U28 , P1_U3448 );
nand NAND2_8829 ( P1_R1162_U29 , P1_U3448 , P1_REG1_REG_0_ );
not NOT1_8830 ( P1_R1162_U30 , P1_REG1_REG_3_ );
not NOT1_8831 ( P1_R1162_U31 , P1_U3460 );
nand NAND2_8832 ( P1_R1162_U32 , P1_U3463 , P1_REG1_REG_4_ );
not NOT1_8833 ( P1_R1162_U33 , P1_REG1_REG_5_ );
not NOT1_8834 ( P1_R1162_U34 , P1_REG1_REG_8_ );
not NOT1_8835 ( P1_R1162_U35 , P1_U3475 );
not NOT1_8836 ( P1_R1162_U36 , P1_U3478 );
not NOT1_8837 ( P1_R1162_U37 , P1_REG1_REG_9_ );
nand NAND2_8838 ( P1_R1162_U38 , P1_R1162_U49 , P1_R1162_U121 );
nand NAND3_8839 ( P1_R1162_U39 , P1_R1162_U110 , P1_R1162_U108 , P1_R1162_U109 );
nand NAND2_8840 ( P1_R1162_U40 , P1_R1162_U98 , P1_R1162_U99 );
nand NAND2_8841 ( P1_R1162_U41 , P1_REG1_REG_1_ , P1_U3454 );
nand NAND3_8842 ( P1_R1162_U42 , P1_R1162_U136 , P1_R1162_U134 , P1_R1162_U135 );
nand NAND2_8843 ( P1_R1162_U43 , P1_R1162_U132 , P1_R1162_U131 );
not NOT1_8844 ( P1_R1162_U44 , P1_REG1_REG_16_ );
not NOT1_8845 ( P1_R1162_U45 , P1_U3499 );
not NOT1_8846 ( P1_R1162_U46 , P1_U3502 );
nand NAND2_8847 ( P1_R1162_U47 , P1_U3499 , P1_REG1_REG_16_ );
not NOT1_8848 ( P1_R1162_U48 , P1_REG1_REG_17_ );
nand NAND2_8849 ( P1_R1162_U49 , P1_U3475 , P1_REG1_REG_8_ );
not NOT1_8850 ( P1_R1162_U50 , P1_REG1_REG_10_ );
not NOT1_8851 ( P1_R1162_U51 , P1_U3481 );
not NOT1_8852 ( P1_R1162_U52 , P1_REG1_REG_12_ );
not NOT1_8853 ( P1_R1162_U53 , P1_U3487 );
not NOT1_8854 ( P1_R1162_U54 , P1_REG1_REG_11_ );
not NOT1_8855 ( P1_R1162_U55 , P1_U3484 );
nand NAND2_8856 ( P1_R1162_U56 , P1_U3484 , P1_REG1_REG_11_ );
not NOT1_8857 ( P1_R1162_U57 , P1_REG1_REG_13_ );
not NOT1_8858 ( P1_R1162_U58 , P1_U3490 );
not NOT1_8859 ( P1_R1162_U59 , P1_REG1_REG_14_ );
not NOT1_8860 ( P1_R1162_U60 , P1_U3493 );
not NOT1_8861 ( P1_R1162_U61 , P1_REG1_REG_15_ );
not NOT1_8862 ( P1_R1162_U62 , P1_U3496 );
not NOT1_8863 ( P1_R1162_U63 , P1_REG1_REG_18_ );
not NOT1_8864 ( P1_R1162_U64 , P1_U3505 );
nand NAND3_8865 ( P1_R1162_U65 , P1_R1162_U186 , P1_R1162_U185 , P1_R1162_U187 );
nand NAND2_8866 ( P1_R1162_U66 , P1_R1162_U179 , P1_R1162_U178 );
nand NAND2_8867 ( P1_R1162_U67 , P1_R1162_U56 , P1_R1162_U204 );
nand NAND2_8868 ( P1_R1162_U68 , P1_R1162_U259 , P1_R1162_U258 );
nand NAND2_8869 ( P1_R1162_U69 , P1_R1162_U308 , P1_R1162_U307 );
nand NAND2_8870 ( P1_R1162_U70 , P1_R1162_U231 , P1_R1162_U230 );
nand NAND2_8871 ( P1_R1162_U71 , P1_R1162_U236 , P1_R1162_U235 );
nand NAND2_8872 ( P1_R1162_U72 , P1_R1162_U243 , P1_R1162_U242 );
nand NAND2_8873 ( P1_R1162_U73 , P1_R1162_U250 , P1_R1162_U249 );
nand NAND2_8874 ( P1_R1162_U74 , P1_R1162_U255 , P1_R1162_U254 );
nand NAND2_8875 ( P1_R1162_U75 , P1_R1162_U271 , P1_R1162_U270 );
nand NAND2_8876 ( P1_R1162_U76 , P1_R1162_U278 , P1_R1162_U277 );
nand NAND2_8877 ( P1_R1162_U77 , P1_R1162_U285 , P1_R1162_U284 );
nand NAND2_8878 ( P1_R1162_U78 , P1_R1162_U292 , P1_R1162_U291 );
nand NAND2_8879 ( P1_R1162_U79 , P1_R1162_U299 , P1_R1162_U298 );
nand NAND2_8880 ( P1_R1162_U80 , P1_R1162_U304 , P1_R1162_U303 );
nand NAND3_8881 ( P1_R1162_U81 , P1_R1162_U117 , P1_R1162_U116 , P1_R1162_U118 );
nand NAND2_8882 ( P1_R1162_U82 , P1_R1162_U133 , P1_R1162_U145 );
nand NAND2_8883 ( P1_R1162_U83 , P1_R1162_U41 , P1_R1162_U152 );
not NOT1_8884 ( P1_R1162_U84 , P1_U3442 );
not NOT1_8885 ( P1_R1162_U85 , P1_REG1_REG_19_ );
nand NAND2_8886 ( P1_R1162_U86 , P1_R1162_U175 , P1_R1162_U174 );
nand NAND2_8887 ( P1_R1162_U87 , P1_R1162_U171 , P1_R1162_U170 );
nand NAND2_8888 ( P1_R1162_U88 , P1_R1162_U161 , P1_R1162_U160 );
not NOT1_8889 ( P1_R1162_U89 , P1_R1162_U32 );
nand NAND2_8890 ( P1_R1162_U90 , P1_REG1_REG_9_ , P1_U3478 );
nand NAND2_8891 ( P1_R1162_U91 , P1_U3487 , P1_REG1_REG_12_ );
not NOT1_8892 ( P1_R1162_U92 , P1_R1162_U56 );
not NOT1_8893 ( P1_R1162_U93 , P1_R1162_U49 );
or OR2_8894 ( P1_R1162_U94 , P1_U3466 , P1_REG1_REG_5_ );
or OR2_8895 ( P1_R1162_U95 , P1_U3463 , P1_REG1_REG_4_ );
or OR2_8896 ( P1_R1162_U96 , P1_REG1_REG_3_ , P1_U3460 );
or OR2_8897 ( P1_R1162_U97 , P1_REG1_REG_2_ , P1_U3457 );
not NOT1_8898 ( P1_R1162_U98 , P1_R1162_U29 );
or OR2_8899 ( P1_R1162_U99 , P1_REG1_REG_1_ , P1_U3454 );
not NOT1_8900 ( P1_R1162_U100 , P1_R1162_U40 );
not NOT1_8901 ( P1_R1162_U101 , P1_R1162_U41 );
nand NAND2_8902 ( P1_R1162_U102 , P1_R1162_U40 , P1_R1162_U41 );
nand NAND3_8903 ( P1_R1162_U103 , P1_REG1_REG_2_ , P1_U3457 , P1_R1162_U96 );
nand NAND2_8904 ( P1_R1162_U104 , P1_R1162_U5 , P1_R1162_U102 );
nand NAND2_8905 ( P1_R1162_U105 , P1_U3460 , P1_REG1_REG_3_ );
nand NAND3_8906 ( P1_R1162_U106 , P1_R1162_U105 , P1_R1162_U103 , P1_R1162_U104 );
nand NAND2_8907 ( P1_R1162_U107 , P1_R1162_U33 , P1_R1162_U32 );
nand NAND2_8908 ( P1_R1162_U108 , P1_U3466 , P1_R1162_U107 );
nand NAND2_8909 ( P1_R1162_U109 , P1_R1162_U4 , P1_R1162_U106 );
nand NAND2_8910 ( P1_R1162_U110 , P1_REG1_REG_5_ , P1_R1162_U89 );
not NOT1_8911 ( P1_R1162_U111 , P1_R1162_U39 );
or OR2_8912 ( P1_R1162_U112 , P1_U3472 , P1_REG1_REG_7_ );
or OR2_8913 ( P1_R1162_U113 , P1_U3469 , P1_REG1_REG_6_ );
not NOT1_8914 ( P1_R1162_U114 , P1_R1162_U20 );
nand NAND2_8915 ( P1_R1162_U115 , P1_R1162_U21 , P1_R1162_U20 );
nand NAND2_8916 ( P1_R1162_U116 , P1_U3472 , P1_R1162_U115 );
nand NAND2_8917 ( P1_R1162_U117 , P1_REG1_REG_7_ , P1_R1162_U114 );
nand NAND2_8918 ( P1_R1162_U118 , P1_R1162_U6 , P1_R1162_U39 );
not NOT1_8919 ( P1_R1162_U119 , P1_R1162_U81 );
or OR2_8920 ( P1_R1162_U120 , P1_REG1_REG_8_ , P1_U3475 );
nand NAND2_8921 ( P1_R1162_U121 , P1_R1162_U120 , P1_R1162_U81 );
not NOT1_8922 ( P1_R1162_U122 , P1_R1162_U38 );
or OR2_8923 ( P1_R1162_U123 , P1_U3478 , P1_REG1_REG_9_ );
or OR2_8924 ( P1_R1162_U124 , P1_REG1_REG_6_ , P1_U3469 );
nand NAND2_8925 ( P1_R1162_U125 , P1_R1162_U124 , P1_R1162_U39 );
nand NAND4_8926 ( P1_R1162_U126 , P1_R1162_U238 , P1_R1162_U237 , P1_R1162_U20 , P1_R1162_U125 );
nand NAND2_8927 ( P1_R1162_U127 , P1_R1162_U111 , P1_R1162_U20 );
nand NAND2_8928 ( P1_R1162_U128 , P1_REG1_REG_7_ , P1_U3472 );
nand NAND3_8929 ( P1_R1162_U129 , P1_R1162_U128 , P1_R1162_U6 , P1_R1162_U127 );
or OR2_8930 ( P1_R1162_U130 , P1_U3469 , P1_REG1_REG_6_ );
nand NAND2_8931 ( P1_R1162_U131 , P1_R1162_U101 , P1_R1162_U97 );
nand NAND2_8932 ( P1_R1162_U132 , P1_U3457 , P1_REG1_REG_2_ );
not NOT1_8933 ( P1_R1162_U133 , P1_R1162_U43 );
nand NAND2_8934 ( P1_R1162_U134 , P1_R1162_U100 , P1_R1162_U5 );
nand NAND2_8935 ( P1_R1162_U135 , P1_R1162_U43 , P1_R1162_U96 );
nand NAND2_8936 ( P1_R1162_U136 , P1_U3460 , P1_REG1_REG_3_ );
not NOT1_8937 ( P1_R1162_U137 , P1_R1162_U42 );
or OR2_8938 ( P1_R1162_U138 , P1_REG1_REG_4_ , P1_U3463 );
nand NAND2_8939 ( P1_R1162_U139 , P1_R1162_U138 , P1_R1162_U42 );
nand NAND4_8940 ( P1_R1162_U140 , P1_R1162_U245 , P1_R1162_U244 , P1_R1162_U32 , P1_R1162_U139 );
nand NAND2_8941 ( P1_R1162_U141 , P1_R1162_U137 , P1_R1162_U32 );
nand NAND2_8942 ( P1_R1162_U142 , P1_REG1_REG_5_ , P1_U3466 );
nand NAND3_8943 ( P1_R1162_U143 , P1_R1162_U142 , P1_R1162_U4 , P1_R1162_U141 );
or OR2_8944 ( P1_R1162_U144 , P1_U3463 , P1_REG1_REG_4_ );
nand NAND2_8945 ( P1_R1162_U145 , P1_R1162_U100 , P1_R1162_U97 );
not NOT1_8946 ( P1_R1162_U146 , P1_R1162_U82 );
nand NAND2_8947 ( P1_R1162_U147 , P1_U3460 , P1_REG1_REG_3_ );
nand NAND4_8948 ( P1_R1162_U148 , P1_R1162_U257 , P1_R1162_U256 , P1_R1162_U41 , P1_R1162_U40 );
nand NAND2_8949 ( P1_R1162_U149 , P1_R1162_U41 , P1_R1162_U40 );
nand NAND2_8950 ( P1_R1162_U150 , P1_U3457 , P1_REG1_REG_2_ );
nand NAND3_8951 ( P1_R1162_U151 , P1_R1162_U150 , P1_R1162_U97 , P1_R1162_U149 );
or OR2_8952 ( P1_R1162_U152 , P1_REG1_REG_1_ , P1_U3454 );
not NOT1_8953 ( P1_R1162_U153 , P1_R1162_U83 );
or OR2_8954 ( P1_R1162_U154 , P1_U3478 , P1_REG1_REG_9_ );
or OR2_8955 ( P1_R1162_U155 , P1_U3481 , P1_REG1_REG_10_ );
nand NAND2_8956 ( P1_R1162_U156 , P1_R1162_U93 , P1_R1162_U7 );
nand NAND2_8957 ( P1_R1162_U157 , P1_U3481 , P1_REG1_REG_10_ );
nand NAND3_8958 ( P1_R1162_U158 , P1_R1162_U157 , P1_R1162_U90 , P1_R1162_U156 );
or OR2_8959 ( P1_R1162_U159 , P1_REG1_REG_10_ , P1_U3481 );
nand NAND3_8960 ( P1_R1162_U160 , P1_R1162_U120 , P1_R1162_U7 , P1_R1162_U81 );
nand NAND2_8961 ( P1_R1162_U161 , P1_R1162_U159 , P1_R1162_U158 );
not NOT1_8962 ( P1_R1162_U162 , P1_R1162_U88 );
or OR2_8963 ( P1_R1162_U163 , P1_U3490 , P1_REG1_REG_13_ );
or OR2_8964 ( P1_R1162_U164 , P1_U3487 , P1_REG1_REG_12_ );
nand NAND2_8965 ( P1_R1162_U165 , P1_R1162_U92 , P1_R1162_U8 );
nand NAND2_8966 ( P1_R1162_U166 , P1_U3490 , P1_REG1_REG_13_ );
nand NAND3_8967 ( P1_R1162_U167 , P1_R1162_U166 , P1_R1162_U91 , P1_R1162_U165 );
or OR2_8968 ( P1_R1162_U168 , P1_REG1_REG_11_ , P1_U3484 );
or OR2_8969 ( P1_R1162_U169 , P1_REG1_REG_13_ , P1_U3490 );
nand NAND3_8970 ( P1_R1162_U170 , P1_R1162_U168 , P1_R1162_U8 , P1_R1162_U88 );
nand NAND2_8971 ( P1_R1162_U171 , P1_R1162_U169 , P1_R1162_U167 );
not NOT1_8972 ( P1_R1162_U172 , P1_R1162_U87 );
or OR2_8973 ( P1_R1162_U173 , P1_REG1_REG_14_ , P1_U3493 );
nand NAND2_8974 ( P1_R1162_U174 , P1_R1162_U173 , P1_R1162_U87 );
nand NAND2_8975 ( P1_R1162_U175 , P1_U3493 , P1_REG1_REG_14_ );
not NOT1_8976 ( P1_R1162_U176 , P1_R1162_U86 );
or OR2_8977 ( P1_R1162_U177 , P1_REG1_REG_15_ , P1_U3496 );
nand NAND2_8978 ( P1_R1162_U178 , P1_R1162_U177 , P1_R1162_U86 );
nand NAND2_8979 ( P1_R1162_U179 , P1_U3496 , P1_REG1_REG_15_ );
not NOT1_8980 ( P1_R1162_U180 , P1_R1162_U66 );
or OR2_8981 ( P1_R1162_U181 , P1_U3502 , P1_REG1_REG_17_ );
or OR2_8982 ( P1_R1162_U182 , P1_U3499 , P1_REG1_REG_16_ );
not NOT1_8983 ( P1_R1162_U183 , P1_R1162_U47 );
nand NAND2_8984 ( P1_R1162_U184 , P1_R1162_U48 , P1_R1162_U47 );
nand NAND2_8985 ( P1_R1162_U185 , P1_U3502 , P1_R1162_U184 );
nand NAND2_8986 ( P1_R1162_U186 , P1_REG1_REG_17_ , P1_R1162_U183 );
nand NAND2_8987 ( P1_R1162_U187 , P1_R1162_U9 , P1_R1162_U66 );
not NOT1_8988 ( P1_R1162_U188 , P1_R1162_U65 );
or OR2_8989 ( P1_R1162_U189 , P1_REG1_REG_18_ , P1_U3505 );
nand NAND2_8990 ( P1_R1162_U190 , P1_R1162_U189 , P1_R1162_U65 );
nand NAND2_8991 ( P1_R1162_U191 , P1_U3505 , P1_REG1_REG_18_ );
nand NAND4_8992 ( P1_R1162_U192 , P1_R1162_U261 , P1_R1162_U260 , P1_R1162_U191 , P1_R1162_U190 );
nand NAND2_8993 ( P1_R1162_U193 , P1_U3505 , P1_REG1_REG_18_ );
nand NAND2_8994 ( P1_R1162_U194 , P1_R1162_U188 , P1_R1162_U193 );
or OR2_8995 ( P1_R1162_U195 , P1_U3505 , P1_REG1_REG_18_ );
nand NAND3_8996 ( P1_R1162_U196 , P1_R1162_U195 , P1_R1162_U264 , P1_R1162_U194 );
or OR2_8997 ( P1_R1162_U197 , P1_REG1_REG_16_ , P1_U3499 );
nand NAND2_8998 ( P1_R1162_U198 , P1_R1162_U197 , P1_R1162_U66 );
nand NAND4_8999 ( P1_R1162_U199 , P1_R1162_U273 , P1_R1162_U272 , P1_R1162_U47 , P1_R1162_U198 );
nand NAND2_9000 ( P1_R1162_U200 , P1_R1162_U180 , P1_R1162_U47 );
nand NAND2_9001 ( P1_R1162_U201 , P1_REG1_REG_17_ , P1_U3502 );
nand NAND3_9002 ( P1_R1162_U202 , P1_R1162_U201 , P1_R1162_U9 , P1_R1162_U200 );
or OR2_9003 ( P1_R1162_U203 , P1_U3499 , P1_REG1_REG_16_ );
nand NAND2_9004 ( P1_R1162_U204 , P1_R1162_U168 , P1_R1162_U88 );
not NOT1_9005 ( P1_R1162_U205 , P1_R1162_U67 );
or OR2_9006 ( P1_R1162_U206 , P1_REG1_REG_12_ , P1_U3487 );
nand NAND2_9007 ( P1_R1162_U207 , P1_R1162_U206 , P1_R1162_U67 );
nand NAND4_9008 ( P1_R1162_U208 , P1_R1162_U294 , P1_R1162_U293 , P1_R1162_U91 , P1_R1162_U207 );
nand NAND2_9009 ( P1_R1162_U209 , P1_R1162_U205 , P1_R1162_U91 );
nand NAND2_9010 ( P1_R1162_U210 , P1_U3490 , P1_REG1_REG_13_ );
nand NAND3_9011 ( P1_R1162_U211 , P1_R1162_U210 , P1_R1162_U8 , P1_R1162_U209 );
or OR2_9012 ( P1_R1162_U212 , P1_U3487 , P1_REG1_REG_12_ );
or OR2_9013 ( P1_R1162_U213 , P1_REG1_REG_9_ , P1_U3478 );
nand NAND2_9014 ( P1_R1162_U214 , P1_R1162_U213 , P1_R1162_U38 );
nand NAND4_9015 ( P1_R1162_U215 , P1_R1162_U306 , P1_R1162_U305 , P1_R1162_U90 , P1_R1162_U214 );
nand NAND2_9016 ( P1_R1162_U216 , P1_R1162_U122 , P1_R1162_U90 );
nand NAND2_9017 ( P1_R1162_U217 , P1_U3481 , P1_REG1_REG_10_ );
nand NAND3_9018 ( P1_R1162_U218 , P1_R1162_U217 , P1_R1162_U7 , P1_R1162_U216 );
nand NAND2_9019 ( P1_R1162_U219 , P1_R1162_U123 , P1_R1162_U90 );
nand NAND2_9020 ( P1_R1162_U220 , P1_R1162_U120 , P1_R1162_U49 );
nand NAND2_9021 ( P1_R1162_U221 , P1_R1162_U130 , P1_R1162_U20 );
nand NAND2_9022 ( P1_R1162_U222 , P1_R1162_U144 , P1_R1162_U32 );
nand NAND2_9023 ( P1_R1162_U223 , P1_R1162_U147 , P1_R1162_U96 );
nand NAND2_9024 ( P1_R1162_U224 , P1_R1162_U203 , P1_R1162_U47 );
nand NAND2_9025 ( P1_R1162_U225 , P1_R1162_U212 , P1_R1162_U91 );
nand NAND2_9026 ( P1_R1162_U226 , P1_R1162_U168 , P1_R1162_U56 );
nand NAND2_9027 ( P1_R1162_U227 , P1_U3478 , P1_R1162_U37 );
nand NAND2_9028 ( P1_R1162_U228 , P1_REG1_REG_9_ , P1_R1162_U36 );
nand NAND2_9029 ( P1_R1162_U229 , P1_R1162_U228 , P1_R1162_U227 );
nand NAND2_9030 ( P1_R1162_U230 , P1_R1162_U219 , P1_R1162_U38 );
nand NAND2_9031 ( P1_R1162_U231 , P1_R1162_U229 , P1_R1162_U122 );
nand NAND2_9032 ( P1_R1162_U232 , P1_U3475 , P1_R1162_U34 );
nand NAND2_9033 ( P1_R1162_U233 , P1_REG1_REG_8_ , P1_R1162_U35 );
nand NAND2_9034 ( P1_R1162_U234 , P1_R1162_U233 , P1_R1162_U232 );
nand NAND2_9035 ( P1_R1162_U235 , P1_R1162_U220 , P1_R1162_U81 );
nand NAND2_9036 ( P1_R1162_U236 , P1_R1162_U119 , P1_R1162_U234 );
nand NAND2_9037 ( P1_R1162_U237 , P1_U3472 , P1_R1162_U21 );
nand NAND2_9038 ( P1_R1162_U238 , P1_REG1_REG_7_ , P1_R1162_U19 );
nand NAND2_9039 ( P1_R1162_U239 , P1_U3469 , P1_R1162_U17 );
nand NAND2_9040 ( P1_R1162_U240 , P1_REG1_REG_6_ , P1_R1162_U18 );
nand NAND2_9041 ( P1_R1162_U241 , P1_R1162_U240 , P1_R1162_U239 );
nand NAND2_9042 ( P1_R1162_U242 , P1_R1162_U221 , P1_R1162_U39 );
nand NAND2_9043 ( P1_R1162_U243 , P1_R1162_U241 , P1_R1162_U111 );
nand NAND2_9044 ( P1_R1162_U244 , P1_U3466 , P1_R1162_U33 );
nand NAND2_9045 ( P1_R1162_U245 , P1_REG1_REG_5_ , P1_R1162_U24 );
nand NAND2_9046 ( P1_R1162_U246 , P1_U3463 , P1_R1162_U22 );
nand NAND2_9047 ( P1_R1162_U247 , P1_REG1_REG_4_ , P1_R1162_U23 );
nand NAND2_9048 ( P1_R1162_U248 , P1_R1162_U247 , P1_R1162_U246 );
nand NAND2_9049 ( P1_R1162_U249 , P1_R1162_U222 , P1_R1162_U42 );
nand NAND2_9050 ( P1_R1162_U250 , P1_R1162_U248 , P1_R1162_U137 );
nand NAND2_9051 ( P1_R1162_U251 , P1_U3460 , P1_R1162_U30 );
nand NAND2_9052 ( P1_R1162_U252 , P1_REG1_REG_3_ , P1_R1162_U31 );
nand NAND2_9053 ( P1_R1162_U253 , P1_R1162_U252 , P1_R1162_U251 );
nand NAND2_9054 ( P1_R1162_U254 , P1_R1162_U223 , P1_R1162_U82 );
nand NAND2_9055 ( P1_R1162_U255 , P1_R1162_U146 , P1_R1162_U253 );
nand NAND2_9056 ( P1_R1162_U256 , P1_U3457 , P1_R1162_U25 );
nand NAND2_9057 ( P1_R1162_U257 , P1_REG1_REG_2_ , P1_R1162_U26 );
nand NAND2_9058 ( P1_R1162_U258 , P1_R1162_U98 , P1_R1162_U83 );
nand NAND2_9059 ( P1_R1162_U259 , P1_R1162_U153 , P1_R1162_U29 );
nand NAND2_9060 ( P1_R1162_U260 , P1_U3442 , P1_R1162_U85 );
nand NAND2_9061 ( P1_R1162_U261 , P1_REG1_REG_19_ , P1_R1162_U84 );
nand NAND2_9062 ( P1_R1162_U262 , P1_U3442 , P1_R1162_U85 );
nand NAND2_9063 ( P1_R1162_U263 , P1_REG1_REG_19_ , P1_R1162_U84 );
nand NAND2_9064 ( P1_R1162_U264 , P1_R1162_U263 , P1_R1162_U262 );
nand NAND2_9065 ( P1_R1162_U265 , P1_U3505 , P1_R1162_U63 );
nand NAND2_9066 ( P1_R1162_U266 , P1_REG1_REG_18_ , P1_R1162_U64 );
nand NAND2_9067 ( P1_R1162_U267 , P1_U3505 , P1_R1162_U63 );
nand NAND2_9068 ( P1_R1162_U268 , P1_REG1_REG_18_ , P1_R1162_U64 );
nand NAND2_9069 ( P1_R1162_U269 , P1_R1162_U268 , P1_R1162_U267 );
nand NAND3_9070 ( P1_R1162_U270 , P1_R1162_U266 , P1_R1162_U265 , P1_R1162_U65 );
nand NAND2_9071 ( P1_R1162_U271 , P1_R1162_U269 , P1_R1162_U188 );
nand NAND2_9072 ( P1_R1162_U272 , P1_U3502 , P1_R1162_U48 );
nand NAND2_9073 ( P1_R1162_U273 , P1_REG1_REG_17_ , P1_R1162_U46 );
nand NAND2_9074 ( P1_R1162_U274 , P1_U3499 , P1_R1162_U44 );
nand NAND2_9075 ( P1_R1162_U275 , P1_REG1_REG_16_ , P1_R1162_U45 );
nand NAND2_9076 ( P1_R1162_U276 , P1_R1162_U275 , P1_R1162_U274 );
nand NAND2_9077 ( P1_R1162_U277 , P1_R1162_U224 , P1_R1162_U66 );
nand NAND2_9078 ( P1_R1162_U278 , P1_R1162_U276 , P1_R1162_U180 );
nand NAND2_9079 ( P1_R1162_U279 , P1_U3496 , P1_R1162_U61 );
nand NAND2_9080 ( P1_R1162_U280 , P1_REG1_REG_15_ , P1_R1162_U62 );
nand NAND2_9081 ( P1_R1162_U281 , P1_U3496 , P1_R1162_U61 );
nand NAND2_9082 ( P1_R1162_U282 , P1_REG1_REG_15_ , P1_R1162_U62 );
nand NAND2_9083 ( P1_R1162_U283 , P1_R1162_U282 , P1_R1162_U281 );
nand NAND3_9084 ( P1_R1162_U284 , P1_R1162_U280 , P1_R1162_U279 , P1_R1162_U86 );
nand NAND2_9085 ( P1_R1162_U285 , P1_R1162_U176 , P1_R1162_U283 );
nand NAND2_9086 ( P1_R1162_U286 , P1_U3493 , P1_R1162_U59 );
nand NAND2_9087 ( P1_R1162_U287 , P1_REG1_REG_14_ , P1_R1162_U60 );
nand NAND2_9088 ( P1_R1162_U288 , P1_U3493 , P1_R1162_U59 );
nand NAND2_9089 ( P1_R1162_U289 , P1_REG1_REG_14_ , P1_R1162_U60 );
nand NAND2_9090 ( P1_R1162_U290 , P1_R1162_U289 , P1_R1162_U288 );
nand NAND3_9091 ( P1_R1162_U291 , P1_R1162_U287 , P1_R1162_U286 , P1_R1162_U87 );
nand NAND2_9092 ( P1_R1162_U292 , P1_R1162_U172 , P1_R1162_U290 );
nand NAND2_9093 ( P1_R1162_U293 , P1_U3490 , P1_R1162_U57 );
nand NAND2_9094 ( P1_R1162_U294 , P1_REG1_REG_13_ , P1_R1162_U58 );
nand NAND2_9095 ( P1_R1162_U295 , P1_U3487 , P1_R1162_U52 );
nand NAND2_9096 ( P1_R1162_U296 , P1_REG1_REG_12_ , P1_R1162_U53 );
nand NAND2_9097 ( P1_R1162_U297 , P1_R1162_U296 , P1_R1162_U295 );
nand NAND2_9098 ( P1_R1162_U298 , P1_R1162_U225 , P1_R1162_U67 );
nand NAND2_9099 ( P1_R1162_U299 , P1_R1162_U297 , P1_R1162_U205 );
nand NAND2_9100 ( P1_R1162_U300 , P1_U3484 , P1_R1162_U54 );
nand NAND2_9101 ( P1_R1162_U301 , P1_REG1_REG_11_ , P1_R1162_U55 );
nand NAND2_9102 ( P1_R1162_U302 , P1_R1162_U301 , P1_R1162_U300 );
nand NAND2_9103 ( P1_R1162_U303 , P1_R1162_U226 , P1_R1162_U88 );
nand NAND2_9104 ( P1_R1162_U304 , P1_R1162_U162 , P1_R1162_U302 );
nand NAND2_9105 ( P1_R1162_U305 , P1_U3481 , P1_R1162_U50 );
nand NAND2_9106 ( P1_R1162_U306 , P1_REG1_REG_10_ , P1_R1162_U51 );
nand NAND2_9107 ( P1_R1162_U307 , P1_U3448 , P1_R1162_U27 );
nand NAND2_9108 ( P1_R1162_U308 , P1_REG1_REG_0_ , P1_R1162_U28 );
and AND2_9109 ( P1_R1117_U6 , P1_R1117_U198 , P1_R1117_U197 );
and AND2_9110 ( P1_R1117_U7 , P1_R1117_U237 , P1_R1117_U236 );
and AND2_9111 ( P1_R1117_U8 , P1_R1117_U254 , P1_R1117_U253 );
and AND2_9112 ( P1_R1117_U9 , P1_R1117_U280 , P1_R1117_U279 );
nand NAND2_9113 ( P1_R1117_U10 , P1_R1117_U340 , P1_R1117_U343 );
nand NAND2_9114 ( P1_R1117_U11 , P1_R1117_U329 , P1_R1117_U332 );
nand NAND2_9115 ( P1_R1117_U12 , P1_R1117_U318 , P1_R1117_U321 );
nand NAND2_9116 ( P1_R1117_U13 , P1_R1117_U310 , P1_R1117_U312 );
nand NAND2_9117 ( P1_R1117_U14 , P1_R1117_U347 , P1_R1117_U308 );
nand NAND2_9118 ( P1_R1117_U15 , P1_R1117_U231 , P1_R1117_U233 );
nand NAND2_9119 ( P1_R1117_U16 , P1_R1117_U223 , P1_R1117_U226 );
nand NAND2_9120 ( P1_R1117_U17 , P1_R1117_U215 , P1_R1117_U217 );
nand NAND2_9121 ( P1_R1117_U18 , P1_R1117_U23 , P1_R1117_U346 );
not NOT1_9122 ( P1_R1117_U19 , P1_U3473 );
not NOT1_9123 ( P1_R1117_U20 , P1_U3467 );
not NOT1_9124 ( P1_R1117_U21 , P1_U3458 );
not NOT1_9125 ( P1_R1117_U22 , P1_U3450 );
nand NAND2_9126 ( P1_R1117_U23 , P1_U3450 , P1_R1117_U91 );
not NOT1_9127 ( P1_R1117_U24 , P1_U3078 );
not NOT1_9128 ( P1_R1117_U25 , P1_U3461 );
not NOT1_9129 ( P1_R1117_U26 , P1_U3068 );
nand NAND2_9130 ( P1_R1117_U27 , P1_U3068 , P1_R1117_U21 );
not NOT1_9131 ( P1_R1117_U28 , P1_U3064 );
not NOT1_9132 ( P1_R1117_U29 , P1_U3470 );
not NOT1_9133 ( P1_R1117_U30 , P1_U3464 );
not NOT1_9134 ( P1_R1117_U31 , P1_U3071 );
not NOT1_9135 ( P1_R1117_U32 , P1_U3067 );
not NOT1_9136 ( P1_R1117_U33 , P1_U3060 );
nand NAND2_9137 ( P1_R1117_U34 , P1_U3060 , P1_R1117_U30 );
not NOT1_9138 ( P1_R1117_U35 , P1_U3476 );
not NOT1_9139 ( P1_R1117_U36 , P1_U3070 );
nand NAND2_9140 ( P1_R1117_U37 , P1_U3070 , P1_R1117_U19 );
not NOT1_9141 ( P1_R1117_U38 , P1_U3084 );
not NOT1_9142 ( P1_R1117_U39 , P1_U3479 );
not NOT1_9143 ( P1_R1117_U40 , P1_U3083 );
nand NAND2_9144 ( P1_R1117_U41 , P1_R1117_U204 , P1_R1117_U203 );
nand NAND2_9145 ( P1_R1117_U42 , P1_R1117_U34 , P1_R1117_U219 );
nand NAND2_9146 ( P1_R1117_U43 , P1_R1117_U188 , P1_R1117_U187 );
not NOT1_9147 ( P1_R1117_U44 , P1_U3976 );
not NOT1_9148 ( P1_R1117_U45 , P1_U3980 );
not NOT1_9149 ( P1_R1117_U46 , P1_U3497 );
not NOT1_9150 ( P1_R1117_U47 , P1_U3482 );
not NOT1_9151 ( P1_R1117_U48 , P1_U3485 );
not NOT1_9152 ( P1_R1117_U49 , P1_U3063 );
not NOT1_9153 ( P1_R1117_U50 , P1_U3062 );
nand NAND2_9154 ( P1_R1117_U51 , P1_U3083 , P1_R1117_U39 );
not NOT1_9155 ( P1_R1117_U52 , P1_U3488 );
not NOT1_9156 ( P1_R1117_U53 , P1_U3072 );
not NOT1_9157 ( P1_R1117_U54 , P1_U3491 );
not NOT1_9158 ( P1_R1117_U55 , P1_U3080 );
not NOT1_9159 ( P1_R1117_U56 , P1_U3500 );
not NOT1_9160 ( P1_R1117_U57 , P1_U3494 );
not NOT1_9161 ( P1_R1117_U58 , P1_U3073 );
not NOT1_9162 ( P1_R1117_U59 , P1_U3074 );
not NOT1_9163 ( P1_R1117_U60 , P1_U3079 );
nand NAND2_9164 ( P1_R1117_U61 , P1_U3079 , P1_R1117_U57 );
not NOT1_9165 ( P1_R1117_U62 , P1_U3503 );
not NOT1_9166 ( P1_R1117_U63 , P1_U3069 );
nand NAND2_9167 ( P1_R1117_U64 , P1_R1117_U264 , P1_R1117_U263 );
not NOT1_9168 ( P1_R1117_U65 , P1_U3082 );
not NOT1_9169 ( P1_R1117_U66 , P1_U3508 );
not NOT1_9170 ( P1_R1117_U67 , P1_U3081 );
not NOT1_9171 ( P1_R1117_U68 , P1_U3982 );
not NOT1_9172 ( P1_R1117_U69 , P1_U3076 );
not NOT1_9173 ( P1_R1117_U70 , P1_U3979 );
not NOT1_9174 ( P1_R1117_U71 , P1_U3981 );
not NOT1_9175 ( P1_R1117_U72 , P1_U3066 );
not NOT1_9176 ( P1_R1117_U73 , P1_U3061 );
not NOT1_9177 ( P1_R1117_U74 , P1_U3075 );
nand NAND2_9178 ( P1_R1117_U75 , P1_U3075 , P1_R1117_U71 );
not NOT1_9179 ( P1_R1117_U76 , P1_U3978 );
not NOT1_9180 ( P1_R1117_U77 , P1_U3065 );
not NOT1_9181 ( P1_R1117_U78 , P1_U3977 );
not NOT1_9182 ( P1_R1117_U79 , P1_U3058 );
not NOT1_9183 ( P1_R1117_U80 , P1_U3975 );
not NOT1_9184 ( P1_R1117_U81 , P1_U3057 );
nand NAND2_9185 ( P1_R1117_U82 , P1_U3057 , P1_R1117_U44 );
not NOT1_9186 ( P1_R1117_U83 , P1_U3053 );
not NOT1_9187 ( P1_R1117_U84 , P1_U3974 );
not NOT1_9188 ( P1_R1117_U85 , P1_U3054 );
nand NAND2_9189 ( P1_R1117_U86 , P1_R1117_U126 , P1_R1117_U297 );
nand NAND2_9190 ( P1_R1117_U87 , P1_R1117_U294 , P1_R1117_U293 );
nand NAND2_9191 ( P1_R1117_U88 , P1_R1117_U75 , P1_R1117_U314 );
nand NAND2_9192 ( P1_R1117_U89 , P1_R1117_U61 , P1_R1117_U325 );
nand NAND2_9193 ( P1_R1117_U90 , P1_R1117_U51 , P1_R1117_U336 );
not NOT1_9194 ( P1_R1117_U91 , P1_U3077 );
nand NAND2_9195 ( P1_R1117_U92 , P1_R1117_U390 , P1_R1117_U389 );
nand NAND2_9196 ( P1_R1117_U93 , P1_R1117_U404 , P1_R1117_U403 );
nand NAND2_9197 ( P1_R1117_U94 , P1_R1117_U409 , P1_R1117_U408 );
nand NAND2_9198 ( P1_R1117_U95 , P1_R1117_U425 , P1_R1117_U424 );
nand NAND2_9199 ( P1_R1117_U96 , P1_R1117_U430 , P1_R1117_U429 );
nand NAND2_9200 ( P1_R1117_U97 , P1_R1117_U435 , P1_R1117_U434 );
nand NAND2_9201 ( P1_R1117_U98 , P1_R1117_U440 , P1_R1117_U439 );
nand NAND2_9202 ( P1_R1117_U99 , P1_R1117_U445 , P1_R1117_U444 );
nand NAND2_9203 ( P1_R1117_U100 , P1_R1117_U461 , P1_R1117_U460 );
nand NAND2_9204 ( P1_R1117_U101 , P1_R1117_U466 , P1_R1117_U465 );
nand NAND2_9205 ( P1_R1117_U102 , P1_R1117_U351 , P1_R1117_U350 );
nand NAND2_9206 ( P1_R1117_U103 , P1_R1117_U360 , P1_R1117_U359 );
nand NAND2_9207 ( P1_R1117_U104 , P1_R1117_U367 , P1_R1117_U366 );
nand NAND2_9208 ( P1_R1117_U105 , P1_R1117_U371 , P1_R1117_U370 );
nand NAND2_9209 ( P1_R1117_U106 , P1_R1117_U380 , P1_R1117_U379 );
nand NAND2_9210 ( P1_R1117_U107 , P1_R1117_U399 , P1_R1117_U398 );
nand NAND2_9211 ( P1_R1117_U108 , P1_R1117_U416 , P1_R1117_U415 );
nand NAND2_9212 ( P1_R1117_U109 , P1_R1117_U420 , P1_R1117_U419 );
nand NAND2_9213 ( P1_R1117_U110 , P1_R1117_U452 , P1_R1117_U451 );
nand NAND2_9214 ( P1_R1117_U111 , P1_R1117_U456 , P1_R1117_U455 );
nand NAND2_9215 ( P1_R1117_U112 , P1_R1117_U473 , P1_R1117_U472 );
and AND2_9216 ( P1_R1117_U113 , P1_R1117_U193 , P1_R1117_U194 );
and AND2_9217 ( P1_R1117_U114 , P1_R1117_U201 , P1_R1117_U196 );
and AND2_9218 ( P1_R1117_U115 , P1_R1117_U206 , P1_R1117_U180 );
and AND2_9219 ( P1_R1117_U116 , P1_R1117_U209 , P1_R1117_U210 );
and AND3_9220 ( P1_R1117_U117 , P1_R1117_U353 , P1_R1117_U352 , P1_R1117_U37 );
and AND2_9221 ( P1_R1117_U118 , P1_R1117_U356 , P1_R1117_U180 );
and AND2_9222 ( P1_R1117_U119 , P1_R1117_U225 , P1_R1117_U6 );
and AND2_9223 ( P1_R1117_U120 , P1_R1117_U363 , P1_R1117_U179 );
and AND3_9224 ( P1_R1117_U121 , P1_R1117_U373 , P1_R1117_U372 , P1_R1117_U27 );
and AND2_9225 ( P1_R1117_U122 , P1_R1117_U376 , P1_R1117_U178 );
and AND3_9226 ( P1_R1117_U123 , P1_R1117_U235 , P1_R1117_U212 , P1_R1117_U174 );
and AND3_9227 ( P1_R1117_U124 , P1_R1117_U257 , P1_R1117_U175 , P1_R1117_U252 );
and AND2_9228 ( P1_R1117_U125 , P1_R1117_U283 , P1_R1117_U176 );
and AND2_9229 ( P1_R1117_U126 , P1_R1117_U299 , P1_R1117_U300 );
nand NAND2_9230 ( P1_R1117_U127 , P1_R1117_U387 , P1_R1117_U386 );
and AND3_9231 ( P1_R1117_U128 , P1_R1117_U392 , P1_R1117_U391 , P1_R1117_U82 );
and AND2_9232 ( P1_R1117_U129 , P1_R1117_U395 , P1_R1117_U177 );
nand NAND2_9233 ( P1_R1117_U130 , P1_R1117_U401 , P1_R1117_U400 );
nand NAND2_9234 ( P1_R1117_U131 , P1_R1117_U406 , P1_R1117_U405 );
and AND2_9235 ( P1_R1117_U132 , P1_R1117_U412 , P1_R1117_U176 );
nand NAND2_9236 ( P1_R1117_U133 , P1_R1117_U422 , P1_R1117_U421 );
nand NAND2_9237 ( P1_R1117_U134 , P1_R1117_U427 , P1_R1117_U426 );
nand NAND2_9238 ( P1_R1117_U135 , P1_R1117_U432 , P1_R1117_U431 );
nand NAND2_9239 ( P1_R1117_U136 , P1_R1117_U437 , P1_R1117_U436 );
nand NAND2_9240 ( P1_R1117_U137 , P1_R1117_U442 , P1_R1117_U441 );
and AND2_9241 ( P1_R1117_U138 , P1_R1117_U331 , P1_R1117_U8 );
and AND2_9242 ( P1_R1117_U139 , P1_R1117_U448 , P1_R1117_U175 );
nand NAND2_9243 ( P1_R1117_U140 , P1_R1117_U458 , P1_R1117_U457 );
nand NAND2_9244 ( P1_R1117_U141 , P1_R1117_U463 , P1_R1117_U462 );
and AND2_9245 ( P1_R1117_U142 , P1_R1117_U342 , P1_R1117_U7 );
and AND2_9246 ( P1_R1117_U143 , P1_R1117_U469 , P1_R1117_U174 );
and AND2_9247 ( P1_R1117_U144 , P1_R1117_U349 , P1_R1117_U348 );
nand NAND2_9248 ( P1_R1117_U145 , P1_R1117_U116 , P1_R1117_U207 );
and AND2_9249 ( P1_R1117_U146 , P1_R1117_U358 , P1_R1117_U357 );
and AND2_9250 ( P1_R1117_U147 , P1_R1117_U365 , P1_R1117_U364 );
and AND2_9251 ( P1_R1117_U148 , P1_R1117_U369 , P1_R1117_U368 );
nand NAND2_9252 ( P1_R1117_U149 , P1_R1117_U113 , P1_R1117_U191 );
and AND2_9253 ( P1_R1117_U150 , P1_R1117_U378 , P1_R1117_U377 );
not NOT1_9254 ( P1_R1117_U151 , P1_U3985 );
not NOT1_9255 ( P1_R1117_U152 , P1_U3055 );
and AND2_9256 ( P1_R1117_U153 , P1_R1117_U382 , P1_R1117_U381 );
and AND2_9257 ( P1_R1117_U154 , P1_R1117_U397 , P1_R1117_U396 );
nand NAND2_9258 ( P1_R1117_U155 , P1_R1117_U290 , P1_R1117_U289 );
nand NAND2_9259 ( P1_R1117_U156 , P1_R1117_U286 , P1_R1117_U285 );
and AND2_9260 ( P1_R1117_U157 , P1_R1117_U414 , P1_R1117_U413 );
and AND2_9261 ( P1_R1117_U158 , P1_R1117_U418 , P1_R1117_U417 );
nand NAND2_9262 ( P1_R1117_U159 , P1_R1117_U276 , P1_R1117_U275 );
nand NAND2_9263 ( P1_R1117_U160 , P1_R1117_U272 , P1_R1117_U271 );
not NOT1_9264 ( P1_R1117_U161 , P1_U3455 );
nand NAND2_9265 ( P1_R1117_U162 , P1_R1117_U268 , P1_R1117_U267 );
not NOT1_9266 ( P1_R1117_U163 , P1_U3506 );
nand NAND2_9267 ( P1_R1117_U164 , P1_R1117_U260 , P1_R1117_U259 );
and AND2_9268 ( P1_R1117_U165 , P1_R1117_U450 , P1_R1117_U449 );
and AND2_9269 ( P1_R1117_U166 , P1_R1117_U454 , P1_R1117_U453 );
nand NAND2_9270 ( P1_R1117_U167 , P1_R1117_U250 , P1_R1117_U249 );
nand NAND2_9271 ( P1_R1117_U168 , P1_R1117_U246 , P1_R1117_U245 );
nand NAND2_9272 ( P1_R1117_U169 , P1_R1117_U242 , P1_R1117_U241 );
and AND2_9273 ( P1_R1117_U170 , P1_R1117_U471 , P1_R1117_U470 );
not NOT1_9274 ( P1_R1117_U171 , P1_R1117_U82 );
not NOT1_9275 ( P1_R1117_U172 , P1_R1117_U27 );
not NOT1_9276 ( P1_R1117_U173 , P1_R1117_U37 );
nand NAND2_9277 ( P1_R1117_U174 , P1_U3482 , P1_R1117_U50 );
nand NAND2_9278 ( P1_R1117_U175 , P1_U3497 , P1_R1117_U59 );
nand NAND2_9279 ( P1_R1117_U176 , P1_U3980 , P1_R1117_U73 );
nand NAND2_9280 ( P1_R1117_U177 , P1_U3976 , P1_R1117_U81 );
nand NAND2_9281 ( P1_R1117_U178 , P1_U3458 , P1_R1117_U26 );
nand NAND2_9282 ( P1_R1117_U179 , P1_U3467 , P1_R1117_U32 );
nand NAND2_9283 ( P1_R1117_U180 , P1_U3473 , P1_R1117_U36 );
not NOT1_9284 ( P1_R1117_U181 , P1_R1117_U61 );
not NOT1_9285 ( P1_R1117_U182 , P1_R1117_U75 );
not NOT1_9286 ( P1_R1117_U183 , P1_R1117_U34 );
not NOT1_9287 ( P1_R1117_U184 , P1_R1117_U51 );
not NOT1_9288 ( P1_R1117_U185 , P1_R1117_U23 );
nand NAND2_9289 ( P1_R1117_U186 , P1_R1117_U185 , P1_R1117_U24 );
nand NAND2_9290 ( P1_R1117_U187 , P1_R1117_U186 , P1_R1117_U161 );
nand NAND2_9291 ( P1_R1117_U188 , P1_U3078 , P1_R1117_U23 );
not NOT1_9292 ( P1_R1117_U189 , P1_R1117_U43 );
nand NAND2_9293 ( P1_R1117_U190 , P1_U3461 , P1_R1117_U28 );
nand NAND3_9294 ( P1_R1117_U191 , P1_R1117_U43 , P1_R1117_U178 , P1_R1117_U190 );
nand NAND2_9295 ( P1_R1117_U192 , P1_R1117_U28 , P1_R1117_U27 );
nand NAND2_9296 ( P1_R1117_U193 , P1_R1117_U192 , P1_R1117_U25 );
nand NAND2_9297 ( P1_R1117_U194 , P1_U3064 , P1_R1117_U172 );
not NOT1_9298 ( P1_R1117_U195 , P1_R1117_U149 );
nand NAND2_9299 ( P1_R1117_U196 , P1_U3470 , P1_R1117_U31 );
nand NAND2_9300 ( P1_R1117_U197 , P1_U3071 , P1_R1117_U29 );
nand NAND2_9301 ( P1_R1117_U198 , P1_U3067 , P1_R1117_U20 );
nand NAND2_9302 ( P1_R1117_U199 , P1_R1117_U183 , P1_R1117_U179 );
nand NAND2_9303 ( P1_R1117_U200 , P1_R1117_U6 , P1_R1117_U199 );
nand NAND2_9304 ( P1_R1117_U201 , P1_U3464 , P1_R1117_U33 );
nand NAND2_9305 ( P1_R1117_U202 , P1_U3470 , P1_R1117_U31 );
nand NAND3_9306 ( P1_R1117_U203 , P1_R1117_U149 , P1_R1117_U179 , P1_R1117_U114 );
nand NAND2_9307 ( P1_R1117_U204 , P1_R1117_U202 , P1_R1117_U200 );
not NOT1_9308 ( P1_R1117_U205 , P1_R1117_U41 );
nand NAND2_9309 ( P1_R1117_U206 , P1_U3476 , P1_R1117_U38 );
nand NAND2_9310 ( P1_R1117_U207 , P1_R1117_U115 , P1_R1117_U41 );
nand NAND2_9311 ( P1_R1117_U208 , P1_R1117_U38 , P1_R1117_U37 );
nand NAND2_9312 ( P1_R1117_U209 , P1_R1117_U208 , P1_R1117_U35 );
nand NAND2_9313 ( P1_R1117_U210 , P1_U3084 , P1_R1117_U173 );
not NOT1_9314 ( P1_R1117_U211 , P1_R1117_U145 );
nand NAND2_9315 ( P1_R1117_U212 , P1_U3479 , P1_R1117_U40 );
nand NAND2_9316 ( P1_R1117_U213 , P1_R1117_U212 , P1_R1117_U51 );
nand NAND2_9317 ( P1_R1117_U214 , P1_R1117_U205 , P1_R1117_U37 );
nand NAND2_9318 ( P1_R1117_U215 , P1_R1117_U118 , P1_R1117_U214 );
nand NAND2_9319 ( P1_R1117_U216 , P1_R1117_U41 , P1_R1117_U180 );
nand NAND2_9320 ( P1_R1117_U217 , P1_R1117_U117 , P1_R1117_U216 );
nand NAND2_9321 ( P1_R1117_U218 , P1_R1117_U37 , P1_R1117_U180 );
nand NAND2_9322 ( P1_R1117_U219 , P1_R1117_U201 , P1_R1117_U149 );
not NOT1_9323 ( P1_R1117_U220 , P1_R1117_U42 );
nand NAND2_9324 ( P1_R1117_U221 , P1_U3067 , P1_R1117_U20 );
nand NAND2_9325 ( P1_R1117_U222 , P1_R1117_U220 , P1_R1117_U221 );
nand NAND2_9326 ( P1_R1117_U223 , P1_R1117_U120 , P1_R1117_U222 );
nand NAND2_9327 ( P1_R1117_U224 , P1_R1117_U42 , P1_R1117_U179 );
nand NAND2_9328 ( P1_R1117_U225 , P1_U3470 , P1_R1117_U31 );
nand NAND2_9329 ( P1_R1117_U226 , P1_R1117_U119 , P1_R1117_U224 );
nand NAND2_9330 ( P1_R1117_U227 , P1_U3067 , P1_R1117_U20 );
nand NAND2_9331 ( P1_R1117_U228 , P1_R1117_U179 , P1_R1117_U227 );
nand NAND2_9332 ( P1_R1117_U229 , P1_R1117_U201 , P1_R1117_U34 );
nand NAND2_9333 ( P1_R1117_U230 , P1_R1117_U189 , P1_R1117_U27 );
nand NAND2_9334 ( P1_R1117_U231 , P1_R1117_U122 , P1_R1117_U230 );
nand NAND2_9335 ( P1_R1117_U232 , P1_R1117_U43 , P1_R1117_U178 );
nand NAND2_9336 ( P1_R1117_U233 , P1_R1117_U121 , P1_R1117_U232 );
nand NAND2_9337 ( P1_R1117_U234 , P1_R1117_U27 , P1_R1117_U178 );
nand NAND2_9338 ( P1_R1117_U235 , P1_U3485 , P1_R1117_U49 );
nand NAND2_9339 ( P1_R1117_U236 , P1_U3063 , P1_R1117_U48 );
nand NAND2_9340 ( P1_R1117_U237 , P1_U3062 , P1_R1117_U47 );
nand NAND2_9341 ( P1_R1117_U238 , P1_R1117_U184 , P1_R1117_U174 );
nand NAND2_9342 ( P1_R1117_U239 , P1_R1117_U7 , P1_R1117_U238 );
nand NAND2_9343 ( P1_R1117_U240 , P1_U3485 , P1_R1117_U49 );
nand NAND2_9344 ( P1_R1117_U241 , P1_R1117_U145 , P1_R1117_U123 );
nand NAND2_9345 ( P1_R1117_U242 , P1_R1117_U240 , P1_R1117_U239 );
not NOT1_9346 ( P1_R1117_U243 , P1_R1117_U169 );
nand NAND2_9347 ( P1_R1117_U244 , P1_U3488 , P1_R1117_U53 );
nand NAND2_9348 ( P1_R1117_U245 , P1_R1117_U244 , P1_R1117_U169 );
nand NAND2_9349 ( P1_R1117_U246 , P1_U3072 , P1_R1117_U52 );
not NOT1_9350 ( P1_R1117_U247 , P1_R1117_U168 );
nand NAND2_9351 ( P1_R1117_U248 , P1_U3491 , P1_R1117_U55 );
nand NAND2_9352 ( P1_R1117_U249 , P1_R1117_U248 , P1_R1117_U168 );
nand NAND2_9353 ( P1_R1117_U250 , P1_U3080 , P1_R1117_U54 );
not NOT1_9354 ( P1_R1117_U251 , P1_R1117_U167 );
nand NAND2_9355 ( P1_R1117_U252 , P1_U3500 , P1_R1117_U58 );
nand NAND2_9356 ( P1_R1117_U253 , P1_U3073 , P1_R1117_U56 );
nand NAND2_9357 ( P1_R1117_U254 , P1_U3074 , P1_R1117_U46 );
nand NAND2_9358 ( P1_R1117_U255 , P1_R1117_U181 , P1_R1117_U175 );
nand NAND2_9359 ( P1_R1117_U256 , P1_R1117_U8 , P1_R1117_U255 );
nand NAND2_9360 ( P1_R1117_U257 , P1_U3494 , P1_R1117_U60 );
nand NAND2_9361 ( P1_R1117_U258 , P1_U3500 , P1_R1117_U58 );
nand NAND2_9362 ( P1_R1117_U259 , P1_R1117_U167 , P1_R1117_U124 );
nand NAND2_9363 ( P1_R1117_U260 , P1_R1117_U258 , P1_R1117_U256 );
not NOT1_9364 ( P1_R1117_U261 , P1_R1117_U164 );
nand NAND2_9365 ( P1_R1117_U262 , P1_U3503 , P1_R1117_U63 );
nand NAND2_9366 ( P1_R1117_U263 , P1_R1117_U262 , P1_R1117_U164 );
nand NAND2_9367 ( P1_R1117_U264 , P1_U3069 , P1_R1117_U62 );
not NOT1_9368 ( P1_R1117_U265 , P1_R1117_U64 );
nand NAND2_9369 ( P1_R1117_U266 , P1_R1117_U265 , P1_R1117_U65 );
nand NAND2_9370 ( P1_R1117_U267 , P1_R1117_U266 , P1_R1117_U163 );
nand NAND2_9371 ( P1_R1117_U268 , P1_U3082 , P1_R1117_U64 );
not NOT1_9372 ( P1_R1117_U269 , P1_R1117_U162 );
nand NAND2_9373 ( P1_R1117_U270 , P1_U3508 , P1_R1117_U67 );
nand NAND2_9374 ( P1_R1117_U271 , P1_R1117_U270 , P1_R1117_U162 );
nand NAND2_9375 ( P1_R1117_U272 , P1_U3081 , P1_R1117_U66 );
not NOT1_9376 ( P1_R1117_U273 , P1_R1117_U160 );
nand NAND2_9377 ( P1_R1117_U274 , P1_U3982 , P1_R1117_U69 );
nand NAND2_9378 ( P1_R1117_U275 , P1_R1117_U274 , P1_R1117_U160 );
nand NAND2_9379 ( P1_R1117_U276 , P1_U3076 , P1_R1117_U68 );
not NOT1_9380 ( P1_R1117_U277 , P1_R1117_U159 );
nand NAND2_9381 ( P1_R1117_U278 , P1_U3979 , P1_R1117_U72 );
nand NAND2_9382 ( P1_R1117_U279 , P1_U3066 , P1_R1117_U70 );
nand NAND2_9383 ( P1_R1117_U280 , P1_U3061 , P1_R1117_U45 );
nand NAND2_9384 ( P1_R1117_U281 , P1_R1117_U182 , P1_R1117_U176 );
nand NAND2_9385 ( P1_R1117_U282 , P1_R1117_U9 , P1_R1117_U281 );
nand NAND2_9386 ( P1_R1117_U283 , P1_U3981 , P1_R1117_U74 );
nand NAND2_9387 ( P1_R1117_U284 , P1_U3979 , P1_R1117_U72 );
nand NAND3_9388 ( P1_R1117_U285 , P1_R1117_U159 , P1_R1117_U125 , P1_R1117_U278 );
nand NAND2_9389 ( P1_R1117_U286 , P1_R1117_U284 , P1_R1117_U282 );
not NOT1_9390 ( P1_R1117_U287 , P1_R1117_U156 );
nand NAND2_9391 ( P1_R1117_U288 , P1_U3978 , P1_R1117_U77 );
nand NAND2_9392 ( P1_R1117_U289 , P1_R1117_U288 , P1_R1117_U156 );
nand NAND2_9393 ( P1_R1117_U290 , P1_U3065 , P1_R1117_U76 );
not NOT1_9394 ( P1_R1117_U291 , P1_R1117_U155 );
nand NAND2_9395 ( P1_R1117_U292 , P1_U3977 , P1_R1117_U79 );
nand NAND2_9396 ( P1_R1117_U293 , P1_R1117_U292 , P1_R1117_U155 );
nand NAND2_9397 ( P1_R1117_U294 , P1_U3058 , P1_R1117_U78 );
not NOT1_9398 ( P1_R1117_U295 , P1_R1117_U87 );
nand NAND2_9399 ( P1_R1117_U296 , P1_U3975 , P1_R1117_U83 );
nand NAND3_9400 ( P1_R1117_U297 , P1_R1117_U87 , P1_R1117_U177 , P1_R1117_U296 );
nand NAND2_9401 ( P1_R1117_U298 , P1_R1117_U83 , P1_R1117_U82 );
nand NAND2_9402 ( P1_R1117_U299 , P1_R1117_U298 , P1_R1117_U80 );
nand NAND2_9403 ( P1_R1117_U300 , P1_U3053 , P1_R1117_U171 );
not NOT1_9404 ( P1_R1117_U301 , P1_R1117_U86 );
nand NAND2_9405 ( P1_R1117_U302 , P1_U3054 , P1_R1117_U84 );
nand NAND2_9406 ( P1_R1117_U303 , P1_R1117_U301 , P1_R1117_U302 );
nand NAND2_9407 ( P1_R1117_U304 , P1_U3974 , P1_R1117_U85 );
nand NAND2_9408 ( P1_R1117_U305 , P1_U3974 , P1_R1117_U85 );
nand NAND2_9409 ( P1_R1117_U306 , P1_R1117_U305 , P1_R1117_U86 );
nand NAND2_9410 ( P1_R1117_U307 , P1_U3054 , P1_R1117_U84 );
nand NAND3_9411 ( P1_R1117_U308 , P1_R1117_U307 , P1_R1117_U306 , P1_R1117_U153 );
nand NAND2_9412 ( P1_R1117_U309 , P1_R1117_U295 , P1_R1117_U82 );
nand NAND2_9413 ( P1_R1117_U310 , P1_R1117_U129 , P1_R1117_U309 );
nand NAND2_9414 ( P1_R1117_U311 , P1_R1117_U87 , P1_R1117_U177 );
nand NAND2_9415 ( P1_R1117_U312 , P1_R1117_U128 , P1_R1117_U311 );
nand NAND2_9416 ( P1_R1117_U313 , P1_R1117_U82 , P1_R1117_U177 );
nand NAND2_9417 ( P1_R1117_U314 , P1_R1117_U283 , P1_R1117_U159 );
not NOT1_9418 ( P1_R1117_U315 , P1_R1117_U88 );
nand NAND2_9419 ( P1_R1117_U316 , P1_U3061 , P1_R1117_U45 );
nand NAND2_9420 ( P1_R1117_U317 , P1_R1117_U315 , P1_R1117_U316 );
nand NAND2_9421 ( P1_R1117_U318 , P1_R1117_U132 , P1_R1117_U317 );
nand NAND2_9422 ( P1_R1117_U319 , P1_R1117_U88 , P1_R1117_U176 );
nand NAND2_9423 ( P1_R1117_U320 , P1_U3979 , P1_R1117_U72 );
nand NAND3_9424 ( P1_R1117_U321 , P1_R1117_U320 , P1_R1117_U319 , P1_R1117_U9 );
nand NAND2_9425 ( P1_R1117_U322 , P1_U3061 , P1_R1117_U45 );
nand NAND2_9426 ( P1_R1117_U323 , P1_R1117_U176 , P1_R1117_U322 );
nand NAND2_9427 ( P1_R1117_U324 , P1_R1117_U283 , P1_R1117_U75 );
nand NAND2_9428 ( P1_R1117_U325 , P1_R1117_U257 , P1_R1117_U167 );
not NOT1_9429 ( P1_R1117_U326 , P1_R1117_U89 );
nand NAND2_9430 ( P1_R1117_U327 , P1_U3074 , P1_R1117_U46 );
nand NAND2_9431 ( P1_R1117_U328 , P1_R1117_U326 , P1_R1117_U327 );
nand NAND2_9432 ( P1_R1117_U329 , P1_R1117_U139 , P1_R1117_U328 );
nand NAND2_9433 ( P1_R1117_U330 , P1_R1117_U89 , P1_R1117_U175 );
nand NAND2_9434 ( P1_R1117_U331 , P1_U3500 , P1_R1117_U58 );
nand NAND2_9435 ( P1_R1117_U332 , P1_R1117_U138 , P1_R1117_U330 );
nand NAND2_9436 ( P1_R1117_U333 , P1_U3074 , P1_R1117_U46 );
nand NAND2_9437 ( P1_R1117_U334 , P1_R1117_U175 , P1_R1117_U333 );
nand NAND2_9438 ( P1_R1117_U335 , P1_R1117_U257 , P1_R1117_U61 );
nand NAND2_9439 ( P1_R1117_U336 , P1_R1117_U212 , P1_R1117_U145 );
not NOT1_9440 ( P1_R1117_U337 , P1_R1117_U90 );
nand NAND2_9441 ( P1_R1117_U338 , P1_U3062 , P1_R1117_U47 );
nand NAND2_9442 ( P1_R1117_U339 , P1_R1117_U337 , P1_R1117_U338 );
nand NAND2_9443 ( P1_R1117_U340 , P1_R1117_U143 , P1_R1117_U339 );
nand NAND2_9444 ( P1_R1117_U341 , P1_R1117_U90 , P1_R1117_U174 );
nand NAND2_9445 ( P1_R1117_U342 , P1_U3485 , P1_R1117_U49 );
nand NAND2_9446 ( P1_R1117_U343 , P1_R1117_U142 , P1_R1117_U341 );
nand NAND2_9447 ( P1_R1117_U344 , P1_U3062 , P1_R1117_U47 );
nand NAND2_9448 ( P1_R1117_U345 , P1_R1117_U174 , P1_R1117_U344 );
nand NAND2_9449 ( P1_R1117_U346 , P1_U3077 , P1_R1117_U22 );
nand NAND3_9450 ( P1_R1117_U347 , P1_R1117_U304 , P1_R1117_U303 , P1_R1117_U385 );
nand NAND2_9451 ( P1_R1117_U348 , P1_U3479 , P1_R1117_U40 );
nand NAND2_9452 ( P1_R1117_U349 , P1_U3083 , P1_R1117_U39 );
nand NAND2_9453 ( P1_R1117_U350 , P1_R1117_U213 , P1_R1117_U145 );
nand NAND2_9454 ( P1_R1117_U351 , P1_R1117_U211 , P1_R1117_U144 );
nand NAND2_9455 ( P1_R1117_U352 , P1_U3476 , P1_R1117_U38 );
nand NAND2_9456 ( P1_R1117_U353 , P1_U3084 , P1_R1117_U35 );
nand NAND2_9457 ( P1_R1117_U354 , P1_U3476 , P1_R1117_U38 );
nand NAND2_9458 ( P1_R1117_U355 , P1_U3084 , P1_R1117_U35 );
nand NAND2_9459 ( P1_R1117_U356 , P1_R1117_U355 , P1_R1117_U354 );
nand NAND2_9460 ( P1_R1117_U357 , P1_U3473 , P1_R1117_U36 );
nand NAND2_9461 ( P1_R1117_U358 , P1_U3070 , P1_R1117_U19 );
nand NAND2_9462 ( P1_R1117_U359 , P1_R1117_U218 , P1_R1117_U41 );
nand NAND2_9463 ( P1_R1117_U360 , P1_R1117_U146 , P1_R1117_U205 );
nand NAND2_9464 ( P1_R1117_U361 , P1_U3470 , P1_R1117_U31 );
nand NAND2_9465 ( P1_R1117_U362 , P1_U3071 , P1_R1117_U29 );
nand NAND2_9466 ( P1_R1117_U363 , P1_R1117_U362 , P1_R1117_U361 );
nand NAND2_9467 ( P1_R1117_U364 , P1_U3467 , P1_R1117_U32 );
nand NAND2_9468 ( P1_R1117_U365 , P1_U3067 , P1_R1117_U20 );
nand NAND2_9469 ( P1_R1117_U366 , P1_R1117_U228 , P1_R1117_U42 );
nand NAND2_9470 ( P1_R1117_U367 , P1_R1117_U147 , P1_R1117_U220 );
nand NAND2_9471 ( P1_R1117_U368 , P1_U3464 , P1_R1117_U33 );
nand NAND2_9472 ( P1_R1117_U369 , P1_U3060 , P1_R1117_U30 );
nand NAND2_9473 ( P1_R1117_U370 , P1_R1117_U229 , P1_R1117_U149 );
nand NAND2_9474 ( P1_R1117_U371 , P1_R1117_U195 , P1_R1117_U148 );
nand NAND2_9475 ( P1_R1117_U372 , P1_U3461 , P1_R1117_U28 );
nand NAND2_9476 ( P1_R1117_U373 , P1_U3064 , P1_R1117_U25 );
nand NAND2_9477 ( P1_R1117_U374 , P1_U3461 , P1_R1117_U28 );
nand NAND2_9478 ( P1_R1117_U375 , P1_U3064 , P1_R1117_U25 );
nand NAND2_9479 ( P1_R1117_U376 , P1_R1117_U375 , P1_R1117_U374 );
nand NAND2_9480 ( P1_R1117_U377 , P1_U3458 , P1_R1117_U26 );
nand NAND2_9481 ( P1_R1117_U378 , P1_U3068 , P1_R1117_U21 );
nand NAND2_9482 ( P1_R1117_U379 , P1_R1117_U234 , P1_R1117_U43 );
nand NAND2_9483 ( P1_R1117_U380 , P1_R1117_U150 , P1_R1117_U189 );
nand NAND2_9484 ( P1_R1117_U381 , P1_U3985 , P1_R1117_U152 );
nand NAND2_9485 ( P1_R1117_U382 , P1_U3055 , P1_R1117_U151 );
nand NAND2_9486 ( P1_R1117_U383 , P1_U3985 , P1_R1117_U152 );
nand NAND2_9487 ( P1_R1117_U384 , P1_U3055 , P1_R1117_U151 );
nand NAND2_9488 ( P1_R1117_U385 , P1_R1117_U384 , P1_R1117_U383 );
nand NAND2_9489 ( P1_R1117_U386 , P1_U3974 , P1_R1117_U85 );
nand NAND2_9490 ( P1_R1117_U387 , P1_U3054 , P1_R1117_U84 );
not NOT1_9491 ( P1_R1117_U388 , P1_R1117_U127 );
nand NAND2_9492 ( P1_R1117_U389 , P1_R1117_U388 , P1_R1117_U301 );
nand NAND2_9493 ( P1_R1117_U390 , P1_R1117_U127 , P1_R1117_U86 );
nand NAND2_9494 ( P1_R1117_U391 , P1_U3975 , P1_R1117_U83 );
nand NAND2_9495 ( P1_R1117_U392 , P1_U3053 , P1_R1117_U80 );
nand NAND2_9496 ( P1_R1117_U393 , P1_U3975 , P1_R1117_U83 );
nand NAND2_9497 ( P1_R1117_U394 , P1_U3053 , P1_R1117_U80 );
nand NAND2_9498 ( P1_R1117_U395 , P1_R1117_U394 , P1_R1117_U393 );
nand NAND2_9499 ( P1_R1117_U396 , P1_U3976 , P1_R1117_U81 );
nand NAND2_9500 ( P1_R1117_U397 , P1_U3057 , P1_R1117_U44 );
nand NAND2_9501 ( P1_R1117_U398 , P1_R1117_U313 , P1_R1117_U87 );
nand NAND2_9502 ( P1_R1117_U399 , P1_R1117_U154 , P1_R1117_U295 );
nand NAND2_9503 ( P1_R1117_U400 , P1_U3977 , P1_R1117_U79 );
nand NAND2_9504 ( P1_R1117_U401 , P1_U3058 , P1_R1117_U78 );
not NOT1_9505 ( P1_R1117_U402 , P1_R1117_U130 );
nand NAND2_9506 ( P1_R1117_U403 , P1_R1117_U291 , P1_R1117_U402 );
nand NAND2_9507 ( P1_R1117_U404 , P1_R1117_U130 , P1_R1117_U155 );
nand NAND2_9508 ( P1_R1117_U405 , P1_U3978 , P1_R1117_U77 );
nand NAND2_9509 ( P1_R1117_U406 , P1_U3065 , P1_R1117_U76 );
not NOT1_9510 ( P1_R1117_U407 , P1_R1117_U131 );
nand NAND2_9511 ( P1_R1117_U408 , P1_R1117_U287 , P1_R1117_U407 );
nand NAND2_9512 ( P1_R1117_U409 , P1_R1117_U131 , P1_R1117_U156 );
nand NAND2_9513 ( P1_R1117_U410 , P1_U3979 , P1_R1117_U72 );
nand NAND2_9514 ( P1_R1117_U411 , P1_U3066 , P1_R1117_U70 );
nand NAND2_9515 ( P1_R1117_U412 , P1_R1117_U411 , P1_R1117_U410 );
nand NAND2_9516 ( P1_R1117_U413 , P1_U3980 , P1_R1117_U73 );
nand NAND2_9517 ( P1_R1117_U414 , P1_U3061 , P1_R1117_U45 );
nand NAND2_9518 ( P1_R1117_U415 , P1_R1117_U323 , P1_R1117_U88 );
nand NAND2_9519 ( P1_R1117_U416 , P1_R1117_U157 , P1_R1117_U315 );
nand NAND2_9520 ( P1_R1117_U417 , P1_U3981 , P1_R1117_U74 );
nand NAND2_9521 ( P1_R1117_U418 , P1_U3075 , P1_R1117_U71 );
nand NAND2_9522 ( P1_R1117_U419 , P1_R1117_U324 , P1_R1117_U159 );
nand NAND2_9523 ( P1_R1117_U420 , P1_R1117_U277 , P1_R1117_U158 );
nand NAND2_9524 ( P1_R1117_U421 , P1_U3982 , P1_R1117_U69 );
nand NAND2_9525 ( P1_R1117_U422 , P1_U3076 , P1_R1117_U68 );
not NOT1_9526 ( P1_R1117_U423 , P1_R1117_U133 );
nand NAND2_9527 ( P1_R1117_U424 , P1_R1117_U273 , P1_R1117_U423 );
nand NAND2_9528 ( P1_R1117_U425 , P1_R1117_U133 , P1_R1117_U160 );
nand NAND2_9529 ( P1_R1117_U426 , P1_R1117_U185 , P1_R1117_U24 );
nand NAND2_9530 ( P1_R1117_U427 , P1_U3078 , P1_R1117_U23 );
not NOT1_9531 ( P1_R1117_U428 , P1_R1117_U134 );
nand NAND2_9532 ( P1_R1117_U429 , P1_U3455 , P1_R1117_U428 );
nand NAND2_9533 ( P1_R1117_U430 , P1_R1117_U134 , P1_R1117_U161 );
nand NAND2_9534 ( P1_R1117_U431 , P1_U3508 , P1_R1117_U67 );
nand NAND2_9535 ( P1_R1117_U432 , P1_U3081 , P1_R1117_U66 );
not NOT1_9536 ( P1_R1117_U433 , P1_R1117_U135 );
nand NAND2_9537 ( P1_R1117_U434 , P1_R1117_U269 , P1_R1117_U433 );
nand NAND2_9538 ( P1_R1117_U435 , P1_R1117_U135 , P1_R1117_U162 );
nand NAND2_9539 ( P1_R1117_U436 , P1_U3506 , P1_R1117_U65 );
nand NAND2_9540 ( P1_R1117_U437 , P1_U3082 , P1_R1117_U163 );
not NOT1_9541 ( P1_R1117_U438 , P1_R1117_U136 );
nand NAND2_9542 ( P1_R1117_U439 , P1_R1117_U438 , P1_R1117_U265 );
nand NAND2_9543 ( P1_R1117_U440 , P1_R1117_U136 , P1_R1117_U64 );
nand NAND2_9544 ( P1_R1117_U441 , P1_U3503 , P1_R1117_U63 );
nand NAND2_9545 ( P1_R1117_U442 , P1_U3069 , P1_R1117_U62 );
not NOT1_9546 ( P1_R1117_U443 , P1_R1117_U137 );
nand NAND2_9547 ( P1_R1117_U444 , P1_R1117_U261 , P1_R1117_U443 );
nand NAND2_9548 ( P1_R1117_U445 , P1_R1117_U137 , P1_R1117_U164 );
nand NAND2_9549 ( P1_R1117_U446 , P1_U3500 , P1_R1117_U58 );
nand NAND2_9550 ( P1_R1117_U447 , P1_U3073 , P1_R1117_U56 );
nand NAND2_9551 ( P1_R1117_U448 , P1_R1117_U447 , P1_R1117_U446 );
nand NAND2_9552 ( P1_R1117_U449 , P1_U3497 , P1_R1117_U59 );
nand NAND2_9553 ( P1_R1117_U450 , P1_U3074 , P1_R1117_U46 );
nand NAND2_9554 ( P1_R1117_U451 , P1_R1117_U334 , P1_R1117_U89 );
nand NAND2_9555 ( P1_R1117_U452 , P1_R1117_U165 , P1_R1117_U326 );
nand NAND2_9556 ( P1_R1117_U453 , P1_U3494 , P1_R1117_U60 );
nand NAND2_9557 ( P1_R1117_U454 , P1_U3079 , P1_R1117_U57 );
nand NAND2_9558 ( P1_R1117_U455 , P1_R1117_U335 , P1_R1117_U167 );
nand NAND2_9559 ( P1_R1117_U456 , P1_R1117_U251 , P1_R1117_U166 );
nand NAND2_9560 ( P1_R1117_U457 , P1_U3491 , P1_R1117_U55 );
nand NAND2_9561 ( P1_R1117_U458 , P1_U3080 , P1_R1117_U54 );
not NOT1_9562 ( P1_R1117_U459 , P1_R1117_U140 );
nand NAND2_9563 ( P1_R1117_U460 , P1_R1117_U247 , P1_R1117_U459 );
nand NAND2_9564 ( P1_R1117_U461 , P1_R1117_U140 , P1_R1117_U168 );
nand NAND2_9565 ( P1_R1117_U462 , P1_U3488 , P1_R1117_U53 );
nand NAND2_9566 ( P1_R1117_U463 , P1_U3072 , P1_R1117_U52 );
not NOT1_9567 ( P1_R1117_U464 , P1_R1117_U141 );
nand NAND2_9568 ( P1_R1117_U465 , P1_R1117_U243 , P1_R1117_U464 );
nand NAND2_9569 ( P1_R1117_U466 , P1_R1117_U141 , P1_R1117_U169 );
nand NAND2_9570 ( P1_R1117_U467 , P1_U3485 , P1_R1117_U49 );
nand NAND2_9571 ( P1_R1117_U468 , P1_U3063 , P1_R1117_U48 );
nand NAND2_9572 ( P1_R1117_U469 , P1_R1117_U468 , P1_R1117_U467 );
nand NAND2_9573 ( P1_R1117_U470 , P1_U3482 , P1_R1117_U50 );
nand NAND2_9574 ( P1_R1117_U471 , P1_U3062 , P1_R1117_U47 );
nand NAND2_9575 ( P1_R1117_U472 , P1_R1117_U345 , P1_R1117_U90 );
nand NAND2_9576 ( P1_R1117_U473 , P1_R1117_U170 , P1_R1117_U337 );
and AND2_9577 ( P1_R1375_U6 , P1_R1375_U119 , P1_R1375_U120 );
and AND2_9578 ( P1_R1375_U7 , P1_R1375_U137 , P1_R1375_U136 );
and AND4_9579 ( P1_R1375_U8 , P1_R1375_U144 , P1_R1375_U143 , P1_R1375_U142 , P1_R1375_U141 );
and AND2_9580 ( P1_R1375_U9 , P1_R1375_U164 , P1_R1375_U163 );
and AND4_9581 ( P1_R1375_U10 , P1_R1375_U197 , P1_R1375_U196 , P1_R1375_U198 , P1_R1375_U6 );
and AND2_9582 ( P1_R1375_U11 , P1_U3985 , P1_R1375_U20 );
and AND4_9583 ( P1_R1375_U12 , P1_R1375_U207 , P1_R1375_U206 , P1_R1375_U118 , P1_R1375_U117 );
and AND2_9584 ( P1_R1375_U13 , P1_U3450 , P1_R1375_U48 );
and AND3_9585 ( P1_R1375_U14 , P1_R1375_U205 , P1_R1375_U115 , P1_R1375_U204 );
not NOT1_9586 ( P1_R1375_U15 , P1_U3983 );
not NOT1_9587 ( P1_R1375_U16 , P1_U3984 );
not NOT1_9588 ( P1_R1375_U17 , P1_U3056 );
not NOT1_9589 ( P1_R1375_U18 , P1_U3985 );
not NOT1_9590 ( P1_R1375_U19 , P1_U3059 );
not NOT1_9591 ( P1_R1375_U20 , P1_U3055 );
not NOT1_9592 ( P1_R1375_U21 , P1_U3054 );
not NOT1_9593 ( P1_R1375_U22 , P1_U3975 );
not NOT1_9594 ( P1_R1375_U23 , P1_U3057 );
not NOT1_9595 ( P1_R1375_U24 , P1_U3977 );
not NOT1_9596 ( P1_R1375_U25 , P1_U3974 );
not NOT1_9597 ( P1_R1375_U26 , P1_U3976 );
not NOT1_9598 ( P1_R1375_U27 , P1_U3978 );
not NOT1_9599 ( P1_R1375_U28 , P1_U3066 );
not NOT1_9600 ( P1_R1375_U29 , P1_U3979 );
not NOT1_9601 ( P1_R1375_U30 , P1_U3061 );
not NOT1_9602 ( P1_R1375_U31 , P1_U3058 );
not NOT1_9603 ( P1_R1375_U32 , P1_U3065 );
not NOT1_9604 ( P1_R1375_U33 , P1_U3075 );
not NOT1_9605 ( P1_R1375_U34 , P1_U3076 );
not NOT1_9606 ( P1_R1375_U35 , P1_U3503 );
not NOT1_9607 ( P1_R1375_U36 , P1_U3506 );
not NOT1_9608 ( P1_R1375_U37 , P1_U3074 );
not NOT1_9609 ( P1_R1375_U38 , P1_U3079 );
not NOT1_9610 ( P1_R1375_U39 , P1_U3470 );
not NOT1_9611 ( P1_R1375_U40 , P1_U3067 );
not NOT1_9612 ( P1_R1375_U41 , P1_U3083 );
not NOT1_9613 ( P1_R1375_U42 , P1_U3084 );
not NOT1_9614 ( P1_R1375_U43 , P1_U3071 );
not NOT1_9615 ( P1_R1375_U44 , P1_U3070 );
not NOT1_9616 ( P1_R1375_U45 , P1_U3060 );
not NOT1_9617 ( P1_R1375_U46 , P1_U3064 );
not NOT1_9618 ( P1_R1375_U47 , P1_U3450 );
not NOT1_9619 ( P1_R1375_U48 , P1_U3077 );
nand NAND2_9620 ( P1_R1375_U49 , P1_R1375_U147 , P1_R1375_U146 );
not NOT1_9621 ( P1_R1375_U50 , P1_U3455 );
not NOT1_9622 ( P1_R1375_U51 , P1_U3068 );
not NOT1_9623 ( P1_R1375_U52 , P1_U3485 );
not NOT1_9624 ( P1_R1375_U53 , P1_U3488 );
not NOT1_9625 ( P1_R1375_U54 , P1_U3458 );
not NOT1_9626 ( P1_R1375_U55 , P1_U3461 );
not NOT1_9627 ( P1_R1375_U56 , P1_U3467 );
not NOT1_9628 ( P1_R1375_U57 , P1_U3464 );
not NOT1_9629 ( P1_R1375_U58 , P1_U3473 );
not NOT1_9630 ( P1_R1375_U59 , P1_U3476 );
not NOT1_9631 ( P1_R1375_U60 , P1_U3479 );
not NOT1_9632 ( P1_R1375_U61 , P1_U3482 );
not NOT1_9633 ( P1_R1375_U62 , P1_U3062 );
not NOT1_9634 ( P1_R1375_U63 , P1_U3072 );
not NOT1_9635 ( P1_R1375_U64 , P1_U3063 );
not NOT1_9636 ( P1_R1375_U65 , P1_U3080 );
not NOT1_9637 ( P1_R1375_U66 , P1_U3491 );
not NOT1_9638 ( P1_R1375_U67 , P1_U3494 );
not NOT1_9639 ( P1_R1375_U68 , P1_U3497 );
not NOT1_9640 ( P1_R1375_U69 , P1_U3500 );
not NOT1_9641 ( P1_R1375_U70 , P1_U3073 );
not NOT1_9642 ( P1_R1375_U71 , P1_U3069 );
not NOT1_9643 ( P1_R1375_U72 , P1_U3082 );
not NOT1_9644 ( P1_R1375_U73 , P1_U3081 );
not NOT1_9645 ( P1_R1375_U74 , P1_U3508 );
not NOT1_9646 ( P1_R1375_U75 , P1_U3982 );
not NOT1_9647 ( P1_R1375_U76 , P1_U3981 );
not NOT1_9648 ( P1_R1375_U77 , P1_U3980 );
nand NAND2_9649 ( P1_R1375_U78 , P1_R1375_U11 , P1_R1375_U125 );
nand NAND4_9650 ( P1_R1375_U79 , P1_R1375_U124 , P1_R1375_U122 , P1_R1375_U87 , P1_R1375_U12 );
nand NAND2_9651 ( P1_R1375_U80 , P1_R1375_U109 , P1_R1375_U195 );
and AND2_9652 ( P1_R1375_U81 , P1_U3975 , P1_R1375_U113 );
and AND2_9653 ( P1_R1375_U82 , P1_U3977 , P1_R1375_U31 );
and AND2_9654 ( P1_R1375_U83 , P1_U3974 , P1_R1375_U21 );
and AND2_9655 ( P1_R1375_U84 , P1_U3976 , P1_R1375_U23 );
and AND2_9656 ( P1_R1375_U85 , P1_U3066 , P1_R1375_U29 );
and AND2_9657 ( P1_R1375_U86 , P1_U3061 , P1_R1375_U77 );
and AND2_9658 ( P1_R1375_U87 , P1_R1375_U123 , P1_R1375_U121 );
and AND2_9659 ( P1_R1375_U88 , P1_R1375_U129 , P1_R1375_U126 );
and AND3_9660 ( P1_R1375_U89 , P1_R1375_U131 , P1_R1375_U201 , P1_R1375_U128 );
and AND2_9661 ( P1_R1375_U90 , P1_U3067 , P1_R1375_U56 );
and AND2_9662 ( P1_R1375_U91 , P1_R1375_U145 , P1_R1375_U149 );
and AND2_9663 ( P1_R1375_U92 , P1_R1375_U91 , P1_R1375_U140 );
and AND3_9664 ( P1_R1375_U93 , P1_R1375_U153 , P1_R1375_U152 , P1_R1375_U8 );
and AND2_9665 ( P1_R1375_U94 , P1_U3458 , P1_R1375_U51 );
and AND3_9666 ( P1_R1375_U95 , P1_R1375_U161 , P1_R1375_U160 , P1_R1375_U159 );
and AND2_9667 ( P1_R1375_U96 , P1_U3473 , P1_R1375_U44 );
and AND2_9668 ( P1_R1375_U97 , P1_R1375_U171 , P1_R1375_U170 );
and AND2_9669 ( P1_R1375_U98 , P1_R1375_U97 , P1_R1375_U9 );
and AND2_9670 ( P1_R1375_U99 , P1_U3062 , P1_R1375_U61 );
and AND2_9671 ( P1_R1375_U100 , P1_U3063 , P1_R1375_U52 );
and AND3_9672 ( P1_R1375_U101 , P1_R1375_U173 , P1_R1375_U174 , P1_R1375_U102 );
and AND2_9673 ( P1_R1375_U102 , P1_R1375_U177 , P1_R1375_U176 );
and AND2_9674 ( P1_R1375_U103 , P1_R1375_U7 , P1_R1375_U104 );
and AND2_9675 ( P1_R1375_U104 , P1_R1375_U185 , P1_R1375_U186 );
and AND2_9676 ( P1_R1375_U105 , P1_U3073 , P1_R1375_U69 );
and AND2_9677 ( P1_R1375_U106 , P1_U3069 , P1_R1375_U35 );
and AND3_9678 ( P1_R1375_U107 , P1_R1375_U188 , P1_R1375_U190 , P1_R1375_U108 );
and AND2_9679 ( P1_R1375_U108 , P1_R1375_U192 , P1_R1375_U191 );
and AND2_9680 ( P1_R1375_U109 , P1_R1375_U134 , P1_R1375_U133 );
and AND2_9681 ( P1_R1375_U110 , P1_U3982 , P1_R1375_U34 );
and AND2_9682 ( P1_R1375_U111 , P1_R1375_U128 , P1_R1375_U127 );
and AND4_9683 ( P1_R1375_U112 , P1_R1375_U10 , P1_R1375_U131 , P1_R1375_U129 , P1_R1375_U130 );
not NOT1_9684 ( P1_R1375_U113 , P1_U3053 );
nand NAND2_9685 ( P1_R1375_U114 , P1_R1375_U200 , P1_R1375_U199 );
nand NAND2_9686 ( P1_R1375_U115 , P1_U3983 , P1_R1375_U17 );
nand NAND2_9687 ( P1_R1375_U116 , P1_U3055 , P1_R1375_U18 );
nand NAND2_9688 ( P1_R1375_U117 , P1_U3054 , P1_R1375_U25 );
nand NAND2_9689 ( P1_R1375_U118 , P1_U3057 , P1_R1375_U26 );
nand NAND2_9690 ( P1_R1375_U119 , P1_U3978 , P1_R1375_U32 );
nand NAND2_9691 ( P1_R1375_U120 , P1_U3979 , P1_R1375_U28 );
nand NAND2_9692 ( P1_R1375_U121 , P1_R1375_U85 , P1_R1375_U119 );
nand NAND2_9693 ( P1_R1375_U122 , P1_R1375_U86 , P1_R1375_U6 );
nand NAND2_9694 ( P1_R1375_U123 , P1_U3058 , P1_R1375_U24 );
nand NAND2_9695 ( P1_R1375_U124 , P1_U3065 , P1_R1375_U27 );
nand NAND2_9696 ( P1_R1375_U125 , P1_U3059 , P1_R1375_U16 );
nand NAND3_9697 ( P1_R1375_U126 , P1_R1375_U81 , P1_R1375_U117 , P1_R1375_U115 );
nand NAND3_9698 ( P1_R1375_U127 , P1_R1375_U82 , P1_R1375_U12 , P1_R1375_U115 );
nand NAND3_9699 ( P1_R1375_U128 , P1_R1375_U115 , P1_R1375_U19 , P1_U3984 );
nand NAND2_9700 ( P1_R1375_U129 , P1_R1375_U83 , P1_R1375_U115 );
nand NAND3_9701 ( P1_R1375_U130 , P1_R1375_U84 , P1_R1375_U12 , P1_R1375_U115 );
nand NAND2_9702 ( P1_R1375_U131 , P1_U3056 , P1_R1375_U15 );
nand NAND4_9703 ( P1_R1375_U132 , P1_R1375_U79 , P1_R1375_U130 , P1_R1375_U88 , P1_R1375_U127 );
nand NAND2_9704 ( P1_R1375_U133 , P1_U3075 , P1_R1375_U76 );
nand NAND2_9705 ( P1_R1375_U134 , P1_U3076 , P1_R1375_U75 );
nand NAND2_9706 ( P1_R1375_U135 , P1_U3074 , P1_R1375_U68 );
nand NAND2_9707 ( P1_R1375_U136 , P1_U3503 , P1_R1375_U71 );
nand NAND2_9708 ( P1_R1375_U137 , P1_U3506 , P1_R1375_U72 );
nand NAND2_9709 ( P1_R1375_U138 , P1_U3079 , P1_R1375_U67 );
nand NAND2_9710 ( P1_R1375_U139 , P1_U3470 , P1_R1375_U43 );
nand NAND2_9711 ( P1_R1375_U140 , P1_R1375_U90 , P1_R1375_U139 );
nand NAND2_9712 ( P1_R1375_U141 , P1_U3083 , P1_R1375_U60 );
nand NAND2_9713 ( P1_R1375_U142 , P1_U3084 , P1_R1375_U59 );
nand NAND2_9714 ( P1_R1375_U143 , P1_U3071 , P1_R1375_U39 );
nand NAND2_9715 ( P1_R1375_U144 , P1_U3070 , P1_R1375_U58 );
nand NAND2_9716 ( P1_R1375_U145 , P1_U3060 , P1_R1375_U57 );
or OR2_9717 ( P1_R1375_U146 , P1_U3447 , P1_R1375_U13 );
nand NAND2_9718 ( P1_R1375_U147 , P1_U3077 , P1_R1375_U47 );
not NOT1_9719 ( P1_R1375_U148 , P1_R1375_U49 );
nand NAND2_9720 ( P1_R1375_U149 , P1_U3064 , P1_R1375_U55 );
nand NAND2_9721 ( P1_R1375_U150 , P1_U3455 , P1_R1375_U148 );
nand NAND2_9722 ( P1_R1375_U151 , P1_U3078 , P1_R1375_U150 );
nand NAND2_9723 ( P1_R1375_U152 , P1_R1375_U49 , P1_R1375_U50 );
nand NAND2_9724 ( P1_R1375_U153 , P1_U3068 , P1_R1375_U54 );
nand NAND3_9725 ( P1_R1375_U154 , P1_R1375_U92 , P1_R1375_U151 , P1_R1375_U93 );
nand NAND2_9726 ( P1_R1375_U155 , P1_R1375_U94 , P1_R1375_U149 );
nand NAND2_9727 ( P1_R1375_U156 , P1_U3461 , P1_R1375_U46 );
nand NAND2_9728 ( P1_R1375_U157 , P1_R1375_U156 , P1_R1375_U155 );
nand NAND2_9729 ( P1_R1375_U158 , P1_R1375_U157 , P1_R1375_U145 );
nand NAND2_9730 ( P1_R1375_U159 , P1_U3467 , P1_R1375_U40 );
nand NAND2_9731 ( P1_R1375_U160 , P1_U3464 , P1_R1375_U45 );
nand NAND2_9732 ( P1_R1375_U161 , P1_U3470 , P1_R1375_U43 );
nand NAND2_9733 ( P1_R1375_U162 , P1_R1375_U158 , P1_R1375_U95 );
nand NAND2_9734 ( P1_R1375_U163 , P1_U3485 , P1_R1375_U64 );
nand NAND2_9735 ( P1_R1375_U164 , P1_U3488 , P1_R1375_U63 );
nand NAND2_9736 ( P1_R1375_U165 , P1_R1375_U96 , P1_R1375_U142 );
nand NAND2_9737 ( P1_R1375_U166 , P1_U3476 , P1_R1375_U42 );
nand NAND2_9738 ( P1_R1375_U167 , P1_R1375_U166 , P1_R1375_U165 );
nand NAND3_9739 ( P1_R1375_U168 , P1_R1375_U162 , P1_R1375_U140 , P1_R1375_U8 );
nand NAND2_9740 ( P1_R1375_U169 , P1_R1375_U167 , P1_R1375_U141 );
nand NAND2_9741 ( P1_R1375_U170 , P1_U3479 , P1_R1375_U41 );
nand NAND2_9742 ( P1_R1375_U171 , P1_U3482 , P1_R1375_U62 );
nand NAND4_9743 ( P1_R1375_U172 , P1_R1375_U168 , P1_R1375_U169 , P1_R1375_U98 , P1_R1375_U154 );
nand NAND2_9744 ( P1_R1375_U173 , P1_R1375_U99 , P1_R1375_U9 );
nand NAND2_9745 ( P1_R1375_U174 , P1_U3072 , P1_R1375_U53 );
nand NAND2_9746 ( P1_R1375_U175 , P1_U3488 , P1_R1375_U63 );
nand NAND2_9747 ( P1_R1375_U176 , P1_R1375_U100 , P1_R1375_U175 );
nand NAND2_9748 ( P1_R1375_U177 , P1_U3080 , P1_R1375_U66 );
nand NAND2_9749 ( P1_R1375_U178 , P1_R1375_U172 , P1_R1375_U101 );
nand NAND2_9750 ( P1_R1375_U179 , P1_U3491 , P1_R1375_U65 );
nand NAND2_9751 ( P1_R1375_U180 , P1_R1375_U179 , P1_R1375_U178 );
nand NAND2_9752 ( P1_R1375_U181 , P1_R1375_U180 , P1_R1375_U138 );
nand NAND2_9753 ( P1_R1375_U182 , P1_U3494 , P1_R1375_U38 );
nand NAND2_9754 ( P1_R1375_U183 , P1_R1375_U182 , P1_R1375_U181 );
nand NAND2_9755 ( P1_R1375_U184 , P1_R1375_U183 , P1_R1375_U135 );
nand NAND2_9756 ( P1_R1375_U185 , P1_U3497 , P1_R1375_U37 );
nand NAND2_9757 ( P1_R1375_U186 , P1_U3500 , P1_R1375_U70 );
nand NAND2_9758 ( P1_R1375_U187 , P1_R1375_U184 , P1_R1375_U103 );
nand NAND2_9759 ( P1_R1375_U188 , P1_R1375_U105 , P1_R1375_U7 );
nand NAND2_9760 ( P1_R1375_U189 , P1_U3506 , P1_R1375_U72 );
nand NAND2_9761 ( P1_R1375_U190 , P1_R1375_U106 , P1_R1375_U189 );
nand NAND2_9762 ( P1_R1375_U191 , P1_U3082 , P1_R1375_U36 );
nand NAND2_9763 ( P1_R1375_U192 , P1_U3081 , P1_R1375_U74 );
nand NAND2_9764 ( P1_R1375_U193 , P1_R1375_U187 , P1_R1375_U107 );
nand NAND2_9765 ( P1_R1375_U194 , P1_U3508 , P1_R1375_U73 );
nand NAND2_9766 ( P1_R1375_U195 , P1_R1375_U194 , P1_R1375_U193 );
nand NAND2_9767 ( P1_R1375_U196 , P1_R1375_U110 , P1_R1375_U133 );
nand NAND2_9768 ( P1_R1375_U197 , P1_U3981 , P1_R1375_U33 );
nand NAND2_9769 ( P1_R1375_U198 , P1_U3980 , P1_R1375_U30 );
nand NAND2_9770 ( P1_R1375_U199 , P1_U3984 , P1_R1375_U116 );
nand NAND2_9771 ( P1_R1375_U200 , P1_R1375_U19 , P1_R1375_U116 );
nand NAND2_9772 ( P1_R1375_U201 , P1_R1375_U11 , P1_R1375_U202 );
nand NAND2_9773 ( P1_R1375_U202 , P1_U3059 , P1_R1375_U16 );
nand NAND2_9774 ( P1_R1375_U203 , P1_R1375_U132 , P1_R1375_U114 );
nand NAND2_9775 ( P1_R1375_U204 , P1_R1375_U89 , P1_R1375_U203 );
nand NAND5_9776 ( P1_R1375_U205 , P1_R1375_U126 , P1_R1375_U80 , P1_R1375_U78 , P1_R1375_U111 , P1_R1375_U112 );
nand NAND2_9777 ( P1_R1375_U206 , P1_U3053 , P1_R1375_U22 );
nand NAND2_9778 ( P1_R1375_U207 , P1_U3975 , P1_R1375_U113 );
and AND2_9779 ( P1_R1352_U6 , P1_U3059 , P1_R1352_U7 );
not NOT1_9780 ( P1_R1352_U7 , P1_U3056 );
and AND2_9781 ( P1_R1207_U6 , P1_R1207_U198 , P1_R1207_U197 );
and AND2_9782 ( P1_R1207_U7 , P1_R1207_U237 , P1_R1207_U236 );
and AND2_9783 ( P1_R1207_U8 , P1_R1207_U254 , P1_R1207_U253 );
and AND2_9784 ( P1_R1207_U9 , P1_R1207_U280 , P1_R1207_U279 );
nand NAND2_9785 ( P1_R1207_U10 , P1_R1207_U340 , P1_R1207_U343 );
nand NAND2_9786 ( P1_R1207_U11 , P1_R1207_U329 , P1_R1207_U332 );
nand NAND2_9787 ( P1_R1207_U12 , P1_R1207_U318 , P1_R1207_U321 );
nand NAND2_9788 ( P1_R1207_U13 , P1_R1207_U310 , P1_R1207_U312 );
nand NAND2_9789 ( P1_R1207_U14 , P1_R1207_U347 , P1_R1207_U308 );
nand NAND2_9790 ( P1_R1207_U15 , P1_R1207_U231 , P1_R1207_U233 );
nand NAND2_9791 ( P1_R1207_U16 , P1_R1207_U223 , P1_R1207_U226 );
nand NAND2_9792 ( P1_R1207_U17 , P1_R1207_U215 , P1_R1207_U217 );
nand NAND2_9793 ( P1_R1207_U18 , P1_R1207_U23 , P1_R1207_U346 );
not NOT1_9794 ( P1_R1207_U19 , P1_U3473 );
not NOT1_9795 ( P1_R1207_U20 , P1_U3467 );
not NOT1_9796 ( P1_R1207_U21 , P1_U3458 );
not NOT1_9797 ( P1_R1207_U22 , P1_U3450 );
nand NAND2_9798 ( P1_R1207_U23 , P1_U3450 , P1_R1207_U91 );
not NOT1_9799 ( P1_R1207_U24 , P1_U3078 );
not NOT1_9800 ( P1_R1207_U25 , P1_U3461 );
not NOT1_9801 ( P1_R1207_U26 , P1_U3068 );
nand NAND2_9802 ( P1_R1207_U27 , P1_U3068 , P1_R1207_U21 );
not NOT1_9803 ( P1_R1207_U28 , P1_U3064 );
not NOT1_9804 ( P1_R1207_U29 , P1_U3470 );
not NOT1_9805 ( P1_R1207_U30 , P1_U3464 );
not NOT1_9806 ( P1_R1207_U31 , P1_U3071 );
not NOT1_9807 ( P1_R1207_U32 , P1_U3067 );
not NOT1_9808 ( P1_R1207_U33 , P1_U3060 );
nand NAND2_9809 ( P1_R1207_U34 , P1_U3060 , P1_R1207_U30 );
not NOT1_9810 ( P1_R1207_U35 , P1_U3476 );
not NOT1_9811 ( P1_R1207_U36 , P1_U3070 );
nand NAND2_9812 ( P1_R1207_U37 , P1_U3070 , P1_R1207_U19 );
not NOT1_9813 ( P1_R1207_U38 , P1_U3084 );
not NOT1_9814 ( P1_R1207_U39 , P1_U3479 );
not NOT1_9815 ( P1_R1207_U40 , P1_U3083 );
nand NAND2_9816 ( P1_R1207_U41 , P1_R1207_U204 , P1_R1207_U203 );
nand NAND2_9817 ( P1_R1207_U42 , P1_R1207_U34 , P1_R1207_U219 );
nand NAND2_9818 ( P1_R1207_U43 , P1_R1207_U188 , P1_R1207_U187 );
not NOT1_9819 ( P1_R1207_U44 , P1_U3976 );
not NOT1_9820 ( P1_R1207_U45 , P1_U3980 );
not NOT1_9821 ( P1_R1207_U46 , P1_U3497 );
not NOT1_9822 ( P1_R1207_U47 , P1_U3482 );
not NOT1_9823 ( P1_R1207_U48 , P1_U3485 );
not NOT1_9824 ( P1_R1207_U49 , P1_U3063 );
not NOT1_9825 ( P1_R1207_U50 , P1_U3062 );
nand NAND2_9826 ( P1_R1207_U51 , P1_U3083 , P1_R1207_U39 );
not NOT1_9827 ( P1_R1207_U52 , P1_U3488 );
not NOT1_9828 ( P1_R1207_U53 , P1_U3072 );
not NOT1_9829 ( P1_R1207_U54 , P1_U3491 );
not NOT1_9830 ( P1_R1207_U55 , P1_U3080 );
not NOT1_9831 ( P1_R1207_U56 , P1_U3500 );
not NOT1_9832 ( P1_R1207_U57 , P1_U3494 );
not NOT1_9833 ( P1_R1207_U58 , P1_U3073 );
not NOT1_9834 ( P1_R1207_U59 , P1_U3074 );
not NOT1_9835 ( P1_R1207_U60 , P1_U3079 );
nand NAND2_9836 ( P1_R1207_U61 , P1_U3079 , P1_R1207_U57 );
not NOT1_9837 ( P1_R1207_U62 , P1_U3503 );
not NOT1_9838 ( P1_R1207_U63 , P1_U3069 );
nand NAND2_9839 ( P1_R1207_U64 , P1_R1207_U264 , P1_R1207_U263 );
not NOT1_9840 ( P1_R1207_U65 , P1_U3082 );
not NOT1_9841 ( P1_R1207_U66 , P1_U3508 );
not NOT1_9842 ( P1_R1207_U67 , P1_U3081 );
not NOT1_9843 ( P1_R1207_U68 , P1_U3982 );
not NOT1_9844 ( P1_R1207_U69 , P1_U3076 );
not NOT1_9845 ( P1_R1207_U70 , P1_U3979 );
not NOT1_9846 ( P1_R1207_U71 , P1_U3981 );
not NOT1_9847 ( P1_R1207_U72 , P1_U3066 );
not NOT1_9848 ( P1_R1207_U73 , P1_U3061 );
not NOT1_9849 ( P1_R1207_U74 , P1_U3075 );
nand NAND2_9850 ( P1_R1207_U75 , P1_U3075 , P1_R1207_U71 );
not NOT1_9851 ( P1_R1207_U76 , P1_U3978 );
not NOT1_9852 ( P1_R1207_U77 , P1_U3065 );
not NOT1_9853 ( P1_R1207_U78 , P1_U3977 );
not NOT1_9854 ( P1_R1207_U79 , P1_U3058 );
not NOT1_9855 ( P1_R1207_U80 , P1_U3975 );
not NOT1_9856 ( P1_R1207_U81 , P1_U3057 );
nand NAND2_9857 ( P1_R1207_U82 , P1_U3057 , P1_R1207_U44 );
not NOT1_9858 ( P1_R1207_U83 , P1_U3053 );
not NOT1_9859 ( P1_R1207_U84 , P1_U3974 );
not NOT1_9860 ( P1_R1207_U85 , P1_U3054 );
nand NAND2_9861 ( P1_R1207_U86 , P1_R1207_U126 , P1_R1207_U297 );
nand NAND2_9862 ( P1_R1207_U87 , P1_R1207_U294 , P1_R1207_U293 );
nand NAND2_9863 ( P1_R1207_U88 , P1_R1207_U75 , P1_R1207_U314 );
nand NAND2_9864 ( P1_R1207_U89 , P1_R1207_U61 , P1_R1207_U325 );
nand NAND2_9865 ( P1_R1207_U90 , P1_R1207_U51 , P1_R1207_U336 );
not NOT1_9866 ( P1_R1207_U91 , P1_U3077 );
nand NAND2_9867 ( P1_R1207_U92 , P1_R1207_U390 , P1_R1207_U389 );
nand NAND2_9868 ( P1_R1207_U93 , P1_R1207_U404 , P1_R1207_U403 );
nand NAND2_9869 ( P1_R1207_U94 , P1_R1207_U409 , P1_R1207_U408 );
nand NAND2_9870 ( P1_R1207_U95 , P1_R1207_U425 , P1_R1207_U424 );
nand NAND2_9871 ( P1_R1207_U96 , P1_R1207_U430 , P1_R1207_U429 );
nand NAND2_9872 ( P1_R1207_U97 , P1_R1207_U435 , P1_R1207_U434 );
nand NAND2_9873 ( P1_R1207_U98 , P1_R1207_U440 , P1_R1207_U439 );
nand NAND2_9874 ( P1_R1207_U99 , P1_R1207_U445 , P1_R1207_U444 );
nand NAND2_9875 ( P1_R1207_U100 , P1_R1207_U461 , P1_R1207_U460 );
nand NAND2_9876 ( P1_R1207_U101 , P1_R1207_U466 , P1_R1207_U465 );
nand NAND2_9877 ( P1_R1207_U102 , P1_R1207_U351 , P1_R1207_U350 );
nand NAND2_9878 ( P1_R1207_U103 , P1_R1207_U360 , P1_R1207_U359 );
nand NAND2_9879 ( P1_R1207_U104 , P1_R1207_U367 , P1_R1207_U366 );
nand NAND2_9880 ( P1_R1207_U105 , P1_R1207_U371 , P1_R1207_U370 );
nand NAND2_9881 ( P1_R1207_U106 , P1_R1207_U380 , P1_R1207_U379 );
nand NAND2_9882 ( P1_R1207_U107 , P1_R1207_U399 , P1_R1207_U398 );
nand NAND2_9883 ( P1_R1207_U108 , P1_R1207_U416 , P1_R1207_U415 );
nand NAND2_9884 ( P1_R1207_U109 , P1_R1207_U420 , P1_R1207_U419 );
nand NAND2_9885 ( P1_R1207_U110 , P1_R1207_U452 , P1_R1207_U451 );
nand NAND2_9886 ( P1_R1207_U111 , P1_R1207_U456 , P1_R1207_U455 );
nand NAND2_9887 ( P1_R1207_U112 , P1_R1207_U473 , P1_R1207_U472 );
and AND2_9888 ( P1_R1207_U113 , P1_R1207_U193 , P1_R1207_U194 );
and AND2_9889 ( P1_R1207_U114 , P1_R1207_U201 , P1_R1207_U196 );
and AND2_9890 ( P1_R1207_U115 , P1_R1207_U206 , P1_R1207_U180 );
and AND2_9891 ( P1_R1207_U116 , P1_R1207_U209 , P1_R1207_U210 );
and AND3_9892 ( P1_R1207_U117 , P1_R1207_U353 , P1_R1207_U352 , P1_R1207_U37 );
and AND2_9893 ( P1_R1207_U118 , P1_R1207_U356 , P1_R1207_U180 );
and AND2_9894 ( P1_R1207_U119 , P1_R1207_U225 , P1_R1207_U6 );
and AND2_9895 ( P1_R1207_U120 , P1_R1207_U363 , P1_R1207_U179 );
and AND3_9896 ( P1_R1207_U121 , P1_R1207_U373 , P1_R1207_U372 , P1_R1207_U27 );
and AND2_9897 ( P1_R1207_U122 , P1_R1207_U376 , P1_R1207_U178 );
and AND3_9898 ( P1_R1207_U123 , P1_R1207_U235 , P1_R1207_U212 , P1_R1207_U174 );
and AND3_9899 ( P1_R1207_U124 , P1_R1207_U257 , P1_R1207_U175 , P1_R1207_U252 );
and AND2_9900 ( P1_R1207_U125 , P1_R1207_U283 , P1_R1207_U176 );
and AND2_9901 ( P1_R1207_U126 , P1_R1207_U299 , P1_R1207_U300 );
nand NAND2_9902 ( P1_R1207_U127 , P1_R1207_U387 , P1_R1207_U386 );
and AND3_9903 ( P1_R1207_U128 , P1_R1207_U392 , P1_R1207_U391 , P1_R1207_U82 );
and AND2_9904 ( P1_R1207_U129 , P1_R1207_U395 , P1_R1207_U177 );
nand NAND2_9905 ( P1_R1207_U130 , P1_R1207_U401 , P1_R1207_U400 );
nand NAND2_9906 ( P1_R1207_U131 , P1_R1207_U406 , P1_R1207_U405 );
and AND2_9907 ( P1_R1207_U132 , P1_R1207_U412 , P1_R1207_U176 );
nand NAND2_9908 ( P1_R1207_U133 , P1_R1207_U422 , P1_R1207_U421 );
nand NAND2_9909 ( P1_R1207_U134 , P1_R1207_U427 , P1_R1207_U426 );
nand NAND2_9910 ( P1_R1207_U135 , P1_R1207_U432 , P1_R1207_U431 );
nand NAND2_9911 ( P1_R1207_U136 , P1_R1207_U437 , P1_R1207_U436 );
nand NAND2_9912 ( P1_R1207_U137 , P1_R1207_U442 , P1_R1207_U441 );
and AND2_9913 ( P1_R1207_U138 , P1_R1207_U331 , P1_R1207_U8 );
and AND2_9914 ( P1_R1207_U139 , P1_R1207_U448 , P1_R1207_U175 );
nand NAND2_9915 ( P1_R1207_U140 , P1_R1207_U458 , P1_R1207_U457 );
nand NAND2_9916 ( P1_R1207_U141 , P1_R1207_U463 , P1_R1207_U462 );
and AND2_9917 ( P1_R1207_U142 , P1_R1207_U342 , P1_R1207_U7 );
and AND2_9918 ( P1_R1207_U143 , P1_R1207_U469 , P1_R1207_U174 );
and AND2_9919 ( P1_R1207_U144 , P1_R1207_U349 , P1_R1207_U348 );
nand NAND2_9920 ( P1_R1207_U145 , P1_R1207_U116 , P1_R1207_U207 );
and AND2_9921 ( P1_R1207_U146 , P1_R1207_U358 , P1_R1207_U357 );
and AND2_9922 ( P1_R1207_U147 , P1_R1207_U365 , P1_R1207_U364 );
and AND2_9923 ( P1_R1207_U148 , P1_R1207_U369 , P1_R1207_U368 );
nand NAND2_9924 ( P1_R1207_U149 , P1_R1207_U113 , P1_R1207_U191 );
and AND2_9925 ( P1_R1207_U150 , P1_R1207_U378 , P1_R1207_U377 );
not NOT1_9926 ( P1_R1207_U151 , P1_U3985 );
not NOT1_9927 ( P1_R1207_U152 , P1_U3055 );
and AND2_9928 ( P1_R1207_U153 , P1_R1207_U382 , P1_R1207_U381 );
and AND2_9929 ( P1_R1207_U154 , P1_R1207_U397 , P1_R1207_U396 );
nand NAND2_9930 ( P1_R1207_U155 , P1_R1207_U290 , P1_R1207_U289 );
nand NAND2_9931 ( P1_R1207_U156 , P1_R1207_U286 , P1_R1207_U285 );
and AND2_9932 ( P1_R1207_U157 , P1_R1207_U414 , P1_R1207_U413 );
and AND2_9933 ( P1_R1207_U158 , P1_R1207_U418 , P1_R1207_U417 );
nand NAND2_9934 ( P1_R1207_U159 , P1_R1207_U276 , P1_R1207_U275 );
nand NAND2_9935 ( P1_R1207_U160 , P1_R1207_U272 , P1_R1207_U271 );
not NOT1_9936 ( P1_R1207_U161 , P1_U3455 );
nand NAND2_9937 ( P1_R1207_U162 , P1_R1207_U268 , P1_R1207_U267 );
not NOT1_9938 ( P1_R1207_U163 , P1_U3506 );
nand NAND2_9939 ( P1_R1207_U164 , P1_R1207_U260 , P1_R1207_U259 );
and AND2_9940 ( P1_R1207_U165 , P1_R1207_U450 , P1_R1207_U449 );
and AND2_9941 ( P1_R1207_U166 , P1_R1207_U454 , P1_R1207_U453 );
nand NAND2_9942 ( P1_R1207_U167 , P1_R1207_U250 , P1_R1207_U249 );
nand NAND2_9943 ( P1_R1207_U168 , P1_R1207_U246 , P1_R1207_U245 );
nand NAND2_9944 ( P1_R1207_U169 , P1_R1207_U242 , P1_R1207_U241 );
and AND2_9945 ( P1_R1207_U170 , P1_R1207_U471 , P1_R1207_U470 );
not NOT1_9946 ( P1_R1207_U171 , P1_R1207_U82 );
not NOT1_9947 ( P1_R1207_U172 , P1_R1207_U27 );
not NOT1_9948 ( P1_R1207_U173 , P1_R1207_U37 );
nand NAND2_9949 ( P1_R1207_U174 , P1_U3482 , P1_R1207_U50 );
nand NAND2_9950 ( P1_R1207_U175 , P1_U3497 , P1_R1207_U59 );
nand NAND2_9951 ( P1_R1207_U176 , P1_U3980 , P1_R1207_U73 );
nand NAND2_9952 ( P1_R1207_U177 , P1_U3976 , P1_R1207_U81 );
nand NAND2_9953 ( P1_R1207_U178 , P1_U3458 , P1_R1207_U26 );
nand NAND2_9954 ( P1_R1207_U179 , P1_U3467 , P1_R1207_U32 );
nand NAND2_9955 ( P1_R1207_U180 , P1_U3473 , P1_R1207_U36 );
not NOT1_9956 ( P1_R1207_U181 , P1_R1207_U61 );
not NOT1_9957 ( P1_R1207_U182 , P1_R1207_U75 );
not NOT1_9958 ( P1_R1207_U183 , P1_R1207_U34 );
not NOT1_9959 ( P1_R1207_U184 , P1_R1207_U51 );
not NOT1_9960 ( P1_R1207_U185 , P1_R1207_U23 );
nand NAND2_9961 ( P1_R1207_U186 , P1_R1207_U185 , P1_R1207_U24 );
nand NAND2_9962 ( P1_R1207_U187 , P1_R1207_U186 , P1_R1207_U161 );
nand NAND2_9963 ( P1_R1207_U188 , P1_U3078 , P1_R1207_U23 );
not NOT1_9964 ( P1_R1207_U189 , P1_R1207_U43 );
nand NAND2_9965 ( P1_R1207_U190 , P1_U3461 , P1_R1207_U28 );
nand NAND3_9966 ( P1_R1207_U191 , P1_R1207_U43 , P1_R1207_U178 , P1_R1207_U190 );
nand NAND2_9967 ( P1_R1207_U192 , P1_R1207_U28 , P1_R1207_U27 );
nand NAND2_9968 ( P1_R1207_U193 , P1_R1207_U192 , P1_R1207_U25 );
nand NAND2_9969 ( P1_R1207_U194 , P1_U3064 , P1_R1207_U172 );
not NOT1_9970 ( P1_R1207_U195 , P1_R1207_U149 );
nand NAND2_9971 ( P1_R1207_U196 , P1_U3470 , P1_R1207_U31 );
nand NAND2_9972 ( P1_R1207_U197 , P1_U3071 , P1_R1207_U29 );
nand NAND2_9973 ( P1_R1207_U198 , P1_U3067 , P1_R1207_U20 );
nand NAND2_9974 ( P1_R1207_U199 , P1_R1207_U183 , P1_R1207_U179 );
nand NAND2_9975 ( P1_R1207_U200 , P1_R1207_U6 , P1_R1207_U199 );
nand NAND2_9976 ( P1_R1207_U201 , P1_U3464 , P1_R1207_U33 );
nand NAND2_9977 ( P1_R1207_U202 , P1_U3470 , P1_R1207_U31 );
nand NAND3_9978 ( P1_R1207_U203 , P1_R1207_U149 , P1_R1207_U179 , P1_R1207_U114 );
nand NAND2_9979 ( P1_R1207_U204 , P1_R1207_U202 , P1_R1207_U200 );
not NOT1_9980 ( P1_R1207_U205 , P1_R1207_U41 );
nand NAND2_9981 ( P1_R1207_U206 , P1_U3476 , P1_R1207_U38 );
nand NAND2_9982 ( P1_R1207_U207 , P1_R1207_U115 , P1_R1207_U41 );
nand NAND2_9983 ( P1_R1207_U208 , P1_R1207_U38 , P1_R1207_U37 );
nand NAND2_9984 ( P1_R1207_U209 , P1_R1207_U208 , P1_R1207_U35 );
nand NAND2_9985 ( P1_R1207_U210 , P1_U3084 , P1_R1207_U173 );
not NOT1_9986 ( P1_R1207_U211 , P1_R1207_U145 );
nand NAND2_9987 ( P1_R1207_U212 , P1_U3479 , P1_R1207_U40 );
nand NAND2_9988 ( P1_R1207_U213 , P1_R1207_U212 , P1_R1207_U51 );
nand NAND2_9989 ( P1_R1207_U214 , P1_R1207_U205 , P1_R1207_U37 );
nand NAND2_9990 ( P1_R1207_U215 , P1_R1207_U118 , P1_R1207_U214 );
nand NAND2_9991 ( P1_R1207_U216 , P1_R1207_U41 , P1_R1207_U180 );
nand NAND2_9992 ( P1_R1207_U217 , P1_R1207_U117 , P1_R1207_U216 );
nand NAND2_9993 ( P1_R1207_U218 , P1_R1207_U37 , P1_R1207_U180 );
nand NAND2_9994 ( P1_R1207_U219 , P1_R1207_U201 , P1_R1207_U149 );
not NOT1_9995 ( P1_R1207_U220 , P1_R1207_U42 );
nand NAND2_9996 ( P1_R1207_U221 , P1_U3067 , P1_R1207_U20 );
nand NAND2_9997 ( P1_R1207_U222 , P1_R1207_U220 , P1_R1207_U221 );
nand NAND2_9998 ( P1_R1207_U223 , P1_R1207_U120 , P1_R1207_U222 );
nand NAND2_9999 ( P1_R1207_U224 , P1_R1207_U42 , P1_R1207_U179 );
nand NAND2_10000 ( P1_R1207_U225 , P1_U3470 , P1_R1207_U31 );
nand NAND2_10001 ( P1_R1207_U226 , P1_R1207_U119 , P1_R1207_U224 );
nand NAND2_10002 ( P1_R1207_U227 , P1_U3067 , P1_R1207_U20 );
nand NAND2_10003 ( P1_R1207_U228 , P1_R1207_U179 , P1_R1207_U227 );
nand NAND2_10004 ( P1_R1207_U229 , P1_R1207_U201 , P1_R1207_U34 );
nand NAND2_10005 ( P1_R1207_U230 , P1_R1207_U189 , P1_R1207_U27 );
nand NAND2_10006 ( P1_R1207_U231 , P1_R1207_U122 , P1_R1207_U230 );
nand NAND2_10007 ( P1_R1207_U232 , P1_R1207_U43 , P1_R1207_U178 );
nand NAND2_10008 ( P1_R1207_U233 , P1_R1207_U121 , P1_R1207_U232 );
nand NAND2_10009 ( P1_R1207_U234 , P1_R1207_U27 , P1_R1207_U178 );
nand NAND2_10010 ( P1_R1207_U235 , P1_U3485 , P1_R1207_U49 );
nand NAND2_10011 ( P1_R1207_U236 , P1_U3063 , P1_R1207_U48 );
nand NAND2_10012 ( P1_R1207_U237 , P1_U3062 , P1_R1207_U47 );
nand NAND2_10013 ( P1_R1207_U238 , P1_R1207_U184 , P1_R1207_U174 );
nand NAND2_10014 ( P1_R1207_U239 , P1_R1207_U7 , P1_R1207_U238 );
nand NAND2_10015 ( P1_R1207_U240 , P1_U3485 , P1_R1207_U49 );
nand NAND2_10016 ( P1_R1207_U241 , P1_R1207_U145 , P1_R1207_U123 );
nand NAND2_10017 ( P1_R1207_U242 , P1_R1207_U240 , P1_R1207_U239 );
not NOT1_10018 ( P1_R1207_U243 , P1_R1207_U169 );
nand NAND2_10019 ( P1_R1207_U244 , P1_U3488 , P1_R1207_U53 );
nand NAND2_10020 ( P1_R1207_U245 , P1_R1207_U244 , P1_R1207_U169 );
nand NAND2_10021 ( P1_R1207_U246 , P1_U3072 , P1_R1207_U52 );
not NOT1_10022 ( P1_R1207_U247 , P1_R1207_U168 );
nand NAND2_10023 ( P1_R1207_U248 , P1_U3491 , P1_R1207_U55 );
nand NAND2_10024 ( P1_R1207_U249 , P1_R1207_U248 , P1_R1207_U168 );
nand NAND2_10025 ( P1_R1207_U250 , P1_U3080 , P1_R1207_U54 );
not NOT1_10026 ( P1_R1207_U251 , P1_R1207_U167 );
nand NAND2_10027 ( P1_R1207_U252 , P1_U3500 , P1_R1207_U58 );
nand NAND2_10028 ( P1_R1207_U253 , P1_U3073 , P1_R1207_U56 );
nand NAND2_10029 ( P1_R1207_U254 , P1_U3074 , P1_R1207_U46 );
nand NAND2_10030 ( P1_R1207_U255 , P1_R1207_U181 , P1_R1207_U175 );
nand NAND2_10031 ( P1_R1207_U256 , P1_R1207_U8 , P1_R1207_U255 );
nand NAND2_10032 ( P1_R1207_U257 , P1_U3494 , P1_R1207_U60 );
nand NAND2_10033 ( P1_R1207_U258 , P1_U3500 , P1_R1207_U58 );
nand NAND2_10034 ( P1_R1207_U259 , P1_R1207_U167 , P1_R1207_U124 );
nand NAND2_10035 ( P1_R1207_U260 , P1_R1207_U258 , P1_R1207_U256 );
not NOT1_10036 ( P1_R1207_U261 , P1_R1207_U164 );
nand NAND2_10037 ( P1_R1207_U262 , P1_U3503 , P1_R1207_U63 );
nand NAND2_10038 ( P1_R1207_U263 , P1_R1207_U262 , P1_R1207_U164 );
nand NAND2_10039 ( P1_R1207_U264 , P1_U3069 , P1_R1207_U62 );
not NOT1_10040 ( P1_R1207_U265 , P1_R1207_U64 );
nand NAND2_10041 ( P1_R1207_U266 , P1_R1207_U265 , P1_R1207_U65 );
nand NAND2_10042 ( P1_R1207_U267 , P1_R1207_U266 , P1_R1207_U163 );
nand NAND2_10043 ( P1_R1207_U268 , P1_U3082 , P1_R1207_U64 );
not NOT1_10044 ( P1_R1207_U269 , P1_R1207_U162 );
nand NAND2_10045 ( P1_R1207_U270 , P1_U3508 , P1_R1207_U67 );
nand NAND2_10046 ( P1_R1207_U271 , P1_R1207_U270 , P1_R1207_U162 );
nand NAND2_10047 ( P1_R1207_U272 , P1_U3081 , P1_R1207_U66 );
not NOT1_10048 ( P1_R1207_U273 , P1_R1207_U160 );
nand NAND2_10049 ( P1_R1207_U274 , P1_U3982 , P1_R1207_U69 );
nand NAND2_10050 ( P1_R1207_U275 , P1_R1207_U274 , P1_R1207_U160 );
nand NAND2_10051 ( P1_R1207_U276 , P1_U3076 , P1_R1207_U68 );
not NOT1_10052 ( P1_R1207_U277 , P1_R1207_U159 );
nand NAND2_10053 ( P1_R1207_U278 , P1_U3979 , P1_R1207_U72 );
nand NAND2_10054 ( P1_R1207_U279 , P1_U3066 , P1_R1207_U70 );
nand NAND2_10055 ( P1_R1207_U280 , P1_U3061 , P1_R1207_U45 );
nand NAND2_10056 ( P1_R1207_U281 , P1_R1207_U182 , P1_R1207_U176 );
nand NAND2_10057 ( P1_R1207_U282 , P1_R1207_U9 , P1_R1207_U281 );
nand NAND2_10058 ( P1_R1207_U283 , P1_U3981 , P1_R1207_U74 );
nand NAND2_10059 ( P1_R1207_U284 , P1_U3979 , P1_R1207_U72 );
nand NAND3_10060 ( P1_R1207_U285 , P1_R1207_U159 , P1_R1207_U125 , P1_R1207_U278 );
nand NAND2_10061 ( P1_R1207_U286 , P1_R1207_U284 , P1_R1207_U282 );
not NOT1_10062 ( P1_R1207_U287 , P1_R1207_U156 );
nand NAND2_10063 ( P1_R1207_U288 , P1_U3978 , P1_R1207_U77 );
nand NAND2_10064 ( P1_R1207_U289 , P1_R1207_U288 , P1_R1207_U156 );
nand NAND2_10065 ( P1_R1207_U290 , P1_U3065 , P1_R1207_U76 );
not NOT1_10066 ( P1_R1207_U291 , P1_R1207_U155 );
nand NAND2_10067 ( P1_R1207_U292 , P1_U3977 , P1_R1207_U79 );
nand NAND2_10068 ( P1_R1207_U293 , P1_R1207_U292 , P1_R1207_U155 );
nand NAND2_10069 ( P1_R1207_U294 , P1_U3058 , P1_R1207_U78 );
not NOT1_10070 ( P1_R1207_U295 , P1_R1207_U87 );
nand NAND2_10071 ( P1_R1207_U296 , P1_U3975 , P1_R1207_U83 );
nand NAND3_10072 ( P1_R1207_U297 , P1_R1207_U87 , P1_R1207_U177 , P1_R1207_U296 );
nand NAND2_10073 ( P1_R1207_U298 , P1_R1207_U83 , P1_R1207_U82 );
nand NAND2_10074 ( P1_R1207_U299 , P1_R1207_U298 , P1_R1207_U80 );
nand NAND2_10075 ( P1_R1207_U300 , P1_U3053 , P1_R1207_U171 );
not NOT1_10076 ( P1_R1207_U301 , P1_R1207_U86 );
nand NAND2_10077 ( P1_R1207_U302 , P1_U3054 , P1_R1207_U84 );
nand NAND2_10078 ( P1_R1207_U303 , P1_R1207_U301 , P1_R1207_U302 );
nand NAND2_10079 ( P1_R1207_U304 , P1_U3974 , P1_R1207_U85 );
nand NAND2_10080 ( P1_R1207_U305 , P1_U3974 , P1_R1207_U85 );
nand NAND2_10081 ( P1_R1207_U306 , P1_R1207_U305 , P1_R1207_U86 );
nand NAND2_10082 ( P1_R1207_U307 , P1_U3054 , P1_R1207_U84 );
nand NAND3_10083 ( P1_R1207_U308 , P1_R1207_U307 , P1_R1207_U306 , P1_R1207_U153 );
nand NAND2_10084 ( P1_R1207_U309 , P1_R1207_U295 , P1_R1207_U82 );
nand NAND2_10085 ( P1_R1207_U310 , P1_R1207_U129 , P1_R1207_U309 );
nand NAND2_10086 ( P1_R1207_U311 , P1_R1207_U87 , P1_R1207_U177 );
nand NAND2_10087 ( P1_R1207_U312 , P1_R1207_U128 , P1_R1207_U311 );
nand NAND2_10088 ( P1_R1207_U313 , P1_R1207_U82 , P1_R1207_U177 );
nand NAND2_10089 ( P1_R1207_U314 , P1_R1207_U283 , P1_R1207_U159 );
not NOT1_10090 ( P1_R1207_U315 , P1_R1207_U88 );
nand NAND2_10091 ( P1_R1207_U316 , P1_U3061 , P1_R1207_U45 );
nand NAND2_10092 ( P1_R1207_U317 , P1_R1207_U315 , P1_R1207_U316 );
nand NAND2_10093 ( P1_R1207_U318 , P1_R1207_U132 , P1_R1207_U317 );
nand NAND2_10094 ( P1_R1207_U319 , P1_R1207_U88 , P1_R1207_U176 );
nand NAND2_10095 ( P1_R1207_U320 , P1_U3979 , P1_R1207_U72 );
nand NAND3_10096 ( P1_R1207_U321 , P1_R1207_U320 , P1_R1207_U319 , P1_R1207_U9 );
nand NAND2_10097 ( P1_R1207_U322 , P1_U3061 , P1_R1207_U45 );
nand NAND2_10098 ( P1_R1207_U323 , P1_R1207_U176 , P1_R1207_U322 );
nand NAND2_10099 ( P1_R1207_U324 , P1_R1207_U283 , P1_R1207_U75 );
nand NAND2_10100 ( P1_R1207_U325 , P1_R1207_U257 , P1_R1207_U167 );
not NOT1_10101 ( P1_R1207_U326 , P1_R1207_U89 );
nand NAND2_10102 ( P1_R1207_U327 , P1_U3074 , P1_R1207_U46 );
nand NAND2_10103 ( P1_R1207_U328 , P1_R1207_U326 , P1_R1207_U327 );
nand NAND2_10104 ( P1_R1207_U329 , P1_R1207_U139 , P1_R1207_U328 );
nand NAND2_10105 ( P1_R1207_U330 , P1_R1207_U89 , P1_R1207_U175 );
nand NAND2_10106 ( P1_R1207_U331 , P1_U3500 , P1_R1207_U58 );
nand NAND2_10107 ( P1_R1207_U332 , P1_R1207_U138 , P1_R1207_U330 );
nand NAND2_10108 ( P1_R1207_U333 , P1_U3074 , P1_R1207_U46 );
nand NAND2_10109 ( P1_R1207_U334 , P1_R1207_U175 , P1_R1207_U333 );
nand NAND2_10110 ( P1_R1207_U335 , P1_R1207_U257 , P1_R1207_U61 );
nand NAND2_10111 ( P1_R1207_U336 , P1_R1207_U212 , P1_R1207_U145 );
not NOT1_10112 ( P1_R1207_U337 , P1_R1207_U90 );
nand NAND2_10113 ( P1_R1207_U338 , P1_U3062 , P1_R1207_U47 );
nand NAND2_10114 ( P1_R1207_U339 , P1_R1207_U337 , P1_R1207_U338 );
nand NAND2_10115 ( P1_R1207_U340 , P1_R1207_U143 , P1_R1207_U339 );
nand NAND2_10116 ( P1_R1207_U341 , P1_R1207_U90 , P1_R1207_U174 );
nand NAND2_10117 ( P1_R1207_U342 , P1_U3485 , P1_R1207_U49 );
nand NAND2_10118 ( P1_R1207_U343 , P1_R1207_U142 , P1_R1207_U341 );
nand NAND2_10119 ( P1_R1207_U344 , P1_U3062 , P1_R1207_U47 );
nand NAND2_10120 ( P1_R1207_U345 , P1_R1207_U174 , P1_R1207_U344 );
nand NAND2_10121 ( P1_R1207_U346 , P1_U3077 , P1_R1207_U22 );
nand NAND3_10122 ( P1_R1207_U347 , P1_R1207_U304 , P1_R1207_U303 , P1_R1207_U385 );
nand NAND2_10123 ( P1_R1207_U348 , P1_U3479 , P1_R1207_U40 );
nand NAND2_10124 ( P1_R1207_U349 , P1_U3083 , P1_R1207_U39 );
nand NAND2_10125 ( P1_R1207_U350 , P1_R1207_U213 , P1_R1207_U145 );
nand NAND2_10126 ( P1_R1207_U351 , P1_R1207_U211 , P1_R1207_U144 );
nand NAND2_10127 ( P1_R1207_U352 , P1_U3476 , P1_R1207_U38 );
nand NAND2_10128 ( P1_R1207_U353 , P1_U3084 , P1_R1207_U35 );
nand NAND2_10129 ( P1_R1207_U354 , P1_U3476 , P1_R1207_U38 );
nand NAND2_10130 ( P1_R1207_U355 , P1_U3084 , P1_R1207_U35 );
nand NAND2_10131 ( P1_R1207_U356 , P1_R1207_U355 , P1_R1207_U354 );
nand NAND2_10132 ( P1_R1207_U357 , P1_U3473 , P1_R1207_U36 );
nand NAND2_10133 ( P1_R1207_U358 , P1_U3070 , P1_R1207_U19 );
nand NAND2_10134 ( P1_R1207_U359 , P1_R1207_U218 , P1_R1207_U41 );
nand NAND2_10135 ( P1_R1207_U360 , P1_R1207_U146 , P1_R1207_U205 );
nand NAND2_10136 ( P1_R1207_U361 , P1_U3470 , P1_R1207_U31 );
nand NAND2_10137 ( P1_R1207_U362 , P1_U3071 , P1_R1207_U29 );
nand NAND2_10138 ( P1_R1207_U363 , P1_R1207_U362 , P1_R1207_U361 );
nand NAND2_10139 ( P1_R1207_U364 , P1_U3467 , P1_R1207_U32 );
nand NAND2_10140 ( P1_R1207_U365 , P1_U3067 , P1_R1207_U20 );
nand NAND2_10141 ( P1_R1207_U366 , P1_R1207_U228 , P1_R1207_U42 );
nand NAND2_10142 ( P1_R1207_U367 , P1_R1207_U147 , P1_R1207_U220 );
nand NAND2_10143 ( P1_R1207_U368 , P1_U3464 , P1_R1207_U33 );
nand NAND2_10144 ( P1_R1207_U369 , P1_U3060 , P1_R1207_U30 );
nand NAND2_10145 ( P1_R1207_U370 , P1_R1207_U229 , P1_R1207_U149 );
nand NAND2_10146 ( P1_R1207_U371 , P1_R1207_U195 , P1_R1207_U148 );
nand NAND2_10147 ( P1_R1207_U372 , P1_U3461 , P1_R1207_U28 );
nand NAND2_10148 ( P1_R1207_U373 , P1_U3064 , P1_R1207_U25 );
nand NAND2_10149 ( P1_R1207_U374 , P1_U3461 , P1_R1207_U28 );
nand NAND2_10150 ( P1_R1207_U375 , P1_U3064 , P1_R1207_U25 );
nand NAND2_10151 ( P1_R1207_U376 , P1_R1207_U375 , P1_R1207_U374 );
nand NAND2_10152 ( P1_R1207_U377 , P1_U3458 , P1_R1207_U26 );
nand NAND2_10153 ( P1_R1207_U378 , P1_U3068 , P1_R1207_U21 );
nand NAND2_10154 ( P1_R1207_U379 , P1_R1207_U234 , P1_R1207_U43 );
nand NAND2_10155 ( P1_R1207_U380 , P1_R1207_U150 , P1_R1207_U189 );
nand NAND2_10156 ( P1_R1207_U381 , P1_U3985 , P1_R1207_U152 );
nand NAND2_10157 ( P1_R1207_U382 , P1_U3055 , P1_R1207_U151 );
nand NAND2_10158 ( P1_R1207_U383 , P1_U3985 , P1_R1207_U152 );
nand NAND2_10159 ( P1_R1207_U384 , P1_U3055 , P1_R1207_U151 );
nand NAND2_10160 ( P1_R1207_U385 , P1_R1207_U384 , P1_R1207_U383 );
nand NAND2_10161 ( P1_R1207_U386 , P1_U3974 , P1_R1207_U85 );
nand NAND2_10162 ( P1_R1207_U387 , P1_U3054 , P1_R1207_U84 );
not NOT1_10163 ( P1_R1207_U388 , P1_R1207_U127 );
nand NAND2_10164 ( P1_R1207_U389 , P1_R1207_U388 , P1_R1207_U301 );
nand NAND2_10165 ( P1_R1207_U390 , P1_R1207_U127 , P1_R1207_U86 );
nand NAND2_10166 ( P1_R1207_U391 , P1_U3975 , P1_R1207_U83 );
nand NAND2_10167 ( P1_R1207_U392 , P1_U3053 , P1_R1207_U80 );
nand NAND2_10168 ( P1_R1207_U393 , P1_U3975 , P1_R1207_U83 );
nand NAND2_10169 ( P1_R1207_U394 , P1_U3053 , P1_R1207_U80 );
nand NAND2_10170 ( P1_R1207_U395 , P1_R1207_U394 , P1_R1207_U393 );
nand NAND2_10171 ( P1_R1207_U396 , P1_U3976 , P1_R1207_U81 );
nand NAND2_10172 ( P1_R1207_U397 , P1_U3057 , P1_R1207_U44 );
nand NAND2_10173 ( P1_R1207_U398 , P1_R1207_U313 , P1_R1207_U87 );
nand NAND2_10174 ( P1_R1207_U399 , P1_R1207_U154 , P1_R1207_U295 );
nand NAND2_10175 ( P1_R1207_U400 , P1_U3977 , P1_R1207_U79 );
nand NAND2_10176 ( P1_R1207_U401 , P1_U3058 , P1_R1207_U78 );
not NOT1_10177 ( P1_R1207_U402 , P1_R1207_U130 );
nand NAND2_10178 ( P1_R1207_U403 , P1_R1207_U291 , P1_R1207_U402 );
nand NAND2_10179 ( P1_R1207_U404 , P1_R1207_U130 , P1_R1207_U155 );
nand NAND2_10180 ( P1_R1207_U405 , P1_U3978 , P1_R1207_U77 );
nand NAND2_10181 ( P1_R1207_U406 , P1_U3065 , P1_R1207_U76 );
not NOT1_10182 ( P1_R1207_U407 , P1_R1207_U131 );
nand NAND2_10183 ( P1_R1207_U408 , P1_R1207_U287 , P1_R1207_U407 );
nand NAND2_10184 ( P1_R1207_U409 , P1_R1207_U131 , P1_R1207_U156 );
nand NAND2_10185 ( P1_R1207_U410 , P1_U3979 , P1_R1207_U72 );
nand NAND2_10186 ( P1_R1207_U411 , P1_U3066 , P1_R1207_U70 );
nand NAND2_10187 ( P1_R1207_U412 , P1_R1207_U411 , P1_R1207_U410 );
nand NAND2_10188 ( P1_R1207_U413 , P1_U3980 , P1_R1207_U73 );
nand NAND2_10189 ( P1_R1207_U414 , P1_U3061 , P1_R1207_U45 );
nand NAND2_10190 ( P1_R1207_U415 , P1_R1207_U323 , P1_R1207_U88 );
nand NAND2_10191 ( P1_R1207_U416 , P1_R1207_U157 , P1_R1207_U315 );
nand NAND2_10192 ( P1_R1207_U417 , P1_U3981 , P1_R1207_U74 );
nand NAND2_10193 ( P1_R1207_U418 , P1_U3075 , P1_R1207_U71 );
nand NAND2_10194 ( P1_R1207_U419 , P1_R1207_U324 , P1_R1207_U159 );
nand NAND2_10195 ( P1_R1207_U420 , P1_R1207_U277 , P1_R1207_U158 );
nand NAND2_10196 ( P1_R1207_U421 , P1_U3982 , P1_R1207_U69 );
nand NAND2_10197 ( P1_R1207_U422 , P1_U3076 , P1_R1207_U68 );
not NOT1_10198 ( P1_R1207_U423 , P1_R1207_U133 );
nand NAND2_10199 ( P1_R1207_U424 , P1_R1207_U273 , P1_R1207_U423 );
nand NAND2_10200 ( P1_R1207_U425 , P1_R1207_U133 , P1_R1207_U160 );
nand NAND2_10201 ( P1_R1207_U426 , P1_R1207_U185 , P1_R1207_U24 );
nand NAND2_10202 ( P1_R1207_U427 , P1_U3078 , P1_R1207_U23 );
not NOT1_10203 ( P1_R1207_U428 , P1_R1207_U134 );
nand NAND2_10204 ( P1_R1207_U429 , P1_U3455 , P1_R1207_U428 );
nand NAND2_10205 ( P1_R1207_U430 , P1_R1207_U134 , P1_R1207_U161 );
nand NAND2_10206 ( P1_R1207_U431 , P1_U3508 , P1_R1207_U67 );
nand NAND2_10207 ( P1_R1207_U432 , P1_U3081 , P1_R1207_U66 );
not NOT1_10208 ( P1_R1207_U433 , P1_R1207_U135 );
nand NAND2_10209 ( P1_R1207_U434 , P1_R1207_U269 , P1_R1207_U433 );
nand NAND2_10210 ( P1_R1207_U435 , P1_R1207_U135 , P1_R1207_U162 );
nand NAND2_10211 ( P1_R1207_U436 , P1_U3506 , P1_R1207_U65 );
nand NAND2_10212 ( P1_R1207_U437 , P1_U3082 , P1_R1207_U163 );
not NOT1_10213 ( P1_R1207_U438 , P1_R1207_U136 );
nand NAND2_10214 ( P1_R1207_U439 , P1_R1207_U438 , P1_R1207_U265 );
nand NAND2_10215 ( P1_R1207_U440 , P1_R1207_U136 , P1_R1207_U64 );
nand NAND2_10216 ( P1_R1207_U441 , P1_U3503 , P1_R1207_U63 );
nand NAND2_10217 ( P1_R1207_U442 , P1_U3069 , P1_R1207_U62 );
not NOT1_10218 ( P1_R1207_U443 , P1_R1207_U137 );
nand NAND2_10219 ( P1_R1207_U444 , P1_R1207_U261 , P1_R1207_U443 );
nand NAND2_10220 ( P1_R1207_U445 , P1_R1207_U137 , P1_R1207_U164 );
nand NAND2_10221 ( P1_R1207_U446 , P1_U3500 , P1_R1207_U58 );
nand NAND2_10222 ( P1_R1207_U447 , P1_U3073 , P1_R1207_U56 );
nand NAND2_10223 ( P1_R1207_U448 , P1_R1207_U447 , P1_R1207_U446 );
nand NAND2_10224 ( P1_R1207_U449 , P1_U3497 , P1_R1207_U59 );
nand NAND2_10225 ( P1_R1207_U450 , P1_U3074 , P1_R1207_U46 );
nand NAND2_10226 ( P1_R1207_U451 , P1_R1207_U334 , P1_R1207_U89 );
nand NAND2_10227 ( P1_R1207_U452 , P1_R1207_U165 , P1_R1207_U326 );
nand NAND2_10228 ( P1_R1207_U453 , P1_U3494 , P1_R1207_U60 );
nand NAND2_10229 ( P1_R1207_U454 , P1_U3079 , P1_R1207_U57 );
nand NAND2_10230 ( P1_R1207_U455 , P1_R1207_U335 , P1_R1207_U167 );
nand NAND2_10231 ( P1_R1207_U456 , P1_R1207_U251 , P1_R1207_U166 );
nand NAND2_10232 ( P1_R1207_U457 , P1_U3491 , P1_R1207_U55 );
nand NAND2_10233 ( P1_R1207_U458 , P1_U3080 , P1_R1207_U54 );
not NOT1_10234 ( P1_R1207_U459 , P1_R1207_U140 );
nand NAND2_10235 ( P1_R1207_U460 , P1_R1207_U247 , P1_R1207_U459 );
nand NAND2_10236 ( P1_R1207_U461 , P1_R1207_U140 , P1_R1207_U168 );
nand NAND2_10237 ( P1_R1207_U462 , P1_U3488 , P1_R1207_U53 );
nand NAND2_10238 ( P1_R1207_U463 , P1_U3072 , P1_R1207_U52 );
not NOT1_10239 ( P1_R1207_U464 , P1_R1207_U141 );
nand NAND2_10240 ( P1_R1207_U465 , P1_R1207_U243 , P1_R1207_U464 );
nand NAND2_10241 ( P1_R1207_U466 , P1_R1207_U141 , P1_R1207_U169 );
nand NAND2_10242 ( P1_R1207_U467 , P1_U3485 , P1_R1207_U49 );
nand NAND2_10243 ( P1_R1207_U468 , P1_U3063 , P1_R1207_U48 );
nand NAND2_10244 ( P1_R1207_U469 , P1_R1207_U468 , P1_R1207_U467 );
nand NAND2_10245 ( P1_R1207_U470 , P1_U3482 , P1_R1207_U50 );
nand NAND2_10246 ( P1_R1207_U471 , P1_U3062 , P1_R1207_U47 );
nand NAND2_10247 ( P1_R1207_U472 , P1_R1207_U345 , P1_R1207_U90 );
nand NAND2_10248 ( P1_R1207_U473 , P1_R1207_U170 , P1_R1207_U337 );
and AND2_10249 ( P1_R1165_U4 , P1_R1165_U210 , P1_R1165_U209 );
and AND2_10250 ( P1_R1165_U5 , P1_R1165_U222 , P1_R1165_U221 );
and AND2_10251 ( P1_R1165_U6 , P1_R1165_U253 , P1_R1165_U252 );
and AND2_10252 ( P1_R1165_U7 , P1_R1165_U271 , P1_R1165_U270 );
and AND2_10253 ( P1_R1165_U8 , P1_R1165_U283 , P1_R1165_U282 );
and AND2_10254 ( P1_R1165_U9 , P1_R1165_U507 , P1_R1165_U506 );
and AND2_10255 ( P1_R1165_U10 , P1_R1165_U339 , P1_R1165_U336 );
and AND2_10256 ( P1_R1165_U11 , P1_R1165_U330 , P1_R1165_U327 );
and AND2_10257 ( P1_R1165_U12 , P1_R1165_U323 , P1_R1165_U320 );
and AND3_10258 ( P1_R1165_U13 , P1_R1165_U360 , P1_R1165_U311 , P1_R1165_U314 );
and AND2_10259 ( P1_R1165_U14 , P1_R1165_U245 , P1_R1165_U242 );
and AND2_10260 ( P1_R1165_U15 , P1_R1165_U238 , P1_R1165_U235 );
not NOT1_10261 ( P1_R1165_U16 , P1_U3211 );
not NOT1_10262 ( P1_R1165_U17 , P1_U3175 );
nand NAND2_10263 ( P1_R1165_U18 , P1_U3175 , P1_R1165_U58 );
not NOT1_10264 ( P1_R1165_U19 , P1_U3174 );
not NOT1_10265 ( P1_R1165_U20 , P1_U3177 );
not NOT1_10266 ( P1_R1165_U21 , P1_U3179 );
nand NAND2_10267 ( P1_R1165_U22 , P1_U3179 , P1_R1165_U61 );
not NOT1_10268 ( P1_R1165_U23 , P1_U3178 );
not NOT1_10269 ( P1_R1165_U24 , P1_U3181 );
not NOT1_10270 ( P1_R1165_U25 , P1_U3180 );
not NOT1_10271 ( P1_R1165_U26 , P1_U3176 );
not NOT1_10272 ( P1_R1165_U27 , P1_U3173 );
not NOT1_10273 ( P1_R1165_U28 , P1_U3172 );
nand NAND2_10274 ( P1_R1165_U29 , P1_R1165_U219 , P1_R1165_U218 );
nand NAND2_10275 ( P1_R1165_U30 , P1_R1165_U207 , P1_R1165_U206 );
not NOT1_10276 ( P1_R1165_U31 , P1_U3154 );
not NOT1_10277 ( P1_R1165_U32 , P1_U3155 );
not NOT1_10278 ( P1_R1165_U33 , P1_U3156 );
not NOT1_10279 ( P1_R1165_U34 , P1_U3157 );
not NOT1_10280 ( P1_R1165_U35 , P1_U3165 );
nand NAND2_10281 ( P1_R1165_U36 , P1_U3165 , P1_R1165_U71 );
not NOT1_10282 ( P1_R1165_U37 , P1_U3164 );
not NOT1_10283 ( P1_R1165_U38 , P1_U3171 );
not NOT1_10284 ( P1_R1165_U39 , P1_U3169 );
not NOT1_10285 ( P1_R1165_U40 , P1_U3170 );
nand NAND2_10286 ( P1_R1165_U41 , P1_U3170 , P1_R1165_U74 );
not NOT1_10287 ( P1_R1165_U42 , P1_U3168 );
not NOT1_10288 ( P1_R1165_U43 , P1_U3167 );
not NOT1_10289 ( P1_R1165_U44 , P1_U3166 );
not NOT1_10290 ( P1_R1165_U45 , P1_U3163 );
not NOT1_10291 ( P1_R1165_U46 , P1_U3161 );
not NOT1_10292 ( P1_R1165_U47 , P1_U3162 );
nand NAND2_10293 ( P1_R1165_U48 , P1_U3162 , P1_R1165_U80 );
not NOT1_10294 ( P1_R1165_U49 , P1_U3160 );
not NOT1_10295 ( P1_R1165_U50 , P1_U3159 );
not NOT1_10296 ( P1_R1165_U51 , P1_U3158 );
nand NAND2_10297 ( P1_R1165_U52 , P1_U3155 , P1_R1165_U69 );
nand NAND2_10298 ( P1_R1165_U53 , P1_R1165_U200 , P1_R1165_U309 );
nand NAND2_10299 ( P1_R1165_U54 , P1_R1165_U48 , P1_R1165_U316 );
nand NAND2_10300 ( P1_R1165_U55 , P1_R1165_U268 , P1_R1165_U267 );
nand NAND2_10301 ( P1_R1165_U56 , P1_R1165_U41 , P1_R1165_U332 );
nand NAND2_10302 ( P1_R1165_U57 , P1_R1165_U366 , P1_R1165_U365 );
nand NAND2_10303 ( P1_R1165_U58 , P1_R1165_U395 , P1_R1165_U394 );
nand NAND2_10304 ( P1_R1165_U59 , P1_R1165_U392 , P1_R1165_U391 );
nand NAND2_10305 ( P1_R1165_U60 , P1_R1165_U374 , P1_R1165_U373 );
nand NAND2_10306 ( P1_R1165_U61 , P1_R1165_U386 , P1_R1165_U385 );
nand NAND2_10307 ( P1_R1165_U62 , P1_R1165_U383 , P1_R1165_U382 );
nand NAND2_10308 ( P1_R1165_U63 , P1_R1165_U377 , P1_R1165_U376 );
nand NAND2_10309 ( P1_R1165_U64 , P1_R1165_U380 , P1_R1165_U379 );
nand NAND2_10310 ( P1_R1165_U65 , P1_R1165_U389 , P1_R1165_U388 );
nand NAND2_10311 ( P1_R1165_U66 , P1_R1165_U398 , P1_R1165_U397 );
nand NAND2_10312 ( P1_R1165_U67 , P1_R1165_U438 , P1_R1165_U437 );
nand NAND2_10313 ( P1_R1165_U68 , P1_R1165_U441 , P1_R1165_U440 );
nand NAND2_10314 ( P1_R1165_U69 , P1_R1165_U444 , P1_R1165_U443 );
nand NAND2_10315 ( P1_R1165_U70 , P1_R1165_U447 , P1_R1165_U446 );
nand NAND2_10316 ( P1_R1165_U71 , P1_R1165_U471 , P1_R1165_U470 );
nand NAND2_10317 ( P1_R1165_U72 , P1_R1165_U468 , P1_R1165_U467 );
nand NAND2_10318 ( P1_R1165_U73 , P1_R1165_U450 , P1_R1165_U449 );
nand NAND2_10319 ( P1_R1165_U74 , P1_R1165_U459 , P1_R1165_U458 );
nand NAND2_10320 ( P1_R1165_U75 , P1_R1165_U453 , P1_R1165_U452 );
nand NAND2_10321 ( P1_R1165_U76 , P1_R1165_U456 , P1_R1165_U455 );
nand NAND2_10322 ( P1_R1165_U77 , P1_R1165_U462 , P1_R1165_U461 );
nand NAND2_10323 ( P1_R1165_U78 , P1_R1165_U465 , P1_R1165_U464 );
nand NAND2_10324 ( P1_R1165_U79 , P1_R1165_U474 , P1_R1165_U473 );
nand NAND2_10325 ( P1_R1165_U80 , P1_R1165_U483 , P1_R1165_U482 );
nand NAND2_10326 ( P1_R1165_U81 , P1_R1165_U477 , P1_R1165_U476 );
nand NAND2_10327 ( P1_R1165_U82 , P1_R1165_U480 , P1_R1165_U479 );
nand NAND2_10328 ( P1_R1165_U83 , P1_R1165_U486 , P1_R1165_U485 );
nand NAND2_10329 ( P1_R1165_U84 , P1_R1165_U489 , P1_R1165_U488 );
nand NAND2_10330 ( P1_R1165_U85 , P1_R1165_U495 , P1_R1165_U494 );
nand NAND2_10331 ( P1_R1165_U86 , P1_R1165_U602 , P1_R1165_U601 );
nand NAND2_10332 ( P1_R1165_U87 , P1_R1165_U401 , P1_R1165_U400 );
nand NAND2_10333 ( P1_R1165_U88 , P1_R1165_U408 , P1_R1165_U407 );
nand NAND2_10334 ( P1_R1165_U89 , P1_R1165_U415 , P1_R1165_U414 );
nand NAND2_10335 ( P1_R1165_U90 , P1_R1165_U422 , P1_R1165_U421 );
nand NAND2_10336 ( P1_R1165_U91 , P1_R1165_U429 , P1_R1165_U428 );
nand NAND2_10337 ( P1_R1165_U92 , P1_R1165_U436 , P1_R1165_U435 );
nand NAND2_10338 ( P1_R1165_U93 , P1_R1165_U498 , P1_R1165_U497 );
nand NAND2_10339 ( P1_R1165_U94 , P1_R1165_U505 , P1_R1165_U504 );
nand NAND2_10340 ( P1_R1165_U95 , P1_R1165_U512 , P1_R1165_U511 );
nand NAND2_10341 ( P1_R1165_U96 , P1_R1165_U517 , P1_R1165_U516 );
nand NAND2_10342 ( P1_R1165_U97 , P1_R1165_U524 , P1_R1165_U523 );
nand NAND2_10343 ( P1_R1165_U98 , P1_R1165_U531 , P1_R1165_U530 );
nand NAND2_10344 ( P1_R1165_U99 , P1_R1165_U538 , P1_R1165_U537 );
nand NAND2_10345 ( P1_R1165_U100 , P1_R1165_U545 , P1_R1165_U544 );
nand NAND2_10346 ( P1_R1165_U101 , P1_R1165_U550 , P1_R1165_U549 );
nand NAND2_10347 ( P1_R1165_U102 , P1_R1165_U557 , P1_R1165_U556 );
nand NAND2_10348 ( P1_R1165_U103 , P1_R1165_U564 , P1_R1165_U563 );
nand NAND2_10349 ( P1_R1165_U104 , P1_R1165_U571 , P1_R1165_U570 );
nand NAND2_10350 ( P1_R1165_U105 , P1_R1165_U578 , P1_R1165_U577 );
nand NAND2_10351 ( P1_R1165_U106 , P1_R1165_U585 , P1_R1165_U584 );
nand NAND2_10352 ( P1_R1165_U107 , P1_R1165_U590 , P1_R1165_U589 );
nand NAND2_10353 ( P1_R1165_U108 , P1_R1165_U597 , P1_R1165_U596 );
and AND2_10354 ( P1_R1165_U109 , P1_R1165_U213 , P1_R1165_U212 );
and AND2_10355 ( P1_R1165_U110 , P1_R1165_U226 , P1_R1165_U225 );
and AND3_10356 ( P1_R1165_U111 , P1_R1165_U410 , P1_R1165_U409 , P1_R1165_U18 );
and AND2_10357 ( P1_R1165_U112 , P1_R1165_U237 , P1_R1165_U5 );
and AND3_10358 ( P1_R1165_U113 , P1_R1165_U431 , P1_R1165_U430 , P1_R1165_U22 );
and AND2_10359 ( P1_R1165_U114 , P1_R1165_U244 , P1_R1165_U4 );
and AND2_10360 ( P1_R1165_U115 , P1_R1165_U257 , P1_R1165_U6 );
and AND2_10361 ( P1_R1165_U116 , P1_R1165_U255 , P1_R1165_U195 );
and AND2_10362 ( P1_R1165_U117 , P1_R1165_U275 , P1_R1165_U274 );
and AND2_10363 ( P1_R1165_U118 , P1_R1165_U287 , P1_R1165_U8 );
and AND2_10364 ( P1_R1165_U119 , P1_R1165_U285 , P1_R1165_U196 );
and AND2_10365 ( P1_R1165_U120 , P1_R1165_U359 , P1_R1165_U52 );
and AND2_10366 ( P1_R1165_U121 , P1_R1165_U308 , P1_R1165_U303 );
and AND2_10367 ( P1_R1165_U122 , P1_R1165_U356 , P1_R1165_U307 );
nand NAND2_10368 ( P1_R1165_U123 , P1_R1165_U492 , P1_R1165_U491 );
and AND2_10369 ( P1_R1165_U124 , P1_R1165_U352 , P1_R1165_U52 );
and AND2_10370 ( P1_R1165_U125 , P1_R1165_U442 , P1_R1165_U33 );
and AND2_10371 ( P1_R1165_U126 , P1_R1165_U200 , P1_R1165_U197 );
and AND2_10372 ( P1_R1165_U127 , P1_R1165_U313 , P1_R1165_U193 );
and AND2_10373 ( P1_R1165_U128 , P1_R1165_U9 , P1_R1165_U197 );
and AND3_10374 ( P1_R1165_U129 , P1_R1165_U533 , P1_R1165_U532 , P1_R1165_U196 );
and AND2_10375 ( P1_R1165_U130 , P1_R1165_U322 , P1_R1165_U8 );
and AND3_10376 ( P1_R1165_U131 , P1_R1165_U559 , P1_R1165_U558 , P1_R1165_U36 );
and AND2_10377 ( P1_R1165_U132 , P1_R1165_U329 , P1_R1165_U7 );
and AND3_10378 ( P1_R1165_U133 , P1_R1165_U580 , P1_R1165_U579 , P1_R1165_U195 );
and AND2_10379 ( P1_R1165_U134 , P1_R1165_U338 , P1_R1165_U6 );
nand NAND2_10380 ( P1_R1165_U135 , P1_R1165_U599 , P1_R1165_U598 );
not NOT1_10381 ( P1_R1165_U136 , P1_U3201 );
and AND2_10382 ( P1_R1165_U137 , P1_R1165_U369 , P1_R1165_U368 );
not NOT1_10383 ( P1_R1165_U138 , P1_U3206 );
not NOT1_10384 ( P1_R1165_U139 , P1_U3210 );
not NOT1_10385 ( P1_R1165_U140 , P1_U3209 );
not NOT1_10386 ( P1_R1165_U141 , P1_U3207 );
not NOT1_10387 ( P1_R1165_U142 , P1_U3208 );
not NOT1_10388 ( P1_R1165_U143 , P1_U3205 );
not NOT1_10389 ( P1_R1165_U144 , P1_U3203 );
not NOT1_10390 ( P1_R1165_U145 , P1_U3204 );
not NOT1_10391 ( P1_R1165_U146 , P1_U3202 );
nand NAND2_10392 ( P1_R1165_U147 , P1_R1165_U231 , P1_R1165_U230 );
and AND2_10393 ( P1_R1165_U148 , P1_R1165_U403 , P1_R1165_U402 );
nand NAND2_10394 ( P1_R1165_U149 , P1_R1165_U110 , P1_R1165_U227 );
and AND2_10395 ( P1_R1165_U150 , P1_R1165_U417 , P1_R1165_U416 );
nand NAND2_10396 ( P1_R1165_U151 , P1_R1165_U361 , P1_R1165_U350 );
and AND2_10397 ( P1_R1165_U152 , P1_R1165_U424 , P1_R1165_U423 );
nand NAND2_10398 ( P1_R1165_U153 , P1_R1165_U109 , P1_R1165_U214 );
not NOT1_10399 ( P1_R1165_U154 , P1_U3183 );
not NOT1_10400 ( P1_R1165_U155 , P1_U3185 );
not NOT1_10401 ( P1_R1165_U156 , P1_U3184 );
not NOT1_10402 ( P1_R1165_U157 , P1_U3186 );
not NOT1_10403 ( P1_R1165_U158 , P1_U3200 );
not NOT1_10404 ( P1_R1165_U159 , P1_U3197 );
not NOT1_10405 ( P1_R1165_U160 , P1_U3198 );
not NOT1_10406 ( P1_R1165_U161 , P1_U3199 );
not NOT1_10407 ( P1_R1165_U162 , P1_U3196 );
not NOT1_10408 ( P1_R1165_U163 , P1_U3195 );
not NOT1_10409 ( P1_R1165_U164 , P1_U3193 );
not NOT1_10410 ( P1_R1165_U165 , P1_U3194 );
not NOT1_10411 ( P1_R1165_U166 , P1_U3192 );
not NOT1_10412 ( P1_R1165_U167 , P1_U3189 );
not NOT1_10413 ( P1_R1165_U168 , P1_U3190 );
not NOT1_10414 ( P1_R1165_U169 , P1_U3191 );
not NOT1_10415 ( P1_R1165_U170 , P1_U3188 );
not NOT1_10416 ( P1_R1165_U171 , P1_U3187 );
not NOT1_10417 ( P1_R1165_U172 , P1_U3153 );
not NOT1_10418 ( P1_R1165_U173 , P1_U3182 );
and AND2_10419 ( P1_R1165_U174 , P1_R1165_U500 , P1_R1165_U499 );
nand NAND2_10420 ( P1_R1165_U175 , P1_R1165_U124 , P1_R1165_U304 );
nand NAND2_10421 ( P1_R1165_U176 , P1_R1165_U298 , P1_R1165_U297 );
and AND2_10422 ( P1_R1165_U177 , P1_R1165_U519 , P1_R1165_U518 );
nand NAND2_10423 ( P1_R1165_U178 , P1_R1165_U294 , P1_R1165_U293 );
and AND2_10424 ( P1_R1165_U179 , P1_R1165_U526 , P1_R1165_U525 );
nand NAND2_10425 ( P1_R1165_U180 , P1_R1165_U290 , P1_R1165_U289 );
and AND2_10426 ( P1_R1165_U181 , P1_R1165_U540 , P1_R1165_U539 );
nand NAND2_10427 ( P1_R1165_U182 , P1_R1165_U203 , P1_R1165_U202 );
nand NAND2_10428 ( P1_R1165_U183 , P1_R1165_U280 , P1_R1165_U279 );
and AND2_10429 ( P1_R1165_U184 , P1_R1165_U552 , P1_R1165_U551 );
nand NAND2_10430 ( P1_R1165_U185 , P1_R1165_U117 , P1_R1165_U276 );
and AND2_10431 ( P1_R1165_U186 , P1_R1165_U566 , P1_R1165_U565 );
nand NAND2_10432 ( P1_R1165_U187 , P1_R1165_U264 , P1_R1165_U263 );
and AND2_10433 ( P1_R1165_U188 , P1_R1165_U573 , P1_R1165_U572 );
nand NAND2_10434 ( P1_R1165_U189 , P1_R1165_U260 , P1_R1165_U259 );
nand NAND2_10435 ( P1_R1165_U190 , P1_R1165_U250 , P1_R1165_U249 );
and AND2_10436 ( P1_R1165_U191 , P1_R1165_U592 , P1_R1165_U591 );
nand NAND2_10437 ( P1_R1165_U192 , P1_R1165_U363 , P1_R1165_U353 );
nand NAND2_10438 ( P1_R1165_U193 , P1_R1165_U355 , P1_R1165_U354 );
not NOT1_10439 ( P1_R1165_U194 , P1_R1165_U22 );
nand NAND2_10440 ( P1_R1165_U195 , P1_U3169 , P1_R1165_U76 );
nand NAND2_10441 ( P1_R1165_U196 , P1_U3161 , P1_R1165_U82 );
nand NAND2_10442 ( P1_R1165_U197 , P1_U3156 , P1_R1165_U68 );
not NOT1_10443 ( P1_R1165_U198 , P1_R1165_U41 );
not NOT1_10444 ( P1_R1165_U199 , P1_R1165_U48 );
nand NAND2_10445 ( P1_R1165_U200 , P1_U3157 , P1_R1165_U70 );
or OR2_10446 ( P1_R1165_U201 , P1_U3211 , P1_U3181 );
nand NAND2_10447 ( P1_R1165_U202 , P1_R1165_U63 , P1_R1165_U201 );
nand NAND2_10448 ( P1_R1165_U203 , P1_U3181 , P1_U3211 );
not NOT1_10449 ( P1_R1165_U204 , P1_R1165_U182 );
nand NAND2_10450 ( P1_R1165_U205 , P1_R1165_U381 , P1_R1165_U25 );
nand NAND2_10451 ( P1_R1165_U206 , P1_R1165_U205 , P1_R1165_U182 );
nand NAND2_10452 ( P1_R1165_U207 , P1_U3180 , P1_R1165_U64 );
not NOT1_10453 ( P1_R1165_U208 , P1_R1165_U30 );
nand NAND2_10454 ( P1_R1165_U209 , P1_R1165_U384 , P1_R1165_U23 );
nand NAND2_10455 ( P1_R1165_U210 , P1_R1165_U387 , P1_R1165_U21 );
nand NAND2_10456 ( P1_R1165_U211 , P1_R1165_U23 , P1_R1165_U22 );
nand NAND2_10457 ( P1_R1165_U212 , P1_R1165_U62 , P1_R1165_U211 );
nand NAND2_10458 ( P1_R1165_U213 , P1_U3178 , P1_R1165_U194 );
nand NAND2_10459 ( P1_R1165_U214 , P1_R1165_U4 , P1_R1165_U30 );
not NOT1_10460 ( P1_R1165_U215 , P1_R1165_U153 );
nand NAND2_10461 ( P1_R1165_U216 , P1_R1165_U375 , P1_R1165_U20 );
nand NAND2_10462 ( P1_R1165_U217 , P1_R1165_U390 , P1_R1165_U26 );
nand NAND2_10463 ( P1_R1165_U218 , P1_R1165_U217 , P1_R1165_U151 );
nand NAND2_10464 ( P1_R1165_U219 , P1_U3176 , P1_R1165_U65 );
not NOT1_10465 ( P1_R1165_U220 , P1_R1165_U29 );
nand NAND2_10466 ( P1_R1165_U221 , P1_R1165_U393 , P1_R1165_U19 );
nand NAND2_10467 ( P1_R1165_U222 , P1_R1165_U396 , P1_R1165_U17 );
not NOT1_10468 ( P1_R1165_U223 , P1_R1165_U18 );
nand NAND2_10469 ( P1_R1165_U224 , P1_R1165_U19 , P1_R1165_U18 );
nand NAND2_10470 ( P1_R1165_U225 , P1_R1165_U59 , P1_R1165_U224 );
nand NAND2_10471 ( P1_R1165_U226 , P1_U3174 , P1_R1165_U223 );
nand NAND2_10472 ( P1_R1165_U227 , P1_R1165_U5 , P1_R1165_U29 );
not NOT1_10473 ( P1_R1165_U228 , P1_R1165_U149 );
nand NAND2_10474 ( P1_R1165_U229 , P1_R1165_U399 , P1_R1165_U27 );
nand NAND2_10475 ( P1_R1165_U230 , P1_R1165_U229 , P1_R1165_U149 );
nand NAND2_10476 ( P1_R1165_U231 , P1_U3173 , P1_R1165_U66 );
not NOT1_10477 ( P1_R1165_U232 , P1_R1165_U147 );
nand NAND2_10478 ( P1_R1165_U233 , P1_R1165_U396 , P1_R1165_U17 );
nand NAND2_10479 ( P1_R1165_U234 , P1_R1165_U233 , P1_R1165_U29 );
nand NAND2_10480 ( P1_R1165_U235 , P1_R1165_U111 , P1_R1165_U234 );
nand NAND2_10481 ( P1_R1165_U236 , P1_R1165_U220 , P1_R1165_U18 );
nand NAND2_10482 ( P1_R1165_U237 , P1_U3174 , P1_R1165_U59 );
nand NAND2_10483 ( P1_R1165_U238 , P1_R1165_U112 , P1_R1165_U236 );
nand NAND2_10484 ( P1_R1165_U239 , P1_R1165_U396 , P1_R1165_U17 );
nand NAND2_10485 ( P1_R1165_U240 , P1_R1165_U387 , P1_R1165_U21 );
nand NAND2_10486 ( P1_R1165_U241 , P1_R1165_U240 , P1_R1165_U30 );
nand NAND2_10487 ( P1_R1165_U242 , P1_R1165_U113 , P1_R1165_U241 );
nand NAND2_10488 ( P1_R1165_U243 , P1_R1165_U208 , P1_R1165_U22 );
nand NAND2_10489 ( P1_R1165_U244 , P1_U3178 , P1_R1165_U62 );
nand NAND2_10490 ( P1_R1165_U245 , P1_R1165_U114 , P1_R1165_U243 );
nand NAND2_10491 ( P1_R1165_U246 , P1_R1165_U387 , P1_R1165_U21 );
nand NAND2_10492 ( P1_R1165_U247 , P1_R1165_U367 , P1_R1165_U28 );
nand NAND2_10493 ( P1_R1165_U248 , P1_R1165_U451 , P1_R1165_U38 );
nand NAND2_10494 ( P1_R1165_U249 , P1_R1165_U248 , P1_R1165_U192 );
nand NAND2_10495 ( P1_R1165_U250 , P1_U3171 , P1_R1165_U73 );
not NOT1_10496 ( P1_R1165_U251 , P1_R1165_U190 );
nand NAND2_10497 ( P1_R1165_U252 , P1_R1165_U454 , P1_R1165_U42 );
nand NAND2_10498 ( P1_R1165_U253 , P1_R1165_U457 , P1_R1165_U39 );
nand NAND2_10499 ( P1_R1165_U254 , P1_R1165_U198 , P1_R1165_U6 );
nand NAND2_10500 ( P1_R1165_U255 , P1_U3168 , P1_R1165_U75 );
nand NAND2_10501 ( P1_R1165_U256 , P1_R1165_U116 , P1_R1165_U254 );
nand NAND2_10502 ( P1_R1165_U257 , P1_R1165_U460 , P1_R1165_U40 );
nand NAND2_10503 ( P1_R1165_U258 , P1_R1165_U454 , P1_R1165_U42 );
nand NAND2_10504 ( P1_R1165_U259 , P1_R1165_U115 , P1_R1165_U190 );
nand NAND2_10505 ( P1_R1165_U260 , P1_R1165_U258 , P1_R1165_U256 );
not NOT1_10506 ( P1_R1165_U261 , P1_R1165_U189 );
nand NAND2_10507 ( P1_R1165_U262 , P1_R1165_U463 , P1_R1165_U43 );
nand NAND2_10508 ( P1_R1165_U263 , P1_R1165_U262 , P1_R1165_U189 );
nand NAND2_10509 ( P1_R1165_U264 , P1_U3167 , P1_R1165_U77 );
not NOT1_10510 ( P1_R1165_U265 , P1_R1165_U187 );
nand NAND2_10511 ( P1_R1165_U266 , P1_R1165_U466 , P1_R1165_U44 );
nand NAND2_10512 ( P1_R1165_U267 , P1_R1165_U266 , P1_R1165_U187 );
nand NAND2_10513 ( P1_R1165_U268 , P1_U3166 , P1_R1165_U78 );
not NOT1_10514 ( P1_R1165_U269 , P1_R1165_U55 );
nand NAND2_10515 ( P1_R1165_U270 , P1_R1165_U469 , P1_R1165_U37 );
nand NAND2_10516 ( P1_R1165_U271 , P1_R1165_U472 , P1_R1165_U35 );
not NOT1_10517 ( P1_R1165_U272 , P1_R1165_U36 );
nand NAND2_10518 ( P1_R1165_U273 , P1_R1165_U37 , P1_R1165_U36 );
nand NAND2_10519 ( P1_R1165_U274 , P1_R1165_U72 , P1_R1165_U273 );
nand NAND2_10520 ( P1_R1165_U275 , P1_U3164 , P1_R1165_U272 );
nand NAND2_10521 ( P1_R1165_U276 , P1_R1165_U7 , P1_R1165_U55 );
not NOT1_10522 ( P1_R1165_U277 , P1_R1165_U185 );
nand NAND2_10523 ( P1_R1165_U278 , P1_R1165_U475 , P1_R1165_U45 );
nand NAND2_10524 ( P1_R1165_U279 , P1_R1165_U278 , P1_R1165_U185 );
nand NAND2_10525 ( P1_R1165_U280 , P1_U3163 , P1_R1165_U79 );
not NOT1_10526 ( P1_R1165_U281 , P1_R1165_U183 );
nand NAND2_10527 ( P1_R1165_U282 , P1_R1165_U478 , P1_R1165_U49 );
nand NAND2_10528 ( P1_R1165_U283 , P1_R1165_U481 , P1_R1165_U46 );
nand NAND2_10529 ( P1_R1165_U284 , P1_R1165_U199 , P1_R1165_U8 );
nand NAND2_10530 ( P1_R1165_U285 , P1_U3160 , P1_R1165_U81 );
nand NAND2_10531 ( P1_R1165_U286 , P1_R1165_U119 , P1_R1165_U284 );
nand NAND2_10532 ( P1_R1165_U287 , P1_R1165_U484 , P1_R1165_U47 );
nand NAND2_10533 ( P1_R1165_U288 , P1_R1165_U478 , P1_R1165_U49 );
nand NAND2_10534 ( P1_R1165_U289 , P1_R1165_U118 , P1_R1165_U183 );
nand NAND2_10535 ( P1_R1165_U290 , P1_R1165_U288 , P1_R1165_U286 );
not NOT1_10536 ( P1_R1165_U291 , P1_R1165_U180 );
nand NAND2_10537 ( P1_R1165_U292 , P1_R1165_U487 , P1_R1165_U50 );
nand NAND2_10538 ( P1_R1165_U293 , P1_R1165_U292 , P1_R1165_U180 );
nand NAND2_10539 ( P1_R1165_U294 , P1_U3159 , P1_R1165_U83 );
not NOT1_10540 ( P1_R1165_U295 , P1_R1165_U178 );
nand NAND2_10541 ( P1_R1165_U296 , P1_R1165_U490 , P1_R1165_U51 );
nand NAND2_10542 ( P1_R1165_U297 , P1_R1165_U296 , P1_R1165_U178 );
nand NAND2_10543 ( P1_R1165_U298 , P1_U3158 , P1_R1165_U84 );
not NOT1_10544 ( P1_R1165_U299 , P1_R1165_U176 );
nand NAND2_10545 ( P1_R1165_U300 , P1_R1165_U442 , P1_R1165_U33 );
nand NAND2_10546 ( P1_R1165_U301 , P1_R1165_U200 , P1_R1165_U197 );
not NOT1_10547 ( P1_R1165_U302 , P1_R1165_U52 );
nand NAND2_10548 ( P1_R1165_U303 , P1_R1165_U448 , P1_R1165_U34 );
nand NAND3_10549 ( P1_R1165_U304 , P1_R1165_U176 , P1_R1165_U303 , P1_R1165_U193 );
not NOT1_10550 ( P1_R1165_U305 , P1_R1165_U175 );
nand NAND2_10551 ( P1_R1165_U306 , P1_R1165_U439 , P1_R1165_U31 );
nand NAND2_10552 ( P1_R1165_U307 , P1_U3154 , P1_R1165_U67 );
nand NAND2_10553 ( P1_R1165_U308 , P1_R1165_U439 , P1_R1165_U31 );
nand NAND2_10554 ( P1_R1165_U309 , P1_R1165_U303 , P1_R1165_U176 );
not NOT1_10555 ( P1_R1165_U310 , P1_R1165_U53 );
nand NAND2_10556 ( P1_R1165_U311 , P1_R1165_U125 , P1_R1165_U9 );
nand NAND2_10557 ( P1_R1165_U312 , P1_R1165_U126 , P1_R1165_U309 );
nand NAND2_10558 ( P1_R1165_U313 , P1_U3155 , P1_R1165_U69 );
nand NAND2_10559 ( P1_R1165_U314 , P1_R1165_U127 , P1_R1165_U312 );
nand NAND2_10560 ( P1_R1165_U315 , P1_R1165_U442 , P1_R1165_U33 );
nand NAND2_10561 ( P1_R1165_U316 , P1_R1165_U287 , P1_R1165_U183 );
not NOT1_10562 ( P1_R1165_U317 , P1_R1165_U54 );
nand NAND2_10563 ( P1_R1165_U318 , P1_R1165_U481 , P1_R1165_U46 );
nand NAND2_10564 ( P1_R1165_U319 , P1_R1165_U318 , P1_R1165_U54 );
nand NAND2_10565 ( P1_R1165_U320 , P1_R1165_U129 , P1_R1165_U319 );
nand NAND2_10566 ( P1_R1165_U321 , P1_R1165_U317 , P1_R1165_U196 );
nand NAND2_10567 ( P1_R1165_U322 , P1_U3160 , P1_R1165_U81 );
nand NAND2_10568 ( P1_R1165_U323 , P1_R1165_U130 , P1_R1165_U321 );
nand NAND2_10569 ( P1_R1165_U324 , P1_R1165_U481 , P1_R1165_U46 );
nand NAND2_10570 ( P1_R1165_U325 , P1_R1165_U472 , P1_R1165_U35 );
nand NAND2_10571 ( P1_R1165_U326 , P1_R1165_U325 , P1_R1165_U55 );
nand NAND2_10572 ( P1_R1165_U327 , P1_R1165_U131 , P1_R1165_U326 );
nand NAND2_10573 ( P1_R1165_U328 , P1_R1165_U269 , P1_R1165_U36 );
nand NAND2_10574 ( P1_R1165_U329 , P1_U3164 , P1_R1165_U72 );
nand NAND2_10575 ( P1_R1165_U330 , P1_R1165_U132 , P1_R1165_U328 );
nand NAND2_10576 ( P1_R1165_U331 , P1_R1165_U472 , P1_R1165_U35 );
nand NAND2_10577 ( P1_R1165_U332 , P1_R1165_U257 , P1_R1165_U190 );
not NOT1_10578 ( P1_R1165_U333 , P1_R1165_U56 );
nand NAND2_10579 ( P1_R1165_U334 , P1_R1165_U457 , P1_R1165_U39 );
nand NAND2_10580 ( P1_R1165_U335 , P1_R1165_U334 , P1_R1165_U56 );
nand NAND2_10581 ( P1_R1165_U336 , P1_R1165_U133 , P1_R1165_U335 );
nand NAND2_10582 ( P1_R1165_U337 , P1_R1165_U333 , P1_R1165_U195 );
nand NAND2_10583 ( P1_R1165_U338 , P1_U3168 , P1_R1165_U75 );
nand NAND2_10584 ( P1_R1165_U339 , P1_R1165_U134 , P1_R1165_U337 );
nand NAND2_10585 ( P1_R1165_U340 , P1_R1165_U457 , P1_R1165_U39 );
nand NAND2_10586 ( P1_R1165_U341 , P1_R1165_U239 , P1_R1165_U18 );
nand NAND2_10587 ( P1_R1165_U342 , P1_R1165_U246 , P1_R1165_U22 );
nand NAND2_10588 ( P1_R1165_U343 , P1_R1165_U315 , P1_R1165_U197 );
nand NAND2_10589 ( P1_R1165_U344 , P1_R1165_U303 , P1_R1165_U200 );
nand NAND2_10590 ( P1_R1165_U345 , P1_R1165_U324 , P1_R1165_U196 );
nand NAND2_10591 ( P1_R1165_U346 , P1_R1165_U287 , P1_R1165_U48 );
nand NAND2_10592 ( P1_R1165_U347 , P1_R1165_U331 , P1_R1165_U36 );
nand NAND2_10593 ( P1_R1165_U348 , P1_R1165_U340 , P1_R1165_U195 );
nand NAND2_10594 ( P1_R1165_U349 , P1_R1165_U257 , P1_R1165_U41 );
nand NAND2_10595 ( P1_R1165_U350 , P1_U3177 , P1_R1165_U60 );
nand NAND3_10596 ( P1_R1165_U351 , P1_R1165_U352 , P1_R1165_U304 , P1_R1165_U120 );
nand NAND2_10597 ( P1_R1165_U352 , P1_R1165_U301 , P1_R1165_U193 );
nand NAND2_10598 ( P1_R1165_U353 , P1_U3172 , P1_R1165_U57 );
nand NAND2_10599 ( P1_R1165_U354 , P1_R1165_U69 , P1_R1165_U300 );
nand NAND2_10600 ( P1_R1165_U355 , P1_U3155 , P1_R1165_U300 );
nand NAND3_10601 ( P1_R1165_U356 , P1_R1165_U301 , P1_R1165_U193 , P1_R1165_U308 );
nand NAND3_10602 ( P1_R1165_U357 , P1_R1165_U176 , P1_R1165_U193 , P1_R1165_U121 );
nand NAND2_10603 ( P1_R1165_U358 , P1_R1165_U302 , P1_R1165_U308 );
nand NAND2_10604 ( P1_R1165_U359 , P1_U3154 , P1_R1165_U67 );
nand NAND2_10605 ( P1_R1165_U360 , P1_R1165_U128 , P1_R1165_U310 );
nand NAND2_10606 ( P1_R1165_U361 , P1_R1165_U216 , P1_R1165_U153 );
not NOT1_10607 ( P1_R1165_U362 , P1_R1165_U151 );
nand NAND2_10608 ( P1_R1165_U363 , P1_R1165_U247 , P1_R1165_U147 );
not NOT1_10609 ( P1_R1165_U364 , P1_R1165_U192 );
nand NAND2_10610 ( P1_R1165_U365 , P1_U3211 , P1_R1165_U136 );
nand NAND2_10611 ( P1_R1165_U366 , P1_U3201 , P1_R1165_U16 );
not NOT1_10612 ( P1_R1165_U367 , P1_R1165_U57 );
nand NAND2_10613 ( P1_R1165_U368 , P1_R1165_U367 , P1_U3172 );
nand NAND2_10614 ( P1_R1165_U369 , P1_R1165_U57 , P1_R1165_U28 );
nand NAND2_10615 ( P1_R1165_U370 , P1_R1165_U367 , P1_U3172 );
nand NAND2_10616 ( P1_R1165_U371 , P1_R1165_U57 , P1_R1165_U28 );
nand NAND2_10617 ( P1_R1165_U372 , P1_R1165_U371 , P1_R1165_U370 );
nand NAND2_10618 ( P1_R1165_U373 , P1_U3211 , P1_R1165_U138 );
nand NAND2_10619 ( P1_R1165_U374 , P1_U3206 , P1_R1165_U16 );
not NOT1_10620 ( P1_R1165_U375 , P1_R1165_U60 );
nand NAND2_10621 ( P1_R1165_U376 , P1_U3211 , P1_R1165_U139 );
nand NAND2_10622 ( P1_R1165_U377 , P1_U3210 , P1_R1165_U16 );
not NOT1_10623 ( P1_R1165_U378 , P1_R1165_U63 );
nand NAND2_10624 ( P1_R1165_U379 , P1_U3211 , P1_R1165_U140 );
nand NAND2_10625 ( P1_R1165_U380 , P1_U3209 , P1_R1165_U16 );
not NOT1_10626 ( P1_R1165_U381 , P1_R1165_U64 );
nand NAND2_10627 ( P1_R1165_U382 , P1_U3211 , P1_R1165_U141 );
nand NAND2_10628 ( P1_R1165_U383 , P1_U3207 , P1_R1165_U16 );
not NOT1_10629 ( P1_R1165_U384 , P1_R1165_U62 );
nand NAND2_10630 ( P1_R1165_U385 , P1_U3211 , P1_R1165_U142 );
nand NAND2_10631 ( P1_R1165_U386 , P1_U3208 , P1_R1165_U16 );
not NOT1_10632 ( P1_R1165_U387 , P1_R1165_U61 );
nand NAND2_10633 ( P1_R1165_U388 , P1_U3211 , P1_R1165_U143 );
nand NAND2_10634 ( P1_R1165_U389 , P1_U3205 , P1_R1165_U16 );
not NOT1_10635 ( P1_R1165_U390 , P1_R1165_U65 );
nand NAND2_10636 ( P1_R1165_U391 , P1_U3211 , P1_R1165_U144 );
nand NAND2_10637 ( P1_R1165_U392 , P1_U3203 , P1_R1165_U16 );
not NOT1_10638 ( P1_R1165_U393 , P1_R1165_U59 );
nand NAND2_10639 ( P1_R1165_U394 , P1_U3211 , P1_R1165_U145 );
nand NAND2_10640 ( P1_R1165_U395 , P1_U3204 , P1_R1165_U16 );
not NOT1_10641 ( P1_R1165_U396 , P1_R1165_U58 );
nand NAND2_10642 ( P1_R1165_U397 , P1_U3211 , P1_R1165_U146 );
nand NAND2_10643 ( P1_R1165_U398 , P1_U3202 , P1_R1165_U16 );
not NOT1_10644 ( P1_R1165_U399 , P1_R1165_U66 );
nand NAND2_10645 ( P1_R1165_U400 , P1_R1165_U137 , P1_R1165_U147 );
nand NAND2_10646 ( P1_R1165_U401 , P1_R1165_U232 , P1_R1165_U372 );
nand NAND2_10647 ( P1_R1165_U402 , P1_R1165_U399 , P1_U3173 );
nand NAND2_10648 ( P1_R1165_U403 , P1_R1165_U66 , P1_R1165_U27 );
nand NAND2_10649 ( P1_R1165_U404 , P1_R1165_U399 , P1_U3173 );
nand NAND2_10650 ( P1_R1165_U405 , P1_R1165_U66 , P1_R1165_U27 );
nand NAND2_10651 ( P1_R1165_U406 , P1_R1165_U405 , P1_R1165_U404 );
nand NAND2_10652 ( P1_R1165_U407 , P1_R1165_U148 , P1_R1165_U149 );
nand NAND2_10653 ( P1_R1165_U408 , P1_R1165_U228 , P1_R1165_U406 );
nand NAND2_10654 ( P1_R1165_U409 , P1_R1165_U393 , P1_U3174 );
nand NAND2_10655 ( P1_R1165_U410 , P1_R1165_U59 , P1_R1165_U19 );
nand NAND2_10656 ( P1_R1165_U411 , P1_R1165_U396 , P1_U3175 );
nand NAND2_10657 ( P1_R1165_U412 , P1_R1165_U58 , P1_R1165_U17 );
nand NAND2_10658 ( P1_R1165_U413 , P1_R1165_U412 , P1_R1165_U411 );
nand NAND2_10659 ( P1_R1165_U414 , P1_R1165_U341 , P1_R1165_U29 );
nand NAND2_10660 ( P1_R1165_U415 , P1_R1165_U413 , P1_R1165_U220 );
nand NAND2_10661 ( P1_R1165_U416 , P1_R1165_U390 , P1_U3176 );
nand NAND2_10662 ( P1_R1165_U417 , P1_R1165_U65 , P1_R1165_U26 );
nand NAND2_10663 ( P1_R1165_U418 , P1_R1165_U390 , P1_U3176 );
nand NAND2_10664 ( P1_R1165_U419 , P1_R1165_U65 , P1_R1165_U26 );
nand NAND2_10665 ( P1_R1165_U420 , P1_R1165_U419 , P1_R1165_U418 );
nand NAND2_10666 ( P1_R1165_U421 , P1_R1165_U150 , P1_R1165_U151 );
nand NAND2_10667 ( P1_R1165_U422 , P1_R1165_U362 , P1_R1165_U420 );
nand NAND2_10668 ( P1_R1165_U423 , P1_R1165_U375 , P1_U3177 );
nand NAND2_10669 ( P1_R1165_U424 , P1_R1165_U60 , P1_R1165_U20 );
nand NAND2_10670 ( P1_R1165_U425 , P1_R1165_U375 , P1_U3177 );
nand NAND2_10671 ( P1_R1165_U426 , P1_R1165_U60 , P1_R1165_U20 );
nand NAND2_10672 ( P1_R1165_U427 , P1_R1165_U426 , P1_R1165_U425 );
nand NAND2_10673 ( P1_R1165_U428 , P1_R1165_U152 , P1_R1165_U153 );
nand NAND2_10674 ( P1_R1165_U429 , P1_R1165_U215 , P1_R1165_U427 );
nand NAND2_10675 ( P1_R1165_U430 , P1_R1165_U384 , P1_U3178 );
nand NAND2_10676 ( P1_R1165_U431 , P1_R1165_U62 , P1_R1165_U23 );
nand NAND2_10677 ( P1_R1165_U432 , P1_R1165_U387 , P1_U3179 );
nand NAND2_10678 ( P1_R1165_U433 , P1_R1165_U61 , P1_R1165_U21 );
nand NAND2_10679 ( P1_R1165_U434 , P1_R1165_U433 , P1_R1165_U432 );
nand NAND2_10680 ( P1_R1165_U435 , P1_R1165_U342 , P1_R1165_U30 );
nand NAND2_10681 ( P1_R1165_U436 , P1_R1165_U434 , P1_R1165_U208 );
nand NAND2_10682 ( P1_R1165_U437 , P1_U3211 , P1_R1165_U154 );
nand NAND2_10683 ( P1_R1165_U438 , P1_U3183 , P1_R1165_U16 );
not NOT1_10684 ( P1_R1165_U439 , P1_R1165_U67 );
nand NAND2_10685 ( P1_R1165_U440 , P1_U3211 , P1_R1165_U155 );
nand NAND2_10686 ( P1_R1165_U441 , P1_U3185 , P1_R1165_U16 );
not NOT1_10687 ( P1_R1165_U442 , P1_R1165_U68 );
nand NAND2_10688 ( P1_R1165_U443 , P1_U3211 , P1_R1165_U156 );
nand NAND2_10689 ( P1_R1165_U444 , P1_U3184 , P1_R1165_U16 );
not NOT1_10690 ( P1_R1165_U445 , P1_R1165_U69 );
nand NAND2_10691 ( P1_R1165_U446 , P1_U3211 , P1_R1165_U157 );
nand NAND2_10692 ( P1_R1165_U447 , P1_U3186 , P1_R1165_U16 );
not NOT1_10693 ( P1_R1165_U448 , P1_R1165_U70 );
nand NAND2_10694 ( P1_R1165_U449 , P1_U3211 , P1_R1165_U158 );
nand NAND2_10695 ( P1_R1165_U450 , P1_U3200 , P1_R1165_U16 );
not NOT1_10696 ( P1_R1165_U451 , P1_R1165_U73 );
nand NAND2_10697 ( P1_R1165_U452 , P1_U3211 , P1_R1165_U159 );
nand NAND2_10698 ( P1_R1165_U453 , P1_U3197 , P1_R1165_U16 );
not NOT1_10699 ( P1_R1165_U454 , P1_R1165_U75 );
nand NAND2_10700 ( P1_R1165_U455 , P1_U3211 , P1_R1165_U160 );
nand NAND2_10701 ( P1_R1165_U456 , P1_U3198 , P1_R1165_U16 );
not NOT1_10702 ( P1_R1165_U457 , P1_R1165_U76 );
nand NAND2_10703 ( P1_R1165_U458 , P1_U3211 , P1_R1165_U161 );
nand NAND2_10704 ( P1_R1165_U459 , P1_U3199 , P1_R1165_U16 );
not NOT1_10705 ( P1_R1165_U460 , P1_R1165_U74 );
nand NAND2_10706 ( P1_R1165_U461 , P1_U3211 , P1_R1165_U162 );
nand NAND2_10707 ( P1_R1165_U462 , P1_U3196 , P1_R1165_U16 );
not NOT1_10708 ( P1_R1165_U463 , P1_R1165_U77 );
nand NAND2_10709 ( P1_R1165_U464 , P1_U3211 , P1_R1165_U163 );
nand NAND2_10710 ( P1_R1165_U465 , P1_U3195 , P1_R1165_U16 );
not NOT1_10711 ( P1_R1165_U466 , P1_R1165_U78 );
nand NAND2_10712 ( P1_R1165_U467 , P1_U3211 , P1_R1165_U164 );
nand NAND2_10713 ( P1_R1165_U468 , P1_U3193 , P1_R1165_U16 );
not NOT1_10714 ( P1_R1165_U469 , P1_R1165_U72 );
nand NAND2_10715 ( P1_R1165_U470 , P1_U3211 , P1_R1165_U165 );
nand NAND2_10716 ( P1_R1165_U471 , P1_U3194 , P1_R1165_U16 );
not NOT1_10717 ( P1_R1165_U472 , P1_R1165_U71 );
nand NAND2_10718 ( P1_R1165_U473 , P1_U3211 , P1_R1165_U166 );
nand NAND2_10719 ( P1_R1165_U474 , P1_U3192 , P1_R1165_U16 );
not NOT1_10720 ( P1_R1165_U475 , P1_R1165_U79 );
nand NAND2_10721 ( P1_R1165_U476 , P1_U3211 , P1_R1165_U167 );
nand NAND2_10722 ( P1_R1165_U477 , P1_U3189 , P1_R1165_U16 );
not NOT1_10723 ( P1_R1165_U478 , P1_R1165_U81 );
nand NAND2_10724 ( P1_R1165_U479 , P1_U3211 , P1_R1165_U168 );
nand NAND2_10725 ( P1_R1165_U480 , P1_U3190 , P1_R1165_U16 );
not NOT1_10726 ( P1_R1165_U481 , P1_R1165_U82 );
nand NAND2_10727 ( P1_R1165_U482 , P1_U3211 , P1_R1165_U169 );
nand NAND2_10728 ( P1_R1165_U483 , P1_U3191 , P1_R1165_U16 );
not NOT1_10729 ( P1_R1165_U484 , P1_R1165_U80 );
nand NAND2_10730 ( P1_R1165_U485 , P1_U3211 , P1_R1165_U170 );
nand NAND2_10731 ( P1_R1165_U486 , P1_U3188 , P1_R1165_U16 );
not NOT1_10732 ( P1_R1165_U487 , P1_R1165_U83 );
nand NAND2_10733 ( P1_R1165_U488 , P1_U3211 , P1_R1165_U171 );
nand NAND2_10734 ( P1_R1165_U489 , P1_U3187 , P1_R1165_U16 );
not NOT1_10735 ( P1_R1165_U490 , P1_R1165_U84 );
nand NAND2_10736 ( P1_R1165_U491 , P1_U3211 , P1_R1165_U172 );
nand NAND2_10737 ( P1_R1165_U492 , P1_U3153 , P1_R1165_U16 );
not NOT1_10738 ( P1_R1165_U493 , P1_R1165_U123 );
nand NAND2_10739 ( P1_R1165_U494 , P1_U3182 , P1_R1165_U493 );
nand NAND2_10740 ( P1_R1165_U495 , P1_R1165_U123 , P1_R1165_U173 );
not NOT1_10741 ( P1_R1165_U496 , P1_R1165_U85 );
nand NAND3_10742 ( P1_R1165_U497 , P1_R1165_U351 , P1_R1165_U306 , P1_R1165_U496 );
nand NAND4_10743 ( P1_R1165_U498 , P1_R1165_U358 , P1_R1165_U357 , P1_R1165_U122 , P1_R1165_U85 );
nand NAND2_10744 ( P1_R1165_U499 , P1_R1165_U439 , P1_U3154 );
nand NAND2_10745 ( P1_R1165_U500 , P1_R1165_U67 , P1_R1165_U31 );
nand NAND2_10746 ( P1_R1165_U501 , P1_R1165_U439 , P1_U3154 );
nand NAND2_10747 ( P1_R1165_U502 , P1_R1165_U67 , P1_R1165_U31 );
nand NAND2_10748 ( P1_R1165_U503 , P1_R1165_U502 , P1_R1165_U501 );
nand NAND2_10749 ( P1_R1165_U504 , P1_R1165_U174 , P1_R1165_U175 );
nand NAND2_10750 ( P1_R1165_U505 , P1_R1165_U305 , P1_R1165_U503 );
nand NAND2_10751 ( P1_R1165_U506 , P1_R1165_U445 , P1_U3155 );
nand NAND2_10752 ( P1_R1165_U507 , P1_R1165_U69 , P1_R1165_U32 );
nand NAND2_10753 ( P1_R1165_U508 , P1_R1165_U442 , P1_U3156 );
nand NAND2_10754 ( P1_R1165_U509 , P1_R1165_U68 , P1_R1165_U33 );
nand NAND2_10755 ( P1_R1165_U510 , P1_R1165_U509 , P1_R1165_U508 );
nand NAND2_10756 ( P1_R1165_U511 , P1_R1165_U343 , P1_R1165_U53 );
nand NAND2_10757 ( P1_R1165_U512 , P1_R1165_U510 , P1_R1165_U310 );
nand NAND2_10758 ( P1_R1165_U513 , P1_R1165_U448 , P1_U3157 );
nand NAND2_10759 ( P1_R1165_U514 , P1_R1165_U70 , P1_R1165_U34 );
nand NAND2_10760 ( P1_R1165_U515 , P1_R1165_U514 , P1_R1165_U513 );
nand NAND2_10761 ( P1_R1165_U516 , P1_R1165_U344 , P1_R1165_U176 );
nand NAND2_10762 ( P1_R1165_U517 , P1_R1165_U299 , P1_R1165_U515 );
nand NAND2_10763 ( P1_R1165_U518 , P1_R1165_U490 , P1_U3158 );
nand NAND2_10764 ( P1_R1165_U519 , P1_R1165_U84 , P1_R1165_U51 );
nand NAND2_10765 ( P1_R1165_U520 , P1_R1165_U490 , P1_U3158 );
nand NAND2_10766 ( P1_R1165_U521 , P1_R1165_U84 , P1_R1165_U51 );
nand NAND2_10767 ( P1_R1165_U522 , P1_R1165_U521 , P1_R1165_U520 );
nand NAND2_10768 ( P1_R1165_U523 , P1_R1165_U177 , P1_R1165_U178 );
nand NAND2_10769 ( P1_R1165_U524 , P1_R1165_U295 , P1_R1165_U522 );
nand NAND2_10770 ( P1_R1165_U525 , P1_R1165_U487 , P1_U3159 );
nand NAND2_10771 ( P1_R1165_U526 , P1_R1165_U83 , P1_R1165_U50 );
nand NAND2_10772 ( P1_R1165_U527 , P1_R1165_U487 , P1_U3159 );
nand NAND2_10773 ( P1_R1165_U528 , P1_R1165_U83 , P1_R1165_U50 );
nand NAND2_10774 ( P1_R1165_U529 , P1_R1165_U528 , P1_R1165_U527 );
nand NAND2_10775 ( P1_R1165_U530 , P1_R1165_U179 , P1_R1165_U180 );
nand NAND2_10776 ( P1_R1165_U531 , P1_R1165_U291 , P1_R1165_U529 );
nand NAND2_10777 ( P1_R1165_U532 , P1_R1165_U478 , P1_U3160 );
nand NAND2_10778 ( P1_R1165_U533 , P1_R1165_U81 , P1_R1165_U49 );
nand NAND2_10779 ( P1_R1165_U534 , P1_R1165_U481 , P1_U3161 );
nand NAND2_10780 ( P1_R1165_U535 , P1_R1165_U82 , P1_R1165_U46 );
nand NAND2_10781 ( P1_R1165_U536 , P1_R1165_U535 , P1_R1165_U534 );
nand NAND2_10782 ( P1_R1165_U537 , P1_R1165_U345 , P1_R1165_U54 );
nand NAND2_10783 ( P1_R1165_U538 , P1_R1165_U536 , P1_R1165_U317 );
nand NAND2_10784 ( P1_R1165_U539 , P1_R1165_U381 , P1_U3180 );
nand NAND2_10785 ( P1_R1165_U540 , P1_R1165_U64 , P1_R1165_U25 );
nand NAND2_10786 ( P1_R1165_U541 , P1_R1165_U381 , P1_U3180 );
nand NAND2_10787 ( P1_R1165_U542 , P1_R1165_U64 , P1_R1165_U25 );
nand NAND2_10788 ( P1_R1165_U543 , P1_R1165_U542 , P1_R1165_U541 );
nand NAND2_10789 ( P1_R1165_U544 , P1_R1165_U181 , P1_R1165_U182 );
nand NAND2_10790 ( P1_R1165_U545 , P1_R1165_U204 , P1_R1165_U543 );
nand NAND2_10791 ( P1_R1165_U546 , P1_R1165_U484 , P1_U3162 );
nand NAND2_10792 ( P1_R1165_U547 , P1_R1165_U80 , P1_R1165_U47 );
nand NAND2_10793 ( P1_R1165_U548 , P1_R1165_U547 , P1_R1165_U546 );
nand NAND2_10794 ( P1_R1165_U549 , P1_R1165_U346 , P1_R1165_U183 );
nand NAND2_10795 ( P1_R1165_U550 , P1_R1165_U281 , P1_R1165_U548 );
nand NAND2_10796 ( P1_R1165_U551 , P1_R1165_U475 , P1_U3163 );
nand NAND2_10797 ( P1_R1165_U552 , P1_R1165_U79 , P1_R1165_U45 );
nand NAND2_10798 ( P1_R1165_U553 , P1_R1165_U475 , P1_U3163 );
nand NAND2_10799 ( P1_R1165_U554 , P1_R1165_U79 , P1_R1165_U45 );
nand NAND2_10800 ( P1_R1165_U555 , P1_R1165_U554 , P1_R1165_U553 );
nand NAND2_10801 ( P1_R1165_U556 , P1_R1165_U184 , P1_R1165_U185 );
nand NAND2_10802 ( P1_R1165_U557 , P1_R1165_U277 , P1_R1165_U555 );
nand NAND2_10803 ( P1_R1165_U558 , P1_R1165_U469 , P1_U3164 );
nand NAND2_10804 ( P1_R1165_U559 , P1_R1165_U72 , P1_R1165_U37 );
nand NAND2_10805 ( P1_R1165_U560 , P1_R1165_U472 , P1_U3165 );
nand NAND2_10806 ( P1_R1165_U561 , P1_R1165_U71 , P1_R1165_U35 );
nand NAND2_10807 ( P1_R1165_U562 , P1_R1165_U561 , P1_R1165_U560 );
nand NAND2_10808 ( P1_R1165_U563 , P1_R1165_U347 , P1_R1165_U55 );
nand NAND2_10809 ( P1_R1165_U564 , P1_R1165_U562 , P1_R1165_U269 );
nand NAND2_10810 ( P1_R1165_U565 , P1_R1165_U466 , P1_U3166 );
nand NAND2_10811 ( P1_R1165_U566 , P1_R1165_U78 , P1_R1165_U44 );
nand NAND2_10812 ( P1_R1165_U567 , P1_R1165_U466 , P1_U3166 );
nand NAND2_10813 ( P1_R1165_U568 , P1_R1165_U78 , P1_R1165_U44 );
nand NAND2_10814 ( P1_R1165_U569 , P1_R1165_U568 , P1_R1165_U567 );
nand NAND2_10815 ( P1_R1165_U570 , P1_R1165_U186 , P1_R1165_U187 );
nand NAND2_10816 ( P1_R1165_U571 , P1_R1165_U265 , P1_R1165_U569 );
nand NAND2_10817 ( P1_R1165_U572 , P1_R1165_U463 , P1_U3167 );
nand NAND2_10818 ( P1_R1165_U573 , P1_R1165_U77 , P1_R1165_U43 );
nand NAND2_10819 ( P1_R1165_U574 , P1_R1165_U463 , P1_U3167 );
nand NAND2_10820 ( P1_R1165_U575 , P1_R1165_U77 , P1_R1165_U43 );
nand NAND2_10821 ( P1_R1165_U576 , P1_R1165_U575 , P1_R1165_U574 );
nand NAND2_10822 ( P1_R1165_U577 , P1_R1165_U188 , P1_R1165_U189 );
nand NAND2_10823 ( P1_R1165_U578 , P1_R1165_U261 , P1_R1165_U576 );
nand NAND2_10824 ( P1_R1165_U579 , P1_R1165_U454 , P1_U3168 );
nand NAND2_10825 ( P1_R1165_U580 , P1_R1165_U75 , P1_R1165_U42 );
nand NAND2_10826 ( P1_R1165_U581 , P1_R1165_U457 , P1_U3169 );
nand NAND2_10827 ( P1_R1165_U582 , P1_R1165_U76 , P1_R1165_U39 );
nand NAND2_10828 ( P1_R1165_U583 , P1_R1165_U582 , P1_R1165_U581 );
nand NAND2_10829 ( P1_R1165_U584 , P1_R1165_U348 , P1_R1165_U56 );
nand NAND2_10830 ( P1_R1165_U585 , P1_R1165_U583 , P1_R1165_U333 );
nand NAND2_10831 ( P1_R1165_U586 , P1_R1165_U460 , P1_U3170 );
nand NAND2_10832 ( P1_R1165_U587 , P1_R1165_U74 , P1_R1165_U40 );
nand NAND2_10833 ( P1_R1165_U588 , P1_R1165_U587 , P1_R1165_U586 );
nand NAND2_10834 ( P1_R1165_U589 , P1_R1165_U349 , P1_R1165_U190 );
nand NAND2_10835 ( P1_R1165_U590 , P1_R1165_U251 , P1_R1165_U588 );
nand NAND2_10836 ( P1_R1165_U591 , P1_R1165_U451 , P1_U3171 );
nand NAND2_10837 ( P1_R1165_U592 , P1_R1165_U73 , P1_R1165_U38 );
nand NAND2_10838 ( P1_R1165_U593 , P1_R1165_U451 , P1_U3171 );
nand NAND2_10839 ( P1_R1165_U594 , P1_R1165_U73 , P1_R1165_U38 );
nand NAND2_10840 ( P1_R1165_U595 , P1_R1165_U594 , P1_R1165_U593 );
nand NAND2_10841 ( P1_R1165_U596 , P1_R1165_U191 , P1_R1165_U192 );
nand NAND2_10842 ( P1_R1165_U597 , P1_R1165_U364 , P1_R1165_U595 );
nand NAND2_10843 ( P1_R1165_U598 , P1_U3181 , P1_R1165_U16 );
nand NAND2_10844 ( P1_R1165_U599 , P1_U3211 , P1_R1165_U24 );
not NOT1_10845 ( P1_R1165_U600 , P1_R1165_U135 );
nand NAND2_10846 ( P1_R1165_U601 , P1_R1165_U63 , P1_R1165_U600 );
nand NAND2_10847 ( P1_R1165_U602 , P1_R1165_U135 , P1_R1165_U378 );
and AND2_10848 ( P1_R1150_U6 , P1_R1150_U198 , P1_R1150_U197 );
and AND2_10849 ( P1_R1150_U7 , P1_R1150_U237 , P1_R1150_U236 );
and AND2_10850 ( P1_R1150_U8 , P1_R1150_U254 , P1_R1150_U253 );
and AND2_10851 ( P1_R1150_U9 , P1_R1150_U280 , P1_R1150_U279 );
nand NAND2_10852 ( P1_R1150_U10 , P1_R1150_U340 , P1_R1150_U343 );
nand NAND2_10853 ( P1_R1150_U11 , P1_R1150_U329 , P1_R1150_U332 );
nand NAND2_10854 ( P1_R1150_U12 , P1_R1150_U318 , P1_R1150_U321 );
nand NAND2_10855 ( P1_R1150_U13 , P1_R1150_U310 , P1_R1150_U312 );
nand NAND2_10856 ( P1_R1150_U14 , P1_R1150_U347 , P1_R1150_U308 );
nand NAND2_10857 ( P1_R1150_U15 , P1_R1150_U231 , P1_R1150_U233 );
nand NAND2_10858 ( P1_R1150_U16 , P1_R1150_U223 , P1_R1150_U226 );
nand NAND2_10859 ( P1_R1150_U17 , P1_R1150_U215 , P1_R1150_U217 );
nand NAND2_10860 ( P1_R1150_U18 , P1_R1150_U23 , P1_R1150_U346 );
not NOT1_10861 ( P1_R1150_U19 , P1_U3473 );
not NOT1_10862 ( P1_R1150_U20 , P1_U3467 );
not NOT1_10863 ( P1_R1150_U21 , P1_U3458 );
not NOT1_10864 ( P1_R1150_U22 , P1_U3450 );
nand NAND2_10865 ( P1_R1150_U23 , P1_U3450 , P1_R1150_U91 );
not NOT1_10866 ( P1_R1150_U24 , P1_U3078 );
not NOT1_10867 ( P1_R1150_U25 , P1_U3461 );
not NOT1_10868 ( P1_R1150_U26 , P1_U3068 );
nand NAND2_10869 ( P1_R1150_U27 , P1_U3068 , P1_R1150_U21 );
not NOT1_10870 ( P1_R1150_U28 , P1_U3064 );
not NOT1_10871 ( P1_R1150_U29 , P1_U3470 );
not NOT1_10872 ( P1_R1150_U30 , P1_U3464 );
not NOT1_10873 ( P1_R1150_U31 , P1_U3071 );
not NOT1_10874 ( P1_R1150_U32 , P1_U3067 );
not NOT1_10875 ( P1_R1150_U33 , P1_U3060 );
nand NAND2_10876 ( P1_R1150_U34 , P1_U3060 , P1_R1150_U30 );
not NOT1_10877 ( P1_R1150_U35 , P1_U3476 );
not NOT1_10878 ( P1_R1150_U36 , P1_U3070 );
nand NAND2_10879 ( P1_R1150_U37 , P1_U3070 , P1_R1150_U19 );
not NOT1_10880 ( P1_R1150_U38 , P1_U3084 );
not NOT1_10881 ( P1_R1150_U39 , P1_U3479 );
not NOT1_10882 ( P1_R1150_U40 , P1_U3083 );
nand NAND2_10883 ( P1_R1150_U41 , P1_R1150_U204 , P1_R1150_U203 );
nand NAND2_10884 ( P1_R1150_U42 , P1_R1150_U34 , P1_R1150_U219 );
nand NAND2_10885 ( P1_R1150_U43 , P1_R1150_U188 , P1_R1150_U187 );
not NOT1_10886 ( P1_R1150_U44 , P1_U3976 );
not NOT1_10887 ( P1_R1150_U45 , P1_U3980 );
not NOT1_10888 ( P1_R1150_U46 , P1_U3497 );
not NOT1_10889 ( P1_R1150_U47 , P1_U3482 );
not NOT1_10890 ( P1_R1150_U48 , P1_U3485 );
not NOT1_10891 ( P1_R1150_U49 , P1_U3063 );
not NOT1_10892 ( P1_R1150_U50 , P1_U3062 );
nand NAND2_10893 ( P1_R1150_U51 , P1_U3083 , P1_R1150_U39 );
not NOT1_10894 ( P1_R1150_U52 , P1_U3488 );
not NOT1_10895 ( P1_R1150_U53 , P1_U3072 );
not NOT1_10896 ( P1_R1150_U54 , P1_U3491 );
not NOT1_10897 ( P1_R1150_U55 , P1_U3080 );
not NOT1_10898 ( P1_R1150_U56 , P1_U3500 );
not NOT1_10899 ( P1_R1150_U57 , P1_U3494 );
not NOT1_10900 ( P1_R1150_U58 , P1_U3073 );
not NOT1_10901 ( P1_R1150_U59 , P1_U3074 );
not NOT1_10902 ( P1_R1150_U60 , P1_U3079 );
nand NAND2_10903 ( P1_R1150_U61 , P1_U3079 , P1_R1150_U57 );
not NOT1_10904 ( P1_R1150_U62 , P1_U3503 );
not NOT1_10905 ( P1_R1150_U63 , P1_U3069 );
nand NAND2_10906 ( P1_R1150_U64 , P1_R1150_U264 , P1_R1150_U263 );
not NOT1_10907 ( P1_R1150_U65 , P1_U3082 );
not NOT1_10908 ( P1_R1150_U66 , P1_U3508 );
not NOT1_10909 ( P1_R1150_U67 , P1_U3081 );
not NOT1_10910 ( P1_R1150_U68 , P1_U3982 );
not NOT1_10911 ( P1_R1150_U69 , P1_U3076 );
not NOT1_10912 ( P1_R1150_U70 , P1_U3979 );
not NOT1_10913 ( P1_R1150_U71 , P1_U3981 );
not NOT1_10914 ( P1_R1150_U72 , P1_U3066 );
not NOT1_10915 ( P1_R1150_U73 , P1_U3061 );
not NOT1_10916 ( P1_R1150_U74 , P1_U3075 );
nand NAND2_10917 ( P1_R1150_U75 , P1_U3075 , P1_R1150_U71 );
not NOT1_10918 ( P1_R1150_U76 , P1_U3978 );
not NOT1_10919 ( P1_R1150_U77 , P1_U3065 );
not NOT1_10920 ( P1_R1150_U78 , P1_U3977 );
not NOT1_10921 ( P1_R1150_U79 , P1_U3058 );
not NOT1_10922 ( P1_R1150_U80 , P1_U3975 );
not NOT1_10923 ( P1_R1150_U81 , P1_U3057 );
nand NAND2_10924 ( P1_R1150_U82 , P1_U3057 , P1_R1150_U44 );
not NOT1_10925 ( P1_R1150_U83 , P1_U3053 );
not NOT1_10926 ( P1_R1150_U84 , P1_U3974 );
not NOT1_10927 ( P1_R1150_U85 , P1_U3054 );
nand NAND2_10928 ( P1_R1150_U86 , P1_R1150_U126 , P1_R1150_U297 );
nand NAND2_10929 ( P1_R1150_U87 , P1_R1150_U294 , P1_R1150_U293 );
nand NAND2_10930 ( P1_R1150_U88 , P1_R1150_U75 , P1_R1150_U314 );
nand NAND2_10931 ( P1_R1150_U89 , P1_R1150_U61 , P1_R1150_U325 );
nand NAND2_10932 ( P1_R1150_U90 , P1_R1150_U51 , P1_R1150_U336 );
not NOT1_10933 ( P1_R1150_U91 , P1_U3077 );
nand NAND2_10934 ( P1_R1150_U92 , P1_R1150_U390 , P1_R1150_U389 );
nand NAND2_10935 ( P1_R1150_U93 , P1_R1150_U404 , P1_R1150_U403 );
nand NAND2_10936 ( P1_R1150_U94 , P1_R1150_U409 , P1_R1150_U408 );
nand NAND2_10937 ( P1_R1150_U95 , P1_R1150_U425 , P1_R1150_U424 );
nand NAND2_10938 ( P1_R1150_U96 , P1_R1150_U430 , P1_R1150_U429 );
nand NAND2_10939 ( P1_R1150_U97 , P1_R1150_U435 , P1_R1150_U434 );
nand NAND2_10940 ( P1_R1150_U98 , P1_R1150_U440 , P1_R1150_U439 );
nand NAND2_10941 ( P1_R1150_U99 , P1_R1150_U445 , P1_R1150_U444 );
nand NAND2_10942 ( P1_R1150_U100 , P1_R1150_U461 , P1_R1150_U460 );
nand NAND2_10943 ( P1_R1150_U101 , P1_R1150_U466 , P1_R1150_U465 );
nand NAND2_10944 ( P1_R1150_U102 , P1_R1150_U351 , P1_R1150_U350 );
nand NAND2_10945 ( P1_R1150_U103 , P1_R1150_U360 , P1_R1150_U359 );
nand NAND2_10946 ( P1_R1150_U104 , P1_R1150_U367 , P1_R1150_U366 );
nand NAND2_10947 ( P1_R1150_U105 , P1_R1150_U371 , P1_R1150_U370 );
nand NAND2_10948 ( P1_R1150_U106 , P1_R1150_U380 , P1_R1150_U379 );
nand NAND2_10949 ( P1_R1150_U107 , P1_R1150_U399 , P1_R1150_U398 );
nand NAND2_10950 ( P1_R1150_U108 , P1_R1150_U416 , P1_R1150_U415 );
nand NAND2_10951 ( P1_R1150_U109 , P1_R1150_U420 , P1_R1150_U419 );
nand NAND2_10952 ( P1_R1150_U110 , P1_R1150_U452 , P1_R1150_U451 );
nand NAND2_10953 ( P1_R1150_U111 , P1_R1150_U456 , P1_R1150_U455 );
nand NAND2_10954 ( P1_R1150_U112 , P1_R1150_U473 , P1_R1150_U472 );
and AND2_10955 ( P1_R1150_U113 , P1_R1150_U193 , P1_R1150_U194 );
and AND2_10956 ( P1_R1150_U114 , P1_R1150_U201 , P1_R1150_U196 );
and AND2_10957 ( P1_R1150_U115 , P1_R1150_U206 , P1_R1150_U180 );
and AND2_10958 ( P1_R1150_U116 , P1_R1150_U209 , P1_R1150_U210 );
and AND3_10959 ( P1_R1150_U117 , P1_R1150_U353 , P1_R1150_U352 , P1_R1150_U37 );
and AND2_10960 ( P1_R1150_U118 , P1_R1150_U356 , P1_R1150_U180 );
and AND2_10961 ( P1_R1150_U119 , P1_R1150_U225 , P1_R1150_U6 );
and AND2_10962 ( P1_R1150_U120 , P1_R1150_U363 , P1_R1150_U179 );
and AND3_10963 ( P1_R1150_U121 , P1_R1150_U373 , P1_R1150_U372 , P1_R1150_U27 );
and AND2_10964 ( P1_R1150_U122 , P1_R1150_U376 , P1_R1150_U178 );
and AND3_10965 ( P1_R1150_U123 , P1_R1150_U235 , P1_R1150_U212 , P1_R1150_U174 );
and AND3_10966 ( P1_R1150_U124 , P1_R1150_U257 , P1_R1150_U175 , P1_R1150_U252 );
and AND2_10967 ( P1_R1150_U125 , P1_R1150_U283 , P1_R1150_U176 );
and AND2_10968 ( P1_R1150_U126 , P1_R1150_U299 , P1_R1150_U300 );
nand NAND2_10969 ( P1_R1150_U127 , P1_R1150_U387 , P1_R1150_U386 );
and AND3_10970 ( P1_R1150_U128 , P1_R1150_U392 , P1_R1150_U391 , P1_R1150_U82 );
and AND2_10971 ( P1_R1150_U129 , P1_R1150_U395 , P1_R1150_U177 );
nand NAND2_10972 ( P1_R1150_U130 , P1_R1150_U401 , P1_R1150_U400 );
nand NAND2_10973 ( P1_R1150_U131 , P1_R1150_U406 , P1_R1150_U405 );
and AND2_10974 ( P1_R1150_U132 , P1_R1150_U412 , P1_R1150_U176 );
nand NAND2_10975 ( P1_R1150_U133 , P1_R1150_U422 , P1_R1150_U421 );
nand NAND2_10976 ( P1_R1150_U134 , P1_R1150_U427 , P1_R1150_U426 );
nand NAND2_10977 ( P1_R1150_U135 , P1_R1150_U432 , P1_R1150_U431 );
nand NAND2_10978 ( P1_R1150_U136 , P1_R1150_U437 , P1_R1150_U436 );
nand NAND2_10979 ( P1_R1150_U137 , P1_R1150_U442 , P1_R1150_U441 );
and AND2_10980 ( P1_R1150_U138 , P1_R1150_U331 , P1_R1150_U8 );
and AND2_10981 ( P1_R1150_U139 , P1_R1150_U448 , P1_R1150_U175 );
nand NAND2_10982 ( P1_R1150_U140 , P1_R1150_U458 , P1_R1150_U457 );
nand NAND2_10983 ( P1_R1150_U141 , P1_R1150_U463 , P1_R1150_U462 );
and AND2_10984 ( P1_R1150_U142 , P1_R1150_U342 , P1_R1150_U7 );
and AND2_10985 ( P1_R1150_U143 , P1_R1150_U469 , P1_R1150_U174 );
and AND2_10986 ( P1_R1150_U144 , P1_R1150_U349 , P1_R1150_U348 );
nand NAND2_10987 ( P1_R1150_U145 , P1_R1150_U116 , P1_R1150_U207 );
and AND2_10988 ( P1_R1150_U146 , P1_R1150_U358 , P1_R1150_U357 );
and AND2_10989 ( P1_R1150_U147 , P1_R1150_U365 , P1_R1150_U364 );
and AND2_10990 ( P1_R1150_U148 , P1_R1150_U369 , P1_R1150_U368 );
nand NAND2_10991 ( P1_R1150_U149 , P1_R1150_U113 , P1_R1150_U191 );
and AND2_10992 ( P1_R1150_U150 , P1_R1150_U378 , P1_R1150_U377 );
not NOT1_10993 ( P1_R1150_U151 , P1_U3985 );
not NOT1_10994 ( P1_R1150_U152 , P1_U3055 );
and AND2_10995 ( P1_R1150_U153 , P1_R1150_U382 , P1_R1150_U381 );
and AND2_10996 ( P1_R1150_U154 , P1_R1150_U397 , P1_R1150_U396 );
nand NAND2_10997 ( P1_R1150_U155 , P1_R1150_U290 , P1_R1150_U289 );
nand NAND2_10998 ( P1_R1150_U156 , P1_R1150_U286 , P1_R1150_U285 );
and AND2_10999 ( P1_R1150_U157 , P1_R1150_U414 , P1_R1150_U413 );
and AND2_11000 ( P1_R1150_U158 , P1_R1150_U418 , P1_R1150_U417 );
nand NAND2_11001 ( P1_R1150_U159 , P1_R1150_U276 , P1_R1150_U275 );
nand NAND2_11002 ( P1_R1150_U160 , P1_R1150_U272 , P1_R1150_U271 );
not NOT1_11003 ( P1_R1150_U161 , P1_U3455 );
nand NAND2_11004 ( P1_R1150_U162 , P1_R1150_U268 , P1_R1150_U267 );
not NOT1_11005 ( P1_R1150_U163 , P1_U3506 );
nand NAND2_11006 ( P1_R1150_U164 , P1_R1150_U260 , P1_R1150_U259 );
and AND2_11007 ( P1_R1150_U165 , P1_R1150_U450 , P1_R1150_U449 );
and AND2_11008 ( P1_R1150_U166 , P1_R1150_U454 , P1_R1150_U453 );
nand NAND2_11009 ( P1_R1150_U167 , P1_R1150_U250 , P1_R1150_U249 );
nand NAND2_11010 ( P1_R1150_U168 , P1_R1150_U246 , P1_R1150_U245 );
nand NAND2_11011 ( P1_R1150_U169 , P1_R1150_U242 , P1_R1150_U241 );
and AND2_11012 ( P1_R1150_U170 , P1_R1150_U471 , P1_R1150_U470 );
not NOT1_11013 ( P1_R1150_U171 , P1_R1150_U82 );
not NOT1_11014 ( P1_R1150_U172 , P1_R1150_U27 );
not NOT1_11015 ( P1_R1150_U173 , P1_R1150_U37 );
nand NAND2_11016 ( P1_R1150_U174 , P1_U3482 , P1_R1150_U50 );
nand NAND2_11017 ( P1_R1150_U175 , P1_U3497 , P1_R1150_U59 );
nand NAND2_11018 ( P1_R1150_U176 , P1_U3980 , P1_R1150_U73 );
nand NAND2_11019 ( P1_R1150_U177 , P1_U3976 , P1_R1150_U81 );
nand NAND2_11020 ( P1_R1150_U178 , P1_U3458 , P1_R1150_U26 );
nand NAND2_11021 ( P1_R1150_U179 , P1_U3467 , P1_R1150_U32 );
nand NAND2_11022 ( P1_R1150_U180 , P1_U3473 , P1_R1150_U36 );
not NOT1_11023 ( P1_R1150_U181 , P1_R1150_U61 );
not NOT1_11024 ( P1_R1150_U182 , P1_R1150_U75 );
not NOT1_11025 ( P1_R1150_U183 , P1_R1150_U34 );
not NOT1_11026 ( P1_R1150_U184 , P1_R1150_U51 );
not NOT1_11027 ( P1_R1150_U185 , P1_R1150_U23 );
nand NAND2_11028 ( P1_R1150_U186 , P1_R1150_U185 , P1_R1150_U24 );
nand NAND2_11029 ( P1_R1150_U187 , P1_R1150_U186 , P1_R1150_U161 );
nand NAND2_11030 ( P1_R1150_U188 , P1_U3078 , P1_R1150_U23 );
not NOT1_11031 ( P1_R1150_U189 , P1_R1150_U43 );
nand NAND2_11032 ( P1_R1150_U190 , P1_U3461 , P1_R1150_U28 );
nand NAND3_11033 ( P1_R1150_U191 , P1_R1150_U43 , P1_R1150_U178 , P1_R1150_U190 );
nand NAND2_11034 ( P1_R1150_U192 , P1_R1150_U28 , P1_R1150_U27 );
nand NAND2_11035 ( P1_R1150_U193 , P1_R1150_U192 , P1_R1150_U25 );
nand NAND2_11036 ( P1_R1150_U194 , P1_U3064 , P1_R1150_U172 );
not NOT1_11037 ( P1_R1150_U195 , P1_R1150_U149 );
nand NAND2_11038 ( P1_R1150_U196 , P1_U3470 , P1_R1150_U31 );
nand NAND2_11039 ( P1_R1150_U197 , P1_U3071 , P1_R1150_U29 );
nand NAND2_11040 ( P1_R1150_U198 , P1_U3067 , P1_R1150_U20 );
nand NAND2_11041 ( P1_R1150_U199 , P1_R1150_U183 , P1_R1150_U179 );
nand NAND2_11042 ( P1_R1150_U200 , P1_R1150_U6 , P1_R1150_U199 );
nand NAND2_11043 ( P1_R1150_U201 , P1_U3464 , P1_R1150_U33 );
nand NAND2_11044 ( P1_R1150_U202 , P1_U3470 , P1_R1150_U31 );
nand NAND3_11045 ( P1_R1150_U203 , P1_R1150_U149 , P1_R1150_U179 , P1_R1150_U114 );
nand NAND2_11046 ( P1_R1150_U204 , P1_R1150_U202 , P1_R1150_U200 );
not NOT1_11047 ( P1_R1150_U205 , P1_R1150_U41 );
nand NAND2_11048 ( P1_R1150_U206 , P1_U3476 , P1_R1150_U38 );
nand NAND2_11049 ( P1_R1150_U207 , P1_R1150_U115 , P1_R1150_U41 );
nand NAND2_11050 ( P1_R1150_U208 , P1_R1150_U38 , P1_R1150_U37 );
nand NAND2_11051 ( P1_R1150_U209 , P1_R1150_U208 , P1_R1150_U35 );
nand NAND2_11052 ( P1_R1150_U210 , P1_U3084 , P1_R1150_U173 );
not NOT1_11053 ( P1_R1150_U211 , P1_R1150_U145 );
nand NAND2_11054 ( P1_R1150_U212 , P1_U3479 , P1_R1150_U40 );
nand NAND2_11055 ( P1_R1150_U213 , P1_R1150_U212 , P1_R1150_U51 );
nand NAND2_11056 ( P1_R1150_U214 , P1_R1150_U205 , P1_R1150_U37 );
nand NAND2_11057 ( P1_R1150_U215 , P1_R1150_U118 , P1_R1150_U214 );
nand NAND2_11058 ( P1_R1150_U216 , P1_R1150_U41 , P1_R1150_U180 );
nand NAND2_11059 ( P1_R1150_U217 , P1_R1150_U117 , P1_R1150_U216 );
nand NAND2_11060 ( P1_R1150_U218 , P1_R1150_U37 , P1_R1150_U180 );
nand NAND2_11061 ( P1_R1150_U219 , P1_R1150_U201 , P1_R1150_U149 );
not NOT1_11062 ( P1_R1150_U220 , P1_R1150_U42 );
nand NAND2_11063 ( P1_R1150_U221 , P1_U3067 , P1_R1150_U20 );
nand NAND2_11064 ( P1_R1150_U222 , P1_R1150_U220 , P1_R1150_U221 );
nand NAND2_11065 ( P1_R1150_U223 , P1_R1150_U120 , P1_R1150_U222 );
nand NAND2_11066 ( P1_R1150_U224 , P1_R1150_U42 , P1_R1150_U179 );
nand NAND2_11067 ( P1_R1150_U225 , P1_U3470 , P1_R1150_U31 );
nand NAND2_11068 ( P1_R1150_U226 , P1_R1150_U119 , P1_R1150_U224 );
nand NAND2_11069 ( P1_R1150_U227 , P1_U3067 , P1_R1150_U20 );
nand NAND2_11070 ( P1_R1150_U228 , P1_R1150_U179 , P1_R1150_U227 );
nand NAND2_11071 ( P1_R1150_U229 , P1_R1150_U201 , P1_R1150_U34 );
nand NAND2_11072 ( P1_R1150_U230 , P1_R1150_U189 , P1_R1150_U27 );
nand NAND2_11073 ( P1_R1150_U231 , P1_R1150_U122 , P1_R1150_U230 );
nand NAND2_11074 ( P1_R1150_U232 , P1_R1150_U43 , P1_R1150_U178 );
nand NAND2_11075 ( P1_R1150_U233 , P1_R1150_U121 , P1_R1150_U232 );
nand NAND2_11076 ( P1_R1150_U234 , P1_R1150_U27 , P1_R1150_U178 );
nand NAND2_11077 ( P1_R1150_U235 , P1_U3485 , P1_R1150_U49 );
nand NAND2_11078 ( P1_R1150_U236 , P1_U3063 , P1_R1150_U48 );
nand NAND2_11079 ( P1_R1150_U237 , P1_U3062 , P1_R1150_U47 );
nand NAND2_11080 ( P1_R1150_U238 , P1_R1150_U184 , P1_R1150_U174 );
nand NAND2_11081 ( P1_R1150_U239 , P1_R1150_U7 , P1_R1150_U238 );
nand NAND2_11082 ( P1_R1150_U240 , P1_U3485 , P1_R1150_U49 );
nand NAND2_11083 ( P1_R1150_U241 , P1_R1150_U145 , P1_R1150_U123 );
nand NAND2_11084 ( P1_R1150_U242 , P1_R1150_U240 , P1_R1150_U239 );
not NOT1_11085 ( P1_R1150_U243 , P1_R1150_U169 );
nand NAND2_11086 ( P1_R1150_U244 , P1_U3488 , P1_R1150_U53 );
nand NAND2_11087 ( P1_R1150_U245 , P1_R1150_U244 , P1_R1150_U169 );
nand NAND2_11088 ( P1_R1150_U246 , P1_U3072 , P1_R1150_U52 );
not NOT1_11089 ( P1_R1150_U247 , P1_R1150_U168 );
nand NAND2_11090 ( P1_R1150_U248 , P1_U3491 , P1_R1150_U55 );
nand NAND2_11091 ( P1_R1150_U249 , P1_R1150_U248 , P1_R1150_U168 );
nand NAND2_11092 ( P1_R1150_U250 , P1_U3080 , P1_R1150_U54 );
not NOT1_11093 ( P1_R1150_U251 , P1_R1150_U167 );
nand NAND2_11094 ( P1_R1150_U252 , P1_U3500 , P1_R1150_U58 );
nand NAND2_11095 ( P1_R1150_U253 , P1_U3073 , P1_R1150_U56 );
nand NAND2_11096 ( P1_R1150_U254 , P1_U3074 , P1_R1150_U46 );
nand NAND2_11097 ( P1_R1150_U255 , P1_R1150_U181 , P1_R1150_U175 );
nand NAND2_11098 ( P1_R1150_U256 , P1_R1150_U8 , P1_R1150_U255 );
nand NAND2_11099 ( P1_R1150_U257 , P1_U3494 , P1_R1150_U60 );
nand NAND2_11100 ( P1_R1150_U258 , P1_U3500 , P1_R1150_U58 );
nand NAND2_11101 ( P1_R1150_U259 , P1_R1150_U167 , P1_R1150_U124 );
nand NAND2_11102 ( P1_R1150_U260 , P1_R1150_U258 , P1_R1150_U256 );
not NOT1_11103 ( P1_R1150_U261 , P1_R1150_U164 );
nand NAND2_11104 ( P1_R1150_U262 , P1_U3503 , P1_R1150_U63 );
nand NAND2_11105 ( P1_R1150_U263 , P1_R1150_U262 , P1_R1150_U164 );
nand NAND2_11106 ( P1_R1150_U264 , P1_U3069 , P1_R1150_U62 );
not NOT1_11107 ( P1_R1150_U265 , P1_R1150_U64 );
nand NAND2_11108 ( P1_R1150_U266 , P1_R1150_U265 , P1_R1150_U65 );
nand NAND2_11109 ( P1_R1150_U267 , P1_R1150_U266 , P1_R1150_U163 );
nand NAND2_11110 ( P1_R1150_U268 , P1_U3082 , P1_R1150_U64 );
not NOT1_11111 ( P1_R1150_U269 , P1_R1150_U162 );
nand NAND2_11112 ( P1_R1150_U270 , P1_U3508 , P1_R1150_U67 );
nand NAND2_11113 ( P1_R1150_U271 , P1_R1150_U270 , P1_R1150_U162 );
nand NAND2_11114 ( P1_R1150_U272 , P1_U3081 , P1_R1150_U66 );
not NOT1_11115 ( P1_R1150_U273 , P1_R1150_U160 );
nand NAND2_11116 ( P1_R1150_U274 , P1_U3982 , P1_R1150_U69 );
nand NAND2_11117 ( P1_R1150_U275 , P1_R1150_U274 , P1_R1150_U160 );
nand NAND2_11118 ( P1_R1150_U276 , P1_U3076 , P1_R1150_U68 );
not NOT1_11119 ( P1_R1150_U277 , P1_R1150_U159 );
nand NAND2_11120 ( P1_R1150_U278 , P1_U3979 , P1_R1150_U72 );
nand NAND2_11121 ( P1_R1150_U279 , P1_U3066 , P1_R1150_U70 );
nand NAND2_11122 ( P1_R1150_U280 , P1_U3061 , P1_R1150_U45 );
nand NAND2_11123 ( P1_R1150_U281 , P1_R1150_U182 , P1_R1150_U176 );
nand NAND2_11124 ( P1_R1150_U282 , P1_R1150_U9 , P1_R1150_U281 );
nand NAND2_11125 ( P1_R1150_U283 , P1_U3981 , P1_R1150_U74 );
nand NAND2_11126 ( P1_R1150_U284 , P1_U3979 , P1_R1150_U72 );
nand NAND3_11127 ( P1_R1150_U285 , P1_R1150_U159 , P1_R1150_U125 , P1_R1150_U278 );
nand NAND2_11128 ( P1_R1150_U286 , P1_R1150_U284 , P1_R1150_U282 );
not NOT1_11129 ( P1_R1150_U287 , P1_R1150_U156 );
nand NAND2_11130 ( P1_R1150_U288 , P1_U3978 , P1_R1150_U77 );
nand NAND2_11131 ( P1_R1150_U289 , P1_R1150_U288 , P1_R1150_U156 );
nand NAND2_11132 ( P1_R1150_U290 , P1_U3065 , P1_R1150_U76 );
not NOT1_11133 ( P1_R1150_U291 , P1_R1150_U155 );
nand NAND2_11134 ( P1_R1150_U292 , P1_U3977 , P1_R1150_U79 );
nand NAND2_11135 ( P1_R1150_U293 , P1_R1150_U292 , P1_R1150_U155 );
nand NAND2_11136 ( P1_R1150_U294 , P1_U3058 , P1_R1150_U78 );
not NOT1_11137 ( P1_R1150_U295 , P1_R1150_U87 );
nand NAND2_11138 ( P1_R1150_U296 , P1_U3975 , P1_R1150_U83 );
nand NAND3_11139 ( P1_R1150_U297 , P1_R1150_U87 , P1_R1150_U177 , P1_R1150_U296 );
nand NAND2_11140 ( P1_R1150_U298 , P1_R1150_U83 , P1_R1150_U82 );
nand NAND2_11141 ( P1_R1150_U299 , P1_R1150_U298 , P1_R1150_U80 );
nand NAND2_11142 ( P1_R1150_U300 , P1_U3053 , P1_R1150_U171 );
not NOT1_11143 ( P1_R1150_U301 , P1_R1150_U86 );
nand NAND2_11144 ( P1_R1150_U302 , P1_U3054 , P1_R1150_U84 );
nand NAND2_11145 ( P1_R1150_U303 , P1_R1150_U301 , P1_R1150_U302 );
nand NAND2_11146 ( P1_R1150_U304 , P1_U3974 , P1_R1150_U85 );
nand NAND2_11147 ( P1_R1150_U305 , P1_U3974 , P1_R1150_U85 );
nand NAND2_11148 ( P1_R1150_U306 , P1_R1150_U305 , P1_R1150_U86 );
nand NAND2_11149 ( P1_R1150_U307 , P1_U3054 , P1_R1150_U84 );
nand NAND3_11150 ( P1_R1150_U308 , P1_R1150_U307 , P1_R1150_U306 , P1_R1150_U153 );
nand NAND2_11151 ( P1_R1150_U309 , P1_R1150_U295 , P1_R1150_U82 );
nand NAND2_11152 ( P1_R1150_U310 , P1_R1150_U129 , P1_R1150_U309 );
nand NAND2_11153 ( P1_R1150_U311 , P1_R1150_U87 , P1_R1150_U177 );
nand NAND2_11154 ( P1_R1150_U312 , P1_R1150_U128 , P1_R1150_U311 );
nand NAND2_11155 ( P1_R1150_U313 , P1_R1150_U82 , P1_R1150_U177 );
nand NAND2_11156 ( P1_R1150_U314 , P1_R1150_U283 , P1_R1150_U159 );
not NOT1_11157 ( P1_R1150_U315 , P1_R1150_U88 );
nand NAND2_11158 ( P1_R1150_U316 , P1_U3061 , P1_R1150_U45 );
nand NAND2_11159 ( P1_R1150_U317 , P1_R1150_U315 , P1_R1150_U316 );
nand NAND2_11160 ( P1_R1150_U318 , P1_R1150_U132 , P1_R1150_U317 );
nand NAND2_11161 ( P1_R1150_U319 , P1_R1150_U88 , P1_R1150_U176 );
nand NAND2_11162 ( P1_R1150_U320 , P1_U3979 , P1_R1150_U72 );
nand NAND3_11163 ( P1_R1150_U321 , P1_R1150_U320 , P1_R1150_U319 , P1_R1150_U9 );
nand NAND2_11164 ( P1_R1150_U322 , P1_U3061 , P1_R1150_U45 );
nand NAND2_11165 ( P1_R1150_U323 , P1_R1150_U176 , P1_R1150_U322 );
nand NAND2_11166 ( P1_R1150_U324 , P1_R1150_U283 , P1_R1150_U75 );
nand NAND2_11167 ( P1_R1150_U325 , P1_R1150_U257 , P1_R1150_U167 );
not NOT1_11168 ( P1_R1150_U326 , P1_R1150_U89 );
nand NAND2_11169 ( P1_R1150_U327 , P1_U3074 , P1_R1150_U46 );
nand NAND2_11170 ( P1_R1150_U328 , P1_R1150_U326 , P1_R1150_U327 );
nand NAND2_11171 ( P1_R1150_U329 , P1_R1150_U139 , P1_R1150_U328 );
nand NAND2_11172 ( P1_R1150_U330 , P1_R1150_U89 , P1_R1150_U175 );
nand NAND2_11173 ( P1_R1150_U331 , P1_U3500 , P1_R1150_U58 );
nand NAND2_11174 ( P1_R1150_U332 , P1_R1150_U138 , P1_R1150_U330 );
nand NAND2_11175 ( P1_R1150_U333 , P1_U3074 , P1_R1150_U46 );
nand NAND2_11176 ( P1_R1150_U334 , P1_R1150_U175 , P1_R1150_U333 );
nand NAND2_11177 ( P1_R1150_U335 , P1_R1150_U257 , P1_R1150_U61 );
nand NAND2_11178 ( P1_R1150_U336 , P1_R1150_U212 , P1_R1150_U145 );
not NOT1_11179 ( P1_R1150_U337 , P1_R1150_U90 );
nand NAND2_11180 ( P1_R1150_U338 , P1_U3062 , P1_R1150_U47 );
nand NAND2_11181 ( P1_R1150_U339 , P1_R1150_U337 , P1_R1150_U338 );
nand NAND2_11182 ( P1_R1150_U340 , P1_R1150_U143 , P1_R1150_U339 );
nand NAND2_11183 ( P1_R1150_U341 , P1_R1150_U90 , P1_R1150_U174 );
nand NAND2_11184 ( P1_R1150_U342 , P1_U3485 , P1_R1150_U49 );
nand NAND2_11185 ( P1_R1150_U343 , P1_R1150_U142 , P1_R1150_U341 );
nand NAND2_11186 ( P1_R1150_U344 , P1_U3062 , P1_R1150_U47 );
nand NAND2_11187 ( P1_R1150_U345 , P1_R1150_U174 , P1_R1150_U344 );
nand NAND2_11188 ( P1_R1150_U346 , P1_U3077 , P1_R1150_U22 );
nand NAND3_11189 ( P1_R1150_U347 , P1_R1150_U304 , P1_R1150_U303 , P1_R1150_U385 );
nand NAND2_11190 ( P1_R1150_U348 , P1_U3479 , P1_R1150_U40 );
nand NAND2_11191 ( P1_R1150_U349 , P1_U3083 , P1_R1150_U39 );
nand NAND2_11192 ( P1_R1150_U350 , P1_R1150_U213 , P1_R1150_U145 );
nand NAND2_11193 ( P1_R1150_U351 , P1_R1150_U211 , P1_R1150_U144 );
nand NAND2_11194 ( P1_R1150_U352 , P1_U3476 , P1_R1150_U38 );
nand NAND2_11195 ( P1_R1150_U353 , P1_U3084 , P1_R1150_U35 );
nand NAND2_11196 ( P1_R1150_U354 , P1_U3476 , P1_R1150_U38 );
nand NAND2_11197 ( P1_R1150_U355 , P1_U3084 , P1_R1150_U35 );
nand NAND2_11198 ( P1_R1150_U356 , P1_R1150_U355 , P1_R1150_U354 );
nand NAND2_11199 ( P1_R1150_U357 , P1_U3473 , P1_R1150_U36 );
nand NAND2_11200 ( P1_R1150_U358 , P1_U3070 , P1_R1150_U19 );
nand NAND2_11201 ( P1_R1150_U359 , P1_R1150_U218 , P1_R1150_U41 );
nand NAND2_11202 ( P1_R1150_U360 , P1_R1150_U146 , P1_R1150_U205 );
nand NAND2_11203 ( P1_R1150_U361 , P1_U3470 , P1_R1150_U31 );
nand NAND2_11204 ( P1_R1150_U362 , P1_U3071 , P1_R1150_U29 );
nand NAND2_11205 ( P1_R1150_U363 , P1_R1150_U362 , P1_R1150_U361 );
nand NAND2_11206 ( P1_R1150_U364 , P1_U3467 , P1_R1150_U32 );
nand NAND2_11207 ( P1_R1150_U365 , P1_U3067 , P1_R1150_U20 );
nand NAND2_11208 ( P1_R1150_U366 , P1_R1150_U228 , P1_R1150_U42 );
nand NAND2_11209 ( P1_R1150_U367 , P1_R1150_U147 , P1_R1150_U220 );
nand NAND2_11210 ( P1_R1150_U368 , P1_U3464 , P1_R1150_U33 );
nand NAND2_11211 ( P1_R1150_U369 , P1_U3060 , P1_R1150_U30 );
nand NAND2_11212 ( P1_R1150_U370 , P1_R1150_U229 , P1_R1150_U149 );
nand NAND2_11213 ( P1_R1150_U371 , P1_R1150_U195 , P1_R1150_U148 );
nand NAND2_11214 ( P1_R1150_U372 , P1_U3461 , P1_R1150_U28 );
nand NAND2_11215 ( P1_R1150_U373 , P1_U3064 , P1_R1150_U25 );
nand NAND2_11216 ( P1_R1150_U374 , P1_U3461 , P1_R1150_U28 );
nand NAND2_11217 ( P1_R1150_U375 , P1_U3064 , P1_R1150_U25 );
nand NAND2_11218 ( P1_R1150_U376 , P1_R1150_U375 , P1_R1150_U374 );
nand NAND2_11219 ( P1_R1150_U377 , P1_U3458 , P1_R1150_U26 );
nand NAND2_11220 ( P1_R1150_U378 , P1_U3068 , P1_R1150_U21 );
nand NAND2_11221 ( P1_R1150_U379 , P1_R1150_U234 , P1_R1150_U43 );
nand NAND2_11222 ( P1_R1150_U380 , P1_R1150_U150 , P1_R1150_U189 );
nand NAND2_11223 ( P1_R1150_U381 , P1_U3985 , P1_R1150_U152 );
nand NAND2_11224 ( P1_R1150_U382 , P1_U3055 , P1_R1150_U151 );
nand NAND2_11225 ( P1_R1150_U383 , P1_U3985 , P1_R1150_U152 );
nand NAND2_11226 ( P1_R1150_U384 , P1_U3055 , P1_R1150_U151 );
nand NAND2_11227 ( P1_R1150_U385 , P1_R1150_U384 , P1_R1150_U383 );
nand NAND2_11228 ( P1_R1150_U386 , P1_U3974 , P1_R1150_U85 );
nand NAND2_11229 ( P1_R1150_U387 , P1_U3054 , P1_R1150_U84 );
not NOT1_11230 ( P1_R1150_U388 , P1_R1150_U127 );
nand NAND2_11231 ( P1_R1150_U389 , P1_R1150_U388 , P1_R1150_U301 );
nand NAND2_11232 ( P1_R1150_U390 , P1_R1150_U127 , P1_R1150_U86 );
nand NAND2_11233 ( P1_R1150_U391 , P1_U3975 , P1_R1150_U83 );
nand NAND2_11234 ( P1_R1150_U392 , P1_U3053 , P1_R1150_U80 );
nand NAND2_11235 ( P1_R1150_U393 , P1_U3975 , P1_R1150_U83 );
nand NAND2_11236 ( P1_R1150_U394 , P1_U3053 , P1_R1150_U80 );
nand NAND2_11237 ( P1_R1150_U395 , P1_R1150_U394 , P1_R1150_U393 );
nand NAND2_11238 ( P1_R1150_U396 , P1_U3976 , P1_R1150_U81 );
nand NAND2_11239 ( P1_R1150_U397 , P1_U3057 , P1_R1150_U44 );
nand NAND2_11240 ( P1_R1150_U398 , P1_R1150_U313 , P1_R1150_U87 );
nand NAND2_11241 ( P1_R1150_U399 , P1_R1150_U154 , P1_R1150_U295 );
nand NAND2_11242 ( P1_R1150_U400 , P1_U3977 , P1_R1150_U79 );
nand NAND2_11243 ( P1_R1150_U401 , P1_U3058 , P1_R1150_U78 );
not NOT1_11244 ( P1_R1150_U402 , P1_R1150_U130 );
nand NAND2_11245 ( P1_R1150_U403 , P1_R1150_U291 , P1_R1150_U402 );
nand NAND2_11246 ( P1_R1150_U404 , P1_R1150_U130 , P1_R1150_U155 );
nand NAND2_11247 ( P1_R1150_U405 , P1_U3978 , P1_R1150_U77 );
nand NAND2_11248 ( P1_R1150_U406 , P1_U3065 , P1_R1150_U76 );
not NOT1_11249 ( P1_R1150_U407 , P1_R1150_U131 );
nand NAND2_11250 ( P1_R1150_U408 , P1_R1150_U287 , P1_R1150_U407 );
nand NAND2_11251 ( P1_R1150_U409 , P1_R1150_U131 , P1_R1150_U156 );
nand NAND2_11252 ( P1_R1150_U410 , P1_U3979 , P1_R1150_U72 );
nand NAND2_11253 ( P1_R1150_U411 , P1_U3066 , P1_R1150_U70 );
nand NAND2_11254 ( P1_R1150_U412 , P1_R1150_U411 , P1_R1150_U410 );
nand NAND2_11255 ( P1_R1150_U413 , P1_U3980 , P1_R1150_U73 );
nand NAND2_11256 ( P1_R1150_U414 , P1_U3061 , P1_R1150_U45 );
nand NAND2_11257 ( P1_R1150_U415 , P1_R1150_U323 , P1_R1150_U88 );
nand NAND2_11258 ( P1_R1150_U416 , P1_R1150_U157 , P1_R1150_U315 );
nand NAND2_11259 ( P1_R1150_U417 , P1_U3981 , P1_R1150_U74 );
nand NAND2_11260 ( P1_R1150_U418 , P1_U3075 , P1_R1150_U71 );
nand NAND2_11261 ( P1_R1150_U419 , P1_R1150_U324 , P1_R1150_U159 );
nand NAND2_11262 ( P1_R1150_U420 , P1_R1150_U277 , P1_R1150_U158 );
nand NAND2_11263 ( P1_R1150_U421 , P1_U3982 , P1_R1150_U69 );
nand NAND2_11264 ( P1_R1150_U422 , P1_U3076 , P1_R1150_U68 );
not NOT1_11265 ( P1_R1150_U423 , P1_R1150_U133 );
nand NAND2_11266 ( P1_R1150_U424 , P1_R1150_U273 , P1_R1150_U423 );
nand NAND2_11267 ( P1_R1150_U425 , P1_R1150_U133 , P1_R1150_U160 );
nand NAND2_11268 ( P1_R1150_U426 , P1_R1150_U185 , P1_R1150_U24 );
nand NAND2_11269 ( P1_R1150_U427 , P1_U3078 , P1_R1150_U23 );
not NOT1_11270 ( P1_R1150_U428 , P1_R1150_U134 );
nand NAND2_11271 ( P1_R1150_U429 , P1_U3455 , P1_R1150_U428 );
nand NAND2_11272 ( P1_R1150_U430 , P1_R1150_U134 , P1_R1150_U161 );
nand NAND2_11273 ( P1_R1150_U431 , P1_U3508 , P1_R1150_U67 );
nand NAND2_11274 ( P1_R1150_U432 , P1_U3081 , P1_R1150_U66 );
not NOT1_11275 ( P1_R1150_U433 , P1_R1150_U135 );
nand NAND2_11276 ( P1_R1150_U434 , P1_R1150_U269 , P1_R1150_U433 );
nand NAND2_11277 ( P1_R1150_U435 , P1_R1150_U135 , P1_R1150_U162 );
nand NAND2_11278 ( P1_R1150_U436 , P1_U3506 , P1_R1150_U65 );
nand NAND2_11279 ( P1_R1150_U437 , P1_U3082 , P1_R1150_U163 );
not NOT1_11280 ( P1_R1150_U438 , P1_R1150_U136 );
nand NAND2_11281 ( P1_R1150_U439 , P1_R1150_U438 , P1_R1150_U265 );
nand NAND2_11282 ( P1_R1150_U440 , P1_R1150_U136 , P1_R1150_U64 );
nand NAND2_11283 ( P1_R1150_U441 , P1_U3503 , P1_R1150_U63 );
nand NAND2_11284 ( P1_R1150_U442 , P1_U3069 , P1_R1150_U62 );
not NOT1_11285 ( P1_R1150_U443 , P1_R1150_U137 );
nand NAND2_11286 ( P1_R1150_U444 , P1_R1150_U261 , P1_R1150_U443 );
nand NAND2_11287 ( P1_R1150_U445 , P1_R1150_U137 , P1_R1150_U164 );
nand NAND2_11288 ( P1_R1150_U446 , P1_U3500 , P1_R1150_U58 );
nand NAND2_11289 ( P1_R1150_U447 , P1_U3073 , P1_R1150_U56 );
nand NAND2_11290 ( P1_R1150_U448 , P1_R1150_U447 , P1_R1150_U446 );
nand NAND2_11291 ( P1_R1150_U449 , P1_U3497 , P1_R1150_U59 );
nand NAND2_11292 ( P1_R1150_U450 , P1_U3074 , P1_R1150_U46 );
nand NAND2_11293 ( P1_R1150_U451 , P1_R1150_U334 , P1_R1150_U89 );
nand NAND2_11294 ( P1_R1150_U452 , P1_R1150_U165 , P1_R1150_U326 );
nand NAND2_11295 ( P1_R1150_U453 , P1_U3494 , P1_R1150_U60 );
nand NAND2_11296 ( P1_R1150_U454 , P1_U3079 , P1_R1150_U57 );
nand NAND2_11297 ( P1_R1150_U455 , P1_R1150_U335 , P1_R1150_U167 );
nand NAND2_11298 ( P1_R1150_U456 , P1_R1150_U251 , P1_R1150_U166 );
nand NAND2_11299 ( P1_R1150_U457 , P1_U3491 , P1_R1150_U55 );
nand NAND2_11300 ( P1_R1150_U458 , P1_U3080 , P1_R1150_U54 );
not NOT1_11301 ( P1_R1150_U459 , P1_R1150_U140 );
nand NAND2_11302 ( P1_R1150_U460 , P1_R1150_U247 , P1_R1150_U459 );
nand NAND2_11303 ( P1_R1150_U461 , P1_R1150_U140 , P1_R1150_U168 );
nand NAND2_11304 ( P1_R1150_U462 , P1_U3488 , P1_R1150_U53 );
nand NAND2_11305 ( P1_R1150_U463 , P1_U3072 , P1_R1150_U52 );
not NOT1_11306 ( P1_R1150_U464 , P1_R1150_U141 );
nand NAND2_11307 ( P1_R1150_U465 , P1_R1150_U243 , P1_R1150_U464 );
nand NAND2_11308 ( P1_R1150_U466 , P1_R1150_U141 , P1_R1150_U169 );
nand NAND2_11309 ( P1_R1150_U467 , P1_U3485 , P1_R1150_U49 );
nand NAND2_11310 ( P1_R1150_U468 , P1_U3063 , P1_R1150_U48 );
nand NAND2_11311 ( P1_R1150_U469 , P1_R1150_U468 , P1_R1150_U467 );
nand NAND2_11312 ( P1_R1150_U470 , P1_U3482 , P1_R1150_U50 );
nand NAND2_11313 ( P1_R1150_U471 , P1_U3062 , P1_R1150_U47 );
nand NAND2_11314 ( P1_R1150_U472 , P1_R1150_U345 , P1_R1150_U90 );
nand NAND2_11315 ( P1_R1150_U473 , P1_R1150_U170 , P1_R1150_U337 );
and AND2_11316 ( P1_R1192_U6 , P1_R1192_U198 , P1_R1192_U197 );
and AND2_11317 ( P1_R1192_U7 , P1_R1192_U237 , P1_R1192_U236 );
and AND2_11318 ( P1_R1192_U8 , P1_R1192_U254 , P1_R1192_U253 );
and AND2_11319 ( P1_R1192_U9 , P1_R1192_U280 , P1_R1192_U279 );
nand NAND2_11320 ( P1_R1192_U10 , P1_R1192_U340 , P1_R1192_U343 );
nand NAND2_11321 ( P1_R1192_U11 , P1_R1192_U329 , P1_R1192_U332 );
nand NAND2_11322 ( P1_R1192_U12 , P1_R1192_U318 , P1_R1192_U321 );
nand NAND2_11323 ( P1_R1192_U13 , P1_R1192_U310 , P1_R1192_U312 );
nand NAND2_11324 ( P1_R1192_U14 , P1_R1192_U347 , P1_R1192_U308 );
nand NAND2_11325 ( P1_R1192_U15 , P1_R1192_U231 , P1_R1192_U233 );
nand NAND2_11326 ( P1_R1192_U16 , P1_R1192_U223 , P1_R1192_U226 );
nand NAND2_11327 ( P1_R1192_U17 , P1_R1192_U215 , P1_R1192_U217 );
nand NAND2_11328 ( P1_R1192_U18 , P1_R1192_U23 , P1_R1192_U346 );
not NOT1_11329 ( P1_R1192_U19 , P1_U3473 );
not NOT1_11330 ( P1_R1192_U20 , P1_U3467 );
not NOT1_11331 ( P1_R1192_U21 , P1_U3458 );
not NOT1_11332 ( P1_R1192_U22 , P1_U3450 );
nand NAND2_11333 ( P1_R1192_U23 , P1_U3450 , P1_R1192_U91 );
not NOT1_11334 ( P1_R1192_U24 , P1_U3078 );
not NOT1_11335 ( P1_R1192_U25 , P1_U3461 );
not NOT1_11336 ( P1_R1192_U26 , P1_U3068 );
nand NAND2_11337 ( P1_R1192_U27 , P1_U3068 , P1_R1192_U21 );
not NOT1_11338 ( P1_R1192_U28 , P1_U3064 );
not NOT1_11339 ( P1_R1192_U29 , P1_U3470 );
not NOT1_11340 ( P1_R1192_U30 , P1_U3464 );
not NOT1_11341 ( P1_R1192_U31 , P1_U3071 );
not NOT1_11342 ( P1_R1192_U32 , P1_U3067 );
not NOT1_11343 ( P1_R1192_U33 , P1_U3060 );
nand NAND2_11344 ( P1_R1192_U34 , P1_U3060 , P1_R1192_U30 );
not NOT1_11345 ( P1_R1192_U35 , P1_U3476 );
not NOT1_11346 ( P1_R1192_U36 , P1_U3070 );
nand NAND2_11347 ( P1_R1192_U37 , P1_U3070 , P1_R1192_U19 );
not NOT1_11348 ( P1_R1192_U38 , P1_U3084 );
not NOT1_11349 ( P1_R1192_U39 , P1_U3479 );
not NOT1_11350 ( P1_R1192_U40 , P1_U3083 );
nand NAND2_11351 ( P1_R1192_U41 , P1_R1192_U204 , P1_R1192_U203 );
nand NAND2_11352 ( P1_R1192_U42 , P1_R1192_U34 , P1_R1192_U219 );
nand NAND2_11353 ( P1_R1192_U43 , P1_R1192_U188 , P1_R1192_U187 );
not NOT1_11354 ( P1_R1192_U44 , P1_U3976 );
not NOT1_11355 ( P1_R1192_U45 , P1_U3980 );
not NOT1_11356 ( P1_R1192_U46 , P1_U3497 );
not NOT1_11357 ( P1_R1192_U47 , P1_U3482 );
not NOT1_11358 ( P1_R1192_U48 , P1_U3485 );
not NOT1_11359 ( P1_R1192_U49 , P1_U3063 );
not NOT1_11360 ( P1_R1192_U50 , P1_U3062 );
nand NAND2_11361 ( P1_R1192_U51 , P1_U3083 , P1_R1192_U39 );
not NOT1_11362 ( P1_R1192_U52 , P1_U3488 );
not NOT1_11363 ( P1_R1192_U53 , P1_U3072 );
not NOT1_11364 ( P1_R1192_U54 , P1_U3491 );
not NOT1_11365 ( P1_R1192_U55 , P1_U3080 );
not NOT1_11366 ( P1_R1192_U56 , P1_U3500 );
not NOT1_11367 ( P1_R1192_U57 , P1_U3494 );
not NOT1_11368 ( P1_R1192_U58 , P1_U3073 );
not NOT1_11369 ( P1_R1192_U59 , P1_U3074 );
not NOT1_11370 ( P1_R1192_U60 , P1_U3079 );
nand NAND2_11371 ( P1_R1192_U61 , P1_U3079 , P1_R1192_U57 );
not NOT1_11372 ( P1_R1192_U62 , P1_U3503 );
not NOT1_11373 ( P1_R1192_U63 , P1_U3069 );
nand NAND2_11374 ( P1_R1192_U64 , P1_R1192_U264 , P1_R1192_U263 );
not NOT1_11375 ( P1_R1192_U65 , P1_U3082 );
not NOT1_11376 ( P1_R1192_U66 , P1_U3508 );
not NOT1_11377 ( P1_R1192_U67 , P1_U3081 );
not NOT1_11378 ( P1_R1192_U68 , P1_U3982 );
not NOT1_11379 ( P1_R1192_U69 , P1_U3076 );
not NOT1_11380 ( P1_R1192_U70 , P1_U3979 );
not NOT1_11381 ( P1_R1192_U71 , P1_U3981 );
not NOT1_11382 ( P1_R1192_U72 , P1_U3066 );
not NOT1_11383 ( P1_R1192_U73 , P1_U3061 );
not NOT1_11384 ( P1_R1192_U74 , P1_U3075 );
nand NAND2_11385 ( P1_R1192_U75 , P1_U3075 , P1_R1192_U71 );
not NOT1_11386 ( P1_R1192_U76 , P1_U3978 );
not NOT1_11387 ( P1_R1192_U77 , P1_U3065 );
not NOT1_11388 ( P1_R1192_U78 , P1_U3977 );
not NOT1_11389 ( P1_R1192_U79 , P1_U3058 );
not NOT1_11390 ( P1_R1192_U80 , P1_U3975 );
not NOT1_11391 ( P1_R1192_U81 , P1_U3057 );
nand NAND2_11392 ( P1_R1192_U82 , P1_U3057 , P1_R1192_U44 );
not NOT1_11393 ( P1_R1192_U83 , P1_U3053 );
not NOT1_11394 ( P1_R1192_U84 , P1_U3974 );
not NOT1_11395 ( P1_R1192_U85 , P1_U3054 );
nand NAND2_11396 ( P1_R1192_U86 , P1_R1192_U126 , P1_R1192_U297 );
nand NAND2_11397 ( P1_R1192_U87 , P1_R1192_U294 , P1_R1192_U293 );
nand NAND2_11398 ( P1_R1192_U88 , P1_R1192_U75 , P1_R1192_U314 );
nand NAND2_11399 ( P1_R1192_U89 , P1_R1192_U61 , P1_R1192_U325 );
nand NAND2_11400 ( P1_R1192_U90 , P1_R1192_U51 , P1_R1192_U336 );
not NOT1_11401 ( P1_R1192_U91 , P1_U3077 );
nand NAND2_11402 ( P1_R1192_U92 , P1_R1192_U390 , P1_R1192_U389 );
nand NAND2_11403 ( P1_R1192_U93 , P1_R1192_U404 , P1_R1192_U403 );
nand NAND2_11404 ( P1_R1192_U94 , P1_R1192_U409 , P1_R1192_U408 );
nand NAND2_11405 ( P1_R1192_U95 , P1_R1192_U425 , P1_R1192_U424 );
nand NAND2_11406 ( P1_R1192_U96 , P1_R1192_U430 , P1_R1192_U429 );
nand NAND2_11407 ( P1_R1192_U97 , P1_R1192_U435 , P1_R1192_U434 );
nand NAND2_11408 ( P1_R1192_U98 , P1_R1192_U440 , P1_R1192_U439 );
nand NAND2_11409 ( P1_R1192_U99 , P1_R1192_U445 , P1_R1192_U444 );
nand NAND2_11410 ( P1_R1192_U100 , P1_R1192_U461 , P1_R1192_U460 );
nand NAND2_11411 ( P1_R1192_U101 , P1_R1192_U466 , P1_R1192_U465 );
nand NAND2_11412 ( P1_R1192_U102 , P1_R1192_U351 , P1_R1192_U350 );
nand NAND2_11413 ( P1_R1192_U103 , P1_R1192_U360 , P1_R1192_U359 );
nand NAND2_11414 ( P1_R1192_U104 , P1_R1192_U367 , P1_R1192_U366 );
nand NAND2_11415 ( P1_R1192_U105 , P1_R1192_U371 , P1_R1192_U370 );
nand NAND2_11416 ( P1_R1192_U106 , P1_R1192_U380 , P1_R1192_U379 );
nand NAND2_11417 ( P1_R1192_U107 , P1_R1192_U399 , P1_R1192_U398 );
nand NAND2_11418 ( P1_R1192_U108 , P1_R1192_U416 , P1_R1192_U415 );
nand NAND2_11419 ( P1_R1192_U109 , P1_R1192_U420 , P1_R1192_U419 );
nand NAND2_11420 ( P1_R1192_U110 , P1_R1192_U452 , P1_R1192_U451 );
nand NAND2_11421 ( P1_R1192_U111 , P1_R1192_U456 , P1_R1192_U455 );
nand NAND2_11422 ( P1_R1192_U112 , P1_R1192_U473 , P1_R1192_U472 );
and AND2_11423 ( P1_R1192_U113 , P1_R1192_U193 , P1_R1192_U194 );
and AND2_11424 ( P1_R1192_U114 , P1_R1192_U201 , P1_R1192_U196 );
and AND2_11425 ( P1_R1192_U115 , P1_R1192_U206 , P1_R1192_U180 );
and AND2_11426 ( P1_R1192_U116 , P1_R1192_U209 , P1_R1192_U210 );
and AND3_11427 ( P1_R1192_U117 , P1_R1192_U353 , P1_R1192_U352 , P1_R1192_U37 );
and AND2_11428 ( P1_R1192_U118 , P1_R1192_U356 , P1_R1192_U180 );
and AND2_11429 ( P1_R1192_U119 , P1_R1192_U225 , P1_R1192_U6 );
and AND2_11430 ( P1_R1192_U120 , P1_R1192_U363 , P1_R1192_U179 );
and AND3_11431 ( P1_R1192_U121 , P1_R1192_U373 , P1_R1192_U372 , P1_R1192_U27 );
and AND2_11432 ( P1_R1192_U122 , P1_R1192_U376 , P1_R1192_U178 );
and AND3_11433 ( P1_R1192_U123 , P1_R1192_U235 , P1_R1192_U212 , P1_R1192_U174 );
and AND3_11434 ( P1_R1192_U124 , P1_R1192_U257 , P1_R1192_U175 , P1_R1192_U252 );
and AND2_11435 ( P1_R1192_U125 , P1_R1192_U283 , P1_R1192_U176 );
and AND2_11436 ( P1_R1192_U126 , P1_R1192_U299 , P1_R1192_U300 );
nand NAND2_11437 ( P1_R1192_U127 , P1_R1192_U387 , P1_R1192_U386 );
and AND3_11438 ( P1_R1192_U128 , P1_R1192_U392 , P1_R1192_U391 , P1_R1192_U82 );
and AND2_11439 ( P1_R1192_U129 , P1_R1192_U395 , P1_R1192_U177 );
nand NAND2_11440 ( P1_R1192_U130 , P1_R1192_U401 , P1_R1192_U400 );
nand NAND2_11441 ( P1_R1192_U131 , P1_R1192_U406 , P1_R1192_U405 );
and AND2_11442 ( P1_R1192_U132 , P1_R1192_U412 , P1_R1192_U176 );
nand NAND2_11443 ( P1_R1192_U133 , P1_R1192_U422 , P1_R1192_U421 );
nand NAND2_11444 ( P1_R1192_U134 , P1_R1192_U427 , P1_R1192_U426 );
nand NAND2_11445 ( P1_R1192_U135 , P1_R1192_U432 , P1_R1192_U431 );
nand NAND2_11446 ( P1_R1192_U136 , P1_R1192_U437 , P1_R1192_U436 );
nand NAND2_11447 ( P1_R1192_U137 , P1_R1192_U442 , P1_R1192_U441 );
and AND2_11448 ( P1_R1192_U138 , P1_R1192_U331 , P1_R1192_U8 );
and AND2_11449 ( P1_R1192_U139 , P1_R1192_U448 , P1_R1192_U175 );
nand NAND2_11450 ( P1_R1192_U140 , P1_R1192_U458 , P1_R1192_U457 );
nand NAND2_11451 ( P1_R1192_U141 , P1_R1192_U463 , P1_R1192_U462 );
and AND2_11452 ( P1_R1192_U142 , P1_R1192_U342 , P1_R1192_U7 );
and AND2_11453 ( P1_R1192_U143 , P1_R1192_U469 , P1_R1192_U174 );
and AND2_11454 ( P1_R1192_U144 , P1_R1192_U349 , P1_R1192_U348 );
nand NAND2_11455 ( P1_R1192_U145 , P1_R1192_U116 , P1_R1192_U207 );
and AND2_11456 ( P1_R1192_U146 , P1_R1192_U358 , P1_R1192_U357 );
and AND2_11457 ( P1_R1192_U147 , P1_R1192_U365 , P1_R1192_U364 );
and AND2_11458 ( P1_R1192_U148 , P1_R1192_U369 , P1_R1192_U368 );
nand NAND2_11459 ( P1_R1192_U149 , P1_R1192_U113 , P1_R1192_U191 );
and AND2_11460 ( P1_R1192_U150 , P1_R1192_U378 , P1_R1192_U377 );
not NOT1_11461 ( P1_R1192_U151 , P1_U3985 );
not NOT1_11462 ( P1_R1192_U152 , P1_U3055 );
and AND2_11463 ( P1_R1192_U153 , P1_R1192_U382 , P1_R1192_U381 );
and AND2_11464 ( P1_R1192_U154 , P1_R1192_U397 , P1_R1192_U396 );
nand NAND2_11465 ( P1_R1192_U155 , P1_R1192_U290 , P1_R1192_U289 );
nand NAND2_11466 ( P1_R1192_U156 , P1_R1192_U286 , P1_R1192_U285 );
and AND2_11467 ( P1_R1192_U157 , P1_R1192_U414 , P1_R1192_U413 );
and AND2_11468 ( P1_R1192_U158 , P1_R1192_U418 , P1_R1192_U417 );
nand NAND2_11469 ( P1_R1192_U159 , P1_R1192_U276 , P1_R1192_U275 );
nand NAND2_11470 ( P1_R1192_U160 , P1_R1192_U272 , P1_R1192_U271 );
not NOT1_11471 ( P1_R1192_U161 , P1_U3455 );
nand NAND2_11472 ( P1_R1192_U162 , P1_R1192_U268 , P1_R1192_U267 );
not NOT1_11473 ( P1_R1192_U163 , P1_U3506 );
nand NAND2_11474 ( P1_R1192_U164 , P1_R1192_U260 , P1_R1192_U259 );
and AND2_11475 ( P1_R1192_U165 , P1_R1192_U450 , P1_R1192_U449 );
and AND2_11476 ( P1_R1192_U166 , P1_R1192_U454 , P1_R1192_U453 );
nand NAND2_11477 ( P1_R1192_U167 , P1_R1192_U250 , P1_R1192_U249 );
nand NAND2_11478 ( P1_R1192_U168 , P1_R1192_U246 , P1_R1192_U245 );
nand NAND2_11479 ( P1_R1192_U169 , P1_R1192_U242 , P1_R1192_U241 );
and AND2_11480 ( P1_R1192_U170 , P1_R1192_U471 , P1_R1192_U470 );
not NOT1_11481 ( P1_R1192_U171 , P1_R1192_U82 );
not NOT1_11482 ( P1_R1192_U172 , P1_R1192_U27 );
not NOT1_11483 ( P1_R1192_U173 , P1_R1192_U37 );
nand NAND2_11484 ( P1_R1192_U174 , P1_U3482 , P1_R1192_U50 );
nand NAND2_11485 ( P1_R1192_U175 , P1_U3497 , P1_R1192_U59 );
nand NAND2_11486 ( P1_R1192_U176 , P1_U3980 , P1_R1192_U73 );
nand NAND2_11487 ( P1_R1192_U177 , P1_U3976 , P1_R1192_U81 );
nand NAND2_11488 ( P1_R1192_U178 , P1_U3458 , P1_R1192_U26 );
nand NAND2_11489 ( P1_R1192_U179 , P1_U3467 , P1_R1192_U32 );
nand NAND2_11490 ( P1_R1192_U180 , P1_U3473 , P1_R1192_U36 );
not NOT1_11491 ( P1_R1192_U181 , P1_R1192_U61 );
not NOT1_11492 ( P1_R1192_U182 , P1_R1192_U75 );
not NOT1_11493 ( P1_R1192_U183 , P1_R1192_U34 );
not NOT1_11494 ( P1_R1192_U184 , P1_R1192_U51 );
not NOT1_11495 ( P1_R1192_U185 , P1_R1192_U23 );
nand NAND2_11496 ( P1_R1192_U186 , P1_R1192_U185 , P1_R1192_U24 );
nand NAND2_11497 ( P1_R1192_U187 , P1_R1192_U186 , P1_R1192_U161 );
nand NAND2_11498 ( P1_R1192_U188 , P1_U3078 , P1_R1192_U23 );
not NOT1_11499 ( P1_R1192_U189 , P1_R1192_U43 );
nand NAND2_11500 ( P1_R1192_U190 , P1_U3461 , P1_R1192_U28 );
nand NAND3_11501 ( P1_R1192_U191 , P1_R1192_U43 , P1_R1192_U178 , P1_R1192_U190 );
nand NAND2_11502 ( P1_R1192_U192 , P1_R1192_U28 , P1_R1192_U27 );
nand NAND2_11503 ( P1_R1192_U193 , P1_R1192_U192 , P1_R1192_U25 );
nand NAND2_11504 ( P1_R1192_U194 , P1_U3064 , P1_R1192_U172 );
not NOT1_11505 ( P1_R1192_U195 , P1_R1192_U149 );
nand NAND2_11506 ( P1_R1192_U196 , P1_U3470 , P1_R1192_U31 );
nand NAND2_11507 ( P1_R1192_U197 , P1_U3071 , P1_R1192_U29 );
nand NAND2_11508 ( P1_R1192_U198 , P1_U3067 , P1_R1192_U20 );
nand NAND2_11509 ( P1_R1192_U199 , P1_R1192_U183 , P1_R1192_U179 );
nand NAND2_11510 ( P1_R1192_U200 , P1_R1192_U6 , P1_R1192_U199 );
nand NAND2_11511 ( P1_R1192_U201 , P1_U3464 , P1_R1192_U33 );
nand NAND2_11512 ( P1_R1192_U202 , P1_U3470 , P1_R1192_U31 );
nand NAND3_11513 ( P1_R1192_U203 , P1_R1192_U149 , P1_R1192_U179 , P1_R1192_U114 );
nand NAND2_11514 ( P1_R1192_U204 , P1_R1192_U202 , P1_R1192_U200 );
not NOT1_11515 ( P1_R1192_U205 , P1_R1192_U41 );
nand NAND2_11516 ( P1_R1192_U206 , P1_U3476 , P1_R1192_U38 );
nand NAND2_11517 ( P1_R1192_U207 , P1_R1192_U115 , P1_R1192_U41 );
nand NAND2_11518 ( P1_R1192_U208 , P1_R1192_U38 , P1_R1192_U37 );
nand NAND2_11519 ( P1_R1192_U209 , P1_R1192_U208 , P1_R1192_U35 );
nand NAND2_11520 ( P1_R1192_U210 , P1_U3084 , P1_R1192_U173 );
not NOT1_11521 ( P1_R1192_U211 , P1_R1192_U145 );
nand NAND2_11522 ( P1_R1192_U212 , P1_U3479 , P1_R1192_U40 );
nand NAND2_11523 ( P1_R1192_U213 , P1_R1192_U212 , P1_R1192_U51 );
nand NAND2_11524 ( P1_R1192_U214 , P1_R1192_U205 , P1_R1192_U37 );
nand NAND2_11525 ( P1_R1192_U215 , P1_R1192_U118 , P1_R1192_U214 );
nand NAND2_11526 ( P1_R1192_U216 , P1_R1192_U41 , P1_R1192_U180 );
nand NAND2_11527 ( P1_R1192_U217 , P1_R1192_U117 , P1_R1192_U216 );
nand NAND2_11528 ( P1_R1192_U218 , P1_R1192_U37 , P1_R1192_U180 );
nand NAND2_11529 ( P1_R1192_U219 , P1_R1192_U201 , P1_R1192_U149 );
not NOT1_11530 ( P1_R1192_U220 , P1_R1192_U42 );
nand NAND2_11531 ( P1_R1192_U221 , P1_U3067 , P1_R1192_U20 );
nand NAND2_11532 ( P1_R1192_U222 , P1_R1192_U220 , P1_R1192_U221 );
nand NAND2_11533 ( P1_R1192_U223 , P1_R1192_U120 , P1_R1192_U222 );
nand NAND2_11534 ( P1_R1192_U224 , P1_R1192_U42 , P1_R1192_U179 );
nand NAND2_11535 ( P1_R1192_U225 , P1_U3470 , P1_R1192_U31 );
nand NAND2_11536 ( P1_R1192_U226 , P1_R1192_U119 , P1_R1192_U224 );
nand NAND2_11537 ( P1_R1192_U227 , P1_U3067 , P1_R1192_U20 );
nand NAND2_11538 ( P1_R1192_U228 , P1_R1192_U179 , P1_R1192_U227 );
nand NAND2_11539 ( P1_R1192_U229 , P1_R1192_U201 , P1_R1192_U34 );
nand NAND2_11540 ( P1_R1192_U230 , P1_R1192_U189 , P1_R1192_U27 );
nand NAND2_11541 ( P1_R1192_U231 , P1_R1192_U122 , P1_R1192_U230 );
nand NAND2_11542 ( P1_R1192_U232 , P1_R1192_U43 , P1_R1192_U178 );
nand NAND2_11543 ( P1_R1192_U233 , P1_R1192_U121 , P1_R1192_U232 );
nand NAND2_11544 ( P1_R1192_U234 , P1_R1192_U27 , P1_R1192_U178 );
nand NAND2_11545 ( P1_R1192_U235 , P1_U3485 , P1_R1192_U49 );
nand NAND2_11546 ( P1_R1192_U236 , P1_U3063 , P1_R1192_U48 );
nand NAND2_11547 ( P1_R1192_U237 , P1_U3062 , P1_R1192_U47 );
nand NAND2_11548 ( P1_R1192_U238 , P1_R1192_U184 , P1_R1192_U174 );
nand NAND2_11549 ( P1_R1192_U239 , P1_R1192_U7 , P1_R1192_U238 );
nand NAND2_11550 ( P1_R1192_U240 , P1_U3485 , P1_R1192_U49 );
nand NAND2_11551 ( P1_R1192_U241 , P1_R1192_U145 , P1_R1192_U123 );
nand NAND2_11552 ( P1_R1192_U242 , P1_R1192_U240 , P1_R1192_U239 );
not NOT1_11553 ( P1_R1192_U243 , P1_R1192_U169 );
nand NAND2_11554 ( P1_R1192_U244 , P1_U3488 , P1_R1192_U53 );
nand NAND2_11555 ( P1_R1192_U245 , P1_R1192_U244 , P1_R1192_U169 );
nand NAND2_11556 ( P1_R1192_U246 , P1_U3072 , P1_R1192_U52 );
not NOT1_11557 ( P1_R1192_U247 , P1_R1192_U168 );
nand NAND2_11558 ( P1_R1192_U248 , P1_U3491 , P1_R1192_U55 );
nand NAND2_11559 ( P1_R1192_U249 , P1_R1192_U248 , P1_R1192_U168 );
nand NAND2_11560 ( P1_R1192_U250 , P1_U3080 , P1_R1192_U54 );
not NOT1_11561 ( P1_R1192_U251 , P1_R1192_U167 );
nand NAND2_11562 ( P1_R1192_U252 , P1_U3500 , P1_R1192_U58 );
nand NAND2_11563 ( P1_R1192_U253 , P1_U3073 , P1_R1192_U56 );
nand NAND2_11564 ( P1_R1192_U254 , P1_U3074 , P1_R1192_U46 );
nand NAND2_11565 ( P1_R1192_U255 , P1_R1192_U181 , P1_R1192_U175 );
nand NAND2_11566 ( P1_R1192_U256 , P1_R1192_U8 , P1_R1192_U255 );
nand NAND2_11567 ( P1_R1192_U257 , P1_U3494 , P1_R1192_U60 );
nand NAND2_11568 ( P1_R1192_U258 , P1_U3500 , P1_R1192_U58 );
nand NAND2_11569 ( P1_R1192_U259 , P1_R1192_U167 , P1_R1192_U124 );
nand NAND2_11570 ( P1_R1192_U260 , P1_R1192_U258 , P1_R1192_U256 );
not NOT1_11571 ( P1_R1192_U261 , P1_R1192_U164 );
nand NAND2_11572 ( P1_R1192_U262 , P1_U3503 , P1_R1192_U63 );
nand NAND2_11573 ( P1_R1192_U263 , P1_R1192_U262 , P1_R1192_U164 );
nand NAND2_11574 ( P1_R1192_U264 , P1_U3069 , P1_R1192_U62 );
not NOT1_11575 ( P1_R1192_U265 , P1_R1192_U64 );
nand NAND2_11576 ( P1_R1192_U266 , P1_R1192_U265 , P1_R1192_U65 );
nand NAND2_11577 ( P1_R1192_U267 , P1_R1192_U266 , P1_R1192_U163 );
nand NAND2_11578 ( P1_R1192_U268 , P1_U3082 , P1_R1192_U64 );
not NOT1_11579 ( P1_R1192_U269 , P1_R1192_U162 );
nand NAND2_11580 ( P1_R1192_U270 , P1_U3508 , P1_R1192_U67 );
nand NAND2_11581 ( P1_R1192_U271 , P1_R1192_U270 , P1_R1192_U162 );
nand NAND2_11582 ( P1_R1192_U272 , P1_U3081 , P1_R1192_U66 );
not NOT1_11583 ( P1_R1192_U273 , P1_R1192_U160 );
nand NAND2_11584 ( P1_R1192_U274 , P1_U3982 , P1_R1192_U69 );
nand NAND2_11585 ( P1_R1192_U275 , P1_R1192_U274 , P1_R1192_U160 );
nand NAND2_11586 ( P1_R1192_U276 , P1_U3076 , P1_R1192_U68 );
not NOT1_11587 ( P1_R1192_U277 , P1_R1192_U159 );
nand NAND2_11588 ( P1_R1192_U278 , P1_U3979 , P1_R1192_U72 );
nand NAND2_11589 ( P1_R1192_U279 , P1_U3066 , P1_R1192_U70 );
nand NAND2_11590 ( P1_R1192_U280 , P1_U3061 , P1_R1192_U45 );
nand NAND2_11591 ( P1_R1192_U281 , P1_R1192_U182 , P1_R1192_U176 );
nand NAND2_11592 ( P1_R1192_U282 , P1_R1192_U9 , P1_R1192_U281 );
nand NAND2_11593 ( P1_R1192_U283 , P1_U3981 , P1_R1192_U74 );
nand NAND2_11594 ( P1_R1192_U284 , P1_U3979 , P1_R1192_U72 );
nand NAND3_11595 ( P1_R1192_U285 , P1_R1192_U159 , P1_R1192_U125 , P1_R1192_U278 );
nand NAND2_11596 ( P1_R1192_U286 , P1_R1192_U284 , P1_R1192_U282 );
not NOT1_11597 ( P1_R1192_U287 , P1_R1192_U156 );
nand NAND2_11598 ( P1_R1192_U288 , P1_U3978 , P1_R1192_U77 );
nand NAND2_11599 ( P1_R1192_U289 , P1_R1192_U288 , P1_R1192_U156 );
nand NAND2_11600 ( P1_R1192_U290 , P1_U3065 , P1_R1192_U76 );
not NOT1_11601 ( P1_R1192_U291 , P1_R1192_U155 );
nand NAND2_11602 ( P1_R1192_U292 , P1_U3977 , P1_R1192_U79 );
nand NAND2_11603 ( P1_R1192_U293 , P1_R1192_U292 , P1_R1192_U155 );
nand NAND2_11604 ( P1_R1192_U294 , P1_U3058 , P1_R1192_U78 );
not NOT1_11605 ( P1_R1192_U295 , P1_R1192_U87 );
nand NAND2_11606 ( P1_R1192_U296 , P1_U3975 , P1_R1192_U83 );
nand NAND3_11607 ( P1_R1192_U297 , P1_R1192_U87 , P1_R1192_U177 , P1_R1192_U296 );
nand NAND2_11608 ( P1_R1192_U298 , P1_R1192_U83 , P1_R1192_U82 );
nand NAND2_11609 ( P1_R1192_U299 , P1_R1192_U298 , P1_R1192_U80 );
nand NAND2_11610 ( P1_R1192_U300 , P1_U3053 , P1_R1192_U171 );
not NOT1_11611 ( P1_R1192_U301 , P1_R1192_U86 );
nand NAND2_11612 ( P1_R1192_U302 , P1_U3054 , P1_R1192_U84 );
nand NAND2_11613 ( P1_R1192_U303 , P1_R1192_U301 , P1_R1192_U302 );
nand NAND2_11614 ( P1_R1192_U304 , P1_U3974 , P1_R1192_U85 );
nand NAND2_11615 ( P1_R1192_U305 , P1_U3974 , P1_R1192_U85 );
nand NAND2_11616 ( P1_R1192_U306 , P1_R1192_U305 , P1_R1192_U86 );
nand NAND2_11617 ( P1_R1192_U307 , P1_U3054 , P1_R1192_U84 );
nand NAND3_11618 ( P1_R1192_U308 , P1_R1192_U307 , P1_R1192_U306 , P1_R1192_U153 );
nand NAND2_11619 ( P1_R1192_U309 , P1_R1192_U295 , P1_R1192_U82 );
nand NAND2_11620 ( P1_R1192_U310 , P1_R1192_U129 , P1_R1192_U309 );
nand NAND2_11621 ( P1_R1192_U311 , P1_R1192_U87 , P1_R1192_U177 );
nand NAND2_11622 ( P1_R1192_U312 , P1_R1192_U128 , P1_R1192_U311 );
nand NAND2_11623 ( P1_R1192_U313 , P1_R1192_U82 , P1_R1192_U177 );
nand NAND2_11624 ( P1_R1192_U314 , P1_R1192_U283 , P1_R1192_U159 );
not NOT1_11625 ( P1_R1192_U315 , P1_R1192_U88 );
nand NAND2_11626 ( P1_R1192_U316 , P1_U3061 , P1_R1192_U45 );
nand NAND2_11627 ( P1_R1192_U317 , P1_R1192_U315 , P1_R1192_U316 );
nand NAND2_11628 ( P1_R1192_U318 , P1_R1192_U132 , P1_R1192_U317 );
nand NAND2_11629 ( P1_R1192_U319 , P1_R1192_U88 , P1_R1192_U176 );
nand NAND2_11630 ( P1_R1192_U320 , P1_U3979 , P1_R1192_U72 );
nand NAND3_11631 ( P1_R1192_U321 , P1_R1192_U320 , P1_R1192_U319 , P1_R1192_U9 );
nand NAND2_11632 ( P1_R1192_U322 , P1_U3061 , P1_R1192_U45 );
nand NAND2_11633 ( P1_R1192_U323 , P1_R1192_U176 , P1_R1192_U322 );
nand NAND2_11634 ( P1_R1192_U324 , P1_R1192_U283 , P1_R1192_U75 );
nand NAND2_11635 ( P1_R1192_U325 , P1_R1192_U257 , P1_R1192_U167 );
not NOT1_11636 ( P1_R1192_U326 , P1_R1192_U89 );
nand NAND2_11637 ( P1_R1192_U327 , P1_U3074 , P1_R1192_U46 );
nand NAND2_11638 ( P1_R1192_U328 , P1_R1192_U326 , P1_R1192_U327 );
nand NAND2_11639 ( P1_R1192_U329 , P1_R1192_U139 , P1_R1192_U328 );
nand NAND2_11640 ( P1_R1192_U330 , P1_R1192_U89 , P1_R1192_U175 );
nand NAND2_11641 ( P1_R1192_U331 , P1_U3500 , P1_R1192_U58 );
nand NAND2_11642 ( P1_R1192_U332 , P1_R1192_U138 , P1_R1192_U330 );
nand NAND2_11643 ( P1_R1192_U333 , P1_U3074 , P1_R1192_U46 );
nand NAND2_11644 ( P1_R1192_U334 , P1_R1192_U175 , P1_R1192_U333 );
nand NAND2_11645 ( P1_R1192_U335 , P1_R1192_U257 , P1_R1192_U61 );
nand NAND2_11646 ( P1_R1192_U336 , P1_R1192_U212 , P1_R1192_U145 );
not NOT1_11647 ( P1_R1192_U337 , P1_R1192_U90 );
nand NAND2_11648 ( P1_R1192_U338 , P1_U3062 , P1_R1192_U47 );
nand NAND2_11649 ( P1_R1192_U339 , P1_R1192_U337 , P1_R1192_U338 );
nand NAND2_11650 ( P1_R1192_U340 , P1_R1192_U143 , P1_R1192_U339 );
nand NAND2_11651 ( P1_R1192_U341 , P1_R1192_U90 , P1_R1192_U174 );
nand NAND2_11652 ( P1_R1192_U342 , P1_U3485 , P1_R1192_U49 );
nand NAND2_11653 ( P1_R1192_U343 , P1_R1192_U142 , P1_R1192_U341 );
nand NAND2_11654 ( P1_R1192_U344 , P1_U3062 , P1_R1192_U47 );
nand NAND2_11655 ( P1_R1192_U345 , P1_R1192_U174 , P1_R1192_U344 );
nand NAND2_11656 ( P1_R1192_U346 , P1_U3077 , P1_R1192_U22 );
nand NAND3_11657 ( P1_R1192_U347 , P1_R1192_U304 , P1_R1192_U303 , P1_R1192_U385 );
nand NAND2_11658 ( P1_R1192_U348 , P1_U3479 , P1_R1192_U40 );
nand NAND2_11659 ( P1_R1192_U349 , P1_U3083 , P1_R1192_U39 );
nand NAND2_11660 ( P1_R1192_U350 , P1_R1192_U213 , P1_R1192_U145 );
nand NAND2_11661 ( P1_R1192_U351 , P1_R1192_U211 , P1_R1192_U144 );
nand NAND2_11662 ( P1_R1192_U352 , P1_U3476 , P1_R1192_U38 );
nand NAND2_11663 ( P1_R1192_U353 , P1_U3084 , P1_R1192_U35 );
nand NAND2_11664 ( P1_R1192_U354 , P1_U3476 , P1_R1192_U38 );
nand NAND2_11665 ( P1_R1192_U355 , P1_U3084 , P1_R1192_U35 );
nand NAND2_11666 ( P1_R1192_U356 , P1_R1192_U355 , P1_R1192_U354 );
nand NAND2_11667 ( P1_R1192_U357 , P1_U3473 , P1_R1192_U36 );
nand NAND2_11668 ( P1_R1192_U358 , P1_U3070 , P1_R1192_U19 );
nand NAND2_11669 ( P1_R1192_U359 , P1_R1192_U218 , P1_R1192_U41 );
nand NAND2_11670 ( P1_R1192_U360 , P1_R1192_U146 , P1_R1192_U205 );
nand NAND2_11671 ( P1_R1192_U361 , P1_U3470 , P1_R1192_U31 );
nand NAND2_11672 ( P1_R1192_U362 , P1_U3071 , P1_R1192_U29 );
nand NAND2_11673 ( P1_R1192_U363 , P1_R1192_U362 , P1_R1192_U361 );
nand NAND2_11674 ( P1_R1192_U364 , P1_U3467 , P1_R1192_U32 );
nand NAND2_11675 ( P1_R1192_U365 , P1_U3067 , P1_R1192_U20 );
nand NAND2_11676 ( P1_R1192_U366 , P1_R1192_U228 , P1_R1192_U42 );
nand NAND2_11677 ( P1_R1192_U367 , P1_R1192_U147 , P1_R1192_U220 );
nand NAND2_11678 ( P1_R1192_U368 , P1_U3464 , P1_R1192_U33 );
nand NAND2_11679 ( P1_R1192_U369 , P1_U3060 , P1_R1192_U30 );
nand NAND2_11680 ( P1_R1192_U370 , P1_R1192_U229 , P1_R1192_U149 );
nand NAND2_11681 ( P1_R1192_U371 , P1_R1192_U195 , P1_R1192_U148 );
nand NAND2_11682 ( P1_R1192_U372 , P1_U3461 , P1_R1192_U28 );
nand NAND2_11683 ( P1_R1192_U373 , P1_U3064 , P1_R1192_U25 );
nand NAND2_11684 ( P1_R1192_U374 , P1_U3461 , P1_R1192_U28 );
nand NAND2_11685 ( P1_R1192_U375 , P1_U3064 , P1_R1192_U25 );
nand NAND2_11686 ( P1_R1192_U376 , P1_R1192_U375 , P1_R1192_U374 );
nand NAND2_11687 ( P1_R1192_U377 , P1_U3458 , P1_R1192_U26 );
nand NAND2_11688 ( P1_R1192_U378 , P1_U3068 , P1_R1192_U21 );
nand NAND2_11689 ( P1_R1192_U379 , P1_R1192_U234 , P1_R1192_U43 );
nand NAND2_11690 ( P1_R1192_U380 , P1_R1192_U150 , P1_R1192_U189 );
nand NAND2_11691 ( P1_R1192_U381 , P1_U3985 , P1_R1192_U152 );
nand NAND2_11692 ( P1_R1192_U382 , P1_U3055 , P1_R1192_U151 );
nand NAND2_11693 ( P1_R1192_U383 , P1_U3985 , P1_R1192_U152 );
nand NAND2_11694 ( P1_R1192_U384 , P1_U3055 , P1_R1192_U151 );
nand NAND2_11695 ( P1_R1192_U385 , P1_R1192_U384 , P1_R1192_U383 );
nand NAND2_11696 ( P1_R1192_U386 , P1_U3974 , P1_R1192_U85 );
nand NAND2_11697 ( P1_R1192_U387 , P1_U3054 , P1_R1192_U84 );
not NOT1_11698 ( P1_R1192_U388 , P1_R1192_U127 );
nand NAND2_11699 ( P1_R1192_U389 , P1_R1192_U388 , P1_R1192_U301 );
nand NAND2_11700 ( P1_R1192_U390 , P1_R1192_U127 , P1_R1192_U86 );
nand NAND2_11701 ( P1_R1192_U391 , P1_U3975 , P1_R1192_U83 );
nand NAND2_11702 ( P1_R1192_U392 , P1_U3053 , P1_R1192_U80 );
nand NAND2_11703 ( P1_R1192_U393 , P1_U3975 , P1_R1192_U83 );
nand NAND2_11704 ( P1_R1192_U394 , P1_U3053 , P1_R1192_U80 );
nand NAND2_11705 ( P1_R1192_U395 , P1_R1192_U394 , P1_R1192_U393 );
nand NAND2_11706 ( P1_R1192_U396 , P1_U3976 , P1_R1192_U81 );
nand NAND2_11707 ( P1_R1192_U397 , P1_U3057 , P1_R1192_U44 );
nand NAND2_11708 ( P1_R1192_U398 , P1_R1192_U313 , P1_R1192_U87 );
nand NAND2_11709 ( P1_R1192_U399 , P1_R1192_U154 , P1_R1192_U295 );
nand NAND2_11710 ( P1_R1192_U400 , P1_U3977 , P1_R1192_U79 );
nand NAND2_11711 ( P1_R1192_U401 , P1_U3058 , P1_R1192_U78 );
not NOT1_11712 ( P1_R1192_U402 , P1_R1192_U130 );
nand NAND2_11713 ( P1_R1192_U403 , P1_R1192_U291 , P1_R1192_U402 );
nand NAND2_11714 ( P1_R1192_U404 , P1_R1192_U130 , P1_R1192_U155 );
nand NAND2_11715 ( P1_R1192_U405 , P1_U3978 , P1_R1192_U77 );
nand NAND2_11716 ( P1_R1192_U406 , P1_U3065 , P1_R1192_U76 );
not NOT1_11717 ( P1_R1192_U407 , P1_R1192_U131 );
nand NAND2_11718 ( P1_R1192_U408 , P1_R1192_U287 , P1_R1192_U407 );
nand NAND2_11719 ( P1_R1192_U409 , P1_R1192_U131 , P1_R1192_U156 );
nand NAND2_11720 ( P1_R1192_U410 , P1_U3979 , P1_R1192_U72 );
nand NAND2_11721 ( P1_R1192_U411 , P1_U3066 , P1_R1192_U70 );
nand NAND2_11722 ( P1_R1192_U412 , P1_R1192_U411 , P1_R1192_U410 );
nand NAND2_11723 ( P1_R1192_U413 , P1_U3980 , P1_R1192_U73 );
nand NAND2_11724 ( P1_R1192_U414 , P1_U3061 , P1_R1192_U45 );
nand NAND2_11725 ( P1_R1192_U415 , P1_R1192_U323 , P1_R1192_U88 );
nand NAND2_11726 ( P1_R1192_U416 , P1_R1192_U157 , P1_R1192_U315 );
nand NAND2_11727 ( P1_R1192_U417 , P1_U3981 , P1_R1192_U74 );
nand NAND2_11728 ( P1_R1192_U418 , P1_U3075 , P1_R1192_U71 );
nand NAND2_11729 ( P1_R1192_U419 , P1_R1192_U324 , P1_R1192_U159 );
nand NAND2_11730 ( P1_R1192_U420 , P1_R1192_U277 , P1_R1192_U158 );
nand NAND2_11731 ( P1_R1192_U421 , P1_U3982 , P1_R1192_U69 );
nand NAND2_11732 ( P1_R1192_U422 , P1_U3076 , P1_R1192_U68 );
not NOT1_11733 ( P1_R1192_U423 , P1_R1192_U133 );
nand NAND2_11734 ( P1_R1192_U424 , P1_R1192_U273 , P1_R1192_U423 );
nand NAND2_11735 ( P1_R1192_U425 , P1_R1192_U133 , P1_R1192_U160 );
nand NAND2_11736 ( P1_R1192_U426 , P1_R1192_U185 , P1_R1192_U24 );
nand NAND2_11737 ( P1_R1192_U427 , P1_U3078 , P1_R1192_U23 );
not NOT1_11738 ( P1_R1192_U428 , P1_R1192_U134 );
nand NAND2_11739 ( P1_R1192_U429 , P1_U3455 , P1_R1192_U428 );
nand NAND2_11740 ( P1_R1192_U430 , P1_R1192_U134 , P1_R1192_U161 );
nand NAND2_11741 ( P1_R1192_U431 , P1_U3508 , P1_R1192_U67 );
nand NAND2_11742 ( P1_R1192_U432 , P1_U3081 , P1_R1192_U66 );
not NOT1_11743 ( P1_R1192_U433 , P1_R1192_U135 );
nand NAND2_11744 ( P1_R1192_U434 , P1_R1192_U269 , P1_R1192_U433 );
nand NAND2_11745 ( P1_R1192_U435 , P1_R1192_U135 , P1_R1192_U162 );
nand NAND2_11746 ( P1_R1192_U436 , P1_U3506 , P1_R1192_U65 );
nand NAND2_11747 ( P1_R1192_U437 , P1_U3082 , P1_R1192_U163 );
not NOT1_11748 ( P1_R1192_U438 , P1_R1192_U136 );
nand NAND2_11749 ( P1_R1192_U439 , P1_R1192_U438 , P1_R1192_U265 );
nand NAND2_11750 ( P1_R1192_U440 , P1_R1192_U136 , P1_R1192_U64 );
nand NAND2_11751 ( P1_R1192_U441 , P1_U3503 , P1_R1192_U63 );
nand NAND2_11752 ( P1_R1192_U442 , P1_U3069 , P1_R1192_U62 );
not NOT1_11753 ( P1_R1192_U443 , P1_R1192_U137 );
nand NAND2_11754 ( P1_R1192_U444 , P1_R1192_U261 , P1_R1192_U443 );
nand NAND2_11755 ( P1_R1192_U445 , P1_R1192_U137 , P1_R1192_U164 );
nand NAND2_11756 ( P1_R1192_U446 , P1_U3500 , P1_R1192_U58 );
nand NAND2_11757 ( P1_R1192_U447 , P1_U3073 , P1_R1192_U56 );
nand NAND2_11758 ( P1_R1192_U448 , P1_R1192_U447 , P1_R1192_U446 );
nand NAND2_11759 ( P1_R1192_U449 , P1_U3497 , P1_R1192_U59 );
nand NAND2_11760 ( P1_R1192_U450 , P1_U3074 , P1_R1192_U46 );
nand NAND2_11761 ( P1_R1192_U451 , P1_R1192_U334 , P1_R1192_U89 );
nand NAND2_11762 ( P1_R1192_U452 , P1_R1192_U165 , P1_R1192_U326 );
nand NAND2_11763 ( P1_R1192_U453 , P1_U3494 , P1_R1192_U60 );
nand NAND2_11764 ( P1_R1192_U454 , P1_U3079 , P1_R1192_U57 );
nand NAND2_11765 ( P1_R1192_U455 , P1_R1192_U335 , P1_R1192_U167 );
nand NAND2_11766 ( P1_R1192_U456 , P1_R1192_U251 , P1_R1192_U166 );
nand NAND2_11767 ( P1_R1192_U457 , P1_U3491 , P1_R1192_U55 );
nand NAND2_11768 ( P1_R1192_U458 , P1_U3080 , P1_R1192_U54 );
not NOT1_11769 ( P1_R1192_U459 , P1_R1192_U140 );
nand NAND2_11770 ( P1_R1192_U460 , P1_R1192_U247 , P1_R1192_U459 );
nand NAND2_11771 ( P1_R1192_U461 , P1_R1192_U140 , P1_R1192_U168 );
nand NAND2_11772 ( P1_R1192_U462 , P1_U3488 , P1_R1192_U53 );
nand NAND2_11773 ( P1_R1192_U463 , P1_U3072 , P1_R1192_U52 );
not NOT1_11774 ( P1_R1192_U464 , P1_R1192_U141 );
nand NAND2_11775 ( P1_R1192_U465 , P1_R1192_U243 , P1_R1192_U464 );
nand NAND2_11776 ( P1_R1192_U466 , P1_R1192_U141 , P1_R1192_U169 );
nand NAND2_11777 ( P1_R1192_U467 , P1_U3485 , P1_R1192_U49 );
nand NAND2_11778 ( P1_R1192_U468 , P1_U3063 , P1_R1192_U48 );
nand NAND2_11779 ( P1_R1192_U469 , P1_R1192_U468 , P1_R1192_U467 );
nand NAND2_11780 ( P1_R1192_U470 , P1_U3482 , P1_R1192_U50 );
nand NAND2_11781 ( P1_R1192_U471 , P1_U3062 , P1_R1192_U47 );
nand NAND2_11782 ( P1_R1192_U472 , P1_R1192_U345 , P1_R1192_U90 );
nand NAND2_11783 ( P1_R1192_U473 , P1_R1192_U170 , P1_R1192_U337 );
and AND2_11784 ( P1_LT_197_U6 , P1_LT_197_U115 , P1_LT_197_U116 );
and AND2_11785 ( P1_LT_197_U7 , P1_LT_197_U117 , P1_LT_197_U118 );
and AND4_11786 ( P1_LT_197_U8 , P1_LT_197_U81 , P1_LT_197_U120 , P1_LT_197_U122 , P1_LT_197_U7 );
and AND2_11787 ( P1_LT_197_U9 , P1_LT_197_U130 , P1_LT_197_U129 );
and AND4_11788 ( P1_LT_197_U10 , P1_LT_197_U131 , P1_LT_197_U128 , P1_LT_197_U84 , P1_LT_197_U85 );
and AND2_11789 ( P1_LT_197_U11 , P1_LT_197_U145 , P1_LT_197_U144 );
and AND2_11790 ( P1_LT_197_U12 , P1_LT_197_U193 , P1_LT_197_U72 );
and AND2_11791 ( P1_LT_197_U13 , P1_LT_197_U200 , P1_LT_197_U199 );
not NOT1_11792 ( P1_LT_197_U14 , P1_U3983 );
not NOT1_11793 ( P1_LT_197_U15 , P1_U3593 );
not NOT1_11794 ( P1_LT_197_U16 , P1_U3594 );
not NOT1_11795 ( P1_LT_197_U17 , P1_U3598 );
not NOT1_11796 ( P1_LT_197_U18 , P1_U3599 );
not NOT1_11797 ( P1_LT_197_U19 , P1_U3977 );
not NOT1_11798 ( P1_LT_197_U20 , P1_U3978 );
not NOT1_11799 ( P1_LT_197_U21 , P1_U3603 );
not NOT1_11800 ( P1_LT_197_U22 , P1_U3981 );
not NOT1_11801 ( P1_LT_197_U23 , P1_U3604 );
not NOT1_11802 ( P1_LT_197_U24 , P1_U3982 );
not NOT1_11803 ( P1_LT_197_U25 , P1_U3508 );
not NOT1_11804 ( P1_LT_197_U26 , P1_U3608 );
not NOT1_11805 ( P1_LT_197_U27 , P1_U3506 );
not NOT1_11806 ( P1_LT_197_U28 , P1_U3609 );
not NOT1_11807 ( P1_LT_197_U29 , P1_U3607 );
not NOT1_11808 ( P1_LT_197_U30 , P1_U3605 );
not NOT1_11809 ( P1_LT_197_U31 , P1_U3503 );
not NOT1_11810 ( P1_LT_197_U32 , P1_U3500 );
not NOT1_11811 ( P1_LT_197_U33 , P1_U3610 );
not NOT1_11812 ( P1_LT_197_U34 , P1_U3611 );
not NOT1_11813 ( P1_LT_197_U35 , P1_U3473 );
not NOT1_11814 ( P1_LT_197_U36 , P1_U3589 );
not NOT1_11815 ( P1_LT_197_U37 , P1_U3470 );
not NOT1_11816 ( P1_LT_197_U38 , P1_U3590 );
not NOT1_11817 ( P1_LT_197_U39 , P1_U3586 );
not NOT1_11818 ( P1_LT_197_U40 , P1_U3616 );
not NOT1_11819 ( P1_LT_197_U41 , P1_U3587 );
not NOT1_11820 ( P1_LT_197_U42 , P1_U3588 );
not NOT1_11821 ( P1_LT_197_U43 , P1_U3591 );
not NOT1_11822 ( P1_LT_197_U44 , P1_U3592 );
nand NAND2_11823 ( P1_LT_197_U45 , P1_U3450 , P1_LT_197_U108 );
not NOT1_11824 ( P1_LT_197_U46 , P1_U3455 );
not NOT1_11825 ( P1_LT_197_U47 , P1_U3595 );
not NOT1_11826 ( P1_LT_197_U48 , P1_U3488 );
not NOT1_11827 ( P1_LT_197_U49 , P1_U3491 );
not NOT1_11828 ( P1_LT_197_U50 , P1_U3458 );
not NOT1_11829 ( P1_LT_197_U51 , P1_U3461 );
not NOT1_11830 ( P1_LT_197_U52 , P1_U3464 );
not NOT1_11831 ( P1_LT_197_U53 , P1_U3467 );
not NOT1_11832 ( P1_LT_197_U54 , P1_U3476 );
not NOT1_11833 ( P1_LT_197_U55 , P1_U3479 );
not NOT1_11834 ( P1_LT_197_U56 , P1_U3482 );
not NOT1_11835 ( P1_LT_197_U57 , P1_U3485 );
not NOT1_11836 ( P1_LT_197_U58 , P1_U3614 );
not NOT1_11837 ( P1_LT_197_U59 , P1_U3615 );
not NOT1_11838 ( P1_LT_197_U60 , P1_U3612 );
not NOT1_11839 ( P1_LT_197_U61 , P1_U3613 );
not NOT1_11840 ( P1_LT_197_U62 , P1_U3494 );
not NOT1_11841 ( P1_LT_197_U63 , P1_U3497 );
not NOT1_11842 ( P1_LT_197_U64 , P1_U3980 );
not NOT1_11843 ( P1_LT_197_U65 , P1_U3979 );
not NOT1_11844 ( P1_LT_197_U66 , P1_U3602 );
not NOT1_11845 ( P1_LT_197_U67 , P1_U3601 );
not NOT1_11846 ( P1_LT_197_U68 , P1_U3600 );
not NOT1_11847 ( P1_LT_197_U69 , P1_U3976 );
not NOT1_11848 ( P1_LT_197_U70 , P1_U3975 );
nand NAND2_11849 ( P1_LT_197_U71 , P1_LT_197_U192 , P1_LT_197_U191 );
not NOT1_11850 ( P1_LT_197_U72 , P1_U3974 );
not NOT1_11851 ( P1_LT_197_U73 , P1_U3985 );
not NOT1_11852 ( P1_LT_197_U74 , P1_U3596 );
not NOT1_11853 ( P1_LT_197_U75 , P1_U3984 );
and AND2_11854 ( P1_LT_197_U76 , P1_U3981 , P1_LT_197_U23 );
and AND2_11855 ( P1_LT_197_U77 , P1_U3982 , P1_LT_197_U30 );
and AND2_11856 ( P1_LT_197_U78 , P1_LT_197_U175 , P1_LT_197_U174 );
and AND2_11857 ( P1_LT_197_U79 , P1_U3608 , P1_LT_197_U27 );
and AND2_11858 ( P1_LT_197_U80 , P1_U3609 , P1_LT_197_U31 );
and AND2_11859 ( P1_LT_197_U81 , P1_LT_197_U121 , P1_LT_197_U119 );
and AND2_11860 ( P1_LT_197_U82 , P1_U3589 , P1_LT_197_U37 );
and AND2_11861 ( P1_LT_197_U83 , P1_U3590 , P1_LT_197_U53 );
and AND2_11862 ( P1_LT_197_U84 , P1_LT_197_U133 , P1_LT_197_U132 );
and AND4_11863 ( P1_LT_197_U85 , P1_LT_197_U137 , P1_LT_197_U136 , P1_LT_197_U135 , P1_LT_197_U134 );
and AND2_11864 ( P1_LT_197_U86 , P1_LT_197_U141 , P1_LT_197_U142 );
and AND2_11865 ( P1_LT_197_U87 , P1_LT_197_U86 , P1_LT_197_U140 );
and AND2_11866 ( P1_LT_197_U88 , P1_U3458 , P1_LT_197_U47 );
and AND2_11867 ( P1_LT_197_U89 , P1_U3461 , P1_LT_197_U44 );
and AND3_11868 ( P1_LT_197_U90 , P1_LT_197_U135 , P1_LT_197_U128 , P1_LT_197_U134 );
and AND3_11869 ( P1_LT_197_U91 , P1_LT_197_U158 , P1_LT_197_U143 , P1_LT_197_U93 );
and AND2_11870 ( P1_LT_197_U92 , P1_LT_197_U161 , P1_LT_197_U160 );
and AND2_11871 ( P1_LT_197_U93 , P1_LT_197_U92 , P1_LT_197_U11 );
and AND2_11872 ( P1_LT_197_U94 , P1_U3614 , P1_LT_197_U48 );
and AND2_11873 ( P1_LT_197_U95 , P1_U3615 , P1_LT_197_U57 );
and AND2_11874 ( P1_LT_197_U96 , P1_LT_197_U164 , P1_LT_197_U98 );
and AND2_11875 ( P1_LT_197_U97 , P1_LT_197_U96 , P1_LT_197_U165 );
and AND2_11876 ( P1_LT_197_U98 , P1_LT_197_U167 , P1_LT_197_U166 );
and AND2_11877 ( P1_LT_197_U99 , P1_LT_197_U177 , P1_LT_197_U124 );
and AND2_11878 ( P1_LT_197_U100 , P1_LT_197_U179 , P1_LT_197_U178 );
and AND2_11879 ( P1_LT_197_U101 , P1_LT_197_U181 , P1_LT_197_U182 );
and AND2_11880 ( P1_LT_197_U102 , P1_U3602 , P1_LT_197_U65 );
and AND2_11881 ( P1_LT_197_U103 , P1_LT_197_U186 , P1_LT_197_U185 );
and AND2_11882 ( P1_LT_197_U104 , P1_LT_197_U189 , P1_LT_197_U125 );
and AND2_11883 ( P1_LT_197_U105 , P1_LT_197_U196 , P1_LT_197_U195 );
and AND2_11884 ( P1_LT_197_U106 , P1_U3596 , P1_LT_197_U73 );
and AND2_11885 ( P1_LT_197_U107 , P1_LT_197_U198 , P1_LT_197_U112 );
not NOT1_11886 ( P1_LT_197_U108 , P1_U3617 );
nand NAND2_11887 ( P1_LT_197_U109 , P1_LT_197_U107 , P1_LT_197_U197 );
nand NAND2_11888 ( P1_LT_197_U110 , P1_U3984 , P1_LT_197_U16 );
nand NAND2_11889 ( P1_LT_197_U111 , P1_U3593 , P1_LT_197_U14 );
nand NAND3_11890 ( P1_LT_197_U112 , P1_LT_197_U111 , P1_U3594 , P1_LT_197_U75 );
nand NAND2_11891 ( P1_LT_197_U113 , P1_U3593 , P1_LT_197_U14 );
nand NAND2_11892 ( P1_LT_197_U114 , P1_U3598 , P1_LT_197_U70 );
nand NAND2_11893 ( P1_LT_197_U115 , P1_U3508 , P1_LT_197_U29 );
nand NAND2_11894 ( P1_LT_197_U116 , P1_U3506 , P1_LT_197_U26 );
nand NAND2_11895 ( P1_LT_197_U117 , P1_U3603 , P1_LT_197_U64 );
nand NAND2_11896 ( P1_LT_197_U118 , P1_U3604 , P1_LT_197_U22 );
nand NAND2_11897 ( P1_LT_197_U119 , P1_LT_197_U79 , P1_LT_197_U115 );
nand NAND2_11898 ( P1_LT_197_U120 , P1_LT_197_U80 , P1_LT_197_U6 );
nand NAND2_11899 ( P1_LT_197_U121 , P1_U3607 , P1_LT_197_U25 );
nand NAND2_11900 ( P1_LT_197_U122 , P1_U3605 , P1_LT_197_U24 );
nand NAND2_11901 ( P1_LT_197_U123 , P1_U3610 , P1_LT_197_U32 );
nand NAND2_11902 ( P1_LT_197_U124 , P1_U3978 , P1_LT_197_U67 );
nand NAND2_11903 ( P1_LT_197_U125 , P1_U3977 , P1_LT_197_U68 );
nand NAND2_11904 ( P1_LT_197_U126 , P1_U3611 , P1_LT_197_U63 );
nand NAND2_11905 ( P1_LT_197_U127 , P1_U3473 , P1_LT_197_U42 );
nand NAND2_11906 ( P1_LT_197_U128 , P1_LT_197_U82 , P1_LT_197_U127 );
nand NAND2_11907 ( P1_LT_197_U129 , P1_U3470 , P1_LT_197_U36 );
nand NAND2_11908 ( P1_LT_197_U130 , P1_U3473 , P1_LT_197_U42 );
nand NAND2_11909 ( P1_LT_197_U131 , P1_LT_197_U83 , P1_LT_197_U9 );
nand NAND2_11910 ( P1_LT_197_U132 , P1_U3586 , P1_LT_197_U55 );
nand NAND2_11911 ( P1_LT_197_U133 , P1_U3616 , P1_LT_197_U56 );
nand NAND2_11912 ( P1_LT_197_U134 , P1_U3587 , P1_LT_197_U54 );
nand NAND2_11913 ( P1_LT_197_U135 , P1_U3588 , P1_LT_197_U35 );
nand NAND2_11914 ( P1_LT_197_U136 , P1_U3591 , P1_LT_197_U52 );
nand NAND2_11915 ( P1_LT_197_U137 , P1_U3592 , P1_LT_197_U51 );
not NOT1_11916 ( P1_LT_197_U138 , P1_LT_197_U45 );
nand NAND2_11917 ( P1_LT_197_U139 , P1_U3455 , P1_LT_197_U138 );
nand NAND2_11918 ( P1_LT_197_U140 , P1_U3606 , P1_LT_197_U139 );
nand NAND2_11919 ( P1_LT_197_U141 , P1_LT_197_U45 , P1_LT_197_U46 );
nand NAND2_11920 ( P1_LT_197_U142 , P1_U3595 , P1_LT_197_U50 );
nand NAND2_11921 ( P1_LT_197_U143 , P1_LT_197_U87 , P1_LT_197_U10 );
nand NAND2_11922 ( P1_LT_197_U144 , P1_U3488 , P1_LT_197_U58 );
nand NAND2_11923 ( P1_LT_197_U145 , P1_U3491 , P1_LT_197_U61 );
nand NAND2_11924 ( P1_LT_197_U146 , P1_LT_197_U89 , P1_LT_197_U136 );
nand NAND2_11925 ( P1_LT_197_U147 , P1_U3464 , P1_LT_197_U43 );
nand NAND3_11926 ( P1_LT_197_U148 , P1_LT_197_U147 , P1_LT_197_U146 , P1_LT_197_U9 );
nand NAND2_11927 ( P1_LT_197_U149 , P1_LT_197_U148 , P1_LT_197_U131 );
nand NAND2_11928 ( P1_LT_197_U150 , P1_U3467 , P1_LT_197_U38 );
nand NAND2_11929 ( P1_LT_197_U151 , P1_LT_197_U150 , P1_LT_197_U149 );
nand NAND2_11930 ( P1_LT_197_U152 , P1_LT_197_U90 , P1_LT_197_U151 );
nand NAND2_11931 ( P1_LT_197_U153 , P1_U3476 , P1_LT_197_U41 );
nand NAND2_11932 ( P1_LT_197_U154 , P1_LT_197_U153 , P1_LT_197_U152 );
nand NAND2_11933 ( P1_LT_197_U155 , P1_LT_197_U154 , P1_LT_197_U132 );
nand NAND2_11934 ( P1_LT_197_U156 , P1_U3479 , P1_LT_197_U39 );
nand NAND2_11935 ( P1_LT_197_U157 , P1_LT_197_U156 , P1_LT_197_U155 );
nand NAND2_11936 ( P1_LT_197_U158 , P1_LT_197_U88 , P1_LT_197_U10 );
nand NAND2_11937 ( P1_LT_197_U159 , P1_LT_197_U157 , P1_LT_197_U133 );
nand NAND2_11938 ( P1_LT_197_U160 , P1_U3482 , P1_LT_197_U40 );
nand NAND2_11939 ( P1_LT_197_U161 , P1_U3485 , P1_LT_197_U59 );
nand NAND2_11940 ( P1_LT_197_U162 , P1_LT_197_U159 , P1_LT_197_U91 );
nand NAND2_11941 ( P1_LT_197_U163 , P1_U3491 , P1_LT_197_U61 );
nand NAND2_11942 ( P1_LT_197_U164 , P1_LT_197_U94 , P1_LT_197_U163 );
nand NAND2_11943 ( P1_LT_197_U165 , P1_LT_197_U95 , P1_LT_197_U11 );
nand NAND2_11944 ( P1_LT_197_U166 , P1_U3612 , P1_LT_197_U62 );
nand NAND2_11945 ( P1_LT_197_U167 , P1_U3613 , P1_LT_197_U49 );
nand NAND2_11946 ( P1_LT_197_U168 , P1_LT_197_U162 , P1_LT_197_U97 );
nand NAND2_11947 ( P1_LT_197_U169 , P1_U3494 , P1_LT_197_U60 );
nand NAND2_11948 ( P1_LT_197_U170 , P1_LT_197_U169 , P1_LT_197_U168 );
nand NAND2_11949 ( P1_LT_197_U171 , P1_LT_197_U170 , P1_LT_197_U126 );
nand NAND2_11950 ( P1_LT_197_U172 , P1_U3497 , P1_LT_197_U34 );
nand NAND2_11951 ( P1_LT_197_U173 , P1_LT_197_U172 , P1_LT_197_U171 );
nand NAND2_11952 ( P1_LT_197_U174 , P1_U3503 , P1_LT_197_U28 );
nand NAND2_11953 ( P1_LT_197_U175 , P1_U3500 , P1_LT_197_U33 );
nand NAND2_11954 ( P1_LT_197_U176 , P1_LT_197_U78 , P1_LT_197_U6 );
nand NAND2_11955 ( P1_LT_197_U177 , P1_LT_197_U76 , P1_LT_197_U117 );
nand NAND2_11956 ( P1_LT_197_U178 , P1_LT_197_U77 , P1_LT_197_U7 );
nand NAND2_11957 ( P1_LT_197_U179 , P1_LT_197_U8 , P1_LT_197_U176 );
nand NAND3_11958 ( P1_LT_197_U180 , P1_LT_197_U173 , P1_LT_197_U123 , P1_LT_197_U8 );
nand NAND2_11959 ( P1_LT_197_U181 , P1_U3980 , P1_LT_197_U21 );
nand NAND2_11960 ( P1_LT_197_U182 , P1_U3979 , P1_LT_197_U66 );
nand NAND4_11961 ( P1_LT_197_U183 , P1_LT_197_U101 , P1_LT_197_U180 , P1_LT_197_U100 , P1_LT_197_U99 );
nand NAND2_11962 ( P1_LT_197_U184 , P1_LT_197_U102 , P1_LT_197_U124 );
nand NAND2_11963 ( P1_LT_197_U185 , P1_U3601 , P1_LT_197_U20 );
nand NAND2_11964 ( P1_LT_197_U186 , P1_U3600 , P1_LT_197_U19 );
nand NAND2_11965 ( P1_LT_197_U187 , P1_U3599 , P1_LT_197_U69 );
nand NAND3_11966 ( P1_LT_197_U188 , P1_LT_197_U184 , P1_LT_197_U183 , P1_LT_197_U103 );
nand NAND2_11967 ( P1_LT_197_U189 , P1_U3976 , P1_LT_197_U18 );
nand NAND2_11968 ( P1_LT_197_U190 , P1_LT_197_U104 , P1_LT_197_U188 );
nand NAND3_11969 ( P1_LT_197_U191 , P1_LT_197_U187 , P1_LT_197_U190 , P1_LT_197_U114 );
nand NAND2_11970 ( P1_LT_197_U192 , P1_U3975 , P1_LT_197_U17 );
not NOT1_11971 ( P1_LT_197_U193 , P1_LT_197_U71 );
or OR2_11972 ( P1_LT_197_U194 , P1_U3597 , P1_LT_197_U12 );
nand NAND2_11973 ( P1_LT_197_U195 , P1_U3974 , P1_LT_197_U71 );
nand NAND2_11974 ( P1_LT_197_U196 , P1_U3985 , P1_LT_197_U74 );
nand NAND3_11975 ( P1_LT_197_U197 , P1_LT_197_U194 , P1_LT_197_U113 , P1_LT_197_U105 );
nand NAND2_11976 ( P1_LT_197_U198 , P1_LT_197_U106 , P1_LT_197_U113 );
nand NAND2_11977 ( P1_LT_197_U199 , P1_U3983 , P1_LT_197_U15 );
nand NAND2_11978 ( P1_LT_197_U200 , P1_LT_197_U110 , P1_LT_197_U109 );
and AND2_11979 ( P1_R1360_U6 , P1_R1360_U111 , P1_R1360_U112 );
and AND2_11980 ( P1_R1360_U7 , P1_R1360_U116 , P1_R1360_U115 );
and AND2_11981 ( P1_R1360_U8 , P1_R1360_U118 , P1_R1360_U119 );
and AND2_11982 ( P1_R1360_U9 , P1_R1360_U123 , P1_R1360_U122 );
and AND5_11983 ( P1_R1360_U10 , P1_R1360_U199 , P1_R1360_U185 , P1_R1360_U186 , P1_R1360_U184 , P1_R1360_U183 );
and AND2_11984 ( P1_R1360_U11 , P1_R1360_U183 , P1_R1360_U104 );
and AND2_11985 ( P1_R1360_U12 , P1_R1360_U203 , P1_R1360_U202 );
and AND2_11986 ( P1_R1360_U13 , P1_R1360_U205 , P1_R1360_U204 );
nand NAND3_11987 ( P1_R1360_U14 , P1_R1360_U108 , P1_R1360_U200 , P1_R1360_U107 );
not NOT1_11988 ( P1_R1360_U15 , P1_U3088 );
not NOT1_11989 ( P1_R1360_U16 , P1_U3087 );
not NOT1_11990 ( P1_R1360_U17 , P1_U3121 );
not NOT1_11991 ( P1_R1360_U18 , P1_U3089 );
not NOT1_11992 ( P1_R1360_U19 , P1_U3090 );
not NOT1_11993 ( P1_R1360_U20 , P1_U3123 );
not NOT1_11994 ( P1_R1360_U21 , P1_U3122 );
not NOT1_11995 ( P1_R1360_U22 , P1_U3120 );
not NOT1_11996 ( P1_R1360_U23 , P1_U3127 );
not NOT1_11997 ( P1_R1360_U24 , P1_U3126 );
not NOT1_11998 ( P1_R1360_U25 , P1_U3097 );
not NOT1_11999 ( P1_R1360_U26 , P1_U3098 );
not NOT1_12000 ( P1_R1360_U27 , P1_U3133 );
not NOT1_12001 ( P1_R1360_U28 , P1_U3132 );
not NOT1_12002 ( P1_R1360_U29 , P1_U3103 );
not NOT1_12003 ( P1_R1360_U30 , P1_U3104 );
not NOT1_12004 ( P1_R1360_U31 , P1_U3139 );
not NOT1_12005 ( P1_R1360_U32 , P1_U3138 );
not NOT1_12006 ( P1_R1360_U33 , P1_U3109 );
not NOT1_12007 ( P1_R1360_U34 , P1_U3142 );
not NOT1_12008 ( P1_R1360_U35 , P1_U3110 );
not NOT1_12009 ( P1_R1360_U36 , P1_U3143 );
not NOT1_12010 ( P1_R1360_U37 , P1_U3112 );
not NOT1_12011 ( P1_R1360_U38 , P1_U3111 );
not NOT1_12012 ( P1_R1360_U39 , P1_U3114 );
not NOT1_12013 ( P1_R1360_U40 , P1_U3113 );
not NOT1_12014 ( P1_R1360_U41 , P1_U3116 );
not NOT1_12015 ( P1_R1360_U42 , P1_U3115 );
not NOT1_12016 ( P1_R1360_U43 , P1_U3117 );
not NOT1_12017 ( P1_R1360_U44 , P1_U3149 );
not NOT1_12018 ( P1_R1360_U45 , P1_U3148 );
not NOT1_12019 ( P1_R1360_U46 , P1_U3147 );
not NOT1_12020 ( P1_R1360_U47 , P1_U3146 );
not NOT1_12021 ( P1_R1360_U48 , P1_U3145 );
not NOT1_12022 ( P1_R1360_U49 , P1_U3144 );
not NOT1_12023 ( P1_R1360_U50 , P1_U3141 );
not NOT1_12024 ( P1_R1360_U51 , P1_U3140 );
not NOT1_12025 ( P1_R1360_U52 , P1_U3108 );
not NOT1_12026 ( P1_R1360_U53 , P1_U3106 );
not NOT1_12027 ( P1_R1360_U54 , P1_U3107 );
not NOT1_12028 ( P1_R1360_U55 , P1_U3105 );
not NOT1_12029 ( P1_R1360_U56 , P1_U3137 );
not NOT1_12030 ( P1_R1360_U57 , P1_U3136 );
not NOT1_12031 ( P1_R1360_U58 , P1_U3135 );
not NOT1_12032 ( P1_R1360_U59 , P1_U3134 );
not NOT1_12033 ( P1_R1360_U60 , P1_U3102 );
not NOT1_12034 ( P1_R1360_U61 , P1_U3101 );
not NOT1_12035 ( P1_R1360_U62 , P1_U3100 );
not NOT1_12036 ( P1_R1360_U63 , P1_U3099 );
not NOT1_12037 ( P1_R1360_U64 , P1_U3131 );
not NOT1_12038 ( P1_R1360_U65 , P1_U3130 );
not NOT1_12039 ( P1_R1360_U66 , P1_U3129 );
not NOT1_12040 ( P1_R1360_U67 , P1_U3128 );
not NOT1_12041 ( P1_R1360_U68 , P1_U3092 );
not NOT1_12042 ( P1_R1360_U69 , P1_U3091 );
not NOT1_12043 ( P1_R1360_U70 , P1_U3095 );
not NOT1_12044 ( P1_R1360_U71 , P1_U3096 );
not NOT1_12045 ( P1_R1360_U72 , P1_U3093 );
not NOT1_12046 ( P1_R1360_U73 , P1_U3094 );
not NOT1_12047 ( P1_R1360_U74 , P1_U3124 );
not NOT1_12048 ( P1_R1360_U75 , P1_U3125 );
not NOT1_12049 ( P1_R1360_U76 , P1_U3152 );
and AND2_12050 ( P1_R1360_U77 , P1_R1360_U18 , P1_U3121 );
and AND2_12051 ( P1_R1360_U78 , P1_R1360_U183 , P1_R1360_U184 );
and AND2_12052 ( P1_R1360_U79 , P1_U3142 , P1_R1360_U35 );
and AND2_12053 ( P1_R1360_U80 , P1_U3143 , P1_R1360_U38 );
and AND4_12054 ( P1_R1360_U81 , P1_R1360_U127 , P1_R1360_U126 , P1_R1360_U125 , P1_R1360_U124 );
and AND3_12055 ( P1_R1360_U82 , P1_R1360_U130 , P1_R1360_U131 , P1_R1360_U129 );
and AND2_12056 ( P1_R1360_U83 , P1_U3149 , P1_R1360_U43 );
and AND2_12057 ( P1_R1360_U84 , P1_R1360_U85 , P1_R1360_U132 );
and AND2_12058 ( P1_R1360_U85 , P1_R1360_U144 , P1_R1360_U143 );
and AND2_12059 ( P1_R1360_U86 , P1_R1360_U121 , P1_R1360_U120 );
and AND2_12060 ( P1_R1360_U87 , P1_R1360_U8 , P1_R1360_U86 );
and AND3_12061 ( P1_R1360_U88 , P1_R1360_U147 , P1_R1360_U146 , P1_R1360_U90 );
and AND2_12062 ( P1_R1360_U89 , P1_R1360_U150 , P1_R1360_U149 );
and AND2_12063 ( P1_R1360_U90 , P1_R1360_U89 , P1_R1360_U9 );
and AND2_12064 ( P1_R1360_U91 , P1_U3108 , P1_R1360_U51 );
and AND2_12065 ( P1_R1360_U92 , P1_U3107 , P1_R1360_U31 );
and AND3_12066 ( P1_R1360_U93 , P1_R1360_U152 , P1_R1360_U153 , P1_R1360_U94 );
and AND2_12067 ( P1_R1360_U94 , P1_R1360_U156 , P1_R1360_U155 );
and AND2_12068 ( P1_R1360_U95 , P1_R1360_U7 , P1_R1360_U96 );
and AND2_12069 ( P1_R1360_U96 , P1_R1360_U164 , P1_R1360_U165 );
and AND2_12070 ( P1_R1360_U97 , P1_U3102 , P1_R1360_U59 );
and AND2_12071 ( P1_R1360_U98 , P1_U3101 , P1_R1360_U27 );
and AND3_12072 ( P1_R1360_U99 , P1_R1360_U167 , P1_R1360_U169 , P1_R1360_U100 );
and AND2_12073 ( P1_R1360_U100 , P1_R1360_U171 , P1_R1360_U170 );
and AND2_12074 ( P1_R1360_U101 , P1_R1360_U179 , P1_R1360_U180 );
and AND2_12075 ( P1_R1360_U102 , P1_U3095 , P1_R1360_U23 );
and AND2_12076 ( P1_R1360_U103 , P1_U3096 , P1_R1360_U67 );
and AND5_12077 ( P1_R1360_U104 , P1_R1360_U181 , P1_R1360_U185 , P1_R1360_U186 , P1_R1360_U106 , P1_R1360_U184 );
and AND2_12078 ( P1_R1360_U105 , P1_R1360_U190 , P1_R1360_U189 );
and AND3_12079 ( P1_R1360_U106 , P1_R1360_U188 , P1_R1360_U187 , P1_R1360_U105 );
and AND3_12080 ( P1_R1360_U107 , P1_R1360_U196 , P1_R1360_U194 , P1_R1360_U195 );
and AND2_12081 ( P1_R1360_U108 , P1_R1360_U201 , P1_R1360_U13 );
not NOT1_12082 ( P1_R1360_U109 , P1_U3119 );
nand NAND2_12083 ( P1_R1360_U110 , P1_U3097 , P1_R1360_U66 );
nand NAND2_12084 ( P1_R1360_U111 , P1_U3126 , P1_R1360_U73 );
nand NAND2_12085 ( P1_R1360_U112 , P1_U3127 , P1_R1360_U70 );
nand NAND2_12086 ( P1_R1360_U113 , P1_U3098 , P1_R1360_U65 );
nand NAND2_12087 ( P1_R1360_U114 , P1_U3103 , P1_R1360_U58 );
nand NAND2_12088 ( P1_R1360_U115 , P1_U3133 , P1_R1360_U61 );
nand NAND2_12089 ( P1_R1360_U116 , P1_U3132 , P1_R1360_U62 );
nand NAND2_12090 ( P1_R1360_U117 , P1_U3104 , P1_R1360_U57 );
nand NAND2_12091 ( P1_R1360_U118 , P1_U3109 , P1_R1360_U50 );
nand NAND2_12092 ( P1_R1360_U119 , P1_U3110 , P1_R1360_U34 );
nand NAND2_12093 ( P1_R1360_U120 , P1_U3112 , P1_R1360_U49 );
nand NAND2_12094 ( P1_R1360_U121 , P1_U3111 , P1_R1360_U36 );
nand NAND2_12095 ( P1_R1360_U122 , P1_U3139 , P1_R1360_U54 );
nand NAND2_12096 ( P1_R1360_U123 , P1_U3138 , P1_R1360_U53 );
nand NAND2_12097 ( P1_R1360_U124 , P1_U3114 , P1_R1360_U47 );
nand NAND2_12098 ( P1_R1360_U125 , P1_U3113 , P1_R1360_U48 );
nand NAND2_12099 ( P1_R1360_U126 , P1_U3116 , P1_R1360_U45 );
nand NAND2_12100 ( P1_R1360_U127 , P1_U3115 , P1_R1360_U46 );
nand NAND2_12101 ( P1_R1360_U128 , P1_U3150 , P1_U3151 );
nand NAND2_12102 ( P1_R1360_U129 , P1_U3118 , P1_R1360_U128 );
or OR2_12103 ( P1_R1360_U130 , P1_U3150 , P1_U3151 );
nand NAND2_12104 ( P1_R1360_U131 , P1_U3117 , P1_R1360_U44 );
nand NAND2_12105 ( P1_R1360_U132 , P1_R1360_U82 , P1_R1360_U81 );
nand NAND2_12106 ( P1_R1360_U133 , P1_R1360_U83 , P1_R1360_U126 );
nand NAND2_12107 ( P1_R1360_U134 , P1_U3148 , P1_R1360_U41 );
nand NAND2_12108 ( P1_R1360_U135 , P1_R1360_U134 , P1_R1360_U133 );
nand NAND2_12109 ( P1_R1360_U136 , P1_R1360_U135 , P1_R1360_U127 );
nand NAND2_12110 ( P1_R1360_U137 , P1_U3147 , P1_R1360_U42 );
nand NAND2_12111 ( P1_R1360_U138 , P1_R1360_U137 , P1_R1360_U136 );
nand NAND2_12112 ( P1_R1360_U139 , P1_R1360_U138 , P1_R1360_U124 );
nand NAND2_12113 ( P1_R1360_U140 , P1_U3146 , P1_R1360_U39 );
nand NAND2_12114 ( P1_R1360_U141 , P1_R1360_U140 , P1_R1360_U139 );
nand NAND2_12115 ( P1_R1360_U142 , P1_R1360_U141 , P1_R1360_U125 );
nand NAND2_12116 ( P1_R1360_U143 , P1_U3145 , P1_R1360_U40 );
nand NAND2_12117 ( P1_R1360_U144 , P1_U3144 , P1_R1360_U37 );
nand NAND2_12118 ( P1_R1360_U145 , P1_R1360_U142 , P1_R1360_U84 );
nand NAND2_12119 ( P1_R1360_U146 , P1_R1360_U79 , P1_R1360_U118 );
nand NAND2_12120 ( P1_R1360_U147 , P1_R1360_U80 , P1_R1360_U8 );
nand NAND2_12121 ( P1_R1360_U148 , P1_R1360_U87 , P1_R1360_U145 );
nand NAND2_12122 ( P1_R1360_U149 , P1_U3141 , P1_R1360_U33 );
nand NAND2_12123 ( P1_R1360_U150 , P1_U3140 , P1_R1360_U52 );
nand NAND2_12124 ( P1_R1360_U151 , P1_R1360_U148 , P1_R1360_U88 );
nand NAND2_12125 ( P1_R1360_U152 , P1_R1360_U91 , P1_R1360_U9 );
nand NAND2_12126 ( P1_R1360_U153 , P1_U3106 , P1_R1360_U32 );
nand NAND2_12127 ( P1_R1360_U154 , P1_U3138 , P1_R1360_U53 );
nand NAND2_12128 ( P1_R1360_U155 , P1_R1360_U92 , P1_R1360_U154 );
nand NAND2_12129 ( P1_R1360_U156 , P1_U3105 , P1_R1360_U56 );
nand NAND2_12130 ( P1_R1360_U157 , P1_R1360_U151 , P1_R1360_U93 );
nand NAND2_12131 ( P1_R1360_U158 , P1_U3137 , P1_R1360_U55 );
nand NAND2_12132 ( P1_R1360_U159 , P1_R1360_U158 , P1_R1360_U157 );
nand NAND2_12133 ( P1_R1360_U160 , P1_R1360_U159 , P1_R1360_U117 );
nand NAND2_12134 ( P1_R1360_U161 , P1_U3136 , P1_R1360_U30 );
nand NAND2_12135 ( P1_R1360_U162 , P1_R1360_U161 , P1_R1360_U160 );
nand NAND2_12136 ( P1_R1360_U163 , P1_R1360_U162 , P1_R1360_U114 );
nand NAND2_12137 ( P1_R1360_U164 , P1_U3135 , P1_R1360_U29 );
nand NAND2_12138 ( P1_R1360_U165 , P1_U3134 , P1_R1360_U60 );
nand NAND2_12139 ( P1_R1360_U166 , P1_R1360_U163 , P1_R1360_U95 );
nand NAND2_12140 ( P1_R1360_U167 , P1_R1360_U97 , P1_R1360_U7 );
nand NAND2_12141 ( P1_R1360_U168 , P1_U3132 , P1_R1360_U62 );
nand NAND2_12142 ( P1_R1360_U169 , P1_R1360_U98 , P1_R1360_U168 );
nand NAND2_12143 ( P1_R1360_U170 , P1_U3100 , P1_R1360_U28 );
nand NAND2_12144 ( P1_R1360_U171 , P1_U3099 , P1_R1360_U64 );
nand NAND2_12145 ( P1_R1360_U172 , P1_R1360_U166 , P1_R1360_U99 );
nand NAND2_12146 ( P1_R1360_U173 , P1_U3131 , P1_R1360_U63 );
nand NAND2_12147 ( P1_R1360_U174 , P1_R1360_U173 , P1_R1360_U172 );
nand NAND2_12148 ( P1_R1360_U175 , P1_R1360_U174 , P1_R1360_U113 );
nand NAND2_12149 ( P1_R1360_U176 , P1_U3130 , P1_R1360_U26 );
nand NAND2_12150 ( P1_R1360_U177 , P1_R1360_U176 , P1_R1360_U175 );
nand NAND2_12151 ( P1_R1360_U178 , P1_R1360_U177 , P1_R1360_U110 );
nand NAND2_12152 ( P1_R1360_U179 , P1_U3129 , P1_R1360_U25 );
nand NAND2_12153 ( P1_R1360_U180 , P1_U3128 , P1_R1360_U71 );
nand NAND3_12154 ( P1_R1360_U181 , P1_R1360_U101 , P1_R1360_U178 , P1_R1360_U6 );
nand NAND2_12155 ( P1_R1360_U182 , P1_U3088 , P1_R1360_U22 );
nand NAND2_12156 ( P1_R1360_U183 , P1_U3089 , P1_R1360_U17 );
nand NAND2_12157 ( P1_R1360_U184 , P1_U3090 , P1_R1360_U21 );
nand NAND2_12158 ( P1_R1360_U185 , P1_U3092 , P1_R1360_U74 );
nand NAND2_12159 ( P1_R1360_U186 , P1_U3091 , P1_R1360_U20 );
nand NAND2_12160 ( P1_R1360_U187 , P1_R1360_U102 , P1_R1360_U111 );
nand NAND2_12161 ( P1_R1360_U188 , P1_R1360_U103 , P1_R1360_U6 );
nand NAND2_12162 ( P1_R1360_U189 , P1_U3093 , P1_R1360_U75 );
nand NAND2_12163 ( P1_R1360_U190 , P1_U3094 , P1_R1360_U24 );
nand NAND2_12164 ( P1_R1360_U191 , P1_U3123 , P1_R1360_U69 );
nand NAND2_12165 ( P1_R1360_U192 , P1_U3122 , P1_R1360_U19 );
nand NAND2_12166 ( P1_R1360_U193 , P1_R1360_U192 , P1_R1360_U191 );
nand NAND3_12167 ( P1_R1360_U194 , P1_R1360_U77 , P1_R1360_U12 , P1_R1360_U182 );
nand NAND4_12168 ( P1_R1360_U195 , P1_R1360_U12 , P1_R1360_U193 , P1_R1360_U78 , P1_R1360_U182 );
nand NAND3_12169 ( P1_R1360_U196 , P1_R1360_U12 , P1_R1360_U15 , P1_U3120 );
nand NAND2_12170 ( P1_R1360_U197 , P1_U3124 , P1_R1360_U68 );
nand NAND2_12171 ( P1_R1360_U198 , P1_U3125 , P1_R1360_U72 );
nand NAND2_12172 ( P1_R1360_U199 , P1_R1360_U198 , P1_R1360_U197 );
nand NAND3_12173 ( P1_R1360_U200 , P1_R1360_U12 , P1_R1360_U11 , P1_R1360_U182 );
nand NAND3_12174 ( P1_R1360_U201 , P1_R1360_U12 , P1_R1360_U10 , P1_R1360_U182 );
nand NAND2_12175 ( P1_R1360_U202 , P1_U3087 , P1_R1360_U109 );
nand NAND2_12176 ( P1_R1360_U203 , P1_U3119 , P1_R1360_U16 );
nand NAND3_12177 ( P1_R1360_U204 , P1_U3152 , P1_U3087 , P1_R1360_U109 );
nand NAND3_12178 ( P1_R1360_U205 , P1_R1360_U76 , P1_R1360_U16 , P1_U3119 );
and AND2_12179 ( P1_R1171_U4 , P1_R1171_U178 , P1_R1171_U177 );
and AND2_12180 ( P1_R1171_U5 , P1_R1171_U179 , P1_R1171_U180 );
and AND2_12181 ( P1_R1171_U6 , P1_R1171_U196 , P1_R1171_U195 );
and AND2_12182 ( P1_R1171_U7 , P1_R1171_U236 , P1_R1171_U235 );
and AND2_12183 ( P1_R1171_U8 , P1_R1171_U245 , P1_R1171_U244 );
and AND2_12184 ( P1_R1171_U9 , P1_R1171_U263 , P1_R1171_U262 );
and AND2_12185 ( P1_R1171_U10 , P1_R1171_U271 , P1_R1171_U270 );
and AND2_12186 ( P1_R1171_U11 , P1_R1171_U350 , P1_R1171_U347 );
and AND2_12187 ( P1_R1171_U12 , P1_R1171_U343 , P1_R1171_U340 );
and AND2_12188 ( P1_R1171_U13 , P1_R1171_U334 , P1_R1171_U331 );
and AND2_12189 ( P1_R1171_U14 , P1_R1171_U325 , P1_R1171_U322 );
and AND2_12190 ( P1_R1171_U15 , P1_R1171_U319 , P1_R1171_U317 );
and AND2_12191 ( P1_R1171_U16 , P1_R1171_U312 , P1_R1171_U309 );
and AND2_12192 ( P1_R1171_U17 , P1_R1171_U234 , P1_R1171_U231 );
and AND2_12193 ( P1_R1171_U18 , P1_R1171_U226 , P1_R1171_U223 );
and AND2_12194 ( P1_R1171_U19 , P1_R1171_U212 , P1_R1171_U209 );
not NOT1_12195 ( P1_R1171_U20 , P1_U3470 );
not NOT1_12196 ( P1_R1171_U21 , P1_U3071 );
not NOT1_12197 ( P1_R1171_U22 , P1_U3070 );
nand NAND2_12198 ( P1_R1171_U23 , P1_U3071 , P1_U3470 );
not NOT1_12199 ( P1_R1171_U24 , P1_U3473 );
not NOT1_12200 ( P1_R1171_U25 , P1_U3464 );
not NOT1_12201 ( P1_R1171_U26 , P1_U3060 );
not NOT1_12202 ( P1_R1171_U27 , P1_U3067 );
not NOT1_12203 ( P1_R1171_U28 , P1_U3458 );
not NOT1_12204 ( P1_R1171_U29 , P1_U3068 );
not NOT1_12205 ( P1_R1171_U30 , P1_U3450 );
not NOT1_12206 ( P1_R1171_U31 , P1_U3077 );
nand NAND2_12207 ( P1_R1171_U32 , P1_U3077 , P1_U3450 );
not NOT1_12208 ( P1_R1171_U33 , P1_U3461 );
not NOT1_12209 ( P1_R1171_U34 , P1_U3064 );
nand NAND2_12210 ( P1_R1171_U35 , P1_U3060 , P1_U3464 );
not NOT1_12211 ( P1_R1171_U36 , P1_U3467 );
not NOT1_12212 ( P1_R1171_U37 , P1_U3476 );
not NOT1_12213 ( P1_R1171_U38 , P1_U3084 );
not NOT1_12214 ( P1_R1171_U39 , P1_U3083 );
not NOT1_12215 ( P1_R1171_U40 , P1_U3479 );
nand NAND2_12216 ( P1_R1171_U41 , P1_R1171_U62 , P1_R1171_U204 );
nand NAND2_12217 ( P1_R1171_U42 , P1_R1171_U118 , P1_R1171_U192 );
nand NAND2_12218 ( P1_R1171_U43 , P1_R1171_U181 , P1_R1171_U182 );
nand NAND2_12219 ( P1_R1171_U44 , P1_U3455 , P1_U3078 );
nand NAND2_12220 ( P1_R1171_U45 , P1_R1171_U122 , P1_R1171_U218 );
nand NAND2_12221 ( P1_R1171_U46 , P1_R1171_U215 , P1_R1171_U214 );
not NOT1_12222 ( P1_R1171_U47 , P1_U3975 );
not NOT1_12223 ( P1_R1171_U48 , P1_U3053 );
not NOT1_12224 ( P1_R1171_U49 , P1_U3057 );
not NOT1_12225 ( P1_R1171_U50 , P1_U3976 );
not NOT1_12226 ( P1_R1171_U51 , P1_U3977 );
not NOT1_12227 ( P1_R1171_U52 , P1_U3058 );
not NOT1_12228 ( P1_R1171_U53 , P1_U3978 );
not NOT1_12229 ( P1_R1171_U54 , P1_U3065 );
not NOT1_12230 ( P1_R1171_U55 , P1_U3981 );
not NOT1_12231 ( P1_R1171_U56 , P1_U3075 );
not NOT1_12232 ( P1_R1171_U57 , P1_U3500 );
not NOT1_12233 ( P1_R1171_U58 , P1_U3073 );
not NOT1_12234 ( P1_R1171_U59 , P1_U3069 );
nand NAND2_12235 ( P1_R1171_U60 , P1_U3073 , P1_U3500 );
not NOT1_12236 ( P1_R1171_U61 , P1_U3503 );
nand NAND2_12237 ( P1_R1171_U62 , P1_U3084 , P1_U3476 );
not NOT1_12238 ( P1_R1171_U63 , P1_U3482 );
not NOT1_12239 ( P1_R1171_U64 , P1_U3062 );
not NOT1_12240 ( P1_R1171_U65 , P1_U3488 );
not NOT1_12241 ( P1_R1171_U66 , P1_U3072 );
not NOT1_12242 ( P1_R1171_U67 , P1_U3485 );
not NOT1_12243 ( P1_R1171_U68 , P1_U3063 );
nand NAND2_12244 ( P1_R1171_U69 , P1_U3063 , P1_U3485 );
not NOT1_12245 ( P1_R1171_U70 , P1_U3491 );
not NOT1_12246 ( P1_R1171_U71 , P1_U3080 );
not NOT1_12247 ( P1_R1171_U72 , P1_U3494 );
not NOT1_12248 ( P1_R1171_U73 , P1_U3079 );
not NOT1_12249 ( P1_R1171_U74 , P1_U3497 );
not NOT1_12250 ( P1_R1171_U75 , P1_U3074 );
not NOT1_12251 ( P1_R1171_U76 , P1_U3506 );
not NOT1_12252 ( P1_R1171_U77 , P1_U3082 );
nand NAND2_12253 ( P1_R1171_U78 , P1_U3082 , P1_U3506 );
not NOT1_12254 ( P1_R1171_U79 , P1_U3508 );
not NOT1_12255 ( P1_R1171_U80 , P1_U3081 );
nand NAND2_12256 ( P1_R1171_U81 , P1_U3081 , P1_U3508 );
not NOT1_12257 ( P1_R1171_U82 , P1_U3982 );
not NOT1_12258 ( P1_R1171_U83 , P1_U3980 );
not NOT1_12259 ( P1_R1171_U84 , P1_U3061 );
not NOT1_12260 ( P1_R1171_U85 , P1_U3979 );
not NOT1_12261 ( P1_R1171_U86 , P1_U3066 );
nand NAND2_12262 ( P1_R1171_U87 , P1_U3976 , P1_U3057 );
not NOT1_12263 ( P1_R1171_U88 , P1_U3054 );
not NOT1_12264 ( P1_R1171_U89 , P1_U3974 );
nand NAND2_12265 ( P1_R1171_U90 , P1_R1171_U305 , P1_R1171_U175 );
not NOT1_12266 ( P1_R1171_U91 , P1_U3076 );
nand NAND2_12267 ( P1_R1171_U92 , P1_R1171_U78 , P1_R1171_U314 );
nand NAND2_12268 ( P1_R1171_U93 , P1_R1171_U260 , P1_R1171_U259 );
nand NAND2_12269 ( P1_R1171_U94 , P1_R1171_U69 , P1_R1171_U336 );
nand NAND2_12270 ( P1_R1171_U95 , P1_R1171_U456 , P1_R1171_U455 );
nand NAND2_12271 ( P1_R1171_U96 , P1_R1171_U503 , P1_R1171_U502 );
nand NAND2_12272 ( P1_R1171_U97 , P1_R1171_U374 , P1_R1171_U373 );
nand NAND2_12273 ( P1_R1171_U98 , P1_R1171_U379 , P1_R1171_U378 );
nand NAND2_12274 ( P1_R1171_U99 , P1_R1171_U386 , P1_R1171_U385 );
nand NAND2_12275 ( P1_R1171_U100 , P1_R1171_U393 , P1_R1171_U392 );
nand NAND2_12276 ( P1_R1171_U101 , P1_R1171_U398 , P1_R1171_U397 );
nand NAND2_12277 ( P1_R1171_U102 , P1_R1171_U407 , P1_R1171_U406 );
nand NAND2_12278 ( P1_R1171_U103 , P1_R1171_U414 , P1_R1171_U413 );
nand NAND2_12279 ( P1_R1171_U104 , P1_R1171_U421 , P1_R1171_U420 );
nand NAND2_12280 ( P1_R1171_U105 , P1_R1171_U428 , P1_R1171_U427 );
nand NAND2_12281 ( P1_R1171_U106 , P1_R1171_U433 , P1_R1171_U432 );
nand NAND2_12282 ( P1_R1171_U107 , P1_R1171_U440 , P1_R1171_U439 );
nand NAND2_12283 ( P1_R1171_U108 , P1_R1171_U447 , P1_R1171_U446 );
nand NAND2_12284 ( P1_R1171_U109 , P1_R1171_U461 , P1_R1171_U460 );
nand NAND2_12285 ( P1_R1171_U110 , P1_R1171_U466 , P1_R1171_U465 );
nand NAND2_12286 ( P1_R1171_U111 , P1_R1171_U473 , P1_R1171_U472 );
nand NAND2_12287 ( P1_R1171_U112 , P1_R1171_U480 , P1_R1171_U479 );
nand NAND2_12288 ( P1_R1171_U113 , P1_R1171_U487 , P1_R1171_U486 );
nand NAND2_12289 ( P1_R1171_U114 , P1_R1171_U494 , P1_R1171_U493 );
nand NAND2_12290 ( P1_R1171_U115 , P1_R1171_U499 , P1_R1171_U498 );
and AND2_12291 ( P1_R1171_U116 , P1_U3458 , P1_U3068 );
and AND2_12292 ( P1_R1171_U117 , P1_R1171_U188 , P1_R1171_U186 );
and AND2_12293 ( P1_R1171_U118 , P1_R1171_U193 , P1_R1171_U191 );
and AND2_12294 ( P1_R1171_U119 , P1_R1171_U200 , P1_R1171_U199 );
and AND3_12295 ( P1_R1171_U120 , P1_R1171_U381 , P1_R1171_U380 , P1_R1171_U23 );
and AND2_12296 ( P1_R1171_U121 , P1_R1171_U211 , P1_R1171_U6 );
and AND2_12297 ( P1_R1171_U122 , P1_R1171_U219 , P1_R1171_U217 );
and AND3_12298 ( P1_R1171_U123 , P1_R1171_U388 , P1_R1171_U387 , P1_R1171_U35 );
and AND2_12299 ( P1_R1171_U124 , P1_R1171_U225 , P1_R1171_U4 );
and AND2_12300 ( P1_R1171_U125 , P1_R1171_U233 , P1_R1171_U180 );
and AND2_12301 ( P1_R1171_U126 , P1_R1171_U203 , P1_R1171_U7 );
and AND2_12302 ( P1_R1171_U127 , P1_R1171_U238 , P1_R1171_U170 );
and AND2_12303 ( P1_R1171_U128 , P1_R1171_U249 , P1_R1171_U8 );
and AND2_12304 ( P1_R1171_U129 , P1_R1171_U247 , P1_R1171_U171 );
and AND2_12305 ( P1_R1171_U130 , P1_R1171_U267 , P1_R1171_U266 );
and AND2_12306 ( P1_R1171_U131 , P1_R1171_U10 , P1_R1171_U281 );
and AND2_12307 ( P1_R1171_U132 , P1_R1171_U284 , P1_R1171_U279 );
and AND2_12308 ( P1_R1171_U133 , P1_R1171_U300 , P1_R1171_U297 );
and AND2_12309 ( P1_R1171_U134 , P1_R1171_U367 , P1_R1171_U301 );
and AND2_12310 ( P1_R1171_U135 , P1_R1171_U159 , P1_R1171_U277 );
and AND3_12311 ( P1_R1171_U136 , P1_R1171_U454 , P1_R1171_U453 , P1_R1171_U81 );
and AND3_12312 ( P1_R1171_U137 , P1_R1171_U468 , P1_R1171_U467 , P1_R1171_U60 );
and AND2_12313 ( P1_R1171_U138 , P1_R1171_U333 , P1_R1171_U9 );
and AND3_12314 ( P1_R1171_U139 , P1_R1171_U489 , P1_R1171_U488 , P1_R1171_U171 );
and AND2_12315 ( P1_R1171_U140 , P1_R1171_U342 , P1_R1171_U8 );
and AND3_12316 ( P1_R1171_U141 , P1_R1171_U501 , P1_R1171_U500 , P1_R1171_U170 );
and AND2_12317 ( P1_R1171_U142 , P1_R1171_U349 , P1_R1171_U7 );
nand NAND2_12318 ( P1_R1171_U143 , P1_R1171_U119 , P1_R1171_U201 );
nand NAND2_12319 ( P1_R1171_U144 , P1_R1171_U216 , P1_R1171_U228 );
not NOT1_12320 ( P1_R1171_U145 , P1_U3055 );
not NOT1_12321 ( P1_R1171_U146 , P1_U3985 );
and AND2_12322 ( P1_R1171_U147 , P1_R1171_U402 , P1_R1171_U401 );
nand NAND3_12323 ( P1_R1171_U148 , P1_R1171_U303 , P1_R1171_U168 , P1_R1171_U363 );
and AND2_12324 ( P1_R1171_U149 , P1_R1171_U409 , P1_R1171_U408 );
nand NAND3_12325 ( P1_R1171_U150 , P1_R1171_U369 , P1_R1171_U368 , P1_R1171_U134 );
and AND2_12326 ( P1_R1171_U151 , P1_R1171_U416 , P1_R1171_U415 );
nand NAND3_12327 ( P1_R1171_U152 , P1_R1171_U364 , P1_R1171_U298 , P1_R1171_U87 );
and AND2_12328 ( P1_R1171_U153 , P1_R1171_U423 , P1_R1171_U422 );
nand NAND2_12329 ( P1_R1171_U154 , P1_R1171_U292 , P1_R1171_U291 );
and AND2_12330 ( P1_R1171_U155 , P1_R1171_U435 , P1_R1171_U434 );
nand NAND2_12331 ( P1_R1171_U156 , P1_R1171_U288 , P1_R1171_U287 );
and AND2_12332 ( P1_R1171_U157 , P1_R1171_U442 , P1_R1171_U441 );
nand NAND2_12333 ( P1_R1171_U158 , P1_R1171_U132 , P1_R1171_U283 );
and AND2_12334 ( P1_R1171_U159 , P1_R1171_U449 , P1_R1171_U448 );
nand NAND2_12335 ( P1_R1171_U160 , P1_R1171_U44 , P1_R1171_U326 );
nand NAND2_12336 ( P1_R1171_U161 , P1_R1171_U130 , P1_R1171_U268 );
and AND2_12337 ( P1_R1171_U162 , P1_R1171_U475 , P1_R1171_U474 );
nand NAND2_12338 ( P1_R1171_U163 , P1_R1171_U256 , P1_R1171_U255 );
and AND2_12339 ( P1_R1171_U164 , P1_R1171_U482 , P1_R1171_U481 );
nand NAND2_12340 ( P1_R1171_U165 , P1_R1171_U252 , P1_R1171_U251 );
nand NAND2_12341 ( P1_R1171_U166 , P1_R1171_U242 , P1_R1171_U241 );
nand NAND2_12342 ( P1_R1171_U167 , P1_R1171_U366 , P1_R1171_U365 );
nand NAND2_12343 ( P1_R1171_U168 , P1_U3054 , P1_R1171_U150 );
not NOT1_12344 ( P1_R1171_U169 , P1_R1171_U35 );
nand NAND2_12345 ( P1_R1171_U170 , P1_U3479 , P1_U3083 );
nand NAND2_12346 ( P1_R1171_U171 , P1_U3072 , P1_U3488 );
nand NAND2_12347 ( P1_R1171_U172 , P1_U3058 , P1_U3977 );
not NOT1_12348 ( P1_R1171_U173 , P1_R1171_U69 );
not NOT1_12349 ( P1_R1171_U174 , P1_R1171_U78 );
nand NAND2_12350 ( P1_R1171_U175 , P1_U3065 , P1_U3978 );
not NOT1_12351 ( P1_R1171_U176 , P1_R1171_U62 );
or OR2_12352 ( P1_R1171_U177 , P1_U3067 , P1_U3467 );
or OR2_12353 ( P1_R1171_U178 , P1_U3060 , P1_U3464 );
or OR2_12354 ( P1_R1171_U179 , P1_U3461 , P1_U3064 );
or OR2_12355 ( P1_R1171_U180 , P1_U3458 , P1_U3068 );
not NOT1_12356 ( P1_R1171_U181 , P1_R1171_U32 );
or OR2_12357 ( P1_R1171_U182 , P1_U3455 , P1_U3078 );
not NOT1_12358 ( P1_R1171_U183 , P1_R1171_U43 );
not NOT1_12359 ( P1_R1171_U184 , P1_R1171_U44 );
nand NAND2_12360 ( P1_R1171_U185 , P1_R1171_U43 , P1_R1171_U44 );
nand NAND2_12361 ( P1_R1171_U186 , P1_R1171_U116 , P1_R1171_U179 );
nand NAND2_12362 ( P1_R1171_U187 , P1_R1171_U5 , P1_R1171_U185 );
nand NAND2_12363 ( P1_R1171_U188 , P1_U3064 , P1_U3461 );
nand NAND2_12364 ( P1_R1171_U189 , P1_R1171_U117 , P1_R1171_U187 );
nand NAND2_12365 ( P1_R1171_U190 , P1_R1171_U36 , P1_R1171_U35 );
nand NAND2_12366 ( P1_R1171_U191 , P1_U3067 , P1_R1171_U190 );
nand NAND2_12367 ( P1_R1171_U192 , P1_R1171_U4 , P1_R1171_U189 );
nand NAND2_12368 ( P1_R1171_U193 , P1_U3467 , P1_R1171_U169 );
not NOT1_12369 ( P1_R1171_U194 , P1_R1171_U42 );
or OR2_12370 ( P1_R1171_U195 , P1_U3070 , P1_U3473 );
or OR2_12371 ( P1_R1171_U196 , P1_U3071 , P1_U3470 );
not NOT1_12372 ( P1_R1171_U197 , P1_R1171_U23 );
nand NAND2_12373 ( P1_R1171_U198 , P1_R1171_U24 , P1_R1171_U23 );
nand NAND2_12374 ( P1_R1171_U199 , P1_U3070 , P1_R1171_U198 );
nand NAND2_12375 ( P1_R1171_U200 , P1_U3473 , P1_R1171_U197 );
nand NAND2_12376 ( P1_R1171_U201 , P1_R1171_U6 , P1_R1171_U42 );
not NOT1_12377 ( P1_R1171_U202 , P1_R1171_U143 );
or OR2_12378 ( P1_R1171_U203 , P1_U3476 , P1_U3084 );
nand NAND2_12379 ( P1_R1171_U204 , P1_R1171_U203 , P1_R1171_U143 );
not NOT1_12380 ( P1_R1171_U205 , P1_R1171_U41 );
or OR2_12381 ( P1_R1171_U206 , P1_U3083 , P1_U3479 );
or OR2_12382 ( P1_R1171_U207 , P1_U3470 , P1_U3071 );
nand NAND2_12383 ( P1_R1171_U208 , P1_R1171_U207 , P1_R1171_U42 );
nand NAND2_12384 ( P1_R1171_U209 , P1_R1171_U120 , P1_R1171_U208 );
nand NAND2_12385 ( P1_R1171_U210 , P1_R1171_U194 , P1_R1171_U23 );
nand NAND2_12386 ( P1_R1171_U211 , P1_U3473 , P1_U3070 );
nand NAND2_12387 ( P1_R1171_U212 , P1_R1171_U121 , P1_R1171_U210 );
or OR2_12388 ( P1_R1171_U213 , P1_U3071 , P1_U3470 );
nand NAND2_12389 ( P1_R1171_U214 , P1_R1171_U184 , P1_R1171_U180 );
nand NAND2_12390 ( P1_R1171_U215 , P1_U3068 , P1_U3458 );
not NOT1_12391 ( P1_R1171_U216 , P1_R1171_U46 );
nand NAND2_12392 ( P1_R1171_U217 , P1_R1171_U183 , P1_R1171_U5 );
nand NAND2_12393 ( P1_R1171_U218 , P1_R1171_U46 , P1_R1171_U179 );
nand NAND2_12394 ( P1_R1171_U219 , P1_U3064 , P1_U3461 );
not NOT1_12395 ( P1_R1171_U220 , P1_R1171_U45 );
or OR2_12396 ( P1_R1171_U221 , P1_U3464 , P1_U3060 );
nand NAND2_12397 ( P1_R1171_U222 , P1_R1171_U221 , P1_R1171_U45 );
nand NAND2_12398 ( P1_R1171_U223 , P1_R1171_U123 , P1_R1171_U222 );
nand NAND2_12399 ( P1_R1171_U224 , P1_R1171_U220 , P1_R1171_U35 );
nand NAND2_12400 ( P1_R1171_U225 , P1_U3467 , P1_U3067 );
nand NAND2_12401 ( P1_R1171_U226 , P1_R1171_U124 , P1_R1171_U224 );
or OR2_12402 ( P1_R1171_U227 , P1_U3060 , P1_U3464 );
nand NAND2_12403 ( P1_R1171_U228 , P1_R1171_U183 , P1_R1171_U180 );
not NOT1_12404 ( P1_R1171_U229 , P1_R1171_U144 );
nand NAND2_12405 ( P1_R1171_U230 , P1_U3064 , P1_U3461 );
nand NAND4_12406 ( P1_R1171_U231 , P1_R1171_U400 , P1_R1171_U399 , P1_R1171_U44 , P1_R1171_U43 );
nand NAND2_12407 ( P1_R1171_U232 , P1_R1171_U44 , P1_R1171_U43 );
nand NAND2_12408 ( P1_R1171_U233 , P1_U3068 , P1_U3458 );
nand NAND2_12409 ( P1_R1171_U234 , P1_R1171_U125 , P1_R1171_U232 );
or OR2_12410 ( P1_R1171_U235 , P1_U3083 , P1_U3479 );
or OR2_12411 ( P1_R1171_U236 , P1_U3062 , P1_U3482 );
nand NAND2_12412 ( P1_R1171_U237 , P1_R1171_U176 , P1_R1171_U7 );
nand NAND2_12413 ( P1_R1171_U238 , P1_U3062 , P1_U3482 );
nand NAND2_12414 ( P1_R1171_U239 , P1_R1171_U127 , P1_R1171_U237 );
or OR2_12415 ( P1_R1171_U240 , P1_U3482 , P1_U3062 );
nand NAND2_12416 ( P1_R1171_U241 , P1_R1171_U126 , P1_R1171_U143 );
nand NAND2_12417 ( P1_R1171_U242 , P1_R1171_U240 , P1_R1171_U239 );
not NOT1_12418 ( P1_R1171_U243 , P1_R1171_U166 );
or OR2_12419 ( P1_R1171_U244 , P1_U3080 , P1_U3491 );
or OR2_12420 ( P1_R1171_U245 , P1_U3072 , P1_U3488 );
nand NAND2_12421 ( P1_R1171_U246 , P1_R1171_U173 , P1_R1171_U8 );
nand NAND2_12422 ( P1_R1171_U247 , P1_U3080 , P1_U3491 );
nand NAND2_12423 ( P1_R1171_U248 , P1_R1171_U129 , P1_R1171_U246 );
or OR2_12424 ( P1_R1171_U249 , P1_U3485 , P1_U3063 );
or OR2_12425 ( P1_R1171_U250 , P1_U3491 , P1_U3080 );
nand NAND2_12426 ( P1_R1171_U251 , P1_R1171_U128 , P1_R1171_U166 );
nand NAND2_12427 ( P1_R1171_U252 , P1_R1171_U250 , P1_R1171_U248 );
not NOT1_12428 ( P1_R1171_U253 , P1_R1171_U165 );
or OR2_12429 ( P1_R1171_U254 , P1_U3494 , P1_U3079 );
nand NAND2_12430 ( P1_R1171_U255 , P1_R1171_U254 , P1_R1171_U165 );
nand NAND2_12431 ( P1_R1171_U256 , P1_U3079 , P1_U3494 );
not NOT1_12432 ( P1_R1171_U257 , P1_R1171_U163 );
or OR2_12433 ( P1_R1171_U258 , P1_U3497 , P1_U3074 );
nand NAND2_12434 ( P1_R1171_U259 , P1_R1171_U258 , P1_R1171_U163 );
nand NAND2_12435 ( P1_R1171_U260 , P1_U3074 , P1_U3497 );
not NOT1_12436 ( P1_R1171_U261 , P1_R1171_U93 );
or OR2_12437 ( P1_R1171_U262 , P1_U3069 , P1_U3503 );
or OR2_12438 ( P1_R1171_U263 , P1_U3073 , P1_U3500 );
not NOT1_12439 ( P1_R1171_U264 , P1_R1171_U60 );
nand NAND2_12440 ( P1_R1171_U265 , P1_R1171_U61 , P1_R1171_U60 );
nand NAND2_12441 ( P1_R1171_U266 , P1_U3069 , P1_R1171_U265 );
nand NAND2_12442 ( P1_R1171_U267 , P1_U3503 , P1_R1171_U264 );
nand NAND2_12443 ( P1_R1171_U268 , P1_R1171_U9 , P1_R1171_U93 );
not NOT1_12444 ( P1_R1171_U269 , P1_R1171_U161 );
or OR2_12445 ( P1_R1171_U270 , P1_U3076 , P1_U3982 );
or OR2_12446 ( P1_R1171_U271 , P1_U3081 , P1_U3508 );
or OR2_12447 ( P1_R1171_U272 , P1_U3075 , P1_U3981 );
not NOT1_12448 ( P1_R1171_U273 , P1_R1171_U81 );
nand NAND2_12449 ( P1_R1171_U274 , P1_U3982 , P1_R1171_U273 );
nand NAND2_12450 ( P1_R1171_U275 , P1_R1171_U274 , P1_R1171_U91 );
nand NAND2_12451 ( P1_R1171_U276 , P1_R1171_U81 , P1_R1171_U82 );
nand NAND2_12452 ( P1_R1171_U277 , P1_R1171_U276 , P1_R1171_U275 );
nand NAND2_12453 ( P1_R1171_U278 , P1_R1171_U174 , P1_R1171_U10 );
nand NAND2_12454 ( P1_R1171_U279 , P1_U3075 , P1_U3981 );
nand NAND2_12455 ( P1_R1171_U280 , P1_R1171_U277 , P1_R1171_U278 );
or OR2_12456 ( P1_R1171_U281 , P1_U3506 , P1_U3082 );
or OR2_12457 ( P1_R1171_U282 , P1_U3981 , P1_U3075 );
nand NAND3_12458 ( P1_R1171_U283 , P1_R1171_U272 , P1_R1171_U161 , P1_R1171_U131 );
nand NAND2_12459 ( P1_R1171_U284 , P1_R1171_U282 , P1_R1171_U280 );
not NOT1_12460 ( P1_R1171_U285 , P1_R1171_U158 );
or OR2_12461 ( P1_R1171_U286 , P1_U3980 , P1_U3061 );
nand NAND2_12462 ( P1_R1171_U287 , P1_R1171_U286 , P1_R1171_U158 );
nand NAND2_12463 ( P1_R1171_U288 , P1_U3061 , P1_U3980 );
not NOT1_12464 ( P1_R1171_U289 , P1_R1171_U156 );
or OR2_12465 ( P1_R1171_U290 , P1_U3979 , P1_U3066 );
nand NAND2_12466 ( P1_R1171_U291 , P1_R1171_U290 , P1_R1171_U156 );
nand NAND2_12467 ( P1_R1171_U292 , P1_U3066 , P1_U3979 );
not NOT1_12468 ( P1_R1171_U293 , P1_R1171_U154 );
or OR2_12469 ( P1_R1171_U294 , P1_U3058 , P1_U3977 );
nand NAND2_12470 ( P1_R1171_U295 , P1_R1171_U175 , P1_R1171_U172 );
not NOT1_12471 ( P1_R1171_U296 , P1_R1171_U87 );
or OR2_12472 ( P1_R1171_U297 , P1_U3978 , P1_U3065 );
nand NAND3_12473 ( P1_R1171_U298 , P1_R1171_U154 , P1_R1171_U297 , P1_R1171_U167 );
not NOT1_12474 ( P1_R1171_U299 , P1_R1171_U152 );
or OR2_12475 ( P1_R1171_U300 , P1_U3975 , P1_U3053 );
nand NAND2_12476 ( P1_R1171_U301 , P1_U3053 , P1_U3975 );
not NOT1_12477 ( P1_R1171_U302 , P1_R1171_U150 );
nand NAND2_12478 ( P1_R1171_U303 , P1_U3974 , P1_R1171_U150 );
not NOT1_12479 ( P1_R1171_U304 , P1_R1171_U148 );
nand NAND2_12480 ( P1_R1171_U305 , P1_R1171_U297 , P1_R1171_U154 );
not NOT1_12481 ( P1_R1171_U306 , P1_R1171_U90 );
or OR2_12482 ( P1_R1171_U307 , P1_U3977 , P1_U3058 );
nand NAND2_12483 ( P1_R1171_U308 , P1_R1171_U307 , P1_R1171_U90 );
nand NAND3_12484 ( P1_R1171_U309 , P1_R1171_U308 , P1_R1171_U172 , P1_R1171_U153 );
nand NAND2_12485 ( P1_R1171_U310 , P1_R1171_U306 , P1_R1171_U172 );
nand NAND2_12486 ( P1_R1171_U311 , P1_U3976 , P1_U3057 );
nand NAND3_12487 ( P1_R1171_U312 , P1_R1171_U310 , P1_R1171_U311 , P1_R1171_U167 );
or OR2_12488 ( P1_R1171_U313 , P1_U3058 , P1_U3977 );
nand NAND2_12489 ( P1_R1171_U314 , P1_R1171_U281 , P1_R1171_U161 );
not NOT1_12490 ( P1_R1171_U315 , P1_R1171_U92 );
nand NAND2_12491 ( P1_R1171_U316 , P1_R1171_U10 , P1_R1171_U92 );
nand NAND2_12492 ( P1_R1171_U317 , P1_R1171_U135 , P1_R1171_U316 );
nand NAND2_12493 ( P1_R1171_U318 , P1_R1171_U316 , P1_R1171_U277 );
nand NAND2_12494 ( P1_R1171_U319 , P1_R1171_U452 , P1_R1171_U318 );
or OR2_12495 ( P1_R1171_U320 , P1_U3508 , P1_U3081 );
nand NAND2_12496 ( P1_R1171_U321 , P1_R1171_U320 , P1_R1171_U92 );
nand NAND2_12497 ( P1_R1171_U322 , P1_R1171_U136 , P1_R1171_U321 );
nand NAND2_12498 ( P1_R1171_U323 , P1_R1171_U315 , P1_R1171_U81 );
nand NAND2_12499 ( P1_R1171_U324 , P1_U3076 , P1_U3982 );
nand NAND3_12500 ( P1_R1171_U325 , P1_R1171_U324 , P1_R1171_U323 , P1_R1171_U10 );
or OR2_12501 ( P1_R1171_U326 , P1_U3455 , P1_U3078 );
not NOT1_12502 ( P1_R1171_U327 , P1_R1171_U160 );
or OR2_12503 ( P1_R1171_U328 , P1_U3081 , P1_U3508 );
or OR2_12504 ( P1_R1171_U329 , P1_U3500 , P1_U3073 );
nand NAND2_12505 ( P1_R1171_U330 , P1_R1171_U329 , P1_R1171_U93 );
nand NAND2_12506 ( P1_R1171_U331 , P1_R1171_U137 , P1_R1171_U330 );
nand NAND2_12507 ( P1_R1171_U332 , P1_R1171_U261 , P1_R1171_U60 );
nand NAND2_12508 ( P1_R1171_U333 , P1_U3503 , P1_U3069 );
nand NAND2_12509 ( P1_R1171_U334 , P1_R1171_U138 , P1_R1171_U332 );
or OR2_12510 ( P1_R1171_U335 , P1_U3073 , P1_U3500 );
nand NAND2_12511 ( P1_R1171_U336 , P1_R1171_U249 , P1_R1171_U166 );
not NOT1_12512 ( P1_R1171_U337 , P1_R1171_U94 );
or OR2_12513 ( P1_R1171_U338 , P1_U3488 , P1_U3072 );
nand NAND2_12514 ( P1_R1171_U339 , P1_R1171_U338 , P1_R1171_U94 );
nand NAND2_12515 ( P1_R1171_U340 , P1_R1171_U139 , P1_R1171_U339 );
nand NAND2_12516 ( P1_R1171_U341 , P1_R1171_U337 , P1_R1171_U171 );
nand NAND2_12517 ( P1_R1171_U342 , P1_U3080 , P1_U3491 );
nand NAND2_12518 ( P1_R1171_U343 , P1_R1171_U140 , P1_R1171_U341 );
or OR2_12519 ( P1_R1171_U344 , P1_U3072 , P1_U3488 );
or OR2_12520 ( P1_R1171_U345 , P1_U3479 , P1_U3083 );
nand NAND2_12521 ( P1_R1171_U346 , P1_R1171_U345 , P1_R1171_U41 );
nand NAND2_12522 ( P1_R1171_U347 , P1_R1171_U141 , P1_R1171_U346 );
nand NAND2_12523 ( P1_R1171_U348 , P1_R1171_U205 , P1_R1171_U170 );
nand NAND2_12524 ( P1_R1171_U349 , P1_U3062 , P1_U3482 );
nand NAND2_12525 ( P1_R1171_U350 , P1_R1171_U142 , P1_R1171_U348 );
nand NAND2_12526 ( P1_R1171_U351 , P1_R1171_U206 , P1_R1171_U170 );
nand NAND2_12527 ( P1_R1171_U352 , P1_R1171_U203 , P1_R1171_U62 );
nand NAND2_12528 ( P1_R1171_U353 , P1_R1171_U213 , P1_R1171_U23 );
nand NAND2_12529 ( P1_R1171_U354 , P1_R1171_U227 , P1_R1171_U35 );
nand NAND2_12530 ( P1_R1171_U355 , P1_R1171_U230 , P1_R1171_U179 );
nand NAND2_12531 ( P1_R1171_U356 , P1_R1171_U313 , P1_R1171_U172 );
nand NAND2_12532 ( P1_R1171_U357 , P1_R1171_U297 , P1_R1171_U175 );
nand NAND2_12533 ( P1_R1171_U358 , P1_R1171_U328 , P1_R1171_U81 );
nand NAND2_12534 ( P1_R1171_U359 , P1_R1171_U281 , P1_R1171_U78 );
nand NAND2_12535 ( P1_R1171_U360 , P1_R1171_U335 , P1_R1171_U60 );
nand NAND2_12536 ( P1_R1171_U361 , P1_R1171_U344 , P1_R1171_U171 );
nand NAND2_12537 ( P1_R1171_U362 , P1_R1171_U249 , P1_R1171_U69 );
nand NAND2_12538 ( P1_R1171_U363 , P1_U3974 , P1_U3054 );
nand NAND2_12539 ( P1_R1171_U364 , P1_R1171_U295 , P1_R1171_U167 );
nand NAND2_12540 ( P1_R1171_U365 , P1_U3057 , P1_R1171_U294 );
nand NAND2_12541 ( P1_R1171_U366 , P1_U3976 , P1_R1171_U294 );
nand NAND3_12542 ( P1_R1171_U367 , P1_R1171_U295 , P1_R1171_U167 , P1_R1171_U300 );
nand NAND3_12543 ( P1_R1171_U368 , P1_R1171_U154 , P1_R1171_U167 , P1_R1171_U133 );
nand NAND2_12544 ( P1_R1171_U369 , P1_R1171_U296 , P1_R1171_U300 );
nand NAND2_12545 ( P1_R1171_U370 , P1_U3083 , P1_R1171_U40 );
nand NAND2_12546 ( P1_R1171_U371 , P1_U3479 , P1_R1171_U39 );
nand NAND2_12547 ( P1_R1171_U372 , P1_R1171_U371 , P1_R1171_U370 );
nand NAND2_12548 ( P1_R1171_U373 , P1_R1171_U351 , P1_R1171_U41 );
nand NAND2_12549 ( P1_R1171_U374 , P1_R1171_U372 , P1_R1171_U205 );
nand NAND2_12550 ( P1_R1171_U375 , P1_U3084 , P1_R1171_U37 );
nand NAND2_12551 ( P1_R1171_U376 , P1_U3476 , P1_R1171_U38 );
nand NAND2_12552 ( P1_R1171_U377 , P1_R1171_U376 , P1_R1171_U375 );
nand NAND2_12553 ( P1_R1171_U378 , P1_R1171_U352 , P1_R1171_U143 );
nand NAND2_12554 ( P1_R1171_U379 , P1_R1171_U202 , P1_R1171_U377 );
nand NAND2_12555 ( P1_R1171_U380 , P1_U3070 , P1_R1171_U24 );
nand NAND2_12556 ( P1_R1171_U381 , P1_U3473 , P1_R1171_U22 );
nand NAND2_12557 ( P1_R1171_U382 , P1_U3071 , P1_R1171_U20 );
nand NAND2_12558 ( P1_R1171_U383 , P1_U3470 , P1_R1171_U21 );
nand NAND2_12559 ( P1_R1171_U384 , P1_R1171_U383 , P1_R1171_U382 );
nand NAND2_12560 ( P1_R1171_U385 , P1_R1171_U353 , P1_R1171_U42 );
nand NAND2_12561 ( P1_R1171_U386 , P1_R1171_U384 , P1_R1171_U194 );
nand NAND2_12562 ( P1_R1171_U387 , P1_U3067 , P1_R1171_U36 );
nand NAND2_12563 ( P1_R1171_U388 , P1_U3467 , P1_R1171_U27 );
nand NAND2_12564 ( P1_R1171_U389 , P1_U3060 , P1_R1171_U25 );
nand NAND2_12565 ( P1_R1171_U390 , P1_U3464 , P1_R1171_U26 );
nand NAND2_12566 ( P1_R1171_U391 , P1_R1171_U390 , P1_R1171_U389 );
nand NAND2_12567 ( P1_R1171_U392 , P1_R1171_U354 , P1_R1171_U45 );
nand NAND2_12568 ( P1_R1171_U393 , P1_R1171_U391 , P1_R1171_U220 );
nand NAND2_12569 ( P1_R1171_U394 , P1_U3064 , P1_R1171_U33 );
nand NAND2_12570 ( P1_R1171_U395 , P1_U3461 , P1_R1171_U34 );
nand NAND2_12571 ( P1_R1171_U396 , P1_R1171_U395 , P1_R1171_U394 );
nand NAND2_12572 ( P1_R1171_U397 , P1_R1171_U355 , P1_R1171_U144 );
nand NAND2_12573 ( P1_R1171_U398 , P1_R1171_U229 , P1_R1171_U396 );
nand NAND2_12574 ( P1_R1171_U399 , P1_U3068 , P1_R1171_U28 );
nand NAND2_12575 ( P1_R1171_U400 , P1_U3458 , P1_R1171_U29 );
nand NAND2_12576 ( P1_R1171_U401 , P1_U3055 , P1_R1171_U146 );
nand NAND2_12577 ( P1_R1171_U402 , P1_U3985 , P1_R1171_U145 );
nand NAND2_12578 ( P1_R1171_U403 , P1_U3055 , P1_R1171_U146 );
nand NAND2_12579 ( P1_R1171_U404 , P1_U3985 , P1_R1171_U145 );
nand NAND2_12580 ( P1_R1171_U405 , P1_R1171_U404 , P1_R1171_U403 );
nand NAND2_12581 ( P1_R1171_U406 , P1_R1171_U147 , P1_R1171_U148 );
nand NAND2_12582 ( P1_R1171_U407 , P1_R1171_U304 , P1_R1171_U405 );
nand NAND2_12583 ( P1_R1171_U408 , P1_U3054 , P1_R1171_U89 );
nand NAND2_12584 ( P1_R1171_U409 , P1_U3974 , P1_R1171_U88 );
nand NAND2_12585 ( P1_R1171_U410 , P1_U3054 , P1_R1171_U89 );
nand NAND2_12586 ( P1_R1171_U411 , P1_U3974 , P1_R1171_U88 );
nand NAND2_12587 ( P1_R1171_U412 , P1_R1171_U411 , P1_R1171_U410 );
nand NAND2_12588 ( P1_R1171_U413 , P1_R1171_U149 , P1_R1171_U150 );
nand NAND2_12589 ( P1_R1171_U414 , P1_R1171_U302 , P1_R1171_U412 );
nand NAND2_12590 ( P1_R1171_U415 , P1_U3053 , P1_R1171_U47 );
nand NAND2_12591 ( P1_R1171_U416 , P1_U3975 , P1_R1171_U48 );
nand NAND2_12592 ( P1_R1171_U417 , P1_U3053 , P1_R1171_U47 );
nand NAND2_12593 ( P1_R1171_U418 , P1_U3975 , P1_R1171_U48 );
nand NAND2_12594 ( P1_R1171_U419 , P1_R1171_U418 , P1_R1171_U417 );
nand NAND2_12595 ( P1_R1171_U420 , P1_R1171_U151 , P1_R1171_U152 );
nand NAND2_12596 ( P1_R1171_U421 , P1_R1171_U299 , P1_R1171_U419 );
nand NAND2_12597 ( P1_R1171_U422 , P1_U3057 , P1_R1171_U50 );
nand NAND2_12598 ( P1_R1171_U423 , P1_U3976 , P1_R1171_U49 );
nand NAND2_12599 ( P1_R1171_U424 , P1_U3058 , P1_R1171_U51 );
nand NAND2_12600 ( P1_R1171_U425 , P1_U3977 , P1_R1171_U52 );
nand NAND2_12601 ( P1_R1171_U426 , P1_R1171_U425 , P1_R1171_U424 );
nand NAND2_12602 ( P1_R1171_U427 , P1_R1171_U356 , P1_R1171_U90 );
nand NAND2_12603 ( P1_R1171_U428 , P1_R1171_U426 , P1_R1171_U306 );
nand NAND2_12604 ( P1_R1171_U429 , P1_U3065 , P1_R1171_U53 );
nand NAND2_12605 ( P1_R1171_U430 , P1_U3978 , P1_R1171_U54 );
nand NAND2_12606 ( P1_R1171_U431 , P1_R1171_U430 , P1_R1171_U429 );
nand NAND2_12607 ( P1_R1171_U432 , P1_R1171_U357 , P1_R1171_U154 );
nand NAND2_12608 ( P1_R1171_U433 , P1_R1171_U293 , P1_R1171_U431 );
nand NAND2_12609 ( P1_R1171_U434 , P1_U3066 , P1_R1171_U85 );
nand NAND2_12610 ( P1_R1171_U435 , P1_U3979 , P1_R1171_U86 );
nand NAND2_12611 ( P1_R1171_U436 , P1_U3066 , P1_R1171_U85 );
nand NAND2_12612 ( P1_R1171_U437 , P1_U3979 , P1_R1171_U86 );
nand NAND2_12613 ( P1_R1171_U438 , P1_R1171_U437 , P1_R1171_U436 );
nand NAND2_12614 ( P1_R1171_U439 , P1_R1171_U155 , P1_R1171_U156 );
nand NAND2_12615 ( P1_R1171_U440 , P1_R1171_U289 , P1_R1171_U438 );
nand NAND2_12616 ( P1_R1171_U441 , P1_U3061 , P1_R1171_U83 );
nand NAND2_12617 ( P1_R1171_U442 , P1_U3980 , P1_R1171_U84 );
nand NAND2_12618 ( P1_R1171_U443 , P1_U3061 , P1_R1171_U83 );
nand NAND2_12619 ( P1_R1171_U444 , P1_U3980 , P1_R1171_U84 );
nand NAND2_12620 ( P1_R1171_U445 , P1_R1171_U444 , P1_R1171_U443 );
nand NAND2_12621 ( P1_R1171_U446 , P1_R1171_U157 , P1_R1171_U158 );
nand NAND2_12622 ( P1_R1171_U447 , P1_R1171_U285 , P1_R1171_U445 );
nand NAND2_12623 ( P1_R1171_U448 , P1_U3075 , P1_R1171_U55 );
nand NAND2_12624 ( P1_R1171_U449 , P1_U3981 , P1_R1171_U56 );
nand NAND2_12625 ( P1_R1171_U450 , P1_U3075 , P1_R1171_U55 );
nand NAND2_12626 ( P1_R1171_U451 , P1_U3981 , P1_R1171_U56 );
nand NAND2_12627 ( P1_R1171_U452 , P1_R1171_U451 , P1_R1171_U450 );
nand NAND2_12628 ( P1_R1171_U453 , P1_U3076 , P1_R1171_U82 );
nand NAND2_12629 ( P1_R1171_U454 , P1_U3982 , P1_R1171_U91 );
nand NAND2_12630 ( P1_R1171_U455 , P1_R1171_U181 , P1_R1171_U160 );
nand NAND2_12631 ( P1_R1171_U456 , P1_R1171_U327 , P1_R1171_U32 );
nand NAND2_12632 ( P1_R1171_U457 , P1_U3081 , P1_R1171_U79 );
nand NAND2_12633 ( P1_R1171_U458 , P1_U3508 , P1_R1171_U80 );
nand NAND2_12634 ( P1_R1171_U459 , P1_R1171_U458 , P1_R1171_U457 );
nand NAND2_12635 ( P1_R1171_U460 , P1_R1171_U358 , P1_R1171_U92 );
nand NAND2_12636 ( P1_R1171_U461 , P1_R1171_U459 , P1_R1171_U315 );
nand NAND2_12637 ( P1_R1171_U462 , P1_U3082 , P1_R1171_U76 );
nand NAND2_12638 ( P1_R1171_U463 , P1_U3506 , P1_R1171_U77 );
nand NAND2_12639 ( P1_R1171_U464 , P1_R1171_U463 , P1_R1171_U462 );
nand NAND2_12640 ( P1_R1171_U465 , P1_R1171_U359 , P1_R1171_U161 );
nand NAND2_12641 ( P1_R1171_U466 , P1_R1171_U269 , P1_R1171_U464 );
nand NAND2_12642 ( P1_R1171_U467 , P1_U3069 , P1_R1171_U61 );
nand NAND2_12643 ( P1_R1171_U468 , P1_U3503 , P1_R1171_U59 );
nand NAND2_12644 ( P1_R1171_U469 , P1_U3073 , P1_R1171_U57 );
nand NAND2_12645 ( P1_R1171_U470 , P1_U3500 , P1_R1171_U58 );
nand NAND2_12646 ( P1_R1171_U471 , P1_R1171_U470 , P1_R1171_U469 );
nand NAND2_12647 ( P1_R1171_U472 , P1_R1171_U360 , P1_R1171_U93 );
nand NAND2_12648 ( P1_R1171_U473 , P1_R1171_U471 , P1_R1171_U261 );
nand NAND2_12649 ( P1_R1171_U474 , P1_U3074 , P1_R1171_U74 );
nand NAND2_12650 ( P1_R1171_U475 , P1_U3497 , P1_R1171_U75 );
nand NAND2_12651 ( P1_R1171_U476 , P1_U3074 , P1_R1171_U74 );
nand NAND2_12652 ( P1_R1171_U477 , P1_U3497 , P1_R1171_U75 );
nand NAND2_12653 ( P1_R1171_U478 , P1_R1171_U477 , P1_R1171_U476 );
nand NAND2_12654 ( P1_R1171_U479 , P1_R1171_U162 , P1_R1171_U163 );
nand NAND2_12655 ( P1_R1171_U480 , P1_R1171_U257 , P1_R1171_U478 );
nand NAND2_12656 ( P1_R1171_U481 , P1_U3079 , P1_R1171_U72 );
nand NAND2_12657 ( P1_R1171_U482 , P1_U3494 , P1_R1171_U73 );
nand NAND2_12658 ( P1_R1171_U483 , P1_U3079 , P1_R1171_U72 );
nand NAND2_12659 ( P1_R1171_U484 , P1_U3494 , P1_R1171_U73 );
nand NAND2_12660 ( P1_R1171_U485 , P1_R1171_U484 , P1_R1171_U483 );
nand NAND2_12661 ( P1_R1171_U486 , P1_R1171_U164 , P1_R1171_U165 );
nand NAND2_12662 ( P1_R1171_U487 , P1_R1171_U253 , P1_R1171_U485 );
nand NAND2_12663 ( P1_R1171_U488 , P1_U3080 , P1_R1171_U70 );
nand NAND2_12664 ( P1_R1171_U489 , P1_U3491 , P1_R1171_U71 );
nand NAND2_12665 ( P1_R1171_U490 , P1_U3072 , P1_R1171_U65 );
nand NAND2_12666 ( P1_R1171_U491 , P1_U3488 , P1_R1171_U66 );
nand NAND2_12667 ( P1_R1171_U492 , P1_R1171_U491 , P1_R1171_U490 );
nand NAND2_12668 ( P1_R1171_U493 , P1_R1171_U361 , P1_R1171_U94 );
nand NAND2_12669 ( P1_R1171_U494 , P1_R1171_U492 , P1_R1171_U337 );
nand NAND2_12670 ( P1_R1171_U495 , P1_U3063 , P1_R1171_U67 );
nand NAND2_12671 ( P1_R1171_U496 , P1_U3485 , P1_R1171_U68 );
nand NAND2_12672 ( P1_R1171_U497 , P1_R1171_U496 , P1_R1171_U495 );
nand NAND2_12673 ( P1_R1171_U498 , P1_R1171_U362 , P1_R1171_U166 );
nand NAND2_12674 ( P1_R1171_U499 , P1_R1171_U243 , P1_R1171_U497 );
nand NAND2_12675 ( P1_R1171_U500 , P1_U3062 , P1_R1171_U63 );
nand NAND2_12676 ( P1_R1171_U501 , P1_U3482 , P1_R1171_U64 );
nand NAND2_12677 ( P1_R1171_U502 , P1_U3077 , P1_R1171_U30 );
nand NAND2_12678 ( P1_R1171_U503 , P1_U3450 , P1_R1171_U31 );
and AND2_12679 ( P1_R1138_U4 , P1_R1138_U178 , P1_R1138_U177 );
and AND2_12680 ( P1_R1138_U5 , P1_R1138_U179 , P1_R1138_U180 );
and AND2_12681 ( P1_R1138_U6 , P1_R1138_U196 , P1_R1138_U195 );
and AND2_12682 ( P1_R1138_U7 , P1_R1138_U236 , P1_R1138_U235 );
and AND2_12683 ( P1_R1138_U8 , P1_R1138_U245 , P1_R1138_U244 );
and AND2_12684 ( P1_R1138_U9 , P1_R1138_U263 , P1_R1138_U262 );
and AND2_12685 ( P1_R1138_U10 , P1_R1138_U271 , P1_R1138_U270 );
and AND2_12686 ( P1_R1138_U11 , P1_R1138_U350 , P1_R1138_U347 );
and AND2_12687 ( P1_R1138_U12 , P1_R1138_U343 , P1_R1138_U340 );
and AND2_12688 ( P1_R1138_U13 , P1_R1138_U334 , P1_R1138_U331 );
and AND2_12689 ( P1_R1138_U14 , P1_R1138_U325 , P1_R1138_U322 );
and AND2_12690 ( P1_R1138_U15 , P1_R1138_U319 , P1_R1138_U317 );
and AND2_12691 ( P1_R1138_U16 , P1_R1138_U312 , P1_R1138_U309 );
and AND2_12692 ( P1_R1138_U17 , P1_R1138_U234 , P1_R1138_U231 );
and AND2_12693 ( P1_R1138_U18 , P1_R1138_U226 , P1_R1138_U223 );
and AND2_12694 ( P1_R1138_U19 , P1_R1138_U212 , P1_R1138_U209 );
not NOT1_12695 ( P1_R1138_U20 , P1_U3470 );
not NOT1_12696 ( P1_R1138_U21 , P1_U3071 );
not NOT1_12697 ( P1_R1138_U22 , P1_U3070 );
nand NAND2_12698 ( P1_R1138_U23 , P1_U3071 , P1_U3470 );
not NOT1_12699 ( P1_R1138_U24 , P1_U3473 );
not NOT1_12700 ( P1_R1138_U25 , P1_U3464 );
not NOT1_12701 ( P1_R1138_U26 , P1_U3060 );
not NOT1_12702 ( P1_R1138_U27 , P1_U3067 );
not NOT1_12703 ( P1_R1138_U28 , P1_U3458 );
not NOT1_12704 ( P1_R1138_U29 , P1_U3068 );
not NOT1_12705 ( P1_R1138_U30 , P1_U3450 );
not NOT1_12706 ( P1_R1138_U31 , P1_U3077 );
nand NAND2_12707 ( P1_R1138_U32 , P1_U3077 , P1_U3450 );
not NOT1_12708 ( P1_R1138_U33 , P1_U3461 );
not NOT1_12709 ( P1_R1138_U34 , P1_U3064 );
nand NAND2_12710 ( P1_R1138_U35 , P1_U3060 , P1_U3464 );
not NOT1_12711 ( P1_R1138_U36 , P1_U3467 );
not NOT1_12712 ( P1_R1138_U37 , P1_U3476 );
not NOT1_12713 ( P1_R1138_U38 , P1_U3084 );
not NOT1_12714 ( P1_R1138_U39 , P1_U3083 );
not NOT1_12715 ( P1_R1138_U40 , P1_U3479 );
nand NAND2_12716 ( P1_R1138_U41 , P1_R1138_U62 , P1_R1138_U204 );
nand NAND2_12717 ( P1_R1138_U42 , P1_R1138_U118 , P1_R1138_U192 );
nand NAND2_12718 ( P1_R1138_U43 , P1_R1138_U181 , P1_R1138_U182 );
nand NAND2_12719 ( P1_R1138_U44 , P1_U3455 , P1_U3078 );
nand NAND2_12720 ( P1_R1138_U45 , P1_R1138_U122 , P1_R1138_U218 );
nand NAND2_12721 ( P1_R1138_U46 , P1_R1138_U215 , P1_R1138_U214 );
not NOT1_12722 ( P1_R1138_U47 , P1_U3975 );
not NOT1_12723 ( P1_R1138_U48 , P1_U3053 );
not NOT1_12724 ( P1_R1138_U49 , P1_U3057 );
not NOT1_12725 ( P1_R1138_U50 , P1_U3976 );
not NOT1_12726 ( P1_R1138_U51 , P1_U3977 );
not NOT1_12727 ( P1_R1138_U52 , P1_U3058 );
not NOT1_12728 ( P1_R1138_U53 , P1_U3978 );
not NOT1_12729 ( P1_R1138_U54 , P1_U3065 );
not NOT1_12730 ( P1_R1138_U55 , P1_U3981 );
not NOT1_12731 ( P1_R1138_U56 , P1_U3075 );
not NOT1_12732 ( P1_R1138_U57 , P1_U3500 );
not NOT1_12733 ( P1_R1138_U58 , P1_U3073 );
not NOT1_12734 ( P1_R1138_U59 , P1_U3069 );
nand NAND2_12735 ( P1_R1138_U60 , P1_U3073 , P1_U3500 );
not NOT1_12736 ( P1_R1138_U61 , P1_U3503 );
nand NAND2_12737 ( P1_R1138_U62 , P1_U3084 , P1_U3476 );
not NOT1_12738 ( P1_R1138_U63 , P1_U3482 );
not NOT1_12739 ( P1_R1138_U64 , P1_U3062 );
not NOT1_12740 ( P1_R1138_U65 , P1_U3488 );
not NOT1_12741 ( P1_R1138_U66 , P1_U3072 );
not NOT1_12742 ( P1_R1138_U67 , P1_U3485 );
not NOT1_12743 ( P1_R1138_U68 , P1_U3063 );
nand NAND2_12744 ( P1_R1138_U69 , P1_U3063 , P1_U3485 );
not NOT1_12745 ( P1_R1138_U70 , P1_U3491 );
not NOT1_12746 ( P1_R1138_U71 , P1_U3080 );
not NOT1_12747 ( P1_R1138_U72 , P1_U3494 );
not NOT1_12748 ( P1_R1138_U73 , P1_U3079 );
not NOT1_12749 ( P1_R1138_U74 , P1_U3497 );
not NOT1_12750 ( P1_R1138_U75 , P1_U3074 );
not NOT1_12751 ( P1_R1138_U76 , P1_U3506 );
not NOT1_12752 ( P1_R1138_U77 , P1_U3082 );
nand NAND2_12753 ( P1_R1138_U78 , P1_U3082 , P1_U3506 );
not NOT1_12754 ( P1_R1138_U79 , P1_U3508 );
not NOT1_12755 ( P1_R1138_U80 , P1_U3081 );
nand NAND2_12756 ( P1_R1138_U81 , P1_U3081 , P1_U3508 );
not NOT1_12757 ( P1_R1138_U82 , P1_U3982 );
not NOT1_12758 ( P1_R1138_U83 , P1_U3980 );
not NOT1_12759 ( P1_R1138_U84 , P1_U3061 );
not NOT1_12760 ( P1_R1138_U85 , P1_U3979 );
not NOT1_12761 ( P1_R1138_U86 , P1_U3066 );
nand NAND2_12762 ( P1_R1138_U87 , P1_U3976 , P1_U3057 );
not NOT1_12763 ( P1_R1138_U88 , P1_U3054 );
not NOT1_12764 ( P1_R1138_U89 , P1_U3974 );
nand NAND2_12765 ( P1_R1138_U90 , P1_R1138_U305 , P1_R1138_U175 );
not NOT1_12766 ( P1_R1138_U91 , P1_U3076 );
nand NAND2_12767 ( P1_R1138_U92 , P1_R1138_U78 , P1_R1138_U314 );
nand NAND2_12768 ( P1_R1138_U93 , P1_R1138_U260 , P1_R1138_U259 );
nand NAND2_12769 ( P1_R1138_U94 , P1_R1138_U69 , P1_R1138_U336 );
nand NAND2_12770 ( P1_R1138_U95 , P1_R1138_U456 , P1_R1138_U455 );
nand NAND2_12771 ( P1_R1138_U96 , P1_R1138_U503 , P1_R1138_U502 );
nand NAND2_12772 ( P1_R1138_U97 , P1_R1138_U374 , P1_R1138_U373 );
nand NAND2_12773 ( P1_R1138_U98 , P1_R1138_U379 , P1_R1138_U378 );
nand NAND2_12774 ( P1_R1138_U99 , P1_R1138_U386 , P1_R1138_U385 );
nand NAND2_12775 ( P1_R1138_U100 , P1_R1138_U393 , P1_R1138_U392 );
nand NAND2_12776 ( P1_R1138_U101 , P1_R1138_U398 , P1_R1138_U397 );
nand NAND2_12777 ( P1_R1138_U102 , P1_R1138_U407 , P1_R1138_U406 );
nand NAND2_12778 ( P1_R1138_U103 , P1_R1138_U414 , P1_R1138_U413 );
nand NAND2_12779 ( P1_R1138_U104 , P1_R1138_U421 , P1_R1138_U420 );
nand NAND2_12780 ( P1_R1138_U105 , P1_R1138_U428 , P1_R1138_U427 );
nand NAND2_12781 ( P1_R1138_U106 , P1_R1138_U433 , P1_R1138_U432 );
nand NAND2_12782 ( P1_R1138_U107 , P1_R1138_U440 , P1_R1138_U439 );
nand NAND2_12783 ( P1_R1138_U108 , P1_R1138_U447 , P1_R1138_U446 );
nand NAND2_12784 ( P1_R1138_U109 , P1_R1138_U461 , P1_R1138_U460 );
nand NAND2_12785 ( P1_R1138_U110 , P1_R1138_U466 , P1_R1138_U465 );
nand NAND2_12786 ( P1_R1138_U111 , P1_R1138_U473 , P1_R1138_U472 );
nand NAND2_12787 ( P1_R1138_U112 , P1_R1138_U480 , P1_R1138_U479 );
nand NAND2_12788 ( P1_R1138_U113 , P1_R1138_U487 , P1_R1138_U486 );
nand NAND2_12789 ( P1_R1138_U114 , P1_R1138_U494 , P1_R1138_U493 );
nand NAND2_12790 ( P1_R1138_U115 , P1_R1138_U499 , P1_R1138_U498 );
and AND2_12791 ( P1_R1138_U116 , P1_U3458 , P1_U3068 );
and AND2_12792 ( P1_R1138_U117 , P1_R1138_U188 , P1_R1138_U186 );
and AND2_12793 ( P1_R1138_U118 , P1_R1138_U193 , P1_R1138_U191 );
and AND2_12794 ( P1_R1138_U119 , P1_R1138_U200 , P1_R1138_U199 );
and AND3_12795 ( P1_R1138_U120 , P1_R1138_U381 , P1_R1138_U380 , P1_R1138_U23 );
and AND2_12796 ( P1_R1138_U121 , P1_R1138_U211 , P1_R1138_U6 );
and AND2_12797 ( P1_R1138_U122 , P1_R1138_U219 , P1_R1138_U217 );
and AND3_12798 ( P1_R1138_U123 , P1_R1138_U388 , P1_R1138_U387 , P1_R1138_U35 );
and AND2_12799 ( P1_R1138_U124 , P1_R1138_U225 , P1_R1138_U4 );
and AND2_12800 ( P1_R1138_U125 , P1_R1138_U233 , P1_R1138_U180 );
and AND2_12801 ( P1_R1138_U126 , P1_R1138_U203 , P1_R1138_U7 );
and AND2_12802 ( P1_R1138_U127 , P1_R1138_U238 , P1_R1138_U170 );
and AND2_12803 ( P1_R1138_U128 , P1_R1138_U249 , P1_R1138_U8 );
and AND2_12804 ( P1_R1138_U129 , P1_R1138_U247 , P1_R1138_U171 );
and AND2_12805 ( P1_R1138_U130 , P1_R1138_U267 , P1_R1138_U266 );
and AND2_12806 ( P1_R1138_U131 , P1_R1138_U10 , P1_R1138_U281 );
and AND2_12807 ( P1_R1138_U132 , P1_R1138_U284 , P1_R1138_U279 );
and AND2_12808 ( P1_R1138_U133 , P1_R1138_U300 , P1_R1138_U297 );
and AND2_12809 ( P1_R1138_U134 , P1_R1138_U367 , P1_R1138_U301 );
and AND2_12810 ( P1_R1138_U135 , P1_R1138_U159 , P1_R1138_U277 );
and AND3_12811 ( P1_R1138_U136 , P1_R1138_U454 , P1_R1138_U453 , P1_R1138_U81 );
and AND3_12812 ( P1_R1138_U137 , P1_R1138_U468 , P1_R1138_U467 , P1_R1138_U60 );
and AND2_12813 ( P1_R1138_U138 , P1_R1138_U333 , P1_R1138_U9 );
and AND3_12814 ( P1_R1138_U139 , P1_R1138_U489 , P1_R1138_U488 , P1_R1138_U171 );
and AND2_12815 ( P1_R1138_U140 , P1_R1138_U342 , P1_R1138_U8 );
and AND3_12816 ( P1_R1138_U141 , P1_R1138_U501 , P1_R1138_U500 , P1_R1138_U170 );
and AND2_12817 ( P1_R1138_U142 , P1_R1138_U349 , P1_R1138_U7 );
nand NAND2_12818 ( P1_R1138_U143 , P1_R1138_U119 , P1_R1138_U201 );
nand NAND2_12819 ( P1_R1138_U144 , P1_R1138_U216 , P1_R1138_U228 );
not NOT1_12820 ( P1_R1138_U145 , P1_U3055 );
not NOT1_12821 ( P1_R1138_U146 , P1_U3985 );
and AND2_12822 ( P1_R1138_U147 , P1_R1138_U402 , P1_R1138_U401 );
nand NAND3_12823 ( P1_R1138_U148 , P1_R1138_U303 , P1_R1138_U168 , P1_R1138_U363 );
and AND2_12824 ( P1_R1138_U149 , P1_R1138_U409 , P1_R1138_U408 );
nand NAND3_12825 ( P1_R1138_U150 , P1_R1138_U369 , P1_R1138_U368 , P1_R1138_U134 );
and AND2_12826 ( P1_R1138_U151 , P1_R1138_U416 , P1_R1138_U415 );
nand NAND3_12827 ( P1_R1138_U152 , P1_R1138_U364 , P1_R1138_U298 , P1_R1138_U87 );
and AND2_12828 ( P1_R1138_U153 , P1_R1138_U423 , P1_R1138_U422 );
nand NAND2_12829 ( P1_R1138_U154 , P1_R1138_U292 , P1_R1138_U291 );
and AND2_12830 ( P1_R1138_U155 , P1_R1138_U435 , P1_R1138_U434 );
nand NAND2_12831 ( P1_R1138_U156 , P1_R1138_U288 , P1_R1138_U287 );
and AND2_12832 ( P1_R1138_U157 , P1_R1138_U442 , P1_R1138_U441 );
nand NAND2_12833 ( P1_R1138_U158 , P1_R1138_U132 , P1_R1138_U283 );
and AND2_12834 ( P1_R1138_U159 , P1_R1138_U449 , P1_R1138_U448 );
nand NAND2_12835 ( P1_R1138_U160 , P1_R1138_U44 , P1_R1138_U326 );
nand NAND2_12836 ( P1_R1138_U161 , P1_R1138_U130 , P1_R1138_U268 );
and AND2_12837 ( P1_R1138_U162 , P1_R1138_U475 , P1_R1138_U474 );
nand NAND2_12838 ( P1_R1138_U163 , P1_R1138_U256 , P1_R1138_U255 );
and AND2_12839 ( P1_R1138_U164 , P1_R1138_U482 , P1_R1138_U481 );
nand NAND2_12840 ( P1_R1138_U165 , P1_R1138_U252 , P1_R1138_U251 );
nand NAND2_12841 ( P1_R1138_U166 , P1_R1138_U242 , P1_R1138_U241 );
nand NAND2_12842 ( P1_R1138_U167 , P1_R1138_U366 , P1_R1138_U365 );
nand NAND2_12843 ( P1_R1138_U168 , P1_U3054 , P1_R1138_U150 );
not NOT1_12844 ( P1_R1138_U169 , P1_R1138_U35 );
nand NAND2_12845 ( P1_R1138_U170 , P1_U3479 , P1_U3083 );
nand NAND2_12846 ( P1_R1138_U171 , P1_U3072 , P1_U3488 );
nand NAND2_12847 ( P1_R1138_U172 , P1_U3058 , P1_U3977 );
not NOT1_12848 ( P1_R1138_U173 , P1_R1138_U69 );
not NOT1_12849 ( P1_R1138_U174 , P1_R1138_U78 );
nand NAND2_12850 ( P1_R1138_U175 , P1_U3065 , P1_U3978 );
not NOT1_12851 ( P1_R1138_U176 , P1_R1138_U62 );
or OR2_12852 ( P1_R1138_U177 , P1_U3067 , P1_U3467 );
or OR2_12853 ( P1_R1138_U178 , P1_U3060 , P1_U3464 );
or OR2_12854 ( P1_R1138_U179 , P1_U3461 , P1_U3064 );
or OR2_12855 ( P1_R1138_U180 , P1_U3458 , P1_U3068 );
not NOT1_12856 ( P1_R1138_U181 , P1_R1138_U32 );
or OR2_12857 ( P1_R1138_U182 , P1_U3455 , P1_U3078 );
not NOT1_12858 ( P1_R1138_U183 , P1_R1138_U43 );
not NOT1_12859 ( P1_R1138_U184 , P1_R1138_U44 );
nand NAND2_12860 ( P1_R1138_U185 , P1_R1138_U43 , P1_R1138_U44 );
nand NAND2_12861 ( P1_R1138_U186 , P1_R1138_U116 , P1_R1138_U179 );
nand NAND2_12862 ( P1_R1138_U187 , P1_R1138_U5 , P1_R1138_U185 );
nand NAND2_12863 ( P1_R1138_U188 , P1_U3064 , P1_U3461 );
nand NAND2_12864 ( P1_R1138_U189 , P1_R1138_U117 , P1_R1138_U187 );
nand NAND2_12865 ( P1_R1138_U190 , P1_R1138_U36 , P1_R1138_U35 );
nand NAND2_12866 ( P1_R1138_U191 , P1_U3067 , P1_R1138_U190 );
nand NAND2_12867 ( P1_R1138_U192 , P1_R1138_U4 , P1_R1138_U189 );
nand NAND2_12868 ( P1_R1138_U193 , P1_U3467 , P1_R1138_U169 );
not NOT1_12869 ( P1_R1138_U194 , P1_R1138_U42 );
or OR2_12870 ( P1_R1138_U195 , P1_U3070 , P1_U3473 );
or OR2_12871 ( P1_R1138_U196 , P1_U3071 , P1_U3470 );
not NOT1_12872 ( P1_R1138_U197 , P1_R1138_U23 );
nand NAND2_12873 ( P1_R1138_U198 , P1_R1138_U24 , P1_R1138_U23 );
nand NAND2_12874 ( P1_R1138_U199 , P1_U3070 , P1_R1138_U198 );
nand NAND2_12875 ( P1_R1138_U200 , P1_U3473 , P1_R1138_U197 );
nand NAND2_12876 ( P1_R1138_U201 , P1_R1138_U6 , P1_R1138_U42 );
not NOT1_12877 ( P1_R1138_U202 , P1_R1138_U143 );
or OR2_12878 ( P1_R1138_U203 , P1_U3476 , P1_U3084 );
nand NAND2_12879 ( P1_R1138_U204 , P1_R1138_U203 , P1_R1138_U143 );
not NOT1_12880 ( P1_R1138_U205 , P1_R1138_U41 );
or OR2_12881 ( P1_R1138_U206 , P1_U3083 , P1_U3479 );
or OR2_12882 ( P1_R1138_U207 , P1_U3470 , P1_U3071 );
nand NAND2_12883 ( P1_R1138_U208 , P1_R1138_U207 , P1_R1138_U42 );
nand NAND2_12884 ( P1_R1138_U209 , P1_R1138_U120 , P1_R1138_U208 );
nand NAND2_12885 ( P1_R1138_U210 , P1_R1138_U194 , P1_R1138_U23 );
nand NAND2_12886 ( P1_R1138_U211 , P1_U3473 , P1_U3070 );
nand NAND2_12887 ( P1_R1138_U212 , P1_R1138_U121 , P1_R1138_U210 );
or OR2_12888 ( P1_R1138_U213 , P1_U3071 , P1_U3470 );
nand NAND2_12889 ( P1_R1138_U214 , P1_R1138_U184 , P1_R1138_U180 );
nand NAND2_12890 ( P1_R1138_U215 , P1_U3068 , P1_U3458 );
not NOT1_12891 ( P1_R1138_U216 , P1_R1138_U46 );
nand NAND2_12892 ( P1_R1138_U217 , P1_R1138_U183 , P1_R1138_U5 );
nand NAND2_12893 ( P1_R1138_U218 , P1_R1138_U46 , P1_R1138_U179 );
nand NAND2_12894 ( P1_R1138_U219 , P1_U3064 , P1_U3461 );
not NOT1_12895 ( P1_R1138_U220 , P1_R1138_U45 );
or OR2_12896 ( P1_R1138_U221 , P1_U3464 , P1_U3060 );
nand NAND2_12897 ( P1_R1138_U222 , P1_R1138_U221 , P1_R1138_U45 );
nand NAND2_12898 ( P1_R1138_U223 , P1_R1138_U123 , P1_R1138_U222 );
nand NAND2_12899 ( P1_R1138_U224 , P1_R1138_U220 , P1_R1138_U35 );
nand NAND2_12900 ( P1_R1138_U225 , P1_U3467 , P1_U3067 );
nand NAND2_12901 ( P1_R1138_U226 , P1_R1138_U124 , P1_R1138_U224 );
or OR2_12902 ( P1_R1138_U227 , P1_U3060 , P1_U3464 );
nand NAND2_12903 ( P1_R1138_U228 , P1_R1138_U183 , P1_R1138_U180 );
not NOT1_12904 ( P1_R1138_U229 , P1_R1138_U144 );
nand NAND2_12905 ( P1_R1138_U230 , P1_U3064 , P1_U3461 );
nand NAND4_12906 ( P1_R1138_U231 , P1_R1138_U400 , P1_R1138_U399 , P1_R1138_U44 , P1_R1138_U43 );
nand NAND2_12907 ( P1_R1138_U232 , P1_R1138_U44 , P1_R1138_U43 );
nand NAND2_12908 ( P1_R1138_U233 , P1_U3068 , P1_U3458 );
nand NAND2_12909 ( P1_R1138_U234 , P1_R1138_U125 , P1_R1138_U232 );
or OR2_12910 ( P1_R1138_U235 , P1_U3083 , P1_U3479 );
or OR2_12911 ( P1_R1138_U236 , P1_U3062 , P1_U3482 );
nand NAND2_12912 ( P1_R1138_U237 , P1_R1138_U176 , P1_R1138_U7 );
nand NAND2_12913 ( P1_R1138_U238 , P1_U3062 , P1_U3482 );
nand NAND2_12914 ( P1_R1138_U239 , P1_R1138_U127 , P1_R1138_U237 );
or OR2_12915 ( P1_R1138_U240 , P1_U3482 , P1_U3062 );
nand NAND2_12916 ( P1_R1138_U241 , P1_R1138_U126 , P1_R1138_U143 );
nand NAND2_12917 ( P1_R1138_U242 , P1_R1138_U240 , P1_R1138_U239 );
not NOT1_12918 ( P1_R1138_U243 , P1_R1138_U166 );
or OR2_12919 ( P1_R1138_U244 , P1_U3080 , P1_U3491 );
or OR2_12920 ( P1_R1138_U245 , P1_U3072 , P1_U3488 );
nand NAND2_12921 ( P1_R1138_U246 , P1_R1138_U173 , P1_R1138_U8 );
nand NAND2_12922 ( P1_R1138_U247 , P1_U3080 , P1_U3491 );
nand NAND2_12923 ( P1_R1138_U248 , P1_R1138_U129 , P1_R1138_U246 );
or OR2_12924 ( P1_R1138_U249 , P1_U3485 , P1_U3063 );
or OR2_12925 ( P1_R1138_U250 , P1_U3491 , P1_U3080 );
nand NAND2_12926 ( P1_R1138_U251 , P1_R1138_U128 , P1_R1138_U166 );
nand NAND2_12927 ( P1_R1138_U252 , P1_R1138_U250 , P1_R1138_U248 );
not NOT1_12928 ( P1_R1138_U253 , P1_R1138_U165 );
or OR2_12929 ( P1_R1138_U254 , P1_U3494 , P1_U3079 );
nand NAND2_12930 ( P1_R1138_U255 , P1_R1138_U254 , P1_R1138_U165 );
nand NAND2_12931 ( P1_R1138_U256 , P1_U3079 , P1_U3494 );
not NOT1_12932 ( P1_R1138_U257 , P1_R1138_U163 );
or OR2_12933 ( P1_R1138_U258 , P1_U3497 , P1_U3074 );
nand NAND2_12934 ( P1_R1138_U259 , P1_R1138_U258 , P1_R1138_U163 );
nand NAND2_12935 ( P1_R1138_U260 , P1_U3074 , P1_U3497 );
not NOT1_12936 ( P1_R1138_U261 , P1_R1138_U93 );
or OR2_12937 ( P1_R1138_U262 , P1_U3069 , P1_U3503 );
or OR2_12938 ( P1_R1138_U263 , P1_U3073 , P1_U3500 );
not NOT1_12939 ( P1_R1138_U264 , P1_R1138_U60 );
nand NAND2_12940 ( P1_R1138_U265 , P1_R1138_U61 , P1_R1138_U60 );
nand NAND2_12941 ( P1_R1138_U266 , P1_U3069 , P1_R1138_U265 );
nand NAND2_12942 ( P1_R1138_U267 , P1_U3503 , P1_R1138_U264 );
nand NAND2_12943 ( P1_R1138_U268 , P1_R1138_U9 , P1_R1138_U93 );
not NOT1_12944 ( P1_R1138_U269 , P1_R1138_U161 );
or OR2_12945 ( P1_R1138_U270 , P1_U3076 , P1_U3982 );
or OR2_12946 ( P1_R1138_U271 , P1_U3081 , P1_U3508 );
or OR2_12947 ( P1_R1138_U272 , P1_U3075 , P1_U3981 );
not NOT1_12948 ( P1_R1138_U273 , P1_R1138_U81 );
nand NAND2_12949 ( P1_R1138_U274 , P1_U3982 , P1_R1138_U273 );
nand NAND2_12950 ( P1_R1138_U275 , P1_R1138_U274 , P1_R1138_U91 );
nand NAND2_12951 ( P1_R1138_U276 , P1_R1138_U81 , P1_R1138_U82 );
nand NAND2_12952 ( P1_R1138_U277 , P1_R1138_U276 , P1_R1138_U275 );
nand NAND2_12953 ( P1_R1138_U278 , P1_R1138_U174 , P1_R1138_U10 );
nand NAND2_12954 ( P1_R1138_U279 , P1_U3075 , P1_U3981 );
nand NAND2_12955 ( P1_R1138_U280 , P1_R1138_U277 , P1_R1138_U278 );
or OR2_12956 ( P1_R1138_U281 , P1_U3506 , P1_U3082 );
or OR2_12957 ( P1_R1138_U282 , P1_U3981 , P1_U3075 );
nand NAND3_12958 ( P1_R1138_U283 , P1_R1138_U272 , P1_R1138_U161 , P1_R1138_U131 );
nand NAND2_12959 ( P1_R1138_U284 , P1_R1138_U282 , P1_R1138_U280 );
not NOT1_12960 ( P1_R1138_U285 , P1_R1138_U158 );
or OR2_12961 ( P1_R1138_U286 , P1_U3980 , P1_U3061 );
nand NAND2_12962 ( P1_R1138_U287 , P1_R1138_U286 , P1_R1138_U158 );
nand NAND2_12963 ( P1_R1138_U288 , P1_U3061 , P1_U3980 );
not NOT1_12964 ( P1_R1138_U289 , P1_R1138_U156 );
or OR2_12965 ( P1_R1138_U290 , P1_U3979 , P1_U3066 );
nand NAND2_12966 ( P1_R1138_U291 , P1_R1138_U290 , P1_R1138_U156 );
nand NAND2_12967 ( P1_R1138_U292 , P1_U3066 , P1_U3979 );
not NOT1_12968 ( P1_R1138_U293 , P1_R1138_U154 );
or OR2_12969 ( P1_R1138_U294 , P1_U3058 , P1_U3977 );
nand NAND2_12970 ( P1_R1138_U295 , P1_R1138_U175 , P1_R1138_U172 );
not NOT1_12971 ( P1_R1138_U296 , P1_R1138_U87 );
or OR2_12972 ( P1_R1138_U297 , P1_U3978 , P1_U3065 );
nand NAND3_12973 ( P1_R1138_U298 , P1_R1138_U154 , P1_R1138_U297 , P1_R1138_U167 );
not NOT1_12974 ( P1_R1138_U299 , P1_R1138_U152 );
or OR2_12975 ( P1_R1138_U300 , P1_U3975 , P1_U3053 );
nand NAND2_12976 ( P1_R1138_U301 , P1_U3053 , P1_U3975 );
not NOT1_12977 ( P1_R1138_U302 , P1_R1138_U150 );
nand NAND2_12978 ( P1_R1138_U303 , P1_U3974 , P1_R1138_U150 );
not NOT1_12979 ( P1_R1138_U304 , P1_R1138_U148 );
nand NAND2_12980 ( P1_R1138_U305 , P1_R1138_U297 , P1_R1138_U154 );
not NOT1_12981 ( P1_R1138_U306 , P1_R1138_U90 );
or OR2_12982 ( P1_R1138_U307 , P1_U3977 , P1_U3058 );
nand NAND2_12983 ( P1_R1138_U308 , P1_R1138_U307 , P1_R1138_U90 );
nand NAND3_12984 ( P1_R1138_U309 , P1_R1138_U308 , P1_R1138_U172 , P1_R1138_U153 );
nand NAND2_12985 ( P1_R1138_U310 , P1_R1138_U306 , P1_R1138_U172 );
nand NAND2_12986 ( P1_R1138_U311 , P1_U3976 , P1_U3057 );
nand NAND3_12987 ( P1_R1138_U312 , P1_R1138_U310 , P1_R1138_U311 , P1_R1138_U167 );
or OR2_12988 ( P1_R1138_U313 , P1_U3058 , P1_U3977 );
nand NAND2_12989 ( P1_R1138_U314 , P1_R1138_U281 , P1_R1138_U161 );
not NOT1_12990 ( P1_R1138_U315 , P1_R1138_U92 );
nand NAND2_12991 ( P1_R1138_U316 , P1_R1138_U10 , P1_R1138_U92 );
nand NAND2_12992 ( P1_R1138_U317 , P1_R1138_U135 , P1_R1138_U316 );
nand NAND2_12993 ( P1_R1138_U318 , P1_R1138_U316 , P1_R1138_U277 );
nand NAND2_12994 ( P1_R1138_U319 , P1_R1138_U452 , P1_R1138_U318 );
or OR2_12995 ( P1_R1138_U320 , P1_U3508 , P1_U3081 );
nand NAND2_12996 ( P1_R1138_U321 , P1_R1138_U320 , P1_R1138_U92 );
nand NAND2_12997 ( P1_R1138_U322 , P1_R1138_U136 , P1_R1138_U321 );
nand NAND2_12998 ( P1_R1138_U323 , P1_R1138_U315 , P1_R1138_U81 );
nand NAND2_12999 ( P1_R1138_U324 , P1_U3076 , P1_U3982 );
nand NAND3_13000 ( P1_R1138_U325 , P1_R1138_U324 , P1_R1138_U323 , P1_R1138_U10 );
or OR2_13001 ( P1_R1138_U326 , P1_U3455 , P1_U3078 );
not NOT1_13002 ( P1_R1138_U327 , P1_R1138_U160 );
or OR2_13003 ( P1_R1138_U328 , P1_U3081 , P1_U3508 );
or OR2_13004 ( P1_R1138_U329 , P1_U3500 , P1_U3073 );
nand NAND2_13005 ( P1_R1138_U330 , P1_R1138_U329 , P1_R1138_U93 );
nand NAND2_13006 ( P1_R1138_U331 , P1_R1138_U137 , P1_R1138_U330 );
nand NAND2_13007 ( P1_R1138_U332 , P1_R1138_U261 , P1_R1138_U60 );
nand NAND2_13008 ( P1_R1138_U333 , P1_U3503 , P1_U3069 );
nand NAND2_13009 ( P1_R1138_U334 , P1_R1138_U138 , P1_R1138_U332 );
or OR2_13010 ( P1_R1138_U335 , P1_U3073 , P1_U3500 );
nand NAND2_13011 ( P1_R1138_U336 , P1_R1138_U249 , P1_R1138_U166 );
not NOT1_13012 ( P1_R1138_U337 , P1_R1138_U94 );
or OR2_13013 ( P1_R1138_U338 , P1_U3488 , P1_U3072 );
nand NAND2_13014 ( P1_R1138_U339 , P1_R1138_U338 , P1_R1138_U94 );
nand NAND2_13015 ( P1_R1138_U340 , P1_R1138_U139 , P1_R1138_U339 );
nand NAND2_13016 ( P1_R1138_U341 , P1_R1138_U337 , P1_R1138_U171 );
nand NAND2_13017 ( P1_R1138_U342 , P1_U3080 , P1_U3491 );
nand NAND2_13018 ( P1_R1138_U343 , P1_R1138_U140 , P1_R1138_U341 );
or OR2_13019 ( P1_R1138_U344 , P1_U3072 , P1_U3488 );
or OR2_13020 ( P1_R1138_U345 , P1_U3479 , P1_U3083 );
nand NAND2_13021 ( P1_R1138_U346 , P1_R1138_U345 , P1_R1138_U41 );
nand NAND2_13022 ( P1_R1138_U347 , P1_R1138_U141 , P1_R1138_U346 );
nand NAND2_13023 ( P1_R1138_U348 , P1_R1138_U205 , P1_R1138_U170 );
nand NAND2_13024 ( P1_R1138_U349 , P1_U3062 , P1_U3482 );
nand NAND2_13025 ( P1_R1138_U350 , P1_R1138_U142 , P1_R1138_U348 );
nand NAND2_13026 ( P1_R1138_U351 , P1_R1138_U206 , P1_R1138_U170 );
nand NAND2_13027 ( P1_R1138_U352 , P1_R1138_U203 , P1_R1138_U62 );
nand NAND2_13028 ( P1_R1138_U353 , P1_R1138_U213 , P1_R1138_U23 );
nand NAND2_13029 ( P1_R1138_U354 , P1_R1138_U227 , P1_R1138_U35 );
nand NAND2_13030 ( P1_R1138_U355 , P1_R1138_U230 , P1_R1138_U179 );
nand NAND2_13031 ( P1_R1138_U356 , P1_R1138_U313 , P1_R1138_U172 );
nand NAND2_13032 ( P1_R1138_U357 , P1_R1138_U297 , P1_R1138_U175 );
nand NAND2_13033 ( P1_R1138_U358 , P1_R1138_U328 , P1_R1138_U81 );
nand NAND2_13034 ( P1_R1138_U359 , P1_R1138_U281 , P1_R1138_U78 );
nand NAND2_13035 ( P1_R1138_U360 , P1_R1138_U335 , P1_R1138_U60 );
nand NAND2_13036 ( P1_R1138_U361 , P1_R1138_U344 , P1_R1138_U171 );
nand NAND2_13037 ( P1_R1138_U362 , P1_R1138_U249 , P1_R1138_U69 );
nand NAND2_13038 ( P1_R1138_U363 , P1_U3974 , P1_U3054 );
nand NAND2_13039 ( P1_R1138_U364 , P1_R1138_U295 , P1_R1138_U167 );
nand NAND2_13040 ( P1_R1138_U365 , P1_U3057 , P1_R1138_U294 );
nand NAND2_13041 ( P1_R1138_U366 , P1_U3976 , P1_R1138_U294 );
nand NAND3_13042 ( P1_R1138_U367 , P1_R1138_U295 , P1_R1138_U167 , P1_R1138_U300 );
nand NAND3_13043 ( P1_R1138_U368 , P1_R1138_U154 , P1_R1138_U167 , P1_R1138_U133 );
nand NAND2_13044 ( P1_R1138_U369 , P1_R1138_U296 , P1_R1138_U300 );
nand NAND2_13045 ( P1_R1138_U370 , P1_U3083 , P1_R1138_U40 );
nand NAND2_13046 ( P1_R1138_U371 , P1_U3479 , P1_R1138_U39 );
nand NAND2_13047 ( P1_R1138_U372 , P1_R1138_U371 , P1_R1138_U370 );
nand NAND2_13048 ( P1_R1138_U373 , P1_R1138_U351 , P1_R1138_U41 );
nand NAND2_13049 ( P1_R1138_U374 , P1_R1138_U372 , P1_R1138_U205 );
nand NAND2_13050 ( P1_R1138_U375 , P1_U3084 , P1_R1138_U37 );
nand NAND2_13051 ( P1_R1138_U376 , P1_U3476 , P1_R1138_U38 );
nand NAND2_13052 ( P1_R1138_U377 , P1_R1138_U376 , P1_R1138_U375 );
nand NAND2_13053 ( P1_R1138_U378 , P1_R1138_U352 , P1_R1138_U143 );
nand NAND2_13054 ( P1_R1138_U379 , P1_R1138_U202 , P1_R1138_U377 );
nand NAND2_13055 ( P1_R1138_U380 , P1_U3070 , P1_R1138_U24 );
nand NAND2_13056 ( P1_R1138_U381 , P1_U3473 , P1_R1138_U22 );
nand NAND2_13057 ( P1_R1138_U382 , P1_U3071 , P1_R1138_U20 );
nand NAND2_13058 ( P1_R1138_U383 , P1_U3470 , P1_R1138_U21 );
nand NAND2_13059 ( P1_R1138_U384 , P1_R1138_U383 , P1_R1138_U382 );
nand NAND2_13060 ( P1_R1138_U385 , P1_R1138_U353 , P1_R1138_U42 );
nand NAND2_13061 ( P1_R1138_U386 , P1_R1138_U384 , P1_R1138_U194 );
nand NAND2_13062 ( P1_R1138_U387 , P1_U3067 , P1_R1138_U36 );
nand NAND2_13063 ( P1_R1138_U388 , P1_U3467 , P1_R1138_U27 );
nand NAND2_13064 ( P1_R1138_U389 , P1_U3060 , P1_R1138_U25 );
nand NAND2_13065 ( P1_R1138_U390 , P1_U3464 , P1_R1138_U26 );
nand NAND2_13066 ( P1_R1138_U391 , P1_R1138_U390 , P1_R1138_U389 );
nand NAND2_13067 ( P1_R1138_U392 , P1_R1138_U354 , P1_R1138_U45 );
nand NAND2_13068 ( P1_R1138_U393 , P1_R1138_U391 , P1_R1138_U220 );
nand NAND2_13069 ( P1_R1138_U394 , P1_U3064 , P1_R1138_U33 );
nand NAND2_13070 ( P1_R1138_U395 , P1_U3461 , P1_R1138_U34 );
nand NAND2_13071 ( P1_R1138_U396 , P1_R1138_U395 , P1_R1138_U394 );
nand NAND2_13072 ( P1_R1138_U397 , P1_R1138_U355 , P1_R1138_U144 );
nand NAND2_13073 ( P1_R1138_U398 , P1_R1138_U229 , P1_R1138_U396 );
nand NAND2_13074 ( P1_R1138_U399 , P1_U3068 , P1_R1138_U28 );
nand NAND2_13075 ( P1_R1138_U400 , P1_U3458 , P1_R1138_U29 );
nand NAND2_13076 ( P1_R1138_U401 , P1_U3055 , P1_R1138_U146 );
nand NAND2_13077 ( P1_R1138_U402 , P1_U3985 , P1_R1138_U145 );
nand NAND2_13078 ( P1_R1138_U403 , P1_U3055 , P1_R1138_U146 );
nand NAND2_13079 ( P1_R1138_U404 , P1_U3985 , P1_R1138_U145 );
nand NAND2_13080 ( P1_R1138_U405 , P1_R1138_U404 , P1_R1138_U403 );
nand NAND2_13081 ( P1_R1138_U406 , P1_R1138_U147 , P1_R1138_U148 );
nand NAND2_13082 ( P1_R1138_U407 , P1_R1138_U304 , P1_R1138_U405 );
nand NAND2_13083 ( P1_R1138_U408 , P1_U3054 , P1_R1138_U89 );
nand NAND2_13084 ( P1_R1138_U409 , P1_U3974 , P1_R1138_U88 );
nand NAND2_13085 ( P1_R1138_U410 , P1_U3054 , P1_R1138_U89 );
nand NAND2_13086 ( P1_R1138_U411 , P1_U3974 , P1_R1138_U88 );
nand NAND2_13087 ( P1_R1138_U412 , P1_R1138_U411 , P1_R1138_U410 );
nand NAND2_13088 ( P1_R1138_U413 , P1_R1138_U149 , P1_R1138_U150 );
nand NAND2_13089 ( P1_R1138_U414 , P1_R1138_U302 , P1_R1138_U412 );
nand NAND2_13090 ( P1_R1138_U415 , P1_U3053 , P1_R1138_U47 );
nand NAND2_13091 ( P1_R1138_U416 , P1_U3975 , P1_R1138_U48 );
nand NAND2_13092 ( P1_R1138_U417 , P1_U3053 , P1_R1138_U47 );
nand NAND2_13093 ( P1_R1138_U418 , P1_U3975 , P1_R1138_U48 );
nand NAND2_13094 ( P1_R1138_U419 , P1_R1138_U418 , P1_R1138_U417 );
nand NAND2_13095 ( P1_R1138_U420 , P1_R1138_U151 , P1_R1138_U152 );
nand NAND2_13096 ( P1_R1138_U421 , P1_R1138_U299 , P1_R1138_U419 );
nand NAND2_13097 ( P1_R1138_U422 , P1_U3057 , P1_R1138_U50 );
nand NAND2_13098 ( P1_R1138_U423 , P1_U3976 , P1_R1138_U49 );
nand NAND2_13099 ( P1_R1138_U424 , P1_U3058 , P1_R1138_U51 );
nand NAND2_13100 ( P1_R1138_U425 , P1_U3977 , P1_R1138_U52 );
nand NAND2_13101 ( P1_R1138_U426 , P1_R1138_U425 , P1_R1138_U424 );
nand NAND2_13102 ( P1_R1138_U427 , P1_R1138_U356 , P1_R1138_U90 );
nand NAND2_13103 ( P1_R1138_U428 , P1_R1138_U426 , P1_R1138_U306 );
nand NAND2_13104 ( P1_R1138_U429 , P1_U3065 , P1_R1138_U53 );
nand NAND2_13105 ( P1_R1138_U430 , P1_U3978 , P1_R1138_U54 );
nand NAND2_13106 ( P1_R1138_U431 , P1_R1138_U430 , P1_R1138_U429 );
nand NAND2_13107 ( P1_R1138_U432 , P1_R1138_U357 , P1_R1138_U154 );
nand NAND2_13108 ( P1_R1138_U433 , P1_R1138_U293 , P1_R1138_U431 );
nand NAND2_13109 ( P1_R1138_U434 , P1_U3066 , P1_R1138_U85 );
nand NAND2_13110 ( P1_R1138_U435 , P1_U3979 , P1_R1138_U86 );
nand NAND2_13111 ( P1_R1138_U436 , P1_U3066 , P1_R1138_U85 );
nand NAND2_13112 ( P1_R1138_U437 , P1_U3979 , P1_R1138_U86 );
nand NAND2_13113 ( P1_R1138_U438 , P1_R1138_U437 , P1_R1138_U436 );
nand NAND2_13114 ( P1_R1138_U439 , P1_R1138_U155 , P1_R1138_U156 );
nand NAND2_13115 ( P1_R1138_U440 , P1_R1138_U289 , P1_R1138_U438 );
nand NAND2_13116 ( P1_R1138_U441 , P1_U3061 , P1_R1138_U83 );
nand NAND2_13117 ( P1_R1138_U442 , P1_U3980 , P1_R1138_U84 );
nand NAND2_13118 ( P1_R1138_U443 , P1_U3061 , P1_R1138_U83 );
nand NAND2_13119 ( P1_R1138_U444 , P1_U3980 , P1_R1138_U84 );
nand NAND2_13120 ( P1_R1138_U445 , P1_R1138_U444 , P1_R1138_U443 );
nand NAND2_13121 ( P1_R1138_U446 , P1_R1138_U157 , P1_R1138_U158 );
nand NAND2_13122 ( P1_R1138_U447 , P1_R1138_U285 , P1_R1138_U445 );
nand NAND2_13123 ( P1_R1138_U448 , P1_U3075 , P1_R1138_U55 );
nand NAND2_13124 ( P1_R1138_U449 , P1_U3981 , P1_R1138_U56 );
nand NAND2_13125 ( P1_R1138_U450 , P1_U3075 , P1_R1138_U55 );
nand NAND2_13126 ( P1_R1138_U451 , P1_U3981 , P1_R1138_U56 );
nand NAND2_13127 ( P1_R1138_U452 , P1_R1138_U451 , P1_R1138_U450 );
nand NAND2_13128 ( P1_R1138_U453 , P1_U3076 , P1_R1138_U82 );
nand NAND2_13129 ( P1_R1138_U454 , P1_U3982 , P1_R1138_U91 );
nand NAND2_13130 ( P1_R1138_U455 , P1_R1138_U181 , P1_R1138_U160 );
nand NAND2_13131 ( P1_R1138_U456 , P1_R1138_U327 , P1_R1138_U32 );
nand NAND2_13132 ( P1_R1138_U457 , P1_U3081 , P1_R1138_U79 );
nand NAND2_13133 ( P1_R1138_U458 , P1_U3508 , P1_R1138_U80 );
nand NAND2_13134 ( P1_R1138_U459 , P1_R1138_U458 , P1_R1138_U457 );
nand NAND2_13135 ( P1_R1138_U460 , P1_R1138_U358 , P1_R1138_U92 );
nand NAND2_13136 ( P1_R1138_U461 , P1_R1138_U459 , P1_R1138_U315 );
nand NAND2_13137 ( P1_R1138_U462 , P1_U3082 , P1_R1138_U76 );
nand NAND2_13138 ( P1_R1138_U463 , P1_U3506 , P1_R1138_U77 );
nand NAND2_13139 ( P1_R1138_U464 , P1_R1138_U463 , P1_R1138_U462 );
nand NAND2_13140 ( P1_R1138_U465 , P1_R1138_U359 , P1_R1138_U161 );
nand NAND2_13141 ( P1_R1138_U466 , P1_R1138_U269 , P1_R1138_U464 );
nand NAND2_13142 ( P1_R1138_U467 , P1_U3069 , P1_R1138_U61 );
nand NAND2_13143 ( P1_R1138_U468 , P1_U3503 , P1_R1138_U59 );
nand NAND2_13144 ( P1_R1138_U469 , P1_U3073 , P1_R1138_U57 );
nand NAND2_13145 ( P1_R1138_U470 , P1_U3500 , P1_R1138_U58 );
nand NAND2_13146 ( P1_R1138_U471 , P1_R1138_U470 , P1_R1138_U469 );
nand NAND2_13147 ( P1_R1138_U472 , P1_R1138_U360 , P1_R1138_U93 );
nand NAND2_13148 ( P1_R1138_U473 , P1_R1138_U471 , P1_R1138_U261 );
nand NAND2_13149 ( P1_R1138_U474 , P1_U3074 , P1_R1138_U74 );
nand NAND2_13150 ( P1_R1138_U475 , P1_U3497 , P1_R1138_U75 );
nand NAND2_13151 ( P1_R1138_U476 , P1_U3074 , P1_R1138_U74 );
nand NAND2_13152 ( P1_R1138_U477 , P1_U3497 , P1_R1138_U75 );
nand NAND2_13153 ( P1_R1138_U478 , P1_R1138_U477 , P1_R1138_U476 );
nand NAND2_13154 ( P1_R1138_U479 , P1_R1138_U162 , P1_R1138_U163 );
nand NAND2_13155 ( P1_R1138_U480 , P1_R1138_U257 , P1_R1138_U478 );
nand NAND2_13156 ( P1_R1138_U481 , P1_U3079 , P1_R1138_U72 );
nand NAND2_13157 ( P1_R1138_U482 , P1_U3494 , P1_R1138_U73 );
nand NAND2_13158 ( P1_R1138_U483 , P1_U3079 , P1_R1138_U72 );
nand NAND2_13159 ( P1_R1138_U484 , P1_U3494 , P1_R1138_U73 );
nand NAND2_13160 ( P1_R1138_U485 , P1_R1138_U484 , P1_R1138_U483 );
nand NAND2_13161 ( P1_R1138_U486 , P1_R1138_U164 , P1_R1138_U165 );
nand NAND2_13162 ( P1_R1138_U487 , P1_R1138_U253 , P1_R1138_U485 );
nand NAND2_13163 ( P1_R1138_U488 , P1_U3080 , P1_R1138_U70 );
nand NAND2_13164 ( P1_R1138_U489 , P1_U3491 , P1_R1138_U71 );
nand NAND2_13165 ( P1_R1138_U490 , P1_U3072 , P1_R1138_U65 );
nand NAND2_13166 ( P1_R1138_U491 , P1_U3488 , P1_R1138_U66 );
nand NAND2_13167 ( P1_R1138_U492 , P1_R1138_U491 , P1_R1138_U490 );
nand NAND2_13168 ( P1_R1138_U493 , P1_R1138_U361 , P1_R1138_U94 );
nand NAND2_13169 ( P1_R1138_U494 , P1_R1138_U492 , P1_R1138_U337 );
nand NAND2_13170 ( P1_R1138_U495 , P1_U3063 , P1_R1138_U67 );
nand NAND2_13171 ( P1_R1138_U496 , P1_U3485 , P1_R1138_U68 );
nand NAND2_13172 ( P1_R1138_U497 , P1_R1138_U496 , P1_R1138_U495 );
nand NAND2_13173 ( P1_R1138_U498 , P1_R1138_U362 , P1_R1138_U166 );
nand NAND2_13174 ( P1_R1138_U499 , P1_R1138_U243 , P1_R1138_U497 );
nand NAND2_13175 ( P1_R1138_U500 , P1_U3062 , P1_R1138_U63 );
nand NAND2_13176 ( P1_R1138_U501 , P1_U3482 , P1_R1138_U64 );
nand NAND2_13177 ( P1_R1138_U502 , P1_U3077 , P1_R1138_U30 );
nand NAND2_13178 ( P1_R1138_U503 , P1_U3450 , P1_R1138_U31 );
and AND2_13179 ( P1_R1222_U4 , P1_R1222_U178 , P1_R1222_U177 );
and AND2_13180 ( P1_R1222_U5 , P1_R1222_U179 , P1_R1222_U180 );
and AND2_13181 ( P1_R1222_U6 , P1_R1222_U196 , P1_R1222_U195 );
and AND2_13182 ( P1_R1222_U7 , P1_R1222_U236 , P1_R1222_U235 );
and AND2_13183 ( P1_R1222_U8 , P1_R1222_U245 , P1_R1222_U244 );
and AND2_13184 ( P1_R1222_U9 , P1_R1222_U263 , P1_R1222_U262 );
and AND2_13185 ( P1_R1222_U10 , P1_R1222_U271 , P1_R1222_U270 );
and AND2_13186 ( P1_R1222_U11 , P1_R1222_U350 , P1_R1222_U347 );
and AND2_13187 ( P1_R1222_U12 , P1_R1222_U343 , P1_R1222_U340 );
and AND2_13188 ( P1_R1222_U13 , P1_R1222_U334 , P1_R1222_U331 );
and AND2_13189 ( P1_R1222_U14 , P1_R1222_U325 , P1_R1222_U322 );
and AND2_13190 ( P1_R1222_U15 , P1_R1222_U319 , P1_R1222_U317 );
and AND2_13191 ( P1_R1222_U16 , P1_R1222_U312 , P1_R1222_U309 );
and AND2_13192 ( P1_R1222_U17 , P1_R1222_U234 , P1_R1222_U231 );
and AND2_13193 ( P1_R1222_U18 , P1_R1222_U226 , P1_R1222_U223 );
and AND2_13194 ( P1_R1222_U19 , P1_R1222_U212 , P1_R1222_U209 );
not NOT1_13195 ( P1_R1222_U20 , P1_U3470 );
not NOT1_13196 ( P1_R1222_U21 , P1_U3071 );
not NOT1_13197 ( P1_R1222_U22 , P1_U3070 );
nand NAND2_13198 ( P1_R1222_U23 , P1_U3071 , P1_U3470 );
not NOT1_13199 ( P1_R1222_U24 , P1_U3473 );
not NOT1_13200 ( P1_R1222_U25 , P1_U3464 );
not NOT1_13201 ( P1_R1222_U26 , P1_U3060 );
not NOT1_13202 ( P1_R1222_U27 , P1_U3067 );
not NOT1_13203 ( P1_R1222_U28 , P1_U3458 );
not NOT1_13204 ( P1_R1222_U29 , P1_U3068 );
not NOT1_13205 ( P1_R1222_U30 , P1_U3450 );
not NOT1_13206 ( P1_R1222_U31 , P1_U3077 );
nand NAND2_13207 ( P1_R1222_U32 , P1_U3077 , P1_U3450 );
not NOT1_13208 ( P1_R1222_U33 , P1_U3461 );
not NOT1_13209 ( P1_R1222_U34 , P1_U3064 );
nand NAND2_13210 ( P1_R1222_U35 , P1_U3060 , P1_U3464 );
not NOT1_13211 ( P1_R1222_U36 , P1_U3467 );
not NOT1_13212 ( P1_R1222_U37 , P1_U3476 );
not NOT1_13213 ( P1_R1222_U38 , P1_U3084 );
not NOT1_13214 ( P1_R1222_U39 , P1_U3083 );
not NOT1_13215 ( P1_R1222_U40 , P1_U3479 );
nand NAND2_13216 ( P1_R1222_U41 , P1_R1222_U62 , P1_R1222_U204 );
nand NAND2_13217 ( P1_R1222_U42 , P1_R1222_U118 , P1_R1222_U192 );
nand NAND2_13218 ( P1_R1222_U43 , P1_R1222_U181 , P1_R1222_U182 );
nand NAND2_13219 ( P1_R1222_U44 , P1_U3455 , P1_U3078 );
nand NAND2_13220 ( P1_R1222_U45 , P1_R1222_U122 , P1_R1222_U218 );
nand NAND2_13221 ( P1_R1222_U46 , P1_R1222_U215 , P1_R1222_U214 );
not NOT1_13222 ( P1_R1222_U47 , P1_U3975 );
not NOT1_13223 ( P1_R1222_U48 , P1_U3053 );
not NOT1_13224 ( P1_R1222_U49 , P1_U3057 );
not NOT1_13225 ( P1_R1222_U50 , P1_U3976 );
not NOT1_13226 ( P1_R1222_U51 , P1_U3977 );
not NOT1_13227 ( P1_R1222_U52 , P1_U3058 );
not NOT1_13228 ( P1_R1222_U53 , P1_U3978 );
not NOT1_13229 ( P1_R1222_U54 , P1_U3065 );
not NOT1_13230 ( P1_R1222_U55 , P1_U3981 );
not NOT1_13231 ( P1_R1222_U56 , P1_U3075 );
not NOT1_13232 ( P1_R1222_U57 , P1_U3500 );
not NOT1_13233 ( P1_R1222_U58 , P1_U3073 );
not NOT1_13234 ( P1_R1222_U59 , P1_U3069 );
nand NAND2_13235 ( P1_R1222_U60 , P1_U3073 , P1_U3500 );
not NOT1_13236 ( P1_R1222_U61 , P1_U3503 );
nand NAND2_13237 ( P1_R1222_U62 , P1_U3084 , P1_U3476 );
not NOT1_13238 ( P1_R1222_U63 , P1_U3482 );
not NOT1_13239 ( P1_R1222_U64 , P1_U3062 );
not NOT1_13240 ( P1_R1222_U65 , P1_U3488 );
not NOT1_13241 ( P1_R1222_U66 , P1_U3072 );
not NOT1_13242 ( P1_R1222_U67 , P1_U3485 );
not NOT1_13243 ( P1_R1222_U68 , P1_U3063 );
nand NAND2_13244 ( P1_R1222_U69 , P1_U3063 , P1_U3485 );
not NOT1_13245 ( P1_R1222_U70 , P1_U3491 );
not NOT1_13246 ( P1_R1222_U71 , P1_U3080 );
not NOT1_13247 ( P1_R1222_U72 , P1_U3494 );
not NOT1_13248 ( P1_R1222_U73 , P1_U3079 );
not NOT1_13249 ( P1_R1222_U74 , P1_U3497 );
not NOT1_13250 ( P1_R1222_U75 , P1_U3074 );
not NOT1_13251 ( P1_R1222_U76 , P1_U3506 );
not NOT1_13252 ( P1_R1222_U77 , P1_U3082 );
nand NAND2_13253 ( P1_R1222_U78 , P1_U3082 , P1_U3506 );
not NOT1_13254 ( P1_R1222_U79 , P1_U3508 );
not NOT1_13255 ( P1_R1222_U80 , P1_U3081 );
nand NAND2_13256 ( P1_R1222_U81 , P1_U3081 , P1_U3508 );
not NOT1_13257 ( P1_R1222_U82 , P1_U3982 );
not NOT1_13258 ( P1_R1222_U83 , P1_U3980 );
not NOT1_13259 ( P1_R1222_U84 , P1_U3061 );
not NOT1_13260 ( P1_R1222_U85 , P1_U3979 );
not NOT1_13261 ( P1_R1222_U86 , P1_U3066 );
nand NAND2_13262 ( P1_R1222_U87 , P1_U3976 , P1_U3057 );
not NOT1_13263 ( P1_R1222_U88 , P1_U3054 );
not NOT1_13264 ( P1_R1222_U89 , P1_U3974 );
nand NAND2_13265 ( P1_R1222_U90 , P1_R1222_U305 , P1_R1222_U175 );
not NOT1_13266 ( P1_R1222_U91 , P1_U3076 );
nand NAND2_13267 ( P1_R1222_U92 , P1_R1222_U78 , P1_R1222_U314 );
nand NAND2_13268 ( P1_R1222_U93 , P1_R1222_U260 , P1_R1222_U259 );
nand NAND2_13269 ( P1_R1222_U94 , P1_R1222_U69 , P1_R1222_U336 );
nand NAND2_13270 ( P1_R1222_U95 , P1_R1222_U456 , P1_R1222_U455 );
nand NAND2_13271 ( P1_R1222_U96 , P1_R1222_U503 , P1_R1222_U502 );
nand NAND2_13272 ( P1_R1222_U97 , P1_R1222_U374 , P1_R1222_U373 );
nand NAND2_13273 ( P1_R1222_U98 , P1_R1222_U379 , P1_R1222_U378 );
nand NAND2_13274 ( P1_R1222_U99 , P1_R1222_U386 , P1_R1222_U385 );
nand NAND2_13275 ( P1_R1222_U100 , P1_R1222_U393 , P1_R1222_U392 );
nand NAND2_13276 ( P1_R1222_U101 , P1_R1222_U398 , P1_R1222_U397 );
nand NAND2_13277 ( P1_R1222_U102 , P1_R1222_U407 , P1_R1222_U406 );
nand NAND2_13278 ( P1_R1222_U103 , P1_R1222_U414 , P1_R1222_U413 );
nand NAND2_13279 ( P1_R1222_U104 , P1_R1222_U421 , P1_R1222_U420 );
nand NAND2_13280 ( P1_R1222_U105 , P1_R1222_U428 , P1_R1222_U427 );
nand NAND2_13281 ( P1_R1222_U106 , P1_R1222_U433 , P1_R1222_U432 );
nand NAND2_13282 ( P1_R1222_U107 , P1_R1222_U440 , P1_R1222_U439 );
nand NAND2_13283 ( P1_R1222_U108 , P1_R1222_U447 , P1_R1222_U446 );
nand NAND2_13284 ( P1_R1222_U109 , P1_R1222_U461 , P1_R1222_U460 );
nand NAND2_13285 ( P1_R1222_U110 , P1_R1222_U466 , P1_R1222_U465 );
nand NAND2_13286 ( P1_R1222_U111 , P1_R1222_U473 , P1_R1222_U472 );
nand NAND2_13287 ( P1_R1222_U112 , P1_R1222_U480 , P1_R1222_U479 );
nand NAND2_13288 ( P1_R1222_U113 , P1_R1222_U487 , P1_R1222_U486 );
nand NAND2_13289 ( P1_R1222_U114 , P1_R1222_U494 , P1_R1222_U493 );
nand NAND2_13290 ( P1_R1222_U115 , P1_R1222_U499 , P1_R1222_U498 );
and AND2_13291 ( P1_R1222_U116 , P1_U3458 , P1_U3068 );
and AND2_13292 ( P1_R1222_U117 , P1_R1222_U188 , P1_R1222_U186 );
and AND2_13293 ( P1_R1222_U118 , P1_R1222_U193 , P1_R1222_U191 );
and AND2_13294 ( P1_R1222_U119 , P1_R1222_U200 , P1_R1222_U199 );
and AND3_13295 ( P1_R1222_U120 , P1_R1222_U381 , P1_R1222_U380 , P1_R1222_U23 );
and AND2_13296 ( P1_R1222_U121 , P1_R1222_U211 , P1_R1222_U6 );
and AND2_13297 ( P1_R1222_U122 , P1_R1222_U219 , P1_R1222_U217 );
and AND3_13298 ( P1_R1222_U123 , P1_R1222_U388 , P1_R1222_U387 , P1_R1222_U35 );
and AND2_13299 ( P1_R1222_U124 , P1_R1222_U225 , P1_R1222_U4 );
and AND2_13300 ( P1_R1222_U125 , P1_R1222_U233 , P1_R1222_U180 );
and AND2_13301 ( P1_R1222_U126 , P1_R1222_U203 , P1_R1222_U7 );
and AND2_13302 ( P1_R1222_U127 , P1_R1222_U238 , P1_R1222_U170 );
and AND2_13303 ( P1_R1222_U128 , P1_R1222_U249 , P1_R1222_U8 );
and AND2_13304 ( P1_R1222_U129 , P1_R1222_U247 , P1_R1222_U171 );
and AND2_13305 ( P1_R1222_U130 , P1_R1222_U267 , P1_R1222_U266 );
and AND2_13306 ( P1_R1222_U131 , P1_R1222_U10 , P1_R1222_U281 );
and AND2_13307 ( P1_R1222_U132 , P1_R1222_U284 , P1_R1222_U279 );
and AND2_13308 ( P1_R1222_U133 , P1_R1222_U300 , P1_R1222_U297 );
and AND2_13309 ( P1_R1222_U134 , P1_R1222_U367 , P1_R1222_U301 );
and AND2_13310 ( P1_R1222_U135 , P1_R1222_U159 , P1_R1222_U277 );
and AND3_13311 ( P1_R1222_U136 , P1_R1222_U454 , P1_R1222_U453 , P1_R1222_U81 );
and AND3_13312 ( P1_R1222_U137 , P1_R1222_U468 , P1_R1222_U467 , P1_R1222_U60 );
and AND2_13313 ( P1_R1222_U138 , P1_R1222_U333 , P1_R1222_U9 );
and AND3_13314 ( P1_R1222_U139 , P1_R1222_U489 , P1_R1222_U488 , P1_R1222_U171 );
and AND2_13315 ( P1_R1222_U140 , P1_R1222_U342 , P1_R1222_U8 );
and AND3_13316 ( P1_R1222_U141 , P1_R1222_U501 , P1_R1222_U500 , P1_R1222_U170 );
and AND2_13317 ( P1_R1222_U142 , P1_R1222_U349 , P1_R1222_U7 );
nand NAND2_13318 ( P1_R1222_U143 , P1_R1222_U119 , P1_R1222_U201 );
nand NAND2_13319 ( P1_R1222_U144 , P1_R1222_U216 , P1_R1222_U228 );
not NOT1_13320 ( P1_R1222_U145 , P1_U3055 );
not NOT1_13321 ( P1_R1222_U146 , P1_U3985 );
and AND2_13322 ( P1_R1222_U147 , P1_R1222_U402 , P1_R1222_U401 );
nand NAND3_13323 ( P1_R1222_U148 , P1_R1222_U303 , P1_R1222_U168 , P1_R1222_U363 );
and AND2_13324 ( P1_R1222_U149 , P1_R1222_U409 , P1_R1222_U408 );
nand NAND3_13325 ( P1_R1222_U150 , P1_R1222_U369 , P1_R1222_U368 , P1_R1222_U134 );
and AND2_13326 ( P1_R1222_U151 , P1_R1222_U416 , P1_R1222_U415 );
nand NAND3_13327 ( P1_R1222_U152 , P1_R1222_U364 , P1_R1222_U298 , P1_R1222_U87 );
and AND2_13328 ( P1_R1222_U153 , P1_R1222_U423 , P1_R1222_U422 );
nand NAND2_13329 ( P1_R1222_U154 , P1_R1222_U292 , P1_R1222_U291 );
and AND2_13330 ( P1_R1222_U155 , P1_R1222_U435 , P1_R1222_U434 );
nand NAND2_13331 ( P1_R1222_U156 , P1_R1222_U288 , P1_R1222_U287 );
and AND2_13332 ( P1_R1222_U157 , P1_R1222_U442 , P1_R1222_U441 );
nand NAND2_13333 ( P1_R1222_U158 , P1_R1222_U132 , P1_R1222_U283 );
and AND2_13334 ( P1_R1222_U159 , P1_R1222_U449 , P1_R1222_U448 );
nand NAND2_13335 ( P1_R1222_U160 , P1_R1222_U44 , P1_R1222_U326 );
nand NAND2_13336 ( P1_R1222_U161 , P1_R1222_U130 , P1_R1222_U268 );
and AND2_13337 ( P1_R1222_U162 , P1_R1222_U475 , P1_R1222_U474 );
nand NAND2_13338 ( P1_R1222_U163 , P1_R1222_U256 , P1_R1222_U255 );
and AND2_13339 ( P1_R1222_U164 , P1_R1222_U482 , P1_R1222_U481 );
nand NAND2_13340 ( P1_R1222_U165 , P1_R1222_U252 , P1_R1222_U251 );
nand NAND2_13341 ( P1_R1222_U166 , P1_R1222_U242 , P1_R1222_U241 );
nand NAND2_13342 ( P1_R1222_U167 , P1_R1222_U366 , P1_R1222_U365 );
nand NAND2_13343 ( P1_R1222_U168 , P1_U3054 , P1_R1222_U150 );
not NOT1_13344 ( P1_R1222_U169 , P1_R1222_U35 );
nand NAND2_13345 ( P1_R1222_U170 , P1_U3479 , P1_U3083 );
nand NAND2_13346 ( P1_R1222_U171 , P1_U3072 , P1_U3488 );
nand NAND2_13347 ( P1_R1222_U172 , P1_U3058 , P1_U3977 );
not NOT1_13348 ( P1_R1222_U173 , P1_R1222_U69 );
not NOT1_13349 ( P1_R1222_U174 , P1_R1222_U78 );
nand NAND2_13350 ( P1_R1222_U175 , P1_U3065 , P1_U3978 );
not NOT1_13351 ( P1_R1222_U176 , P1_R1222_U62 );
or OR2_13352 ( P1_R1222_U177 , P1_U3067 , P1_U3467 );
or OR2_13353 ( P1_R1222_U178 , P1_U3060 , P1_U3464 );
or OR2_13354 ( P1_R1222_U179 , P1_U3461 , P1_U3064 );
or OR2_13355 ( P1_R1222_U180 , P1_U3458 , P1_U3068 );
not NOT1_13356 ( P1_R1222_U181 , P1_R1222_U32 );
or OR2_13357 ( P1_R1222_U182 , P1_U3455 , P1_U3078 );
not NOT1_13358 ( P1_R1222_U183 , P1_R1222_U43 );
not NOT1_13359 ( P1_R1222_U184 , P1_R1222_U44 );
nand NAND2_13360 ( P1_R1222_U185 , P1_R1222_U43 , P1_R1222_U44 );
nand NAND2_13361 ( P1_R1222_U186 , P1_R1222_U116 , P1_R1222_U179 );
nand NAND2_13362 ( P1_R1222_U187 , P1_R1222_U5 , P1_R1222_U185 );
nand NAND2_13363 ( P1_R1222_U188 , P1_U3064 , P1_U3461 );
nand NAND2_13364 ( P1_R1222_U189 , P1_R1222_U117 , P1_R1222_U187 );
nand NAND2_13365 ( P1_R1222_U190 , P1_R1222_U36 , P1_R1222_U35 );
nand NAND2_13366 ( P1_R1222_U191 , P1_U3067 , P1_R1222_U190 );
nand NAND2_13367 ( P1_R1222_U192 , P1_R1222_U4 , P1_R1222_U189 );
nand NAND2_13368 ( P1_R1222_U193 , P1_U3467 , P1_R1222_U169 );
not NOT1_13369 ( P1_R1222_U194 , P1_R1222_U42 );
or OR2_13370 ( P1_R1222_U195 , P1_U3070 , P1_U3473 );
or OR2_13371 ( P1_R1222_U196 , P1_U3071 , P1_U3470 );
not NOT1_13372 ( P1_R1222_U197 , P1_R1222_U23 );
nand NAND2_13373 ( P1_R1222_U198 , P1_R1222_U24 , P1_R1222_U23 );
nand NAND2_13374 ( P1_R1222_U199 , P1_U3070 , P1_R1222_U198 );
nand NAND2_13375 ( P1_R1222_U200 , P1_U3473 , P1_R1222_U197 );
nand NAND2_13376 ( P1_R1222_U201 , P1_R1222_U6 , P1_R1222_U42 );
not NOT1_13377 ( P1_R1222_U202 , P1_R1222_U143 );
or OR2_13378 ( P1_R1222_U203 , P1_U3476 , P1_U3084 );
nand NAND2_13379 ( P1_R1222_U204 , P1_R1222_U203 , P1_R1222_U143 );
not NOT1_13380 ( P1_R1222_U205 , P1_R1222_U41 );
or OR2_13381 ( P1_R1222_U206 , P1_U3083 , P1_U3479 );
or OR2_13382 ( P1_R1222_U207 , P1_U3470 , P1_U3071 );
nand NAND2_13383 ( P1_R1222_U208 , P1_R1222_U207 , P1_R1222_U42 );
nand NAND2_13384 ( P1_R1222_U209 , P1_R1222_U120 , P1_R1222_U208 );
nand NAND2_13385 ( P1_R1222_U210 , P1_R1222_U194 , P1_R1222_U23 );
nand NAND2_13386 ( P1_R1222_U211 , P1_U3473 , P1_U3070 );
nand NAND2_13387 ( P1_R1222_U212 , P1_R1222_U121 , P1_R1222_U210 );
or OR2_13388 ( P1_R1222_U213 , P1_U3071 , P1_U3470 );
nand NAND2_13389 ( P1_R1222_U214 , P1_R1222_U184 , P1_R1222_U180 );
nand NAND2_13390 ( P1_R1222_U215 , P1_U3068 , P1_U3458 );
not NOT1_13391 ( P1_R1222_U216 , P1_R1222_U46 );
nand NAND2_13392 ( P1_R1222_U217 , P1_R1222_U183 , P1_R1222_U5 );
nand NAND2_13393 ( P1_R1222_U218 , P1_R1222_U46 , P1_R1222_U179 );
nand NAND2_13394 ( P1_R1222_U219 , P1_U3064 , P1_U3461 );
not NOT1_13395 ( P1_R1222_U220 , P1_R1222_U45 );
or OR2_13396 ( P1_R1222_U221 , P1_U3464 , P1_U3060 );
nand NAND2_13397 ( P1_R1222_U222 , P1_R1222_U221 , P1_R1222_U45 );
nand NAND2_13398 ( P1_R1222_U223 , P1_R1222_U123 , P1_R1222_U222 );
nand NAND2_13399 ( P1_R1222_U224 , P1_R1222_U220 , P1_R1222_U35 );
nand NAND2_13400 ( P1_R1222_U225 , P1_U3467 , P1_U3067 );
nand NAND2_13401 ( P1_R1222_U226 , P1_R1222_U124 , P1_R1222_U224 );
or OR2_13402 ( P1_R1222_U227 , P1_U3060 , P1_U3464 );
nand NAND2_13403 ( P1_R1222_U228 , P1_R1222_U183 , P1_R1222_U180 );
not NOT1_13404 ( P1_R1222_U229 , P1_R1222_U144 );
nand NAND2_13405 ( P1_R1222_U230 , P1_U3064 , P1_U3461 );
nand NAND4_13406 ( P1_R1222_U231 , P1_R1222_U400 , P1_R1222_U399 , P1_R1222_U44 , P1_R1222_U43 );
nand NAND2_13407 ( P1_R1222_U232 , P1_R1222_U44 , P1_R1222_U43 );
nand NAND2_13408 ( P1_R1222_U233 , P1_U3068 , P1_U3458 );
nand NAND2_13409 ( P1_R1222_U234 , P1_R1222_U125 , P1_R1222_U232 );
or OR2_13410 ( P1_R1222_U235 , P1_U3083 , P1_U3479 );
or OR2_13411 ( P1_R1222_U236 , P1_U3062 , P1_U3482 );
nand NAND2_13412 ( P1_R1222_U237 , P1_R1222_U176 , P1_R1222_U7 );
nand NAND2_13413 ( P1_R1222_U238 , P1_U3062 , P1_U3482 );
nand NAND2_13414 ( P1_R1222_U239 , P1_R1222_U127 , P1_R1222_U237 );
or OR2_13415 ( P1_R1222_U240 , P1_U3482 , P1_U3062 );
nand NAND2_13416 ( P1_R1222_U241 , P1_R1222_U126 , P1_R1222_U143 );
nand NAND2_13417 ( P1_R1222_U242 , P1_R1222_U240 , P1_R1222_U239 );
not NOT1_13418 ( P1_R1222_U243 , P1_R1222_U166 );
or OR2_13419 ( P1_R1222_U244 , P1_U3080 , P1_U3491 );
or OR2_13420 ( P1_R1222_U245 , P1_U3072 , P1_U3488 );
nand NAND2_13421 ( P1_R1222_U246 , P1_R1222_U173 , P1_R1222_U8 );
nand NAND2_13422 ( P1_R1222_U247 , P1_U3080 , P1_U3491 );
nand NAND2_13423 ( P1_R1222_U248 , P1_R1222_U129 , P1_R1222_U246 );
or OR2_13424 ( P1_R1222_U249 , P1_U3485 , P1_U3063 );
or OR2_13425 ( P1_R1222_U250 , P1_U3491 , P1_U3080 );
nand NAND2_13426 ( P1_R1222_U251 , P1_R1222_U128 , P1_R1222_U166 );
nand NAND2_13427 ( P1_R1222_U252 , P1_R1222_U250 , P1_R1222_U248 );
not NOT1_13428 ( P1_R1222_U253 , P1_R1222_U165 );
or OR2_13429 ( P1_R1222_U254 , P1_U3494 , P1_U3079 );
nand NAND2_13430 ( P1_R1222_U255 , P1_R1222_U254 , P1_R1222_U165 );
nand NAND2_13431 ( P1_R1222_U256 , P1_U3079 , P1_U3494 );
not NOT1_13432 ( P1_R1222_U257 , P1_R1222_U163 );
or OR2_13433 ( P1_R1222_U258 , P1_U3497 , P1_U3074 );
nand NAND2_13434 ( P1_R1222_U259 , P1_R1222_U258 , P1_R1222_U163 );
nand NAND2_13435 ( P1_R1222_U260 , P1_U3074 , P1_U3497 );
not NOT1_13436 ( P1_R1222_U261 , P1_R1222_U93 );
or OR2_13437 ( P1_R1222_U262 , P1_U3069 , P1_U3503 );
or OR2_13438 ( P1_R1222_U263 , P1_U3073 , P1_U3500 );
not NOT1_13439 ( P1_R1222_U264 , P1_R1222_U60 );
nand NAND2_13440 ( P1_R1222_U265 , P1_R1222_U61 , P1_R1222_U60 );
nand NAND2_13441 ( P1_R1222_U266 , P1_U3069 , P1_R1222_U265 );
nand NAND2_13442 ( P1_R1222_U267 , P1_U3503 , P1_R1222_U264 );
nand NAND2_13443 ( P1_R1222_U268 , P1_R1222_U9 , P1_R1222_U93 );
not NOT1_13444 ( P1_R1222_U269 , P1_R1222_U161 );
or OR2_13445 ( P1_R1222_U270 , P1_U3076 , P1_U3982 );
or OR2_13446 ( P1_R1222_U271 , P1_U3081 , P1_U3508 );
or OR2_13447 ( P1_R1222_U272 , P1_U3075 , P1_U3981 );
not NOT1_13448 ( P1_R1222_U273 , P1_R1222_U81 );
nand NAND2_13449 ( P1_R1222_U274 , P1_U3982 , P1_R1222_U273 );
nand NAND2_13450 ( P1_R1222_U275 , P1_R1222_U274 , P1_R1222_U91 );
nand NAND2_13451 ( P1_R1222_U276 , P1_R1222_U81 , P1_R1222_U82 );
nand NAND2_13452 ( P1_R1222_U277 , P1_R1222_U276 , P1_R1222_U275 );
nand NAND2_13453 ( P1_R1222_U278 , P1_R1222_U174 , P1_R1222_U10 );
nand NAND2_13454 ( P1_R1222_U279 , P1_U3075 , P1_U3981 );
nand NAND2_13455 ( P1_R1222_U280 , P1_R1222_U277 , P1_R1222_U278 );
or OR2_13456 ( P1_R1222_U281 , P1_U3506 , P1_U3082 );
or OR2_13457 ( P1_R1222_U282 , P1_U3981 , P1_U3075 );
nand NAND3_13458 ( P1_R1222_U283 , P1_R1222_U272 , P1_R1222_U161 , P1_R1222_U131 );
nand NAND2_13459 ( P1_R1222_U284 , P1_R1222_U282 , P1_R1222_U280 );
not NOT1_13460 ( P1_R1222_U285 , P1_R1222_U158 );
or OR2_13461 ( P1_R1222_U286 , P1_U3980 , P1_U3061 );
nand NAND2_13462 ( P1_R1222_U287 , P1_R1222_U286 , P1_R1222_U158 );
nand NAND2_13463 ( P1_R1222_U288 , P1_U3061 , P1_U3980 );
not NOT1_13464 ( P1_R1222_U289 , P1_R1222_U156 );
or OR2_13465 ( P1_R1222_U290 , P1_U3979 , P1_U3066 );
nand NAND2_13466 ( P1_R1222_U291 , P1_R1222_U290 , P1_R1222_U156 );
nand NAND2_13467 ( P1_R1222_U292 , P1_U3066 , P1_U3979 );
not NOT1_13468 ( P1_R1222_U293 , P1_R1222_U154 );
or OR2_13469 ( P1_R1222_U294 , P1_U3058 , P1_U3977 );
nand NAND2_13470 ( P1_R1222_U295 , P1_R1222_U175 , P1_R1222_U172 );
not NOT1_13471 ( P1_R1222_U296 , P1_R1222_U87 );
or OR2_13472 ( P1_R1222_U297 , P1_U3978 , P1_U3065 );
nand NAND3_13473 ( P1_R1222_U298 , P1_R1222_U154 , P1_R1222_U297 , P1_R1222_U167 );
not NOT1_13474 ( P1_R1222_U299 , P1_R1222_U152 );
or OR2_13475 ( P1_R1222_U300 , P1_U3975 , P1_U3053 );
nand NAND2_13476 ( P1_R1222_U301 , P1_U3053 , P1_U3975 );
not NOT1_13477 ( P1_R1222_U302 , P1_R1222_U150 );
nand NAND2_13478 ( P1_R1222_U303 , P1_U3974 , P1_R1222_U150 );
not NOT1_13479 ( P1_R1222_U304 , P1_R1222_U148 );
nand NAND2_13480 ( P1_R1222_U305 , P1_R1222_U297 , P1_R1222_U154 );
not NOT1_13481 ( P1_R1222_U306 , P1_R1222_U90 );
or OR2_13482 ( P1_R1222_U307 , P1_U3977 , P1_U3058 );
nand NAND2_13483 ( P1_R1222_U308 , P1_R1222_U307 , P1_R1222_U90 );
nand NAND3_13484 ( P1_R1222_U309 , P1_R1222_U308 , P1_R1222_U172 , P1_R1222_U153 );
nand NAND2_13485 ( P1_R1222_U310 , P1_R1222_U306 , P1_R1222_U172 );
nand NAND2_13486 ( P1_R1222_U311 , P1_U3976 , P1_U3057 );
nand NAND3_13487 ( P1_R1222_U312 , P1_R1222_U310 , P1_R1222_U311 , P1_R1222_U167 );
or OR2_13488 ( P1_R1222_U313 , P1_U3058 , P1_U3977 );
nand NAND2_13489 ( P1_R1222_U314 , P1_R1222_U281 , P1_R1222_U161 );
not NOT1_13490 ( P1_R1222_U315 , P1_R1222_U92 );
nand NAND2_13491 ( P1_R1222_U316 , P1_R1222_U10 , P1_R1222_U92 );
nand NAND2_13492 ( P1_R1222_U317 , P1_R1222_U135 , P1_R1222_U316 );
nand NAND2_13493 ( P1_R1222_U318 , P1_R1222_U316 , P1_R1222_U277 );
nand NAND2_13494 ( P1_R1222_U319 , P1_R1222_U452 , P1_R1222_U318 );
or OR2_13495 ( P1_R1222_U320 , P1_U3508 , P1_U3081 );
nand NAND2_13496 ( P1_R1222_U321 , P1_R1222_U320 , P1_R1222_U92 );
nand NAND2_13497 ( P1_R1222_U322 , P1_R1222_U136 , P1_R1222_U321 );
nand NAND2_13498 ( P1_R1222_U323 , P1_R1222_U315 , P1_R1222_U81 );
nand NAND2_13499 ( P1_R1222_U324 , P1_U3076 , P1_U3982 );
nand NAND3_13500 ( P1_R1222_U325 , P1_R1222_U324 , P1_R1222_U323 , P1_R1222_U10 );
or OR2_13501 ( P1_R1222_U326 , P1_U3455 , P1_U3078 );
not NOT1_13502 ( P1_R1222_U327 , P1_R1222_U160 );
or OR2_13503 ( P1_R1222_U328 , P1_U3081 , P1_U3508 );
or OR2_13504 ( P1_R1222_U329 , P1_U3500 , P1_U3073 );
nand NAND2_13505 ( P1_R1222_U330 , P1_R1222_U329 , P1_R1222_U93 );
nand NAND2_13506 ( P1_R1222_U331 , P1_R1222_U137 , P1_R1222_U330 );
nand NAND2_13507 ( P1_R1222_U332 , P1_R1222_U261 , P1_R1222_U60 );
nand NAND2_13508 ( P1_R1222_U333 , P1_U3503 , P1_U3069 );
nand NAND2_13509 ( P1_R1222_U334 , P1_R1222_U138 , P1_R1222_U332 );
or OR2_13510 ( P1_R1222_U335 , P1_U3073 , P1_U3500 );
nand NAND2_13511 ( P1_R1222_U336 , P1_R1222_U249 , P1_R1222_U166 );
not NOT1_13512 ( P1_R1222_U337 , P1_R1222_U94 );
or OR2_13513 ( P1_R1222_U338 , P1_U3488 , P1_U3072 );
nand NAND2_13514 ( P1_R1222_U339 , P1_R1222_U338 , P1_R1222_U94 );
nand NAND2_13515 ( P1_R1222_U340 , P1_R1222_U139 , P1_R1222_U339 );
nand NAND2_13516 ( P1_R1222_U341 , P1_R1222_U337 , P1_R1222_U171 );
nand NAND2_13517 ( P1_R1222_U342 , P1_U3080 , P1_U3491 );
nand NAND2_13518 ( P1_R1222_U343 , P1_R1222_U140 , P1_R1222_U341 );
or OR2_13519 ( P1_R1222_U344 , P1_U3072 , P1_U3488 );
or OR2_13520 ( P1_R1222_U345 , P1_U3479 , P1_U3083 );
nand NAND2_13521 ( P1_R1222_U346 , P1_R1222_U345 , P1_R1222_U41 );
nand NAND2_13522 ( P1_R1222_U347 , P1_R1222_U141 , P1_R1222_U346 );
nand NAND2_13523 ( P1_R1222_U348 , P1_R1222_U205 , P1_R1222_U170 );
nand NAND2_13524 ( P1_R1222_U349 , P1_U3062 , P1_U3482 );
nand NAND2_13525 ( P1_R1222_U350 , P1_R1222_U142 , P1_R1222_U348 );
nand NAND2_13526 ( P1_R1222_U351 , P1_R1222_U206 , P1_R1222_U170 );
nand NAND2_13527 ( P1_R1222_U352 , P1_R1222_U203 , P1_R1222_U62 );
nand NAND2_13528 ( P1_R1222_U353 , P1_R1222_U213 , P1_R1222_U23 );
nand NAND2_13529 ( P1_R1222_U354 , P1_R1222_U227 , P1_R1222_U35 );
nand NAND2_13530 ( P1_R1222_U355 , P1_R1222_U230 , P1_R1222_U179 );
nand NAND2_13531 ( P1_R1222_U356 , P1_R1222_U313 , P1_R1222_U172 );
nand NAND2_13532 ( P1_R1222_U357 , P1_R1222_U297 , P1_R1222_U175 );
nand NAND2_13533 ( P1_R1222_U358 , P1_R1222_U328 , P1_R1222_U81 );
nand NAND2_13534 ( P1_R1222_U359 , P1_R1222_U281 , P1_R1222_U78 );
nand NAND2_13535 ( P1_R1222_U360 , P1_R1222_U335 , P1_R1222_U60 );
nand NAND2_13536 ( P1_R1222_U361 , P1_R1222_U344 , P1_R1222_U171 );
nand NAND2_13537 ( P1_R1222_U362 , P1_R1222_U249 , P1_R1222_U69 );
nand NAND2_13538 ( P1_R1222_U363 , P1_U3974 , P1_U3054 );
nand NAND2_13539 ( P1_R1222_U364 , P1_R1222_U295 , P1_R1222_U167 );
nand NAND2_13540 ( P1_R1222_U365 , P1_U3057 , P1_R1222_U294 );
nand NAND2_13541 ( P1_R1222_U366 , P1_U3976 , P1_R1222_U294 );
nand NAND3_13542 ( P1_R1222_U367 , P1_R1222_U295 , P1_R1222_U167 , P1_R1222_U300 );
nand NAND3_13543 ( P1_R1222_U368 , P1_R1222_U154 , P1_R1222_U167 , P1_R1222_U133 );
nand NAND2_13544 ( P1_R1222_U369 , P1_R1222_U296 , P1_R1222_U300 );
nand NAND2_13545 ( P1_R1222_U370 , P1_U3083 , P1_R1222_U40 );
nand NAND2_13546 ( P1_R1222_U371 , P1_U3479 , P1_R1222_U39 );
nand NAND2_13547 ( P1_R1222_U372 , P1_R1222_U371 , P1_R1222_U370 );
nand NAND2_13548 ( P1_R1222_U373 , P1_R1222_U351 , P1_R1222_U41 );
nand NAND2_13549 ( P1_R1222_U374 , P1_R1222_U372 , P1_R1222_U205 );
nand NAND2_13550 ( P1_R1222_U375 , P1_U3084 , P1_R1222_U37 );
nand NAND2_13551 ( P1_R1222_U376 , P1_U3476 , P1_R1222_U38 );
nand NAND2_13552 ( P1_R1222_U377 , P1_R1222_U376 , P1_R1222_U375 );
nand NAND2_13553 ( P1_R1222_U378 , P1_R1222_U352 , P1_R1222_U143 );
nand NAND2_13554 ( P1_R1222_U379 , P1_R1222_U202 , P1_R1222_U377 );
nand NAND2_13555 ( P1_R1222_U380 , P1_U3070 , P1_R1222_U24 );
nand NAND2_13556 ( P1_R1222_U381 , P1_U3473 , P1_R1222_U22 );
nand NAND2_13557 ( P1_R1222_U382 , P1_U3071 , P1_R1222_U20 );
nand NAND2_13558 ( P1_R1222_U383 , P1_U3470 , P1_R1222_U21 );
nand NAND2_13559 ( P1_R1222_U384 , P1_R1222_U383 , P1_R1222_U382 );
nand NAND2_13560 ( P1_R1222_U385 , P1_R1222_U353 , P1_R1222_U42 );
nand NAND2_13561 ( P1_R1222_U386 , P1_R1222_U384 , P1_R1222_U194 );
nand NAND2_13562 ( P1_R1222_U387 , P1_U3067 , P1_R1222_U36 );
nand NAND2_13563 ( P1_R1222_U388 , P1_U3467 , P1_R1222_U27 );
nand NAND2_13564 ( P1_R1222_U389 , P1_U3060 , P1_R1222_U25 );
nand NAND2_13565 ( P1_R1222_U390 , P1_U3464 , P1_R1222_U26 );
nand NAND2_13566 ( P1_R1222_U391 , P1_R1222_U390 , P1_R1222_U389 );
nand NAND2_13567 ( P1_R1222_U392 , P1_R1222_U354 , P1_R1222_U45 );
nand NAND2_13568 ( P1_R1222_U393 , P1_R1222_U391 , P1_R1222_U220 );
nand NAND2_13569 ( P1_R1222_U394 , P1_U3064 , P1_R1222_U33 );
nand NAND2_13570 ( P1_R1222_U395 , P1_U3461 , P1_R1222_U34 );
nand NAND2_13571 ( P1_R1222_U396 , P1_R1222_U395 , P1_R1222_U394 );
nand NAND2_13572 ( P1_R1222_U397 , P1_R1222_U355 , P1_R1222_U144 );
nand NAND2_13573 ( P1_R1222_U398 , P1_R1222_U229 , P1_R1222_U396 );
nand NAND2_13574 ( P1_R1222_U399 , P1_U3068 , P1_R1222_U28 );
nand NAND2_13575 ( P1_R1222_U400 , P1_U3458 , P1_R1222_U29 );
nand NAND2_13576 ( P1_R1222_U401 , P1_U3055 , P1_R1222_U146 );
nand NAND2_13577 ( P1_R1222_U402 , P1_U3985 , P1_R1222_U145 );
nand NAND2_13578 ( P1_R1222_U403 , P1_U3055 , P1_R1222_U146 );
nand NAND2_13579 ( P1_R1222_U404 , P1_U3985 , P1_R1222_U145 );
nand NAND2_13580 ( P1_R1222_U405 , P1_R1222_U404 , P1_R1222_U403 );
nand NAND2_13581 ( P1_R1222_U406 , P1_R1222_U147 , P1_R1222_U148 );
nand NAND2_13582 ( P1_R1222_U407 , P1_R1222_U304 , P1_R1222_U405 );
nand NAND2_13583 ( P1_R1222_U408 , P1_U3054 , P1_R1222_U89 );
nand NAND2_13584 ( P1_R1222_U409 , P1_U3974 , P1_R1222_U88 );
nand NAND2_13585 ( P1_R1222_U410 , P1_U3054 , P1_R1222_U89 );
nand NAND2_13586 ( P1_R1222_U411 , P1_U3974 , P1_R1222_U88 );
nand NAND2_13587 ( P1_R1222_U412 , P1_R1222_U411 , P1_R1222_U410 );
nand NAND2_13588 ( P1_R1222_U413 , P1_R1222_U149 , P1_R1222_U150 );
nand NAND2_13589 ( P1_R1222_U414 , P1_R1222_U302 , P1_R1222_U412 );
nand NAND2_13590 ( P1_R1222_U415 , P1_U3053 , P1_R1222_U47 );
nand NAND2_13591 ( P1_R1222_U416 , P1_U3975 , P1_R1222_U48 );
nand NAND2_13592 ( P1_R1222_U417 , P1_U3053 , P1_R1222_U47 );
nand NAND2_13593 ( P1_R1222_U418 , P1_U3975 , P1_R1222_U48 );
nand NAND2_13594 ( P1_R1222_U419 , P1_R1222_U418 , P1_R1222_U417 );
nand NAND2_13595 ( P1_R1222_U420 , P1_R1222_U151 , P1_R1222_U152 );
nand NAND2_13596 ( P1_R1222_U421 , P1_R1222_U299 , P1_R1222_U419 );
nand NAND2_13597 ( P1_R1222_U422 , P1_U3057 , P1_R1222_U50 );
nand NAND2_13598 ( P1_R1222_U423 , P1_U3976 , P1_R1222_U49 );
nand NAND2_13599 ( P1_R1222_U424 , P1_U3058 , P1_R1222_U51 );
nand NAND2_13600 ( P1_R1222_U425 , P1_U3977 , P1_R1222_U52 );
nand NAND2_13601 ( P1_R1222_U426 , P1_R1222_U425 , P1_R1222_U424 );
nand NAND2_13602 ( P1_R1222_U427 , P1_R1222_U356 , P1_R1222_U90 );
nand NAND2_13603 ( P1_R1222_U428 , P1_R1222_U426 , P1_R1222_U306 );
nand NAND2_13604 ( P1_R1222_U429 , P1_U3065 , P1_R1222_U53 );
nand NAND2_13605 ( P1_R1222_U430 , P1_U3978 , P1_R1222_U54 );
nand NAND2_13606 ( P1_R1222_U431 , P1_R1222_U430 , P1_R1222_U429 );
nand NAND2_13607 ( P1_R1222_U432 , P1_R1222_U357 , P1_R1222_U154 );
nand NAND2_13608 ( P1_R1222_U433 , P1_R1222_U293 , P1_R1222_U431 );
nand NAND2_13609 ( P1_R1222_U434 , P1_U3066 , P1_R1222_U85 );
nand NAND2_13610 ( P1_R1222_U435 , P1_U3979 , P1_R1222_U86 );
nand NAND2_13611 ( P1_R1222_U436 , P1_U3066 , P1_R1222_U85 );
nand NAND2_13612 ( P1_R1222_U437 , P1_U3979 , P1_R1222_U86 );
nand NAND2_13613 ( P1_R1222_U438 , P1_R1222_U437 , P1_R1222_U436 );
nand NAND2_13614 ( P1_R1222_U439 , P1_R1222_U155 , P1_R1222_U156 );
nand NAND2_13615 ( P1_R1222_U440 , P1_R1222_U289 , P1_R1222_U438 );
nand NAND2_13616 ( P1_R1222_U441 , P1_U3061 , P1_R1222_U83 );
nand NAND2_13617 ( P1_R1222_U442 , P1_U3980 , P1_R1222_U84 );
nand NAND2_13618 ( P1_R1222_U443 , P1_U3061 , P1_R1222_U83 );
nand NAND2_13619 ( P1_R1222_U444 , P1_U3980 , P1_R1222_U84 );
nand NAND2_13620 ( P1_R1222_U445 , P1_R1222_U444 , P1_R1222_U443 );
nand NAND2_13621 ( P1_R1222_U446 , P1_R1222_U157 , P1_R1222_U158 );
nand NAND2_13622 ( P1_R1222_U447 , P1_R1222_U285 , P1_R1222_U445 );
nand NAND2_13623 ( P1_R1222_U448 , P1_U3075 , P1_R1222_U55 );
nand NAND2_13624 ( P1_R1222_U449 , P1_U3981 , P1_R1222_U56 );
nand NAND2_13625 ( P1_R1222_U450 , P1_U3075 , P1_R1222_U55 );
nand NAND2_13626 ( P1_R1222_U451 , P1_U3981 , P1_R1222_U56 );
nand NAND2_13627 ( P1_R1222_U452 , P1_R1222_U451 , P1_R1222_U450 );
nand NAND2_13628 ( P1_R1222_U453 , P1_U3076 , P1_R1222_U82 );
nand NAND2_13629 ( P1_R1222_U454 , P1_U3982 , P1_R1222_U91 );
nand NAND2_13630 ( P1_R1222_U455 , P1_R1222_U181 , P1_R1222_U160 );
nand NAND2_13631 ( P1_R1222_U456 , P1_R1222_U327 , P1_R1222_U32 );
nand NAND2_13632 ( P1_R1222_U457 , P1_U3081 , P1_R1222_U79 );
nand NAND2_13633 ( P1_R1222_U458 , P1_U3508 , P1_R1222_U80 );
nand NAND2_13634 ( P1_R1222_U459 , P1_R1222_U458 , P1_R1222_U457 );
nand NAND2_13635 ( P1_R1222_U460 , P1_R1222_U358 , P1_R1222_U92 );
nand NAND2_13636 ( P1_R1222_U461 , P1_R1222_U459 , P1_R1222_U315 );
nand NAND2_13637 ( P1_R1222_U462 , P1_U3082 , P1_R1222_U76 );
nand NAND2_13638 ( P1_R1222_U463 , P1_U3506 , P1_R1222_U77 );
nand NAND2_13639 ( P1_R1222_U464 , P1_R1222_U463 , P1_R1222_U462 );
nand NAND2_13640 ( P1_R1222_U465 , P1_R1222_U359 , P1_R1222_U161 );
nand NAND2_13641 ( P1_R1222_U466 , P1_R1222_U269 , P1_R1222_U464 );
nand NAND2_13642 ( P1_R1222_U467 , P1_U3069 , P1_R1222_U61 );
nand NAND2_13643 ( P1_R1222_U468 , P1_U3503 , P1_R1222_U59 );
nand NAND2_13644 ( P1_R1222_U469 , P1_U3073 , P1_R1222_U57 );
nand NAND2_13645 ( P1_R1222_U470 , P1_U3500 , P1_R1222_U58 );
nand NAND2_13646 ( P1_R1222_U471 , P1_R1222_U470 , P1_R1222_U469 );
nand NAND2_13647 ( P1_R1222_U472 , P1_R1222_U360 , P1_R1222_U93 );
nand NAND2_13648 ( P1_R1222_U473 , P1_R1222_U471 , P1_R1222_U261 );
nand NAND2_13649 ( P1_R1222_U474 , P1_U3074 , P1_R1222_U74 );
nand NAND2_13650 ( P1_R1222_U475 , P1_U3497 , P1_R1222_U75 );
nand NAND2_13651 ( P1_R1222_U476 , P1_U3074 , P1_R1222_U74 );
nand NAND2_13652 ( P1_R1222_U477 , P1_U3497 , P1_R1222_U75 );
nand NAND2_13653 ( P1_R1222_U478 , P1_R1222_U477 , P1_R1222_U476 );
nand NAND2_13654 ( P1_R1222_U479 , P1_R1222_U162 , P1_R1222_U163 );
nand NAND2_13655 ( P1_R1222_U480 , P1_R1222_U257 , P1_R1222_U478 );
nand NAND2_13656 ( P1_R1222_U481 , P1_U3079 , P1_R1222_U72 );
nand NAND2_13657 ( P1_R1222_U482 , P1_U3494 , P1_R1222_U73 );
nand NAND2_13658 ( P1_R1222_U483 , P1_U3079 , P1_R1222_U72 );
nand NAND2_13659 ( P1_R1222_U484 , P1_U3494 , P1_R1222_U73 );
nand NAND2_13660 ( P1_R1222_U485 , P1_R1222_U484 , P1_R1222_U483 );
nand NAND2_13661 ( P1_R1222_U486 , P1_R1222_U164 , P1_R1222_U165 );
nand NAND2_13662 ( P1_R1222_U487 , P1_R1222_U253 , P1_R1222_U485 );
nand NAND2_13663 ( P1_R1222_U488 , P1_U3080 , P1_R1222_U70 );
nand NAND2_13664 ( P1_R1222_U489 , P1_U3491 , P1_R1222_U71 );
nand NAND2_13665 ( P1_R1222_U490 , P1_U3072 , P1_R1222_U65 );
nand NAND2_13666 ( P1_R1222_U491 , P1_U3488 , P1_R1222_U66 );
nand NAND2_13667 ( P1_R1222_U492 , P1_R1222_U491 , P1_R1222_U490 );
nand NAND2_13668 ( P1_R1222_U493 , P1_R1222_U361 , P1_R1222_U94 );
nand NAND2_13669 ( P1_R1222_U494 , P1_R1222_U492 , P1_R1222_U337 );
nand NAND2_13670 ( P1_R1222_U495 , P1_U3063 , P1_R1222_U67 );
nand NAND2_13671 ( P1_R1222_U496 , P1_U3485 , P1_R1222_U68 );
nand NAND2_13672 ( P1_R1222_U497 , P1_R1222_U496 , P1_R1222_U495 );
nand NAND2_13673 ( P1_R1222_U498 , P1_R1222_U362 , P1_R1222_U166 );
nand NAND2_13674 ( P1_R1222_U499 , P1_R1222_U243 , P1_R1222_U497 );
nand NAND2_13675 ( P1_R1222_U500 , P1_U3062 , P1_R1222_U63 );
nand NAND2_13676 ( P1_R1222_U501 , P1_U3482 , P1_R1222_U64 );
nand NAND2_13677 ( P1_R1222_U502 , P1_U3077 , P1_R1222_U30 );
nand NAND2_13678 ( P1_R1222_U503 , P1_U3450 , P1_R1222_U31 );
nor nor_13679 ( P2_SUB_594_U6 , P2_IR_REG_12_ , P2_IR_REG_9_ , P2_IR_REG_10_ , P2_IR_REG_11_ );
nor nor_13680 ( P2_SUB_594_U7 , P2_IR_REG_19_ , P2_IR_REG_20_ , P2_IR_REG_17_ , P2_IR_REG_18_ );
and AND2_13681 ( P2_SUB_594_U8 , P2_SUB_594_U135 , P2_SUB_594_U51 );
and AND2_13682 ( P2_SUB_594_U9 , P2_SUB_594_U133 , P2_SUB_594_U101 );
and AND2_13683 ( P2_SUB_594_U10 , P2_SUB_594_U132 , P2_SUB_594_U47 );
and AND2_13684 ( P2_SUB_594_U11 , P2_SUB_594_U131 , P2_SUB_594_U48 );
and AND2_13685 ( P2_SUB_594_U12 , P2_SUB_594_U129 , P2_SUB_594_U104 );
and AND2_13686 ( P2_SUB_594_U13 , P2_SUB_594_U128 , P2_SUB_594_U35 );
and AND2_13687 ( P2_SUB_594_U14 , P2_SUB_594_U127 , P2_SUB_594_U45 );
and AND2_13688 ( P2_SUB_594_U15 , P2_SUB_594_U125 , P2_SUB_594_U107 );
and AND2_13689 ( P2_SUB_594_U16 , P2_SUB_594_U124 , P2_SUB_594_U41 );
and AND2_13690 ( P2_SUB_594_U17 , P2_SUB_594_U123 , P2_SUB_594_U42 );
and AND2_13691 ( P2_SUB_594_U18 , P2_SUB_594_U121 , P2_SUB_594_U110 );
and AND2_13692 ( P2_SUB_594_U19 , P2_SUB_594_U120 , P2_SUB_594_U36 );
and AND2_13693 ( P2_SUB_594_U20 , P2_SUB_594_U119 , P2_SUB_594_U76 );
and AND2_13694 ( P2_SUB_594_U21 , P2_SUB_594_U64 , P2_SUB_594_U138 );
and AND2_13695 ( P2_SUB_594_U22 , P2_SUB_594_U117 , P2_SUB_594_U38 );
and AND2_13696 ( P2_SUB_594_U23 , P2_SUB_594_U116 , P2_SUB_594_U33 );
and AND2_13697 ( P2_SUB_594_U24 , P2_SUB_594_U99 , P2_SUB_594_U89 );
and AND2_13698 ( P2_SUB_594_U25 , P2_SUB_594_U98 , P2_SUB_594_U30 );
and AND2_13699 ( P2_SUB_594_U26 , P2_SUB_594_U97 , P2_SUB_594_U31 );
and AND2_13700 ( P2_SUB_594_U27 , P2_SUB_594_U95 , P2_SUB_594_U92 );
and AND2_13701 ( P2_SUB_594_U28 , P2_SUB_594_U94 , P2_SUB_594_U29 );
nand NAND2_13702 ( P2_SUB_594_U29 , P2_SUB_594_U56 , P2_SUB_594_U55 );
or OR5_13703 ( P2_SUB_594_U30 , P2_IR_REG_1_ , P2_IR_REG_0_ , P2_IR_REG_2_ , P2_IR_REG_3_ , P2_IR_REG_4_ );
nand NAND2_13704 ( P2_SUB_594_U31 , P2_SUB_594_U57 , P2_SUB_594_U90 );
not NOT1_13705 ( P2_SUB_594_U32 , P2_IR_REG_7_ );
or OR3_13706 ( P2_SUB_594_U33 , P2_IR_REG_1_ , P2_IR_REG_0_ , P2_IR_REG_2_ );
not NOT1_13707 ( P2_SUB_594_U34 , P2_IR_REG_3_ );
nand NAND2_13708 ( P2_SUB_594_U35 , P2_SUB_594_U59 , P2_SUB_594_U93 );
nand NAND2_13709 ( P2_SUB_594_U36 , P2_SUB_594_U61 , P2_SUB_594_U105 );
nand NAND2_13710 ( P2_SUB_594_U37 , P2_SUB_594_U62 , P2_SUB_594_U111 );
nand NAND2_13711 ( P2_SUB_594_U38 , P2_SUB_594_U113 , P2_SUB_594_U39 );
not NOT1_13712 ( P2_SUB_594_U39 , P2_IR_REG_29_ );
not NOT1_13713 ( P2_SUB_594_U40 , P2_IR_REG_27_ );
nand NAND2_13714 ( P2_SUB_594_U41 , P2_SUB_594_U105 , P2_SUB_594_U7 );
nand NAND2_13715 ( P2_SUB_594_U42 , P2_SUB_594_U65 , P2_SUB_594_U108 );
not NOT1_13716 ( P2_SUB_594_U43 , P2_IR_REG_24_ );
not NOT1_13717 ( P2_SUB_594_U44 , P2_IR_REG_23_ );
nand NAND2_13718 ( P2_SUB_594_U45 , P2_SUB_594_U66 , P2_SUB_594_U105 );
not NOT1_13719 ( P2_SUB_594_U46 , P2_IR_REG_19_ );
nand NAND2_13720 ( P2_SUB_594_U47 , P2_SUB_594_U6 , P2_SUB_594_U93 );
nand NAND2_13721 ( P2_SUB_594_U48 , P2_SUB_594_U67 , P2_SUB_594_U102 );
not NOT1_13722 ( P2_SUB_594_U49 , P2_IR_REG_16_ );
not NOT1_13723 ( P2_SUB_594_U50 , P2_IR_REG_15_ );
nand NAND2_13724 ( P2_SUB_594_U51 , P2_SUB_594_U68 , P2_SUB_594_U93 );
not NOT1_13725 ( P2_SUB_594_U52 , P2_IR_REG_11_ );
nand NAND2_13726 ( P2_SUB_594_U53 , P2_SUB_594_U154 , P2_SUB_594_U153 );
nand NAND2_13727 ( P2_SUB_594_U54 , P2_SUB_594_U144 , P2_SUB_594_U143 );
nor nor_13728 ( P2_SUB_594_U55 , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_2_ , P2_IR_REG_1_ , P2_IR_REG_0_ );
nor nor_13729 ( P2_SUB_594_U56 , P2_IR_REG_5_ , P2_IR_REG_6_ , P2_IR_REG_7_ , P2_IR_REG_8_ );
nor nor_13730 ( P2_SUB_594_U57 , P2_IR_REG_5_ , P2_IR_REG_6_ );
nor nor_13731 ( P2_SUB_594_U58 , P2_IR_REG_15_ , P2_IR_REG_13_ , P2_IR_REG_14_ );
and AND3_13732 ( P2_SUB_594_U59 , P2_SUB_594_U6 , P2_SUB_594_U49 , P2_SUB_594_U58 );
nor nor_13733 ( P2_SUB_594_U60 , P2_IR_REG_23_ , P2_IR_REG_21_ , P2_IR_REG_22_ );
and AND3_13734 ( P2_SUB_594_U61 , P2_SUB_594_U7 , P2_SUB_594_U43 , P2_SUB_594_U60 );
nor nor_13735 ( P2_SUB_594_U62 , P2_IR_REG_25_ , P2_IR_REG_26_ , P2_IR_REG_27_ , P2_IR_REG_28_ );
nor nor_13736 ( P2_SUB_594_U63 , P2_IR_REG_25_ , P2_IR_REG_26_ );
and AND2_13737 ( P2_SUB_594_U64 , P2_SUB_594_U137 , P2_SUB_594_U37 );
nor nor_13738 ( P2_SUB_594_U65 , P2_IR_REG_21_ , P2_IR_REG_22_ );
nor nor_13739 ( P2_SUB_594_U66 , P2_IR_REG_17_ , P2_IR_REG_18_ );
nor nor_13740 ( P2_SUB_594_U67 , P2_IR_REG_13_ , P2_IR_REG_14_ );
nor nor_13741 ( P2_SUB_594_U68 , P2_IR_REG_10_ , P2_IR_REG_9_ );
not NOT1_13742 ( P2_SUB_594_U69 , P2_IR_REG_9_ );
and AND2_13743 ( P2_SUB_594_U70 , P2_SUB_594_U140 , P2_SUB_594_U139 );
not NOT1_13744 ( P2_SUB_594_U71 , P2_IR_REG_5_ );
and AND2_13745 ( P2_SUB_594_U72 , P2_SUB_594_U142 , P2_SUB_594_U141 );
not NOT1_13746 ( P2_SUB_594_U73 , P2_IR_REG_31_ );
not NOT1_13747 ( P2_SUB_594_U74 , P2_IR_REG_30_ );
and AND2_13748 ( P2_SUB_594_U75 , P2_SUB_594_U146 , P2_SUB_594_U145 );
nand NAND2_13749 ( P2_SUB_594_U76 , P2_SUB_594_U63 , P2_SUB_594_U111 );
and AND2_13750 ( P2_SUB_594_U77 , P2_SUB_594_U148 , P2_SUB_594_U147 );
not NOT1_13751 ( P2_SUB_594_U78 , P2_IR_REG_25_ );
and AND2_13752 ( P2_SUB_594_U79 , P2_SUB_594_U150 , P2_SUB_594_U149 );
not NOT1_13753 ( P2_SUB_594_U80 , P2_IR_REG_21_ );
and AND2_13754 ( P2_SUB_594_U81 , P2_SUB_594_U152 , P2_SUB_594_U151 );
not NOT1_13755 ( P2_SUB_594_U82 , P2_IR_REG_1_ );
not NOT1_13756 ( P2_SUB_594_U83 , P2_IR_REG_0_ );
not NOT1_13757 ( P2_SUB_594_U84 , P2_IR_REG_17_ );
and AND2_13758 ( P2_SUB_594_U85 , P2_SUB_594_U156 , P2_SUB_594_U155 );
not NOT1_13759 ( P2_SUB_594_U86 , P2_IR_REG_13_ );
and AND2_13760 ( P2_SUB_594_U87 , P2_SUB_594_U158 , P2_SUB_594_U157 );
not NOT1_13761 ( P2_SUB_594_U88 , P2_SUB_594_U33 );
nand NAND2_13762 ( P2_SUB_594_U89 , P2_SUB_594_U88 , P2_SUB_594_U34 );
not NOT1_13763 ( P2_SUB_594_U90 , P2_SUB_594_U30 );
not NOT1_13764 ( P2_SUB_594_U91 , P2_SUB_594_U31 );
nand NAND2_13765 ( P2_SUB_594_U92 , P2_SUB_594_U91 , P2_SUB_594_U32 );
not NOT1_13766 ( P2_SUB_594_U93 , P2_SUB_594_U29 );
nand NAND2_13767 ( P2_SUB_594_U94 , P2_IR_REG_8_ , P2_SUB_594_U92 );
nand NAND2_13768 ( P2_SUB_594_U95 , P2_IR_REG_7_ , P2_SUB_594_U31 );
nand NAND2_13769 ( P2_SUB_594_U96 , P2_SUB_594_U90 , P2_SUB_594_U71 );
nand NAND2_13770 ( P2_SUB_594_U97 , P2_IR_REG_6_ , P2_SUB_594_U96 );
nand NAND2_13771 ( P2_SUB_594_U98 , P2_IR_REG_4_ , P2_SUB_594_U89 );
nand NAND2_13772 ( P2_SUB_594_U99 , P2_IR_REG_3_ , P2_SUB_594_U33 );
not NOT1_13773 ( P2_SUB_594_U100 , P2_SUB_594_U51 );
nand NAND2_13774 ( P2_SUB_594_U101 , P2_SUB_594_U100 , P2_SUB_594_U52 );
not NOT1_13775 ( P2_SUB_594_U102 , P2_SUB_594_U47 );
not NOT1_13776 ( P2_SUB_594_U103 , P2_SUB_594_U48 );
nand NAND2_13777 ( P2_SUB_594_U104 , P2_SUB_594_U103 , P2_SUB_594_U50 );
not NOT1_13778 ( P2_SUB_594_U105 , P2_SUB_594_U35 );
not NOT1_13779 ( P2_SUB_594_U106 , P2_SUB_594_U45 );
nand NAND2_13780 ( P2_SUB_594_U107 , P2_SUB_594_U106 , P2_SUB_594_U46 );
not NOT1_13781 ( P2_SUB_594_U108 , P2_SUB_594_U41 );
not NOT1_13782 ( P2_SUB_594_U109 , P2_SUB_594_U42 );
nand NAND2_13783 ( P2_SUB_594_U110 , P2_SUB_594_U109 , P2_SUB_594_U44 );
not NOT1_13784 ( P2_SUB_594_U111 , P2_SUB_594_U36 );
not NOT1_13785 ( P2_SUB_594_U112 , P2_SUB_594_U76 );
not NOT1_13786 ( P2_SUB_594_U113 , P2_SUB_594_U37 );
not NOT1_13787 ( P2_SUB_594_U114 , P2_SUB_594_U38 );
or OR2_13788 ( P2_SUB_594_U115 , P2_IR_REG_1_ , P2_IR_REG_0_ );
nand NAND2_13789 ( P2_SUB_594_U116 , P2_IR_REG_2_ , P2_SUB_594_U115 );
nand NAND2_13790 ( P2_SUB_594_U117 , P2_IR_REG_29_ , P2_SUB_594_U37 );
nand NAND2_13791 ( P2_SUB_594_U118 , P2_SUB_594_U111 , P2_SUB_594_U78 );
nand NAND2_13792 ( P2_SUB_594_U119 , P2_IR_REG_26_ , P2_SUB_594_U118 );
nand NAND2_13793 ( P2_SUB_594_U120 , P2_IR_REG_24_ , P2_SUB_594_U110 );
nand NAND2_13794 ( P2_SUB_594_U121 , P2_IR_REG_23_ , P2_SUB_594_U42 );
nand NAND2_13795 ( P2_SUB_594_U122 , P2_SUB_594_U108 , P2_SUB_594_U80 );
nand NAND2_13796 ( P2_SUB_594_U123 , P2_IR_REG_22_ , P2_SUB_594_U122 );
nand NAND2_13797 ( P2_SUB_594_U124 , P2_IR_REG_20_ , P2_SUB_594_U107 );
nand NAND2_13798 ( P2_SUB_594_U125 , P2_IR_REG_19_ , P2_SUB_594_U45 );
nand NAND2_13799 ( P2_SUB_594_U126 , P2_SUB_594_U105 , P2_SUB_594_U84 );
nand NAND2_13800 ( P2_SUB_594_U127 , P2_IR_REG_18_ , P2_SUB_594_U126 );
nand NAND2_13801 ( P2_SUB_594_U128 , P2_IR_REG_16_ , P2_SUB_594_U104 );
nand NAND2_13802 ( P2_SUB_594_U129 , P2_IR_REG_15_ , P2_SUB_594_U48 );
nand NAND2_13803 ( P2_SUB_594_U130 , P2_SUB_594_U102 , P2_SUB_594_U86 );
nand NAND2_13804 ( P2_SUB_594_U131 , P2_IR_REG_14_ , P2_SUB_594_U130 );
nand NAND2_13805 ( P2_SUB_594_U132 , P2_IR_REG_12_ , P2_SUB_594_U101 );
nand NAND2_13806 ( P2_SUB_594_U133 , P2_IR_REG_11_ , P2_SUB_594_U51 );
nand NAND2_13807 ( P2_SUB_594_U134 , P2_SUB_594_U93 , P2_SUB_594_U69 );
nand NAND2_13808 ( P2_SUB_594_U135 , P2_IR_REG_10_ , P2_SUB_594_U134 );
nand NAND2_13809 ( P2_SUB_594_U136 , P2_SUB_594_U114 , P2_SUB_594_U74 );
nand NAND2_13810 ( P2_SUB_594_U137 , P2_IR_REG_27_ , P2_IR_REG_28_ );
nand NAND2_13811 ( P2_SUB_594_U138 , P2_IR_REG_28_ , P2_SUB_594_U76 );
nand NAND2_13812 ( P2_SUB_594_U139 , P2_IR_REG_9_ , P2_SUB_594_U29 );
nand NAND2_13813 ( P2_SUB_594_U140 , P2_SUB_594_U93 , P2_SUB_594_U69 );
nand NAND2_13814 ( P2_SUB_594_U141 , P2_IR_REG_5_ , P2_SUB_594_U30 );
nand NAND2_13815 ( P2_SUB_594_U142 , P2_SUB_594_U90 , P2_SUB_594_U71 );
nand NAND2_13816 ( P2_SUB_594_U143 , P2_SUB_594_U136 , P2_SUB_594_U73 );
nand NAND3_13817 ( P2_SUB_594_U144 , P2_SUB_594_U114 , P2_SUB_594_U74 , P2_IR_REG_31_ );
nand NAND2_13818 ( P2_SUB_594_U145 , P2_IR_REG_30_ , P2_SUB_594_U38 );
nand NAND2_13819 ( P2_SUB_594_U146 , P2_SUB_594_U114 , P2_SUB_594_U74 );
nand NAND2_13820 ( P2_SUB_594_U147 , P2_IR_REG_27_ , P2_SUB_594_U76 );
nand NAND2_13821 ( P2_SUB_594_U148 , P2_SUB_594_U112 , P2_SUB_594_U40 );
nand NAND2_13822 ( P2_SUB_594_U149 , P2_IR_REG_25_ , P2_SUB_594_U36 );
nand NAND2_13823 ( P2_SUB_594_U150 , P2_SUB_594_U111 , P2_SUB_594_U78 );
nand NAND2_13824 ( P2_SUB_594_U151 , P2_IR_REG_21_ , P2_SUB_594_U41 );
nand NAND2_13825 ( P2_SUB_594_U152 , P2_SUB_594_U108 , P2_SUB_594_U80 );
nand NAND2_13826 ( P2_SUB_594_U153 , P2_IR_REG_1_ , P2_SUB_594_U83 );
nand NAND2_13827 ( P2_SUB_594_U154 , P2_IR_REG_0_ , P2_SUB_594_U82 );
nand NAND2_13828 ( P2_SUB_594_U155 , P2_IR_REG_17_ , P2_SUB_594_U35 );
nand NAND2_13829 ( P2_SUB_594_U156 , P2_SUB_594_U105 , P2_SUB_594_U84 );
nand NAND2_13830 ( P2_SUB_594_U157 , P2_IR_REG_13_ , P2_SUB_594_U47 );
nand NAND2_13831 ( P2_SUB_594_U158 , P2_SUB_594_U102 , P2_SUB_594_U86 );
and AND3_13832 ( P2_R693_U6 , P2_R693_U110 , P2_R693_U111 , P2_R693_U109 );
and AND2_13833 ( P2_R693_U7 , P2_R693_U118 , P2_R693_U119 );
and AND2_13834 ( P2_R693_U8 , P2_R693_U120 , P2_R693_U121 );
and AND4_13835 ( P2_R693_U9 , P2_R693_U81 , P2_R693_U123 , P2_R693_U125 , P2_R693_U8 );
and AND4_13836 ( P2_R693_U10 , P2_R693_U134 , P2_R693_U133 , P2_R693_U132 , P2_R693_U130 );
and AND2_13837 ( P2_R693_U11 , P2_R693_U83 , P2_R693_U10 );
and AND2_13838 ( P2_R693_U12 , P2_R693_U11 , P2_R693_U138 );
and AND2_13839 ( P2_R693_U13 , P2_R693_U144 , P2_R693_U143 );
and AND3_13840 ( P2_R693_U14 , P2_R693_U105 , P2_R693_U189 , P2_R693_U104 );
not NOT1_13841 ( P2_R693_U15 , P2_U3529 );
not NOT1_13842 ( P2_R693_U16 , P2_U3904 );
not NOT1_13843 ( P2_R693_U17 , P2_U3896 );
not NOT1_13844 ( P2_R693_U18 , P2_U3895 );
not NOT1_13845 ( P2_R693_U19 , P2_U3535 );
not NOT1_13846 ( P2_R693_U20 , P2_U3532 );
not NOT1_13847 ( P2_R693_U21 , P2_U3534 );
not NOT1_13848 ( P2_R693_U22 , P2_U3537 );
not NOT1_13849 ( P2_R693_U23 , P2_U3536 );
not NOT1_13850 ( P2_R693_U24 , P2_U3901 );
not NOT1_13851 ( P2_R693_U25 , P2_U3540 );
not NOT1_13852 ( P2_R693_U26 , P2_U3902 );
not NOT1_13853 ( P2_R693_U27 , P2_U3541 );
not NOT1_13854 ( P2_R693_U28 , P2_U3543 );
not NOT1_13855 ( P2_R693_U29 , P2_U3443 );
not NOT1_13856 ( P2_R693_U30 , P2_U3544 );
not NOT1_13857 ( P2_R693_U31 , P2_U3440 );
not NOT1_13858 ( P2_R693_U32 , P2_U3445 );
not NOT1_13859 ( P2_R693_U33 , P2_U3903 );
not NOT1_13860 ( P2_R693_U34 , P2_U3545 );
not NOT1_13861 ( P2_R693_U35 , P2_U3546 );
not NOT1_13862 ( P2_R693_U36 , P2_U3437 );
not NOT1_13863 ( P2_R693_U37 , P2_U3434 );
not NOT1_13864 ( P2_R693_U38 , P2_U3419 );
not NOT1_13865 ( P2_R693_U39 , P2_U3416 );
not NOT1_13866 ( P2_R693_U40 , P2_U3410 );
not NOT1_13867 ( P2_R693_U41 , P2_U3413 );
not NOT1_13868 ( P2_R693_U42 , P2_U3407 );
not NOT1_13869 ( P2_R693_U43 , P2_U3404 );
not NOT1_13870 ( P2_R693_U44 , P2_U3401 );
not NOT1_13871 ( P2_R693_U45 , P2_U3398 );
not NOT1_13872 ( P2_R693_U46 , P2_U3553 );
not NOT1_13873 ( P2_R693_U47 , P2_U3395 );
not NOT1_13874 ( P2_R693_U48 , P2_U3392 );
not NOT1_13875 ( P2_R693_U49 , P2_U3550 );
not NOT1_13876 ( P2_R693_U50 , P2_U3549 );
not NOT1_13877 ( P2_R693_U51 , P2_U3542 );
not NOT1_13878 ( P2_R693_U52 , P2_U3531 );
not NOT1_13879 ( P2_R693_U53 , P2_U3528 );
not NOT1_13880 ( P2_R693_U54 , P2_U3527 );
not NOT1_13881 ( P2_R693_U55 , P2_U3526 );
not NOT1_13882 ( P2_R693_U56 , P2_U3525 );
not NOT1_13883 ( P2_R693_U57 , P2_U3524 );
not NOT1_13884 ( P2_R693_U58 , P2_U3523 );
not NOT1_13885 ( P2_R693_U59 , P2_U3552 );
not NOT1_13886 ( P2_R693_U60 , P2_U3551 );
not NOT1_13887 ( P2_R693_U61 , P2_U3425 );
not NOT1_13888 ( P2_R693_U62 , P2_U3422 );
not NOT1_13889 ( P2_R693_U63 , P2_U3431 );
not NOT1_13890 ( P2_R693_U64 , P2_U3428 );
not NOT1_13891 ( P2_R693_U65 , P2_U3548 );
not NOT1_13892 ( P2_R693_U66 , P2_U3547 );
not NOT1_13893 ( P2_R693_U67 , P2_U3539 );
not NOT1_13894 ( P2_R693_U68 , P2_U3538 );
not NOT1_13895 ( P2_R693_U69 , P2_U3900 );
not NOT1_13896 ( P2_R693_U70 , P2_U3899 );
not NOT1_13897 ( P2_R693_U71 , P2_U3898 );
not NOT1_13898 ( P2_R693_U72 , P2_U3897 );
not NOT1_13899 ( P2_R693_U73 , P2_U3868 );
not NOT1_13900 ( P2_R693_U74 , P2_U3533 );
and AND2_13901 ( P2_R693_U75 , P2_U3532 , P2_R693_U16 );
and AND2_13902 ( P2_R693_U76 , P2_U3540 , P2_R693_U26 );
and AND2_13903 ( P2_R693_U77 , P2_U3541 , P2_R693_U33 );
and AND2_13904 ( P2_R693_U78 , P2_R693_U174 , P2_R693_U173 );
and AND2_13905 ( P2_R693_U79 , P2_U3443 , P2_R693_U30 );
and AND2_13906 ( P2_R693_U80 , P2_U3440 , P2_R693_U34 );
and AND2_13907 ( P2_R693_U81 , P2_R693_U124 , P2_R693_U122 );
and AND2_13908 ( P2_R693_U82 , P2_U3387 , P2_R693_U107 );
and AND3_13909 ( P2_R693_U83 , P2_R693_U136 , P2_R693_U135 , P2_R693_U137 );
and AND2_13910 ( P2_R693_U84 , P2_R693_U140 , P2_R693_U141 );
and AND2_13911 ( P2_R693_U85 , P2_R693_U84 , P2_R693_U139 );
and AND2_13912 ( P2_R693_U86 , P2_U3542 , P2_R693_U47 );
and AND2_13913 ( P2_R693_U87 , P2_U3531 , P2_R693_U45 );
and AND2_13914 ( P2_R693_U88 , P2_R693_U136 , P2_R693_U135 );
and AND2_13915 ( P2_R693_U89 , P2_R693_U152 , P2_R693_U153 );
and AND2_13916 ( P2_R693_U90 , P2_R693_U132 , P2_R693_U130 );
and AND2_13917 ( P2_R693_U91 , P2_R693_U13 , P2_R693_U160 );
and AND3_13918 ( P2_R693_U92 , P2_R693_U159 , P2_R693_U158 , P2_R693_U91 );
and AND2_13919 ( P2_R693_U93 , P2_U3425 , P2_R693_U49 );
and AND2_13920 ( P2_R693_U94 , P2_U3422 , P2_R693_U60 );
and AND2_13921 ( P2_R693_U95 , P2_R693_U163 , P2_R693_U97 );
and AND2_13922 ( P2_R693_U96 , P2_R693_U95 , P2_R693_U164 );
and AND2_13923 ( P2_R693_U97 , P2_R693_U166 , P2_R693_U165 );
and AND4_13924 ( P2_R693_U98 , P2_R693_U177 , P2_R693_U176 , P2_R693_U127 , P2_R693_U128 );
and AND2_13925 ( P2_R693_U99 , P2_R693_U181 , P2_R693_U180 );
and AND2_13926 ( P2_R693_U100 , P2_R693_U188 , P2_R693_U187 );
and AND2_13927 ( P2_R693_U101 , P2_R693_U100 , P2_R693_U6 );
and AND2_13928 ( P2_R693_U102 , P2_R693_U103 , P2_R693_U191 );
and AND2_13929 ( P2_R693_U103 , P2_U3533 , P2_R693_U18 );
and AND4_13930 ( P2_R693_U104 , P2_R693_U117 , P2_R693_U116 , P2_R693_U115 , P2_R693_U114 );
and AND2_13931 ( P2_R693_U105 , P2_R693_U190 , P2_R693_U192 );
not NOT1_13932 ( P2_R693_U106 , P2_U3869 );
not NOT1_13933 ( P2_R693_U107 , P2_U3554 );
nand NAND2_13934 ( P2_R693_U108 , P2_R693_U113 , P2_R693_U193 );
nand NAND2_13935 ( P2_R693_U109 , P2_U3904 , P2_R693_U20 );
nand NAND2_13936 ( P2_R693_U110 , P2_U3896 , P2_R693_U21 );
nand NAND2_13937 ( P2_R693_U111 , P2_U3895 , P2_R693_U74 );
nand NAND2_13938 ( P2_R693_U112 , P2_U3529 , P2_R693_U73 );
nand NAND2_13939 ( P2_R693_U113 , P2_R693_U112 , P2_R693_U106 );
nand NAND4_13940 ( P2_R693_U114 , P2_U3535 , P2_R693_U6 , P2_R693_U108 , P2_R693_U72 );
nand NAND3_13941 ( P2_R693_U115 , P2_R693_U112 , P2_U3530 , P2_R693_U106 );
nand NAND2_13942 ( P2_R693_U116 , P2_R693_U75 , P2_R693_U108 );
nand NAND4_13943 ( P2_R693_U117 , P2_U3534 , P2_R693_U6 , P2_R693_U108 , P2_R693_U17 );
nand NAND2_13944 ( P2_R693_U118 , P2_U3543 , P2_R693_U32 );
nand NAND2_13945 ( P2_R693_U119 , P2_U3544 , P2_R693_U29 );
nand NAND2_13946 ( P2_R693_U120 , P2_U3901 , P2_R693_U67 );
nand NAND2_13947 ( P2_R693_U121 , P2_U3902 , P2_R693_U25 );
nand NAND2_13948 ( P2_R693_U122 , P2_R693_U79 , P2_R693_U118 );
nand NAND2_13949 ( P2_R693_U123 , P2_R693_U80 , P2_R693_U7 );
nand NAND2_13950 ( P2_R693_U124 , P2_U3445 , P2_R693_U28 );
nand NAND2_13951 ( P2_R693_U125 , P2_U3903 , P2_R693_U27 );
nand NAND2_13952 ( P2_R693_U126 , P2_U3437 , P2_R693_U35 );
nand NAND2_13953 ( P2_R693_U127 , P2_U3537 , P2_R693_U70 );
nand NAND2_13954 ( P2_R693_U128 , P2_U3536 , P2_R693_U71 );
nand NAND2_13955 ( P2_R693_U129 , P2_U3434 , P2_R693_U66 );
nand NAND2_13956 ( P2_R693_U130 , P2_U3419 , P2_R693_U59 );
nand NAND2_13957 ( P2_R693_U131 , P2_U3553 , P2_R693_U48 );
nand NAND2_13958 ( P2_R693_U132 , P2_U3416 , P2_R693_U58 );
nand NAND2_13959 ( P2_R693_U133 , P2_U3410 , P2_R693_U56 );
nand NAND2_13960 ( P2_R693_U134 , P2_U3413 , P2_R693_U57 );
nand NAND2_13961 ( P2_R693_U135 , P2_U3407 , P2_R693_U55 );
nand NAND2_13962 ( P2_R693_U136 , P2_U3404 , P2_R693_U54 );
nand NAND2_13963 ( P2_R693_U137 , P2_U3401 , P2_R693_U53 );
nand NAND2_13964 ( P2_R693_U138 , P2_U3398 , P2_R693_U52 );
nand NAND2_13965 ( P2_R693_U139 , P2_R693_U82 , P2_R693_U131 );
nand NAND2_13966 ( P2_R693_U140 , P2_U3395 , P2_R693_U51 );
nand NAND2_13967 ( P2_R693_U141 , P2_U3392 , P2_R693_U46 );
nand NAND2_13968 ( P2_R693_U142 , P2_R693_U85 , P2_R693_U12 );
nand NAND2_13969 ( P2_R693_U143 , P2_U3550 , P2_R693_U61 );
nand NAND2_13970 ( P2_R693_U144 , P2_U3549 , P2_R693_U64 );
nand NAND2_13971 ( P2_R693_U145 , P2_U3524 , P2_R693_U41 );
nand NAND2_13972 ( P2_R693_U146 , P2_U3523 , P2_R693_U39 );
nand NAND2_13973 ( P2_R693_U147 , P2_R693_U146 , P2_R693_U145 );
nand NAND2_13974 ( P2_R693_U148 , P2_U3528 , P2_R693_U44 );
nand NAND2_13975 ( P2_R693_U149 , P2_U3527 , P2_R693_U43 );
nand NAND2_13976 ( P2_R693_U150 , P2_R693_U149 , P2_R693_U148 );
nand NAND2_13977 ( P2_R693_U151 , P2_R693_U88 , P2_R693_U150 );
nand NAND2_13978 ( P2_R693_U152 , P2_U3526 , P2_R693_U42 );
nand NAND2_13979 ( P2_R693_U153 , P2_U3525 , P2_R693_U40 );
nand NAND2_13980 ( P2_R693_U154 , P2_R693_U89 , P2_R693_U151 );
nand NAND2_13981 ( P2_R693_U155 , P2_R693_U86 , P2_R693_U12 );
nand NAND2_13982 ( P2_R693_U156 , P2_R693_U87 , P2_R693_U11 );
nand NAND2_13983 ( P2_R693_U157 , P2_R693_U10 , P2_R693_U154 );
nand NAND2_13984 ( P2_R693_U158 , P2_R693_U90 , P2_R693_U147 );
nand NAND2_13985 ( P2_R693_U159 , P2_U3552 , P2_R693_U38 );
nand NAND2_13986 ( P2_R693_U160 , P2_U3551 , P2_R693_U62 );
nand NAND5_13987 ( P2_R693_U161 , P2_R693_U157 , P2_R693_U156 , P2_R693_U92 , P2_R693_U155 , P2_R693_U142 );
nand NAND2_13988 ( P2_R693_U162 , P2_U3549 , P2_R693_U64 );
nand NAND2_13989 ( P2_R693_U163 , P2_R693_U93 , P2_R693_U162 );
nand NAND2_13990 ( P2_R693_U164 , P2_R693_U94 , P2_R693_U13 );
nand NAND2_13991 ( P2_R693_U165 , P2_U3431 , P2_R693_U65 );
nand NAND2_13992 ( P2_R693_U166 , P2_U3428 , P2_R693_U50 );
nand NAND2_13993 ( P2_R693_U167 , P2_R693_U161 , P2_R693_U96 );
nand NAND2_13994 ( P2_R693_U168 , P2_U3548 , P2_R693_U63 );
nand NAND2_13995 ( P2_R693_U169 , P2_R693_U168 , P2_R693_U167 );
nand NAND2_13996 ( P2_R693_U170 , P2_R693_U169 , P2_R693_U129 );
nand NAND2_13997 ( P2_R693_U171 , P2_U3547 , P2_R693_U37 );
nand NAND2_13998 ( P2_R693_U172 , P2_R693_U171 , P2_R693_U170 );
nand NAND2_13999 ( P2_R693_U173 , P2_U3545 , P2_R693_U31 );
nand NAND2_14000 ( P2_R693_U174 , P2_U3546 , P2_R693_U36 );
nand NAND2_14001 ( P2_R693_U175 , P2_R693_U78 , P2_R693_U7 );
nand NAND2_14002 ( P2_R693_U176 , P2_R693_U76 , P2_R693_U120 );
nand NAND2_14003 ( P2_R693_U177 , P2_R693_U77 , P2_R693_U8 );
nand NAND2_14004 ( P2_R693_U178 , P2_R693_U9 , P2_R693_U175 );
nand NAND3_14005 ( P2_R693_U179 , P2_R693_U172 , P2_R693_U126 , P2_R693_U9 );
nand NAND2_14006 ( P2_R693_U180 , P2_U3539 , P2_R693_U24 );
nand NAND2_14007 ( P2_R693_U181 , P2_U3538 , P2_R693_U69 );
nand NAND4_14008 ( P2_R693_U182 , P2_R693_U179 , P2_R693_U178 , P2_R693_U99 , P2_R693_U98 );
nand NAND2_14009 ( P2_R693_U183 , P2_U3900 , P2_R693_U68 );
nand NAND2_14010 ( P2_R693_U184 , P2_U3899 , P2_R693_U22 );
nand NAND2_14011 ( P2_R693_U185 , P2_R693_U184 , P2_R693_U183 );
nand NAND3_14012 ( P2_R693_U186 , P2_R693_U185 , P2_R693_U127 , P2_R693_U128 );
nand NAND2_14013 ( P2_R693_U187 , P2_U3898 , P2_R693_U23 );
nand NAND2_14014 ( P2_R693_U188 , P2_U3897 , P2_R693_U19 );
nand NAND4_14015 ( P2_R693_U189 , P2_R693_U182 , P2_R693_U186 , P2_R693_U108 , P2_R693_U101 );
nand NAND2_14016 ( P2_R693_U190 , P2_U3868 , P2_R693_U15 );
nand NAND2_14017 ( P2_R693_U191 , P2_U3904 , P2_R693_U20 );
nand NAND2_14018 ( P2_R693_U192 , P2_R693_U108 , P2_R693_U102 );
nand NAND2_14019 ( P2_R693_U193 , P2_U3530 , P2_R693_U112 );
nand NAND2_14020 ( P2_SUB_605_U6 , P2_SUB_605_U39 , P2_SUB_605_U100 );
nand NAND2_14021 ( P2_SUB_605_U7 , P2_SUB_605_U81 , P2_SUB_605_U107 );
nand NAND2_14022 ( P2_SUB_605_U8 , P2_SUB_605_U65 , P2_SUB_605_U72 );
nand NAND2_14023 ( P2_SUB_605_U9 , P2_SUB_605_U34 , P2_SUB_605_U112 );
nand NAND2_14024 ( P2_SUB_605_U10 , P2_SUB_605_U89 , P2_SUB_605_U99 );
nand NAND2_14025 ( P2_SUB_605_U11 , P2_SUB_605_U83 , P2_SUB_605_U105 );
nand NAND2_14026 ( P2_SUB_605_U12 , P2_SUB_605_U67 , P2_SUB_605_U70 );
nand NAND2_14027 ( P2_SUB_605_U13 , P2_SUB_605_U75 , P2_SUB_605_U113 );
nand NAND2_14028 ( P2_SUB_605_U14 , P2_SUB_605_U68 , P2_SUB_605_U69 );
nand NAND2_14029 ( P2_SUB_605_U15 , P2_SUB_605_U37 , P2_SUB_605_U104 );
nand NAND2_14030 ( P2_SUB_605_U16 , P2_SUB_605_U40 , P2_SUB_605_U98 );
nand NAND2_14031 ( P2_SUB_605_U17 , P2_SUB_605_U87 , P2_SUB_605_U101 );
nand NAND2_14032 ( P2_SUB_605_U18 , P2_SUB_605_U32 , P2_SUB_605_U71 );
nand NAND2_14033 ( P2_SUB_605_U19 , P2_SUB_605_U36 , P2_SUB_605_U106 );
nand NAND2_14034 ( P2_SUB_605_U20 , P2_SUB_605_U85 , P2_SUB_605_U103 );
nand NAND2_14035 ( P2_SUB_605_U21 , P2_SUB_605_U35 , P2_SUB_605_U108 );
nand NAND2_14036 ( P2_SUB_605_U22 , P2_SUB_605_U64 , P2_SUB_605_U73 );
nand NAND2_14037 ( P2_SUB_605_U23 , P2_SUB_605_U41 , P2_SUB_605_U96 );
nand NAND2_14038 ( P2_SUB_605_U24 , P2_SUB_605_U77 , P2_SUB_605_U111 );
nand NAND2_14039 ( P2_SUB_605_U25 , P2_SUB_605_U49 , P2_SUB_605_U110 );
not NOT1_14040 ( P2_SUB_605_U26 , P2_REG3_REG_3_ );
nand NAND2_14041 ( P2_SUB_605_U27 , P2_SUB_605_U91 , P2_SUB_605_U97 );
nand NAND2_14042 ( P2_SUB_605_U28 , P2_SUB_605_U38 , P2_SUB_605_U102 );
nand NAND2_14043 ( P2_SUB_605_U29 , P2_SUB_605_U93 , P2_SUB_605_U95 );
nand NAND2_14044 ( P2_SUB_605_U30 , P2_SUB_605_U63 , P2_SUB_605_U74 );
nand NAND2_14045 ( P2_SUB_605_U31 , P2_SUB_605_U79 , P2_SUB_605_U109 );
or OR5_14046 ( P2_SUB_605_U32 , P2_REG3_REG_4_ , P2_REG3_REG_3_ , P2_REG3_REG_5_ , P2_REG3_REG_6_ , P2_REG3_REG_7_ );
not NOT1_14047 ( P2_SUB_605_U33 , P2_REG3_REG_8_ );
nand NAND2_14048 ( P2_SUB_605_U34 , P2_SUB_605_U53 , P2_SUB_605_U66 );
nand NAND2_14049 ( P2_SUB_605_U35 , P2_SUB_605_U54 , P2_SUB_605_U76 );
nand NAND2_14050 ( P2_SUB_605_U36 , P2_SUB_605_U55 , P2_SUB_605_U80 );
nand NAND2_14051 ( P2_SUB_605_U37 , P2_SUB_605_U56 , P2_SUB_605_U82 );
nand NAND2_14052 ( P2_SUB_605_U38 , P2_SUB_605_U57 , P2_SUB_605_U84 );
nand NAND2_14053 ( P2_SUB_605_U39 , P2_SUB_605_U58 , P2_SUB_605_U86 );
nand NAND2_14054 ( P2_SUB_605_U40 , P2_SUB_605_U59 , P2_SUB_605_U88 );
nand NAND2_14055 ( P2_SUB_605_U41 , P2_SUB_605_U60 , P2_SUB_605_U90 );
not NOT1_14056 ( P2_SUB_605_U42 , P2_REG3_REG_28_ );
not NOT1_14057 ( P2_SUB_605_U43 , P2_REG3_REG_26_ );
not NOT1_14058 ( P2_SUB_605_U44 , P2_REG3_REG_24_ );
not NOT1_14059 ( P2_SUB_605_U45 , P2_REG3_REG_22_ );
not NOT1_14060 ( P2_SUB_605_U46 , P2_REG3_REG_20_ );
not NOT1_14061 ( P2_SUB_605_U47 , P2_REG3_REG_18_ );
not NOT1_14062 ( P2_SUB_605_U48 , P2_REG3_REG_16_ );
nand NAND2_14063 ( P2_SUB_605_U49 , P2_SUB_605_U61 , P2_SUB_605_U76 );
not NOT1_14064 ( P2_SUB_605_U50 , P2_REG3_REG_14_ );
not NOT1_14065 ( P2_SUB_605_U51 , P2_REG3_REG_12_ );
nor nor_14066 ( P2_SUB_605_U52 , P2_REG3_REG_8_ , P2_REG3_REG_9_ );
nor nor_14067 ( P2_SUB_605_U53 , P2_REG3_REG_10_ , P2_REG3_REG_11_ , P2_REG3_REG_8_ , P2_REG3_REG_9_ );
nor nor_14068 ( P2_SUB_605_U54 , P2_REG3_REG_12_ , P2_REG3_REG_13_ , P2_REG3_REG_14_ , P2_REG3_REG_15_ );
nor nor_14069 ( P2_SUB_605_U55 , P2_REG3_REG_16_ , P2_REG3_REG_17_ );
nor nor_14070 ( P2_SUB_605_U56 , P2_REG3_REG_18_ , P2_REG3_REG_19_ );
nor nor_14071 ( P2_SUB_605_U57 , P2_REG3_REG_20_ , P2_REG3_REG_21_ );
nor nor_14072 ( P2_SUB_605_U58 , P2_REG3_REG_22_ , P2_REG3_REG_23_ );
nor nor_14073 ( P2_SUB_605_U59 , P2_REG3_REG_24_ , P2_REG3_REG_25_ );
nor nor_14074 ( P2_SUB_605_U60 , P2_REG3_REG_26_ , P2_REG3_REG_27_ );
nor nor_14075 ( P2_SUB_605_U61 , P2_REG3_REG_12_ , P2_REG3_REG_13_ );
nor nor_14076 ( P2_SUB_605_U62 , P2_REG3_REG_9_ , P2_REG3_REG_10_ , P2_REG3_REG_8_ );
or OR2_14077 ( P2_SUB_605_U63 , P2_REG3_REG_3_ , P2_REG3_REG_4_ );
or OR3_14078 ( P2_SUB_605_U64 , P2_REG3_REG_4_ , P2_REG3_REG_3_ , P2_REG3_REG_5_ );
or OR4_14079 ( P2_SUB_605_U65 , P2_REG3_REG_5_ , P2_REG3_REG_6_ , P2_REG3_REG_4_ , P2_REG3_REG_3_ );
not NOT1_14080 ( P2_SUB_605_U66 , P2_SUB_605_U32 );
nand NAND2_14081 ( P2_SUB_605_U67 , P2_SUB_605_U66 , P2_SUB_605_U33 );
nand NAND2_14082 ( P2_SUB_605_U68 , P2_SUB_605_U52 , P2_SUB_605_U66 );
nand NAND2_14083 ( P2_SUB_605_U69 , P2_REG3_REG_9_ , P2_SUB_605_U67 );
nand NAND2_14084 ( P2_SUB_605_U70 , P2_REG3_REG_8_ , P2_SUB_605_U32 );
nand NAND2_14085 ( P2_SUB_605_U71 , P2_REG3_REG_7_ , P2_SUB_605_U65 );
nand NAND2_14086 ( P2_SUB_605_U72 , P2_REG3_REG_6_ , P2_SUB_605_U64 );
nand NAND2_14087 ( P2_SUB_605_U73 , P2_REG3_REG_5_ , P2_SUB_605_U63 );
nand NAND2_14088 ( P2_SUB_605_U74 , P2_REG3_REG_4_ , P2_REG3_REG_3_ );
nand NAND2_14089 ( P2_SUB_605_U75 , P2_SUB_605_U62 , P2_SUB_605_U66 );
not NOT1_14090 ( P2_SUB_605_U76 , P2_SUB_605_U34 );
nand NAND2_14091 ( P2_SUB_605_U77 , P2_SUB_605_U76 , P2_SUB_605_U51 );
not NOT1_14092 ( P2_SUB_605_U78 , P2_SUB_605_U49 );
nand NAND2_14093 ( P2_SUB_605_U79 , P2_SUB_605_U78 , P2_SUB_605_U50 );
not NOT1_14094 ( P2_SUB_605_U80 , P2_SUB_605_U35 );
nand NAND2_14095 ( P2_SUB_605_U81 , P2_SUB_605_U80 , P2_SUB_605_U48 );
not NOT1_14096 ( P2_SUB_605_U82 , P2_SUB_605_U36 );
nand NAND2_14097 ( P2_SUB_605_U83 , P2_SUB_605_U82 , P2_SUB_605_U47 );
not NOT1_14098 ( P2_SUB_605_U84 , P2_SUB_605_U37 );
nand NAND2_14099 ( P2_SUB_605_U85 , P2_SUB_605_U84 , P2_SUB_605_U46 );
not NOT1_14100 ( P2_SUB_605_U86 , P2_SUB_605_U38 );
nand NAND2_14101 ( P2_SUB_605_U87 , P2_SUB_605_U86 , P2_SUB_605_U45 );
not NOT1_14102 ( P2_SUB_605_U88 , P2_SUB_605_U39 );
nand NAND2_14103 ( P2_SUB_605_U89 , P2_SUB_605_U88 , P2_SUB_605_U44 );
not NOT1_14104 ( P2_SUB_605_U90 , P2_SUB_605_U40 );
nand NAND2_14105 ( P2_SUB_605_U91 , P2_SUB_605_U90 , P2_SUB_605_U43 );
not NOT1_14106 ( P2_SUB_605_U92 , P2_SUB_605_U41 );
nand NAND2_14107 ( P2_SUB_605_U93 , P2_SUB_605_U92 , P2_SUB_605_U42 );
not NOT1_14108 ( P2_SUB_605_U94 , P2_SUB_605_U93 );
nand NAND2_14109 ( P2_SUB_605_U95 , P2_REG3_REG_28_ , P2_SUB_605_U41 );
nand NAND2_14110 ( P2_SUB_605_U96 , P2_REG3_REG_27_ , P2_SUB_605_U91 );
nand NAND2_14111 ( P2_SUB_605_U97 , P2_REG3_REG_26_ , P2_SUB_605_U40 );
nand NAND2_14112 ( P2_SUB_605_U98 , P2_REG3_REG_25_ , P2_SUB_605_U89 );
nand NAND2_14113 ( P2_SUB_605_U99 , P2_REG3_REG_24_ , P2_SUB_605_U39 );
nand NAND2_14114 ( P2_SUB_605_U100 , P2_REG3_REG_23_ , P2_SUB_605_U87 );
nand NAND2_14115 ( P2_SUB_605_U101 , P2_REG3_REG_22_ , P2_SUB_605_U38 );
nand NAND2_14116 ( P2_SUB_605_U102 , P2_REG3_REG_21_ , P2_SUB_605_U85 );
nand NAND2_14117 ( P2_SUB_605_U103 , P2_REG3_REG_20_ , P2_SUB_605_U37 );
nand NAND2_14118 ( P2_SUB_605_U104 , P2_REG3_REG_19_ , P2_SUB_605_U83 );
nand NAND2_14119 ( P2_SUB_605_U105 , P2_REG3_REG_18_ , P2_SUB_605_U36 );
nand NAND2_14120 ( P2_SUB_605_U106 , P2_REG3_REG_17_ , P2_SUB_605_U81 );
nand NAND2_14121 ( P2_SUB_605_U107 , P2_REG3_REG_16_ , P2_SUB_605_U35 );
nand NAND2_14122 ( P2_SUB_605_U108 , P2_REG3_REG_15_ , P2_SUB_605_U79 );
nand NAND2_14123 ( P2_SUB_605_U109 , P2_REG3_REG_14_ , P2_SUB_605_U49 );
nand NAND2_14124 ( P2_SUB_605_U110 , P2_REG3_REG_13_ , P2_SUB_605_U77 );
nand NAND2_14125 ( P2_SUB_605_U111 , P2_REG3_REG_12_ , P2_SUB_605_U34 );
nand NAND2_14126 ( P2_SUB_605_U112 , P2_REG3_REG_11_ , P2_SUB_605_U75 );
nand NAND2_14127 ( P2_SUB_605_U113 , P2_REG3_REG_10_ , P2_SUB_605_U68 );
and AND2_14128 ( P2_R1095_U6 , P2_R1095_U212 , P2_R1095_U211 );
and AND2_14129 ( P2_R1095_U7 , P2_R1095_U246 , P2_R1095_U245 );
and AND2_14130 ( P2_R1095_U8 , P2_R1095_U193 , P2_R1095_U257 );
and AND2_14131 ( P2_R1095_U9 , P2_R1095_U259 , P2_R1095_U258 );
and AND2_14132 ( P2_R1095_U10 , P2_R1095_U194 , P2_R1095_U281 );
and AND2_14133 ( P2_R1095_U11 , P2_R1095_U283 , P2_R1095_U282 );
and AND2_14134 ( P2_R1095_U12 , P2_R1095_U299 , P2_R1095_U195 );
and AND3_14135 ( P2_R1095_U13 , P2_R1095_U210 , P2_R1095_U197 , P2_R1095_U215 );
and AND2_14136 ( P2_R1095_U14 , P2_R1095_U220 , P2_R1095_U198 );
and AND3_14137 ( P2_R1095_U15 , P2_R1095_U224 , P2_R1095_U192 , P2_R1095_U244 );
and AND2_14138 ( P2_R1095_U16 , P2_R1095_U399 , P2_R1095_U398 );
nand NAND2_14139 ( P2_R1095_U17 , P2_R1095_U331 , P2_R1095_U334 );
nand NAND2_14140 ( P2_R1095_U18 , P2_R1095_U322 , P2_R1095_U325 );
nand NAND2_14141 ( P2_R1095_U19 , P2_R1095_U311 , P2_R1095_U314 );
nand NAND2_14142 ( P2_R1095_U20 , P2_R1095_U305 , P2_R1095_U357 );
nand NAND2_14143 ( P2_R1095_U21 , P2_R1095_U137 , P2_R1095_U186 );
nand NAND2_14144 ( P2_R1095_U22 , P2_R1095_U242 , P2_R1095_U347 );
nand NAND2_14145 ( P2_R1095_U23 , P2_R1095_U235 , P2_R1095_U238 );
nand NAND2_14146 ( P2_R1095_U24 , P2_R1095_U227 , P2_R1095_U229 );
nand NAND2_14147 ( P2_R1095_U25 , P2_R1095_U175 , P2_R1095_U337 );
not NOT1_14148 ( P2_R1095_U26 , P2_U3069 );
nand NAND2_14149 ( P2_R1095_U27 , P2_U3069 , P2_R1095_U32 );
not NOT1_14150 ( P2_R1095_U28 , P2_U3083 );
not NOT1_14151 ( P2_R1095_U29 , P2_U3404 );
not NOT1_14152 ( P2_R1095_U30 , P2_U3407 );
not NOT1_14153 ( P2_R1095_U31 , P2_U3401 );
not NOT1_14154 ( P2_R1095_U32 , P2_U3410 );
not NOT1_14155 ( P2_R1095_U33 , P2_U3413 );
not NOT1_14156 ( P2_R1095_U34 , P2_U3067 );
nand NAND2_14157 ( P2_R1095_U35 , P2_U3067 , P2_R1095_U37 );
not NOT1_14158 ( P2_R1095_U36 , P2_U3063 );
not NOT1_14159 ( P2_R1095_U37 , P2_U3395 );
not NOT1_14160 ( P2_R1095_U38 , P2_U3387 );
not NOT1_14161 ( P2_R1095_U39 , P2_U3077 );
not NOT1_14162 ( P2_R1095_U40 , P2_U3398 );
not NOT1_14163 ( P2_R1095_U41 , P2_U3070 );
not NOT1_14164 ( P2_R1095_U42 , P2_U3066 );
not NOT1_14165 ( P2_R1095_U43 , P2_U3059 );
nand NAND2_14166 ( P2_R1095_U44 , P2_U3059 , P2_R1095_U31 );
nand NAND2_14167 ( P2_R1095_U45 , P2_R1095_U216 , P2_R1095_U214 );
not NOT1_14168 ( P2_R1095_U46 , P2_U3416 );
not NOT1_14169 ( P2_R1095_U47 , P2_U3082 );
nand NAND2_14170 ( P2_R1095_U48 , P2_R1095_U45 , P2_R1095_U217 );
nand NAND2_14171 ( P2_R1095_U49 , P2_R1095_U44 , P2_R1095_U231 );
nand NAND3_14172 ( P2_R1095_U50 , P2_R1095_U204 , P2_R1095_U188 , P2_R1095_U338 );
not NOT1_14173 ( P2_R1095_U51 , P2_U3895 );
not NOT1_14174 ( P2_R1095_U52 , P2_U3056 );
nand NAND2_14175 ( P2_R1095_U53 , P2_U3056 , P2_R1095_U90 );
not NOT1_14176 ( P2_R1095_U54 , P2_U3052 );
not NOT1_14177 ( P2_R1095_U55 , P2_U3071 );
not NOT1_14178 ( P2_R1095_U56 , P2_U3062 );
not NOT1_14179 ( P2_R1095_U57 , P2_U3061 );
not NOT1_14180 ( P2_R1095_U58 , P2_U3419 );
nand NAND2_14181 ( P2_R1095_U59 , P2_U3082 , P2_R1095_U46 );
not NOT1_14182 ( P2_R1095_U60 , P2_U3422 );
not NOT1_14183 ( P2_R1095_U61 , P2_U3425 );
nand NAND2_14184 ( P2_R1095_U62 , P2_R1095_U249 , P2_R1095_U248 );
not NOT1_14185 ( P2_R1095_U63 , P2_U3428 );
not NOT1_14186 ( P2_R1095_U64 , P2_U3079 );
not NOT1_14187 ( P2_R1095_U65 , P2_U3437 );
not NOT1_14188 ( P2_R1095_U66 , P2_U3434 );
not NOT1_14189 ( P2_R1095_U67 , P2_U3431 );
not NOT1_14190 ( P2_R1095_U68 , P2_U3072 );
not NOT1_14191 ( P2_R1095_U69 , P2_U3073 );
not NOT1_14192 ( P2_R1095_U70 , P2_U3078 );
nand NAND2_14193 ( P2_R1095_U71 , P2_U3078 , P2_R1095_U67 );
not NOT1_14194 ( P2_R1095_U72 , P2_U3440 );
not NOT1_14195 ( P2_R1095_U73 , P2_U3068 );
not NOT1_14196 ( P2_R1095_U74 , P2_U3081 );
not NOT1_14197 ( P2_R1095_U75 , P2_U3445 );
not NOT1_14198 ( P2_R1095_U76 , P2_U3080 );
not NOT1_14199 ( P2_R1095_U77 , P2_U3903 );
not NOT1_14200 ( P2_R1095_U78 , P2_U3075 );
not NOT1_14201 ( P2_R1095_U79 , P2_U3900 );
not NOT1_14202 ( P2_R1095_U80 , P2_U3901 );
not NOT1_14203 ( P2_R1095_U81 , P2_U3902 );
not NOT1_14204 ( P2_R1095_U82 , P2_U3065 );
not NOT1_14205 ( P2_R1095_U83 , P2_U3060 );
not NOT1_14206 ( P2_R1095_U84 , P2_U3074 );
nand NAND2_14207 ( P2_R1095_U85 , P2_U3074 , P2_R1095_U81 );
not NOT1_14208 ( P2_R1095_U86 , P2_U3899 );
not NOT1_14209 ( P2_R1095_U87 , P2_U3064 );
not NOT1_14210 ( P2_R1095_U88 , P2_U3898 );
not NOT1_14211 ( P2_R1095_U89 , P2_U3057 );
not NOT1_14212 ( P2_R1095_U90 , P2_U3897 );
not NOT1_14213 ( P2_R1095_U91 , P2_U3896 );
not NOT1_14214 ( P2_R1095_U92 , P2_U3053 );
nand NAND2_14215 ( P2_R1095_U93 , P2_R1095_U297 , P2_R1095_U296 );
nand NAND2_14216 ( P2_R1095_U94 , P2_R1095_U85 , P2_R1095_U307 );
nand NAND2_14217 ( P2_R1095_U95 , P2_R1095_U71 , P2_R1095_U318 );
nand NAND2_14218 ( P2_R1095_U96 , P2_R1095_U349 , P2_R1095_U59 );
not NOT1_14219 ( P2_R1095_U97 , P2_U3076 );
nand NAND2_14220 ( P2_R1095_U98 , P2_R1095_U406 , P2_R1095_U405 );
nand NAND2_14221 ( P2_R1095_U99 , P2_R1095_U420 , P2_R1095_U419 );
nand NAND2_14222 ( P2_R1095_U100 , P2_R1095_U425 , P2_R1095_U424 );
nand NAND2_14223 ( P2_R1095_U101 , P2_R1095_U441 , P2_R1095_U440 );
nand NAND2_14224 ( P2_R1095_U102 , P2_R1095_U446 , P2_R1095_U445 );
nand NAND2_14225 ( P2_R1095_U103 , P2_R1095_U451 , P2_R1095_U450 );
nand NAND2_14226 ( P2_R1095_U104 , P2_R1095_U456 , P2_R1095_U455 );
nand NAND2_14227 ( P2_R1095_U105 , P2_R1095_U461 , P2_R1095_U460 );
nand NAND2_14228 ( P2_R1095_U106 , P2_R1095_U477 , P2_R1095_U476 );
nand NAND2_14229 ( P2_R1095_U107 , P2_R1095_U482 , P2_R1095_U481 );
nand NAND2_14230 ( P2_R1095_U108 , P2_R1095_U365 , P2_R1095_U364 );
nand NAND2_14231 ( P2_R1095_U109 , P2_R1095_U374 , P2_R1095_U373 );
nand NAND2_14232 ( P2_R1095_U110 , P2_R1095_U381 , P2_R1095_U380 );
nand NAND2_14233 ( P2_R1095_U111 , P2_R1095_U385 , P2_R1095_U384 );
nand NAND2_14234 ( P2_R1095_U112 , P2_R1095_U394 , P2_R1095_U393 );
nand NAND2_14235 ( P2_R1095_U113 , P2_R1095_U415 , P2_R1095_U414 );
nand NAND2_14236 ( P2_R1095_U114 , P2_R1095_U432 , P2_R1095_U431 );
nand NAND2_14237 ( P2_R1095_U115 , P2_R1095_U436 , P2_R1095_U435 );
nand NAND2_14238 ( P2_R1095_U116 , P2_R1095_U468 , P2_R1095_U467 );
nand NAND2_14239 ( P2_R1095_U117 , P2_R1095_U472 , P2_R1095_U471 );
nand NAND2_14240 ( P2_R1095_U118 , P2_R1095_U489 , P2_R1095_U488 );
and AND2_14241 ( P2_R1095_U119 , P2_R1095_U206 , P2_R1095_U196 );
and AND2_14242 ( P2_R1095_U120 , P2_R1095_U209 , P2_R1095_U208 );
and AND2_14243 ( P2_R1095_U121 , P2_R1095_U14 , P2_R1095_U13 );
and AND2_14244 ( P2_R1095_U122 , P2_R1095_U340 , P2_R1095_U222 );
and AND2_14245 ( P2_R1095_U123 , P2_R1095_U342 , P2_R1095_U122 );
and AND3_14246 ( P2_R1095_U124 , P2_R1095_U367 , P2_R1095_U366 , P2_R1095_U27 );
and AND2_14247 ( P2_R1095_U125 , P2_R1095_U370 , P2_R1095_U198 );
and AND2_14248 ( P2_R1095_U126 , P2_R1095_U237 , P2_R1095_U6 );
and AND2_14249 ( P2_R1095_U127 , P2_R1095_U377 , P2_R1095_U197 );
and AND3_14250 ( P2_R1095_U128 , P2_R1095_U387 , P2_R1095_U386 , P2_R1095_U35 );
and AND2_14251 ( P2_R1095_U129 , P2_R1095_U390 , P2_R1095_U196 );
and AND2_14252 ( P2_R1095_U130 , P2_R1095_U251 , P2_R1095_U15 );
and AND2_14253 ( P2_R1095_U131 , P2_R1095_U343 , P2_R1095_U252 );
and AND2_14254 ( P2_R1095_U132 , P2_R1095_U262 , P2_R1095_U8 );
and AND2_14255 ( P2_R1095_U133 , P2_R1095_U286 , P2_R1095_U10 );
and AND2_14256 ( P2_R1095_U134 , P2_R1095_U302 , P2_R1095_U301 );
and AND2_14257 ( P2_R1095_U135 , P2_R1095_U397 , P2_R1095_U303 );
and AND4_14258 ( P2_R1095_U136 , P2_R1095_U302 , P2_R1095_U301 , P2_R1095_U304 , P2_R1095_U16 );
and AND2_14259 ( P2_R1095_U137 , P2_R1095_U359 , P2_R1095_U165 );
nand NAND2_14260 ( P2_R1095_U138 , P2_R1095_U403 , P2_R1095_U402 );
and AND3_14261 ( P2_R1095_U139 , P2_R1095_U408 , P2_R1095_U407 , P2_R1095_U53 );
and AND2_14262 ( P2_R1095_U140 , P2_R1095_U411 , P2_R1095_U195 );
nand NAND2_14263 ( P2_R1095_U141 , P2_R1095_U417 , P2_R1095_U416 );
nand NAND2_14264 ( P2_R1095_U142 , P2_R1095_U422 , P2_R1095_U421 );
and AND2_14265 ( P2_R1095_U143 , P2_R1095_U313 , P2_R1095_U11 );
and AND2_14266 ( P2_R1095_U144 , P2_R1095_U428 , P2_R1095_U194 );
nand NAND2_14267 ( P2_R1095_U145 , P2_R1095_U438 , P2_R1095_U437 );
nand NAND2_14268 ( P2_R1095_U146 , P2_R1095_U443 , P2_R1095_U442 );
nand NAND2_14269 ( P2_R1095_U147 , P2_R1095_U448 , P2_R1095_U447 );
nand NAND2_14270 ( P2_R1095_U148 , P2_R1095_U453 , P2_R1095_U452 );
nand NAND2_14271 ( P2_R1095_U149 , P2_R1095_U458 , P2_R1095_U457 );
and AND2_14272 ( P2_R1095_U150 , P2_R1095_U324 , P2_R1095_U9 );
and AND2_14273 ( P2_R1095_U151 , P2_R1095_U464 , P2_R1095_U193 );
nand NAND2_14274 ( P2_R1095_U152 , P2_R1095_U474 , P2_R1095_U473 );
nand NAND2_14275 ( P2_R1095_U153 , P2_R1095_U479 , P2_R1095_U478 );
and AND2_14276 ( P2_R1095_U154 , P2_R1095_U333 , P2_R1095_U7 );
and AND2_14277 ( P2_R1095_U155 , P2_R1095_U485 , P2_R1095_U192 );
and AND2_14278 ( P2_R1095_U156 , P2_R1095_U363 , P2_R1095_U362 );
nand NAND2_14279 ( P2_R1095_U157 , P2_R1095_U123 , P2_R1095_U341 );
and AND2_14280 ( P2_R1095_U158 , P2_R1095_U372 , P2_R1095_U371 );
and AND2_14281 ( P2_R1095_U159 , P2_R1095_U379 , P2_R1095_U378 );
and AND2_14282 ( P2_R1095_U160 , P2_R1095_U383 , P2_R1095_U382 );
nand NAND2_14283 ( P2_R1095_U161 , P2_R1095_U120 , P2_R1095_U344 );
and AND2_14284 ( P2_R1095_U162 , P2_R1095_U392 , P2_R1095_U391 );
not NOT1_14285 ( P2_R1095_U163 , P2_U3904 );
not NOT1_14286 ( P2_R1095_U164 , P2_U3054 );
and AND2_14287 ( P2_R1095_U165 , P2_R1095_U401 , P2_R1095_U400 );
nand NAND2_14288 ( P2_R1095_U166 , P2_R1095_U134 , P2_R1095_U360 );
and AND2_14289 ( P2_R1095_U167 , P2_R1095_U413 , P2_R1095_U412 );
nand NAND2_14290 ( P2_R1095_U168 , P2_R1095_U293 , P2_R1095_U292 );
nand NAND2_14291 ( P2_R1095_U169 , P2_R1095_U289 , P2_R1095_U288 );
and AND2_14292 ( P2_R1095_U170 , P2_R1095_U430 , P2_R1095_U429 );
and AND2_14293 ( P2_R1095_U171 , P2_R1095_U434 , P2_R1095_U433 );
nand NAND2_14294 ( P2_R1095_U172 , P2_R1095_U279 , P2_R1095_U278 );
nand NAND2_14295 ( P2_R1095_U173 , P2_R1095_U275 , P2_R1095_U274 );
not NOT1_14296 ( P2_R1095_U174 , P2_U3392 );
nand NAND2_14297 ( P2_R1095_U175 , P2_U3387 , P2_R1095_U97 );
nand NAND3_14298 ( P2_R1095_U176 , P2_R1095_U271 , P2_R1095_U187 , P2_R1095_U339 );
not NOT1_14299 ( P2_R1095_U177 , P2_U3443 );
nand NAND2_14300 ( P2_R1095_U178 , P2_R1095_U269 , P2_R1095_U268 );
nand NAND2_14301 ( P2_R1095_U179 , P2_R1095_U265 , P2_R1095_U264 );
and AND2_14302 ( P2_R1095_U180 , P2_R1095_U466 , P2_R1095_U465 );
and AND2_14303 ( P2_R1095_U181 , P2_R1095_U470 , P2_R1095_U469 );
nand NAND2_14304 ( P2_R1095_U182 , P2_R1095_U255 , P2_R1095_U254 );
nand NAND2_14305 ( P2_R1095_U183 , P2_R1095_U131 , P2_R1095_U353 );
nand NAND2_14306 ( P2_R1095_U184 , P2_R1095_U351 , P2_R1095_U62 );
and AND2_14307 ( P2_R1095_U185 , P2_R1095_U487 , P2_R1095_U486 );
nand NAND2_14308 ( P2_R1095_U186 , P2_R1095_U135 , P2_R1095_U166 );
nand NAND2_14309 ( P2_R1095_U187 , P2_R1095_U178 , P2_R1095_U177 );
nand NAND2_14310 ( P2_R1095_U188 , P2_R1095_U175 , P2_R1095_U174 );
not NOT1_14311 ( P2_R1095_U189 , P2_R1095_U53 );
not NOT1_14312 ( P2_R1095_U190 , P2_R1095_U35 );
not NOT1_14313 ( P2_R1095_U191 , P2_R1095_U27 );
nand NAND2_14314 ( P2_R1095_U192 , P2_U3419 , P2_R1095_U57 );
nand NAND2_14315 ( P2_R1095_U193 , P2_U3434 , P2_R1095_U69 );
nand NAND2_14316 ( P2_R1095_U194 , P2_U3901 , P2_R1095_U83 );
nand NAND2_14317 ( P2_R1095_U195 , P2_U3897 , P2_R1095_U52 );
nand NAND2_14318 ( P2_R1095_U196 , P2_U3395 , P2_R1095_U34 );
nand NAND2_14319 ( P2_R1095_U197 , P2_U3404 , P2_R1095_U42 );
nand NAND2_14320 ( P2_R1095_U198 , P2_U3410 , P2_R1095_U26 );
not NOT1_14321 ( P2_R1095_U199 , P2_R1095_U71 );
not NOT1_14322 ( P2_R1095_U200 , P2_R1095_U85 );
not NOT1_14323 ( P2_R1095_U201 , P2_R1095_U44 );
not NOT1_14324 ( P2_R1095_U202 , P2_R1095_U59 );
not NOT1_14325 ( P2_R1095_U203 , P2_R1095_U175 );
nand NAND2_14326 ( P2_R1095_U204 , P2_U3077 , P2_R1095_U175 );
not NOT1_14327 ( P2_R1095_U205 , P2_R1095_U50 );
nand NAND2_14328 ( P2_R1095_U206 , P2_U3398 , P2_R1095_U36 );
nand NAND2_14329 ( P2_R1095_U207 , P2_R1095_U36 , P2_R1095_U35 );
nand NAND2_14330 ( P2_R1095_U208 , P2_R1095_U207 , P2_R1095_U40 );
nand NAND2_14331 ( P2_R1095_U209 , P2_U3063 , P2_R1095_U190 );
nand NAND2_14332 ( P2_R1095_U210 , P2_U3407 , P2_R1095_U41 );
nand NAND2_14333 ( P2_R1095_U211 , P2_U3070 , P2_R1095_U30 );
nand NAND2_14334 ( P2_R1095_U212 , P2_U3066 , P2_R1095_U29 );
nand NAND2_14335 ( P2_R1095_U213 , P2_R1095_U201 , P2_R1095_U197 );
nand NAND2_14336 ( P2_R1095_U214 , P2_R1095_U6 , P2_R1095_U213 );
nand NAND2_14337 ( P2_R1095_U215 , P2_U3401 , P2_R1095_U43 );
nand NAND2_14338 ( P2_R1095_U216 , P2_U3407 , P2_R1095_U41 );
nand NAND2_14339 ( P2_R1095_U217 , P2_R1095_U13 , P2_R1095_U161 );
not NOT1_14340 ( P2_R1095_U218 , P2_R1095_U45 );
not NOT1_14341 ( P2_R1095_U219 , P2_R1095_U48 );
nand NAND2_14342 ( P2_R1095_U220 , P2_U3413 , P2_R1095_U28 );
nand NAND2_14343 ( P2_R1095_U221 , P2_R1095_U28 , P2_R1095_U27 );
nand NAND2_14344 ( P2_R1095_U222 , P2_U3083 , P2_R1095_U191 );
not NOT1_14345 ( P2_R1095_U223 , P2_R1095_U157 );
nand NAND2_14346 ( P2_R1095_U224 , P2_U3416 , P2_R1095_U47 );
nand NAND2_14347 ( P2_R1095_U225 , P2_R1095_U224 , P2_R1095_U59 );
nand NAND2_14348 ( P2_R1095_U226 , P2_R1095_U219 , P2_R1095_U27 );
nand NAND2_14349 ( P2_R1095_U227 , P2_R1095_U125 , P2_R1095_U226 );
nand NAND2_14350 ( P2_R1095_U228 , P2_R1095_U48 , P2_R1095_U198 );
nand NAND2_14351 ( P2_R1095_U229 , P2_R1095_U124 , P2_R1095_U228 );
nand NAND2_14352 ( P2_R1095_U230 , P2_R1095_U27 , P2_R1095_U198 );
nand NAND2_14353 ( P2_R1095_U231 , P2_R1095_U215 , P2_R1095_U161 );
not NOT1_14354 ( P2_R1095_U232 , P2_R1095_U49 );
nand NAND2_14355 ( P2_R1095_U233 , P2_U3066 , P2_R1095_U29 );
nand NAND2_14356 ( P2_R1095_U234 , P2_R1095_U232 , P2_R1095_U233 );
nand NAND2_14357 ( P2_R1095_U235 , P2_R1095_U127 , P2_R1095_U234 );
nand NAND2_14358 ( P2_R1095_U236 , P2_R1095_U49 , P2_R1095_U197 );
nand NAND2_14359 ( P2_R1095_U237 , P2_U3407 , P2_R1095_U41 );
nand NAND2_14360 ( P2_R1095_U238 , P2_R1095_U126 , P2_R1095_U236 );
nand NAND2_14361 ( P2_R1095_U239 , P2_U3066 , P2_R1095_U29 );
nand NAND2_14362 ( P2_R1095_U240 , P2_R1095_U239 , P2_R1095_U197 );
nand NAND2_14363 ( P2_R1095_U241 , P2_R1095_U215 , P2_R1095_U44 );
nand NAND2_14364 ( P2_R1095_U242 , P2_R1095_U129 , P2_R1095_U348 );
nand NAND2_14365 ( P2_R1095_U243 , P2_R1095_U35 , P2_R1095_U196 );
nand NAND2_14366 ( P2_R1095_U244 , P2_U3422 , P2_R1095_U56 );
nand NAND2_14367 ( P2_R1095_U245 , P2_U3062 , P2_R1095_U60 );
nand NAND2_14368 ( P2_R1095_U246 , P2_U3061 , P2_R1095_U58 );
nand NAND2_14369 ( P2_R1095_U247 , P2_R1095_U202 , P2_R1095_U192 );
nand NAND2_14370 ( P2_R1095_U248 , P2_R1095_U7 , P2_R1095_U247 );
nand NAND2_14371 ( P2_R1095_U249 , P2_U3422 , P2_R1095_U56 );
not NOT1_14372 ( P2_R1095_U250 , P2_R1095_U62 );
nand NAND2_14373 ( P2_R1095_U251 , P2_U3425 , P2_R1095_U55 );
nand NAND2_14374 ( P2_R1095_U252 , P2_U3071 , P2_R1095_U61 );
nand NAND2_14375 ( P2_R1095_U253 , P2_U3428 , P2_R1095_U64 );
nand NAND2_14376 ( P2_R1095_U254 , P2_R1095_U253 , P2_R1095_U183 );
nand NAND2_14377 ( P2_R1095_U255 , P2_U3079 , P2_R1095_U63 );
not NOT1_14378 ( P2_R1095_U256 , P2_R1095_U182 );
nand NAND2_14379 ( P2_R1095_U257 , P2_U3437 , P2_R1095_U68 );
nand NAND2_14380 ( P2_R1095_U258 , P2_U3072 , P2_R1095_U65 );
nand NAND2_14381 ( P2_R1095_U259 , P2_U3073 , P2_R1095_U66 );
nand NAND2_14382 ( P2_R1095_U260 , P2_R1095_U199 , P2_R1095_U8 );
nand NAND2_14383 ( P2_R1095_U261 , P2_R1095_U9 , P2_R1095_U260 );
nand NAND2_14384 ( P2_R1095_U262 , P2_U3431 , P2_R1095_U70 );
nand NAND2_14385 ( P2_R1095_U263 , P2_U3437 , P2_R1095_U68 );
nand NAND2_14386 ( P2_R1095_U264 , P2_R1095_U132 , P2_R1095_U182 );
nand NAND2_14387 ( P2_R1095_U265 , P2_R1095_U263 , P2_R1095_U261 );
not NOT1_14388 ( P2_R1095_U266 , P2_R1095_U179 );
nand NAND2_14389 ( P2_R1095_U267 , P2_U3440 , P2_R1095_U73 );
nand NAND2_14390 ( P2_R1095_U268 , P2_R1095_U267 , P2_R1095_U179 );
nand NAND2_14391 ( P2_R1095_U269 , P2_U3068 , P2_R1095_U72 );
not NOT1_14392 ( P2_R1095_U270 , P2_R1095_U178 );
nand NAND2_14393 ( P2_R1095_U271 , P2_U3081 , P2_R1095_U178 );
not NOT1_14394 ( P2_R1095_U272 , P2_R1095_U176 );
nand NAND2_14395 ( P2_R1095_U273 , P2_U3445 , P2_R1095_U76 );
nand NAND2_14396 ( P2_R1095_U274 , P2_R1095_U273 , P2_R1095_U176 );
nand NAND2_14397 ( P2_R1095_U275 , P2_U3080 , P2_R1095_U75 );
not NOT1_14398 ( P2_R1095_U276 , P2_R1095_U173 );
nand NAND2_14399 ( P2_R1095_U277 , P2_U3903 , P2_R1095_U78 );
nand NAND2_14400 ( P2_R1095_U278 , P2_R1095_U277 , P2_R1095_U173 );
nand NAND2_14401 ( P2_R1095_U279 , P2_U3075 , P2_R1095_U77 );
not NOT1_14402 ( P2_R1095_U280 , P2_R1095_U172 );
nand NAND2_14403 ( P2_R1095_U281 , P2_U3900 , P2_R1095_U82 );
nand NAND2_14404 ( P2_R1095_U282 , P2_U3065 , P2_R1095_U79 );
nand NAND2_14405 ( P2_R1095_U283 , P2_U3060 , P2_R1095_U80 );
nand NAND2_14406 ( P2_R1095_U284 , P2_R1095_U200 , P2_R1095_U10 );
nand NAND2_14407 ( P2_R1095_U285 , P2_R1095_U11 , P2_R1095_U284 );
nand NAND2_14408 ( P2_R1095_U286 , P2_U3902 , P2_R1095_U84 );
nand NAND2_14409 ( P2_R1095_U287 , P2_U3900 , P2_R1095_U82 );
nand NAND2_14410 ( P2_R1095_U288 , P2_R1095_U133 , P2_R1095_U172 );
nand NAND2_14411 ( P2_R1095_U289 , P2_R1095_U287 , P2_R1095_U285 );
not NOT1_14412 ( P2_R1095_U290 , P2_R1095_U169 );
nand NAND2_14413 ( P2_R1095_U291 , P2_U3899 , P2_R1095_U87 );
nand NAND2_14414 ( P2_R1095_U292 , P2_R1095_U291 , P2_R1095_U169 );
nand NAND2_14415 ( P2_R1095_U293 , P2_U3064 , P2_R1095_U86 );
not NOT1_14416 ( P2_R1095_U294 , P2_R1095_U168 );
nand NAND2_14417 ( P2_R1095_U295 , P2_U3898 , P2_R1095_U89 );
nand NAND2_14418 ( P2_R1095_U296 , P2_R1095_U295 , P2_R1095_U168 );
nand NAND2_14419 ( P2_R1095_U297 , P2_U3057 , P2_R1095_U88 );
not NOT1_14420 ( P2_R1095_U298 , P2_R1095_U93 );
nand NAND2_14421 ( P2_R1095_U299 , P2_U3896 , P2_R1095_U54 );
nand NAND2_14422 ( P2_R1095_U300 , P2_R1095_U54 , P2_R1095_U53 );
nand NAND2_14423 ( P2_R1095_U301 , P2_R1095_U300 , P2_R1095_U91 );
nand NAND2_14424 ( P2_R1095_U302 , P2_U3052 , P2_R1095_U189 );
nand NAND2_14425 ( P2_R1095_U303 , P2_U3895 , P2_R1095_U92 );
nand NAND2_14426 ( P2_R1095_U304 , P2_U3053 , P2_R1095_U51 );
nand NAND2_14427 ( P2_R1095_U305 , P2_R1095_U140 , P2_R1095_U355 );
nand NAND2_14428 ( P2_R1095_U306 , P2_R1095_U53 , P2_R1095_U195 );
nand NAND2_14429 ( P2_R1095_U307 , P2_R1095_U286 , P2_R1095_U172 );
not NOT1_14430 ( P2_R1095_U308 , P2_R1095_U94 );
nand NAND2_14431 ( P2_R1095_U309 , P2_U3060 , P2_R1095_U80 );
nand NAND2_14432 ( P2_R1095_U310 , P2_R1095_U308 , P2_R1095_U309 );
nand NAND2_14433 ( P2_R1095_U311 , P2_R1095_U144 , P2_R1095_U310 );
nand NAND2_14434 ( P2_R1095_U312 , P2_R1095_U94 , P2_R1095_U194 );
nand NAND2_14435 ( P2_R1095_U313 , P2_U3900 , P2_R1095_U82 );
nand NAND2_14436 ( P2_R1095_U314 , P2_R1095_U143 , P2_R1095_U312 );
nand NAND2_14437 ( P2_R1095_U315 , P2_U3060 , P2_R1095_U80 );
nand NAND2_14438 ( P2_R1095_U316 , P2_R1095_U194 , P2_R1095_U315 );
nand NAND2_14439 ( P2_R1095_U317 , P2_R1095_U286 , P2_R1095_U85 );
nand NAND2_14440 ( P2_R1095_U318 , P2_R1095_U262 , P2_R1095_U182 );
not NOT1_14441 ( P2_R1095_U319 , P2_R1095_U95 );
nand NAND2_14442 ( P2_R1095_U320 , P2_U3073 , P2_R1095_U66 );
nand NAND2_14443 ( P2_R1095_U321 , P2_R1095_U319 , P2_R1095_U320 );
nand NAND2_14444 ( P2_R1095_U322 , P2_R1095_U151 , P2_R1095_U321 );
nand NAND2_14445 ( P2_R1095_U323 , P2_R1095_U95 , P2_R1095_U193 );
nand NAND2_14446 ( P2_R1095_U324 , P2_U3437 , P2_R1095_U68 );
nand NAND2_14447 ( P2_R1095_U325 , P2_R1095_U150 , P2_R1095_U323 );
nand NAND2_14448 ( P2_R1095_U326 , P2_U3073 , P2_R1095_U66 );
nand NAND2_14449 ( P2_R1095_U327 , P2_R1095_U193 , P2_R1095_U326 );
nand NAND2_14450 ( P2_R1095_U328 , P2_R1095_U262 , P2_R1095_U71 );
nand NAND2_14451 ( P2_R1095_U329 , P2_U3061 , P2_R1095_U58 );
nand NAND2_14452 ( P2_R1095_U330 , P2_R1095_U350 , P2_R1095_U329 );
nand NAND2_14453 ( P2_R1095_U331 , P2_R1095_U155 , P2_R1095_U330 );
nand NAND2_14454 ( P2_R1095_U332 , P2_R1095_U96 , P2_R1095_U192 );
nand NAND2_14455 ( P2_R1095_U333 , P2_U3422 , P2_R1095_U56 );
nand NAND2_14456 ( P2_R1095_U334 , P2_R1095_U154 , P2_R1095_U332 );
nand NAND2_14457 ( P2_R1095_U335 , P2_U3061 , P2_R1095_U58 );
nand NAND2_14458 ( P2_R1095_U336 , P2_R1095_U192 , P2_R1095_U335 );
nand NAND2_14459 ( P2_R1095_U337 , P2_U3076 , P2_R1095_U38 );
nand NAND2_14460 ( P2_R1095_U338 , P2_U3077 , P2_R1095_U174 );
nand NAND2_14461 ( P2_R1095_U339 , P2_U3081 , P2_R1095_U177 );
nand NAND2_14462 ( P2_R1095_U340 , P2_R1095_U33 , P2_R1095_U221 );
nand NAND2_14463 ( P2_R1095_U341 , P2_R1095_U121 , P2_R1095_U161 );
nand NAND2_14464 ( P2_R1095_U342 , P2_R1095_U218 , P2_R1095_U14 );
nand NAND2_14465 ( P2_R1095_U343 , P2_R1095_U250 , P2_R1095_U251 );
nand NAND2_14466 ( P2_R1095_U344 , P2_R1095_U119 , P2_R1095_U50 );
not NOT1_14467 ( P2_R1095_U345 , P2_R1095_U161 );
nand NAND2_14468 ( P2_R1095_U346 , P2_R1095_U196 , P2_R1095_U50 );
nand NAND2_14469 ( P2_R1095_U347 , P2_R1095_U128 , P2_R1095_U346 );
nand NAND2_14470 ( P2_R1095_U348 , P2_R1095_U205 , P2_R1095_U35 );
nand NAND2_14471 ( P2_R1095_U349 , P2_R1095_U224 , P2_R1095_U157 );
not NOT1_14472 ( P2_R1095_U350 , P2_R1095_U96 );
nand NAND2_14473 ( P2_R1095_U351 , P2_R1095_U15 , P2_R1095_U157 );
not NOT1_14474 ( P2_R1095_U352 , P2_R1095_U184 );
nand NAND2_14475 ( P2_R1095_U353 , P2_R1095_U130 , P2_R1095_U157 );
not NOT1_14476 ( P2_R1095_U354 , P2_R1095_U183 );
nand NAND2_14477 ( P2_R1095_U355 , P2_R1095_U298 , P2_R1095_U53 );
nand NAND2_14478 ( P2_R1095_U356 , P2_R1095_U195 , P2_R1095_U93 );
nand NAND2_14479 ( P2_R1095_U357 , P2_R1095_U139 , P2_R1095_U356 );
nand NAND2_14480 ( P2_R1095_U358 , P2_R1095_U12 , P2_R1095_U93 );
nand NAND2_14481 ( P2_R1095_U359 , P2_R1095_U136 , P2_R1095_U358 );
nand NAND2_14482 ( P2_R1095_U360 , P2_R1095_U12 , P2_R1095_U93 );
not NOT1_14483 ( P2_R1095_U361 , P2_R1095_U166 );
nand NAND2_14484 ( P2_R1095_U362 , P2_U3416 , P2_R1095_U47 );
nand NAND2_14485 ( P2_R1095_U363 , P2_U3082 , P2_R1095_U46 );
nand NAND2_14486 ( P2_R1095_U364 , P2_R1095_U225 , P2_R1095_U157 );
nand NAND2_14487 ( P2_R1095_U365 , P2_R1095_U223 , P2_R1095_U156 );
nand NAND2_14488 ( P2_R1095_U366 , P2_U3413 , P2_R1095_U28 );
nand NAND2_14489 ( P2_R1095_U367 , P2_U3083 , P2_R1095_U33 );
nand NAND2_14490 ( P2_R1095_U368 , P2_U3413 , P2_R1095_U28 );
nand NAND2_14491 ( P2_R1095_U369 , P2_U3083 , P2_R1095_U33 );
nand NAND2_14492 ( P2_R1095_U370 , P2_R1095_U369 , P2_R1095_U368 );
nand NAND2_14493 ( P2_R1095_U371 , P2_U3410 , P2_R1095_U26 );
nand NAND2_14494 ( P2_R1095_U372 , P2_U3069 , P2_R1095_U32 );
nand NAND2_14495 ( P2_R1095_U373 , P2_R1095_U230 , P2_R1095_U48 );
nand NAND2_14496 ( P2_R1095_U374 , P2_R1095_U158 , P2_R1095_U219 );
nand NAND2_14497 ( P2_R1095_U375 , P2_U3407 , P2_R1095_U41 );
nand NAND2_14498 ( P2_R1095_U376 , P2_U3070 , P2_R1095_U30 );
nand NAND2_14499 ( P2_R1095_U377 , P2_R1095_U376 , P2_R1095_U375 );
nand NAND2_14500 ( P2_R1095_U378 , P2_U3404 , P2_R1095_U42 );
nand NAND2_14501 ( P2_R1095_U379 , P2_U3066 , P2_R1095_U29 );
nand NAND2_14502 ( P2_R1095_U380 , P2_R1095_U240 , P2_R1095_U49 );
nand NAND2_14503 ( P2_R1095_U381 , P2_R1095_U159 , P2_R1095_U232 );
nand NAND2_14504 ( P2_R1095_U382 , P2_U3401 , P2_R1095_U43 );
nand NAND2_14505 ( P2_R1095_U383 , P2_U3059 , P2_R1095_U31 );
nand NAND2_14506 ( P2_R1095_U384 , P2_R1095_U161 , P2_R1095_U241 );
nand NAND2_14507 ( P2_R1095_U385 , P2_R1095_U345 , P2_R1095_U160 );
nand NAND2_14508 ( P2_R1095_U386 , P2_U3398 , P2_R1095_U36 );
nand NAND2_14509 ( P2_R1095_U387 , P2_U3063 , P2_R1095_U40 );
nand NAND2_14510 ( P2_R1095_U388 , P2_U3398 , P2_R1095_U36 );
nand NAND2_14511 ( P2_R1095_U389 , P2_U3063 , P2_R1095_U40 );
nand NAND2_14512 ( P2_R1095_U390 , P2_R1095_U389 , P2_R1095_U388 );
nand NAND2_14513 ( P2_R1095_U391 , P2_U3395 , P2_R1095_U34 );
nand NAND2_14514 ( P2_R1095_U392 , P2_U3067 , P2_R1095_U37 );
nand NAND2_14515 ( P2_R1095_U393 , P2_R1095_U243 , P2_R1095_U50 );
nand NAND2_14516 ( P2_R1095_U394 , P2_R1095_U162 , P2_R1095_U205 );
nand NAND2_14517 ( P2_R1095_U395 , P2_U3904 , P2_R1095_U164 );
nand NAND2_14518 ( P2_R1095_U396 , P2_U3054 , P2_R1095_U163 );
nand NAND2_14519 ( P2_R1095_U397 , P2_R1095_U396 , P2_R1095_U395 );
nand NAND2_14520 ( P2_R1095_U398 , P2_U3904 , P2_R1095_U164 );
nand NAND2_14521 ( P2_R1095_U399 , P2_U3054 , P2_R1095_U163 );
nand NAND3_14522 ( P2_R1095_U400 , P2_U3053 , P2_R1095_U397 , P2_R1095_U51 );
nand NAND3_14523 ( P2_R1095_U401 , P2_R1095_U16 , P2_R1095_U92 , P2_U3895 );
nand NAND2_14524 ( P2_R1095_U402 , P2_U3895 , P2_R1095_U92 );
nand NAND2_14525 ( P2_R1095_U403 , P2_U3053 , P2_R1095_U51 );
not NOT1_14526 ( P2_R1095_U404 , P2_R1095_U138 );
nand NAND2_14527 ( P2_R1095_U405 , P2_R1095_U361 , P2_R1095_U404 );
nand NAND2_14528 ( P2_R1095_U406 , P2_R1095_U138 , P2_R1095_U166 );
nand NAND2_14529 ( P2_R1095_U407 , P2_U3896 , P2_R1095_U54 );
nand NAND2_14530 ( P2_R1095_U408 , P2_U3052 , P2_R1095_U91 );
nand NAND2_14531 ( P2_R1095_U409 , P2_U3896 , P2_R1095_U54 );
nand NAND2_14532 ( P2_R1095_U410 , P2_U3052 , P2_R1095_U91 );
nand NAND2_14533 ( P2_R1095_U411 , P2_R1095_U410 , P2_R1095_U409 );
nand NAND2_14534 ( P2_R1095_U412 , P2_U3897 , P2_R1095_U52 );
nand NAND2_14535 ( P2_R1095_U413 , P2_U3056 , P2_R1095_U90 );
nand NAND2_14536 ( P2_R1095_U414 , P2_R1095_U306 , P2_R1095_U93 );
nand NAND2_14537 ( P2_R1095_U415 , P2_R1095_U167 , P2_R1095_U298 );
nand NAND2_14538 ( P2_R1095_U416 , P2_U3898 , P2_R1095_U89 );
nand NAND2_14539 ( P2_R1095_U417 , P2_U3057 , P2_R1095_U88 );
not NOT1_14540 ( P2_R1095_U418 , P2_R1095_U141 );
nand NAND2_14541 ( P2_R1095_U419 , P2_R1095_U294 , P2_R1095_U418 );
nand NAND2_14542 ( P2_R1095_U420 , P2_R1095_U141 , P2_R1095_U168 );
nand NAND2_14543 ( P2_R1095_U421 , P2_U3899 , P2_R1095_U87 );
nand NAND2_14544 ( P2_R1095_U422 , P2_U3064 , P2_R1095_U86 );
not NOT1_14545 ( P2_R1095_U423 , P2_R1095_U142 );
nand NAND2_14546 ( P2_R1095_U424 , P2_R1095_U290 , P2_R1095_U423 );
nand NAND2_14547 ( P2_R1095_U425 , P2_R1095_U142 , P2_R1095_U169 );
nand NAND2_14548 ( P2_R1095_U426 , P2_U3900 , P2_R1095_U82 );
nand NAND2_14549 ( P2_R1095_U427 , P2_U3065 , P2_R1095_U79 );
nand NAND2_14550 ( P2_R1095_U428 , P2_R1095_U427 , P2_R1095_U426 );
nand NAND2_14551 ( P2_R1095_U429 , P2_U3901 , P2_R1095_U83 );
nand NAND2_14552 ( P2_R1095_U430 , P2_U3060 , P2_R1095_U80 );
nand NAND2_14553 ( P2_R1095_U431 , P2_R1095_U316 , P2_R1095_U94 );
nand NAND2_14554 ( P2_R1095_U432 , P2_R1095_U170 , P2_R1095_U308 );
nand NAND2_14555 ( P2_R1095_U433 , P2_U3902 , P2_R1095_U84 );
nand NAND2_14556 ( P2_R1095_U434 , P2_U3074 , P2_R1095_U81 );
nand NAND2_14557 ( P2_R1095_U435 , P2_R1095_U317 , P2_R1095_U172 );
nand NAND2_14558 ( P2_R1095_U436 , P2_R1095_U280 , P2_R1095_U171 );
nand NAND2_14559 ( P2_R1095_U437 , P2_U3903 , P2_R1095_U78 );
nand NAND2_14560 ( P2_R1095_U438 , P2_U3075 , P2_R1095_U77 );
not NOT1_14561 ( P2_R1095_U439 , P2_R1095_U145 );
nand NAND2_14562 ( P2_R1095_U440 , P2_R1095_U276 , P2_R1095_U439 );
nand NAND2_14563 ( P2_R1095_U441 , P2_R1095_U145 , P2_R1095_U173 );
nand NAND2_14564 ( P2_R1095_U442 , P2_U3392 , P2_R1095_U39 );
nand NAND2_14565 ( P2_R1095_U443 , P2_U3077 , P2_R1095_U174 );
not NOT1_14566 ( P2_R1095_U444 , P2_R1095_U146 );
nand NAND2_14567 ( P2_R1095_U445 , P2_R1095_U203 , P2_R1095_U444 );
nand NAND2_14568 ( P2_R1095_U446 , P2_R1095_U146 , P2_R1095_U175 );
nand NAND2_14569 ( P2_R1095_U447 , P2_U3445 , P2_R1095_U76 );
nand NAND2_14570 ( P2_R1095_U448 , P2_U3080 , P2_R1095_U75 );
not NOT1_14571 ( P2_R1095_U449 , P2_R1095_U147 );
nand NAND2_14572 ( P2_R1095_U450 , P2_R1095_U272 , P2_R1095_U449 );
nand NAND2_14573 ( P2_R1095_U451 , P2_R1095_U147 , P2_R1095_U176 );
nand NAND2_14574 ( P2_R1095_U452 , P2_U3443 , P2_R1095_U74 );
nand NAND2_14575 ( P2_R1095_U453 , P2_U3081 , P2_R1095_U177 );
not NOT1_14576 ( P2_R1095_U454 , P2_R1095_U148 );
nand NAND2_14577 ( P2_R1095_U455 , P2_R1095_U270 , P2_R1095_U454 );
nand NAND2_14578 ( P2_R1095_U456 , P2_R1095_U148 , P2_R1095_U178 );
nand NAND2_14579 ( P2_R1095_U457 , P2_U3440 , P2_R1095_U73 );
nand NAND2_14580 ( P2_R1095_U458 , P2_U3068 , P2_R1095_U72 );
not NOT1_14581 ( P2_R1095_U459 , P2_R1095_U149 );
nand NAND2_14582 ( P2_R1095_U460 , P2_R1095_U266 , P2_R1095_U459 );
nand NAND2_14583 ( P2_R1095_U461 , P2_R1095_U149 , P2_R1095_U179 );
nand NAND2_14584 ( P2_R1095_U462 , P2_U3437 , P2_R1095_U68 );
nand NAND2_14585 ( P2_R1095_U463 , P2_U3072 , P2_R1095_U65 );
nand NAND2_14586 ( P2_R1095_U464 , P2_R1095_U463 , P2_R1095_U462 );
nand NAND2_14587 ( P2_R1095_U465 , P2_U3434 , P2_R1095_U69 );
nand NAND2_14588 ( P2_R1095_U466 , P2_U3073 , P2_R1095_U66 );
nand NAND2_14589 ( P2_R1095_U467 , P2_R1095_U327 , P2_R1095_U95 );
nand NAND2_14590 ( P2_R1095_U468 , P2_R1095_U180 , P2_R1095_U319 );
nand NAND2_14591 ( P2_R1095_U469 , P2_U3431 , P2_R1095_U70 );
nand NAND2_14592 ( P2_R1095_U470 , P2_U3078 , P2_R1095_U67 );
nand NAND2_14593 ( P2_R1095_U471 , P2_R1095_U328 , P2_R1095_U182 );
nand NAND2_14594 ( P2_R1095_U472 , P2_R1095_U256 , P2_R1095_U181 );
nand NAND2_14595 ( P2_R1095_U473 , P2_U3428 , P2_R1095_U64 );
nand NAND2_14596 ( P2_R1095_U474 , P2_U3079 , P2_R1095_U63 );
not NOT1_14597 ( P2_R1095_U475 , P2_R1095_U152 );
nand NAND2_14598 ( P2_R1095_U476 , P2_R1095_U354 , P2_R1095_U475 );
nand NAND2_14599 ( P2_R1095_U477 , P2_R1095_U152 , P2_R1095_U183 );
nand NAND2_14600 ( P2_R1095_U478 , P2_U3425 , P2_R1095_U55 );
nand NAND2_14601 ( P2_R1095_U479 , P2_U3071 , P2_R1095_U61 );
not NOT1_14602 ( P2_R1095_U480 , P2_R1095_U153 );
nand NAND2_14603 ( P2_R1095_U481 , P2_R1095_U352 , P2_R1095_U480 );
nand NAND2_14604 ( P2_R1095_U482 , P2_R1095_U153 , P2_R1095_U184 );
nand NAND2_14605 ( P2_R1095_U483 , P2_U3422 , P2_R1095_U56 );
nand NAND2_14606 ( P2_R1095_U484 , P2_U3062 , P2_R1095_U60 );
nand NAND2_14607 ( P2_R1095_U485 , P2_R1095_U484 , P2_R1095_U483 );
nand NAND2_14608 ( P2_R1095_U486 , P2_U3419 , P2_R1095_U57 );
nand NAND2_14609 ( P2_R1095_U487 , P2_U3061 , P2_R1095_U58 );
nand NAND2_14610 ( P2_R1095_U488 , P2_R1095_U96 , P2_R1095_U336 );
nand NAND2_14611 ( P2_R1095_U489 , P2_R1095_U185 , P2_R1095_U350 );
nand NAND2_14612 ( P2_R1212_U6 , P2_R1212_U176 , P2_R1212_U180 );
nand NAND2_14613 ( P2_R1212_U7 , P2_R1212_U9 , P2_R1212_U181 );
not NOT1_14614 ( P2_R1212_U8 , P2_REG2_REG_0_ );
nand NAND2_14615 ( P2_R1212_U9 , P2_REG2_REG_0_ , P2_R1212_U48 );
not NOT1_14616 ( P2_R1212_U10 , P2_REG2_REG_1_ );
not NOT1_14617 ( P2_R1212_U11 , P2_U3391 );
not NOT1_14618 ( P2_R1212_U12 , P2_REG2_REG_2_ );
not NOT1_14619 ( P2_R1212_U13 , P2_U3394 );
not NOT1_14620 ( P2_R1212_U14 , P2_REG2_REG_3_ );
not NOT1_14621 ( P2_R1212_U15 , P2_U3397 );
not NOT1_14622 ( P2_R1212_U16 , P2_REG2_REG_4_ );
not NOT1_14623 ( P2_R1212_U17 , P2_U3400 );
not NOT1_14624 ( P2_R1212_U18 , P2_REG2_REG_5_ );
not NOT1_14625 ( P2_R1212_U19 , P2_U3403 );
not NOT1_14626 ( P2_R1212_U20 , P2_REG2_REG_6_ );
not NOT1_14627 ( P2_R1212_U21 , P2_U3406 );
not NOT1_14628 ( P2_R1212_U22 , P2_REG2_REG_7_ );
not NOT1_14629 ( P2_R1212_U23 , P2_U3409 );
not NOT1_14630 ( P2_R1212_U24 , P2_REG2_REG_8_ );
not NOT1_14631 ( P2_R1212_U25 , P2_U3412 );
not NOT1_14632 ( P2_R1212_U26 , P2_REG2_REG_9_ );
not NOT1_14633 ( P2_R1212_U27 , P2_U3415 );
not NOT1_14634 ( P2_R1212_U28 , P2_REG2_REG_10_ );
not NOT1_14635 ( P2_R1212_U29 , P2_U3418 );
not NOT1_14636 ( P2_R1212_U30 , P2_REG2_REG_11_ );
not NOT1_14637 ( P2_R1212_U31 , P2_U3421 );
not NOT1_14638 ( P2_R1212_U32 , P2_REG2_REG_12_ );
not NOT1_14639 ( P2_R1212_U33 , P2_U3424 );
not NOT1_14640 ( P2_R1212_U34 , P2_REG2_REG_13_ );
not NOT1_14641 ( P2_R1212_U35 , P2_U3427 );
not NOT1_14642 ( P2_R1212_U36 , P2_REG2_REG_14_ );
not NOT1_14643 ( P2_R1212_U37 , P2_U3430 );
nand NAND2_14644 ( P2_R1212_U38 , P2_R1212_U159 , P2_R1212_U158 );
not NOT1_14645 ( P2_R1212_U39 , P2_REG2_REG_15_ );
not NOT1_14646 ( P2_R1212_U40 , P2_U3433 );
not NOT1_14647 ( P2_R1212_U41 , P2_REG2_REG_16_ );
not NOT1_14648 ( P2_R1212_U42 , P2_U3436 );
not NOT1_14649 ( P2_R1212_U43 , P2_REG2_REG_17_ );
not NOT1_14650 ( P2_R1212_U44 , P2_U3439 );
not NOT1_14651 ( P2_R1212_U45 , P2_REG2_REG_18_ );
not NOT1_14652 ( P2_R1212_U46 , P2_U3442 );
nand NAND2_14653 ( P2_R1212_U47 , P2_R1212_U171 , P2_R1212_U170 );
not NOT1_14654 ( P2_R1212_U48 , P2_U3386 );
nand NAND2_14655 ( P2_R1212_U49 , P2_R1212_U186 , P2_R1212_U185 );
nand NAND2_14656 ( P2_R1212_U50 , P2_R1212_U191 , P2_R1212_U190 );
nand NAND2_14657 ( P2_R1212_U51 , P2_R1212_U196 , P2_R1212_U195 );
nand NAND2_14658 ( P2_R1212_U52 , P2_R1212_U201 , P2_R1212_U200 );
nand NAND2_14659 ( P2_R1212_U53 , P2_R1212_U206 , P2_R1212_U205 );
nand NAND2_14660 ( P2_R1212_U54 , P2_R1212_U211 , P2_R1212_U210 );
nand NAND2_14661 ( P2_R1212_U55 , P2_R1212_U216 , P2_R1212_U215 );
nand NAND2_14662 ( P2_R1212_U56 , P2_R1212_U221 , P2_R1212_U220 );
nand NAND2_14663 ( P2_R1212_U57 , P2_R1212_U226 , P2_R1212_U225 );
nand NAND2_14664 ( P2_R1212_U58 , P2_R1212_U236 , P2_R1212_U235 );
nand NAND2_14665 ( P2_R1212_U59 , P2_R1212_U241 , P2_R1212_U240 );
nand NAND2_14666 ( P2_R1212_U60 , P2_R1212_U246 , P2_R1212_U245 );
nand NAND2_14667 ( P2_R1212_U61 , P2_R1212_U251 , P2_R1212_U250 );
nand NAND2_14668 ( P2_R1212_U62 , P2_R1212_U256 , P2_R1212_U255 );
nand NAND2_14669 ( P2_R1212_U63 , P2_R1212_U261 , P2_R1212_U260 );
nand NAND2_14670 ( P2_R1212_U64 , P2_R1212_U266 , P2_R1212_U265 );
nand NAND2_14671 ( P2_R1212_U65 , P2_R1212_U271 , P2_R1212_U270 );
nand NAND2_14672 ( P2_R1212_U66 , P2_R1212_U276 , P2_R1212_U275 );
nand NAND2_14673 ( P2_R1212_U67 , P2_R1212_U183 , P2_R1212_U182 );
nand NAND2_14674 ( P2_R1212_U68 , P2_R1212_U188 , P2_R1212_U187 );
nand NAND2_14675 ( P2_R1212_U69 , P2_R1212_U193 , P2_R1212_U192 );
nand NAND2_14676 ( P2_R1212_U70 , P2_R1212_U198 , P2_R1212_U197 );
nand NAND2_14677 ( P2_R1212_U71 , P2_R1212_U203 , P2_R1212_U202 );
nand NAND2_14678 ( P2_R1212_U72 , P2_R1212_U208 , P2_R1212_U207 );
nand NAND2_14679 ( P2_R1212_U73 , P2_R1212_U213 , P2_R1212_U212 );
nand NAND2_14680 ( P2_R1212_U74 , P2_R1212_U218 , P2_R1212_U217 );
nand NAND2_14681 ( P2_R1212_U75 , P2_R1212_U223 , P2_R1212_U222 );
and AND3_14682 ( P2_R1212_U76 , P2_R1212_U228 , P2_R1212_U227 , P2_R1212_U179 );
and AND2_14683 ( P2_R1212_U77 , P2_R1212_U175 , P2_R1212_U231 );
nand NAND2_14684 ( P2_R1212_U78 , P2_R1212_U233 , P2_R1212_U232 );
nand NAND2_14685 ( P2_R1212_U79 , P2_R1212_U238 , P2_R1212_U237 );
nand NAND2_14686 ( P2_R1212_U80 , P2_R1212_U243 , P2_R1212_U242 );
nand NAND2_14687 ( P2_R1212_U81 , P2_R1212_U248 , P2_R1212_U247 );
nand NAND2_14688 ( P2_R1212_U82 , P2_R1212_U253 , P2_R1212_U252 );
nand NAND2_14689 ( P2_R1212_U83 , P2_R1212_U258 , P2_R1212_U257 );
nand NAND2_14690 ( P2_R1212_U84 , P2_R1212_U263 , P2_R1212_U262 );
nand NAND2_14691 ( P2_R1212_U85 , P2_R1212_U268 , P2_R1212_U267 );
nand NAND2_14692 ( P2_R1212_U86 , P2_R1212_U273 , P2_R1212_U272 );
nand NAND2_14693 ( P2_R1212_U87 , P2_R1212_U135 , P2_R1212_U134 );
nand NAND2_14694 ( P2_R1212_U88 , P2_R1212_U131 , P2_R1212_U130 );
nand NAND2_14695 ( P2_R1212_U89 , P2_R1212_U127 , P2_R1212_U126 );
nand NAND2_14696 ( P2_R1212_U90 , P2_R1212_U123 , P2_R1212_U122 );
nand NAND2_14697 ( P2_R1212_U91 , P2_R1212_U119 , P2_R1212_U118 );
nand NAND2_14698 ( P2_R1212_U92 , P2_R1212_U115 , P2_R1212_U114 );
nand NAND2_14699 ( P2_R1212_U93 , P2_R1212_U111 , P2_R1212_U110 );
nand NAND2_14700 ( P2_R1212_U94 , P2_R1212_U107 , P2_R1212_U106 );
not NOT1_14701 ( P2_R1212_U95 , P2_REG2_REG_19_ );
not NOT1_14702 ( P2_R1212_U96 , P2_U3379 );
nand NAND2_14703 ( P2_R1212_U97 , P2_R1212_U167 , P2_R1212_U166 );
nand NAND2_14704 ( P2_R1212_U98 , P2_R1212_U163 , P2_R1212_U162 );
nand NAND2_14705 ( P2_R1212_U99 , P2_R1212_U155 , P2_R1212_U154 );
nand NAND2_14706 ( P2_R1212_U100 , P2_R1212_U151 , P2_R1212_U150 );
nand NAND2_14707 ( P2_R1212_U101 , P2_R1212_U147 , P2_R1212_U146 );
nand NAND2_14708 ( P2_R1212_U102 , P2_R1212_U143 , P2_R1212_U142 );
nand NAND2_14709 ( P2_R1212_U103 , P2_R1212_U139 , P2_R1212_U138 );
not NOT1_14710 ( P2_R1212_U104 , P2_R1212_U9 );
nand NAND2_14711 ( P2_R1212_U105 , P2_REG2_REG_1_ , P2_R1212_U104 );
nand NAND2_14712 ( P2_R1212_U106 , P2_U3391 , P2_R1212_U105 );
nand NAND2_14713 ( P2_R1212_U107 , P2_R1212_U9 , P2_R1212_U10 );
not NOT1_14714 ( P2_R1212_U108 , P2_R1212_U94 );
nand NAND2_14715 ( P2_R1212_U109 , P2_REG2_REG_2_ , P2_R1212_U13 );
nand NAND2_14716 ( P2_R1212_U110 , P2_R1212_U109 , P2_R1212_U94 );
nand NAND2_14717 ( P2_R1212_U111 , P2_U3394 , P2_R1212_U12 );
not NOT1_14718 ( P2_R1212_U112 , P2_R1212_U93 );
nand NAND2_14719 ( P2_R1212_U113 , P2_REG2_REG_3_ , P2_R1212_U15 );
nand NAND2_14720 ( P2_R1212_U114 , P2_R1212_U113 , P2_R1212_U93 );
nand NAND2_14721 ( P2_R1212_U115 , P2_U3397 , P2_R1212_U14 );
not NOT1_14722 ( P2_R1212_U116 , P2_R1212_U92 );
nand NAND2_14723 ( P2_R1212_U117 , P2_REG2_REG_4_ , P2_R1212_U17 );
nand NAND2_14724 ( P2_R1212_U118 , P2_R1212_U117 , P2_R1212_U92 );
nand NAND2_14725 ( P2_R1212_U119 , P2_U3400 , P2_R1212_U16 );
not NOT1_14726 ( P2_R1212_U120 , P2_R1212_U91 );
nand NAND2_14727 ( P2_R1212_U121 , P2_REG2_REG_5_ , P2_R1212_U19 );
nand NAND2_14728 ( P2_R1212_U122 , P2_R1212_U121 , P2_R1212_U91 );
nand NAND2_14729 ( P2_R1212_U123 , P2_U3403 , P2_R1212_U18 );
not NOT1_14730 ( P2_R1212_U124 , P2_R1212_U90 );
nand NAND2_14731 ( P2_R1212_U125 , P2_REG2_REG_6_ , P2_R1212_U21 );
nand NAND2_14732 ( P2_R1212_U126 , P2_R1212_U125 , P2_R1212_U90 );
nand NAND2_14733 ( P2_R1212_U127 , P2_U3406 , P2_R1212_U20 );
not NOT1_14734 ( P2_R1212_U128 , P2_R1212_U89 );
nand NAND2_14735 ( P2_R1212_U129 , P2_REG2_REG_7_ , P2_R1212_U23 );
nand NAND2_14736 ( P2_R1212_U130 , P2_R1212_U129 , P2_R1212_U89 );
nand NAND2_14737 ( P2_R1212_U131 , P2_U3409 , P2_R1212_U22 );
not NOT1_14738 ( P2_R1212_U132 , P2_R1212_U88 );
nand NAND2_14739 ( P2_R1212_U133 , P2_REG2_REG_8_ , P2_R1212_U25 );
nand NAND2_14740 ( P2_R1212_U134 , P2_R1212_U133 , P2_R1212_U88 );
nand NAND2_14741 ( P2_R1212_U135 , P2_U3412 , P2_R1212_U24 );
not NOT1_14742 ( P2_R1212_U136 , P2_R1212_U87 );
nand NAND2_14743 ( P2_R1212_U137 , P2_REG2_REG_9_ , P2_R1212_U27 );
nand NAND2_14744 ( P2_R1212_U138 , P2_R1212_U137 , P2_R1212_U87 );
nand NAND2_14745 ( P2_R1212_U139 , P2_U3415 , P2_R1212_U26 );
not NOT1_14746 ( P2_R1212_U140 , P2_R1212_U103 );
nand NAND2_14747 ( P2_R1212_U141 , P2_REG2_REG_10_ , P2_R1212_U29 );
nand NAND2_14748 ( P2_R1212_U142 , P2_R1212_U141 , P2_R1212_U103 );
nand NAND2_14749 ( P2_R1212_U143 , P2_U3418 , P2_R1212_U28 );
not NOT1_14750 ( P2_R1212_U144 , P2_R1212_U102 );
nand NAND2_14751 ( P2_R1212_U145 , P2_REG2_REG_11_ , P2_R1212_U31 );
nand NAND2_14752 ( P2_R1212_U146 , P2_R1212_U145 , P2_R1212_U102 );
nand NAND2_14753 ( P2_R1212_U147 , P2_U3421 , P2_R1212_U30 );
not NOT1_14754 ( P2_R1212_U148 , P2_R1212_U101 );
nand NAND2_14755 ( P2_R1212_U149 , P2_REG2_REG_12_ , P2_R1212_U33 );
nand NAND2_14756 ( P2_R1212_U150 , P2_R1212_U149 , P2_R1212_U101 );
nand NAND2_14757 ( P2_R1212_U151 , P2_U3424 , P2_R1212_U32 );
not NOT1_14758 ( P2_R1212_U152 , P2_R1212_U100 );
nand NAND2_14759 ( P2_R1212_U153 , P2_REG2_REG_13_ , P2_R1212_U35 );
nand NAND2_14760 ( P2_R1212_U154 , P2_R1212_U153 , P2_R1212_U100 );
nand NAND2_14761 ( P2_R1212_U155 , P2_U3427 , P2_R1212_U34 );
not NOT1_14762 ( P2_R1212_U156 , P2_R1212_U99 );
nand NAND2_14763 ( P2_R1212_U157 , P2_REG2_REG_14_ , P2_R1212_U37 );
nand NAND2_14764 ( P2_R1212_U158 , P2_R1212_U157 , P2_R1212_U99 );
nand NAND2_14765 ( P2_R1212_U159 , P2_U3430 , P2_R1212_U36 );
not NOT1_14766 ( P2_R1212_U160 , P2_R1212_U38 );
nand NAND2_14767 ( P2_R1212_U161 , P2_REG2_REG_15_ , P2_R1212_U160 );
nand NAND2_14768 ( P2_R1212_U162 , P2_U3433 , P2_R1212_U161 );
nand NAND2_14769 ( P2_R1212_U163 , P2_R1212_U38 , P2_R1212_U39 );
not NOT1_14770 ( P2_R1212_U164 , P2_R1212_U98 );
nand NAND2_14771 ( P2_R1212_U165 , P2_REG2_REG_16_ , P2_R1212_U42 );
nand NAND2_14772 ( P2_R1212_U166 , P2_R1212_U165 , P2_R1212_U98 );
nand NAND2_14773 ( P2_R1212_U167 , P2_U3436 , P2_R1212_U41 );
not NOT1_14774 ( P2_R1212_U168 , P2_R1212_U97 );
nand NAND2_14775 ( P2_R1212_U169 , P2_REG2_REG_17_ , P2_R1212_U44 );
nand NAND2_14776 ( P2_R1212_U170 , P2_R1212_U169 , P2_R1212_U97 );
nand NAND2_14777 ( P2_R1212_U171 , P2_U3439 , P2_R1212_U43 );
not NOT1_14778 ( P2_R1212_U172 , P2_R1212_U47 );
nand NAND2_14779 ( P2_R1212_U173 , P2_U3442 , P2_R1212_U45 );
nand NAND2_14780 ( P2_R1212_U174 , P2_R1212_U172 , P2_R1212_U173 );
nand NAND2_14781 ( P2_R1212_U175 , P2_REG2_REG_18_ , P2_R1212_U46 );
nand NAND2_14782 ( P2_R1212_U176 , P2_R1212_U77 , P2_R1212_U174 );
nand NAND2_14783 ( P2_R1212_U177 , P2_REG2_REG_18_ , P2_R1212_U46 );
nand NAND2_14784 ( P2_R1212_U178 , P2_R1212_U177 , P2_R1212_U47 );
nand NAND2_14785 ( P2_R1212_U179 , P2_U3442 , P2_R1212_U45 );
nand NAND2_14786 ( P2_R1212_U180 , P2_R1212_U76 , P2_R1212_U178 );
nand NAND2_14787 ( P2_R1212_U181 , P2_U3386 , P2_R1212_U8 );
nand NAND2_14788 ( P2_R1212_U182 , P2_REG2_REG_9_ , P2_R1212_U27 );
nand NAND2_14789 ( P2_R1212_U183 , P2_U3415 , P2_R1212_U26 );
not NOT1_14790 ( P2_R1212_U184 , P2_R1212_U67 );
nand NAND2_14791 ( P2_R1212_U185 , P2_R1212_U136 , P2_R1212_U184 );
nand NAND2_14792 ( P2_R1212_U186 , P2_R1212_U67 , P2_R1212_U87 );
nand NAND2_14793 ( P2_R1212_U187 , P2_REG2_REG_8_ , P2_R1212_U25 );
nand NAND2_14794 ( P2_R1212_U188 , P2_U3412 , P2_R1212_U24 );
not NOT1_14795 ( P2_R1212_U189 , P2_R1212_U68 );
nand NAND2_14796 ( P2_R1212_U190 , P2_R1212_U132 , P2_R1212_U189 );
nand NAND2_14797 ( P2_R1212_U191 , P2_R1212_U68 , P2_R1212_U88 );
nand NAND2_14798 ( P2_R1212_U192 , P2_REG2_REG_7_ , P2_R1212_U23 );
nand NAND2_14799 ( P2_R1212_U193 , P2_U3409 , P2_R1212_U22 );
not NOT1_14800 ( P2_R1212_U194 , P2_R1212_U69 );
nand NAND2_14801 ( P2_R1212_U195 , P2_R1212_U128 , P2_R1212_U194 );
nand NAND2_14802 ( P2_R1212_U196 , P2_R1212_U69 , P2_R1212_U89 );
nand NAND2_14803 ( P2_R1212_U197 , P2_REG2_REG_6_ , P2_R1212_U21 );
nand NAND2_14804 ( P2_R1212_U198 , P2_U3406 , P2_R1212_U20 );
not NOT1_14805 ( P2_R1212_U199 , P2_R1212_U70 );
nand NAND2_14806 ( P2_R1212_U200 , P2_R1212_U124 , P2_R1212_U199 );
nand NAND2_14807 ( P2_R1212_U201 , P2_R1212_U70 , P2_R1212_U90 );
nand NAND2_14808 ( P2_R1212_U202 , P2_REG2_REG_5_ , P2_R1212_U19 );
nand NAND2_14809 ( P2_R1212_U203 , P2_U3403 , P2_R1212_U18 );
not NOT1_14810 ( P2_R1212_U204 , P2_R1212_U71 );
nand NAND2_14811 ( P2_R1212_U205 , P2_R1212_U120 , P2_R1212_U204 );
nand NAND2_14812 ( P2_R1212_U206 , P2_R1212_U71 , P2_R1212_U91 );
nand NAND2_14813 ( P2_R1212_U207 , P2_REG2_REG_4_ , P2_R1212_U17 );
nand NAND2_14814 ( P2_R1212_U208 , P2_U3400 , P2_R1212_U16 );
not NOT1_14815 ( P2_R1212_U209 , P2_R1212_U72 );
nand NAND2_14816 ( P2_R1212_U210 , P2_R1212_U116 , P2_R1212_U209 );
nand NAND2_14817 ( P2_R1212_U211 , P2_R1212_U72 , P2_R1212_U92 );
nand NAND2_14818 ( P2_R1212_U212 , P2_REG2_REG_3_ , P2_R1212_U15 );
nand NAND2_14819 ( P2_R1212_U213 , P2_U3397 , P2_R1212_U14 );
not NOT1_14820 ( P2_R1212_U214 , P2_R1212_U73 );
nand NAND2_14821 ( P2_R1212_U215 , P2_R1212_U112 , P2_R1212_U214 );
nand NAND2_14822 ( P2_R1212_U216 , P2_R1212_U73 , P2_R1212_U93 );
nand NAND2_14823 ( P2_R1212_U217 , P2_REG2_REG_2_ , P2_R1212_U13 );
nand NAND2_14824 ( P2_R1212_U218 , P2_U3394 , P2_R1212_U12 );
not NOT1_14825 ( P2_R1212_U219 , P2_R1212_U74 );
nand NAND2_14826 ( P2_R1212_U220 , P2_R1212_U108 , P2_R1212_U219 );
nand NAND2_14827 ( P2_R1212_U221 , P2_R1212_U74 , P2_R1212_U94 );
nand NAND2_14828 ( P2_R1212_U222 , P2_R1212_U104 , P2_R1212_U10 );
nand NAND2_14829 ( P2_R1212_U223 , P2_REG2_REG_1_ , P2_R1212_U9 );
not NOT1_14830 ( P2_R1212_U224 , P2_R1212_U75 );
nand NAND2_14831 ( P2_R1212_U225 , P2_R1212_U224 , P2_U3391 );
nand NAND2_14832 ( P2_R1212_U226 , P2_R1212_U75 , P2_R1212_U11 );
nand NAND2_14833 ( P2_R1212_U227 , P2_REG2_REG_19_ , P2_R1212_U96 );
nand NAND2_14834 ( P2_R1212_U228 , P2_U3379 , P2_R1212_U95 );
nand NAND2_14835 ( P2_R1212_U229 , P2_REG2_REG_19_ , P2_R1212_U96 );
nand NAND2_14836 ( P2_R1212_U230 , P2_U3379 , P2_R1212_U95 );
nand NAND2_14837 ( P2_R1212_U231 , P2_R1212_U230 , P2_R1212_U229 );
nand NAND2_14838 ( P2_R1212_U232 , P2_REG2_REG_18_ , P2_R1212_U46 );
nand NAND2_14839 ( P2_R1212_U233 , P2_U3442 , P2_R1212_U45 );
not NOT1_14840 ( P2_R1212_U234 , P2_R1212_U78 );
nand NAND2_14841 ( P2_R1212_U235 , P2_R1212_U234 , P2_R1212_U172 );
nand NAND2_14842 ( P2_R1212_U236 , P2_R1212_U78 , P2_R1212_U47 );
nand NAND2_14843 ( P2_R1212_U237 , P2_REG2_REG_17_ , P2_R1212_U44 );
nand NAND2_14844 ( P2_R1212_U238 , P2_U3439 , P2_R1212_U43 );
not NOT1_14845 ( P2_R1212_U239 , P2_R1212_U79 );
nand NAND2_14846 ( P2_R1212_U240 , P2_R1212_U168 , P2_R1212_U239 );
nand NAND2_14847 ( P2_R1212_U241 , P2_R1212_U79 , P2_R1212_U97 );
nand NAND2_14848 ( P2_R1212_U242 , P2_REG2_REG_16_ , P2_R1212_U42 );
nand NAND2_14849 ( P2_R1212_U243 , P2_U3436 , P2_R1212_U41 );
not NOT1_14850 ( P2_R1212_U244 , P2_R1212_U80 );
nand NAND2_14851 ( P2_R1212_U245 , P2_R1212_U164 , P2_R1212_U244 );
nand NAND2_14852 ( P2_R1212_U246 , P2_R1212_U80 , P2_R1212_U98 );
nand NAND2_14853 ( P2_R1212_U247 , P2_U3433 , P2_R1212_U39 );
nand NAND2_14854 ( P2_R1212_U248 , P2_REG2_REG_15_ , P2_R1212_U40 );
not NOT1_14855 ( P2_R1212_U249 , P2_R1212_U81 );
nand NAND2_14856 ( P2_R1212_U250 , P2_R1212_U249 , P2_R1212_U160 );
nand NAND2_14857 ( P2_R1212_U251 , P2_R1212_U81 , P2_R1212_U38 );
nand NAND2_14858 ( P2_R1212_U252 , P2_REG2_REG_14_ , P2_R1212_U37 );
nand NAND2_14859 ( P2_R1212_U253 , P2_U3430 , P2_R1212_U36 );
not NOT1_14860 ( P2_R1212_U254 , P2_R1212_U82 );
nand NAND2_14861 ( P2_R1212_U255 , P2_R1212_U156 , P2_R1212_U254 );
nand NAND2_14862 ( P2_R1212_U256 , P2_R1212_U82 , P2_R1212_U99 );
nand NAND2_14863 ( P2_R1212_U257 , P2_REG2_REG_13_ , P2_R1212_U35 );
nand NAND2_14864 ( P2_R1212_U258 , P2_U3427 , P2_R1212_U34 );
not NOT1_14865 ( P2_R1212_U259 , P2_R1212_U83 );
nand NAND2_14866 ( P2_R1212_U260 , P2_R1212_U152 , P2_R1212_U259 );
nand NAND2_14867 ( P2_R1212_U261 , P2_R1212_U83 , P2_R1212_U100 );
nand NAND2_14868 ( P2_R1212_U262 , P2_REG2_REG_12_ , P2_R1212_U33 );
nand NAND2_14869 ( P2_R1212_U263 , P2_U3424 , P2_R1212_U32 );
not NOT1_14870 ( P2_R1212_U264 , P2_R1212_U84 );
nand NAND2_14871 ( P2_R1212_U265 , P2_R1212_U148 , P2_R1212_U264 );
nand NAND2_14872 ( P2_R1212_U266 , P2_R1212_U84 , P2_R1212_U101 );
nand NAND2_14873 ( P2_R1212_U267 , P2_REG2_REG_11_ , P2_R1212_U31 );
nand NAND2_14874 ( P2_R1212_U268 , P2_U3421 , P2_R1212_U30 );
not NOT1_14875 ( P2_R1212_U269 , P2_R1212_U85 );
nand NAND2_14876 ( P2_R1212_U270 , P2_R1212_U144 , P2_R1212_U269 );
nand NAND2_14877 ( P2_R1212_U271 , P2_R1212_U85 , P2_R1212_U102 );
nand NAND2_14878 ( P2_R1212_U272 , P2_REG2_REG_10_ , P2_R1212_U29 );
nand NAND2_14879 ( P2_R1212_U273 , P2_U3418 , P2_R1212_U28 );
not NOT1_14880 ( P2_R1212_U274 , P2_R1212_U86 );
nand NAND2_14881 ( P2_R1212_U275 , P2_R1212_U140 , P2_R1212_U274 );
nand NAND2_14882 ( P2_R1212_U276 , P2_R1212_U86 , P2_R1212_U103 );
nand NAND2_14883 ( P2_R1209_U6 , P2_R1209_U176 , P2_R1209_U180 );
nand NAND2_14884 ( P2_R1209_U7 , P2_R1209_U9 , P2_R1209_U181 );
not NOT1_14885 ( P2_R1209_U8 , P2_REG1_REG_0_ );
nand NAND2_14886 ( P2_R1209_U9 , P2_REG1_REG_0_ , P2_R1209_U48 );
not NOT1_14887 ( P2_R1209_U10 , P2_REG1_REG_1_ );
not NOT1_14888 ( P2_R1209_U11 , P2_U3391 );
not NOT1_14889 ( P2_R1209_U12 , P2_REG1_REG_2_ );
not NOT1_14890 ( P2_R1209_U13 , P2_U3394 );
not NOT1_14891 ( P2_R1209_U14 , P2_REG1_REG_3_ );
not NOT1_14892 ( P2_R1209_U15 , P2_U3397 );
not NOT1_14893 ( P2_R1209_U16 , P2_REG1_REG_4_ );
not NOT1_14894 ( P2_R1209_U17 , P2_U3400 );
not NOT1_14895 ( P2_R1209_U18 , P2_REG1_REG_5_ );
not NOT1_14896 ( P2_R1209_U19 , P2_U3403 );
not NOT1_14897 ( P2_R1209_U20 , P2_REG1_REG_6_ );
not NOT1_14898 ( P2_R1209_U21 , P2_U3406 );
not NOT1_14899 ( P2_R1209_U22 , P2_REG1_REG_7_ );
not NOT1_14900 ( P2_R1209_U23 , P2_U3409 );
not NOT1_14901 ( P2_R1209_U24 , P2_REG1_REG_8_ );
not NOT1_14902 ( P2_R1209_U25 , P2_U3412 );
not NOT1_14903 ( P2_R1209_U26 , P2_REG1_REG_9_ );
not NOT1_14904 ( P2_R1209_U27 , P2_U3415 );
not NOT1_14905 ( P2_R1209_U28 , P2_REG1_REG_10_ );
not NOT1_14906 ( P2_R1209_U29 , P2_U3418 );
not NOT1_14907 ( P2_R1209_U30 , P2_REG1_REG_11_ );
not NOT1_14908 ( P2_R1209_U31 , P2_U3421 );
not NOT1_14909 ( P2_R1209_U32 , P2_REG1_REG_12_ );
not NOT1_14910 ( P2_R1209_U33 , P2_U3424 );
not NOT1_14911 ( P2_R1209_U34 , P2_REG1_REG_13_ );
not NOT1_14912 ( P2_R1209_U35 , P2_U3427 );
not NOT1_14913 ( P2_R1209_U36 , P2_REG1_REG_14_ );
not NOT1_14914 ( P2_R1209_U37 , P2_U3430 );
nand NAND2_14915 ( P2_R1209_U38 , P2_R1209_U159 , P2_R1209_U158 );
not NOT1_14916 ( P2_R1209_U39 , P2_REG1_REG_15_ );
not NOT1_14917 ( P2_R1209_U40 , P2_U3433 );
not NOT1_14918 ( P2_R1209_U41 , P2_REG1_REG_16_ );
not NOT1_14919 ( P2_R1209_U42 , P2_U3436 );
not NOT1_14920 ( P2_R1209_U43 , P2_REG1_REG_17_ );
not NOT1_14921 ( P2_R1209_U44 , P2_U3439 );
not NOT1_14922 ( P2_R1209_U45 , P2_REG1_REG_18_ );
not NOT1_14923 ( P2_R1209_U46 , P2_U3442 );
nand NAND2_14924 ( P2_R1209_U47 , P2_R1209_U171 , P2_R1209_U170 );
not NOT1_14925 ( P2_R1209_U48 , P2_U3386 );
nand NAND2_14926 ( P2_R1209_U49 , P2_R1209_U186 , P2_R1209_U185 );
nand NAND2_14927 ( P2_R1209_U50 , P2_R1209_U191 , P2_R1209_U190 );
nand NAND2_14928 ( P2_R1209_U51 , P2_R1209_U196 , P2_R1209_U195 );
nand NAND2_14929 ( P2_R1209_U52 , P2_R1209_U201 , P2_R1209_U200 );
nand NAND2_14930 ( P2_R1209_U53 , P2_R1209_U206 , P2_R1209_U205 );
nand NAND2_14931 ( P2_R1209_U54 , P2_R1209_U211 , P2_R1209_U210 );
nand NAND2_14932 ( P2_R1209_U55 , P2_R1209_U216 , P2_R1209_U215 );
nand NAND2_14933 ( P2_R1209_U56 , P2_R1209_U221 , P2_R1209_U220 );
nand NAND2_14934 ( P2_R1209_U57 , P2_R1209_U226 , P2_R1209_U225 );
nand NAND2_14935 ( P2_R1209_U58 , P2_R1209_U236 , P2_R1209_U235 );
nand NAND2_14936 ( P2_R1209_U59 , P2_R1209_U241 , P2_R1209_U240 );
nand NAND2_14937 ( P2_R1209_U60 , P2_R1209_U246 , P2_R1209_U245 );
nand NAND2_14938 ( P2_R1209_U61 , P2_R1209_U251 , P2_R1209_U250 );
nand NAND2_14939 ( P2_R1209_U62 , P2_R1209_U256 , P2_R1209_U255 );
nand NAND2_14940 ( P2_R1209_U63 , P2_R1209_U261 , P2_R1209_U260 );
nand NAND2_14941 ( P2_R1209_U64 , P2_R1209_U266 , P2_R1209_U265 );
nand NAND2_14942 ( P2_R1209_U65 , P2_R1209_U271 , P2_R1209_U270 );
nand NAND2_14943 ( P2_R1209_U66 , P2_R1209_U276 , P2_R1209_U275 );
nand NAND2_14944 ( P2_R1209_U67 , P2_R1209_U183 , P2_R1209_U182 );
nand NAND2_14945 ( P2_R1209_U68 , P2_R1209_U188 , P2_R1209_U187 );
nand NAND2_14946 ( P2_R1209_U69 , P2_R1209_U193 , P2_R1209_U192 );
nand NAND2_14947 ( P2_R1209_U70 , P2_R1209_U198 , P2_R1209_U197 );
nand NAND2_14948 ( P2_R1209_U71 , P2_R1209_U203 , P2_R1209_U202 );
nand NAND2_14949 ( P2_R1209_U72 , P2_R1209_U208 , P2_R1209_U207 );
nand NAND2_14950 ( P2_R1209_U73 , P2_R1209_U213 , P2_R1209_U212 );
nand NAND2_14951 ( P2_R1209_U74 , P2_R1209_U218 , P2_R1209_U217 );
nand NAND2_14952 ( P2_R1209_U75 , P2_R1209_U223 , P2_R1209_U222 );
and AND3_14953 ( P2_R1209_U76 , P2_R1209_U228 , P2_R1209_U227 , P2_R1209_U179 );
and AND2_14954 ( P2_R1209_U77 , P2_R1209_U175 , P2_R1209_U231 );
nand NAND2_14955 ( P2_R1209_U78 , P2_R1209_U233 , P2_R1209_U232 );
nand NAND2_14956 ( P2_R1209_U79 , P2_R1209_U238 , P2_R1209_U237 );
nand NAND2_14957 ( P2_R1209_U80 , P2_R1209_U243 , P2_R1209_U242 );
nand NAND2_14958 ( P2_R1209_U81 , P2_R1209_U248 , P2_R1209_U247 );
nand NAND2_14959 ( P2_R1209_U82 , P2_R1209_U253 , P2_R1209_U252 );
nand NAND2_14960 ( P2_R1209_U83 , P2_R1209_U258 , P2_R1209_U257 );
nand NAND2_14961 ( P2_R1209_U84 , P2_R1209_U263 , P2_R1209_U262 );
nand NAND2_14962 ( P2_R1209_U85 , P2_R1209_U268 , P2_R1209_U267 );
nand NAND2_14963 ( P2_R1209_U86 , P2_R1209_U273 , P2_R1209_U272 );
nand NAND2_14964 ( P2_R1209_U87 , P2_R1209_U135 , P2_R1209_U134 );
nand NAND2_14965 ( P2_R1209_U88 , P2_R1209_U131 , P2_R1209_U130 );
nand NAND2_14966 ( P2_R1209_U89 , P2_R1209_U127 , P2_R1209_U126 );
nand NAND2_14967 ( P2_R1209_U90 , P2_R1209_U123 , P2_R1209_U122 );
nand NAND2_14968 ( P2_R1209_U91 , P2_R1209_U119 , P2_R1209_U118 );
nand NAND2_14969 ( P2_R1209_U92 , P2_R1209_U115 , P2_R1209_U114 );
nand NAND2_14970 ( P2_R1209_U93 , P2_R1209_U111 , P2_R1209_U110 );
nand NAND2_14971 ( P2_R1209_U94 , P2_R1209_U107 , P2_R1209_U106 );
not NOT1_14972 ( P2_R1209_U95 , P2_REG1_REG_19_ );
not NOT1_14973 ( P2_R1209_U96 , P2_U3379 );
nand NAND2_14974 ( P2_R1209_U97 , P2_R1209_U167 , P2_R1209_U166 );
nand NAND2_14975 ( P2_R1209_U98 , P2_R1209_U163 , P2_R1209_U162 );
nand NAND2_14976 ( P2_R1209_U99 , P2_R1209_U155 , P2_R1209_U154 );
nand NAND2_14977 ( P2_R1209_U100 , P2_R1209_U151 , P2_R1209_U150 );
nand NAND2_14978 ( P2_R1209_U101 , P2_R1209_U147 , P2_R1209_U146 );
nand NAND2_14979 ( P2_R1209_U102 , P2_R1209_U143 , P2_R1209_U142 );
nand NAND2_14980 ( P2_R1209_U103 , P2_R1209_U139 , P2_R1209_U138 );
not NOT1_14981 ( P2_R1209_U104 , P2_R1209_U9 );
nand NAND2_14982 ( P2_R1209_U105 , P2_REG1_REG_1_ , P2_R1209_U104 );
nand NAND2_14983 ( P2_R1209_U106 , P2_U3391 , P2_R1209_U105 );
nand NAND2_14984 ( P2_R1209_U107 , P2_R1209_U9 , P2_R1209_U10 );
not NOT1_14985 ( P2_R1209_U108 , P2_R1209_U94 );
nand NAND2_14986 ( P2_R1209_U109 , P2_REG1_REG_2_ , P2_R1209_U13 );
nand NAND2_14987 ( P2_R1209_U110 , P2_R1209_U109 , P2_R1209_U94 );
nand NAND2_14988 ( P2_R1209_U111 , P2_U3394 , P2_R1209_U12 );
not NOT1_14989 ( P2_R1209_U112 , P2_R1209_U93 );
nand NAND2_14990 ( P2_R1209_U113 , P2_REG1_REG_3_ , P2_R1209_U15 );
nand NAND2_14991 ( P2_R1209_U114 , P2_R1209_U113 , P2_R1209_U93 );
nand NAND2_14992 ( P2_R1209_U115 , P2_U3397 , P2_R1209_U14 );
not NOT1_14993 ( P2_R1209_U116 , P2_R1209_U92 );
nand NAND2_14994 ( P2_R1209_U117 , P2_REG1_REG_4_ , P2_R1209_U17 );
nand NAND2_14995 ( P2_R1209_U118 , P2_R1209_U117 , P2_R1209_U92 );
nand NAND2_14996 ( P2_R1209_U119 , P2_U3400 , P2_R1209_U16 );
not NOT1_14997 ( P2_R1209_U120 , P2_R1209_U91 );
nand NAND2_14998 ( P2_R1209_U121 , P2_REG1_REG_5_ , P2_R1209_U19 );
nand NAND2_14999 ( P2_R1209_U122 , P2_R1209_U121 , P2_R1209_U91 );
nand NAND2_15000 ( P2_R1209_U123 , P2_U3403 , P2_R1209_U18 );
not NOT1_15001 ( P2_R1209_U124 , P2_R1209_U90 );
nand NAND2_15002 ( P2_R1209_U125 , P2_REG1_REG_6_ , P2_R1209_U21 );
nand NAND2_15003 ( P2_R1209_U126 , P2_R1209_U125 , P2_R1209_U90 );
nand NAND2_15004 ( P2_R1209_U127 , P2_U3406 , P2_R1209_U20 );
not NOT1_15005 ( P2_R1209_U128 , P2_R1209_U89 );
nand NAND2_15006 ( P2_R1209_U129 , P2_REG1_REG_7_ , P2_R1209_U23 );
nand NAND2_15007 ( P2_R1209_U130 , P2_R1209_U129 , P2_R1209_U89 );
nand NAND2_15008 ( P2_R1209_U131 , P2_U3409 , P2_R1209_U22 );
not NOT1_15009 ( P2_R1209_U132 , P2_R1209_U88 );
nand NAND2_15010 ( P2_R1209_U133 , P2_REG1_REG_8_ , P2_R1209_U25 );
nand NAND2_15011 ( P2_R1209_U134 , P2_R1209_U133 , P2_R1209_U88 );
nand NAND2_15012 ( P2_R1209_U135 , P2_U3412 , P2_R1209_U24 );
not NOT1_15013 ( P2_R1209_U136 , P2_R1209_U87 );
nand NAND2_15014 ( P2_R1209_U137 , P2_REG1_REG_9_ , P2_R1209_U27 );
nand NAND2_15015 ( P2_R1209_U138 , P2_R1209_U137 , P2_R1209_U87 );
nand NAND2_15016 ( P2_R1209_U139 , P2_U3415 , P2_R1209_U26 );
not NOT1_15017 ( P2_R1209_U140 , P2_R1209_U103 );
nand NAND2_15018 ( P2_R1209_U141 , P2_REG1_REG_10_ , P2_R1209_U29 );
nand NAND2_15019 ( P2_R1209_U142 , P2_R1209_U141 , P2_R1209_U103 );
nand NAND2_15020 ( P2_R1209_U143 , P2_U3418 , P2_R1209_U28 );
not NOT1_15021 ( P2_R1209_U144 , P2_R1209_U102 );
nand NAND2_15022 ( P2_R1209_U145 , P2_REG1_REG_11_ , P2_R1209_U31 );
nand NAND2_15023 ( P2_R1209_U146 , P2_R1209_U145 , P2_R1209_U102 );
nand NAND2_15024 ( P2_R1209_U147 , P2_U3421 , P2_R1209_U30 );
not NOT1_15025 ( P2_R1209_U148 , P2_R1209_U101 );
nand NAND2_15026 ( P2_R1209_U149 , P2_REG1_REG_12_ , P2_R1209_U33 );
nand NAND2_15027 ( P2_R1209_U150 , P2_R1209_U149 , P2_R1209_U101 );
nand NAND2_15028 ( P2_R1209_U151 , P2_U3424 , P2_R1209_U32 );
not NOT1_15029 ( P2_R1209_U152 , P2_R1209_U100 );
nand NAND2_15030 ( P2_R1209_U153 , P2_REG1_REG_13_ , P2_R1209_U35 );
nand NAND2_15031 ( P2_R1209_U154 , P2_R1209_U153 , P2_R1209_U100 );
nand NAND2_15032 ( P2_R1209_U155 , P2_U3427 , P2_R1209_U34 );
not NOT1_15033 ( P2_R1209_U156 , P2_R1209_U99 );
nand NAND2_15034 ( P2_R1209_U157 , P2_REG1_REG_14_ , P2_R1209_U37 );
nand NAND2_15035 ( P2_R1209_U158 , P2_R1209_U157 , P2_R1209_U99 );
nand NAND2_15036 ( P2_R1209_U159 , P2_U3430 , P2_R1209_U36 );
not NOT1_15037 ( P2_R1209_U160 , P2_R1209_U38 );
nand NAND2_15038 ( P2_R1209_U161 , P2_REG1_REG_15_ , P2_R1209_U160 );
nand NAND2_15039 ( P2_R1209_U162 , P2_U3433 , P2_R1209_U161 );
nand NAND2_15040 ( P2_R1209_U163 , P2_R1209_U38 , P2_R1209_U39 );
not NOT1_15041 ( P2_R1209_U164 , P2_R1209_U98 );
nand NAND2_15042 ( P2_R1209_U165 , P2_REG1_REG_16_ , P2_R1209_U42 );
nand NAND2_15043 ( P2_R1209_U166 , P2_R1209_U165 , P2_R1209_U98 );
nand NAND2_15044 ( P2_R1209_U167 , P2_U3436 , P2_R1209_U41 );
not NOT1_15045 ( P2_R1209_U168 , P2_R1209_U97 );
nand NAND2_15046 ( P2_R1209_U169 , P2_REG1_REG_17_ , P2_R1209_U44 );
nand NAND2_15047 ( P2_R1209_U170 , P2_R1209_U169 , P2_R1209_U97 );
nand NAND2_15048 ( P2_R1209_U171 , P2_U3439 , P2_R1209_U43 );
not NOT1_15049 ( P2_R1209_U172 , P2_R1209_U47 );
nand NAND2_15050 ( P2_R1209_U173 , P2_U3442 , P2_R1209_U45 );
nand NAND2_15051 ( P2_R1209_U174 , P2_R1209_U172 , P2_R1209_U173 );
nand NAND2_15052 ( P2_R1209_U175 , P2_REG1_REG_18_ , P2_R1209_U46 );
nand NAND2_15053 ( P2_R1209_U176 , P2_R1209_U77 , P2_R1209_U174 );
nand NAND2_15054 ( P2_R1209_U177 , P2_REG1_REG_18_ , P2_R1209_U46 );
nand NAND2_15055 ( P2_R1209_U178 , P2_R1209_U177 , P2_R1209_U47 );
nand NAND2_15056 ( P2_R1209_U179 , P2_U3442 , P2_R1209_U45 );
nand NAND2_15057 ( P2_R1209_U180 , P2_R1209_U76 , P2_R1209_U178 );
nand NAND2_15058 ( P2_R1209_U181 , P2_U3386 , P2_R1209_U8 );
nand NAND2_15059 ( P2_R1209_U182 , P2_REG1_REG_9_ , P2_R1209_U27 );
nand NAND2_15060 ( P2_R1209_U183 , P2_U3415 , P2_R1209_U26 );
not NOT1_15061 ( P2_R1209_U184 , P2_R1209_U67 );
nand NAND2_15062 ( P2_R1209_U185 , P2_R1209_U136 , P2_R1209_U184 );
nand NAND2_15063 ( P2_R1209_U186 , P2_R1209_U67 , P2_R1209_U87 );
nand NAND2_15064 ( P2_R1209_U187 , P2_REG1_REG_8_ , P2_R1209_U25 );
nand NAND2_15065 ( P2_R1209_U188 , P2_U3412 , P2_R1209_U24 );
not NOT1_15066 ( P2_R1209_U189 , P2_R1209_U68 );
nand NAND2_15067 ( P2_R1209_U190 , P2_R1209_U132 , P2_R1209_U189 );
nand NAND2_15068 ( P2_R1209_U191 , P2_R1209_U68 , P2_R1209_U88 );
nand NAND2_15069 ( P2_R1209_U192 , P2_REG1_REG_7_ , P2_R1209_U23 );
nand NAND2_15070 ( P2_R1209_U193 , P2_U3409 , P2_R1209_U22 );
not NOT1_15071 ( P2_R1209_U194 , P2_R1209_U69 );
nand NAND2_15072 ( P2_R1209_U195 , P2_R1209_U128 , P2_R1209_U194 );
nand NAND2_15073 ( P2_R1209_U196 , P2_R1209_U69 , P2_R1209_U89 );
nand NAND2_15074 ( P2_R1209_U197 , P2_REG1_REG_6_ , P2_R1209_U21 );
nand NAND2_15075 ( P2_R1209_U198 , P2_U3406 , P2_R1209_U20 );
not NOT1_15076 ( P2_R1209_U199 , P2_R1209_U70 );
nand NAND2_15077 ( P2_R1209_U200 , P2_R1209_U124 , P2_R1209_U199 );
nand NAND2_15078 ( P2_R1209_U201 , P2_R1209_U70 , P2_R1209_U90 );
nand NAND2_15079 ( P2_R1209_U202 , P2_REG1_REG_5_ , P2_R1209_U19 );
nand NAND2_15080 ( P2_R1209_U203 , P2_U3403 , P2_R1209_U18 );
not NOT1_15081 ( P2_R1209_U204 , P2_R1209_U71 );
nand NAND2_15082 ( P2_R1209_U205 , P2_R1209_U120 , P2_R1209_U204 );
nand NAND2_15083 ( P2_R1209_U206 , P2_R1209_U71 , P2_R1209_U91 );
nand NAND2_15084 ( P2_R1209_U207 , P2_REG1_REG_4_ , P2_R1209_U17 );
nand NAND2_15085 ( P2_R1209_U208 , P2_U3400 , P2_R1209_U16 );
not NOT1_15086 ( P2_R1209_U209 , P2_R1209_U72 );
nand NAND2_15087 ( P2_R1209_U210 , P2_R1209_U116 , P2_R1209_U209 );
nand NAND2_15088 ( P2_R1209_U211 , P2_R1209_U72 , P2_R1209_U92 );
nand NAND2_15089 ( P2_R1209_U212 , P2_REG1_REG_3_ , P2_R1209_U15 );
nand NAND2_15090 ( P2_R1209_U213 , P2_U3397 , P2_R1209_U14 );
not NOT1_15091 ( P2_R1209_U214 , P2_R1209_U73 );
nand NAND2_15092 ( P2_R1209_U215 , P2_R1209_U112 , P2_R1209_U214 );
nand NAND2_15093 ( P2_R1209_U216 , P2_R1209_U73 , P2_R1209_U93 );
nand NAND2_15094 ( P2_R1209_U217 , P2_REG1_REG_2_ , P2_R1209_U13 );
nand NAND2_15095 ( P2_R1209_U218 , P2_U3394 , P2_R1209_U12 );
not NOT1_15096 ( P2_R1209_U219 , P2_R1209_U74 );
nand NAND2_15097 ( P2_R1209_U220 , P2_R1209_U108 , P2_R1209_U219 );
nand NAND2_15098 ( P2_R1209_U221 , P2_R1209_U74 , P2_R1209_U94 );
nand NAND2_15099 ( P2_R1209_U222 , P2_R1209_U104 , P2_R1209_U10 );
nand NAND2_15100 ( P2_R1209_U223 , P2_REG1_REG_1_ , P2_R1209_U9 );
not NOT1_15101 ( P2_R1209_U224 , P2_R1209_U75 );
nand NAND2_15102 ( P2_R1209_U225 , P2_R1209_U224 , P2_U3391 );
nand NAND2_15103 ( P2_R1209_U226 , P2_R1209_U75 , P2_R1209_U11 );
nand NAND2_15104 ( P2_R1209_U227 , P2_REG1_REG_19_ , P2_R1209_U96 );
nand NAND2_15105 ( P2_R1209_U228 , P2_U3379 , P2_R1209_U95 );
nand NAND2_15106 ( P2_R1209_U229 , P2_REG1_REG_19_ , P2_R1209_U96 );
nand NAND2_15107 ( P2_R1209_U230 , P2_U3379 , P2_R1209_U95 );
nand NAND2_15108 ( P2_R1209_U231 , P2_R1209_U230 , P2_R1209_U229 );
nand NAND2_15109 ( P2_R1209_U232 , P2_REG1_REG_18_ , P2_R1209_U46 );
nand NAND2_15110 ( P2_R1209_U233 , P2_U3442 , P2_R1209_U45 );
not NOT1_15111 ( P2_R1209_U234 , P2_R1209_U78 );
nand NAND2_15112 ( P2_R1209_U235 , P2_R1209_U234 , P2_R1209_U172 );
nand NAND2_15113 ( P2_R1209_U236 , P2_R1209_U78 , P2_R1209_U47 );
nand NAND2_15114 ( P2_R1209_U237 , P2_REG1_REG_17_ , P2_R1209_U44 );
nand NAND2_15115 ( P2_R1209_U238 , P2_U3439 , P2_R1209_U43 );
not NOT1_15116 ( P2_R1209_U239 , P2_R1209_U79 );
nand NAND2_15117 ( P2_R1209_U240 , P2_R1209_U168 , P2_R1209_U239 );
nand NAND2_15118 ( P2_R1209_U241 , P2_R1209_U79 , P2_R1209_U97 );
nand NAND2_15119 ( P2_R1209_U242 , P2_REG1_REG_16_ , P2_R1209_U42 );
nand NAND2_15120 ( P2_R1209_U243 , P2_U3436 , P2_R1209_U41 );
not NOT1_15121 ( P2_R1209_U244 , P2_R1209_U80 );
nand NAND2_15122 ( P2_R1209_U245 , P2_R1209_U164 , P2_R1209_U244 );
nand NAND2_15123 ( P2_R1209_U246 , P2_R1209_U80 , P2_R1209_U98 );
nand NAND2_15124 ( P2_R1209_U247 , P2_U3433 , P2_R1209_U39 );
nand NAND2_15125 ( P2_R1209_U248 , P2_REG1_REG_15_ , P2_R1209_U40 );
not NOT1_15126 ( P2_R1209_U249 , P2_R1209_U81 );
nand NAND2_15127 ( P2_R1209_U250 , P2_R1209_U249 , P2_R1209_U160 );
nand NAND2_15128 ( P2_R1209_U251 , P2_R1209_U81 , P2_R1209_U38 );
nand NAND2_15129 ( P2_R1209_U252 , P2_REG1_REG_14_ , P2_R1209_U37 );
nand NAND2_15130 ( P2_R1209_U253 , P2_U3430 , P2_R1209_U36 );
not NOT1_15131 ( P2_R1209_U254 , P2_R1209_U82 );
nand NAND2_15132 ( P2_R1209_U255 , P2_R1209_U156 , P2_R1209_U254 );
nand NAND2_15133 ( P2_R1209_U256 , P2_R1209_U82 , P2_R1209_U99 );
nand NAND2_15134 ( P2_R1209_U257 , P2_REG1_REG_13_ , P2_R1209_U35 );
nand NAND2_15135 ( P2_R1209_U258 , P2_U3427 , P2_R1209_U34 );
not NOT1_15136 ( P2_R1209_U259 , P2_R1209_U83 );
nand NAND2_15137 ( P2_R1209_U260 , P2_R1209_U152 , P2_R1209_U259 );
nand NAND2_15138 ( P2_R1209_U261 , P2_R1209_U83 , P2_R1209_U100 );
nand NAND2_15139 ( P2_R1209_U262 , P2_REG1_REG_12_ , P2_R1209_U33 );
nand NAND2_15140 ( P2_R1209_U263 , P2_U3424 , P2_R1209_U32 );
not NOT1_15141 ( P2_R1209_U264 , P2_R1209_U84 );
nand NAND2_15142 ( P2_R1209_U265 , P2_R1209_U148 , P2_R1209_U264 );
nand NAND2_15143 ( P2_R1209_U266 , P2_R1209_U84 , P2_R1209_U101 );
nand NAND2_15144 ( P2_R1209_U267 , P2_REG1_REG_11_ , P2_R1209_U31 );
nand NAND2_15145 ( P2_R1209_U268 , P2_U3421 , P2_R1209_U30 );
not NOT1_15146 ( P2_R1209_U269 , P2_R1209_U85 );
nand NAND2_15147 ( P2_R1209_U270 , P2_R1209_U144 , P2_R1209_U269 );
nand NAND2_15148 ( P2_R1209_U271 , P2_R1209_U85 , P2_R1209_U102 );
nand NAND2_15149 ( P2_R1209_U272 , P2_REG1_REG_10_ , P2_R1209_U29 );
nand NAND2_15150 ( P2_R1209_U273 , P2_U3418 , P2_R1209_U28 );
not NOT1_15151 ( P2_R1209_U274 , P2_R1209_U86 );
nand NAND2_15152 ( P2_R1209_U275 , P2_R1209_U140 , P2_R1209_U274 );
nand NAND2_15153 ( P2_R1209_U276 , P2_R1209_U86 , P2_R1209_U103 );
not NOT1_15154 ( P2_R1300_U6 , P2_U3058 );
not NOT1_15155 ( P2_R1300_U7 , P2_U3055 );
and AND2_15156 ( P2_R1300_U8 , P2_R1300_U10 , P2_R1300_U9 );
nand NAND2_15157 ( P2_R1300_U9 , P2_U3055 , P2_R1300_U6 );
nand NAND2_15158 ( P2_R1300_U10 , P2_U3058 , P2_R1300_U7 );
and AND2_15159 ( P2_R1200_U6 , P2_R1200_U212 , P2_R1200_U211 );
and AND2_15160 ( P2_R1200_U7 , P2_R1200_U246 , P2_R1200_U245 );
and AND2_15161 ( P2_R1200_U8 , P2_R1200_U193 , P2_R1200_U257 );
and AND2_15162 ( P2_R1200_U9 , P2_R1200_U259 , P2_R1200_U258 );
and AND2_15163 ( P2_R1200_U10 , P2_R1200_U194 , P2_R1200_U281 );
and AND2_15164 ( P2_R1200_U11 , P2_R1200_U283 , P2_R1200_U282 );
and AND2_15165 ( P2_R1200_U12 , P2_R1200_U299 , P2_R1200_U195 );
and AND3_15166 ( P2_R1200_U13 , P2_R1200_U210 , P2_R1200_U197 , P2_R1200_U215 );
and AND2_15167 ( P2_R1200_U14 , P2_R1200_U220 , P2_R1200_U198 );
and AND3_15168 ( P2_R1200_U15 , P2_R1200_U224 , P2_R1200_U192 , P2_R1200_U244 );
and AND2_15169 ( P2_R1200_U16 , P2_R1200_U399 , P2_R1200_U398 );
nand NAND2_15170 ( P2_R1200_U17 , P2_R1200_U331 , P2_R1200_U334 );
nand NAND2_15171 ( P2_R1200_U18 , P2_R1200_U322 , P2_R1200_U325 );
nand NAND2_15172 ( P2_R1200_U19 , P2_R1200_U311 , P2_R1200_U314 );
nand NAND2_15173 ( P2_R1200_U20 , P2_R1200_U305 , P2_R1200_U357 );
nand NAND2_15174 ( P2_R1200_U21 , P2_R1200_U137 , P2_R1200_U186 );
nand NAND2_15175 ( P2_R1200_U22 , P2_R1200_U242 , P2_R1200_U347 );
nand NAND2_15176 ( P2_R1200_U23 , P2_R1200_U235 , P2_R1200_U238 );
nand NAND2_15177 ( P2_R1200_U24 , P2_R1200_U227 , P2_R1200_U229 );
nand NAND2_15178 ( P2_R1200_U25 , P2_R1200_U175 , P2_R1200_U337 );
not NOT1_15179 ( P2_R1200_U26 , P2_U3069 );
nand NAND2_15180 ( P2_R1200_U27 , P2_U3069 , P2_R1200_U32 );
not NOT1_15181 ( P2_R1200_U28 , P2_U3083 );
not NOT1_15182 ( P2_R1200_U29 , P2_U3404 );
not NOT1_15183 ( P2_R1200_U30 , P2_U3407 );
not NOT1_15184 ( P2_R1200_U31 , P2_U3401 );
not NOT1_15185 ( P2_R1200_U32 , P2_U3410 );
not NOT1_15186 ( P2_R1200_U33 , P2_U3413 );
not NOT1_15187 ( P2_R1200_U34 , P2_U3067 );
nand NAND2_15188 ( P2_R1200_U35 , P2_U3067 , P2_R1200_U37 );
not NOT1_15189 ( P2_R1200_U36 , P2_U3063 );
not NOT1_15190 ( P2_R1200_U37 , P2_U3395 );
not NOT1_15191 ( P2_R1200_U38 , P2_U3387 );
not NOT1_15192 ( P2_R1200_U39 , P2_U3077 );
not NOT1_15193 ( P2_R1200_U40 , P2_U3398 );
not NOT1_15194 ( P2_R1200_U41 , P2_U3070 );
not NOT1_15195 ( P2_R1200_U42 , P2_U3066 );
not NOT1_15196 ( P2_R1200_U43 , P2_U3059 );
nand NAND2_15197 ( P2_R1200_U44 , P2_U3059 , P2_R1200_U31 );
nand NAND2_15198 ( P2_R1200_U45 , P2_R1200_U216 , P2_R1200_U214 );
not NOT1_15199 ( P2_R1200_U46 , P2_U3416 );
not NOT1_15200 ( P2_R1200_U47 , P2_U3082 );
nand NAND2_15201 ( P2_R1200_U48 , P2_R1200_U45 , P2_R1200_U217 );
nand NAND2_15202 ( P2_R1200_U49 , P2_R1200_U44 , P2_R1200_U231 );
nand NAND3_15203 ( P2_R1200_U50 , P2_R1200_U204 , P2_R1200_U188 , P2_R1200_U338 );
not NOT1_15204 ( P2_R1200_U51 , P2_U3895 );
not NOT1_15205 ( P2_R1200_U52 , P2_U3056 );
nand NAND2_15206 ( P2_R1200_U53 , P2_U3056 , P2_R1200_U90 );
not NOT1_15207 ( P2_R1200_U54 , P2_U3052 );
not NOT1_15208 ( P2_R1200_U55 , P2_U3071 );
not NOT1_15209 ( P2_R1200_U56 , P2_U3062 );
not NOT1_15210 ( P2_R1200_U57 , P2_U3061 );
not NOT1_15211 ( P2_R1200_U58 , P2_U3419 );
nand NAND2_15212 ( P2_R1200_U59 , P2_U3082 , P2_R1200_U46 );
not NOT1_15213 ( P2_R1200_U60 , P2_U3422 );
not NOT1_15214 ( P2_R1200_U61 , P2_U3425 );
nand NAND2_15215 ( P2_R1200_U62 , P2_R1200_U249 , P2_R1200_U248 );
not NOT1_15216 ( P2_R1200_U63 , P2_U3428 );
not NOT1_15217 ( P2_R1200_U64 , P2_U3079 );
not NOT1_15218 ( P2_R1200_U65 , P2_U3437 );
not NOT1_15219 ( P2_R1200_U66 , P2_U3434 );
not NOT1_15220 ( P2_R1200_U67 , P2_U3431 );
not NOT1_15221 ( P2_R1200_U68 , P2_U3072 );
not NOT1_15222 ( P2_R1200_U69 , P2_U3073 );
not NOT1_15223 ( P2_R1200_U70 , P2_U3078 );
nand NAND2_15224 ( P2_R1200_U71 , P2_U3078 , P2_R1200_U67 );
not NOT1_15225 ( P2_R1200_U72 , P2_U3440 );
not NOT1_15226 ( P2_R1200_U73 , P2_U3068 );
not NOT1_15227 ( P2_R1200_U74 , P2_U3081 );
not NOT1_15228 ( P2_R1200_U75 , P2_U3445 );
not NOT1_15229 ( P2_R1200_U76 , P2_U3080 );
not NOT1_15230 ( P2_R1200_U77 , P2_U3903 );
not NOT1_15231 ( P2_R1200_U78 , P2_U3075 );
not NOT1_15232 ( P2_R1200_U79 , P2_U3900 );
not NOT1_15233 ( P2_R1200_U80 , P2_U3901 );
not NOT1_15234 ( P2_R1200_U81 , P2_U3902 );
not NOT1_15235 ( P2_R1200_U82 , P2_U3065 );
not NOT1_15236 ( P2_R1200_U83 , P2_U3060 );
not NOT1_15237 ( P2_R1200_U84 , P2_U3074 );
nand NAND2_15238 ( P2_R1200_U85 , P2_U3074 , P2_R1200_U81 );
not NOT1_15239 ( P2_R1200_U86 , P2_U3899 );
not NOT1_15240 ( P2_R1200_U87 , P2_U3064 );
not NOT1_15241 ( P2_R1200_U88 , P2_U3898 );
not NOT1_15242 ( P2_R1200_U89 , P2_U3057 );
not NOT1_15243 ( P2_R1200_U90 , P2_U3897 );
not NOT1_15244 ( P2_R1200_U91 , P2_U3896 );
not NOT1_15245 ( P2_R1200_U92 , P2_U3053 );
nand NAND2_15246 ( P2_R1200_U93 , P2_R1200_U297 , P2_R1200_U296 );
nand NAND2_15247 ( P2_R1200_U94 , P2_R1200_U85 , P2_R1200_U307 );
nand NAND2_15248 ( P2_R1200_U95 , P2_R1200_U71 , P2_R1200_U318 );
nand NAND2_15249 ( P2_R1200_U96 , P2_R1200_U349 , P2_R1200_U59 );
not NOT1_15250 ( P2_R1200_U97 , P2_U3076 );
nand NAND2_15251 ( P2_R1200_U98 , P2_R1200_U406 , P2_R1200_U405 );
nand NAND2_15252 ( P2_R1200_U99 , P2_R1200_U420 , P2_R1200_U419 );
nand NAND2_15253 ( P2_R1200_U100 , P2_R1200_U425 , P2_R1200_U424 );
nand NAND2_15254 ( P2_R1200_U101 , P2_R1200_U441 , P2_R1200_U440 );
nand NAND2_15255 ( P2_R1200_U102 , P2_R1200_U446 , P2_R1200_U445 );
nand NAND2_15256 ( P2_R1200_U103 , P2_R1200_U451 , P2_R1200_U450 );
nand NAND2_15257 ( P2_R1200_U104 , P2_R1200_U456 , P2_R1200_U455 );
nand NAND2_15258 ( P2_R1200_U105 , P2_R1200_U461 , P2_R1200_U460 );
nand NAND2_15259 ( P2_R1200_U106 , P2_R1200_U477 , P2_R1200_U476 );
nand NAND2_15260 ( P2_R1200_U107 , P2_R1200_U482 , P2_R1200_U481 );
nand NAND2_15261 ( P2_R1200_U108 , P2_R1200_U365 , P2_R1200_U364 );
nand NAND2_15262 ( P2_R1200_U109 , P2_R1200_U374 , P2_R1200_U373 );
nand NAND2_15263 ( P2_R1200_U110 , P2_R1200_U381 , P2_R1200_U380 );
nand NAND2_15264 ( P2_R1200_U111 , P2_R1200_U385 , P2_R1200_U384 );
nand NAND2_15265 ( P2_R1200_U112 , P2_R1200_U394 , P2_R1200_U393 );
nand NAND2_15266 ( P2_R1200_U113 , P2_R1200_U415 , P2_R1200_U414 );
nand NAND2_15267 ( P2_R1200_U114 , P2_R1200_U432 , P2_R1200_U431 );
nand NAND2_15268 ( P2_R1200_U115 , P2_R1200_U436 , P2_R1200_U435 );
nand NAND2_15269 ( P2_R1200_U116 , P2_R1200_U468 , P2_R1200_U467 );
nand NAND2_15270 ( P2_R1200_U117 , P2_R1200_U472 , P2_R1200_U471 );
nand NAND2_15271 ( P2_R1200_U118 , P2_R1200_U489 , P2_R1200_U488 );
and AND2_15272 ( P2_R1200_U119 , P2_R1200_U206 , P2_R1200_U196 );
and AND2_15273 ( P2_R1200_U120 , P2_R1200_U209 , P2_R1200_U208 );
and AND2_15274 ( P2_R1200_U121 , P2_R1200_U14 , P2_R1200_U13 );
and AND2_15275 ( P2_R1200_U122 , P2_R1200_U340 , P2_R1200_U222 );
and AND2_15276 ( P2_R1200_U123 , P2_R1200_U342 , P2_R1200_U122 );
and AND3_15277 ( P2_R1200_U124 , P2_R1200_U367 , P2_R1200_U366 , P2_R1200_U27 );
and AND2_15278 ( P2_R1200_U125 , P2_R1200_U370 , P2_R1200_U198 );
and AND2_15279 ( P2_R1200_U126 , P2_R1200_U237 , P2_R1200_U6 );
and AND2_15280 ( P2_R1200_U127 , P2_R1200_U377 , P2_R1200_U197 );
and AND3_15281 ( P2_R1200_U128 , P2_R1200_U387 , P2_R1200_U386 , P2_R1200_U35 );
and AND2_15282 ( P2_R1200_U129 , P2_R1200_U390 , P2_R1200_U196 );
and AND2_15283 ( P2_R1200_U130 , P2_R1200_U251 , P2_R1200_U15 );
and AND2_15284 ( P2_R1200_U131 , P2_R1200_U343 , P2_R1200_U252 );
and AND2_15285 ( P2_R1200_U132 , P2_R1200_U262 , P2_R1200_U8 );
and AND2_15286 ( P2_R1200_U133 , P2_R1200_U286 , P2_R1200_U10 );
and AND2_15287 ( P2_R1200_U134 , P2_R1200_U302 , P2_R1200_U301 );
and AND2_15288 ( P2_R1200_U135 , P2_R1200_U397 , P2_R1200_U303 );
and AND4_15289 ( P2_R1200_U136 , P2_R1200_U302 , P2_R1200_U301 , P2_R1200_U304 , P2_R1200_U16 );
and AND2_15290 ( P2_R1200_U137 , P2_R1200_U359 , P2_R1200_U165 );
nand NAND2_15291 ( P2_R1200_U138 , P2_R1200_U403 , P2_R1200_U402 );
and AND3_15292 ( P2_R1200_U139 , P2_R1200_U408 , P2_R1200_U407 , P2_R1200_U53 );
and AND2_15293 ( P2_R1200_U140 , P2_R1200_U411 , P2_R1200_U195 );
nand NAND2_15294 ( P2_R1200_U141 , P2_R1200_U417 , P2_R1200_U416 );
nand NAND2_15295 ( P2_R1200_U142 , P2_R1200_U422 , P2_R1200_U421 );
and AND2_15296 ( P2_R1200_U143 , P2_R1200_U313 , P2_R1200_U11 );
and AND2_15297 ( P2_R1200_U144 , P2_R1200_U428 , P2_R1200_U194 );
nand NAND2_15298 ( P2_R1200_U145 , P2_R1200_U438 , P2_R1200_U437 );
nand NAND2_15299 ( P2_R1200_U146 , P2_R1200_U443 , P2_R1200_U442 );
nand NAND2_15300 ( P2_R1200_U147 , P2_R1200_U448 , P2_R1200_U447 );
nand NAND2_15301 ( P2_R1200_U148 , P2_R1200_U453 , P2_R1200_U452 );
nand NAND2_15302 ( P2_R1200_U149 , P2_R1200_U458 , P2_R1200_U457 );
and AND2_15303 ( P2_R1200_U150 , P2_R1200_U324 , P2_R1200_U9 );
and AND2_15304 ( P2_R1200_U151 , P2_R1200_U464 , P2_R1200_U193 );
nand NAND2_15305 ( P2_R1200_U152 , P2_R1200_U474 , P2_R1200_U473 );
nand NAND2_15306 ( P2_R1200_U153 , P2_R1200_U479 , P2_R1200_U478 );
and AND2_15307 ( P2_R1200_U154 , P2_R1200_U333 , P2_R1200_U7 );
and AND2_15308 ( P2_R1200_U155 , P2_R1200_U485 , P2_R1200_U192 );
and AND2_15309 ( P2_R1200_U156 , P2_R1200_U363 , P2_R1200_U362 );
nand NAND2_15310 ( P2_R1200_U157 , P2_R1200_U123 , P2_R1200_U341 );
and AND2_15311 ( P2_R1200_U158 , P2_R1200_U372 , P2_R1200_U371 );
and AND2_15312 ( P2_R1200_U159 , P2_R1200_U379 , P2_R1200_U378 );
and AND2_15313 ( P2_R1200_U160 , P2_R1200_U383 , P2_R1200_U382 );
nand NAND2_15314 ( P2_R1200_U161 , P2_R1200_U120 , P2_R1200_U344 );
and AND2_15315 ( P2_R1200_U162 , P2_R1200_U392 , P2_R1200_U391 );
not NOT1_15316 ( P2_R1200_U163 , P2_U3904 );
not NOT1_15317 ( P2_R1200_U164 , P2_U3054 );
and AND2_15318 ( P2_R1200_U165 , P2_R1200_U401 , P2_R1200_U400 );
nand NAND2_15319 ( P2_R1200_U166 , P2_R1200_U134 , P2_R1200_U360 );
and AND2_15320 ( P2_R1200_U167 , P2_R1200_U413 , P2_R1200_U412 );
nand NAND2_15321 ( P2_R1200_U168 , P2_R1200_U293 , P2_R1200_U292 );
nand NAND2_15322 ( P2_R1200_U169 , P2_R1200_U289 , P2_R1200_U288 );
and AND2_15323 ( P2_R1200_U170 , P2_R1200_U430 , P2_R1200_U429 );
and AND2_15324 ( P2_R1200_U171 , P2_R1200_U434 , P2_R1200_U433 );
nand NAND2_15325 ( P2_R1200_U172 , P2_R1200_U279 , P2_R1200_U278 );
nand NAND2_15326 ( P2_R1200_U173 , P2_R1200_U275 , P2_R1200_U274 );
not NOT1_15327 ( P2_R1200_U174 , P2_U3392 );
nand NAND2_15328 ( P2_R1200_U175 , P2_U3387 , P2_R1200_U97 );
nand NAND3_15329 ( P2_R1200_U176 , P2_R1200_U271 , P2_R1200_U187 , P2_R1200_U339 );
not NOT1_15330 ( P2_R1200_U177 , P2_U3443 );
nand NAND2_15331 ( P2_R1200_U178 , P2_R1200_U269 , P2_R1200_U268 );
nand NAND2_15332 ( P2_R1200_U179 , P2_R1200_U265 , P2_R1200_U264 );
and AND2_15333 ( P2_R1200_U180 , P2_R1200_U466 , P2_R1200_U465 );
and AND2_15334 ( P2_R1200_U181 , P2_R1200_U470 , P2_R1200_U469 );
nand NAND2_15335 ( P2_R1200_U182 , P2_R1200_U255 , P2_R1200_U254 );
nand NAND2_15336 ( P2_R1200_U183 , P2_R1200_U131 , P2_R1200_U353 );
nand NAND2_15337 ( P2_R1200_U184 , P2_R1200_U351 , P2_R1200_U62 );
and AND2_15338 ( P2_R1200_U185 , P2_R1200_U487 , P2_R1200_U486 );
nand NAND2_15339 ( P2_R1200_U186 , P2_R1200_U135 , P2_R1200_U166 );
nand NAND2_15340 ( P2_R1200_U187 , P2_R1200_U178 , P2_R1200_U177 );
nand NAND2_15341 ( P2_R1200_U188 , P2_R1200_U175 , P2_R1200_U174 );
not NOT1_15342 ( P2_R1200_U189 , P2_R1200_U53 );
not NOT1_15343 ( P2_R1200_U190 , P2_R1200_U35 );
not NOT1_15344 ( P2_R1200_U191 , P2_R1200_U27 );
nand NAND2_15345 ( P2_R1200_U192 , P2_U3419 , P2_R1200_U57 );
nand NAND2_15346 ( P2_R1200_U193 , P2_U3434 , P2_R1200_U69 );
nand NAND2_15347 ( P2_R1200_U194 , P2_U3901 , P2_R1200_U83 );
nand NAND2_15348 ( P2_R1200_U195 , P2_U3897 , P2_R1200_U52 );
nand NAND2_15349 ( P2_R1200_U196 , P2_U3395 , P2_R1200_U34 );
nand NAND2_15350 ( P2_R1200_U197 , P2_U3404 , P2_R1200_U42 );
nand NAND2_15351 ( P2_R1200_U198 , P2_U3410 , P2_R1200_U26 );
not NOT1_15352 ( P2_R1200_U199 , P2_R1200_U71 );
not NOT1_15353 ( P2_R1200_U200 , P2_R1200_U85 );
not NOT1_15354 ( P2_R1200_U201 , P2_R1200_U44 );
not NOT1_15355 ( P2_R1200_U202 , P2_R1200_U59 );
not NOT1_15356 ( P2_R1200_U203 , P2_R1200_U175 );
nand NAND2_15357 ( P2_R1200_U204 , P2_U3077 , P2_R1200_U175 );
not NOT1_15358 ( P2_R1200_U205 , P2_R1200_U50 );
nand NAND2_15359 ( P2_R1200_U206 , P2_U3398 , P2_R1200_U36 );
nand NAND2_15360 ( P2_R1200_U207 , P2_R1200_U36 , P2_R1200_U35 );
nand NAND2_15361 ( P2_R1200_U208 , P2_R1200_U207 , P2_R1200_U40 );
nand NAND2_15362 ( P2_R1200_U209 , P2_U3063 , P2_R1200_U190 );
nand NAND2_15363 ( P2_R1200_U210 , P2_U3407 , P2_R1200_U41 );
nand NAND2_15364 ( P2_R1200_U211 , P2_U3070 , P2_R1200_U30 );
nand NAND2_15365 ( P2_R1200_U212 , P2_U3066 , P2_R1200_U29 );
nand NAND2_15366 ( P2_R1200_U213 , P2_R1200_U201 , P2_R1200_U197 );
nand NAND2_15367 ( P2_R1200_U214 , P2_R1200_U6 , P2_R1200_U213 );
nand NAND2_15368 ( P2_R1200_U215 , P2_U3401 , P2_R1200_U43 );
nand NAND2_15369 ( P2_R1200_U216 , P2_U3407 , P2_R1200_U41 );
nand NAND2_15370 ( P2_R1200_U217 , P2_R1200_U13 , P2_R1200_U161 );
not NOT1_15371 ( P2_R1200_U218 , P2_R1200_U45 );
not NOT1_15372 ( P2_R1200_U219 , P2_R1200_U48 );
nand NAND2_15373 ( P2_R1200_U220 , P2_U3413 , P2_R1200_U28 );
nand NAND2_15374 ( P2_R1200_U221 , P2_R1200_U28 , P2_R1200_U27 );
nand NAND2_15375 ( P2_R1200_U222 , P2_U3083 , P2_R1200_U191 );
not NOT1_15376 ( P2_R1200_U223 , P2_R1200_U157 );
nand NAND2_15377 ( P2_R1200_U224 , P2_U3416 , P2_R1200_U47 );
nand NAND2_15378 ( P2_R1200_U225 , P2_R1200_U224 , P2_R1200_U59 );
nand NAND2_15379 ( P2_R1200_U226 , P2_R1200_U219 , P2_R1200_U27 );
nand NAND2_15380 ( P2_R1200_U227 , P2_R1200_U125 , P2_R1200_U226 );
nand NAND2_15381 ( P2_R1200_U228 , P2_R1200_U48 , P2_R1200_U198 );
nand NAND2_15382 ( P2_R1200_U229 , P2_R1200_U124 , P2_R1200_U228 );
nand NAND2_15383 ( P2_R1200_U230 , P2_R1200_U27 , P2_R1200_U198 );
nand NAND2_15384 ( P2_R1200_U231 , P2_R1200_U215 , P2_R1200_U161 );
not NOT1_15385 ( P2_R1200_U232 , P2_R1200_U49 );
nand NAND2_15386 ( P2_R1200_U233 , P2_U3066 , P2_R1200_U29 );
nand NAND2_15387 ( P2_R1200_U234 , P2_R1200_U232 , P2_R1200_U233 );
nand NAND2_15388 ( P2_R1200_U235 , P2_R1200_U127 , P2_R1200_U234 );
nand NAND2_15389 ( P2_R1200_U236 , P2_R1200_U49 , P2_R1200_U197 );
nand NAND2_15390 ( P2_R1200_U237 , P2_U3407 , P2_R1200_U41 );
nand NAND2_15391 ( P2_R1200_U238 , P2_R1200_U126 , P2_R1200_U236 );
nand NAND2_15392 ( P2_R1200_U239 , P2_U3066 , P2_R1200_U29 );
nand NAND2_15393 ( P2_R1200_U240 , P2_R1200_U239 , P2_R1200_U197 );
nand NAND2_15394 ( P2_R1200_U241 , P2_R1200_U215 , P2_R1200_U44 );
nand NAND2_15395 ( P2_R1200_U242 , P2_R1200_U129 , P2_R1200_U348 );
nand NAND2_15396 ( P2_R1200_U243 , P2_R1200_U35 , P2_R1200_U196 );
nand NAND2_15397 ( P2_R1200_U244 , P2_U3422 , P2_R1200_U56 );
nand NAND2_15398 ( P2_R1200_U245 , P2_U3062 , P2_R1200_U60 );
nand NAND2_15399 ( P2_R1200_U246 , P2_U3061 , P2_R1200_U58 );
nand NAND2_15400 ( P2_R1200_U247 , P2_R1200_U202 , P2_R1200_U192 );
nand NAND2_15401 ( P2_R1200_U248 , P2_R1200_U7 , P2_R1200_U247 );
nand NAND2_15402 ( P2_R1200_U249 , P2_U3422 , P2_R1200_U56 );
not NOT1_15403 ( P2_R1200_U250 , P2_R1200_U62 );
nand NAND2_15404 ( P2_R1200_U251 , P2_U3425 , P2_R1200_U55 );
nand NAND2_15405 ( P2_R1200_U252 , P2_U3071 , P2_R1200_U61 );
nand NAND2_15406 ( P2_R1200_U253 , P2_U3428 , P2_R1200_U64 );
nand NAND2_15407 ( P2_R1200_U254 , P2_R1200_U253 , P2_R1200_U183 );
nand NAND2_15408 ( P2_R1200_U255 , P2_U3079 , P2_R1200_U63 );
not NOT1_15409 ( P2_R1200_U256 , P2_R1200_U182 );
nand NAND2_15410 ( P2_R1200_U257 , P2_U3437 , P2_R1200_U68 );
nand NAND2_15411 ( P2_R1200_U258 , P2_U3072 , P2_R1200_U65 );
nand NAND2_15412 ( P2_R1200_U259 , P2_U3073 , P2_R1200_U66 );
nand NAND2_15413 ( P2_R1200_U260 , P2_R1200_U199 , P2_R1200_U8 );
nand NAND2_15414 ( P2_R1200_U261 , P2_R1200_U9 , P2_R1200_U260 );
nand NAND2_15415 ( P2_R1200_U262 , P2_U3431 , P2_R1200_U70 );
nand NAND2_15416 ( P2_R1200_U263 , P2_U3437 , P2_R1200_U68 );
nand NAND2_15417 ( P2_R1200_U264 , P2_R1200_U132 , P2_R1200_U182 );
nand NAND2_15418 ( P2_R1200_U265 , P2_R1200_U263 , P2_R1200_U261 );
not NOT1_15419 ( P2_R1200_U266 , P2_R1200_U179 );
nand NAND2_15420 ( P2_R1200_U267 , P2_U3440 , P2_R1200_U73 );
nand NAND2_15421 ( P2_R1200_U268 , P2_R1200_U267 , P2_R1200_U179 );
nand NAND2_15422 ( P2_R1200_U269 , P2_U3068 , P2_R1200_U72 );
not NOT1_15423 ( P2_R1200_U270 , P2_R1200_U178 );
nand NAND2_15424 ( P2_R1200_U271 , P2_U3081 , P2_R1200_U178 );
not NOT1_15425 ( P2_R1200_U272 , P2_R1200_U176 );
nand NAND2_15426 ( P2_R1200_U273 , P2_U3445 , P2_R1200_U76 );
nand NAND2_15427 ( P2_R1200_U274 , P2_R1200_U273 , P2_R1200_U176 );
nand NAND2_15428 ( P2_R1200_U275 , P2_U3080 , P2_R1200_U75 );
not NOT1_15429 ( P2_R1200_U276 , P2_R1200_U173 );
nand NAND2_15430 ( P2_R1200_U277 , P2_U3903 , P2_R1200_U78 );
nand NAND2_15431 ( P2_R1200_U278 , P2_R1200_U277 , P2_R1200_U173 );
nand NAND2_15432 ( P2_R1200_U279 , P2_U3075 , P2_R1200_U77 );
not NOT1_15433 ( P2_R1200_U280 , P2_R1200_U172 );
nand NAND2_15434 ( P2_R1200_U281 , P2_U3900 , P2_R1200_U82 );
nand NAND2_15435 ( P2_R1200_U282 , P2_U3065 , P2_R1200_U79 );
nand NAND2_15436 ( P2_R1200_U283 , P2_U3060 , P2_R1200_U80 );
nand NAND2_15437 ( P2_R1200_U284 , P2_R1200_U200 , P2_R1200_U10 );
nand NAND2_15438 ( P2_R1200_U285 , P2_R1200_U11 , P2_R1200_U284 );
nand NAND2_15439 ( P2_R1200_U286 , P2_U3902 , P2_R1200_U84 );
nand NAND2_15440 ( P2_R1200_U287 , P2_U3900 , P2_R1200_U82 );
nand NAND2_15441 ( P2_R1200_U288 , P2_R1200_U133 , P2_R1200_U172 );
nand NAND2_15442 ( P2_R1200_U289 , P2_R1200_U287 , P2_R1200_U285 );
not NOT1_15443 ( P2_R1200_U290 , P2_R1200_U169 );
nand NAND2_15444 ( P2_R1200_U291 , P2_U3899 , P2_R1200_U87 );
nand NAND2_15445 ( P2_R1200_U292 , P2_R1200_U291 , P2_R1200_U169 );
nand NAND2_15446 ( P2_R1200_U293 , P2_U3064 , P2_R1200_U86 );
not NOT1_15447 ( P2_R1200_U294 , P2_R1200_U168 );
nand NAND2_15448 ( P2_R1200_U295 , P2_U3898 , P2_R1200_U89 );
nand NAND2_15449 ( P2_R1200_U296 , P2_R1200_U295 , P2_R1200_U168 );
nand NAND2_15450 ( P2_R1200_U297 , P2_U3057 , P2_R1200_U88 );
not NOT1_15451 ( P2_R1200_U298 , P2_R1200_U93 );
nand NAND2_15452 ( P2_R1200_U299 , P2_U3896 , P2_R1200_U54 );
nand NAND2_15453 ( P2_R1200_U300 , P2_R1200_U54 , P2_R1200_U53 );
nand NAND2_15454 ( P2_R1200_U301 , P2_R1200_U300 , P2_R1200_U91 );
nand NAND2_15455 ( P2_R1200_U302 , P2_U3052 , P2_R1200_U189 );
nand NAND2_15456 ( P2_R1200_U303 , P2_U3895 , P2_R1200_U92 );
nand NAND2_15457 ( P2_R1200_U304 , P2_U3053 , P2_R1200_U51 );
nand NAND2_15458 ( P2_R1200_U305 , P2_R1200_U140 , P2_R1200_U355 );
nand NAND2_15459 ( P2_R1200_U306 , P2_R1200_U53 , P2_R1200_U195 );
nand NAND2_15460 ( P2_R1200_U307 , P2_R1200_U286 , P2_R1200_U172 );
not NOT1_15461 ( P2_R1200_U308 , P2_R1200_U94 );
nand NAND2_15462 ( P2_R1200_U309 , P2_U3060 , P2_R1200_U80 );
nand NAND2_15463 ( P2_R1200_U310 , P2_R1200_U308 , P2_R1200_U309 );
nand NAND2_15464 ( P2_R1200_U311 , P2_R1200_U144 , P2_R1200_U310 );
nand NAND2_15465 ( P2_R1200_U312 , P2_R1200_U94 , P2_R1200_U194 );
nand NAND2_15466 ( P2_R1200_U313 , P2_U3900 , P2_R1200_U82 );
nand NAND2_15467 ( P2_R1200_U314 , P2_R1200_U143 , P2_R1200_U312 );
nand NAND2_15468 ( P2_R1200_U315 , P2_U3060 , P2_R1200_U80 );
nand NAND2_15469 ( P2_R1200_U316 , P2_R1200_U194 , P2_R1200_U315 );
nand NAND2_15470 ( P2_R1200_U317 , P2_R1200_U286 , P2_R1200_U85 );
nand NAND2_15471 ( P2_R1200_U318 , P2_R1200_U262 , P2_R1200_U182 );
not NOT1_15472 ( P2_R1200_U319 , P2_R1200_U95 );
nand NAND2_15473 ( P2_R1200_U320 , P2_U3073 , P2_R1200_U66 );
nand NAND2_15474 ( P2_R1200_U321 , P2_R1200_U319 , P2_R1200_U320 );
nand NAND2_15475 ( P2_R1200_U322 , P2_R1200_U151 , P2_R1200_U321 );
nand NAND2_15476 ( P2_R1200_U323 , P2_R1200_U95 , P2_R1200_U193 );
nand NAND2_15477 ( P2_R1200_U324 , P2_U3437 , P2_R1200_U68 );
nand NAND2_15478 ( P2_R1200_U325 , P2_R1200_U150 , P2_R1200_U323 );
nand NAND2_15479 ( P2_R1200_U326 , P2_U3073 , P2_R1200_U66 );
nand NAND2_15480 ( P2_R1200_U327 , P2_R1200_U193 , P2_R1200_U326 );
nand NAND2_15481 ( P2_R1200_U328 , P2_R1200_U262 , P2_R1200_U71 );
nand NAND2_15482 ( P2_R1200_U329 , P2_U3061 , P2_R1200_U58 );
nand NAND2_15483 ( P2_R1200_U330 , P2_R1200_U350 , P2_R1200_U329 );
nand NAND2_15484 ( P2_R1200_U331 , P2_R1200_U155 , P2_R1200_U330 );
nand NAND2_15485 ( P2_R1200_U332 , P2_R1200_U96 , P2_R1200_U192 );
nand NAND2_15486 ( P2_R1200_U333 , P2_U3422 , P2_R1200_U56 );
nand NAND2_15487 ( P2_R1200_U334 , P2_R1200_U154 , P2_R1200_U332 );
nand NAND2_15488 ( P2_R1200_U335 , P2_U3061 , P2_R1200_U58 );
nand NAND2_15489 ( P2_R1200_U336 , P2_R1200_U192 , P2_R1200_U335 );
nand NAND2_15490 ( P2_R1200_U337 , P2_U3076 , P2_R1200_U38 );
nand NAND2_15491 ( P2_R1200_U338 , P2_U3077 , P2_R1200_U174 );
nand NAND2_15492 ( P2_R1200_U339 , P2_U3081 , P2_R1200_U177 );
nand NAND2_15493 ( P2_R1200_U340 , P2_R1200_U33 , P2_R1200_U221 );
nand NAND2_15494 ( P2_R1200_U341 , P2_R1200_U121 , P2_R1200_U161 );
nand NAND2_15495 ( P2_R1200_U342 , P2_R1200_U218 , P2_R1200_U14 );
nand NAND2_15496 ( P2_R1200_U343 , P2_R1200_U250 , P2_R1200_U251 );
nand NAND2_15497 ( P2_R1200_U344 , P2_R1200_U119 , P2_R1200_U50 );
not NOT1_15498 ( P2_R1200_U345 , P2_R1200_U161 );
nand NAND2_15499 ( P2_R1200_U346 , P2_R1200_U196 , P2_R1200_U50 );
nand NAND2_15500 ( P2_R1200_U347 , P2_R1200_U128 , P2_R1200_U346 );
nand NAND2_15501 ( P2_R1200_U348 , P2_R1200_U205 , P2_R1200_U35 );
nand NAND2_15502 ( P2_R1200_U349 , P2_R1200_U224 , P2_R1200_U157 );
not NOT1_15503 ( P2_R1200_U350 , P2_R1200_U96 );
nand NAND2_15504 ( P2_R1200_U351 , P2_R1200_U15 , P2_R1200_U157 );
not NOT1_15505 ( P2_R1200_U352 , P2_R1200_U184 );
nand NAND2_15506 ( P2_R1200_U353 , P2_R1200_U130 , P2_R1200_U157 );
not NOT1_15507 ( P2_R1200_U354 , P2_R1200_U183 );
nand NAND2_15508 ( P2_R1200_U355 , P2_R1200_U298 , P2_R1200_U53 );
nand NAND2_15509 ( P2_R1200_U356 , P2_R1200_U195 , P2_R1200_U93 );
nand NAND2_15510 ( P2_R1200_U357 , P2_R1200_U139 , P2_R1200_U356 );
nand NAND2_15511 ( P2_R1200_U358 , P2_R1200_U12 , P2_R1200_U93 );
nand NAND2_15512 ( P2_R1200_U359 , P2_R1200_U136 , P2_R1200_U358 );
nand NAND2_15513 ( P2_R1200_U360 , P2_R1200_U12 , P2_R1200_U93 );
not NOT1_15514 ( P2_R1200_U361 , P2_R1200_U166 );
nand NAND2_15515 ( P2_R1200_U362 , P2_U3416 , P2_R1200_U47 );
nand NAND2_15516 ( P2_R1200_U363 , P2_U3082 , P2_R1200_U46 );
nand NAND2_15517 ( P2_R1200_U364 , P2_R1200_U225 , P2_R1200_U157 );
nand NAND2_15518 ( P2_R1200_U365 , P2_R1200_U223 , P2_R1200_U156 );
nand NAND2_15519 ( P2_R1200_U366 , P2_U3413 , P2_R1200_U28 );
nand NAND2_15520 ( P2_R1200_U367 , P2_U3083 , P2_R1200_U33 );
nand NAND2_15521 ( P2_R1200_U368 , P2_U3413 , P2_R1200_U28 );
nand NAND2_15522 ( P2_R1200_U369 , P2_U3083 , P2_R1200_U33 );
nand NAND2_15523 ( P2_R1200_U370 , P2_R1200_U369 , P2_R1200_U368 );
nand NAND2_15524 ( P2_R1200_U371 , P2_U3410 , P2_R1200_U26 );
nand NAND2_15525 ( P2_R1200_U372 , P2_U3069 , P2_R1200_U32 );
nand NAND2_15526 ( P2_R1200_U373 , P2_R1200_U230 , P2_R1200_U48 );
nand NAND2_15527 ( P2_R1200_U374 , P2_R1200_U158 , P2_R1200_U219 );
nand NAND2_15528 ( P2_R1200_U375 , P2_U3407 , P2_R1200_U41 );
nand NAND2_15529 ( P2_R1200_U376 , P2_U3070 , P2_R1200_U30 );
nand NAND2_15530 ( P2_R1200_U377 , P2_R1200_U376 , P2_R1200_U375 );
nand NAND2_15531 ( P2_R1200_U378 , P2_U3404 , P2_R1200_U42 );
nand NAND2_15532 ( P2_R1200_U379 , P2_U3066 , P2_R1200_U29 );
nand NAND2_15533 ( P2_R1200_U380 , P2_R1200_U240 , P2_R1200_U49 );
nand NAND2_15534 ( P2_R1200_U381 , P2_R1200_U159 , P2_R1200_U232 );
nand NAND2_15535 ( P2_R1200_U382 , P2_U3401 , P2_R1200_U43 );
nand NAND2_15536 ( P2_R1200_U383 , P2_U3059 , P2_R1200_U31 );
nand NAND2_15537 ( P2_R1200_U384 , P2_R1200_U161 , P2_R1200_U241 );
nand NAND2_15538 ( P2_R1200_U385 , P2_R1200_U345 , P2_R1200_U160 );
nand NAND2_15539 ( P2_R1200_U386 , P2_U3398 , P2_R1200_U36 );
nand NAND2_15540 ( P2_R1200_U387 , P2_U3063 , P2_R1200_U40 );
nand NAND2_15541 ( P2_R1200_U388 , P2_U3398 , P2_R1200_U36 );
nand NAND2_15542 ( P2_R1200_U389 , P2_U3063 , P2_R1200_U40 );
nand NAND2_15543 ( P2_R1200_U390 , P2_R1200_U389 , P2_R1200_U388 );
nand NAND2_15544 ( P2_R1200_U391 , P2_U3395 , P2_R1200_U34 );
nand NAND2_15545 ( P2_R1200_U392 , P2_U3067 , P2_R1200_U37 );
nand NAND2_15546 ( P2_R1200_U393 , P2_R1200_U243 , P2_R1200_U50 );
nand NAND2_15547 ( P2_R1200_U394 , P2_R1200_U162 , P2_R1200_U205 );
nand NAND2_15548 ( P2_R1200_U395 , P2_U3904 , P2_R1200_U164 );
nand NAND2_15549 ( P2_R1200_U396 , P2_U3054 , P2_R1200_U163 );
nand NAND2_15550 ( P2_R1200_U397 , P2_R1200_U396 , P2_R1200_U395 );
nand NAND2_15551 ( P2_R1200_U398 , P2_U3904 , P2_R1200_U164 );
nand NAND2_15552 ( P2_R1200_U399 , P2_U3054 , P2_R1200_U163 );
nand NAND3_15553 ( P2_R1200_U400 , P2_U3053 , P2_R1200_U397 , P2_R1200_U51 );
nand NAND3_15554 ( P2_R1200_U401 , P2_R1200_U16 , P2_R1200_U92 , P2_U3895 );
nand NAND2_15555 ( P2_R1200_U402 , P2_U3895 , P2_R1200_U92 );
nand NAND2_15556 ( P2_R1200_U403 , P2_U3053 , P2_R1200_U51 );
not NOT1_15557 ( P2_R1200_U404 , P2_R1200_U138 );
nand NAND2_15558 ( P2_R1200_U405 , P2_R1200_U361 , P2_R1200_U404 );
nand NAND2_15559 ( P2_R1200_U406 , P2_R1200_U138 , P2_R1200_U166 );
nand NAND2_15560 ( P2_R1200_U407 , P2_U3896 , P2_R1200_U54 );
nand NAND2_15561 ( P2_R1200_U408 , P2_U3052 , P2_R1200_U91 );
nand NAND2_15562 ( P2_R1200_U409 , P2_U3896 , P2_R1200_U54 );
nand NAND2_15563 ( P2_R1200_U410 , P2_U3052 , P2_R1200_U91 );
nand NAND2_15564 ( P2_R1200_U411 , P2_R1200_U410 , P2_R1200_U409 );
nand NAND2_15565 ( P2_R1200_U412 , P2_U3897 , P2_R1200_U52 );
nand NAND2_15566 ( P2_R1200_U413 , P2_U3056 , P2_R1200_U90 );
nand NAND2_15567 ( P2_R1200_U414 , P2_R1200_U306 , P2_R1200_U93 );
nand NAND2_15568 ( P2_R1200_U415 , P2_R1200_U167 , P2_R1200_U298 );
nand NAND2_15569 ( P2_R1200_U416 , P2_U3898 , P2_R1200_U89 );
nand NAND2_15570 ( P2_R1200_U417 , P2_U3057 , P2_R1200_U88 );
not NOT1_15571 ( P2_R1200_U418 , P2_R1200_U141 );
nand NAND2_15572 ( P2_R1200_U419 , P2_R1200_U294 , P2_R1200_U418 );
nand NAND2_15573 ( P2_R1200_U420 , P2_R1200_U141 , P2_R1200_U168 );
nand NAND2_15574 ( P2_R1200_U421 , P2_U3899 , P2_R1200_U87 );
nand NAND2_15575 ( P2_R1200_U422 , P2_U3064 , P2_R1200_U86 );
not NOT1_15576 ( P2_R1200_U423 , P2_R1200_U142 );
nand NAND2_15577 ( P2_R1200_U424 , P2_R1200_U290 , P2_R1200_U423 );
nand NAND2_15578 ( P2_R1200_U425 , P2_R1200_U142 , P2_R1200_U169 );
nand NAND2_15579 ( P2_R1200_U426 , P2_U3900 , P2_R1200_U82 );
nand NAND2_15580 ( P2_R1200_U427 , P2_U3065 , P2_R1200_U79 );
nand NAND2_15581 ( P2_R1200_U428 , P2_R1200_U427 , P2_R1200_U426 );
nand NAND2_15582 ( P2_R1200_U429 , P2_U3901 , P2_R1200_U83 );
nand NAND2_15583 ( P2_R1200_U430 , P2_U3060 , P2_R1200_U80 );
nand NAND2_15584 ( P2_R1200_U431 , P2_R1200_U316 , P2_R1200_U94 );
nand NAND2_15585 ( P2_R1200_U432 , P2_R1200_U170 , P2_R1200_U308 );
nand NAND2_15586 ( P2_R1200_U433 , P2_U3902 , P2_R1200_U84 );
nand NAND2_15587 ( P2_R1200_U434 , P2_U3074 , P2_R1200_U81 );
nand NAND2_15588 ( P2_R1200_U435 , P2_R1200_U317 , P2_R1200_U172 );
nand NAND2_15589 ( P2_R1200_U436 , P2_R1200_U280 , P2_R1200_U171 );
nand NAND2_15590 ( P2_R1200_U437 , P2_U3903 , P2_R1200_U78 );
nand NAND2_15591 ( P2_R1200_U438 , P2_U3075 , P2_R1200_U77 );
not NOT1_15592 ( P2_R1200_U439 , P2_R1200_U145 );
nand NAND2_15593 ( P2_R1200_U440 , P2_R1200_U276 , P2_R1200_U439 );
nand NAND2_15594 ( P2_R1200_U441 , P2_R1200_U145 , P2_R1200_U173 );
nand NAND2_15595 ( P2_R1200_U442 , P2_U3392 , P2_R1200_U39 );
nand NAND2_15596 ( P2_R1200_U443 , P2_U3077 , P2_R1200_U174 );
not NOT1_15597 ( P2_R1200_U444 , P2_R1200_U146 );
nand NAND2_15598 ( P2_R1200_U445 , P2_R1200_U203 , P2_R1200_U444 );
nand NAND2_15599 ( P2_R1200_U446 , P2_R1200_U146 , P2_R1200_U175 );
nand NAND2_15600 ( P2_R1200_U447 , P2_U3445 , P2_R1200_U76 );
nand NAND2_15601 ( P2_R1200_U448 , P2_U3080 , P2_R1200_U75 );
not NOT1_15602 ( P2_R1200_U449 , P2_R1200_U147 );
nand NAND2_15603 ( P2_R1200_U450 , P2_R1200_U272 , P2_R1200_U449 );
nand NAND2_15604 ( P2_R1200_U451 , P2_R1200_U147 , P2_R1200_U176 );
nand NAND2_15605 ( P2_R1200_U452 , P2_U3443 , P2_R1200_U74 );
nand NAND2_15606 ( P2_R1200_U453 , P2_U3081 , P2_R1200_U177 );
not NOT1_15607 ( P2_R1200_U454 , P2_R1200_U148 );
nand NAND2_15608 ( P2_R1200_U455 , P2_R1200_U270 , P2_R1200_U454 );
nand NAND2_15609 ( P2_R1200_U456 , P2_R1200_U148 , P2_R1200_U178 );
nand NAND2_15610 ( P2_R1200_U457 , P2_U3440 , P2_R1200_U73 );
nand NAND2_15611 ( P2_R1200_U458 , P2_U3068 , P2_R1200_U72 );
not NOT1_15612 ( P2_R1200_U459 , P2_R1200_U149 );
nand NAND2_15613 ( P2_R1200_U460 , P2_R1200_U266 , P2_R1200_U459 );
nand NAND2_15614 ( P2_R1200_U461 , P2_R1200_U149 , P2_R1200_U179 );
nand NAND2_15615 ( P2_R1200_U462 , P2_U3437 , P2_R1200_U68 );
nand NAND2_15616 ( P2_R1200_U463 , P2_U3072 , P2_R1200_U65 );
nand NAND2_15617 ( P2_R1200_U464 , P2_R1200_U463 , P2_R1200_U462 );
nand NAND2_15618 ( P2_R1200_U465 , P2_U3434 , P2_R1200_U69 );
nand NAND2_15619 ( P2_R1200_U466 , P2_U3073 , P2_R1200_U66 );
nand NAND2_15620 ( P2_R1200_U467 , P2_R1200_U327 , P2_R1200_U95 );
nand NAND2_15621 ( P2_R1200_U468 , P2_R1200_U180 , P2_R1200_U319 );
nand NAND2_15622 ( P2_R1200_U469 , P2_U3431 , P2_R1200_U70 );
nand NAND2_15623 ( P2_R1200_U470 , P2_U3078 , P2_R1200_U67 );
nand NAND2_15624 ( P2_R1200_U471 , P2_R1200_U328 , P2_R1200_U182 );
nand NAND2_15625 ( P2_R1200_U472 , P2_R1200_U256 , P2_R1200_U181 );
nand NAND2_15626 ( P2_R1200_U473 , P2_U3428 , P2_R1200_U64 );
nand NAND2_15627 ( P2_R1200_U474 , P2_U3079 , P2_R1200_U63 );
not NOT1_15628 ( P2_R1200_U475 , P2_R1200_U152 );
nand NAND2_15629 ( P2_R1200_U476 , P2_R1200_U354 , P2_R1200_U475 );
nand NAND2_15630 ( P2_R1200_U477 , P2_R1200_U152 , P2_R1200_U183 );
nand NAND2_15631 ( P2_R1200_U478 , P2_U3425 , P2_R1200_U55 );
nand NAND2_15632 ( P2_R1200_U479 , P2_U3071 , P2_R1200_U61 );
not NOT1_15633 ( P2_R1200_U480 , P2_R1200_U153 );
nand NAND2_15634 ( P2_R1200_U481 , P2_R1200_U352 , P2_R1200_U480 );
nand NAND2_15635 ( P2_R1200_U482 , P2_R1200_U153 , P2_R1200_U184 );
nand NAND2_15636 ( P2_R1200_U483 , P2_U3422 , P2_R1200_U56 );
nand NAND2_15637 ( P2_R1200_U484 , P2_U3062 , P2_R1200_U60 );
nand NAND2_15638 ( P2_R1200_U485 , P2_R1200_U484 , P2_R1200_U483 );
nand NAND2_15639 ( P2_R1200_U486 , P2_U3419 , P2_R1200_U57 );
nand NAND2_15640 ( P2_R1200_U487 , P2_U3061 , P2_R1200_U58 );
nand NAND2_15641 ( P2_R1200_U488 , P2_R1200_U96 , P2_R1200_U336 );
nand NAND2_15642 ( P2_R1200_U489 , P2_R1200_U185 , P2_R1200_U350 );
and AND2_15643 ( P2_R1179_U6 , P2_R1179_U212 , P2_R1179_U211 );
and AND2_15644 ( P2_R1179_U7 , P2_R1179_U246 , P2_R1179_U245 );
and AND2_15645 ( P2_R1179_U8 , P2_R1179_U193 , P2_R1179_U257 );
and AND2_15646 ( P2_R1179_U9 , P2_R1179_U259 , P2_R1179_U258 );
and AND2_15647 ( P2_R1179_U10 , P2_R1179_U194 , P2_R1179_U281 );
and AND2_15648 ( P2_R1179_U11 , P2_R1179_U283 , P2_R1179_U282 );
and AND2_15649 ( P2_R1179_U12 , P2_R1179_U299 , P2_R1179_U195 );
and AND3_15650 ( P2_R1179_U13 , P2_R1179_U210 , P2_R1179_U197 , P2_R1179_U215 );
and AND2_15651 ( P2_R1179_U14 , P2_R1179_U220 , P2_R1179_U198 );
and AND3_15652 ( P2_R1179_U15 , P2_R1179_U224 , P2_R1179_U192 , P2_R1179_U244 );
and AND2_15653 ( P2_R1179_U16 , P2_R1179_U399 , P2_R1179_U398 );
nand NAND2_15654 ( P2_R1179_U17 , P2_R1179_U331 , P2_R1179_U334 );
nand NAND2_15655 ( P2_R1179_U18 , P2_R1179_U322 , P2_R1179_U325 );
nand NAND2_15656 ( P2_R1179_U19 , P2_R1179_U311 , P2_R1179_U314 );
nand NAND2_15657 ( P2_R1179_U20 , P2_R1179_U305 , P2_R1179_U357 );
nand NAND2_15658 ( P2_R1179_U21 , P2_R1179_U137 , P2_R1179_U186 );
nand NAND2_15659 ( P2_R1179_U22 , P2_R1179_U242 , P2_R1179_U347 );
nand NAND2_15660 ( P2_R1179_U23 , P2_R1179_U235 , P2_R1179_U238 );
nand NAND2_15661 ( P2_R1179_U24 , P2_R1179_U227 , P2_R1179_U229 );
nand NAND2_15662 ( P2_R1179_U25 , P2_R1179_U175 , P2_R1179_U337 );
not NOT1_15663 ( P2_R1179_U26 , P2_U3069 );
nand NAND2_15664 ( P2_R1179_U27 , P2_U3069 , P2_R1179_U32 );
not NOT1_15665 ( P2_R1179_U28 , P2_U3083 );
not NOT1_15666 ( P2_R1179_U29 , P2_U3404 );
not NOT1_15667 ( P2_R1179_U30 , P2_U3407 );
not NOT1_15668 ( P2_R1179_U31 , P2_U3401 );
not NOT1_15669 ( P2_R1179_U32 , P2_U3410 );
not NOT1_15670 ( P2_R1179_U33 , P2_U3413 );
not NOT1_15671 ( P2_R1179_U34 , P2_U3067 );
nand NAND2_15672 ( P2_R1179_U35 , P2_U3067 , P2_R1179_U37 );
not NOT1_15673 ( P2_R1179_U36 , P2_U3063 );
not NOT1_15674 ( P2_R1179_U37 , P2_U3395 );
not NOT1_15675 ( P2_R1179_U38 , P2_U3387 );
not NOT1_15676 ( P2_R1179_U39 , P2_U3077 );
not NOT1_15677 ( P2_R1179_U40 , P2_U3398 );
not NOT1_15678 ( P2_R1179_U41 , P2_U3070 );
not NOT1_15679 ( P2_R1179_U42 , P2_U3066 );
not NOT1_15680 ( P2_R1179_U43 , P2_U3059 );
nand NAND2_15681 ( P2_R1179_U44 , P2_U3059 , P2_R1179_U31 );
nand NAND2_15682 ( P2_R1179_U45 , P2_R1179_U216 , P2_R1179_U214 );
not NOT1_15683 ( P2_R1179_U46 , P2_U3416 );
not NOT1_15684 ( P2_R1179_U47 , P2_U3082 );
nand NAND2_15685 ( P2_R1179_U48 , P2_R1179_U45 , P2_R1179_U217 );
nand NAND2_15686 ( P2_R1179_U49 , P2_R1179_U44 , P2_R1179_U231 );
nand NAND3_15687 ( P2_R1179_U50 , P2_R1179_U204 , P2_R1179_U188 , P2_R1179_U338 );
not NOT1_15688 ( P2_R1179_U51 , P2_U3895 );
not NOT1_15689 ( P2_R1179_U52 , P2_U3056 );
nand NAND2_15690 ( P2_R1179_U53 , P2_U3056 , P2_R1179_U90 );
not NOT1_15691 ( P2_R1179_U54 , P2_U3052 );
not NOT1_15692 ( P2_R1179_U55 , P2_U3071 );
not NOT1_15693 ( P2_R1179_U56 , P2_U3062 );
not NOT1_15694 ( P2_R1179_U57 , P2_U3061 );
not NOT1_15695 ( P2_R1179_U58 , P2_U3419 );
nand NAND2_15696 ( P2_R1179_U59 , P2_U3082 , P2_R1179_U46 );
not NOT1_15697 ( P2_R1179_U60 , P2_U3422 );
not NOT1_15698 ( P2_R1179_U61 , P2_U3425 );
nand NAND2_15699 ( P2_R1179_U62 , P2_R1179_U249 , P2_R1179_U248 );
not NOT1_15700 ( P2_R1179_U63 , P2_U3428 );
not NOT1_15701 ( P2_R1179_U64 , P2_U3079 );
not NOT1_15702 ( P2_R1179_U65 , P2_U3437 );
not NOT1_15703 ( P2_R1179_U66 , P2_U3434 );
not NOT1_15704 ( P2_R1179_U67 , P2_U3431 );
not NOT1_15705 ( P2_R1179_U68 , P2_U3072 );
not NOT1_15706 ( P2_R1179_U69 , P2_U3073 );
not NOT1_15707 ( P2_R1179_U70 , P2_U3078 );
nand NAND2_15708 ( P2_R1179_U71 , P2_U3078 , P2_R1179_U67 );
not NOT1_15709 ( P2_R1179_U72 , P2_U3440 );
not NOT1_15710 ( P2_R1179_U73 , P2_U3068 );
not NOT1_15711 ( P2_R1179_U74 , P2_U3081 );
not NOT1_15712 ( P2_R1179_U75 , P2_U3445 );
not NOT1_15713 ( P2_R1179_U76 , P2_U3080 );
not NOT1_15714 ( P2_R1179_U77 , P2_U3903 );
not NOT1_15715 ( P2_R1179_U78 , P2_U3075 );
not NOT1_15716 ( P2_R1179_U79 , P2_U3900 );
not NOT1_15717 ( P2_R1179_U80 , P2_U3901 );
not NOT1_15718 ( P2_R1179_U81 , P2_U3902 );
not NOT1_15719 ( P2_R1179_U82 , P2_U3065 );
not NOT1_15720 ( P2_R1179_U83 , P2_U3060 );
not NOT1_15721 ( P2_R1179_U84 , P2_U3074 );
nand NAND2_15722 ( P2_R1179_U85 , P2_U3074 , P2_R1179_U81 );
not NOT1_15723 ( P2_R1179_U86 , P2_U3899 );
not NOT1_15724 ( P2_R1179_U87 , P2_U3064 );
not NOT1_15725 ( P2_R1179_U88 , P2_U3898 );
not NOT1_15726 ( P2_R1179_U89 , P2_U3057 );
not NOT1_15727 ( P2_R1179_U90 , P2_U3897 );
not NOT1_15728 ( P2_R1179_U91 , P2_U3896 );
not NOT1_15729 ( P2_R1179_U92 , P2_U3053 );
nand NAND2_15730 ( P2_R1179_U93 , P2_R1179_U297 , P2_R1179_U296 );
nand NAND2_15731 ( P2_R1179_U94 , P2_R1179_U85 , P2_R1179_U307 );
nand NAND2_15732 ( P2_R1179_U95 , P2_R1179_U71 , P2_R1179_U318 );
nand NAND2_15733 ( P2_R1179_U96 , P2_R1179_U349 , P2_R1179_U59 );
not NOT1_15734 ( P2_R1179_U97 , P2_U3076 );
nand NAND2_15735 ( P2_R1179_U98 , P2_R1179_U406 , P2_R1179_U405 );
nand NAND2_15736 ( P2_R1179_U99 , P2_R1179_U420 , P2_R1179_U419 );
nand NAND2_15737 ( P2_R1179_U100 , P2_R1179_U425 , P2_R1179_U424 );
nand NAND2_15738 ( P2_R1179_U101 , P2_R1179_U441 , P2_R1179_U440 );
nand NAND2_15739 ( P2_R1179_U102 , P2_R1179_U446 , P2_R1179_U445 );
nand NAND2_15740 ( P2_R1179_U103 , P2_R1179_U451 , P2_R1179_U450 );
nand NAND2_15741 ( P2_R1179_U104 , P2_R1179_U456 , P2_R1179_U455 );
nand NAND2_15742 ( P2_R1179_U105 , P2_R1179_U461 , P2_R1179_U460 );
nand NAND2_15743 ( P2_R1179_U106 , P2_R1179_U477 , P2_R1179_U476 );
nand NAND2_15744 ( P2_R1179_U107 , P2_R1179_U482 , P2_R1179_U481 );
nand NAND2_15745 ( P2_R1179_U108 , P2_R1179_U365 , P2_R1179_U364 );
nand NAND2_15746 ( P2_R1179_U109 , P2_R1179_U374 , P2_R1179_U373 );
nand NAND2_15747 ( P2_R1179_U110 , P2_R1179_U381 , P2_R1179_U380 );
nand NAND2_15748 ( P2_R1179_U111 , P2_R1179_U385 , P2_R1179_U384 );
nand NAND2_15749 ( P2_R1179_U112 , P2_R1179_U394 , P2_R1179_U393 );
nand NAND2_15750 ( P2_R1179_U113 , P2_R1179_U415 , P2_R1179_U414 );
nand NAND2_15751 ( P2_R1179_U114 , P2_R1179_U432 , P2_R1179_U431 );
nand NAND2_15752 ( P2_R1179_U115 , P2_R1179_U436 , P2_R1179_U435 );
nand NAND2_15753 ( P2_R1179_U116 , P2_R1179_U468 , P2_R1179_U467 );
nand NAND2_15754 ( P2_R1179_U117 , P2_R1179_U472 , P2_R1179_U471 );
nand NAND2_15755 ( P2_R1179_U118 , P2_R1179_U489 , P2_R1179_U488 );
and AND2_15756 ( P2_R1179_U119 , P2_R1179_U206 , P2_R1179_U196 );
and AND2_15757 ( P2_R1179_U120 , P2_R1179_U209 , P2_R1179_U208 );
and AND2_15758 ( P2_R1179_U121 , P2_R1179_U14 , P2_R1179_U13 );
and AND2_15759 ( P2_R1179_U122 , P2_R1179_U340 , P2_R1179_U222 );
and AND2_15760 ( P2_R1179_U123 , P2_R1179_U342 , P2_R1179_U122 );
and AND3_15761 ( P2_R1179_U124 , P2_R1179_U367 , P2_R1179_U366 , P2_R1179_U27 );
and AND2_15762 ( P2_R1179_U125 , P2_R1179_U370 , P2_R1179_U198 );
and AND2_15763 ( P2_R1179_U126 , P2_R1179_U237 , P2_R1179_U6 );
and AND2_15764 ( P2_R1179_U127 , P2_R1179_U377 , P2_R1179_U197 );
and AND3_15765 ( P2_R1179_U128 , P2_R1179_U387 , P2_R1179_U386 , P2_R1179_U35 );
and AND2_15766 ( P2_R1179_U129 , P2_R1179_U390 , P2_R1179_U196 );
and AND2_15767 ( P2_R1179_U130 , P2_R1179_U251 , P2_R1179_U15 );
and AND2_15768 ( P2_R1179_U131 , P2_R1179_U343 , P2_R1179_U252 );
and AND2_15769 ( P2_R1179_U132 , P2_R1179_U262 , P2_R1179_U8 );
and AND2_15770 ( P2_R1179_U133 , P2_R1179_U286 , P2_R1179_U10 );
and AND2_15771 ( P2_R1179_U134 , P2_R1179_U302 , P2_R1179_U301 );
and AND2_15772 ( P2_R1179_U135 , P2_R1179_U397 , P2_R1179_U303 );
and AND4_15773 ( P2_R1179_U136 , P2_R1179_U302 , P2_R1179_U301 , P2_R1179_U304 , P2_R1179_U16 );
and AND2_15774 ( P2_R1179_U137 , P2_R1179_U359 , P2_R1179_U165 );
nand NAND2_15775 ( P2_R1179_U138 , P2_R1179_U403 , P2_R1179_U402 );
and AND3_15776 ( P2_R1179_U139 , P2_R1179_U408 , P2_R1179_U407 , P2_R1179_U53 );
and AND2_15777 ( P2_R1179_U140 , P2_R1179_U411 , P2_R1179_U195 );
nand NAND2_15778 ( P2_R1179_U141 , P2_R1179_U417 , P2_R1179_U416 );
nand NAND2_15779 ( P2_R1179_U142 , P2_R1179_U422 , P2_R1179_U421 );
and AND2_15780 ( P2_R1179_U143 , P2_R1179_U313 , P2_R1179_U11 );
and AND2_15781 ( P2_R1179_U144 , P2_R1179_U428 , P2_R1179_U194 );
nand NAND2_15782 ( P2_R1179_U145 , P2_R1179_U438 , P2_R1179_U437 );
nand NAND2_15783 ( P2_R1179_U146 , P2_R1179_U443 , P2_R1179_U442 );
nand NAND2_15784 ( P2_R1179_U147 , P2_R1179_U448 , P2_R1179_U447 );
nand NAND2_15785 ( P2_R1179_U148 , P2_R1179_U453 , P2_R1179_U452 );
nand NAND2_15786 ( P2_R1179_U149 , P2_R1179_U458 , P2_R1179_U457 );
and AND2_15787 ( P2_R1179_U150 , P2_R1179_U324 , P2_R1179_U9 );
and AND2_15788 ( P2_R1179_U151 , P2_R1179_U464 , P2_R1179_U193 );
nand NAND2_15789 ( P2_R1179_U152 , P2_R1179_U474 , P2_R1179_U473 );
nand NAND2_15790 ( P2_R1179_U153 , P2_R1179_U479 , P2_R1179_U478 );
and AND2_15791 ( P2_R1179_U154 , P2_R1179_U333 , P2_R1179_U7 );
and AND2_15792 ( P2_R1179_U155 , P2_R1179_U485 , P2_R1179_U192 );
and AND2_15793 ( P2_R1179_U156 , P2_R1179_U363 , P2_R1179_U362 );
nand NAND2_15794 ( P2_R1179_U157 , P2_R1179_U123 , P2_R1179_U341 );
and AND2_15795 ( P2_R1179_U158 , P2_R1179_U372 , P2_R1179_U371 );
and AND2_15796 ( P2_R1179_U159 , P2_R1179_U379 , P2_R1179_U378 );
and AND2_15797 ( P2_R1179_U160 , P2_R1179_U383 , P2_R1179_U382 );
nand NAND2_15798 ( P2_R1179_U161 , P2_R1179_U120 , P2_R1179_U344 );
and AND2_15799 ( P2_R1179_U162 , P2_R1179_U392 , P2_R1179_U391 );
not NOT1_15800 ( P2_R1179_U163 , P2_U3904 );
not NOT1_15801 ( P2_R1179_U164 , P2_U3054 );
and AND2_15802 ( P2_R1179_U165 , P2_R1179_U401 , P2_R1179_U400 );
nand NAND2_15803 ( P2_R1179_U166 , P2_R1179_U134 , P2_R1179_U360 );
and AND2_15804 ( P2_R1179_U167 , P2_R1179_U413 , P2_R1179_U412 );
nand NAND2_15805 ( P2_R1179_U168 , P2_R1179_U293 , P2_R1179_U292 );
nand NAND2_15806 ( P2_R1179_U169 , P2_R1179_U289 , P2_R1179_U288 );
and AND2_15807 ( P2_R1179_U170 , P2_R1179_U430 , P2_R1179_U429 );
and AND2_15808 ( P2_R1179_U171 , P2_R1179_U434 , P2_R1179_U433 );
nand NAND2_15809 ( P2_R1179_U172 , P2_R1179_U279 , P2_R1179_U278 );
nand NAND2_15810 ( P2_R1179_U173 , P2_R1179_U275 , P2_R1179_U274 );
not NOT1_15811 ( P2_R1179_U174 , P2_U3392 );
nand NAND2_15812 ( P2_R1179_U175 , P2_U3387 , P2_R1179_U97 );
nand NAND3_15813 ( P2_R1179_U176 , P2_R1179_U271 , P2_R1179_U187 , P2_R1179_U339 );
not NOT1_15814 ( P2_R1179_U177 , P2_U3443 );
nand NAND2_15815 ( P2_R1179_U178 , P2_R1179_U269 , P2_R1179_U268 );
nand NAND2_15816 ( P2_R1179_U179 , P2_R1179_U265 , P2_R1179_U264 );
and AND2_15817 ( P2_R1179_U180 , P2_R1179_U466 , P2_R1179_U465 );
and AND2_15818 ( P2_R1179_U181 , P2_R1179_U470 , P2_R1179_U469 );
nand NAND2_15819 ( P2_R1179_U182 , P2_R1179_U255 , P2_R1179_U254 );
nand NAND2_15820 ( P2_R1179_U183 , P2_R1179_U131 , P2_R1179_U353 );
nand NAND2_15821 ( P2_R1179_U184 , P2_R1179_U351 , P2_R1179_U62 );
and AND2_15822 ( P2_R1179_U185 , P2_R1179_U487 , P2_R1179_U486 );
nand NAND2_15823 ( P2_R1179_U186 , P2_R1179_U135 , P2_R1179_U166 );
nand NAND2_15824 ( P2_R1179_U187 , P2_R1179_U178 , P2_R1179_U177 );
nand NAND2_15825 ( P2_R1179_U188 , P2_R1179_U175 , P2_R1179_U174 );
not NOT1_15826 ( P2_R1179_U189 , P2_R1179_U53 );
not NOT1_15827 ( P2_R1179_U190 , P2_R1179_U35 );
not NOT1_15828 ( P2_R1179_U191 , P2_R1179_U27 );
nand NAND2_15829 ( P2_R1179_U192 , P2_U3419 , P2_R1179_U57 );
nand NAND2_15830 ( P2_R1179_U193 , P2_U3434 , P2_R1179_U69 );
nand NAND2_15831 ( P2_R1179_U194 , P2_U3901 , P2_R1179_U83 );
nand NAND2_15832 ( P2_R1179_U195 , P2_U3897 , P2_R1179_U52 );
nand NAND2_15833 ( P2_R1179_U196 , P2_U3395 , P2_R1179_U34 );
nand NAND2_15834 ( P2_R1179_U197 , P2_U3404 , P2_R1179_U42 );
nand NAND2_15835 ( P2_R1179_U198 , P2_U3410 , P2_R1179_U26 );
not NOT1_15836 ( P2_R1179_U199 , P2_R1179_U71 );
not NOT1_15837 ( P2_R1179_U200 , P2_R1179_U85 );
not NOT1_15838 ( P2_R1179_U201 , P2_R1179_U44 );
not NOT1_15839 ( P2_R1179_U202 , P2_R1179_U59 );
not NOT1_15840 ( P2_R1179_U203 , P2_R1179_U175 );
nand NAND2_15841 ( P2_R1179_U204 , P2_U3077 , P2_R1179_U175 );
not NOT1_15842 ( P2_R1179_U205 , P2_R1179_U50 );
nand NAND2_15843 ( P2_R1179_U206 , P2_U3398 , P2_R1179_U36 );
nand NAND2_15844 ( P2_R1179_U207 , P2_R1179_U36 , P2_R1179_U35 );
nand NAND2_15845 ( P2_R1179_U208 , P2_R1179_U207 , P2_R1179_U40 );
nand NAND2_15846 ( P2_R1179_U209 , P2_U3063 , P2_R1179_U190 );
nand NAND2_15847 ( P2_R1179_U210 , P2_U3407 , P2_R1179_U41 );
nand NAND2_15848 ( P2_R1179_U211 , P2_U3070 , P2_R1179_U30 );
nand NAND2_15849 ( P2_R1179_U212 , P2_U3066 , P2_R1179_U29 );
nand NAND2_15850 ( P2_R1179_U213 , P2_R1179_U201 , P2_R1179_U197 );
nand NAND2_15851 ( P2_R1179_U214 , P2_R1179_U6 , P2_R1179_U213 );
nand NAND2_15852 ( P2_R1179_U215 , P2_U3401 , P2_R1179_U43 );
nand NAND2_15853 ( P2_R1179_U216 , P2_U3407 , P2_R1179_U41 );
nand NAND2_15854 ( P2_R1179_U217 , P2_R1179_U13 , P2_R1179_U161 );
not NOT1_15855 ( P2_R1179_U218 , P2_R1179_U45 );
not NOT1_15856 ( P2_R1179_U219 , P2_R1179_U48 );
nand NAND2_15857 ( P2_R1179_U220 , P2_U3413 , P2_R1179_U28 );
nand NAND2_15858 ( P2_R1179_U221 , P2_R1179_U28 , P2_R1179_U27 );
nand NAND2_15859 ( P2_R1179_U222 , P2_U3083 , P2_R1179_U191 );
not NOT1_15860 ( P2_R1179_U223 , P2_R1179_U157 );
nand NAND2_15861 ( P2_R1179_U224 , P2_U3416 , P2_R1179_U47 );
nand NAND2_15862 ( P2_R1179_U225 , P2_R1179_U224 , P2_R1179_U59 );
nand NAND2_15863 ( P2_R1179_U226 , P2_R1179_U219 , P2_R1179_U27 );
nand NAND2_15864 ( P2_R1179_U227 , P2_R1179_U125 , P2_R1179_U226 );
nand NAND2_15865 ( P2_R1179_U228 , P2_R1179_U48 , P2_R1179_U198 );
nand NAND2_15866 ( P2_R1179_U229 , P2_R1179_U124 , P2_R1179_U228 );
nand NAND2_15867 ( P2_R1179_U230 , P2_R1179_U27 , P2_R1179_U198 );
nand NAND2_15868 ( P2_R1179_U231 , P2_R1179_U215 , P2_R1179_U161 );
not NOT1_15869 ( P2_R1179_U232 , P2_R1179_U49 );
nand NAND2_15870 ( P2_R1179_U233 , P2_U3066 , P2_R1179_U29 );
nand NAND2_15871 ( P2_R1179_U234 , P2_R1179_U232 , P2_R1179_U233 );
nand NAND2_15872 ( P2_R1179_U235 , P2_R1179_U127 , P2_R1179_U234 );
nand NAND2_15873 ( P2_R1179_U236 , P2_R1179_U49 , P2_R1179_U197 );
nand NAND2_15874 ( P2_R1179_U237 , P2_U3407 , P2_R1179_U41 );
nand NAND2_15875 ( P2_R1179_U238 , P2_R1179_U126 , P2_R1179_U236 );
nand NAND2_15876 ( P2_R1179_U239 , P2_U3066 , P2_R1179_U29 );
nand NAND2_15877 ( P2_R1179_U240 , P2_R1179_U239 , P2_R1179_U197 );
nand NAND2_15878 ( P2_R1179_U241 , P2_R1179_U215 , P2_R1179_U44 );
nand NAND2_15879 ( P2_R1179_U242 , P2_R1179_U129 , P2_R1179_U348 );
nand NAND2_15880 ( P2_R1179_U243 , P2_R1179_U35 , P2_R1179_U196 );
nand NAND2_15881 ( P2_R1179_U244 , P2_U3422 , P2_R1179_U56 );
nand NAND2_15882 ( P2_R1179_U245 , P2_U3062 , P2_R1179_U60 );
nand NAND2_15883 ( P2_R1179_U246 , P2_U3061 , P2_R1179_U58 );
nand NAND2_15884 ( P2_R1179_U247 , P2_R1179_U202 , P2_R1179_U192 );
nand NAND2_15885 ( P2_R1179_U248 , P2_R1179_U7 , P2_R1179_U247 );
nand NAND2_15886 ( P2_R1179_U249 , P2_U3422 , P2_R1179_U56 );
not NOT1_15887 ( P2_R1179_U250 , P2_R1179_U62 );
nand NAND2_15888 ( P2_R1179_U251 , P2_U3425 , P2_R1179_U55 );
nand NAND2_15889 ( P2_R1179_U252 , P2_U3071 , P2_R1179_U61 );
nand NAND2_15890 ( P2_R1179_U253 , P2_U3428 , P2_R1179_U64 );
nand NAND2_15891 ( P2_R1179_U254 , P2_R1179_U253 , P2_R1179_U183 );
nand NAND2_15892 ( P2_R1179_U255 , P2_U3079 , P2_R1179_U63 );
not NOT1_15893 ( P2_R1179_U256 , P2_R1179_U182 );
nand NAND2_15894 ( P2_R1179_U257 , P2_U3437 , P2_R1179_U68 );
nand NAND2_15895 ( P2_R1179_U258 , P2_U3072 , P2_R1179_U65 );
nand NAND2_15896 ( P2_R1179_U259 , P2_U3073 , P2_R1179_U66 );
nand NAND2_15897 ( P2_R1179_U260 , P2_R1179_U199 , P2_R1179_U8 );
nand NAND2_15898 ( P2_R1179_U261 , P2_R1179_U9 , P2_R1179_U260 );
nand NAND2_15899 ( P2_R1179_U262 , P2_U3431 , P2_R1179_U70 );
nand NAND2_15900 ( P2_R1179_U263 , P2_U3437 , P2_R1179_U68 );
nand NAND2_15901 ( P2_R1179_U264 , P2_R1179_U132 , P2_R1179_U182 );
nand NAND2_15902 ( P2_R1179_U265 , P2_R1179_U263 , P2_R1179_U261 );
not NOT1_15903 ( P2_R1179_U266 , P2_R1179_U179 );
nand NAND2_15904 ( P2_R1179_U267 , P2_U3440 , P2_R1179_U73 );
nand NAND2_15905 ( P2_R1179_U268 , P2_R1179_U267 , P2_R1179_U179 );
nand NAND2_15906 ( P2_R1179_U269 , P2_U3068 , P2_R1179_U72 );
not NOT1_15907 ( P2_R1179_U270 , P2_R1179_U178 );
nand NAND2_15908 ( P2_R1179_U271 , P2_U3081 , P2_R1179_U178 );
not NOT1_15909 ( P2_R1179_U272 , P2_R1179_U176 );
nand NAND2_15910 ( P2_R1179_U273 , P2_U3445 , P2_R1179_U76 );
nand NAND2_15911 ( P2_R1179_U274 , P2_R1179_U273 , P2_R1179_U176 );
nand NAND2_15912 ( P2_R1179_U275 , P2_U3080 , P2_R1179_U75 );
not NOT1_15913 ( P2_R1179_U276 , P2_R1179_U173 );
nand NAND2_15914 ( P2_R1179_U277 , P2_U3903 , P2_R1179_U78 );
nand NAND2_15915 ( P2_R1179_U278 , P2_R1179_U277 , P2_R1179_U173 );
nand NAND2_15916 ( P2_R1179_U279 , P2_U3075 , P2_R1179_U77 );
not NOT1_15917 ( P2_R1179_U280 , P2_R1179_U172 );
nand NAND2_15918 ( P2_R1179_U281 , P2_U3900 , P2_R1179_U82 );
nand NAND2_15919 ( P2_R1179_U282 , P2_U3065 , P2_R1179_U79 );
nand NAND2_15920 ( P2_R1179_U283 , P2_U3060 , P2_R1179_U80 );
nand NAND2_15921 ( P2_R1179_U284 , P2_R1179_U200 , P2_R1179_U10 );
nand NAND2_15922 ( P2_R1179_U285 , P2_R1179_U11 , P2_R1179_U284 );
nand NAND2_15923 ( P2_R1179_U286 , P2_U3902 , P2_R1179_U84 );
nand NAND2_15924 ( P2_R1179_U287 , P2_U3900 , P2_R1179_U82 );
nand NAND2_15925 ( P2_R1179_U288 , P2_R1179_U133 , P2_R1179_U172 );
nand NAND2_15926 ( P2_R1179_U289 , P2_R1179_U287 , P2_R1179_U285 );
not NOT1_15927 ( P2_R1179_U290 , P2_R1179_U169 );
nand NAND2_15928 ( P2_R1179_U291 , P2_U3899 , P2_R1179_U87 );
nand NAND2_15929 ( P2_R1179_U292 , P2_R1179_U291 , P2_R1179_U169 );
nand NAND2_15930 ( P2_R1179_U293 , P2_U3064 , P2_R1179_U86 );
not NOT1_15931 ( P2_R1179_U294 , P2_R1179_U168 );
nand NAND2_15932 ( P2_R1179_U295 , P2_U3898 , P2_R1179_U89 );
nand NAND2_15933 ( P2_R1179_U296 , P2_R1179_U295 , P2_R1179_U168 );
nand NAND2_15934 ( P2_R1179_U297 , P2_U3057 , P2_R1179_U88 );
not NOT1_15935 ( P2_R1179_U298 , P2_R1179_U93 );
nand NAND2_15936 ( P2_R1179_U299 , P2_U3896 , P2_R1179_U54 );
nand NAND2_15937 ( P2_R1179_U300 , P2_R1179_U54 , P2_R1179_U53 );
nand NAND2_15938 ( P2_R1179_U301 , P2_R1179_U300 , P2_R1179_U91 );
nand NAND2_15939 ( P2_R1179_U302 , P2_U3052 , P2_R1179_U189 );
nand NAND2_15940 ( P2_R1179_U303 , P2_U3895 , P2_R1179_U92 );
nand NAND2_15941 ( P2_R1179_U304 , P2_U3053 , P2_R1179_U51 );
nand NAND2_15942 ( P2_R1179_U305 , P2_R1179_U140 , P2_R1179_U355 );
nand NAND2_15943 ( P2_R1179_U306 , P2_R1179_U53 , P2_R1179_U195 );
nand NAND2_15944 ( P2_R1179_U307 , P2_R1179_U286 , P2_R1179_U172 );
not NOT1_15945 ( P2_R1179_U308 , P2_R1179_U94 );
nand NAND2_15946 ( P2_R1179_U309 , P2_U3060 , P2_R1179_U80 );
nand NAND2_15947 ( P2_R1179_U310 , P2_R1179_U308 , P2_R1179_U309 );
nand NAND2_15948 ( P2_R1179_U311 , P2_R1179_U144 , P2_R1179_U310 );
nand NAND2_15949 ( P2_R1179_U312 , P2_R1179_U94 , P2_R1179_U194 );
nand NAND2_15950 ( P2_R1179_U313 , P2_U3900 , P2_R1179_U82 );
nand NAND2_15951 ( P2_R1179_U314 , P2_R1179_U143 , P2_R1179_U312 );
nand NAND2_15952 ( P2_R1179_U315 , P2_U3060 , P2_R1179_U80 );
nand NAND2_15953 ( P2_R1179_U316 , P2_R1179_U194 , P2_R1179_U315 );
nand NAND2_15954 ( P2_R1179_U317 , P2_R1179_U286 , P2_R1179_U85 );
nand NAND2_15955 ( P2_R1179_U318 , P2_R1179_U262 , P2_R1179_U182 );
not NOT1_15956 ( P2_R1179_U319 , P2_R1179_U95 );
nand NAND2_15957 ( P2_R1179_U320 , P2_U3073 , P2_R1179_U66 );
nand NAND2_15958 ( P2_R1179_U321 , P2_R1179_U319 , P2_R1179_U320 );
nand NAND2_15959 ( P2_R1179_U322 , P2_R1179_U151 , P2_R1179_U321 );
nand NAND2_15960 ( P2_R1179_U323 , P2_R1179_U95 , P2_R1179_U193 );
nand NAND2_15961 ( P2_R1179_U324 , P2_U3437 , P2_R1179_U68 );
nand NAND2_15962 ( P2_R1179_U325 , P2_R1179_U150 , P2_R1179_U323 );
nand NAND2_15963 ( P2_R1179_U326 , P2_U3073 , P2_R1179_U66 );
nand NAND2_15964 ( P2_R1179_U327 , P2_R1179_U193 , P2_R1179_U326 );
nand NAND2_15965 ( P2_R1179_U328 , P2_R1179_U262 , P2_R1179_U71 );
nand NAND2_15966 ( P2_R1179_U329 , P2_U3061 , P2_R1179_U58 );
nand NAND2_15967 ( P2_R1179_U330 , P2_R1179_U350 , P2_R1179_U329 );
nand NAND2_15968 ( P2_R1179_U331 , P2_R1179_U155 , P2_R1179_U330 );
nand NAND2_15969 ( P2_R1179_U332 , P2_R1179_U96 , P2_R1179_U192 );
nand NAND2_15970 ( P2_R1179_U333 , P2_U3422 , P2_R1179_U56 );
nand NAND2_15971 ( P2_R1179_U334 , P2_R1179_U154 , P2_R1179_U332 );
nand NAND2_15972 ( P2_R1179_U335 , P2_U3061 , P2_R1179_U58 );
nand NAND2_15973 ( P2_R1179_U336 , P2_R1179_U192 , P2_R1179_U335 );
nand NAND2_15974 ( P2_R1179_U337 , P2_U3076 , P2_R1179_U38 );
nand NAND2_15975 ( P2_R1179_U338 , P2_U3077 , P2_R1179_U174 );
nand NAND2_15976 ( P2_R1179_U339 , P2_U3081 , P2_R1179_U177 );
nand NAND2_15977 ( P2_R1179_U340 , P2_R1179_U33 , P2_R1179_U221 );
nand NAND2_15978 ( P2_R1179_U341 , P2_R1179_U121 , P2_R1179_U161 );
nand NAND2_15979 ( P2_R1179_U342 , P2_R1179_U218 , P2_R1179_U14 );
nand NAND2_15980 ( P2_R1179_U343 , P2_R1179_U250 , P2_R1179_U251 );
nand NAND2_15981 ( P2_R1179_U344 , P2_R1179_U119 , P2_R1179_U50 );
not NOT1_15982 ( P2_R1179_U345 , P2_R1179_U161 );
nand NAND2_15983 ( P2_R1179_U346 , P2_R1179_U196 , P2_R1179_U50 );
nand NAND2_15984 ( P2_R1179_U347 , P2_R1179_U128 , P2_R1179_U346 );
nand NAND2_15985 ( P2_R1179_U348 , P2_R1179_U205 , P2_R1179_U35 );
nand NAND2_15986 ( P2_R1179_U349 , P2_R1179_U224 , P2_R1179_U157 );
not NOT1_15987 ( P2_R1179_U350 , P2_R1179_U96 );
nand NAND2_15988 ( P2_R1179_U351 , P2_R1179_U15 , P2_R1179_U157 );
not NOT1_15989 ( P2_R1179_U352 , P2_R1179_U184 );
nand NAND2_15990 ( P2_R1179_U353 , P2_R1179_U130 , P2_R1179_U157 );
not NOT1_15991 ( P2_R1179_U354 , P2_R1179_U183 );
nand NAND2_15992 ( P2_R1179_U355 , P2_R1179_U298 , P2_R1179_U53 );
nand NAND2_15993 ( P2_R1179_U356 , P2_R1179_U195 , P2_R1179_U93 );
nand NAND2_15994 ( P2_R1179_U357 , P2_R1179_U139 , P2_R1179_U356 );
nand NAND2_15995 ( P2_R1179_U358 , P2_R1179_U12 , P2_R1179_U93 );
nand NAND2_15996 ( P2_R1179_U359 , P2_R1179_U136 , P2_R1179_U358 );
nand NAND2_15997 ( P2_R1179_U360 , P2_R1179_U12 , P2_R1179_U93 );
not NOT1_15998 ( P2_R1179_U361 , P2_R1179_U166 );
nand NAND2_15999 ( P2_R1179_U362 , P2_U3416 , P2_R1179_U47 );
nand NAND2_16000 ( P2_R1179_U363 , P2_U3082 , P2_R1179_U46 );
nand NAND2_16001 ( P2_R1179_U364 , P2_R1179_U225 , P2_R1179_U157 );
nand NAND2_16002 ( P2_R1179_U365 , P2_R1179_U223 , P2_R1179_U156 );
nand NAND2_16003 ( P2_R1179_U366 , P2_U3413 , P2_R1179_U28 );
nand NAND2_16004 ( P2_R1179_U367 , P2_U3083 , P2_R1179_U33 );
nand NAND2_16005 ( P2_R1179_U368 , P2_U3413 , P2_R1179_U28 );
nand NAND2_16006 ( P2_R1179_U369 , P2_U3083 , P2_R1179_U33 );
nand NAND2_16007 ( P2_R1179_U370 , P2_R1179_U369 , P2_R1179_U368 );
nand NAND2_16008 ( P2_R1179_U371 , P2_U3410 , P2_R1179_U26 );
nand NAND2_16009 ( P2_R1179_U372 , P2_U3069 , P2_R1179_U32 );
nand NAND2_16010 ( P2_R1179_U373 , P2_R1179_U230 , P2_R1179_U48 );
nand NAND2_16011 ( P2_R1179_U374 , P2_R1179_U158 , P2_R1179_U219 );
nand NAND2_16012 ( P2_R1179_U375 , P2_U3407 , P2_R1179_U41 );
nand NAND2_16013 ( P2_R1179_U376 , P2_U3070 , P2_R1179_U30 );
nand NAND2_16014 ( P2_R1179_U377 , P2_R1179_U376 , P2_R1179_U375 );
nand NAND2_16015 ( P2_R1179_U378 , P2_U3404 , P2_R1179_U42 );
nand NAND2_16016 ( P2_R1179_U379 , P2_U3066 , P2_R1179_U29 );
nand NAND2_16017 ( P2_R1179_U380 , P2_R1179_U240 , P2_R1179_U49 );
nand NAND2_16018 ( P2_R1179_U381 , P2_R1179_U159 , P2_R1179_U232 );
nand NAND2_16019 ( P2_R1179_U382 , P2_U3401 , P2_R1179_U43 );
nand NAND2_16020 ( P2_R1179_U383 , P2_U3059 , P2_R1179_U31 );
nand NAND2_16021 ( P2_R1179_U384 , P2_R1179_U161 , P2_R1179_U241 );
nand NAND2_16022 ( P2_R1179_U385 , P2_R1179_U345 , P2_R1179_U160 );
nand NAND2_16023 ( P2_R1179_U386 , P2_U3398 , P2_R1179_U36 );
nand NAND2_16024 ( P2_R1179_U387 , P2_U3063 , P2_R1179_U40 );
nand NAND2_16025 ( P2_R1179_U388 , P2_U3398 , P2_R1179_U36 );
nand NAND2_16026 ( P2_R1179_U389 , P2_U3063 , P2_R1179_U40 );
nand NAND2_16027 ( P2_R1179_U390 , P2_R1179_U389 , P2_R1179_U388 );
nand NAND2_16028 ( P2_R1179_U391 , P2_U3395 , P2_R1179_U34 );
nand NAND2_16029 ( P2_R1179_U392 , P2_U3067 , P2_R1179_U37 );
nand NAND2_16030 ( P2_R1179_U393 , P2_R1179_U243 , P2_R1179_U50 );
nand NAND2_16031 ( P2_R1179_U394 , P2_R1179_U162 , P2_R1179_U205 );
nand NAND2_16032 ( P2_R1179_U395 , P2_U3904 , P2_R1179_U164 );
nand NAND2_16033 ( P2_R1179_U396 , P2_U3054 , P2_R1179_U163 );
nand NAND2_16034 ( P2_R1179_U397 , P2_R1179_U396 , P2_R1179_U395 );
nand NAND2_16035 ( P2_R1179_U398 , P2_U3904 , P2_R1179_U164 );
nand NAND2_16036 ( P2_R1179_U399 , P2_U3054 , P2_R1179_U163 );
nand NAND3_16037 ( P2_R1179_U400 , P2_U3053 , P2_R1179_U397 , P2_R1179_U51 );
nand NAND3_16038 ( P2_R1179_U401 , P2_R1179_U16 , P2_R1179_U92 , P2_U3895 );
nand NAND2_16039 ( P2_R1179_U402 , P2_U3895 , P2_R1179_U92 );
nand NAND2_16040 ( P2_R1179_U403 , P2_U3053 , P2_R1179_U51 );
not NOT1_16041 ( P2_R1179_U404 , P2_R1179_U138 );
nand NAND2_16042 ( P2_R1179_U405 , P2_R1179_U361 , P2_R1179_U404 );
nand NAND2_16043 ( P2_R1179_U406 , P2_R1179_U138 , P2_R1179_U166 );
nand NAND2_16044 ( P2_R1179_U407 , P2_U3896 , P2_R1179_U54 );
nand NAND2_16045 ( P2_R1179_U408 , P2_U3052 , P2_R1179_U91 );
nand NAND2_16046 ( P2_R1179_U409 , P2_U3896 , P2_R1179_U54 );
nand NAND2_16047 ( P2_R1179_U410 , P2_U3052 , P2_R1179_U91 );
nand NAND2_16048 ( P2_R1179_U411 , P2_R1179_U410 , P2_R1179_U409 );
nand NAND2_16049 ( P2_R1179_U412 , P2_U3897 , P2_R1179_U52 );
nand NAND2_16050 ( P2_R1179_U413 , P2_U3056 , P2_R1179_U90 );
nand NAND2_16051 ( P2_R1179_U414 , P2_R1179_U306 , P2_R1179_U93 );
nand NAND2_16052 ( P2_R1179_U415 , P2_R1179_U167 , P2_R1179_U298 );
nand NAND2_16053 ( P2_R1179_U416 , P2_U3898 , P2_R1179_U89 );
nand NAND2_16054 ( P2_R1179_U417 , P2_U3057 , P2_R1179_U88 );
not NOT1_16055 ( P2_R1179_U418 , P2_R1179_U141 );
nand NAND2_16056 ( P2_R1179_U419 , P2_R1179_U294 , P2_R1179_U418 );
nand NAND2_16057 ( P2_R1179_U420 , P2_R1179_U141 , P2_R1179_U168 );
nand NAND2_16058 ( P2_R1179_U421 , P2_U3899 , P2_R1179_U87 );
nand NAND2_16059 ( P2_R1179_U422 , P2_U3064 , P2_R1179_U86 );
not NOT1_16060 ( P2_R1179_U423 , P2_R1179_U142 );
nand NAND2_16061 ( P2_R1179_U424 , P2_R1179_U290 , P2_R1179_U423 );
nand NAND2_16062 ( P2_R1179_U425 , P2_R1179_U142 , P2_R1179_U169 );
nand NAND2_16063 ( P2_R1179_U426 , P2_U3900 , P2_R1179_U82 );
nand NAND2_16064 ( P2_R1179_U427 , P2_U3065 , P2_R1179_U79 );
nand NAND2_16065 ( P2_R1179_U428 , P2_R1179_U427 , P2_R1179_U426 );
nand NAND2_16066 ( P2_R1179_U429 , P2_U3901 , P2_R1179_U83 );
nand NAND2_16067 ( P2_R1179_U430 , P2_U3060 , P2_R1179_U80 );
nand NAND2_16068 ( P2_R1179_U431 , P2_R1179_U316 , P2_R1179_U94 );
nand NAND2_16069 ( P2_R1179_U432 , P2_R1179_U170 , P2_R1179_U308 );
nand NAND2_16070 ( P2_R1179_U433 , P2_U3902 , P2_R1179_U84 );
nand NAND2_16071 ( P2_R1179_U434 , P2_U3074 , P2_R1179_U81 );
nand NAND2_16072 ( P2_R1179_U435 , P2_R1179_U317 , P2_R1179_U172 );
nand NAND2_16073 ( P2_R1179_U436 , P2_R1179_U280 , P2_R1179_U171 );
nand NAND2_16074 ( P2_R1179_U437 , P2_U3903 , P2_R1179_U78 );
nand NAND2_16075 ( P2_R1179_U438 , P2_U3075 , P2_R1179_U77 );
not NOT1_16076 ( P2_R1179_U439 , P2_R1179_U145 );
nand NAND2_16077 ( P2_R1179_U440 , P2_R1179_U276 , P2_R1179_U439 );
nand NAND2_16078 ( P2_R1179_U441 , P2_R1179_U145 , P2_R1179_U173 );
nand NAND2_16079 ( P2_R1179_U442 , P2_U3392 , P2_R1179_U39 );
nand NAND2_16080 ( P2_R1179_U443 , P2_U3077 , P2_R1179_U174 );
not NOT1_16081 ( P2_R1179_U444 , P2_R1179_U146 );
nand NAND2_16082 ( P2_R1179_U445 , P2_R1179_U203 , P2_R1179_U444 );
nand NAND2_16083 ( P2_R1179_U446 , P2_R1179_U146 , P2_R1179_U175 );
nand NAND2_16084 ( P2_R1179_U447 , P2_U3445 , P2_R1179_U76 );
nand NAND2_16085 ( P2_R1179_U448 , P2_U3080 , P2_R1179_U75 );
not NOT1_16086 ( P2_R1179_U449 , P2_R1179_U147 );
nand NAND2_16087 ( P2_R1179_U450 , P2_R1179_U272 , P2_R1179_U449 );
nand NAND2_16088 ( P2_R1179_U451 , P2_R1179_U147 , P2_R1179_U176 );
nand NAND2_16089 ( P2_R1179_U452 , P2_U3443 , P2_R1179_U74 );
nand NAND2_16090 ( P2_R1179_U453 , P2_U3081 , P2_R1179_U177 );
not NOT1_16091 ( P2_R1179_U454 , P2_R1179_U148 );
nand NAND2_16092 ( P2_R1179_U455 , P2_R1179_U270 , P2_R1179_U454 );
nand NAND2_16093 ( P2_R1179_U456 , P2_R1179_U148 , P2_R1179_U178 );
nand NAND2_16094 ( P2_R1179_U457 , P2_U3440 , P2_R1179_U73 );
nand NAND2_16095 ( P2_R1179_U458 , P2_U3068 , P2_R1179_U72 );
not NOT1_16096 ( P2_R1179_U459 , P2_R1179_U149 );
nand NAND2_16097 ( P2_R1179_U460 , P2_R1179_U266 , P2_R1179_U459 );
nand NAND2_16098 ( P2_R1179_U461 , P2_R1179_U149 , P2_R1179_U179 );
nand NAND2_16099 ( P2_R1179_U462 , P2_U3437 , P2_R1179_U68 );
nand NAND2_16100 ( P2_R1179_U463 , P2_U3072 , P2_R1179_U65 );
nand NAND2_16101 ( P2_R1179_U464 , P2_R1179_U463 , P2_R1179_U462 );
nand NAND2_16102 ( P2_R1179_U465 , P2_U3434 , P2_R1179_U69 );
nand NAND2_16103 ( P2_R1179_U466 , P2_U3073 , P2_R1179_U66 );
nand NAND2_16104 ( P2_R1179_U467 , P2_R1179_U327 , P2_R1179_U95 );
nand NAND2_16105 ( P2_R1179_U468 , P2_R1179_U180 , P2_R1179_U319 );
nand NAND2_16106 ( P2_R1179_U469 , P2_U3431 , P2_R1179_U70 );
nand NAND2_16107 ( P2_R1179_U470 , P2_U3078 , P2_R1179_U67 );
nand NAND2_16108 ( P2_R1179_U471 , P2_R1179_U328 , P2_R1179_U182 );
nand NAND2_16109 ( P2_R1179_U472 , P2_R1179_U256 , P2_R1179_U181 );
nand NAND2_16110 ( P2_R1179_U473 , P2_U3428 , P2_R1179_U64 );
nand NAND2_16111 ( P2_R1179_U474 , P2_U3079 , P2_R1179_U63 );
not NOT1_16112 ( P2_R1179_U475 , P2_R1179_U152 );
nand NAND2_16113 ( P2_R1179_U476 , P2_R1179_U354 , P2_R1179_U475 );
nand NAND2_16114 ( P2_R1179_U477 , P2_R1179_U152 , P2_R1179_U183 );
nand NAND2_16115 ( P2_R1179_U478 , P2_U3425 , P2_R1179_U55 );
nand NAND2_16116 ( P2_R1179_U479 , P2_U3071 , P2_R1179_U61 );
not NOT1_16117 ( P2_R1179_U480 , P2_R1179_U153 );
nand NAND2_16118 ( P2_R1179_U481 , P2_R1179_U352 , P2_R1179_U480 );
nand NAND2_16119 ( P2_R1179_U482 , P2_R1179_U153 , P2_R1179_U184 );
nand NAND2_16120 ( P2_R1179_U483 , P2_U3422 , P2_R1179_U56 );
nand NAND2_16121 ( P2_R1179_U484 , P2_U3062 , P2_R1179_U60 );
nand NAND2_16122 ( P2_R1179_U485 , P2_R1179_U484 , P2_R1179_U483 );
nand NAND2_16123 ( P2_R1179_U486 , P2_U3419 , P2_R1179_U57 );
nand NAND2_16124 ( P2_R1179_U487 , P2_U3061 , P2_R1179_U58 );
nand NAND2_16125 ( P2_R1179_U488 , P2_R1179_U96 , P2_R1179_U336 );
nand NAND2_16126 ( P2_R1179_U489 , P2_R1179_U185 , P2_R1179_U350 );
and AND2_16127 ( P2_R1269_U6 , P2_R1269_U130 , P2_R1269_U131 );
and AND2_16128 ( P2_R1269_U7 , P2_R1269_U132 , P2_R1269_U133 );
and AND4_16129 ( P2_R1269_U8 , P2_R1269_U91 , P2_R1269_U135 , P2_R1269_U137 , P2_R1269_U7 );
and AND2_16130 ( P2_R1269_U9 , P2_R1269_U144 , P2_R1269_U145 );
and AND2_16131 ( P2_R1269_U10 , P2_R1269_U147 , P2_R1269_U146 );
and AND3_16132 ( P2_R1269_U11 , P2_R1269_U94 , P2_R1269_U148 , P2_R1269_U95 );
and AND2_16133 ( P2_R1269_U12 , P2_R1269_U96 , P2_R1269_U11 );
and AND2_16134 ( P2_R1269_U13 , P2_R1269_U163 , P2_R1269_U162 );
and AND5_16135 ( P2_R1269_U14 , P2_R1269_U195 , P2_R1269_U191 , P2_R1269_U113 , P2_R1269_U20 , P2_R1269_U21 );
and AND2_16136 ( P2_R1269_U15 , P2_R1269_U129 , P2_R1269_U128 );
and AND3_16137 ( P2_R1269_U16 , P2_R1269_U114 , P2_R1269_U20 , P2_R1269_U21 );
and AND3_16138 ( P2_R1269_U17 , P2_R1269_U115 , P2_R1269_U20 , P2_R1269_U21 );
and AND2_16139 ( P2_R1269_U18 , P2_R1269_U117 , P2_R1269_U21 );
and AND2_16140 ( P2_R1269_U19 , P2_R1269_U118 , P2_R1269_U21 );
and AND3_16141 ( P2_R1269_U20 , P2_R1269_U124 , P2_R1269_U125 , P2_R1269_U123 );
and AND2_16142 ( P2_R1269_U21 , P2_R1269_U207 , P2_R1269_U206 );
nand NAND4_16143 ( P2_R1269_U22 , P2_R1269_U200 , P2_R1269_U127 , P2_R1269_U119 , P2_R1269_U120 );
not NOT1_16144 ( P2_R1269_U23 , P2_U3085 );
not NOT1_16145 ( P2_R1269_U24 , P2_U3084 );
not NOT1_16146 ( P2_R1269_U25 , P2_U3116 );
not NOT1_16147 ( P2_R1269_U26 , P2_U3118 );
not NOT1_16148 ( P2_R1269_U27 , P2_U3117 );
not NOT1_16149 ( P2_R1269_U28 , P2_U3086 );
not NOT1_16150 ( P2_R1269_U29 , P2_U3124 );
not NOT1_16151 ( P2_R1269_U30 , P2_U3123 );
not NOT1_16152 ( P2_R1269_U31 , P2_U3094 );
not NOT1_16153 ( P2_R1269_U32 , P2_U3127 );
not NOT1_16154 ( P2_R1269_U33 , P2_U3095 );
not NOT1_16155 ( P2_R1269_U34 , P2_U3128 );
not NOT1_16156 ( P2_R1269_U35 , P2_U3129 );
not NOT1_16157 ( P2_R1269_U36 , P2_U3098 );
not NOT1_16158 ( P2_R1269_U37 , P2_U3130 );
not NOT1_16159 ( P2_R1269_U38 , P2_U3099 );
not NOT1_16160 ( P2_R1269_U39 , P2_U3097 );
not NOT1_16161 ( P2_R1269_U40 , P2_U3096 );
not NOT1_16162 ( P2_R1269_U41 , P2_U3131 );
not NOT1_16163 ( P2_R1269_U42 , P2_U3132 );
not NOT1_16164 ( P2_R1269_U43 , P2_U3100 );
not NOT1_16165 ( P2_R1269_U44 , P2_U3101 );
not NOT1_16166 ( P2_R1269_U45 , P2_U3141 );
not NOT1_16167 ( P2_R1269_U46 , P2_U3110 );
not NOT1_16168 ( P2_R1269_U47 , P2_U3107 );
not NOT1_16169 ( P2_R1269_U48 , P2_U3106 );
not NOT1_16170 ( P2_R1269_U49 , P2_U3142 );
not NOT1_16171 ( P2_R1269_U50 , P2_U3111 );
not NOT1_16172 ( P2_R1269_U51 , P2_U3109 );
not NOT1_16173 ( P2_R1269_U52 , P2_U3108 );
not NOT1_16174 ( P2_R1269_U53 , P2_U3112 );
not NOT1_16175 ( P2_R1269_U54 , P2_U3113 );
not NOT1_16176 ( P2_R1269_U55 , P2_U3114 );
not NOT1_16177 ( P2_R1269_U56 , P2_U3136 );
not NOT1_16178 ( P2_R1269_U57 , P2_U3135 );
not NOT1_16179 ( P2_R1269_U58 , P2_U3139 );
not NOT1_16180 ( P2_R1269_U59 , P2_U3140 );
not NOT1_16181 ( P2_R1269_U60 , P2_U3146 );
not NOT1_16182 ( P2_R1269_U61 , P2_U3145 );
not NOT1_16183 ( P2_R1269_U62 , P2_U3143 );
not NOT1_16184 ( P2_R1269_U63 , P2_U3144 );
not NOT1_16185 ( P2_R1269_U64 , P2_U3138 );
not NOT1_16186 ( P2_R1269_U65 , P2_U3137 );
not NOT1_16187 ( P2_R1269_U66 , P2_U3104 );
not NOT1_16188 ( P2_R1269_U67 , P2_U3105 );
not NOT1_16189 ( P2_R1269_U68 , P2_U3102 );
not NOT1_16190 ( P2_R1269_U69 , P2_U3103 );
not NOT1_16191 ( P2_R1269_U70 , P2_U3134 );
not NOT1_16192 ( P2_R1269_U71 , P2_U3133 );
not NOT1_16193 ( P2_R1269_U72 , P2_U3126 );
not NOT1_16194 ( P2_R1269_U73 , P2_U3125 );
not NOT1_16195 ( P2_R1269_U74 , P2_U3093 );
not NOT1_16196 ( P2_R1269_U75 , P2_U3092 );
not NOT1_16197 ( P2_R1269_U76 , P2_U3090 );
not NOT1_16198 ( P2_R1269_U77 , P2_U3091 );
not NOT1_16199 ( P2_R1269_U78 , P2_U3087 );
not NOT1_16200 ( P2_R1269_U79 , P2_U3089 );
not NOT1_16201 ( P2_R1269_U80 , P2_U3088 );
not NOT1_16202 ( P2_R1269_U81 , P2_U3122 );
not NOT1_16203 ( P2_R1269_U82 , P2_U3121 );
not NOT1_16204 ( P2_R1269_U83 , P2_U3120 );
not NOT1_16205 ( P2_R1269_U84 , P2_U3119 );
and AND2_16206 ( P2_R1269_U85 , P2_R1269_U28 , P2_U3118 );
and AND2_16207 ( P2_R1269_U86 , P2_U3127 , P2_R1269_U33 );
and AND2_16208 ( P2_R1269_U87 , P2_U3128 , P2_R1269_U40 );
and AND2_16209 ( P2_R1269_U88 , P2_R1269_U183 , P2_R1269_U182 );
and AND2_16210 ( P2_R1269_U89 , P2_U3098 , P2_R1269_U37 );
and AND2_16211 ( P2_R1269_U90 , P2_U3099 , P2_R1269_U41 );
and AND2_16212 ( P2_R1269_U91 , P2_R1269_U136 , P2_R1269_U134 );
and AND2_16213 ( P2_R1269_U92 , P2_U3110 , P2_R1269_U49 );
and AND2_16214 ( P2_R1269_U93 , P2_U3111 , P2_R1269_U62 );
and AND2_16215 ( P2_R1269_U94 , P2_R1269_U149 , P2_R1269_U143 );
and AND2_16216 ( P2_R1269_U95 , P2_R1269_U9 , P2_R1269_U150 );
and AND2_16217 ( P2_R1269_U96 , P2_R1269_U152 , P2_R1269_U151 );
and AND3_16218 ( P2_R1269_U97 , P2_R1269_U155 , P2_R1269_U156 , P2_R1269_U154 );
and AND2_16219 ( P2_R1269_U98 , P2_U3139 , P2_R1269_U47 );
and AND2_16220 ( P2_R1269_U99 , P2_U3140 , P2_R1269_U52 );
and AND2_16221 ( P2_R1269_U100 , P2_U3146 , P2_R1269_U55 );
and AND2_16222 ( P2_R1269_U101 , P2_U3145 , P2_R1269_U54 );
and AND2_16223 ( P2_R1269_U102 , P2_R1269_U13 , P2_R1269_U103 );
and AND2_16224 ( P2_R1269_U103 , P2_R1269_U168 , P2_R1269_U169 );
and AND2_16225 ( P2_R1269_U104 , P2_R1269_U167 , P2_R1269_U102 );
and AND2_16226 ( P2_R1269_U105 , P2_U3104 , P2_R1269_U56 );
and AND2_16227 ( P2_R1269_U106 , P2_U3105 , P2_R1269_U65 );
and AND2_16228 ( P2_R1269_U107 , P2_R1269_U172 , P2_R1269_U109 );
and AND2_16229 ( P2_R1269_U108 , P2_R1269_U107 , P2_R1269_U173 );
and AND2_16230 ( P2_R1269_U109 , P2_R1269_U175 , P2_R1269_U174 );
and AND3_16231 ( P2_R1269_U110 , P2_R1269_U186 , P2_R1269_U185 , P2_R1269_U139 );
and AND2_16232 ( P2_R1269_U111 , P2_R1269_U190 , P2_R1269_U189 );
and AND2_16233 ( P2_R1269_U112 , P2_U3093 , P2_R1269_U73 );
and AND2_16234 ( P2_R1269_U113 , P2_R1269_U197 , P2_R1269_U196 );
and AND2_16235 ( P2_R1269_U114 , P2_U3122 , P2_R1269_U76 );
and AND2_16236 ( P2_R1269_U115 , P2_U3121 , P2_R1269_U79 );
and AND2_16237 ( P2_R1269_U116 , P2_U3120 , P2_R1269_U80 );
and AND2_16238 ( P2_R1269_U117 , P2_R1269_U116 , P2_R1269_U123 );
and AND2_16239 ( P2_R1269_U118 , P2_U3119 , P2_R1269_U78 );
and AND2_16240 ( P2_R1269_U119 , P2_R1269_U202 , P2_R1269_U201 );
and AND3_16241 ( P2_R1269_U120 , P2_R1269_U204 , P2_R1269_U203 , P2_R1269_U15 );
nand NAND2_16242 ( P2_R1269_U121 , P2_R1269_U199 , P2_R1269_U198 );
nand NAND2_16243 ( P2_R1269_U122 , P2_U3086 , P2_R1269_U26 );
nand NAND2_16244 ( P2_R1269_U123 , P2_U3087 , P2_R1269_U84 );
nand NAND2_16245 ( P2_R1269_U124 , P2_U3089 , P2_R1269_U82 );
nand NAND2_16246 ( P2_R1269_U125 , P2_U3088 , P2_R1269_U83 );
nand NAND2_16247 ( P2_R1269_U126 , P2_U3085 , P2_R1269_U27 );
nand NAND3_16248 ( P2_R1269_U127 , P2_R1269_U85 , P2_R1269_U21 , P2_R1269_U126 );
nand NAND3_16249 ( P2_R1269_U128 , P2_R1269_U209 , P2_R1269_U208 , P2_R1269_U205 );
nand NAND3_16250 ( P2_R1269_U129 , P2_R1269_U21 , P2_R1269_U23 , P2_U3117 );
nand NAND2_16251 ( P2_R1269_U130 , P2_U3129 , P2_R1269_U39 );
nand NAND2_16252 ( P2_R1269_U131 , P2_U3130 , P2_R1269_U36 );
nand NAND2_16253 ( P2_R1269_U132 , P2_U3094 , P2_R1269_U72 );
nand NAND2_16254 ( P2_R1269_U133 , P2_U3095 , P2_R1269_U32 );
nand NAND2_16255 ( P2_R1269_U134 , P2_R1269_U89 , P2_R1269_U130 );
nand NAND2_16256 ( P2_R1269_U135 , P2_R1269_U90 , P2_R1269_U6 );
nand NAND2_16257 ( P2_R1269_U136 , P2_U3097 , P2_R1269_U35 );
nand NAND2_16258 ( P2_R1269_U137 , P2_U3096 , P2_R1269_U34 );
nand NAND2_16259 ( P2_R1269_U138 , P2_U3100 , P2_R1269_U42 );
nand NAND2_16260 ( P2_R1269_U139 , P2_U3124 , P2_R1269_U75 );
nand NAND2_16261 ( P2_R1269_U140 , P2_U3123 , P2_R1269_U77 );
nand NAND2_16262 ( P2_R1269_U141 , P2_U3101 , P2_R1269_U71 );
nand NAND2_16263 ( P2_R1269_U142 , P2_U3141 , P2_R1269_U51 );
nand NAND2_16264 ( P2_R1269_U143 , P2_R1269_U92 , P2_R1269_U142 );
nand NAND2_16265 ( P2_R1269_U144 , P2_U3106 , P2_R1269_U64 );
nand NAND2_16266 ( P2_R1269_U145 , P2_U3107 , P2_R1269_U58 );
nand NAND2_16267 ( P2_R1269_U146 , P2_U3142 , P2_R1269_U46 );
nand NAND2_16268 ( P2_R1269_U147 , P2_U3141 , P2_R1269_U51 );
nand NAND2_16269 ( P2_R1269_U148 , P2_R1269_U93 , P2_R1269_U10 );
nand NAND2_16270 ( P2_R1269_U149 , P2_U3109 , P2_R1269_U45 );
nand NAND2_16271 ( P2_R1269_U150 , P2_U3108 , P2_R1269_U59 );
nand NAND2_16272 ( P2_R1269_U151 , P2_U3112 , P2_R1269_U63 );
nand NAND2_16273 ( P2_R1269_U152 , P2_U3113 , P2_R1269_U61 );
nand NAND2_16274 ( P2_R1269_U153 , P2_U3147 , P2_U3148 );
nand NAND2_16275 ( P2_R1269_U154 , P2_U3115 , P2_R1269_U153 );
or OR2_16276 ( P2_R1269_U155 , P2_U3147 , P2_U3148 );
nand NAND2_16277 ( P2_R1269_U156 , P2_U3114 , P2_R1269_U60 );
nand NAND2_16278 ( P2_R1269_U157 , P2_R1269_U97 , P2_R1269_U12 );
nand NAND2_16279 ( P2_R1269_U158 , P2_R1269_U101 , P2_R1269_U151 );
nand NAND2_16280 ( P2_R1269_U159 , P2_U3143 , P2_R1269_U50 );
nand NAND2_16281 ( P2_R1269_U160 , P2_U3144 , P2_R1269_U53 );
nand NAND4_16282 ( P2_R1269_U161 , P2_R1269_U10 , P2_R1269_U160 , P2_R1269_U159 , P2_R1269_U158 );
nand NAND2_16283 ( P2_R1269_U162 , P2_U3136 , P2_R1269_U66 );
nand NAND2_16284 ( P2_R1269_U163 , P2_U3135 , P2_R1269_U69 );
nand NAND2_16285 ( P2_R1269_U164 , P2_R1269_U98 , P2_R1269_U144 );
nand NAND2_16286 ( P2_R1269_U165 , P2_R1269_U99 , P2_R1269_U9 );
nand NAND2_16287 ( P2_R1269_U166 , P2_R1269_U100 , P2_R1269_U12 );
nand NAND2_16288 ( P2_R1269_U167 , P2_R1269_U11 , P2_R1269_U161 );
nand NAND2_16289 ( P2_R1269_U168 , P2_U3138 , P2_R1269_U48 );
nand NAND2_16290 ( P2_R1269_U169 , P2_U3137 , P2_R1269_U67 );
nand NAND5_16291 ( P2_R1269_U170 , P2_R1269_U166 , P2_R1269_U165 , P2_R1269_U164 , P2_R1269_U157 , P2_R1269_U104 );
nand NAND2_16292 ( P2_R1269_U171 , P2_U3135 , P2_R1269_U69 );
nand NAND2_16293 ( P2_R1269_U172 , P2_R1269_U105 , P2_R1269_U171 );
nand NAND2_16294 ( P2_R1269_U173 , P2_R1269_U106 , P2_R1269_U13 );
nand NAND2_16295 ( P2_R1269_U174 , P2_U3102 , P2_R1269_U70 );
nand NAND2_16296 ( P2_R1269_U175 , P2_U3103 , P2_R1269_U57 );
nand NAND2_16297 ( P2_R1269_U176 , P2_R1269_U170 , P2_R1269_U108 );
nand NAND2_16298 ( P2_R1269_U177 , P2_U3134 , P2_R1269_U68 );
nand NAND2_16299 ( P2_R1269_U178 , P2_R1269_U177 , P2_R1269_U176 );
nand NAND2_16300 ( P2_R1269_U179 , P2_R1269_U178 , P2_R1269_U141 );
nand NAND2_16301 ( P2_R1269_U180 , P2_U3133 , P2_R1269_U44 );
nand NAND2_16302 ( P2_R1269_U181 , P2_R1269_U180 , P2_R1269_U179 );
nand NAND2_16303 ( P2_R1269_U182 , P2_U3131 , P2_R1269_U38 );
nand NAND2_16304 ( P2_R1269_U183 , P2_U3132 , P2_R1269_U43 );
nand NAND2_16305 ( P2_R1269_U184 , P2_R1269_U88 , P2_R1269_U6 );
nand NAND2_16306 ( P2_R1269_U185 , P2_R1269_U86 , P2_R1269_U132 );
nand NAND2_16307 ( P2_R1269_U186 , P2_R1269_U87 , P2_R1269_U7 );
nand NAND2_16308 ( P2_R1269_U187 , P2_R1269_U8 , P2_R1269_U184 );
nand NAND3_16309 ( P2_R1269_U188 , P2_R1269_U181 , P2_R1269_U138 , P2_R1269_U8 );
nand NAND2_16310 ( P2_R1269_U189 , P2_U3126 , P2_R1269_U31 );
nand NAND2_16311 ( P2_R1269_U190 , P2_U3125 , P2_R1269_U74 );
nand NAND5_16312 ( P2_R1269_U191 , P2_R1269_U188 , P2_R1269_U187 , P2_R1269_U111 , P2_R1269_U110 , P2_R1269_U140 );
nand NAND2_16313 ( P2_R1269_U192 , P2_R1269_U112 , P2_R1269_U139 );
nand NAND2_16314 ( P2_R1269_U193 , P2_U3092 , P2_R1269_U29 );
nand NAND2_16315 ( P2_R1269_U194 , P2_R1269_U193 , P2_R1269_U192 );
nand NAND2_16316 ( P2_R1269_U195 , P2_R1269_U194 , P2_R1269_U140 );
nand NAND2_16317 ( P2_R1269_U196 , P2_U3090 , P2_R1269_U81 );
nand NAND2_16318 ( P2_R1269_U197 , P2_U3091 , P2_R1269_U30 );
nand NAND2_16319 ( P2_R1269_U198 , P2_U3117 , P2_R1269_U122 );
nand NAND2_16320 ( P2_R1269_U199 , P2_R1269_U122 , P2_R1269_U23 );
nand NAND2_16321 ( P2_R1269_U200 , P2_R1269_U14 , P2_R1269_U121 );
nand NAND2_16322 ( P2_R1269_U201 , P2_R1269_U16 , P2_R1269_U121 );
nand NAND2_16323 ( P2_R1269_U202 , P2_R1269_U17 , P2_R1269_U121 );
nand NAND2_16324 ( P2_R1269_U203 , P2_R1269_U18 , P2_R1269_U121 );
nand NAND2_16325 ( P2_R1269_U204 , P2_R1269_U19 , P2_R1269_U121 );
nand NAND2_16326 ( P2_R1269_U205 , P2_U3116 , P2_U3084 );
nand NAND2_16327 ( P2_R1269_U206 , P2_U3084 , P2_R1269_U25 );
nand NAND2_16328 ( P2_R1269_U207 , P2_U3116 , P2_R1269_U24 );
or OR2_16329 ( P2_R1269_U208 , P2_U3149 , P2_U3116 );
nand NAND2_16330 ( P2_R1269_U209 , P2_U3149 , P2_R1269_U24 );
and AND2_16331 ( P2_R1110_U4 , P2_R1110_U179 , P2_R1110_U178 );
and AND2_16332 ( P2_R1110_U5 , P2_R1110_U197 , P2_R1110_U196 );
and AND2_16333 ( P2_R1110_U6 , P2_R1110_U237 , P2_R1110_U236 );
and AND2_16334 ( P2_R1110_U7 , P2_R1110_U246 , P2_R1110_U245 );
and AND2_16335 ( P2_R1110_U8 , P2_R1110_U264 , P2_R1110_U263 );
and AND2_16336 ( P2_R1110_U9 , P2_R1110_U272 , P2_R1110_U271 );
and AND2_16337 ( P2_R1110_U10 , P2_R1110_U351 , P2_R1110_U348 );
and AND2_16338 ( P2_R1110_U11 , P2_R1110_U344 , P2_R1110_U341 );
and AND2_16339 ( P2_R1110_U12 , P2_R1110_U335 , P2_R1110_U332 );
and AND2_16340 ( P2_R1110_U13 , P2_R1110_U326 , P2_R1110_U323 );
and AND2_16341 ( P2_R1110_U14 , P2_R1110_U320 , P2_R1110_U318 );
and AND2_16342 ( P2_R1110_U15 , P2_R1110_U313 , P2_R1110_U310 );
and AND2_16343 ( P2_R1110_U16 , P2_R1110_U235 , P2_R1110_U232 );
and AND2_16344 ( P2_R1110_U17 , P2_R1110_U227 , P2_R1110_U224 );
and AND2_16345 ( P2_R1110_U18 , P2_R1110_U213 , P2_R1110_U210 );
not NOT1_16346 ( P2_R1110_U19 , P2_U3407 );
not NOT1_16347 ( P2_R1110_U20 , P2_U3070 );
not NOT1_16348 ( P2_R1110_U21 , P2_U3069 );
nand NAND2_16349 ( P2_R1110_U22 , P2_U3070 , P2_U3407 );
not NOT1_16350 ( P2_R1110_U23 , P2_U3410 );
not NOT1_16351 ( P2_R1110_U24 , P2_U3401 );
not NOT1_16352 ( P2_R1110_U25 , P2_U3059 );
not NOT1_16353 ( P2_R1110_U26 , P2_U3066 );
not NOT1_16354 ( P2_R1110_U27 , P2_U3395 );
not NOT1_16355 ( P2_R1110_U28 , P2_U3067 );
not NOT1_16356 ( P2_R1110_U29 , P2_U3387 );
not NOT1_16357 ( P2_R1110_U30 , P2_U3076 );
nand NAND2_16358 ( P2_R1110_U31 , P2_U3076 , P2_U3387 );
not NOT1_16359 ( P2_R1110_U32 , P2_U3398 );
not NOT1_16360 ( P2_R1110_U33 , P2_U3063 );
nand NAND2_16361 ( P2_R1110_U34 , P2_U3059 , P2_U3401 );
not NOT1_16362 ( P2_R1110_U35 , P2_U3404 );
not NOT1_16363 ( P2_R1110_U36 , P2_U3413 );
not NOT1_16364 ( P2_R1110_U37 , P2_U3083 );
not NOT1_16365 ( P2_R1110_U38 , P2_U3082 );
not NOT1_16366 ( P2_R1110_U39 , P2_U3416 );
nand NAND2_16367 ( P2_R1110_U40 , P2_R1110_U65 , P2_R1110_U205 );
nand NAND2_16368 ( P2_R1110_U41 , P2_R1110_U117 , P2_R1110_U193 );
nand NAND2_16369 ( P2_R1110_U42 , P2_R1110_U182 , P2_R1110_U183 );
nand NAND2_16370 ( P2_R1110_U43 , P2_U3392 , P2_U3077 );
nand NAND2_16371 ( P2_R1110_U44 , P2_R1110_U122 , P2_R1110_U219 );
nand NAND2_16372 ( P2_R1110_U45 , P2_R1110_U216 , P2_R1110_U215 );
not NOT1_16373 ( P2_R1110_U46 , P2_U3896 );
not NOT1_16374 ( P2_R1110_U47 , P2_U3052 );
not NOT1_16375 ( P2_R1110_U48 , P2_U3056 );
not NOT1_16376 ( P2_R1110_U49 , P2_U3897 );
not NOT1_16377 ( P2_R1110_U50 , P2_U3898 );
not NOT1_16378 ( P2_R1110_U51 , P2_U3057 );
not NOT1_16379 ( P2_R1110_U52 , P2_U3899 );
not NOT1_16380 ( P2_R1110_U53 , P2_U3064 );
not NOT1_16381 ( P2_R1110_U54 , P2_U3902 );
not NOT1_16382 ( P2_R1110_U55 , P2_U3074 );
not NOT1_16383 ( P2_R1110_U56 , P2_U3437 );
not NOT1_16384 ( P2_R1110_U57 , P2_U3072 );
not NOT1_16385 ( P2_R1110_U58 , P2_U3068 );
nand NAND2_16386 ( P2_R1110_U59 , P2_U3072 , P2_U3437 );
not NOT1_16387 ( P2_R1110_U60 , P2_U3440 );
not NOT1_16388 ( P2_R1110_U61 , P2_U3428 );
not NOT1_16389 ( P2_R1110_U62 , P2_U3079 );
not NOT1_16390 ( P2_R1110_U63 , P2_U3419 );
not NOT1_16391 ( P2_R1110_U64 , P2_U3061 );
nand NAND2_16392 ( P2_R1110_U65 , P2_U3083 , P2_U3413 );
not NOT1_16393 ( P2_R1110_U66 , P2_U3422 );
not NOT1_16394 ( P2_R1110_U67 , P2_U3062 );
nand NAND2_16395 ( P2_R1110_U68 , P2_U3062 , P2_U3422 );
not NOT1_16396 ( P2_R1110_U69 , P2_U3425 );
not NOT1_16397 ( P2_R1110_U70 , P2_U3071 );
not NOT1_16398 ( P2_R1110_U71 , P2_U3431 );
not NOT1_16399 ( P2_R1110_U72 , P2_U3078 );
not NOT1_16400 ( P2_R1110_U73 , P2_U3434 );
not NOT1_16401 ( P2_R1110_U74 , P2_U3073 );
not NOT1_16402 ( P2_R1110_U75 , P2_U3443 );
not NOT1_16403 ( P2_R1110_U76 , P2_U3081 );
nand NAND2_16404 ( P2_R1110_U77 , P2_U3081 , P2_U3443 );
not NOT1_16405 ( P2_R1110_U78 , P2_U3445 );
not NOT1_16406 ( P2_R1110_U79 , P2_U3080 );
nand NAND2_16407 ( P2_R1110_U80 , P2_U3080 , P2_U3445 );
not NOT1_16408 ( P2_R1110_U81 , P2_U3903 );
not NOT1_16409 ( P2_R1110_U82 , P2_U3901 );
not NOT1_16410 ( P2_R1110_U83 , P2_U3060 );
not NOT1_16411 ( P2_R1110_U84 , P2_U3900 );
not NOT1_16412 ( P2_R1110_U85 , P2_U3065 );
nand NAND2_16413 ( P2_R1110_U86 , P2_U3897 , P2_U3056 );
not NOT1_16414 ( P2_R1110_U87 , P2_U3053 );
not NOT1_16415 ( P2_R1110_U88 , P2_U3895 );
nand NAND2_16416 ( P2_R1110_U89 , P2_R1110_U306 , P2_R1110_U176 );
not NOT1_16417 ( P2_R1110_U90 , P2_U3075 );
nand NAND2_16418 ( P2_R1110_U91 , P2_R1110_U77 , P2_R1110_U315 );
nand NAND2_16419 ( P2_R1110_U92 , P2_R1110_U261 , P2_R1110_U260 );
nand NAND2_16420 ( P2_R1110_U93 , P2_R1110_U68 , P2_R1110_U337 );
nand NAND2_16421 ( P2_R1110_U94 , P2_R1110_U457 , P2_R1110_U456 );
nand NAND2_16422 ( P2_R1110_U95 , P2_R1110_U504 , P2_R1110_U503 );
nand NAND2_16423 ( P2_R1110_U96 , P2_R1110_U375 , P2_R1110_U374 );
nand NAND2_16424 ( P2_R1110_U97 , P2_R1110_U380 , P2_R1110_U379 );
nand NAND2_16425 ( P2_R1110_U98 , P2_R1110_U387 , P2_R1110_U386 );
nand NAND2_16426 ( P2_R1110_U99 , P2_R1110_U394 , P2_R1110_U393 );
nand NAND2_16427 ( P2_R1110_U100 , P2_R1110_U399 , P2_R1110_U398 );
nand NAND2_16428 ( P2_R1110_U101 , P2_R1110_U408 , P2_R1110_U407 );
nand NAND2_16429 ( P2_R1110_U102 , P2_R1110_U415 , P2_R1110_U414 );
nand NAND2_16430 ( P2_R1110_U103 , P2_R1110_U422 , P2_R1110_U421 );
nand NAND2_16431 ( P2_R1110_U104 , P2_R1110_U429 , P2_R1110_U428 );
nand NAND2_16432 ( P2_R1110_U105 , P2_R1110_U434 , P2_R1110_U433 );
nand NAND2_16433 ( P2_R1110_U106 , P2_R1110_U441 , P2_R1110_U440 );
nand NAND2_16434 ( P2_R1110_U107 , P2_R1110_U448 , P2_R1110_U447 );
nand NAND2_16435 ( P2_R1110_U108 , P2_R1110_U462 , P2_R1110_U461 );
nand NAND2_16436 ( P2_R1110_U109 , P2_R1110_U467 , P2_R1110_U466 );
nand NAND2_16437 ( P2_R1110_U110 , P2_R1110_U474 , P2_R1110_U473 );
nand NAND2_16438 ( P2_R1110_U111 , P2_R1110_U481 , P2_R1110_U480 );
nand NAND2_16439 ( P2_R1110_U112 , P2_R1110_U488 , P2_R1110_U487 );
nand NAND2_16440 ( P2_R1110_U113 , P2_R1110_U495 , P2_R1110_U494 );
nand NAND2_16441 ( P2_R1110_U114 , P2_R1110_U500 , P2_R1110_U499 );
and AND2_16442 ( P2_R1110_U115 , P2_R1110_U189 , P2_R1110_U187 );
and AND2_16443 ( P2_R1110_U116 , P2_R1110_U4 , P2_R1110_U180 );
and AND2_16444 ( P2_R1110_U117 , P2_R1110_U194 , P2_R1110_U192 );
and AND2_16445 ( P2_R1110_U118 , P2_R1110_U201 , P2_R1110_U200 );
and AND3_16446 ( P2_R1110_U119 , P2_R1110_U382 , P2_R1110_U381 , P2_R1110_U22 );
and AND2_16447 ( P2_R1110_U120 , P2_R1110_U212 , P2_R1110_U5 );
and AND2_16448 ( P2_R1110_U121 , P2_R1110_U181 , P2_R1110_U180 );
and AND2_16449 ( P2_R1110_U122 , P2_R1110_U220 , P2_R1110_U218 );
and AND3_16450 ( P2_R1110_U123 , P2_R1110_U389 , P2_R1110_U388 , P2_R1110_U34 );
and AND2_16451 ( P2_R1110_U124 , P2_R1110_U226 , P2_R1110_U4 );
and AND2_16452 ( P2_R1110_U125 , P2_R1110_U234 , P2_R1110_U181 );
and AND2_16453 ( P2_R1110_U126 , P2_R1110_U204 , P2_R1110_U6 );
and AND2_16454 ( P2_R1110_U127 , P2_R1110_U243 , P2_R1110_U239 );
and AND2_16455 ( P2_R1110_U128 , P2_R1110_U250 , P2_R1110_U7 );
and AND2_16456 ( P2_R1110_U129 , P2_R1110_U253 , P2_R1110_U248 );
and AND2_16457 ( P2_R1110_U130 , P2_R1110_U268 , P2_R1110_U267 );
and AND2_16458 ( P2_R1110_U131 , P2_R1110_U9 , P2_R1110_U282 );
and AND2_16459 ( P2_R1110_U132 , P2_R1110_U285 , P2_R1110_U280 );
and AND2_16460 ( P2_R1110_U133 , P2_R1110_U301 , P2_R1110_U298 );
and AND2_16461 ( P2_R1110_U134 , P2_R1110_U368 , P2_R1110_U302 );
and AND2_16462 ( P2_R1110_U135 , P2_R1110_U160 , P2_R1110_U278 );
and AND3_16463 ( P2_R1110_U136 , P2_R1110_U455 , P2_R1110_U454 , P2_R1110_U80 );
and AND2_16464 ( P2_R1110_U137 , P2_R1110_U325 , P2_R1110_U9 );
and AND3_16465 ( P2_R1110_U138 , P2_R1110_U469 , P2_R1110_U468 , P2_R1110_U59 );
and AND2_16466 ( P2_R1110_U139 , P2_R1110_U334 , P2_R1110_U8 );
and AND3_16467 ( P2_R1110_U140 , P2_R1110_U490 , P2_R1110_U489 , P2_R1110_U172 );
and AND2_16468 ( P2_R1110_U141 , P2_R1110_U343 , P2_R1110_U7 );
and AND3_16469 ( P2_R1110_U142 , P2_R1110_U502 , P2_R1110_U501 , P2_R1110_U171 );
and AND2_16470 ( P2_R1110_U143 , P2_R1110_U350 , P2_R1110_U6 );
nand NAND2_16471 ( P2_R1110_U144 , P2_R1110_U118 , P2_R1110_U202 );
nand NAND2_16472 ( P2_R1110_U145 , P2_R1110_U217 , P2_R1110_U229 );
not NOT1_16473 ( P2_R1110_U146 , P2_U3054 );
not NOT1_16474 ( P2_R1110_U147 , P2_U3904 );
and AND2_16475 ( P2_R1110_U148 , P2_R1110_U403 , P2_R1110_U402 );
nand NAND3_16476 ( P2_R1110_U149 , P2_R1110_U304 , P2_R1110_U169 , P2_R1110_U364 );
and AND2_16477 ( P2_R1110_U150 , P2_R1110_U410 , P2_R1110_U409 );
nand NAND3_16478 ( P2_R1110_U151 , P2_R1110_U370 , P2_R1110_U369 , P2_R1110_U134 );
and AND2_16479 ( P2_R1110_U152 , P2_R1110_U417 , P2_R1110_U416 );
nand NAND3_16480 ( P2_R1110_U153 , P2_R1110_U365 , P2_R1110_U299 , P2_R1110_U86 );
and AND2_16481 ( P2_R1110_U154 , P2_R1110_U424 , P2_R1110_U423 );
nand NAND2_16482 ( P2_R1110_U155 , P2_R1110_U293 , P2_R1110_U292 );
and AND2_16483 ( P2_R1110_U156 , P2_R1110_U436 , P2_R1110_U435 );
nand NAND2_16484 ( P2_R1110_U157 , P2_R1110_U289 , P2_R1110_U288 );
and AND2_16485 ( P2_R1110_U158 , P2_R1110_U443 , P2_R1110_U442 );
nand NAND2_16486 ( P2_R1110_U159 , P2_R1110_U132 , P2_R1110_U284 );
and AND2_16487 ( P2_R1110_U160 , P2_R1110_U450 , P2_R1110_U449 );
nand NAND2_16488 ( P2_R1110_U161 , P2_R1110_U43 , P2_R1110_U327 );
nand NAND2_16489 ( P2_R1110_U162 , P2_R1110_U130 , P2_R1110_U269 );
and AND2_16490 ( P2_R1110_U163 , P2_R1110_U476 , P2_R1110_U475 );
nand NAND2_16491 ( P2_R1110_U164 , P2_R1110_U257 , P2_R1110_U256 );
and AND2_16492 ( P2_R1110_U165 , P2_R1110_U483 , P2_R1110_U482 );
nand NAND2_16493 ( P2_R1110_U166 , P2_R1110_U129 , P2_R1110_U252 );
nand NAND2_16494 ( P2_R1110_U167 , P2_R1110_U127 , P2_R1110_U242 );
nand NAND2_16495 ( P2_R1110_U168 , P2_R1110_U367 , P2_R1110_U366 );
nand NAND2_16496 ( P2_R1110_U169 , P2_U3053 , P2_R1110_U151 );
not NOT1_16497 ( P2_R1110_U170 , P2_R1110_U34 );
nand NAND2_16498 ( P2_R1110_U171 , P2_U3416 , P2_U3082 );
nand NAND2_16499 ( P2_R1110_U172 , P2_U3071 , P2_U3425 );
nand NAND2_16500 ( P2_R1110_U173 , P2_U3057 , P2_U3898 );
not NOT1_16501 ( P2_R1110_U174 , P2_R1110_U68 );
not NOT1_16502 ( P2_R1110_U175 , P2_R1110_U77 );
nand NAND2_16503 ( P2_R1110_U176 , P2_U3064 , P2_U3899 );
not NOT1_16504 ( P2_R1110_U177 , P2_R1110_U65 );
or OR2_16505 ( P2_R1110_U178 , P2_U3066 , P2_U3404 );
or OR2_16506 ( P2_R1110_U179 , P2_U3059 , P2_U3401 );
or OR2_16507 ( P2_R1110_U180 , P2_U3398 , P2_U3063 );
or OR2_16508 ( P2_R1110_U181 , P2_U3395 , P2_U3067 );
not NOT1_16509 ( P2_R1110_U182 , P2_R1110_U31 );
or OR2_16510 ( P2_R1110_U183 , P2_U3392 , P2_U3077 );
not NOT1_16511 ( P2_R1110_U184 , P2_R1110_U42 );
not NOT1_16512 ( P2_R1110_U185 , P2_R1110_U43 );
nand NAND2_16513 ( P2_R1110_U186 , P2_R1110_U42 , P2_R1110_U43 );
nand NAND2_16514 ( P2_R1110_U187 , P2_U3067 , P2_U3395 );
nand NAND2_16515 ( P2_R1110_U188 , P2_R1110_U186 , P2_R1110_U181 );
nand NAND2_16516 ( P2_R1110_U189 , P2_U3063 , P2_U3398 );
nand NAND2_16517 ( P2_R1110_U190 , P2_R1110_U115 , P2_R1110_U188 );
nand NAND2_16518 ( P2_R1110_U191 , P2_R1110_U35 , P2_R1110_U34 );
nand NAND2_16519 ( P2_R1110_U192 , P2_U3066 , P2_R1110_U191 );
nand NAND2_16520 ( P2_R1110_U193 , P2_R1110_U116 , P2_R1110_U190 );
nand NAND2_16521 ( P2_R1110_U194 , P2_U3404 , P2_R1110_U170 );
not NOT1_16522 ( P2_R1110_U195 , P2_R1110_U41 );
or OR2_16523 ( P2_R1110_U196 , P2_U3069 , P2_U3410 );
or OR2_16524 ( P2_R1110_U197 , P2_U3070 , P2_U3407 );
not NOT1_16525 ( P2_R1110_U198 , P2_R1110_U22 );
nand NAND2_16526 ( P2_R1110_U199 , P2_R1110_U23 , P2_R1110_U22 );
nand NAND2_16527 ( P2_R1110_U200 , P2_U3069 , P2_R1110_U199 );
nand NAND2_16528 ( P2_R1110_U201 , P2_U3410 , P2_R1110_U198 );
nand NAND2_16529 ( P2_R1110_U202 , P2_R1110_U5 , P2_R1110_U41 );
not NOT1_16530 ( P2_R1110_U203 , P2_R1110_U144 );
or OR2_16531 ( P2_R1110_U204 , P2_U3413 , P2_U3083 );
nand NAND2_16532 ( P2_R1110_U205 , P2_R1110_U204 , P2_R1110_U144 );
not NOT1_16533 ( P2_R1110_U206 , P2_R1110_U40 );
or OR2_16534 ( P2_R1110_U207 , P2_U3082 , P2_U3416 );
or OR2_16535 ( P2_R1110_U208 , P2_U3407 , P2_U3070 );
nand NAND2_16536 ( P2_R1110_U209 , P2_R1110_U208 , P2_R1110_U41 );
nand NAND2_16537 ( P2_R1110_U210 , P2_R1110_U119 , P2_R1110_U209 );
nand NAND2_16538 ( P2_R1110_U211 , P2_R1110_U195 , P2_R1110_U22 );
nand NAND2_16539 ( P2_R1110_U212 , P2_U3410 , P2_U3069 );
nand NAND2_16540 ( P2_R1110_U213 , P2_R1110_U120 , P2_R1110_U211 );
or OR2_16541 ( P2_R1110_U214 , P2_U3070 , P2_U3407 );
nand NAND2_16542 ( P2_R1110_U215 , P2_R1110_U185 , P2_R1110_U181 );
nand NAND2_16543 ( P2_R1110_U216 , P2_U3067 , P2_U3395 );
not NOT1_16544 ( P2_R1110_U217 , P2_R1110_U45 );
nand NAND2_16545 ( P2_R1110_U218 , P2_R1110_U121 , P2_R1110_U184 );
nand NAND2_16546 ( P2_R1110_U219 , P2_R1110_U45 , P2_R1110_U180 );
nand NAND2_16547 ( P2_R1110_U220 , P2_U3063 , P2_U3398 );
not NOT1_16548 ( P2_R1110_U221 , P2_R1110_U44 );
or OR2_16549 ( P2_R1110_U222 , P2_U3401 , P2_U3059 );
nand NAND2_16550 ( P2_R1110_U223 , P2_R1110_U222 , P2_R1110_U44 );
nand NAND2_16551 ( P2_R1110_U224 , P2_R1110_U123 , P2_R1110_U223 );
nand NAND2_16552 ( P2_R1110_U225 , P2_R1110_U221 , P2_R1110_U34 );
nand NAND2_16553 ( P2_R1110_U226 , P2_U3404 , P2_U3066 );
nand NAND2_16554 ( P2_R1110_U227 , P2_R1110_U124 , P2_R1110_U225 );
or OR2_16555 ( P2_R1110_U228 , P2_U3059 , P2_U3401 );
nand NAND2_16556 ( P2_R1110_U229 , P2_R1110_U184 , P2_R1110_U181 );
not NOT1_16557 ( P2_R1110_U230 , P2_R1110_U145 );
nand NAND2_16558 ( P2_R1110_U231 , P2_U3063 , P2_U3398 );
nand NAND4_16559 ( P2_R1110_U232 , P2_R1110_U401 , P2_R1110_U400 , P2_R1110_U43 , P2_R1110_U42 );
nand NAND2_16560 ( P2_R1110_U233 , P2_R1110_U43 , P2_R1110_U42 );
nand NAND2_16561 ( P2_R1110_U234 , P2_U3067 , P2_U3395 );
nand NAND2_16562 ( P2_R1110_U235 , P2_R1110_U125 , P2_R1110_U233 );
or OR2_16563 ( P2_R1110_U236 , P2_U3082 , P2_U3416 );
or OR2_16564 ( P2_R1110_U237 , P2_U3061 , P2_U3419 );
nand NAND2_16565 ( P2_R1110_U238 , P2_R1110_U177 , P2_R1110_U6 );
nand NAND2_16566 ( P2_R1110_U239 , P2_U3061 , P2_U3419 );
nand NAND2_16567 ( P2_R1110_U240 , P2_R1110_U171 , P2_R1110_U238 );
or OR2_16568 ( P2_R1110_U241 , P2_U3419 , P2_U3061 );
nand NAND2_16569 ( P2_R1110_U242 , P2_R1110_U126 , P2_R1110_U144 );
nand NAND2_16570 ( P2_R1110_U243 , P2_R1110_U241 , P2_R1110_U240 );
not NOT1_16571 ( P2_R1110_U244 , P2_R1110_U167 );
or OR2_16572 ( P2_R1110_U245 , P2_U3079 , P2_U3428 );
or OR2_16573 ( P2_R1110_U246 , P2_U3071 , P2_U3425 );
nand NAND2_16574 ( P2_R1110_U247 , P2_R1110_U174 , P2_R1110_U7 );
nand NAND2_16575 ( P2_R1110_U248 , P2_U3079 , P2_U3428 );
nand NAND2_16576 ( P2_R1110_U249 , P2_R1110_U172 , P2_R1110_U247 );
or OR2_16577 ( P2_R1110_U250 , P2_U3422 , P2_U3062 );
or OR2_16578 ( P2_R1110_U251 , P2_U3428 , P2_U3079 );
nand NAND2_16579 ( P2_R1110_U252 , P2_R1110_U128 , P2_R1110_U167 );
nand NAND2_16580 ( P2_R1110_U253 , P2_R1110_U251 , P2_R1110_U249 );
not NOT1_16581 ( P2_R1110_U254 , P2_R1110_U166 );
or OR2_16582 ( P2_R1110_U255 , P2_U3431 , P2_U3078 );
nand NAND2_16583 ( P2_R1110_U256 , P2_R1110_U255 , P2_R1110_U166 );
nand NAND2_16584 ( P2_R1110_U257 , P2_U3078 , P2_U3431 );
not NOT1_16585 ( P2_R1110_U258 , P2_R1110_U164 );
or OR2_16586 ( P2_R1110_U259 , P2_U3434 , P2_U3073 );
nand NAND2_16587 ( P2_R1110_U260 , P2_R1110_U259 , P2_R1110_U164 );
nand NAND2_16588 ( P2_R1110_U261 , P2_U3073 , P2_U3434 );
not NOT1_16589 ( P2_R1110_U262 , P2_R1110_U92 );
or OR2_16590 ( P2_R1110_U263 , P2_U3068 , P2_U3440 );
or OR2_16591 ( P2_R1110_U264 , P2_U3072 , P2_U3437 );
not NOT1_16592 ( P2_R1110_U265 , P2_R1110_U59 );
nand NAND2_16593 ( P2_R1110_U266 , P2_R1110_U60 , P2_R1110_U59 );
nand NAND2_16594 ( P2_R1110_U267 , P2_U3068 , P2_R1110_U266 );
nand NAND2_16595 ( P2_R1110_U268 , P2_U3440 , P2_R1110_U265 );
nand NAND2_16596 ( P2_R1110_U269 , P2_R1110_U8 , P2_R1110_U92 );
not NOT1_16597 ( P2_R1110_U270 , P2_R1110_U162 );
or OR2_16598 ( P2_R1110_U271 , P2_U3075 , P2_U3903 );
or OR2_16599 ( P2_R1110_U272 , P2_U3080 , P2_U3445 );
or OR2_16600 ( P2_R1110_U273 , P2_U3074 , P2_U3902 );
not NOT1_16601 ( P2_R1110_U274 , P2_R1110_U80 );
nand NAND2_16602 ( P2_R1110_U275 , P2_U3903 , P2_R1110_U274 );
nand NAND2_16603 ( P2_R1110_U276 , P2_R1110_U275 , P2_R1110_U90 );
nand NAND2_16604 ( P2_R1110_U277 , P2_R1110_U80 , P2_R1110_U81 );
nand NAND2_16605 ( P2_R1110_U278 , P2_R1110_U277 , P2_R1110_U276 );
nand NAND2_16606 ( P2_R1110_U279 , P2_R1110_U175 , P2_R1110_U9 );
nand NAND2_16607 ( P2_R1110_U280 , P2_U3074 , P2_U3902 );
nand NAND2_16608 ( P2_R1110_U281 , P2_R1110_U278 , P2_R1110_U279 );
or OR2_16609 ( P2_R1110_U282 , P2_U3443 , P2_U3081 );
or OR2_16610 ( P2_R1110_U283 , P2_U3902 , P2_U3074 );
nand NAND3_16611 ( P2_R1110_U284 , P2_R1110_U273 , P2_R1110_U162 , P2_R1110_U131 );
nand NAND2_16612 ( P2_R1110_U285 , P2_R1110_U283 , P2_R1110_U281 );
not NOT1_16613 ( P2_R1110_U286 , P2_R1110_U159 );
or OR2_16614 ( P2_R1110_U287 , P2_U3901 , P2_U3060 );
nand NAND2_16615 ( P2_R1110_U288 , P2_R1110_U287 , P2_R1110_U159 );
nand NAND2_16616 ( P2_R1110_U289 , P2_U3060 , P2_U3901 );
not NOT1_16617 ( P2_R1110_U290 , P2_R1110_U157 );
or OR2_16618 ( P2_R1110_U291 , P2_U3900 , P2_U3065 );
nand NAND2_16619 ( P2_R1110_U292 , P2_R1110_U291 , P2_R1110_U157 );
nand NAND2_16620 ( P2_R1110_U293 , P2_U3065 , P2_U3900 );
not NOT1_16621 ( P2_R1110_U294 , P2_R1110_U155 );
or OR2_16622 ( P2_R1110_U295 , P2_U3057 , P2_U3898 );
nand NAND2_16623 ( P2_R1110_U296 , P2_R1110_U176 , P2_R1110_U173 );
not NOT1_16624 ( P2_R1110_U297 , P2_R1110_U86 );
or OR2_16625 ( P2_R1110_U298 , P2_U3899 , P2_U3064 );
nand NAND3_16626 ( P2_R1110_U299 , P2_R1110_U155 , P2_R1110_U298 , P2_R1110_U168 );
not NOT1_16627 ( P2_R1110_U300 , P2_R1110_U153 );
or OR2_16628 ( P2_R1110_U301 , P2_U3896 , P2_U3052 );
nand NAND2_16629 ( P2_R1110_U302 , P2_U3052 , P2_U3896 );
not NOT1_16630 ( P2_R1110_U303 , P2_R1110_U151 );
nand NAND2_16631 ( P2_R1110_U304 , P2_U3895 , P2_R1110_U151 );
not NOT1_16632 ( P2_R1110_U305 , P2_R1110_U149 );
nand NAND2_16633 ( P2_R1110_U306 , P2_R1110_U298 , P2_R1110_U155 );
not NOT1_16634 ( P2_R1110_U307 , P2_R1110_U89 );
or OR2_16635 ( P2_R1110_U308 , P2_U3898 , P2_U3057 );
nand NAND2_16636 ( P2_R1110_U309 , P2_R1110_U308 , P2_R1110_U89 );
nand NAND3_16637 ( P2_R1110_U310 , P2_R1110_U309 , P2_R1110_U173 , P2_R1110_U154 );
nand NAND2_16638 ( P2_R1110_U311 , P2_R1110_U307 , P2_R1110_U173 );
nand NAND2_16639 ( P2_R1110_U312 , P2_U3897 , P2_U3056 );
nand NAND3_16640 ( P2_R1110_U313 , P2_R1110_U311 , P2_R1110_U312 , P2_R1110_U168 );
or OR2_16641 ( P2_R1110_U314 , P2_U3057 , P2_U3898 );
nand NAND2_16642 ( P2_R1110_U315 , P2_R1110_U282 , P2_R1110_U162 );
not NOT1_16643 ( P2_R1110_U316 , P2_R1110_U91 );
nand NAND2_16644 ( P2_R1110_U317 , P2_R1110_U9 , P2_R1110_U91 );
nand NAND2_16645 ( P2_R1110_U318 , P2_R1110_U135 , P2_R1110_U317 );
nand NAND2_16646 ( P2_R1110_U319 , P2_R1110_U317 , P2_R1110_U278 );
nand NAND2_16647 ( P2_R1110_U320 , P2_R1110_U453 , P2_R1110_U319 );
or OR2_16648 ( P2_R1110_U321 , P2_U3445 , P2_U3080 );
nand NAND2_16649 ( P2_R1110_U322 , P2_R1110_U321 , P2_R1110_U91 );
nand NAND2_16650 ( P2_R1110_U323 , P2_R1110_U136 , P2_R1110_U322 );
nand NAND2_16651 ( P2_R1110_U324 , P2_R1110_U316 , P2_R1110_U80 );
nand NAND2_16652 ( P2_R1110_U325 , P2_U3075 , P2_U3903 );
nand NAND2_16653 ( P2_R1110_U326 , P2_R1110_U137 , P2_R1110_U324 );
or OR2_16654 ( P2_R1110_U327 , P2_U3392 , P2_U3077 );
not NOT1_16655 ( P2_R1110_U328 , P2_R1110_U161 );
or OR2_16656 ( P2_R1110_U329 , P2_U3080 , P2_U3445 );
or OR2_16657 ( P2_R1110_U330 , P2_U3437 , P2_U3072 );
nand NAND2_16658 ( P2_R1110_U331 , P2_R1110_U330 , P2_R1110_U92 );
nand NAND2_16659 ( P2_R1110_U332 , P2_R1110_U138 , P2_R1110_U331 );
nand NAND2_16660 ( P2_R1110_U333 , P2_R1110_U262 , P2_R1110_U59 );
nand NAND2_16661 ( P2_R1110_U334 , P2_U3440 , P2_U3068 );
nand NAND2_16662 ( P2_R1110_U335 , P2_R1110_U139 , P2_R1110_U333 );
or OR2_16663 ( P2_R1110_U336 , P2_U3072 , P2_U3437 );
nand NAND2_16664 ( P2_R1110_U337 , P2_R1110_U250 , P2_R1110_U167 );
not NOT1_16665 ( P2_R1110_U338 , P2_R1110_U93 );
or OR2_16666 ( P2_R1110_U339 , P2_U3425 , P2_U3071 );
nand NAND2_16667 ( P2_R1110_U340 , P2_R1110_U339 , P2_R1110_U93 );
nand NAND2_16668 ( P2_R1110_U341 , P2_R1110_U140 , P2_R1110_U340 );
nand NAND2_16669 ( P2_R1110_U342 , P2_R1110_U338 , P2_R1110_U172 );
nand NAND2_16670 ( P2_R1110_U343 , P2_U3079 , P2_U3428 );
nand NAND2_16671 ( P2_R1110_U344 , P2_R1110_U141 , P2_R1110_U342 );
or OR2_16672 ( P2_R1110_U345 , P2_U3071 , P2_U3425 );
or OR2_16673 ( P2_R1110_U346 , P2_U3416 , P2_U3082 );
nand NAND2_16674 ( P2_R1110_U347 , P2_R1110_U346 , P2_R1110_U40 );
nand NAND2_16675 ( P2_R1110_U348 , P2_R1110_U142 , P2_R1110_U347 );
nand NAND2_16676 ( P2_R1110_U349 , P2_R1110_U206 , P2_R1110_U171 );
nand NAND2_16677 ( P2_R1110_U350 , P2_U3061 , P2_U3419 );
nand NAND2_16678 ( P2_R1110_U351 , P2_R1110_U143 , P2_R1110_U349 );
nand NAND2_16679 ( P2_R1110_U352 , P2_R1110_U207 , P2_R1110_U171 );
nand NAND2_16680 ( P2_R1110_U353 , P2_R1110_U204 , P2_R1110_U65 );
nand NAND2_16681 ( P2_R1110_U354 , P2_R1110_U214 , P2_R1110_U22 );
nand NAND2_16682 ( P2_R1110_U355 , P2_R1110_U228 , P2_R1110_U34 );
nand NAND2_16683 ( P2_R1110_U356 , P2_R1110_U231 , P2_R1110_U180 );
nand NAND2_16684 ( P2_R1110_U357 , P2_R1110_U314 , P2_R1110_U173 );
nand NAND2_16685 ( P2_R1110_U358 , P2_R1110_U298 , P2_R1110_U176 );
nand NAND2_16686 ( P2_R1110_U359 , P2_R1110_U329 , P2_R1110_U80 );
nand NAND2_16687 ( P2_R1110_U360 , P2_R1110_U282 , P2_R1110_U77 );
nand NAND2_16688 ( P2_R1110_U361 , P2_R1110_U336 , P2_R1110_U59 );
nand NAND2_16689 ( P2_R1110_U362 , P2_R1110_U345 , P2_R1110_U172 );
nand NAND2_16690 ( P2_R1110_U363 , P2_R1110_U250 , P2_R1110_U68 );
nand NAND2_16691 ( P2_R1110_U364 , P2_U3895 , P2_U3053 );
nand NAND2_16692 ( P2_R1110_U365 , P2_R1110_U296 , P2_R1110_U168 );
nand NAND2_16693 ( P2_R1110_U366 , P2_U3056 , P2_R1110_U295 );
nand NAND2_16694 ( P2_R1110_U367 , P2_U3897 , P2_R1110_U295 );
nand NAND3_16695 ( P2_R1110_U368 , P2_R1110_U296 , P2_R1110_U168 , P2_R1110_U301 );
nand NAND3_16696 ( P2_R1110_U369 , P2_R1110_U155 , P2_R1110_U168 , P2_R1110_U133 );
nand NAND2_16697 ( P2_R1110_U370 , P2_R1110_U297 , P2_R1110_U301 );
nand NAND2_16698 ( P2_R1110_U371 , P2_U3082 , P2_R1110_U39 );
nand NAND2_16699 ( P2_R1110_U372 , P2_U3416 , P2_R1110_U38 );
nand NAND2_16700 ( P2_R1110_U373 , P2_R1110_U372 , P2_R1110_U371 );
nand NAND2_16701 ( P2_R1110_U374 , P2_R1110_U352 , P2_R1110_U40 );
nand NAND2_16702 ( P2_R1110_U375 , P2_R1110_U373 , P2_R1110_U206 );
nand NAND2_16703 ( P2_R1110_U376 , P2_U3083 , P2_R1110_U36 );
nand NAND2_16704 ( P2_R1110_U377 , P2_U3413 , P2_R1110_U37 );
nand NAND2_16705 ( P2_R1110_U378 , P2_R1110_U377 , P2_R1110_U376 );
nand NAND2_16706 ( P2_R1110_U379 , P2_R1110_U353 , P2_R1110_U144 );
nand NAND2_16707 ( P2_R1110_U380 , P2_R1110_U203 , P2_R1110_U378 );
nand NAND2_16708 ( P2_R1110_U381 , P2_U3069 , P2_R1110_U23 );
nand NAND2_16709 ( P2_R1110_U382 , P2_U3410 , P2_R1110_U21 );
nand NAND2_16710 ( P2_R1110_U383 , P2_U3070 , P2_R1110_U19 );
nand NAND2_16711 ( P2_R1110_U384 , P2_U3407 , P2_R1110_U20 );
nand NAND2_16712 ( P2_R1110_U385 , P2_R1110_U384 , P2_R1110_U383 );
nand NAND2_16713 ( P2_R1110_U386 , P2_R1110_U354 , P2_R1110_U41 );
nand NAND2_16714 ( P2_R1110_U387 , P2_R1110_U385 , P2_R1110_U195 );
nand NAND2_16715 ( P2_R1110_U388 , P2_U3066 , P2_R1110_U35 );
nand NAND2_16716 ( P2_R1110_U389 , P2_U3404 , P2_R1110_U26 );
nand NAND2_16717 ( P2_R1110_U390 , P2_U3059 , P2_R1110_U24 );
nand NAND2_16718 ( P2_R1110_U391 , P2_U3401 , P2_R1110_U25 );
nand NAND2_16719 ( P2_R1110_U392 , P2_R1110_U391 , P2_R1110_U390 );
nand NAND2_16720 ( P2_R1110_U393 , P2_R1110_U355 , P2_R1110_U44 );
nand NAND2_16721 ( P2_R1110_U394 , P2_R1110_U392 , P2_R1110_U221 );
nand NAND2_16722 ( P2_R1110_U395 , P2_U3063 , P2_R1110_U32 );
nand NAND2_16723 ( P2_R1110_U396 , P2_U3398 , P2_R1110_U33 );
nand NAND2_16724 ( P2_R1110_U397 , P2_R1110_U396 , P2_R1110_U395 );
nand NAND2_16725 ( P2_R1110_U398 , P2_R1110_U356 , P2_R1110_U145 );
nand NAND2_16726 ( P2_R1110_U399 , P2_R1110_U230 , P2_R1110_U397 );
nand NAND2_16727 ( P2_R1110_U400 , P2_U3067 , P2_R1110_U27 );
nand NAND2_16728 ( P2_R1110_U401 , P2_U3395 , P2_R1110_U28 );
nand NAND2_16729 ( P2_R1110_U402 , P2_U3054 , P2_R1110_U147 );
nand NAND2_16730 ( P2_R1110_U403 , P2_U3904 , P2_R1110_U146 );
nand NAND2_16731 ( P2_R1110_U404 , P2_U3054 , P2_R1110_U147 );
nand NAND2_16732 ( P2_R1110_U405 , P2_U3904 , P2_R1110_U146 );
nand NAND2_16733 ( P2_R1110_U406 , P2_R1110_U405 , P2_R1110_U404 );
nand NAND2_16734 ( P2_R1110_U407 , P2_R1110_U148 , P2_R1110_U149 );
nand NAND2_16735 ( P2_R1110_U408 , P2_R1110_U305 , P2_R1110_U406 );
nand NAND2_16736 ( P2_R1110_U409 , P2_U3053 , P2_R1110_U88 );
nand NAND2_16737 ( P2_R1110_U410 , P2_U3895 , P2_R1110_U87 );
nand NAND2_16738 ( P2_R1110_U411 , P2_U3053 , P2_R1110_U88 );
nand NAND2_16739 ( P2_R1110_U412 , P2_U3895 , P2_R1110_U87 );
nand NAND2_16740 ( P2_R1110_U413 , P2_R1110_U412 , P2_R1110_U411 );
nand NAND2_16741 ( P2_R1110_U414 , P2_R1110_U150 , P2_R1110_U151 );
nand NAND2_16742 ( P2_R1110_U415 , P2_R1110_U303 , P2_R1110_U413 );
nand NAND2_16743 ( P2_R1110_U416 , P2_U3052 , P2_R1110_U46 );
nand NAND2_16744 ( P2_R1110_U417 , P2_U3896 , P2_R1110_U47 );
nand NAND2_16745 ( P2_R1110_U418 , P2_U3052 , P2_R1110_U46 );
nand NAND2_16746 ( P2_R1110_U419 , P2_U3896 , P2_R1110_U47 );
nand NAND2_16747 ( P2_R1110_U420 , P2_R1110_U419 , P2_R1110_U418 );
nand NAND2_16748 ( P2_R1110_U421 , P2_R1110_U152 , P2_R1110_U153 );
nand NAND2_16749 ( P2_R1110_U422 , P2_R1110_U300 , P2_R1110_U420 );
nand NAND2_16750 ( P2_R1110_U423 , P2_U3056 , P2_R1110_U49 );
nand NAND2_16751 ( P2_R1110_U424 , P2_U3897 , P2_R1110_U48 );
nand NAND2_16752 ( P2_R1110_U425 , P2_U3057 , P2_R1110_U50 );
nand NAND2_16753 ( P2_R1110_U426 , P2_U3898 , P2_R1110_U51 );
nand NAND2_16754 ( P2_R1110_U427 , P2_R1110_U426 , P2_R1110_U425 );
nand NAND2_16755 ( P2_R1110_U428 , P2_R1110_U357 , P2_R1110_U89 );
nand NAND2_16756 ( P2_R1110_U429 , P2_R1110_U427 , P2_R1110_U307 );
nand NAND2_16757 ( P2_R1110_U430 , P2_U3064 , P2_R1110_U52 );
nand NAND2_16758 ( P2_R1110_U431 , P2_U3899 , P2_R1110_U53 );
nand NAND2_16759 ( P2_R1110_U432 , P2_R1110_U431 , P2_R1110_U430 );
nand NAND2_16760 ( P2_R1110_U433 , P2_R1110_U358 , P2_R1110_U155 );
nand NAND2_16761 ( P2_R1110_U434 , P2_R1110_U294 , P2_R1110_U432 );
nand NAND2_16762 ( P2_R1110_U435 , P2_U3065 , P2_R1110_U84 );
nand NAND2_16763 ( P2_R1110_U436 , P2_U3900 , P2_R1110_U85 );
nand NAND2_16764 ( P2_R1110_U437 , P2_U3065 , P2_R1110_U84 );
nand NAND2_16765 ( P2_R1110_U438 , P2_U3900 , P2_R1110_U85 );
nand NAND2_16766 ( P2_R1110_U439 , P2_R1110_U438 , P2_R1110_U437 );
nand NAND2_16767 ( P2_R1110_U440 , P2_R1110_U156 , P2_R1110_U157 );
nand NAND2_16768 ( P2_R1110_U441 , P2_R1110_U290 , P2_R1110_U439 );
nand NAND2_16769 ( P2_R1110_U442 , P2_U3060 , P2_R1110_U82 );
nand NAND2_16770 ( P2_R1110_U443 , P2_U3901 , P2_R1110_U83 );
nand NAND2_16771 ( P2_R1110_U444 , P2_U3060 , P2_R1110_U82 );
nand NAND2_16772 ( P2_R1110_U445 , P2_U3901 , P2_R1110_U83 );
nand NAND2_16773 ( P2_R1110_U446 , P2_R1110_U445 , P2_R1110_U444 );
nand NAND2_16774 ( P2_R1110_U447 , P2_R1110_U158 , P2_R1110_U159 );
nand NAND2_16775 ( P2_R1110_U448 , P2_R1110_U286 , P2_R1110_U446 );
nand NAND2_16776 ( P2_R1110_U449 , P2_U3074 , P2_R1110_U54 );
nand NAND2_16777 ( P2_R1110_U450 , P2_U3902 , P2_R1110_U55 );
nand NAND2_16778 ( P2_R1110_U451 , P2_U3074 , P2_R1110_U54 );
nand NAND2_16779 ( P2_R1110_U452 , P2_U3902 , P2_R1110_U55 );
nand NAND2_16780 ( P2_R1110_U453 , P2_R1110_U452 , P2_R1110_U451 );
nand NAND2_16781 ( P2_R1110_U454 , P2_U3075 , P2_R1110_U81 );
nand NAND2_16782 ( P2_R1110_U455 , P2_U3903 , P2_R1110_U90 );
nand NAND2_16783 ( P2_R1110_U456 , P2_R1110_U182 , P2_R1110_U161 );
nand NAND2_16784 ( P2_R1110_U457 , P2_R1110_U328 , P2_R1110_U31 );
nand NAND2_16785 ( P2_R1110_U458 , P2_U3080 , P2_R1110_U78 );
nand NAND2_16786 ( P2_R1110_U459 , P2_U3445 , P2_R1110_U79 );
nand NAND2_16787 ( P2_R1110_U460 , P2_R1110_U459 , P2_R1110_U458 );
nand NAND2_16788 ( P2_R1110_U461 , P2_R1110_U359 , P2_R1110_U91 );
nand NAND2_16789 ( P2_R1110_U462 , P2_R1110_U460 , P2_R1110_U316 );
nand NAND2_16790 ( P2_R1110_U463 , P2_U3081 , P2_R1110_U75 );
nand NAND2_16791 ( P2_R1110_U464 , P2_U3443 , P2_R1110_U76 );
nand NAND2_16792 ( P2_R1110_U465 , P2_R1110_U464 , P2_R1110_U463 );
nand NAND2_16793 ( P2_R1110_U466 , P2_R1110_U360 , P2_R1110_U162 );
nand NAND2_16794 ( P2_R1110_U467 , P2_R1110_U270 , P2_R1110_U465 );
nand NAND2_16795 ( P2_R1110_U468 , P2_U3068 , P2_R1110_U60 );
nand NAND2_16796 ( P2_R1110_U469 , P2_U3440 , P2_R1110_U58 );
nand NAND2_16797 ( P2_R1110_U470 , P2_U3072 , P2_R1110_U56 );
nand NAND2_16798 ( P2_R1110_U471 , P2_U3437 , P2_R1110_U57 );
nand NAND2_16799 ( P2_R1110_U472 , P2_R1110_U471 , P2_R1110_U470 );
nand NAND2_16800 ( P2_R1110_U473 , P2_R1110_U361 , P2_R1110_U92 );
nand NAND2_16801 ( P2_R1110_U474 , P2_R1110_U472 , P2_R1110_U262 );
nand NAND2_16802 ( P2_R1110_U475 , P2_U3073 , P2_R1110_U73 );
nand NAND2_16803 ( P2_R1110_U476 , P2_U3434 , P2_R1110_U74 );
nand NAND2_16804 ( P2_R1110_U477 , P2_U3073 , P2_R1110_U73 );
nand NAND2_16805 ( P2_R1110_U478 , P2_U3434 , P2_R1110_U74 );
nand NAND2_16806 ( P2_R1110_U479 , P2_R1110_U478 , P2_R1110_U477 );
nand NAND2_16807 ( P2_R1110_U480 , P2_R1110_U163 , P2_R1110_U164 );
nand NAND2_16808 ( P2_R1110_U481 , P2_R1110_U258 , P2_R1110_U479 );
nand NAND2_16809 ( P2_R1110_U482 , P2_U3078 , P2_R1110_U71 );
nand NAND2_16810 ( P2_R1110_U483 , P2_U3431 , P2_R1110_U72 );
nand NAND2_16811 ( P2_R1110_U484 , P2_U3078 , P2_R1110_U71 );
nand NAND2_16812 ( P2_R1110_U485 , P2_U3431 , P2_R1110_U72 );
nand NAND2_16813 ( P2_R1110_U486 , P2_R1110_U485 , P2_R1110_U484 );
nand NAND2_16814 ( P2_R1110_U487 , P2_R1110_U165 , P2_R1110_U166 );
nand NAND2_16815 ( P2_R1110_U488 , P2_R1110_U254 , P2_R1110_U486 );
nand NAND2_16816 ( P2_R1110_U489 , P2_U3079 , P2_R1110_U61 );
nand NAND2_16817 ( P2_R1110_U490 , P2_U3428 , P2_R1110_U62 );
nand NAND2_16818 ( P2_R1110_U491 , P2_U3071 , P2_R1110_U69 );
nand NAND2_16819 ( P2_R1110_U492 , P2_U3425 , P2_R1110_U70 );
nand NAND2_16820 ( P2_R1110_U493 , P2_R1110_U492 , P2_R1110_U491 );
nand NAND2_16821 ( P2_R1110_U494 , P2_R1110_U362 , P2_R1110_U93 );
nand NAND2_16822 ( P2_R1110_U495 , P2_R1110_U493 , P2_R1110_U338 );
nand NAND2_16823 ( P2_R1110_U496 , P2_U3062 , P2_R1110_U66 );
nand NAND2_16824 ( P2_R1110_U497 , P2_U3422 , P2_R1110_U67 );
nand NAND2_16825 ( P2_R1110_U498 , P2_R1110_U497 , P2_R1110_U496 );
nand NAND2_16826 ( P2_R1110_U499 , P2_R1110_U363 , P2_R1110_U167 );
nand NAND2_16827 ( P2_R1110_U500 , P2_R1110_U244 , P2_R1110_U498 );
nand NAND2_16828 ( P2_R1110_U501 , P2_U3061 , P2_R1110_U63 );
nand NAND2_16829 ( P2_R1110_U502 , P2_U3419 , P2_R1110_U64 );
nand NAND2_16830 ( P2_R1110_U503 , P2_U3076 , P2_R1110_U29 );
nand NAND2_16831 ( P2_R1110_U504 , P2_U3387 , P2_R1110_U30 );
and AND2_16832 ( P2_R1297_U6 , P2_U3058 , P2_R1297_U7 );
not NOT1_16833 ( P2_R1297_U7 , P2_U3055 );
and AND2_16834 ( P2_R1077_U4 , P2_R1077_U179 , P2_R1077_U178 );
and AND2_16835 ( P2_R1077_U5 , P2_R1077_U197 , P2_R1077_U196 );
and AND2_16836 ( P2_R1077_U6 , P2_R1077_U237 , P2_R1077_U236 );
and AND2_16837 ( P2_R1077_U7 , P2_R1077_U246 , P2_R1077_U245 );
and AND2_16838 ( P2_R1077_U8 , P2_R1077_U264 , P2_R1077_U263 );
and AND2_16839 ( P2_R1077_U9 , P2_R1077_U272 , P2_R1077_U271 );
and AND2_16840 ( P2_R1077_U10 , P2_R1077_U351 , P2_R1077_U348 );
and AND2_16841 ( P2_R1077_U11 , P2_R1077_U344 , P2_R1077_U341 );
and AND2_16842 ( P2_R1077_U12 , P2_R1077_U335 , P2_R1077_U332 );
and AND2_16843 ( P2_R1077_U13 , P2_R1077_U326 , P2_R1077_U323 );
and AND2_16844 ( P2_R1077_U14 , P2_R1077_U320 , P2_R1077_U318 );
and AND2_16845 ( P2_R1077_U15 , P2_R1077_U313 , P2_R1077_U310 );
and AND2_16846 ( P2_R1077_U16 , P2_R1077_U235 , P2_R1077_U232 );
and AND2_16847 ( P2_R1077_U17 , P2_R1077_U227 , P2_R1077_U224 );
and AND2_16848 ( P2_R1077_U18 , P2_R1077_U213 , P2_R1077_U210 );
not NOT1_16849 ( P2_R1077_U19 , P2_U3407 );
not NOT1_16850 ( P2_R1077_U20 , P2_U3070 );
not NOT1_16851 ( P2_R1077_U21 , P2_U3069 );
nand NAND2_16852 ( P2_R1077_U22 , P2_U3070 , P2_U3407 );
not NOT1_16853 ( P2_R1077_U23 , P2_U3410 );
not NOT1_16854 ( P2_R1077_U24 , P2_U3401 );
not NOT1_16855 ( P2_R1077_U25 , P2_U3059 );
not NOT1_16856 ( P2_R1077_U26 , P2_U3066 );
not NOT1_16857 ( P2_R1077_U27 , P2_U3395 );
not NOT1_16858 ( P2_R1077_U28 , P2_U3067 );
not NOT1_16859 ( P2_R1077_U29 , P2_U3387 );
not NOT1_16860 ( P2_R1077_U30 , P2_U3076 );
nand NAND2_16861 ( P2_R1077_U31 , P2_U3076 , P2_U3387 );
not NOT1_16862 ( P2_R1077_U32 , P2_U3398 );
not NOT1_16863 ( P2_R1077_U33 , P2_U3063 );
nand NAND2_16864 ( P2_R1077_U34 , P2_U3059 , P2_U3401 );
not NOT1_16865 ( P2_R1077_U35 , P2_U3404 );
not NOT1_16866 ( P2_R1077_U36 , P2_U3413 );
not NOT1_16867 ( P2_R1077_U37 , P2_U3083 );
not NOT1_16868 ( P2_R1077_U38 , P2_U3082 );
not NOT1_16869 ( P2_R1077_U39 , P2_U3416 );
nand NAND2_16870 ( P2_R1077_U40 , P2_R1077_U65 , P2_R1077_U205 );
nand NAND2_16871 ( P2_R1077_U41 , P2_R1077_U117 , P2_R1077_U193 );
nand NAND2_16872 ( P2_R1077_U42 , P2_R1077_U182 , P2_R1077_U183 );
nand NAND2_16873 ( P2_R1077_U43 , P2_U3392 , P2_U3077 );
nand NAND2_16874 ( P2_R1077_U44 , P2_R1077_U122 , P2_R1077_U219 );
nand NAND2_16875 ( P2_R1077_U45 , P2_R1077_U216 , P2_R1077_U215 );
not NOT1_16876 ( P2_R1077_U46 , P2_U3896 );
not NOT1_16877 ( P2_R1077_U47 , P2_U3052 );
not NOT1_16878 ( P2_R1077_U48 , P2_U3056 );
not NOT1_16879 ( P2_R1077_U49 , P2_U3897 );
not NOT1_16880 ( P2_R1077_U50 , P2_U3898 );
not NOT1_16881 ( P2_R1077_U51 , P2_U3057 );
not NOT1_16882 ( P2_R1077_U52 , P2_U3899 );
not NOT1_16883 ( P2_R1077_U53 , P2_U3064 );
not NOT1_16884 ( P2_R1077_U54 , P2_U3902 );
not NOT1_16885 ( P2_R1077_U55 , P2_U3074 );
not NOT1_16886 ( P2_R1077_U56 , P2_U3437 );
not NOT1_16887 ( P2_R1077_U57 , P2_U3072 );
not NOT1_16888 ( P2_R1077_U58 , P2_U3068 );
nand NAND2_16889 ( P2_R1077_U59 , P2_U3072 , P2_U3437 );
not NOT1_16890 ( P2_R1077_U60 , P2_U3440 );
not NOT1_16891 ( P2_R1077_U61 , P2_U3428 );
not NOT1_16892 ( P2_R1077_U62 , P2_U3079 );
not NOT1_16893 ( P2_R1077_U63 , P2_U3419 );
not NOT1_16894 ( P2_R1077_U64 , P2_U3061 );
nand NAND2_16895 ( P2_R1077_U65 , P2_U3083 , P2_U3413 );
not NOT1_16896 ( P2_R1077_U66 , P2_U3422 );
not NOT1_16897 ( P2_R1077_U67 , P2_U3062 );
nand NAND2_16898 ( P2_R1077_U68 , P2_U3062 , P2_U3422 );
not NOT1_16899 ( P2_R1077_U69 , P2_U3425 );
not NOT1_16900 ( P2_R1077_U70 , P2_U3071 );
not NOT1_16901 ( P2_R1077_U71 , P2_U3431 );
not NOT1_16902 ( P2_R1077_U72 , P2_U3078 );
not NOT1_16903 ( P2_R1077_U73 , P2_U3434 );
not NOT1_16904 ( P2_R1077_U74 , P2_U3073 );
not NOT1_16905 ( P2_R1077_U75 , P2_U3443 );
not NOT1_16906 ( P2_R1077_U76 , P2_U3081 );
nand NAND2_16907 ( P2_R1077_U77 , P2_U3081 , P2_U3443 );
not NOT1_16908 ( P2_R1077_U78 , P2_U3445 );
not NOT1_16909 ( P2_R1077_U79 , P2_U3080 );
nand NAND2_16910 ( P2_R1077_U80 , P2_U3080 , P2_U3445 );
not NOT1_16911 ( P2_R1077_U81 , P2_U3903 );
not NOT1_16912 ( P2_R1077_U82 , P2_U3901 );
not NOT1_16913 ( P2_R1077_U83 , P2_U3060 );
not NOT1_16914 ( P2_R1077_U84 , P2_U3900 );
not NOT1_16915 ( P2_R1077_U85 , P2_U3065 );
nand NAND2_16916 ( P2_R1077_U86 , P2_U3897 , P2_U3056 );
not NOT1_16917 ( P2_R1077_U87 , P2_U3053 );
not NOT1_16918 ( P2_R1077_U88 , P2_U3895 );
nand NAND2_16919 ( P2_R1077_U89 , P2_R1077_U306 , P2_R1077_U176 );
not NOT1_16920 ( P2_R1077_U90 , P2_U3075 );
nand NAND2_16921 ( P2_R1077_U91 , P2_R1077_U77 , P2_R1077_U315 );
nand NAND2_16922 ( P2_R1077_U92 , P2_R1077_U261 , P2_R1077_U260 );
nand NAND2_16923 ( P2_R1077_U93 , P2_R1077_U68 , P2_R1077_U337 );
nand NAND2_16924 ( P2_R1077_U94 , P2_R1077_U457 , P2_R1077_U456 );
nand NAND2_16925 ( P2_R1077_U95 , P2_R1077_U504 , P2_R1077_U503 );
nand NAND2_16926 ( P2_R1077_U96 , P2_R1077_U375 , P2_R1077_U374 );
nand NAND2_16927 ( P2_R1077_U97 , P2_R1077_U380 , P2_R1077_U379 );
nand NAND2_16928 ( P2_R1077_U98 , P2_R1077_U387 , P2_R1077_U386 );
nand NAND2_16929 ( P2_R1077_U99 , P2_R1077_U394 , P2_R1077_U393 );
nand NAND2_16930 ( P2_R1077_U100 , P2_R1077_U399 , P2_R1077_U398 );
nand NAND2_16931 ( P2_R1077_U101 , P2_R1077_U408 , P2_R1077_U407 );
nand NAND2_16932 ( P2_R1077_U102 , P2_R1077_U415 , P2_R1077_U414 );
nand NAND2_16933 ( P2_R1077_U103 , P2_R1077_U422 , P2_R1077_U421 );
nand NAND2_16934 ( P2_R1077_U104 , P2_R1077_U429 , P2_R1077_U428 );
nand NAND2_16935 ( P2_R1077_U105 , P2_R1077_U434 , P2_R1077_U433 );
nand NAND2_16936 ( P2_R1077_U106 , P2_R1077_U441 , P2_R1077_U440 );
nand NAND2_16937 ( P2_R1077_U107 , P2_R1077_U448 , P2_R1077_U447 );
nand NAND2_16938 ( P2_R1077_U108 , P2_R1077_U462 , P2_R1077_U461 );
nand NAND2_16939 ( P2_R1077_U109 , P2_R1077_U467 , P2_R1077_U466 );
nand NAND2_16940 ( P2_R1077_U110 , P2_R1077_U474 , P2_R1077_U473 );
nand NAND2_16941 ( P2_R1077_U111 , P2_R1077_U481 , P2_R1077_U480 );
nand NAND2_16942 ( P2_R1077_U112 , P2_R1077_U488 , P2_R1077_U487 );
nand NAND2_16943 ( P2_R1077_U113 , P2_R1077_U495 , P2_R1077_U494 );
nand NAND2_16944 ( P2_R1077_U114 , P2_R1077_U500 , P2_R1077_U499 );
and AND2_16945 ( P2_R1077_U115 , P2_R1077_U189 , P2_R1077_U187 );
and AND2_16946 ( P2_R1077_U116 , P2_R1077_U4 , P2_R1077_U180 );
and AND2_16947 ( P2_R1077_U117 , P2_R1077_U194 , P2_R1077_U192 );
and AND2_16948 ( P2_R1077_U118 , P2_R1077_U201 , P2_R1077_U200 );
and AND3_16949 ( P2_R1077_U119 , P2_R1077_U382 , P2_R1077_U381 , P2_R1077_U22 );
and AND2_16950 ( P2_R1077_U120 , P2_R1077_U212 , P2_R1077_U5 );
and AND2_16951 ( P2_R1077_U121 , P2_R1077_U181 , P2_R1077_U180 );
and AND2_16952 ( P2_R1077_U122 , P2_R1077_U220 , P2_R1077_U218 );
and AND3_16953 ( P2_R1077_U123 , P2_R1077_U389 , P2_R1077_U388 , P2_R1077_U34 );
and AND2_16954 ( P2_R1077_U124 , P2_R1077_U226 , P2_R1077_U4 );
and AND2_16955 ( P2_R1077_U125 , P2_R1077_U234 , P2_R1077_U181 );
and AND2_16956 ( P2_R1077_U126 , P2_R1077_U204 , P2_R1077_U6 );
and AND2_16957 ( P2_R1077_U127 , P2_R1077_U243 , P2_R1077_U239 );
and AND2_16958 ( P2_R1077_U128 , P2_R1077_U250 , P2_R1077_U7 );
and AND2_16959 ( P2_R1077_U129 , P2_R1077_U253 , P2_R1077_U248 );
and AND2_16960 ( P2_R1077_U130 , P2_R1077_U268 , P2_R1077_U267 );
and AND2_16961 ( P2_R1077_U131 , P2_R1077_U9 , P2_R1077_U282 );
and AND2_16962 ( P2_R1077_U132 , P2_R1077_U285 , P2_R1077_U280 );
and AND2_16963 ( P2_R1077_U133 , P2_R1077_U301 , P2_R1077_U298 );
and AND2_16964 ( P2_R1077_U134 , P2_R1077_U368 , P2_R1077_U302 );
and AND2_16965 ( P2_R1077_U135 , P2_R1077_U160 , P2_R1077_U278 );
and AND3_16966 ( P2_R1077_U136 , P2_R1077_U455 , P2_R1077_U454 , P2_R1077_U80 );
and AND2_16967 ( P2_R1077_U137 , P2_R1077_U325 , P2_R1077_U9 );
and AND3_16968 ( P2_R1077_U138 , P2_R1077_U469 , P2_R1077_U468 , P2_R1077_U59 );
and AND2_16969 ( P2_R1077_U139 , P2_R1077_U334 , P2_R1077_U8 );
and AND3_16970 ( P2_R1077_U140 , P2_R1077_U490 , P2_R1077_U489 , P2_R1077_U172 );
and AND2_16971 ( P2_R1077_U141 , P2_R1077_U343 , P2_R1077_U7 );
and AND3_16972 ( P2_R1077_U142 , P2_R1077_U502 , P2_R1077_U501 , P2_R1077_U171 );
and AND2_16973 ( P2_R1077_U143 , P2_R1077_U350 , P2_R1077_U6 );
nand NAND2_16974 ( P2_R1077_U144 , P2_R1077_U118 , P2_R1077_U202 );
nand NAND2_16975 ( P2_R1077_U145 , P2_R1077_U217 , P2_R1077_U229 );
not NOT1_16976 ( P2_R1077_U146 , P2_U3054 );
not NOT1_16977 ( P2_R1077_U147 , P2_U3904 );
and AND2_16978 ( P2_R1077_U148 , P2_R1077_U403 , P2_R1077_U402 );
nand NAND3_16979 ( P2_R1077_U149 , P2_R1077_U304 , P2_R1077_U169 , P2_R1077_U364 );
and AND2_16980 ( P2_R1077_U150 , P2_R1077_U410 , P2_R1077_U409 );
nand NAND3_16981 ( P2_R1077_U151 , P2_R1077_U370 , P2_R1077_U369 , P2_R1077_U134 );
and AND2_16982 ( P2_R1077_U152 , P2_R1077_U417 , P2_R1077_U416 );
nand NAND3_16983 ( P2_R1077_U153 , P2_R1077_U365 , P2_R1077_U299 , P2_R1077_U86 );
and AND2_16984 ( P2_R1077_U154 , P2_R1077_U424 , P2_R1077_U423 );
nand NAND2_16985 ( P2_R1077_U155 , P2_R1077_U293 , P2_R1077_U292 );
and AND2_16986 ( P2_R1077_U156 , P2_R1077_U436 , P2_R1077_U435 );
nand NAND2_16987 ( P2_R1077_U157 , P2_R1077_U289 , P2_R1077_U288 );
and AND2_16988 ( P2_R1077_U158 , P2_R1077_U443 , P2_R1077_U442 );
nand NAND2_16989 ( P2_R1077_U159 , P2_R1077_U132 , P2_R1077_U284 );
and AND2_16990 ( P2_R1077_U160 , P2_R1077_U450 , P2_R1077_U449 );
nand NAND2_16991 ( P2_R1077_U161 , P2_R1077_U43 , P2_R1077_U327 );
nand NAND2_16992 ( P2_R1077_U162 , P2_R1077_U130 , P2_R1077_U269 );
and AND2_16993 ( P2_R1077_U163 , P2_R1077_U476 , P2_R1077_U475 );
nand NAND2_16994 ( P2_R1077_U164 , P2_R1077_U257 , P2_R1077_U256 );
and AND2_16995 ( P2_R1077_U165 , P2_R1077_U483 , P2_R1077_U482 );
nand NAND2_16996 ( P2_R1077_U166 , P2_R1077_U129 , P2_R1077_U252 );
nand NAND2_16997 ( P2_R1077_U167 , P2_R1077_U127 , P2_R1077_U242 );
nand NAND2_16998 ( P2_R1077_U168 , P2_R1077_U367 , P2_R1077_U366 );
nand NAND2_16999 ( P2_R1077_U169 , P2_U3053 , P2_R1077_U151 );
not NOT1_17000 ( P2_R1077_U170 , P2_R1077_U34 );
nand NAND2_17001 ( P2_R1077_U171 , P2_U3416 , P2_U3082 );
nand NAND2_17002 ( P2_R1077_U172 , P2_U3071 , P2_U3425 );
nand NAND2_17003 ( P2_R1077_U173 , P2_U3057 , P2_U3898 );
not NOT1_17004 ( P2_R1077_U174 , P2_R1077_U68 );
not NOT1_17005 ( P2_R1077_U175 , P2_R1077_U77 );
nand NAND2_17006 ( P2_R1077_U176 , P2_U3064 , P2_U3899 );
not NOT1_17007 ( P2_R1077_U177 , P2_R1077_U65 );
or OR2_17008 ( P2_R1077_U178 , P2_U3066 , P2_U3404 );
or OR2_17009 ( P2_R1077_U179 , P2_U3059 , P2_U3401 );
or OR2_17010 ( P2_R1077_U180 , P2_U3398 , P2_U3063 );
or OR2_17011 ( P2_R1077_U181 , P2_U3395 , P2_U3067 );
not NOT1_17012 ( P2_R1077_U182 , P2_R1077_U31 );
or OR2_17013 ( P2_R1077_U183 , P2_U3392 , P2_U3077 );
not NOT1_17014 ( P2_R1077_U184 , P2_R1077_U42 );
not NOT1_17015 ( P2_R1077_U185 , P2_R1077_U43 );
nand NAND2_17016 ( P2_R1077_U186 , P2_R1077_U42 , P2_R1077_U43 );
nand NAND2_17017 ( P2_R1077_U187 , P2_U3067 , P2_U3395 );
nand NAND2_17018 ( P2_R1077_U188 , P2_R1077_U186 , P2_R1077_U181 );
nand NAND2_17019 ( P2_R1077_U189 , P2_U3063 , P2_U3398 );
nand NAND2_17020 ( P2_R1077_U190 , P2_R1077_U115 , P2_R1077_U188 );
nand NAND2_17021 ( P2_R1077_U191 , P2_R1077_U35 , P2_R1077_U34 );
nand NAND2_17022 ( P2_R1077_U192 , P2_U3066 , P2_R1077_U191 );
nand NAND2_17023 ( P2_R1077_U193 , P2_R1077_U116 , P2_R1077_U190 );
nand NAND2_17024 ( P2_R1077_U194 , P2_U3404 , P2_R1077_U170 );
not NOT1_17025 ( P2_R1077_U195 , P2_R1077_U41 );
or OR2_17026 ( P2_R1077_U196 , P2_U3069 , P2_U3410 );
or OR2_17027 ( P2_R1077_U197 , P2_U3070 , P2_U3407 );
not NOT1_17028 ( P2_R1077_U198 , P2_R1077_U22 );
nand NAND2_17029 ( P2_R1077_U199 , P2_R1077_U23 , P2_R1077_U22 );
nand NAND2_17030 ( P2_R1077_U200 , P2_U3069 , P2_R1077_U199 );
nand NAND2_17031 ( P2_R1077_U201 , P2_U3410 , P2_R1077_U198 );
nand NAND2_17032 ( P2_R1077_U202 , P2_R1077_U5 , P2_R1077_U41 );
not NOT1_17033 ( P2_R1077_U203 , P2_R1077_U144 );
or OR2_17034 ( P2_R1077_U204 , P2_U3413 , P2_U3083 );
nand NAND2_17035 ( P2_R1077_U205 , P2_R1077_U204 , P2_R1077_U144 );
not NOT1_17036 ( P2_R1077_U206 , P2_R1077_U40 );
or OR2_17037 ( P2_R1077_U207 , P2_U3082 , P2_U3416 );
or OR2_17038 ( P2_R1077_U208 , P2_U3407 , P2_U3070 );
nand NAND2_17039 ( P2_R1077_U209 , P2_R1077_U208 , P2_R1077_U41 );
nand NAND2_17040 ( P2_R1077_U210 , P2_R1077_U119 , P2_R1077_U209 );
nand NAND2_17041 ( P2_R1077_U211 , P2_R1077_U195 , P2_R1077_U22 );
nand NAND2_17042 ( P2_R1077_U212 , P2_U3410 , P2_U3069 );
nand NAND2_17043 ( P2_R1077_U213 , P2_R1077_U120 , P2_R1077_U211 );
or OR2_17044 ( P2_R1077_U214 , P2_U3070 , P2_U3407 );
nand NAND2_17045 ( P2_R1077_U215 , P2_R1077_U185 , P2_R1077_U181 );
nand NAND2_17046 ( P2_R1077_U216 , P2_U3067 , P2_U3395 );
not NOT1_17047 ( P2_R1077_U217 , P2_R1077_U45 );
nand NAND2_17048 ( P2_R1077_U218 , P2_R1077_U121 , P2_R1077_U184 );
nand NAND2_17049 ( P2_R1077_U219 , P2_R1077_U45 , P2_R1077_U180 );
nand NAND2_17050 ( P2_R1077_U220 , P2_U3063 , P2_U3398 );
not NOT1_17051 ( P2_R1077_U221 , P2_R1077_U44 );
or OR2_17052 ( P2_R1077_U222 , P2_U3401 , P2_U3059 );
nand NAND2_17053 ( P2_R1077_U223 , P2_R1077_U222 , P2_R1077_U44 );
nand NAND2_17054 ( P2_R1077_U224 , P2_R1077_U123 , P2_R1077_U223 );
nand NAND2_17055 ( P2_R1077_U225 , P2_R1077_U221 , P2_R1077_U34 );
nand NAND2_17056 ( P2_R1077_U226 , P2_U3404 , P2_U3066 );
nand NAND2_17057 ( P2_R1077_U227 , P2_R1077_U124 , P2_R1077_U225 );
or OR2_17058 ( P2_R1077_U228 , P2_U3059 , P2_U3401 );
nand NAND2_17059 ( P2_R1077_U229 , P2_R1077_U184 , P2_R1077_U181 );
not NOT1_17060 ( P2_R1077_U230 , P2_R1077_U145 );
nand NAND2_17061 ( P2_R1077_U231 , P2_U3063 , P2_U3398 );
nand NAND4_17062 ( P2_R1077_U232 , P2_R1077_U401 , P2_R1077_U400 , P2_R1077_U43 , P2_R1077_U42 );
nand NAND2_17063 ( P2_R1077_U233 , P2_R1077_U43 , P2_R1077_U42 );
nand NAND2_17064 ( P2_R1077_U234 , P2_U3067 , P2_U3395 );
nand NAND2_17065 ( P2_R1077_U235 , P2_R1077_U125 , P2_R1077_U233 );
or OR2_17066 ( P2_R1077_U236 , P2_U3082 , P2_U3416 );
or OR2_17067 ( P2_R1077_U237 , P2_U3061 , P2_U3419 );
nand NAND2_17068 ( P2_R1077_U238 , P2_R1077_U177 , P2_R1077_U6 );
nand NAND2_17069 ( P2_R1077_U239 , P2_U3061 , P2_U3419 );
nand NAND2_17070 ( P2_R1077_U240 , P2_R1077_U171 , P2_R1077_U238 );
or OR2_17071 ( P2_R1077_U241 , P2_U3419 , P2_U3061 );
nand NAND2_17072 ( P2_R1077_U242 , P2_R1077_U126 , P2_R1077_U144 );
nand NAND2_17073 ( P2_R1077_U243 , P2_R1077_U241 , P2_R1077_U240 );
not NOT1_17074 ( P2_R1077_U244 , P2_R1077_U167 );
or OR2_17075 ( P2_R1077_U245 , P2_U3079 , P2_U3428 );
or OR2_17076 ( P2_R1077_U246 , P2_U3071 , P2_U3425 );
nand NAND2_17077 ( P2_R1077_U247 , P2_R1077_U174 , P2_R1077_U7 );
nand NAND2_17078 ( P2_R1077_U248 , P2_U3079 , P2_U3428 );
nand NAND2_17079 ( P2_R1077_U249 , P2_R1077_U172 , P2_R1077_U247 );
or OR2_17080 ( P2_R1077_U250 , P2_U3422 , P2_U3062 );
or OR2_17081 ( P2_R1077_U251 , P2_U3428 , P2_U3079 );
nand NAND2_17082 ( P2_R1077_U252 , P2_R1077_U128 , P2_R1077_U167 );
nand NAND2_17083 ( P2_R1077_U253 , P2_R1077_U251 , P2_R1077_U249 );
not NOT1_17084 ( P2_R1077_U254 , P2_R1077_U166 );
or OR2_17085 ( P2_R1077_U255 , P2_U3431 , P2_U3078 );
nand NAND2_17086 ( P2_R1077_U256 , P2_R1077_U255 , P2_R1077_U166 );
nand NAND2_17087 ( P2_R1077_U257 , P2_U3078 , P2_U3431 );
not NOT1_17088 ( P2_R1077_U258 , P2_R1077_U164 );
or OR2_17089 ( P2_R1077_U259 , P2_U3434 , P2_U3073 );
nand NAND2_17090 ( P2_R1077_U260 , P2_R1077_U259 , P2_R1077_U164 );
nand NAND2_17091 ( P2_R1077_U261 , P2_U3073 , P2_U3434 );
not NOT1_17092 ( P2_R1077_U262 , P2_R1077_U92 );
or OR2_17093 ( P2_R1077_U263 , P2_U3068 , P2_U3440 );
or OR2_17094 ( P2_R1077_U264 , P2_U3072 , P2_U3437 );
not NOT1_17095 ( P2_R1077_U265 , P2_R1077_U59 );
nand NAND2_17096 ( P2_R1077_U266 , P2_R1077_U60 , P2_R1077_U59 );
nand NAND2_17097 ( P2_R1077_U267 , P2_U3068 , P2_R1077_U266 );
nand NAND2_17098 ( P2_R1077_U268 , P2_U3440 , P2_R1077_U265 );
nand NAND2_17099 ( P2_R1077_U269 , P2_R1077_U8 , P2_R1077_U92 );
not NOT1_17100 ( P2_R1077_U270 , P2_R1077_U162 );
or OR2_17101 ( P2_R1077_U271 , P2_U3075 , P2_U3903 );
or OR2_17102 ( P2_R1077_U272 , P2_U3080 , P2_U3445 );
or OR2_17103 ( P2_R1077_U273 , P2_U3074 , P2_U3902 );
not NOT1_17104 ( P2_R1077_U274 , P2_R1077_U80 );
nand NAND2_17105 ( P2_R1077_U275 , P2_U3903 , P2_R1077_U274 );
nand NAND2_17106 ( P2_R1077_U276 , P2_R1077_U275 , P2_R1077_U90 );
nand NAND2_17107 ( P2_R1077_U277 , P2_R1077_U80 , P2_R1077_U81 );
nand NAND2_17108 ( P2_R1077_U278 , P2_R1077_U277 , P2_R1077_U276 );
nand NAND2_17109 ( P2_R1077_U279 , P2_R1077_U175 , P2_R1077_U9 );
nand NAND2_17110 ( P2_R1077_U280 , P2_U3074 , P2_U3902 );
nand NAND2_17111 ( P2_R1077_U281 , P2_R1077_U278 , P2_R1077_U279 );
or OR2_17112 ( P2_R1077_U282 , P2_U3443 , P2_U3081 );
or OR2_17113 ( P2_R1077_U283 , P2_U3902 , P2_U3074 );
nand NAND3_17114 ( P2_R1077_U284 , P2_R1077_U273 , P2_R1077_U162 , P2_R1077_U131 );
nand NAND2_17115 ( P2_R1077_U285 , P2_R1077_U283 , P2_R1077_U281 );
not NOT1_17116 ( P2_R1077_U286 , P2_R1077_U159 );
or OR2_17117 ( P2_R1077_U287 , P2_U3901 , P2_U3060 );
nand NAND2_17118 ( P2_R1077_U288 , P2_R1077_U287 , P2_R1077_U159 );
nand NAND2_17119 ( P2_R1077_U289 , P2_U3060 , P2_U3901 );
not NOT1_17120 ( P2_R1077_U290 , P2_R1077_U157 );
or OR2_17121 ( P2_R1077_U291 , P2_U3900 , P2_U3065 );
nand NAND2_17122 ( P2_R1077_U292 , P2_R1077_U291 , P2_R1077_U157 );
nand NAND2_17123 ( P2_R1077_U293 , P2_U3065 , P2_U3900 );
not NOT1_17124 ( P2_R1077_U294 , P2_R1077_U155 );
or OR2_17125 ( P2_R1077_U295 , P2_U3057 , P2_U3898 );
nand NAND2_17126 ( P2_R1077_U296 , P2_R1077_U176 , P2_R1077_U173 );
not NOT1_17127 ( P2_R1077_U297 , P2_R1077_U86 );
or OR2_17128 ( P2_R1077_U298 , P2_U3899 , P2_U3064 );
nand NAND3_17129 ( P2_R1077_U299 , P2_R1077_U155 , P2_R1077_U298 , P2_R1077_U168 );
not NOT1_17130 ( P2_R1077_U300 , P2_R1077_U153 );
or OR2_17131 ( P2_R1077_U301 , P2_U3896 , P2_U3052 );
nand NAND2_17132 ( P2_R1077_U302 , P2_U3052 , P2_U3896 );
not NOT1_17133 ( P2_R1077_U303 , P2_R1077_U151 );
nand NAND2_17134 ( P2_R1077_U304 , P2_U3895 , P2_R1077_U151 );
not NOT1_17135 ( P2_R1077_U305 , P2_R1077_U149 );
nand NAND2_17136 ( P2_R1077_U306 , P2_R1077_U298 , P2_R1077_U155 );
not NOT1_17137 ( P2_R1077_U307 , P2_R1077_U89 );
or OR2_17138 ( P2_R1077_U308 , P2_U3898 , P2_U3057 );
nand NAND2_17139 ( P2_R1077_U309 , P2_R1077_U308 , P2_R1077_U89 );
nand NAND3_17140 ( P2_R1077_U310 , P2_R1077_U309 , P2_R1077_U173 , P2_R1077_U154 );
nand NAND2_17141 ( P2_R1077_U311 , P2_R1077_U307 , P2_R1077_U173 );
nand NAND2_17142 ( P2_R1077_U312 , P2_U3897 , P2_U3056 );
nand NAND3_17143 ( P2_R1077_U313 , P2_R1077_U311 , P2_R1077_U312 , P2_R1077_U168 );
or OR2_17144 ( P2_R1077_U314 , P2_U3057 , P2_U3898 );
nand NAND2_17145 ( P2_R1077_U315 , P2_R1077_U282 , P2_R1077_U162 );
not NOT1_17146 ( P2_R1077_U316 , P2_R1077_U91 );
nand NAND2_17147 ( P2_R1077_U317 , P2_R1077_U9 , P2_R1077_U91 );
nand NAND2_17148 ( P2_R1077_U318 , P2_R1077_U135 , P2_R1077_U317 );
nand NAND2_17149 ( P2_R1077_U319 , P2_R1077_U317 , P2_R1077_U278 );
nand NAND2_17150 ( P2_R1077_U320 , P2_R1077_U453 , P2_R1077_U319 );
or OR2_17151 ( P2_R1077_U321 , P2_U3445 , P2_U3080 );
nand NAND2_17152 ( P2_R1077_U322 , P2_R1077_U321 , P2_R1077_U91 );
nand NAND2_17153 ( P2_R1077_U323 , P2_R1077_U136 , P2_R1077_U322 );
nand NAND2_17154 ( P2_R1077_U324 , P2_R1077_U316 , P2_R1077_U80 );
nand NAND2_17155 ( P2_R1077_U325 , P2_U3075 , P2_U3903 );
nand NAND2_17156 ( P2_R1077_U326 , P2_R1077_U137 , P2_R1077_U324 );
or OR2_17157 ( P2_R1077_U327 , P2_U3392 , P2_U3077 );
not NOT1_17158 ( P2_R1077_U328 , P2_R1077_U161 );
or OR2_17159 ( P2_R1077_U329 , P2_U3080 , P2_U3445 );
or OR2_17160 ( P2_R1077_U330 , P2_U3437 , P2_U3072 );
nand NAND2_17161 ( P2_R1077_U331 , P2_R1077_U330 , P2_R1077_U92 );
nand NAND2_17162 ( P2_R1077_U332 , P2_R1077_U138 , P2_R1077_U331 );
nand NAND2_17163 ( P2_R1077_U333 , P2_R1077_U262 , P2_R1077_U59 );
nand NAND2_17164 ( P2_R1077_U334 , P2_U3440 , P2_U3068 );
nand NAND2_17165 ( P2_R1077_U335 , P2_R1077_U139 , P2_R1077_U333 );
or OR2_17166 ( P2_R1077_U336 , P2_U3072 , P2_U3437 );
nand NAND2_17167 ( P2_R1077_U337 , P2_R1077_U250 , P2_R1077_U167 );
not NOT1_17168 ( P2_R1077_U338 , P2_R1077_U93 );
or OR2_17169 ( P2_R1077_U339 , P2_U3425 , P2_U3071 );
nand NAND2_17170 ( P2_R1077_U340 , P2_R1077_U339 , P2_R1077_U93 );
nand NAND2_17171 ( P2_R1077_U341 , P2_R1077_U140 , P2_R1077_U340 );
nand NAND2_17172 ( P2_R1077_U342 , P2_R1077_U338 , P2_R1077_U172 );
nand NAND2_17173 ( P2_R1077_U343 , P2_U3079 , P2_U3428 );
nand NAND2_17174 ( P2_R1077_U344 , P2_R1077_U141 , P2_R1077_U342 );
or OR2_17175 ( P2_R1077_U345 , P2_U3071 , P2_U3425 );
or OR2_17176 ( P2_R1077_U346 , P2_U3416 , P2_U3082 );
nand NAND2_17177 ( P2_R1077_U347 , P2_R1077_U346 , P2_R1077_U40 );
nand NAND2_17178 ( P2_R1077_U348 , P2_R1077_U142 , P2_R1077_U347 );
nand NAND2_17179 ( P2_R1077_U349 , P2_R1077_U206 , P2_R1077_U171 );
nand NAND2_17180 ( P2_R1077_U350 , P2_U3061 , P2_U3419 );
nand NAND2_17181 ( P2_R1077_U351 , P2_R1077_U143 , P2_R1077_U349 );
nand NAND2_17182 ( P2_R1077_U352 , P2_R1077_U207 , P2_R1077_U171 );
nand NAND2_17183 ( P2_R1077_U353 , P2_R1077_U204 , P2_R1077_U65 );
nand NAND2_17184 ( P2_R1077_U354 , P2_R1077_U214 , P2_R1077_U22 );
nand NAND2_17185 ( P2_R1077_U355 , P2_R1077_U228 , P2_R1077_U34 );
nand NAND2_17186 ( P2_R1077_U356 , P2_R1077_U231 , P2_R1077_U180 );
nand NAND2_17187 ( P2_R1077_U357 , P2_R1077_U314 , P2_R1077_U173 );
nand NAND2_17188 ( P2_R1077_U358 , P2_R1077_U298 , P2_R1077_U176 );
nand NAND2_17189 ( P2_R1077_U359 , P2_R1077_U329 , P2_R1077_U80 );
nand NAND2_17190 ( P2_R1077_U360 , P2_R1077_U282 , P2_R1077_U77 );
nand NAND2_17191 ( P2_R1077_U361 , P2_R1077_U336 , P2_R1077_U59 );
nand NAND2_17192 ( P2_R1077_U362 , P2_R1077_U345 , P2_R1077_U172 );
nand NAND2_17193 ( P2_R1077_U363 , P2_R1077_U250 , P2_R1077_U68 );
nand NAND2_17194 ( P2_R1077_U364 , P2_U3895 , P2_U3053 );
nand NAND2_17195 ( P2_R1077_U365 , P2_R1077_U296 , P2_R1077_U168 );
nand NAND2_17196 ( P2_R1077_U366 , P2_U3056 , P2_R1077_U295 );
nand NAND2_17197 ( P2_R1077_U367 , P2_U3897 , P2_R1077_U295 );
nand NAND3_17198 ( P2_R1077_U368 , P2_R1077_U296 , P2_R1077_U168 , P2_R1077_U301 );
nand NAND3_17199 ( P2_R1077_U369 , P2_R1077_U155 , P2_R1077_U168 , P2_R1077_U133 );
nand NAND2_17200 ( P2_R1077_U370 , P2_R1077_U297 , P2_R1077_U301 );
nand NAND2_17201 ( P2_R1077_U371 , P2_U3082 , P2_R1077_U39 );
nand NAND2_17202 ( P2_R1077_U372 , P2_U3416 , P2_R1077_U38 );
nand NAND2_17203 ( P2_R1077_U373 , P2_R1077_U372 , P2_R1077_U371 );
nand NAND2_17204 ( P2_R1077_U374 , P2_R1077_U352 , P2_R1077_U40 );
nand NAND2_17205 ( P2_R1077_U375 , P2_R1077_U373 , P2_R1077_U206 );
nand NAND2_17206 ( P2_R1077_U376 , P2_U3083 , P2_R1077_U36 );
nand NAND2_17207 ( P2_R1077_U377 , P2_U3413 , P2_R1077_U37 );
nand NAND2_17208 ( P2_R1077_U378 , P2_R1077_U377 , P2_R1077_U376 );
nand NAND2_17209 ( P2_R1077_U379 , P2_R1077_U353 , P2_R1077_U144 );
nand NAND2_17210 ( P2_R1077_U380 , P2_R1077_U203 , P2_R1077_U378 );
nand NAND2_17211 ( P2_R1077_U381 , P2_U3069 , P2_R1077_U23 );
nand NAND2_17212 ( P2_R1077_U382 , P2_U3410 , P2_R1077_U21 );
nand NAND2_17213 ( P2_R1077_U383 , P2_U3070 , P2_R1077_U19 );
nand NAND2_17214 ( P2_R1077_U384 , P2_U3407 , P2_R1077_U20 );
nand NAND2_17215 ( P2_R1077_U385 , P2_R1077_U384 , P2_R1077_U383 );
nand NAND2_17216 ( P2_R1077_U386 , P2_R1077_U354 , P2_R1077_U41 );
nand NAND2_17217 ( P2_R1077_U387 , P2_R1077_U385 , P2_R1077_U195 );
nand NAND2_17218 ( P2_R1077_U388 , P2_U3066 , P2_R1077_U35 );
nand NAND2_17219 ( P2_R1077_U389 , P2_U3404 , P2_R1077_U26 );
nand NAND2_17220 ( P2_R1077_U390 , P2_U3059 , P2_R1077_U24 );
nand NAND2_17221 ( P2_R1077_U391 , P2_U3401 , P2_R1077_U25 );
nand NAND2_17222 ( P2_R1077_U392 , P2_R1077_U391 , P2_R1077_U390 );
nand NAND2_17223 ( P2_R1077_U393 , P2_R1077_U355 , P2_R1077_U44 );
nand NAND2_17224 ( P2_R1077_U394 , P2_R1077_U392 , P2_R1077_U221 );
nand NAND2_17225 ( P2_R1077_U395 , P2_U3063 , P2_R1077_U32 );
nand NAND2_17226 ( P2_R1077_U396 , P2_U3398 , P2_R1077_U33 );
nand NAND2_17227 ( P2_R1077_U397 , P2_R1077_U396 , P2_R1077_U395 );
nand NAND2_17228 ( P2_R1077_U398 , P2_R1077_U356 , P2_R1077_U145 );
nand NAND2_17229 ( P2_R1077_U399 , P2_R1077_U230 , P2_R1077_U397 );
nand NAND2_17230 ( P2_R1077_U400 , P2_U3067 , P2_R1077_U27 );
nand NAND2_17231 ( P2_R1077_U401 , P2_U3395 , P2_R1077_U28 );
nand NAND2_17232 ( P2_R1077_U402 , P2_U3054 , P2_R1077_U147 );
nand NAND2_17233 ( P2_R1077_U403 , P2_U3904 , P2_R1077_U146 );
nand NAND2_17234 ( P2_R1077_U404 , P2_U3054 , P2_R1077_U147 );
nand NAND2_17235 ( P2_R1077_U405 , P2_U3904 , P2_R1077_U146 );
nand NAND2_17236 ( P2_R1077_U406 , P2_R1077_U405 , P2_R1077_U404 );
nand NAND2_17237 ( P2_R1077_U407 , P2_R1077_U148 , P2_R1077_U149 );
nand NAND2_17238 ( P2_R1077_U408 , P2_R1077_U305 , P2_R1077_U406 );
nand NAND2_17239 ( P2_R1077_U409 , P2_U3053 , P2_R1077_U88 );
nand NAND2_17240 ( P2_R1077_U410 , P2_U3895 , P2_R1077_U87 );
nand NAND2_17241 ( P2_R1077_U411 , P2_U3053 , P2_R1077_U88 );
nand NAND2_17242 ( P2_R1077_U412 , P2_U3895 , P2_R1077_U87 );
nand NAND2_17243 ( P2_R1077_U413 , P2_R1077_U412 , P2_R1077_U411 );
nand NAND2_17244 ( P2_R1077_U414 , P2_R1077_U150 , P2_R1077_U151 );
nand NAND2_17245 ( P2_R1077_U415 , P2_R1077_U303 , P2_R1077_U413 );
nand NAND2_17246 ( P2_R1077_U416 , P2_U3052 , P2_R1077_U46 );
nand NAND2_17247 ( P2_R1077_U417 , P2_U3896 , P2_R1077_U47 );
nand NAND2_17248 ( P2_R1077_U418 , P2_U3052 , P2_R1077_U46 );
nand NAND2_17249 ( P2_R1077_U419 , P2_U3896 , P2_R1077_U47 );
nand NAND2_17250 ( P2_R1077_U420 , P2_R1077_U419 , P2_R1077_U418 );
nand NAND2_17251 ( P2_R1077_U421 , P2_R1077_U152 , P2_R1077_U153 );
nand NAND2_17252 ( P2_R1077_U422 , P2_R1077_U300 , P2_R1077_U420 );
nand NAND2_17253 ( P2_R1077_U423 , P2_U3056 , P2_R1077_U49 );
nand NAND2_17254 ( P2_R1077_U424 , P2_U3897 , P2_R1077_U48 );
nand NAND2_17255 ( P2_R1077_U425 , P2_U3057 , P2_R1077_U50 );
nand NAND2_17256 ( P2_R1077_U426 , P2_U3898 , P2_R1077_U51 );
nand NAND2_17257 ( P2_R1077_U427 , P2_R1077_U426 , P2_R1077_U425 );
nand NAND2_17258 ( P2_R1077_U428 , P2_R1077_U357 , P2_R1077_U89 );
nand NAND2_17259 ( P2_R1077_U429 , P2_R1077_U427 , P2_R1077_U307 );
nand NAND2_17260 ( P2_R1077_U430 , P2_U3064 , P2_R1077_U52 );
nand NAND2_17261 ( P2_R1077_U431 , P2_U3899 , P2_R1077_U53 );
nand NAND2_17262 ( P2_R1077_U432 , P2_R1077_U431 , P2_R1077_U430 );
nand NAND2_17263 ( P2_R1077_U433 , P2_R1077_U358 , P2_R1077_U155 );
nand NAND2_17264 ( P2_R1077_U434 , P2_R1077_U294 , P2_R1077_U432 );
nand NAND2_17265 ( P2_R1077_U435 , P2_U3065 , P2_R1077_U84 );
nand NAND2_17266 ( P2_R1077_U436 , P2_U3900 , P2_R1077_U85 );
nand NAND2_17267 ( P2_R1077_U437 , P2_U3065 , P2_R1077_U84 );
nand NAND2_17268 ( P2_R1077_U438 , P2_U3900 , P2_R1077_U85 );
nand NAND2_17269 ( P2_R1077_U439 , P2_R1077_U438 , P2_R1077_U437 );
nand NAND2_17270 ( P2_R1077_U440 , P2_R1077_U156 , P2_R1077_U157 );
nand NAND2_17271 ( P2_R1077_U441 , P2_R1077_U290 , P2_R1077_U439 );
nand NAND2_17272 ( P2_R1077_U442 , P2_U3060 , P2_R1077_U82 );
nand NAND2_17273 ( P2_R1077_U443 , P2_U3901 , P2_R1077_U83 );
nand NAND2_17274 ( P2_R1077_U444 , P2_U3060 , P2_R1077_U82 );
nand NAND2_17275 ( P2_R1077_U445 , P2_U3901 , P2_R1077_U83 );
nand NAND2_17276 ( P2_R1077_U446 , P2_R1077_U445 , P2_R1077_U444 );
nand NAND2_17277 ( P2_R1077_U447 , P2_R1077_U158 , P2_R1077_U159 );
nand NAND2_17278 ( P2_R1077_U448 , P2_R1077_U286 , P2_R1077_U446 );
nand NAND2_17279 ( P2_R1077_U449 , P2_U3074 , P2_R1077_U54 );
nand NAND2_17280 ( P2_R1077_U450 , P2_U3902 , P2_R1077_U55 );
nand NAND2_17281 ( P2_R1077_U451 , P2_U3074 , P2_R1077_U54 );
nand NAND2_17282 ( P2_R1077_U452 , P2_U3902 , P2_R1077_U55 );
nand NAND2_17283 ( P2_R1077_U453 , P2_R1077_U452 , P2_R1077_U451 );
nand NAND2_17284 ( P2_R1077_U454 , P2_U3075 , P2_R1077_U81 );
nand NAND2_17285 ( P2_R1077_U455 , P2_U3903 , P2_R1077_U90 );
nand NAND2_17286 ( P2_R1077_U456 , P2_R1077_U182 , P2_R1077_U161 );
nand NAND2_17287 ( P2_R1077_U457 , P2_R1077_U328 , P2_R1077_U31 );
nand NAND2_17288 ( P2_R1077_U458 , P2_U3080 , P2_R1077_U78 );
nand NAND2_17289 ( P2_R1077_U459 , P2_U3445 , P2_R1077_U79 );
nand NAND2_17290 ( P2_R1077_U460 , P2_R1077_U459 , P2_R1077_U458 );
nand NAND2_17291 ( P2_R1077_U461 , P2_R1077_U359 , P2_R1077_U91 );
nand NAND2_17292 ( P2_R1077_U462 , P2_R1077_U460 , P2_R1077_U316 );
nand NAND2_17293 ( P2_R1077_U463 , P2_U3081 , P2_R1077_U75 );
nand NAND2_17294 ( P2_R1077_U464 , P2_U3443 , P2_R1077_U76 );
nand NAND2_17295 ( P2_R1077_U465 , P2_R1077_U464 , P2_R1077_U463 );
nand NAND2_17296 ( P2_R1077_U466 , P2_R1077_U360 , P2_R1077_U162 );
nand NAND2_17297 ( P2_R1077_U467 , P2_R1077_U270 , P2_R1077_U465 );
nand NAND2_17298 ( P2_R1077_U468 , P2_U3068 , P2_R1077_U60 );
nand NAND2_17299 ( P2_R1077_U469 , P2_U3440 , P2_R1077_U58 );
nand NAND2_17300 ( P2_R1077_U470 , P2_U3072 , P2_R1077_U56 );
nand NAND2_17301 ( P2_R1077_U471 , P2_U3437 , P2_R1077_U57 );
nand NAND2_17302 ( P2_R1077_U472 , P2_R1077_U471 , P2_R1077_U470 );
nand NAND2_17303 ( P2_R1077_U473 , P2_R1077_U361 , P2_R1077_U92 );
nand NAND2_17304 ( P2_R1077_U474 , P2_R1077_U472 , P2_R1077_U262 );
nand NAND2_17305 ( P2_R1077_U475 , P2_U3073 , P2_R1077_U73 );
nand NAND2_17306 ( P2_R1077_U476 , P2_U3434 , P2_R1077_U74 );
nand NAND2_17307 ( P2_R1077_U477 , P2_U3073 , P2_R1077_U73 );
nand NAND2_17308 ( P2_R1077_U478 , P2_U3434 , P2_R1077_U74 );
nand NAND2_17309 ( P2_R1077_U479 , P2_R1077_U478 , P2_R1077_U477 );
nand NAND2_17310 ( P2_R1077_U480 , P2_R1077_U163 , P2_R1077_U164 );
nand NAND2_17311 ( P2_R1077_U481 , P2_R1077_U258 , P2_R1077_U479 );
nand NAND2_17312 ( P2_R1077_U482 , P2_U3078 , P2_R1077_U71 );
nand NAND2_17313 ( P2_R1077_U483 , P2_U3431 , P2_R1077_U72 );
nand NAND2_17314 ( P2_R1077_U484 , P2_U3078 , P2_R1077_U71 );
nand NAND2_17315 ( P2_R1077_U485 , P2_U3431 , P2_R1077_U72 );
nand NAND2_17316 ( P2_R1077_U486 , P2_R1077_U485 , P2_R1077_U484 );
nand NAND2_17317 ( P2_R1077_U487 , P2_R1077_U165 , P2_R1077_U166 );
nand NAND2_17318 ( P2_R1077_U488 , P2_R1077_U254 , P2_R1077_U486 );
nand NAND2_17319 ( P2_R1077_U489 , P2_U3079 , P2_R1077_U61 );
nand NAND2_17320 ( P2_R1077_U490 , P2_U3428 , P2_R1077_U62 );
nand NAND2_17321 ( P2_R1077_U491 , P2_U3071 , P2_R1077_U69 );
nand NAND2_17322 ( P2_R1077_U492 , P2_U3425 , P2_R1077_U70 );
nand NAND2_17323 ( P2_R1077_U493 , P2_R1077_U492 , P2_R1077_U491 );
nand NAND2_17324 ( P2_R1077_U494 , P2_R1077_U362 , P2_R1077_U93 );
nand NAND2_17325 ( P2_R1077_U495 , P2_R1077_U493 , P2_R1077_U338 );
nand NAND2_17326 ( P2_R1077_U496 , P2_U3062 , P2_R1077_U66 );
nand NAND2_17327 ( P2_R1077_U497 , P2_U3422 , P2_R1077_U67 );
nand NAND2_17328 ( P2_R1077_U498 , P2_R1077_U497 , P2_R1077_U496 );
nand NAND2_17329 ( P2_R1077_U499 , P2_R1077_U363 , P2_R1077_U167 );
nand NAND2_17330 ( P2_R1077_U500 , P2_R1077_U244 , P2_R1077_U498 );
nand NAND2_17331 ( P2_R1077_U501 , P2_U3061 , P2_R1077_U63 );
nand NAND2_17332 ( P2_R1077_U502 , P2_U3419 , P2_R1077_U64 );
nand NAND2_17333 ( P2_R1077_U503 , P2_U3076 , P2_R1077_U29 );
nand NAND2_17334 ( P2_R1077_U504 , P2_U3387 , P2_R1077_U30 );
and AND2_17335 ( P2_R1143_U4 , P2_R1143_U179 , P2_R1143_U178 );
and AND2_17336 ( P2_R1143_U5 , P2_R1143_U197 , P2_R1143_U196 );
and AND2_17337 ( P2_R1143_U6 , P2_R1143_U237 , P2_R1143_U236 );
and AND2_17338 ( P2_R1143_U7 , P2_R1143_U246 , P2_R1143_U245 );
and AND2_17339 ( P2_R1143_U8 , P2_R1143_U264 , P2_R1143_U263 );
and AND2_17340 ( P2_R1143_U9 , P2_R1143_U272 , P2_R1143_U271 );
and AND2_17341 ( P2_R1143_U10 , P2_R1143_U351 , P2_R1143_U348 );
and AND2_17342 ( P2_R1143_U11 , P2_R1143_U344 , P2_R1143_U341 );
and AND2_17343 ( P2_R1143_U12 , P2_R1143_U335 , P2_R1143_U332 );
and AND2_17344 ( P2_R1143_U13 , P2_R1143_U326 , P2_R1143_U323 );
and AND2_17345 ( P2_R1143_U14 , P2_R1143_U320 , P2_R1143_U318 );
and AND2_17346 ( P2_R1143_U15 , P2_R1143_U313 , P2_R1143_U310 );
and AND2_17347 ( P2_R1143_U16 , P2_R1143_U235 , P2_R1143_U232 );
and AND2_17348 ( P2_R1143_U17 , P2_R1143_U227 , P2_R1143_U224 );
and AND2_17349 ( P2_R1143_U18 , P2_R1143_U213 , P2_R1143_U210 );
not NOT1_17350 ( P2_R1143_U19 , P2_U3407 );
not NOT1_17351 ( P2_R1143_U20 , P2_U3070 );
not NOT1_17352 ( P2_R1143_U21 , P2_U3069 );
nand NAND2_17353 ( P2_R1143_U22 , P2_U3070 , P2_U3407 );
not NOT1_17354 ( P2_R1143_U23 , P2_U3410 );
not NOT1_17355 ( P2_R1143_U24 , P2_U3401 );
not NOT1_17356 ( P2_R1143_U25 , P2_U3059 );
not NOT1_17357 ( P2_R1143_U26 , P2_U3066 );
not NOT1_17358 ( P2_R1143_U27 , P2_U3395 );
not NOT1_17359 ( P2_R1143_U28 , P2_U3067 );
not NOT1_17360 ( P2_R1143_U29 , P2_U3387 );
not NOT1_17361 ( P2_R1143_U30 , P2_U3076 );
nand NAND2_17362 ( P2_R1143_U31 , P2_U3076 , P2_U3387 );
not NOT1_17363 ( P2_R1143_U32 , P2_U3398 );
not NOT1_17364 ( P2_R1143_U33 , P2_U3063 );
nand NAND2_17365 ( P2_R1143_U34 , P2_U3059 , P2_U3401 );
not NOT1_17366 ( P2_R1143_U35 , P2_U3404 );
not NOT1_17367 ( P2_R1143_U36 , P2_U3413 );
not NOT1_17368 ( P2_R1143_U37 , P2_U3083 );
not NOT1_17369 ( P2_R1143_U38 , P2_U3082 );
not NOT1_17370 ( P2_R1143_U39 , P2_U3416 );
nand NAND2_17371 ( P2_R1143_U40 , P2_R1143_U65 , P2_R1143_U205 );
nand NAND2_17372 ( P2_R1143_U41 , P2_R1143_U117 , P2_R1143_U193 );
nand NAND2_17373 ( P2_R1143_U42 , P2_R1143_U182 , P2_R1143_U183 );
nand NAND2_17374 ( P2_R1143_U43 , P2_U3392 , P2_U3077 );
nand NAND2_17375 ( P2_R1143_U44 , P2_R1143_U122 , P2_R1143_U219 );
nand NAND2_17376 ( P2_R1143_U45 , P2_R1143_U216 , P2_R1143_U215 );
not NOT1_17377 ( P2_R1143_U46 , P2_U3896 );
not NOT1_17378 ( P2_R1143_U47 , P2_U3052 );
not NOT1_17379 ( P2_R1143_U48 , P2_U3056 );
not NOT1_17380 ( P2_R1143_U49 , P2_U3897 );
not NOT1_17381 ( P2_R1143_U50 , P2_U3898 );
not NOT1_17382 ( P2_R1143_U51 , P2_U3057 );
not NOT1_17383 ( P2_R1143_U52 , P2_U3899 );
not NOT1_17384 ( P2_R1143_U53 , P2_U3064 );
not NOT1_17385 ( P2_R1143_U54 , P2_U3902 );
not NOT1_17386 ( P2_R1143_U55 , P2_U3074 );
not NOT1_17387 ( P2_R1143_U56 , P2_U3437 );
not NOT1_17388 ( P2_R1143_U57 , P2_U3072 );
not NOT1_17389 ( P2_R1143_U58 , P2_U3068 );
nand NAND2_17390 ( P2_R1143_U59 , P2_U3072 , P2_U3437 );
not NOT1_17391 ( P2_R1143_U60 , P2_U3440 );
not NOT1_17392 ( P2_R1143_U61 , P2_U3428 );
not NOT1_17393 ( P2_R1143_U62 , P2_U3079 );
not NOT1_17394 ( P2_R1143_U63 , P2_U3419 );
not NOT1_17395 ( P2_R1143_U64 , P2_U3061 );
nand NAND2_17396 ( P2_R1143_U65 , P2_U3083 , P2_U3413 );
not NOT1_17397 ( P2_R1143_U66 , P2_U3422 );
not NOT1_17398 ( P2_R1143_U67 , P2_U3062 );
nand NAND2_17399 ( P2_R1143_U68 , P2_U3062 , P2_U3422 );
not NOT1_17400 ( P2_R1143_U69 , P2_U3425 );
not NOT1_17401 ( P2_R1143_U70 , P2_U3071 );
not NOT1_17402 ( P2_R1143_U71 , P2_U3431 );
not NOT1_17403 ( P2_R1143_U72 , P2_U3078 );
not NOT1_17404 ( P2_R1143_U73 , P2_U3434 );
not NOT1_17405 ( P2_R1143_U74 , P2_U3073 );
not NOT1_17406 ( P2_R1143_U75 , P2_U3443 );
not NOT1_17407 ( P2_R1143_U76 , P2_U3081 );
nand NAND2_17408 ( P2_R1143_U77 , P2_U3081 , P2_U3443 );
not NOT1_17409 ( P2_R1143_U78 , P2_U3445 );
not NOT1_17410 ( P2_R1143_U79 , P2_U3080 );
nand NAND2_17411 ( P2_R1143_U80 , P2_U3080 , P2_U3445 );
not NOT1_17412 ( P2_R1143_U81 , P2_U3903 );
not NOT1_17413 ( P2_R1143_U82 , P2_U3901 );
not NOT1_17414 ( P2_R1143_U83 , P2_U3060 );
not NOT1_17415 ( P2_R1143_U84 , P2_U3900 );
not NOT1_17416 ( P2_R1143_U85 , P2_U3065 );
nand NAND2_17417 ( P2_R1143_U86 , P2_U3897 , P2_U3056 );
not NOT1_17418 ( P2_R1143_U87 , P2_U3053 );
not NOT1_17419 ( P2_R1143_U88 , P2_U3895 );
nand NAND2_17420 ( P2_R1143_U89 , P2_R1143_U306 , P2_R1143_U176 );
not NOT1_17421 ( P2_R1143_U90 , P2_U3075 );
nand NAND2_17422 ( P2_R1143_U91 , P2_R1143_U77 , P2_R1143_U315 );
nand NAND2_17423 ( P2_R1143_U92 , P2_R1143_U261 , P2_R1143_U260 );
nand NAND2_17424 ( P2_R1143_U93 , P2_R1143_U68 , P2_R1143_U337 );
nand NAND2_17425 ( P2_R1143_U94 , P2_R1143_U457 , P2_R1143_U456 );
nand NAND2_17426 ( P2_R1143_U95 , P2_R1143_U504 , P2_R1143_U503 );
nand NAND2_17427 ( P2_R1143_U96 , P2_R1143_U375 , P2_R1143_U374 );
nand NAND2_17428 ( P2_R1143_U97 , P2_R1143_U380 , P2_R1143_U379 );
nand NAND2_17429 ( P2_R1143_U98 , P2_R1143_U387 , P2_R1143_U386 );
nand NAND2_17430 ( P2_R1143_U99 , P2_R1143_U394 , P2_R1143_U393 );
nand NAND2_17431 ( P2_R1143_U100 , P2_R1143_U399 , P2_R1143_U398 );
nand NAND2_17432 ( P2_R1143_U101 , P2_R1143_U408 , P2_R1143_U407 );
nand NAND2_17433 ( P2_R1143_U102 , P2_R1143_U415 , P2_R1143_U414 );
nand NAND2_17434 ( P2_R1143_U103 , P2_R1143_U422 , P2_R1143_U421 );
nand NAND2_17435 ( P2_R1143_U104 , P2_R1143_U429 , P2_R1143_U428 );
nand NAND2_17436 ( P2_R1143_U105 , P2_R1143_U434 , P2_R1143_U433 );
nand NAND2_17437 ( P2_R1143_U106 , P2_R1143_U441 , P2_R1143_U440 );
nand NAND2_17438 ( P2_R1143_U107 , P2_R1143_U448 , P2_R1143_U447 );
nand NAND2_17439 ( P2_R1143_U108 , P2_R1143_U462 , P2_R1143_U461 );
nand NAND2_17440 ( P2_R1143_U109 , P2_R1143_U467 , P2_R1143_U466 );
nand NAND2_17441 ( P2_R1143_U110 , P2_R1143_U474 , P2_R1143_U473 );
nand NAND2_17442 ( P2_R1143_U111 , P2_R1143_U481 , P2_R1143_U480 );
nand NAND2_17443 ( P2_R1143_U112 , P2_R1143_U488 , P2_R1143_U487 );
nand NAND2_17444 ( P2_R1143_U113 , P2_R1143_U495 , P2_R1143_U494 );
nand NAND2_17445 ( P2_R1143_U114 , P2_R1143_U500 , P2_R1143_U499 );
and AND2_17446 ( P2_R1143_U115 , P2_R1143_U189 , P2_R1143_U187 );
and AND2_17447 ( P2_R1143_U116 , P2_R1143_U4 , P2_R1143_U180 );
and AND2_17448 ( P2_R1143_U117 , P2_R1143_U194 , P2_R1143_U192 );
and AND2_17449 ( P2_R1143_U118 , P2_R1143_U201 , P2_R1143_U200 );
and AND3_17450 ( P2_R1143_U119 , P2_R1143_U382 , P2_R1143_U381 , P2_R1143_U22 );
and AND2_17451 ( P2_R1143_U120 , P2_R1143_U212 , P2_R1143_U5 );
and AND2_17452 ( P2_R1143_U121 , P2_R1143_U181 , P2_R1143_U180 );
and AND2_17453 ( P2_R1143_U122 , P2_R1143_U220 , P2_R1143_U218 );
and AND3_17454 ( P2_R1143_U123 , P2_R1143_U389 , P2_R1143_U388 , P2_R1143_U34 );
and AND2_17455 ( P2_R1143_U124 , P2_R1143_U226 , P2_R1143_U4 );
and AND2_17456 ( P2_R1143_U125 , P2_R1143_U234 , P2_R1143_U181 );
and AND2_17457 ( P2_R1143_U126 , P2_R1143_U204 , P2_R1143_U6 );
and AND2_17458 ( P2_R1143_U127 , P2_R1143_U243 , P2_R1143_U239 );
and AND2_17459 ( P2_R1143_U128 , P2_R1143_U250 , P2_R1143_U7 );
and AND2_17460 ( P2_R1143_U129 , P2_R1143_U253 , P2_R1143_U248 );
and AND2_17461 ( P2_R1143_U130 , P2_R1143_U268 , P2_R1143_U267 );
and AND2_17462 ( P2_R1143_U131 , P2_R1143_U9 , P2_R1143_U282 );
and AND2_17463 ( P2_R1143_U132 , P2_R1143_U285 , P2_R1143_U280 );
and AND2_17464 ( P2_R1143_U133 , P2_R1143_U301 , P2_R1143_U298 );
and AND2_17465 ( P2_R1143_U134 , P2_R1143_U368 , P2_R1143_U302 );
and AND2_17466 ( P2_R1143_U135 , P2_R1143_U160 , P2_R1143_U278 );
and AND3_17467 ( P2_R1143_U136 , P2_R1143_U455 , P2_R1143_U454 , P2_R1143_U80 );
and AND2_17468 ( P2_R1143_U137 , P2_R1143_U325 , P2_R1143_U9 );
and AND3_17469 ( P2_R1143_U138 , P2_R1143_U469 , P2_R1143_U468 , P2_R1143_U59 );
and AND2_17470 ( P2_R1143_U139 , P2_R1143_U334 , P2_R1143_U8 );
and AND3_17471 ( P2_R1143_U140 , P2_R1143_U490 , P2_R1143_U489 , P2_R1143_U172 );
and AND2_17472 ( P2_R1143_U141 , P2_R1143_U343 , P2_R1143_U7 );
and AND3_17473 ( P2_R1143_U142 , P2_R1143_U502 , P2_R1143_U501 , P2_R1143_U171 );
and AND2_17474 ( P2_R1143_U143 , P2_R1143_U350 , P2_R1143_U6 );
nand NAND2_17475 ( P2_R1143_U144 , P2_R1143_U118 , P2_R1143_U202 );
nand NAND2_17476 ( P2_R1143_U145 , P2_R1143_U217 , P2_R1143_U229 );
not NOT1_17477 ( P2_R1143_U146 , P2_U3054 );
not NOT1_17478 ( P2_R1143_U147 , P2_U3904 );
and AND2_17479 ( P2_R1143_U148 , P2_R1143_U403 , P2_R1143_U402 );
nand NAND3_17480 ( P2_R1143_U149 , P2_R1143_U304 , P2_R1143_U169 , P2_R1143_U364 );
and AND2_17481 ( P2_R1143_U150 , P2_R1143_U410 , P2_R1143_U409 );
nand NAND3_17482 ( P2_R1143_U151 , P2_R1143_U370 , P2_R1143_U369 , P2_R1143_U134 );
and AND2_17483 ( P2_R1143_U152 , P2_R1143_U417 , P2_R1143_U416 );
nand NAND3_17484 ( P2_R1143_U153 , P2_R1143_U365 , P2_R1143_U299 , P2_R1143_U86 );
and AND2_17485 ( P2_R1143_U154 , P2_R1143_U424 , P2_R1143_U423 );
nand NAND2_17486 ( P2_R1143_U155 , P2_R1143_U293 , P2_R1143_U292 );
and AND2_17487 ( P2_R1143_U156 , P2_R1143_U436 , P2_R1143_U435 );
nand NAND2_17488 ( P2_R1143_U157 , P2_R1143_U289 , P2_R1143_U288 );
and AND2_17489 ( P2_R1143_U158 , P2_R1143_U443 , P2_R1143_U442 );
nand NAND2_17490 ( P2_R1143_U159 , P2_R1143_U132 , P2_R1143_U284 );
and AND2_17491 ( P2_R1143_U160 , P2_R1143_U450 , P2_R1143_U449 );
nand NAND2_17492 ( P2_R1143_U161 , P2_R1143_U43 , P2_R1143_U327 );
nand NAND2_17493 ( P2_R1143_U162 , P2_R1143_U130 , P2_R1143_U269 );
and AND2_17494 ( P2_R1143_U163 , P2_R1143_U476 , P2_R1143_U475 );
nand NAND2_17495 ( P2_R1143_U164 , P2_R1143_U257 , P2_R1143_U256 );
and AND2_17496 ( P2_R1143_U165 , P2_R1143_U483 , P2_R1143_U482 );
nand NAND2_17497 ( P2_R1143_U166 , P2_R1143_U129 , P2_R1143_U252 );
nand NAND2_17498 ( P2_R1143_U167 , P2_R1143_U127 , P2_R1143_U242 );
nand NAND2_17499 ( P2_R1143_U168 , P2_R1143_U367 , P2_R1143_U366 );
nand NAND2_17500 ( P2_R1143_U169 , P2_U3053 , P2_R1143_U151 );
not NOT1_17501 ( P2_R1143_U170 , P2_R1143_U34 );
nand NAND2_17502 ( P2_R1143_U171 , P2_U3416 , P2_U3082 );
nand NAND2_17503 ( P2_R1143_U172 , P2_U3071 , P2_U3425 );
nand NAND2_17504 ( P2_R1143_U173 , P2_U3057 , P2_U3898 );
not NOT1_17505 ( P2_R1143_U174 , P2_R1143_U68 );
not NOT1_17506 ( P2_R1143_U175 , P2_R1143_U77 );
nand NAND2_17507 ( P2_R1143_U176 , P2_U3064 , P2_U3899 );
not NOT1_17508 ( P2_R1143_U177 , P2_R1143_U65 );
or OR2_17509 ( P2_R1143_U178 , P2_U3066 , P2_U3404 );
or OR2_17510 ( P2_R1143_U179 , P2_U3059 , P2_U3401 );
or OR2_17511 ( P2_R1143_U180 , P2_U3398 , P2_U3063 );
or OR2_17512 ( P2_R1143_U181 , P2_U3395 , P2_U3067 );
not NOT1_17513 ( P2_R1143_U182 , P2_R1143_U31 );
or OR2_17514 ( P2_R1143_U183 , P2_U3392 , P2_U3077 );
not NOT1_17515 ( P2_R1143_U184 , P2_R1143_U42 );
not NOT1_17516 ( P2_R1143_U185 , P2_R1143_U43 );
nand NAND2_17517 ( P2_R1143_U186 , P2_R1143_U42 , P2_R1143_U43 );
nand NAND2_17518 ( P2_R1143_U187 , P2_U3067 , P2_U3395 );
nand NAND2_17519 ( P2_R1143_U188 , P2_R1143_U186 , P2_R1143_U181 );
nand NAND2_17520 ( P2_R1143_U189 , P2_U3063 , P2_U3398 );
nand NAND2_17521 ( P2_R1143_U190 , P2_R1143_U115 , P2_R1143_U188 );
nand NAND2_17522 ( P2_R1143_U191 , P2_R1143_U35 , P2_R1143_U34 );
nand NAND2_17523 ( P2_R1143_U192 , P2_U3066 , P2_R1143_U191 );
nand NAND2_17524 ( P2_R1143_U193 , P2_R1143_U116 , P2_R1143_U190 );
nand NAND2_17525 ( P2_R1143_U194 , P2_U3404 , P2_R1143_U170 );
not NOT1_17526 ( P2_R1143_U195 , P2_R1143_U41 );
or OR2_17527 ( P2_R1143_U196 , P2_U3069 , P2_U3410 );
or OR2_17528 ( P2_R1143_U197 , P2_U3070 , P2_U3407 );
not NOT1_17529 ( P2_R1143_U198 , P2_R1143_U22 );
nand NAND2_17530 ( P2_R1143_U199 , P2_R1143_U23 , P2_R1143_U22 );
nand NAND2_17531 ( P2_R1143_U200 , P2_U3069 , P2_R1143_U199 );
nand NAND2_17532 ( P2_R1143_U201 , P2_U3410 , P2_R1143_U198 );
nand NAND2_17533 ( P2_R1143_U202 , P2_R1143_U5 , P2_R1143_U41 );
not NOT1_17534 ( P2_R1143_U203 , P2_R1143_U144 );
or OR2_17535 ( P2_R1143_U204 , P2_U3413 , P2_U3083 );
nand NAND2_17536 ( P2_R1143_U205 , P2_R1143_U204 , P2_R1143_U144 );
not NOT1_17537 ( P2_R1143_U206 , P2_R1143_U40 );
or OR2_17538 ( P2_R1143_U207 , P2_U3082 , P2_U3416 );
or OR2_17539 ( P2_R1143_U208 , P2_U3407 , P2_U3070 );
nand NAND2_17540 ( P2_R1143_U209 , P2_R1143_U208 , P2_R1143_U41 );
nand NAND2_17541 ( P2_R1143_U210 , P2_R1143_U119 , P2_R1143_U209 );
nand NAND2_17542 ( P2_R1143_U211 , P2_R1143_U195 , P2_R1143_U22 );
nand NAND2_17543 ( P2_R1143_U212 , P2_U3410 , P2_U3069 );
nand NAND2_17544 ( P2_R1143_U213 , P2_R1143_U120 , P2_R1143_U211 );
or OR2_17545 ( P2_R1143_U214 , P2_U3070 , P2_U3407 );
nand NAND2_17546 ( P2_R1143_U215 , P2_R1143_U185 , P2_R1143_U181 );
nand NAND2_17547 ( P2_R1143_U216 , P2_U3067 , P2_U3395 );
not NOT1_17548 ( P2_R1143_U217 , P2_R1143_U45 );
nand NAND2_17549 ( P2_R1143_U218 , P2_R1143_U121 , P2_R1143_U184 );
nand NAND2_17550 ( P2_R1143_U219 , P2_R1143_U45 , P2_R1143_U180 );
nand NAND2_17551 ( P2_R1143_U220 , P2_U3063 , P2_U3398 );
not NOT1_17552 ( P2_R1143_U221 , P2_R1143_U44 );
or OR2_17553 ( P2_R1143_U222 , P2_U3401 , P2_U3059 );
nand NAND2_17554 ( P2_R1143_U223 , P2_R1143_U222 , P2_R1143_U44 );
nand NAND2_17555 ( P2_R1143_U224 , P2_R1143_U123 , P2_R1143_U223 );
nand NAND2_17556 ( P2_R1143_U225 , P2_R1143_U221 , P2_R1143_U34 );
nand NAND2_17557 ( P2_R1143_U226 , P2_U3404 , P2_U3066 );
nand NAND2_17558 ( P2_R1143_U227 , P2_R1143_U124 , P2_R1143_U225 );
or OR2_17559 ( P2_R1143_U228 , P2_U3059 , P2_U3401 );
nand NAND2_17560 ( P2_R1143_U229 , P2_R1143_U184 , P2_R1143_U181 );
not NOT1_17561 ( P2_R1143_U230 , P2_R1143_U145 );
nand NAND2_17562 ( P2_R1143_U231 , P2_U3063 , P2_U3398 );
nand NAND4_17563 ( P2_R1143_U232 , P2_R1143_U401 , P2_R1143_U400 , P2_R1143_U43 , P2_R1143_U42 );
nand NAND2_17564 ( P2_R1143_U233 , P2_R1143_U43 , P2_R1143_U42 );
nand NAND2_17565 ( P2_R1143_U234 , P2_U3067 , P2_U3395 );
nand NAND2_17566 ( P2_R1143_U235 , P2_R1143_U125 , P2_R1143_U233 );
or OR2_17567 ( P2_R1143_U236 , P2_U3082 , P2_U3416 );
or OR2_17568 ( P2_R1143_U237 , P2_U3061 , P2_U3419 );
nand NAND2_17569 ( P2_R1143_U238 , P2_R1143_U177 , P2_R1143_U6 );
nand NAND2_17570 ( P2_R1143_U239 , P2_U3061 , P2_U3419 );
nand NAND2_17571 ( P2_R1143_U240 , P2_R1143_U171 , P2_R1143_U238 );
or OR2_17572 ( P2_R1143_U241 , P2_U3419 , P2_U3061 );
nand NAND2_17573 ( P2_R1143_U242 , P2_R1143_U126 , P2_R1143_U144 );
nand NAND2_17574 ( P2_R1143_U243 , P2_R1143_U241 , P2_R1143_U240 );
not NOT1_17575 ( P2_R1143_U244 , P2_R1143_U167 );
or OR2_17576 ( P2_R1143_U245 , P2_U3079 , P2_U3428 );
or OR2_17577 ( P2_R1143_U246 , P2_U3071 , P2_U3425 );
nand NAND2_17578 ( P2_R1143_U247 , P2_R1143_U174 , P2_R1143_U7 );
nand NAND2_17579 ( P2_R1143_U248 , P2_U3079 , P2_U3428 );
nand NAND2_17580 ( P2_R1143_U249 , P2_R1143_U172 , P2_R1143_U247 );
or OR2_17581 ( P2_R1143_U250 , P2_U3422 , P2_U3062 );
or OR2_17582 ( P2_R1143_U251 , P2_U3428 , P2_U3079 );
nand NAND2_17583 ( P2_R1143_U252 , P2_R1143_U128 , P2_R1143_U167 );
nand NAND2_17584 ( P2_R1143_U253 , P2_R1143_U251 , P2_R1143_U249 );
not NOT1_17585 ( P2_R1143_U254 , P2_R1143_U166 );
or OR2_17586 ( P2_R1143_U255 , P2_U3431 , P2_U3078 );
nand NAND2_17587 ( P2_R1143_U256 , P2_R1143_U255 , P2_R1143_U166 );
nand NAND2_17588 ( P2_R1143_U257 , P2_U3078 , P2_U3431 );
not NOT1_17589 ( P2_R1143_U258 , P2_R1143_U164 );
or OR2_17590 ( P2_R1143_U259 , P2_U3434 , P2_U3073 );
nand NAND2_17591 ( P2_R1143_U260 , P2_R1143_U259 , P2_R1143_U164 );
nand NAND2_17592 ( P2_R1143_U261 , P2_U3073 , P2_U3434 );
not NOT1_17593 ( P2_R1143_U262 , P2_R1143_U92 );
or OR2_17594 ( P2_R1143_U263 , P2_U3068 , P2_U3440 );
or OR2_17595 ( P2_R1143_U264 , P2_U3072 , P2_U3437 );
not NOT1_17596 ( P2_R1143_U265 , P2_R1143_U59 );
nand NAND2_17597 ( P2_R1143_U266 , P2_R1143_U60 , P2_R1143_U59 );
nand NAND2_17598 ( P2_R1143_U267 , P2_U3068 , P2_R1143_U266 );
nand NAND2_17599 ( P2_R1143_U268 , P2_U3440 , P2_R1143_U265 );
nand NAND2_17600 ( P2_R1143_U269 , P2_R1143_U8 , P2_R1143_U92 );
not NOT1_17601 ( P2_R1143_U270 , P2_R1143_U162 );
or OR2_17602 ( P2_R1143_U271 , P2_U3075 , P2_U3903 );
or OR2_17603 ( P2_R1143_U272 , P2_U3080 , P2_U3445 );
or OR2_17604 ( P2_R1143_U273 , P2_U3074 , P2_U3902 );
not NOT1_17605 ( P2_R1143_U274 , P2_R1143_U80 );
nand NAND2_17606 ( P2_R1143_U275 , P2_U3903 , P2_R1143_U274 );
nand NAND2_17607 ( P2_R1143_U276 , P2_R1143_U275 , P2_R1143_U90 );
nand NAND2_17608 ( P2_R1143_U277 , P2_R1143_U80 , P2_R1143_U81 );
nand NAND2_17609 ( P2_R1143_U278 , P2_R1143_U277 , P2_R1143_U276 );
nand NAND2_17610 ( P2_R1143_U279 , P2_R1143_U175 , P2_R1143_U9 );
nand NAND2_17611 ( P2_R1143_U280 , P2_U3074 , P2_U3902 );
nand NAND2_17612 ( P2_R1143_U281 , P2_R1143_U278 , P2_R1143_U279 );
or OR2_17613 ( P2_R1143_U282 , P2_U3443 , P2_U3081 );
or OR2_17614 ( P2_R1143_U283 , P2_U3902 , P2_U3074 );
nand NAND3_17615 ( P2_R1143_U284 , P2_R1143_U273 , P2_R1143_U162 , P2_R1143_U131 );
nand NAND2_17616 ( P2_R1143_U285 , P2_R1143_U283 , P2_R1143_U281 );
not NOT1_17617 ( P2_R1143_U286 , P2_R1143_U159 );
or OR2_17618 ( P2_R1143_U287 , P2_U3901 , P2_U3060 );
nand NAND2_17619 ( P2_R1143_U288 , P2_R1143_U287 , P2_R1143_U159 );
nand NAND2_17620 ( P2_R1143_U289 , P2_U3060 , P2_U3901 );
not NOT1_17621 ( P2_R1143_U290 , P2_R1143_U157 );
or OR2_17622 ( P2_R1143_U291 , P2_U3900 , P2_U3065 );
nand NAND2_17623 ( P2_R1143_U292 , P2_R1143_U291 , P2_R1143_U157 );
nand NAND2_17624 ( P2_R1143_U293 , P2_U3065 , P2_U3900 );
not NOT1_17625 ( P2_R1143_U294 , P2_R1143_U155 );
or OR2_17626 ( P2_R1143_U295 , P2_U3057 , P2_U3898 );
nand NAND2_17627 ( P2_R1143_U296 , P2_R1143_U176 , P2_R1143_U173 );
not NOT1_17628 ( P2_R1143_U297 , P2_R1143_U86 );
or OR2_17629 ( P2_R1143_U298 , P2_U3899 , P2_U3064 );
nand NAND3_17630 ( P2_R1143_U299 , P2_R1143_U155 , P2_R1143_U298 , P2_R1143_U168 );
not NOT1_17631 ( P2_R1143_U300 , P2_R1143_U153 );
or OR2_17632 ( P2_R1143_U301 , P2_U3896 , P2_U3052 );
nand NAND2_17633 ( P2_R1143_U302 , P2_U3052 , P2_U3896 );
not NOT1_17634 ( P2_R1143_U303 , P2_R1143_U151 );
nand NAND2_17635 ( P2_R1143_U304 , P2_U3895 , P2_R1143_U151 );
not NOT1_17636 ( P2_R1143_U305 , P2_R1143_U149 );
nand NAND2_17637 ( P2_R1143_U306 , P2_R1143_U298 , P2_R1143_U155 );
not NOT1_17638 ( P2_R1143_U307 , P2_R1143_U89 );
or OR2_17639 ( P2_R1143_U308 , P2_U3898 , P2_U3057 );
nand NAND2_17640 ( P2_R1143_U309 , P2_R1143_U308 , P2_R1143_U89 );
nand NAND3_17641 ( P2_R1143_U310 , P2_R1143_U309 , P2_R1143_U173 , P2_R1143_U154 );
nand NAND2_17642 ( P2_R1143_U311 , P2_R1143_U307 , P2_R1143_U173 );
nand NAND2_17643 ( P2_R1143_U312 , P2_U3897 , P2_U3056 );
nand NAND3_17644 ( P2_R1143_U313 , P2_R1143_U311 , P2_R1143_U312 , P2_R1143_U168 );
or OR2_17645 ( P2_R1143_U314 , P2_U3057 , P2_U3898 );
nand NAND2_17646 ( P2_R1143_U315 , P2_R1143_U282 , P2_R1143_U162 );
not NOT1_17647 ( P2_R1143_U316 , P2_R1143_U91 );
nand NAND2_17648 ( P2_R1143_U317 , P2_R1143_U9 , P2_R1143_U91 );
nand NAND2_17649 ( P2_R1143_U318 , P2_R1143_U135 , P2_R1143_U317 );
nand NAND2_17650 ( P2_R1143_U319 , P2_R1143_U317 , P2_R1143_U278 );
nand NAND2_17651 ( P2_R1143_U320 , P2_R1143_U453 , P2_R1143_U319 );
or OR2_17652 ( P2_R1143_U321 , P2_U3445 , P2_U3080 );
nand NAND2_17653 ( P2_R1143_U322 , P2_R1143_U321 , P2_R1143_U91 );
nand NAND2_17654 ( P2_R1143_U323 , P2_R1143_U136 , P2_R1143_U322 );
nand NAND2_17655 ( P2_R1143_U324 , P2_R1143_U316 , P2_R1143_U80 );
nand NAND2_17656 ( P2_R1143_U325 , P2_U3075 , P2_U3903 );
nand NAND2_17657 ( P2_R1143_U326 , P2_R1143_U137 , P2_R1143_U324 );
or OR2_17658 ( P2_R1143_U327 , P2_U3392 , P2_U3077 );
not NOT1_17659 ( P2_R1143_U328 , P2_R1143_U161 );
or OR2_17660 ( P2_R1143_U329 , P2_U3080 , P2_U3445 );
or OR2_17661 ( P2_R1143_U330 , P2_U3437 , P2_U3072 );
nand NAND2_17662 ( P2_R1143_U331 , P2_R1143_U330 , P2_R1143_U92 );
nand NAND2_17663 ( P2_R1143_U332 , P2_R1143_U138 , P2_R1143_U331 );
nand NAND2_17664 ( P2_R1143_U333 , P2_R1143_U262 , P2_R1143_U59 );
nand NAND2_17665 ( P2_R1143_U334 , P2_U3440 , P2_U3068 );
nand NAND2_17666 ( P2_R1143_U335 , P2_R1143_U139 , P2_R1143_U333 );
or OR2_17667 ( P2_R1143_U336 , P2_U3072 , P2_U3437 );
nand NAND2_17668 ( P2_R1143_U337 , P2_R1143_U250 , P2_R1143_U167 );
not NOT1_17669 ( P2_R1143_U338 , P2_R1143_U93 );
or OR2_17670 ( P2_R1143_U339 , P2_U3425 , P2_U3071 );
nand NAND2_17671 ( P2_R1143_U340 , P2_R1143_U339 , P2_R1143_U93 );
nand NAND2_17672 ( P2_R1143_U341 , P2_R1143_U140 , P2_R1143_U340 );
nand NAND2_17673 ( P2_R1143_U342 , P2_R1143_U338 , P2_R1143_U172 );
nand NAND2_17674 ( P2_R1143_U343 , P2_U3079 , P2_U3428 );
nand NAND2_17675 ( P2_R1143_U344 , P2_R1143_U141 , P2_R1143_U342 );
or OR2_17676 ( P2_R1143_U345 , P2_U3071 , P2_U3425 );
or OR2_17677 ( P2_R1143_U346 , P2_U3416 , P2_U3082 );
nand NAND2_17678 ( P2_R1143_U347 , P2_R1143_U346 , P2_R1143_U40 );
nand NAND2_17679 ( P2_R1143_U348 , P2_R1143_U142 , P2_R1143_U347 );
nand NAND2_17680 ( P2_R1143_U349 , P2_R1143_U206 , P2_R1143_U171 );
nand NAND2_17681 ( P2_R1143_U350 , P2_U3061 , P2_U3419 );
nand NAND2_17682 ( P2_R1143_U351 , P2_R1143_U143 , P2_R1143_U349 );
nand NAND2_17683 ( P2_R1143_U352 , P2_R1143_U207 , P2_R1143_U171 );
nand NAND2_17684 ( P2_R1143_U353 , P2_R1143_U204 , P2_R1143_U65 );
nand NAND2_17685 ( P2_R1143_U354 , P2_R1143_U214 , P2_R1143_U22 );
nand NAND2_17686 ( P2_R1143_U355 , P2_R1143_U228 , P2_R1143_U34 );
nand NAND2_17687 ( P2_R1143_U356 , P2_R1143_U231 , P2_R1143_U180 );
nand NAND2_17688 ( P2_R1143_U357 , P2_R1143_U314 , P2_R1143_U173 );
nand NAND2_17689 ( P2_R1143_U358 , P2_R1143_U298 , P2_R1143_U176 );
nand NAND2_17690 ( P2_R1143_U359 , P2_R1143_U329 , P2_R1143_U80 );
nand NAND2_17691 ( P2_R1143_U360 , P2_R1143_U282 , P2_R1143_U77 );
nand NAND2_17692 ( P2_R1143_U361 , P2_R1143_U336 , P2_R1143_U59 );
nand NAND2_17693 ( P2_R1143_U362 , P2_R1143_U345 , P2_R1143_U172 );
nand NAND2_17694 ( P2_R1143_U363 , P2_R1143_U250 , P2_R1143_U68 );
nand NAND2_17695 ( P2_R1143_U364 , P2_U3895 , P2_U3053 );
nand NAND2_17696 ( P2_R1143_U365 , P2_R1143_U296 , P2_R1143_U168 );
nand NAND2_17697 ( P2_R1143_U366 , P2_U3056 , P2_R1143_U295 );
nand NAND2_17698 ( P2_R1143_U367 , P2_U3897 , P2_R1143_U295 );
nand NAND3_17699 ( P2_R1143_U368 , P2_R1143_U296 , P2_R1143_U168 , P2_R1143_U301 );
nand NAND3_17700 ( P2_R1143_U369 , P2_R1143_U155 , P2_R1143_U168 , P2_R1143_U133 );
nand NAND2_17701 ( P2_R1143_U370 , P2_R1143_U297 , P2_R1143_U301 );
nand NAND2_17702 ( P2_R1143_U371 , P2_U3082 , P2_R1143_U39 );
nand NAND2_17703 ( P2_R1143_U372 , P2_U3416 , P2_R1143_U38 );
nand NAND2_17704 ( P2_R1143_U373 , P2_R1143_U372 , P2_R1143_U371 );
nand NAND2_17705 ( P2_R1143_U374 , P2_R1143_U352 , P2_R1143_U40 );
nand NAND2_17706 ( P2_R1143_U375 , P2_R1143_U373 , P2_R1143_U206 );
nand NAND2_17707 ( P2_R1143_U376 , P2_U3083 , P2_R1143_U36 );
nand NAND2_17708 ( P2_R1143_U377 , P2_U3413 , P2_R1143_U37 );
nand NAND2_17709 ( P2_R1143_U378 , P2_R1143_U377 , P2_R1143_U376 );
nand NAND2_17710 ( P2_R1143_U379 , P2_R1143_U353 , P2_R1143_U144 );
nand NAND2_17711 ( P2_R1143_U380 , P2_R1143_U203 , P2_R1143_U378 );
nand NAND2_17712 ( P2_R1143_U381 , P2_U3069 , P2_R1143_U23 );
nand NAND2_17713 ( P2_R1143_U382 , P2_U3410 , P2_R1143_U21 );
nand NAND2_17714 ( P2_R1143_U383 , P2_U3070 , P2_R1143_U19 );
nand NAND2_17715 ( P2_R1143_U384 , P2_U3407 , P2_R1143_U20 );
nand NAND2_17716 ( P2_R1143_U385 , P2_R1143_U384 , P2_R1143_U383 );
nand NAND2_17717 ( P2_R1143_U386 , P2_R1143_U354 , P2_R1143_U41 );
nand NAND2_17718 ( P2_R1143_U387 , P2_R1143_U385 , P2_R1143_U195 );
nand NAND2_17719 ( P2_R1143_U388 , P2_U3066 , P2_R1143_U35 );
nand NAND2_17720 ( P2_R1143_U389 , P2_U3404 , P2_R1143_U26 );
nand NAND2_17721 ( P2_R1143_U390 , P2_U3059 , P2_R1143_U24 );
nand NAND2_17722 ( P2_R1143_U391 , P2_U3401 , P2_R1143_U25 );
nand NAND2_17723 ( P2_R1143_U392 , P2_R1143_U391 , P2_R1143_U390 );
nand NAND2_17724 ( P2_R1143_U393 , P2_R1143_U355 , P2_R1143_U44 );
nand NAND2_17725 ( P2_R1143_U394 , P2_R1143_U392 , P2_R1143_U221 );
nand NAND2_17726 ( P2_R1143_U395 , P2_U3063 , P2_R1143_U32 );
nand NAND2_17727 ( P2_R1143_U396 , P2_U3398 , P2_R1143_U33 );
nand NAND2_17728 ( P2_R1143_U397 , P2_R1143_U396 , P2_R1143_U395 );
nand NAND2_17729 ( P2_R1143_U398 , P2_R1143_U356 , P2_R1143_U145 );
nand NAND2_17730 ( P2_R1143_U399 , P2_R1143_U230 , P2_R1143_U397 );
nand NAND2_17731 ( P2_R1143_U400 , P2_U3067 , P2_R1143_U27 );
nand NAND2_17732 ( P2_R1143_U401 , P2_U3395 , P2_R1143_U28 );
nand NAND2_17733 ( P2_R1143_U402 , P2_U3054 , P2_R1143_U147 );
nand NAND2_17734 ( P2_R1143_U403 , P2_U3904 , P2_R1143_U146 );
nand NAND2_17735 ( P2_R1143_U404 , P2_U3054 , P2_R1143_U147 );
nand NAND2_17736 ( P2_R1143_U405 , P2_U3904 , P2_R1143_U146 );
nand NAND2_17737 ( P2_R1143_U406 , P2_R1143_U405 , P2_R1143_U404 );
nand NAND2_17738 ( P2_R1143_U407 , P2_R1143_U148 , P2_R1143_U149 );
nand NAND2_17739 ( P2_R1143_U408 , P2_R1143_U305 , P2_R1143_U406 );
nand NAND2_17740 ( P2_R1143_U409 , P2_U3053 , P2_R1143_U88 );
nand NAND2_17741 ( P2_R1143_U410 , P2_U3895 , P2_R1143_U87 );
nand NAND2_17742 ( P2_R1143_U411 , P2_U3053 , P2_R1143_U88 );
nand NAND2_17743 ( P2_R1143_U412 , P2_U3895 , P2_R1143_U87 );
nand NAND2_17744 ( P2_R1143_U413 , P2_R1143_U412 , P2_R1143_U411 );
nand NAND2_17745 ( P2_R1143_U414 , P2_R1143_U150 , P2_R1143_U151 );
nand NAND2_17746 ( P2_R1143_U415 , P2_R1143_U303 , P2_R1143_U413 );
nand NAND2_17747 ( P2_R1143_U416 , P2_U3052 , P2_R1143_U46 );
nand NAND2_17748 ( P2_R1143_U417 , P2_U3896 , P2_R1143_U47 );
nand NAND2_17749 ( P2_R1143_U418 , P2_U3052 , P2_R1143_U46 );
nand NAND2_17750 ( P2_R1143_U419 , P2_U3896 , P2_R1143_U47 );
nand NAND2_17751 ( P2_R1143_U420 , P2_R1143_U419 , P2_R1143_U418 );
nand NAND2_17752 ( P2_R1143_U421 , P2_R1143_U152 , P2_R1143_U153 );
nand NAND2_17753 ( P2_R1143_U422 , P2_R1143_U300 , P2_R1143_U420 );
nand NAND2_17754 ( P2_R1143_U423 , P2_U3056 , P2_R1143_U49 );
nand NAND2_17755 ( P2_R1143_U424 , P2_U3897 , P2_R1143_U48 );
nand NAND2_17756 ( P2_R1143_U425 , P2_U3057 , P2_R1143_U50 );
nand NAND2_17757 ( P2_R1143_U426 , P2_U3898 , P2_R1143_U51 );
nand NAND2_17758 ( P2_R1143_U427 , P2_R1143_U426 , P2_R1143_U425 );
nand NAND2_17759 ( P2_R1143_U428 , P2_R1143_U357 , P2_R1143_U89 );
nand NAND2_17760 ( P2_R1143_U429 , P2_R1143_U427 , P2_R1143_U307 );
nand NAND2_17761 ( P2_R1143_U430 , P2_U3064 , P2_R1143_U52 );
nand NAND2_17762 ( P2_R1143_U431 , P2_U3899 , P2_R1143_U53 );
nand NAND2_17763 ( P2_R1143_U432 , P2_R1143_U431 , P2_R1143_U430 );
nand NAND2_17764 ( P2_R1143_U433 , P2_R1143_U358 , P2_R1143_U155 );
nand NAND2_17765 ( P2_R1143_U434 , P2_R1143_U294 , P2_R1143_U432 );
nand NAND2_17766 ( P2_R1143_U435 , P2_U3065 , P2_R1143_U84 );
nand NAND2_17767 ( P2_R1143_U436 , P2_U3900 , P2_R1143_U85 );
nand NAND2_17768 ( P2_R1143_U437 , P2_U3065 , P2_R1143_U84 );
nand NAND2_17769 ( P2_R1143_U438 , P2_U3900 , P2_R1143_U85 );
nand NAND2_17770 ( P2_R1143_U439 , P2_R1143_U438 , P2_R1143_U437 );
nand NAND2_17771 ( P2_R1143_U440 , P2_R1143_U156 , P2_R1143_U157 );
nand NAND2_17772 ( P2_R1143_U441 , P2_R1143_U290 , P2_R1143_U439 );
nand NAND2_17773 ( P2_R1143_U442 , P2_U3060 , P2_R1143_U82 );
nand NAND2_17774 ( P2_R1143_U443 , P2_U3901 , P2_R1143_U83 );
nand NAND2_17775 ( P2_R1143_U444 , P2_U3060 , P2_R1143_U82 );
nand NAND2_17776 ( P2_R1143_U445 , P2_U3901 , P2_R1143_U83 );
nand NAND2_17777 ( P2_R1143_U446 , P2_R1143_U445 , P2_R1143_U444 );
nand NAND2_17778 ( P2_R1143_U447 , P2_R1143_U158 , P2_R1143_U159 );
nand NAND2_17779 ( P2_R1143_U448 , P2_R1143_U286 , P2_R1143_U446 );
nand NAND2_17780 ( P2_R1143_U449 , P2_U3074 , P2_R1143_U54 );
nand NAND2_17781 ( P2_R1143_U450 , P2_U3902 , P2_R1143_U55 );
nand NAND2_17782 ( P2_R1143_U451 , P2_U3074 , P2_R1143_U54 );
nand NAND2_17783 ( P2_R1143_U452 , P2_U3902 , P2_R1143_U55 );
nand NAND2_17784 ( P2_R1143_U453 , P2_R1143_U452 , P2_R1143_U451 );
nand NAND2_17785 ( P2_R1143_U454 , P2_U3075 , P2_R1143_U81 );
nand NAND2_17786 ( P2_R1143_U455 , P2_U3903 , P2_R1143_U90 );
nand NAND2_17787 ( P2_R1143_U456 , P2_R1143_U182 , P2_R1143_U161 );
nand NAND2_17788 ( P2_R1143_U457 , P2_R1143_U328 , P2_R1143_U31 );
nand NAND2_17789 ( P2_R1143_U458 , P2_U3080 , P2_R1143_U78 );
nand NAND2_17790 ( P2_R1143_U459 , P2_U3445 , P2_R1143_U79 );
nand NAND2_17791 ( P2_R1143_U460 , P2_R1143_U459 , P2_R1143_U458 );
nand NAND2_17792 ( P2_R1143_U461 , P2_R1143_U359 , P2_R1143_U91 );
nand NAND2_17793 ( P2_R1143_U462 , P2_R1143_U460 , P2_R1143_U316 );
nand NAND2_17794 ( P2_R1143_U463 , P2_U3081 , P2_R1143_U75 );
nand NAND2_17795 ( P2_R1143_U464 , P2_U3443 , P2_R1143_U76 );
nand NAND2_17796 ( P2_R1143_U465 , P2_R1143_U464 , P2_R1143_U463 );
nand NAND2_17797 ( P2_R1143_U466 , P2_R1143_U360 , P2_R1143_U162 );
nand NAND2_17798 ( P2_R1143_U467 , P2_R1143_U270 , P2_R1143_U465 );
nand NAND2_17799 ( P2_R1143_U468 , P2_U3068 , P2_R1143_U60 );
nand NAND2_17800 ( P2_R1143_U469 , P2_U3440 , P2_R1143_U58 );
nand NAND2_17801 ( P2_R1143_U470 , P2_U3072 , P2_R1143_U56 );
nand NAND2_17802 ( P2_R1143_U471 , P2_U3437 , P2_R1143_U57 );
nand NAND2_17803 ( P2_R1143_U472 , P2_R1143_U471 , P2_R1143_U470 );
nand NAND2_17804 ( P2_R1143_U473 , P2_R1143_U361 , P2_R1143_U92 );
nand NAND2_17805 ( P2_R1143_U474 , P2_R1143_U472 , P2_R1143_U262 );
nand NAND2_17806 ( P2_R1143_U475 , P2_U3073 , P2_R1143_U73 );
nand NAND2_17807 ( P2_R1143_U476 , P2_U3434 , P2_R1143_U74 );
nand NAND2_17808 ( P2_R1143_U477 , P2_U3073 , P2_R1143_U73 );
nand NAND2_17809 ( P2_R1143_U478 , P2_U3434 , P2_R1143_U74 );
nand NAND2_17810 ( P2_R1143_U479 , P2_R1143_U478 , P2_R1143_U477 );
nand NAND2_17811 ( P2_R1143_U480 , P2_R1143_U163 , P2_R1143_U164 );
nand NAND2_17812 ( P2_R1143_U481 , P2_R1143_U258 , P2_R1143_U479 );
nand NAND2_17813 ( P2_R1143_U482 , P2_U3078 , P2_R1143_U71 );
nand NAND2_17814 ( P2_R1143_U483 , P2_U3431 , P2_R1143_U72 );
nand NAND2_17815 ( P2_R1143_U484 , P2_U3078 , P2_R1143_U71 );
nand NAND2_17816 ( P2_R1143_U485 , P2_U3431 , P2_R1143_U72 );
nand NAND2_17817 ( P2_R1143_U486 , P2_R1143_U485 , P2_R1143_U484 );
nand NAND2_17818 ( P2_R1143_U487 , P2_R1143_U165 , P2_R1143_U166 );
nand NAND2_17819 ( P2_R1143_U488 , P2_R1143_U254 , P2_R1143_U486 );
nand NAND2_17820 ( P2_R1143_U489 , P2_U3079 , P2_R1143_U61 );
nand NAND2_17821 ( P2_R1143_U490 , P2_U3428 , P2_R1143_U62 );
nand NAND2_17822 ( P2_R1143_U491 , P2_U3071 , P2_R1143_U69 );
nand NAND2_17823 ( P2_R1143_U492 , P2_U3425 , P2_R1143_U70 );
nand NAND2_17824 ( P2_R1143_U493 , P2_R1143_U492 , P2_R1143_U491 );
nand NAND2_17825 ( P2_R1143_U494 , P2_R1143_U362 , P2_R1143_U93 );
nand NAND2_17826 ( P2_R1143_U495 , P2_R1143_U493 , P2_R1143_U338 );
nand NAND2_17827 ( P2_R1143_U496 , P2_U3062 , P2_R1143_U66 );
nand NAND2_17828 ( P2_R1143_U497 , P2_U3422 , P2_R1143_U67 );
nand NAND2_17829 ( P2_R1143_U498 , P2_R1143_U497 , P2_R1143_U496 );
nand NAND2_17830 ( P2_R1143_U499 , P2_R1143_U363 , P2_R1143_U167 );
nand NAND2_17831 ( P2_R1143_U500 , P2_R1143_U244 , P2_R1143_U498 );
nand NAND2_17832 ( P2_R1143_U501 , P2_U3061 , P2_R1143_U63 );
nand NAND2_17833 ( P2_R1143_U502 , P2_U3419 , P2_R1143_U64 );
nand NAND2_17834 ( P2_R1143_U503 , P2_U3076 , P2_R1143_U29 );
nand NAND2_17835 ( P2_R1143_U504 , P2_U3387 , P2_R1143_U30 );
and AND2_17836 ( P2_R1158_U4 , P2_R1158_U227 , P2_R1158_U226 );
and AND2_17837 ( P2_R1158_U5 , P2_R1158_U238 , P2_R1158_U237 );
and AND2_17838 ( P2_R1158_U6 , P2_R1158_U264 , P2_R1158_U263 );
and AND2_17839 ( P2_R1158_U7 , P2_R1158_U276 , P2_R1158_U275 );
and AND2_17840 ( P2_R1158_U8 , P2_R1158_U288 , P2_R1158_U287 );
and AND2_17841 ( P2_R1158_U9 , P2_R1158_U6 , P2_R1158_U268 );
and AND2_17842 ( P2_R1158_U10 , P2_R1158_U5 , P2_R1158_U235 );
and AND2_17843 ( P2_R1158_U11 , P2_R1158_U9 , P2_R1158_U261 );
and AND2_17844 ( P2_R1158_U12 , P2_R1158_U11 , P2_R1158_U271 );
and AND2_17845 ( P2_R1158_U13 , P2_R1158_U537 , P2_R1158_U536 );
and AND2_17846 ( P2_R1158_U14 , P2_R1158_U343 , P2_R1158_U340 );
and AND2_17847 ( P2_R1158_U15 , P2_R1158_U334 , P2_R1158_U331 );
and AND2_17848 ( P2_R1158_U16 , P2_R1158_U327 , P2_R1158_U324 );
and AND4_17849 ( P2_R1158_U17 , P2_R1158_U142 , P2_R1158_U394 , P2_R1158_U539 , P2_R1158_U538 );
and AND2_17850 ( P2_R1158_U18 , P2_R1158_U257 , P2_R1158_U254 );
and AND2_17851 ( P2_R1158_U19 , P2_R1158_U250 , P2_R1158_U247 );
nand NAND2_17852 ( P2_R1158_U20 , P2_U3056 , P2_R1158_U305 );
not NOT1_17853 ( P2_R1158_U21 , P2_U3152 );
not NOT1_17854 ( P2_R1158_U22 , P2_U3083 );
not NOT1_17855 ( P2_R1158_U23 , P2_U3070 );
nand NAND2_17856 ( P2_R1158_U24 , P2_U3070 , P2_R1158_U69 );
not NOT1_17857 ( P2_R1158_U25 , P2_U3069 );
not NOT1_17858 ( P2_R1158_U26 , P2_U3066 );
nand NAND2_17859 ( P2_R1158_U27 , P2_U3066 , P2_R1158_U71 );
not NOT1_17860 ( P2_R1158_U28 , P2_U3067 );
nand NAND2_17861 ( P2_R1158_U29 , P2_U3067 , P2_R1158_U72 );
not NOT1_17862 ( P2_R1158_U30 , P2_U3063 );
not NOT1_17863 ( P2_R1158_U31 , P2_U3077 );
not NOT1_17864 ( P2_R1158_U32 , P2_U3076 );
not NOT1_17865 ( P2_R1158_U33 , P2_U3059 );
not NOT1_17866 ( P2_R1158_U34 , P2_U3082 );
nand NAND3_17867 ( P2_R1158_U35 , P2_R1158_U242 , P2_R1158_U241 , P2_R1158_U359 );
nand NAND2_17868 ( P2_R1158_U36 , P2_R1158_U386 , P2_R1158_U27 );
nand NAND3_17869 ( P2_R1158_U37 , P2_R1158_U358 , P2_R1158_U224 , P2_R1158_U357 );
not NOT1_17870 ( P2_R1158_U38 , P2_U3052 );
not NOT1_17871 ( P2_R1158_U39 , P2_U3057 );
not NOT1_17872 ( P2_R1158_U40 , P2_U3064 );
not NOT1_17873 ( P2_R1158_U41 , P2_U3056 );
not NOT1_17874 ( P2_R1158_U42 , P2_U3072 );
nand NAND2_17875 ( P2_R1158_U43 , P2_U3072 , P2_R1158_U81 );
not NOT1_17876 ( P2_R1158_U44 , P2_U3068 );
not NOT1_17877 ( P2_R1158_U45 , P2_U3073 );
not NOT1_17878 ( P2_R1158_U46 , P2_U3078 );
not NOT1_17879 ( P2_R1158_U47 , P2_U3071 );
not NOT1_17880 ( P2_R1158_U48 , P2_U3062 );
nand NAND2_17881 ( P2_R1158_U49 , P2_U3062 , P2_R1158_U87 );
not NOT1_17882 ( P2_R1158_U50 , P2_U3079 );
not NOT1_17883 ( P2_R1158_U51 , P2_U3061 );
nand NAND2_17884 ( P2_R1158_U52 , P2_U3061 , P2_R1158_U88 );
not NOT1_17885 ( P2_R1158_U53 , P2_U3081 );
not NOT1_17886 ( P2_R1158_U54 , P2_U3075 );
not NOT1_17887 ( P2_R1158_U55 , P2_U3080 );
nand NAND2_17888 ( P2_R1158_U56 , P2_U3080 , P2_R1158_U90 );
not NOT1_17889 ( P2_R1158_U57 , P2_U3074 );
not NOT1_17890 ( P2_R1158_U58 , P2_U3060 );
not NOT1_17891 ( P2_R1158_U59 , P2_U3065 );
nand NAND2_17892 ( P2_R1158_U60 , P2_U3057 , P2_R1158_U78 );
nand NAND2_17893 ( P2_R1158_U61 , P2_R1158_U308 , P2_R1158_U192 );
nand NAND2_17894 ( P2_R1158_U62 , P2_R1158_U56 , P2_R1158_U320 );
nand NAND2_17895 ( P2_R1158_U63 , P2_R1158_U129 , P2_R1158_U384 );
nand NAND2_17896 ( P2_R1158_U64 , P2_R1158_U364 , P2_R1158_U272 );
nand NAND2_17897 ( P2_R1158_U65 , P2_R1158_U362 , P2_R1158_U270 );
nand NAND2_17898 ( P2_R1158_U66 , P2_R1158_U49 , P2_R1158_U336 );
nand NAND2_17899 ( P2_R1158_U67 , P2_R1158_U396 , P2_R1158_U395 );
nand NAND2_17900 ( P2_R1158_U68 , P2_R1158_U428 , P2_R1158_U427 );
nand NAND2_17901 ( P2_R1158_U69 , P2_R1158_U425 , P2_R1158_U424 );
nand NAND2_17902 ( P2_R1158_U70 , P2_R1158_U422 , P2_R1158_U421 );
nand NAND2_17903 ( P2_R1158_U71 , P2_R1158_U419 , P2_R1158_U418 );
nand NAND2_17904 ( P2_R1158_U72 , P2_R1158_U416 , P2_R1158_U415 );
nand NAND2_17905 ( P2_R1158_U73 , P2_R1158_U413 , P2_R1158_U412 );
nand NAND2_17906 ( P2_R1158_U74 , P2_R1158_U407 , P2_R1158_U406 );
nand NAND2_17907 ( P2_R1158_U75 , P2_R1158_U410 , P2_R1158_U409 );
nand NAND2_17908 ( P2_R1158_U76 , P2_R1158_U404 , P2_R1158_U403 );
nand NAND2_17909 ( P2_R1158_U77 , P2_R1158_U468 , P2_R1158_U467 );
nand NAND2_17910 ( P2_R1158_U78 , P2_R1158_U516 , P2_R1158_U515 );
nand NAND2_17911 ( P2_R1158_U79 , P2_R1158_U519 , P2_R1158_U518 );
nand NAND2_17912 ( P2_R1158_U80 , P2_R1158_U513 , P2_R1158_U512 );
nand NAND2_17913 ( P2_R1158_U81 , P2_R1158_U492 , P2_R1158_U491 );
nand NAND2_17914 ( P2_R1158_U82 , P2_R1158_U489 , P2_R1158_U488 );
nand NAND2_17915 ( P2_R1158_U83 , P2_R1158_U486 , P2_R1158_U485 );
nand NAND2_17916 ( P2_R1158_U84 , P2_R1158_U471 , P2_R1158_U470 );
nand NAND2_17917 ( P2_R1158_U85 , P2_R1158_U483 , P2_R1158_U482 );
nand NAND2_17918 ( P2_R1158_U86 , P2_R1158_U480 , P2_R1158_U479 );
nand NAND2_17919 ( P2_R1158_U87 , P2_R1158_U477 , P2_R1158_U476 );
nand NAND2_17920 ( P2_R1158_U88 , P2_R1158_U474 , P2_R1158_U473 );
nand NAND2_17921 ( P2_R1158_U89 , P2_R1158_U495 , P2_R1158_U494 );
nand NAND2_17922 ( P2_R1158_U90 , P2_R1158_U504 , P2_R1158_U503 );
nand NAND2_17923 ( P2_R1158_U91 , P2_R1158_U498 , P2_R1158_U497 );
nand NAND2_17924 ( P2_R1158_U92 , P2_R1158_U501 , P2_R1158_U500 );
nand NAND2_17925 ( P2_R1158_U93 , P2_R1158_U507 , P2_R1158_U506 );
nand NAND2_17926 ( P2_R1158_U94 , P2_R1158_U510 , P2_R1158_U509 );
nand NAND2_17927 ( P2_R1158_U95 , P2_R1158_U525 , P2_R1158_U524 );
nand NAND2_17928 ( P2_R1158_U96 , P2_R1158_U634 , P2_R1158_U633 );
nand NAND2_17929 ( P2_R1158_U97 , P2_R1158_U431 , P2_R1158_U430 );
nand NAND2_17930 ( P2_R1158_U98 , P2_R1158_U438 , P2_R1158_U437 );
nand NAND2_17931 ( P2_R1158_U99 , P2_R1158_U445 , P2_R1158_U444 );
nand NAND2_17932 ( P2_R1158_U100 , P2_R1158_U452 , P2_R1158_U451 );
nand NAND2_17933 ( P2_R1158_U101 , P2_R1158_U459 , P2_R1158_U458 );
nand NAND2_17934 ( P2_R1158_U102 , P2_R1158_U466 , P2_R1158_U465 );
nand NAND2_17935 ( P2_R1158_U103 , P2_R1158_U528 , P2_R1158_U527 );
nand NAND2_17936 ( P2_R1158_U104 , P2_R1158_U535 , P2_R1158_U534 );
nand NAND2_17937 ( P2_R1158_U105 , P2_R1158_U544 , P2_R1158_U543 );
nand NAND2_17938 ( P2_R1158_U106 , P2_R1158_U549 , P2_R1158_U548 );
nand NAND2_17939 ( P2_R1158_U107 , P2_R1158_U556 , P2_R1158_U555 );
nand NAND2_17940 ( P2_R1158_U108 , P2_R1158_U563 , P2_R1158_U562 );
nand NAND2_17941 ( P2_R1158_U109 , P2_R1158_U570 , P2_R1158_U569 );
nand NAND2_17942 ( P2_R1158_U110 , P2_R1158_U577 , P2_R1158_U576 );
nand NAND2_17943 ( P2_R1158_U111 , P2_R1158_U582 , P2_R1158_U581 );
nand NAND2_17944 ( P2_R1158_U112 , P2_R1158_U589 , P2_R1158_U588 );
nand NAND2_17945 ( P2_R1158_U113 , P2_R1158_U596 , P2_R1158_U595 );
nand NAND2_17946 ( P2_R1158_U114 , P2_R1158_U603 , P2_R1158_U602 );
nand NAND2_17947 ( P2_R1158_U115 , P2_R1158_U610 , P2_R1158_U609 );
nand NAND2_17948 ( P2_R1158_U116 , P2_R1158_U617 , P2_R1158_U616 );
nand NAND2_17949 ( P2_R1158_U117 , P2_R1158_U622 , P2_R1158_U621 );
nand NAND2_17950 ( P2_R1158_U118 , P2_R1158_U629 , P2_R1158_U628 );
and AND2_17951 ( P2_R1158_U119 , P2_R1158_U75 , P2_U3152 );
and AND2_17952 ( P2_R1158_U120 , P2_R1158_U230 , P2_R1158_U229 );
and AND2_17953 ( P2_R1158_U121 , P2_R1158_U243 , P2_R1158_U10 );
and AND2_17954 ( P2_R1158_U122 , P2_R1158_U361 , P2_R1158_U244 );
and AND3_17955 ( P2_R1158_U123 , P2_R1158_U440 , P2_R1158_U439 , P2_R1158_U24 );
and AND2_17956 ( P2_R1158_U124 , P2_R1158_U249 , P2_R1158_U5 );
and AND3_17957 ( P2_R1158_U125 , P2_R1158_U461 , P2_R1158_U460 , P2_R1158_U29 );
and AND2_17958 ( P2_R1158_U126 , P2_R1158_U256 , P2_R1158_U4 );
and AND2_17959 ( P2_R1158_U127 , P2_R1158_U266 , P2_R1158_U213 );
and AND2_17960 ( P2_R1158_U128 , P2_R1158_U273 , P2_R1158_U12 );
and AND2_17961 ( P2_R1158_U129 , P2_R1158_U372 , P2_R1158_U274 );
and AND2_17962 ( P2_R1158_U130 , P2_R1158_U280 , P2_R1158_U279 );
and AND2_17963 ( P2_R1158_U131 , P2_R1158_U292 , P2_R1158_U8 );
and AND2_17964 ( P2_R1158_U132 , P2_R1158_U290 , P2_R1158_U214 );
and AND2_17965 ( P2_R1158_U133 , P2_R1158_U313 , P2_R1158_U375 );
and AND2_17966 ( P2_R1158_U134 , P2_R1158_U315 , P2_R1158_U306 );
and AND2_17967 ( P2_R1158_U135 , P2_R1158_U315 , P2_R1158_U369 );
and AND2_17968 ( P2_R1158_U136 , P2_R1158_U373 , P2_R1158_U314 );
nand NAND2_17969 ( P2_R1158_U137 , P2_R1158_U522 , P2_R1158_U521 );
and AND2_17970 ( P2_R1158_U138 , P2_R1158_U318 , P2_R1158_U215 );
and AND2_17971 ( P2_R1158_U139 , P2_R1158_U517 , P2_R1158_U39 );
and AND2_17972 ( P2_R1158_U140 , P2_R1158_U318 , P2_R1158_U209 );
and AND2_17973 ( P2_R1158_U141 , P2_R1158_U13 , P2_R1158_U60 );
and AND2_17974 ( P2_R1158_U142 , P2_R1158_U393 , P2_R1158_U392 );
and AND3_17975 ( P2_R1158_U143 , P2_R1158_U565 , P2_R1158_U564 , P2_R1158_U214 );
and AND2_17976 ( P2_R1158_U144 , P2_R1158_U326 , P2_R1158_U8 );
and AND3_17977 ( P2_R1158_U145 , P2_R1158_U591 , P2_R1158_U590 , P2_R1158_U43 );
and AND2_17978 ( P2_R1158_U146 , P2_R1158_U333 , P2_R1158_U7 );
and AND3_17979 ( P2_R1158_U147 , P2_R1158_U612 , P2_R1158_U611 , P2_R1158_U213 );
and AND2_17980 ( P2_R1158_U148 , P2_R1158_U342 , P2_R1158_U6 );
nand NAND2_17981 ( P2_R1158_U149 , P2_R1158_U631 , P2_R1158_U630 );
not NOT1_17982 ( P2_R1158_U150 , P2_U3416 );
and AND2_17983 ( P2_R1158_U151 , P2_R1158_U399 , P2_R1158_U398 );
not NOT1_17984 ( P2_R1158_U152 , P2_U3401 );
not NOT1_17985 ( P2_R1158_U153 , P2_U3392 );
not NOT1_17986 ( P2_R1158_U154 , P2_U3387 );
not NOT1_17987 ( P2_R1158_U155 , P2_U3398 );
not NOT1_17988 ( P2_R1158_U156 , P2_U3395 );
not NOT1_17989 ( P2_R1158_U157 , P2_U3404 );
not NOT1_17990 ( P2_R1158_U158 , P2_U3410 );
not NOT1_17991 ( P2_R1158_U159 , P2_U3407 );
not NOT1_17992 ( P2_R1158_U160 , P2_U3413 );
nand NAND2_17993 ( P2_R1158_U161 , P2_R1158_U122 , P2_R1158_U390 );
and AND2_17994 ( P2_R1158_U162 , P2_R1158_U433 , P2_R1158_U432 );
nand NAND2_17995 ( P2_R1158_U163 , P2_R1158_U360 , P2_R1158_U388 );
and AND2_17996 ( P2_R1158_U164 , P2_R1158_U447 , P2_R1158_U446 );
nand NAND3_17997 ( P2_R1158_U165 , P2_R1158_U233 , P2_R1158_U211 , P2_R1158_U354 );
and AND2_17998 ( P2_R1158_U166 , P2_R1158_U454 , P2_R1158_U453 );
nand NAND2_17999 ( P2_R1158_U167 , P2_R1158_U120 , P2_R1158_U231 );
not NOT1_18000 ( P2_R1158_U168 , P2_U3896 );
not NOT1_18001 ( P2_R1158_U169 , P2_U3431 );
not NOT1_18002 ( P2_R1158_U170 , P2_U3419 );
not NOT1_18003 ( P2_R1158_U171 , P2_U3422 );
not NOT1_18004 ( P2_R1158_U172 , P2_U3428 );
not NOT1_18005 ( P2_R1158_U173 , P2_U3425 );
not NOT1_18006 ( P2_R1158_U174 , P2_U3434 );
not NOT1_18007 ( P2_R1158_U175 , P2_U3440 );
not NOT1_18008 ( P2_R1158_U176 , P2_U3437 );
not NOT1_18009 ( P2_R1158_U177 , P2_U3443 );
not NOT1_18010 ( P2_R1158_U178 , P2_U3902 );
not NOT1_18011 ( P2_R1158_U179 , P2_U3903 );
not NOT1_18012 ( P2_R1158_U180 , P2_U3445 );
not NOT1_18013 ( P2_R1158_U181 , P2_U3901 );
not NOT1_18014 ( P2_R1158_U182 , P2_U3900 );
not NOT1_18015 ( P2_R1158_U183 , P2_U3897 );
not NOT1_18016 ( P2_R1158_U184 , P2_U3898 );
not NOT1_18017 ( P2_R1158_U185 , P2_U3899 );
not NOT1_18018 ( P2_R1158_U186 , P2_U3053 );
not NOT1_18019 ( P2_R1158_U187 , P2_U3895 );
and AND2_18020 ( P2_R1158_U188 , P2_R1158_U530 , P2_R1158_U529 );
nand NAND2_18021 ( P2_R1158_U189 , P2_R1158_U310 , P2_R1158_U309 );
nand NAND2_18022 ( P2_R1158_U190 , P2_U3064 , P2_R1158_U79 );
nand NAND2_18023 ( P2_R1158_U191 , P2_R1158_U190 , P2_R1158_U61 );
nand NAND2_18024 ( P2_R1158_U192 , P2_R1158_U303 , P2_R1158_U302 );
and AND2_18025 ( P2_R1158_U193 , P2_R1158_U551 , P2_R1158_U550 );
nand NAND2_18026 ( P2_R1158_U194 , P2_R1158_U299 , P2_R1158_U298 );
and AND2_18027 ( P2_R1158_U195 , P2_R1158_U558 , P2_R1158_U557 );
nand NAND2_18028 ( P2_R1158_U196 , P2_R1158_U295 , P2_R1158_U294 );
and AND2_18029 ( P2_R1158_U197 , P2_R1158_U572 , P2_R1158_U571 );
nand NAND2_18030 ( P2_R1158_U198 , P2_R1158_U221 , P2_R1158_U220 );
nand NAND2_18031 ( P2_R1158_U199 , P2_R1158_U285 , P2_R1158_U284 );
and AND2_18032 ( P2_R1158_U200 , P2_R1158_U584 , P2_R1158_U583 );
nand NAND2_18033 ( P2_R1158_U201 , P2_R1158_U130 , P2_R1158_U281 );
and AND2_18034 ( P2_R1158_U202 , P2_R1158_U598 , P2_R1158_U597 );
nand NAND2_18035 ( P2_R1158_U203 , P2_R1158_U368 , P2_R1158_U382 );
and AND2_18036 ( P2_R1158_U204 , P2_R1158_U605 , P2_R1158_U604 );
nand NAND2_18037 ( P2_R1158_U205 , P2_R1158_U363 , P2_R1158_U380 );
nand NAND2_18038 ( P2_R1158_U206 , P2_R1158_U378 , P2_R1158_U52 );
and AND2_18039 ( P2_R1158_U207 , P2_R1158_U624 , P2_R1158_U623 );
nand NAND3_18040 ( P2_R1158_U208 , P2_R1158_U259 , P2_R1158_U210 , P2_R1158_U355 );
nand NAND2_18041 ( P2_R1158_U209 , P2_R1158_U20 , P2_R1158_U366 );
nand NAND2_18042 ( P2_R1158_U210 , P2_R1158_U67 , P2_R1158_U161 );
nand NAND2_18043 ( P2_R1158_U211 , P2_R1158_U76 , P2_R1158_U167 );
not NOT1_18044 ( P2_R1158_U212 , P2_R1158_U29 );
nand NAND2_18045 ( P2_R1158_U213 , P2_U3071 , P2_R1158_U85 );
nand NAND2_18046 ( P2_R1158_U214 , P2_U3075 , P2_R1158_U92 );
not NOT1_18047 ( P2_R1158_U215 , P2_R1158_U60 );
not NOT1_18048 ( P2_R1158_U216 , P2_R1158_U49 );
not NOT1_18049 ( P2_R1158_U217 , P2_R1158_U56 );
not NOT1_18050 ( P2_R1158_U218 , P2_R1158_U190 );
nand NAND2_18051 ( P2_R1158_U219 , P2_R1158_U411 , P2_R1158_U21 );
nand NAND2_18052 ( P2_R1158_U220 , P2_U3076 , P2_R1158_U219 );
nand NAND2_18053 ( P2_R1158_U221 , P2_U3152 , P2_R1158_U75 );
not NOT1_18054 ( P2_R1158_U222 , P2_R1158_U198 );
nand NAND2_18055 ( P2_R1158_U223 , P2_R1158_U408 , P2_R1158_U31 );
nand NAND2_18056 ( P2_R1158_U224 , P2_U3077 , P2_R1158_U74 );
not NOT1_18057 ( P2_R1158_U225 , P2_R1158_U37 );
nand NAND2_18058 ( P2_R1158_U226 , P2_R1158_U414 , P2_R1158_U30 );
nand NAND2_18059 ( P2_R1158_U227 , P2_R1158_U417 , P2_R1158_U28 );
nand NAND2_18060 ( P2_R1158_U228 , P2_R1158_U30 , P2_R1158_U29 );
nand NAND2_18061 ( P2_R1158_U229 , P2_R1158_U73 , P2_R1158_U228 );
nand NAND2_18062 ( P2_R1158_U230 , P2_U3063 , P2_R1158_U212 );
nand NAND2_18063 ( P2_R1158_U231 , P2_R1158_U4 , P2_R1158_U37 );
not NOT1_18064 ( P2_R1158_U232 , P2_R1158_U167 );
nand NAND2_18065 ( P2_R1158_U233 , P2_U3059 , P2_R1158_U167 );
not NOT1_18066 ( P2_R1158_U234 , P2_R1158_U165 );
nand NAND2_18067 ( P2_R1158_U235 , P2_R1158_U420 , P2_R1158_U26 );
not NOT1_18068 ( P2_R1158_U236 , P2_R1158_U27 );
nand NAND2_18069 ( P2_R1158_U237 , P2_R1158_U423 , P2_R1158_U25 );
nand NAND2_18070 ( P2_R1158_U238 , P2_R1158_U426 , P2_R1158_U23 );
not NOT1_18071 ( P2_R1158_U239 , P2_R1158_U24 );
nand NAND2_18072 ( P2_R1158_U240 , P2_R1158_U25 , P2_R1158_U24 );
nand NAND2_18073 ( P2_R1158_U241 , P2_R1158_U70 , P2_R1158_U240 );
nand NAND2_18074 ( P2_R1158_U242 , P2_U3069 , P2_R1158_U239 );
nand NAND2_18075 ( P2_R1158_U243 , P2_R1158_U429 , P2_R1158_U22 );
nand NAND2_18076 ( P2_R1158_U244 , P2_U3083 , P2_R1158_U68 );
nand NAND2_18077 ( P2_R1158_U245 , P2_R1158_U426 , P2_R1158_U23 );
nand NAND2_18078 ( P2_R1158_U246 , P2_R1158_U245 , P2_R1158_U36 );
nand NAND2_18079 ( P2_R1158_U247 , P2_R1158_U123 , P2_R1158_U246 );
nand NAND2_18080 ( P2_R1158_U248 , P2_R1158_U387 , P2_R1158_U24 );
nand NAND2_18081 ( P2_R1158_U249 , P2_U3069 , P2_R1158_U70 );
nand NAND2_18082 ( P2_R1158_U250 , P2_R1158_U124 , P2_R1158_U248 );
nand NAND2_18083 ( P2_R1158_U251 , P2_R1158_U426 , P2_R1158_U23 );
nand NAND2_18084 ( P2_R1158_U252 , P2_R1158_U417 , P2_R1158_U28 );
nand NAND2_18085 ( P2_R1158_U253 , P2_R1158_U252 , P2_R1158_U37 );
nand NAND2_18086 ( P2_R1158_U254 , P2_R1158_U125 , P2_R1158_U253 );
nand NAND2_18087 ( P2_R1158_U255 , P2_R1158_U225 , P2_R1158_U29 );
nand NAND2_18088 ( P2_R1158_U256 , P2_U3063 , P2_R1158_U73 );
nand NAND2_18089 ( P2_R1158_U257 , P2_R1158_U126 , P2_R1158_U255 );
nand NAND2_18090 ( P2_R1158_U258 , P2_R1158_U417 , P2_R1158_U28 );
nand NAND2_18091 ( P2_R1158_U259 , P2_U3082 , P2_R1158_U161 );
not NOT1_18092 ( P2_R1158_U260 , P2_R1158_U208 );
nand NAND2_18093 ( P2_R1158_U261 , P2_R1158_U475 , P2_R1158_U51 );
not NOT1_18094 ( P2_R1158_U262 , P2_R1158_U52 );
nand NAND2_18095 ( P2_R1158_U263 , P2_R1158_U481 , P2_R1158_U50 );
nand NAND2_18096 ( P2_R1158_U264 , P2_R1158_U484 , P2_R1158_U47 );
nand NAND2_18097 ( P2_R1158_U265 , P2_R1158_U216 , P2_R1158_U6 );
nand NAND2_18098 ( P2_R1158_U266 , P2_U3079 , P2_R1158_U86 );
nand NAND2_18099 ( P2_R1158_U267 , P2_R1158_U127 , P2_R1158_U265 );
nand NAND2_18100 ( P2_R1158_U268 , P2_R1158_U478 , P2_R1158_U48 );
nand NAND2_18101 ( P2_R1158_U269 , P2_R1158_U481 , P2_R1158_U50 );
nand NAND2_18102 ( P2_R1158_U270 , P2_R1158_U269 , P2_R1158_U267 );
nand NAND2_18103 ( P2_R1158_U271 , P2_R1158_U472 , P2_R1158_U46 );
nand NAND2_18104 ( P2_R1158_U272 , P2_U3078 , P2_R1158_U84 );
nand NAND2_18105 ( P2_R1158_U273 , P2_R1158_U487 , P2_R1158_U45 );
nand NAND2_18106 ( P2_R1158_U274 , P2_U3073 , P2_R1158_U83 );
nand NAND2_18107 ( P2_R1158_U275 , P2_R1158_U490 , P2_R1158_U44 );
nand NAND2_18108 ( P2_R1158_U276 , P2_R1158_U493 , P2_R1158_U42 );
not NOT1_18109 ( P2_R1158_U277 , P2_R1158_U43 );
nand NAND2_18110 ( P2_R1158_U278 , P2_R1158_U44 , P2_R1158_U43 );
nand NAND2_18111 ( P2_R1158_U279 , P2_R1158_U82 , P2_R1158_U278 );
nand NAND2_18112 ( P2_R1158_U280 , P2_U3068 , P2_R1158_U277 );
nand NAND2_18113 ( P2_R1158_U281 , P2_R1158_U7 , P2_R1158_U63 );
not NOT1_18114 ( P2_R1158_U282 , P2_R1158_U201 );
nand NAND2_18115 ( P2_R1158_U283 , P2_R1158_U496 , P2_R1158_U53 );
nand NAND2_18116 ( P2_R1158_U284 , P2_R1158_U283 , P2_R1158_U201 );
nand NAND2_18117 ( P2_R1158_U285 , P2_U3081 , P2_R1158_U89 );
not NOT1_18118 ( P2_R1158_U286 , P2_R1158_U199 );
nand NAND2_18119 ( P2_R1158_U287 , P2_R1158_U499 , P2_R1158_U57 );
nand NAND2_18120 ( P2_R1158_U288 , P2_R1158_U502 , P2_R1158_U54 );
nand NAND2_18121 ( P2_R1158_U289 , P2_R1158_U217 , P2_R1158_U8 );
nand NAND2_18122 ( P2_R1158_U290 , P2_U3074 , P2_R1158_U91 );
nand NAND2_18123 ( P2_R1158_U291 , P2_R1158_U132 , P2_R1158_U289 );
nand NAND2_18124 ( P2_R1158_U292 , P2_R1158_U505 , P2_R1158_U55 );
nand NAND2_18125 ( P2_R1158_U293 , P2_R1158_U499 , P2_R1158_U57 );
nand NAND2_18126 ( P2_R1158_U294 , P2_R1158_U131 , P2_R1158_U199 );
nand NAND2_18127 ( P2_R1158_U295 , P2_R1158_U293 , P2_R1158_U291 );
not NOT1_18128 ( P2_R1158_U296 , P2_R1158_U196 );
nand NAND2_18129 ( P2_R1158_U297 , P2_R1158_U508 , P2_R1158_U58 );
nand NAND2_18130 ( P2_R1158_U298 , P2_R1158_U297 , P2_R1158_U196 );
nand NAND2_18131 ( P2_R1158_U299 , P2_U3060 , P2_R1158_U93 );
not NOT1_18132 ( P2_R1158_U300 , P2_R1158_U194 );
nand NAND2_18133 ( P2_R1158_U301 , P2_R1158_U511 , P2_R1158_U59 );
nand NAND2_18134 ( P2_R1158_U302 , P2_R1158_U301 , P2_R1158_U194 );
nand NAND2_18135 ( P2_R1158_U303 , P2_U3065 , P2_R1158_U94 );
not NOT1_18136 ( P2_R1158_U304 , P2_R1158_U192 );
nand NAND2_18137 ( P2_R1158_U305 , P2_R1158_U517 , P2_R1158_U39 );
nand NAND3_18138 ( P2_R1158_U306 , P2_R1158_U190 , P2_R1158_U60 , P2_R1158_U307 );
nand NAND2_18139 ( P2_R1158_U307 , P2_U3056 , P2_R1158_U80 );
nand NAND2_18140 ( P2_R1158_U308 , P2_R1158_U520 , P2_R1158_U40 );
nand NAND2_18141 ( P2_R1158_U309 , P2_R1158_U369 , P2_R1158_U192 );
nand NAND2_18142 ( P2_R1158_U310 , P2_R1158_U365 , P2_R1158_U306 );
not NOT1_18143 ( P2_R1158_U311 , P2_R1158_U189 );
nand NAND2_18144 ( P2_R1158_U312 , P2_R1158_U469 , P2_R1158_U38 );
nand NAND2_18145 ( P2_R1158_U313 , P2_U3052 , P2_R1158_U77 );
nand NAND2_18146 ( P2_R1158_U314 , P2_U3052 , P2_R1158_U77 );
nand NAND2_18147 ( P2_R1158_U315 , P2_R1158_U469 , P2_R1158_U38 );
not NOT1_18148 ( P2_R1158_U316 , P2_R1158_U61 );
not NOT1_18149 ( P2_R1158_U317 , P2_R1158_U191 );
nand NAND2_18150 ( P2_R1158_U318 , P2_U3056 , P2_R1158_U80 );
nand NAND2_18151 ( P2_R1158_U319 , P2_R1158_U517 , P2_R1158_U39 );
nand NAND2_18152 ( P2_R1158_U320 , P2_R1158_U292 , P2_R1158_U199 );
not NOT1_18153 ( P2_R1158_U321 , P2_R1158_U62 );
nand NAND2_18154 ( P2_R1158_U322 , P2_R1158_U502 , P2_R1158_U54 );
nand NAND2_18155 ( P2_R1158_U323 , P2_R1158_U322 , P2_R1158_U62 );
nand NAND2_18156 ( P2_R1158_U324 , P2_R1158_U143 , P2_R1158_U323 );
nand NAND2_18157 ( P2_R1158_U325 , P2_R1158_U321 , P2_R1158_U214 );
nand NAND2_18158 ( P2_R1158_U326 , P2_U3074 , P2_R1158_U91 );
nand NAND2_18159 ( P2_R1158_U327 , P2_R1158_U144 , P2_R1158_U325 );
nand NAND2_18160 ( P2_R1158_U328 , P2_R1158_U502 , P2_R1158_U54 );
nand NAND2_18161 ( P2_R1158_U329 , P2_R1158_U493 , P2_R1158_U42 );
nand NAND2_18162 ( P2_R1158_U330 , P2_R1158_U329 , P2_R1158_U63 );
nand NAND2_18163 ( P2_R1158_U331 , P2_R1158_U145 , P2_R1158_U330 );
nand NAND2_18164 ( P2_R1158_U332 , P2_R1158_U385 , P2_R1158_U43 );
nand NAND2_18165 ( P2_R1158_U333 , P2_U3068 , P2_R1158_U82 );
nand NAND2_18166 ( P2_R1158_U334 , P2_R1158_U146 , P2_R1158_U332 );
nand NAND2_18167 ( P2_R1158_U335 , P2_R1158_U493 , P2_R1158_U42 );
nand NAND2_18168 ( P2_R1158_U336 , P2_R1158_U268 , P2_R1158_U206 );
not NOT1_18169 ( P2_R1158_U337 , P2_R1158_U66 );
nand NAND2_18170 ( P2_R1158_U338 , P2_R1158_U484 , P2_R1158_U47 );
nand NAND2_18171 ( P2_R1158_U339 , P2_R1158_U338 , P2_R1158_U66 );
nand NAND2_18172 ( P2_R1158_U340 , P2_R1158_U147 , P2_R1158_U339 );
nand NAND2_18173 ( P2_R1158_U341 , P2_R1158_U337 , P2_R1158_U213 );
nand NAND2_18174 ( P2_R1158_U342 , P2_U3079 , P2_R1158_U86 );
nand NAND2_18175 ( P2_R1158_U343 , P2_R1158_U148 , P2_R1158_U341 );
nand NAND2_18176 ( P2_R1158_U344 , P2_R1158_U484 , P2_R1158_U47 );
nand NAND2_18177 ( P2_R1158_U345 , P2_R1158_U251 , P2_R1158_U24 );
nand NAND2_18178 ( P2_R1158_U346 , P2_R1158_U258 , P2_R1158_U29 );
nand NAND2_18179 ( P2_R1158_U347 , P2_R1158_U319 , P2_R1158_U60 );
nand NAND2_18180 ( P2_R1158_U348 , P2_R1158_U308 , P2_R1158_U190 );
nand NAND2_18181 ( P2_R1158_U349 , P2_R1158_U328 , P2_R1158_U214 );
nand NAND2_18182 ( P2_R1158_U350 , P2_R1158_U292 , P2_R1158_U56 );
nand NAND2_18183 ( P2_R1158_U351 , P2_R1158_U335 , P2_R1158_U43 );
nand NAND2_18184 ( P2_R1158_U352 , P2_R1158_U344 , P2_R1158_U213 );
nand NAND2_18185 ( P2_R1158_U353 , P2_R1158_U268 , P2_R1158_U49 );
nand NAND2_18186 ( P2_R1158_U354 , P2_U3059 , P2_R1158_U76 );
nand NAND2_18187 ( P2_R1158_U355 , P2_U3082 , P2_R1158_U67 );
nand NAND2_18188 ( P2_R1158_U356 , P2_R1158_U133 , P2_R1158_U309 );
nand NAND3_18189 ( P2_R1158_U357 , P2_U3076 , P2_R1158_U219 , P2_R1158_U223 );
nand NAND2_18190 ( P2_R1158_U358 , P2_R1158_U119 , P2_R1158_U223 );
nand NAND2_18191 ( P2_R1158_U359 , P2_R1158_U236 , P2_R1158_U5 );
not NOT1_18192 ( P2_R1158_U360 , P2_R1158_U35 );
nand NAND2_18193 ( P2_R1158_U361 , P2_R1158_U35 , P2_R1158_U243 );
nand NAND2_18194 ( P2_R1158_U362 , P2_R1158_U262 , P2_R1158_U9 );
not NOT1_18195 ( P2_R1158_U363 , P2_R1158_U65 );
nand NAND2_18196 ( P2_R1158_U364 , P2_R1158_U65 , P2_R1158_U271 );
nand NAND3_18197 ( P2_R1158_U365 , P2_R1158_U366 , P2_R1158_U307 , P2_R1158_U20 );
nand NAND2_18198 ( P2_R1158_U366 , P2_R1158_U80 , P2_R1158_U305 );
not NOT1_18199 ( P2_R1158_U367 , P2_R1158_U20 );
not NOT1_18200 ( P2_R1158_U368 , P2_R1158_U64 );
nand NAND2_18201 ( P2_R1158_U369 , P2_R1158_U371 , P2_R1158_U370 );
nand NAND3_18202 ( P2_R1158_U370 , P2_R1158_U308 , P2_R1158_U305 , P2_R1158_U80 );
nand NAND2_18203 ( P2_R1158_U371 , P2_R1158_U367 , P2_R1158_U308 );
nand NAND2_18204 ( P2_R1158_U372 , P2_R1158_U64 , P2_R1158_U273 );
nand NAND2_18205 ( P2_R1158_U373 , P2_R1158_U134 , P2_R1158_U365 );
nand NAND2_18206 ( P2_R1158_U374 , P2_R1158_U135 , P2_R1158_U192 );
nand NAND2_18207 ( P2_R1158_U375 , P2_R1158_U377 , P2_R1158_U376 );
nand NAND3_18208 ( P2_R1158_U376 , P2_R1158_U190 , P2_R1158_U60 , P2_R1158_U307 );
nand NAND3_18209 ( P2_R1158_U377 , P2_R1158_U366 , P2_R1158_U307 , P2_R1158_U20 );
nand NAND2_18210 ( P2_R1158_U378 , P2_R1158_U261 , P2_R1158_U208 );
not NOT1_18211 ( P2_R1158_U379 , P2_R1158_U206 );
nand NAND2_18212 ( P2_R1158_U380 , P2_R1158_U11 , P2_R1158_U208 );
not NOT1_18213 ( P2_R1158_U381 , P2_R1158_U205 );
nand NAND2_18214 ( P2_R1158_U382 , P2_R1158_U12 , P2_R1158_U208 );
not NOT1_18215 ( P2_R1158_U383 , P2_R1158_U203 );
nand NAND2_18216 ( P2_R1158_U384 , P2_R1158_U128 , P2_R1158_U208 );
not NOT1_18217 ( P2_R1158_U385 , P2_R1158_U63 );
nand NAND2_18218 ( P2_R1158_U386 , P2_R1158_U235 , P2_R1158_U165 );
not NOT1_18219 ( P2_R1158_U387 , P2_R1158_U36 );
nand NAND2_18220 ( P2_R1158_U388 , P2_R1158_U10 , P2_R1158_U165 );
not NOT1_18221 ( P2_R1158_U389 , P2_R1158_U163 );
nand NAND2_18222 ( P2_R1158_U390 , P2_R1158_U121 , P2_R1158_U165 );
not NOT1_18223 ( P2_R1158_U391 , P2_R1158_U161 );
nand NAND2_18224 ( P2_R1158_U392 , P2_R1158_U138 , P2_R1158_U209 );
nand NAND2_18225 ( P2_R1158_U393 , P2_R1158_U139 , P2_R1158_U13 );
nand NAND2_18226 ( P2_R1158_U394 , P2_R1158_U140 , P2_R1158_U316 );
nand NAND2_18227 ( P2_R1158_U395 , P2_U3152 , P2_R1158_U150 );
nand NAND2_18228 ( P2_R1158_U396 , P2_U3416 , P2_R1158_U21 );
not NOT1_18229 ( P2_R1158_U397 , P2_R1158_U67 );
nand NAND2_18230 ( P2_R1158_U398 , P2_R1158_U397 , P2_U3082 );
nand NAND2_18231 ( P2_R1158_U399 , P2_R1158_U67 , P2_R1158_U34 );
nand NAND2_18232 ( P2_R1158_U400 , P2_R1158_U397 , P2_U3082 );
nand NAND2_18233 ( P2_R1158_U401 , P2_R1158_U67 , P2_R1158_U34 );
nand NAND2_18234 ( P2_R1158_U402 , P2_R1158_U401 , P2_R1158_U400 );
nand NAND2_18235 ( P2_R1158_U403 , P2_U3152 , P2_R1158_U152 );
nand NAND2_18236 ( P2_R1158_U404 , P2_U3401 , P2_R1158_U21 );
not NOT1_18237 ( P2_R1158_U405 , P2_R1158_U76 );
nand NAND2_18238 ( P2_R1158_U406 , P2_U3152 , P2_R1158_U153 );
nand NAND2_18239 ( P2_R1158_U407 , P2_U3392 , P2_R1158_U21 );
not NOT1_18240 ( P2_R1158_U408 , P2_R1158_U74 );
nand NAND2_18241 ( P2_R1158_U409 , P2_U3152 , P2_R1158_U154 );
nand NAND2_18242 ( P2_R1158_U410 , P2_U3387 , P2_R1158_U21 );
not NOT1_18243 ( P2_R1158_U411 , P2_R1158_U75 );
nand NAND2_18244 ( P2_R1158_U412 , P2_U3152 , P2_R1158_U155 );
nand NAND2_18245 ( P2_R1158_U413 , P2_U3398 , P2_R1158_U21 );
not NOT1_18246 ( P2_R1158_U414 , P2_R1158_U73 );
nand NAND2_18247 ( P2_R1158_U415 , P2_U3152 , P2_R1158_U156 );
nand NAND2_18248 ( P2_R1158_U416 , P2_U3395 , P2_R1158_U21 );
not NOT1_18249 ( P2_R1158_U417 , P2_R1158_U72 );
nand NAND2_18250 ( P2_R1158_U418 , P2_U3152 , P2_R1158_U157 );
nand NAND2_18251 ( P2_R1158_U419 , P2_U3404 , P2_R1158_U21 );
not NOT1_18252 ( P2_R1158_U420 , P2_R1158_U71 );
nand NAND2_18253 ( P2_R1158_U421 , P2_U3152 , P2_R1158_U158 );
nand NAND2_18254 ( P2_R1158_U422 , P2_U3410 , P2_R1158_U21 );
not NOT1_18255 ( P2_R1158_U423 , P2_R1158_U70 );
nand NAND2_18256 ( P2_R1158_U424 , P2_U3152 , P2_R1158_U159 );
nand NAND2_18257 ( P2_R1158_U425 , P2_U3407 , P2_R1158_U21 );
not NOT1_18258 ( P2_R1158_U426 , P2_R1158_U69 );
nand NAND2_18259 ( P2_R1158_U427 , P2_U3152 , P2_R1158_U160 );
nand NAND2_18260 ( P2_R1158_U428 , P2_U3413 , P2_R1158_U21 );
not NOT1_18261 ( P2_R1158_U429 , P2_R1158_U68 );
nand NAND2_18262 ( P2_R1158_U430 , P2_R1158_U151 , P2_R1158_U161 );
nand NAND2_18263 ( P2_R1158_U431 , P2_R1158_U391 , P2_R1158_U402 );
nand NAND2_18264 ( P2_R1158_U432 , P2_R1158_U429 , P2_U3083 );
nand NAND2_18265 ( P2_R1158_U433 , P2_R1158_U68 , P2_R1158_U22 );
nand NAND2_18266 ( P2_R1158_U434 , P2_R1158_U429 , P2_U3083 );
nand NAND2_18267 ( P2_R1158_U435 , P2_R1158_U68 , P2_R1158_U22 );
nand NAND2_18268 ( P2_R1158_U436 , P2_R1158_U435 , P2_R1158_U434 );
nand NAND2_18269 ( P2_R1158_U437 , P2_R1158_U162 , P2_R1158_U163 );
nand NAND2_18270 ( P2_R1158_U438 , P2_R1158_U389 , P2_R1158_U436 );
nand NAND2_18271 ( P2_R1158_U439 , P2_R1158_U423 , P2_U3069 );
nand NAND2_18272 ( P2_R1158_U440 , P2_R1158_U70 , P2_R1158_U25 );
nand NAND2_18273 ( P2_R1158_U441 , P2_R1158_U426 , P2_U3070 );
nand NAND2_18274 ( P2_R1158_U442 , P2_R1158_U69 , P2_R1158_U23 );
nand NAND2_18275 ( P2_R1158_U443 , P2_R1158_U442 , P2_R1158_U441 );
nand NAND2_18276 ( P2_R1158_U444 , P2_R1158_U36 , P2_R1158_U345 );
nand NAND2_18277 ( P2_R1158_U445 , P2_R1158_U443 , P2_R1158_U387 );
nand NAND2_18278 ( P2_R1158_U446 , P2_R1158_U420 , P2_U3066 );
nand NAND2_18279 ( P2_R1158_U447 , P2_R1158_U71 , P2_R1158_U26 );
nand NAND2_18280 ( P2_R1158_U448 , P2_R1158_U420 , P2_U3066 );
nand NAND2_18281 ( P2_R1158_U449 , P2_R1158_U71 , P2_R1158_U26 );
nand NAND2_18282 ( P2_R1158_U450 , P2_R1158_U449 , P2_R1158_U448 );
nand NAND2_18283 ( P2_R1158_U451 , P2_R1158_U164 , P2_R1158_U165 );
nand NAND2_18284 ( P2_R1158_U452 , P2_R1158_U234 , P2_R1158_U450 );
nand NAND2_18285 ( P2_R1158_U453 , P2_R1158_U405 , P2_U3059 );
nand NAND2_18286 ( P2_R1158_U454 , P2_R1158_U76 , P2_R1158_U33 );
nand NAND2_18287 ( P2_R1158_U455 , P2_R1158_U405 , P2_U3059 );
nand NAND2_18288 ( P2_R1158_U456 , P2_R1158_U76 , P2_R1158_U33 );
nand NAND2_18289 ( P2_R1158_U457 , P2_R1158_U456 , P2_R1158_U455 );
nand NAND2_18290 ( P2_R1158_U458 , P2_R1158_U166 , P2_R1158_U167 );
nand NAND2_18291 ( P2_R1158_U459 , P2_R1158_U232 , P2_R1158_U457 );
nand NAND2_18292 ( P2_R1158_U460 , P2_R1158_U414 , P2_U3063 );
nand NAND2_18293 ( P2_R1158_U461 , P2_R1158_U73 , P2_R1158_U30 );
nand NAND2_18294 ( P2_R1158_U462 , P2_R1158_U417 , P2_U3067 );
nand NAND2_18295 ( P2_R1158_U463 , P2_R1158_U72 , P2_R1158_U28 );
nand NAND2_18296 ( P2_R1158_U464 , P2_R1158_U463 , P2_R1158_U462 );
nand NAND2_18297 ( P2_R1158_U465 , P2_R1158_U346 , P2_R1158_U37 );
nand NAND2_18298 ( P2_R1158_U466 , P2_R1158_U464 , P2_R1158_U225 );
nand NAND2_18299 ( P2_R1158_U467 , P2_U3152 , P2_R1158_U168 );
nand NAND2_18300 ( P2_R1158_U468 , P2_U3896 , P2_R1158_U21 );
not NOT1_18301 ( P2_R1158_U469 , P2_R1158_U77 );
nand NAND2_18302 ( P2_R1158_U470 , P2_U3152 , P2_R1158_U169 );
nand NAND2_18303 ( P2_R1158_U471 , P2_U3431 , P2_R1158_U21 );
not NOT1_18304 ( P2_R1158_U472 , P2_R1158_U84 );
nand NAND2_18305 ( P2_R1158_U473 , P2_U3152 , P2_R1158_U170 );
nand NAND2_18306 ( P2_R1158_U474 , P2_U3419 , P2_R1158_U21 );
not NOT1_18307 ( P2_R1158_U475 , P2_R1158_U88 );
nand NAND2_18308 ( P2_R1158_U476 , P2_U3152 , P2_R1158_U171 );
nand NAND2_18309 ( P2_R1158_U477 , P2_U3422 , P2_R1158_U21 );
not NOT1_18310 ( P2_R1158_U478 , P2_R1158_U87 );
nand NAND2_18311 ( P2_R1158_U479 , P2_U3152 , P2_R1158_U172 );
nand NAND2_18312 ( P2_R1158_U480 , P2_U3428 , P2_R1158_U21 );
not NOT1_18313 ( P2_R1158_U481 , P2_R1158_U86 );
nand NAND2_18314 ( P2_R1158_U482 , P2_U3152 , P2_R1158_U173 );
nand NAND2_18315 ( P2_R1158_U483 , P2_U3425 , P2_R1158_U21 );
not NOT1_18316 ( P2_R1158_U484 , P2_R1158_U85 );
nand NAND2_18317 ( P2_R1158_U485 , P2_U3152 , P2_R1158_U174 );
nand NAND2_18318 ( P2_R1158_U486 , P2_U3434 , P2_R1158_U21 );
not NOT1_18319 ( P2_R1158_U487 , P2_R1158_U83 );
nand NAND2_18320 ( P2_R1158_U488 , P2_U3152 , P2_R1158_U175 );
nand NAND2_18321 ( P2_R1158_U489 , P2_U3440 , P2_R1158_U21 );
not NOT1_18322 ( P2_R1158_U490 , P2_R1158_U82 );
nand NAND2_18323 ( P2_R1158_U491 , P2_U3152 , P2_R1158_U176 );
nand NAND2_18324 ( P2_R1158_U492 , P2_U3437 , P2_R1158_U21 );
not NOT1_18325 ( P2_R1158_U493 , P2_R1158_U81 );
nand NAND2_18326 ( P2_R1158_U494 , P2_U3152 , P2_R1158_U177 );
nand NAND2_18327 ( P2_R1158_U495 , P2_U3443 , P2_R1158_U21 );
not NOT1_18328 ( P2_R1158_U496 , P2_R1158_U89 );
nand NAND2_18329 ( P2_R1158_U497 , P2_U3152 , P2_R1158_U178 );
nand NAND2_18330 ( P2_R1158_U498 , P2_U3902 , P2_R1158_U21 );
not NOT1_18331 ( P2_R1158_U499 , P2_R1158_U91 );
nand NAND2_18332 ( P2_R1158_U500 , P2_U3152 , P2_R1158_U179 );
nand NAND2_18333 ( P2_R1158_U501 , P2_U3903 , P2_R1158_U21 );
not NOT1_18334 ( P2_R1158_U502 , P2_R1158_U92 );
nand NAND2_18335 ( P2_R1158_U503 , P2_U3152 , P2_R1158_U180 );
nand NAND2_18336 ( P2_R1158_U504 , P2_U3445 , P2_R1158_U21 );
not NOT1_18337 ( P2_R1158_U505 , P2_R1158_U90 );
nand NAND2_18338 ( P2_R1158_U506 , P2_U3152 , P2_R1158_U181 );
nand NAND2_18339 ( P2_R1158_U507 , P2_U3901 , P2_R1158_U21 );
not NOT1_18340 ( P2_R1158_U508 , P2_R1158_U93 );
nand NAND2_18341 ( P2_R1158_U509 , P2_U3152 , P2_R1158_U182 );
nand NAND2_18342 ( P2_R1158_U510 , P2_U3900 , P2_R1158_U21 );
not NOT1_18343 ( P2_R1158_U511 , P2_R1158_U94 );
nand NAND2_18344 ( P2_R1158_U512 , P2_U3152 , P2_R1158_U183 );
nand NAND2_18345 ( P2_R1158_U513 , P2_U3897 , P2_R1158_U21 );
not NOT1_18346 ( P2_R1158_U514 , P2_R1158_U80 );
nand NAND2_18347 ( P2_R1158_U515 , P2_U3152 , P2_R1158_U184 );
nand NAND2_18348 ( P2_R1158_U516 , P2_U3898 , P2_R1158_U21 );
not NOT1_18349 ( P2_R1158_U517 , P2_R1158_U78 );
nand NAND2_18350 ( P2_R1158_U518 , P2_U3152 , P2_R1158_U185 );
nand NAND2_18351 ( P2_R1158_U519 , P2_U3899 , P2_R1158_U21 );
not NOT1_18352 ( P2_R1158_U520 , P2_R1158_U79 );
nand NAND2_18353 ( P2_R1158_U521 , P2_U3152 , P2_R1158_U186 );
nand NAND2_18354 ( P2_R1158_U522 , P2_U3053 , P2_R1158_U21 );
not NOT1_18355 ( P2_R1158_U523 , P2_R1158_U137 );
nand NAND2_18356 ( P2_R1158_U524 , P2_U3895 , P2_R1158_U523 );
nand NAND2_18357 ( P2_R1158_U525 , P2_R1158_U137 , P2_R1158_U187 );
not NOT1_18358 ( P2_R1158_U526 , P2_R1158_U95 );
nand NAND3_18359 ( P2_R1158_U527 , P2_R1158_U356 , P2_R1158_U312 , P2_R1158_U526 );
nand NAND3_18360 ( P2_R1158_U528 , P2_R1158_U136 , P2_R1158_U374 , P2_R1158_U95 );
nand NAND2_18361 ( P2_R1158_U529 , P2_R1158_U469 , P2_U3052 );
nand NAND2_18362 ( P2_R1158_U530 , P2_R1158_U77 , P2_R1158_U38 );
nand NAND2_18363 ( P2_R1158_U531 , P2_R1158_U469 , P2_U3052 );
nand NAND2_18364 ( P2_R1158_U532 , P2_R1158_U77 , P2_R1158_U38 );
nand NAND2_18365 ( P2_R1158_U533 , P2_R1158_U532 , P2_R1158_U531 );
nand NAND2_18366 ( P2_R1158_U534 , P2_R1158_U188 , P2_R1158_U189 );
nand NAND2_18367 ( P2_R1158_U535 , P2_R1158_U311 , P2_R1158_U533 );
nand NAND2_18368 ( P2_R1158_U536 , P2_R1158_U514 , P2_U3056 );
nand NAND2_18369 ( P2_R1158_U537 , P2_R1158_U80 , P2_R1158_U41 );
nand NAND3_18370 ( P2_R1158_U538 , P2_R1158_U141 , P2_R1158_U61 , P2_R1158_U190 );
nand NAND3_18371 ( P2_R1158_U539 , P2_R1158_U318 , P2_R1158_U209 , P2_R1158_U218 );
nand NAND2_18372 ( P2_R1158_U540 , P2_R1158_U517 , P2_U3057 );
nand NAND2_18373 ( P2_R1158_U541 , P2_R1158_U78 , P2_R1158_U39 );
nand NAND2_18374 ( P2_R1158_U542 , P2_R1158_U541 , P2_R1158_U540 );
nand NAND2_18375 ( P2_R1158_U543 , P2_R1158_U347 , P2_R1158_U191 );
nand NAND2_18376 ( P2_R1158_U544 , P2_R1158_U317 , P2_R1158_U542 );
nand NAND2_18377 ( P2_R1158_U545 , P2_R1158_U520 , P2_U3064 );
nand NAND2_18378 ( P2_R1158_U546 , P2_R1158_U79 , P2_R1158_U40 );
nand NAND2_18379 ( P2_R1158_U547 , P2_R1158_U546 , P2_R1158_U545 );
nand NAND2_18380 ( P2_R1158_U548 , P2_R1158_U348 , P2_R1158_U192 );
nand NAND2_18381 ( P2_R1158_U549 , P2_R1158_U304 , P2_R1158_U547 );
nand NAND2_18382 ( P2_R1158_U550 , P2_R1158_U511 , P2_U3065 );
nand NAND2_18383 ( P2_R1158_U551 , P2_R1158_U94 , P2_R1158_U59 );
nand NAND2_18384 ( P2_R1158_U552 , P2_R1158_U511 , P2_U3065 );
nand NAND2_18385 ( P2_R1158_U553 , P2_R1158_U94 , P2_R1158_U59 );
nand NAND2_18386 ( P2_R1158_U554 , P2_R1158_U553 , P2_R1158_U552 );
nand NAND2_18387 ( P2_R1158_U555 , P2_R1158_U193 , P2_R1158_U194 );
nand NAND2_18388 ( P2_R1158_U556 , P2_R1158_U300 , P2_R1158_U554 );
nand NAND2_18389 ( P2_R1158_U557 , P2_R1158_U508 , P2_U3060 );
nand NAND2_18390 ( P2_R1158_U558 , P2_R1158_U93 , P2_R1158_U58 );
nand NAND2_18391 ( P2_R1158_U559 , P2_R1158_U508 , P2_U3060 );
nand NAND2_18392 ( P2_R1158_U560 , P2_R1158_U93 , P2_R1158_U58 );
nand NAND2_18393 ( P2_R1158_U561 , P2_R1158_U560 , P2_R1158_U559 );
nand NAND2_18394 ( P2_R1158_U562 , P2_R1158_U195 , P2_R1158_U196 );
nand NAND2_18395 ( P2_R1158_U563 , P2_R1158_U296 , P2_R1158_U561 );
nand NAND2_18396 ( P2_R1158_U564 , P2_R1158_U499 , P2_U3074 );
nand NAND2_18397 ( P2_R1158_U565 , P2_R1158_U91 , P2_R1158_U57 );
nand NAND2_18398 ( P2_R1158_U566 , P2_R1158_U502 , P2_U3075 );
nand NAND2_18399 ( P2_R1158_U567 , P2_R1158_U92 , P2_R1158_U54 );
nand NAND2_18400 ( P2_R1158_U568 , P2_R1158_U567 , P2_R1158_U566 );
nand NAND2_18401 ( P2_R1158_U569 , P2_R1158_U349 , P2_R1158_U62 );
nand NAND2_18402 ( P2_R1158_U570 , P2_R1158_U568 , P2_R1158_U321 );
nand NAND2_18403 ( P2_R1158_U571 , P2_R1158_U408 , P2_U3077 );
nand NAND2_18404 ( P2_R1158_U572 , P2_R1158_U74 , P2_R1158_U31 );
nand NAND2_18405 ( P2_R1158_U573 , P2_R1158_U408 , P2_U3077 );
nand NAND2_18406 ( P2_R1158_U574 , P2_R1158_U74 , P2_R1158_U31 );
nand NAND2_18407 ( P2_R1158_U575 , P2_R1158_U574 , P2_R1158_U573 );
nand NAND2_18408 ( P2_R1158_U576 , P2_R1158_U197 , P2_R1158_U198 );
nand NAND2_18409 ( P2_R1158_U577 , P2_R1158_U222 , P2_R1158_U575 );
nand NAND2_18410 ( P2_R1158_U578 , P2_R1158_U505 , P2_U3080 );
nand NAND2_18411 ( P2_R1158_U579 , P2_R1158_U90 , P2_R1158_U55 );
nand NAND2_18412 ( P2_R1158_U580 , P2_R1158_U579 , P2_R1158_U578 );
nand NAND2_18413 ( P2_R1158_U581 , P2_R1158_U350 , P2_R1158_U199 );
nand NAND2_18414 ( P2_R1158_U582 , P2_R1158_U286 , P2_R1158_U580 );
nand NAND2_18415 ( P2_R1158_U583 , P2_R1158_U496 , P2_U3081 );
nand NAND2_18416 ( P2_R1158_U584 , P2_R1158_U89 , P2_R1158_U53 );
nand NAND2_18417 ( P2_R1158_U585 , P2_R1158_U496 , P2_U3081 );
nand NAND2_18418 ( P2_R1158_U586 , P2_R1158_U89 , P2_R1158_U53 );
nand NAND2_18419 ( P2_R1158_U587 , P2_R1158_U586 , P2_R1158_U585 );
nand NAND2_18420 ( P2_R1158_U588 , P2_R1158_U200 , P2_R1158_U201 );
nand NAND2_18421 ( P2_R1158_U589 , P2_R1158_U282 , P2_R1158_U587 );
nand NAND2_18422 ( P2_R1158_U590 , P2_R1158_U490 , P2_U3068 );
nand NAND2_18423 ( P2_R1158_U591 , P2_R1158_U82 , P2_R1158_U44 );
nand NAND2_18424 ( P2_R1158_U592 , P2_R1158_U493 , P2_U3072 );
nand NAND2_18425 ( P2_R1158_U593 , P2_R1158_U81 , P2_R1158_U42 );
nand NAND2_18426 ( P2_R1158_U594 , P2_R1158_U593 , P2_R1158_U592 );
nand NAND2_18427 ( P2_R1158_U595 , P2_R1158_U63 , P2_R1158_U351 );
nand NAND2_18428 ( P2_R1158_U596 , P2_R1158_U594 , P2_R1158_U385 );
nand NAND2_18429 ( P2_R1158_U597 , P2_R1158_U487 , P2_U3073 );
nand NAND2_18430 ( P2_R1158_U598 , P2_R1158_U83 , P2_R1158_U45 );
nand NAND2_18431 ( P2_R1158_U599 , P2_R1158_U487 , P2_U3073 );
nand NAND2_18432 ( P2_R1158_U600 , P2_R1158_U83 , P2_R1158_U45 );
nand NAND2_18433 ( P2_R1158_U601 , P2_R1158_U600 , P2_R1158_U599 );
nand NAND2_18434 ( P2_R1158_U602 , P2_R1158_U202 , P2_R1158_U203 );
nand NAND2_18435 ( P2_R1158_U603 , P2_R1158_U383 , P2_R1158_U601 );
nand NAND2_18436 ( P2_R1158_U604 , P2_R1158_U472 , P2_U3078 );
nand NAND2_18437 ( P2_R1158_U605 , P2_R1158_U84 , P2_R1158_U46 );
nand NAND2_18438 ( P2_R1158_U606 , P2_R1158_U472 , P2_U3078 );
nand NAND2_18439 ( P2_R1158_U607 , P2_R1158_U84 , P2_R1158_U46 );
nand NAND2_18440 ( P2_R1158_U608 , P2_R1158_U607 , P2_R1158_U606 );
nand NAND2_18441 ( P2_R1158_U609 , P2_R1158_U204 , P2_R1158_U205 );
nand NAND2_18442 ( P2_R1158_U610 , P2_R1158_U381 , P2_R1158_U608 );
nand NAND2_18443 ( P2_R1158_U611 , P2_R1158_U481 , P2_U3079 );
nand NAND2_18444 ( P2_R1158_U612 , P2_R1158_U86 , P2_R1158_U50 );
nand NAND2_18445 ( P2_R1158_U613 , P2_R1158_U484 , P2_U3071 );
nand NAND2_18446 ( P2_R1158_U614 , P2_R1158_U85 , P2_R1158_U47 );
nand NAND2_18447 ( P2_R1158_U615 , P2_R1158_U614 , P2_R1158_U613 );
nand NAND2_18448 ( P2_R1158_U616 , P2_R1158_U352 , P2_R1158_U66 );
nand NAND2_18449 ( P2_R1158_U617 , P2_R1158_U615 , P2_R1158_U337 );
nand NAND2_18450 ( P2_R1158_U618 , P2_R1158_U478 , P2_U3062 );
nand NAND2_18451 ( P2_R1158_U619 , P2_R1158_U87 , P2_R1158_U48 );
nand NAND2_18452 ( P2_R1158_U620 , P2_R1158_U619 , P2_R1158_U618 );
nand NAND2_18453 ( P2_R1158_U621 , P2_R1158_U206 , P2_R1158_U353 );
nand NAND2_18454 ( P2_R1158_U622 , P2_R1158_U379 , P2_R1158_U620 );
nand NAND2_18455 ( P2_R1158_U623 , P2_R1158_U475 , P2_U3061 );
nand NAND2_18456 ( P2_R1158_U624 , P2_R1158_U88 , P2_R1158_U51 );
nand NAND2_18457 ( P2_R1158_U625 , P2_R1158_U475 , P2_U3061 );
nand NAND2_18458 ( P2_R1158_U626 , P2_R1158_U88 , P2_R1158_U51 );
nand NAND2_18459 ( P2_R1158_U627 , P2_R1158_U626 , P2_R1158_U625 );
nand NAND2_18460 ( P2_R1158_U628 , P2_R1158_U207 , P2_R1158_U208 );
nand NAND2_18461 ( P2_R1158_U629 , P2_R1158_U260 , P2_R1158_U627 );
nand NAND2_18462 ( P2_R1158_U630 , P2_R1158_U75 , P2_R1158_U21 );
nand NAND2_18463 ( P2_R1158_U631 , P2_R1158_U411 , P2_U3152 );
not NOT1_18464 ( P2_R1158_U632 , P2_R1158_U149 );
nand NAND2_18465 ( P2_R1158_U633 , P2_R1158_U632 , P2_U3076 );
nand NAND2_18466 ( P2_R1158_U634 , P2_R1158_U149 , P2_R1158_U32 );
and AND2_18467 ( P2_R1131_U6 , P2_R1131_U212 , P2_R1131_U211 );
and AND2_18468 ( P2_R1131_U7 , P2_R1131_U246 , P2_R1131_U245 );
and AND2_18469 ( P2_R1131_U8 , P2_R1131_U193 , P2_R1131_U257 );
and AND2_18470 ( P2_R1131_U9 , P2_R1131_U259 , P2_R1131_U258 );
and AND2_18471 ( P2_R1131_U10 , P2_R1131_U194 , P2_R1131_U281 );
and AND2_18472 ( P2_R1131_U11 , P2_R1131_U283 , P2_R1131_U282 );
and AND2_18473 ( P2_R1131_U12 , P2_R1131_U299 , P2_R1131_U195 );
and AND3_18474 ( P2_R1131_U13 , P2_R1131_U210 , P2_R1131_U197 , P2_R1131_U215 );
and AND2_18475 ( P2_R1131_U14 , P2_R1131_U220 , P2_R1131_U198 );
and AND3_18476 ( P2_R1131_U15 , P2_R1131_U224 , P2_R1131_U192 , P2_R1131_U244 );
and AND2_18477 ( P2_R1131_U16 , P2_R1131_U399 , P2_R1131_U398 );
nand NAND2_18478 ( P2_R1131_U17 , P2_R1131_U331 , P2_R1131_U334 );
nand NAND2_18479 ( P2_R1131_U18 , P2_R1131_U322 , P2_R1131_U325 );
nand NAND2_18480 ( P2_R1131_U19 , P2_R1131_U311 , P2_R1131_U314 );
nand NAND2_18481 ( P2_R1131_U20 , P2_R1131_U305 , P2_R1131_U357 );
nand NAND2_18482 ( P2_R1131_U21 , P2_R1131_U137 , P2_R1131_U186 );
nand NAND2_18483 ( P2_R1131_U22 , P2_R1131_U242 , P2_R1131_U347 );
nand NAND2_18484 ( P2_R1131_U23 , P2_R1131_U235 , P2_R1131_U238 );
nand NAND2_18485 ( P2_R1131_U24 , P2_R1131_U227 , P2_R1131_U229 );
nand NAND2_18486 ( P2_R1131_U25 , P2_R1131_U175 , P2_R1131_U337 );
not NOT1_18487 ( P2_R1131_U26 , P2_U3069 );
nand NAND2_18488 ( P2_R1131_U27 , P2_U3069 , P2_R1131_U32 );
not NOT1_18489 ( P2_R1131_U28 , P2_U3083 );
not NOT1_18490 ( P2_R1131_U29 , P2_U3404 );
not NOT1_18491 ( P2_R1131_U30 , P2_U3407 );
not NOT1_18492 ( P2_R1131_U31 , P2_U3401 );
not NOT1_18493 ( P2_R1131_U32 , P2_U3410 );
not NOT1_18494 ( P2_R1131_U33 , P2_U3413 );
not NOT1_18495 ( P2_R1131_U34 , P2_U3067 );
nand NAND2_18496 ( P2_R1131_U35 , P2_U3067 , P2_R1131_U37 );
not NOT1_18497 ( P2_R1131_U36 , P2_U3063 );
not NOT1_18498 ( P2_R1131_U37 , P2_U3395 );
not NOT1_18499 ( P2_R1131_U38 , P2_U3387 );
not NOT1_18500 ( P2_R1131_U39 , P2_U3077 );
not NOT1_18501 ( P2_R1131_U40 , P2_U3398 );
not NOT1_18502 ( P2_R1131_U41 , P2_U3070 );
not NOT1_18503 ( P2_R1131_U42 , P2_U3066 );
not NOT1_18504 ( P2_R1131_U43 , P2_U3059 );
nand NAND2_18505 ( P2_R1131_U44 , P2_U3059 , P2_R1131_U31 );
nand NAND2_18506 ( P2_R1131_U45 , P2_R1131_U216 , P2_R1131_U214 );
not NOT1_18507 ( P2_R1131_U46 , P2_U3416 );
not NOT1_18508 ( P2_R1131_U47 , P2_U3082 );
nand NAND2_18509 ( P2_R1131_U48 , P2_R1131_U45 , P2_R1131_U217 );
nand NAND2_18510 ( P2_R1131_U49 , P2_R1131_U44 , P2_R1131_U231 );
nand NAND3_18511 ( P2_R1131_U50 , P2_R1131_U204 , P2_R1131_U188 , P2_R1131_U338 );
not NOT1_18512 ( P2_R1131_U51 , P2_U3895 );
not NOT1_18513 ( P2_R1131_U52 , P2_U3056 );
nand NAND2_18514 ( P2_R1131_U53 , P2_U3056 , P2_R1131_U90 );
not NOT1_18515 ( P2_R1131_U54 , P2_U3052 );
not NOT1_18516 ( P2_R1131_U55 , P2_U3071 );
not NOT1_18517 ( P2_R1131_U56 , P2_U3062 );
not NOT1_18518 ( P2_R1131_U57 , P2_U3061 );
not NOT1_18519 ( P2_R1131_U58 , P2_U3419 );
nand NAND2_18520 ( P2_R1131_U59 , P2_U3082 , P2_R1131_U46 );
not NOT1_18521 ( P2_R1131_U60 , P2_U3422 );
not NOT1_18522 ( P2_R1131_U61 , P2_U3425 );
nand NAND2_18523 ( P2_R1131_U62 , P2_R1131_U249 , P2_R1131_U248 );
not NOT1_18524 ( P2_R1131_U63 , P2_U3428 );
not NOT1_18525 ( P2_R1131_U64 , P2_U3079 );
not NOT1_18526 ( P2_R1131_U65 , P2_U3437 );
not NOT1_18527 ( P2_R1131_U66 , P2_U3434 );
not NOT1_18528 ( P2_R1131_U67 , P2_U3431 );
not NOT1_18529 ( P2_R1131_U68 , P2_U3072 );
not NOT1_18530 ( P2_R1131_U69 , P2_U3073 );
not NOT1_18531 ( P2_R1131_U70 , P2_U3078 );
nand NAND2_18532 ( P2_R1131_U71 , P2_U3078 , P2_R1131_U67 );
not NOT1_18533 ( P2_R1131_U72 , P2_U3440 );
not NOT1_18534 ( P2_R1131_U73 , P2_U3068 );
not NOT1_18535 ( P2_R1131_U74 , P2_U3081 );
not NOT1_18536 ( P2_R1131_U75 , P2_U3445 );
not NOT1_18537 ( P2_R1131_U76 , P2_U3080 );
not NOT1_18538 ( P2_R1131_U77 , P2_U3903 );
not NOT1_18539 ( P2_R1131_U78 , P2_U3075 );
not NOT1_18540 ( P2_R1131_U79 , P2_U3900 );
not NOT1_18541 ( P2_R1131_U80 , P2_U3901 );
not NOT1_18542 ( P2_R1131_U81 , P2_U3902 );
not NOT1_18543 ( P2_R1131_U82 , P2_U3065 );
not NOT1_18544 ( P2_R1131_U83 , P2_U3060 );
not NOT1_18545 ( P2_R1131_U84 , P2_U3074 );
nand NAND2_18546 ( P2_R1131_U85 , P2_U3074 , P2_R1131_U81 );
not NOT1_18547 ( P2_R1131_U86 , P2_U3899 );
not NOT1_18548 ( P2_R1131_U87 , P2_U3064 );
not NOT1_18549 ( P2_R1131_U88 , P2_U3898 );
not NOT1_18550 ( P2_R1131_U89 , P2_U3057 );
not NOT1_18551 ( P2_R1131_U90 , P2_U3897 );
not NOT1_18552 ( P2_R1131_U91 , P2_U3896 );
not NOT1_18553 ( P2_R1131_U92 , P2_U3053 );
nand NAND2_18554 ( P2_R1131_U93 , P2_R1131_U297 , P2_R1131_U296 );
nand NAND2_18555 ( P2_R1131_U94 , P2_R1131_U85 , P2_R1131_U307 );
nand NAND2_18556 ( P2_R1131_U95 , P2_R1131_U71 , P2_R1131_U318 );
nand NAND2_18557 ( P2_R1131_U96 , P2_R1131_U349 , P2_R1131_U59 );
not NOT1_18558 ( P2_R1131_U97 , P2_U3076 );
nand NAND2_18559 ( P2_R1131_U98 , P2_R1131_U406 , P2_R1131_U405 );
nand NAND2_18560 ( P2_R1131_U99 , P2_R1131_U420 , P2_R1131_U419 );
nand NAND2_18561 ( P2_R1131_U100 , P2_R1131_U425 , P2_R1131_U424 );
nand NAND2_18562 ( P2_R1131_U101 , P2_R1131_U441 , P2_R1131_U440 );
nand NAND2_18563 ( P2_R1131_U102 , P2_R1131_U446 , P2_R1131_U445 );
nand NAND2_18564 ( P2_R1131_U103 , P2_R1131_U451 , P2_R1131_U450 );
nand NAND2_18565 ( P2_R1131_U104 , P2_R1131_U456 , P2_R1131_U455 );
nand NAND2_18566 ( P2_R1131_U105 , P2_R1131_U461 , P2_R1131_U460 );
nand NAND2_18567 ( P2_R1131_U106 , P2_R1131_U477 , P2_R1131_U476 );
nand NAND2_18568 ( P2_R1131_U107 , P2_R1131_U482 , P2_R1131_U481 );
nand NAND2_18569 ( P2_R1131_U108 , P2_R1131_U365 , P2_R1131_U364 );
nand NAND2_18570 ( P2_R1131_U109 , P2_R1131_U374 , P2_R1131_U373 );
nand NAND2_18571 ( P2_R1131_U110 , P2_R1131_U381 , P2_R1131_U380 );
nand NAND2_18572 ( P2_R1131_U111 , P2_R1131_U385 , P2_R1131_U384 );
nand NAND2_18573 ( P2_R1131_U112 , P2_R1131_U394 , P2_R1131_U393 );
nand NAND2_18574 ( P2_R1131_U113 , P2_R1131_U415 , P2_R1131_U414 );
nand NAND2_18575 ( P2_R1131_U114 , P2_R1131_U432 , P2_R1131_U431 );
nand NAND2_18576 ( P2_R1131_U115 , P2_R1131_U436 , P2_R1131_U435 );
nand NAND2_18577 ( P2_R1131_U116 , P2_R1131_U468 , P2_R1131_U467 );
nand NAND2_18578 ( P2_R1131_U117 , P2_R1131_U472 , P2_R1131_U471 );
nand NAND2_18579 ( P2_R1131_U118 , P2_R1131_U489 , P2_R1131_U488 );
and AND2_18580 ( P2_R1131_U119 , P2_R1131_U206 , P2_R1131_U196 );
and AND2_18581 ( P2_R1131_U120 , P2_R1131_U209 , P2_R1131_U208 );
and AND2_18582 ( P2_R1131_U121 , P2_R1131_U14 , P2_R1131_U13 );
and AND2_18583 ( P2_R1131_U122 , P2_R1131_U340 , P2_R1131_U222 );
and AND2_18584 ( P2_R1131_U123 , P2_R1131_U342 , P2_R1131_U122 );
and AND3_18585 ( P2_R1131_U124 , P2_R1131_U367 , P2_R1131_U366 , P2_R1131_U27 );
and AND2_18586 ( P2_R1131_U125 , P2_R1131_U370 , P2_R1131_U198 );
and AND2_18587 ( P2_R1131_U126 , P2_R1131_U237 , P2_R1131_U6 );
and AND2_18588 ( P2_R1131_U127 , P2_R1131_U377 , P2_R1131_U197 );
and AND3_18589 ( P2_R1131_U128 , P2_R1131_U387 , P2_R1131_U386 , P2_R1131_U35 );
and AND2_18590 ( P2_R1131_U129 , P2_R1131_U390 , P2_R1131_U196 );
and AND2_18591 ( P2_R1131_U130 , P2_R1131_U251 , P2_R1131_U15 );
and AND2_18592 ( P2_R1131_U131 , P2_R1131_U343 , P2_R1131_U252 );
and AND2_18593 ( P2_R1131_U132 , P2_R1131_U262 , P2_R1131_U8 );
and AND2_18594 ( P2_R1131_U133 , P2_R1131_U286 , P2_R1131_U10 );
and AND2_18595 ( P2_R1131_U134 , P2_R1131_U302 , P2_R1131_U301 );
and AND2_18596 ( P2_R1131_U135 , P2_R1131_U397 , P2_R1131_U303 );
and AND4_18597 ( P2_R1131_U136 , P2_R1131_U302 , P2_R1131_U301 , P2_R1131_U304 , P2_R1131_U16 );
and AND2_18598 ( P2_R1131_U137 , P2_R1131_U359 , P2_R1131_U165 );
nand NAND2_18599 ( P2_R1131_U138 , P2_R1131_U403 , P2_R1131_U402 );
and AND3_18600 ( P2_R1131_U139 , P2_R1131_U408 , P2_R1131_U407 , P2_R1131_U53 );
and AND2_18601 ( P2_R1131_U140 , P2_R1131_U411 , P2_R1131_U195 );
nand NAND2_18602 ( P2_R1131_U141 , P2_R1131_U417 , P2_R1131_U416 );
nand NAND2_18603 ( P2_R1131_U142 , P2_R1131_U422 , P2_R1131_U421 );
and AND2_18604 ( P2_R1131_U143 , P2_R1131_U313 , P2_R1131_U11 );
and AND2_18605 ( P2_R1131_U144 , P2_R1131_U428 , P2_R1131_U194 );
nand NAND2_18606 ( P2_R1131_U145 , P2_R1131_U438 , P2_R1131_U437 );
nand NAND2_18607 ( P2_R1131_U146 , P2_R1131_U443 , P2_R1131_U442 );
nand NAND2_18608 ( P2_R1131_U147 , P2_R1131_U448 , P2_R1131_U447 );
nand NAND2_18609 ( P2_R1131_U148 , P2_R1131_U453 , P2_R1131_U452 );
nand NAND2_18610 ( P2_R1131_U149 , P2_R1131_U458 , P2_R1131_U457 );
and AND2_18611 ( P2_R1131_U150 , P2_R1131_U324 , P2_R1131_U9 );
and AND2_18612 ( P2_R1131_U151 , P2_R1131_U464 , P2_R1131_U193 );
nand NAND2_18613 ( P2_R1131_U152 , P2_R1131_U474 , P2_R1131_U473 );
nand NAND2_18614 ( P2_R1131_U153 , P2_R1131_U479 , P2_R1131_U478 );
and AND2_18615 ( P2_R1131_U154 , P2_R1131_U333 , P2_R1131_U7 );
and AND2_18616 ( P2_R1131_U155 , P2_R1131_U485 , P2_R1131_U192 );
and AND2_18617 ( P2_R1131_U156 , P2_R1131_U363 , P2_R1131_U362 );
nand NAND2_18618 ( P2_R1131_U157 , P2_R1131_U123 , P2_R1131_U341 );
and AND2_18619 ( P2_R1131_U158 , P2_R1131_U372 , P2_R1131_U371 );
and AND2_18620 ( P2_R1131_U159 , P2_R1131_U379 , P2_R1131_U378 );
and AND2_18621 ( P2_R1131_U160 , P2_R1131_U383 , P2_R1131_U382 );
nand NAND2_18622 ( P2_R1131_U161 , P2_R1131_U120 , P2_R1131_U344 );
and AND2_18623 ( P2_R1131_U162 , P2_R1131_U392 , P2_R1131_U391 );
not NOT1_18624 ( P2_R1131_U163 , P2_U3904 );
not NOT1_18625 ( P2_R1131_U164 , P2_U3054 );
and AND2_18626 ( P2_R1131_U165 , P2_R1131_U401 , P2_R1131_U400 );
nand NAND2_18627 ( P2_R1131_U166 , P2_R1131_U134 , P2_R1131_U360 );
and AND2_18628 ( P2_R1131_U167 , P2_R1131_U413 , P2_R1131_U412 );
nand NAND2_18629 ( P2_R1131_U168 , P2_R1131_U293 , P2_R1131_U292 );
nand NAND2_18630 ( P2_R1131_U169 , P2_R1131_U289 , P2_R1131_U288 );
and AND2_18631 ( P2_R1131_U170 , P2_R1131_U430 , P2_R1131_U429 );
and AND2_18632 ( P2_R1131_U171 , P2_R1131_U434 , P2_R1131_U433 );
nand NAND2_18633 ( P2_R1131_U172 , P2_R1131_U279 , P2_R1131_U278 );
nand NAND2_18634 ( P2_R1131_U173 , P2_R1131_U275 , P2_R1131_U274 );
not NOT1_18635 ( P2_R1131_U174 , P2_U3392 );
nand NAND2_18636 ( P2_R1131_U175 , P2_U3387 , P2_R1131_U97 );
nand NAND3_18637 ( P2_R1131_U176 , P2_R1131_U271 , P2_R1131_U187 , P2_R1131_U339 );
not NOT1_18638 ( P2_R1131_U177 , P2_U3443 );
nand NAND2_18639 ( P2_R1131_U178 , P2_R1131_U269 , P2_R1131_U268 );
nand NAND2_18640 ( P2_R1131_U179 , P2_R1131_U265 , P2_R1131_U264 );
and AND2_18641 ( P2_R1131_U180 , P2_R1131_U466 , P2_R1131_U465 );
and AND2_18642 ( P2_R1131_U181 , P2_R1131_U470 , P2_R1131_U469 );
nand NAND2_18643 ( P2_R1131_U182 , P2_R1131_U255 , P2_R1131_U254 );
nand NAND2_18644 ( P2_R1131_U183 , P2_R1131_U131 , P2_R1131_U353 );
nand NAND2_18645 ( P2_R1131_U184 , P2_R1131_U351 , P2_R1131_U62 );
and AND2_18646 ( P2_R1131_U185 , P2_R1131_U487 , P2_R1131_U486 );
nand NAND2_18647 ( P2_R1131_U186 , P2_R1131_U135 , P2_R1131_U166 );
nand NAND2_18648 ( P2_R1131_U187 , P2_R1131_U178 , P2_R1131_U177 );
nand NAND2_18649 ( P2_R1131_U188 , P2_R1131_U175 , P2_R1131_U174 );
not NOT1_18650 ( P2_R1131_U189 , P2_R1131_U53 );
not NOT1_18651 ( P2_R1131_U190 , P2_R1131_U35 );
not NOT1_18652 ( P2_R1131_U191 , P2_R1131_U27 );
nand NAND2_18653 ( P2_R1131_U192 , P2_U3419 , P2_R1131_U57 );
nand NAND2_18654 ( P2_R1131_U193 , P2_U3434 , P2_R1131_U69 );
nand NAND2_18655 ( P2_R1131_U194 , P2_U3901 , P2_R1131_U83 );
nand NAND2_18656 ( P2_R1131_U195 , P2_U3897 , P2_R1131_U52 );
nand NAND2_18657 ( P2_R1131_U196 , P2_U3395 , P2_R1131_U34 );
nand NAND2_18658 ( P2_R1131_U197 , P2_U3404 , P2_R1131_U42 );
nand NAND2_18659 ( P2_R1131_U198 , P2_U3410 , P2_R1131_U26 );
not NOT1_18660 ( P2_R1131_U199 , P2_R1131_U71 );
not NOT1_18661 ( P2_R1131_U200 , P2_R1131_U85 );
not NOT1_18662 ( P2_R1131_U201 , P2_R1131_U44 );
not NOT1_18663 ( P2_R1131_U202 , P2_R1131_U59 );
not NOT1_18664 ( P2_R1131_U203 , P2_R1131_U175 );
nand NAND2_18665 ( P2_R1131_U204 , P2_U3077 , P2_R1131_U175 );
not NOT1_18666 ( P2_R1131_U205 , P2_R1131_U50 );
nand NAND2_18667 ( P2_R1131_U206 , P2_U3398 , P2_R1131_U36 );
nand NAND2_18668 ( P2_R1131_U207 , P2_R1131_U36 , P2_R1131_U35 );
nand NAND2_18669 ( P2_R1131_U208 , P2_R1131_U207 , P2_R1131_U40 );
nand NAND2_18670 ( P2_R1131_U209 , P2_U3063 , P2_R1131_U190 );
nand NAND2_18671 ( P2_R1131_U210 , P2_U3407 , P2_R1131_U41 );
nand NAND2_18672 ( P2_R1131_U211 , P2_U3070 , P2_R1131_U30 );
nand NAND2_18673 ( P2_R1131_U212 , P2_U3066 , P2_R1131_U29 );
nand NAND2_18674 ( P2_R1131_U213 , P2_R1131_U201 , P2_R1131_U197 );
nand NAND2_18675 ( P2_R1131_U214 , P2_R1131_U6 , P2_R1131_U213 );
nand NAND2_18676 ( P2_R1131_U215 , P2_U3401 , P2_R1131_U43 );
nand NAND2_18677 ( P2_R1131_U216 , P2_U3407 , P2_R1131_U41 );
nand NAND2_18678 ( P2_R1131_U217 , P2_R1131_U13 , P2_R1131_U161 );
not NOT1_18679 ( P2_R1131_U218 , P2_R1131_U45 );
not NOT1_18680 ( P2_R1131_U219 , P2_R1131_U48 );
nand NAND2_18681 ( P2_R1131_U220 , P2_U3413 , P2_R1131_U28 );
nand NAND2_18682 ( P2_R1131_U221 , P2_R1131_U28 , P2_R1131_U27 );
nand NAND2_18683 ( P2_R1131_U222 , P2_U3083 , P2_R1131_U191 );
not NOT1_18684 ( P2_R1131_U223 , P2_R1131_U157 );
nand NAND2_18685 ( P2_R1131_U224 , P2_U3416 , P2_R1131_U47 );
nand NAND2_18686 ( P2_R1131_U225 , P2_R1131_U224 , P2_R1131_U59 );
nand NAND2_18687 ( P2_R1131_U226 , P2_R1131_U219 , P2_R1131_U27 );
nand NAND2_18688 ( P2_R1131_U227 , P2_R1131_U125 , P2_R1131_U226 );
nand NAND2_18689 ( P2_R1131_U228 , P2_R1131_U48 , P2_R1131_U198 );
nand NAND2_18690 ( P2_R1131_U229 , P2_R1131_U124 , P2_R1131_U228 );
nand NAND2_18691 ( P2_R1131_U230 , P2_R1131_U27 , P2_R1131_U198 );
nand NAND2_18692 ( P2_R1131_U231 , P2_R1131_U215 , P2_R1131_U161 );
not NOT1_18693 ( P2_R1131_U232 , P2_R1131_U49 );
nand NAND2_18694 ( P2_R1131_U233 , P2_U3066 , P2_R1131_U29 );
nand NAND2_18695 ( P2_R1131_U234 , P2_R1131_U232 , P2_R1131_U233 );
nand NAND2_18696 ( P2_R1131_U235 , P2_R1131_U127 , P2_R1131_U234 );
nand NAND2_18697 ( P2_R1131_U236 , P2_R1131_U49 , P2_R1131_U197 );
nand NAND2_18698 ( P2_R1131_U237 , P2_U3407 , P2_R1131_U41 );
nand NAND2_18699 ( P2_R1131_U238 , P2_R1131_U126 , P2_R1131_U236 );
nand NAND2_18700 ( P2_R1131_U239 , P2_U3066 , P2_R1131_U29 );
nand NAND2_18701 ( P2_R1131_U240 , P2_R1131_U239 , P2_R1131_U197 );
nand NAND2_18702 ( P2_R1131_U241 , P2_R1131_U215 , P2_R1131_U44 );
nand NAND2_18703 ( P2_R1131_U242 , P2_R1131_U129 , P2_R1131_U348 );
nand NAND2_18704 ( P2_R1131_U243 , P2_R1131_U35 , P2_R1131_U196 );
nand NAND2_18705 ( P2_R1131_U244 , P2_U3422 , P2_R1131_U56 );
nand NAND2_18706 ( P2_R1131_U245 , P2_U3062 , P2_R1131_U60 );
nand NAND2_18707 ( P2_R1131_U246 , P2_U3061 , P2_R1131_U58 );
nand NAND2_18708 ( P2_R1131_U247 , P2_R1131_U202 , P2_R1131_U192 );
nand NAND2_18709 ( P2_R1131_U248 , P2_R1131_U7 , P2_R1131_U247 );
nand NAND2_18710 ( P2_R1131_U249 , P2_U3422 , P2_R1131_U56 );
not NOT1_18711 ( P2_R1131_U250 , P2_R1131_U62 );
nand NAND2_18712 ( P2_R1131_U251 , P2_U3425 , P2_R1131_U55 );
nand NAND2_18713 ( P2_R1131_U252 , P2_U3071 , P2_R1131_U61 );
nand NAND2_18714 ( P2_R1131_U253 , P2_U3428 , P2_R1131_U64 );
nand NAND2_18715 ( P2_R1131_U254 , P2_R1131_U253 , P2_R1131_U183 );
nand NAND2_18716 ( P2_R1131_U255 , P2_U3079 , P2_R1131_U63 );
not NOT1_18717 ( P2_R1131_U256 , P2_R1131_U182 );
nand NAND2_18718 ( P2_R1131_U257 , P2_U3437 , P2_R1131_U68 );
nand NAND2_18719 ( P2_R1131_U258 , P2_U3072 , P2_R1131_U65 );
nand NAND2_18720 ( P2_R1131_U259 , P2_U3073 , P2_R1131_U66 );
nand NAND2_18721 ( P2_R1131_U260 , P2_R1131_U199 , P2_R1131_U8 );
nand NAND2_18722 ( P2_R1131_U261 , P2_R1131_U9 , P2_R1131_U260 );
nand NAND2_18723 ( P2_R1131_U262 , P2_U3431 , P2_R1131_U70 );
nand NAND2_18724 ( P2_R1131_U263 , P2_U3437 , P2_R1131_U68 );
nand NAND2_18725 ( P2_R1131_U264 , P2_R1131_U132 , P2_R1131_U182 );
nand NAND2_18726 ( P2_R1131_U265 , P2_R1131_U263 , P2_R1131_U261 );
not NOT1_18727 ( P2_R1131_U266 , P2_R1131_U179 );
nand NAND2_18728 ( P2_R1131_U267 , P2_U3440 , P2_R1131_U73 );
nand NAND2_18729 ( P2_R1131_U268 , P2_R1131_U267 , P2_R1131_U179 );
nand NAND2_18730 ( P2_R1131_U269 , P2_U3068 , P2_R1131_U72 );
not NOT1_18731 ( P2_R1131_U270 , P2_R1131_U178 );
nand NAND2_18732 ( P2_R1131_U271 , P2_U3081 , P2_R1131_U178 );
not NOT1_18733 ( P2_R1131_U272 , P2_R1131_U176 );
nand NAND2_18734 ( P2_R1131_U273 , P2_U3445 , P2_R1131_U76 );
nand NAND2_18735 ( P2_R1131_U274 , P2_R1131_U273 , P2_R1131_U176 );
nand NAND2_18736 ( P2_R1131_U275 , P2_U3080 , P2_R1131_U75 );
not NOT1_18737 ( P2_R1131_U276 , P2_R1131_U173 );
nand NAND2_18738 ( P2_R1131_U277 , P2_U3903 , P2_R1131_U78 );
nand NAND2_18739 ( P2_R1131_U278 , P2_R1131_U277 , P2_R1131_U173 );
nand NAND2_18740 ( P2_R1131_U279 , P2_U3075 , P2_R1131_U77 );
not NOT1_18741 ( P2_R1131_U280 , P2_R1131_U172 );
nand NAND2_18742 ( P2_R1131_U281 , P2_U3900 , P2_R1131_U82 );
nand NAND2_18743 ( P2_R1131_U282 , P2_U3065 , P2_R1131_U79 );
nand NAND2_18744 ( P2_R1131_U283 , P2_U3060 , P2_R1131_U80 );
nand NAND2_18745 ( P2_R1131_U284 , P2_R1131_U200 , P2_R1131_U10 );
nand NAND2_18746 ( P2_R1131_U285 , P2_R1131_U11 , P2_R1131_U284 );
nand NAND2_18747 ( P2_R1131_U286 , P2_U3902 , P2_R1131_U84 );
nand NAND2_18748 ( P2_R1131_U287 , P2_U3900 , P2_R1131_U82 );
nand NAND2_18749 ( P2_R1131_U288 , P2_R1131_U133 , P2_R1131_U172 );
nand NAND2_18750 ( P2_R1131_U289 , P2_R1131_U287 , P2_R1131_U285 );
not NOT1_18751 ( P2_R1131_U290 , P2_R1131_U169 );
nand NAND2_18752 ( P2_R1131_U291 , P2_U3899 , P2_R1131_U87 );
nand NAND2_18753 ( P2_R1131_U292 , P2_R1131_U291 , P2_R1131_U169 );
nand NAND2_18754 ( P2_R1131_U293 , P2_U3064 , P2_R1131_U86 );
not NOT1_18755 ( P2_R1131_U294 , P2_R1131_U168 );
nand NAND2_18756 ( P2_R1131_U295 , P2_U3898 , P2_R1131_U89 );
nand NAND2_18757 ( P2_R1131_U296 , P2_R1131_U295 , P2_R1131_U168 );
nand NAND2_18758 ( P2_R1131_U297 , P2_U3057 , P2_R1131_U88 );
not NOT1_18759 ( P2_R1131_U298 , P2_R1131_U93 );
nand NAND2_18760 ( P2_R1131_U299 , P2_U3896 , P2_R1131_U54 );
nand NAND2_18761 ( P2_R1131_U300 , P2_R1131_U54 , P2_R1131_U53 );
nand NAND2_18762 ( P2_R1131_U301 , P2_R1131_U300 , P2_R1131_U91 );
nand NAND2_18763 ( P2_R1131_U302 , P2_U3052 , P2_R1131_U189 );
nand NAND2_18764 ( P2_R1131_U303 , P2_U3895 , P2_R1131_U92 );
nand NAND2_18765 ( P2_R1131_U304 , P2_U3053 , P2_R1131_U51 );
nand NAND2_18766 ( P2_R1131_U305 , P2_R1131_U140 , P2_R1131_U355 );
nand NAND2_18767 ( P2_R1131_U306 , P2_R1131_U53 , P2_R1131_U195 );
nand NAND2_18768 ( P2_R1131_U307 , P2_R1131_U286 , P2_R1131_U172 );
not NOT1_18769 ( P2_R1131_U308 , P2_R1131_U94 );
nand NAND2_18770 ( P2_R1131_U309 , P2_U3060 , P2_R1131_U80 );
nand NAND2_18771 ( P2_R1131_U310 , P2_R1131_U308 , P2_R1131_U309 );
nand NAND2_18772 ( P2_R1131_U311 , P2_R1131_U144 , P2_R1131_U310 );
nand NAND2_18773 ( P2_R1131_U312 , P2_R1131_U94 , P2_R1131_U194 );
nand NAND2_18774 ( P2_R1131_U313 , P2_U3900 , P2_R1131_U82 );
nand NAND2_18775 ( P2_R1131_U314 , P2_R1131_U143 , P2_R1131_U312 );
nand NAND2_18776 ( P2_R1131_U315 , P2_U3060 , P2_R1131_U80 );
nand NAND2_18777 ( P2_R1131_U316 , P2_R1131_U194 , P2_R1131_U315 );
nand NAND2_18778 ( P2_R1131_U317 , P2_R1131_U286 , P2_R1131_U85 );
nand NAND2_18779 ( P2_R1131_U318 , P2_R1131_U262 , P2_R1131_U182 );
not NOT1_18780 ( P2_R1131_U319 , P2_R1131_U95 );
nand NAND2_18781 ( P2_R1131_U320 , P2_U3073 , P2_R1131_U66 );
nand NAND2_18782 ( P2_R1131_U321 , P2_R1131_U319 , P2_R1131_U320 );
nand NAND2_18783 ( P2_R1131_U322 , P2_R1131_U151 , P2_R1131_U321 );
nand NAND2_18784 ( P2_R1131_U323 , P2_R1131_U95 , P2_R1131_U193 );
nand NAND2_18785 ( P2_R1131_U324 , P2_U3437 , P2_R1131_U68 );
nand NAND2_18786 ( P2_R1131_U325 , P2_R1131_U150 , P2_R1131_U323 );
nand NAND2_18787 ( P2_R1131_U326 , P2_U3073 , P2_R1131_U66 );
nand NAND2_18788 ( P2_R1131_U327 , P2_R1131_U193 , P2_R1131_U326 );
nand NAND2_18789 ( P2_R1131_U328 , P2_R1131_U262 , P2_R1131_U71 );
nand NAND2_18790 ( P2_R1131_U329 , P2_U3061 , P2_R1131_U58 );
nand NAND2_18791 ( P2_R1131_U330 , P2_R1131_U350 , P2_R1131_U329 );
nand NAND2_18792 ( P2_R1131_U331 , P2_R1131_U155 , P2_R1131_U330 );
nand NAND2_18793 ( P2_R1131_U332 , P2_R1131_U96 , P2_R1131_U192 );
nand NAND2_18794 ( P2_R1131_U333 , P2_U3422 , P2_R1131_U56 );
nand NAND2_18795 ( P2_R1131_U334 , P2_R1131_U154 , P2_R1131_U332 );
nand NAND2_18796 ( P2_R1131_U335 , P2_U3061 , P2_R1131_U58 );
nand NAND2_18797 ( P2_R1131_U336 , P2_R1131_U192 , P2_R1131_U335 );
nand NAND2_18798 ( P2_R1131_U337 , P2_U3076 , P2_R1131_U38 );
nand NAND2_18799 ( P2_R1131_U338 , P2_U3077 , P2_R1131_U174 );
nand NAND2_18800 ( P2_R1131_U339 , P2_U3081 , P2_R1131_U177 );
nand NAND2_18801 ( P2_R1131_U340 , P2_R1131_U33 , P2_R1131_U221 );
nand NAND2_18802 ( P2_R1131_U341 , P2_R1131_U121 , P2_R1131_U161 );
nand NAND2_18803 ( P2_R1131_U342 , P2_R1131_U218 , P2_R1131_U14 );
nand NAND2_18804 ( P2_R1131_U343 , P2_R1131_U250 , P2_R1131_U251 );
nand NAND2_18805 ( P2_R1131_U344 , P2_R1131_U119 , P2_R1131_U50 );
not NOT1_18806 ( P2_R1131_U345 , P2_R1131_U161 );
nand NAND2_18807 ( P2_R1131_U346 , P2_R1131_U196 , P2_R1131_U50 );
nand NAND2_18808 ( P2_R1131_U347 , P2_R1131_U128 , P2_R1131_U346 );
nand NAND2_18809 ( P2_R1131_U348 , P2_R1131_U205 , P2_R1131_U35 );
nand NAND2_18810 ( P2_R1131_U349 , P2_R1131_U224 , P2_R1131_U157 );
not NOT1_18811 ( P2_R1131_U350 , P2_R1131_U96 );
nand NAND2_18812 ( P2_R1131_U351 , P2_R1131_U15 , P2_R1131_U157 );
not NOT1_18813 ( P2_R1131_U352 , P2_R1131_U184 );
nand NAND2_18814 ( P2_R1131_U353 , P2_R1131_U130 , P2_R1131_U157 );
not NOT1_18815 ( P2_R1131_U354 , P2_R1131_U183 );
nand NAND2_18816 ( P2_R1131_U355 , P2_R1131_U298 , P2_R1131_U53 );
nand NAND2_18817 ( P2_R1131_U356 , P2_R1131_U195 , P2_R1131_U93 );
nand NAND2_18818 ( P2_R1131_U357 , P2_R1131_U139 , P2_R1131_U356 );
nand NAND2_18819 ( P2_R1131_U358 , P2_R1131_U12 , P2_R1131_U93 );
nand NAND2_18820 ( P2_R1131_U359 , P2_R1131_U136 , P2_R1131_U358 );
nand NAND2_18821 ( P2_R1131_U360 , P2_R1131_U12 , P2_R1131_U93 );
not NOT1_18822 ( P2_R1131_U361 , P2_R1131_U166 );
nand NAND2_18823 ( P2_R1131_U362 , P2_U3416 , P2_R1131_U47 );
nand NAND2_18824 ( P2_R1131_U363 , P2_U3082 , P2_R1131_U46 );
nand NAND2_18825 ( P2_R1131_U364 , P2_R1131_U225 , P2_R1131_U157 );
nand NAND2_18826 ( P2_R1131_U365 , P2_R1131_U223 , P2_R1131_U156 );
nand NAND2_18827 ( P2_R1131_U366 , P2_U3413 , P2_R1131_U28 );
nand NAND2_18828 ( P2_R1131_U367 , P2_U3083 , P2_R1131_U33 );
nand NAND2_18829 ( P2_R1131_U368 , P2_U3413 , P2_R1131_U28 );
nand NAND2_18830 ( P2_R1131_U369 , P2_U3083 , P2_R1131_U33 );
nand NAND2_18831 ( P2_R1131_U370 , P2_R1131_U369 , P2_R1131_U368 );
nand NAND2_18832 ( P2_R1131_U371 , P2_U3410 , P2_R1131_U26 );
nand NAND2_18833 ( P2_R1131_U372 , P2_U3069 , P2_R1131_U32 );
nand NAND2_18834 ( P2_R1131_U373 , P2_R1131_U230 , P2_R1131_U48 );
nand NAND2_18835 ( P2_R1131_U374 , P2_R1131_U158 , P2_R1131_U219 );
nand NAND2_18836 ( P2_R1131_U375 , P2_U3407 , P2_R1131_U41 );
nand NAND2_18837 ( P2_R1131_U376 , P2_U3070 , P2_R1131_U30 );
nand NAND2_18838 ( P2_R1131_U377 , P2_R1131_U376 , P2_R1131_U375 );
nand NAND2_18839 ( P2_R1131_U378 , P2_U3404 , P2_R1131_U42 );
nand NAND2_18840 ( P2_R1131_U379 , P2_U3066 , P2_R1131_U29 );
nand NAND2_18841 ( P2_R1131_U380 , P2_R1131_U240 , P2_R1131_U49 );
nand NAND2_18842 ( P2_R1131_U381 , P2_R1131_U159 , P2_R1131_U232 );
nand NAND2_18843 ( P2_R1131_U382 , P2_U3401 , P2_R1131_U43 );
nand NAND2_18844 ( P2_R1131_U383 , P2_U3059 , P2_R1131_U31 );
nand NAND2_18845 ( P2_R1131_U384 , P2_R1131_U161 , P2_R1131_U241 );
nand NAND2_18846 ( P2_R1131_U385 , P2_R1131_U345 , P2_R1131_U160 );
nand NAND2_18847 ( P2_R1131_U386 , P2_U3398 , P2_R1131_U36 );
nand NAND2_18848 ( P2_R1131_U387 , P2_U3063 , P2_R1131_U40 );
nand NAND2_18849 ( P2_R1131_U388 , P2_U3398 , P2_R1131_U36 );
nand NAND2_18850 ( P2_R1131_U389 , P2_U3063 , P2_R1131_U40 );
nand NAND2_18851 ( P2_R1131_U390 , P2_R1131_U389 , P2_R1131_U388 );
nand NAND2_18852 ( P2_R1131_U391 , P2_U3395 , P2_R1131_U34 );
nand NAND2_18853 ( P2_R1131_U392 , P2_U3067 , P2_R1131_U37 );
nand NAND2_18854 ( P2_R1131_U393 , P2_R1131_U243 , P2_R1131_U50 );
nand NAND2_18855 ( P2_R1131_U394 , P2_R1131_U162 , P2_R1131_U205 );
nand NAND2_18856 ( P2_R1131_U395 , P2_U3904 , P2_R1131_U164 );
nand NAND2_18857 ( P2_R1131_U396 , P2_U3054 , P2_R1131_U163 );
nand NAND2_18858 ( P2_R1131_U397 , P2_R1131_U396 , P2_R1131_U395 );
nand NAND2_18859 ( P2_R1131_U398 , P2_U3904 , P2_R1131_U164 );
nand NAND2_18860 ( P2_R1131_U399 , P2_U3054 , P2_R1131_U163 );
nand NAND3_18861 ( P2_R1131_U400 , P2_U3053 , P2_R1131_U397 , P2_R1131_U51 );
nand NAND3_18862 ( P2_R1131_U401 , P2_R1131_U16 , P2_R1131_U92 , P2_U3895 );
nand NAND2_18863 ( P2_R1131_U402 , P2_U3895 , P2_R1131_U92 );
nand NAND2_18864 ( P2_R1131_U403 , P2_U3053 , P2_R1131_U51 );
not NOT1_18865 ( P2_R1131_U404 , P2_R1131_U138 );
nand NAND2_18866 ( P2_R1131_U405 , P2_R1131_U361 , P2_R1131_U404 );
nand NAND2_18867 ( P2_R1131_U406 , P2_R1131_U138 , P2_R1131_U166 );
nand NAND2_18868 ( P2_R1131_U407 , P2_U3896 , P2_R1131_U54 );
nand NAND2_18869 ( P2_R1131_U408 , P2_U3052 , P2_R1131_U91 );
nand NAND2_18870 ( P2_R1131_U409 , P2_U3896 , P2_R1131_U54 );
nand NAND2_18871 ( P2_R1131_U410 , P2_U3052 , P2_R1131_U91 );
nand NAND2_18872 ( P2_R1131_U411 , P2_R1131_U410 , P2_R1131_U409 );
nand NAND2_18873 ( P2_R1131_U412 , P2_U3897 , P2_R1131_U52 );
nand NAND2_18874 ( P2_R1131_U413 , P2_U3056 , P2_R1131_U90 );
nand NAND2_18875 ( P2_R1131_U414 , P2_R1131_U306 , P2_R1131_U93 );
nand NAND2_18876 ( P2_R1131_U415 , P2_R1131_U167 , P2_R1131_U298 );
nand NAND2_18877 ( P2_R1131_U416 , P2_U3898 , P2_R1131_U89 );
nand NAND2_18878 ( P2_R1131_U417 , P2_U3057 , P2_R1131_U88 );
not NOT1_18879 ( P2_R1131_U418 , P2_R1131_U141 );
nand NAND2_18880 ( P2_R1131_U419 , P2_R1131_U294 , P2_R1131_U418 );
nand NAND2_18881 ( P2_R1131_U420 , P2_R1131_U141 , P2_R1131_U168 );
nand NAND2_18882 ( P2_R1131_U421 , P2_U3899 , P2_R1131_U87 );
nand NAND2_18883 ( P2_R1131_U422 , P2_U3064 , P2_R1131_U86 );
not NOT1_18884 ( P2_R1131_U423 , P2_R1131_U142 );
nand NAND2_18885 ( P2_R1131_U424 , P2_R1131_U290 , P2_R1131_U423 );
nand NAND2_18886 ( P2_R1131_U425 , P2_R1131_U142 , P2_R1131_U169 );
nand NAND2_18887 ( P2_R1131_U426 , P2_U3900 , P2_R1131_U82 );
nand NAND2_18888 ( P2_R1131_U427 , P2_U3065 , P2_R1131_U79 );
nand NAND2_18889 ( P2_R1131_U428 , P2_R1131_U427 , P2_R1131_U426 );
nand NAND2_18890 ( P2_R1131_U429 , P2_U3901 , P2_R1131_U83 );
nand NAND2_18891 ( P2_R1131_U430 , P2_U3060 , P2_R1131_U80 );
nand NAND2_18892 ( P2_R1131_U431 , P2_R1131_U316 , P2_R1131_U94 );
nand NAND2_18893 ( P2_R1131_U432 , P2_R1131_U170 , P2_R1131_U308 );
nand NAND2_18894 ( P2_R1131_U433 , P2_U3902 , P2_R1131_U84 );
nand NAND2_18895 ( P2_R1131_U434 , P2_U3074 , P2_R1131_U81 );
nand NAND2_18896 ( P2_R1131_U435 , P2_R1131_U317 , P2_R1131_U172 );
nand NAND2_18897 ( P2_R1131_U436 , P2_R1131_U280 , P2_R1131_U171 );
nand NAND2_18898 ( P2_R1131_U437 , P2_U3903 , P2_R1131_U78 );
nand NAND2_18899 ( P2_R1131_U438 , P2_U3075 , P2_R1131_U77 );
not NOT1_18900 ( P2_R1131_U439 , P2_R1131_U145 );
nand NAND2_18901 ( P2_R1131_U440 , P2_R1131_U276 , P2_R1131_U439 );
nand NAND2_18902 ( P2_R1131_U441 , P2_R1131_U145 , P2_R1131_U173 );
nand NAND2_18903 ( P2_R1131_U442 , P2_U3392 , P2_R1131_U39 );
nand NAND2_18904 ( P2_R1131_U443 , P2_U3077 , P2_R1131_U174 );
not NOT1_18905 ( P2_R1131_U444 , P2_R1131_U146 );
nand NAND2_18906 ( P2_R1131_U445 , P2_R1131_U203 , P2_R1131_U444 );
nand NAND2_18907 ( P2_R1131_U446 , P2_R1131_U146 , P2_R1131_U175 );
nand NAND2_18908 ( P2_R1131_U447 , P2_U3445 , P2_R1131_U76 );
nand NAND2_18909 ( P2_R1131_U448 , P2_U3080 , P2_R1131_U75 );
not NOT1_18910 ( P2_R1131_U449 , P2_R1131_U147 );
nand NAND2_18911 ( P2_R1131_U450 , P2_R1131_U272 , P2_R1131_U449 );
nand NAND2_18912 ( P2_R1131_U451 , P2_R1131_U147 , P2_R1131_U176 );
nand NAND2_18913 ( P2_R1131_U452 , P2_U3443 , P2_R1131_U74 );
nand NAND2_18914 ( P2_R1131_U453 , P2_U3081 , P2_R1131_U177 );
not NOT1_18915 ( P2_R1131_U454 , P2_R1131_U148 );
nand NAND2_18916 ( P2_R1131_U455 , P2_R1131_U270 , P2_R1131_U454 );
nand NAND2_18917 ( P2_R1131_U456 , P2_R1131_U148 , P2_R1131_U178 );
nand NAND2_18918 ( P2_R1131_U457 , P2_U3440 , P2_R1131_U73 );
nand NAND2_18919 ( P2_R1131_U458 , P2_U3068 , P2_R1131_U72 );
not NOT1_18920 ( P2_R1131_U459 , P2_R1131_U149 );
nand NAND2_18921 ( P2_R1131_U460 , P2_R1131_U266 , P2_R1131_U459 );
nand NAND2_18922 ( P2_R1131_U461 , P2_R1131_U149 , P2_R1131_U179 );
nand NAND2_18923 ( P2_R1131_U462 , P2_U3437 , P2_R1131_U68 );
nand NAND2_18924 ( P2_R1131_U463 , P2_U3072 , P2_R1131_U65 );
nand NAND2_18925 ( P2_R1131_U464 , P2_R1131_U463 , P2_R1131_U462 );
nand NAND2_18926 ( P2_R1131_U465 , P2_U3434 , P2_R1131_U69 );
nand NAND2_18927 ( P2_R1131_U466 , P2_U3073 , P2_R1131_U66 );
nand NAND2_18928 ( P2_R1131_U467 , P2_R1131_U327 , P2_R1131_U95 );
nand NAND2_18929 ( P2_R1131_U468 , P2_R1131_U180 , P2_R1131_U319 );
nand NAND2_18930 ( P2_R1131_U469 , P2_U3431 , P2_R1131_U70 );
nand NAND2_18931 ( P2_R1131_U470 , P2_U3078 , P2_R1131_U67 );
nand NAND2_18932 ( P2_R1131_U471 , P2_R1131_U328 , P2_R1131_U182 );
nand NAND2_18933 ( P2_R1131_U472 , P2_R1131_U256 , P2_R1131_U181 );
nand NAND2_18934 ( P2_R1131_U473 , P2_U3428 , P2_R1131_U64 );
nand NAND2_18935 ( P2_R1131_U474 , P2_U3079 , P2_R1131_U63 );
not NOT1_18936 ( P2_R1131_U475 , P2_R1131_U152 );
nand NAND2_18937 ( P2_R1131_U476 , P2_R1131_U354 , P2_R1131_U475 );
nand NAND2_18938 ( P2_R1131_U477 , P2_R1131_U152 , P2_R1131_U183 );
nand NAND2_18939 ( P2_R1131_U478 , P2_U3425 , P2_R1131_U55 );
nand NAND2_18940 ( P2_R1131_U479 , P2_U3071 , P2_R1131_U61 );
not NOT1_18941 ( P2_R1131_U480 , P2_R1131_U153 );
nand NAND2_18942 ( P2_R1131_U481 , P2_R1131_U352 , P2_R1131_U480 );
nand NAND2_18943 ( P2_R1131_U482 , P2_R1131_U153 , P2_R1131_U184 );
nand NAND2_18944 ( P2_R1131_U483 , P2_U3422 , P2_R1131_U56 );
nand NAND2_18945 ( P2_R1131_U484 , P2_U3062 , P2_R1131_U60 );
nand NAND2_18946 ( P2_R1131_U485 , P2_R1131_U484 , P2_R1131_U483 );
nand NAND2_18947 ( P2_R1131_U486 , P2_U3419 , P2_R1131_U57 );
nand NAND2_18948 ( P2_R1131_U487 , P2_U3061 , P2_R1131_U58 );
nand NAND2_18949 ( P2_R1131_U488 , P2_R1131_U96 , P2_R1131_U336 );
nand NAND2_18950 ( P2_R1131_U489 , P2_R1131_U185 , P2_R1131_U350 );
and AND2_18951 ( P2_R1054_U6 , P2_R1054_U102 , P2_R1054_U118 );
and AND2_18952 ( P2_R1054_U7 , P2_R1054_U120 , P2_R1054_U119 );
and AND2_18953 ( P2_R1054_U8 , P2_R1054_U99 , P2_R1054_U157 );
and AND2_18954 ( P2_R1054_U9 , P2_R1054_U159 , P2_R1054_U158 );
and AND2_18955 ( P2_R1054_U10 , P2_R1054_U100 , P2_R1054_U174 );
and AND2_18956 ( P2_R1054_U11 , P2_R1054_U176 , P2_R1054_U175 );
nand NAND2_18957 ( P2_R1054_U12 , P2_R1054_U207 , P2_R1054_U210 );
nand NAND2_18958 ( P2_R1054_U13 , P2_R1054_U196 , P2_R1054_U199 );
nand NAND2_18959 ( P2_R1054_U14 , P2_R1054_U153 , P2_R1054_U155 );
nand NAND2_18960 ( P2_R1054_U15 , P2_R1054_U145 , P2_R1054_U148 );
nand NAND2_18961 ( P2_R1054_U16 , P2_R1054_U137 , P2_R1054_U139 );
nand NAND2_18962 ( P2_R1054_U17 , P2_R1054_U21 , P2_R1054_U213 );
not NOT1_18963 ( P2_R1054_U18 , P2_U3409 );
not NOT1_18964 ( P2_R1054_U19 , P2_U3394 );
not NOT1_18965 ( P2_R1054_U20 , P2_U3386 );
nand NAND2_18966 ( P2_R1054_U21 , P2_U3386 , P2_R1054_U65 );
not NOT1_18967 ( P2_R1054_U22 , P2_U3573 );
not NOT1_18968 ( P2_R1054_U23 , P2_U3397 );
not NOT1_18969 ( P2_R1054_U24 , P2_U3562 );
nand NAND2_18970 ( P2_R1054_U25 , P2_U3562 , P2_R1054_U19 );
not NOT1_18971 ( P2_R1054_U26 , P2_U3561 );
not NOT1_18972 ( P2_R1054_U27 , P2_U3406 );
not NOT1_18973 ( P2_R1054_U28 , P2_U3403 );
not NOT1_18974 ( P2_R1054_U29 , P2_U3400 );
not NOT1_18975 ( P2_R1054_U30 , P2_U3558 );
not NOT1_18976 ( P2_R1054_U31 , P2_U3559 );
not NOT1_18977 ( P2_R1054_U32 , P2_U3560 );
nand NAND2_18978 ( P2_R1054_U33 , P2_U3560 , P2_R1054_U29 );
not NOT1_18979 ( P2_R1054_U34 , P2_U3412 );
not NOT1_18980 ( P2_R1054_U35 , P2_U3557 );
nand NAND2_18981 ( P2_R1054_U36 , P2_U3557 , P2_R1054_U18 );
not NOT1_18982 ( P2_R1054_U37 , P2_U3556 );
not NOT1_18983 ( P2_R1054_U38 , P2_U3415 );
not NOT1_18984 ( P2_R1054_U39 , P2_U3555 );
nand NAND2_18985 ( P2_R1054_U40 , P2_R1054_U126 , P2_R1054_U125 );
nand NAND2_18986 ( P2_R1054_U41 , P2_R1054_U33 , P2_R1054_U141 );
nand NAND2_18987 ( P2_R1054_U42 , P2_R1054_U110 , P2_R1054_U109 );
not NOT1_18988 ( P2_R1054_U43 , P2_U3421 );
not NOT1_18989 ( P2_R1054_U44 , P2_U3418 );
not NOT1_18990 ( P2_R1054_U45 , P2_U3571 );
not NOT1_18991 ( P2_R1054_U46 , P2_U3572 );
nand NAND2_18992 ( P2_R1054_U47 , P2_U3555 , P2_R1054_U38 );
not NOT1_18993 ( P2_R1054_U48 , P2_U3424 );
not NOT1_18994 ( P2_R1054_U49 , P2_U3570 );
not NOT1_18995 ( P2_R1054_U50 , P2_U3427 );
not NOT1_18996 ( P2_R1054_U51 , P2_U3569 );
not NOT1_18997 ( P2_R1054_U52 , P2_U3436 );
not NOT1_18998 ( P2_R1054_U53 , P2_U3433 );
not NOT1_18999 ( P2_R1054_U54 , P2_U3430 );
not NOT1_19000 ( P2_R1054_U55 , P2_U3566 );
not NOT1_19001 ( P2_R1054_U56 , P2_U3567 );
not NOT1_19002 ( P2_R1054_U57 , P2_U3568 );
nand NAND2_19003 ( P2_R1054_U58 , P2_U3568 , P2_R1054_U54 );
not NOT1_19004 ( P2_R1054_U59 , P2_U3439 );
not NOT1_19005 ( P2_R1054_U60 , P2_U3565 );
nand NAND2_19006 ( P2_R1054_U61 , P2_R1054_U186 , P2_R1054_U185 );
not NOT1_19007 ( P2_R1054_U62 , P2_U3564 );
nand NAND2_19008 ( P2_R1054_U63 , P2_R1054_U58 , P2_R1054_U192 );
nand NAND2_19009 ( P2_R1054_U64 , P2_R1054_U47 , P2_R1054_U203 );
not NOT1_19010 ( P2_R1054_U65 , P2_U3574 );
nand NAND2_19011 ( P2_R1054_U66 , P2_R1054_U251 , P2_R1054_U250 );
nand NAND2_19012 ( P2_R1054_U67 , P2_R1054_U256 , P2_R1054_U255 );
nand NAND2_19013 ( P2_R1054_U68 , P2_R1054_U261 , P2_R1054_U260 );
nand NAND2_19014 ( P2_R1054_U69 , P2_R1054_U266 , P2_R1054_U265 );
nand NAND2_19015 ( P2_R1054_U70 , P2_R1054_U282 , P2_R1054_U281 );
nand NAND2_19016 ( P2_R1054_U71 , P2_R1054_U287 , P2_R1054_U286 );
nand NAND2_19017 ( P2_R1054_U72 , P2_R1054_U217 , P2_R1054_U216 );
nand NAND2_19018 ( P2_R1054_U73 , P2_R1054_U226 , P2_R1054_U225 );
nand NAND2_19019 ( P2_R1054_U74 , P2_R1054_U233 , P2_R1054_U232 );
nand NAND2_19020 ( P2_R1054_U75 , P2_R1054_U237 , P2_R1054_U236 );
nand NAND2_19021 ( P2_R1054_U76 , P2_R1054_U246 , P2_R1054_U245 );
nand NAND2_19022 ( P2_R1054_U77 , P2_R1054_U273 , P2_R1054_U272 );
nand NAND2_19023 ( P2_R1054_U78 , P2_R1054_U277 , P2_R1054_U276 );
nand NAND2_19024 ( P2_R1054_U79 , P2_R1054_U294 , P2_R1054_U293 );
nand NAND2_19025 ( P2_R1054_U80 , P2_R1054_U248 , P2_R1054_U247 );
nand NAND2_19026 ( P2_R1054_U81 , P2_R1054_U253 , P2_R1054_U252 );
nand NAND2_19027 ( P2_R1054_U82 , P2_R1054_U258 , P2_R1054_U257 );
nand NAND2_19028 ( P2_R1054_U83 , P2_R1054_U263 , P2_R1054_U262 );
nand NAND2_19029 ( P2_R1054_U84 , P2_R1054_U279 , P2_R1054_U278 );
nand NAND2_19030 ( P2_R1054_U85 , P2_R1054_U284 , P2_R1054_U283 );
nand NAND3_19031 ( P2_R1054_U86 , P2_R1054_U131 , P2_R1054_U132 , P2_R1054_U129 );
nand NAND3_19032 ( P2_R1054_U87 , P2_R1054_U115 , P2_R1054_U116 , P2_R1054_U113 );
not NOT1_19033 ( P2_R1054_U88 , P2_U3391 );
not NOT1_19034 ( P2_R1054_U89 , P2_U3379 );
not NOT1_19035 ( P2_R1054_U90 , P2_U3563 );
nand NAND2_19036 ( P2_R1054_U91 , P2_R1054_U190 , P2_R1054_U189 );
not NOT1_19037 ( P2_R1054_U92 , P2_U3442 );
nand NAND2_19038 ( P2_R1054_U93 , P2_R1054_U182 , P2_R1054_U181 );
nand NAND2_19039 ( P2_R1054_U94 , P2_R1054_U172 , P2_R1054_U171 );
nand NAND2_19040 ( P2_R1054_U95 , P2_R1054_U168 , P2_R1054_U167 );
nand NAND2_19041 ( P2_R1054_U96 , P2_R1054_U164 , P2_R1054_U163 );
not NOT1_19042 ( P2_R1054_U97 , P2_R1054_U25 );
not NOT1_19043 ( P2_R1054_U98 , P2_R1054_U36 );
nand NAND2_19044 ( P2_R1054_U99 , P2_U3418 , P2_R1054_U46 );
nand NAND2_19045 ( P2_R1054_U100 , P2_U3433 , P2_R1054_U56 );
nand NAND2_19046 ( P2_R1054_U101 , P2_U3394 , P2_R1054_U24 );
nand NAND2_19047 ( P2_R1054_U102 , P2_U3403 , P2_R1054_U31 );
nand NAND2_19048 ( P2_R1054_U103 , P2_U3409 , P2_R1054_U35 );
not NOT1_19049 ( P2_R1054_U104 , P2_R1054_U58 );
not NOT1_19050 ( P2_R1054_U105 , P2_R1054_U33 );
not NOT1_19051 ( P2_R1054_U106 , P2_R1054_U47 );
not NOT1_19052 ( P2_R1054_U107 , P2_R1054_U21 );
nand NAND2_19053 ( P2_R1054_U108 , P2_R1054_U107 , P2_R1054_U22 );
nand NAND2_19054 ( P2_R1054_U109 , P2_R1054_U108 , P2_R1054_U88 );
nand NAND2_19055 ( P2_R1054_U110 , P2_U3573 , P2_R1054_U21 );
not NOT1_19056 ( P2_R1054_U111 , P2_R1054_U42 );
nand NAND2_19057 ( P2_R1054_U112 , P2_U3397 , P2_R1054_U26 );
nand NAND3_19058 ( P2_R1054_U113 , P2_R1054_U112 , P2_R1054_U101 , P2_R1054_U42 );
nand NAND2_19059 ( P2_R1054_U114 , P2_R1054_U26 , P2_R1054_U25 );
nand NAND2_19060 ( P2_R1054_U115 , P2_R1054_U114 , P2_R1054_U23 );
nand NAND2_19061 ( P2_R1054_U116 , P2_U3561 , P2_R1054_U97 );
not NOT1_19062 ( P2_R1054_U117 , P2_R1054_U87 );
nand NAND2_19063 ( P2_R1054_U118 , P2_U3406 , P2_R1054_U30 );
nand NAND2_19064 ( P2_R1054_U119 , P2_U3558 , P2_R1054_U27 );
nand NAND2_19065 ( P2_R1054_U120 , P2_U3559 , P2_R1054_U28 );
nand NAND2_19066 ( P2_R1054_U121 , P2_R1054_U105 , P2_R1054_U6 );
nand NAND2_19067 ( P2_R1054_U122 , P2_R1054_U7 , P2_R1054_U121 );
nand NAND2_19068 ( P2_R1054_U123 , P2_U3400 , P2_R1054_U32 );
nand NAND2_19069 ( P2_R1054_U124 , P2_U3406 , P2_R1054_U30 );
nand NAND3_19070 ( P2_R1054_U125 , P2_R1054_U123 , P2_R1054_U6 , P2_R1054_U87 );
nand NAND2_19071 ( P2_R1054_U126 , P2_R1054_U124 , P2_R1054_U122 );
not NOT1_19072 ( P2_R1054_U127 , P2_R1054_U40 );
nand NAND2_19073 ( P2_R1054_U128 , P2_U3412 , P2_R1054_U37 );
nand NAND3_19074 ( P2_R1054_U129 , P2_R1054_U128 , P2_R1054_U103 , P2_R1054_U40 );
nand NAND2_19075 ( P2_R1054_U130 , P2_R1054_U37 , P2_R1054_U36 );
nand NAND2_19076 ( P2_R1054_U131 , P2_R1054_U130 , P2_R1054_U34 );
nand NAND2_19077 ( P2_R1054_U132 , P2_U3556 , P2_R1054_U98 );
not NOT1_19078 ( P2_R1054_U133 , P2_R1054_U86 );
nand NAND2_19079 ( P2_R1054_U134 , P2_U3415 , P2_R1054_U39 );
nand NAND2_19080 ( P2_R1054_U135 , P2_R1054_U134 , P2_R1054_U47 );
nand NAND2_19081 ( P2_R1054_U136 , P2_R1054_U127 , P2_R1054_U36 );
nand NAND3_19082 ( P2_R1054_U137 , P2_R1054_U222 , P2_R1054_U103 , P2_R1054_U136 );
nand NAND2_19083 ( P2_R1054_U138 , P2_R1054_U40 , P2_R1054_U103 );
nand NAND4_19084 ( P2_R1054_U139 , P2_R1054_U219 , P2_R1054_U218 , P2_R1054_U36 , P2_R1054_U138 );
nand NAND2_19085 ( P2_R1054_U140 , P2_R1054_U36 , P2_R1054_U103 );
nand NAND2_19086 ( P2_R1054_U141 , P2_R1054_U123 , P2_R1054_U87 );
not NOT1_19087 ( P2_R1054_U142 , P2_R1054_U41 );
nand NAND2_19088 ( P2_R1054_U143 , P2_U3559 , P2_R1054_U28 );
nand NAND2_19089 ( P2_R1054_U144 , P2_R1054_U142 , P2_R1054_U143 );
nand NAND3_19090 ( P2_R1054_U145 , P2_R1054_U229 , P2_R1054_U102 , P2_R1054_U144 );
nand NAND2_19091 ( P2_R1054_U146 , P2_R1054_U41 , P2_R1054_U102 );
nand NAND2_19092 ( P2_R1054_U147 , P2_U3406 , P2_R1054_U30 );
nand NAND3_19093 ( P2_R1054_U148 , P2_R1054_U147 , P2_R1054_U7 , P2_R1054_U146 );
nand NAND2_19094 ( P2_R1054_U149 , P2_U3559 , P2_R1054_U28 );
nand NAND2_19095 ( P2_R1054_U150 , P2_R1054_U102 , P2_R1054_U149 );
nand NAND2_19096 ( P2_R1054_U151 , P2_R1054_U123 , P2_R1054_U33 );
nand NAND2_19097 ( P2_R1054_U152 , P2_R1054_U111 , P2_R1054_U25 );
nand NAND3_19098 ( P2_R1054_U153 , P2_R1054_U242 , P2_R1054_U101 , P2_R1054_U152 );
nand NAND2_19099 ( P2_R1054_U154 , P2_R1054_U42 , P2_R1054_U101 );
nand NAND4_19100 ( P2_R1054_U155 , P2_R1054_U239 , P2_R1054_U238 , P2_R1054_U25 , P2_R1054_U154 );
nand NAND2_19101 ( P2_R1054_U156 , P2_R1054_U25 , P2_R1054_U101 );
nand NAND2_19102 ( P2_R1054_U157 , P2_U3421 , P2_R1054_U45 );
nand NAND2_19103 ( P2_R1054_U158 , P2_U3571 , P2_R1054_U43 );
nand NAND2_19104 ( P2_R1054_U159 , P2_U3572 , P2_R1054_U44 );
nand NAND2_19105 ( P2_R1054_U160 , P2_R1054_U106 , P2_R1054_U8 );
nand NAND2_19106 ( P2_R1054_U161 , P2_R1054_U9 , P2_R1054_U160 );
nand NAND2_19107 ( P2_R1054_U162 , P2_U3421 , P2_R1054_U45 );
nand NAND3_19108 ( P2_R1054_U163 , P2_R1054_U134 , P2_R1054_U8 , P2_R1054_U86 );
nand NAND2_19109 ( P2_R1054_U164 , P2_R1054_U162 , P2_R1054_U161 );
not NOT1_19110 ( P2_R1054_U165 , P2_R1054_U96 );
nand NAND2_19111 ( P2_R1054_U166 , P2_U3424 , P2_R1054_U49 );
nand NAND2_19112 ( P2_R1054_U167 , P2_R1054_U166 , P2_R1054_U96 );
nand NAND2_19113 ( P2_R1054_U168 , P2_U3570 , P2_R1054_U48 );
not NOT1_19114 ( P2_R1054_U169 , P2_R1054_U95 );
nand NAND2_19115 ( P2_R1054_U170 , P2_U3427 , P2_R1054_U51 );
nand NAND2_19116 ( P2_R1054_U171 , P2_R1054_U170 , P2_R1054_U95 );
nand NAND2_19117 ( P2_R1054_U172 , P2_U3569 , P2_R1054_U50 );
not NOT1_19118 ( P2_R1054_U173 , P2_R1054_U94 );
nand NAND2_19119 ( P2_R1054_U174 , P2_U3436 , P2_R1054_U55 );
nand NAND2_19120 ( P2_R1054_U175 , P2_U3566 , P2_R1054_U52 );
nand NAND2_19121 ( P2_R1054_U176 , P2_U3567 , P2_R1054_U53 );
nand NAND2_19122 ( P2_R1054_U177 , P2_R1054_U104 , P2_R1054_U10 );
nand NAND2_19123 ( P2_R1054_U178 , P2_R1054_U11 , P2_R1054_U177 );
nand NAND2_19124 ( P2_R1054_U179 , P2_U3430 , P2_R1054_U57 );
nand NAND2_19125 ( P2_R1054_U180 , P2_U3436 , P2_R1054_U55 );
nand NAND3_19126 ( P2_R1054_U181 , P2_R1054_U179 , P2_R1054_U10 , P2_R1054_U94 );
nand NAND2_19127 ( P2_R1054_U182 , P2_R1054_U180 , P2_R1054_U178 );
not NOT1_19128 ( P2_R1054_U183 , P2_R1054_U93 );
nand NAND2_19129 ( P2_R1054_U184 , P2_U3439 , P2_R1054_U60 );
nand NAND2_19130 ( P2_R1054_U185 , P2_R1054_U184 , P2_R1054_U93 );
nand NAND2_19131 ( P2_R1054_U186 , P2_U3565 , P2_R1054_U59 );
not NOT1_19132 ( P2_R1054_U187 , P2_R1054_U61 );
nand NAND2_19133 ( P2_R1054_U188 , P2_R1054_U187 , P2_R1054_U62 );
nand NAND2_19134 ( P2_R1054_U189 , P2_R1054_U188 , P2_R1054_U92 );
nand NAND2_19135 ( P2_R1054_U190 , P2_U3564 , P2_R1054_U61 );
not NOT1_19136 ( P2_R1054_U191 , P2_R1054_U91 );
nand NAND2_19137 ( P2_R1054_U192 , P2_R1054_U179 , P2_R1054_U94 );
not NOT1_19138 ( P2_R1054_U193 , P2_R1054_U63 );
nand NAND2_19139 ( P2_R1054_U194 , P2_U3567 , P2_R1054_U53 );
nand NAND2_19140 ( P2_R1054_U195 , P2_R1054_U193 , P2_R1054_U194 );
nand NAND3_19141 ( P2_R1054_U196 , P2_R1054_U269 , P2_R1054_U100 , P2_R1054_U195 );
nand NAND2_19142 ( P2_R1054_U197 , P2_R1054_U63 , P2_R1054_U100 );
nand NAND2_19143 ( P2_R1054_U198 , P2_U3436 , P2_R1054_U55 );
nand NAND3_19144 ( P2_R1054_U199 , P2_R1054_U198 , P2_R1054_U11 , P2_R1054_U197 );
nand NAND2_19145 ( P2_R1054_U200 , P2_U3567 , P2_R1054_U53 );
nand NAND2_19146 ( P2_R1054_U201 , P2_R1054_U100 , P2_R1054_U200 );
nand NAND2_19147 ( P2_R1054_U202 , P2_R1054_U179 , P2_R1054_U58 );
nand NAND2_19148 ( P2_R1054_U203 , P2_R1054_U134 , P2_R1054_U86 );
not NOT1_19149 ( P2_R1054_U204 , P2_R1054_U64 );
nand NAND2_19150 ( P2_R1054_U205 , P2_U3572 , P2_R1054_U44 );
nand NAND2_19151 ( P2_R1054_U206 , P2_R1054_U204 , P2_R1054_U205 );
nand NAND3_19152 ( P2_R1054_U207 , P2_R1054_U290 , P2_R1054_U99 , P2_R1054_U206 );
nand NAND2_19153 ( P2_R1054_U208 , P2_R1054_U64 , P2_R1054_U99 );
nand NAND2_19154 ( P2_R1054_U209 , P2_U3421 , P2_R1054_U45 );
nand NAND3_19155 ( P2_R1054_U210 , P2_R1054_U209 , P2_R1054_U9 , P2_R1054_U208 );
nand NAND2_19156 ( P2_R1054_U211 , P2_U3572 , P2_R1054_U44 );
nand NAND2_19157 ( P2_R1054_U212 , P2_R1054_U99 , P2_R1054_U211 );
nand NAND2_19158 ( P2_R1054_U213 , P2_U3574 , P2_R1054_U20 );
nand NAND2_19159 ( P2_R1054_U214 , P2_U3415 , P2_R1054_U39 );
nand NAND2_19160 ( P2_R1054_U215 , P2_U3555 , P2_R1054_U38 );
nand NAND2_19161 ( P2_R1054_U216 , P2_R1054_U135 , P2_R1054_U86 );
nand NAND3_19162 ( P2_R1054_U217 , P2_R1054_U215 , P2_R1054_U214 , P2_R1054_U133 );
nand NAND2_19163 ( P2_R1054_U218 , P2_U3412 , P2_R1054_U37 );
nand NAND2_19164 ( P2_R1054_U219 , P2_U3556 , P2_R1054_U34 );
nand NAND2_19165 ( P2_R1054_U220 , P2_U3412 , P2_R1054_U37 );
nand NAND2_19166 ( P2_R1054_U221 , P2_U3556 , P2_R1054_U34 );
nand NAND2_19167 ( P2_R1054_U222 , P2_R1054_U221 , P2_R1054_U220 );
nand NAND2_19168 ( P2_R1054_U223 , P2_U3409 , P2_R1054_U35 );
nand NAND2_19169 ( P2_R1054_U224 , P2_U3557 , P2_R1054_U18 );
nand NAND2_19170 ( P2_R1054_U225 , P2_R1054_U140 , P2_R1054_U40 );
nand NAND3_19171 ( P2_R1054_U226 , P2_R1054_U224 , P2_R1054_U223 , P2_R1054_U127 );
nand NAND2_19172 ( P2_R1054_U227 , P2_U3406 , P2_R1054_U30 );
nand NAND2_19173 ( P2_R1054_U228 , P2_U3558 , P2_R1054_U27 );
nand NAND2_19174 ( P2_R1054_U229 , P2_R1054_U228 , P2_R1054_U227 );
nand NAND2_19175 ( P2_R1054_U230 , P2_U3403 , P2_R1054_U31 );
nand NAND2_19176 ( P2_R1054_U231 , P2_U3559 , P2_R1054_U28 );
nand NAND2_19177 ( P2_R1054_U232 , P2_R1054_U150 , P2_R1054_U41 );
nand NAND3_19178 ( P2_R1054_U233 , P2_R1054_U231 , P2_R1054_U230 , P2_R1054_U142 );
nand NAND2_19179 ( P2_R1054_U234 , P2_U3400 , P2_R1054_U32 );
nand NAND2_19180 ( P2_R1054_U235 , P2_U3560 , P2_R1054_U29 );
nand NAND2_19181 ( P2_R1054_U236 , P2_R1054_U151 , P2_R1054_U87 );
nand NAND3_19182 ( P2_R1054_U237 , P2_R1054_U235 , P2_R1054_U234 , P2_R1054_U117 );
nand NAND2_19183 ( P2_R1054_U238 , P2_U3397 , P2_R1054_U26 );
nand NAND2_19184 ( P2_R1054_U239 , P2_U3561 , P2_R1054_U23 );
nand NAND2_19185 ( P2_R1054_U240 , P2_U3397 , P2_R1054_U26 );
nand NAND2_19186 ( P2_R1054_U241 , P2_U3561 , P2_R1054_U23 );
nand NAND2_19187 ( P2_R1054_U242 , P2_R1054_U241 , P2_R1054_U240 );
nand NAND2_19188 ( P2_R1054_U243 , P2_U3394 , P2_R1054_U24 );
nand NAND2_19189 ( P2_R1054_U244 , P2_U3562 , P2_R1054_U19 );
nand NAND2_19190 ( P2_R1054_U245 , P2_R1054_U156 , P2_R1054_U42 );
nand NAND3_19191 ( P2_R1054_U246 , P2_R1054_U244 , P2_R1054_U243 , P2_R1054_U111 );
nand NAND2_19192 ( P2_R1054_U247 , P2_U3391 , P2_R1054_U22 );
nand NAND2_19193 ( P2_R1054_U248 , P2_U3573 , P2_R1054_U88 );
not NOT1_19194 ( P2_R1054_U249 , P2_R1054_U80 );
nand NAND2_19195 ( P2_R1054_U250 , P2_R1054_U249 , P2_R1054_U107 );
nand NAND2_19196 ( P2_R1054_U251 , P2_R1054_U80 , P2_R1054_U21 );
nand NAND2_19197 ( P2_R1054_U252 , P2_U3379 , P2_R1054_U90 );
nand NAND2_19198 ( P2_R1054_U253 , P2_U3563 , P2_R1054_U89 );
not NOT1_19199 ( P2_R1054_U254 , P2_R1054_U81 );
nand NAND2_19200 ( P2_R1054_U255 , P2_R1054_U191 , P2_R1054_U254 );
nand NAND2_19201 ( P2_R1054_U256 , P2_R1054_U81 , P2_R1054_U91 );
nand NAND2_19202 ( P2_R1054_U257 , P2_U3442 , P2_R1054_U62 );
nand NAND2_19203 ( P2_R1054_U258 , P2_U3564 , P2_R1054_U92 );
not NOT1_19204 ( P2_R1054_U259 , P2_R1054_U82 );
nand NAND2_19205 ( P2_R1054_U260 , P2_R1054_U259 , P2_R1054_U187 );
nand NAND2_19206 ( P2_R1054_U261 , P2_R1054_U82 , P2_R1054_U61 );
nand NAND2_19207 ( P2_R1054_U262 , P2_U3439 , P2_R1054_U60 );
nand NAND2_19208 ( P2_R1054_U263 , P2_U3565 , P2_R1054_U59 );
not NOT1_19209 ( P2_R1054_U264 , P2_R1054_U83 );
nand NAND2_19210 ( P2_R1054_U265 , P2_R1054_U183 , P2_R1054_U264 );
nand NAND2_19211 ( P2_R1054_U266 , P2_R1054_U83 , P2_R1054_U93 );
nand NAND2_19212 ( P2_R1054_U267 , P2_U3436 , P2_R1054_U55 );
nand NAND2_19213 ( P2_R1054_U268 , P2_U3566 , P2_R1054_U52 );
nand NAND2_19214 ( P2_R1054_U269 , P2_R1054_U268 , P2_R1054_U267 );
nand NAND2_19215 ( P2_R1054_U270 , P2_U3433 , P2_R1054_U56 );
nand NAND2_19216 ( P2_R1054_U271 , P2_U3567 , P2_R1054_U53 );
nand NAND2_19217 ( P2_R1054_U272 , P2_R1054_U201 , P2_R1054_U63 );
nand NAND3_19218 ( P2_R1054_U273 , P2_R1054_U271 , P2_R1054_U270 , P2_R1054_U193 );
nand NAND2_19219 ( P2_R1054_U274 , P2_U3430 , P2_R1054_U57 );
nand NAND2_19220 ( P2_R1054_U275 , P2_U3568 , P2_R1054_U54 );
nand NAND2_19221 ( P2_R1054_U276 , P2_R1054_U202 , P2_R1054_U94 );
nand NAND3_19222 ( P2_R1054_U277 , P2_R1054_U275 , P2_R1054_U274 , P2_R1054_U173 );
nand NAND2_19223 ( P2_R1054_U278 , P2_U3427 , P2_R1054_U51 );
nand NAND2_19224 ( P2_R1054_U279 , P2_U3569 , P2_R1054_U50 );
not NOT1_19225 ( P2_R1054_U280 , P2_R1054_U84 );
nand NAND2_19226 ( P2_R1054_U281 , P2_R1054_U169 , P2_R1054_U280 );
nand NAND2_19227 ( P2_R1054_U282 , P2_R1054_U84 , P2_R1054_U95 );
nand NAND2_19228 ( P2_R1054_U283 , P2_U3424 , P2_R1054_U49 );
nand NAND2_19229 ( P2_R1054_U284 , P2_U3570 , P2_R1054_U48 );
not NOT1_19230 ( P2_R1054_U285 , P2_R1054_U85 );
nand NAND2_19231 ( P2_R1054_U286 , P2_R1054_U165 , P2_R1054_U285 );
nand NAND2_19232 ( P2_R1054_U287 , P2_R1054_U85 , P2_R1054_U96 );
nand NAND2_19233 ( P2_R1054_U288 , P2_U3421 , P2_R1054_U45 );
nand NAND2_19234 ( P2_R1054_U289 , P2_U3571 , P2_R1054_U43 );
nand NAND2_19235 ( P2_R1054_U290 , P2_R1054_U289 , P2_R1054_U288 );
nand NAND2_19236 ( P2_R1054_U291 , P2_U3418 , P2_R1054_U46 );
nand NAND2_19237 ( P2_R1054_U292 , P2_U3572 , P2_R1054_U44 );
nand NAND2_19238 ( P2_R1054_U293 , P2_R1054_U212 , P2_R1054_U64 );
nand NAND3_19239 ( P2_R1054_U294 , P2_R1054_U292 , P2_R1054_U291 , P2_R1054_U204 );
and AND2_19240 ( P2_R1161_U4 , P2_R1161_U179 , P2_R1161_U178 );
and AND2_19241 ( P2_R1161_U5 , P2_R1161_U197 , P2_R1161_U196 );
and AND2_19242 ( P2_R1161_U6 , P2_R1161_U237 , P2_R1161_U236 );
and AND2_19243 ( P2_R1161_U7 , P2_R1161_U246 , P2_R1161_U245 );
and AND2_19244 ( P2_R1161_U8 , P2_R1161_U264 , P2_R1161_U263 );
and AND2_19245 ( P2_R1161_U9 , P2_R1161_U272 , P2_R1161_U271 );
and AND2_19246 ( P2_R1161_U10 , P2_R1161_U351 , P2_R1161_U348 );
and AND2_19247 ( P2_R1161_U11 , P2_R1161_U344 , P2_R1161_U341 );
and AND2_19248 ( P2_R1161_U12 , P2_R1161_U335 , P2_R1161_U332 );
and AND2_19249 ( P2_R1161_U13 , P2_R1161_U326 , P2_R1161_U323 );
and AND2_19250 ( P2_R1161_U14 , P2_R1161_U320 , P2_R1161_U318 );
and AND2_19251 ( P2_R1161_U15 , P2_R1161_U313 , P2_R1161_U310 );
and AND2_19252 ( P2_R1161_U16 , P2_R1161_U235 , P2_R1161_U232 );
and AND2_19253 ( P2_R1161_U17 , P2_R1161_U227 , P2_R1161_U224 );
and AND2_19254 ( P2_R1161_U18 , P2_R1161_U213 , P2_R1161_U210 );
not NOT1_19255 ( P2_R1161_U19 , P2_U3407 );
not NOT1_19256 ( P2_R1161_U20 , P2_U3070 );
not NOT1_19257 ( P2_R1161_U21 , P2_U3069 );
nand NAND2_19258 ( P2_R1161_U22 , P2_U3070 , P2_U3407 );
not NOT1_19259 ( P2_R1161_U23 , P2_U3410 );
not NOT1_19260 ( P2_R1161_U24 , P2_U3401 );
not NOT1_19261 ( P2_R1161_U25 , P2_U3059 );
not NOT1_19262 ( P2_R1161_U26 , P2_U3066 );
not NOT1_19263 ( P2_R1161_U27 , P2_U3395 );
not NOT1_19264 ( P2_R1161_U28 , P2_U3067 );
not NOT1_19265 ( P2_R1161_U29 , P2_U3387 );
not NOT1_19266 ( P2_R1161_U30 , P2_U3076 );
nand NAND2_19267 ( P2_R1161_U31 , P2_U3076 , P2_U3387 );
not NOT1_19268 ( P2_R1161_U32 , P2_U3398 );
not NOT1_19269 ( P2_R1161_U33 , P2_U3063 );
nand NAND2_19270 ( P2_R1161_U34 , P2_U3059 , P2_U3401 );
not NOT1_19271 ( P2_R1161_U35 , P2_U3404 );
not NOT1_19272 ( P2_R1161_U36 , P2_U3413 );
not NOT1_19273 ( P2_R1161_U37 , P2_U3083 );
not NOT1_19274 ( P2_R1161_U38 , P2_U3082 );
not NOT1_19275 ( P2_R1161_U39 , P2_U3416 );
nand NAND2_19276 ( P2_R1161_U40 , P2_R1161_U65 , P2_R1161_U205 );
nand NAND2_19277 ( P2_R1161_U41 , P2_R1161_U117 , P2_R1161_U193 );
nand NAND2_19278 ( P2_R1161_U42 , P2_R1161_U182 , P2_R1161_U183 );
nand NAND2_19279 ( P2_R1161_U43 , P2_U3392 , P2_U3077 );
nand NAND2_19280 ( P2_R1161_U44 , P2_R1161_U122 , P2_R1161_U219 );
nand NAND2_19281 ( P2_R1161_U45 , P2_R1161_U216 , P2_R1161_U215 );
not NOT1_19282 ( P2_R1161_U46 , P2_U3896 );
not NOT1_19283 ( P2_R1161_U47 , P2_U3052 );
not NOT1_19284 ( P2_R1161_U48 , P2_U3056 );
not NOT1_19285 ( P2_R1161_U49 , P2_U3897 );
not NOT1_19286 ( P2_R1161_U50 , P2_U3898 );
not NOT1_19287 ( P2_R1161_U51 , P2_U3057 );
not NOT1_19288 ( P2_R1161_U52 , P2_U3899 );
not NOT1_19289 ( P2_R1161_U53 , P2_U3064 );
not NOT1_19290 ( P2_R1161_U54 , P2_U3902 );
not NOT1_19291 ( P2_R1161_U55 , P2_U3074 );
not NOT1_19292 ( P2_R1161_U56 , P2_U3437 );
not NOT1_19293 ( P2_R1161_U57 , P2_U3072 );
not NOT1_19294 ( P2_R1161_U58 , P2_U3068 );
nand NAND2_19295 ( P2_R1161_U59 , P2_U3072 , P2_U3437 );
not NOT1_19296 ( P2_R1161_U60 , P2_U3440 );
not NOT1_19297 ( P2_R1161_U61 , P2_U3428 );
not NOT1_19298 ( P2_R1161_U62 , P2_U3079 );
not NOT1_19299 ( P2_R1161_U63 , P2_U3419 );
not NOT1_19300 ( P2_R1161_U64 , P2_U3061 );
nand NAND2_19301 ( P2_R1161_U65 , P2_U3083 , P2_U3413 );
not NOT1_19302 ( P2_R1161_U66 , P2_U3422 );
not NOT1_19303 ( P2_R1161_U67 , P2_U3062 );
nand NAND2_19304 ( P2_R1161_U68 , P2_U3062 , P2_U3422 );
not NOT1_19305 ( P2_R1161_U69 , P2_U3425 );
not NOT1_19306 ( P2_R1161_U70 , P2_U3071 );
not NOT1_19307 ( P2_R1161_U71 , P2_U3431 );
not NOT1_19308 ( P2_R1161_U72 , P2_U3078 );
not NOT1_19309 ( P2_R1161_U73 , P2_U3434 );
not NOT1_19310 ( P2_R1161_U74 , P2_U3073 );
not NOT1_19311 ( P2_R1161_U75 , P2_U3443 );
not NOT1_19312 ( P2_R1161_U76 , P2_U3081 );
nand NAND2_19313 ( P2_R1161_U77 , P2_U3081 , P2_U3443 );
not NOT1_19314 ( P2_R1161_U78 , P2_U3445 );
not NOT1_19315 ( P2_R1161_U79 , P2_U3080 );
nand NAND2_19316 ( P2_R1161_U80 , P2_U3080 , P2_U3445 );
not NOT1_19317 ( P2_R1161_U81 , P2_U3903 );
not NOT1_19318 ( P2_R1161_U82 , P2_U3901 );
not NOT1_19319 ( P2_R1161_U83 , P2_U3060 );
not NOT1_19320 ( P2_R1161_U84 , P2_U3900 );
not NOT1_19321 ( P2_R1161_U85 , P2_U3065 );
nand NAND2_19322 ( P2_R1161_U86 , P2_U3897 , P2_U3056 );
not NOT1_19323 ( P2_R1161_U87 , P2_U3053 );
not NOT1_19324 ( P2_R1161_U88 , P2_U3895 );
nand NAND2_19325 ( P2_R1161_U89 , P2_R1161_U306 , P2_R1161_U176 );
not NOT1_19326 ( P2_R1161_U90 , P2_U3075 );
nand NAND2_19327 ( P2_R1161_U91 , P2_R1161_U77 , P2_R1161_U315 );
nand NAND2_19328 ( P2_R1161_U92 , P2_R1161_U261 , P2_R1161_U260 );
nand NAND2_19329 ( P2_R1161_U93 , P2_R1161_U68 , P2_R1161_U337 );
nand NAND2_19330 ( P2_R1161_U94 , P2_R1161_U457 , P2_R1161_U456 );
nand NAND2_19331 ( P2_R1161_U95 , P2_R1161_U504 , P2_R1161_U503 );
nand NAND2_19332 ( P2_R1161_U96 , P2_R1161_U375 , P2_R1161_U374 );
nand NAND2_19333 ( P2_R1161_U97 , P2_R1161_U380 , P2_R1161_U379 );
nand NAND2_19334 ( P2_R1161_U98 , P2_R1161_U387 , P2_R1161_U386 );
nand NAND2_19335 ( P2_R1161_U99 , P2_R1161_U394 , P2_R1161_U393 );
nand NAND2_19336 ( P2_R1161_U100 , P2_R1161_U399 , P2_R1161_U398 );
nand NAND2_19337 ( P2_R1161_U101 , P2_R1161_U408 , P2_R1161_U407 );
nand NAND2_19338 ( P2_R1161_U102 , P2_R1161_U415 , P2_R1161_U414 );
nand NAND2_19339 ( P2_R1161_U103 , P2_R1161_U422 , P2_R1161_U421 );
nand NAND2_19340 ( P2_R1161_U104 , P2_R1161_U429 , P2_R1161_U428 );
nand NAND2_19341 ( P2_R1161_U105 , P2_R1161_U434 , P2_R1161_U433 );
nand NAND2_19342 ( P2_R1161_U106 , P2_R1161_U441 , P2_R1161_U440 );
nand NAND2_19343 ( P2_R1161_U107 , P2_R1161_U448 , P2_R1161_U447 );
nand NAND2_19344 ( P2_R1161_U108 , P2_R1161_U462 , P2_R1161_U461 );
nand NAND2_19345 ( P2_R1161_U109 , P2_R1161_U467 , P2_R1161_U466 );
nand NAND2_19346 ( P2_R1161_U110 , P2_R1161_U474 , P2_R1161_U473 );
nand NAND2_19347 ( P2_R1161_U111 , P2_R1161_U481 , P2_R1161_U480 );
nand NAND2_19348 ( P2_R1161_U112 , P2_R1161_U488 , P2_R1161_U487 );
nand NAND2_19349 ( P2_R1161_U113 , P2_R1161_U495 , P2_R1161_U494 );
nand NAND2_19350 ( P2_R1161_U114 , P2_R1161_U500 , P2_R1161_U499 );
and AND2_19351 ( P2_R1161_U115 , P2_R1161_U189 , P2_R1161_U187 );
and AND2_19352 ( P2_R1161_U116 , P2_R1161_U4 , P2_R1161_U180 );
and AND2_19353 ( P2_R1161_U117 , P2_R1161_U194 , P2_R1161_U192 );
and AND2_19354 ( P2_R1161_U118 , P2_R1161_U201 , P2_R1161_U200 );
and AND3_19355 ( P2_R1161_U119 , P2_R1161_U382 , P2_R1161_U381 , P2_R1161_U22 );
and AND2_19356 ( P2_R1161_U120 , P2_R1161_U212 , P2_R1161_U5 );
and AND2_19357 ( P2_R1161_U121 , P2_R1161_U181 , P2_R1161_U180 );
and AND2_19358 ( P2_R1161_U122 , P2_R1161_U220 , P2_R1161_U218 );
and AND3_19359 ( P2_R1161_U123 , P2_R1161_U389 , P2_R1161_U388 , P2_R1161_U34 );
and AND2_19360 ( P2_R1161_U124 , P2_R1161_U226 , P2_R1161_U4 );
and AND2_19361 ( P2_R1161_U125 , P2_R1161_U234 , P2_R1161_U181 );
and AND2_19362 ( P2_R1161_U126 , P2_R1161_U204 , P2_R1161_U6 );
and AND2_19363 ( P2_R1161_U127 , P2_R1161_U243 , P2_R1161_U239 );
and AND2_19364 ( P2_R1161_U128 , P2_R1161_U250 , P2_R1161_U7 );
and AND2_19365 ( P2_R1161_U129 , P2_R1161_U253 , P2_R1161_U248 );
and AND2_19366 ( P2_R1161_U130 , P2_R1161_U268 , P2_R1161_U267 );
and AND2_19367 ( P2_R1161_U131 , P2_R1161_U9 , P2_R1161_U282 );
and AND2_19368 ( P2_R1161_U132 , P2_R1161_U285 , P2_R1161_U280 );
and AND2_19369 ( P2_R1161_U133 , P2_R1161_U301 , P2_R1161_U298 );
and AND2_19370 ( P2_R1161_U134 , P2_R1161_U368 , P2_R1161_U302 );
and AND2_19371 ( P2_R1161_U135 , P2_R1161_U160 , P2_R1161_U278 );
and AND3_19372 ( P2_R1161_U136 , P2_R1161_U455 , P2_R1161_U454 , P2_R1161_U80 );
and AND2_19373 ( P2_R1161_U137 , P2_R1161_U325 , P2_R1161_U9 );
and AND3_19374 ( P2_R1161_U138 , P2_R1161_U469 , P2_R1161_U468 , P2_R1161_U59 );
and AND2_19375 ( P2_R1161_U139 , P2_R1161_U334 , P2_R1161_U8 );
and AND3_19376 ( P2_R1161_U140 , P2_R1161_U490 , P2_R1161_U489 , P2_R1161_U172 );
and AND2_19377 ( P2_R1161_U141 , P2_R1161_U343 , P2_R1161_U7 );
and AND3_19378 ( P2_R1161_U142 , P2_R1161_U502 , P2_R1161_U501 , P2_R1161_U171 );
and AND2_19379 ( P2_R1161_U143 , P2_R1161_U350 , P2_R1161_U6 );
nand NAND2_19380 ( P2_R1161_U144 , P2_R1161_U118 , P2_R1161_U202 );
nand NAND2_19381 ( P2_R1161_U145 , P2_R1161_U217 , P2_R1161_U229 );
not NOT1_19382 ( P2_R1161_U146 , P2_U3054 );
not NOT1_19383 ( P2_R1161_U147 , P2_U3904 );
and AND2_19384 ( P2_R1161_U148 , P2_R1161_U403 , P2_R1161_U402 );
nand NAND3_19385 ( P2_R1161_U149 , P2_R1161_U304 , P2_R1161_U169 , P2_R1161_U364 );
and AND2_19386 ( P2_R1161_U150 , P2_R1161_U410 , P2_R1161_U409 );
nand NAND3_19387 ( P2_R1161_U151 , P2_R1161_U370 , P2_R1161_U369 , P2_R1161_U134 );
and AND2_19388 ( P2_R1161_U152 , P2_R1161_U417 , P2_R1161_U416 );
nand NAND3_19389 ( P2_R1161_U153 , P2_R1161_U365 , P2_R1161_U299 , P2_R1161_U86 );
and AND2_19390 ( P2_R1161_U154 , P2_R1161_U424 , P2_R1161_U423 );
nand NAND2_19391 ( P2_R1161_U155 , P2_R1161_U293 , P2_R1161_U292 );
and AND2_19392 ( P2_R1161_U156 , P2_R1161_U436 , P2_R1161_U435 );
nand NAND2_19393 ( P2_R1161_U157 , P2_R1161_U289 , P2_R1161_U288 );
and AND2_19394 ( P2_R1161_U158 , P2_R1161_U443 , P2_R1161_U442 );
nand NAND2_19395 ( P2_R1161_U159 , P2_R1161_U132 , P2_R1161_U284 );
and AND2_19396 ( P2_R1161_U160 , P2_R1161_U450 , P2_R1161_U449 );
nand NAND2_19397 ( P2_R1161_U161 , P2_R1161_U43 , P2_R1161_U327 );
nand NAND2_19398 ( P2_R1161_U162 , P2_R1161_U130 , P2_R1161_U269 );
and AND2_19399 ( P2_R1161_U163 , P2_R1161_U476 , P2_R1161_U475 );
nand NAND2_19400 ( P2_R1161_U164 , P2_R1161_U257 , P2_R1161_U256 );
and AND2_19401 ( P2_R1161_U165 , P2_R1161_U483 , P2_R1161_U482 );
nand NAND2_19402 ( P2_R1161_U166 , P2_R1161_U129 , P2_R1161_U252 );
nand NAND2_19403 ( P2_R1161_U167 , P2_R1161_U127 , P2_R1161_U242 );
nand NAND2_19404 ( P2_R1161_U168 , P2_R1161_U367 , P2_R1161_U366 );
nand NAND2_19405 ( P2_R1161_U169 , P2_U3053 , P2_R1161_U151 );
not NOT1_19406 ( P2_R1161_U170 , P2_R1161_U34 );
nand NAND2_19407 ( P2_R1161_U171 , P2_U3416 , P2_U3082 );
nand NAND2_19408 ( P2_R1161_U172 , P2_U3071 , P2_U3425 );
nand NAND2_19409 ( P2_R1161_U173 , P2_U3057 , P2_U3898 );
not NOT1_19410 ( P2_R1161_U174 , P2_R1161_U68 );
not NOT1_19411 ( P2_R1161_U175 , P2_R1161_U77 );
nand NAND2_19412 ( P2_R1161_U176 , P2_U3064 , P2_U3899 );
not NOT1_19413 ( P2_R1161_U177 , P2_R1161_U65 );
or OR2_19414 ( P2_R1161_U178 , P2_U3066 , P2_U3404 );
or OR2_19415 ( P2_R1161_U179 , P2_U3059 , P2_U3401 );
or OR2_19416 ( P2_R1161_U180 , P2_U3398 , P2_U3063 );
or OR2_19417 ( P2_R1161_U181 , P2_U3395 , P2_U3067 );
not NOT1_19418 ( P2_R1161_U182 , P2_R1161_U31 );
or OR2_19419 ( P2_R1161_U183 , P2_U3392 , P2_U3077 );
not NOT1_19420 ( P2_R1161_U184 , P2_R1161_U42 );
not NOT1_19421 ( P2_R1161_U185 , P2_R1161_U43 );
nand NAND2_19422 ( P2_R1161_U186 , P2_R1161_U42 , P2_R1161_U43 );
nand NAND2_19423 ( P2_R1161_U187 , P2_U3067 , P2_U3395 );
nand NAND2_19424 ( P2_R1161_U188 , P2_R1161_U186 , P2_R1161_U181 );
nand NAND2_19425 ( P2_R1161_U189 , P2_U3063 , P2_U3398 );
nand NAND2_19426 ( P2_R1161_U190 , P2_R1161_U115 , P2_R1161_U188 );
nand NAND2_19427 ( P2_R1161_U191 , P2_R1161_U35 , P2_R1161_U34 );
nand NAND2_19428 ( P2_R1161_U192 , P2_U3066 , P2_R1161_U191 );
nand NAND2_19429 ( P2_R1161_U193 , P2_R1161_U116 , P2_R1161_U190 );
nand NAND2_19430 ( P2_R1161_U194 , P2_U3404 , P2_R1161_U170 );
not NOT1_19431 ( P2_R1161_U195 , P2_R1161_U41 );
or OR2_19432 ( P2_R1161_U196 , P2_U3069 , P2_U3410 );
or OR2_19433 ( P2_R1161_U197 , P2_U3070 , P2_U3407 );
not NOT1_19434 ( P2_R1161_U198 , P2_R1161_U22 );
nand NAND2_19435 ( P2_R1161_U199 , P2_R1161_U23 , P2_R1161_U22 );
nand NAND2_19436 ( P2_R1161_U200 , P2_U3069 , P2_R1161_U199 );
nand NAND2_19437 ( P2_R1161_U201 , P2_U3410 , P2_R1161_U198 );
nand NAND2_19438 ( P2_R1161_U202 , P2_R1161_U5 , P2_R1161_U41 );
not NOT1_19439 ( P2_R1161_U203 , P2_R1161_U144 );
or OR2_19440 ( P2_R1161_U204 , P2_U3413 , P2_U3083 );
nand NAND2_19441 ( P2_R1161_U205 , P2_R1161_U204 , P2_R1161_U144 );
not NOT1_19442 ( P2_R1161_U206 , P2_R1161_U40 );
or OR2_19443 ( P2_R1161_U207 , P2_U3082 , P2_U3416 );
or OR2_19444 ( P2_R1161_U208 , P2_U3407 , P2_U3070 );
nand NAND2_19445 ( P2_R1161_U209 , P2_R1161_U208 , P2_R1161_U41 );
nand NAND2_19446 ( P2_R1161_U210 , P2_R1161_U119 , P2_R1161_U209 );
nand NAND2_19447 ( P2_R1161_U211 , P2_R1161_U195 , P2_R1161_U22 );
nand NAND2_19448 ( P2_R1161_U212 , P2_U3410 , P2_U3069 );
nand NAND2_19449 ( P2_R1161_U213 , P2_R1161_U120 , P2_R1161_U211 );
or OR2_19450 ( P2_R1161_U214 , P2_U3070 , P2_U3407 );
nand NAND2_19451 ( P2_R1161_U215 , P2_R1161_U185 , P2_R1161_U181 );
nand NAND2_19452 ( P2_R1161_U216 , P2_U3067 , P2_U3395 );
not NOT1_19453 ( P2_R1161_U217 , P2_R1161_U45 );
nand NAND2_19454 ( P2_R1161_U218 , P2_R1161_U121 , P2_R1161_U184 );
nand NAND2_19455 ( P2_R1161_U219 , P2_R1161_U45 , P2_R1161_U180 );
nand NAND2_19456 ( P2_R1161_U220 , P2_U3063 , P2_U3398 );
not NOT1_19457 ( P2_R1161_U221 , P2_R1161_U44 );
or OR2_19458 ( P2_R1161_U222 , P2_U3401 , P2_U3059 );
nand NAND2_19459 ( P2_R1161_U223 , P2_R1161_U222 , P2_R1161_U44 );
nand NAND2_19460 ( P2_R1161_U224 , P2_R1161_U123 , P2_R1161_U223 );
nand NAND2_19461 ( P2_R1161_U225 , P2_R1161_U221 , P2_R1161_U34 );
nand NAND2_19462 ( P2_R1161_U226 , P2_U3404 , P2_U3066 );
nand NAND2_19463 ( P2_R1161_U227 , P2_R1161_U124 , P2_R1161_U225 );
or OR2_19464 ( P2_R1161_U228 , P2_U3059 , P2_U3401 );
nand NAND2_19465 ( P2_R1161_U229 , P2_R1161_U184 , P2_R1161_U181 );
not NOT1_19466 ( P2_R1161_U230 , P2_R1161_U145 );
nand NAND2_19467 ( P2_R1161_U231 , P2_U3063 , P2_U3398 );
nand NAND4_19468 ( P2_R1161_U232 , P2_R1161_U401 , P2_R1161_U400 , P2_R1161_U43 , P2_R1161_U42 );
nand NAND2_19469 ( P2_R1161_U233 , P2_R1161_U43 , P2_R1161_U42 );
nand NAND2_19470 ( P2_R1161_U234 , P2_U3067 , P2_U3395 );
nand NAND2_19471 ( P2_R1161_U235 , P2_R1161_U125 , P2_R1161_U233 );
or OR2_19472 ( P2_R1161_U236 , P2_U3082 , P2_U3416 );
or OR2_19473 ( P2_R1161_U237 , P2_U3061 , P2_U3419 );
nand NAND2_19474 ( P2_R1161_U238 , P2_R1161_U177 , P2_R1161_U6 );
nand NAND2_19475 ( P2_R1161_U239 , P2_U3061 , P2_U3419 );
nand NAND2_19476 ( P2_R1161_U240 , P2_R1161_U171 , P2_R1161_U238 );
or OR2_19477 ( P2_R1161_U241 , P2_U3419 , P2_U3061 );
nand NAND2_19478 ( P2_R1161_U242 , P2_R1161_U126 , P2_R1161_U144 );
nand NAND2_19479 ( P2_R1161_U243 , P2_R1161_U241 , P2_R1161_U240 );
not NOT1_19480 ( P2_R1161_U244 , P2_R1161_U167 );
or OR2_19481 ( P2_R1161_U245 , P2_U3079 , P2_U3428 );
or OR2_19482 ( P2_R1161_U246 , P2_U3071 , P2_U3425 );
nand NAND2_19483 ( P2_R1161_U247 , P2_R1161_U174 , P2_R1161_U7 );
nand NAND2_19484 ( P2_R1161_U248 , P2_U3079 , P2_U3428 );
nand NAND2_19485 ( P2_R1161_U249 , P2_R1161_U172 , P2_R1161_U247 );
or OR2_19486 ( P2_R1161_U250 , P2_U3422 , P2_U3062 );
or OR2_19487 ( P2_R1161_U251 , P2_U3428 , P2_U3079 );
nand NAND2_19488 ( P2_R1161_U252 , P2_R1161_U128 , P2_R1161_U167 );
nand NAND2_19489 ( P2_R1161_U253 , P2_R1161_U251 , P2_R1161_U249 );
not NOT1_19490 ( P2_R1161_U254 , P2_R1161_U166 );
or OR2_19491 ( P2_R1161_U255 , P2_U3431 , P2_U3078 );
nand NAND2_19492 ( P2_R1161_U256 , P2_R1161_U255 , P2_R1161_U166 );
nand NAND2_19493 ( P2_R1161_U257 , P2_U3078 , P2_U3431 );
not NOT1_19494 ( P2_R1161_U258 , P2_R1161_U164 );
or OR2_19495 ( P2_R1161_U259 , P2_U3434 , P2_U3073 );
nand NAND2_19496 ( P2_R1161_U260 , P2_R1161_U259 , P2_R1161_U164 );
nand NAND2_19497 ( P2_R1161_U261 , P2_U3073 , P2_U3434 );
not NOT1_19498 ( P2_R1161_U262 , P2_R1161_U92 );
or OR2_19499 ( P2_R1161_U263 , P2_U3068 , P2_U3440 );
or OR2_19500 ( P2_R1161_U264 , P2_U3072 , P2_U3437 );
not NOT1_19501 ( P2_R1161_U265 , P2_R1161_U59 );
nand NAND2_19502 ( P2_R1161_U266 , P2_R1161_U60 , P2_R1161_U59 );
nand NAND2_19503 ( P2_R1161_U267 , P2_U3068 , P2_R1161_U266 );
nand NAND2_19504 ( P2_R1161_U268 , P2_U3440 , P2_R1161_U265 );
nand NAND2_19505 ( P2_R1161_U269 , P2_R1161_U8 , P2_R1161_U92 );
not NOT1_19506 ( P2_R1161_U270 , P2_R1161_U162 );
or OR2_19507 ( P2_R1161_U271 , P2_U3075 , P2_U3903 );
or OR2_19508 ( P2_R1161_U272 , P2_U3080 , P2_U3445 );
or OR2_19509 ( P2_R1161_U273 , P2_U3074 , P2_U3902 );
not NOT1_19510 ( P2_R1161_U274 , P2_R1161_U80 );
nand NAND2_19511 ( P2_R1161_U275 , P2_U3903 , P2_R1161_U274 );
nand NAND2_19512 ( P2_R1161_U276 , P2_R1161_U275 , P2_R1161_U90 );
nand NAND2_19513 ( P2_R1161_U277 , P2_R1161_U80 , P2_R1161_U81 );
nand NAND2_19514 ( P2_R1161_U278 , P2_R1161_U277 , P2_R1161_U276 );
nand NAND2_19515 ( P2_R1161_U279 , P2_R1161_U175 , P2_R1161_U9 );
nand NAND2_19516 ( P2_R1161_U280 , P2_U3074 , P2_U3902 );
nand NAND2_19517 ( P2_R1161_U281 , P2_R1161_U278 , P2_R1161_U279 );
or OR2_19518 ( P2_R1161_U282 , P2_U3443 , P2_U3081 );
or OR2_19519 ( P2_R1161_U283 , P2_U3902 , P2_U3074 );
nand NAND3_19520 ( P2_R1161_U284 , P2_R1161_U273 , P2_R1161_U162 , P2_R1161_U131 );
nand NAND2_19521 ( P2_R1161_U285 , P2_R1161_U283 , P2_R1161_U281 );
not NOT1_19522 ( P2_R1161_U286 , P2_R1161_U159 );
or OR2_19523 ( P2_R1161_U287 , P2_U3901 , P2_U3060 );
nand NAND2_19524 ( P2_R1161_U288 , P2_R1161_U287 , P2_R1161_U159 );
nand NAND2_19525 ( P2_R1161_U289 , P2_U3060 , P2_U3901 );
not NOT1_19526 ( P2_R1161_U290 , P2_R1161_U157 );
or OR2_19527 ( P2_R1161_U291 , P2_U3900 , P2_U3065 );
nand NAND2_19528 ( P2_R1161_U292 , P2_R1161_U291 , P2_R1161_U157 );
nand NAND2_19529 ( P2_R1161_U293 , P2_U3065 , P2_U3900 );
not NOT1_19530 ( P2_R1161_U294 , P2_R1161_U155 );
or OR2_19531 ( P2_R1161_U295 , P2_U3057 , P2_U3898 );
nand NAND2_19532 ( P2_R1161_U296 , P2_R1161_U176 , P2_R1161_U173 );
not NOT1_19533 ( P2_R1161_U297 , P2_R1161_U86 );
or OR2_19534 ( P2_R1161_U298 , P2_U3899 , P2_U3064 );
nand NAND3_19535 ( P2_R1161_U299 , P2_R1161_U155 , P2_R1161_U298 , P2_R1161_U168 );
not NOT1_19536 ( P2_R1161_U300 , P2_R1161_U153 );
or OR2_19537 ( P2_R1161_U301 , P2_U3896 , P2_U3052 );
nand NAND2_19538 ( P2_R1161_U302 , P2_U3052 , P2_U3896 );
not NOT1_19539 ( P2_R1161_U303 , P2_R1161_U151 );
nand NAND2_19540 ( P2_R1161_U304 , P2_U3895 , P2_R1161_U151 );
not NOT1_19541 ( P2_R1161_U305 , P2_R1161_U149 );
nand NAND2_19542 ( P2_R1161_U306 , P2_R1161_U298 , P2_R1161_U155 );
not NOT1_19543 ( P2_R1161_U307 , P2_R1161_U89 );
or OR2_19544 ( P2_R1161_U308 , P2_U3898 , P2_U3057 );
nand NAND2_19545 ( P2_R1161_U309 , P2_R1161_U308 , P2_R1161_U89 );
nand NAND3_19546 ( P2_R1161_U310 , P2_R1161_U309 , P2_R1161_U173 , P2_R1161_U154 );
nand NAND2_19547 ( P2_R1161_U311 , P2_R1161_U307 , P2_R1161_U173 );
nand NAND2_19548 ( P2_R1161_U312 , P2_U3897 , P2_U3056 );
nand NAND3_19549 ( P2_R1161_U313 , P2_R1161_U311 , P2_R1161_U312 , P2_R1161_U168 );
or OR2_19550 ( P2_R1161_U314 , P2_U3057 , P2_U3898 );
nand NAND2_19551 ( P2_R1161_U315 , P2_R1161_U282 , P2_R1161_U162 );
not NOT1_19552 ( P2_R1161_U316 , P2_R1161_U91 );
nand NAND2_19553 ( P2_R1161_U317 , P2_R1161_U9 , P2_R1161_U91 );
nand NAND2_19554 ( P2_R1161_U318 , P2_R1161_U135 , P2_R1161_U317 );
nand NAND2_19555 ( P2_R1161_U319 , P2_R1161_U317 , P2_R1161_U278 );
nand NAND2_19556 ( P2_R1161_U320 , P2_R1161_U453 , P2_R1161_U319 );
or OR2_19557 ( P2_R1161_U321 , P2_U3445 , P2_U3080 );
nand NAND2_19558 ( P2_R1161_U322 , P2_R1161_U321 , P2_R1161_U91 );
nand NAND2_19559 ( P2_R1161_U323 , P2_R1161_U136 , P2_R1161_U322 );
nand NAND2_19560 ( P2_R1161_U324 , P2_R1161_U316 , P2_R1161_U80 );
nand NAND2_19561 ( P2_R1161_U325 , P2_U3075 , P2_U3903 );
nand NAND2_19562 ( P2_R1161_U326 , P2_R1161_U137 , P2_R1161_U324 );
or OR2_19563 ( P2_R1161_U327 , P2_U3392 , P2_U3077 );
not NOT1_19564 ( P2_R1161_U328 , P2_R1161_U161 );
or OR2_19565 ( P2_R1161_U329 , P2_U3080 , P2_U3445 );
or OR2_19566 ( P2_R1161_U330 , P2_U3437 , P2_U3072 );
nand NAND2_19567 ( P2_R1161_U331 , P2_R1161_U330 , P2_R1161_U92 );
nand NAND2_19568 ( P2_R1161_U332 , P2_R1161_U138 , P2_R1161_U331 );
nand NAND2_19569 ( P2_R1161_U333 , P2_R1161_U262 , P2_R1161_U59 );
nand NAND2_19570 ( P2_R1161_U334 , P2_U3440 , P2_U3068 );
nand NAND2_19571 ( P2_R1161_U335 , P2_R1161_U139 , P2_R1161_U333 );
or OR2_19572 ( P2_R1161_U336 , P2_U3072 , P2_U3437 );
nand NAND2_19573 ( P2_R1161_U337 , P2_R1161_U250 , P2_R1161_U167 );
not NOT1_19574 ( P2_R1161_U338 , P2_R1161_U93 );
or OR2_19575 ( P2_R1161_U339 , P2_U3425 , P2_U3071 );
nand NAND2_19576 ( P2_R1161_U340 , P2_R1161_U339 , P2_R1161_U93 );
nand NAND2_19577 ( P2_R1161_U341 , P2_R1161_U140 , P2_R1161_U340 );
nand NAND2_19578 ( P2_R1161_U342 , P2_R1161_U338 , P2_R1161_U172 );
nand NAND2_19579 ( P2_R1161_U343 , P2_U3079 , P2_U3428 );
nand NAND2_19580 ( P2_R1161_U344 , P2_R1161_U141 , P2_R1161_U342 );
or OR2_19581 ( P2_R1161_U345 , P2_U3071 , P2_U3425 );
or OR2_19582 ( P2_R1161_U346 , P2_U3416 , P2_U3082 );
nand NAND2_19583 ( P2_R1161_U347 , P2_R1161_U346 , P2_R1161_U40 );
nand NAND2_19584 ( P2_R1161_U348 , P2_R1161_U142 , P2_R1161_U347 );
nand NAND2_19585 ( P2_R1161_U349 , P2_R1161_U206 , P2_R1161_U171 );
nand NAND2_19586 ( P2_R1161_U350 , P2_U3061 , P2_U3419 );
nand NAND2_19587 ( P2_R1161_U351 , P2_R1161_U143 , P2_R1161_U349 );
nand NAND2_19588 ( P2_R1161_U352 , P2_R1161_U207 , P2_R1161_U171 );
nand NAND2_19589 ( P2_R1161_U353 , P2_R1161_U204 , P2_R1161_U65 );
nand NAND2_19590 ( P2_R1161_U354 , P2_R1161_U214 , P2_R1161_U22 );
nand NAND2_19591 ( P2_R1161_U355 , P2_R1161_U228 , P2_R1161_U34 );
nand NAND2_19592 ( P2_R1161_U356 , P2_R1161_U231 , P2_R1161_U180 );
nand NAND2_19593 ( P2_R1161_U357 , P2_R1161_U314 , P2_R1161_U173 );
nand NAND2_19594 ( P2_R1161_U358 , P2_R1161_U298 , P2_R1161_U176 );
nand NAND2_19595 ( P2_R1161_U359 , P2_R1161_U329 , P2_R1161_U80 );
nand NAND2_19596 ( P2_R1161_U360 , P2_R1161_U282 , P2_R1161_U77 );
nand NAND2_19597 ( P2_R1161_U361 , P2_R1161_U336 , P2_R1161_U59 );
nand NAND2_19598 ( P2_R1161_U362 , P2_R1161_U345 , P2_R1161_U172 );
nand NAND2_19599 ( P2_R1161_U363 , P2_R1161_U250 , P2_R1161_U68 );
nand NAND2_19600 ( P2_R1161_U364 , P2_U3895 , P2_U3053 );
nand NAND2_19601 ( P2_R1161_U365 , P2_R1161_U296 , P2_R1161_U168 );
nand NAND2_19602 ( P2_R1161_U366 , P2_U3056 , P2_R1161_U295 );
nand NAND2_19603 ( P2_R1161_U367 , P2_U3897 , P2_R1161_U295 );
nand NAND3_19604 ( P2_R1161_U368 , P2_R1161_U296 , P2_R1161_U168 , P2_R1161_U301 );
nand NAND3_19605 ( P2_R1161_U369 , P2_R1161_U155 , P2_R1161_U168 , P2_R1161_U133 );
nand NAND2_19606 ( P2_R1161_U370 , P2_R1161_U297 , P2_R1161_U301 );
nand NAND2_19607 ( P2_R1161_U371 , P2_U3082 , P2_R1161_U39 );
nand NAND2_19608 ( P2_R1161_U372 , P2_U3416 , P2_R1161_U38 );
nand NAND2_19609 ( P2_R1161_U373 , P2_R1161_U372 , P2_R1161_U371 );
nand NAND2_19610 ( P2_R1161_U374 , P2_R1161_U352 , P2_R1161_U40 );
nand NAND2_19611 ( P2_R1161_U375 , P2_R1161_U373 , P2_R1161_U206 );
nand NAND2_19612 ( P2_R1161_U376 , P2_U3083 , P2_R1161_U36 );
nand NAND2_19613 ( P2_R1161_U377 , P2_U3413 , P2_R1161_U37 );
nand NAND2_19614 ( P2_R1161_U378 , P2_R1161_U377 , P2_R1161_U376 );
nand NAND2_19615 ( P2_R1161_U379 , P2_R1161_U353 , P2_R1161_U144 );
nand NAND2_19616 ( P2_R1161_U380 , P2_R1161_U203 , P2_R1161_U378 );
nand NAND2_19617 ( P2_R1161_U381 , P2_U3069 , P2_R1161_U23 );
nand NAND2_19618 ( P2_R1161_U382 , P2_U3410 , P2_R1161_U21 );
nand NAND2_19619 ( P2_R1161_U383 , P2_U3070 , P2_R1161_U19 );
nand NAND2_19620 ( P2_R1161_U384 , P2_U3407 , P2_R1161_U20 );
nand NAND2_19621 ( P2_R1161_U385 , P2_R1161_U384 , P2_R1161_U383 );
nand NAND2_19622 ( P2_R1161_U386 , P2_R1161_U354 , P2_R1161_U41 );
nand NAND2_19623 ( P2_R1161_U387 , P2_R1161_U385 , P2_R1161_U195 );
nand NAND2_19624 ( P2_R1161_U388 , P2_U3066 , P2_R1161_U35 );
nand NAND2_19625 ( P2_R1161_U389 , P2_U3404 , P2_R1161_U26 );
nand NAND2_19626 ( P2_R1161_U390 , P2_U3059 , P2_R1161_U24 );
nand NAND2_19627 ( P2_R1161_U391 , P2_U3401 , P2_R1161_U25 );
nand NAND2_19628 ( P2_R1161_U392 , P2_R1161_U391 , P2_R1161_U390 );
nand NAND2_19629 ( P2_R1161_U393 , P2_R1161_U355 , P2_R1161_U44 );
nand NAND2_19630 ( P2_R1161_U394 , P2_R1161_U392 , P2_R1161_U221 );
nand NAND2_19631 ( P2_R1161_U395 , P2_U3063 , P2_R1161_U32 );
nand NAND2_19632 ( P2_R1161_U396 , P2_U3398 , P2_R1161_U33 );
nand NAND2_19633 ( P2_R1161_U397 , P2_R1161_U396 , P2_R1161_U395 );
nand NAND2_19634 ( P2_R1161_U398 , P2_R1161_U356 , P2_R1161_U145 );
nand NAND2_19635 ( P2_R1161_U399 , P2_R1161_U230 , P2_R1161_U397 );
nand NAND2_19636 ( P2_R1161_U400 , P2_U3067 , P2_R1161_U27 );
nand NAND2_19637 ( P2_R1161_U401 , P2_U3395 , P2_R1161_U28 );
nand NAND2_19638 ( P2_R1161_U402 , P2_U3054 , P2_R1161_U147 );
nand NAND2_19639 ( P2_R1161_U403 , P2_U3904 , P2_R1161_U146 );
nand NAND2_19640 ( P2_R1161_U404 , P2_U3054 , P2_R1161_U147 );
nand NAND2_19641 ( P2_R1161_U405 , P2_U3904 , P2_R1161_U146 );
nand NAND2_19642 ( P2_R1161_U406 , P2_R1161_U405 , P2_R1161_U404 );
nand NAND2_19643 ( P2_R1161_U407 , P2_R1161_U148 , P2_R1161_U149 );
nand NAND2_19644 ( P2_R1161_U408 , P2_R1161_U305 , P2_R1161_U406 );
nand NAND2_19645 ( P2_R1161_U409 , P2_U3053 , P2_R1161_U88 );
nand NAND2_19646 ( P2_R1161_U410 , P2_U3895 , P2_R1161_U87 );
nand NAND2_19647 ( P2_R1161_U411 , P2_U3053 , P2_R1161_U88 );
nand NAND2_19648 ( P2_R1161_U412 , P2_U3895 , P2_R1161_U87 );
nand NAND2_19649 ( P2_R1161_U413 , P2_R1161_U412 , P2_R1161_U411 );
nand NAND2_19650 ( P2_R1161_U414 , P2_R1161_U150 , P2_R1161_U151 );
nand NAND2_19651 ( P2_R1161_U415 , P2_R1161_U303 , P2_R1161_U413 );
nand NAND2_19652 ( P2_R1161_U416 , P2_U3052 , P2_R1161_U46 );
nand NAND2_19653 ( P2_R1161_U417 , P2_U3896 , P2_R1161_U47 );
nand NAND2_19654 ( P2_R1161_U418 , P2_U3052 , P2_R1161_U46 );
nand NAND2_19655 ( P2_R1161_U419 , P2_U3896 , P2_R1161_U47 );
nand NAND2_19656 ( P2_R1161_U420 , P2_R1161_U419 , P2_R1161_U418 );
nand NAND2_19657 ( P2_R1161_U421 , P2_R1161_U152 , P2_R1161_U153 );
nand NAND2_19658 ( P2_R1161_U422 , P2_R1161_U300 , P2_R1161_U420 );
nand NAND2_19659 ( P2_R1161_U423 , P2_U3056 , P2_R1161_U49 );
nand NAND2_19660 ( P2_R1161_U424 , P2_U3897 , P2_R1161_U48 );
nand NAND2_19661 ( P2_R1161_U425 , P2_U3057 , P2_R1161_U50 );
nand NAND2_19662 ( P2_R1161_U426 , P2_U3898 , P2_R1161_U51 );
nand NAND2_19663 ( P2_R1161_U427 , P2_R1161_U426 , P2_R1161_U425 );
nand NAND2_19664 ( P2_R1161_U428 , P2_R1161_U357 , P2_R1161_U89 );
nand NAND2_19665 ( P2_R1161_U429 , P2_R1161_U427 , P2_R1161_U307 );
nand NAND2_19666 ( P2_R1161_U430 , P2_U3064 , P2_R1161_U52 );
nand NAND2_19667 ( P2_R1161_U431 , P2_U3899 , P2_R1161_U53 );
nand NAND2_19668 ( P2_R1161_U432 , P2_R1161_U431 , P2_R1161_U430 );
nand NAND2_19669 ( P2_R1161_U433 , P2_R1161_U358 , P2_R1161_U155 );
nand NAND2_19670 ( P2_R1161_U434 , P2_R1161_U294 , P2_R1161_U432 );
nand NAND2_19671 ( P2_R1161_U435 , P2_U3065 , P2_R1161_U84 );
nand NAND2_19672 ( P2_R1161_U436 , P2_U3900 , P2_R1161_U85 );
nand NAND2_19673 ( P2_R1161_U437 , P2_U3065 , P2_R1161_U84 );
nand NAND2_19674 ( P2_R1161_U438 , P2_U3900 , P2_R1161_U85 );
nand NAND2_19675 ( P2_R1161_U439 , P2_R1161_U438 , P2_R1161_U437 );
nand NAND2_19676 ( P2_R1161_U440 , P2_R1161_U156 , P2_R1161_U157 );
nand NAND2_19677 ( P2_R1161_U441 , P2_R1161_U290 , P2_R1161_U439 );
nand NAND2_19678 ( P2_R1161_U442 , P2_U3060 , P2_R1161_U82 );
nand NAND2_19679 ( P2_R1161_U443 , P2_U3901 , P2_R1161_U83 );
nand NAND2_19680 ( P2_R1161_U444 , P2_U3060 , P2_R1161_U82 );
nand NAND2_19681 ( P2_R1161_U445 , P2_U3901 , P2_R1161_U83 );
nand NAND2_19682 ( P2_R1161_U446 , P2_R1161_U445 , P2_R1161_U444 );

endmodule
