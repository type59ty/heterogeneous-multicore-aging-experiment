// b22
// 767 inputs  (32 PIs + 735 PPIs)
// 757 outputs (22 POs + 735 PPOs)
// 29162 gates (24671 gates + 4491 inverters + 0 buffers )
// ( 3092 AND + 716 OR + 20682 NAND + 181 NOR )
// Time: Wed Mar 25 17:47:22 2009
// All copyrigh from NCKU EE TestLAB, Taiwan. [2008.12. WCL]

module b22_ras ( P1_U3355 , P1_U3354 , P1_U3353 , P1_U3352 , P1_U3351 , P1_U3350 ,
             P1_U3349 , P1_U3348 , P1_U3347 , P1_U3346 , P1_U3345 , P1_U3344 ,
             P1_U3343 , P1_U3342 , P1_U3341 , P1_U3340 , P1_U3339 , P1_U3338 ,
             P1_U3337 , P1_U3336 , P1_U3335 , P1_U3334 , P1_U3333 , P1_U3332 ,
             P1_U3331 , P1_U3330 , P1_U3329 , P1_U3328 , P1_U3327 , P1_U3326 ,
             P1_U3325 , P1_U3324 , P1_U3445 , P1_U3446 , P1_U3323 , P1_U3322 ,
             P1_U3321 , P1_U3320 , P1_U3319 , P1_U3318 , P1_U3317 , P1_U3316 ,
             P1_U3315 , P1_U3314 , P1_U3313 , P1_U3312 , P1_U3311 , P1_U3310 ,
             P1_U3309 , P1_U3308 , P1_U3307 , P1_U3306 , P1_U3305 , P1_U3304 ,
             P1_U3303 , P1_U3302 , P1_U3301 , P1_U3300 , P1_U3299 , P1_U3298 ,
             P1_U3297 , P1_U3296 , P1_U3295 , P1_U3294 , P1_U3459 , P1_U3462 ,
             P1_U3465 , P1_U3468 , P1_U3471 , P1_U3474 , P1_U3477 , P1_U3480 ,
             P1_U3483 , P1_U3486 , P1_U3489 , P1_U3492 , P1_U3495 , P1_U3498 ,
             P1_U3501 , P1_U3504 , P1_U3507 , P1_U3510 , P1_U3513 , P1_U3515 ,
             P1_U3516 , P1_U3517 , P1_U3518 , P1_U3519 , P1_U3520 , P1_U3521 ,
             P1_U3522 , P1_U3523 , P1_U3524 , P1_U3525 , P1_U3526 , P1_U3527 ,
             P1_U3528 , P1_U3529 , P1_U3530 , P1_U3531 , P1_U3532 , P1_U3533 ,
             P1_U3534 , P1_U3535 , P1_U3536 , P1_U3537 , P1_U3538 , P1_U3539 ,
             P1_U3540 , P1_U3541 , P1_U3542 , P1_U3543 , P1_U3544 , P1_U3545 ,
             P1_U3546 , P1_U3547 , P1_U3548 , P1_U3549 , P1_U3550 , P1_U3551 ,
             P1_U3552 , P1_U3553 , P1_U3554 , P1_U3555 , P1_U3556 , P1_U3557 ,
             P1_U3558 , P1_U3559 , P1_U3293 , P1_U3292 , P1_U3291 , P1_U3290 ,
             P1_U3289 , P1_U3288 , P1_U3287 , P1_U3286 , P1_U3285 , P1_U3284 ,
             P1_U3283 , P1_U3282 , P1_U3281 , P1_U3280 , P1_U3279 , P1_U3278 ,
             P1_U3277 , P1_U3276 , P1_U3275 , P1_U3274 , P1_U3273 , P1_U3272 ,
             P1_U3271 , P1_U3270 , P1_U3269 , P1_U3268 , P1_U3267 , P1_U3266 ,
             P1_U3265 , P1_U3356 , P1_U3264 , P1_U3263 , P1_U3262 , P1_U3261 ,
             P1_U3260 , P1_U3259 , P1_U3258 , P1_U3257 , P1_U3256 , P1_U3255 ,
             P1_U3254 , P1_U3253 , P1_U3252 , P1_U3251 , P1_U3250 , P1_U3249 ,
             P1_U3248 , P1_U3247 , P1_U3246 , P1_U3245 , P1_U3244 , P1_U3243 ,
             P1_U3560 , P1_U3561 , P1_U3562 , P1_U3563 , P1_U3564 , P1_U3565 ,
             P1_U3566 , P1_U3567 , P1_U3568 , P1_U3569 , P1_U3570 , P1_U3571 ,
             P1_U3572 , P1_U3573 , P1_U3574 , P1_U3575 , P1_U3576 , P1_U3577 ,
             P1_U3578 , P1_U3579 , P1_U3580 , P1_U3581 , P1_U3582 , P1_U3583 ,
             P1_U3584 , P1_U3585 , P1_U3586 , P1_U3587 , P1_U3588 , P1_U3589 ,
             P1_U3590 , P1_U3591 , P1_U3242 , P1_U3241 , P1_U3240 , P1_U3239 ,
             P1_U3238 , P1_U3237 , P1_U3236 , P1_U3235 , P1_U3234 , P1_U3233 ,
             P1_U3232 , P1_U3231 , P1_U3230 , P1_U3229 , P1_U3228 , P1_U3227 ,
             P1_U3226 , P1_U3225 , P1_U3224 , P1_U3223 , P1_U3222 , P1_U3221 ,
             P1_U3220 , P1_U3219 , P1_U3218 , P1_U3217 , P1_U3216 , P1_U3215 ,
             P1_U3214 , P1_U3213 , P1_U3086 , P1_U3085 , P1_U4016 , P2_U3327 ,
             P2_U3326 , P2_U3325 , P2_U3324 , P2_U3323 , P2_U3322 , P2_U3321 ,
             P2_U3320 , P2_U3319 , P2_U3318 , P2_U3317 , P2_U3316 , P2_U3315 ,
             P2_U3314 , P2_U3313 , P2_U3312 , P2_U3311 , P2_U3310 , P2_U3309 ,
             P2_U3308 , P2_U3307 , P2_U3306 , P2_U3305 , P2_U3304 , P2_U3303 ,
             P2_U3302 , P2_U3301 , P2_U3300 , P2_U3299 , P2_U3298 , P2_U3297 ,
             P2_U3296 , P2_U3416 , P2_U3417 , P2_U3295 , P2_U3294 , P2_U3293 ,
             P2_U3292 , P2_U3291 , P2_U3290 , P2_U3289 , P2_U3288 , P2_U3287 ,
             P2_U3286 , P2_U3285 , P2_U3284 , P2_U3283 , P2_U3282 , P2_U3281 ,
             P2_U3280 , P2_U3279 , P2_U3278 , P2_U3277 , P2_U3276 , P2_U3275 ,
             P2_U3274 , P2_U3273 , P2_U3272 , P2_U3271 , P2_U3270 , P2_U3269 ,
             P2_U3268 , P2_U3267 , P2_U3266 , P2_U3430 , P2_U3433 , P2_U3436 ,
             P2_U3439 , P2_U3442 , P2_U3445 , P2_U3448 , P2_U3451 , P2_U3454 ,
             P2_U3457 , P2_U3460 , P2_U3463 , P2_U3466 , P2_U3469 , P2_U3472 ,
             P2_U3475 , P2_U3478 , P2_U3481 , P2_U3484 , P2_U3486 , P2_U3487 ,
             P2_U3488 , P2_U3489 , P2_U3490 , P2_U3491 , P2_U3492 , P2_U3493 ,
             P2_U3494 , P2_U3495 , P2_U3496 , P2_U3497 , P2_U3498 , P2_U3499 ,
             P2_U3500 , P2_U3501 , P2_U3502 , P2_U3503 , P2_U3504 , P2_U3505 ,
             P2_U3506 , P2_U3507 , P2_U3508 , P2_U3509 , P2_U3510 , P2_U3511 ,
             P2_U3512 , P2_U3513 , P2_U3514 , P2_U3515 , P2_U3516 , P2_U3517 ,
             P2_U3518 , P2_U3519 , P2_U3520 , P2_U3521 , P2_U3522 , P2_U3523 ,
             P2_U3524 , P2_U3525 , P2_U3526 , P2_U3527 , P2_U3528 , P2_U3529 ,
             P2_U3530 , P2_U3265 , P2_U3264 , P2_U3263 , P2_U3262 , P2_U3261 ,
             P2_U3260 , P2_U3259 , P2_U3258 , P2_U3257 , P2_U3256 , P2_U3255 ,
             P2_U3254 , P2_U3253 , P2_U3252 , P2_U3251 , P2_U3250 , P2_U3249 ,
             P2_U3248 , P2_U3247 , P2_U3246 , P2_U3245 , P2_U3244 , P2_U3243 ,
             P2_U3242 , P2_U3241 , P2_U3240 , P2_U3239 , P2_U3238 , P2_U3237 ,
             P2_U3236 , P2_U3235 , P2_U3234 , P2_U3233 , P2_U3232 , P2_U3231 ,
             P2_U3230 , P2_U3229 , P2_U3228 , P2_U3227 , P2_U3226 , P2_U3225 ,
             P2_U3224 , P2_U3223 , P2_U3222 , P2_U3221 , P2_U3220 , P2_U3219 ,
             P2_U3218 , P2_U3217 , P2_U3216 , P2_U3215 , P2_U3214 , P2_U3531 ,
             P2_U3532 , P2_U3533 , P2_U3534 , P2_U3535 , P2_U3536 , P2_U3537 ,
             P2_U3538 , P2_U3539 , P2_U3540 , P2_U3541 , P2_U3542 , P2_U3543 ,
             P2_U3544 , P2_U3545 , P2_U3546 , P2_U3547 , P2_U3548 , P2_U3549 ,
             P2_U3550 , P2_U3551 , P2_U3552 , P2_U3553 , P2_U3554 , P2_U3555 ,
             P2_U3556 , P2_U3557 , P2_U3558 , P2_U3559 , P2_U3560 , P2_U3561 ,
             P2_U3562 , P2_U3328 , P2_U3213 , P2_U3212 , P2_U3211 , P2_U3210 ,
             P2_U3209 , P2_U3208 , P2_U3207 , P2_U3206 , P2_U3205 , P2_U3204 ,
             P2_U3203 , P2_U3202 , P2_U3201 , P2_U3200 , P2_U3199 , P2_U3198 ,
             P2_U3197 , P2_U3196 , P2_U3195 , P2_U3194 , P2_U3193 , P2_U3192 ,
             P2_U3191 , P2_U3190 , P2_U3189 , P2_U3188 , P2_U3187 , P2_U3186 ,
             P2_U3185 , P2_U3088 , P2_U3087 , P2_U3947 , P3_U3295 , P3_U3294 ,
             P3_U3293 , P3_U3292 , P3_U3291 , P3_U3290 , P3_U3289 , P3_U3288 ,
             P3_U3287 , P3_U3286 , P3_U3285 , P3_U3284 , P3_U3283 , P3_U3282 ,
             P3_U3281 , P3_U3280 , P3_U3279 , P3_U3278 , P3_U3277 , P3_U3276 ,
             P3_U3275 , P3_U3274 , P3_U3273 , P3_U3272 , P3_U3271 , P3_U3270 ,
             P3_U3269 , P3_U3268 , P3_U3267 , P3_U3266 , P3_U3265 , P3_U3264 ,
             P3_U3376 , P3_U3377 , P3_U3263 , P3_U3262 , P3_U3261 , P3_U3260 ,
             P3_U3259 , P3_U3258 , P3_U3257 , P3_U3256 , P3_U3255 , P3_U3254 ,
             P3_U3253 , P3_U3252 , P3_U3251 , P3_U3250 , P3_U3249 , P3_U3248 ,
             P3_U3247 , P3_U3246 , P3_U3245 , P3_U3244 , P3_U3243 , P3_U3242 ,
             P3_U3241 , P3_U3240 , P3_U3239 , P3_U3238 , P3_U3237 , P3_U3236 ,
             P3_U3235 , P3_U3234 , P3_U3390 , P3_U3393 , P3_U3396 , P3_U3399 ,
             P3_U3402 , P3_U3405 , P3_U3408 , P3_U3411 , P3_U3414 , P3_U3417 ,
             P3_U3420 , P3_U3423 , P3_U3426 , P3_U3429 , P3_U3432 , P3_U3435 ,
             P3_U3438 , P3_U3441 , P3_U3444 , P3_U3446 , P3_U3447 , P3_U3448 ,
             P3_U3449 , P3_U3450 , P3_U3451 , P3_U3452 , P3_U3453 , P3_U3454 ,
             P3_U3455 , P3_U3456 , P3_U3457 , P3_U3458 , P3_U3459 , P3_U3460 ,
             P3_U3461 , P3_U3462 , P3_U3463 , P3_U3464 , P3_U3465 , P3_U3466 ,
             P3_U3467 , P3_U3468 , P3_U3469 , P3_U3470 , P3_U3471 , P3_U3472 ,
             P3_U3473 , P3_U3474 , P3_U3475 , P3_U3476 , P3_U3477 , P3_U3478 ,
             P3_U3479 , P3_U3480 , P3_U3481 , P3_U3482 , P3_U3483 , P3_U3484 ,
             P3_U3485 , P3_U3486 , P3_U3487 , P3_U3488 , P3_U3489 , P3_U3490 ,
             P3_U3233 , P3_U3232 , P3_U3231 , P3_U3230 , P3_U3229 , P3_U3228 ,
             P3_U3227 , P3_U3226 , P3_U3225 , P3_U3224 , P3_U3223 , P3_U3222 ,
             P3_U3221 , P3_U3220 , P3_U3219 , P3_U3218 , P3_U3217 , P3_U3216 ,
             P3_U3215 , P3_U3214 , P3_U3213 , P3_U3212 , P3_U3211 , P3_U3210 ,
             P3_U3209 , P3_U3208 , P3_U3207 , P3_U3206 , P3_U3205 , P3_U3204 ,
             P3_U3203 , P3_U3202 , P3_U3201 , P3_U3200 , P3_U3199 , P3_U3198 ,
             P3_U3197 , P3_U3196 , P3_U3195 , P3_U3194 , P3_U3193 , P3_U3192 ,
             P3_U3191 , P3_U3190 , P3_U3189 , P3_U3188 , P3_U3187 , P3_U3186 ,
             P3_U3185 , P3_U3184 , P3_U3183 , P3_U3182 , P3_U3491 , P3_U3492 ,
             P3_U3493 , P3_U3494 , P3_U3495 , P3_U3496 , P3_U3497 , P3_U3498 ,
             P3_U3499 , P3_U3500 , P3_U3501 , P3_U3502 , P3_U3503 , P3_U3504 ,
             P3_U3505 , P3_U3506 , P3_U3507 , P3_U3508 , P3_U3509 , P3_U3510 ,
             P3_U3511 , P3_U3512 , P3_U3513 , P3_U3514 , P3_U3515 , P3_U3516 ,
             P3_U3517 , P3_U3518 , P3_U3519 , P3_U3520 , P3_U3521 , P3_U3522 ,
             P3_U3296 , P3_U3181 , P3_U3180 , P3_U3179 , P3_U3178 , P3_U3177 ,
             P3_U3176 , P3_U3175 , P3_U3174 , P3_U3173 , P3_U3172 , P3_U3171 ,
             P3_U3170 , P3_U3169 , P3_U3168 , P3_U3167 , P3_U3166 , P3_U3165 ,
             P3_U3164 , P3_U3163 , P3_U3162 , P3_U3161 , P3_U3160 , P3_U3159 ,
             P3_U3158 , P3_U3157 , P3_U3156 , P3_U3155 , P3_U3154 , P3_U3153 ,
             P3_U3151 , P3_U3150 , P3_U3897 , SUB_1596_U4 , SUB_1596_U62 , SUB_1596_U63 ,
             SUB_1596_U64 , SUB_1596_U65 , SUB_1596_U66 , SUB_1596_U67 , SUB_1596_U68 , SUB_1596_U69 ,
             SUB_1596_U70 , SUB_1596_U54 , SUB_1596_U55 , SUB_1596_U56 , SUB_1596_U57 , SUB_1596_U58 ,
             SUB_1596_U59 , SUB_1596_U60 , SUB_1596_U61 , SUB_1596_U5 , SUB_1596_U53 , U29 ,
             U28 ,
             P1_IR_REG_0_ , P1_IR_REG_1_ , P1_IR_REG_2_ , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ ,
             P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_10_ , P1_IR_REG_11_ ,
             P1_IR_REG_12_ , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_ ,
             P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_20_ , P1_IR_REG_21_ , P1_IR_REG_22_ , P1_IR_REG_23_ ,
             P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ , P1_IR_REG_27_ , P1_IR_REG_28_ , P1_IR_REG_29_ ,
             P1_IR_REG_30_ , P1_IR_REG_31_ , P1_D_REG_0_ , P1_D_REG_1_ , P1_D_REG_2_ , P1_D_REG_3_ ,
             P1_D_REG_4_ , P1_D_REG_5_ , P1_D_REG_6_ , P1_D_REG_7_ , P1_D_REG_8_ , P1_D_REG_9_ ,
             P1_D_REG_10_ , P1_D_REG_11_ , P1_D_REG_12_ , P1_D_REG_13_ , P1_D_REG_14_ , P1_D_REG_15_ ,
             P1_D_REG_16_ , P1_D_REG_17_ , P1_D_REG_18_ , P1_D_REG_19_ , P1_D_REG_20_ , P1_D_REG_21_ ,
             P1_D_REG_22_ , P1_D_REG_23_ , P1_D_REG_24_ , P1_D_REG_25_ , P1_D_REG_26_ , P1_D_REG_27_ ,
             P1_D_REG_28_ , P1_D_REG_29_ , P1_D_REG_30_ , P1_D_REG_31_ , P1_REG0_REG_0_ , P1_REG0_REG_1_ ,
             P1_REG0_REG_2_ , P1_REG0_REG_3_ , P1_REG0_REG_4_ , P1_REG0_REG_5_ , P1_REG0_REG_6_ , P1_REG0_REG_7_ ,
             P1_REG0_REG_8_ , P1_REG0_REG_9_ , P1_REG0_REG_10_ , P1_REG0_REG_11_ , P1_REG0_REG_12_ , P1_REG0_REG_13_ ,
             P1_REG0_REG_14_ , P1_REG0_REG_15_ , P1_REG0_REG_16_ , P1_REG0_REG_17_ , P1_REG0_REG_18_ , P1_REG0_REG_19_ ,
             P1_REG0_REG_20_ , P1_REG0_REG_21_ , P1_REG0_REG_22_ , P1_REG0_REG_23_ , P1_REG0_REG_24_ , P1_REG0_REG_25_ ,
             P1_REG0_REG_26_ , P1_REG0_REG_27_ , P1_REG0_REG_28_ , P1_REG0_REG_29_ , P1_REG0_REG_30_ , P1_REG0_REG_31_ ,
             P1_REG1_REG_0_ , P1_REG1_REG_1_ , P1_REG1_REG_2_ , P1_REG1_REG_3_ , P1_REG1_REG_4_ , P1_REG1_REG_5_ ,
             P1_REG1_REG_6_ , P1_REG1_REG_7_ , P1_REG1_REG_8_ , P1_REG1_REG_9_ , P1_REG1_REG_10_ , P1_REG1_REG_11_ ,
             P1_REG1_REG_12_ , P1_REG1_REG_13_ , P1_REG1_REG_14_ , P1_REG1_REG_15_ , P1_REG1_REG_16_ , P1_REG1_REG_17_ ,
             P1_REG1_REG_18_ , P1_REG1_REG_19_ , P1_REG1_REG_20_ , P1_REG1_REG_21_ , P1_REG1_REG_22_ , P1_REG1_REG_23_ ,
             P1_REG1_REG_24_ , P1_REG1_REG_25_ , P1_REG1_REG_26_ , P1_REG1_REG_27_ , P1_REG1_REG_28_ , P1_REG1_REG_29_ ,
             P1_REG1_REG_30_ , P1_REG1_REG_31_ , P1_REG2_REG_0_ , P1_REG2_REG_1_ , P1_REG2_REG_2_ , P1_REG2_REG_3_ ,
             P1_REG2_REG_4_ , P1_REG2_REG_5_ , P1_REG2_REG_6_ , P1_REG2_REG_7_ , P1_REG2_REG_8_ , P1_REG2_REG_9_ ,
             P1_REG2_REG_10_ , P1_REG2_REG_11_ , P1_REG2_REG_12_ , P1_REG2_REG_13_ , P1_REG2_REG_14_ , P1_REG2_REG_15_ ,
             P1_REG2_REG_16_ , P1_REG2_REG_17_ , P1_REG2_REG_18_ , P1_REG2_REG_19_ , P1_REG2_REG_20_ , P1_REG2_REG_21_ ,
             P1_REG2_REG_22_ , P1_REG2_REG_23_ , P1_REG2_REG_24_ , P1_REG2_REG_25_ , P1_REG2_REG_26_ , P1_REG2_REG_27_ ,
             P1_REG2_REG_28_ , P1_REG2_REG_29_ , P1_REG2_REG_30_ , P1_REG2_REG_31_ , P1_ADDR_REG_19_ , P1_ADDR_REG_18_ ,
             P1_ADDR_REG_17_ , P1_ADDR_REG_16_ , P1_ADDR_REG_15_ , P1_ADDR_REG_14_ , P1_ADDR_REG_13_ , P1_ADDR_REG_12_ ,
             P1_ADDR_REG_11_ , P1_ADDR_REG_10_ , P1_ADDR_REG_9_ , P1_ADDR_REG_8_ , P1_ADDR_REG_7_ , P1_ADDR_REG_6_ ,
             P1_ADDR_REG_5_ , P1_ADDR_REG_4_ , P1_ADDR_REG_3_ , P1_ADDR_REG_2_ , P1_ADDR_REG_1_ , P1_ADDR_REG_0_ ,
             P1_DATAO_REG_0_ , P1_DATAO_REG_1_ , P1_DATAO_REG_2_ , P1_DATAO_REG_3_ , P1_DATAO_REG_4_ , P1_DATAO_REG_5_ ,
             P1_DATAO_REG_6_ , P1_DATAO_REG_7_ , P1_DATAO_REG_8_ , P1_DATAO_REG_9_ , P1_DATAO_REG_10_ , P1_DATAO_REG_11_ ,
             P1_DATAO_REG_12_ , P1_DATAO_REG_13_ , P1_DATAO_REG_14_ , P1_DATAO_REG_15_ , P1_DATAO_REG_16_ , P1_DATAO_REG_17_ ,
             P1_DATAO_REG_18_ , P1_DATAO_REG_19_ , P1_DATAO_REG_20_ , P1_DATAO_REG_21_ , P1_DATAO_REG_22_ , P1_DATAO_REG_23_ ,
             P1_DATAO_REG_24_ , P1_DATAO_REG_25_ , P1_DATAO_REG_26_ , P1_DATAO_REG_27_ , P1_DATAO_REG_28_ , P1_DATAO_REG_29_ ,
             P1_DATAO_REG_30_ , P1_DATAO_REG_31_ , P1_B_REG , P1_REG3_REG_15_ , P1_REG3_REG_26_ , P1_REG3_REG_6_ ,
             P1_REG3_REG_18_ , P1_REG3_REG_2_ , P1_REG3_REG_11_ , P1_REG3_REG_22_ , P1_REG3_REG_13_ , P1_REG3_REG_20_ ,
             P1_REG3_REG_0_ , P1_REG3_REG_9_ , P1_REG3_REG_4_ , P1_REG3_REG_24_ , P1_REG3_REG_17_ , P1_REG3_REG_5_ ,
             P1_REG3_REG_16_ , P1_REG3_REG_25_ , P1_REG3_REG_12_ , P1_REG3_REG_21_ , P1_REG3_REG_1_ , P1_REG3_REG_8_ ,
             P1_REG3_REG_28_ , P1_REG3_REG_19_ , P1_REG3_REG_3_ , P1_REG3_REG_10_ , P1_REG3_REG_23_ , P1_REG3_REG_14_ ,
             P1_REG3_REG_27_ , P1_REG3_REG_7_ , P1_STATE_REG , P1_RD_REG , P1_WR_REG , P2_IR_REG_0_ ,
             P2_IR_REG_1_ , P2_IR_REG_2_ , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ , P2_IR_REG_6_ ,
             P2_IR_REG_7_ , P2_IR_REG_8_ , P2_IR_REG_9_ , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_ ,
             P2_IR_REG_13_ , P2_IR_REG_14_ , P2_IR_REG_15_ , P2_IR_REG_16_ , P2_IR_REG_17_ , P2_IR_REG_18_ ,
             P2_IR_REG_19_ , P2_IR_REG_20_ , P2_IR_REG_21_ , P2_IR_REG_22_ , P2_IR_REG_23_ , P2_IR_REG_24_ ,
             P2_IR_REG_25_ , P2_IR_REG_26_ , P2_IR_REG_27_ , P2_IR_REG_28_ , P2_IR_REG_29_ , P2_IR_REG_30_ ,
             P2_IR_REG_31_ , P2_D_REG_0_ , P2_D_REG_1_ , P2_D_REG_2_ , P2_D_REG_3_ , P2_D_REG_4_ ,
             P2_D_REG_5_ , P2_D_REG_6_ , P2_D_REG_7_ , P2_D_REG_8_ , P2_D_REG_9_ , P2_D_REG_10_ ,
             P2_D_REG_11_ , P2_D_REG_12_ , P2_D_REG_13_ , P2_D_REG_14_ , P2_D_REG_15_ , P2_D_REG_16_ ,
             P2_D_REG_17_ , P2_D_REG_18_ , P2_D_REG_19_ , P2_D_REG_20_ , P2_D_REG_21_ , P2_D_REG_22_ ,
             P2_D_REG_23_ , P2_D_REG_24_ , P2_D_REG_25_ , P2_D_REG_26_ , P2_D_REG_27_ , P2_D_REG_28_ ,
             P2_D_REG_29_ , P2_D_REG_30_ , P2_D_REG_31_ , P2_REG0_REG_0_ , P2_REG0_REG_1_ , P2_REG0_REG_2_ ,
             P2_REG0_REG_3_ , P2_REG0_REG_4_ , P2_REG0_REG_5_ , P2_REG0_REG_6_ , P2_REG0_REG_7_ , P2_REG0_REG_8_ ,
             P2_REG0_REG_9_ , P2_REG0_REG_10_ , P2_REG0_REG_11_ , P2_REG0_REG_12_ , P2_REG0_REG_13_ , P2_REG0_REG_14_ ,
             P2_REG0_REG_15_ , P2_REG0_REG_16_ , P2_REG0_REG_17_ , P2_REG0_REG_18_ , P2_REG0_REG_19_ , P2_REG0_REG_20_ ,
             P2_REG0_REG_21_ , P2_REG0_REG_22_ , P2_REG0_REG_23_ , P2_REG0_REG_24_ , P2_REG0_REG_25_ , P2_REG0_REG_26_ ,
             P2_REG0_REG_27_ , P2_REG0_REG_28_ , P2_REG0_REG_29_ , P2_REG0_REG_30_ , P2_REG0_REG_31_ , P2_REG1_REG_0_ ,
             P2_REG1_REG_1_ , P2_REG1_REG_2_ , P2_REG1_REG_3_ , P2_REG1_REG_4_ , P2_REG1_REG_5_ , P2_REG1_REG_6_ ,
             P2_REG1_REG_7_ , P2_REG1_REG_8_ , P2_REG1_REG_9_ , P2_REG1_REG_10_ , P2_REG1_REG_11_ , P2_REG1_REG_12_ ,
             P2_REG1_REG_13_ , P2_REG1_REG_14_ , P2_REG1_REG_15_ , P2_REG1_REG_16_ , P2_REG1_REG_17_ , P2_REG1_REG_18_ ,
             P2_REG1_REG_19_ , P2_REG1_REG_20_ , P2_REG1_REG_21_ , P2_REG1_REG_22_ , P2_REG1_REG_23_ , P2_REG1_REG_24_ ,
             P2_REG1_REG_25_ , P2_REG1_REG_26_ , P2_REG1_REG_27_ , P2_REG1_REG_28_ , P2_REG1_REG_29_ , P2_REG1_REG_30_ ,
             P2_REG1_REG_31_ , P2_REG2_REG_0_ , P2_REG2_REG_1_ , P2_REG2_REG_2_ , P2_REG2_REG_3_ , P2_REG2_REG_4_ ,
             P2_REG2_REG_5_ , P2_REG2_REG_6_ , P2_REG2_REG_7_ , P2_REG2_REG_8_ , P2_REG2_REG_9_ , P2_REG2_REG_10_ ,
             P2_REG2_REG_11_ , P2_REG2_REG_12_ , P2_REG2_REG_13_ , P2_REG2_REG_14_ , P2_REG2_REG_15_ , P2_REG2_REG_16_ ,
             P2_REG2_REG_17_ , P2_REG2_REG_18_ , P2_REG2_REG_19_ , P2_REG2_REG_20_ , P2_REG2_REG_21_ , P2_REG2_REG_22_ ,
             P2_REG2_REG_23_ , P2_REG2_REG_24_ , P2_REG2_REG_25_ , P2_REG2_REG_26_ , P2_REG2_REG_27_ , P2_REG2_REG_28_ ,
             P2_REG2_REG_29_ , P2_REG2_REG_30_ , P2_REG2_REG_31_ , P2_ADDR_REG_19_ , P2_ADDR_REG_18_ , P2_ADDR_REG_17_ ,
             P2_ADDR_REG_16_ , P2_ADDR_REG_15_ , P2_ADDR_REG_14_ , P2_ADDR_REG_13_ , P2_ADDR_REG_12_ , P2_ADDR_REG_11_ ,
             P2_ADDR_REG_10_ , P2_ADDR_REG_9_ , P2_ADDR_REG_8_ , P2_ADDR_REG_7_ , P2_ADDR_REG_6_ , P2_ADDR_REG_5_ ,
             P2_ADDR_REG_4_ , P2_ADDR_REG_3_ , P2_ADDR_REG_2_ , P2_ADDR_REG_1_ , P2_ADDR_REG_0_ , P2_DATAO_REG_0_ ,
             P2_DATAO_REG_1_ , P2_DATAO_REG_2_ , P2_DATAO_REG_3_ , P2_DATAO_REG_4_ , P2_DATAO_REG_5_ , P2_DATAO_REG_6_ ,
             P2_DATAO_REG_7_ , P2_DATAO_REG_8_ , P2_DATAO_REG_9_ , P2_DATAO_REG_10_ , P2_DATAO_REG_11_ , P2_DATAO_REG_12_ ,
             P2_DATAO_REG_13_ , P2_DATAO_REG_14_ , P2_DATAO_REG_15_ , P2_DATAO_REG_16_ , P2_DATAO_REG_17_ , P2_DATAO_REG_18_ ,
             P2_DATAO_REG_19_ , P2_DATAO_REG_20_ , P2_DATAO_REG_21_ , P2_DATAO_REG_22_ , P2_DATAO_REG_23_ , P2_DATAO_REG_24_ ,
             P2_DATAO_REG_25_ , P2_DATAO_REG_26_ , P2_DATAO_REG_27_ , P2_DATAO_REG_28_ , P2_DATAO_REG_29_ , P2_DATAO_REG_30_ ,
             P2_DATAO_REG_31_ , P2_B_REG , P2_REG3_REG_15_ , P2_REG3_REG_26_ , P2_REG3_REG_6_ , P2_REG3_REG_18_ ,
             P2_REG3_REG_2_ , P2_REG3_REG_11_ , P2_REG3_REG_22_ , P2_REG3_REG_13_ , P2_REG3_REG_20_ , P2_REG3_REG_0_ ,
             P2_REG3_REG_9_ , P2_REG3_REG_4_ , P2_REG3_REG_24_ , P2_REG3_REG_17_ , P2_REG3_REG_5_ , P2_REG3_REG_16_ ,
             P2_REG3_REG_25_ , P2_REG3_REG_12_ , P2_REG3_REG_21_ , P2_REG3_REG_1_ , P2_REG3_REG_8_ , P2_REG3_REG_28_ ,
             P2_REG3_REG_19_ , P2_REG3_REG_3_ , P2_REG3_REG_10_ , P2_REG3_REG_23_ , P2_REG3_REG_14_ , P2_REG3_REG_27_ ,
             P2_REG3_REG_7_ , P2_STATE_REG , P2_RD_REG , P2_WR_REG , P3_IR_REG_0_ , P3_IR_REG_1_ ,
             P3_IR_REG_2_ , P3_IR_REG_3_ , P3_IR_REG_4_ , P3_IR_REG_5_ , P3_IR_REG_6_ , P3_IR_REG_7_ ,
             P3_IR_REG_8_ , P3_IR_REG_9_ , P3_IR_REG_10_ , P3_IR_REG_11_ , P3_IR_REG_12_ , P3_IR_REG_13_ ,
             P3_IR_REG_14_ , P3_IR_REG_15_ , P3_IR_REG_16_ , P3_IR_REG_17_ , P3_IR_REG_18_ , P3_IR_REG_19_ ,
             P3_IR_REG_20_ , P3_IR_REG_21_ , P3_IR_REG_22_ , P3_IR_REG_23_ , P3_IR_REG_24_ , P3_IR_REG_25_ ,
             P3_IR_REG_26_ , P3_IR_REG_27_ , P3_IR_REG_28_ , P3_IR_REG_29_ , P3_IR_REG_30_ , P3_IR_REG_31_ ,
             P3_D_REG_0_ , P3_D_REG_1_ , P3_D_REG_2_ , P3_D_REG_3_ , P3_D_REG_4_ , P3_D_REG_5_ ,
             P3_D_REG_6_ , P3_D_REG_7_ , P3_D_REG_8_ , P3_D_REG_9_ , P3_D_REG_10_ , P3_D_REG_11_ ,
             P3_D_REG_12_ , P3_D_REG_13_ , P3_D_REG_14_ , P3_D_REG_15_ , P3_D_REG_16_ , P3_D_REG_17_ ,
             P3_D_REG_18_ , P3_D_REG_19_ , P3_D_REG_20_ , P3_D_REG_21_ , P3_D_REG_22_ , P3_D_REG_23_ ,
             P3_D_REG_24_ , P3_D_REG_25_ , P3_D_REG_26_ , P3_D_REG_27_ , P3_D_REG_28_ , P3_D_REG_29_ ,
             P3_D_REG_30_ , P3_D_REG_31_ , P3_REG0_REG_0_ , P3_REG0_REG_1_ , P3_REG0_REG_2_ , P3_REG0_REG_3_ ,
             P3_REG0_REG_4_ , P3_REG0_REG_5_ , P3_REG0_REG_6_ , P3_REG0_REG_7_ , P3_REG0_REG_8_ , P3_REG0_REG_9_ ,
             P3_REG0_REG_10_ , P3_REG0_REG_11_ , P3_REG0_REG_12_ , P3_REG0_REG_13_ , P3_REG0_REG_14_ , P3_REG0_REG_15_ ,
             P3_REG0_REG_16_ , P3_REG0_REG_17_ , P3_REG0_REG_18_ , P3_REG0_REG_19_ , P3_REG0_REG_20_ , P3_REG0_REG_21_ ,
             P3_REG0_REG_22_ , P3_REG0_REG_23_ , P3_REG0_REG_24_ , P3_REG0_REG_25_ , P3_REG0_REG_26_ , P3_REG0_REG_27_ ,
             P3_REG0_REG_28_ , P3_REG0_REG_29_ , P3_REG0_REG_30_ , P3_REG0_REG_31_ , P3_REG1_REG_0_ , P3_REG1_REG_1_ ,
             P3_REG1_REG_2_ , P3_REG1_REG_3_ , P3_REG1_REG_4_ , P3_REG1_REG_5_ , P3_REG1_REG_6_ , P3_REG1_REG_7_ ,
             P3_REG1_REG_8_ , P3_REG1_REG_9_ , P3_REG1_REG_10_ , P3_REG1_REG_11_ , P3_REG1_REG_12_ , P3_REG1_REG_13_ ,
             P3_REG1_REG_14_ , P3_REG1_REG_15_ , P3_REG1_REG_16_ , P3_REG1_REG_17_ , P3_REG1_REG_18_ , P3_REG1_REG_19_ ,
             P3_REG1_REG_20_ , P3_REG1_REG_21_ , P3_REG1_REG_22_ , P3_REG1_REG_23_ , P3_REG1_REG_24_ , P3_REG1_REG_25_ ,
             P3_REG1_REG_26_ , P3_REG1_REG_27_ , P3_REG1_REG_28_ , P3_REG1_REG_29_ , P3_REG1_REG_30_ , P3_REG1_REG_31_ ,
             P3_REG2_REG_0_ , P3_REG2_REG_1_ , P3_REG2_REG_2_ , P3_REG2_REG_3_ , P3_REG2_REG_4_ , P3_REG2_REG_5_ ,
             P3_REG2_REG_6_ , P3_REG2_REG_7_ , P3_REG2_REG_8_ , P3_REG2_REG_9_ , P3_REG2_REG_10_ , P3_REG2_REG_11_ ,
             P3_REG2_REG_12_ , P3_REG2_REG_13_ , P3_REG2_REG_14_ , P3_REG2_REG_15_ , P3_REG2_REG_16_ , P3_REG2_REG_17_ ,
             P3_REG2_REG_18_ , P3_REG2_REG_19_ , P3_REG2_REG_20_ , P3_REG2_REG_21_ , P3_REG2_REG_22_ , P3_REG2_REG_23_ ,
             P3_REG2_REG_24_ , P3_REG2_REG_25_ , P3_REG2_REG_26_ , P3_REG2_REG_27_ , P3_REG2_REG_28_ , P3_REG2_REG_29_ ,
             P3_REG2_REG_30_ , P3_REG2_REG_31_ , P3_ADDR_REG_19_ , P3_ADDR_REG_18_ , P3_ADDR_REG_17_ , P3_ADDR_REG_16_ ,
             P3_ADDR_REG_15_ , P3_ADDR_REG_14_ , P3_ADDR_REG_13_ , P3_ADDR_REG_12_ , P3_ADDR_REG_11_ , P3_ADDR_REG_10_ ,
             P3_ADDR_REG_9_ , P3_ADDR_REG_8_ , P3_ADDR_REG_7_ , P3_ADDR_REG_6_ , P3_ADDR_REG_5_ , P3_ADDR_REG_4_ ,
             P3_ADDR_REG_3_ , P3_ADDR_REG_2_ , P3_ADDR_REG_1_ , P3_ADDR_REG_0_ , P3_DATAO_REG_0_ , P3_DATAO_REG_1_ ,
             P3_DATAO_REG_2_ , P3_DATAO_REG_3_ , P3_DATAO_REG_4_ , P3_DATAO_REG_5_ , P3_DATAO_REG_6_ , P3_DATAO_REG_7_ ,
             P3_DATAO_REG_8_ , P3_DATAO_REG_9_ , P3_DATAO_REG_10_ , P3_DATAO_REG_11_ , P3_DATAO_REG_12_ , P3_DATAO_REG_13_ ,
             P3_DATAO_REG_14_ , P3_DATAO_REG_15_ , P3_DATAO_REG_16_ , P3_DATAO_REG_17_ , P3_DATAO_REG_18_ , P3_DATAO_REG_19_ ,
             P3_DATAO_REG_20_ , P3_DATAO_REG_21_ , P3_DATAO_REG_22_ , P3_DATAO_REG_23_ , P3_DATAO_REG_24_ , P3_DATAO_REG_25_ ,
             P3_DATAO_REG_26_ , P3_DATAO_REG_27_ , P3_DATAO_REG_28_ , P3_DATAO_REG_29_ , P3_DATAO_REG_30_ , P3_DATAO_REG_31_ ,
             P3_B_REG , P3_REG3_REG_15_ , P3_REG3_REG_26_ , P3_REG3_REG_6_ , P3_REG3_REG_18_ , P3_REG3_REG_2_ ,
             P3_REG3_REG_11_ , P3_REG3_REG_22_ , P3_REG3_REG_13_ , P3_REG3_REG_20_ , P3_REG3_REG_0_ , P3_REG3_REG_9_ ,
             P3_REG3_REG_4_ , P3_REG3_REG_24_ , P3_REG3_REG_17_ , P3_REG3_REG_5_ , P3_REG3_REG_16_ , P3_REG3_REG_25_ ,
             P3_REG3_REG_12_ , P3_REG3_REG_21_ , P3_REG3_REG_1_ , P3_REG3_REG_8_ , P3_REG3_REG_28_ , P3_REG3_REG_19_ ,
             P3_REG3_REG_3_ , P3_REG3_REG_10_ , P3_REG3_REG_23_ , P3_REG3_REG_14_ , P3_REG3_REG_27_ , P3_REG3_REG_7_ ,
             P3_STATE_REG , P3_RD_REG , P3_WR_REG , SI_31_ , SI_30_ , SI_29_ ,
             SI_28_ , SI_27_ , SI_26_ , SI_25_ , SI_24_ , SI_23_ ,
             SI_22_ , SI_21_ , SI_20_ , SI_19_ , SI_18_ , SI_17_ ,
             SI_16_ , SI_15_ , SI_14_ , SI_13_ , SI_12_ , SI_11_ ,
             SI_10_ , SI_9_ , SI_8_ , SI_7_ , SI_6_ , SI_5_ ,
             SI_4_ , SI_3_ , SI_2_ , SI_1_ , SI_0_ );

output SUB_1596_U4 , SUB_1596_U62 , SUB_1596_U63 , SUB_1596_U64 , SUB_1596_U65 , SUB_1596_U66;
output SUB_1596_U67 , SUB_1596_U68 , SUB_1596_U69 , SUB_1596_U70 , SUB_1596_U54 , SUB_1596_U55;
output SUB_1596_U56 , SUB_1596_U57 , SUB_1596_U58 , SUB_1596_U59 , SUB_1596_U60 , SUB_1596_U61;
output SUB_1596_U5 , SUB_1596_U53 , U29 , U28;
output P1_U3355 , P1_U3354 , P1_U3353 , P1_U3352 , P1_U3351 , P1_U3350 , P1_U3349;
output P1_U3348 , P1_U3347 , P1_U3346 , P1_U3345 , P1_U3344 , P1_U3343 , P1_U3342;
output P1_U3341 , P1_U3340 , P1_U3339 , P1_U3338 , P1_U3337 , P1_U3336 , P1_U3335;
output P1_U3334 , P1_U3333 , P1_U3332 , P1_U3331 , P1_U3330 , P1_U3329 , P1_U3328;
output P1_U3327 , P1_U3326 , P1_U3325 , P1_U3324 , P1_U3445 , P1_U3446 , P1_U3323;
output P1_U3322 , P1_U3321 , P1_U3320 , P1_U3319 , P1_U3318 , P1_U3317 , P1_U3316;
output P1_U3315 , P1_U3314 , P1_U3313 , P1_U3312 , P1_U3311 , P1_U3310 , P1_U3309;
output P1_U3308 , P1_U3307 , P1_U3306 , P1_U3305 , P1_U3304 , P1_U3303 , P1_U3302;
output P1_U3301 , P1_U3300 , P1_U3299 , P1_U3298 , P1_U3297 , P1_U3296 , P1_U3295;
output P1_U3294 , P1_U3459 , P1_U3462 , P1_U3465 , P1_U3468 , P1_U3471 , P1_U3474;
output P1_U3477 , P1_U3480 , P1_U3483 , P1_U3486 , P1_U3489 , P1_U3492 , P1_U3495;
output P1_U3498 , P1_U3501 , P1_U3504 , P1_U3507 , P1_U3510 , P1_U3513 , P1_U3515;
output P1_U3516 , P1_U3517 , P1_U3518 , P1_U3519 , P1_U3520 , P1_U3521 , P1_U3522;
output P1_U3523 , P1_U3524 , P1_U3525 , P1_U3526 , P1_U3527 , P1_U3528 , P1_U3529;
output P1_U3530 , P1_U3531 , P1_U3532 , P1_U3533 , P1_U3534 , P1_U3535 , P1_U3536;
output P1_U3537 , P1_U3538 , P1_U3539 , P1_U3540 , P1_U3541 , P1_U3542 , P1_U3543;
output P1_U3544 , P1_U3545 , P1_U3546 , P1_U3547 , P1_U3548 , P1_U3549 , P1_U3550;
output P1_U3551 , P1_U3552 , P1_U3553 , P1_U3554 , P1_U3555 , P1_U3556 , P1_U3557;
output P1_U3558 , P1_U3559 , P1_U3293 , P1_U3292 , P1_U3291 , P1_U3290 , P1_U3289;
output P1_U3288 , P1_U3287 , P1_U3286 , P1_U3285 , P1_U3284 , P1_U3283 , P1_U3282;
output P1_U3281 , P1_U3280 , P1_U3279 , P1_U3278 , P1_U3277 , P1_U3276 , P1_U3275;
output P1_U3274 , P1_U3273 , P1_U3272 , P1_U3271 , P1_U3270 , P1_U3269 , P1_U3268;
output P1_U3267 , P1_U3266 , P1_U3265 , P1_U3356 , P1_U3264 , P1_U3263 , P1_U3262;
output P1_U3261 , P1_U3260 , P1_U3259 , P1_U3258 , P1_U3257 , P1_U3256 , P1_U3255;
output P1_U3254 , P1_U3253 , P1_U3252 , P1_U3251 , P1_U3250 , P1_U3249 , P1_U3248;
output P1_U3247 , P1_U3246 , P1_U3245 , P1_U3244 , P1_U3243 , P1_U3560 , P1_U3561;
output P1_U3562 , P1_U3563 , P1_U3564 , P1_U3565 , P1_U3566 , P1_U3567 , P1_U3568;
output P1_U3569 , P1_U3570 , P1_U3571 , P1_U3572 , P1_U3573 , P1_U3574 , P1_U3575;
output P1_U3576 , P1_U3577 , P1_U3578 , P1_U3579 , P1_U3580 , P1_U3581 , P1_U3582;
output P1_U3583 , P1_U3584 , P1_U3585 , P1_U3586 , P1_U3587 , P1_U3588 , P1_U3589;
output P1_U3590 , P1_U3591 , P1_U3242 , P1_U3241 , P1_U3240 , P1_U3239 , P1_U3238;
output P1_U3237 , P1_U3236 , P1_U3235 , P1_U3234 , P1_U3233 , P1_U3232 , P1_U3231;
output P1_U3230 , P1_U3229 , P1_U3228 , P1_U3227 , P1_U3226 , P1_U3225 , P1_U3224;
output P1_U3223 , P1_U3222 , P1_U3221 , P1_U3220 , P1_U3219 , P1_U3218 , P1_U3217;
output P1_U3216 , P1_U3215 , P1_U3214 , P1_U3213 , P1_U3086 , P1_U3085 , P1_U4016;
output P2_U3327 , P2_U3326 , P2_U3325 , P2_U3324 , P2_U3323 , P2_U3322 , P2_U3321;
output P2_U3320 , P2_U3319 , P2_U3318 , P2_U3317 , P2_U3316 , P2_U3315 , P2_U3314;
output P2_U3313 , P2_U3312 , P2_U3311 , P2_U3310 , P2_U3309 , P2_U3308 , P2_U3307;
output P2_U3306 , P2_U3305 , P2_U3304 , P2_U3303 , P2_U3302 , P2_U3301 , P2_U3300;
output P2_U3299 , P2_U3298 , P2_U3297 , P2_U3296 , P2_U3416 , P2_U3417 , P2_U3295;
output P2_U3294 , P2_U3293 , P2_U3292 , P2_U3291 , P2_U3290 , P2_U3289 , P2_U3288;
output P2_U3287 , P2_U3286 , P2_U3285 , P2_U3284 , P2_U3283 , P2_U3282 , P2_U3281;
output P2_U3280 , P2_U3279 , P2_U3278 , P2_U3277 , P2_U3276 , P2_U3275 , P2_U3274;
output P2_U3273 , P2_U3272 , P2_U3271 , P2_U3270 , P2_U3269 , P2_U3268 , P2_U3267;
output P2_U3266 , P2_U3430 , P2_U3433 , P2_U3436 , P2_U3439 , P2_U3442 , P2_U3445;
output P2_U3448 , P2_U3451 , P2_U3454 , P2_U3457 , P2_U3460 , P2_U3463 , P2_U3466;
output P2_U3469 , P2_U3472 , P2_U3475 , P2_U3478 , P2_U3481 , P2_U3484 , P2_U3486;
output P2_U3487 , P2_U3488 , P2_U3489 , P2_U3490 , P2_U3491 , P2_U3492 , P2_U3493;
output P2_U3494 , P2_U3495 , P2_U3496 , P2_U3497 , P2_U3498 , P2_U3499 , P2_U3500;
output P2_U3501 , P2_U3502 , P2_U3503 , P2_U3504 , P2_U3505 , P2_U3506 , P2_U3507;
output P2_U3508 , P2_U3509 , P2_U3510 , P2_U3511 , P2_U3512 , P2_U3513 , P2_U3514;
output P2_U3515 , P2_U3516 , P2_U3517 , P2_U3518 , P2_U3519 , P2_U3520 , P2_U3521;
output P2_U3522 , P2_U3523 , P2_U3524 , P2_U3525 , P2_U3526 , P2_U3527 , P2_U3528;
output P2_U3529 , P2_U3530 , P2_U3265 , P2_U3264 , P2_U3263 , P2_U3262 , P2_U3261;
output P2_U3260 , P2_U3259 , P2_U3258 , P2_U3257 , P2_U3256 , P2_U3255 , P2_U3254;
output P2_U3253 , P2_U3252 , P2_U3251 , P2_U3250 , P2_U3249 , P2_U3248 , P2_U3247;
output P2_U3246 , P2_U3245 , P2_U3244 , P2_U3243 , P2_U3242 , P2_U3241 , P2_U3240;
output P2_U3239 , P2_U3238 , P2_U3237 , P2_U3236 , P2_U3235 , P2_U3234 , P2_U3233;
output P2_U3232 , P2_U3231 , P2_U3230 , P2_U3229 , P2_U3228 , P2_U3227 , P2_U3226;
output P2_U3225 , P2_U3224 , P2_U3223 , P2_U3222 , P2_U3221 , P2_U3220 , P2_U3219;
output P2_U3218 , P2_U3217 , P2_U3216 , P2_U3215 , P2_U3214 , P2_U3531 , P2_U3532;
output P2_U3533 , P2_U3534 , P2_U3535 , P2_U3536 , P2_U3537 , P2_U3538 , P2_U3539;
output P2_U3540 , P2_U3541 , P2_U3542 , P2_U3543 , P2_U3544 , P2_U3545 , P2_U3546;
output P2_U3547 , P2_U3548 , P2_U3549 , P2_U3550 , P2_U3551 , P2_U3552 , P2_U3553;
output P2_U3554 , P2_U3555 , P2_U3556 , P2_U3557 , P2_U3558 , P2_U3559 , P2_U3560;
output P2_U3561 , P2_U3562 , P2_U3328 , P2_U3213 , P2_U3212 , P2_U3211 , P2_U3210;
output P2_U3209 , P2_U3208 , P2_U3207 , P2_U3206 , P2_U3205 , P2_U3204 , P2_U3203;
output P2_U3202 , P2_U3201 , P2_U3200 , P2_U3199 , P2_U3198 , P2_U3197 , P2_U3196;
output P2_U3195 , P2_U3194 , P2_U3193 , P2_U3192 , P2_U3191 , P2_U3190 , P2_U3189;
output P2_U3188 , P2_U3187 , P2_U3186 , P2_U3185 , P2_U3088 , P2_U3087 , P2_U3947;
output P3_U3295 , P3_U3294 , P3_U3293 , P3_U3292 , P3_U3291 , P3_U3290 , P3_U3289;
output P3_U3288 , P3_U3287 , P3_U3286 , P3_U3285 , P3_U3284 , P3_U3283 , P3_U3282;
output P3_U3281 , P3_U3280 , P3_U3279 , P3_U3278 , P3_U3277 , P3_U3276 , P3_U3275;
output P3_U3274 , P3_U3273 , P3_U3272 , P3_U3271 , P3_U3270 , P3_U3269 , P3_U3268;
output P3_U3267 , P3_U3266 , P3_U3265 , P3_U3264 , P3_U3376 , P3_U3377 , P3_U3263;
output P3_U3262 , P3_U3261 , P3_U3260 , P3_U3259 , P3_U3258 , P3_U3257 , P3_U3256;
output P3_U3255 , P3_U3254 , P3_U3253 , P3_U3252 , P3_U3251 , P3_U3250 , P3_U3249;
output P3_U3248 , P3_U3247 , P3_U3246 , P3_U3245 , P3_U3244 , P3_U3243 , P3_U3242;
output P3_U3241 , P3_U3240 , P3_U3239 , P3_U3238 , P3_U3237 , P3_U3236 , P3_U3235;
output P3_U3234 , P3_U3390 , P3_U3393 , P3_U3396 , P3_U3399 , P3_U3402 , P3_U3405;
output P3_U3408 , P3_U3411 , P3_U3414 , P3_U3417 , P3_U3420 , P3_U3423 , P3_U3426;
output P3_U3429 , P3_U3432 , P3_U3435 , P3_U3438 , P3_U3441 , P3_U3444 , P3_U3446;
output P3_U3447 , P3_U3448 , P3_U3449 , P3_U3450 , P3_U3451 , P3_U3452 , P3_U3453;
output P3_U3454 , P3_U3455 , P3_U3456 , P3_U3457 , P3_U3458 , P3_U3459 , P3_U3460;
output P3_U3461 , P3_U3462 , P3_U3463 , P3_U3464 , P3_U3465 , P3_U3466 , P3_U3467;
output P3_U3468 , P3_U3469 , P3_U3470 , P3_U3471 , P3_U3472 , P3_U3473 , P3_U3474;
output P3_U3475 , P3_U3476 , P3_U3477 , P3_U3478 , P3_U3479 , P3_U3480 , P3_U3481;
output P3_U3482 , P3_U3483 , P3_U3484 , P3_U3485 , P3_U3486 , P3_U3487 , P3_U3488;
output P3_U3489 , P3_U3490 , P3_U3233 , P3_U3232 , P3_U3231 , P3_U3230 , P3_U3229;
output P3_U3228 , P3_U3227 , P3_U3226 , P3_U3225 , P3_U3224 , P3_U3223 , P3_U3222;
output P3_U3221 , P3_U3220 , P3_U3219 , P3_U3218 , P3_U3217 , P3_U3216 , P3_U3215;
output P3_U3214 , P3_U3213 , P3_U3212 , P3_U3211 , P3_U3210 , P3_U3209 , P3_U3208;
output P3_U3207 , P3_U3206 , P3_U3205 , P3_U3204 , P3_U3203 , P3_U3202 , P3_U3201;
output P3_U3200 , P3_U3199 , P3_U3198 , P3_U3197 , P3_U3196 , P3_U3195 , P3_U3194;
output P3_U3193 , P3_U3192 , P3_U3191 , P3_U3190 , P3_U3189 , P3_U3188 , P3_U3187;
output P3_U3186 , P3_U3185 , P3_U3184 , P3_U3183 , P3_U3182 , P3_U3491 , P3_U3492;
output P3_U3493 , P3_U3494 , P3_U3495 , P3_U3496 , P3_U3497 , P3_U3498 , P3_U3499;
output P3_U3500 , P3_U3501 , P3_U3502 , P3_U3503 , P3_U3504 , P3_U3505 , P3_U3506;
output P3_U3507 , P3_U3508 , P3_U3509 , P3_U3510 , P3_U3511 , P3_U3512 , P3_U3513;
output P3_U3514 , P3_U3515 , P3_U3516 , P3_U3517 , P3_U3518 , P3_U3519 , P3_U3520;
output P3_U3521 , P3_U3522 , P3_U3296 , P3_U3181 , P3_U3180 , P3_U3179 , P3_U3178;
output P3_U3177 , P3_U3176 , P3_U3175 , P3_U3174 , P3_U3173 , P3_U3172 , P3_U3171;
output P3_U3170 , P3_U3169 , P3_U3168 , P3_U3167 , P3_U3166 , P3_U3165 , P3_U3164;
output P3_U3163 , P3_U3162 , P3_U3161 , P3_U3160 , P3_U3159 , P3_U3158 , P3_U3157;
output P3_U3156 , P3_U3155 , P3_U3154 , P3_U3153 , P3_U3151 , P3_U3150 , P3_U3897;

input SI_31_ , SI_30_ , SI_29_ , SI_28_ , SI_27_ , SI_26_;
input SI_25_ , SI_24_ , SI_23_ , SI_22_ , SI_21_ , SI_20_;
input SI_19_ , SI_18_ , SI_17_ , SI_16_ , SI_15_ , SI_14_;
input SI_13_ , SI_12_ , SI_11_ , SI_10_ , SI_9_ , SI_8_;
input SI_7_ , SI_6_ , SI_5_ , SI_4_ , SI_3_ , SI_2_;
input SI_1_ , SI_0_;
input P1_IR_REG_0_ , P1_IR_REG_1_ , P1_IR_REG_2_ , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_;
input P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_10_ , P1_IR_REG_11_;
input P1_IR_REG_12_ , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_;
input P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_20_ , P1_IR_REG_21_ , P1_IR_REG_22_ , P1_IR_REG_23_;
input P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ , P1_IR_REG_27_ , P1_IR_REG_28_ , P1_IR_REG_29_;
input P1_IR_REG_30_ , P1_IR_REG_31_ , P1_D_REG_0_ , P1_D_REG_1_ , P1_D_REG_2_ , P1_D_REG_3_;
input P1_D_REG_4_ , P1_D_REG_5_ , P1_D_REG_6_ , P1_D_REG_7_ , P1_D_REG_8_ , P1_D_REG_9_;
input P1_D_REG_10_ , P1_D_REG_11_ , P1_D_REG_12_ , P1_D_REG_13_ , P1_D_REG_14_ , P1_D_REG_15_;
input P1_D_REG_16_ , P1_D_REG_17_ , P1_D_REG_18_ , P1_D_REG_19_ , P1_D_REG_20_ , P1_D_REG_21_;
input P1_D_REG_22_ , P1_D_REG_23_ , P1_D_REG_24_ , P1_D_REG_25_ , P1_D_REG_26_ , P1_D_REG_27_;
input P1_D_REG_28_ , P1_D_REG_29_ , P1_D_REG_30_ , P1_D_REG_31_ , P1_REG0_REG_0_ , P1_REG0_REG_1_;
input P1_REG0_REG_2_ , P1_REG0_REG_3_ , P1_REG0_REG_4_ , P1_REG0_REG_5_ , P1_REG0_REG_6_ , P1_REG0_REG_7_;
input P1_REG0_REG_8_ , P1_REG0_REG_9_ , P1_REG0_REG_10_ , P1_REG0_REG_11_ , P1_REG0_REG_12_ , P1_REG0_REG_13_;
input P1_REG0_REG_14_ , P1_REG0_REG_15_ , P1_REG0_REG_16_ , P1_REG0_REG_17_ , P1_REG0_REG_18_ , P1_REG0_REG_19_;
input P1_REG0_REG_20_ , P1_REG0_REG_21_ , P1_REG0_REG_22_ , P1_REG0_REG_23_ , P1_REG0_REG_24_ , P1_REG0_REG_25_;
input P1_REG0_REG_26_ , P1_REG0_REG_27_ , P1_REG0_REG_28_ , P1_REG0_REG_29_ , P1_REG0_REG_30_ , P1_REG0_REG_31_;
input P1_REG1_REG_0_ , P1_REG1_REG_1_ , P1_REG1_REG_2_ , P1_REG1_REG_3_ , P1_REG1_REG_4_ , P1_REG1_REG_5_;
input P1_REG1_REG_6_ , P1_REG1_REG_7_ , P1_REG1_REG_8_ , P1_REG1_REG_9_ , P1_REG1_REG_10_ , P1_REG1_REG_11_;
input P1_REG1_REG_12_ , P1_REG1_REG_13_ , P1_REG1_REG_14_ , P1_REG1_REG_15_ , P1_REG1_REG_16_ , P1_REG1_REG_17_;
input P1_REG1_REG_18_ , P1_REG1_REG_19_ , P1_REG1_REG_20_ , P1_REG1_REG_21_ , P1_REG1_REG_22_ , P1_REG1_REG_23_;
input P1_REG1_REG_24_ , P1_REG1_REG_25_ , P1_REG1_REG_26_ , P1_REG1_REG_27_ , P1_REG1_REG_28_ , P1_REG1_REG_29_;
input P1_REG1_REG_30_ , P1_REG1_REG_31_ , P1_REG2_REG_0_ , P1_REG2_REG_1_ , P1_REG2_REG_2_ , P1_REG2_REG_3_;
input P1_REG2_REG_4_ , P1_REG2_REG_5_ , P1_REG2_REG_6_ , P1_REG2_REG_7_ , P1_REG2_REG_8_ , P1_REG2_REG_9_;
input P1_REG2_REG_10_ , P1_REG2_REG_11_ , P1_REG2_REG_12_ , P1_REG2_REG_13_ , P1_REG2_REG_14_ , P1_REG2_REG_15_;
input P1_REG2_REG_16_ , P1_REG2_REG_17_ , P1_REG2_REG_18_ , P1_REG2_REG_19_ , P1_REG2_REG_20_ , P1_REG2_REG_21_;
input P1_REG2_REG_22_ , P1_REG2_REG_23_ , P1_REG2_REG_24_ , P1_REG2_REG_25_ , P1_REG2_REG_26_ , P1_REG2_REG_27_;
input P1_REG2_REG_28_ , P1_REG2_REG_29_ , P1_REG2_REG_30_ , P1_REG2_REG_31_ , P1_ADDR_REG_19_ , P1_ADDR_REG_18_;
input P1_ADDR_REG_17_ , P1_ADDR_REG_16_ , P1_ADDR_REG_15_ , P1_ADDR_REG_14_ , P1_ADDR_REG_13_ , P1_ADDR_REG_12_;
input P1_ADDR_REG_11_ , P1_ADDR_REG_10_ , P1_ADDR_REG_9_ , P1_ADDR_REG_8_ , P1_ADDR_REG_7_ , P1_ADDR_REG_6_;
input P1_ADDR_REG_5_ , P1_ADDR_REG_4_ , P1_ADDR_REG_3_ , P1_ADDR_REG_2_ , P1_ADDR_REG_1_ , P1_ADDR_REG_0_;
input P1_DATAO_REG_0_ , P1_DATAO_REG_1_ , P1_DATAO_REG_2_ , P1_DATAO_REG_3_ , P1_DATAO_REG_4_ , P1_DATAO_REG_5_;
input P1_DATAO_REG_6_ , P1_DATAO_REG_7_ , P1_DATAO_REG_8_ , P1_DATAO_REG_9_ , P1_DATAO_REG_10_ , P1_DATAO_REG_11_;
input P1_DATAO_REG_12_ , P1_DATAO_REG_13_ , P1_DATAO_REG_14_ , P1_DATAO_REG_15_ , P1_DATAO_REG_16_ , P1_DATAO_REG_17_;
input P1_DATAO_REG_18_ , P1_DATAO_REG_19_ , P1_DATAO_REG_20_ , P1_DATAO_REG_21_ , P1_DATAO_REG_22_ , P1_DATAO_REG_23_;
input P1_DATAO_REG_24_ , P1_DATAO_REG_25_ , P1_DATAO_REG_26_ , P1_DATAO_REG_27_ , P1_DATAO_REG_28_ , P1_DATAO_REG_29_;
input P1_DATAO_REG_30_ , P1_DATAO_REG_31_ , P1_B_REG , P1_REG3_REG_15_ , P1_REG3_REG_26_ , P1_REG3_REG_6_;
input P1_REG3_REG_18_ , P1_REG3_REG_2_ , P1_REG3_REG_11_ , P1_REG3_REG_22_ , P1_REG3_REG_13_ , P1_REG3_REG_20_;
input P1_REG3_REG_0_ , P1_REG3_REG_9_ , P1_REG3_REG_4_ , P1_REG3_REG_24_ , P1_REG3_REG_17_ , P1_REG3_REG_5_;
input P1_REG3_REG_16_ , P1_REG3_REG_25_ , P1_REG3_REG_12_ , P1_REG3_REG_21_ , P1_REG3_REG_1_ , P1_REG3_REG_8_;
input P1_REG3_REG_28_ , P1_REG3_REG_19_ , P1_REG3_REG_3_ , P1_REG3_REG_10_ , P1_REG3_REG_23_ , P1_REG3_REG_14_;
input P1_REG3_REG_27_ , P1_REG3_REG_7_ , P1_STATE_REG , P1_RD_REG , P1_WR_REG , P2_IR_REG_0_;
input P2_IR_REG_1_ , P2_IR_REG_2_ , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ , P2_IR_REG_6_;
input P2_IR_REG_7_ , P2_IR_REG_8_ , P2_IR_REG_9_ , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_;
input P2_IR_REG_13_ , P2_IR_REG_14_ , P2_IR_REG_15_ , P2_IR_REG_16_ , P2_IR_REG_17_ , P2_IR_REG_18_;
input P2_IR_REG_19_ , P2_IR_REG_20_ , P2_IR_REG_21_ , P2_IR_REG_22_ , P2_IR_REG_23_ , P2_IR_REG_24_;
input P2_IR_REG_25_ , P2_IR_REG_26_ , P2_IR_REG_27_ , P2_IR_REG_28_ , P2_IR_REG_29_ , P2_IR_REG_30_;
input P2_IR_REG_31_ , P2_D_REG_0_ , P2_D_REG_1_ , P2_D_REG_2_ , P2_D_REG_3_ , P2_D_REG_4_;
input P2_D_REG_5_ , P2_D_REG_6_ , P2_D_REG_7_ , P2_D_REG_8_ , P2_D_REG_9_ , P2_D_REG_10_;
input P2_D_REG_11_ , P2_D_REG_12_ , P2_D_REG_13_ , P2_D_REG_14_ , P2_D_REG_15_ , P2_D_REG_16_;
input P2_D_REG_17_ , P2_D_REG_18_ , P2_D_REG_19_ , P2_D_REG_20_ , P2_D_REG_21_ , P2_D_REG_22_;
input P2_D_REG_23_ , P2_D_REG_24_ , P2_D_REG_25_ , P2_D_REG_26_ , P2_D_REG_27_ , P2_D_REG_28_;
input P2_D_REG_29_ , P2_D_REG_30_ , P2_D_REG_31_ , P2_REG0_REG_0_ , P2_REG0_REG_1_ , P2_REG0_REG_2_;
input P2_REG0_REG_3_ , P2_REG0_REG_4_ , P2_REG0_REG_5_ , P2_REG0_REG_6_ , P2_REG0_REG_7_ , P2_REG0_REG_8_;
input P2_REG0_REG_9_ , P2_REG0_REG_10_ , P2_REG0_REG_11_ , P2_REG0_REG_12_ , P2_REG0_REG_13_ , P2_REG0_REG_14_;
input P2_REG0_REG_15_ , P2_REG0_REG_16_ , P2_REG0_REG_17_ , P2_REG0_REG_18_ , P2_REG0_REG_19_ , P2_REG0_REG_20_;
input P2_REG0_REG_21_ , P2_REG0_REG_22_ , P2_REG0_REG_23_ , P2_REG0_REG_24_ , P2_REG0_REG_25_ , P2_REG0_REG_26_;
input P2_REG0_REG_27_ , P2_REG0_REG_28_ , P2_REG0_REG_29_ , P2_REG0_REG_30_ , P2_REG0_REG_31_ , P2_REG1_REG_0_;
input P2_REG1_REG_1_ , P2_REG1_REG_2_ , P2_REG1_REG_3_ , P2_REG1_REG_4_ , P2_REG1_REG_5_ , P2_REG1_REG_6_;
input P2_REG1_REG_7_ , P2_REG1_REG_8_ , P2_REG1_REG_9_ , P2_REG1_REG_10_ , P2_REG1_REG_11_ , P2_REG1_REG_12_;
input P2_REG1_REG_13_ , P2_REG1_REG_14_ , P2_REG1_REG_15_ , P2_REG1_REG_16_ , P2_REG1_REG_17_ , P2_REG1_REG_18_;
input P2_REG1_REG_19_ , P2_REG1_REG_20_ , P2_REG1_REG_21_ , P2_REG1_REG_22_ , P2_REG1_REG_23_ , P2_REG1_REG_24_;
input P2_REG1_REG_25_ , P2_REG1_REG_26_ , P2_REG1_REG_27_ , P2_REG1_REG_28_ , P2_REG1_REG_29_ , P2_REG1_REG_30_;
input P2_REG1_REG_31_ , P2_REG2_REG_0_ , P2_REG2_REG_1_ , P2_REG2_REG_2_ , P2_REG2_REG_3_ , P2_REG2_REG_4_;
input P2_REG2_REG_5_ , P2_REG2_REG_6_ , P2_REG2_REG_7_ , P2_REG2_REG_8_ , P2_REG2_REG_9_ , P2_REG2_REG_10_;
input P2_REG2_REG_11_ , P2_REG2_REG_12_ , P2_REG2_REG_13_ , P2_REG2_REG_14_ , P2_REG2_REG_15_ , P2_REG2_REG_16_;
input P2_REG2_REG_17_ , P2_REG2_REG_18_ , P2_REG2_REG_19_ , P2_REG2_REG_20_ , P2_REG2_REG_21_ , P2_REG2_REG_22_;
input P2_REG2_REG_23_ , P2_REG2_REG_24_ , P2_REG2_REG_25_ , P2_REG2_REG_26_ , P2_REG2_REG_27_ , P2_REG2_REG_28_;
input P2_REG2_REG_29_ , P2_REG2_REG_30_ , P2_REG2_REG_31_ , P2_ADDR_REG_19_ , P2_ADDR_REG_18_ , P2_ADDR_REG_17_;
input P2_ADDR_REG_16_ , P2_ADDR_REG_15_ , P2_ADDR_REG_14_ , P2_ADDR_REG_13_ , P2_ADDR_REG_12_ , P2_ADDR_REG_11_;
input P2_ADDR_REG_10_ , P2_ADDR_REG_9_ , P2_ADDR_REG_8_ , P2_ADDR_REG_7_ , P2_ADDR_REG_6_ , P2_ADDR_REG_5_;
input P2_ADDR_REG_4_ , P2_ADDR_REG_3_ , P2_ADDR_REG_2_ , P2_ADDR_REG_1_ , P2_ADDR_REG_0_ , P2_DATAO_REG_0_;
input P2_DATAO_REG_1_ , P2_DATAO_REG_2_ , P2_DATAO_REG_3_ , P2_DATAO_REG_4_ , P2_DATAO_REG_5_ , P2_DATAO_REG_6_;
input P2_DATAO_REG_7_ , P2_DATAO_REG_8_ , P2_DATAO_REG_9_ , P2_DATAO_REG_10_ , P2_DATAO_REG_11_ , P2_DATAO_REG_12_;
input P2_DATAO_REG_13_ , P2_DATAO_REG_14_ , P2_DATAO_REG_15_ , P2_DATAO_REG_16_ , P2_DATAO_REG_17_ , P2_DATAO_REG_18_;
input P2_DATAO_REG_19_ , P2_DATAO_REG_20_ , P2_DATAO_REG_21_ , P2_DATAO_REG_22_ , P2_DATAO_REG_23_ , P2_DATAO_REG_24_;
input P2_DATAO_REG_25_ , P2_DATAO_REG_26_ , P2_DATAO_REG_27_ , P2_DATAO_REG_28_ , P2_DATAO_REG_29_ , P2_DATAO_REG_30_;
input P2_DATAO_REG_31_ , P2_B_REG , P2_REG3_REG_15_ , P2_REG3_REG_26_ , P2_REG3_REG_6_ , P2_REG3_REG_18_;
input P2_REG3_REG_2_ , P2_REG3_REG_11_ , P2_REG3_REG_22_ , P2_REG3_REG_13_ , P2_REG3_REG_20_ , P2_REG3_REG_0_;
input P2_REG3_REG_9_ , P2_REG3_REG_4_ , P2_REG3_REG_24_ , P2_REG3_REG_17_ , P2_REG3_REG_5_ , P2_REG3_REG_16_;
input P2_REG3_REG_25_ , P2_REG3_REG_12_ , P2_REG3_REG_21_ , P2_REG3_REG_1_ , P2_REG3_REG_8_ , P2_REG3_REG_28_;
input P2_REG3_REG_19_ , P2_REG3_REG_3_ , P2_REG3_REG_10_ , P2_REG3_REG_23_ , P2_REG3_REG_14_ , P2_REG3_REG_27_;
input P2_REG3_REG_7_ , P2_STATE_REG , P2_RD_REG , P2_WR_REG , P3_IR_REG_0_ , P3_IR_REG_1_;
input P3_IR_REG_2_ , P3_IR_REG_3_ , P3_IR_REG_4_ , P3_IR_REG_5_ , P3_IR_REG_6_ , P3_IR_REG_7_;
input P3_IR_REG_8_ , P3_IR_REG_9_ , P3_IR_REG_10_ , P3_IR_REG_11_ , P3_IR_REG_12_ , P3_IR_REG_13_;
input P3_IR_REG_14_ , P3_IR_REG_15_ , P3_IR_REG_16_ , P3_IR_REG_17_ , P3_IR_REG_18_ , P3_IR_REG_19_;
input P3_IR_REG_20_ , P3_IR_REG_21_ , P3_IR_REG_22_ , P3_IR_REG_23_ , P3_IR_REG_24_ , P3_IR_REG_25_;
input P3_IR_REG_26_ , P3_IR_REG_27_ , P3_IR_REG_28_ , P3_IR_REG_29_ , P3_IR_REG_30_ , P3_IR_REG_31_;
input P3_D_REG_0_ , P3_D_REG_1_ , P3_D_REG_2_ , P3_D_REG_3_ , P3_D_REG_4_ , P3_D_REG_5_;
input P3_D_REG_6_ , P3_D_REG_7_ , P3_D_REG_8_ , P3_D_REG_9_ , P3_D_REG_10_ , P3_D_REG_11_;
input P3_D_REG_12_ , P3_D_REG_13_ , P3_D_REG_14_ , P3_D_REG_15_ , P3_D_REG_16_ , P3_D_REG_17_;
input P3_D_REG_18_ , P3_D_REG_19_ , P3_D_REG_20_ , P3_D_REG_21_ , P3_D_REG_22_ , P3_D_REG_23_;
input P3_D_REG_24_ , P3_D_REG_25_ , P3_D_REG_26_ , P3_D_REG_27_ , P3_D_REG_28_ , P3_D_REG_29_;
input P3_D_REG_30_ , P3_D_REG_31_ , P3_REG0_REG_0_ , P3_REG0_REG_1_ , P3_REG0_REG_2_ , P3_REG0_REG_3_;
input P3_REG0_REG_4_ , P3_REG0_REG_5_ , P3_REG0_REG_6_ , P3_REG0_REG_7_ , P3_REG0_REG_8_ , P3_REG0_REG_9_;
input P3_REG0_REG_10_ , P3_REG0_REG_11_ , P3_REG0_REG_12_ , P3_REG0_REG_13_ , P3_REG0_REG_14_ , P3_REG0_REG_15_;
input P3_REG0_REG_16_ , P3_REG0_REG_17_ , P3_REG0_REG_18_ , P3_REG0_REG_19_ , P3_REG0_REG_20_ , P3_REG0_REG_21_;
input P3_REG0_REG_22_ , P3_REG0_REG_23_ , P3_REG0_REG_24_ , P3_REG0_REG_25_ , P3_REG0_REG_26_ , P3_REG0_REG_27_;
input P3_REG0_REG_28_ , P3_REG0_REG_29_ , P3_REG0_REG_30_ , P3_REG0_REG_31_ , P3_REG1_REG_0_ , P3_REG1_REG_1_;
input P3_REG1_REG_2_ , P3_REG1_REG_3_ , P3_REG1_REG_4_ , P3_REG1_REG_5_ , P3_REG1_REG_6_ , P3_REG1_REG_7_;
input P3_REG1_REG_8_ , P3_REG1_REG_9_ , P3_REG1_REG_10_ , P3_REG1_REG_11_ , P3_REG1_REG_12_ , P3_REG1_REG_13_;
input P3_REG1_REG_14_ , P3_REG1_REG_15_ , P3_REG1_REG_16_ , P3_REG1_REG_17_ , P3_REG1_REG_18_ , P3_REG1_REG_19_;
input P3_REG1_REG_20_ , P3_REG1_REG_21_ , P3_REG1_REG_22_ , P3_REG1_REG_23_ , P3_REG1_REG_24_ , P3_REG1_REG_25_;
input P3_REG1_REG_26_ , P3_REG1_REG_27_ , P3_REG1_REG_28_ , P3_REG1_REG_29_ , P3_REG1_REG_30_ , P3_REG1_REG_31_;
input P3_REG2_REG_0_ , P3_REG2_REG_1_ , P3_REG2_REG_2_ , P3_REG2_REG_3_ , P3_REG2_REG_4_ , P3_REG2_REG_5_;
input P3_REG2_REG_6_ , P3_REG2_REG_7_ , P3_REG2_REG_8_ , P3_REG2_REG_9_ , P3_REG2_REG_10_ , P3_REG2_REG_11_;
input P3_REG2_REG_12_ , P3_REG2_REG_13_ , P3_REG2_REG_14_ , P3_REG2_REG_15_ , P3_REG2_REG_16_ , P3_REG2_REG_17_;
input P3_REG2_REG_18_ , P3_REG2_REG_19_ , P3_REG2_REG_20_ , P3_REG2_REG_21_ , P3_REG2_REG_22_ , P3_REG2_REG_23_;
input P3_REG2_REG_24_ , P3_REG2_REG_25_ , P3_REG2_REG_26_ , P3_REG2_REG_27_ , P3_REG2_REG_28_ , P3_REG2_REG_29_;
input P3_REG2_REG_30_ , P3_REG2_REG_31_ , P3_ADDR_REG_19_ , P3_ADDR_REG_18_ , P3_ADDR_REG_17_ , P3_ADDR_REG_16_;
input P3_ADDR_REG_15_ , P3_ADDR_REG_14_ , P3_ADDR_REG_13_ , P3_ADDR_REG_12_ , P3_ADDR_REG_11_ , P3_ADDR_REG_10_;
input P3_ADDR_REG_9_ , P3_ADDR_REG_8_ , P3_ADDR_REG_7_ , P3_ADDR_REG_6_ , P3_ADDR_REG_5_ , P3_ADDR_REG_4_;
input P3_ADDR_REG_3_ , P3_ADDR_REG_2_ , P3_ADDR_REG_1_ , P3_ADDR_REG_0_ , P3_DATAO_REG_0_ , P3_DATAO_REG_1_;
input P3_DATAO_REG_2_ , P3_DATAO_REG_3_ , P3_DATAO_REG_4_ , P3_DATAO_REG_5_ , P3_DATAO_REG_6_ , P3_DATAO_REG_7_;
input P3_DATAO_REG_8_ , P3_DATAO_REG_9_ , P3_DATAO_REG_10_ , P3_DATAO_REG_11_ , P3_DATAO_REG_12_ , P3_DATAO_REG_13_;
input P3_DATAO_REG_14_ , P3_DATAO_REG_15_ , P3_DATAO_REG_16_ , P3_DATAO_REG_17_ , P3_DATAO_REG_18_ , P3_DATAO_REG_19_;
input P3_DATAO_REG_20_ , P3_DATAO_REG_21_ , P3_DATAO_REG_22_ , P3_DATAO_REG_23_ , P3_DATAO_REG_24_ , P3_DATAO_REG_25_;
input P3_DATAO_REG_26_ , P3_DATAO_REG_27_ , P3_DATAO_REG_28_ , P3_DATAO_REG_29_ , P3_DATAO_REG_30_ , P3_DATAO_REG_31_;
input P3_B_REG , P3_REG3_REG_15_ , P3_REG3_REG_26_ , P3_REG3_REG_6_ , P3_REG3_REG_18_ , P3_REG3_REG_2_;
input P3_REG3_REG_11_ , P3_REG3_REG_22_ , P3_REG3_REG_13_ , P3_REG3_REG_20_ , P3_REG3_REG_0_ , P3_REG3_REG_9_;
input P3_REG3_REG_4_ , P3_REG3_REG_24_ , P3_REG3_REG_17_ , P3_REG3_REG_5_ , P3_REG3_REG_16_ , P3_REG3_REG_25_;
input P3_REG3_REG_12_ , P3_REG3_REG_21_ , P3_REG3_REG_1_ , P3_REG3_REG_8_ , P3_REG3_REG_28_ , P3_REG3_REG_19_;
input P3_REG3_REG_3_ , P3_REG3_REG_10_ , P3_REG3_REG_23_ , P3_REG3_REG_14_ , P3_REG3_REG_27_ , P3_REG3_REG_7_;
input P3_STATE_REG , P3_RD_REG , P3_WR_REG;

wire P3_R1161_U504 , P3_R1161_U503 , P3_R1161_U502 , U30 , U31 , U32 , U33 , U34 , U35 , U36;
wire U37 , U38 , U39 , U40 , U41 , U42 , U43 , U44 , U45 , U46;
wire U47 , U48 , U49 , U50 , U51 , U52 , U53 , U54 , U55 , U56;
wire U57 , U58 , U59 , U60 , U61 , U62 , U63 , U64 , U65 , U66;
wire U67 , U68 , U69 , U70 , U71 , U72 , U73 , U74 , U75 , U76;
wire U77 , U78 , U79 , U80 , U81 , U82 , U83 , U84 , U85 , U86;
wire U87 , U88 , U89 , U90 , U91 , U92 , U93 , U94 , U95 , U96;
wire U97 , U98 , U99 , U100 , U101 , U102 , U103 , U104 , U105 , U106;
wire U107 , U108 , U109 , U110 , U111 , U112 , U113 , U114 , U115 , U116;
wire U117 , U118 , U119 , U120 , U121 , U122 , U123 , U124 , U125 , U126;
wire U127 , U128 , U129 , U130 , U131 , U132 , U133 , U134 , U135 , U136;
wire U137 , U138 , U139 , U140 , U141 , U142 , U143 , U144 , U145 , U146;
wire U147 , U148 , U149 , U150 , U151 , U152 , U153 , U154 , U155 , U156;
wire U157 , U158 , U159 , U160 , U161 , U162 , U163 , U164 , U165 , U166;
wire U167 , U168 , U169 , U170 , U171 , U172 , U173 , U174 , U175 , U176;
wire U177 , U178 , U179 , U180 , U181 , U182 , U183 , U184 , U185 , U186;
wire U187 , U188 , U189 , U190 , U191 , U192 , U193 , U194 , U195 , U196;
wire U197 , U198 , U199 , U200 , U201 , U202 , U203 , U204 , U205 , U206;
wire U207 , U208 , U209 , U210 , U211 , U212 , U213 , U214 , U215 , U216;
wire U217 , U218 , U219 , U220 , U221 , U222 , U223 , U224 , U225 , U226;
wire U227 , U228 , U229 , U230 , U231 , U232 , U233 , U234 , U235 , U236;
wire U237 , U238 , U239 , U240 , U241 , U242 , U243 , U244 , U245 , U246;
wire U247 , U248 , U249 , U250 , U251 , U252 , U253 , U254 , U255 , U256;
wire U257 , U258 , U259 , U260 , U261 , U262 , U263 , U264 , U265 , U266;
wire U267 , U268 , U269 , U270 , U271 , U272 , U273 , U274 , U275 , U276;
wire U277 , U278 , U279 , U280 , U281 , U282 , U283 , U284 , U285 , U286;
wire U287 , U288 , U289 , U290 , U291 , U292 , U293 , U294 , U295 , U296;
wire U297 , U298 , U299 , U300 , U301 , U302 , U303 , U304 , U305 , U306;
wire U307 , U308 , U309 , U310 , U311 , U312 , U313 , U314 , U315 , U316;
wire U317 , U318 , U319 , U320 , U321 , U322 , U323 , U324 , U325 , U326;
wire U327 , U328 , U329 , U330 , U331 , U332 , U333 , U334 , U335 , U336;
wire U337 , U338 , U339 , U340 , U341 , U342 , U343 , U344 , U345 , U346;
wire U347 , U348 , U349 , U350 , U351 , U352 , U353 , U354 , U355 , U356;
wire U357 , U358 , U359 , U360 , U361 , U362 , U363 , U364 , U365 , U366;
wire U367 , U368 , U369 , U370 , U371 , U372 , U373 , U374 , U375 , U376;
wire U377 , U378 , U379 , U380 , U381 , U382 , U383 , U384 , U385 , U386;
wire U387 , U388 , U389 , U390 , U391 , U392 , U393 , U394 , U395 , U396;
wire U397 , U398 , U399 , U400 , U401 , U402 , U403 , U404 , U405 , U406;
wire U407 , U408 , U409 , U410 , U411 , U412 , U413 , U414 , U415 , U416;
wire U417 , U418 , U419 , U420 , U421 , U422 , U423 , U424 , U425 , U426;
wire U427 , P3_R1161_U501 , P3_R1161_U500 , P3_R1161_U499 , P3_R1161_U498 , P3_R1161_U497 , P3_R1161_U496 , P3_R1161_U495 , P3_R1161_U494 , P3_R1161_U493;
wire P3_R1161_U492 , P3_R1161_U491 , P3_R1161_U490 , P1_U3014 , P1_U3015 , P1_U3016 , P1_U3017 , P1_U3018 , P1_U3019 , P1_U3020;
wire P1_U3021 , P1_U3022 , P1_U3023 , P1_U3024 , P1_U3025 , P1_U3026 , P1_U3027 , P1_U3028 , P1_U3029 , P1_U3030;
wire P1_U3031 , P1_U3032 , P1_U3033 , P1_U3034 , P1_U3035 , P1_U3036 , P1_U3037 , P1_U3038 , P1_U3039 , P1_U3040;
wire P1_U3041 , P1_U3042 , P1_U3043 , P1_U3044 , P1_U3045 , P1_U3046 , P1_U3047 , P1_U3048 , P1_U3049 , P1_U3050;
wire P1_U3051 , P1_U3052 , P1_U3053 , P1_U3054 , P1_U3055 , P1_U3056 , P1_U3057 , P1_U3058 , P1_U3059 , P1_U3060;
wire P1_U3061 , P1_U3062 , P1_U3063 , P1_U3064 , P1_U3065 , P1_U3066 , P1_U3067 , P1_U3068 , P1_U3069 , P1_U3070;
wire P1_U3071 , P1_U3072 , P1_U3073 , P1_U3074 , P1_U3075 , P1_U3076 , P1_U3077 , P1_U3078 , P1_U3079 , P1_U3080;
wire P1_U3081 , P1_U3082 , P1_U3083 , P1_U3084 , P1_U3087 , P1_U3088 , P1_U3089 , P1_U3090 , P1_U3091 , P1_U3092;
wire P1_U3093 , P1_U3094 , P1_U3095 , P1_U3096 , P1_U3097 , P1_U3098 , P1_U3099 , P1_U3100 , P1_U3101 , P1_U3102;
wire P1_U3103 , P1_U3104 , P1_U3105 , P1_U3106 , P1_U3107 , P1_U3108 , P1_U3109 , P1_U3110 , P1_U3111 , P1_U3112;
wire P1_U3113 , P1_U3114 , P1_U3115 , P1_U3116 , P1_U3117 , P1_U3118 , P1_U3119 , P1_U3120 , P1_U3121 , P1_U3122;
wire P1_U3123 , P1_U3124 , P1_U3125 , P1_U3126 , P1_U3127 , P1_U3128 , P1_U3129 , P1_U3130 , P1_U3131 , P1_U3132;
wire P1_U3133 , P1_U3134 , P1_U3135 , P1_U3136 , P1_U3137 , P1_U3138 , P1_U3139 , P1_U3140 , P1_U3141 , P1_U3142;
wire P1_U3143 , P1_U3144 , P1_U3145 , P1_U3146 , P1_U3147 , P1_U3148 , P1_U3149 , P1_U3150 , P1_U3151 , P1_U3152;
wire P1_U3153 , P1_U3154 , P1_U3155 , P1_U3156 , P1_U3157 , P1_U3158 , P1_U3159 , P1_U3160 , P1_U3161 , P1_U3162;
wire P1_U3163 , P1_U3164 , P1_U3165 , P1_U3166 , P1_U3167 , P1_U3168 , P1_U3169 , P1_U3170 , P1_U3171 , P1_U3172;
wire P1_U3173 , P1_U3174 , P1_U3175 , P1_U3176 , P1_U3177 , P1_U3178 , P1_U3179 , P1_U3180 , P1_U3181 , P1_U3182;
wire P1_U3183 , P1_U3184 , P1_U3185 , P1_U3186 , P1_U3187 , P1_U3188 , P1_U3189 , P1_U3190 , P1_U3191 , P1_U3192;
wire P1_U3193 , P1_U3194 , P1_U3195 , P1_U3196 , P1_U3197 , P1_U3198 , P1_U3199 , P1_U3200 , P1_U3201 , P1_U3202;
wire P1_U3203 , P1_U3204 , P1_U3205 , P1_U3206 , P1_U3207 , P1_U3208 , P1_U3209 , P1_U3210 , P1_U3211 , P1_U3212;
wire P1_U3357 , P1_U3358 , P1_U3359 , P1_U3360 , P1_U3361 , P1_U3362 , P1_U3363 , P1_U3364 , P1_U3365 , P1_U3366;
wire P1_U3367 , P1_U3368 , P1_U3369 , P1_U3370 , P1_U3371 , P1_U3372 , P1_U3373 , P1_U3374 , P1_U3375 , P1_U3376;
wire P1_U3377 , P1_U3378 , P1_U3379 , P1_U3380 , P1_U3381 , P1_U3382 , P1_U3383 , P1_U3384 , P1_U3385 , P1_U3386;
wire P1_U3387 , P1_U3388 , P1_U3389 , P1_U3390 , P1_U3391 , P1_U3392 , P1_U3393 , P1_U3394 , P1_U3395 , P1_U3396;
wire P1_U3397 , P1_U3398 , P1_U3399 , P1_U3400 , P1_U3401 , P1_U3402 , P1_U3403 , P1_U3404 , P1_U3405 , P1_U3406;
wire P1_U3407 , P1_U3408 , P1_U3409 , P1_U3410 , P1_U3411 , P1_U3412 , P1_U3413 , P1_U3414 , P1_U3415 , P1_U3416;
wire P1_U3417 , P1_U3418 , P1_U3419 , P1_U3420 , P1_U3421 , P1_U3422 , P1_U3423 , P1_U3424 , P1_U3425 , P1_U3426;
wire P1_U3427 , P1_U3428 , P1_U3429 , P1_U3430 , P1_U3431 , P1_U3432 , P1_U3433 , P1_U3434 , P1_U3435 , P1_U3436;
wire P1_U3437 , P1_U3438 , P1_U3439 , P1_U3440 , P1_U3441 , P1_U3442 , P1_U3443 , P1_U3444 , P1_U3447 , P1_U3448;
wire P1_U3449 , P1_U3450 , P1_U3451 , P1_U3452 , P1_U3453 , P1_U3454 , P1_U3455 , P1_U3456 , P1_U3457 , P1_U3458;
wire P1_U3460 , P1_U3461 , P1_U3463 , P1_U3464 , P1_U3466 , P1_U3467 , P1_U3469 , P1_U3470 , P1_U3472 , P1_U3473;
wire P1_U3475 , P1_U3476 , P1_U3478 , P1_U3479 , P1_U3481 , P1_U3482 , P1_U3484 , P1_U3485 , P1_U3487 , P1_U3488;
wire P1_U3490 , P1_U3491 , P1_U3493 , P1_U3494 , P1_U3496 , P1_U3497 , P1_U3499 , P1_U3500 , P1_U3502 , P1_U3503;
wire P1_U3505 , P1_U3506 , P1_U3508 , P1_U3509 , P1_U3511 , P1_U3512 , P1_U3514 , P1_U3592 , P1_U3593 , P1_U3594;
wire P1_U3595 , P1_U3596 , P1_U3597 , P1_U3598 , P1_U3599 , P1_U3600 , P1_U3601 , P1_U3602 , P1_U3603 , P1_U3604;
wire P1_U3605 , P1_U3606 , P1_U3607 , P1_U3608 , P1_U3609 , P1_U3610 , P1_U3611 , P1_U3612 , P1_U3613 , P1_U3614;
wire P1_U3615 , P1_U3616 , P1_U3617 , P1_U3618 , P1_U3619 , P1_U3620 , P1_U3621 , P1_U3622 , P1_U3623 , P1_U3624;
wire P1_U3625 , P1_U3626 , P1_U3627 , P1_U3628 , P1_U3629 , P1_U3630 , P1_U3631 , P1_U3632 , P1_U3633 , P1_U3634;
wire P1_U3635 , P1_U3636 , P1_U3637 , P1_U3638 , P1_U3639 , P1_U3640 , P1_U3641 , P1_U3642 , P1_U3643 , P1_U3644;
wire P1_U3645 , P1_U3646 , P1_U3647 , P1_U3648 , P1_U3649 , P1_U3650 , P1_U3651 , P1_U3652 , P1_U3653 , P1_U3654;
wire P1_U3655 , P1_U3656 , P1_U3657 , P1_U3658 , P1_U3659 , P1_U3660 , P1_U3661 , P1_U3662 , P1_U3663 , P1_U3664;
wire P1_U3665 , P1_U3666 , P1_U3667 , P1_U3668 , P1_U3669 , P1_U3670 , P1_U3671 , P1_U3672 , P1_U3673 , P1_U3674;
wire P1_U3675 , P1_U3676 , P1_U3677 , P1_U3678 , P1_U3679 , P1_U3680 , P1_U3681 , P1_U3682 , P1_U3683 , P1_U3684;
wire P1_U3685 , P1_U3686 , P1_U3687 , P1_U3688 , P1_U3689 , P1_U3690 , P1_U3691 , P1_U3692 , P1_U3693 , P1_U3694;
wire P1_U3695 , P1_U3696 , P1_U3697 , P1_U3698 , P1_U3699 , P1_U3700 , P1_U3701 , P1_U3702 , P1_U3703 , P1_U3704;
wire P1_U3705 , P1_U3706 , P1_U3707 , P1_U3708 , P1_U3709 , P1_U3710 , P1_U3711 , P1_U3712 , P1_U3713 , P1_U3714;
wire P1_U3715 , P1_U3716 , P1_U3717 , P1_U3718 , P1_U3719 , P1_U3720 , P1_U3721 , P1_U3722 , P1_U3723 , P1_U3724;
wire P1_U3725 , P1_U3726 , P1_U3727 , P1_U3728 , P1_U3729 , P1_U3730 , P1_U3731 , P1_U3732 , P1_U3733 , P1_U3734;
wire P1_U3735 , P1_U3736 , P1_U3737 , P1_U3738 , P1_U3739 , P1_U3740 , P1_U3741 , P1_U3742 , P1_U3743 , P1_U3744;
wire P1_U3745 , P1_U3746 , P1_U3747 , P1_U3748 , P1_U3749 , P1_U3750 , P1_U3751 , P1_U3752 , P1_U3753 , P1_U3754;
wire P1_U3755 , P1_U3756 , P1_U3757 , P1_U3758 , P1_U3759 , P1_U3760 , P1_U3761 , P1_U3762 , P1_U3763 , P1_U3764;
wire P1_U3765 , P1_U3766 , P1_U3767 , P1_U3768 , P1_U3769 , P1_U3770 , P1_U3771 , P1_U3772 , P1_U3773 , P1_U3774;
wire P1_U3775 , P1_U3776 , P1_U3777 , P1_U3778 , P1_U3779 , P1_U3780 , P1_U3781 , P1_U3782 , P1_U3783 , P1_U3784;
wire P1_U3785 , P1_U3786 , P1_U3787 , P1_U3788 , P1_U3789 , P1_U3790 , P1_U3791 , P1_U3792 , P1_U3793 , P1_U3794;
wire P1_U3795 , P1_U3796 , P1_U3797 , P1_U3798 , P1_U3799 , P1_U3800 , P1_U3801 , P1_U3802 , P1_U3803 , P1_U3804;
wire P1_U3805 , P1_U3806 , P1_U3807 , P1_U3808 , P1_U3809 , P1_U3810 , P1_U3811 , P1_U3812 , P1_U3813 , P1_U3814;
wire P1_U3815 , P1_U3816 , P1_U3817 , P1_U3818 , P1_U3819 , P1_U3820 , P1_U3821 , P1_U3822 , P1_U3823 , P1_U3824;
wire P1_U3825 , P1_U3826 , P1_U3827 , P1_U3828 , P1_U3829 , P1_U3830 , P1_U3831 , P1_U3832 , P1_U3833 , P1_U3834;
wire P1_U3835 , P1_U3836 , P1_U3837 , P1_U3838 , P1_U3839 , P1_U3840 , P1_U3841 , P1_U3842 , P1_U3843 , P1_U3844;
wire P1_U3845 , P1_U3846 , P1_U3847 , P1_U3848 , P1_U3849 , P1_U3850 , P1_U3851 , P1_U3852 , P1_U3853 , P1_U3854;
wire P1_U3855 , P1_U3856 , P1_U3857 , P1_U3858 , P1_U3859 , P1_U3860 , P1_U3861 , P1_U3862 , P1_U3863 , P1_U3864;
wire P1_U3865 , P1_U3866 , P1_U3867 , P1_U3868 , P1_U3869 , P1_U3870 , P1_U3871 , P1_U3872 , P1_U3873 , P1_U3874;
wire P1_U3875 , P1_U3876 , P1_U3877 , P1_U3878 , P1_U3879 , P1_U3880 , P1_U3881 , P1_U3882 , P1_U3883 , P1_U3884;
wire P1_U3885 , P1_U3886 , P1_U3887 , P1_U3888 , P1_U3889 , P1_U3890 , P1_U3891 , P1_U3892 , P1_U3893 , P1_U3894;
wire P1_U3895 , P1_U3896 , P1_U3897 , P1_U3898 , P1_U3899 , P1_U3900 , P1_U3901 , P1_U3902 , P1_U3903 , P1_U3904;
wire P1_U3905 , P1_U3906 , P1_U3907 , P1_U3908 , P1_U3909 , P1_U3910 , P1_U3911 , P1_U3912 , P1_U3913 , P1_U3914;
wire P1_U3915 , P1_U3916 , P1_U3917 , P1_U3918 , P1_U3919 , P1_U3920 , P1_U3921 , P1_U3922 , P1_U3923 , P1_U3924;
wire P1_U3925 , P1_U3926 , P1_U3927 , P1_U3928 , P1_U3929 , P1_U3930 , P1_U3931 , P1_U3932 , P1_U3933 , P1_U3934;
wire P1_U3935 , P1_U3936 , P1_U3937 , P1_U3938 , P1_U3939 , P1_U3940 , P1_U3941 , P1_U3942 , P1_U3943 , P1_U3944;
wire P1_U3945 , P1_U3946 , P1_U3947 , P1_U3948 , P1_U3949 , P1_U3950 , P1_U3951 , P1_U3952 , P1_U3953 , P1_U3954;
wire P1_U3955 , P1_U3956 , P1_U3957 , P1_U3958 , P1_U3959 , P1_U3960 , P1_U3961 , P1_U3962 , P1_U3963 , P1_U3964;
wire P1_U3965 , P1_U3966 , P1_U3967 , P1_U3968 , P1_U3969 , P1_U3970 , P1_U3971 , P1_U3972 , P1_U3973 , P1_U3974;
wire P1_U3975 , P1_U3976 , P1_U3977 , P1_U3978 , P1_U3979 , P1_U3980 , P1_U3981 , P1_U3982 , P1_U3983 , P1_U3984;
wire P1_U3985 , P1_U3986 , P1_U3987 , P1_U3988 , P1_U3989 , P1_U3990 , P1_U3991 , P1_U3992 , P1_U3993 , P1_U3994;
wire P1_U3995 , P1_U3996 , P1_U3997 , P1_U3998 , P1_U3999 , P1_U4000 , P1_U4001 , P1_U4002 , P1_U4003 , P1_U4004;
wire P1_U4005 , P1_U4006 , P1_U4007 , P1_U4008 , P1_U4009 , P1_U4010 , P1_U4011 , P1_U4012 , P1_U4013 , P1_U4014;
wire P1_U4015 , P1_U4017 , P1_U4018 , P1_U4019 , P1_U4020 , P1_U4021 , P1_U4022 , P1_U4023 , P1_U4024 , P1_U4025;
wire P1_U4026 , P1_U4027 , P1_U4028 , P1_U4029 , P1_U4030 , P1_U4031 , P1_U4032 , P1_U4033 , P1_U4034 , P1_U4035;
wire P1_U4036 , P1_U4037 , P1_U4038 , P1_U4039 , P1_U4040 , P1_U4041 , P1_U4042 , P1_U4043 , P1_U4044 , P1_U4045;
wire P1_U4046 , P1_U4047 , P1_U4048 , P1_U4049 , P1_U4050 , P1_U4051 , P1_U4052 , P1_U4053 , P1_U4054 , P1_U4055;
wire P1_U4056 , P1_U4057 , P1_U4058 , P1_U4059 , P1_U4060 , P1_U4061 , P1_U4062 , P1_U4063 , P1_U4064 , P1_U4065;
wire P1_U4066 , P1_U4067 , P1_U4068 , P1_U4069 , P1_U4070 , P1_U4071 , P1_U4072 , P1_U4073 , P1_U4074 , P1_U4075;
wire P1_U4076 , P1_U4077 , P1_U4078 , P1_U4079 , P1_U4080 , P1_U4081 , P1_U4082 , P1_U4083 , P1_U4084 , P1_U4085;
wire P1_U4086 , P1_U4087 , P1_U4088 , P1_U4089 , P1_U4090 , P1_U4091 , P1_U4092 , P1_U4093 , P1_U4094 , P1_U4095;
wire P1_U4096 , P1_U4097 , P1_U4098 , P1_U4099 , P1_U4100 , P1_U4101 , P1_U4102 , P1_U4103 , P1_U4104 , P1_U4105;
wire P1_U4106 , P1_U4107 , P1_U4108 , P1_U4109 , P1_U4110 , P1_U4111 , P1_U4112 , P1_U4113 , P1_U4114 , P1_U4115;
wire P1_U4116 , P1_U4117 , P1_U4118 , P1_U4119 , P1_U4120 , P1_U4121 , P1_U4122 , P1_U4123 , P1_U4124 , P1_U4125;
wire P1_U4126 , P1_U4127 , P1_U4128 , P1_U4129 , P1_U4130 , P1_U4131 , P1_U4132 , P1_U4133 , P1_U4134 , P1_U4135;
wire P1_U4136 , P1_U4137 , P1_U4138 , P1_U4139 , P1_U4140 , P1_U4141 , P1_U4142 , P1_U4143 , P1_U4144 , P1_U4145;
wire P1_U4146 , P1_U4147 , P1_U4148 , P1_U4149 , P1_U4150 , P1_U4151 , P1_U4152 , P1_U4153 , P1_U4154 , P1_U4155;
wire P1_U4156 , P1_U4157 , P1_U4158 , P1_U4159 , P1_U4160 , P1_U4161 , P1_U4162 , P1_U4163 , P1_U4164 , P1_U4165;
wire P1_U4166 , P1_U4167 , P1_U4168 , P1_U4169 , P1_U4170 , P1_U4171 , P1_U4172 , P1_U4173 , P1_U4174 , P1_U4175;
wire P1_U4176 , P1_U4177 , P1_U4178 , P1_U4179 , P1_U4180 , P1_U4181 , P1_U4182 , P1_U4183 , P1_U4184 , P1_U4185;
wire P1_U4186 , P1_U4187 , P1_U4188 , P1_U4189 , P1_U4190 , P1_U4191 , P1_U4192 , P1_U4193 , P1_U4194 , P1_U4195;
wire P1_U4196 , P1_U4197 , P1_U4198 , P1_U4199 , P1_U4200 , P1_U4201 , P1_U4202 , P1_U4203 , P1_U4204 , P1_U4205;
wire P1_U4206 , P1_U4207 , P1_U4208 , P1_U4209 , P1_U4210 , P1_U4211 , P1_U4212 , P1_U4213 , P1_U4214 , P1_U4215;
wire P1_U4216 , P1_U4217 , P1_U4218 , P1_U4219 , P1_U4220 , P1_U4221 , P1_U4222 , P1_U4223 , P1_U4224 , P1_U4225;
wire P1_U4226 , P1_U4227 , P1_U4228 , P1_U4229 , P1_U4230 , P1_U4231 , P1_U4232 , P1_U4233 , P1_U4234 , P1_U4235;
wire P1_U4236 , P1_U4237 , P1_U4238 , P1_U4239 , P1_U4240 , P1_U4241 , P1_U4242 , P1_U4243 , P1_U4244 , P1_U4245;
wire P1_U4246 , P1_U4247 , P1_U4248 , P1_U4249 , P1_U4250 , P1_U4251 , P1_U4252 , P1_U4253 , P1_U4254 , P1_U4255;
wire P1_U4256 , P1_U4257 , P1_U4258 , P1_U4259 , P1_U4260 , P1_U4261 , P1_U4262 , P1_U4263 , P1_U4264 , P1_U4265;
wire P1_U4266 , P1_U4267 , P1_U4268 , P1_U4269 , P1_U4270 , P1_U4271 , P1_U4272 , P1_U4273 , P1_U4274 , P1_U4275;
wire P1_U4276 , P1_U4277 , P1_U4278 , P1_U4279 , P1_U4280 , P1_U4281 , P1_U4282 , P1_U4283 , P1_U4284 , P1_U4285;
wire P1_U4286 , P1_U4287 , P1_U4288 , P1_U4289 , P1_U4290 , P1_U4291 , P1_U4292 , P1_U4293 , P1_U4294 , P1_U4295;
wire P1_U4296 , P1_U4297 , P1_U4298 , P1_U4299 , P1_U4300 , P1_U4301 , P1_U4302 , P1_U4303 , P1_U4304 , P1_U4305;
wire P1_U4306 , P1_U4307 , P1_U4308 , P1_U4309 , P1_U4310 , P1_U4311 , P1_U4312 , P1_U4313 , P1_U4314 , P1_U4315;
wire P1_U4316 , P1_U4317 , P1_U4318 , P1_U4319 , P1_U4320 , P1_U4321 , P1_U4322 , P1_U4323 , P1_U4324 , P1_U4325;
wire P1_U4326 , P1_U4327 , P1_U4328 , P1_U4329 , P1_U4330 , P1_U4331 , P1_U4332 , P1_U4333 , P1_U4334 , P1_U4335;
wire P1_U4336 , P1_U4337 , P1_U4338 , P1_U4339 , P1_U4340 , P1_U4341 , P1_U4342 , P1_U4343 , P1_U4344 , P1_U4345;
wire P1_U4346 , P1_U4347 , P1_U4348 , P1_U4349 , P1_U4350 , P1_U4351 , P1_U4352 , P1_U4353 , P1_U4354 , P1_U4355;
wire P1_U4356 , P1_U4357 , P1_U4358 , P1_U4359 , P1_U4360 , P1_U4361 , P1_U4362 , P1_U4363 , P1_U4364 , P1_U4365;
wire P1_U4366 , P1_U4367 , P1_U4368 , P1_U4369 , P1_U4370 , P1_U4371 , P1_U4372 , P1_U4373 , P1_U4374 , P1_U4375;
wire P1_U4376 , P1_U4377 , P1_U4378 , P1_U4379 , P1_U4380 , P1_U4381 , P1_U4382 , P1_U4383 , P1_U4384 , P1_U4385;
wire P1_U4386 , P1_U4387 , P1_U4388 , P1_U4389 , P1_U4390 , P1_U4391 , P1_U4392 , P1_U4393 , P1_U4394 , P1_U4395;
wire P1_U4396 , P1_U4397 , P1_U4398 , P1_U4399 , P1_U4400 , P1_U4401 , P1_U4402 , P1_U4403 , P1_U4404 , P1_U4405;
wire P1_U4406 , P1_U4407 , P1_U4408 , P1_U4409 , P1_U4410 , P1_U4411 , P1_U4412 , P1_U4413 , P1_U4414 , P1_U4415;
wire P1_U4416 , P1_U4417 , P1_U4418 , P1_U4419 , P1_U4420 , P1_U4421 , P1_U4422 , P1_U4423 , P1_U4424 , P1_U4425;
wire P1_U4426 , P1_U4427 , P1_U4428 , P1_U4429 , P1_U4430 , P1_U4431 , P1_U4432 , P1_U4433 , P1_U4434 , P1_U4435;
wire P1_U4436 , P1_U4437 , P1_U4438 , P1_U4439 , P1_U4440 , P1_U4441 , P1_U4442 , P1_U4443 , P1_U4444 , P1_U4445;
wire P1_U4446 , P1_U4447 , P1_U4448 , P1_U4449 , P1_U4450 , P1_U4451 , P1_U4452 , P1_U4453 , P1_U4454 , P1_U4455;
wire P1_U4456 , P1_U4457 , P1_U4458 , P1_U4459 , P1_U4460 , P1_U4461 , P1_U4462 , P1_U4463 , P1_U4464 , P1_U4465;
wire P1_U4466 , P1_U4467 , P1_U4468 , P1_U4469 , P1_U4470 , P1_U4471 , P1_U4472 , P1_U4473 , P1_U4474 , P1_U4475;
wire P1_U4476 , P1_U4477 , P1_U4478 , P1_U4479 , P1_U4480 , P1_U4481 , P1_U4482 , P1_U4483 , P1_U4484 , P1_U4485;
wire P1_U4486 , P1_U4487 , P1_U4488 , P1_U4489 , P1_U4490 , P1_U4491 , P1_U4492 , P1_U4493 , P1_U4494 , P1_U4495;
wire P1_U4496 , P1_U4497 , P1_U4498 , P1_U4499 , P1_U4500 , P1_U4501 , P1_U4502 , P1_U4503 , P1_U4504 , P1_U4505;
wire P1_U4506 , P1_U4507 , P1_U4508 , P1_U4509 , P1_U4510 , P1_U4511 , P1_U4512 , P1_U4513 , P1_U4514 , P1_U4515;
wire P1_U4516 , P1_U4517 , P1_U4518 , P1_U4519 , P1_U4520 , P1_U4521 , P1_U4522 , P1_U4523 , P1_U4524 , P1_U4525;
wire P1_U4526 , P1_U4527 , P1_U4528 , P1_U4529 , P1_U4530 , P1_U4531 , P1_U4532 , P1_U4533 , P1_U4534 , P1_U4535;
wire P1_U4536 , P1_U4537 , P1_U4538 , P1_U4539 , P1_U4540 , P1_U4541 , P1_U4542 , P1_U4543 , P1_U4544 , P1_U4545;
wire P1_U4546 , P1_U4547 , P1_U4548 , P1_U4549 , P1_U4550 , P1_U4551 , P1_U4552 , P1_U4553 , P1_U4554 , P1_U4555;
wire P1_U4556 , P1_U4557 , P1_U4558 , P1_U4559 , P1_U4560 , P1_U4561 , P1_U4562 , P1_U4563 , P1_U4564 , P1_U4565;
wire P1_U4566 , P1_U4567 , P1_U4568 , P1_U4569 , P1_U4570 , P1_U4571 , P1_U4572 , P1_U4573 , P1_U4574 , P1_U4575;
wire P1_U4576 , P1_U4577 , P1_U4578 , P1_U4579 , P1_U4580 , P1_U4581 , P1_U4582 , P1_U4583 , P1_U4584 , P1_U4585;
wire P1_U4586 , P1_U4587 , P1_U4588 , P1_U4589 , P1_U4590 , P1_U4591 , P1_U4592 , P1_U4593 , P1_U4594 , P1_U4595;
wire P1_U4596 , P1_U4597 , P1_U4598 , P1_U4599 , P1_U4600 , P1_U4601 , P1_U4602 , P1_U4603 , P1_U4604 , P1_U4605;
wire P1_U4606 , P1_U4607 , P1_U4608 , P1_U4609 , P1_U4610 , P1_U4611 , P1_U4612 , P1_U4613 , P1_U4614 , P1_U4615;
wire P1_U4616 , P1_U4617 , P1_U4618 , P1_U4619 , P1_U4620 , P1_U4621 , P1_U4622 , P1_U4623 , P1_U4624 , P1_U4625;
wire P1_U4626 , P1_U4627 , P1_U4628 , P1_U4629 , P1_U4630 , P1_U4631 , P1_U4632 , P1_U4633 , P1_U4634 , P1_U4635;
wire P1_U4636 , P1_U4637 , P1_U4638 , P1_U4639 , P1_U4640 , P1_U4641 , P1_U4642 , P1_U4643 , P1_U4644 , P1_U4645;
wire P1_U4646 , P1_U4647 , P1_U4648 , P1_U4649 , P1_U4650 , P1_U4651 , P1_U4652 , P1_U4653 , P1_U4654 , P1_U4655;
wire P1_U4656 , P1_U4657 , P1_U4658 , P1_U4659 , P1_U4660 , P1_U4661 , P1_U4662 , P1_U4663 , P1_U4664 , P1_U4665;
wire P1_U4666 , P1_U4667 , P1_U4668 , P1_U4669 , P1_U4670 , P1_U4671 , P1_U4672 , P1_U4673 , P1_U4674 , P1_U4675;
wire P1_U4676 , P1_U4677 , P1_U4678 , P1_U4679 , P1_U4680 , P1_U4681 , P1_U4682 , P1_U4683 , P1_U4684 , P1_U4685;
wire P1_U4686 , P1_U4687 , P1_U4688 , P1_U4689 , P1_U4690 , P1_U4691 , P1_U4692 , P1_U4693 , P1_U4694 , P1_U4695;
wire P1_U4696 , P1_U4697 , P1_U4698 , P1_U4699 , P1_U4700 , P1_U4701 , P1_U4702 , P1_U4703 , P1_U4704 , P1_U4705;
wire P1_U4706 , P1_U4707 , P1_U4708 , P1_U4709 , P1_U4710 , P1_U4711 , P1_U4712 , P1_U4713 , P1_U4714 , P1_U4715;
wire P1_U4716 , P1_U4717 , P1_U4718 , P1_U4719 , P1_U4720 , P1_U4721 , P1_U4722 , P1_U4723 , P1_U4724 , P1_U4725;
wire P1_U4726 , P1_U4727 , P1_U4728 , P1_U4729 , P1_U4730 , P1_U4731 , P1_U4732 , P1_U4733 , P1_U4734 , P1_U4735;
wire P1_U4736 , P1_U4737 , P1_U4738 , P1_U4739 , P1_U4740 , P1_U4741 , P1_U4742 , P1_U4743 , P1_U4744 , P1_U4745;
wire P1_U4746 , P1_U4747 , P1_U4748 , P1_U4749 , P1_U4750 , P1_U4751 , P1_U4752 , P1_U4753 , P1_U4754 , P1_U4755;
wire P1_U4756 , P1_U4757 , P1_U4758 , P1_U4759 , P1_U4760 , P1_U4761 , P1_U4762 , P1_U4763 , P1_U4764 , P1_U4765;
wire P1_U4766 , P1_U4767 , P1_U4768 , P1_U4769 , P1_U4770 , P1_U4771 , P1_U4772 , P1_U4773 , P1_U4774 , P1_U4775;
wire P1_U4776 , P1_U4777 , P1_U4778 , P1_U4779 , P1_U4780 , P1_U4781 , P1_U4782 , P1_U4783 , P1_U4784 , P1_U4785;
wire P1_U4786 , P1_U4787 , P1_U4788 , P1_U4789 , P1_U4790 , P1_U4791 , P1_U4792 , P1_U4793 , P1_U4794 , P1_U4795;
wire P1_U4796 , P1_U4797 , P1_U4798 , P1_U4799 , P1_U4800 , P1_U4801 , P1_U4802 , P1_U4803 , P1_U4804 , P1_U4805;
wire P1_U4806 , P1_U4807 , P1_U4808 , P1_U4809 , P1_U4810 , P1_U4811 , P1_U4812 , P1_U4813 , P1_U4814 , P1_U4815;
wire P1_U4816 , P1_U4817 , P1_U4818 , P1_U4819 , P1_U4820 , P1_U4821 , P1_U4822 , P1_U4823 , P1_U4824 , P1_U4825;
wire P1_U4826 , P1_U4827 , P1_U4828 , P1_U4829 , P1_U4830 , P1_U4831 , P1_U4832 , P1_U4833 , P1_U4834 , P1_U4835;
wire P1_U4836 , P1_U4837 , P1_U4838 , P1_U4839 , P1_U4840 , P1_U4841 , P1_U4842 , P1_U4843 , P1_U4844 , P1_U4845;
wire P1_U4846 , P1_U4847 , P1_U4848 , P1_U4849 , P1_U4850 , P1_U4851 , P1_U4852 , P1_U4853 , P1_U4854 , P1_U4855;
wire P1_U4856 , P1_U4857 , P1_U4858 , P1_U4859 , P1_U4860 , P1_U4861 , P1_U4862 , P1_U4863 , P1_U4864 , P1_U4865;
wire P1_U4866 , P1_U4867 , P1_U4868 , P1_U4869 , P1_U4870 , P1_U4871 , P1_U4872 , P1_U4873 , P1_U4874 , P1_U4875;
wire P1_U4876 , P1_U4877 , P1_U4878 , P1_U4879 , P1_U4880 , P1_U4881 , P1_U4882 , P1_U4883 , P1_U4884 , P1_U4885;
wire P1_U4886 , P1_U4887 , P1_U4888 , P1_U4889 , P1_U4890 , P1_U4891 , P1_U4892 , P1_U4893 , P1_U4894 , P1_U4895;
wire P1_U4896 , P1_U4897 , P1_U4898 , P1_U4899 , P1_U4900 , P1_U4901 , P1_U4902 , P1_U4903 , P1_U4904 , P1_U4905;
wire P1_U4906 , P1_U4907 , P1_U4908 , P1_U4909 , P1_U4910 , P1_U4911 , P1_U4912 , P1_U4913 , P1_U4914 , P1_U4915;
wire P1_U4916 , P1_U4917 , P1_U4918 , P1_U4919 , P1_U4920 , P1_U4921 , P1_U4922 , P1_U4923 , P1_U4924 , P1_U4925;
wire P1_U4926 , P1_U4927 , P1_U4928 , P1_U4929 , P1_U4930 , P1_U4931 , P1_U4932 , P1_U4933 , P1_U4934 , P1_U4935;
wire P1_U4936 , P1_U4937 , P1_U4938 , P1_U4939 , P1_U4940 , P1_U4941 , P1_U4942 , P1_U4943 , P1_U4944 , P1_U4945;
wire P1_U4946 , P1_U4947 , P1_U4948 , P1_U4949 , P1_U4950 , P1_U4951 , P1_U4952 , P1_U4953 , P1_U4954 , P1_U4955;
wire P1_U4956 , P1_U4957 , P1_U4958 , P1_U4959 , P1_U4960 , P1_U4961 , P1_U4962 , P1_U4963 , P1_U4964 , P1_U4965;
wire P1_U4966 , P1_U4967 , P1_U4968 , P1_U4969 , P1_U4970 , P1_U4971 , P1_U4972 , P1_U4973 , P1_U4974 , P1_U4975;
wire P1_U4976 , P1_U4977 , P1_U4978 , P1_U4979 , P1_U4980 , P1_U4981 , P1_U4982 , P1_U4983 , P1_U4984 , P1_U4985;
wire P1_U4986 , P1_U4987 , P1_U4988 , P1_U4989 , P1_U4990 , P1_U4991 , P1_U4992 , P1_U4993 , P1_U4994 , P1_U4995;
wire P1_U4996 , P1_U4997 , P1_U4998 , P1_U4999 , P1_U5000 , P1_U5001 , P1_U5002 , P1_U5003 , P1_U5004 , P1_U5005;
wire P1_U5006 , P1_U5007 , P1_U5008 , P1_U5009 , P1_U5010 , P1_U5011 , P1_U5012 , P1_U5013 , P1_U5014 , P1_U5015;
wire P1_U5016 , P1_U5017 , P1_U5018 , P1_U5019 , P1_U5020 , P1_U5021 , P1_U5022 , P1_U5023 , P1_U5024 , P1_U5025;
wire P1_U5026 , P1_U5027 , P1_U5028 , P1_U5029 , P1_U5030 , P1_U5031 , P1_U5032 , P1_U5033 , P1_U5034 , P1_U5035;
wire P1_U5036 , P1_U5037 , P1_U5038 , P1_U5039 , P1_U5040 , P1_U5041 , P1_U5042 , P1_U5043 , P1_U5044 , P1_U5045;
wire P1_U5046 , P1_U5047 , P1_U5048 , P1_U5049 , P1_U5050 , P1_U5051 , P1_U5052 , P1_U5053 , P1_U5054 , P1_U5055;
wire P1_U5056 , P1_U5057 , P1_U5058 , P1_U5059 , P1_U5060 , P1_U5061 , P1_U5062 , P1_U5063 , P1_U5064 , P1_U5065;
wire P1_U5066 , P1_U5067 , P1_U5068 , P1_U5069 , P1_U5070 , P1_U5071 , P1_U5072 , P1_U5073 , P1_U5074 , P1_U5075;
wire P1_U5076 , P1_U5077 , P1_U5078 , P1_U5079 , P1_U5080 , P1_U5081 , P1_U5082 , P1_U5083 , P1_U5084 , P1_U5085;
wire P1_U5086 , P1_U5087 , P1_U5088 , P1_U5089 , P1_U5090 , P1_U5091 , P1_U5092 , P1_U5093 , P1_U5094 , P1_U5095;
wire P1_U5096 , P1_U5097 , P1_U5098 , P1_U5099 , P1_U5100 , P1_U5101 , P1_U5102 , P1_U5103 , P1_U5104 , P1_U5105;
wire P1_U5106 , P1_U5107 , P1_U5108 , P1_U5109 , P1_U5110 , P1_U5111 , P1_U5112 , P1_U5113 , P1_U5114 , P1_U5115;
wire P1_U5116 , P1_U5117 , P1_U5118 , P1_U5119 , P1_U5120 , P1_U5121 , P1_U5122 , P1_U5123 , P1_U5124 , P1_U5125;
wire P1_U5126 , P1_U5127 , P1_U5128 , P1_U5129 , P1_U5130 , P1_U5131 , P1_U5132 , P1_U5133 , P1_U5134 , P1_U5135;
wire P1_U5136 , P1_U5137 , P1_U5138 , P1_U5139 , P1_U5140 , P1_U5141 , P1_U5142 , P1_U5143 , P1_U5144 , P1_U5145;
wire P1_U5146 , P1_U5147 , P1_U5148 , P1_U5149 , P1_U5150 , P1_U5151 , P1_U5152 , P1_U5153 , P1_U5154 , P1_U5155;
wire P1_U5156 , P1_U5157 , P1_U5158 , P1_U5159 , P1_U5160 , P1_U5161 , P1_U5162 , P1_U5163 , P1_U5164 , P1_U5165;
wire P1_U5166 , P1_U5167 , P1_U5168 , P1_U5169 , P1_U5170 , P1_U5171 , P1_U5172 , P1_U5173 , P1_U5174 , P1_U5175;
wire P1_U5176 , P1_U5177 , P1_U5178 , P1_U5179 , P1_U5180 , P1_U5181 , P1_U5182 , P1_U5183 , P1_U5184 , P1_U5185;
wire P1_U5186 , P1_U5187 , P1_U5188 , P1_U5189 , P1_U5190 , P1_U5191 , P1_U5192 , P1_U5193 , P1_U5194 , P1_U5195;
wire P1_U5196 , P1_U5197 , P1_U5198 , P1_U5199 , P1_U5200 , P1_U5201 , P1_U5202 , P1_U5203 , P1_U5204 , P1_U5205;
wire P1_U5206 , P1_U5207 , P1_U5208 , P1_U5209 , P1_U5210 , P1_U5211 , P1_U5212 , P1_U5213 , P1_U5214 , P1_U5215;
wire P1_U5216 , P1_U5217 , P1_U5218 , P1_U5219 , P1_U5220 , P1_U5221 , P1_U5222 , P1_U5223 , P1_U5224 , P1_U5225;
wire P1_U5226 , P1_U5227 , P1_U5228 , P1_U5229 , P1_U5230 , P1_U5231 , P1_U5232 , P1_U5233 , P1_U5234 , P1_U5235;
wire P1_U5236 , P1_U5237 , P1_U5238 , P1_U5239 , P1_U5240 , P1_U5241 , P1_U5242 , P1_U5243 , P1_U5244 , P1_U5245;
wire P1_U5246 , P1_U5247 , P1_U5248 , P1_U5249 , P1_U5250 , P1_U5251 , P1_U5252 , P1_U5253 , P1_U5254 , P1_U5255;
wire P1_U5256 , P1_U5257 , P1_U5258 , P1_U5259 , P1_U5260 , P1_U5261 , P1_U5262 , P1_U5263 , P1_U5264 , P1_U5265;
wire P1_U5266 , P1_U5267 , P1_U5268 , P1_U5269 , P1_U5270 , P1_U5271 , P1_U5272 , P1_U5273 , P1_U5274 , P1_U5275;
wire P1_U5276 , P1_U5277 , P1_U5278 , P1_U5279 , P1_U5280 , P1_U5281 , P1_U5282 , P1_U5283 , P1_U5284 , P1_U5285;
wire P1_U5286 , P1_U5287 , P1_U5288 , P1_U5289 , P1_U5290 , P1_U5291 , P1_U5292 , P1_U5293 , P1_U5294 , P1_U5295;
wire P1_U5296 , P1_U5297 , P1_U5298 , P1_U5299 , P1_U5300 , P1_U5301 , P1_U5302 , P1_U5303 , P1_U5304 , P1_U5305;
wire P1_U5306 , P1_U5307 , P1_U5308 , P1_U5309 , P1_U5310 , P1_U5311 , P1_U5312 , P1_U5313 , P1_U5314 , P1_U5315;
wire P1_U5316 , P1_U5317 , P1_U5318 , P1_U5319 , P1_U5320 , P1_U5321 , P1_U5322 , P1_U5323 , P1_U5324 , P1_U5325;
wire P1_U5326 , P1_U5327 , P1_U5328 , P1_U5329 , P1_U5330 , P1_U5331 , P1_U5332 , P1_U5333 , P1_U5334 , P1_U5335;
wire P1_U5336 , P1_U5337 , P1_U5338 , P1_U5339 , P1_U5340 , P1_U5341 , P1_U5342 , P1_U5343 , P1_U5344 , P1_U5345;
wire P1_U5346 , P1_U5347 , P1_U5348 , P1_U5349 , P1_U5350 , P1_U5351 , P1_U5352 , P1_U5353 , P1_U5354 , P1_U5355;
wire P1_U5356 , P1_U5357 , P1_U5358 , P1_U5359 , P1_U5360 , P1_U5361 , P1_U5362 , P1_U5363 , P1_U5364 , P1_U5365;
wire P1_U5366 , P1_U5367 , P1_U5368 , P1_U5369 , P1_U5370 , P1_U5371 , P1_U5372 , P1_U5373 , P1_U5374 , P1_U5375;
wire P1_U5376 , P1_U5377 , P1_U5378 , P1_U5379 , P1_U5380 , P1_U5381 , P1_U5382 , P1_U5383 , P1_U5384 , P1_U5385;
wire P1_U5386 , P1_U5387 , P1_U5388 , P1_U5389 , P1_U5390 , P1_U5391 , P1_U5392 , P1_U5393 , P1_U5394 , P1_U5395;
wire P1_U5396 , P1_U5397 , P1_U5398 , P1_U5399 , P1_U5400 , P1_U5401 , P1_U5402 , P1_U5403 , P1_U5404 , P1_U5405;
wire P1_U5406 , P1_U5407 , P1_U5408 , P1_U5409 , P1_U5410 , P1_U5411 , P1_U5412 , P1_U5413 , P1_U5414 , P1_U5415;
wire P1_U5416 , P1_U5417 , P1_U5418 , P1_U5419 , P1_U5420 , P1_U5421 , P1_U5422 , P1_U5423 , P1_U5424 , P1_U5425;
wire P1_U5426 , P1_U5427 , P1_U5428 , P1_U5429 , P1_U5430 , P1_U5431 , P1_U5432 , P1_U5433 , P1_U5434 , P1_U5435;
wire P1_U5436 , P1_U5437 , P1_U5438 , P1_U5439 , P1_U5440 , P1_U5441 , P1_U5442 , P1_U5443 , P1_U5444 , P1_U5445;
wire P1_U5446 , P1_U5447 , P1_U5448 , P1_U5449 , P1_U5450 , P1_U5451 , P1_U5452 , P1_U5453 , P1_U5454 , P1_U5455;
wire P1_U5456 , P1_U5457 , P1_U5458 , P1_U5459 , P1_U5460 , P1_U5461 , P1_U5462 , P1_U5463 , P1_U5464 , P1_U5465;
wire P1_U5466 , P1_U5467 , P1_U5468 , P1_U5469 , P1_U5470 , P1_U5471 , P1_U5472 , P1_U5473 , P1_U5474 , P1_U5475;
wire P1_U5476 , P1_U5477 , P1_U5478 , P1_U5479 , P1_U5480 , P1_U5481 , P1_U5482 , P1_U5483 , P1_U5484 , P1_U5485;
wire P1_U5486 , P1_U5487 , P1_U5488 , P1_U5489 , P1_U5490 , P1_U5491 , P1_U5492 , P1_U5493 , P1_U5494 , P1_U5495;
wire P1_U5496 , P1_U5497 , P1_U5498 , P1_U5499 , P1_U5500 , P1_U5501 , P1_U5502 , P1_U5503 , P1_U5504 , P1_U5505;
wire P1_U5506 , P1_U5507 , P1_U5508 , P1_U5509 , P1_U5510 , P1_U5511 , P1_U5512 , P1_U5513 , P1_U5514 , P1_U5515;
wire P1_U5516 , P1_U5517 , P1_U5518 , P1_U5519 , P1_U5520 , P1_U5521 , P1_U5522 , P1_U5523 , P1_U5524 , P1_U5525;
wire P1_U5526 , P1_U5527 , P1_U5528 , P1_U5529 , P1_U5530 , P1_U5531 , P1_U5532 , P1_U5533 , P1_U5534 , P1_U5535;
wire P1_U5536 , P1_U5537 , P1_U5538 , P1_U5539 , P1_U5540 , P1_U5541 , P1_U5542 , P1_U5543 , P1_U5544 , P1_U5545;
wire P1_U5546 , P1_U5547 , P1_U5548 , P1_U5549 , P1_U5550 , P1_U5551 , P1_U5552 , P1_U5553 , P1_U5554 , P1_U5555;
wire P1_U5556 , P1_U5557 , P1_U5558 , P1_U5559 , P1_U5560 , P1_U5561 , P1_U5562 , P1_U5563 , P1_U5564 , P1_U5565;
wire P1_U5566 , P1_U5567 , P1_U5568 , P1_U5569 , P1_U5570 , P1_U5571 , P1_U5572 , P1_U5573 , P1_U5574 , P1_U5575;
wire P1_U5576 , P1_U5577 , P1_U5578 , P1_U5579 , P1_U5580 , P1_U5581 , P1_U5582 , P1_U5583 , P1_U5584 , P1_U5585;
wire P1_U5586 , P1_U5587 , P1_U5588 , P1_U5589 , P1_U5590 , P1_U5591 , P1_U5592 , P1_U5593 , P1_U5594 , P1_U5595;
wire P1_U5596 , P1_U5597 , P1_U5598 , P1_U5599 , P1_U5600 , P1_U5601 , P1_U5602 , P1_U5603 , P1_U5604 , P1_U5605;
wire P1_U5606 , P1_U5607 , P1_U5608 , P1_U5609 , P1_U5610 , P1_U5611 , P1_U5612 , P1_U5613 , P1_U5614 , P1_U5615;
wire P1_U5616 , P1_U5617 , P1_U5618 , P1_U5619 , P1_U5620 , P1_U5621 , P1_U5622 , P1_U5623 , P1_U5624 , P1_U5625;
wire P1_U5626 , P1_U5627 , P1_U5628 , P1_U5629 , P1_U5630 , P1_U5631 , P1_U5632 , P1_U5633 , P1_U5634 , P1_U5635;
wire P1_U5636 , P1_U5637 , P1_U5638 , P1_U5639 , P1_U5640 , P1_U5641 , P1_U5642 , P1_U5643 , P1_U5644 , P1_U5645;
wire P1_U5646 , P1_U5647 , P1_U5648 , P1_U5649 , P1_U5650 , P1_U5651 , P1_U5652 , P1_U5653 , P1_U5654 , P1_U5655;
wire P1_U5656 , P1_U5657 , P1_U5658 , P1_U5659 , P1_U5660 , P1_U5661 , P1_U5662 , P1_U5663 , P1_U5664 , P1_U5665;
wire P1_U5666 , P1_U5667 , P1_U5668 , P1_U5669 , P1_U5670 , P1_U5671 , P1_U5672 , P1_U5673 , P1_U5674 , P1_U5675;
wire P1_U5676 , P1_U5677 , P1_U5678 , P1_U5679 , P1_U5680 , P1_U5681 , P1_U5682 , P1_U5683 , P1_U5684 , P1_U5685;
wire P1_U5686 , P1_U5687 , P1_U5688 , P1_U5689 , P1_U5690 , P1_U5691 , P1_U5692 , P1_U5693 , P1_U5694 , P1_U5695;
wire P1_U5696 , P1_U5697 , P1_U5698 , P1_U5699 , P1_U5700 , P1_U5701 , P1_U5702 , P1_U5703 , P1_U5704 , P1_U5705;
wire P1_U5706 , P1_U5707 , P1_U5708 , P1_U5709 , P1_U5710 , P1_U5711 , P1_U5712 , P1_U5713 , P1_U5714 , P1_U5715;
wire P1_U5716 , P1_U5717 , P1_U5718 , P1_U5719 , P1_U5720 , P1_U5721 , P1_U5722 , P1_U5723 , P1_U5724 , P1_U5725;
wire P1_U5726 , P1_U5727 , P1_U5728 , P1_U5729 , P1_U5730 , P1_U5731 , P1_U5732 , P1_U5733 , P1_U5734 , P1_U5735;
wire P1_U5736 , P1_U5737 , P1_U5738 , P1_U5739 , P1_U5740 , P1_U5741 , P1_U5742 , P1_U5743 , P1_U5744 , P1_U5745;
wire P1_U5746 , P1_U5747 , P1_U5748 , P1_U5749 , P1_U5750 , P1_U5751 , P1_U5752 , P1_U5753 , P1_U5754 , P1_U5755;
wire P1_U5756 , P1_U5757 , P1_U5758 , P1_U5759 , P1_U5760 , P1_U5761 , P1_U5762 , P1_U5763 , P1_U5764 , P1_U5765;
wire P1_U5766 , P1_U5767 , P1_U5768 , P1_U5769 , P1_U5770 , P1_U5771 , P1_U5772 , P1_U5773 , P1_U5774 , P1_U5775;
wire P1_U5776 , P1_U5777 , P1_U5778 , P1_U5779 , P1_U5780 , P1_U5781 , P1_U5782 , P1_U5783 , P1_U5784 , P1_U5785;
wire P1_U5786 , P1_U5787 , P1_U5788 , P1_U5789 , P1_U5790 , P1_U5791 , P1_U5792 , P1_U5793 , P1_U5794 , P1_U5795;
wire P1_U5796 , P1_U5797 , P1_U5798 , P1_U5799 , P1_U5800 , P1_U5801 , P1_U5802 , P1_U5803 , P1_U5804 , P1_U5805;
wire P1_U5806 , P1_U5807 , P1_U5808 , P1_U5809 , P1_U5810 , P1_U5811 , P1_U5812 , P1_U5813 , P1_U5814 , P1_U5815;
wire P1_U5816 , P1_U5817 , P1_U5818 , P1_U5819 , P1_U5820 , P1_U5821 , P1_U5822 , P1_U5823 , P1_U5824 , P1_U5825;
wire P1_U5826 , P1_U5827 , P1_U5828 , P1_U5829 , P1_U5830 , P1_U5831 , P1_U5832 , P1_U5833 , P1_U5834 , P1_U5835;
wire P1_U5836 , P1_U5837 , P1_U5838 , P1_U5839 , P1_U5840 , P1_U5841 , P1_U5842 , P1_U5843 , P1_U5844 , P1_U5845;
wire P1_U5846 , P1_U5847 , P1_U5848 , P1_U5849 , P1_U5850 , P1_U5851 , P1_U5852 , P1_U5853 , P1_U5854 , P1_U5855;
wire P1_U5856 , P1_U5857 , P1_U5858 , P1_U5859 , P1_U5860 , P1_U5861 , P1_U5862 , P1_U5863 , P1_U5864 , P1_U5865;
wire P1_U5866 , P1_U5867 , P1_U5868 , P1_U5869 , P1_U5870 , P1_U5871 , P1_U5872 , P1_U5873 , P1_U5874 , P1_U5875;
wire P1_U5876 , P1_U5877 , P1_U5878 , P1_U5879 , P1_U5880 , P1_U5881 , P1_U5882 , P1_U5883 , P1_U5884 , P1_U5885;
wire P1_U5886 , P1_U5887 , P1_U5888 , P1_U5889 , P1_U5890 , P1_U5891 , P1_U5892 , P1_U5893 , P1_U5894 , P1_U5895;
wire P1_U5896 , P1_U5897 , P1_U5898 , P1_U5899 , P1_U5900 , P1_U5901 , P1_U5902 , P1_U5903 , P1_U5904 , P1_U5905;
wire P1_U5906 , P1_U5907 , P1_U5908 , P1_U5909 , P1_U5910 , P1_U5911 , P1_U5912 , P1_U5913 , P1_U5914 , P1_U5915;
wire P1_U5916 , P1_U5917 , P1_U5918 , P1_U5919 , P1_U5920 , P1_U5921 , P1_U5922 , P1_U5923 , P1_U5924 , P1_U5925;
wire P1_U5926 , P1_U5927 , P1_U5928 , P1_U5929 , P1_U5930 , P1_U5931 , P1_U5932 , P1_U5933 , P1_U5934 , P1_U5935;
wire P1_U5936 , P1_U5937 , P1_U5938 , P1_U5939 , P1_U5940 , P1_U5941 , P1_U5942 , P1_U5943 , P1_U5944 , P1_U5945;
wire P1_U5946 , P1_U5947 , P1_U5948 , P1_U5949 , P1_U5950 , P1_U5951 , P1_U5952 , P1_U5953 , P1_U5954 , P1_U5955;
wire P1_U5956 , P1_U5957 , P1_U5958 , P1_U5959 , P1_U5960 , P1_U5961 , P1_U5962 , P1_U5963 , P1_U5964 , P1_U5965;
wire P1_U5966 , P1_U5967 , P1_U5968 , P1_U5969 , P1_U5970 , P1_U5971 , P1_U5972 , P1_U5973 , P1_U5974 , P1_U5975;
wire P1_U5976 , P1_U5977 , P1_U5978 , P1_U5979 , P1_U5980 , P1_U5981 , P1_U5982 , P1_U5983 , P1_U5984 , P1_U5985;
wire P1_U5986 , P1_U5987 , P1_U5988 , P1_U5989 , P1_U5990 , P1_U5991 , P1_U5992 , P1_U5993 , P1_U5994 , P1_U5995;
wire P1_U5996 , P1_U5997 , P1_U5998 , P1_U5999 , P1_U6000 , P1_U6001 , P1_U6002 , P1_U6003 , P1_U6004 , P1_U6005;
wire P1_U6006 , P1_U6007 , P1_U6008 , P1_U6009 , P1_U6010 , P1_U6011 , P1_U6012 , P1_U6013 , P1_U6014 , P1_U6015;
wire P1_U6016 , P1_U6017 , P1_U6018 , P1_U6019 , P1_U6020 , P1_U6021 , P1_U6022 , P1_U6023 , P1_U6024 , P1_U6025;
wire P1_U6026 , P1_U6027 , P1_U6028 , P1_U6029 , P1_U6030 , P1_U6031 , P1_U6032 , P1_U6033 , P1_U6034 , P1_U6035;
wire P1_U6036 , P1_U6037 , P1_U6038 , P1_U6039 , P1_U6040 , P1_U6041 , P1_U6042 , P1_U6043 , P1_U6044 , P1_U6045;
wire P1_U6046 , P1_U6047 , P1_U6048 , P1_U6049 , P1_U6050 , P1_U6051 , P1_U6052 , P1_U6053 , P1_U6054 , P1_U6055;
wire P1_U6056 , P1_U6057 , P1_U6058 , P1_U6059 , P1_U6060 , P1_U6061 , P1_U6062 , P1_U6063 , P1_U6064 , P1_U6065;
wire P1_U6066 , P1_U6067 , P1_U6068 , P1_U6069 , P1_U6070 , P1_U6071 , P1_U6072 , P1_U6073 , P1_U6074 , P1_U6075;
wire P1_U6076 , P1_U6077 , P1_U6078 , P1_U6079 , P1_U6080 , P1_U6081 , P1_U6082 , P1_U6083 , P1_U6084 , P1_U6085;
wire P1_U6086 , P1_U6087 , P1_U6088 , P1_U6089 , P1_U6090 , P1_U6091 , P1_U6092 , P1_U6093 , P1_U6094 , P1_U6095;
wire P1_U6096 , P1_U6097 , P1_U6098 , P1_U6099 , P1_U6100 , P1_U6101 , P1_U6102 , P1_U6103 , P1_U6104 , P1_U6105;
wire P1_U6106 , P1_U6107 , P1_U6108 , P1_U6109 , P1_U6110 , P1_U6111 , P1_U6112 , P1_U6113 , P1_U6114 , P1_U6115;
wire P1_U6116 , P1_U6117 , P1_U6118 , P1_U6119 , P1_U6120 , P1_U6121 , P1_U6122 , P1_U6123 , P1_U6124 , P1_U6125;
wire P1_U6126 , P1_U6127 , P1_U6128 , P1_U6129 , P1_U6130 , P1_U6131 , P1_U6132 , P1_U6133 , P1_U6134 , P1_U6135;
wire P1_U6136 , P1_U6137 , P1_U6138 , P1_U6139 , P1_U6140 , P1_U6141 , P1_U6142 , P1_U6143 , P1_U6144 , P1_U6145;
wire P1_U6146 , P1_U6147 , P1_U6148 , P1_U6149 , P1_U6150 , P1_U6151 , P1_U6152 , P1_U6153 , P1_U6154 , P1_U6155;
wire P1_U6156 , P1_U6157 , P1_U6158 , P1_U6159 , P1_U6160 , P1_U6161 , P1_U6162 , P1_U6163 , P1_U6164 , P1_U6165;
wire P1_U6166 , P1_U6167 , P1_U6168 , P1_U6169 , P1_U6170 , P1_U6171 , P1_U6172 , P1_U6173 , P1_U6174 , P1_U6175;
wire P1_U6176 , P1_U6177 , P1_U6178 , P1_U6179 , P1_U6180 , P1_U6181 , P1_U6182 , P1_U6183 , P1_U6184 , P1_U6185;
wire P1_U6186 , P1_U6187 , P1_U6188 , P1_U6189 , P1_U6190 , P1_U6191 , P1_U6192 , P1_U6193 , P1_U6194 , P1_U6195;
wire P1_U6196 , P1_U6197 , P1_U6198 , P1_U6199 , P1_U6200 , P1_U6201 , P1_U6202 , P1_U6203 , P1_U6204 , P1_U6205;
wire P1_U6206 , P1_U6207 , P1_U6208 , P1_U6209 , P1_U6210 , P1_U6211 , P1_U6212 , P1_U6213 , P1_U6214 , P1_U6215;
wire P1_U6216 , P1_U6217 , P1_U6218 , P1_U6219 , P1_U6220 , P1_U6221 , P1_U6222 , P1_U6223 , P1_U6224 , P1_U6225;
wire P1_U6226 , P1_U6227 , P1_U6228 , P1_U6229 , P1_U6230 , P1_U6231 , P1_U6232 , P1_U6233 , P1_U6234 , P1_U6235;
wire P1_U6236 , P1_U6237 , P1_U6238 , P1_U6239 , P1_U6240 , P1_U6241 , P1_U6242 , P1_U6243 , P1_U6244 , P1_U6245;
wire P1_U6246 , P1_U6247 , P1_U6248 , P1_U6249 , P1_U6250 , P1_U6251 , P1_U6252 , P1_U6253 , P1_U6254 , P1_U6255;
wire P1_U6256 , P1_U6257 , P1_U6258 , P1_U6259 , P1_U6260 , P1_U6261 , P1_U6262 , P1_U6263 , P1_U6264 , P1_U6265;
wire P1_U6266 , P1_U6267 , P1_U6268 , P1_U6269 , P1_U6270 , P1_U6271 , P1_U6272 , P1_U6273 , P1_U6274 , P1_U6275;
wire P1_U6276 , P1_U6277 , P1_U6278 , P1_U6279 , P1_U6280 , P1_U6281 , P1_U6282 , P1_U6283 , P1_U6284 , P1_U6285;
wire P3_R1161_U489 , P3_R1161_U488 , P3_R1161_U487 , P3_R1161_U486 , P3_R1161_U485 , P3_R1161_U484 , P3_R1161_U483 , P3_R1161_U482 , P3_R1161_U481 , P3_R1161_U480;
wire P3_R1161_U479 , P3_R1161_U478 , P3_R1161_U477 , P3_R1161_U476 , P3_R1161_U475 , P3_R1161_U474 , P3_R1161_U473 , P3_R1161_U472 , P3_R1161_U471 , P3_R1161_U470;
wire P3_R1161_U469 , P2_U3014 , P2_U3015 , P2_U3016 , P2_U3017 , P2_U3018 , P2_U3019 , P2_U3020 , P2_U3021 , P2_U3022;
wire P2_U3023 , P2_U3024 , P2_U3025 , P2_U3026 , P2_U3027 , P2_U3028 , P2_U3029 , P2_U3030 , P2_U3031 , P2_U3032;
wire P2_U3033 , P2_U3034 , P2_U3035 , P2_U3036 , P2_U3037 , P2_U3038 , P2_U3039 , P2_U3040 , P2_U3041 , P2_U3042;
wire P2_U3043 , P2_U3044 , P2_U3045 , P2_U3046 , P2_U3047 , P2_U3048 , P2_U3049 , P2_U3050 , P2_U3051 , P2_U3052;
wire P2_U3053 , P2_U3054 , P2_U3055 , P2_U3056 , P2_U3057 , P2_U3058 , P2_U3059 , P2_U3060 , P2_U3061 , P2_U3062;
wire P2_U3063 , P2_U3064 , P2_U3065 , P2_U3066 , P2_U3067 , P2_U3068 , P2_U3069 , P2_U3070 , P2_U3071 , P2_U3072;
wire P2_U3073 , P2_U3074 , P2_U3075 , P2_U3076 , P2_U3077 , P2_U3078 , P2_U3079 , P2_U3080 , P2_U3081 , P2_U3082;
wire P2_U3083 , P2_U3084 , P2_U3085 , P2_U3086 , P2_U3089 , P2_U3090 , P2_U3091 , P2_U3092 , P2_U3093 , P2_U3094;
wire P2_U3095 , P2_U3096 , P2_U3097 , P2_U3098 , P2_U3099 , P2_U3100 , P2_U3101 , P2_U3102 , P2_U3103 , P2_U3104;
wire P2_U3105 , P2_U3106 , P2_U3107 , P2_U3108 , P2_U3109 , P2_U3110 , P2_U3111 , P2_U3112 , P2_U3113 , P2_U3114;
wire P2_U3115 , P2_U3116 , P2_U3117 , P2_U3118 , P2_U3119 , P2_U3120 , P2_U3121 , P2_U3122 , P2_U3123 , P2_U3124;
wire P2_U3125 , P2_U3126 , P2_U3127 , P2_U3128 , P2_U3129 , P2_U3130 , P2_U3131 , P2_U3132 , P2_U3133 , P2_U3134;
wire P2_U3135 , P2_U3136 , P2_U3137 , P2_U3138 , P2_U3139 , P2_U3140 , P2_U3141 , P2_U3142 , P2_U3143 , P2_U3144;
wire P2_U3145 , P2_U3146 , P2_U3147 , P2_U3148 , P2_U3149 , P2_U3150 , P2_U3151 , P2_U3152 , P2_U3153 , P2_U3154;
wire P2_U3155 , P2_U3156 , P2_U3157 , P2_U3158 , P2_U3159 , P2_U3160 , P2_U3161 , P2_U3162 , P2_U3163 , P2_U3164;
wire P2_U3165 , P2_U3166 , P2_U3167 , P2_U3168 , P2_U3169 , P2_U3170 , P2_U3171 , P2_U3172 , P2_U3173 , P2_U3174;
wire P2_U3175 , P2_U3176 , P2_U3177 , P2_U3178 , P2_U3179 , P2_U3180 , P2_U3181 , P2_U3182 , P2_U3183 , P2_U3184;
wire P2_U3329 , P2_U3330 , P2_U3331 , P2_U3332 , P2_U3333 , P2_U3334 , P2_U3335 , P2_U3336 , P2_U3337 , P2_U3338;
wire P2_U3339 , P2_U3340 , P2_U3341 , P2_U3342 , P2_U3343 , P2_U3344 , P2_U3345 , P2_U3346 , P2_U3347 , P2_U3348;
wire P2_U3349 , P2_U3350 , P2_U3351 , P2_U3352 , P2_U3353 , P2_U3354 , P2_U3355 , P2_U3356 , P2_U3357 , P2_U3358;
wire P2_U3359 , P2_U3360 , P2_U3361 , P2_U3362 , P2_U3363 , P2_U3364 , P2_U3365 , P2_U3366 , P2_U3367 , P2_U3368;
wire P2_U3369 , P2_U3370 , P2_U3371 , P2_U3372 , P2_U3373 , P2_U3374 , P2_U3375 , P2_U3376 , P2_U3377 , P2_U3378;
wire P2_U3379 , P2_U3380 , P2_U3381 , P2_U3382 , P2_U3383 , P2_U3384 , P2_U3385 , P2_U3386 , P2_U3387 , P2_U3388;
wire P2_U3389 , P2_U3390 , P2_U3391 , P2_U3392 , P2_U3393 , P2_U3394 , P2_U3395 , P2_U3396 , P2_U3397 , P2_U3398;
wire P2_U3399 , P2_U3400 , P2_U3401 , P2_U3402 , P2_U3403 , P2_U3404 , P2_U3405 , P2_U3406 , P2_U3407 , P2_U3408;
wire P2_U3409 , P2_U3410 , P2_U3411 , P2_U3412 , P2_U3413 , P2_U3414 , P2_U3415 , P2_U3418 , P2_U3419 , P2_U3420;
wire P2_U3421 , P2_U3422 , P2_U3423 , P2_U3424 , P2_U3425 , P2_U3426 , P2_U3427 , P2_U3428 , P2_U3429 , P2_U3431;
wire P2_U3432 , P2_U3434 , P2_U3435 , P2_U3437 , P2_U3438 , P2_U3440 , P2_U3441 , P2_U3443 , P2_U3444 , P2_U3446;
wire P2_U3447 , P2_U3449 , P2_U3450 , P2_U3452 , P2_U3453 , P2_U3455 , P2_U3456 , P2_U3458 , P2_U3459 , P2_U3461;
wire P2_U3462 , P2_U3464 , P2_U3465 , P2_U3467 , P2_U3468 , P2_U3470 , P2_U3471 , P2_U3473 , P2_U3474 , P2_U3476;
wire P2_U3477 , P2_U3479 , P2_U3480 , P2_U3482 , P2_U3483 , P2_U3485 , P2_U3563 , P2_U3564 , P2_U3565 , P2_U3566;
wire P2_U3567 , P2_U3568 , P2_U3569 , P2_U3570 , P2_U3571 , P2_U3572 , P2_U3573 , P2_U3574 , P2_U3575 , P2_U3576;
wire P2_U3577 , P2_U3578 , P2_U3579 , P2_U3580 , P2_U3581 , P2_U3582 , P2_U3583 , P2_U3584 , P2_U3585 , P2_U3586;
wire P2_U3587 , P2_U3588 , P2_U3589 , P2_U3590 , P2_U3591 , P2_U3592 , P2_U3593 , P2_U3594 , P2_U3595 , P2_U3596;
wire P2_U3597 , P2_U3598 , P2_U3599 , P2_U3600 , P2_U3601 , P2_U3602 , P2_U3603 , P2_U3604 , P2_U3605 , P2_U3606;
wire P2_U3607 , P2_U3608 , P2_U3609 , P2_U3610 , P2_U3611 , P2_U3612 , P2_U3613 , P2_U3614 , P2_U3615 , P2_U3616;
wire P2_U3617 , P2_U3618 , P2_U3619 , P2_U3620 , P2_U3621 , P2_U3622 , P2_U3623 , P2_U3624 , P2_U3625 , P2_U3626;
wire P2_U3627 , P2_U3628 , P2_U3629 , P2_U3630 , P2_U3631 , P2_U3632 , P2_U3633 , P2_U3634 , P2_U3635 , P2_U3636;
wire P2_U3637 , P2_U3638 , P2_U3639 , P2_U3640 , P2_U3641 , P2_U3642 , P2_U3643 , P2_U3644 , P2_U3645 , P2_U3646;
wire P2_U3647 , P2_U3648 , P2_U3649 , P2_U3650 , P2_U3651 , P2_U3652 , P2_U3653 , P2_U3654 , P2_U3655 , P2_U3656;
wire P2_U3657 , P2_U3658 , P2_U3659 , P2_U3660 , P2_U3661 , P2_U3662 , P2_U3663 , P2_U3664 , P2_U3665 , P2_U3666;
wire P2_U3667 , P2_U3668 , P2_U3669 , P2_U3670 , P2_U3671 , P2_U3672 , P2_U3673 , P2_U3674 , P2_U3675 , P2_U3676;
wire P2_U3677 , P2_U3678 , P2_U3679 , P2_U3680 , P2_U3681 , P2_U3682 , P2_U3683 , P2_U3684 , P2_U3685 , P2_U3686;
wire P2_U3687 , P2_U3688 , P2_U3689 , P2_U3690 , P2_U3691 , P2_U3692 , P2_U3693 , P2_U3694 , P2_U3695 , P2_U3696;
wire P2_U3697 , P2_U3698 , P2_U3699 , P2_U3700 , P2_U3701 , P2_U3702 , P2_U3703 , P2_U3704 , P2_U3705 , P2_U3706;
wire P2_U3707 , P2_U3708 , P2_U3709 , P2_U3710 , P2_U3711 , P2_U3712 , P2_U3713 , P2_U3714 , P2_U3715 , P2_U3716;
wire P2_U3717 , P2_U3718 , P2_U3719 , P2_U3720 , P2_U3721 , P2_U3722 , P2_U3723 , P2_U3724 , P2_U3725 , P2_U3726;
wire P2_U3727 , P2_U3728 , P2_U3729 , P2_U3730 , P2_U3731 , P2_U3732 , P2_U3733 , P2_U3734 , P2_U3735 , P2_U3736;
wire P2_U3737 , P2_U3738 , P2_U3739 , P2_U3740 , P2_U3741 , P2_U3742 , P2_U3743 , P2_U3744 , P2_U3745 , P2_U3746;
wire P2_U3747 , P2_U3748 , P2_U3749 , P2_U3750 , P2_U3751 , P2_U3752 , P2_U3753 , P2_U3754 , P2_U3755 , P2_U3756;
wire P2_U3757 , P2_U3758 , P2_U3759 , P2_U3760 , P2_U3761 , P2_U3762 , P2_U3763 , P2_U3764 , P2_U3765 , P2_U3766;
wire P2_U3767 , P2_U3768 , P2_U3769 , P2_U3770 , P2_U3771 , P2_U3772 , P2_U3773 , P2_U3774 , P2_U3775 , P2_U3776;
wire P2_U3777 , P2_U3778 , P2_U3779 , P2_U3780 , P2_U3781 , P2_U3782 , P2_U3783 , P2_U3784 , P2_U3785 , P2_U3786;
wire P2_U3787 , P2_U3788 , P2_U3789 , P2_U3790 , P2_U3791 , P2_U3792 , P2_U3793 , P2_U3794 , P2_U3795 , P2_U3796;
wire P2_U3797 , P2_U3798 , P2_U3799 , P2_U3800 , P2_U3801 , P2_U3802 , P2_U3803 , P2_U3804 , P2_U3805 , P2_U3806;
wire P2_U3807 , P2_U3808 , P2_U3809 , P2_U3810 , P2_U3811 , P2_U3812 , P2_U3813 , P2_U3814 , P2_U3815 , P2_U3816;
wire P2_U3817 , P2_U3818 , P2_U3819 , P2_U3820 , P2_U3821 , P2_U3822 , P2_U3823 , P2_U3824 , P2_U3825 , P2_U3826;
wire P2_U3827 , P2_U3828 , P2_U3829 , P2_U3830 , P2_U3831 , P2_U3832 , P2_U3833 , P2_U3834 , P2_U3835 , P2_U3836;
wire P2_U3837 , P2_U3838 , P2_U3839 , P2_U3840 , P2_U3841 , P2_U3842 , P2_U3843 , P2_U3844 , P2_U3845 , P2_U3846;
wire P2_U3847 , P2_U3848 , P2_U3849 , P2_U3850 , P2_U3851 , P2_U3852 , P2_U3853 , P2_U3854 , P2_U3855 , P2_U3856;
wire P2_U3857 , P2_U3858 , P2_U3859 , P2_U3860 , P2_U3861 , P2_U3862 , P2_U3863 , P2_U3864 , P2_U3865 , P2_U3866;
wire P2_U3867 , P2_U3868 , P2_U3869 , P2_U3870 , P2_U3871 , P2_U3872 , P2_U3873 , P2_U3874 , P2_U3875 , P2_U3876;
wire P2_U3877 , P2_U3878 , P2_U3879 , P2_U3880 , P2_U3881 , P2_U3882 , P2_U3883 , P2_U3884 , P2_U3885 , P2_U3886;
wire P2_U3887 , P2_U3888 , P2_U3889 , P2_U3890 , P2_U3891 , P2_U3892 , P2_U3893 , P2_U3894 , P2_U3895 , P2_U3896;
wire P2_U3897 , P2_U3898 , P2_U3899 , P2_U3900 , P2_U3901 , P2_U3902 , P2_U3903 , P2_U3904 , P2_U3905 , P2_U3906;
wire P2_U3907 , P2_U3908 , P2_U3909 , P2_U3910 , P2_U3911 , P2_U3912 , P2_U3913 , P2_U3914 , P2_U3915 , P2_U3916;
wire P2_U3917 , P2_U3918 , P2_U3919 , P2_U3920 , P2_U3921 , P2_U3922 , P2_U3923 , P2_U3924 , P2_U3925 , P2_U3926;
wire P2_U3927 , P2_U3928 , P2_U3929 , P2_U3930 , P2_U3931 , P2_U3932 , P2_U3933 , P2_U3934 , P2_U3935 , P2_U3936;
wire P2_U3937 , P2_U3938 , P2_U3939 , P2_U3940 , P2_U3941 , P2_U3942 , P2_U3943 , P2_U3944 , P2_U3945 , P2_U3946;
wire P2_U3948 , P2_U3949 , P2_U3950 , P2_U3951 , P2_U3952 , P2_U3953 , P2_U3954 , P2_U3955 , P2_U3956 , P2_U3957;
wire P2_U3958 , P2_U3959 , P2_U3960 , P2_U3961 , P2_U3962 , P2_U3963 , P2_U3964 , P2_U3965 , P2_U3966 , P2_U3967;
wire P2_U3968 , P2_U3969 , P2_U3970 , P2_U3971 , P2_U3972 , P2_U3973 , P2_U3974 , P2_U3975 , P2_U3976 , P2_U3977;
wire P2_U3978 , P2_U3979 , P2_U3980 , P2_U3981 , P2_U3982 , P2_U3983 , P2_U3984 , P2_U3985 , P2_U3986 , P2_U3987;
wire P2_U3988 , P2_U3989 , P2_U3990 , P2_U3991 , P2_U3992 , P2_U3993 , P2_U3994 , P2_U3995 , P2_U3996 , P2_U3997;
wire P2_U3998 , P2_U3999 , P2_U4000 , P2_U4001 , P2_U4002 , P2_U4003 , P2_U4004 , P2_U4005 , P2_U4006 , P2_U4007;
wire P2_U4008 , P2_U4009 , P2_U4010 , P2_U4011 , P2_U4012 , P2_U4013 , P2_U4014 , P2_U4015 , P2_U4016 , P2_U4017;
wire P2_U4018 , P2_U4019 , P2_U4020 , P2_U4021 , P2_U4022 , P2_U4023 , P2_U4024 , P2_U4025 , P2_U4026 , P2_U4027;
wire P2_U4028 , P2_U4029 , P2_U4030 , P2_U4031 , P2_U4032 , P2_U4033 , P2_U4034 , P2_U4035 , P2_U4036 , P2_U4037;
wire P2_U4038 , P2_U4039 , P2_U4040 , P2_U4041 , P2_U4042 , P2_U4043 , P2_U4044 , P2_U4045 , P2_U4046 , P2_U4047;
wire P2_U4048 , P2_U4049 , P2_U4050 , P2_U4051 , P2_U4052 , P2_U4053 , P2_U4054 , P2_U4055 , P2_U4056 , P2_U4057;
wire P2_U4058 , P2_U4059 , P2_U4060 , P2_U4061 , P2_U4062 , P2_U4063 , P2_U4064 , P2_U4065 , P2_U4066 , P2_U4067;
wire P2_U4068 , P2_U4069 , P2_U4070 , P2_U4071 , P2_U4072 , P2_U4073 , P2_U4074 , P2_U4075 , P2_U4076 , P2_U4077;
wire P2_U4078 , P2_U4079 , P2_U4080 , P2_U4081 , P2_U4082 , P2_U4083 , P2_U4084 , P2_U4085 , P2_U4086 , P2_U4087;
wire P2_U4088 , P2_U4089 , P2_U4090 , P2_U4091 , P2_U4092 , P2_U4093 , P2_U4094 , P2_U4095 , P2_U4096 , P2_U4097;
wire P2_U4098 , P2_U4099 , P2_U4100 , P2_U4101 , P2_U4102 , P2_U4103 , P2_U4104 , P2_U4105 , P2_U4106 , P2_U4107;
wire P2_U4108 , P2_U4109 , P2_U4110 , P2_U4111 , P2_U4112 , P2_U4113 , P2_U4114 , P2_U4115 , P2_U4116 , P2_U4117;
wire P2_U4118 , P2_U4119 , P2_U4120 , P2_U4121 , P2_U4122 , P2_U4123 , P2_U4124 , P2_U4125 , P2_U4126 , P2_U4127;
wire P2_U4128 , P2_U4129 , P2_U4130 , P2_U4131 , P2_U4132 , P2_U4133 , P2_U4134 , P2_U4135 , P2_U4136 , P2_U4137;
wire P2_U4138 , P2_U4139 , P2_U4140 , P2_U4141 , P2_U4142 , P2_U4143 , P2_U4144 , P2_U4145 , P2_U4146 , P2_U4147;
wire P2_U4148 , P2_U4149 , P2_U4150 , P2_U4151 , P2_U4152 , P2_U4153 , P2_U4154 , P2_U4155 , P2_U4156 , P2_U4157;
wire P2_U4158 , P2_U4159 , P2_U4160 , P2_U4161 , P2_U4162 , P2_U4163 , P2_U4164 , P2_U4165 , P2_U4166 , P2_U4167;
wire P2_U4168 , P2_U4169 , P2_U4170 , P2_U4171 , P2_U4172 , P2_U4173 , P2_U4174 , P2_U4175 , P2_U4176 , P2_U4177;
wire P2_U4178 , P2_U4179 , P2_U4180 , P2_U4181 , P2_U4182 , P2_U4183 , P2_U4184 , P2_U4185 , P2_U4186 , P2_U4187;
wire P2_U4188 , P2_U4189 , P2_U4190 , P2_U4191 , P2_U4192 , P2_U4193 , P2_U4194 , P2_U4195 , P2_U4196 , P2_U4197;
wire P2_U4198 , P2_U4199 , P2_U4200 , P2_U4201 , P2_U4202 , P2_U4203 , P2_U4204 , P2_U4205 , P2_U4206 , P2_U4207;
wire P2_U4208 , P2_U4209 , P2_U4210 , P2_U4211 , P2_U4212 , P2_U4213 , P2_U4214 , P2_U4215 , P2_U4216 , P2_U4217;
wire P2_U4218 , P2_U4219 , P2_U4220 , P2_U4221 , P2_U4222 , P2_U4223 , P2_U4224 , P2_U4225 , P2_U4226 , P2_U4227;
wire P2_U4228 , P2_U4229 , P2_U4230 , P2_U4231 , P2_U4232 , P2_U4233 , P2_U4234 , P2_U4235 , P2_U4236 , P2_U4237;
wire P2_U4238 , P2_U4239 , P2_U4240 , P2_U4241 , P2_U4242 , P2_U4243 , P2_U4244 , P2_U4245 , P2_U4246 , P2_U4247;
wire P2_U4248 , P2_U4249 , P2_U4250 , P2_U4251 , P2_U4252 , P2_U4253 , P2_U4254 , P2_U4255 , P2_U4256 , P2_U4257;
wire P2_U4258 , P2_U4259 , P2_U4260 , P2_U4261 , P2_U4262 , P2_U4263 , P2_U4264 , P2_U4265 , P2_U4266 , P2_U4267;
wire P2_U4268 , P2_U4269 , P2_U4270 , P2_U4271 , P2_U4272 , P2_U4273 , P2_U4274 , P2_U4275 , P2_U4276 , P2_U4277;
wire P2_U4278 , P2_U4279 , P2_U4280 , P2_U4281 , P2_U4282 , P2_U4283 , P2_U4284 , P2_U4285 , P2_U4286 , P2_U4287;
wire P2_U4288 , P2_U4289 , P2_U4290 , P2_U4291 , P2_U4292 , P2_U4293 , P2_U4294 , P2_U4295 , P2_U4296 , P2_U4297;
wire P2_U4298 , P2_U4299 , P2_U4300 , P2_U4301 , P2_U4302 , P2_U4303 , P2_U4304 , P2_U4305 , P2_U4306 , P2_U4307;
wire P2_U4308 , P2_U4309 , P2_U4310 , P2_U4311 , P2_U4312 , P2_U4313 , P2_U4314 , P2_U4315 , P2_U4316 , P2_U4317;
wire P2_U4318 , P2_U4319 , P2_U4320 , P2_U4321 , P2_U4322 , P2_U4323 , P2_U4324 , P2_U4325 , P2_U4326 , P2_U4327;
wire P2_U4328 , P2_U4329 , P2_U4330 , P2_U4331 , P2_U4332 , P2_U4333 , P2_U4334 , P2_U4335 , P2_U4336 , P2_U4337;
wire P2_U4338 , P2_U4339 , P2_U4340 , P2_U4341 , P2_U4342 , P2_U4343 , P2_U4344 , P2_U4345 , P2_U4346 , P2_U4347;
wire P2_U4348 , P2_U4349 , P2_U4350 , P2_U4351 , P2_U4352 , P2_U4353 , P2_U4354 , P2_U4355 , P2_U4356 , P2_U4357;
wire P2_U4358 , P2_U4359 , P2_U4360 , P2_U4361 , P2_U4362 , P2_U4363 , P2_U4364 , P2_U4365 , P2_U4366 , P2_U4367;
wire P2_U4368 , P2_U4369 , P2_U4370 , P2_U4371 , P2_U4372 , P2_U4373 , P2_U4374 , P2_U4375 , P2_U4376 , P2_U4377;
wire P2_U4378 , P2_U4379 , P2_U4380 , P2_U4381 , P2_U4382 , P2_U4383 , P2_U4384 , P2_U4385 , P2_U4386 , P2_U4387;
wire P2_U4388 , P2_U4389 , P2_U4390 , P2_U4391 , P2_U4392 , P2_U4393 , P2_U4394 , P2_U4395 , P2_U4396 , P2_U4397;
wire P2_U4398 , P2_U4399 , P2_U4400 , P2_U4401 , P2_U4402 , P2_U4403 , P2_U4404 , P2_U4405 , P2_U4406 , P2_U4407;
wire P2_U4408 , P2_U4409 , P2_U4410 , P2_U4411 , P2_U4412 , P2_U4413 , P2_U4414 , P2_U4415 , P2_U4416 , P2_U4417;
wire P2_U4418 , P2_U4419 , P2_U4420 , P2_U4421 , P2_U4422 , P2_U4423 , P2_U4424 , P2_U4425 , P2_U4426 , P2_U4427;
wire P2_U4428 , P2_U4429 , P2_U4430 , P2_U4431 , P2_U4432 , P2_U4433 , P2_U4434 , P2_U4435 , P2_U4436 , P2_U4437;
wire P2_U4438 , P2_U4439 , P2_U4440 , P2_U4441 , P2_U4442 , P2_U4443 , P2_U4444 , P2_U4445 , P2_U4446 , P2_U4447;
wire P2_U4448 , P2_U4449 , P2_U4450 , P2_U4451 , P2_U4452 , P2_U4453 , P2_U4454 , P2_U4455 , P2_U4456 , P2_U4457;
wire P2_U4458 , P2_U4459 , P2_U4460 , P2_U4461 , P2_U4462 , P2_U4463 , P2_U4464 , P2_U4465 , P2_U4466 , P2_U4467;
wire P2_U4468 , P2_U4469 , P2_U4470 , P2_U4471 , P2_U4472 , P2_U4473 , P2_U4474 , P2_U4475 , P2_U4476 , P2_U4477;
wire P2_U4478 , P2_U4479 , P2_U4480 , P2_U4481 , P2_U4482 , P2_U4483 , P2_U4484 , P2_U4485 , P2_U4486 , P2_U4487;
wire P2_U4488 , P2_U4489 , P2_U4490 , P2_U4491 , P2_U4492 , P2_U4493 , P2_U4494 , P2_U4495 , P2_U4496 , P2_U4497;
wire P2_U4498 , P2_U4499 , P2_U4500 , P2_U4501 , P2_U4502 , P2_U4503 , P2_U4504 , P2_U4505 , P2_U4506 , P2_U4507;
wire P2_U4508 , P2_U4509 , P2_U4510 , P2_U4511 , P2_U4512 , P2_U4513 , P2_U4514 , P2_U4515 , P2_U4516 , P2_U4517;
wire P2_U4518 , P2_U4519 , P2_U4520 , P2_U4521 , P2_U4522 , P2_U4523 , P2_U4524 , P2_U4525 , P2_U4526 , P2_U4527;
wire P2_U4528 , P2_U4529 , P2_U4530 , P2_U4531 , P2_U4532 , P2_U4533 , P2_U4534 , P2_U4535 , P2_U4536 , P2_U4537;
wire P2_U4538 , P2_U4539 , P2_U4540 , P2_U4541 , P2_U4542 , P2_U4543 , P2_U4544 , P2_U4545 , P2_U4546 , P2_U4547;
wire P2_U4548 , P2_U4549 , P2_U4550 , P2_U4551 , P2_U4552 , P2_U4553 , P2_U4554 , P2_U4555 , P2_U4556 , P2_U4557;
wire P2_U4558 , P2_U4559 , P2_U4560 , P2_U4561 , P2_U4562 , P2_U4563 , P2_U4564 , P2_U4565 , P2_U4566 , P2_U4567;
wire P2_U4568 , P2_U4569 , P2_U4570 , P2_U4571 , P2_U4572 , P2_U4573 , P2_U4574 , P2_U4575 , P2_U4576 , P2_U4577;
wire P2_U4578 , P2_U4579 , P2_U4580 , P2_U4581 , P2_U4582 , P2_U4583 , P2_U4584 , P2_U4585 , P2_U4586 , P2_U4587;
wire P2_U4588 , P2_U4589 , P2_U4590 , P2_U4591 , P2_U4592 , P2_U4593 , P2_U4594 , P2_U4595 , P2_U4596 , P2_U4597;
wire P2_U4598 , P2_U4599 , P2_U4600 , P2_U4601 , P2_U4602 , P2_U4603 , P2_U4604 , P2_U4605 , P2_U4606 , P2_U4607;
wire P2_U4608 , P2_U4609 , P2_U4610 , P2_U4611 , P2_U4612 , P2_U4613 , P2_U4614 , P2_U4615 , P2_U4616 , P2_U4617;
wire P2_U4618 , P2_U4619 , P2_U4620 , P2_U4621 , P2_U4622 , P2_U4623 , P2_U4624 , P2_U4625 , P2_U4626 , P2_U4627;
wire P2_U4628 , P2_U4629 , P2_U4630 , P2_U4631 , P2_U4632 , P2_U4633 , P2_U4634 , P2_U4635 , P2_U4636 , P2_U4637;
wire P2_U4638 , P2_U4639 , P2_U4640 , P2_U4641 , P2_U4642 , P2_U4643 , P2_U4644 , P2_U4645 , P2_U4646 , P2_U4647;
wire P2_U4648 , P2_U4649 , P2_U4650 , P2_U4651 , P2_U4652 , P2_U4653 , P2_U4654 , P2_U4655 , P2_U4656 , P2_U4657;
wire P2_U4658 , P2_U4659 , P2_U4660 , P2_U4661 , P2_U4662 , P2_U4663 , P2_U4664 , P2_U4665 , P2_U4666 , P2_U4667;
wire P2_U4668 , P2_U4669 , P2_U4670 , P2_U4671 , P2_U4672 , P2_U4673 , P2_U4674 , P2_U4675 , P2_U4676 , P2_U4677;
wire P2_U4678 , P2_U4679 , P2_U4680 , P2_U4681 , P2_U4682 , P2_U4683 , P2_U4684 , P2_U4685 , P2_U4686 , P2_U4687;
wire P2_U4688 , P2_U4689 , P2_U4690 , P2_U4691 , P2_U4692 , P2_U4693 , P2_U4694 , P2_U4695 , P2_U4696 , P2_U4697;
wire P2_U4698 , P2_U4699 , P2_U4700 , P2_U4701 , P2_U4702 , P2_U4703 , P2_U4704 , P2_U4705 , P2_U4706 , P2_U4707;
wire P2_U4708 , P2_U4709 , P2_U4710 , P2_U4711 , P2_U4712 , P2_U4713 , P2_U4714 , P2_U4715 , P2_U4716 , P2_U4717;
wire P2_U4718 , P2_U4719 , P2_U4720 , P2_U4721 , P2_U4722 , P2_U4723 , P2_U4724 , P2_U4725 , P2_U4726 , P2_U4727;
wire P2_U4728 , P2_U4729 , P2_U4730 , P2_U4731 , P2_U4732 , P2_U4733 , P2_U4734 , P2_U4735 , P2_U4736 , P2_U4737;
wire P2_U4738 , P2_U4739 , P2_U4740 , P2_U4741 , P2_U4742 , P2_U4743 , P2_U4744 , P2_U4745 , P2_U4746 , P2_U4747;
wire P2_U4748 , P2_U4749 , P2_U4750 , P2_U4751 , P2_U4752 , P2_U4753 , P2_U4754 , P2_U4755 , P2_U4756 , P2_U4757;
wire P2_U4758 , P2_U4759 , P2_U4760 , P2_U4761 , P2_U4762 , P2_U4763 , P2_U4764 , P2_U4765 , P2_U4766 , P2_U4767;
wire P2_U4768 , P2_U4769 , P2_U4770 , P2_U4771 , P2_U4772 , P2_U4773 , P2_U4774 , P2_U4775 , P2_U4776 , P2_U4777;
wire P2_U4778 , P2_U4779 , P2_U4780 , P2_U4781 , P2_U4782 , P2_U4783 , P2_U4784 , P2_U4785 , P2_U4786 , P2_U4787;
wire P2_U4788 , P2_U4789 , P2_U4790 , P2_U4791 , P2_U4792 , P2_U4793 , P2_U4794 , P2_U4795 , P2_U4796 , P2_U4797;
wire P2_U4798 , P2_U4799 , P2_U4800 , P2_U4801 , P2_U4802 , P2_U4803 , P2_U4804 , P2_U4805 , P2_U4806 , P2_U4807;
wire P2_U4808 , P2_U4809 , P2_U4810 , P2_U4811 , P2_U4812 , P2_U4813 , P2_U4814 , P2_U4815 , P2_U4816 , P2_U4817;
wire P2_U4818 , P2_U4819 , P2_U4820 , P2_U4821 , P2_U4822 , P2_U4823 , P2_U4824 , P2_U4825 , P2_U4826 , P2_U4827;
wire P2_U4828 , P2_U4829 , P2_U4830 , P2_U4831 , P2_U4832 , P2_U4833 , P2_U4834 , P2_U4835 , P2_U4836 , P2_U4837;
wire P2_U4838 , P2_U4839 , P2_U4840 , P2_U4841 , P2_U4842 , P2_U4843 , P2_U4844 , P2_U4845 , P2_U4846 , P2_U4847;
wire P2_U4848 , P2_U4849 , P2_U4850 , P2_U4851 , P2_U4852 , P2_U4853 , P2_U4854 , P2_U4855 , P2_U4856 , P2_U4857;
wire P2_U4858 , P2_U4859 , P2_U4860 , P2_U4861 , P2_U4862 , P2_U4863 , P2_U4864 , P2_U4865 , P2_U4866 , P2_U4867;
wire P2_U4868 , P2_U4869 , P2_U4870 , P2_U4871 , P2_U4872 , P2_U4873 , P2_U4874 , P2_U4875 , P2_U4876 , P2_U4877;
wire P2_U4878 , P2_U4879 , P2_U4880 , P2_U4881 , P2_U4882 , P2_U4883 , P2_U4884 , P2_U4885 , P2_U4886 , P2_U4887;
wire P2_U4888 , P2_U4889 , P2_U4890 , P2_U4891 , P2_U4892 , P2_U4893 , P2_U4894 , P2_U4895 , P2_U4896 , P2_U4897;
wire P2_U4898 , P2_U4899 , P2_U4900 , P2_U4901 , P2_U4902 , P2_U4903 , P2_U4904 , P2_U4905 , P2_U4906 , P2_U4907;
wire P2_U4908 , P2_U4909 , P2_U4910 , P2_U4911 , P2_U4912 , P2_U4913 , P2_U4914 , P2_U4915 , P2_U4916 , P2_U4917;
wire P2_U4918 , P2_U4919 , P2_U4920 , P2_U4921 , P2_U4922 , P2_U4923 , P2_U4924 , P2_U4925 , P2_U4926 , P2_U4927;
wire P2_U4928 , P2_U4929 , P2_U4930 , P2_U4931 , P2_U4932 , P2_U4933 , P2_U4934 , P2_U4935 , P2_U4936 , P2_U4937;
wire P2_U4938 , P2_U4939 , P2_U4940 , P2_U4941 , P2_U4942 , P2_U4943 , P2_U4944 , P2_U4945 , P2_U4946 , P2_U4947;
wire P2_U4948 , P2_U4949 , P2_U4950 , P2_U4951 , P2_U4952 , P2_U4953 , P2_U4954 , P2_U4955 , P2_U4956 , P2_U4957;
wire P2_U4958 , P2_U4959 , P2_U4960 , P2_U4961 , P2_U4962 , P2_U4963 , P2_U4964 , P2_U4965 , P2_U4966 , P2_U4967;
wire P2_U4968 , P2_U4969 , P2_U4970 , P2_U4971 , P2_U4972 , P2_U4973 , P2_U4974 , P2_U4975 , P2_U4976 , P2_U4977;
wire P2_U4978 , P2_U4979 , P2_U4980 , P2_U4981 , P2_U4982 , P2_U4983 , P2_U4984 , P2_U4985 , P2_U4986 , P2_U4987;
wire P2_U4988 , P2_U4989 , P2_U4990 , P2_U4991 , P2_U4992 , P2_U4993 , P2_U4994 , P2_U4995 , P2_U4996 , P2_U4997;
wire P2_U4998 , P2_U4999 , P2_U5000 , P2_U5001 , P2_U5002 , P2_U5003 , P2_U5004 , P2_U5005 , P2_U5006 , P2_U5007;
wire P2_U5008 , P2_U5009 , P2_U5010 , P2_U5011 , P2_U5012 , P2_U5013 , P2_U5014 , P2_U5015 , P2_U5016 , P2_U5017;
wire P2_U5018 , P2_U5019 , P2_U5020 , P2_U5021 , P2_U5022 , P2_U5023 , P2_U5024 , P2_U5025 , P2_U5026 , P2_U5027;
wire P2_U5028 , P2_U5029 , P2_U5030 , P2_U5031 , P2_U5032 , P2_U5033 , P2_U5034 , P2_U5035 , P2_U5036 , P2_U5037;
wire P2_U5038 , P2_U5039 , P2_U5040 , P2_U5041 , P2_U5042 , P2_U5043 , P2_U5044 , P2_U5045 , P2_U5046 , P2_U5047;
wire P2_U5048 , P2_U5049 , P2_U5050 , P2_U5051 , P2_U5052 , P2_U5053 , P2_U5054 , P2_U5055 , P2_U5056 , P2_U5057;
wire P2_U5058 , P2_U5059 , P2_U5060 , P2_U5061 , P2_U5062 , P2_U5063 , P2_U5064 , P2_U5065 , P2_U5066 , P2_U5067;
wire P2_U5068 , P2_U5069 , P2_U5070 , P2_U5071 , P2_U5072 , P2_U5073 , P2_U5074 , P2_U5075 , P2_U5076 , P2_U5077;
wire P2_U5078 , P2_U5079 , P2_U5080 , P2_U5081 , P2_U5082 , P2_U5083 , P2_U5084 , P2_U5085 , P2_U5086 , P2_U5087;
wire P2_U5088 , P2_U5089 , P2_U5090 , P2_U5091 , P2_U5092 , P2_U5093 , P2_U5094 , P2_U5095 , P2_U5096 , P2_U5097;
wire P2_U5098 , P2_U5099 , P2_U5100 , P2_U5101 , P2_U5102 , P2_U5103 , P2_U5104 , P2_U5105 , P2_U5106 , P2_U5107;
wire P2_U5108 , P2_U5109 , P2_U5110 , P2_U5111 , P2_U5112 , P2_U5113 , P2_U5114 , P2_U5115 , P2_U5116 , P2_U5117;
wire P2_U5118 , P2_U5119 , P2_U5120 , P2_U5121 , P2_U5122 , P2_U5123 , P2_U5124 , P2_U5125 , P2_U5126 , P2_U5127;
wire P2_U5128 , P2_U5129 , P2_U5130 , P2_U5131 , P2_U5132 , P2_U5133 , P2_U5134 , P2_U5135 , P2_U5136 , P2_U5137;
wire P2_U5138 , P2_U5139 , P2_U5140 , P2_U5141 , P2_U5142 , P2_U5143 , P2_U5144 , P2_U5145 , P2_U5146 , P2_U5147;
wire P2_U5148 , P2_U5149 , P2_U5150 , P2_U5151 , P2_U5152 , P2_U5153 , P2_U5154 , P2_U5155 , P2_U5156 , P2_U5157;
wire P2_U5158 , P2_U5159 , P2_U5160 , P2_U5161 , P2_U5162 , P2_U5163 , P2_U5164 , P2_U5165 , P2_U5166 , P2_U5167;
wire P2_U5168 , P2_U5169 , P2_U5170 , P2_U5171 , P2_U5172 , P2_U5173 , P2_U5174 , P2_U5175 , P2_U5176 , P2_U5177;
wire P2_U5178 , P2_U5179 , P2_U5180 , P2_U5181 , P2_U5182 , P2_U5183 , P2_U5184 , P2_U5185 , P2_U5186 , P2_U5187;
wire P2_U5188 , P2_U5189 , P2_U5190 , P2_U5191 , P2_U5192 , P2_U5193 , P2_U5194 , P2_U5195 , P2_U5196 , P2_U5197;
wire P2_U5198 , P2_U5199 , P2_U5200 , P2_U5201 , P2_U5202 , P2_U5203 , P2_U5204 , P2_U5205 , P2_U5206 , P2_U5207;
wire P2_U5208 , P2_U5209 , P2_U5210 , P2_U5211 , P2_U5212 , P2_U5213 , P2_U5214 , P2_U5215 , P2_U5216 , P2_U5217;
wire P2_U5218 , P2_U5219 , P2_U5220 , P2_U5221 , P2_U5222 , P2_U5223 , P2_U5224 , P2_U5225 , P2_U5226 , P2_U5227;
wire P2_U5228 , P2_U5229 , P2_U5230 , P2_U5231 , P2_U5232 , P2_U5233 , P2_U5234 , P2_U5235 , P2_U5236 , P2_U5237;
wire P2_U5238 , P2_U5239 , P2_U5240 , P2_U5241 , P2_U5242 , P2_U5243 , P2_U5244 , P2_U5245 , P2_U5246 , P2_U5247;
wire P2_U5248 , P2_U5249 , P2_U5250 , P2_U5251 , P2_U5252 , P2_U5253 , P2_U5254 , P2_U5255 , P2_U5256 , P2_U5257;
wire P2_U5258 , P2_U5259 , P2_U5260 , P2_U5261 , P2_U5262 , P2_U5263 , P2_U5264 , P2_U5265 , P2_U5266 , P2_U5267;
wire P2_U5268 , P2_U5269 , P2_U5270 , P2_U5271 , P2_U5272 , P2_U5273 , P2_U5274 , P2_U5275 , P2_U5276 , P2_U5277;
wire P2_U5278 , P2_U5279 , P2_U5280 , P2_U5281 , P2_U5282 , P2_U5283 , P2_U5284 , P2_U5285 , P2_U5286 , P2_U5287;
wire P2_U5288 , P2_U5289 , P2_U5290 , P2_U5291 , P2_U5292 , P2_U5293 , P2_U5294 , P2_U5295 , P2_U5296 , P2_U5297;
wire P2_U5298 , P2_U5299 , P2_U5300 , P2_U5301 , P2_U5302 , P2_U5303 , P2_U5304 , P2_U5305 , P2_U5306 , P2_U5307;
wire P2_U5308 , P2_U5309 , P2_U5310 , P2_U5311 , P2_U5312 , P2_U5313 , P2_U5314 , P2_U5315 , P2_U5316 , P2_U5317;
wire P2_U5318 , P2_U5319 , P2_U5320 , P2_U5321 , P2_U5322 , P2_U5323 , P2_U5324 , P2_U5325 , P2_U5326 , P2_U5327;
wire P2_U5328 , P2_U5329 , P2_U5330 , P2_U5331 , P2_U5332 , P2_U5333 , P2_U5334 , P2_U5335 , P2_U5336 , P2_U5337;
wire P2_U5338 , P2_U5339 , P2_U5340 , P2_U5341 , P2_U5342 , P2_U5343 , P2_U5344 , P2_U5345 , P2_U5346 , P2_U5347;
wire P2_U5348 , P2_U5349 , P2_U5350 , P2_U5351 , P2_U5352 , P2_U5353 , P2_U5354 , P2_U5355 , P2_U5356 , P2_U5357;
wire P2_U5358 , P2_U5359 , P2_U5360 , P2_U5361 , P2_U5362 , P2_U5363 , P2_U5364 , P2_U5365 , P2_U5366 , P2_U5367;
wire P2_U5368 , P2_U5369 , P2_U5370 , P2_U5371 , P2_U5372 , P2_U5373 , P2_U5374 , P2_U5375 , P2_U5376 , P2_U5377;
wire P2_U5378 , P2_U5379 , P2_U5380 , P2_U5381 , P2_U5382 , P2_U5383 , P2_U5384 , P2_U5385 , P2_U5386 , P2_U5387;
wire P2_U5388 , P2_U5389 , P2_U5390 , P2_U5391 , P2_U5392 , P2_U5393 , P2_U5394 , P2_U5395 , P2_U5396 , P2_U5397;
wire P2_U5398 , P2_U5399 , P2_U5400 , P2_U5401 , P2_U5402 , P2_U5403 , P2_U5404 , P2_U5405 , P2_U5406 , P2_U5407;
wire P2_U5408 , P2_U5409 , P2_U5410 , P2_U5411 , P2_U5412 , P2_U5413 , P2_U5414 , P2_U5415 , P2_U5416 , P2_U5417;
wire P2_U5418 , P2_U5419 , P2_U5420 , P2_U5421 , P2_U5422 , P2_U5423 , P2_U5424 , P2_U5425 , P2_U5426 , P2_U5427;
wire P2_U5428 , P2_U5429 , P2_U5430 , P2_U5431 , P2_U5432 , P2_U5433 , P2_U5434 , P2_U5435 , P2_U5436 , P2_U5437;
wire P2_U5438 , P2_U5439 , P2_U5440 , P2_U5441 , P2_U5442 , P2_U5443 , P2_U5444 , P2_U5445 , P2_U5446 , P2_U5447;
wire P2_U5448 , P2_U5449 , P2_U5450 , P2_U5451 , P2_U5452 , P2_U5453 , P2_U5454 , P2_U5455 , P2_U5456 , P2_U5457;
wire P2_U5458 , P2_U5459 , P2_U5460 , P2_U5461 , P2_U5462 , P2_U5463 , P2_U5464 , P2_U5465 , P2_U5466 , P2_U5467;
wire P2_U5468 , P2_U5469 , P2_U5470 , P2_U5471 , P2_U5472 , P2_U5473 , P2_U5474 , P2_U5475 , P2_U5476 , P2_U5477;
wire P2_U5478 , P2_U5479 , P2_U5480 , P2_U5481 , P2_U5482 , P2_U5483 , P2_U5484 , P2_U5485 , P2_U5486 , P2_U5487;
wire P2_U5488 , P2_U5489 , P2_U5490 , P2_U5491 , P2_U5492 , P2_U5493 , P2_U5494 , P2_U5495 , P2_U5496 , P2_U5497;
wire P2_U5498 , P2_U5499 , P2_U5500 , P2_U5501 , P2_U5502 , P2_U5503 , P2_U5504 , P2_U5505 , P2_U5506 , P2_U5507;
wire P2_U5508 , P2_U5509 , P2_U5510 , P2_U5511 , P2_U5512 , P2_U5513 , P2_U5514 , P2_U5515 , P2_U5516 , P2_U5517;
wire P2_U5518 , P2_U5519 , P2_U5520 , P2_U5521 , P2_U5522 , P2_U5523 , P2_U5524 , P2_U5525 , P2_U5526 , P2_U5527;
wire P2_U5528 , P2_U5529 , P2_U5530 , P2_U5531 , P2_U5532 , P2_U5533 , P2_U5534 , P2_U5535 , P2_U5536 , P2_U5537;
wire P2_U5538 , P2_U5539 , P2_U5540 , P2_U5541 , P2_U5542 , P2_U5543 , P2_U5544 , P2_U5545 , P2_U5546 , P2_U5547;
wire P2_U5548 , P2_U5549 , P2_U5550 , P2_U5551 , P2_U5552 , P2_U5553 , P2_U5554 , P2_U5555 , P2_U5556 , P2_U5557;
wire P2_U5558 , P2_U5559 , P2_U5560 , P2_U5561 , P2_U5562 , P2_U5563 , P2_U5564 , P2_U5565 , P2_U5566 , P2_U5567;
wire P2_U5568 , P2_U5569 , P2_U5570 , P2_U5571 , P2_U5572 , P2_U5573 , P2_U5574 , P2_U5575 , P2_U5576 , P2_U5577;
wire P2_U5578 , P2_U5579 , P2_U5580 , P2_U5581 , P2_U5582 , P2_U5583 , P2_U5584 , P2_U5585 , P2_U5586 , P2_U5587;
wire P2_U5588 , P2_U5589 , P2_U5590 , P2_U5591 , P2_U5592 , P2_U5593 , P2_U5594 , P2_U5595 , P2_U5596 , P2_U5597;
wire P2_U5598 , P2_U5599 , P2_U5600 , P2_U5601 , P2_U5602 , P2_U5603 , P2_U5604 , P2_U5605 , P2_U5606 , P2_U5607;
wire P2_U5608 , P2_U5609 , P2_U5610 , P2_U5611 , P2_U5612 , P2_U5613 , P2_U5614 , P2_U5615 , P2_U5616 , P2_U5617;
wire P2_U5618 , P2_U5619 , P2_U5620 , P2_U5621 , P2_U5622 , P2_U5623 , P2_U5624 , P2_U5625 , P2_U5626 , P2_U5627;
wire P2_U5628 , P2_U5629 , P2_U5630 , P2_U5631 , P2_U5632 , P2_U5633 , P2_U5634 , P2_U5635 , P2_U5636 , P2_U5637;
wire P2_U5638 , P2_U5639 , P2_U5640 , P2_U5641 , P2_U5642 , P2_U5643 , P2_U5644 , P2_U5645 , P2_U5646 , P2_U5647;
wire P2_U5648 , P2_U5649 , P2_U5650 , P2_U5651 , P2_U5652 , P2_U5653 , P2_U5654 , P2_U5655 , P2_U5656 , P2_U5657;
wire P2_U5658 , P2_U5659 , P2_U5660 , P2_U5661 , P2_U5662 , P2_U5663 , P2_U5664 , P2_U5665 , P2_U5666 , P2_U5667;
wire P2_U5668 , P2_U5669 , P2_U5670 , P2_U5671 , P2_U5672 , P2_U5673 , P2_U5674 , P2_U5675 , P2_U5676 , P2_U5677;
wire P2_U5678 , P2_U5679 , P2_U5680 , P2_U5681 , P2_U5682 , P2_U5683 , P2_U5684 , P2_U5685 , P2_U5686 , P2_U5687;
wire P2_U5688 , P2_U5689 , P2_U5690 , P2_U5691 , P2_U5692 , P2_U5693 , P2_U5694 , P2_U5695 , P2_U5696 , P2_U5697;
wire P2_U5698 , P2_U5699 , P2_U5700 , P2_U5701 , P2_U5702 , P2_U5703 , P2_U5704 , P2_U5705 , P2_U5706 , P2_U5707;
wire P2_U5708 , P2_U5709 , P2_U5710 , P2_U5711 , P2_U5712 , P2_U5713 , P2_U5714 , P2_U5715 , P2_U5716 , P2_U5717;
wire P2_U5718 , P2_U5719 , P2_U5720 , P2_U5721 , P2_U5722 , P2_U5723 , P2_U5724 , P2_U5725 , P2_U5726 , P2_U5727;
wire P2_U5728 , P2_U5729 , P2_U5730 , P2_U5731 , P2_U5732 , P2_U5733 , P2_U5734 , P2_U5735 , P2_U5736 , P2_U5737;
wire P2_U5738 , P2_U5739 , P2_U5740 , P2_U5741 , P2_U5742 , P2_U5743 , P2_U5744 , P2_U5745 , P2_U5746 , P2_U5747;
wire P2_U5748 , P2_U5749 , P2_U5750 , P2_U5751 , P2_U5752 , P2_U5753 , P2_U5754 , P2_U5755 , P2_U5756 , P2_U5757;
wire P2_U5758 , P2_U5759 , P2_U5760 , P2_U5761 , P2_U5762 , P2_U5763 , P2_U5764 , P2_U5765 , P2_U5766 , P2_U5767;
wire P2_U5768 , P2_U5769 , P2_U5770 , P2_U5771 , P2_U5772 , P2_U5773 , P2_U5774 , P2_U5775 , P2_U5776 , P2_U5777;
wire P2_U5778 , P2_U5779 , P2_U5780 , P2_U5781 , P2_U5782 , P2_U5783 , P2_U5784 , P2_U5785 , P2_U5786 , P2_U5787;
wire P2_U5788 , P2_U5789 , P2_U5790 , P2_U5791 , P2_U5792 , P2_U5793 , P2_U5794 , P2_U5795 , P2_U5796 , P2_U5797;
wire P2_U5798 , P2_U5799 , P2_U5800 , P2_U5801 , P2_U5802 , P2_U5803 , P2_U5804 , P2_U5805 , P2_U5806 , P2_U5807;
wire P2_U5808 , P2_U5809 , P2_U5810 , P2_U5811 , P2_U5812 , P2_U5813 , P2_U5814 , P2_U5815 , P2_U5816 , P2_U5817;
wire P2_U5818 , P2_U5819 , P2_U5820 , P2_U5821 , P2_U5822 , P2_U5823 , P2_U5824 , P2_U5825 , P2_U5826 , P2_U5827;
wire P2_U5828 , P2_U5829 , P2_U5830 , P2_U5831 , P2_U5832 , P2_U5833 , P2_U5834 , P2_U5835 , P2_U5836 , P2_U5837;
wire P2_U5838 , P2_U5839 , P2_U5840 , P2_U5841 , P2_U5842 , P2_U5843 , P2_U5844 , P2_U5845 , P2_U5846 , P2_U5847;
wire P2_U5848 , P2_U5849 , P2_U5850 , P2_U5851 , P2_U5852 , P2_U5853 , P2_U5854 , P2_U5855 , P2_U5856 , P2_U5857;
wire P2_U5858 , P2_U5859 , P2_U5860 , P2_U5861 , P2_U5862 , P2_U5863 , P2_U5864 , P2_U5865 , P2_U5866 , P2_U5867;
wire P2_U5868 , P2_U5869 , P2_U5870 , P2_U5871 , P2_U5872 , P2_U5873 , P2_U5874 , P2_U5875 , P2_U5876 , P2_U5877;
wire P2_U5878 , P2_U5879 , P2_U5880 , P2_U5881 , P2_U5882 , P2_U5883 , P2_U5884 , P2_U5885 , P2_U5886 , P2_U5887;
wire P2_U5888 , P2_U5889 , P2_U5890 , P2_U5891 , P2_U5892 , P2_U5893 , P2_U5894 , P2_U5895 , P2_U5896 , P2_U5897;
wire P2_U5898 , P2_U5899 , P2_U5900 , P2_U5901 , P2_U5902 , P2_U5903 , P2_U5904 , P2_U5905 , P2_U5906 , P2_U5907;
wire P2_U5908 , P2_U5909 , P2_U5910 , P2_U5911 , P2_U5912 , P2_U5913 , P2_U5914 , P2_U5915 , P2_U5916 , P2_U5917;
wire P2_U5918 , P2_U5919 , P2_U5920 , P2_U5921 , P2_U5922 , P2_U5923 , P2_U5924 , P2_U5925 , P2_U5926 , P2_U5927;
wire P2_U5928 , P2_U5929 , P2_U5930 , P2_U5931 , P2_U5932 , P2_U5933 , P2_U5934 , P2_U5935 , P2_U5936 , P2_U5937;
wire P2_U5938 , P2_U5939 , P2_U5940 , P2_U5941 , P2_U5942 , P2_U5943 , P2_U5944 , P2_U5945 , P2_U5946 , P2_U5947;
wire P2_U5948 , P2_U5949 , P2_U5950 , P2_U5951 , P2_U5952 , P2_U5953 , P2_U5954 , P2_U5955 , P2_U5956 , P2_U5957;
wire P2_U5958 , P2_U5959 , P2_U5960 , P2_U5961 , P2_U5962 , P2_U5963 , P2_U5964 , P2_U5965 , P2_U5966 , P2_U5967;
wire P2_U5968 , P2_U5969 , P2_U5970 , P2_U5971 , P2_U5972 , P2_U5973 , P2_U5974 , P2_U5975 , P2_U5976 , P2_U5977;
wire P2_U5978 , P2_U5979 , P2_U5980 , P2_U5981 , P2_U5982 , P2_U5983 , P2_U5984 , P2_U5985 , P2_U5986 , P2_U5987;
wire P2_U5988 , P2_U5989 , P2_U5990 , P2_U5991 , P2_U5992 , P2_U5993 , P2_U5994 , P2_U5995 , P2_U5996 , P2_U5997;
wire P2_U5998 , P2_U5999 , P2_U6000 , P2_U6001 , P2_U6002 , P2_U6003 , P2_U6004 , P2_U6005 , P2_U6006 , P2_U6007;
wire P2_U6008 , P2_U6009 , P2_U6010 , P2_U6011 , P2_U6012 , P2_U6013 , P2_U6014 , P2_U6015 , P2_U6016 , P2_U6017;
wire P2_U6018 , P2_U6019 , P2_U6020 , P2_U6021 , P2_U6022 , P2_U6023 , P2_U6024 , P2_U6025 , P2_U6026 , P2_U6027;
wire P2_U6028 , P2_U6029 , P2_U6030 , P2_U6031 , P2_U6032 , P2_U6033 , P2_U6034 , P2_U6035 , P2_U6036 , P2_U6037;
wire P2_U6038 , P2_U6039 , P2_U6040 , P2_U6041 , P2_U6042 , P2_U6043 , P2_U6044 , P2_U6045 , P2_U6046 , P2_U6047;
wire P2_U6048 , P2_U6049 , P2_U6050 , P2_U6051 , P2_U6052 , P2_U6053 , P2_U6054 , P2_U6055 , P2_U6056 , P2_U6057;
wire P2_U6058 , P2_U6059 , P2_U6060 , P2_U6061 , P2_U6062 , P2_U6063 , P2_U6064 , P2_U6065 , P2_U6066 , P2_U6067;
wire P2_U6068 , P2_U6069 , P2_U6070 , P2_U6071 , P2_U6072 , P2_U6073 , P2_U6074 , P2_U6075 , P2_U6076 , P2_U6077;
wire P2_U6078 , P2_U6079 , P2_U6080 , P2_U6081 , P2_U6082 , P2_U6083 , P2_U6084 , P2_U6085 , P2_U6086 , P2_U6087;
wire P2_U6088 , P2_U6089 , P2_U6090 , P2_U6091 , P2_U6092 , P2_U6093 , P2_U6094 , P2_U6095 , P2_U6096 , P2_U6097;
wire P2_U6098 , P2_U6099 , P2_U6100 , P2_U6101 , P2_U6102 , P2_U6103 , P2_U6104 , P2_U6105 , P2_U6106 , P2_U6107;
wire P2_U6108 , P2_U6109 , P2_U6110 , P2_U6111 , P2_U6112 , P2_U6113 , P2_U6114 , P2_U6115 , P2_U6116 , P2_U6117;
wire P2_U6118 , P2_U6119 , P2_U6120 , P2_U6121 , P2_U6122 , P2_U6123 , P2_U6124 , P2_U6125 , P2_U6126 , P2_U6127;
wire P2_U6128 , P2_U6129 , P2_U6130 , P2_U6131 , P2_U6132 , P2_U6133 , P2_U6134 , P2_U6135 , P2_U6136 , P2_U6137;
wire P2_U6138 , P2_U6139 , P2_U6140 , P2_U6141 , P2_U6142 , P2_U6143 , P2_U6144 , P2_U6145 , P2_U6146 , P2_U6147;
wire P2_U6148 , P2_U6149 , P2_U6150 , P3_R1161_U468 , P3_R1161_U467 , P3_R1161_U466 , P3_R1161_U465 , P3_R1161_U464 , P3_R1161_U463 , P3_R1161_U462;
wire P3_R1161_U461 , P3_R1161_U460 , P3_R1161_U459 , P3_R1161_U458 , P3_R1161_U457 , P3_R1161_U456 , P3_R1161_U455 , P3_R1161_U454 , P3_R1161_U453 , P3_R1161_U452;
wire P3_R1161_U451 , P3_R1161_U450 , P3_R1161_U449 , P3_U3013 , P3_U3014 , P3_U3015 , P3_U3016 , P3_U3017 , P3_U3018 , P3_U3019;
wire P3_U3020 , P3_U3021 , P3_U3022 , P3_U3023 , P3_U3024 , P3_U3025 , P3_U3026 , P3_U3027 , P3_U3028 , P3_U3029;
wire P3_U3030 , P3_U3031 , P3_U3032 , P3_U3033 , P3_U3034 , P3_U3035 , P3_U3036 , P3_U3037 , P3_U3038 , P3_U3039;
wire P3_U3040 , P3_U3041 , P3_U3042 , P3_U3043 , P3_U3044 , P3_U3045 , P3_U3046 , P3_U3047 , P3_U3048 , P3_U3049;
wire P3_U3050 , P3_U3051 , P3_U3052 , P3_U3053 , P3_U3054 , P3_U3055 , P3_U3056 , P3_U3057 , P3_U3058 , P3_U3059;
wire P3_U3060 , P3_U3061 , P3_U3062 , P3_U3063 , P3_U3064 , P3_U3065 , P3_U3066 , P3_U3067 , P3_U3068 , P3_U3069;
wire P3_U3070 , P3_U3071 , P3_U3072 , P3_U3073 , P3_U3074 , P3_U3075 , P3_U3076 , P3_U3077 , P3_U3078 , P3_U3079;
wire P3_U3080 , P3_U3081 , P3_U3082 , P3_U3083 , P3_U3084 , P3_U3085 , P3_U3086 , P3_U3087 , P3_U3088 , P3_U3089;
wire P3_U3090 , P3_U3091 , P3_U3092 , P3_U3093 , P3_U3094 , P3_U3095 , P3_U3096 , P3_U3097 , P3_U3098 , P3_U3099;
wire P3_U3100 , P3_U3101 , P3_U3102 , P3_U3103 , P3_U3104 , P3_U3105 , P3_U3106 , P3_U3107 , P3_U3108 , P3_U3109;
wire P3_U3110 , P3_U3111 , P3_U3112 , P3_U3113 , P3_U3114 , P3_U3115 , P3_U3116 , P3_U3117 , P3_U3118 , P3_U3119;
wire P3_U3120 , P3_U3121 , P3_U3122 , P3_U3123 , P3_U3124 , P3_U3125 , P3_U3126 , P3_U3127 , P3_U3128 , P3_U3129;
wire P3_U3130 , P3_U3131 , P3_U3132 , P3_U3133 , P3_U3134 , P3_U3135 , P3_U3136 , P3_U3137 , P3_U3138 , P3_U3139;
wire P3_U3140 , P3_U3141 , P3_U3142 , P3_U3143 , P3_U3144 , P3_U3145 , P3_U3146 , P3_U3147 , P3_U3148 , P3_U3149;
wire P3_U3152 , P3_U3297 , P3_U3298 , P3_U3299 , P3_U3300 , P3_U3301 , P3_U3302 , P3_U3303 , P3_U3304 , P3_U3305;
wire P3_U3306 , P3_U3307 , P3_U3308 , P3_U3309 , P3_U3310 , P3_U3311 , P3_U3312 , P3_U3313 , P3_U3314 , P3_U3315;
wire P3_U3316 , P3_U3317 , P3_U3318 , P3_U3319 , P3_U3320 , P3_U3321 , P3_U3322 , P3_U3323 , P3_U3324 , P3_U3325;
wire P3_U3326 , P3_U3327 , P3_U3328 , P3_U3329 , P3_U3330 , P3_U3331 , P3_U3332 , P3_U3333 , P3_U3334 , P3_U3335;
wire P3_U3336 , P3_U3337 , P3_U3338 , P3_U3339 , P3_U3340 , P3_U3341 , P3_U3342 , P3_U3343 , P3_U3344 , P3_U3345;
wire P3_U3346 , P3_U3347 , P3_U3348 , P3_U3349 , P3_U3350 , P3_U3351 , P3_U3352 , P3_U3353 , P3_U3354 , P3_U3355;
wire P3_U3356 , P3_U3357 , P3_U3358 , P3_U3359 , P3_U3360 , P3_U3361 , P3_U3362 , P3_U3363 , P3_U3364 , P3_U3365;
wire P3_U3366 , P3_U3367 , P3_U3368 , P3_U3369 , P3_U3370 , P3_U3371 , P3_U3372 , P3_U3373 , P3_U3374 , P3_U3375;
wire P3_U3378 , P3_U3379 , P3_U3380 , P3_U3381 , P3_U3382 , P3_U3383 , P3_U3384 , P3_U3385 , P3_U3386 , P3_U3387;
wire P3_U3388 , P3_U3389 , P3_U3391 , P3_U3392 , P3_U3394 , P3_U3395 , P3_U3397 , P3_U3398 , P3_U3400 , P3_U3401;
wire P3_U3403 , P3_U3404 , P3_U3406 , P3_U3407 , P3_U3409 , P3_U3410 , P3_U3412 , P3_U3413 , P3_U3415 , P3_U3416;
wire P3_U3418 , P3_U3419 , P3_U3421 , P3_U3422 , P3_U3424 , P3_U3425 , P3_U3427 , P3_U3428 , P3_U3430 , P3_U3431;
wire P3_U3433 , P3_U3434 , P3_U3436 , P3_U3437 , P3_U3439 , P3_U3440 , P3_U3442 , P3_U3443 , P3_U3445 , P3_U3523;
wire P3_U3524 , P3_U3525 , P3_U3526 , P3_U3527 , P3_U3528 , P3_U3529 , P3_U3530 , P3_U3531 , P3_U3532 , P3_U3533;
wire P3_U3534 , P3_U3535 , P3_U3536 , P3_U3537 , P3_U3538 , P3_U3539 , P3_U3540 , P3_U3541 , P3_U3542 , P3_U3543;
wire P3_U3544 , P3_U3545 , P3_U3546 , P3_U3547 , P3_U3548 , P3_U3549 , P3_U3550 , P3_U3551 , P3_U3552 , P3_U3553;
wire P3_U3554 , P3_U3555 , P3_U3556 , P3_U3557 , P3_U3558 , P3_U3559 , P3_U3560 , P3_U3561 , P3_U3562 , P3_U3563;
wire P3_U3564 , P3_U3565 , P3_U3566 , P3_U3567 , P3_U3568 , P3_U3569 , P3_U3570 , P3_U3571 , P3_U3572 , P3_U3573;
wire P3_U3574 , P3_U3575 , P3_U3576 , P3_U3577 , P3_U3578 , P3_U3579 , P3_U3580 , P3_U3581 , P3_U3582 , P3_U3583;
wire P3_U3584 , P3_U3585 , P3_U3586 , P3_U3587 , P3_U3588 , P3_U3589 , P3_U3590 , P3_U3591 , P3_U3592 , P3_U3593;
wire P3_U3594 , P3_U3595 , P3_U3596 , P3_U3597 , P3_U3598 , P3_U3599 , P3_U3600 , P3_U3601 , P3_U3602 , P3_U3603;
wire P3_U3604 , P3_U3605 , P3_U3606 , P3_U3607 , P3_U3608 , P3_U3609 , P3_U3610 , P3_U3611 , P3_U3612 , P3_U3613;
wire P3_U3614 , P3_U3615 , P3_U3616 , P3_U3617 , P3_U3618 , P3_U3619 , P3_U3620 , P3_U3621 , P3_U3622 , P3_U3623;
wire P3_U3624 , P3_U3625 , P3_U3626 , P3_U3627 , P3_U3628 , P3_U3629 , P3_U3630 , P3_U3631 , P3_U3632 , P3_U3633;
wire P3_U3634 , P3_U3635 , P3_U3636 , P3_U3637 , P3_U3638 , P3_U3639 , P3_U3640 , P3_U3641 , P3_U3642 , P3_U3643;
wire P3_U3644 , P3_U3645 , P3_U3646 , P3_U3647 , P3_U3648 , P3_U3649 , P3_U3650 , P3_U3651 , P3_U3652 , P3_U3653;
wire P3_U3654 , P3_U3655 , P3_U3656 , P3_U3657 , P3_U3658 , P3_U3659 , P3_U3660 , P3_U3661 , P3_U3662 , P3_U3663;
wire P3_U3664 , P3_U3665 , P3_U3666 , P3_U3667 , P3_U3668 , P3_U3669 , P3_U3670 , P3_U3671 , P3_U3672 , P3_U3673;
wire P3_U3674 , P3_U3675 , P3_U3676 , P3_U3677 , P3_U3678 , P3_U3679 , P3_U3680 , P3_U3681 , P3_U3682 , P3_U3683;
wire P3_U3684 , P3_U3685 , P3_U3686 , P3_U3687 , P3_U3688 , P3_U3689 , P3_U3690 , P3_U3691 , P3_U3692 , P3_U3693;
wire P3_U3694 , P3_U3695 , P3_U3696 , P3_U3697 , P3_U3698 , P3_U3699 , P3_U3700 , P3_U3701 , P3_U3702 , P3_U3703;
wire P3_U3704 , P3_U3705 , P3_U3706 , P3_U3707 , P3_U3708 , P3_U3709 , P3_U3710 , P3_U3711 , P3_U3712 , P3_U3713;
wire P3_U3714 , P3_U3715 , P3_U3716 , P3_U3717 , P3_U3718 , P3_U3719 , P3_U3720 , P3_U3721 , P3_U3722 , P3_U3723;
wire P3_U3724 , P3_U3725 , P3_U3726 , P3_U3727 , P3_U3728 , P3_U3729 , P3_U3730 , P3_U3731 , P3_U3732 , P3_U3733;
wire P3_U3734 , P3_U3735 , P3_U3736 , P3_U3737 , P3_U3738 , P3_U3739 , P3_U3740 , P3_U3741 , P3_U3742 , P3_U3743;
wire P3_U3744 , P3_U3745 , P3_U3746 , P3_U3747 , P3_U3748 , P3_U3749 , P3_U3750 , P3_U3751 , P3_U3752 , P3_U3753;
wire P3_U3754 , P3_U3755 , P3_U3756 , P3_U3757 , P3_U3758 , P3_U3759 , P3_U3760 , P3_U3761 , P3_U3762 , P3_U3763;
wire P3_U3764 , P3_U3765 , P3_U3766 , P3_U3767 , P3_U3768 , P3_U3769 , P3_U3770 , P3_U3771 , P3_U3772 , P3_U3773;
wire P3_U3774 , P3_U3775 , P3_U3776 , P3_U3777 , P3_U3778 , P3_U3779 , P3_U3780 , P3_U3781 , P3_U3782 , P3_U3783;
wire P3_U3784 , P3_U3785 , P3_U3786 , P3_U3787 , P3_U3788 , P3_U3789 , P3_U3790 , P3_U3791 , P3_U3792 , P3_U3793;
wire P3_U3794 , P3_U3795 , P3_U3796 , P3_U3797 , P3_U3798 , P3_U3799 , P3_U3800 , P3_U3801 , P3_U3802 , P3_U3803;
wire P3_U3804 , P3_U3805 , P3_U3806 , P3_U3807 , P3_U3808 , P3_U3809 , P3_U3810 , P3_U3811 , P3_U3812 , P3_U3813;
wire P3_U3814 , P3_U3815 , P3_U3816 , P3_U3817 , P3_U3818 , P3_U3819 , P3_U3820 , P3_U3821 , P3_U3822 , P3_U3823;
wire P3_U3824 , P3_U3825 , P3_U3826 , P3_U3827 , P3_U3828 , P3_U3829 , P3_U3830 , P3_U3831 , P3_U3832 , P3_U3833;
wire P3_U3834 , P3_U3835 , P3_U3836 , P3_U3837 , P3_U3838 , P3_U3839 , P3_U3840 , P3_U3841 , P3_U3842 , P3_U3843;
wire P3_U3844 , P3_U3845 , P3_U3846 , P3_U3847 , P3_U3848 , P3_U3849 , P3_U3850 , P3_U3851 , P3_U3852 , P3_U3853;
wire P3_U3854 , P3_U3855 , P3_U3856 , P3_U3857 , P3_U3858 , P3_U3859 , P3_U3860 , P3_U3861 , P3_U3862 , P3_U3863;
wire P3_U3864 , P3_U3865 , P3_U3866 , P3_U3867 , P3_U3868 , P3_U3869 , P3_U3870 , P3_U3871 , P3_U3872 , P3_U3873;
wire P3_U3874 , P3_U3875 , P3_U3876 , P3_U3877 , P3_U3878 , P3_U3879 , P3_U3880 , P3_U3881 , P3_U3882 , P3_U3883;
wire P3_U3884 , P3_U3885 , P3_U3886 , P3_U3887 , P3_U3888 , P3_U3889 , P3_U3890 , P3_U3891 , P3_U3892 , P3_U3893;
wire P3_U3894 , P3_U3895 , P3_U3896 , P3_U3898 , P3_U3899 , P3_U3900 , P3_U3901 , P3_U3902 , P3_U3903 , P3_U3904;
wire P3_U3905 , P3_U3906 , P3_U3907 , P3_U3908 , P3_U3909 , P3_U3910 , P3_U3911 , P3_U3912 , P3_U3913 , P3_U3914;
wire P3_U3915 , P3_U3916 , P3_U3917 , P3_U3918 , P3_U3919 , P3_U3920 , P3_U3921 , P3_U3922 , P3_U3923 , P3_U3924;
wire P3_U3925 , P3_U3926 , P3_U3927 , P3_U3928 , P3_U3929 , P3_U3930 , P3_U3931 , P3_U3932 , P3_U3933 , P3_U3934;
wire P3_U3935 , P3_U3936 , P3_U3937 , P3_U3938 , P3_U3939 , P3_U3940 , P3_U3941 , P3_U3942 , P3_U3943 , P3_U3944;
wire P3_U3945 , P3_U3946 , P3_U3947 , P3_U3948 , P3_U3949 , P3_U3950 , P3_U3951 , P3_U3952 , P3_U3953 , P3_U3954;
wire P3_U3955 , P3_U3956 , P3_U3957 , P3_U3958 , P3_U3959 , P3_U3960 , P3_U3961 , P3_U3962 , P3_U3963 , P3_U3964;
wire P3_U3965 , P3_U3966 , P3_U3967 , P3_U3968 , P3_U3969 , P3_U3970 , P3_U3971 , P3_U3972 , P3_U3973 , P3_U3974;
wire P3_U3975 , P3_U3976 , P3_U3977 , P3_U3978 , P3_U3979 , P3_U3980 , P3_U3981 , P3_U3982 , P3_U3983 , P3_U3984;
wire P3_U3985 , P3_U3986 , P3_U3987 , P3_U3988 , P3_U3989 , P3_U3990 , P3_U3991 , P3_U3992 , P3_U3993 , P3_U3994;
wire P3_U3995 , P3_U3996 , P3_U3997 , P3_U3998 , P3_U3999 , P3_U4000 , P3_U4001 , P3_U4002 , P3_U4003 , P3_U4004;
wire P3_U4005 , P3_U4006 , P3_U4007 , P3_U4008 , P3_U4009 , P3_U4010 , P3_U4011 , P3_U4012 , P3_U4013 , P3_U4014;
wire P3_U4015 , P3_U4016 , P3_U4017 , P3_U4018 , P3_U4019 , P3_U4020 , P3_U4021 , P3_U4022 , P3_U4023 , P3_U4024;
wire P3_U4025 , P3_U4026 , P3_U4027 , P3_U4028 , P3_U4029 , P3_U4030 , P3_U4031 , P3_U4032 , P3_U4033 , P3_U4034;
wire P3_U4035 , P3_U4036 , P3_U4037 , P3_U4038 , P3_U4039 , P3_U4040 , P3_U4041 , P3_U4042 , P3_U4043 , P3_U4044;
wire P3_U4045 , P3_U4046 , P3_U4047 , P3_U4048 , P3_U4049 , P3_U4050 , P3_U4051 , P3_U4052 , P3_U4053 , P3_U4054;
wire P3_U4055 , P3_U4056 , P3_U4057 , P3_U4058 , P3_U4059 , P3_U4060 , P3_U4061 , P3_U4062 , P3_U4063 , P3_U4064;
wire P3_U4065 , P3_U4066 , P3_U4067 , P3_U4068 , P3_U4069 , P3_U4070 , P3_U4071 , P3_U4072 , P3_U4073 , P3_U4074;
wire P3_U4075 , P3_U4076 , P3_U4077 , P3_U4078 , P3_U4079 , P3_U4080 , P3_U4081 , P3_U4082 , P3_U4083 , P3_U4084;
wire P3_U4085 , P3_U4086 , P3_U4087 , P3_U4088 , P3_U4089 , P3_U4090 , P3_U4091 , P3_U4092 , P3_U4093 , P3_U4094;
wire P3_U4095 , P3_U4096 , P3_U4097 , P3_U4098 , P3_U4099 , P3_U4100 , P3_U4101 , P3_U4102 , P3_U4103 , P3_U4104;
wire P3_U4105 , P3_U4106 , P3_U4107 , P3_U4108 , P3_U4109 , P3_U4110 , P3_U4111 , P3_U4112 , P3_U4113 , P3_U4114;
wire P3_U4115 , P3_U4116 , P3_U4117 , P3_U4118 , P3_U4119 , P3_U4120 , P3_U4121 , P3_U4122 , P3_U4123 , P3_U4124;
wire P3_U4125 , P3_U4126 , P3_U4127 , P3_U4128 , P3_U4129 , P3_U4130 , P3_U4131 , P3_U4132 , P3_U4133 , P3_U4134;
wire P3_U4135 , P3_U4136 , P3_U4137 , P3_U4138 , P3_U4139 , P3_U4140 , P3_U4141 , P3_U4142 , P3_U4143 , P3_U4144;
wire P3_U4145 , P3_U4146 , P3_U4147 , P3_U4148 , P3_U4149 , P3_U4150 , P3_U4151 , P3_U4152 , P3_U4153 , P3_U4154;
wire P3_U4155 , P3_U4156 , P3_U4157 , P3_U4158 , P3_U4159 , P3_U4160 , P3_U4161 , P3_U4162 , P3_U4163 , P3_U4164;
wire P3_U4165 , P3_U4166 , P3_U4167 , P3_U4168 , P3_U4169 , P3_U4170 , P3_U4171 , P3_U4172 , P3_U4173 , P3_U4174;
wire P3_U4175 , P3_U4176 , P3_U4177 , P3_U4178 , P3_U4179 , P3_U4180 , P3_U4181 , P3_U4182 , P3_U4183 , P3_U4184;
wire P3_U4185 , P3_U4186 , P3_U4187 , P3_U4188 , P3_U4189 , P3_U4190 , P3_U4191 , P3_U4192 , P3_U4193 , P3_U4194;
wire P3_U4195 , P3_U4196 , P3_U4197 , P3_U4198 , P3_U4199 , P3_U4200 , P3_U4201 , P3_U4202 , P3_U4203 , P3_U4204;
wire P3_U4205 , P3_U4206 , P3_U4207 , P3_U4208 , P3_U4209 , P3_U4210 , P3_U4211 , P3_U4212 , P3_U4213 , P3_U4214;
wire P3_U4215 , P3_U4216 , P3_U4217 , P3_U4218 , P3_U4219 , P3_U4220 , P3_U4221 , P3_U4222 , P3_U4223 , P3_U4224;
wire P3_U4225 , P3_U4226 , P3_U4227 , P3_U4228 , P3_U4229 , P3_U4230 , P3_U4231 , P3_U4232 , P3_U4233 , P3_U4234;
wire P3_U4235 , P3_U4236 , P3_U4237 , P3_U4238 , P3_U4239 , P3_U4240 , P3_U4241 , P3_U4242 , P3_U4243 , P3_U4244;
wire P3_U4245 , P3_U4246 , P3_U4247 , P3_U4248 , P3_U4249 , P3_U4250 , P3_U4251 , P3_U4252 , P3_U4253 , P3_U4254;
wire P3_U4255 , P3_U4256 , P3_U4257 , P3_U4258 , P3_U4259 , P3_U4260 , P3_U4261 , P3_U4262 , P3_U4263 , P3_U4264;
wire P3_U4265 , P3_U4266 , P3_U4267 , P3_U4268 , P3_U4269 , P3_U4270 , P3_U4271 , P3_U4272 , P3_U4273 , P3_U4274;
wire P3_U4275 , P3_U4276 , P3_U4277 , P3_U4278 , P3_U4279 , P3_U4280 , P3_U4281 , P3_U4282 , P3_U4283 , P3_U4284;
wire P3_U4285 , P3_U4286 , P3_U4287 , P3_U4288 , P3_U4289 , P3_U4290 , P3_U4291 , P3_U4292 , P3_U4293 , P3_U4294;
wire P3_U4295 , P3_U4296 , P3_U4297 , P3_U4298 , P3_U4299 , P3_U4300 , P3_U4301 , P3_U4302 , P3_U4303 , P3_U4304;
wire P3_U4305 , P3_U4306 , P3_U4307 , P3_U4308 , P3_U4309 , P3_U4310 , P3_U4311 , P3_U4312 , P3_U4313 , P3_U4314;
wire P3_U4315 , P3_U4316 , P3_U4317 , P3_U4318 , P3_U4319 , P3_U4320 , P3_U4321 , P3_U4322 , P3_U4323 , P3_U4324;
wire P3_U4325 , P3_U4326 , P3_U4327 , P3_U4328 , P3_U4329 , P3_U4330 , P3_U4331 , P3_U4332 , P3_U4333 , P3_U4334;
wire P3_U4335 , P3_U4336 , P3_U4337 , P3_U4338 , P3_U4339 , P3_U4340 , P3_U4341 , P3_U4342 , P3_U4343 , P3_U4344;
wire P3_U4345 , P3_U4346 , P3_U4347 , P3_U4348 , P3_U4349 , P3_U4350 , P3_U4351 , P3_U4352 , P3_U4353 , P3_U4354;
wire P3_U4355 , P3_U4356 , P3_U4357 , P3_U4358 , P3_U4359 , P3_U4360 , P3_U4361 , P3_U4362 , P3_U4363 , P3_U4364;
wire P3_U4365 , P3_U4366 , P3_U4367 , P3_U4368 , P3_U4369 , P3_U4370 , P3_U4371 , P3_U4372 , P3_U4373 , P3_U4374;
wire P3_U4375 , P3_U4376 , P3_U4377 , P3_U4378 , P3_U4379 , P3_U4380 , P3_U4381 , P3_U4382 , P3_U4383 , P3_U4384;
wire P3_U4385 , P3_U4386 , P3_U4387 , P3_U4388 , P3_U4389 , P3_U4390 , P3_U4391 , P3_U4392 , P3_U4393 , P3_U4394;
wire P3_U4395 , P3_U4396 , P3_U4397 , P3_U4398 , P3_U4399 , P3_U4400 , P3_U4401 , P3_U4402 , P3_U4403 , P3_U4404;
wire P3_U4405 , P3_U4406 , P3_U4407 , P3_U4408 , P3_U4409 , P3_U4410 , P3_U4411 , P3_U4412 , P3_U4413 , P3_U4414;
wire P3_U4415 , P3_U4416 , P3_U4417 , P3_U4418 , P3_U4419 , P3_U4420 , P3_U4421 , P3_U4422 , P3_U4423 , P3_U4424;
wire P3_U4425 , P3_U4426 , P3_U4427 , P3_U4428 , P3_U4429 , P3_U4430 , P3_U4431 , P3_U4432 , P3_U4433 , P3_U4434;
wire P3_U4435 , P3_U4436 , P3_U4437 , P3_U4438 , P3_U4439 , P3_U4440 , P3_U4441 , P3_U4442 , P3_U4443 , P3_U4444;
wire P3_U4445 , P3_U4446 , P3_U4447 , P3_U4448 , P3_U4449 , P3_U4450 , P3_U4451 , P3_U4452 , P3_U4453 , P3_U4454;
wire P3_U4455 , P3_U4456 , P3_U4457 , P3_U4458 , P3_U4459 , P3_U4460 , P3_U4461 , P3_U4462 , P3_U4463 , P3_U4464;
wire P3_U4465 , P3_U4466 , P3_U4467 , P3_U4468 , P3_U4469 , P3_U4470 , P3_U4471 , P3_U4472 , P3_U4473 , P3_U4474;
wire P3_U4475 , P3_U4476 , P3_U4477 , P3_U4478 , P3_U4479 , P3_U4480 , P3_U4481 , P3_U4482 , P3_U4483 , P3_U4484;
wire P3_U4485 , P3_U4486 , P3_U4487 , P3_U4488 , P3_U4489 , P3_U4490 , P3_U4491 , P3_U4492 , P3_U4493 , P3_U4494;
wire P3_U4495 , P3_U4496 , P3_U4497 , P3_U4498 , P3_U4499 , P3_U4500 , P3_U4501 , P3_U4502 , P3_U4503 , P3_U4504;
wire P3_U4505 , P3_U4506 , P3_U4507 , P3_U4508 , P3_U4509 , P3_U4510 , P3_U4511 , P3_U4512 , P3_U4513 , P3_U4514;
wire P3_U4515 , P3_U4516 , P3_U4517 , P3_U4518 , P3_U4519 , P3_U4520 , P3_U4521 , P3_U4522 , P3_U4523 , P3_U4524;
wire P3_U4525 , P3_U4526 , P3_U4527 , P3_U4528 , P3_U4529 , P3_U4530 , P3_U4531 , P3_U4532 , P3_U4533 , P3_U4534;
wire P3_U4535 , P3_U4536 , P3_U4537 , P3_U4538 , P3_U4539 , P3_U4540 , P3_U4541 , P3_U4542 , P3_U4543 , P3_U4544;
wire P3_U4545 , P3_U4546 , P3_U4547 , P3_U4548 , P3_U4549 , P3_U4550 , P3_U4551 , P3_U4552 , P3_U4553 , P3_U4554;
wire P3_U4555 , P3_U4556 , P3_U4557 , P3_U4558 , P3_U4559 , P3_U4560 , P3_U4561 , P3_U4562 , P3_U4563 , P3_U4564;
wire P3_U4565 , P3_U4566 , P3_U4567 , P3_U4568 , P3_U4569 , P3_U4570 , P3_U4571 , P3_U4572 , P3_U4573 , P3_U4574;
wire P3_U4575 , P3_U4576 , P3_U4577 , P3_U4578 , P3_U4579 , P3_U4580 , P3_U4581 , P3_U4582 , P3_U4583 , P3_U4584;
wire P3_U4585 , P3_U4586 , P3_U4587 , P3_U4588 , P3_U4589 , P3_U4590 , P3_U4591 , P3_U4592 , P3_U4593 , P3_U4594;
wire P3_U4595 , P3_U4596 , P3_U4597 , P3_U4598 , P3_U4599 , P3_U4600 , P3_U4601 , P3_U4602 , P3_U4603 , P3_U4604;
wire P3_U4605 , P3_U4606 , P3_U4607 , P3_U4608 , P3_U4609 , P3_U4610 , P3_U4611 , P3_U4612 , P3_U4613 , P3_U4614;
wire P3_U4615 , P3_U4616 , P3_U4617 , P3_U4618 , P3_U4619 , P3_U4620 , P3_U4621 , P3_U4622 , P3_U4623 , P3_U4624;
wire P3_U4625 , P3_U4626 , P3_U4627 , P3_U4628 , P3_U4629 , P3_U4630 , P3_U4631 , P3_U4632 , P3_U4633 , P3_U4634;
wire P3_U4635 , P3_U4636 , P3_U4637 , P3_U4638 , P3_U4639 , P3_U4640 , P3_U4641 , P3_U4642 , P3_U4643 , P3_U4644;
wire P3_U4645 , P3_U4646 , P3_U4647 , P3_U4648 , P3_U4649 , P3_U4650 , P3_U4651 , P3_U4652 , P3_U4653 , P3_U4654;
wire P3_U4655 , P3_U4656 , P3_U4657 , P3_U4658 , P3_U4659 , P3_U4660 , P3_U4661 , P3_U4662 , P3_U4663 , P3_U4664;
wire P3_U4665 , P3_U4666 , P3_U4667 , P3_U4668 , P3_U4669 , P3_U4670 , P3_U4671 , P3_U4672 , P3_U4673 , P3_U4674;
wire P3_U4675 , P3_U4676 , P3_U4677 , P3_U4678 , P3_U4679 , P3_U4680 , P3_U4681 , P3_U4682 , P3_U4683 , P3_U4684;
wire P3_U4685 , P3_U4686 , P3_U4687 , P3_U4688 , P3_U4689 , P3_U4690 , P3_U4691 , P3_U4692 , P3_U4693 , P3_U4694;
wire P3_U4695 , P3_U4696 , P3_U4697 , P3_U4698 , P3_U4699 , P3_U4700 , P3_U4701 , P3_U4702 , P3_U4703 , P3_U4704;
wire P3_U4705 , P3_U4706 , P3_U4707 , P3_U4708 , P3_U4709 , P3_U4710 , P3_U4711 , P3_U4712 , P3_U4713 , P3_U4714;
wire P3_U4715 , P3_U4716 , P3_U4717 , P3_U4718 , P3_U4719 , P3_U4720 , P3_U4721 , P3_U4722 , P3_U4723 , P3_U4724;
wire P3_U4725 , P3_U4726 , P3_U4727 , P3_U4728 , P3_U4729 , P3_U4730 , P3_U4731 , P3_U4732 , P3_U4733 , P3_U4734;
wire P3_U4735 , P3_U4736 , P3_U4737 , P3_U4738 , P3_U4739 , P3_U4740 , P3_U4741 , P3_U4742 , P3_U4743 , P3_U4744;
wire P3_U4745 , P3_U4746 , P3_U4747 , P3_U4748 , P3_U4749 , P3_U4750 , P3_U4751 , P3_U4752 , P3_U4753 , P3_U4754;
wire P3_U4755 , P3_U4756 , P3_U4757 , P3_U4758 , P3_U4759 , P3_U4760 , P3_U4761 , P3_U4762 , P3_U4763 , P3_U4764;
wire P3_U4765 , P3_U4766 , P3_U4767 , P3_U4768 , P3_U4769 , P3_U4770 , P3_U4771 , P3_U4772 , P3_U4773 , P3_U4774;
wire P3_U4775 , P3_U4776 , P3_U4777 , P3_U4778 , P3_U4779 , P3_U4780 , P3_U4781 , P3_U4782 , P3_U4783 , P3_U4784;
wire P3_U4785 , P3_U4786 , P3_U4787 , P3_U4788 , P3_U4789 , P3_U4790 , P3_U4791 , P3_U4792 , P3_U4793 , P3_U4794;
wire P3_U4795 , P3_U4796 , P3_U4797 , P3_U4798 , P3_U4799 , P3_U4800 , P3_U4801 , P3_U4802 , P3_U4803 , P3_U4804;
wire P3_U4805 , P3_U4806 , P3_U4807 , P3_U4808 , P3_U4809 , P3_U4810 , P3_U4811 , P3_U4812 , P3_U4813 , P3_U4814;
wire P3_U4815 , P3_U4816 , P3_U4817 , P3_U4818 , P3_U4819 , P3_U4820 , P3_U4821 , P3_U4822 , P3_U4823 , P3_U4824;
wire P3_U4825 , P3_U4826 , P3_U4827 , P3_U4828 , P3_U4829 , P3_U4830 , P3_U4831 , P3_U4832 , P3_U4833 , P3_U4834;
wire P3_U4835 , P3_U4836 , P3_U4837 , P3_U4838 , P3_U4839 , P3_U4840 , P3_U4841 , P3_U4842 , P3_U4843 , P3_U4844;
wire P3_U4845 , P3_U4846 , P3_U4847 , P3_U4848 , P3_U4849 , P3_U4850 , P3_U4851 , P3_U4852 , P3_U4853 , P3_U4854;
wire P3_U4855 , P3_U4856 , P3_U4857 , P3_U4858 , P3_U4859 , P3_U4860 , P3_U4861 , P3_U4862 , P3_U4863 , P3_U4864;
wire P3_U4865 , P3_U4866 , P3_U4867 , P3_U4868 , P3_U4869 , P3_U4870 , P3_U4871 , P3_U4872 , P3_U4873 , P3_U4874;
wire P3_U4875 , P3_U4876 , P3_U4877 , P3_U4878 , P3_U4879 , P3_U4880 , P3_U4881 , P3_U4882 , P3_U4883 , P3_U4884;
wire P3_U4885 , P3_U4886 , P3_U4887 , P3_U4888 , P3_U4889 , P3_U4890 , P3_U4891 , P3_U4892 , P3_U4893 , P3_U4894;
wire P3_U4895 , P3_U4896 , P3_U4897 , P3_U4898 , P3_U4899 , P3_U4900 , P3_U4901 , P3_U4902 , P3_U4903 , P3_U4904;
wire P3_U4905 , P3_U4906 , P3_U4907 , P3_U4908 , P3_U4909 , P3_U4910 , P3_U4911 , P3_U4912 , P3_U4913 , P3_U4914;
wire P3_U4915 , P3_U4916 , P3_U4917 , P3_U4918 , P3_U4919 , P3_U4920 , P3_U4921 , P3_U4922 , P3_U4923 , P3_U4924;
wire P3_U4925 , P3_U4926 , P3_U4927 , P3_U4928 , P3_U4929 , P3_U4930 , P3_U4931 , P3_U4932 , P3_U4933 , P3_U4934;
wire P3_U4935 , P3_U4936 , P3_U4937 , P3_U4938 , P3_U4939 , P3_U4940 , P3_U4941 , P3_U4942 , P3_U4943 , P3_U4944;
wire P3_U4945 , P3_U4946 , P3_U4947 , P3_U4948 , P3_U4949 , P3_U4950 , P3_U4951 , P3_U4952 , P3_U4953 , P3_U4954;
wire P3_U4955 , P3_U4956 , P3_U4957 , P3_U4958 , P3_U4959 , P3_U4960 , P3_U4961 , P3_U4962 , P3_U4963 , P3_U4964;
wire P3_U4965 , P3_U4966 , P3_U4967 , P3_U4968 , P3_U4969 , P3_U4970 , P3_U4971 , P3_U4972 , P3_U4973 , P3_U4974;
wire P3_U4975 , P3_U4976 , P3_U4977 , P3_U4978 , P3_U4979 , P3_U4980 , P3_U4981 , P3_U4982 , P3_U4983 , P3_U4984;
wire P3_U4985 , P3_U4986 , P3_U4987 , P3_U4988 , P3_U4989 , P3_U4990 , P3_U4991 , P3_U4992 , P3_U4993 , P3_U4994;
wire P3_U4995 , P3_U4996 , P3_U4997 , P3_U4998 , P3_U4999 , P3_U5000 , P3_U5001 , P3_U5002 , P3_U5003 , P3_U5004;
wire P3_U5005 , P3_U5006 , P3_U5007 , P3_U5008 , P3_U5009 , P3_U5010 , P3_U5011 , P3_U5012 , P3_U5013 , P3_U5014;
wire P3_U5015 , P3_U5016 , P3_U5017 , P3_U5018 , P3_U5019 , P3_U5020 , P3_U5021 , P3_U5022 , P3_U5023 , P3_U5024;
wire P3_U5025 , P3_U5026 , P3_U5027 , P3_U5028 , P3_U5029 , P3_U5030 , P3_U5031 , P3_U5032 , P3_U5033 , P3_U5034;
wire P3_U5035 , P3_U5036 , P3_U5037 , P3_U5038 , P3_U5039 , P3_U5040 , P3_U5041 , P3_U5042 , P3_U5043 , P3_U5044;
wire P3_U5045 , P3_U5046 , P3_U5047 , P3_U5048 , P3_U5049 , P3_U5050 , P3_U5051 , P3_U5052 , P3_U5053 , P3_U5054;
wire P3_U5055 , P3_U5056 , P3_U5057 , P3_U5058 , P3_U5059 , P3_U5060 , P3_U5061 , P3_U5062 , P3_U5063 , P3_U5064;
wire P3_U5065 , P3_U5066 , P3_U5067 , P3_U5068 , P3_U5069 , P3_U5070 , P3_U5071 , P3_U5072 , P3_U5073 , P3_U5074;
wire P3_U5075 , P3_U5076 , P3_U5077 , P3_U5078 , P3_U5079 , P3_U5080 , P3_U5081 , P3_U5082 , P3_U5083 , P3_U5084;
wire P3_U5085 , P3_U5086 , P3_U5087 , P3_U5088 , P3_U5089 , P3_U5090 , P3_U5091 , P3_U5092 , P3_U5093 , P3_U5094;
wire P3_U5095 , P3_U5096 , P3_U5097 , P3_U5098 , P3_U5099 , P3_U5100 , P3_U5101 , P3_U5102 , P3_U5103 , P3_U5104;
wire P3_U5105 , P3_U5106 , P3_U5107 , P3_U5108 , P3_U5109 , P3_U5110 , P3_U5111 , P3_U5112 , P3_U5113 , P3_U5114;
wire P3_U5115 , P3_U5116 , P3_U5117 , P3_U5118 , P3_U5119 , P3_U5120 , P3_U5121 , P3_U5122 , P3_U5123 , P3_U5124;
wire P3_U5125 , P3_U5126 , P3_U5127 , P3_U5128 , P3_U5129 , P3_U5130 , P3_U5131 , P3_U5132 , P3_U5133 , P3_U5134;
wire P3_U5135 , P3_U5136 , P3_U5137 , P3_U5138 , P3_U5139 , P3_U5140 , P3_U5141 , P3_U5142 , P3_U5143 , P3_U5144;
wire P3_U5145 , P3_U5146 , P3_U5147 , P3_U5148 , P3_U5149 , P3_U5150 , P3_U5151 , P3_U5152 , P3_U5153 , P3_U5154;
wire P3_U5155 , P3_U5156 , P3_U5157 , P3_U5158 , P3_U5159 , P3_U5160 , P3_U5161 , P3_U5162 , P3_U5163 , P3_U5164;
wire P3_U5165 , P3_U5166 , P3_U5167 , P3_U5168 , P3_U5169 , P3_U5170 , P3_U5171 , P3_U5172 , P3_U5173 , P3_U5174;
wire P3_U5175 , P3_U5176 , P3_U5177 , P3_U5178 , P3_U5179 , P3_U5180 , P3_U5181 , P3_U5182 , P3_U5183 , P3_U5184;
wire P3_U5185 , P3_U5186 , P3_U5187 , P3_U5188 , P3_U5189 , P3_U5190 , P3_U5191 , P3_U5192 , P3_U5193 , P3_U5194;
wire P3_U5195 , P3_U5196 , P3_U5197 , P3_U5198 , P3_U5199 , P3_U5200 , P3_U5201 , P3_U5202 , P3_U5203 , P3_U5204;
wire P3_U5205 , P3_U5206 , P3_U5207 , P3_U5208 , P3_U5209 , P3_U5210 , P3_U5211 , P3_U5212 , P3_U5213 , P3_U5214;
wire P3_U5215 , P3_U5216 , P3_U5217 , P3_U5218 , P3_U5219 , P3_U5220 , P3_U5221 , P3_U5222 , P3_U5223 , P3_U5224;
wire P3_U5225 , P3_U5226 , P3_U5227 , P3_U5228 , P3_U5229 , P3_U5230 , P3_U5231 , P3_U5232 , P3_U5233 , P3_U5234;
wire P3_U5235 , P3_U5236 , P3_U5237 , P3_U5238 , P3_U5239 , P3_U5240 , P3_U5241 , P3_U5242 , P3_U5243 , P3_U5244;
wire P3_U5245 , P3_U5246 , P3_U5247 , P3_U5248 , P3_U5249 , P3_U5250 , P3_U5251 , P3_U5252 , P3_U5253 , P3_U5254;
wire P3_U5255 , P3_U5256 , P3_U5257 , P3_U5258 , P3_U5259 , P3_U5260 , P3_U5261 , P3_U5262 , P3_U5263 , P3_U5264;
wire P3_U5265 , P3_U5266 , P3_U5267 , P3_U5268 , P3_U5269 , P3_U5270 , P3_U5271 , P3_U5272 , P3_U5273 , P3_U5274;
wire P3_U5275 , P3_U5276 , P3_U5277 , P3_U5278 , P3_U5279 , P3_U5280 , P3_U5281 , P3_U5282 , P3_U5283 , P3_U5284;
wire P3_U5285 , P3_U5286 , P3_U5287 , P3_U5288 , P3_U5289 , P3_U5290 , P3_U5291 , P3_U5292 , P3_U5293 , P3_U5294;
wire P3_U5295 , P3_U5296 , P3_U5297 , P3_U5298 , P3_U5299 , P3_U5300 , P3_U5301 , P3_U5302 , P3_U5303 , P3_U5304;
wire P3_U5305 , P3_U5306 , P3_U5307 , P3_U5308 , P3_U5309 , P3_U5310 , P3_U5311 , P3_U5312 , P3_U5313 , P3_U5314;
wire P3_U5315 , P3_U5316 , P3_U5317 , P3_U5318 , P3_U5319 , P3_U5320 , P3_U5321 , P3_U5322 , P3_U5323 , P3_U5324;
wire P3_U5325 , P3_U5326 , P3_U5327 , P3_U5328 , P3_U5329 , P3_U5330 , P3_U5331 , P3_U5332 , P3_U5333 , P3_U5334;
wire P3_U5335 , P3_U5336 , P3_U5337 , P3_U5338 , P3_U5339 , P3_U5340 , P3_U5341 , P3_U5342 , P3_U5343 , P3_U5344;
wire P3_U5345 , P3_U5346 , P3_U5347 , P3_U5348 , P3_U5349 , P3_U5350 , P3_U5351 , P3_U5352 , P3_U5353 , P3_U5354;
wire P3_U5355 , P3_U5356 , P3_U5357 , P3_U5358 , P3_U5359 , P3_U5360 , P3_U5361 , P3_U5362 , P3_U5363 , P3_U5364;
wire P3_U5365 , P3_U5366 , P3_U5367 , P3_U5368 , P3_U5369 , P3_U5370 , P3_U5371 , P3_U5372 , P3_U5373 , P3_U5374;
wire P3_U5375 , P3_U5376 , P3_U5377 , P3_U5378 , P3_U5379 , P3_U5380 , P3_U5381 , P3_U5382 , P3_U5383 , P3_U5384;
wire P3_U5385 , P3_U5386 , P3_U5387 , P3_U5388 , P3_U5389 , P3_U5390 , P3_U5391 , P3_U5392 , P3_U5393 , P3_U5394;
wire P3_U5395 , P3_U5396 , P3_U5397 , P3_U5398 , P3_U5399 , P3_U5400 , P3_U5401 , P3_U5402 , P3_U5403 , P3_U5404;
wire P3_U5405 , P3_U5406 , P3_U5407 , P3_U5408 , P3_U5409 , P3_U5410 , P3_U5411 , P3_U5412 , P3_U5413 , P3_U5414;
wire P3_U5415 , P3_U5416 , P3_U5417 , P3_U5418 , P3_U5419 , P3_U5420 , P3_U5421 , P3_U5422 , P3_U5423 , P3_U5424;
wire P3_U5425 , P3_U5426 , P3_U5427 , P3_U5428 , P3_U5429 , P3_U5430 , P3_U5431 , P3_U5432 , P3_U5433 , P3_U5434;
wire P3_U5435 , P3_U5436 , P3_U5437 , P3_U5438 , P3_U5439 , P3_U5440 , P3_U5441 , P3_U5442 , P3_U5443 , P3_U5444;
wire P3_U5445 , P3_U5446 , P3_U5447 , P3_U5448 , P3_U5449 , P3_U5450 , P3_U5451 , P3_U5452 , P3_U5453 , P3_U5454;
wire P3_U5455 , P3_U5456 , P3_U5457 , P3_U5458 , P3_U5459 , P3_U5460 , P3_U5461 , P3_U5462 , P3_U5463 , P3_U5464;
wire P3_U5465 , P3_U5466 , P3_U5467 , P3_U5468 , P3_U5469 , P3_U5470 , P3_U5471 , P3_U5472 , P3_U5473 , P3_U5474;
wire P3_U5475 , P3_U5476 , P3_U5477 , P3_U5478 , P3_U5479 , P3_U5480 , P3_U5481 , P3_U5482 , P3_U5483 , P3_U5484;
wire P3_U5485 , P3_U5486 , P3_U5487 , P3_U5488 , P3_U5489 , P3_U5490 , P3_U5491 , P3_U5492 , P3_U5493 , P3_U5494;
wire P3_U5495 , P3_U5496 , P3_U5497 , P3_U5498 , P3_U5499 , P3_U5500 , P3_U5501 , P3_U5502 , P3_U5503 , P3_U5504;
wire P3_U5505 , P3_U5506 , P3_U5507 , P3_U5508 , P3_U5509 , P3_U5510 , P3_U5511 , P3_U5512 , P3_U5513 , P3_U5514;
wire P3_U5515 , P3_U5516 , P3_U5517 , P3_U5518 , P3_U5519 , P3_U5520 , P3_U5521 , P3_U5522 , P3_U5523 , P3_U5524;
wire P3_U5525 , P3_U5526 , P3_U5527 , P3_U5528 , P3_U5529 , P3_U5530 , P3_U5531 , P3_U5532 , P3_U5533 , P3_U5534;
wire P3_U5535 , P3_U5536 , P3_U5537 , P3_U5538 , P3_U5539 , P3_U5540 , P3_U5541 , P3_U5542 , P3_U5543 , P3_U5544;
wire P3_U5545 , P3_U5546 , P3_U5547 , P3_U5548 , P3_U5549 , P3_U5550 , P3_U5551 , P3_U5552 , P3_U5553 , P3_U5554;
wire P3_U5555 , P3_U5556 , P3_U5557 , P3_U5558 , P3_U5559 , P3_U5560 , P3_U5561 , P3_U5562 , P3_U5563 , P3_U5564;
wire P3_U5565 , P3_U5566 , P3_U5567 , P3_U5568 , P3_U5569 , P3_U5570 , P3_U5571 , P3_U5572 , P3_U5573 , P3_U5574;
wire P3_U5575 , P3_U5576 , P3_U5577 , P3_U5578 , P3_U5579 , P3_U5580 , P3_U5581 , P3_U5582 , P3_U5583 , P3_U5584;
wire P3_U5585 , P3_U5586 , P3_U5587 , P3_U5588 , P3_U5589 , P3_U5590 , P3_U5591 , P3_U5592 , P3_U5593 , P3_U5594;
wire P3_U5595 , P3_U5596 , P3_U5597 , P3_U5598 , P3_U5599 , P3_U5600 , P3_U5601 , P3_U5602 , P3_U5603 , P3_U5604;
wire P3_U5605 , P3_U5606 , P3_U5607 , P3_U5608 , P3_U5609 , P3_U5610 , P3_U5611 , P3_U5612 , P3_U5613 , P3_U5614;
wire P3_U5615 , P3_U5616 , P3_U5617 , P3_U5618 , P3_U5619 , P3_U5620 , P3_U5621 , P3_U5622 , P3_U5623 , P3_U5624;
wire P3_U5625 , P3_U5626 , P3_U5627 , P3_U5628 , P3_U5629 , P3_U5630 , P3_U5631 , P3_U5632 , P3_U5633 , P3_U5634;
wire P3_U5635 , P3_U5636 , P3_U5637 , P3_U5638 , P3_U5639 , P3_U5640 , P3_U5641 , P3_U5642 , P3_U5643 , P3_U5644;
wire P3_U5645 , P3_U5646 , P3_U5647 , P3_U5648 , P3_U5649 , P3_U5650 , P3_U5651 , P3_U5652 , P3_U5653 , P3_U5654;
wire P3_U5655 , P3_U5656 , P3_U5657 , P3_U5658 , P3_U5659 , P3_U5660 , P3_U5661 , P3_U5662 , P3_U5663 , P3_U5664;
wire P3_U5665 , P3_U5666 , P3_U5667 , P3_U5668 , P3_U5669 , P3_U5670 , P3_U5671 , P3_U5672 , P3_U5673 , P3_U5674;
wire P3_U5675 , P3_U5676 , P3_U5677 , P3_U5678 , P3_U5679 , P3_U5680 , P3_U5681 , P3_U5682 , P3_U5683 , P3_U5684;
wire P3_U5685 , P3_U5686 , P3_U5687 , P3_U5688 , P3_U5689 , P3_U5690 , P3_U5691 , P3_U5692 , P3_U5693 , P3_U5694;
wire P3_U5695 , P3_U5696 , P3_U5697 , P3_U5698 , P3_U5699 , P3_U5700 , P3_U5701 , P3_U5702 , P3_U5703 , P3_U5704;
wire P3_U5705 , P3_U5706 , P3_U5707 , P3_U5708 , P3_U5709 , P3_U5710 , P3_U5711 , P3_U5712 , P3_U5713 , P3_U5714;
wire P3_U5715 , P3_U5716 , P3_U5717 , P3_U5718 , P3_U5719 , P3_U5720 , P3_U5721 , P3_U5722 , P3_U5723 , P3_U5724;
wire P3_U5725 , P3_U5726 , P3_U5727 , P3_U5728 , P3_U5729 , P3_U5730 , P3_U5731 , P3_U5732 , P3_U5733 , P3_U5734;
wire P3_U5735 , P3_U5736 , P3_U5737 , P3_U5738 , P3_U5739 , P3_U5740 , P3_U5741 , P3_U5742 , P3_U5743 , P3_U5744;
wire P3_U5745 , P3_U5746 , P3_U5747 , P3_U5748 , P3_U5749 , P3_U5750 , P3_U5751 , P3_U5752 , P3_U5753 , P3_U5754;
wire P3_U5755 , P3_U5756 , P3_U5757 , P3_U5758 , P3_U5759 , P3_U5760 , P3_U5761 , P3_U5762 , P3_U5763 , P3_U5764;
wire P3_U5765 , P3_U5766 , P3_U5767 , P3_U5768 , P3_U5769 , P3_U5770 , P3_U5771 , P3_U5772 , P3_U5773 , P3_U5774;
wire P3_U5775 , P3_U5776 , P3_U5777 , P3_U5778 , P3_U5779 , P3_U5780 , P3_U5781 , P3_U5782 , P3_U5783 , P3_U5784;
wire P3_U5785 , P3_U5786 , P3_U5787 , P3_U5788 , P3_U5789 , P3_U5790 , P3_U5791 , P3_U5792 , P3_U5793 , P3_U5794;
wire P3_U5795 , P3_U5796 , P3_U5797 , P3_U5798 , P3_U5799 , P3_U5800 , P3_U5801 , P3_U5802 , P3_U5803 , P3_U5804;
wire P3_U5805 , P3_U5806 , P3_U5807 , P3_U5808 , P3_U5809 , P3_U5810 , P3_U5811 , P3_U5812 , P3_U5813 , P3_U5814;
wire P3_U5815 , P3_U5816 , P3_U5817 , P3_U5818 , P3_U5819 , P3_U5820 , P3_U5821 , P3_U5822 , P3_U5823 , P3_U5824;
wire P3_U5825 , P3_U5826 , P3_U5827 , P3_U5828 , P3_U5829 , P3_U5830 , P3_U5831 , P3_U5832 , P3_U5833 , P3_U5834;
wire P3_U5835 , P3_U5836 , P3_U5837 , P3_U5838 , P3_U5839 , P3_U5840 , P3_U5841 , P3_U5842 , P3_U5843 , P3_U5844;
wire P3_U5845 , P3_U5846 , P3_U5847 , P3_U5848 , P3_U5849 , P3_U5850 , P3_U5851 , P3_U5852 , P3_U5853 , P3_U5854;
wire P3_U5855 , P3_U5856 , P3_U5857 , P3_U5858 , P3_U5859 , P3_U5860 , P3_U5861 , P3_U5862 , P3_U5863 , P3_U5864;
wire P3_U5865 , P3_U5866 , P3_U5867 , P3_U5868 , P3_U5869 , P3_U5870 , P3_U5871 , P3_U5872 , P3_U5873 , P3_U5874;
wire P3_U5875 , P3_U5876 , P3_U5877 , P3_U5878 , P3_U5879 , P3_U5880 , P3_U5881 , P3_U5882 , P3_U5883 , P3_U5884;
wire P3_U5885 , P3_U5886 , P3_U5887 , P3_U5888 , P3_U5889 , P3_U5890 , P3_U5891 , P3_U5892 , P3_U5893 , P3_U5894;
wire P3_U5895 , P3_U5896 , P3_U5897 , P3_U5898 , P3_U5899 , P3_U5900 , P3_U5901 , P3_U5902 , P3_U5903 , P3_U5904;
wire P3_U5905 , P3_U5906 , P3_U5907 , P3_U5908 , P3_U5909 , P3_U5910 , P3_U5911 , P3_U5912 , P3_U5913 , P3_U5914;
wire P3_U5915 , P3_U5916 , P3_U5917 , P3_U5918 , P3_U5919 , P3_U5920 , P3_U5921 , P3_U5922 , P3_U5923 , P3_U5924;
wire P3_U5925 , P3_U5926 , P3_U5927 , P3_U5928 , P3_U5929 , P3_U5930 , P3_U5931 , P3_U5932 , P3_U5933 , P3_U5934;
wire P3_U5935 , P3_U5936 , P3_U5937 , P3_U5938 , P3_U5939 , P3_U5940 , P3_U5941 , P3_U5942 , P3_U5943 , P3_U5944;
wire P3_U5945 , P3_U5946 , P3_U5947 , P3_U5948 , P3_U5949 , P3_U5950 , P3_U5951 , P3_U5952 , P3_U5953 , P3_U5954;
wire P3_U5955 , P3_U5956 , P3_U5957 , P3_U5958 , P3_U5959 , P3_U5960 , P3_U5961 , P3_U5962 , P3_U5963 , P3_U5964;
wire P3_U5965 , P3_U5966 , P3_U5967 , P3_U5968 , P3_U5969 , P3_U5970 , P3_U5971 , P3_U5972 , P3_U5973 , P3_U5974;
wire P3_U5975 , P3_U5976 , P3_U5977 , P3_U5978 , P3_U5979 , P3_U5980 , P3_U5981 , P3_U5982 , P3_U5983 , P3_U5984;
wire P3_U5985 , P3_U5986 , P3_U5987 , P3_U5988 , P3_U5989 , P3_U5990 , P3_U5991 , P3_U5992 , P3_U5993 , P3_U5994;
wire P3_U5995 , P3_U5996 , P3_U5997 , P3_U5998 , P3_U5999 , P3_U6000 , P3_U6001 , P3_U6002 , P3_U6003 , P3_U6004;
wire P3_U6005 , P3_U6006 , P3_U6007 , P3_U6008 , P3_U6009 , P3_U6010 , P3_U6011 , P3_U6012 , P3_U6013 , P3_U6014;
wire P3_U6015 , P3_U6016 , P3_U6017 , P3_U6018 , P3_U6019 , P3_U6020 , P3_U6021 , P3_U6022 , P3_U6023 , P3_U6024;
wire P3_U6025 , P3_U6026 , P3_U6027 , P3_U6028 , P3_U6029 , P3_U6030 , P3_U6031 , P3_U6032 , P3_U6033 , P3_U6034;
wire P3_U6035 , P3_U6036 , P3_U6037 , P3_U6038 , P3_U6039 , P3_U6040 , P3_U6041 , P3_U6042 , P3_U6043 , P3_U6044;
wire P3_U6045 , P3_U6046 , P3_U6047 , P3_U6048 , P3_R1161_U448 , P3_R1161_U447 , P3_R1161_U446 , P3_R1161_U445 , P3_R1161_U444 , P3_R1161_U443;
wire P3_R1161_U442 , P3_R1161_U441 , P3_R1161_U440 , P3_R1161_U439 , P3_R1161_U438 , P3_R1161_U437 , P3_R1161_U436 , P3_R1161_U435 , P3_R1161_U434 , P3_R1161_U433;
wire P3_R1161_U432 , P3_R1161_U431 , P3_R1161_U430 , SUB_1605_U6 , SUB_1605_U7 , SUB_1605_U8 , SUB_1605_U9 , SUB_1605_U10 , SUB_1605_U11 , SUB_1605_U12;
wire SUB_1605_U13 , SUB_1605_U14 , SUB_1605_U15 , SUB_1605_U16 , SUB_1605_U17 , SUB_1605_U18 , SUB_1605_U19 , SUB_1605_U20 , SUB_1605_U21 , SUB_1605_U22;
wire SUB_1605_U23 , SUB_1605_U24 , SUB_1605_U25 , SUB_1605_U26 , SUB_1605_U27 , SUB_1605_U28 , SUB_1605_U29 , SUB_1605_U30 , SUB_1605_U31 , SUB_1605_U32;
wire SUB_1605_U33 , SUB_1605_U34 , SUB_1605_U35 , SUB_1605_U36 , SUB_1605_U37 , SUB_1605_U38 , SUB_1605_U39 , SUB_1605_U40 , SUB_1605_U41 , SUB_1605_U42;
wire SUB_1605_U43 , SUB_1605_U44 , SUB_1605_U45 , SUB_1605_U46 , SUB_1605_U47 , SUB_1605_U48 , SUB_1605_U49 , SUB_1605_U50 , SUB_1605_U51 , SUB_1605_U52;
wire SUB_1605_U53 , SUB_1605_U54 , SUB_1605_U55 , SUB_1605_U56 , SUB_1605_U57 , SUB_1605_U58 , SUB_1605_U59 , SUB_1605_U60 , SUB_1605_U61 , SUB_1605_U62;
wire SUB_1605_U63 , SUB_1605_U64 , SUB_1605_U65 , SUB_1605_U66 , SUB_1605_U67 , SUB_1605_U68 , SUB_1605_U69 , SUB_1605_U70 , SUB_1605_U71 , SUB_1605_U72;
wire SUB_1605_U73 , SUB_1605_U74 , SUB_1605_U75 , SUB_1605_U76 , SUB_1605_U77 , SUB_1605_U78 , SUB_1605_U79 , SUB_1605_U80 , SUB_1605_U81 , SUB_1605_U82;
wire SUB_1605_U83 , SUB_1605_U84 , SUB_1605_U85 , SUB_1605_U86 , SUB_1605_U87 , SUB_1605_U88 , SUB_1605_U89 , SUB_1605_U90 , SUB_1605_U91 , SUB_1605_U92;
wire SUB_1605_U93 , SUB_1605_U94 , SUB_1605_U95 , SUB_1605_U96 , SUB_1605_U97 , SUB_1605_U98 , SUB_1605_U99 , SUB_1605_U100 , SUB_1605_U101 , SUB_1605_U102;
wire SUB_1605_U103 , SUB_1605_U104 , SUB_1605_U105 , SUB_1605_U106 , SUB_1605_U107 , SUB_1605_U108 , SUB_1605_U109 , SUB_1605_U110 , SUB_1605_U111 , SUB_1605_U112;
wire SUB_1605_U113 , SUB_1605_U114 , SUB_1605_U115 , SUB_1605_U116 , SUB_1605_U117 , SUB_1605_U118 , SUB_1605_U119 , SUB_1605_U120 , SUB_1605_U121 , SUB_1605_U122;
wire SUB_1605_U123 , SUB_1605_U124 , SUB_1605_U125 , SUB_1605_U126 , SUB_1605_U127 , SUB_1605_U128 , SUB_1605_U129 , SUB_1605_U130 , SUB_1605_U131 , SUB_1605_U132;
wire SUB_1605_U133 , SUB_1605_U134 , SUB_1605_U135 , SUB_1605_U136 , SUB_1605_U137 , SUB_1605_U138 , SUB_1605_U139 , SUB_1605_U140 , SUB_1605_U141 , SUB_1605_U142;
wire SUB_1605_U143 , SUB_1605_U144 , SUB_1605_U145 , SUB_1605_U146 , SUB_1605_U147 , SUB_1605_U148 , SUB_1605_U149 , SUB_1605_U150 , SUB_1605_U151 , SUB_1605_U152;
wire SUB_1605_U153 , SUB_1605_U154 , SUB_1605_U155 , SUB_1605_U156 , SUB_1605_U157 , SUB_1605_U158 , SUB_1605_U159 , SUB_1605_U160 , SUB_1605_U161 , SUB_1605_U162;
wire SUB_1605_U163 , SUB_1605_U164 , SUB_1605_U165 , SUB_1605_U166 , SUB_1605_U167 , SUB_1605_U168 , SUB_1605_U169 , SUB_1605_U170 , SUB_1605_U171 , SUB_1605_U172;
wire SUB_1605_U173 , SUB_1605_U174 , SUB_1605_U175 , SUB_1605_U176 , SUB_1605_U177 , SUB_1605_U178 , SUB_1605_U179 , SUB_1605_U180 , SUB_1605_U181 , SUB_1605_U182;
wire SUB_1605_U183 , SUB_1605_U184 , SUB_1605_U185 , SUB_1605_U186 , SUB_1605_U187 , SUB_1605_U188 , SUB_1605_U189 , SUB_1605_U190 , SUB_1605_U191 , SUB_1605_U192;
wire SUB_1605_U193 , SUB_1605_U194 , SUB_1605_U195 , SUB_1605_U196 , SUB_1605_U197 , SUB_1605_U198 , SUB_1605_U199 , SUB_1605_U200 , SUB_1605_U201 , SUB_1605_U202;
wire SUB_1605_U203 , SUB_1605_U204 , SUB_1605_U205 , SUB_1605_U206 , SUB_1605_U207 , SUB_1605_U208 , SUB_1605_U209 , SUB_1605_U210 , SUB_1605_U211 , SUB_1605_U212;
wire SUB_1605_U213 , SUB_1605_U214 , SUB_1605_U215 , SUB_1605_U216 , SUB_1605_U217 , SUB_1605_U218 , SUB_1605_U219 , SUB_1605_U220 , SUB_1605_U221 , SUB_1605_U222;
wire SUB_1605_U223 , SUB_1605_U224 , SUB_1605_U225 , SUB_1605_U226 , SUB_1605_U227 , SUB_1605_U228 , SUB_1605_U229 , SUB_1605_U230 , SUB_1605_U231 , SUB_1605_U232;
wire SUB_1605_U233 , SUB_1605_U234 , SUB_1605_U235 , SUB_1605_U236 , SUB_1605_U237 , SUB_1605_U238 , SUB_1605_U239 , SUB_1605_U240 , SUB_1605_U241 , SUB_1605_U242;
wire SUB_1605_U243 , SUB_1605_U244 , SUB_1605_U245 , SUB_1605_U246 , SUB_1605_U247 , SUB_1605_U248 , SUB_1605_U249 , SUB_1605_U250 , SUB_1605_U251 , SUB_1605_U252;
wire SUB_1605_U253 , SUB_1605_U254 , SUB_1605_U255 , SUB_1605_U256 , SUB_1605_U257 , SUB_1605_U258 , SUB_1605_U259 , SUB_1605_U260 , SUB_1605_U261 , SUB_1605_U262;
wire SUB_1605_U263 , SUB_1605_U264 , SUB_1605_U265 , SUB_1605_U266 , SUB_1605_U267 , SUB_1605_U268 , SUB_1605_U269 , SUB_1605_U270 , SUB_1605_U271 , SUB_1605_U272;
wire SUB_1605_U273 , SUB_1605_U274 , SUB_1605_U275 , SUB_1605_U276 , SUB_1605_U277 , SUB_1605_U278 , SUB_1605_U279 , SUB_1605_U280 , SUB_1605_U281 , SUB_1605_U282;
wire SUB_1605_U283 , SUB_1605_U284 , SUB_1605_U285 , SUB_1605_U286 , SUB_1605_U287 , SUB_1605_U288 , SUB_1605_U289 , SUB_1605_U290 , SUB_1605_U291 , SUB_1605_U292;
wire SUB_1605_U293 , SUB_1605_U294 , SUB_1605_U295 , SUB_1605_U296 , SUB_1605_U297 , SUB_1605_U298 , SUB_1605_U299 , SUB_1605_U300 , SUB_1605_U301 , SUB_1605_U302;
wire SUB_1605_U303 , SUB_1605_U304 , SUB_1605_U305 , SUB_1605_U306 , SUB_1605_U307 , SUB_1605_U308 , SUB_1605_U309 , SUB_1605_U310 , SUB_1605_U311 , SUB_1605_U312;
wire SUB_1605_U313 , SUB_1605_U314 , SUB_1605_U315 , SUB_1605_U316 , SUB_1605_U317 , SUB_1605_U318 , SUB_1605_U319 , SUB_1605_U320 , SUB_1605_U321 , SUB_1605_U322;
wire SUB_1605_U323 , SUB_1605_U324 , SUB_1605_U325 , SUB_1605_U326 , SUB_1605_U327 , SUB_1605_U328 , SUB_1605_U329 , SUB_1605_U330 , SUB_1605_U331 , SUB_1605_U332;
wire SUB_1605_U333 , SUB_1605_U334 , SUB_1605_U335 , SUB_1605_U336 , SUB_1605_U337 , SUB_1605_U338 , SUB_1605_U339 , SUB_1605_U340 , SUB_1605_U341 , SUB_1605_U342;
wire SUB_1605_U343 , SUB_1605_U344 , SUB_1605_U345 , SUB_1605_U346 , SUB_1605_U347 , SUB_1605_U348 , SUB_1605_U349 , SUB_1605_U350 , SUB_1605_U351 , SUB_1605_U352;
wire SUB_1605_U353 , SUB_1605_U354 , SUB_1605_U355 , SUB_1605_U356 , SUB_1605_U357 , SUB_1605_U358 , SUB_1605_U359 , SUB_1605_U360 , SUB_1605_U361 , SUB_1605_U362;
wire SUB_1605_U363 , SUB_1605_U364 , SUB_1605_U365 , SUB_1605_U366 , SUB_1605_U367 , SUB_1605_U368 , SUB_1605_U369 , SUB_1605_U370 , SUB_1605_U371 , SUB_1605_U372;
wire SUB_1605_U373 , SUB_1605_U374 , SUB_1605_U375 , SUB_1605_U376 , SUB_1605_U377 , SUB_1605_U378 , SUB_1605_U379 , SUB_1605_U380 , SUB_1605_U381 , SUB_1605_U382;
wire SUB_1605_U383 , SUB_1605_U384 , SUB_1605_U385 , SUB_1605_U386 , SUB_1605_U387 , SUB_1605_U388 , SUB_1605_U389 , SUB_1605_U390 , SUB_1605_U391 , SUB_1605_U392;
wire SUB_1605_U393 , SUB_1605_U394 , SUB_1605_U395 , SUB_1605_U396 , SUB_1605_U397 , SUB_1605_U398 , SUB_1605_U399 , SUB_1605_U400 , SUB_1605_U401 , SUB_1605_U402;
wire SUB_1605_U403 , SUB_1605_U404 , SUB_1605_U405 , SUB_1605_U406 , SUB_1605_U407 , SUB_1605_U408 , SUB_1605_U409 , SUB_1605_U410 , SUB_1605_U411 , SUB_1605_U412;
wire SUB_1605_U413 , SUB_1605_U414 , SUB_1605_U415 , SUB_1605_U416 , SUB_1605_U417 , SUB_1605_U418 , SUB_1605_U419 , SUB_1605_U420 , SUB_1605_U421 , SUB_1605_U422;
wire SUB_1605_U423 , SUB_1605_U424 , SUB_1605_U425 , SUB_1605_U426 , SUB_1605_U427 , SUB_1605_U428 , SUB_1605_U429 , SUB_1605_U430 , SUB_1605_U431 , SUB_1605_U432;
wire SUB_1605_U433 , SUB_1605_U434 , SUB_1605_U435 , SUB_1605_U436 , SUB_1605_U437 , SUB_1605_U438 , SUB_1605_U439 , SUB_1605_U440 , SUB_1605_U441 , SUB_1605_U442;
wire SUB_1605_U443 , SUB_1605_U444 , SUB_1605_U445 , SUB_1605_U446 , SUB_1605_U447 , SUB_1605_U448 , SUB_1605_U449 , SUB_1605_U450 , SUB_1605_U451 , SUB_1605_U452;
wire SUB_1605_U453 , SUB_1605_U454 , SUB_1605_U455 , SUB_1605_U456 , SUB_1605_U457 , SUB_1605_U458 , SUB_1605_U459 , SUB_1605_U460 , SUB_1605_U461 , SUB_1605_U462;
wire SUB_1605_U463 , SUB_1605_U464 , SUB_1605_U465 , SUB_1605_U466 , SUB_1605_U467 , SUB_1605_U468 , SUB_1605_U469 , SUB_1605_U470 , SUB_1605_U471 , SUB_1605_U472;
wire SUB_1605_U473 , SUB_1605_U474 , SUB_1605_U475 , SUB_1605_U476 , SUB_1605_U477 , SUB_1605_U478 , SUB_1605_U479 , SUB_1605_U480 , R152_U4 , R152_U5;
wire R152_U6 , R152_U7 , R152_U8 , R152_U9 , R152_U10 , R152_U11 , R152_U12 , R152_U13 , R152_U14 , R152_U15;
wire R152_U16 , R152_U17 , R152_U18 , R152_U19 , R152_U20 , R152_U21 , R152_U22 , R152_U23 , R152_U24 , R152_U25;
wire R152_U26 , R152_U27 , R152_U28 , R152_U29 , R152_U30 , R152_U31 , R152_U32 , R152_U33 , R152_U34 , R152_U35;
wire R152_U36 , R152_U37 , R152_U38 , R152_U39 , R152_U40 , R152_U41 , R152_U42 , R152_U43 , R152_U44 , R152_U45;
wire R152_U46 , R152_U47 , R152_U48 , R152_U49 , R152_U50 , R152_U51 , R152_U52 , R152_U53 , R152_U54 , R152_U55;
wire R152_U56 , R152_U57 , R152_U58 , R152_U59 , R152_U60 , R152_U61 , R152_U62 , R152_U63 , R152_U64 , R152_U65;
wire R152_U66 , R152_U67 , R152_U68 , R152_U69 , R152_U70 , R152_U71 , R152_U72 , R152_U73 , R152_U74 , R152_U75;
wire R152_U76 , R152_U77 , R152_U78 , R152_U79 , R152_U80 , R152_U81 , R152_U82 , R152_U83 , R152_U84 , R152_U85;
wire R152_U86 , R152_U87 , R152_U88 , R152_U89 , R152_U90 , R152_U91 , R152_U92 , R152_U93 , R152_U94 , R152_U95;
wire R152_U96 , R152_U97 , R152_U98 , R152_U99 , R152_U100 , R152_U101 , R152_U102 , R152_U103 , R152_U104 , R152_U105;
wire R152_U106 , R152_U107 , R152_U108 , R152_U109 , R152_U110 , R152_U111 , R152_U112 , R152_U113 , R152_U114 , R152_U115;
wire R152_U116 , R152_U117 , R152_U118 , R152_U119 , R152_U120 , R152_U121 , R152_U122 , R152_U123 , R152_U124 , R152_U125;
wire R152_U126 , R152_U127 , R152_U128 , R152_U129 , R152_U130 , R152_U131 , R152_U132 , R152_U133 , R152_U134 , R152_U135;
wire R152_U136 , R152_U137 , R152_U138 , R152_U139 , R152_U140 , R152_U141 , R152_U142 , R152_U143 , R152_U144 , R152_U145;
wire R152_U146 , R152_U147 , R152_U148 , R152_U149 , R152_U150 , R152_U151 , R152_U152 , R152_U153 , R152_U154 , R152_U155;
wire R152_U156 , R152_U157 , R152_U158 , R152_U159 , R152_U160 , R152_U161 , R152_U162 , R152_U163 , R152_U164 , R152_U165;
wire R152_U166 , R152_U167 , R152_U168 , R152_U169 , R152_U170 , R152_U171 , R152_U172 , R152_U173 , R152_U174 , R152_U175;
wire R152_U176 , R152_U177 , R152_U178 , R152_U179 , R152_U180 , R152_U181 , R152_U182 , R152_U183 , R152_U184 , R152_U185;
wire R152_U186 , R152_U187 , R152_U188 , R152_U189 , R152_U190 , R152_U191 , R152_U192 , R152_U193 , R152_U194 , R152_U195;
wire R152_U196 , R152_U197 , R152_U198 , R152_U199 , R152_U200 , R152_U201 , R152_U202 , R152_U203 , R152_U204 , R152_U205;
wire R152_U206 , R152_U207 , R152_U208 , R152_U209 , R152_U210 , R152_U211 , R152_U212 , R152_U213 , R152_U214 , R152_U215;
wire R152_U216 , R152_U217 , R152_U218 , R152_U219 , R152_U220 , R152_U221 , R152_U222 , R152_U223 , R152_U224 , R152_U225;
wire R152_U226 , R152_U227 , R152_U228 , R152_U229 , R152_U230 , R152_U231 , R152_U232 , R152_U233 , R152_U234 , R152_U235;
wire R152_U236 , R152_U237 , R152_U238 , R152_U239 , R152_U240 , R152_U241 , R152_U242 , R152_U243 , R152_U244 , R152_U245;
wire R152_U246 , R152_U247 , R152_U248 , R152_U249 , R152_U250 , R152_U251 , R152_U252 , R152_U253 , R152_U254 , R152_U255;
wire R152_U256 , R152_U257 , R152_U258 , R152_U259 , R152_U260 , R152_U261 , R152_U262 , R152_U263 , R152_U264 , R152_U265;
wire R152_U266 , R152_U267 , R152_U268 , R152_U269 , R152_U270 , R152_U271 , R152_U272 , R152_U273 , R152_U274 , R152_U275;
wire R152_U276 , R152_U277 , R152_U278 , R152_U279 , R152_U280 , R152_U281 , R152_U282 , R152_U283 , R152_U284 , R152_U285;
wire R152_U286 , R152_U287 , R152_U288 , R152_U289 , R152_U290 , R152_U291 , R152_U292 , R152_U293 , R152_U294 , R152_U295;
wire R152_U296 , R152_U297 , R152_U298 , R152_U299 , R152_U300 , R152_U301 , R152_U302 , R152_U303 , R152_U304 , R152_U305;
wire R152_U306 , R152_U307 , R152_U308 , R152_U309 , R152_U310 , R152_U311 , R152_U312 , R152_U313 , R152_U314 , R152_U315;
wire R152_U316 , R152_U317 , R152_U318 , R152_U319 , R152_U320 , R152_U321 , R152_U322 , R152_U323 , R152_U324 , R152_U325;
wire R152_U326 , R152_U327 , R152_U328 , R152_U329 , R152_U330 , R152_U331 , R152_U332 , R152_U333 , R152_U334 , R152_U335;
wire R152_U336 , R152_U337 , R152_U338 , R152_U339 , R152_U340 , R152_U341 , R152_U342 , R152_U343 , R152_U344 , R152_U345;
wire R152_U346 , R152_U347 , R152_U348 , R152_U349 , R152_U350 , R152_U351 , R152_U352 , R152_U353 , R152_U354 , R152_U355;
wire R152_U356 , R152_U357 , R152_U358 , R152_U359 , R152_U360 , R152_U361 , R152_U362 , R152_U363 , R152_U364 , R152_U365;
wire R152_U366 , R152_U367 , R152_U368 , R152_U369 , R152_U370 , R152_U371 , R152_U372 , R152_U373 , R152_U374 , R152_U375;
wire R152_U376 , R152_U377 , R152_U378 , R152_U379 , R152_U380 , R152_U381 , R152_U382 , R152_U383 , R152_U384 , R152_U385;
wire R152_U386 , R152_U387 , R152_U388 , R152_U389 , R152_U390 , R152_U391 , R152_U392 , R152_U393 , R152_U394 , R152_U395;
wire R152_U396 , R152_U397 , R152_U398 , R152_U399 , R152_U400 , R152_U401 , R152_U402 , R152_U403 , R152_U404 , R152_U405;
wire R152_U406 , R152_U407 , R152_U408 , R152_U409 , R152_U410 , R152_U411 , R152_U412 , R152_U413 , R152_U414 , R152_U415;
wire R152_U416 , R152_U417 , R152_U418 , R152_U419 , R152_U420 , R152_U421 , R152_U422 , R152_U423 , R152_U424 , R152_U425;
wire R152_U426 , R152_U427 , R152_U428 , R152_U429 , R152_U430 , R152_U431 , R152_U432 , R152_U433 , R152_U434 , R152_U435;
wire R152_U436 , R152_U437 , R152_U438 , R152_U439 , R152_U440 , R152_U441 , R152_U442 , R152_U443 , R152_U444 , R152_U445;
wire R152_U446 , R152_U447 , R152_U448 , R152_U449 , R152_U450 , R152_U451 , R152_U452 , R152_U453 , R152_U454 , R152_U455;
wire R152_U456 , R152_U457 , R152_U458 , R152_U459 , R152_U460 , R152_U461 , R152_U462 , R152_U463 , R152_U464 , R152_U465;
wire R152_U466 , R152_U467 , R152_U468 , R152_U469 , R152_U470 , R152_U471 , R152_U472 , R152_U473 , R152_U474 , R152_U475;
wire R152_U476 , R152_U477 , R152_U478 , R152_U479 , R152_U480 , R152_U481 , R152_U482 , R152_U483 , R152_U484 , R152_U485;
wire R152_U486 , R152_U487 , R152_U488 , R152_U489 , R152_U490 , R152_U491 , R152_U492 , R152_U493 , R152_U494 , R152_U495;
wire R152_U496 , R152_U497 , R152_U498 , R152_U499 , R152_U500 , R152_U501 , R152_U502 , R152_U503 , R152_U504 , R152_U505;
wire R152_U506 , R152_U507 , R152_U508 , R152_U509 , R152_U510 , R152_U511 , R152_U512 , R152_U513 , R152_U514 , R152_U515;
wire R152_U516 , R152_U517 , R152_U518 , R152_U519 , R152_U520 , R152_U521 , R152_U522 , R152_U523 , R152_U524 , R152_U525;
wire R152_U526 , R152_U527 , R152_U528 , R152_U529 , R152_U530 , R152_U531 , R152_U532 , R152_U533 , R152_U534 , R152_U535;
wire R152_U536 , R152_U537 , R152_U538 , R152_U539 , R152_U540 , R152_U541 , R152_U542 , R152_U543 , R152_U544 , R152_U545;
wire R152_U546 , R152_U547 , R152_U548 , R152_U549 , R152_U550 , R152_U551 , R152_U552 , R152_U553 , R152_U554 , LT_1602_U6;
wire LT_1601_U6 , SUB_1596_U6 , SUB_1596_U7 , SUB_1596_U8 , SUB_1596_U9 , SUB_1596_U10 , SUB_1596_U11 , SUB_1596_U12 , SUB_1596_U13 , SUB_1596_U14;
wire SUB_1596_U15 , SUB_1596_U16 , SUB_1596_U17 , SUB_1596_U18 , SUB_1596_U19 , SUB_1596_U20 , SUB_1596_U21 , SUB_1596_U22 , SUB_1596_U23 , SUB_1596_U24;
wire SUB_1596_U25 , SUB_1596_U26 , SUB_1596_U27 , SUB_1596_U28 , SUB_1596_U29 , SUB_1596_U30 , SUB_1596_U31 , SUB_1596_U32 , SUB_1596_U33 , SUB_1596_U34;
wire SUB_1596_U35 , SUB_1596_U36 , SUB_1596_U37 , SUB_1596_U38 , SUB_1596_U39 , SUB_1596_U40 , SUB_1596_U41 , SUB_1596_U42 , SUB_1596_U43 , SUB_1596_U44;
wire SUB_1596_U45 , SUB_1596_U46 , SUB_1596_U47 , SUB_1596_U48 , SUB_1596_U49 , SUB_1596_U50 , SUB_1596_U51 , SUB_1596_U52 , SUB_1596_U71 , SUB_1596_U72;
wire SUB_1596_U73 , SUB_1596_U74 , SUB_1596_U75 , SUB_1596_U76 , SUB_1596_U77 , SUB_1596_U78 , SUB_1596_U79 , SUB_1596_U80 , SUB_1596_U81 , SUB_1596_U82;
wire SUB_1596_U83 , SUB_1596_U84 , SUB_1596_U85 , SUB_1596_U86 , SUB_1596_U87 , SUB_1596_U88 , SUB_1596_U89 , SUB_1596_U90 , SUB_1596_U91 , SUB_1596_U92;
wire SUB_1596_U93 , SUB_1596_U94 , SUB_1596_U95 , SUB_1596_U96 , SUB_1596_U97 , SUB_1596_U98 , SUB_1596_U99 , SUB_1596_U100 , SUB_1596_U101 , SUB_1596_U102;
wire SUB_1596_U103 , SUB_1596_U104 , SUB_1596_U105 , SUB_1596_U106 , SUB_1596_U107 , SUB_1596_U108 , SUB_1596_U109 , SUB_1596_U110 , SUB_1596_U111 , SUB_1596_U112;
wire SUB_1596_U113 , SUB_1596_U114 , SUB_1596_U115 , SUB_1596_U116 , SUB_1596_U117 , SUB_1596_U118 , SUB_1596_U119 , SUB_1596_U120 , SUB_1596_U121 , SUB_1596_U122;
wire SUB_1596_U123 , SUB_1596_U124 , SUB_1596_U125 , SUB_1596_U126 , SUB_1596_U127 , SUB_1596_U128 , SUB_1596_U129 , SUB_1596_U130 , SUB_1596_U131 , SUB_1596_U132;
wire SUB_1596_U133 , SUB_1596_U134 , SUB_1596_U135 , SUB_1596_U136 , SUB_1596_U137 , SUB_1596_U138 , SUB_1596_U139 , SUB_1596_U140 , SUB_1596_U141 , SUB_1596_U142;
wire SUB_1596_U143 , SUB_1596_U144 , SUB_1596_U145 , SUB_1596_U146 , SUB_1596_U147 , SUB_1596_U148 , SUB_1596_U149 , SUB_1596_U150 , SUB_1596_U151 , SUB_1596_U152;
wire SUB_1596_U153 , SUB_1596_U154 , SUB_1596_U155 , SUB_1596_U156 , SUB_1596_U157 , SUB_1596_U158 , SUB_1596_U159 , SUB_1596_U160 , SUB_1596_U161 , SUB_1596_U162;
wire SUB_1596_U163 , SUB_1596_U164 , SUB_1596_U165 , SUB_1596_U166 , SUB_1596_U167 , SUB_1596_U168 , SUB_1596_U169 , SUB_1596_U170 , SUB_1596_U171 , SUB_1596_U172;
wire SUB_1596_U173 , SUB_1596_U174 , SUB_1596_U175 , SUB_1596_U176 , SUB_1596_U177 , SUB_1596_U178 , SUB_1596_U179 , SUB_1596_U180 , SUB_1596_U181 , SUB_1596_U182;
wire SUB_1596_U183 , SUB_1596_U184 , SUB_1596_U185 , SUB_1596_U186 , SUB_1596_U187 , SUB_1596_U188 , SUB_1596_U189 , SUB_1596_U190 , SUB_1596_U191 , SUB_1596_U192;
wire SUB_1596_U193 , SUB_1596_U194 , SUB_1596_U195 , SUB_1596_U196 , SUB_1596_U197 , SUB_1596_U198 , SUB_1596_U199 , SUB_1596_U200 , SUB_1596_U201 , SUB_1596_U202;
wire SUB_1596_U203 , SUB_1596_U204 , SUB_1596_U205 , SUB_1596_U206 , SUB_1596_U207 , SUB_1596_U208 , SUB_1596_U209 , SUB_1596_U210 , SUB_1596_U211 , SUB_1596_U212;
wire SUB_1596_U213 , SUB_1596_U214 , SUB_1596_U215 , SUB_1596_U216 , SUB_1596_U217 , SUB_1596_U218 , SUB_1596_U219 , SUB_1596_U220 , SUB_1596_U221 , SUB_1596_U222;
wire SUB_1596_U223 , SUB_1596_U224 , SUB_1596_U225 , SUB_1596_U226 , SUB_1596_U227 , SUB_1596_U228 , SUB_1596_U229 , SUB_1596_U230 , SUB_1596_U231 , SUB_1596_U232;
wire SUB_1596_U233 , SUB_1596_U234 , SUB_1596_U235 , SUB_1596_U236 , SUB_1596_U237 , SUB_1596_U238 , SUB_1596_U239 , SUB_1596_U240 , SUB_1596_U241 , SUB_1596_U242;
wire SUB_1596_U243 , SUB_1596_U244 , SUB_1596_U245 , SUB_1596_U246 , SUB_1596_U247 , SUB_1596_U248 , SUB_1596_U249 , SUB_1596_U250 , SUB_1596_U251 , SUB_1596_U252;
wire SUB_1596_U253 , SUB_1596_U254 , SUB_1596_U255 , SUB_1596_U256 , SUB_1596_U257 , SUB_1596_U258 , SUB_1596_U259 , SUB_1596_U260 , SUB_1596_U261 , SUB_1596_U262;
wire SUB_1596_U263 , SUB_1596_U264 , SUB_1596_U265 , SUB_1596_U266 , SUB_1596_U267 , SUB_1596_U268 , SUB_1596_U269 , SUB_1596_U270 , SUB_1596_U271 , SUB_1596_U272;
wire SUB_1596_U273 , SUB_1596_U274 , SUB_1596_U275 , SUB_1596_U276 , SUB_1596_U277 , SUB_1596_U278 , SUB_1596_U279 , SUB_1596_U280 , SUB_1596_U281 , SUB_1596_U282;
wire SUB_1596_U283 , SUB_1596_U284 , SUB_1596_U285 , SUB_1596_U286 , SUB_1596_U287 , SUB_1596_U288 , SUB_1596_U289 , SUB_1596_U290 , SUB_1596_U291 , ADD_1596_U6;
wire ADD_1596_U7 , ADD_1596_U8 , ADD_1596_U9 , ADD_1596_U10 , ADD_1596_U11 , ADD_1596_U12 , ADD_1596_U13 , ADD_1596_U14 , ADD_1596_U15 , ADD_1596_U16;
wire ADD_1596_U17 , ADD_1596_U18 , ADD_1596_U19 , ADD_1596_U20 , ADD_1596_U21 , ADD_1596_U22 , ADD_1596_U23 , ADD_1596_U24 , ADD_1596_U25 , ADD_1596_U26;
wire ADD_1596_U27 , ADD_1596_U28 , ADD_1596_U29 , ADD_1596_U30 , ADD_1596_U31 , ADD_1596_U32 , ADD_1596_U33 , ADD_1596_U34 , ADD_1596_U35 , ADD_1596_U36;
wire ADD_1596_U37 , ADD_1596_U38 , ADD_1596_U39 , ADD_1596_U40 , ADD_1596_U41 , ADD_1596_U42 , ADD_1596_U43 , ADD_1596_U44 , ADD_1596_U45 , ADD_1596_U46;
wire ADD_1596_U47 , ADD_1596_U48 , ADD_1596_U49 , ADD_1596_U50 , ADD_1596_U51 , ADD_1596_U52 , ADD_1596_U53 , ADD_1596_U54 , ADD_1596_U55 , ADD_1596_U56;
wire ADD_1596_U57 , ADD_1596_U58 , ADD_1596_U59 , ADD_1596_U60 , ADD_1596_U61 , ADD_1596_U62 , ADD_1596_U63 , ADD_1596_U64 , ADD_1596_U65 , ADD_1596_U66;
wire ADD_1596_U67 , ADD_1596_U68 , ADD_1596_U69 , ADD_1596_U70 , ADD_1596_U71 , ADD_1596_U72 , ADD_1596_U73 , ADD_1596_U74 , ADD_1596_U75 , ADD_1596_U76;
wire ADD_1596_U77 , ADD_1596_U78 , ADD_1596_U79 , ADD_1596_U80 , ADD_1596_U81 , ADD_1596_U82 , ADD_1596_U83 , ADD_1596_U84 , ADD_1596_U85 , ADD_1596_U86;
wire ADD_1596_U87 , ADD_1596_U88 , ADD_1596_U89 , ADD_1596_U90 , ADD_1596_U91 , ADD_1596_U92 , ADD_1596_U93 , ADD_1596_U94 , ADD_1596_U95 , ADD_1596_U96;
wire ADD_1596_U97 , ADD_1596_U98 , ADD_1596_U99 , ADD_1596_U100 , ADD_1596_U101 , ADD_1596_U102 , ADD_1596_U103 , ADD_1596_U104 , ADD_1596_U105 , ADD_1596_U106;
wire ADD_1596_U107 , ADD_1596_U108 , ADD_1596_U109 , ADD_1596_U110 , ADD_1596_U111 , ADD_1596_U112 , ADD_1596_U113 , ADD_1596_U114 , ADD_1596_U115 , ADD_1596_U116;
wire ADD_1596_U117 , ADD_1596_U118 , ADD_1596_U119 , ADD_1596_U120 , ADD_1596_U121 , ADD_1596_U122 , ADD_1596_U123 , ADD_1596_U124 , ADD_1596_U125 , ADD_1596_U126;
wire ADD_1596_U127 , ADD_1596_U128 , ADD_1596_U129 , ADD_1596_U130 , ADD_1596_U131 , ADD_1596_U132 , ADD_1596_U133 , ADD_1596_U134 , ADD_1596_U135 , ADD_1596_U136;
wire ADD_1596_U137 , ADD_1596_U138 , ADD_1596_U139 , ADD_1596_U140 , ADD_1596_U141 , ADD_1596_U142 , ADD_1596_U143 , ADD_1596_U144 , ADD_1596_U145 , ADD_1596_U146;
wire ADD_1596_U147 , ADD_1596_U148 , ADD_1596_U149 , ADD_1596_U150 , ADD_1596_U151 , ADD_1596_U152 , ADD_1596_U153 , ADD_1596_U154 , ADD_1596_U155 , ADD_1596_U156;
wire ADD_1596_U157 , ADD_1596_U158 , ADD_1596_U159 , ADD_1596_U160 , ADD_1596_U161 , ADD_1596_U162 , ADD_1596_U163 , ADD_1596_U164 , ADD_1596_U165 , ADD_1596_U166;
wire ADD_1596_U167 , ADD_1596_U168 , ADD_1596_U169 , ADD_1596_U170 , ADD_1596_U171 , ADD_1596_U172 , ADD_1596_U173 , ADD_1596_U174 , ADD_1596_U175 , ADD_1596_U176;
wire ADD_1596_U177 , ADD_1596_U178 , ADD_1596_U179 , ADD_1596_U180 , ADD_1596_U181 , ADD_1596_U182 , ADD_1596_U183 , ADD_1596_U184 , ADD_1596_U185 , ADD_1596_U186;
wire ADD_1596_U187 , ADD_1596_U188 , ADD_1596_U189 , ADD_1596_U190 , ADD_1596_U191 , ADD_1596_U192 , ADD_1596_U193 , ADD_1596_U194 , ADD_1596_U195 , ADD_1596_U196;
wire ADD_1596_U197 , ADD_1596_U198 , ADD_1596_U199 , ADD_1596_U200 , ADD_1596_U201 , ADD_1596_U202 , ADD_1596_U203 , ADD_1596_U204 , ADD_1596_U205 , ADD_1596_U206;
wire ADD_1596_U207 , ADD_1596_U208 , ADD_1596_U209 , ADD_1596_U210 , ADD_1596_U211 , ADD_1596_U212 , ADD_1596_U213 , ADD_1596_U214 , ADD_1596_U215 , ADD_1596_U216;
wire ADD_1596_U217 , ADD_1596_U218 , ADD_1596_U219 , ADD_1596_U220 , ADD_1596_U221 , ADD_1596_U222 , ADD_1596_U223 , ADD_1596_U224 , ADD_1596_U225 , ADD_1596_U226;
wire ADD_1596_U227 , ADD_1596_U228 , ADD_1596_U229 , ADD_1596_U230 , ADD_1596_U231 , ADD_1596_U232 , ADD_1596_U233 , ADD_1596_U234 , ADD_1596_U235 , ADD_1596_U236;
wire ADD_1596_U237 , ADD_1596_U238 , ADD_1596_U239 , ADD_1596_U240 , ADD_1596_U241 , ADD_1596_U242 , ADD_1596_U243 , ADD_1596_U244 , ADD_1596_U245 , ADD_1596_U246;
wire ADD_1596_U247 , ADD_1596_U248 , ADD_1596_U249 , ADD_1596_U250 , ADD_1596_U251 , ADD_1596_U252 , ADD_1596_U253 , ADD_1596_U254 , ADD_1596_U255 , ADD_1596_U256;
wire ADD_1596_U257 , ADD_1596_U258 , ADD_1596_U259 , ADD_1596_U260 , ADD_1596_U261 , ADD_1596_U262 , ADD_1596_U263 , ADD_1596_U264 , ADD_1596_U265 , ADD_1596_U266;
wire ADD_1596_U267 , ADD_1596_U268 , ADD_1596_U269 , ADD_1596_U270 , ADD_1596_U271 , ADD_1596_U272 , ADD_1596_U273 , ADD_1596_U274 , LT_1601_21_U6 , P1_ADD_99_U4;
wire P1_ADD_99_U5 , P1_ADD_99_U6 , P1_ADD_99_U7 , P1_ADD_99_U8 , P1_ADD_99_U9 , P1_ADD_99_U10 , P1_ADD_99_U11 , P1_ADD_99_U12 , P1_ADD_99_U13 , P1_ADD_99_U14;
wire P1_ADD_99_U15 , P1_ADD_99_U16 , P1_ADD_99_U17 , P1_ADD_99_U18 , P1_ADD_99_U19 , P1_ADD_99_U20 , P1_ADD_99_U21 , P1_ADD_99_U22 , P1_ADD_99_U23 , P1_ADD_99_U24;
wire P1_ADD_99_U25 , P1_ADD_99_U26 , P1_ADD_99_U27 , P1_ADD_99_U28 , P1_ADD_99_U29 , P1_ADD_99_U30 , P1_ADD_99_U31 , P1_ADD_99_U32 , P1_ADD_99_U33 , P1_ADD_99_U34;
wire P1_ADD_99_U35 , P1_ADD_99_U36 , P1_ADD_99_U37 , P1_ADD_99_U38 , P1_ADD_99_U39 , P1_ADD_99_U40 , P1_ADD_99_U41 , P1_ADD_99_U42 , P1_ADD_99_U43 , P1_ADD_99_U44;
wire P1_ADD_99_U45 , P1_ADD_99_U46 , P1_ADD_99_U47 , P1_ADD_99_U48 , P1_ADD_99_U49 , P1_ADD_99_U50 , P1_ADD_99_U51 , P1_ADD_99_U52 , P1_ADD_99_U53 , P1_ADD_99_U54;
wire P1_ADD_99_U55 , P1_ADD_99_U56 , P1_ADD_99_U57 , P1_ADD_99_U58 , P1_ADD_99_U59 , P1_ADD_99_U60 , P1_ADD_99_U61 , P1_ADD_99_U62 , P1_ADD_99_U63 , P1_ADD_99_U64;
wire P1_ADD_99_U65 , P1_ADD_99_U66 , P1_ADD_99_U67 , P1_ADD_99_U68 , P1_ADD_99_U69 , P1_ADD_99_U70 , P1_ADD_99_U71 , P1_ADD_99_U72 , P1_ADD_99_U73 , P1_ADD_99_U74;
wire P1_ADD_99_U75 , P1_ADD_99_U76 , P1_ADD_99_U77 , P1_ADD_99_U78 , P1_ADD_99_U79 , P1_ADD_99_U80 , P1_ADD_99_U81 , P1_ADD_99_U82 , P1_ADD_99_U83 , P1_ADD_99_U84;
wire P1_ADD_99_U85 , P1_ADD_99_U86 , P1_ADD_99_U87 , P1_ADD_99_U88 , P1_ADD_99_U89 , P1_ADD_99_U90 , P1_ADD_99_U91 , P1_ADD_99_U92 , P1_ADD_99_U93 , P1_ADD_99_U94;
wire P1_ADD_99_U95 , P1_ADD_99_U96 , P1_ADD_99_U97 , P1_ADD_99_U98 , P1_ADD_99_U99 , P1_ADD_99_U100 , P1_ADD_99_U101 , P1_ADD_99_U102 , P1_ADD_99_U103 , P1_ADD_99_U104;
wire P1_ADD_99_U105 , P1_ADD_99_U106 , P1_ADD_99_U107 , P1_ADD_99_U108 , P1_ADD_99_U109 , P1_ADD_99_U110 , P1_ADD_99_U111 , P1_ADD_99_U112 , P1_ADD_99_U113 , P1_ADD_99_U114;
wire P1_ADD_99_U115 , P1_ADD_99_U116 , P1_ADD_99_U117 , P1_ADD_99_U118 , P1_ADD_99_U119 , P1_ADD_99_U120 , P1_ADD_99_U121 , P1_ADD_99_U122 , P1_ADD_99_U123 , P1_ADD_99_U124;
wire P1_ADD_99_U125 , P1_ADD_99_U126 , P1_ADD_99_U127 , P1_ADD_99_U128 , P1_ADD_99_U129 , P1_ADD_99_U130 , P1_ADD_99_U131 , P1_ADD_99_U132 , P1_ADD_99_U133 , P1_ADD_99_U134;
wire P1_ADD_99_U135 , P1_ADD_99_U136 , P1_ADD_99_U137 , P1_ADD_99_U138 , P1_ADD_99_U139 , P1_ADD_99_U140 , P1_ADD_99_U141 , P1_ADD_99_U142 , P1_ADD_99_U143 , P1_ADD_99_U144;
wire P1_ADD_99_U145 , P1_ADD_99_U146 , P1_ADD_99_U147 , P1_ADD_99_U148 , P1_ADD_99_U149 , P1_ADD_99_U150 , P1_ADD_99_U151 , P1_ADD_99_U152 , P1_ADD_99_U153 , P1_R1105_U4;
wire P1_R1105_U5 , P1_R1105_U6 , P1_R1105_U7 , P1_R1105_U8 , P1_R1105_U9 , P1_R1105_U10 , P1_R1105_U11 , P1_R1105_U12 , P1_R1105_U13 , P1_R1105_U14;
wire P1_R1105_U15 , P1_R1105_U16 , P1_R1105_U17 , P1_R1105_U18 , P1_R1105_U19 , P1_R1105_U20 , P1_R1105_U21 , P1_R1105_U22 , P1_R1105_U23 , P1_R1105_U24;
wire P1_R1105_U25 , P1_R1105_U26 , P1_R1105_U27 , P1_R1105_U28 , P1_R1105_U29 , P1_R1105_U30 , P1_R1105_U31 , P1_R1105_U32 , P1_R1105_U33 , P1_R1105_U34;
wire P1_R1105_U35 , P1_R1105_U36 , P1_R1105_U37 , P1_R1105_U38 , P1_R1105_U39 , P1_R1105_U40 , P1_R1105_U41 , P1_R1105_U42 , P1_R1105_U43 , P1_R1105_U44;
wire P1_R1105_U45 , P1_R1105_U46 , P1_R1105_U47 , P1_R1105_U48 , P1_R1105_U49 , P1_R1105_U50 , P1_R1105_U51 , P1_R1105_U52 , P1_R1105_U53 , P1_R1105_U54;
wire P1_R1105_U55 , P1_R1105_U56 , P1_R1105_U57 , P1_R1105_U58 , P1_R1105_U59 , P1_R1105_U60 , P1_R1105_U61 , P1_R1105_U62 , P1_R1105_U63 , P1_R1105_U64;
wire P1_R1105_U65 , P1_R1105_U66 , P1_R1105_U67 , P1_R1105_U68 , P1_R1105_U69 , P1_R1105_U70 , P1_R1105_U71 , P1_R1105_U72 , P1_R1105_U73 , P1_R1105_U74;
wire P1_R1105_U75 , P1_R1105_U76 , P1_R1105_U77 , P1_R1105_U78 , P1_R1105_U79 , P1_R1105_U80 , P1_R1105_U81 , P1_R1105_U82 , P1_R1105_U83 , P1_R1105_U84;
wire P1_R1105_U85 , P1_R1105_U86 , P1_R1105_U87 , P1_R1105_U88 , P1_R1105_U89 , P1_R1105_U90 , P1_R1105_U91 , P1_R1105_U92 , P1_R1105_U93 , P1_R1105_U94;
wire P1_R1105_U95 , P1_R1105_U96 , P1_R1105_U97 , P1_R1105_U98 , P1_R1105_U99 , P1_R1105_U100 , P1_R1105_U101 , P1_R1105_U102 , P1_R1105_U103 , P1_R1105_U104;
wire P1_R1105_U105 , P1_R1105_U106 , P1_R1105_U107 , P1_R1105_U108 , P1_R1105_U109 , P1_R1105_U110 , P1_R1105_U111 , P1_R1105_U112 , P1_R1105_U113 , P1_R1105_U114;
wire P1_R1105_U115 , P1_R1105_U116 , P1_R1105_U117 , P1_R1105_U118 , P1_R1105_U119 , P1_R1105_U120 , P1_R1105_U121 , P1_R1105_U122 , P1_R1105_U123 , P1_R1105_U124;
wire P1_R1105_U125 , P1_R1105_U126 , P1_R1105_U127 , P1_R1105_U128 , P1_R1105_U129 , P1_R1105_U130 , P1_R1105_U131 , P1_R1105_U132 , P1_R1105_U133 , P1_R1105_U134;
wire P1_R1105_U135 , P1_R1105_U136 , P1_R1105_U137 , P1_R1105_U138 , P1_R1105_U139 , P1_R1105_U140 , P1_R1105_U141 , P1_R1105_U142 , P1_R1105_U143 , P1_R1105_U144;
wire P1_R1105_U145 , P1_R1105_U146 , P1_R1105_U147 , P1_R1105_U148 , P1_R1105_U149 , P1_R1105_U150 , P1_R1105_U151 , P1_R1105_U152 , P1_R1105_U153 , P1_R1105_U154;
wire P1_R1105_U155 , P1_R1105_U156 , P1_R1105_U157 , P1_R1105_U158 , P1_R1105_U159 , P1_R1105_U160 , P1_R1105_U161 , P1_R1105_U162 , P1_R1105_U163 , P1_R1105_U164;
wire P1_R1105_U165 , P1_R1105_U166 , P1_R1105_U167 , P1_R1105_U168 , P1_R1105_U169 , P1_R1105_U170 , P1_R1105_U171 , P1_R1105_U172 , P1_R1105_U173 , P1_R1105_U174;
wire P1_R1105_U175 , P1_R1105_U176 , P1_R1105_U177 , P1_R1105_U178 , P1_R1105_U179 , P1_R1105_U180 , P1_R1105_U181 , P1_R1105_U182 , P1_R1105_U183 , P1_R1105_U184;
wire P1_R1105_U185 , P1_R1105_U186 , P1_R1105_U187 , P1_R1105_U188 , P1_R1105_U189 , P1_R1105_U190 , P1_R1105_U191 , P1_R1105_U192 , P1_R1105_U193 , P1_R1105_U194;
wire P1_R1105_U195 , P1_R1105_U196 , P1_R1105_U197 , P1_R1105_U198 , P1_R1105_U199 , P1_R1105_U200 , P1_R1105_U201 , P1_R1105_U202 , P1_R1105_U203 , P1_R1105_U204;
wire P1_R1105_U205 , P1_R1105_U206 , P1_R1105_U207 , P1_R1105_U208 , P1_R1105_U209 , P1_R1105_U210 , P1_R1105_U211 , P1_R1105_U212 , P1_R1105_U213 , P1_R1105_U214;
wire P1_R1105_U215 , P1_R1105_U216 , P1_R1105_U217 , P1_R1105_U218 , P1_R1105_U219 , P1_R1105_U220 , P1_R1105_U221 , P1_R1105_U222 , P1_R1105_U223 , P1_R1105_U224;
wire P1_R1105_U225 , P1_R1105_U226 , P1_R1105_U227 , P1_R1105_U228 , P1_R1105_U229 , P1_R1105_U230 , P1_R1105_U231 , P1_R1105_U232 , P1_R1105_U233 , P1_R1105_U234;
wire P1_R1105_U235 , P1_R1105_U236 , P1_R1105_U237 , P1_R1105_U238 , P1_R1105_U239 , P1_R1105_U240 , P1_R1105_U241 , P1_R1105_U242 , P1_R1105_U243 , P1_R1105_U244;
wire P1_R1105_U245 , P1_R1105_U246 , P1_R1105_U247 , P1_R1105_U248 , P1_R1105_U249 , P1_R1105_U250 , P1_R1105_U251 , P1_R1105_U252 , P1_R1105_U253 , P1_R1105_U254;
wire P1_R1105_U255 , P1_R1105_U256 , P1_R1105_U257 , P1_R1105_U258 , P1_R1105_U259 , P1_R1105_U260 , P1_R1105_U261 , P1_R1105_U262 , P1_R1105_U263 , P1_R1105_U264;
wire P1_R1105_U265 , P1_R1105_U266 , P1_R1105_U267 , P1_R1105_U268 , P1_R1105_U269 , P1_R1105_U270 , P1_R1105_U271 , P1_R1105_U272 , P1_R1105_U273 , P1_R1105_U274;
wire P1_R1105_U275 , P1_R1105_U276 , P1_R1105_U277 , P1_R1105_U278 , P1_R1105_U279 , P1_R1105_U280 , P1_R1105_U281 , P1_R1105_U282 , P1_R1105_U283 , P1_R1105_U284;
wire P1_R1105_U285 , P1_R1105_U286 , P1_R1105_U287 , P1_R1105_U288 , P1_R1105_U289 , P1_R1105_U290 , P1_R1105_U291 , P1_R1105_U292 , P1_R1105_U293 , P1_R1105_U294;
wire P1_R1105_U295 , P1_R1105_U296 , P1_R1105_U297 , P1_R1105_U298 , P1_R1105_U299 , P1_R1105_U300 , P1_R1105_U301 , P1_R1105_U302 , P1_R1105_U303 , P1_R1105_U304;
wire P1_R1105_U305 , P1_R1105_U306 , P1_R1105_U307 , P1_R1105_U308 , P1_SUB_88_U6 , P1_SUB_88_U7 , P1_SUB_88_U8 , P1_SUB_88_U9 , P1_SUB_88_U10 , P1_SUB_88_U11;
wire P1_SUB_88_U12 , P1_SUB_88_U13 , P1_SUB_88_U14 , P1_SUB_88_U15 , P1_SUB_88_U16 , P1_SUB_88_U17 , P1_SUB_88_U18 , P1_SUB_88_U19 , P1_SUB_88_U20 , P1_SUB_88_U21;
wire P1_SUB_88_U22 , P1_SUB_88_U23 , P1_SUB_88_U24 , P1_SUB_88_U25 , P1_SUB_88_U26 , P1_SUB_88_U27 , P1_SUB_88_U28 , P1_SUB_88_U29 , P1_SUB_88_U30 , P1_SUB_88_U31;
wire P1_SUB_88_U32 , P1_SUB_88_U33 , P1_SUB_88_U34 , P1_SUB_88_U35 , P1_SUB_88_U36 , P1_SUB_88_U37 , P1_SUB_88_U38 , P1_SUB_88_U39 , P1_SUB_88_U40 , P1_SUB_88_U41;
wire P1_SUB_88_U42 , P1_SUB_88_U43 , P1_SUB_88_U44 , P1_SUB_88_U45 , P1_SUB_88_U46 , P1_SUB_88_U47 , P1_SUB_88_U48 , P1_SUB_88_U49 , P1_SUB_88_U50 , P1_SUB_88_U51;
wire P1_SUB_88_U52 , P1_SUB_88_U53 , P1_SUB_88_U54 , P1_SUB_88_U55 , P1_SUB_88_U56 , P1_SUB_88_U57 , P1_SUB_88_U58 , P1_SUB_88_U59 , P1_SUB_88_U60 , P1_SUB_88_U61;
wire P1_SUB_88_U62 , P1_SUB_88_U63 , P1_SUB_88_U64 , P1_SUB_88_U65 , P1_SUB_88_U66 , P1_SUB_88_U67 , P1_SUB_88_U68 , P1_SUB_88_U69 , P1_SUB_88_U70 , P1_SUB_88_U71;
wire P1_SUB_88_U72 , P1_SUB_88_U73 , P1_SUB_88_U74 , P1_SUB_88_U75 , P1_SUB_88_U76 , P1_SUB_88_U77 , P1_SUB_88_U78 , P1_SUB_88_U79 , P1_SUB_88_U80 , P1_SUB_88_U81;
wire P1_SUB_88_U82 , P1_SUB_88_U83 , P1_SUB_88_U84 , P1_SUB_88_U85 , P1_SUB_88_U86 , P1_SUB_88_U87 , P1_SUB_88_U88 , P1_SUB_88_U89 , P1_SUB_88_U90 , P1_SUB_88_U91;
wire P1_SUB_88_U92 , P1_SUB_88_U93 , P1_SUB_88_U94 , P1_SUB_88_U95 , P1_SUB_88_U96 , P1_SUB_88_U97 , P1_SUB_88_U98 , P1_SUB_88_U99 , P1_SUB_88_U100 , P1_SUB_88_U101;
wire P1_SUB_88_U102 , P1_SUB_88_U103 , P1_SUB_88_U104 , P1_SUB_88_U105 , P1_SUB_88_U106 , P1_SUB_88_U107 , P1_SUB_88_U108 , P1_SUB_88_U109 , P1_SUB_88_U110 , P1_SUB_88_U111;
wire P1_SUB_88_U112 , P1_SUB_88_U113 , P1_SUB_88_U114 , P1_SUB_88_U115 , P1_SUB_88_U116 , P1_SUB_88_U117 , P1_SUB_88_U118 , P1_SUB_88_U119 , P1_SUB_88_U120 , P1_SUB_88_U121;
wire P1_SUB_88_U122 , P1_SUB_88_U123 , P1_SUB_88_U124 , P1_SUB_88_U125 , P1_SUB_88_U126 , P1_SUB_88_U127 , P1_SUB_88_U128 , P1_SUB_88_U129 , P1_SUB_88_U130 , P1_SUB_88_U131;
wire P1_SUB_88_U132 , P1_SUB_88_U133 , P1_SUB_88_U134 , P1_SUB_88_U135 , P1_SUB_88_U136 , P1_SUB_88_U137 , P1_SUB_88_U138 , P1_SUB_88_U139 , P1_SUB_88_U140 , P1_SUB_88_U141;
wire P1_SUB_88_U142 , P1_SUB_88_U143 , P1_SUB_88_U144 , P1_SUB_88_U145 , P1_SUB_88_U146 , P1_SUB_88_U147 , P1_SUB_88_U148 , P1_SUB_88_U149 , P1_SUB_88_U150 , P1_SUB_88_U151;
wire P1_SUB_88_U152 , P1_SUB_88_U153 , P1_SUB_88_U154 , P1_SUB_88_U155 , P1_SUB_88_U156 , P1_SUB_88_U157 , P1_SUB_88_U158 , P1_SUB_88_U159 , P1_SUB_88_U160 , P1_SUB_88_U161;
wire P1_SUB_88_U162 , P1_SUB_88_U163 , P1_SUB_88_U164 , P1_SUB_88_U165 , P1_SUB_88_U166 , P1_SUB_88_U167 , P1_SUB_88_U168 , P1_SUB_88_U169 , P1_SUB_88_U170 , P1_SUB_88_U171;
wire P1_SUB_88_U172 , P1_SUB_88_U173 , P1_SUB_88_U174 , P1_SUB_88_U175 , P1_SUB_88_U176 , P1_SUB_88_U177 , P1_SUB_88_U178 , P1_SUB_88_U179 , P1_SUB_88_U180 , P1_SUB_88_U181;
wire P1_SUB_88_U182 , P1_SUB_88_U183 , P1_SUB_88_U184 , P1_SUB_88_U185 , P1_SUB_88_U186 , P1_SUB_88_U187 , P1_SUB_88_U188 , P1_SUB_88_U189 , P1_SUB_88_U190 , P1_SUB_88_U191;
wire P1_SUB_88_U192 , P1_SUB_88_U193 , P1_SUB_88_U194 , P1_SUB_88_U195 , P1_SUB_88_U196 , P1_SUB_88_U197 , P1_SUB_88_U198 , P1_SUB_88_U199 , P1_SUB_88_U200 , P1_SUB_88_U201;
wire P1_SUB_88_U202 , P1_SUB_88_U203 , P1_SUB_88_U204 , P1_SUB_88_U205 , P1_SUB_88_U206 , P1_SUB_88_U207 , P1_SUB_88_U208 , P1_SUB_88_U209 , P1_SUB_88_U210 , P1_SUB_88_U211;
wire P1_SUB_88_U212 , P1_SUB_88_U213 , P1_SUB_88_U214 , P1_SUB_88_U215 , P1_SUB_88_U216 , P1_SUB_88_U217 , P1_SUB_88_U218 , P1_SUB_88_U219 , P1_SUB_88_U220 , P1_SUB_88_U221;
wire P1_SUB_88_U222 , P1_SUB_88_U223 , P1_SUB_88_U224 , P1_SUB_88_U225 , P1_SUB_88_U226 , P1_SUB_88_U227 , P1_SUB_88_U228 , P1_SUB_88_U229 , P1_SUB_88_U230 , P1_SUB_88_U231;
wire P1_SUB_88_U232 , P1_SUB_88_U233 , P1_SUB_88_U234 , P1_SUB_88_U235 , P1_SUB_88_U236 , P1_SUB_88_U237 , P1_SUB_88_U238 , P1_SUB_88_U239 , P1_SUB_88_U240 , P1_SUB_88_U241;
wire P1_SUB_88_U242 , P1_SUB_88_U243 , P1_SUB_88_U244 , P1_SUB_88_U245 , P1_SUB_88_U246 , P1_SUB_88_U247 , P1_SUB_88_U248 , P1_SUB_88_U249 , P1_SUB_88_U250 , P1_SUB_88_U251;
wire P1_R1309_U6 , P1_R1309_U7 , P1_R1309_U8 , P1_R1309_U9 , P1_R1309_U10 , P1_R1282_U6 , P1_R1282_U7 , P1_R1282_U8 , P1_R1282_U9 , P1_R1282_U10;
wire P1_R1282_U11 , P1_R1282_U12 , P1_R1282_U13 , P1_R1282_U14 , P1_R1282_U15 , P1_R1282_U16 , P1_R1282_U17 , P1_R1282_U18 , P1_R1282_U19 , P1_R1282_U20;
wire P1_R1282_U21 , P1_R1282_U22 , P1_R1282_U23 , P1_R1282_U24 , P1_R1282_U25 , P1_R1282_U26 , P1_R1282_U27 , P1_R1282_U28 , P1_R1282_U29 , P1_R1282_U30;
wire P1_R1282_U31 , P1_R1282_U32 , P1_R1282_U33 , P1_R1282_U34 , P1_R1282_U35 , P1_R1282_U36 , P1_R1282_U37 , P1_R1282_U38 , P1_R1282_U39 , P1_R1282_U40;
wire P1_R1282_U41 , P1_R1282_U42 , P1_R1282_U43 , P1_R1282_U44 , P1_R1282_U45 , P1_R1282_U46 , P1_R1282_U47 , P1_R1282_U48 , P1_R1282_U49 , P1_R1282_U50;
wire P1_R1282_U51 , P1_R1282_U52 , P1_R1282_U53 , P1_R1282_U54 , P1_R1282_U55 , P1_R1282_U56 , P1_R1282_U57 , P1_R1282_U58 , P1_R1282_U59 , P1_R1282_U60;
wire P1_R1282_U61 , P1_R1282_U62 , P1_R1282_U63 , P1_R1282_U64 , P1_R1282_U65 , P1_R1282_U66 , P1_R1282_U67 , P1_R1282_U68 , P1_R1282_U69 , P1_R1282_U70;
wire P1_R1282_U71 , P1_R1282_U72 , P1_R1282_U73 , P1_R1282_U74 , P1_R1282_U75 , P1_R1282_U76 , P1_R1282_U77 , P1_R1282_U78 , P1_R1282_U79 , P1_R1282_U80;
wire P1_R1282_U81 , P1_R1282_U82 , P1_R1282_U83 , P1_R1282_U84 , P1_R1282_U85 , P1_R1282_U86 , P1_R1282_U87 , P1_R1282_U88 , P1_R1282_U89 , P1_R1282_U90;
wire P1_R1282_U91 , P1_R1282_U92 , P1_R1282_U93 , P1_R1282_U94 , P1_R1282_U95 , P1_R1282_U96 , P1_R1282_U97 , P1_R1282_U98 , P1_R1282_U99 , P1_R1282_U100;
wire P1_R1282_U101 , P1_R1282_U102 , P1_R1282_U103 , P1_R1282_U104 , P1_R1282_U105 , P1_R1282_U106 , P1_R1282_U107 , P1_R1282_U108 , P1_R1282_U109 , P1_R1282_U110;
wire P1_R1282_U111 , P1_R1282_U112 , P1_R1282_U113 , P1_R1282_U114 , P1_R1282_U115 , P1_R1282_U116 , P1_R1282_U117 , P1_R1282_U118 , P1_R1282_U119 , P1_R1282_U120;
wire P1_R1282_U121 , P1_R1282_U122 , P1_R1282_U123 , P1_R1282_U124 , P1_R1282_U125 , P1_R1282_U126 , P1_R1282_U127 , P1_R1282_U128 , P1_R1282_U129 , P1_R1282_U130;
wire P1_R1282_U131 , P1_R1282_U132 , P1_R1282_U133 , P1_R1282_U134 , P1_R1282_U135 , P1_R1282_U136 , P1_R1282_U137 , P1_R1282_U138 , P1_R1282_U139 , P1_R1282_U140;
wire P1_R1282_U141 , P1_R1282_U142 , P1_R1282_U143 , P1_R1282_U144 , P1_R1282_U145 , P1_R1282_U146 , P1_R1282_U147 , P1_R1282_U148 , P1_R1282_U149 , P1_R1282_U150;
wire P1_R1282_U151 , P1_R1282_U152 , P1_R1282_U153 , P1_R1282_U154 , P1_R1282_U155 , P1_R1282_U156 , P1_R1282_U157 , P1_R1282_U158 , P1_R1282_U159 , P1_R1240_U4;
wire P1_R1240_U5 , P1_R1240_U6 , P1_R1240_U7 , P1_R1240_U8 , P1_R1240_U9 , P1_R1240_U10 , P1_R1240_U11 , P1_R1240_U12 , P1_R1240_U13 , P1_R1240_U14;
wire P1_R1240_U15 , P1_R1240_U16 , P1_R1240_U17 , P1_R1240_U18 , P1_R1240_U19 , P1_R1240_U20 , P1_R1240_U21 , P1_R1240_U22 , P1_R1240_U23 , P1_R1240_U24;
wire P1_R1240_U25 , P1_R1240_U26 , P1_R1240_U27 , P1_R1240_U28 , P1_R1240_U29 , P1_R1240_U30 , P1_R1240_U31 , P1_R1240_U32 , P1_R1240_U33 , P1_R1240_U34;
wire P1_R1240_U35 , P1_R1240_U36 , P1_R1240_U37 , P1_R1240_U38 , P1_R1240_U39 , P1_R1240_U40 , P1_R1240_U41 , P1_R1240_U42 , P1_R1240_U43 , P1_R1240_U44;
wire P1_R1240_U45 , P1_R1240_U46 , P1_R1240_U47 , P1_R1240_U48 , P1_R1240_U49 , P1_R1240_U50 , P1_R1240_U51 , P1_R1240_U52 , P1_R1240_U53 , P1_R1240_U54;
wire P1_R1240_U55 , P1_R1240_U56 , P1_R1240_U57 , P1_R1240_U58 , P1_R1240_U59 , P1_R1240_U60 , P1_R1240_U61 , P1_R1240_U62 , P1_R1240_U63 , P1_R1240_U64;
wire P1_R1240_U65 , P1_R1240_U66 , P1_R1240_U67 , P1_R1240_U68 , P1_R1240_U69 , P1_R1240_U70 , P1_R1240_U71 , P1_R1240_U72 , P1_R1240_U73 , P1_R1240_U74;
wire P1_R1240_U75 , P1_R1240_U76 , P1_R1240_U77 , P1_R1240_U78 , P1_R1240_U79 , P1_R1240_U80 , P1_R1240_U81 , P1_R1240_U82 , P1_R1240_U83 , P1_R1240_U84;
wire P1_R1240_U85 , P1_R1240_U86 , P1_R1240_U87 , P1_R1240_U88 , P1_R1240_U89 , P1_R1240_U90 , P1_R1240_U91 , P1_R1240_U92 , P1_R1240_U93 , P1_R1240_U94;
wire P1_R1240_U95 , P1_R1240_U96 , P1_R1240_U97 , P1_R1240_U98 , P1_R1240_U99 , P1_R1240_U100 , P1_R1240_U101 , P1_R1240_U102 , P1_R1240_U103 , P1_R1240_U104;
wire P1_R1240_U105 , P1_R1240_U106 , P1_R1240_U107 , P1_R1240_U108 , P1_R1240_U109 , P1_R1240_U110 , P1_R1240_U111 , P1_R1240_U112 , P1_R1240_U113 , P1_R1240_U114;
wire P1_R1240_U115 , P1_R1240_U116 , P1_R1240_U117 , P1_R1240_U118 , P1_R1240_U119 , P1_R1240_U120 , P1_R1240_U121 , P1_R1240_U122 , P1_R1240_U123 , P1_R1240_U124;
wire P1_R1240_U125 , P1_R1240_U126 , P1_R1240_U127 , P1_R1240_U128 , P1_R1240_U129 , P1_R1240_U130 , P1_R1240_U131 , P1_R1240_U132 , P1_R1240_U133 , P1_R1240_U134;
wire P1_R1240_U135 , P1_R1240_U136 , P1_R1240_U137 , P1_R1240_U138 , P1_R1240_U139 , P1_R1240_U140 , P1_R1240_U141 , P1_R1240_U142 , P1_R1240_U143 , P1_R1240_U144;
wire P1_R1240_U145 , P1_R1240_U146 , P1_R1240_U147 , P1_R1240_U148 , P1_R1240_U149 , P1_R1240_U150 , P1_R1240_U151 , P1_R1240_U152 , P1_R1240_U153 , P1_R1240_U154;
wire P1_R1240_U155 , P1_R1240_U156 , P1_R1240_U157 , P1_R1240_U158 , P1_R1240_U159 , P1_R1240_U160 , P1_R1240_U161 , P1_R1240_U162 , P1_R1240_U163 , P1_R1240_U164;
wire P1_R1240_U165 , P1_R1240_U166 , P1_R1240_U167 , P1_R1240_U168 , P1_R1240_U169 , P1_R1240_U170 , P1_R1240_U171 , P1_R1240_U172 , P1_R1240_U173 , P1_R1240_U174;
wire P1_R1240_U175 , P1_R1240_U176 , P1_R1240_U177 , P1_R1240_U178 , P1_R1240_U179 , P1_R1240_U180 , P1_R1240_U181 , P1_R1240_U182 , P1_R1240_U183 , P1_R1240_U184;
wire P1_R1240_U185 , P1_R1240_U186 , P1_R1240_U187 , P1_R1240_U188 , P1_R1240_U189 , P1_R1240_U190 , P1_R1240_U191 , P1_R1240_U192 , P1_R1240_U193 , P1_R1240_U194;
wire P1_R1240_U195 , P1_R1240_U196 , P1_R1240_U197 , P1_R1240_U198 , P1_R1240_U199 , P1_R1240_U200 , P1_R1240_U201 , P1_R1240_U202 , P1_R1240_U203 , P1_R1240_U204;
wire P1_R1240_U205 , P1_R1240_U206 , P1_R1240_U207 , P1_R1240_U208 , P1_R1240_U209 , P1_R1240_U210 , P1_R1240_U211 , P1_R1240_U212 , P1_R1240_U213 , P1_R1240_U214;
wire P1_R1240_U215 , P1_R1240_U216 , P1_R1240_U217 , P1_R1240_U218 , P1_R1240_U219 , P1_R1240_U220 , P1_R1240_U221 , P1_R1240_U222 , P1_R1240_U223 , P1_R1240_U224;
wire P1_R1240_U225 , P1_R1240_U226 , P1_R1240_U227 , P1_R1240_U228 , P1_R1240_U229 , P1_R1240_U230 , P1_R1240_U231 , P1_R1240_U232 , P1_R1240_U233 , P1_R1240_U234;
wire P1_R1240_U235 , P1_R1240_U236 , P1_R1240_U237 , P1_R1240_U238 , P1_R1240_U239 , P1_R1240_U240 , P1_R1240_U241 , P1_R1240_U242 , P1_R1240_U243 , P1_R1240_U244;
wire P1_R1240_U245 , P1_R1240_U246 , P1_R1240_U247 , P1_R1240_U248 , P1_R1240_U249 , P1_R1240_U250 , P1_R1240_U251 , P1_R1240_U252 , P1_R1240_U253 , P1_R1240_U254;
wire P1_R1240_U255 , P1_R1240_U256 , P1_R1240_U257 , P1_R1240_U258 , P1_R1240_U259 , P1_R1240_U260 , P1_R1240_U261 , P1_R1240_U262 , P1_R1240_U263 , P1_R1240_U264;
wire P1_R1240_U265 , P1_R1240_U266 , P1_R1240_U267 , P1_R1240_U268 , P1_R1240_U269 , P1_R1240_U270 , P1_R1240_U271 , P1_R1240_U272 , P1_R1240_U273 , P1_R1240_U274;
wire P1_R1240_U275 , P1_R1240_U276 , P1_R1240_U277 , P1_R1240_U278 , P1_R1240_U279 , P1_R1240_U280 , P1_R1240_U281 , P1_R1240_U282 , P1_R1240_U283 , P1_R1240_U284;
wire P1_R1240_U285 , P1_R1240_U286 , P1_R1240_U287 , P1_R1240_U288 , P1_R1240_U289 , P1_R1240_U290 , P1_R1240_U291 , P1_R1240_U292 , P1_R1240_U293 , P1_R1240_U294;
wire P1_R1240_U295 , P1_R1240_U296 , P1_R1240_U297 , P1_R1240_U298 , P1_R1240_U299 , P1_R1240_U300 , P1_R1240_U301 , P1_R1240_U302 , P1_R1240_U303 , P1_R1240_U304;
wire P1_R1240_U305 , P1_R1240_U306 , P1_R1240_U307 , P1_R1240_U308 , P1_R1240_U309 , P1_R1240_U310 , P1_R1240_U311 , P1_R1240_U312 , P1_R1240_U313 , P1_R1240_U314;
wire P1_R1240_U315 , P1_R1240_U316 , P1_R1240_U317 , P1_R1240_U318 , P1_R1240_U319 , P1_R1240_U320 , P1_R1240_U321 , P1_R1240_U322 , P1_R1240_U323 , P1_R1240_U324;
wire P1_R1240_U325 , P1_R1240_U326 , P1_R1240_U327 , P1_R1240_U328 , P1_R1240_U329 , P1_R1240_U330 , P1_R1240_U331 , P1_R1240_U332 , P1_R1240_U333 , P1_R1240_U334;
wire P1_R1240_U335 , P1_R1240_U336 , P1_R1240_U337 , P1_R1240_U338 , P1_R1240_U339 , P1_R1240_U340 , P1_R1240_U341 , P1_R1240_U342 , P1_R1240_U343 , P1_R1240_U344;
wire P1_R1240_U345 , P1_R1240_U346 , P1_R1240_U347 , P1_R1240_U348 , P1_R1240_U349 , P1_R1240_U350 , P1_R1240_U351 , P1_R1240_U352 , P1_R1240_U353 , P1_R1240_U354;
wire P1_R1240_U355 , P1_R1240_U356 , P1_R1240_U357 , P1_R1240_U358 , P1_R1240_U359 , P1_R1240_U360 , P1_R1240_U361 , P1_R1240_U362 , P1_R1240_U363 , P1_R1240_U364;
wire P1_R1240_U365 , P1_R1240_U366 , P1_R1240_U367 , P1_R1240_U368 , P1_R1240_U369 , P1_R1240_U370 , P1_R1240_U371 , P1_R1240_U372 , P1_R1240_U373 , P1_R1240_U374;
wire P1_R1240_U375 , P1_R1240_U376 , P1_R1240_U377 , P1_R1240_U378 , P1_R1240_U379 , P1_R1240_U380 , P1_R1240_U381 , P1_R1240_U382 , P1_R1240_U383 , P1_R1240_U384;
wire P1_R1240_U385 , P1_R1240_U386 , P1_R1240_U387 , P1_R1240_U388 , P1_R1240_U389 , P1_R1240_U390 , P1_R1240_U391 , P1_R1240_U392 , P1_R1240_U393 , P1_R1240_U394;
wire P1_R1240_U395 , P1_R1240_U396 , P1_R1240_U397 , P1_R1240_U398 , P1_R1240_U399 , P1_R1240_U400 , P1_R1240_U401 , P1_R1240_U402 , P1_R1240_U403 , P1_R1240_U404;
wire P1_R1240_U405 , P1_R1240_U406 , P1_R1240_U407 , P1_R1240_U408 , P1_R1240_U409 , P1_R1240_U410 , P1_R1240_U411 , P1_R1240_U412 , P1_R1240_U413 , P1_R1240_U414;
wire P1_R1240_U415 , P1_R1240_U416 , P1_R1240_U417 , P1_R1240_U418 , P1_R1240_U419 , P1_R1240_U420 , P1_R1240_U421 , P1_R1240_U422 , P1_R1240_U423 , P1_R1240_U424;
wire P1_R1240_U425 , P1_R1240_U426 , P1_R1240_U427 , P1_R1240_U428 , P1_R1240_U429 , P1_R1240_U430 , P1_R1240_U431 , P1_R1240_U432 , P1_R1240_U433 , P1_R1240_U434;
wire P1_R1240_U435 , P1_R1240_U436 , P1_R1240_U437 , P1_R1240_U438 , P1_R1240_U439 , P1_R1240_U440 , P1_R1240_U441 , P1_R1240_U442 , P1_R1240_U443 , P1_R1240_U444;
wire P1_R1240_U445 , P1_R1240_U446 , P1_R1240_U447 , P1_R1240_U448 , P1_R1240_U449 , P1_R1240_U450 , P1_R1240_U451 , P1_R1240_U452 , P1_R1240_U453 , P1_R1240_U454;
wire P1_R1240_U455 , P1_R1240_U456 , P1_R1240_U457 , P1_R1240_U458 , P1_R1240_U459 , P1_R1240_U460 , P1_R1240_U461 , P1_R1240_U462 , P1_R1240_U463 , P1_R1240_U464;
wire P1_R1240_U465 , P1_R1240_U466 , P1_R1240_U467 , P1_R1240_U468 , P1_R1240_U469 , P1_R1240_U470 , P1_R1240_U471 , P1_R1240_U472 , P1_R1240_U473 , P1_R1240_U474;
wire P1_R1240_U475 , P1_R1240_U476 , P1_R1240_U477 , P1_R1240_U478 , P1_R1240_U479 , P1_R1240_U480 , P1_R1240_U481 , P1_R1240_U482 , P1_R1240_U483 , P1_R1240_U484;
wire P1_R1240_U485 , P1_R1240_U486 , P1_R1240_U487 , P1_R1240_U488 , P1_R1240_U489 , P1_R1240_U490 , P1_R1240_U491 , P1_R1240_U492 , P1_R1240_U493 , P1_R1240_U494;
wire P1_R1240_U495 , P1_R1240_U496 , P1_R1240_U497 , P1_R1240_U498 , P1_R1240_U499 , P1_R1240_U500 , P1_R1240_U501 , P1_R1162_U4 , P1_R1162_U5 , P1_R1162_U6;
wire P1_R1162_U7 , P1_R1162_U8 , P1_R1162_U9 , P1_R1162_U10 , P1_R1162_U11 , P1_R1162_U12 , P1_R1162_U13 , P1_R1162_U14 , P1_R1162_U15 , P1_R1162_U16;
wire P1_R1162_U17 , P1_R1162_U18 , P1_R1162_U19 , P1_R1162_U20 , P1_R1162_U21 , P1_R1162_U22 , P1_R1162_U23 , P1_R1162_U24 , P1_R1162_U25 , P1_R1162_U26;
wire P1_R1162_U27 , P1_R1162_U28 , P1_R1162_U29 , P1_R1162_U30 , P1_R1162_U31 , P1_R1162_U32 , P1_R1162_U33 , P1_R1162_U34 , P1_R1162_U35 , P1_R1162_U36;
wire P1_R1162_U37 , P1_R1162_U38 , P1_R1162_U39 , P1_R1162_U40 , P1_R1162_U41 , P1_R1162_U42 , P1_R1162_U43 , P1_R1162_U44 , P1_R1162_U45 , P1_R1162_U46;
wire P1_R1162_U47 , P1_R1162_U48 , P1_R1162_U49 , P1_R1162_U50 , P1_R1162_U51 , P1_R1162_U52 , P1_R1162_U53 , P1_R1162_U54 , P1_R1162_U55 , P1_R1162_U56;
wire P1_R1162_U57 , P1_R1162_U58 , P1_R1162_U59 , P1_R1162_U60 , P1_R1162_U61 , P1_R1162_U62 , P1_R1162_U63 , P1_R1162_U64 , P1_R1162_U65 , P1_R1162_U66;
wire P1_R1162_U67 , P1_R1162_U68 , P1_R1162_U69 , P1_R1162_U70 , P1_R1162_U71 , P1_R1162_U72 , P1_R1162_U73 , P1_R1162_U74 , P1_R1162_U75 , P1_R1162_U76;
wire P1_R1162_U77 , P1_R1162_U78 , P1_R1162_U79 , P1_R1162_U80 , P1_R1162_U81 , P1_R1162_U82 , P1_R1162_U83 , P1_R1162_U84 , P1_R1162_U85 , P1_R1162_U86;
wire P1_R1162_U87 , P1_R1162_U88 , P1_R1162_U89 , P1_R1162_U90 , P1_R1162_U91 , P1_R1162_U92 , P1_R1162_U93 , P1_R1162_U94 , P1_R1162_U95 , P1_R1162_U96;
wire P1_R1162_U97 , P1_R1162_U98 , P1_R1162_U99 , P1_R1162_U100 , P1_R1162_U101 , P1_R1162_U102 , P1_R1162_U103 , P1_R1162_U104 , P1_R1162_U105 , P1_R1162_U106;
wire P1_R1162_U107 , P1_R1162_U108 , P1_R1162_U109 , P1_R1162_U110 , P1_R1162_U111 , P1_R1162_U112 , P1_R1162_U113 , P1_R1162_U114 , P1_R1162_U115 , P1_R1162_U116;
wire P1_R1162_U117 , P1_R1162_U118 , P1_R1162_U119 , P1_R1162_U120 , P1_R1162_U121 , P1_R1162_U122 , P1_R1162_U123 , P1_R1162_U124 , P1_R1162_U125 , P1_R1162_U126;
wire P1_R1162_U127 , P1_R1162_U128 , P1_R1162_U129 , P1_R1162_U130 , P1_R1162_U131 , P1_R1162_U132 , P1_R1162_U133 , P1_R1162_U134 , P1_R1162_U135 , P1_R1162_U136;
wire P1_R1162_U137 , P1_R1162_U138 , P1_R1162_U139 , P1_R1162_U140 , P1_R1162_U141 , P1_R1162_U142 , P1_R1162_U143 , P1_R1162_U144 , P1_R1162_U145 , P1_R1162_U146;
wire P1_R1162_U147 , P1_R1162_U148 , P1_R1162_U149 , P1_R1162_U150 , P1_R1162_U151 , P1_R1162_U152 , P1_R1162_U153 , P1_R1162_U154 , P1_R1162_U155 , P1_R1162_U156;
wire P1_R1162_U157 , P1_R1162_U158 , P1_R1162_U159 , P1_R1162_U160 , P1_R1162_U161 , P1_R1162_U162 , P1_R1162_U163 , P1_R1162_U164 , P1_R1162_U165 , P1_R1162_U166;
wire P1_R1162_U167 , P1_R1162_U168 , P1_R1162_U169 , P1_R1162_U170 , P1_R1162_U171 , P1_R1162_U172 , P1_R1162_U173 , P1_R1162_U174 , P1_R1162_U175 , P1_R1162_U176;
wire P1_R1162_U177 , P1_R1162_U178 , P1_R1162_U179 , P1_R1162_U180 , P1_R1162_U181 , P1_R1162_U182 , P1_R1162_U183 , P1_R1162_U184 , P1_R1162_U185 , P1_R1162_U186;
wire P1_R1162_U187 , P1_R1162_U188 , P1_R1162_U189 , P1_R1162_U190 , P1_R1162_U191 , P1_R1162_U192 , P1_R1162_U193 , P1_R1162_U194 , P1_R1162_U195 , P1_R1162_U196;
wire P1_R1162_U197 , P1_R1162_U198 , P1_R1162_U199 , P1_R1162_U200 , P1_R1162_U201 , P1_R1162_U202 , P1_R1162_U203 , P1_R1162_U204 , P1_R1162_U205 , P1_R1162_U206;
wire P1_R1162_U207 , P1_R1162_U208 , P1_R1162_U209 , P1_R1162_U210 , P1_R1162_U211 , P1_R1162_U212 , P1_R1162_U213 , P1_R1162_U214 , P1_R1162_U215 , P1_R1162_U216;
wire P1_R1162_U217 , P1_R1162_U218 , P1_R1162_U219 , P1_R1162_U220 , P1_R1162_U221 , P1_R1162_U222 , P1_R1162_U223 , P1_R1162_U224 , P1_R1162_U225 , P1_R1162_U226;
wire P1_R1162_U227 , P1_R1162_U228 , P1_R1162_U229 , P1_R1162_U230 , P1_R1162_U231 , P1_R1162_U232 , P1_R1162_U233 , P1_R1162_U234 , P1_R1162_U235 , P1_R1162_U236;
wire P1_R1162_U237 , P1_R1162_U238 , P1_R1162_U239 , P1_R1162_U240 , P1_R1162_U241 , P1_R1162_U242 , P1_R1162_U243 , P1_R1162_U244 , P1_R1162_U245 , P1_R1162_U246;
wire P1_R1162_U247 , P1_R1162_U248 , P1_R1162_U249 , P1_R1162_U250 , P1_R1162_U251 , P1_R1162_U252 , P1_R1162_U253 , P1_R1162_U254 , P1_R1162_U255 , P1_R1162_U256;
wire P1_R1162_U257 , P1_R1162_U258 , P1_R1162_U259 , P1_R1162_U260 , P1_R1162_U261 , P1_R1162_U262 , P1_R1162_U263 , P1_R1162_U264 , P1_R1162_U265 , P1_R1162_U266;
wire P1_R1162_U267 , P1_R1162_U268 , P1_R1162_U269 , P1_R1162_U270 , P1_R1162_U271 , P1_R1162_U272 , P1_R1162_U273 , P1_R1162_U274 , P1_R1162_U275 , P1_R1162_U276;
wire P1_R1162_U277 , P1_R1162_U278 , P1_R1162_U279 , P1_R1162_U280 , P1_R1162_U281 , P1_R1162_U282 , P1_R1162_U283 , P1_R1162_U284 , P1_R1162_U285 , P1_R1162_U286;
wire P1_R1162_U287 , P1_R1162_U288 , P1_R1162_U289 , P1_R1162_U290 , P1_R1162_U291 , P1_R1162_U292 , P1_R1162_U293 , P1_R1162_U294 , P1_R1162_U295 , P1_R1162_U296;
wire P1_R1162_U297 , P1_R1162_U298 , P1_R1162_U299 , P1_R1162_U300 , P1_R1162_U301 , P1_R1162_U302 , P1_R1162_U303 , P1_R1162_U304 , P1_R1162_U305 , P1_R1162_U306;
wire P1_R1162_U307 , P1_R1162_U308 , P1_R1117_U6 , P1_R1117_U7 , P1_R1117_U8 , P1_R1117_U9 , P1_R1117_U10 , P1_R1117_U11 , P1_R1117_U12 , P1_R1117_U13;
wire P1_R1117_U14 , P1_R1117_U15 , P1_R1117_U16 , P1_R1117_U17 , P1_R1117_U18 , P1_R1117_U19 , P1_R1117_U20 , P1_R1117_U21 , P1_R1117_U22 , P1_R1117_U23;
wire P1_R1117_U24 , P1_R1117_U25 , P1_R1117_U26 , P1_R1117_U27 , P1_R1117_U28 , P1_R1117_U29 , P1_R1117_U30 , P1_R1117_U31 , P1_R1117_U32 , P1_R1117_U33;
wire P1_R1117_U34 , P1_R1117_U35 , P1_R1117_U36 , P1_R1117_U37 , P1_R1117_U38 , P1_R1117_U39 , P1_R1117_U40 , P1_R1117_U41 , P1_R1117_U42 , P1_R1117_U43;
wire P1_R1117_U44 , P1_R1117_U45 , P1_R1117_U46 , P1_R1117_U47 , P1_R1117_U48 , P1_R1117_U49 , P1_R1117_U50 , P1_R1117_U51 , P1_R1117_U52 , P1_R1117_U53;
wire P1_R1117_U54 , P1_R1117_U55 , P1_R1117_U56 , P1_R1117_U57 , P1_R1117_U58 , P1_R1117_U59 , P1_R1117_U60 , P1_R1117_U61 , P1_R1117_U62 , P1_R1117_U63;
wire P1_R1117_U64 , P1_R1117_U65 , P1_R1117_U66 , P1_R1117_U67 , P1_R1117_U68 , P1_R1117_U69 , P1_R1117_U70 , P1_R1117_U71 , P1_R1117_U72 , P1_R1117_U73;
wire P1_R1117_U74 , P1_R1117_U75 , P1_R1117_U76 , P1_R1117_U77 , P1_R1117_U78 , P1_R1117_U79 , P1_R1117_U80 , P1_R1117_U81 , P1_R1117_U82 , P1_R1117_U83;
wire P1_R1117_U84 , P1_R1117_U85 , P1_R1117_U86 , P1_R1117_U87 , P1_R1117_U88 , P1_R1117_U89 , P1_R1117_U90 , P1_R1117_U91 , P1_R1117_U92 , P1_R1117_U93;
wire P1_R1117_U94 , P1_R1117_U95 , P1_R1117_U96 , P1_R1117_U97 , P1_R1117_U98 , P1_R1117_U99 , P1_R1117_U100 , P1_R1117_U101 , P1_R1117_U102 , P1_R1117_U103;
wire P1_R1117_U104 , P1_R1117_U105 , P1_R1117_U106 , P1_R1117_U107 , P1_R1117_U108 , P1_R1117_U109 , P1_R1117_U110 , P1_R1117_U111 , P1_R1117_U112 , P1_R1117_U113;
wire P1_R1117_U114 , P1_R1117_U115 , P1_R1117_U116 , P1_R1117_U117 , P1_R1117_U118 , P1_R1117_U119 , P1_R1117_U120 , P1_R1117_U121 , P1_R1117_U122 , P1_R1117_U123;
wire P1_R1117_U124 , P1_R1117_U125 , P1_R1117_U126 , P1_R1117_U127 , P1_R1117_U128 , P1_R1117_U129 , P1_R1117_U130 , P1_R1117_U131 , P1_R1117_U132 , P1_R1117_U133;
wire P1_R1117_U134 , P1_R1117_U135 , P1_R1117_U136 , P1_R1117_U137 , P1_R1117_U138 , P1_R1117_U139 , P1_R1117_U140 , P1_R1117_U141 , P1_R1117_U142 , P1_R1117_U143;
wire P1_R1117_U144 , P1_R1117_U145 , P1_R1117_U146 , P1_R1117_U147 , P1_R1117_U148 , P1_R1117_U149 , P1_R1117_U150 , P1_R1117_U151 , P1_R1117_U152 , P1_R1117_U153;
wire P1_R1117_U154 , P1_R1117_U155 , P1_R1117_U156 , P1_R1117_U157 , P1_R1117_U158 , P1_R1117_U159 , P1_R1117_U160 , P1_R1117_U161 , P1_R1117_U162 , P1_R1117_U163;
wire P1_R1117_U164 , P1_R1117_U165 , P1_R1117_U166 , P1_R1117_U167 , P1_R1117_U168 , P1_R1117_U169 , P1_R1117_U170 , P1_R1117_U171 , P1_R1117_U172 , P1_R1117_U173;
wire P1_R1117_U174 , P1_R1117_U175 , P1_R1117_U176 , P1_R1117_U177 , P1_R1117_U178 , P1_R1117_U179 , P1_R1117_U180 , P1_R1117_U181 , P1_R1117_U182 , P1_R1117_U183;
wire P1_R1117_U184 , P1_R1117_U185 , P1_R1117_U186 , P1_R1117_U187 , P1_R1117_U188 , P1_R1117_U189 , P1_R1117_U190 , P1_R1117_U191 , P1_R1117_U192 , P1_R1117_U193;
wire P1_R1117_U194 , P1_R1117_U195 , P1_R1117_U196 , P1_R1117_U197 , P1_R1117_U198 , P1_R1117_U199 , P1_R1117_U200 , P1_R1117_U201 , P1_R1117_U202 , P1_R1117_U203;
wire P1_R1117_U204 , P1_R1117_U205 , P1_R1117_U206 , P1_R1117_U207 , P1_R1117_U208 , P1_R1117_U209 , P1_R1117_U210 , P1_R1117_U211 , P1_R1117_U212 , P1_R1117_U213;
wire P1_R1117_U214 , P1_R1117_U215 , P1_R1117_U216 , P1_R1117_U217 , P1_R1117_U218 , P1_R1117_U219 , P1_R1117_U220 , P1_R1117_U221 , P1_R1117_U222 , P1_R1117_U223;
wire P1_R1117_U224 , P1_R1117_U225 , P1_R1117_U226 , P1_R1117_U227 , P1_R1117_U228 , P1_R1117_U229 , P1_R1117_U230 , P1_R1117_U231 , P1_R1117_U232 , P1_R1117_U233;
wire P1_R1117_U234 , P1_R1117_U235 , P1_R1117_U236 , P1_R1117_U237 , P1_R1117_U238 , P1_R1117_U239 , P1_R1117_U240 , P1_R1117_U241 , P1_R1117_U242 , P1_R1117_U243;
wire P1_R1117_U244 , P1_R1117_U245 , P1_R1117_U246 , P1_R1117_U247 , P1_R1117_U248 , P1_R1117_U249 , P1_R1117_U250 , P1_R1117_U251 , P1_R1117_U252 , P1_R1117_U253;
wire P1_R1117_U254 , P1_R1117_U255 , P1_R1117_U256 , P1_R1117_U257 , P1_R1117_U258 , P1_R1117_U259 , P1_R1117_U260 , P1_R1117_U261 , P1_R1117_U262 , P1_R1117_U263;
wire P1_R1117_U264 , P1_R1117_U265 , P1_R1117_U266 , P1_R1117_U267 , P1_R1117_U268 , P1_R1117_U269 , P1_R1117_U270 , P1_R1117_U271 , P1_R1117_U272 , P1_R1117_U273;
wire P1_R1117_U274 , P1_R1117_U275 , P1_R1117_U276 , P1_R1117_U277 , P1_R1117_U278 , P1_R1117_U279 , P1_R1117_U280 , P1_R1117_U281 , P1_R1117_U282 , P1_R1117_U283;
wire P1_R1117_U284 , P1_R1117_U285 , P1_R1117_U286 , P1_R1117_U287 , P1_R1117_U288 , P1_R1117_U289 , P1_R1117_U290 , P1_R1117_U291 , P1_R1117_U292 , P1_R1117_U293;
wire P1_R1117_U294 , P1_R1117_U295 , P1_R1117_U296 , P1_R1117_U297 , P1_R1117_U298 , P1_R1117_U299 , P1_R1117_U300 , P1_R1117_U301 , P1_R1117_U302 , P1_R1117_U303;
wire P1_R1117_U304 , P1_R1117_U305 , P1_R1117_U306 , P1_R1117_U307 , P1_R1117_U308 , P1_R1117_U309 , P1_R1117_U310 , P1_R1117_U311 , P1_R1117_U312 , P1_R1117_U313;
wire P1_R1117_U314 , P1_R1117_U315 , P1_R1117_U316 , P1_R1117_U317 , P1_R1117_U318 , P1_R1117_U319 , P1_R1117_U320 , P1_R1117_U321 , P1_R1117_U322 , P1_R1117_U323;
wire P1_R1117_U324 , P1_R1117_U325 , P1_R1117_U326 , P1_R1117_U327 , P1_R1117_U328 , P1_R1117_U329 , P1_R1117_U330 , P1_R1117_U331 , P1_R1117_U332 , P1_R1117_U333;
wire P1_R1117_U334 , P1_R1117_U335 , P1_R1117_U336 , P1_R1117_U337 , P1_R1117_U338 , P1_R1117_U339 , P1_R1117_U340 , P1_R1117_U341 , P1_R1117_U342 , P1_R1117_U343;
wire P1_R1117_U344 , P1_R1117_U345 , P1_R1117_U346 , P1_R1117_U347 , P1_R1117_U348 , P1_R1117_U349 , P1_R1117_U350 , P1_R1117_U351 , P1_R1117_U352 , P1_R1117_U353;
wire P1_R1117_U354 , P1_R1117_U355 , P1_R1117_U356 , P1_R1117_U357 , P1_R1117_U358 , P1_R1117_U359 , P1_R1117_U360 , P1_R1117_U361 , P1_R1117_U362 , P1_R1117_U363;
wire P1_R1117_U364 , P1_R1117_U365 , P1_R1117_U366 , P1_R1117_U367 , P1_R1117_U368 , P1_R1117_U369 , P1_R1117_U370 , P1_R1117_U371 , P1_R1117_U372 , P1_R1117_U373;
wire P1_R1117_U374 , P1_R1117_U375 , P1_R1117_U376 , P1_R1117_U377 , P1_R1117_U378 , P1_R1117_U379 , P1_R1117_U380 , P1_R1117_U381 , P1_R1117_U382 , P1_R1117_U383;
wire P1_R1117_U384 , P1_R1117_U385 , P1_R1117_U386 , P1_R1117_U387 , P1_R1117_U388 , P1_R1117_U389 , P1_R1117_U390 , P1_R1117_U391 , P1_R1117_U392 , P1_R1117_U393;
wire P1_R1117_U394 , P1_R1117_U395 , P1_R1117_U396 , P1_R1117_U397 , P1_R1117_U398 , P1_R1117_U399 , P1_R1117_U400 , P1_R1117_U401 , P1_R1117_U402 , P1_R1117_U403;
wire P1_R1117_U404 , P1_R1117_U405 , P1_R1117_U406 , P1_R1117_U407 , P1_R1117_U408 , P1_R1117_U409 , P1_R1117_U410 , P1_R1117_U411 , P1_R1117_U412 , P1_R1117_U413;
wire P1_R1117_U414 , P1_R1117_U415 , P1_R1117_U416 , P1_R1117_U417 , P1_R1117_U418 , P1_R1117_U419 , P1_R1117_U420 , P1_R1117_U421 , P1_R1117_U422 , P1_R1117_U423;
wire P1_R1117_U424 , P1_R1117_U425 , P1_R1117_U426 , P1_R1117_U427 , P1_R1117_U428 , P1_R1117_U429 , P1_R1117_U430 , P1_R1117_U431 , P1_R1117_U432 , P1_R1117_U433;
wire P1_R1117_U434 , P1_R1117_U435 , P1_R1117_U436 , P1_R1117_U437 , P1_R1117_U438 , P1_R1117_U439 , P1_R1117_U440 , P1_R1117_U441 , P1_R1117_U442 , P1_R1117_U443;
wire P1_R1117_U444 , P1_R1117_U445 , P1_R1117_U446 , P1_R1117_U447 , P1_R1117_U448 , P1_R1117_U449 , P1_R1117_U450 , P1_R1117_U451 , P1_R1117_U452 , P1_R1117_U453;
wire P1_R1117_U454 , P1_R1117_U455 , P1_R1117_U456 , P1_R1117_U457 , P1_R1117_U458 , P1_R1117_U459 , P1_R1117_U460 , P1_R1117_U461 , P1_R1117_U462 , P1_R1117_U463;
wire P1_R1117_U464 , P1_R1117_U465 , P1_R1117_U466 , P1_R1117_U467 , P1_R1117_U468 , P1_R1117_U469 , P1_R1117_U470 , P1_R1117_U471 , P1_R1117_U472 , P1_R1117_U473;
wire P1_R1117_U474 , P1_R1117_U475 , P1_R1117_U476 , P1_R1375_U6 , P1_R1375_U7 , P1_R1375_U8 , P1_R1375_U9 , P1_R1375_U10 , P1_R1375_U11 , P1_R1375_U12;
wire P1_R1375_U13 , P1_R1375_U14 , P1_R1375_U15 , P1_R1375_U16 , P1_R1375_U17 , P1_R1375_U18 , P1_R1375_U19 , P1_R1375_U20 , P1_R1375_U21 , P1_R1375_U22;
wire P1_R1375_U23 , P1_R1375_U24 , P1_R1375_U25 , P1_R1375_U26 , P1_R1375_U27 , P1_R1375_U28 , P1_R1375_U29 , P1_R1375_U30 , P1_R1375_U31 , P1_R1375_U32;
wire P1_R1375_U33 , P1_R1375_U34 , P1_R1375_U35 , P1_R1375_U36 , P1_R1375_U37 , P1_R1375_U38 , P1_R1375_U39 , P1_R1375_U40 , P1_R1375_U41 , P1_R1375_U42;
wire P1_R1375_U43 , P1_R1375_U44 , P1_R1375_U45 , P1_R1375_U46 , P1_R1375_U47 , P1_R1375_U48 , P1_R1375_U49 , P1_R1375_U50 , P1_R1375_U51 , P1_R1375_U52;
wire P1_R1375_U53 , P1_R1375_U54 , P1_R1375_U55 , P1_R1375_U56 , P1_R1375_U57 , P1_R1375_U58 , P1_R1375_U59 , P1_R1375_U60 , P1_R1375_U61 , P1_R1375_U62;
wire P1_R1375_U63 , P1_R1375_U64 , P1_R1375_U65 , P1_R1375_U66 , P1_R1375_U67 , P1_R1375_U68 , P1_R1375_U69 , P1_R1375_U70 , P1_R1375_U71 , P1_R1375_U72;
wire P1_R1375_U73 , P1_R1375_U74 , P1_R1375_U75 , P1_R1375_U76 , P1_R1375_U77 , P1_R1375_U78 , P1_R1375_U79 , P1_R1375_U80 , P1_R1375_U81 , P1_R1375_U82;
wire P1_R1375_U83 , P1_R1375_U84 , P1_R1375_U85 , P1_R1375_U86 , P1_R1375_U87 , P1_R1375_U88 , P1_R1375_U89 , P1_R1375_U90 , P1_R1375_U91 , P1_R1375_U92;
wire P1_R1375_U93 , P1_R1375_U94 , P1_R1375_U95 , P1_R1375_U96 , P1_R1375_U97 , P1_R1375_U98 , P1_R1375_U99 , P1_R1375_U100 , P1_R1375_U101 , P1_R1375_U102;
wire P1_R1375_U103 , P1_R1375_U104 , P1_R1375_U105 , P1_R1375_U106 , P1_R1375_U107 , P1_R1375_U108 , P1_R1375_U109 , P1_R1375_U110 , P1_R1375_U111 , P1_R1375_U112;
wire P1_R1375_U113 , P1_R1375_U114 , P1_R1375_U115 , P1_R1375_U116 , P1_R1375_U117 , P1_R1375_U118 , P1_R1375_U119 , P1_R1375_U120 , P1_R1375_U121 , P1_R1375_U122;
wire P1_R1375_U123 , P1_R1375_U124 , P1_R1375_U125 , P1_R1375_U126 , P1_R1375_U127 , P1_R1375_U128 , P1_R1375_U129 , P1_R1375_U130 , P1_R1375_U131 , P1_R1375_U132;
wire P1_R1375_U133 , P1_R1375_U134 , P1_R1375_U135 , P1_R1375_U136 , P1_R1375_U137 , P1_R1375_U138 , P1_R1375_U139 , P1_R1375_U140 , P1_R1375_U141 , P1_R1375_U142;
wire P1_R1375_U143 , P1_R1375_U144 , P1_R1375_U145 , P1_R1375_U146 , P1_R1375_U147 , P1_R1375_U148 , P1_R1375_U149 , P1_R1375_U150 , P1_R1375_U151 , P1_R1375_U152;
wire P1_R1375_U153 , P1_R1375_U154 , P1_R1375_U155 , P1_R1375_U156 , P1_R1375_U157 , P1_R1375_U158 , P1_R1375_U159 , P1_R1375_U160 , P1_R1375_U161 , P1_R1375_U162;
wire P1_R1375_U163 , P1_R1375_U164 , P1_R1375_U165 , P1_R1375_U166 , P1_R1375_U167 , P1_R1375_U168 , P1_R1375_U169 , P1_R1375_U170 , P1_R1375_U171 , P1_R1375_U172;
wire P1_R1375_U173 , P1_R1375_U174 , P1_R1375_U175 , P1_R1375_U176 , P1_R1375_U177 , P1_R1375_U178 , P1_R1375_U179 , P1_R1375_U180 , P1_R1375_U181 , P1_R1375_U182;
wire P1_R1375_U183 , P1_R1375_U184 , P1_R1375_U185 , P1_R1375_U186 , P1_R1375_U187 , P1_R1375_U188 , P1_R1375_U189 , P1_R1375_U190 , P1_R1375_U191 , P1_R1375_U192;
wire P1_R1375_U193 , P1_R1375_U194 , P1_R1375_U195 , P1_R1375_U196 , P1_R1375_U197 , P1_R1352_U6 , P1_R1352_U7 , P1_R1207_U6 , P1_R1207_U7 , P1_R1207_U8;
wire P1_R1207_U9 , P1_R1207_U10 , P1_R1207_U11 , P1_R1207_U12 , P1_R1207_U13 , P1_R1207_U14 , P1_R1207_U15 , P1_R1207_U16 , P1_R1207_U17 , P1_R1207_U18;
wire P1_R1207_U19 , P1_R1207_U20 , P1_R1207_U21 , P1_R1207_U22 , P1_R1207_U23 , P1_R1207_U24 , P1_R1207_U25 , P1_R1207_U26 , P1_R1207_U27 , P1_R1207_U28;
wire P1_R1207_U29 , P1_R1207_U30 , P1_R1207_U31 , P1_R1207_U32 , P1_R1207_U33 , P1_R1207_U34 , P1_R1207_U35 , P1_R1207_U36 , P1_R1207_U37 , P1_R1207_U38;
wire P1_R1207_U39 , P1_R1207_U40 , P1_R1207_U41 , P1_R1207_U42 , P1_R1207_U43 , P1_R1207_U44 , P1_R1207_U45 , P1_R1207_U46 , P1_R1207_U47 , P1_R1207_U48;
wire P1_R1207_U49 , P1_R1207_U50 , P1_R1207_U51 , P1_R1207_U52 , P1_R1207_U53 , P1_R1207_U54 , P1_R1207_U55 , P1_R1207_U56 , P1_R1207_U57 , P1_R1207_U58;
wire P1_R1207_U59 , P1_R1207_U60 , P1_R1207_U61 , P1_R1207_U62 , P1_R1207_U63 , P1_R1207_U64 , P1_R1207_U65 , P1_R1207_U66 , P1_R1207_U67 , P1_R1207_U68;
wire P1_R1207_U69 , P1_R1207_U70 , P1_R1207_U71 , P1_R1207_U72 , P1_R1207_U73 , P1_R1207_U74 , P1_R1207_U75 , P1_R1207_U76 , P1_R1207_U77 , P1_R1207_U78;
wire P1_R1207_U79 , P1_R1207_U80 , P1_R1207_U81 , P1_R1207_U82 , P1_R1207_U83 , P1_R1207_U84 , P1_R1207_U85 , P1_R1207_U86 , P1_R1207_U87 , P1_R1207_U88;
wire P1_R1207_U89 , P1_R1207_U90 , P1_R1207_U91 , P1_R1207_U92 , P1_R1207_U93 , P1_R1207_U94 , P1_R1207_U95 , P1_R1207_U96 , P1_R1207_U97 , P1_R1207_U98;
wire P1_R1207_U99 , P1_R1207_U100 , P1_R1207_U101 , P1_R1207_U102 , P1_R1207_U103 , P1_R1207_U104 , P1_R1207_U105 , P1_R1207_U106 , P1_R1207_U107 , P1_R1207_U108;
wire P1_R1207_U109 , P1_R1207_U110 , P1_R1207_U111 , P1_R1207_U112 , P1_R1207_U113 , P1_R1207_U114 , P1_R1207_U115 , P1_R1207_U116 , P1_R1207_U117 , P1_R1207_U118;
wire P1_R1207_U119 , P1_R1207_U120 , P1_R1207_U121 , P1_R1207_U122 , P1_R1207_U123 , P1_R1207_U124 , P1_R1207_U125 , P1_R1207_U126 , P1_R1207_U127 , P1_R1207_U128;
wire P1_R1207_U129 , P1_R1207_U130 , P1_R1207_U131 , P1_R1207_U132 , P1_R1207_U133 , P1_R1207_U134 , P1_R1207_U135 , P1_R1207_U136 , P1_R1207_U137 , P1_R1207_U138;
wire P1_R1207_U139 , P1_R1207_U140 , P1_R1207_U141 , P1_R1207_U142 , P1_R1207_U143 , P1_R1207_U144 , P1_R1207_U145 , P1_R1207_U146 , P1_R1207_U147 , P1_R1207_U148;
wire P1_R1207_U149 , P1_R1207_U150 , P1_R1207_U151 , P1_R1207_U152 , P1_R1207_U153 , P1_R1207_U154 , P1_R1207_U155 , P1_R1207_U156 , P1_R1207_U157 , P1_R1207_U158;
wire P1_R1207_U159 , P1_R1207_U160 , P1_R1207_U161 , P1_R1207_U162 , P1_R1207_U163 , P1_R1207_U164 , P1_R1207_U165 , P1_R1207_U166 , P1_R1207_U167 , P1_R1207_U168;
wire P1_R1207_U169 , P1_R1207_U170 , P1_R1207_U171 , P1_R1207_U172 , P1_R1207_U173 , P1_R1207_U174 , P1_R1207_U175 , P1_R1207_U176 , P1_R1207_U177 , P1_R1207_U178;
wire P1_R1207_U179 , P1_R1207_U180 , P1_R1207_U181 , P1_R1207_U182 , P1_R1207_U183 , P1_R1207_U184 , P1_R1207_U185 , P1_R1207_U186 , P1_R1207_U187 , P1_R1207_U188;
wire P1_R1207_U189 , P1_R1207_U190 , P1_R1207_U191 , P1_R1207_U192 , P1_R1207_U193 , P1_R1207_U194 , P1_R1207_U195 , P1_R1207_U196 , P1_R1207_U197 , P1_R1207_U198;
wire P1_R1207_U199 , P1_R1207_U200 , P1_R1207_U201 , P1_R1207_U202 , P1_R1207_U203 , P1_R1207_U204 , P1_R1207_U205 , P1_R1207_U206 , P1_R1207_U207 , P1_R1207_U208;
wire P1_R1207_U209 , P1_R1207_U210 , P1_R1207_U211 , P1_R1207_U212 , P1_R1207_U213 , P1_R1207_U214 , P1_R1207_U215 , P1_R1207_U216 , P1_R1207_U217 , P1_R1207_U218;
wire P1_R1207_U219 , P1_R1207_U220 , P1_R1207_U221 , P1_R1207_U222 , P1_R1207_U223 , P1_R1207_U224 , P1_R1207_U225 , P1_R1207_U226 , P1_R1207_U227 , P1_R1207_U228;
wire P1_R1207_U229 , P1_R1207_U230 , P1_R1207_U231 , P1_R1207_U232 , P1_R1207_U233 , P1_R1207_U234 , P1_R1207_U235 , P1_R1207_U236 , P1_R1207_U237 , P1_R1207_U238;
wire P1_R1207_U239 , P1_R1207_U240 , P1_R1207_U241 , P1_R1207_U242 , P1_R1207_U243 , P1_R1207_U244 , P1_R1207_U245 , P1_R1207_U246 , P1_R1207_U247 , P1_R1207_U248;
wire P1_R1207_U249 , P1_R1207_U250 , P1_R1207_U251 , P1_R1207_U252 , P1_R1207_U253 , P1_R1207_U254 , P1_R1207_U255 , P1_R1207_U256 , P1_R1207_U257 , P1_R1207_U258;
wire P1_R1207_U259 , P1_R1207_U260 , P1_R1207_U261 , P1_R1207_U262 , P1_R1207_U263 , P1_R1207_U264 , P1_R1207_U265 , P1_R1207_U266 , P1_R1207_U267 , P1_R1207_U268;
wire P1_R1207_U269 , P1_R1207_U270 , P1_R1207_U271 , P1_R1207_U272 , P1_R1207_U273 , P1_R1207_U274 , P1_R1207_U275 , P1_R1207_U276 , P1_R1207_U277 , P1_R1207_U278;
wire P1_R1207_U279 , P1_R1207_U280 , P1_R1207_U281 , P1_R1207_U282 , P1_R1207_U283 , P1_R1207_U284 , P1_R1207_U285 , P1_R1207_U286 , P1_R1207_U287 , P1_R1207_U288;
wire P1_R1207_U289 , P1_R1207_U290 , P1_R1207_U291 , P1_R1207_U292 , P1_R1207_U293 , P1_R1207_U294 , P1_R1207_U295 , P1_R1207_U296 , P1_R1207_U297 , P1_R1207_U298;
wire P1_R1207_U299 , P1_R1207_U300 , P1_R1207_U301 , P1_R1207_U302 , P1_R1207_U303 , P1_R1207_U304 , P1_R1207_U305 , P1_R1207_U306 , P1_R1207_U307 , P1_R1207_U308;
wire P1_R1207_U309 , P1_R1207_U310 , P1_R1207_U311 , P1_R1207_U312 , P1_R1207_U313 , P1_R1207_U314 , P1_R1207_U315 , P1_R1207_U316 , P1_R1207_U317 , P1_R1207_U318;
wire P1_R1207_U319 , P1_R1207_U320 , P1_R1207_U321 , P1_R1207_U322 , P1_R1207_U323 , P1_R1207_U324 , P1_R1207_U325 , P1_R1207_U326 , P1_R1207_U327 , P1_R1207_U328;
wire P1_R1207_U329 , P1_R1207_U330 , P1_R1207_U331 , P1_R1207_U332 , P1_R1207_U333 , P1_R1207_U334 , P1_R1207_U335 , P1_R1207_U336 , P1_R1207_U337 , P1_R1207_U338;
wire P1_R1207_U339 , P1_R1207_U340 , P1_R1207_U341 , P1_R1207_U342 , P1_R1207_U343 , P1_R1207_U344 , P1_R1207_U345 , P1_R1207_U346 , P1_R1207_U347 , P1_R1207_U348;
wire P1_R1207_U349 , P1_R1207_U350 , P1_R1207_U351 , P1_R1207_U352 , P1_R1207_U353 , P1_R1207_U354 , P1_R1207_U355 , P1_R1207_U356 , P1_R1207_U357 , P1_R1207_U358;
wire P1_R1207_U359 , P1_R1207_U360 , P1_R1207_U361 , P1_R1207_U362 , P1_R1207_U363 , P1_R1207_U364 , P1_R1207_U365 , P1_R1207_U366 , P1_R1207_U367 , P1_R1207_U368;
wire P1_R1207_U369 , P1_R1207_U370 , P1_R1207_U371 , P1_R1207_U372 , P1_R1207_U373 , P1_R1207_U374 , P1_R1207_U375 , P1_R1207_U376 , P1_R1207_U377 , P1_R1207_U378;
wire P1_R1207_U379 , P1_R1207_U380 , P1_R1207_U381 , P1_R1207_U382 , P1_R1207_U383 , P1_R1207_U384 , P1_R1207_U385 , P1_R1207_U386 , P1_R1207_U387 , P1_R1207_U388;
wire P1_R1207_U389 , P1_R1207_U390 , P1_R1207_U391 , P1_R1207_U392 , P1_R1207_U393 , P1_R1207_U394 , P1_R1207_U395 , P1_R1207_U396 , P1_R1207_U397 , P1_R1207_U398;
wire P1_R1207_U399 , P1_R1207_U400 , P1_R1207_U401 , P1_R1207_U402 , P1_R1207_U403 , P1_R1207_U404 , P1_R1207_U405 , P1_R1207_U406 , P1_R1207_U407 , P1_R1207_U408;
wire P1_R1207_U409 , P1_R1207_U410 , P1_R1207_U411 , P1_R1207_U412 , P1_R1207_U413 , P1_R1207_U414 , P1_R1207_U415 , P1_R1207_U416 , P1_R1207_U417 , P1_R1207_U418;
wire P1_R1207_U419 , P1_R1207_U420 , P1_R1207_U421 , P1_R1207_U422 , P1_R1207_U423 , P1_R1207_U424 , P1_R1207_U425 , P1_R1207_U426 , P1_R1207_U427 , P1_R1207_U428;
wire P1_R1207_U429 , P1_R1207_U430 , P1_R1207_U431 , P1_R1207_U432 , P1_R1207_U433 , P1_R1207_U434 , P1_R1207_U435 , P1_R1207_U436 , P1_R1207_U437 , P1_R1207_U438;
wire P1_R1207_U439 , P1_R1207_U440 , P1_R1207_U441 , P1_R1207_U442 , P1_R1207_U443 , P1_R1207_U444 , P1_R1207_U445 , P1_R1207_U446 , P1_R1207_U447 , P1_R1207_U448;
wire P1_R1207_U449 , P1_R1207_U450 , P1_R1207_U451 , P1_R1207_U452 , P1_R1207_U453 , P1_R1207_U454 , P1_R1207_U455 , P1_R1207_U456 , P1_R1207_U457 , P1_R1207_U458;
wire P1_R1207_U459 , P1_R1207_U460 , P1_R1207_U461 , P1_R1207_U462 , P1_R1207_U463 , P1_R1207_U464 , P1_R1207_U465 , P1_R1207_U466 , P1_R1207_U467 , P1_R1207_U468;
wire P1_R1207_U469 , P1_R1207_U470 , P1_R1207_U471 , P1_R1207_U472 , P1_R1207_U473 , P1_R1207_U474 , P1_R1207_U475 , P1_R1207_U476 , P1_R1165_U4 , P1_R1165_U5;
wire P1_R1165_U6 , P1_R1165_U7 , P1_R1165_U8 , P1_R1165_U9 , P1_R1165_U10 , P1_R1165_U11 , P1_R1165_U12 , P1_R1165_U13 , P1_R1165_U14 , P1_R1165_U15;
wire P1_R1165_U16 , P1_R1165_U17 , P1_R1165_U18 , P1_R1165_U19 , P1_R1165_U20 , P1_R1165_U21 , P1_R1165_U22 , P1_R1165_U23 , P1_R1165_U24 , P1_R1165_U25;
wire P1_R1165_U26 , P1_R1165_U27 , P1_R1165_U28 , P1_R1165_U29 , P1_R1165_U30 , P1_R1165_U31 , P1_R1165_U32 , P1_R1165_U33 , P1_R1165_U34 , P1_R1165_U35;
wire P1_R1165_U36 , P1_R1165_U37 , P1_R1165_U38 , P1_R1165_U39 , P1_R1165_U40 , P1_R1165_U41 , P1_R1165_U42 , P1_R1165_U43 , P1_R1165_U44 , P1_R1165_U45;
wire P1_R1165_U46 , P1_R1165_U47 , P1_R1165_U48 , P1_R1165_U49 , P1_R1165_U50 , P1_R1165_U51 , P1_R1165_U52 , P1_R1165_U53 , P1_R1165_U54 , P1_R1165_U55;
wire P1_R1165_U56 , P1_R1165_U57 , P1_R1165_U58 , P1_R1165_U59 , P1_R1165_U60 , P1_R1165_U61 , P1_R1165_U62 , P1_R1165_U63 , P1_R1165_U64 , P1_R1165_U65;
wire P1_R1165_U66 , P1_R1165_U67 , P1_R1165_U68 , P1_R1165_U69 , P1_R1165_U70 , P1_R1165_U71 , P1_R1165_U72 , P1_R1165_U73 , P1_R1165_U74 , P1_R1165_U75;
wire P1_R1165_U76 , P1_R1165_U77 , P1_R1165_U78 , P1_R1165_U79 , P1_R1165_U80 , P1_R1165_U81 , P1_R1165_U82 , P1_R1165_U83 , P1_R1165_U84 , P1_R1165_U85;
wire P1_R1165_U86 , P1_R1165_U87 , P1_R1165_U88 , P1_R1165_U89 , P1_R1165_U90 , P1_R1165_U91 , P1_R1165_U92 , P1_R1165_U93 , P1_R1165_U94 , P1_R1165_U95;
wire P1_R1165_U96 , P1_R1165_U97 , P1_R1165_U98 , P1_R1165_U99 , P1_R1165_U100 , P1_R1165_U101 , P1_R1165_U102 , P1_R1165_U103 , P1_R1165_U104 , P1_R1165_U105;
wire P1_R1165_U106 , P1_R1165_U107 , P1_R1165_U108 , P1_R1165_U109 , P1_R1165_U110 , P1_R1165_U111 , P1_R1165_U112 , P1_R1165_U113 , P1_R1165_U114 , P1_R1165_U115;
wire P1_R1165_U116 , P1_R1165_U117 , P1_R1165_U118 , P1_R1165_U119 , P1_R1165_U120 , P1_R1165_U121 , P1_R1165_U122 , P1_R1165_U123 , P1_R1165_U124 , P1_R1165_U125;
wire P1_R1165_U126 , P1_R1165_U127 , P1_R1165_U128 , P1_R1165_U129 , P1_R1165_U130 , P1_R1165_U131 , P1_R1165_U132 , P1_R1165_U133 , P1_R1165_U134 , P1_R1165_U135;
wire P1_R1165_U136 , P1_R1165_U137 , P1_R1165_U138 , P1_R1165_U139 , P1_R1165_U140 , P1_R1165_U141 , P1_R1165_U142 , P1_R1165_U143 , P1_R1165_U144 , P1_R1165_U145;
wire P1_R1165_U146 , P1_R1165_U147 , P1_R1165_U148 , P1_R1165_U149 , P1_R1165_U150 , P1_R1165_U151 , P1_R1165_U152 , P1_R1165_U153 , P1_R1165_U154 , P1_R1165_U155;
wire P1_R1165_U156 , P1_R1165_U157 , P1_R1165_U158 , P1_R1165_U159 , P1_R1165_U160 , P1_R1165_U161 , P1_R1165_U162 , P1_R1165_U163 , P1_R1165_U164 , P1_R1165_U165;
wire P1_R1165_U166 , P1_R1165_U167 , P1_R1165_U168 , P1_R1165_U169 , P1_R1165_U170 , P1_R1165_U171 , P1_R1165_U172 , P1_R1165_U173 , P1_R1165_U174 , P1_R1165_U175;
wire P1_R1165_U176 , P1_R1165_U177 , P1_R1165_U178 , P1_R1165_U179 , P1_R1165_U180 , P1_R1165_U181 , P1_R1165_U182 , P1_R1165_U183 , P1_R1165_U184 , P1_R1165_U185;
wire P1_R1165_U186 , P1_R1165_U187 , P1_R1165_U188 , P1_R1165_U189 , P1_R1165_U190 , P1_R1165_U191 , P1_R1165_U192 , P1_R1165_U193 , P1_R1165_U194 , P1_R1165_U195;
wire P1_R1165_U196 , P1_R1165_U197 , P1_R1165_U198 , P1_R1165_U199 , P1_R1165_U200 , P1_R1165_U201 , P1_R1165_U202 , P1_R1165_U203 , P1_R1165_U204 , P1_R1165_U205;
wire P1_R1165_U206 , P1_R1165_U207 , P1_R1165_U208 , P1_R1165_U209 , P1_R1165_U210 , P1_R1165_U211 , P1_R1165_U212 , P1_R1165_U213 , P1_R1165_U214 , P1_R1165_U215;
wire P1_R1165_U216 , P1_R1165_U217 , P1_R1165_U218 , P1_R1165_U219 , P1_R1165_U220 , P1_R1165_U221 , P1_R1165_U222 , P1_R1165_U223 , P1_R1165_U224 , P1_R1165_U225;
wire P1_R1165_U226 , P1_R1165_U227 , P1_R1165_U228 , P1_R1165_U229 , P1_R1165_U230 , P1_R1165_U231 , P1_R1165_U232 , P1_R1165_U233 , P1_R1165_U234 , P1_R1165_U235;
wire P1_R1165_U236 , P1_R1165_U237 , P1_R1165_U238 , P1_R1165_U239 , P1_R1165_U240 , P1_R1165_U241 , P1_R1165_U242 , P1_R1165_U243 , P1_R1165_U244 , P1_R1165_U245;
wire P1_R1165_U246 , P1_R1165_U247 , P1_R1165_U248 , P1_R1165_U249 , P1_R1165_U250 , P1_R1165_U251 , P1_R1165_U252 , P1_R1165_U253 , P1_R1165_U254 , P1_R1165_U255;
wire P1_R1165_U256 , P1_R1165_U257 , P1_R1165_U258 , P1_R1165_U259 , P1_R1165_U260 , P1_R1165_U261 , P1_R1165_U262 , P1_R1165_U263 , P1_R1165_U264 , P1_R1165_U265;
wire P1_R1165_U266 , P1_R1165_U267 , P1_R1165_U268 , P1_R1165_U269 , P1_R1165_U270 , P1_R1165_U271 , P1_R1165_U272 , P1_R1165_U273 , P1_R1165_U274 , P1_R1165_U275;
wire P1_R1165_U276 , P1_R1165_U277 , P1_R1165_U278 , P1_R1165_U279 , P1_R1165_U280 , P1_R1165_U281 , P1_R1165_U282 , P1_R1165_U283 , P1_R1165_U284 , P1_R1165_U285;
wire P1_R1165_U286 , P1_R1165_U287 , P1_R1165_U288 , P1_R1165_U289 , P1_R1165_U290 , P1_R1165_U291 , P1_R1165_U292 , P1_R1165_U293 , P1_R1165_U294 , P1_R1165_U295;
wire P1_R1165_U296 , P1_R1165_U297 , P1_R1165_U298 , P1_R1165_U299 , P1_R1165_U300 , P1_R1165_U301 , P1_R1165_U302 , P1_R1165_U303 , P1_R1165_U304 , P1_R1165_U305;
wire P1_R1165_U306 , P1_R1165_U307 , P1_R1165_U308 , P1_R1165_U309 , P1_R1165_U310 , P1_R1165_U311 , P1_R1165_U312 , P1_R1165_U313 , P1_R1165_U314 , P1_R1165_U315;
wire P1_R1165_U316 , P1_R1165_U317 , P1_R1165_U318 , P1_R1165_U319 , P1_R1165_U320 , P1_R1165_U321 , P1_R1165_U322 , P1_R1165_U323 , P1_R1165_U324 , P1_R1165_U325;
wire P1_R1165_U326 , P1_R1165_U327 , P1_R1165_U328 , P1_R1165_U329 , P1_R1165_U330 , P1_R1165_U331 , P1_R1165_U332 , P1_R1165_U333 , P1_R1165_U334 , P1_R1165_U335;
wire P1_R1165_U336 , P1_R1165_U337 , P1_R1165_U338 , P1_R1165_U339 , P1_R1165_U340 , P1_R1165_U341 , P1_R1165_U342 , P1_R1165_U343 , P1_R1165_U344 , P1_R1165_U345;
wire P1_R1165_U346 , P1_R1165_U347 , P1_R1165_U348 , P1_R1165_U349 , P1_R1165_U350 , P1_R1165_U351 , P1_R1165_U352 , P1_R1165_U353 , P1_R1165_U354 , P1_R1165_U355;
wire P1_R1165_U356 , P1_R1165_U357 , P1_R1165_U358 , P1_R1165_U359 , P1_R1165_U360 , P1_R1165_U361 , P1_R1165_U362 , P1_R1165_U363 , P1_R1165_U364 , P1_R1165_U365;
wire P1_R1165_U366 , P1_R1165_U367 , P1_R1165_U368 , P1_R1165_U369 , P1_R1165_U370 , P1_R1165_U371 , P1_R1165_U372 , P1_R1165_U373 , P1_R1165_U374 , P1_R1165_U375;
wire P1_R1165_U376 , P1_R1165_U377 , P1_R1165_U378 , P1_R1165_U379 , P1_R1165_U380 , P1_R1165_U381 , P1_R1165_U382 , P1_R1165_U383 , P1_R1165_U384 , P1_R1165_U385;
wire P1_R1165_U386 , P1_R1165_U387 , P1_R1165_U388 , P1_R1165_U389 , P1_R1165_U390 , P1_R1165_U391 , P1_R1165_U392 , P1_R1165_U393 , P1_R1165_U394 , P1_R1165_U395;
wire P1_R1165_U396 , P1_R1165_U397 , P1_R1165_U398 , P1_R1165_U399 , P1_R1165_U400 , P1_R1165_U401 , P1_R1165_U402 , P1_R1165_U403 , P1_R1165_U404 , P1_R1165_U405;
wire P1_R1165_U406 , P1_R1165_U407 , P1_R1165_U408 , P1_R1165_U409 , P1_R1165_U410 , P1_R1165_U411 , P1_R1165_U412 , P1_R1165_U413 , P1_R1165_U414 , P1_R1165_U415;
wire P1_R1165_U416 , P1_R1165_U417 , P1_R1165_U418 , P1_R1165_U419 , P1_R1165_U420 , P1_R1165_U421 , P1_R1165_U422 , P1_R1165_U423 , P1_R1165_U424 , P1_R1165_U425;
wire P1_R1165_U426 , P1_R1165_U427 , P1_R1165_U428 , P1_R1165_U429 , P1_R1165_U430 , P1_R1165_U431 , P1_R1165_U432 , P1_R1165_U433 , P1_R1165_U434 , P1_R1165_U435;
wire P1_R1165_U436 , P1_R1165_U437 , P1_R1165_U438 , P1_R1165_U439 , P1_R1165_U440 , P1_R1165_U441 , P1_R1165_U442 , P1_R1165_U443 , P1_R1165_U444 , P1_R1165_U445;
wire P1_R1165_U446 , P1_R1165_U447 , P1_R1165_U448 , P1_R1165_U449 , P1_R1165_U450 , P1_R1165_U451 , P1_R1165_U452 , P1_R1165_U453 , P1_R1165_U454 , P1_R1165_U455;
wire P1_R1165_U456 , P1_R1165_U457 , P1_R1165_U458 , P1_R1165_U459 , P1_R1165_U460 , P1_R1165_U461 , P1_R1165_U462 , P1_R1165_U463 , P1_R1165_U464 , P1_R1165_U465;
wire P1_R1165_U466 , P1_R1165_U467 , P1_R1165_U468 , P1_R1165_U469 , P1_R1165_U470 , P1_R1165_U471 , P1_R1165_U472 , P1_R1165_U473 , P1_R1165_U474 , P1_R1165_U475;
wire P1_R1165_U476 , P1_R1165_U477 , P1_R1165_U478 , P1_R1165_U479 , P1_R1165_U480 , P1_R1165_U481 , P1_R1165_U482 , P1_R1165_U483 , P1_R1165_U484 , P1_R1165_U485;
wire P1_R1165_U486 , P1_R1165_U487 , P1_R1165_U488 , P1_R1165_U489 , P1_R1165_U490 , P1_R1165_U491 , P1_R1165_U492 , P1_R1165_U493 , P1_R1165_U494 , P1_R1165_U495;
wire P1_R1165_U496 , P1_R1165_U497 , P1_R1165_U498 , P1_R1165_U499 , P1_R1165_U500 , P1_R1165_U501 , P1_R1165_U502 , P1_R1165_U503 , P1_R1165_U504 , P1_R1165_U505;
wire P1_R1165_U506 , P1_R1165_U507 , P1_R1165_U508 , P1_R1165_U509 , P1_R1165_U510 , P1_R1165_U511 , P1_R1165_U512 , P1_R1165_U513 , P1_R1165_U514 , P1_R1165_U515;
wire P1_R1165_U516 , P1_R1165_U517 , P1_R1165_U518 , P1_R1165_U519 , P1_R1165_U520 , P1_R1165_U521 , P1_R1165_U522 , P1_R1165_U523 , P1_R1165_U524 , P1_R1165_U525;
wire P1_R1165_U526 , P1_R1165_U527 , P1_R1165_U528 , P1_R1165_U529 , P1_R1165_U530 , P1_R1165_U531 , P1_R1165_U532 , P1_R1165_U533 , P1_R1165_U534 , P1_R1165_U535;
wire P1_R1165_U536 , P1_R1165_U537 , P1_R1165_U538 , P1_R1165_U539 , P1_R1165_U540 , P1_R1165_U541 , P1_R1165_U542 , P1_R1165_U543 , P1_R1165_U544 , P1_R1165_U545;
wire P1_R1165_U546 , P1_R1165_U547 , P1_R1165_U548 , P1_R1165_U549 , P1_R1165_U550 , P1_R1165_U551 , P1_R1165_U552 , P1_R1165_U553 , P1_R1165_U554 , P1_R1165_U555;
wire P1_R1165_U556 , P1_R1165_U557 , P1_R1165_U558 , P1_R1165_U559 , P1_R1165_U560 , P1_R1165_U561 , P1_R1165_U562 , P1_R1165_U563 , P1_R1165_U564 , P1_R1165_U565;
wire P1_R1165_U566 , P1_R1165_U567 , P1_R1165_U568 , P1_R1165_U569 , P1_R1165_U570 , P1_R1165_U571 , P1_R1165_U572 , P1_R1165_U573 , P1_R1165_U574 , P1_R1165_U575;
wire P1_R1165_U576 , P1_R1165_U577 , P1_R1165_U578 , P1_R1165_U579 , P1_R1165_U580 , P1_R1165_U581 , P1_R1165_U582 , P1_R1165_U583 , P1_R1165_U584 , P1_R1165_U585;
wire P1_R1165_U586 , P1_R1165_U587 , P1_R1165_U588 , P1_R1165_U589 , P1_R1165_U590 , P1_R1165_U591 , P1_R1165_U592 , P1_R1165_U593 , P1_R1165_U594 , P1_R1165_U595;
wire P1_R1150_U6 , P1_R1150_U7 , P1_R1150_U8 , P1_R1150_U9 , P1_R1150_U10 , P1_R1150_U11 , P1_R1150_U12 , P1_R1150_U13 , P1_R1150_U14 , P1_R1150_U15;
wire P1_R1150_U16 , P1_R1150_U17 , P1_R1150_U18 , P1_R1150_U19 , P1_R1150_U20 , P1_R1150_U21 , P1_R1150_U22 , P1_R1150_U23 , P1_R1150_U24 , P1_R1150_U25;
wire P1_R1150_U26 , P1_R1150_U27 , P1_R1150_U28 , P1_R1150_U29 , P1_R1150_U30 , P1_R1150_U31 , P1_R1150_U32 , P1_R1150_U33 , P1_R1150_U34 , P1_R1150_U35;
wire P1_R1150_U36 , P1_R1150_U37 , P1_R1150_U38 , P1_R1150_U39 , P1_R1150_U40 , P1_R1150_U41 , P1_R1150_U42 , P1_R1150_U43 , P1_R1150_U44 , P1_R1150_U45;
wire P1_R1150_U46 , P1_R1150_U47 , P1_R1150_U48 , P1_R1150_U49 , P1_R1150_U50 , P1_R1150_U51 , P1_R1150_U52 , P1_R1150_U53 , P1_R1150_U54 , P1_R1150_U55;
wire P1_R1150_U56 , P1_R1150_U57 , P1_R1150_U58 , P1_R1150_U59 , P1_R1150_U60 , P1_R1150_U61 , P1_R1150_U62 , P1_R1150_U63 , P1_R1150_U64 , P1_R1150_U65;
wire P1_R1150_U66 , P1_R1150_U67 , P1_R1150_U68 , P1_R1150_U69 , P1_R1150_U70 , P1_R1150_U71 , P1_R1150_U72 , P1_R1150_U73 , P1_R1150_U74 , P1_R1150_U75;
wire P1_R1150_U76 , P1_R1150_U77 , P1_R1150_U78 , P1_R1150_U79 , P1_R1150_U80 , P1_R1150_U81 , P1_R1150_U82 , P1_R1150_U83 , P1_R1150_U84 , P1_R1150_U85;
wire P1_R1150_U86 , P1_R1150_U87 , P1_R1150_U88 , P1_R1150_U89 , P1_R1150_U90 , P1_R1150_U91 , P1_R1150_U92 , P1_R1150_U93 , P1_R1150_U94 , P1_R1150_U95;
wire P1_R1150_U96 , P1_R1150_U97 , P1_R1150_U98 , P1_R1150_U99 , P1_R1150_U100 , P1_R1150_U101 , P1_R1150_U102 , P1_R1150_U103 , P1_R1150_U104 , P1_R1150_U105;
wire P1_R1150_U106 , P1_R1150_U107 , P1_R1150_U108 , P1_R1150_U109 , P1_R1150_U110 , P1_R1150_U111 , P1_R1150_U112 , P1_R1150_U113 , P1_R1150_U114 , P1_R1150_U115;
wire P1_R1150_U116 , P1_R1150_U117 , P1_R1150_U118 , P1_R1150_U119 , P1_R1150_U120 , P1_R1150_U121 , P1_R1150_U122 , P1_R1150_U123 , P1_R1150_U124 , P1_R1150_U125;
wire P1_R1150_U126 , P1_R1150_U127 , P1_R1150_U128 , P1_R1150_U129 , P1_R1150_U130 , P1_R1150_U131 , P1_R1150_U132 , P1_R1150_U133 , P1_R1150_U134 , P1_R1150_U135;
wire P1_R1150_U136 , P1_R1150_U137 , P1_R1150_U138 , P1_R1150_U139 , P1_R1150_U140 , P1_R1150_U141 , P1_R1150_U142 , P1_R1150_U143 , P1_R1150_U144 , P1_R1150_U145;
wire P1_R1150_U146 , P1_R1150_U147 , P1_R1150_U148 , P1_R1150_U149 , P1_R1150_U150 , P1_R1150_U151 , P1_R1150_U152 , P1_R1150_U153 , P1_R1150_U154 , P1_R1150_U155;
wire P1_R1150_U156 , P1_R1150_U157 , P1_R1150_U158 , P1_R1150_U159 , P1_R1150_U160 , P1_R1150_U161 , P1_R1150_U162 , P1_R1150_U163 , P1_R1150_U164 , P1_R1150_U165;
wire P1_R1150_U166 , P1_R1150_U167 , P1_R1150_U168 , P1_R1150_U169 , P1_R1150_U170 , P1_R1150_U171 , P1_R1150_U172 , P1_R1150_U173 , P1_R1150_U174 , P1_R1150_U175;
wire P1_R1150_U176 , P1_R1150_U177 , P1_R1150_U178 , P1_R1150_U179 , P1_R1150_U180 , P1_R1150_U181 , P1_R1150_U182 , P1_R1150_U183 , P1_R1150_U184 , P1_R1150_U185;
wire P1_R1150_U186 , P1_R1150_U187 , P1_R1150_U188 , P1_R1150_U189 , P1_R1150_U190 , P1_R1150_U191 , P1_R1150_U192 , P1_R1150_U193 , P1_R1150_U194 , P1_R1150_U195;
wire P1_R1150_U196 , P1_R1150_U197 , P1_R1150_U198 , P1_R1150_U199 , P1_R1150_U200 , P1_R1150_U201 , P1_R1150_U202 , P1_R1150_U203 , P1_R1150_U204 , P1_R1150_U205;
wire P1_R1150_U206 , P1_R1150_U207 , P1_R1150_U208 , P1_R1150_U209 , P1_R1150_U210 , P1_R1150_U211 , P1_R1150_U212 , P1_R1150_U213 , P1_R1150_U214 , P1_R1150_U215;
wire P1_R1150_U216 , P1_R1150_U217 , P1_R1150_U218 , P1_R1150_U219 , P1_R1150_U220 , P1_R1150_U221 , P1_R1150_U222 , P1_R1150_U223 , P1_R1150_U224 , P1_R1150_U225;
wire P1_R1150_U226 , P1_R1150_U227 , P1_R1150_U228 , P1_R1150_U229 , P1_R1150_U230 , P1_R1150_U231 , P1_R1150_U232 , P1_R1150_U233 , P1_R1150_U234 , P1_R1150_U235;
wire P1_R1150_U236 , P1_R1150_U237 , P1_R1150_U238 , P1_R1150_U239 , P1_R1150_U240 , P1_R1150_U241 , P1_R1150_U242 , P1_R1150_U243 , P1_R1150_U244 , P1_R1150_U245;
wire P1_R1150_U246 , P1_R1150_U247 , P1_R1150_U248 , P1_R1150_U249 , P1_R1150_U250 , P1_R1150_U251 , P1_R1150_U252 , P1_R1150_U253 , P1_R1150_U254 , P1_R1150_U255;
wire P1_R1150_U256 , P1_R1150_U257 , P1_R1150_U258 , P1_R1150_U259 , P1_R1150_U260 , P1_R1150_U261 , P1_R1150_U262 , P1_R1150_U263 , P1_R1150_U264 , P1_R1150_U265;
wire P1_R1150_U266 , P1_R1150_U267 , P1_R1150_U268 , P1_R1150_U269 , P1_R1150_U270 , P1_R1150_U271 , P1_R1150_U272 , P1_R1150_U273 , P1_R1150_U274 , P1_R1150_U275;
wire P1_R1150_U276 , P1_R1150_U277 , P1_R1150_U278 , P1_R1150_U279 , P1_R1150_U280 , P1_R1150_U281 , P1_R1150_U282 , P1_R1150_U283 , P1_R1150_U284 , P1_R1150_U285;
wire P1_R1150_U286 , P1_R1150_U287 , P1_R1150_U288 , P1_R1150_U289 , P1_R1150_U290 , P1_R1150_U291 , P1_R1150_U292 , P1_R1150_U293 , P1_R1150_U294 , P1_R1150_U295;
wire P1_R1150_U296 , P1_R1150_U297 , P1_R1150_U298 , P1_R1150_U299 , P1_R1150_U300 , P1_R1150_U301 , P1_R1150_U302 , P1_R1150_U303 , P1_R1150_U304 , P1_R1150_U305;
wire P1_R1150_U306 , P1_R1150_U307 , P1_R1150_U308 , P1_R1150_U309 , P1_R1150_U310 , P1_R1150_U311 , P1_R1150_U312 , P1_R1150_U313 , P1_R1150_U314 , P1_R1150_U315;
wire P1_R1150_U316 , P1_R1150_U317 , P1_R1150_U318 , P1_R1150_U319 , P1_R1150_U320 , P1_R1150_U321 , P1_R1150_U322 , P1_R1150_U323 , P1_R1150_U324 , P1_R1150_U325;
wire P1_R1150_U326 , P1_R1150_U327 , P1_R1150_U328 , P1_R1150_U329 , P1_R1150_U330 , P1_R1150_U331 , P1_R1150_U332 , P1_R1150_U333 , P1_R1150_U334 , P1_R1150_U335;
wire P1_R1150_U336 , P1_R1150_U337 , P1_R1150_U338 , P1_R1150_U339 , P1_R1150_U340 , P1_R1150_U341 , P1_R1150_U342 , P1_R1150_U343 , P1_R1150_U344 , P1_R1150_U345;
wire P1_R1150_U346 , P1_R1150_U347 , P1_R1150_U348 , P1_R1150_U349 , P1_R1150_U350 , P1_R1150_U351 , P1_R1150_U352 , P1_R1150_U353 , P1_R1150_U354 , P1_R1150_U355;
wire P1_R1150_U356 , P1_R1150_U357 , P1_R1150_U358 , P1_R1150_U359 , P1_R1150_U360 , P1_R1150_U361 , P1_R1150_U362 , P1_R1150_U363 , P1_R1150_U364 , P1_R1150_U365;
wire P1_R1150_U366 , P1_R1150_U367 , P1_R1150_U368 , P1_R1150_U369 , P1_R1150_U370 , P1_R1150_U371 , P1_R1150_U372 , P1_R1150_U373 , P1_R1150_U374 , P1_R1150_U375;
wire P1_R1150_U376 , P1_R1150_U377 , P1_R1150_U378 , P1_R1150_U379 , P1_R1150_U380 , P1_R1150_U381 , P1_R1150_U382 , P1_R1150_U383 , P1_R1150_U384 , P1_R1150_U385;
wire P1_R1150_U386 , P1_R1150_U387 , P1_R1150_U388 , P1_R1150_U389 , P1_R1150_U390 , P1_R1150_U391 , P1_R1150_U392 , P1_R1150_U393 , P1_R1150_U394 , P1_R1150_U395;
wire P1_R1150_U396 , P1_R1150_U397 , P1_R1150_U398 , P1_R1150_U399 , P1_R1150_U400 , P1_R1150_U401 , P1_R1150_U402 , P1_R1150_U403 , P1_R1150_U404 , P1_R1150_U405;
wire P1_R1150_U406 , P1_R1150_U407 , P1_R1150_U408 , P1_R1150_U409 , P1_R1150_U410 , P1_R1150_U411 , P1_R1150_U412 , P1_R1150_U413 , P1_R1150_U414 , P1_R1150_U415;
wire P1_R1150_U416 , P1_R1150_U417 , P1_R1150_U418 , P1_R1150_U419 , P1_R1150_U420 , P1_R1150_U421 , P1_R1150_U422 , P1_R1150_U423 , P1_R1150_U424 , P1_R1150_U425;
wire P1_R1150_U426 , P1_R1150_U427 , P1_R1150_U428 , P1_R1150_U429 , P1_R1150_U430 , P1_R1150_U431 , P1_R1150_U432 , P1_R1150_U433 , P1_R1150_U434 , P1_R1150_U435;
wire P1_R1150_U436 , P1_R1150_U437 , P1_R1150_U438 , P1_R1150_U439 , P1_R1150_U440 , P1_R1150_U441 , P1_R1150_U442 , P1_R1150_U443 , P1_R1150_U444 , P1_R1150_U445;
wire P1_R1150_U446 , P1_R1150_U447 , P1_R1150_U448 , P1_R1150_U449 , P1_R1150_U450 , P1_R1150_U451 , P1_R1150_U452 , P1_R1150_U453 , P1_R1150_U454 , P1_R1150_U455;
wire P1_R1150_U456 , P1_R1150_U457 , P1_R1150_U458 , P1_R1150_U459 , P1_R1150_U460 , P1_R1150_U461 , P1_R1150_U462 , P1_R1150_U463 , P1_R1150_U464 , P1_R1150_U465;
wire P1_R1150_U466 , P1_R1150_U467 , P1_R1150_U468 , P1_R1150_U469 , P1_R1150_U470 , P1_R1150_U471 , P1_R1150_U472 , P1_R1150_U473 , P1_R1150_U474 , P1_R1150_U475;
wire P1_R1150_U476 , P1_R1192_U6 , P1_R1192_U7 , P1_R1192_U8 , P1_R1192_U9 , P1_R1192_U10 , P1_R1192_U11 , P1_R1192_U12 , P1_R1192_U13 , P1_R1192_U14;
wire P1_R1192_U15 , P1_R1192_U16 , P1_R1192_U17 , P1_R1192_U18 , P1_R1192_U19 , P1_R1192_U20 , P1_R1192_U21 , P1_R1192_U22 , P1_R1192_U23 , P1_R1192_U24;
wire P1_R1192_U25 , P1_R1192_U26 , P1_R1192_U27 , P1_R1192_U28 , P1_R1192_U29 , P1_R1192_U30 , P1_R1192_U31 , P1_R1192_U32 , P1_R1192_U33 , P1_R1192_U34;
wire P1_R1192_U35 , P1_R1192_U36 , P1_R1192_U37 , P1_R1192_U38 , P1_R1192_U39 , P1_R1192_U40 , P1_R1192_U41 , P1_R1192_U42 , P1_R1192_U43 , P1_R1192_U44;
wire P1_R1192_U45 , P1_R1192_U46 , P1_R1192_U47 , P1_R1192_U48 , P1_R1192_U49 , P1_R1192_U50 , P1_R1192_U51 , P1_R1192_U52 , P1_R1192_U53 , P1_R1192_U54;
wire P1_R1192_U55 , P1_R1192_U56 , P1_R1192_U57 , P1_R1192_U58 , P1_R1192_U59 , P1_R1192_U60 , P1_R1192_U61 , P1_R1192_U62 , P1_R1192_U63 , P1_R1192_U64;
wire P1_R1192_U65 , P1_R1192_U66 , P1_R1192_U67 , P1_R1192_U68 , P1_R1192_U69 , P1_R1192_U70 , P1_R1192_U71 , P1_R1192_U72 , P1_R1192_U73 , P1_R1192_U74;
wire P1_R1192_U75 , P1_R1192_U76 , P1_R1192_U77 , P1_R1192_U78 , P1_R1192_U79 , P1_R1192_U80 , P1_R1192_U81 , P1_R1192_U82 , P1_R1192_U83 , P1_R1192_U84;
wire P1_R1192_U85 , P1_R1192_U86 , P1_R1192_U87 , P1_R1192_U88 , P1_R1192_U89 , P1_R1192_U90 , P1_R1192_U91 , P1_R1192_U92 , P1_R1192_U93 , P1_R1192_U94;
wire P1_R1192_U95 , P1_R1192_U96 , P1_R1192_U97 , P1_R1192_U98 , P1_R1192_U99 , P1_R1192_U100 , P1_R1192_U101 , P1_R1192_U102 , P1_R1192_U103 , P1_R1192_U104;
wire P1_R1192_U105 , P1_R1192_U106 , P1_R1192_U107 , P1_R1192_U108 , P1_R1192_U109 , P1_R1192_U110 , P1_R1192_U111 , P1_R1192_U112 , P1_R1192_U113 , P1_R1192_U114;
wire P1_R1192_U115 , P1_R1192_U116 , P1_R1192_U117 , P1_R1192_U118 , P1_R1192_U119 , P1_R1192_U120 , P1_R1192_U121 , P1_R1192_U122 , P1_R1192_U123 , P1_R1192_U124;
wire P1_R1192_U125 , P1_R1192_U126 , P1_R1192_U127 , P1_R1192_U128 , P1_R1192_U129 , P1_R1192_U130 , P1_R1192_U131 , P1_R1192_U132 , P1_R1192_U133 , P1_R1192_U134;
wire P1_R1192_U135 , P1_R1192_U136 , P1_R1192_U137 , P1_R1192_U138 , P1_R1192_U139 , P1_R1192_U140 , P1_R1192_U141 , P1_R1192_U142 , P1_R1192_U143 , P1_R1192_U144;
wire P1_R1192_U145 , P1_R1192_U146 , P1_R1192_U147 , P1_R1192_U148 , P1_R1192_U149 , P1_R1192_U150 , P1_R1192_U151 , P1_R1192_U152 , P1_R1192_U153 , P1_R1192_U154;
wire P1_R1192_U155 , P1_R1192_U156 , P1_R1192_U157 , P1_R1192_U158 , P1_R1192_U159 , P1_R1192_U160 , P1_R1192_U161 , P1_R1192_U162 , P1_R1192_U163 , P1_R1192_U164;
wire P1_R1192_U165 , P1_R1192_U166 , P1_R1192_U167 , P1_R1192_U168 , P1_R1192_U169 , P1_R1192_U170 , P1_R1192_U171 , P1_R1192_U172 , P1_R1192_U173 , P1_R1192_U174;
wire P1_R1192_U175 , P1_R1192_U176 , P1_R1192_U177 , P1_R1192_U178 , P1_R1192_U179 , P1_R1192_U180 , P1_R1192_U181 , P1_R1192_U182 , P1_R1192_U183 , P1_R1192_U184;
wire P1_R1192_U185 , P1_R1192_U186 , P1_R1192_U187 , P1_R1192_U188 , P1_R1192_U189 , P1_R1192_U190 , P1_R1192_U191 , P1_R1192_U192 , P1_R1192_U193 , P1_R1192_U194;
wire P1_R1192_U195 , P1_R1192_U196 , P1_R1192_U197 , P1_R1192_U198 , P1_R1192_U199 , P1_R1192_U200 , P1_R1192_U201 , P1_R1192_U202 , P1_R1192_U203 , P1_R1192_U204;
wire P1_R1192_U205 , P1_R1192_U206 , P1_R1192_U207 , P1_R1192_U208 , P1_R1192_U209 , P1_R1192_U210 , P1_R1192_U211 , P1_R1192_U212 , P1_R1192_U213 , P1_R1192_U214;
wire P1_R1192_U215 , P1_R1192_U216 , P1_R1192_U217 , P1_R1192_U218 , P1_R1192_U219 , P1_R1192_U220 , P1_R1192_U221 , P1_R1192_U222 , P1_R1192_U223 , P1_R1192_U224;
wire P1_R1192_U225 , P1_R1192_U226 , P1_R1192_U227 , P1_R1192_U228 , P1_R1192_U229 , P1_R1192_U230 , P1_R1192_U231 , P1_R1192_U232 , P1_R1192_U233 , P1_R1192_U234;
wire P1_R1192_U235 , P1_R1192_U236 , P1_R1192_U237 , P1_R1192_U238 , P1_R1192_U239 , P1_R1192_U240 , P1_R1192_U241 , P1_R1192_U242 , P1_R1192_U243 , P1_R1192_U244;
wire P1_R1192_U245 , P1_R1192_U246 , P1_R1192_U247 , P1_R1192_U248 , P1_R1192_U249 , P1_R1192_U250 , P1_R1192_U251 , P1_R1192_U252 , P1_R1192_U253 , P1_R1192_U254;
wire P1_R1192_U255 , P1_R1192_U256 , P1_R1192_U257 , P1_R1192_U258 , P1_R1192_U259 , P1_R1192_U260 , P1_R1192_U261 , P1_R1192_U262 , P1_R1192_U263 , P1_R1192_U264;
wire P1_R1192_U265 , P1_R1192_U266 , P1_R1192_U267 , P1_R1192_U268 , P1_R1192_U269 , P1_R1192_U270 , P1_R1192_U271 , P1_R1192_U272 , P1_R1192_U273 , P1_R1192_U274;
wire P1_R1192_U275 , P1_R1192_U276 , P1_R1192_U277 , P1_R1192_U278 , P1_R1192_U279 , P1_R1192_U280 , P1_R1192_U281 , P1_R1192_U282 , P1_R1192_U283 , P1_R1192_U284;
wire P1_R1192_U285 , P1_R1192_U286 , P1_R1192_U287 , P1_R1192_U288 , P1_R1192_U289 , P1_R1192_U290 , P1_R1192_U291 , P1_R1192_U292 , P1_R1192_U293 , P1_R1192_U294;
wire P1_R1192_U295 , P1_R1192_U296 , P1_R1192_U297 , P1_R1192_U298 , P1_R1192_U299 , P1_R1192_U300 , P1_R1192_U301 , P1_R1192_U302 , P1_R1192_U303 , P1_R1192_U304;
wire P1_R1192_U305 , P1_R1192_U306 , P1_R1192_U307 , P1_R1192_U308 , P1_R1192_U309 , P1_R1192_U310 , P1_R1192_U311 , P1_R1192_U312 , P1_R1192_U313 , P1_R1192_U314;
wire P1_R1192_U315 , P1_R1192_U316 , P1_R1192_U317 , P1_R1192_U318 , P1_R1192_U319 , P1_R1192_U320 , P1_R1192_U321 , P1_R1192_U322 , P1_R1192_U323 , P1_R1192_U324;
wire P1_R1192_U325 , P1_R1192_U326 , P1_R1192_U327 , P1_R1192_U328 , P1_R1192_U329 , P1_R1192_U330 , P1_R1192_U331 , P1_R1192_U332 , P1_R1192_U333 , P1_R1192_U334;
wire P1_R1192_U335 , P1_R1192_U336 , P1_R1192_U337 , P1_R1192_U338 , P1_R1192_U339 , P1_R1192_U340 , P1_R1192_U341 , P1_R1192_U342 , P1_R1192_U343 , P1_R1192_U344;
wire P1_R1192_U345 , P1_R1192_U346 , P1_R1192_U347 , P1_R1192_U348 , P1_R1192_U349 , P1_R1192_U350 , P1_R1192_U351 , P1_R1192_U352 , P1_R1192_U353 , P1_R1192_U354;
wire P1_R1192_U355 , P1_R1192_U356 , P1_R1192_U357 , P1_R1192_U358 , P1_R1192_U359 , P1_R1192_U360 , P1_R1192_U361 , P1_R1192_U362 , P1_R1192_U363 , P1_R1192_U364;
wire P1_R1192_U365 , P1_R1192_U366 , P1_R1192_U367 , P1_R1192_U368 , P1_R1192_U369 , P1_R1192_U370 , P1_R1192_U371 , P1_R1192_U372 , P1_R1192_U373 , P1_R1192_U374;
wire P1_R1192_U375 , P1_R1192_U376 , P1_R1192_U377 , P1_R1192_U378 , P1_R1192_U379 , P1_R1192_U380 , P1_R1192_U381 , P1_R1192_U382 , P1_R1192_U383 , P1_R1192_U384;
wire P1_R1192_U385 , P1_R1192_U386 , P1_R1192_U387 , P1_R1192_U388 , P1_R1192_U389 , P1_R1192_U390 , P1_R1192_U391 , P1_R1192_U392 , P1_R1192_U393 , P1_R1192_U394;
wire P1_R1192_U395 , P1_R1192_U396 , P1_R1192_U397 , P1_R1192_U398 , P1_R1192_U399 , P1_R1192_U400 , P1_R1192_U401 , P1_R1192_U402 , P1_R1192_U403 , P1_R1192_U404;
wire P1_R1192_U405 , P1_R1192_U406 , P1_R1192_U407 , P1_R1192_U408 , P1_R1192_U409 , P1_R1192_U410 , P1_R1192_U411 , P1_R1192_U412 , P1_R1192_U413 , P1_R1192_U414;
wire P1_R1192_U415 , P1_R1192_U416 , P1_R1192_U417 , P1_R1192_U418 , P1_R1192_U419 , P1_R1192_U420 , P1_R1192_U421 , P1_R1192_U422 , P1_R1192_U423 , P1_R1192_U424;
wire P1_R1192_U425 , P1_R1192_U426 , P1_R1192_U427 , P1_R1192_U428 , P1_R1192_U429 , P1_R1192_U430 , P1_R1192_U431 , P1_R1192_U432 , P1_R1192_U433 , P1_R1192_U434;
wire P1_R1192_U435 , P1_R1192_U436 , P1_R1192_U437 , P1_R1192_U438 , P1_R1192_U439 , P1_R1192_U440 , P1_R1192_U441 , P1_R1192_U442 , P1_R1192_U443 , P1_R1192_U444;
wire P1_R1192_U445 , P1_R1192_U446 , P1_R1192_U447 , P1_R1192_U448 , P1_R1192_U449 , P1_R1192_U450 , P1_R1192_U451 , P1_R1192_U452 , P1_R1192_U453 , P1_R1192_U454;
wire P1_R1192_U455 , P1_R1192_U456 , P1_R1192_U457 , P1_R1192_U458 , P1_R1192_U459 , P1_R1192_U460 , P1_R1192_U461 , P1_R1192_U462 , P1_R1192_U463 , P1_R1192_U464;
wire P1_R1192_U465 , P1_R1192_U466 , P1_R1192_U467 , P1_R1192_U468 , P1_R1192_U469 , P1_R1192_U470 , P1_R1192_U471 , P1_R1192_U472 , P1_R1192_U473 , P1_R1192_U474;
wire P1_R1192_U475 , P1_R1192_U476 , P1_R1171_U4 , P1_R1171_U5 , P1_R1171_U6 , P1_R1171_U7 , P1_R1171_U8 , P1_R1171_U9 , P1_R1171_U10 , P1_R1171_U11;
wire P1_R1171_U12 , P1_R1171_U13 , P1_R1171_U14 , P1_R1171_U15 , P1_R1171_U16 , P1_R1171_U17 , P1_R1171_U18 , P1_R1171_U19 , P1_R1171_U20 , P1_R1171_U21;
wire P1_R1171_U22 , P1_R1171_U23 , P1_R1171_U24 , P1_R1171_U25 , P1_R1171_U26 , P1_R1171_U27 , P1_R1171_U28 , P1_R1171_U29 , P1_R1171_U30 , P1_R1171_U31;
wire P1_R1171_U32 , P1_R1171_U33 , P1_R1171_U34 , P1_R1171_U35 , P1_R1171_U36 , P1_R1171_U37 , P1_R1171_U38 , P1_R1171_U39 , P1_R1171_U40 , P1_R1171_U41;
wire P1_R1171_U42 , P1_R1171_U43 , P1_R1171_U44 , P1_R1171_U45 , P1_R1171_U46 , P1_R1171_U47 , P1_R1171_U48 , P1_R1171_U49 , P1_R1171_U50 , P1_R1171_U51;
wire P1_R1171_U52 , P1_R1171_U53 , P1_R1171_U54 , P1_R1171_U55 , P1_R1171_U56 , P1_R1171_U57 , P1_R1171_U58 , P1_R1171_U59 , P1_R1171_U60 , P1_R1171_U61;
wire P1_R1171_U62 , P1_R1171_U63 , P1_R1171_U64 , P1_R1171_U65 , P1_R1171_U66 , P1_R1171_U67 , P1_R1171_U68 , P1_R1171_U69 , P1_R1171_U70 , P1_R1171_U71;
wire P1_R1171_U72 , P1_R1171_U73 , P1_R1171_U74 , P1_R1171_U75 , P1_R1171_U76 , P1_R1171_U77 , P1_R1171_U78 , P1_R1171_U79 , P1_R1171_U80 , P1_R1171_U81;
wire P1_R1171_U82 , P1_R1171_U83 , P1_R1171_U84 , P1_R1171_U85 , P1_R1171_U86 , P1_R1171_U87 , P1_R1171_U88 , P1_R1171_U89 , P1_R1171_U90 , P1_R1171_U91;
wire P1_R1171_U92 , P1_R1171_U93 , P1_R1171_U94 , P1_R1171_U95 , P1_R1171_U96 , P1_R1171_U97 , P1_R1171_U98 , P1_R1171_U99 , P1_R1171_U100 , P1_R1171_U101;
wire P1_R1171_U102 , P1_R1171_U103 , P1_R1171_U104 , P1_R1171_U105 , P1_R1171_U106 , P1_R1171_U107 , P1_R1171_U108 , P1_R1171_U109 , P1_R1171_U110 , P1_R1171_U111;
wire P1_R1171_U112 , P1_R1171_U113 , P1_R1171_U114 , P1_R1171_U115 , P1_R1171_U116 , P1_R1171_U117 , P1_R1171_U118 , P1_R1171_U119 , P1_R1171_U120 , P1_R1171_U121;
wire P1_R1171_U122 , P1_R1171_U123 , P1_R1171_U124 , P1_R1171_U125 , P1_R1171_U126 , P1_R1171_U127 , P1_R1171_U128 , P1_R1171_U129 , P1_R1171_U130 , P1_R1171_U131;
wire P1_R1171_U132 , P1_R1171_U133 , P1_R1171_U134 , P1_R1171_U135 , P1_R1171_U136 , P1_R1171_U137 , P1_R1171_U138 , P1_R1171_U139 , P1_R1171_U140 , P1_R1171_U141;
wire P1_R1171_U142 , P1_R1171_U143 , P1_R1171_U144 , P1_R1171_U145 , P1_R1171_U146 , P1_R1171_U147 , P1_R1171_U148 , P1_R1171_U149 , P1_R1171_U150 , P1_R1171_U151;
wire P1_R1171_U152 , P1_R1171_U153 , P1_R1171_U154 , P1_R1171_U155 , P1_R1171_U156 , P1_R1171_U157 , P1_R1171_U158 , P1_R1171_U159 , P1_R1171_U160 , P1_R1171_U161;
wire P1_R1171_U162 , P1_R1171_U163 , P1_R1171_U164 , P1_R1171_U165 , P1_R1171_U166 , P1_R1171_U167 , P1_R1171_U168 , P1_R1171_U169 , P1_R1171_U170 , P1_R1171_U171;
wire P1_R1171_U172 , P1_R1171_U173 , P1_R1171_U174 , P1_R1171_U175 , P1_R1171_U176 , P1_R1171_U177 , P1_R1171_U178 , P1_R1171_U179 , P1_R1171_U180 , P1_R1171_U181;
wire P1_R1171_U182 , P1_R1171_U183 , P1_R1171_U184 , P1_R1171_U185 , P1_R1171_U186 , P1_R1171_U187 , P1_R1171_U188 , P1_R1171_U189 , P1_R1171_U190 , P1_R1171_U191;
wire P1_R1171_U192 , P1_R1171_U193 , P1_R1171_U194 , P1_R1171_U195 , P1_R1171_U196 , P1_R1171_U197 , P1_R1171_U198 , P1_R1171_U199 , P1_R1171_U200 , P1_R1171_U201;
wire P1_R1171_U202 , P1_R1171_U203 , P1_R1171_U204 , P1_R1171_U205 , P1_R1171_U206 , P1_R1171_U207 , P1_R1171_U208 , P1_R1171_U209 , P1_R1171_U210 , P1_R1171_U211;
wire P1_R1171_U212 , P1_R1171_U213 , P1_R1171_U214 , P1_R1171_U215 , P1_R1171_U216 , P1_R1171_U217 , P1_R1171_U218 , P1_R1171_U219 , P1_R1171_U220 , P1_R1171_U221;
wire P1_R1171_U222 , P1_R1171_U223 , P1_R1171_U224 , P1_R1171_U225 , P1_R1171_U226 , P1_R1171_U227 , P1_R1171_U228 , P1_R1171_U229 , P1_R1171_U230 , P1_R1171_U231;
wire P1_R1171_U232 , P1_R1171_U233 , P1_R1171_U234 , P1_R1171_U235 , P1_R1171_U236 , P1_R1171_U237 , P1_R1171_U238 , P1_R1171_U239 , P1_R1171_U240 , P1_R1171_U241;
wire P1_R1171_U242 , P1_R1171_U243 , P1_R1171_U244 , P1_R1171_U245 , P1_R1171_U246 , P1_R1171_U247 , P1_R1171_U248 , P1_R1171_U249 , P1_R1171_U250 , P1_R1171_U251;
wire P1_R1171_U252 , P1_R1171_U253 , P1_R1171_U254 , P1_R1171_U255 , P1_R1171_U256 , P1_R1171_U257 , P1_R1171_U258 , P1_R1171_U259 , P1_R1171_U260 , P1_R1171_U261;
wire P1_R1171_U262 , P1_R1171_U263 , P1_R1171_U264 , P1_R1171_U265 , P1_R1171_U266 , P1_R1171_U267 , P1_R1171_U268 , P1_R1171_U269 , P1_R1171_U270 , P1_R1171_U271;
wire P1_R1171_U272 , P1_R1171_U273 , P1_R1171_U274 , P1_R1171_U275 , P1_R1171_U276 , P1_R1171_U277 , P1_R1171_U278 , P1_R1171_U279 , P1_R1171_U280 , P1_R1171_U281;
wire P1_R1171_U282 , P1_R1171_U283 , P1_R1171_U284 , P1_R1171_U285 , P1_R1171_U286 , P1_R1171_U287 , P1_R1171_U288 , P1_R1171_U289 , P1_R1171_U290 , P1_R1171_U291;
wire P1_R1171_U292 , P1_R1171_U293 , P1_R1171_U294 , P1_R1171_U295 , P1_R1171_U296 , P1_R1171_U297 , P1_R1171_U298 , P1_R1171_U299 , P1_R1171_U300 , P1_R1171_U301;
wire P1_R1171_U302 , P1_R1171_U303 , P1_R1171_U304 , P1_R1171_U305 , P1_R1171_U306 , P1_R1171_U307 , P1_R1171_U308 , P1_R1171_U309 , P1_R1171_U310 , P1_R1171_U311;
wire P1_R1171_U312 , P1_R1171_U313 , P1_R1171_U314 , P1_R1171_U315 , P1_R1171_U316 , P1_R1171_U317 , P1_R1171_U318 , P1_R1171_U319 , P1_R1171_U320 , P1_R1171_U321;
wire P1_R1171_U322 , P1_R1171_U323 , P1_R1171_U324 , P1_R1171_U325 , P1_R1171_U326 , P1_R1171_U327 , P1_R1171_U328 , P1_R1171_U329 , P1_R1171_U330 , P1_R1171_U331;
wire P1_R1171_U332 , P1_R1171_U333 , P1_R1171_U334 , P1_R1171_U335 , P1_R1171_U336 , P1_R1171_U337 , P1_R1171_U338 , P1_R1171_U339 , P1_R1171_U340 , P1_R1171_U341;
wire P1_R1171_U342 , P1_R1171_U343 , P1_R1171_U344 , P1_R1171_U345 , P1_R1171_U346 , P1_R1171_U347 , P1_R1171_U348 , P1_R1171_U349 , P1_R1171_U350 , P1_R1171_U351;
wire P1_R1171_U352 , P1_R1171_U353 , P1_R1171_U354 , P1_R1171_U355 , P1_R1171_U356 , P1_R1171_U357 , P1_R1171_U358 , P1_R1171_U359 , P1_R1171_U360 , P1_R1171_U361;
wire P1_R1171_U362 , P1_R1171_U363 , P1_R1171_U364 , P1_R1171_U365 , P1_R1171_U366 , P1_R1171_U367 , P1_R1171_U368 , P1_R1171_U369 , P1_R1171_U370 , P1_R1171_U371;
wire P1_R1171_U372 , P1_R1171_U373 , P1_R1171_U374 , P1_R1171_U375 , P1_R1171_U376 , P1_R1171_U377 , P1_R1171_U378 , P1_R1171_U379 , P1_R1171_U380 , P1_R1171_U381;
wire P1_R1171_U382 , P1_R1171_U383 , P1_R1171_U384 , P1_R1171_U385 , P1_R1171_U386 , P1_R1171_U387 , P1_R1171_U388 , P1_R1171_U389 , P1_R1171_U390 , P1_R1171_U391;
wire P1_R1171_U392 , P1_R1171_U393 , P1_R1171_U394 , P1_R1171_U395 , P1_R1171_U396 , P1_R1171_U397 , P1_R1171_U398 , P1_R1171_U399 , P1_R1171_U400 , P1_R1171_U401;
wire P1_R1171_U402 , P1_R1171_U403 , P1_R1171_U404 , P1_R1171_U405 , P1_R1171_U406 , P1_R1171_U407 , P1_R1171_U408 , P1_R1171_U409 , P1_R1171_U410 , P1_R1171_U411;
wire P1_R1171_U412 , P1_R1171_U413 , P1_R1171_U414 , P1_R1171_U415 , P1_R1171_U416 , P1_R1171_U417 , P1_R1171_U418 , P1_R1171_U419 , P1_R1171_U420 , P1_R1171_U421;
wire P1_R1171_U422 , P1_R1171_U423 , P1_R1171_U424 , P1_R1171_U425 , P1_R1171_U426 , P1_R1171_U427 , P1_R1171_U428 , P1_R1171_U429 , P1_R1171_U430 , P1_R1171_U431;
wire P1_R1171_U432 , P1_R1171_U433 , P1_R1171_U434 , P1_R1171_U435 , P1_R1171_U436 , P1_R1171_U437 , P1_R1171_U438 , P1_R1171_U439 , P1_R1171_U440 , P1_R1171_U441;
wire P1_R1171_U442 , P1_R1171_U443 , P1_R1171_U444 , P1_R1171_U445 , P1_R1171_U446 , P1_R1171_U447 , P1_R1171_U448 , P1_R1171_U449 , P1_R1171_U450 , P1_R1171_U451;
wire P1_R1171_U452 , P1_R1171_U453 , P1_R1171_U454 , P1_R1171_U455 , P1_R1171_U456 , P1_R1171_U457 , P1_R1171_U458 , P1_R1171_U459 , P1_R1171_U460 , P1_R1171_U461;
wire P1_R1171_U462 , P1_R1171_U463 , P1_R1171_U464 , P1_R1171_U465 , P1_R1171_U466 , P1_R1171_U467 , P1_R1171_U468 , P1_R1171_U469 , P1_R1171_U470 , P1_R1171_U471;
wire P1_R1171_U472 , P1_R1171_U473 , P1_R1171_U474 , P1_R1171_U475 , P1_R1171_U476 , P1_R1171_U477 , P1_R1171_U478 , P1_R1171_U479 , P1_R1171_U480 , P1_R1171_U481;
wire P1_R1171_U482 , P1_R1171_U483 , P1_R1171_U484 , P1_R1171_U485 , P1_R1171_U486 , P1_R1171_U487 , P1_R1171_U488 , P1_R1171_U489 , P1_R1171_U490 , P1_R1171_U491;
wire P1_R1171_U492 , P1_R1171_U493 , P1_R1171_U494 , P1_R1171_U495 , P1_R1171_U496 , P1_R1171_U497 , P1_R1171_U498 , P1_R1171_U499 , P1_R1171_U500 , P1_R1171_U501;
wire P1_R1138_U4 , P1_R1138_U5 , P1_R1138_U6 , P1_R1138_U7 , P1_R1138_U8 , P1_R1138_U9 , P1_R1138_U10 , P1_R1138_U11 , P1_R1138_U12 , P1_R1138_U13;
wire P1_R1138_U14 , P1_R1138_U15 , P1_R1138_U16 , P1_R1138_U17 , P1_R1138_U18 , P1_R1138_U19 , P1_R1138_U20 , P1_R1138_U21 , P1_R1138_U22 , P1_R1138_U23;
wire P1_R1138_U24 , P1_R1138_U25 , P1_R1138_U26 , P1_R1138_U27 , P1_R1138_U28 , P1_R1138_U29 , P1_R1138_U30 , P1_R1138_U31 , P1_R1138_U32 , P1_R1138_U33;
wire P1_R1138_U34 , P1_R1138_U35 , P1_R1138_U36 , P1_R1138_U37 , P1_R1138_U38 , P1_R1138_U39 , P1_R1138_U40 , P1_R1138_U41 , P1_R1138_U42 , P1_R1138_U43;
wire P1_R1138_U44 , P1_R1138_U45 , P1_R1138_U46 , P1_R1138_U47 , P1_R1138_U48 , P1_R1138_U49 , P1_R1138_U50 , P1_R1138_U51 , P1_R1138_U52 , P1_R1138_U53;
wire P1_R1138_U54 , P1_R1138_U55 , P1_R1138_U56 , P1_R1138_U57 , P1_R1138_U58 , P1_R1138_U59 , P1_R1138_U60 , P1_R1138_U61 , P1_R1138_U62 , P1_R1138_U63;
wire P1_R1138_U64 , P1_R1138_U65 , P1_R1138_U66 , P1_R1138_U67 , P1_R1138_U68 , P1_R1138_U69 , P1_R1138_U70 , P1_R1138_U71 , P1_R1138_U72 , P1_R1138_U73;
wire P1_R1138_U74 , P1_R1138_U75 , P1_R1138_U76 , P1_R1138_U77 , P1_R1138_U78 , P1_R1138_U79 , P1_R1138_U80 , P1_R1138_U81 , P1_R1138_U82 , P1_R1138_U83;
wire P1_R1138_U84 , P1_R1138_U85 , P1_R1138_U86 , P1_R1138_U87 , P1_R1138_U88 , P1_R1138_U89 , P1_R1138_U90 , P1_R1138_U91 , P1_R1138_U92 , P1_R1138_U93;
wire P1_R1138_U94 , P1_R1138_U95 , P1_R1138_U96 , P1_R1138_U97 , P1_R1138_U98 , P1_R1138_U99 , P1_R1138_U100 , P1_R1138_U101 , P1_R1138_U102 , P1_R1138_U103;
wire P1_R1138_U104 , P1_R1138_U105 , P1_R1138_U106 , P1_R1138_U107 , P1_R1138_U108 , P1_R1138_U109 , P1_R1138_U110 , P1_R1138_U111 , P1_R1138_U112 , P1_R1138_U113;
wire P1_R1138_U114 , P1_R1138_U115 , P1_R1138_U116 , P1_R1138_U117 , P1_R1138_U118 , P1_R1138_U119 , P1_R1138_U120 , P1_R1138_U121 , P1_R1138_U122 , P1_R1138_U123;
wire P1_R1138_U124 , P1_R1138_U125 , P1_R1138_U126 , P1_R1138_U127 , P1_R1138_U128 , P1_R1138_U129 , P1_R1138_U130 , P1_R1138_U131 , P1_R1138_U132 , P1_R1138_U133;
wire P1_R1138_U134 , P1_R1138_U135 , P1_R1138_U136 , P1_R1138_U137 , P1_R1138_U138 , P1_R1138_U139 , P1_R1138_U140 , P1_R1138_U141 , P1_R1138_U142 , P1_R1138_U143;
wire P1_R1138_U144 , P1_R1138_U145 , P1_R1138_U146 , P1_R1138_U147 , P1_R1138_U148 , P1_R1138_U149 , P1_R1138_U150 , P1_R1138_U151 , P1_R1138_U152 , P1_R1138_U153;
wire P1_R1138_U154 , P1_R1138_U155 , P1_R1138_U156 , P1_R1138_U157 , P1_R1138_U158 , P1_R1138_U159 , P1_R1138_U160 , P1_R1138_U161 , P1_R1138_U162 , P1_R1138_U163;
wire P1_R1138_U164 , P1_R1138_U165 , P1_R1138_U166 , P1_R1138_U167 , P1_R1138_U168 , P1_R1138_U169 , P1_R1138_U170 , P1_R1138_U171 , P1_R1138_U172 , P1_R1138_U173;
wire P1_R1138_U174 , P1_R1138_U175 , P1_R1138_U176 , P1_R1138_U177 , P1_R1138_U178 , P1_R1138_U179 , P1_R1138_U180 , P1_R1138_U181 , P1_R1138_U182 , P1_R1138_U183;
wire P1_R1138_U184 , P1_R1138_U185 , P1_R1138_U186 , P1_R1138_U187 , P1_R1138_U188 , P1_R1138_U189 , P1_R1138_U190 , P1_R1138_U191 , P1_R1138_U192 , P1_R1138_U193;
wire P1_R1138_U194 , P1_R1138_U195 , P1_R1138_U196 , P1_R1138_U197 , P1_R1138_U198 , P1_R1138_U199 , P1_R1138_U200 , P1_R1138_U201 , P1_R1138_U202 , P1_R1138_U203;
wire P1_R1138_U204 , P1_R1138_U205 , P1_R1138_U206 , P1_R1138_U207 , P1_R1138_U208 , P1_R1138_U209 , P1_R1138_U210 , P1_R1138_U211 , P1_R1138_U212 , P1_R1138_U213;
wire P1_R1138_U214 , P1_R1138_U215 , P1_R1138_U216 , P1_R1138_U217 , P1_R1138_U218 , P1_R1138_U219 , P1_R1138_U220 , P1_R1138_U221 , P1_R1138_U222 , P1_R1138_U223;
wire P1_R1138_U224 , P1_R1138_U225 , P1_R1138_U226 , P1_R1138_U227 , P1_R1138_U228 , P1_R1138_U229 , P1_R1138_U230 , P1_R1138_U231 , P1_R1138_U232 , P1_R1138_U233;
wire P1_R1138_U234 , P1_R1138_U235 , P1_R1138_U236 , P1_R1138_U237 , P1_R1138_U238 , P1_R1138_U239 , P1_R1138_U240 , P1_R1138_U241 , P1_R1138_U242 , P1_R1138_U243;
wire P1_R1138_U244 , P1_R1138_U245 , P1_R1138_U246 , P1_R1138_U247 , P1_R1138_U248 , P1_R1138_U249 , P1_R1138_U250 , P1_R1138_U251 , P1_R1138_U252 , P1_R1138_U253;
wire P1_R1138_U254 , P1_R1138_U255 , P1_R1138_U256 , P1_R1138_U257 , P1_R1138_U258 , P1_R1138_U259 , P1_R1138_U260 , P1_R1138_U261 , P1_R1138_U262 , P1_R1138_U263;
wire P1_R1138_U264 , P1_R1138_U265 , P1_R1138_U266 , P1_R1138_U267 , P1_R1138_U268 , P1_R1138_U269 , P1_R1138_U270 , P1_R1138_U271 , P1_R1138_U272 , P1_R1138_U273;
wire P1_R1138_U274 , P1_R1138_U275 , P1_R1138_U276 , P1_R1138_U277 , P1_R1138_U278 , P1_R1138_U279 , P1_R1138_U280 , P1_R1138_U281 , P1_R1138_U282 , P1_R1138_U283;
wire P1_R1138_U284 , P1_R1138_U285 , P1_R1138_U286 , P1_R1138_U287 , P1_R1138_U288 , P1_R1138_U289 , P1_R1138_U290 , P1_R1138_U291 , P1_R1138_U292 , P1_R1138_U293;
wire P1_R1138_U294 , P1_R1138_U295 , P1_R1138_U296 , P1_R1138_U297 , P1_R1138_U298 , P1_R1138_U299 , P1_R1138_U300 , P1_R1138_U301 , P1_R1138_U302 , P1_R1138_U303;
wire P1_R1138_U304 , P1_R1138_U305 , P1_R1138_U306 , P1_R1138_U307 , P1_R1138_U308 , P1_R1138_U309 , P1_R1138_U310 , P1_R1138_U311 , P1_R1138_U312 , P1_R1138_U313;
wire P1_R1138_U314 , P1_R1138_U315 , P1_R1138_U316 , P1_R1138_U317 , P1_R1138_U318 , P1_R1138_U319 , P1_R1138_U320 , P1_R1138_U321 , P1_R1138_U322 , P1_R1138_U323;
wire P1_R1138_U324 , P1_R1138_U325 , P1_R1138_U326 , P1_R1138_U327 , P1_R1138_U328 , P1_R1138_U329 , P1_R1138_U330 , P1_R1138_U331 , P1_R1138_U332 , P1_R1138_U333;
wire P1_R1138_U334 , P1_R1138_U335 , P1_R1138_U336 , P1_R1138_U337 , P1_R1138_U338 , P1_R1138_U339 , P1_R1138_U340 , P1_R1138_U341 , P1_R1138_U342 , P1_R1138_U343;
wire P1_R1138_U344 , P1_R1138_U345 , P1_R1138_U346 , P1_R1138_U347 , P1_R1138_U348 , P1_R1138_U349 , P1_R1138_U350 , P1_R1138_U351 , P1_R1138_U352 , P1_R1138_U353;
wire P1_R1138_U354 , P1_R1138_U355 , P1_R1138_U356 , P1_R1138_U357 , P1_R1138_U358 , P1_R1138_U359 , P1_R1138_U360 , P1_R1138_U361 , P1_R1138_U362 , P1_R1138_U363;
wire P1_R1138_U364 , P1_R1138_U365 , P1_R1138_U366 , P1_R1138_U367 , P1_R1138_U368 , P1_R1138_U369 , P1_R1138_U370 , P1_R1138_U371 , P1_R1138_U372 , P1_R1138_U373;
wire P1_R1138_U374 , P1_R1138_U375 , P1_R1138_U376 , P1_R1138_U377 , P1_R1138_U378 , P1_R1138_U379 , P1_R1138_U380 , P1_R1138_U381 , P1_R1138_U382 , P1_R1138_U383;
wire P1_R1138_U384 , P1_R1138_U385 , P1_R1138_U386 , P1_R1138_U387 , P1_R1138_U388 , P1_R1138_U389 , P1_R1138_U390 , P1_R1138_U391 , P1_R1138_U392 , P1_R1138_U393;
wire P1_R1138_U394 , P1_R1138_U395 , P1_R1138_U396 , P1_R1138_U397 , P1_R1138_U398 , P1_R1138_U399 , P1_R1138_U400 , P1_R1138_U401 , P1_R1138_U402 , P1_R1138_U403;
wire P1_R1138_U404 , P1_R1138_U405 , P1_R1138_U406 , P1_R1138_U407 , P1_R1138_U408 , P1_R1138_U409 , P1_R1138_U410 , P1_R1138_U411 , P1_R1138_U412 , P1_R1138_U413;
wire P1_R1138_U414 , P1_R1138_U415 , P1_R1138_U416 , P1_R1138_U417 , P1_R1138_U418 , P1_R1138_U419 , P1_R1138_U420 , P1_R1138_U421 , P1_R1138_U422 , P1_R1138_U423;
wire P1_R1138_U424 , P1_R1138_U425 , P1_R1138_U426 , P1_R1138_U427 , P1_R1138_U428 , P1_R1138_U429 , P1_R1138_U430 , P1_R1138_U431 , P1_R1138_U432 , P1_R1138_U433;
wire P1_R1138_U434 , P1_R1138_U435 , P1_R1138_U436 , P1_R1138_U437 , P1_R1138_U438 , P1_R1138_U439 , P1_R1138_U440 , P1_R1138_U441 , P1_R1138_U442 , P1_R1138_U443;
wire P1_R1138_U444 , P1_R1138_U445 , P1_R1138_U446 , P1_R1138_U447 , P1_R1138_U448 , P1_R1138_U449 , P1_R1138_U450 , P1_R1138_U451 , P1_R1138_U452 , P1_R1138_U453;
wire P1_R1138_U454 , P1_R1138_U455 , P1_R1138_U456 , P1_R1138_U457 , P1_R1138_U458 , P1_R1138_U459 , P1_R1138_U460 , P1_R1138_U461 , P1_R1138_U462 , P1_R1138_U463;
wire P1_R1138_U464 , P1_R1138_U465 , P1_R1138_U466 , P1_R1138_U467 , P1_R1138_U468 , P1_R1138_U469 , P1_R1138_U470 , P1_R1138_U471 , P1_R1138_U472 , P1_R1138_U473;
wire P1_R1138_U474 , P1_R1138_U475 , P1_R1138_U476 , P1_R1138_U477 , P1_R1138_U478 , P1_R1138_U479 , P1_R1138_U480 , P1_R1138_U481 , P1_R1138_U482 , P1_R1138_U483;
wire P1_R1138_U484 , P1_R1138_U485 , P1_R1138_U486 , P1_R1138_U487 , P1_R1138_U488 , P1_R1138_U489 , P1_R1138_U490 , P1_R1138_U491 , P1_R1138_U492 , P1_R1138_U493;
wire P1_R1138_U494 , P1_R1138_U495 , P1_R1138_U496 , P1_R1138_U497 , P1_R1138_U498 , P1_R1138_U499 , P1_R1138_U500 , P1_R1138_U501 , P1_R1222_U4 , P1_R1222_U5;
wire P1_R1222_U6 , P1_R1222_U7 , P1_R1222_U8 , P1_R1222_U9 , P1_R1222_U10 , P1_R1222_U11 , P1_R1222_U12 , P1_R1222_U13 , P1_R1222_U14 , P1_R1222_U15;
wire P1_R1222_U16 , P1_R1222_U17 , P1_R1222_U18 , P1_R1222_U19 , P1_R1222_U20 , P1_R1222_U21 , P1_R1222_U22 , P1_R1222_U23 , P1_R1222_U24 , P1_R1222_U25;
wire P1_R1222_U26 , P1_R1222_U27 , P1_R1222_U28 , P1_R1222_U29 , P1_R1222_U30 , P1_R1222_U31 , P1_R1222_U32 , P1_R1222_U33 , P1_R1222_U34 , P1_R1222_U35;
wire P1_R1222_U36 , P1_R1222_U37 , P1_R1222_U38 , P1_R1222_U39 , P1_R1222_U40 , P1_R1222_U41 , P1_R1222_U42 , P1_R1222_U43 , P1_R1222_U44 , P1_R1222_U45;
wire P1_R1222_U46 , P1_R1222_U47 , P1_R1222_U48 , P1_R1222_U49 , P1_R1222_U50 , P1_R1222_U51 , P1_R1222_U52 , P1_R1222_U53 , P1_R1222_U54 , P1_R1222_U55;
wire P1_R1222_U56 , P1_R1222_U57 , P1_R1222_U58 , P1_R1222_U59 , P1_R1222_U60 , P1_R1222_U61 , P1_R1222_U62 , P1_R1222_U63 , P1_R1222_U64 , P1_R1222_U65;
wire P1_R1222_U66 , P1_R1222_U67 , P1_R1222_U68 , P1_R1222_U69 , P1_R1222_U70 , P1_R1222_U71 , P1_R1222_U72 , P1_R1222_U73 , P1_R1222_U74 , P1_R1222_U75;
wire P1_R1222_U76 , P1_R1222_U77 , P1_R1222_U78 , P1_R1222_U79 , P1_R1222_U80 , P1_R1222_U81 , P1_R1222_U82 , P1_R1222_U83 , P1_R1222_U84 , P1_R1222_U85;
wire P1_R1222_U86 , P1_R1222_U87 , P1_R1222_U88 , P1_R1222_U89 , P1_R1222_U90 , P1_R1222_U91 , P1_R1222_U92 , P1_R1222_U93 , P1_R1222_U94 , P1_R1222_U95;
wire P1_R1222_U96 , P1_R1222_U97 , P1_R1222_U98 , P1_R1222_U99 , P1_R1222_U100 , P1_R1222_U101 , P1_R1222_U102 , P1_R1222_U103 , P1_R1222_U104 , P1_R1222_U105;
wire P1_R1222_U106 , P1_R1222_U107 , P1_R1222_U108 , P1_R1222_U109 , P1_R1222_U110 , P1_R1222_U111 , P1_R1222_U112 , P1_R1222_U113 , P1_R1222_U114 , P1_R1222_U115;
wire P1_R1222_U116 , P1_R1222_U117 , P1_R1222_U118 , P1_R1222_U119 , P1_R1222_U120 , P1_R1222_U121 , P1_R1222_U122 , P1_R1222_U123 , P1_R1222_U124 , P1_R1222_U125;
wire P1_R1222_U126 , P1_R1222_U127 , P1_R1222_U128 , P1_R1222_U129 , P1_R1222_U130 , P1_R1222_U131 , P1_R1222_U132 , P1_R1222_U133 , P1_R1222_U134 , P1_R1222_U135;
wire P1_R1222_U136 , P1_R1222_U137 , P1_R1222_U138 , P1_R1222_U139 , P1_R1222_U140 , P1_R1222_U141 , P1_R1222_U142 , P1_R1222_U143 , P1_R1222_U144 , P1_R1222_U145;
wire P1_R1222_U146 , P1_R1222_U147 , P1_R1222_U148 , P1_R1222_U149 , P1_R1222_U150 , P1_R1222_U151 , P1_R1222_U152 , P1_R1222_U153 , P1_R1222_U154 , P1_R1222_U155;
wire P1_R1222_U156 , P1_R1222_U157 , P1_R1222_U158 , P1_R1222_U159 , P1_R1222_U160 , P1_R1222_U161 , P1_R1222_U162 , P1_R1222_U163 , P1_R1222_U164 , P1_R1222_U165;
wire P1_R1222_U166 , P1_R1222_U167 , P1_R1222_U168 , P1_R1222_U169 , P1_R1222_U170 , P1_R1222_U171 , P1_R1222_U172 , P1_R1222_U173 , P1_R1222_U174 , P1_R1222_U175;
wire P1_R1222_U176 , P1_R1222_U177 , P1_R1222_U178 , P1_R1222_U179 , P1_R1222_U180 , P1_R1222_U181 , P1_R1222_U182 , P1_R1222_U183 , P1_R1222_U184 , P1_R1222_U185;
wire P1_R1222_U186 , P1_R1222_U187 , P1_R1222_U188 , P1_R1222_U189 , P1_R1222_U190 , P1_R1222_U191 , P1_R1222_U192 , P1_R1222_U193 , P1_R1222_U194 , P1_R1222_U195;
wire P1_R1222_U196 , P1_R1222_U197 , P1_R1222_U198 , P1_R1222_U199 , P1_R1222_U200 , P1_R1222_U201 , P1_R1222_U202 , P1_R1222_U203 , P1_R1222_U204 , P1_R1222_U205;
wire P1_R1222_U206 , P1_R1222_U207 , P1_R1222_U208 , P1_R1222_U209 , P1_R1222_U210 , P1_R1222_U211 , P1_R1222_U212 , P1_R1222_U213 , P1_R1222_U214 , P1_R1222_U215;
wire P1_R1222_U216 , P1_R1222_U217 , P1_R1222_U218 , P1_R1222_U219 , P1_R1222_U220 , P1_R1222_U221 , P1_R1222_U222 , P1_R1222_U223 , P1_R1222_U224 , P1_R1222_U225;
wire P1_R1222_U226 , P1_R1222_U227 , P1_R1222_U228 , P1_R1222_U229 , P1_R1222_U230 , P1_R1222_U231 , P1_R1222_U232 , P1_R1222_U233 , P1_R1222_U234 , P1_R1222_U235;
wire P1_R1222_U236 , P1_R1222_U237 , P1_R1222_U238 , P1_R1222_U239 , P1_R1222_U240 , P1_R1222_U241 , P1_R1222_U242 , P1_R1222_U243 , P1_R1222_U244 , P1_R1222_U245;
wire P1_R1222_U246 , P1_R1222_U247 , P1_R1222_U248 , P1_R1222_U249 , P1_R1222_U250 , P1_R1222_U251 , P1_R1222_U252 , P1_R1222_U253 , P1_R1222_U254 , P1_R1222_U255;
wire P1_R1222_U256 , P1_R1222_U257 , P1_R1222_U258 , P1_R1222_U259 , P1_R1222_U260 , P1_R1222_U261 , P1_R1222_U262 , P1_R1222_U263 , P1_R1222_U264 , P1_R1222_U265;
wire P1_R1222_U266 , P1_R1222_U267 , P1_R1222_U268 , P1_R1222_U269 , P1_R1222_U270 , P1_R1222_U271 , P1_R1222_U272 , P1_R1222_U273 , P1_R1222_U274 , P1_R1222_U275;
wire P1_R1222_U276 , P1_R1222_U277 , P1_R1222_U278 , P1_R1222_U279 , P1_R1222_U280 , P1_R1222_U281 , P1_R1222_U282 , P1_R1222_U283 , P1_R1222_U284 , P1_R1222_U285;
wire P1_R1222_U286 , P1_R1222_U287 , P1_R1222_U288 , P1_R1222_U289 , P1_R1222_U290 , P1_R1222_U291 , P1_R1222_U292 , P1_R1222_U293 , P1_R1222_U294 , P1_R1222_U295;
wire P1_R1222_U296 , P1_R1222_U297 , P1_R1222_U298 , P1_R1222_U299 , P1_R1222_U300 , P1_R1222_U301 , P1_R1222_U302 , P1_R1222_U303 , P1_R1222_U304 , P1_R1222_U305;
wire P1_R1222_U306 , P1_R1222_U307 , P1_R1222_U308 , P1_R1222_U309 , P1_R1222_U310 , P1_R1222_U311 , P1_R1222_U312 , P1_R1222_U313 , P1_R1222_U314 , P1_R1222_U315;
wire P1_R1222_U316 , P1_R1222_U317 , P1_R1222_U318 , P1_R1222_U319 , P1_R1222_U320 , P1_R1222_U321 , P1_R1222_U322 , P1_R1222_U323 , P1_R1222_U324 , P1_R1222_U325;
wire P1_R1222_U326 , P1_R1222_U327 , P1_R1222_U328 , P1_R1222_U329 , P1_R1222_U330 , P1_R1222_U331 , P1_R1222_U332 , P1_R1222_U333 , P1_R1222_U334 , P1_R1222_U335;
wire P1_R1222_U336 , P1_R1222_U337 , P1_R1222_U338 , P1_R1222_U339 , P1_R1222_U340 , P1_R1222_U341 , P1_R1222_U342 , P1_R1222_U343 , P1_R1222_U344 , P1_R1222_U345;
wire P1_R1222_U346 , P1_R1222_U347 , P1_R1222_U348 , P1_R1222_U349 , P1_R1222_U350 , P1_R1222_U351 , P1_R1222_U352 , P1_R1222_U353 , P1_R1222_U354 , P1_R1222_U355;
wire P1_R1222_U356 , P1_R1222_U357 , P1_R1222_U358 , P1_R1222_U359 , P1_R1222_U360 , P1_R1222_U361 , P1_R1222_U362 , P1_R1222_U363 , P1_R1222_U364 , P1_R1222_U365;
wire P1_R1222_U366 , P1_R1222_U367 , P1_R1222_U368 , P1_R1222_U369 , P1_R1222_U370 , P1_R1222_U371 , P1_R1222_U372 , P1_R1222_U373 , P1_R1222_U374 , P1_R1222_U375;
wire P1_R1222_U376 , P1_R1222_U377 , P1_R1222_U378 , P1_R1222_U379 , P1_R1222_U380 , P1_R1222_U381 , P1_R1222_U382 , P1_R1222_U383 , P1_R1222_U384 , P1_R1222_U385;
wire P1_R1222_U386 , P1_R1222_U387 , P1_R1222_U388 , P1_R1222_U389 , P1_R1222_U390 , P1_R1222_U391 , P1_R1222_U392 , P1_R1222_U393 , P1_R1222_U394 , P1_R1222_U395;
wire P1_R1222_U396 , P1_R1222_U397 , P1_R1222_U398 , P1_R1222_U399 , P1_R1222_U400 , P1_R1222_U401 , P1_R1222_U402 , P1_R1222_U403 , P1_R1222_U404 , P1_R1222_U405;
wire P1_R1222_U406 , P1_R1222_U407 , P1_R1222_U408 , P1_R1222_U409 , P1_R1222_U410 , P1_R1222_U411 , P1_R1222_U412 , P1_R1222_U413 , P1_R1222_U414 , P1_R1222_U415;
wire P1_R1222_U416 , P1_R1222_U417 , P1_R1222_U418 , P1_R1222_U419 , P1_R1222_U420 , P1_R1222_U421 , P1_R1222_U422 , P1_R1222_U423 , P1_R1222_U424 , P1_R1222_U425;
wire P1_R1222_U426 , P1_R1222_U427 , P1_R1222_U428 , P1_R1222_U429 , P1_R1222_U430 , P1_R1222_U431 , P1_R1222_U432 , P1_R1222_U433 , P1_R1222_U434 , P1_R1222_U435;
wire P1_R1222_U436 , P1_R1222_U437 , P1_R1222_U438 , P1_R1222_U439 , P1_R1222_U440 , P1_R1222_U441 , P1_R1222_U442 , P1_R1222_U443 , P1_R1222_U444 , P1_R1222_U445;
wire P1_R1222_U446 , P1_R1222_U447 , P1_R1222_U448 , P1_R1222_U449 , P1_R1222_U450 , P1_R1222_U451 , P1_R1222_U452 , P1_R1222_U453 , P1_R1222_U454 , P1_R1222_U455;
wire P1_R1222_U456 , P1_R1222_U457 , P1_R1222_U458 , P1_R1222_U459 , P1_R1222_U460 , P1_R1222_U461 , P1_R1222_U462 , P1_R1222_U463 , P1_R1222_U464 , P1_R1222_U465;
wire P1_R1222_U466 , P1_R1222_U467 , P1_R1222_U468 , P1_R1222_U469 , P1_R1222_U470 , P1_R1222_U471 , P1_R1222_U472 , P1_R1222_U473 , P1_R1222_U474 , P1_R1222_U475;
wire P1_R1222_U476 , P1_R1222_U477 , P1_R1222_U478 , P1_R1222_U479 , P1_R1222_U480 , P1_R1222_U481 , P1_R1222_U482 , P1_R1222_U483 , P1_R1222_U484 , P1_R1222_U485;
wire P1_R1222_U486 , P1_R1222_U487 , P1_R1222_U488 , P1_R1222_U489 , P1_R1222_U490 , P1_R1222_U491 , P1_R1222_U492 , P1_R1222_U493 , P1_R1222_U494 , P1_R1222_U495;
wire P1_R1222_U496 , P1_R1222_U497 , P1_R1222_U498 , P1_R1222_U499 , P1_R1222_U500 , P1_R1222_U501 , P2_ADD_1119_U4 , P2_ADD_1119_U5 , P2_ADD_1119_U6 , P2_ADD_1119_U7;
wire P2_ADD_1119_U8 , P2_ADD_1119_U9 , P2_ADD_1119_U10 , P2_ADD_1119_U11 , P2_ADD_1119_U12 , P2_ADD_1119_U13 , P2_ADD_1119_U14 , P2_ADD_1119_U15 , P2_ADD_1119_U16 , P2_ADD_1119_U17;
wire P2_ADD_1119_U18 , P2_ADD_1119_U19 , P2_ADD_1119_U20 , P2_ADD_1119_U21 , P2_ADD_1119_U22 , P2_ADD_1119_U23 , P2_ADD_1119_U24 , P2_ADD_1119_U25 , P2_ADD_1119_U26 , P2_ADD_1119_U27;
wire P2_ADD_1119_U28 , P2_ADD_1119_U29 , P2_ADD_1119_U30 , P2_ADD_1119_U31 , P2_ADD_1119_U32 , P2_ADD_1119_U33 , P2_ADD_1119_U34 , P2_ADD_1119_U35 , P2_ADD_1119_U36 , P2_ADD_1119_U37;
wire P2_ADD_1119_U38 , P2_ADD_1119_U39 , P2_ADD_1119_U40 , P2_ADD_1119_U41 , P2_ADD_1119_U42 , P2_ADD_1119_U43 , P2_ADD_1119_U44 , P2_ADD_1119_U45 , P2_ADD_1119_U46 , P2_ADD_1119_U47;
wire P2_ADD_1119_U48 , P2_ADD_1119_U49 , P2_ADD_1119_U50 , P2_ADD_1119_U51 , P2_ADD_1119_U52 , P2_ADD_1119_U53 , P2_ADD_1119_U54 , P2_ADD_1119_U55 , P2_ADD_1119_U56 , P2_ADD_1119_U57;
wire P2_ADD_1119_U58 , P2_ADD_1119_U59 , P2_ADD_1119_U60 , P2_ADD_1119_U61 , P2_ADD_1119_U62 , P2_ADD_1119_U63 , P2_ADD_1119_U64 , P2_ADD_1119_U65 , P2_ADD_1119_U66 , P2_ADD_1119_U67;
wire P2_ADD_1119_U68 , P2_ADD_1119_U69 , P2_ADD_1119_U70 , P2_ADD_1119_U71 , P2_ADD_1119_U72 , P2_ADD_1119_U73 , P2_ADD_1119_U74 , P2_ADD_1119_U75 , P2_ADD_1119_U76 , P2_ADD_1119_U77;
wire P2_ADD_1119_U78 , P2_ADD_1119_U79 , P2_ADD_1119_U80 , P2_ADD_1119_U81 , P2_ADD_1119_U82 , P2_ADD_1119_U83 , P2_ADD_1119_U84 , P2_ADD_1119_U85 , P2_ADD_1119_U86 , P2_ADD_1119_U87;
wire P2_ADD_1119_U88 , P2_ADD_1119_U89 , P2_ADD_1119_U90 , P2_ADD_1119_U91 , P2_ADD_1119_U92 , P2_ADD_1119_U93 , P2_ADD_1119_U94 , P2_ADD_1119_U95 , P2_ADD_1119_U96 , P2_ADD_1119_U97;
wire P2_ADD_1119_U98 , P2_ADD_1119_U99 , P2_ADD_1119_U100 , P2_ADD_1119_U101 , P2_ADD_1119_U102 , P2_ADD_1119_U103 , P2_ADD_1119_U104 , P2_ADD_1119_U105 , P2_ADD_1119_U106 , P2_ADD_1119_U107;
wire P2_ADD_1119_U108 , P2_ADD_1119_U109 , P2_ADD_1119_U110 , P2_ADD_1119_U111 , P2_ADD_1119_U112 , P2_ADD_1119_U113 , P2_ADD_1119_U114 , P2_ADD_1119_U115 , P2_ADD_1119_U116 , P2_ADD_1119_U117;
wire P2_ADD_1119_U118 , P2_ADD_1119_U119 , P2_ADD_1119_U120 , P2_ADD_1119_U121 , P2_ADD_1119_U122 , P2_ADD_1119_U123 , P2_ADD_1119_U124 , P2_ADD_1119_U125 , P2_ADD_1119_U126 , P2_ADD_1119_U127;
wire P2_ADD_1119_U128 , P2_ADD_1119_U129 , P2_ADD_1119_U130 , P2_ADD_1119_U131 , P2_ADD_1119_U132 , P2_ADD_1119_U133 , P2_ADD_1119_U134 , P2_ADD_1119_U135 , P2_ADD_1119_U136 , P2_ADD_1119_U137;
wire P2_ADD_1119_U138 , P2_ADD_1119_U139 , P2_ADD_1119_U140 , P2_ADD_1119_U141 , P2_ADD_1119_U142 , P2_ADD_1119_U143 , P2_ADD_1119_U144 , P2_ADD_1119_U145 , P2_ADD_1119_U146 , P2_ADD_1119_U147;
wire P2_ADD_1119_U148 , P2_ADD_1119_U149 , P2_ADD_1119_U150 , P2_ADD_1119_U151 , P2_ADD_1119_U152 , P2_ADD_1119_U153 , P2_ADD_1119_U154 , P2_ADD_1119_U155 , P2_ADD_1119_U156 , P2_ADD_1119_U157;
wire P2_SUB_1108_U6 , P2_SUB_1108_U7 , P2_SUB_1108_U8 , P2_SUB_1108_U9 , P2_SUB_1108_U10 , P2_SUB_1108_U11 , P2_SUB_1108_U12 , P2_SUB_1108_U13 , P2_SUB_1108_U14 , P2_SUB_1108_U15;
wire P2_SUB_1108_U16 , P2_SUB_1108_U17 , P2_SUB_1108_U18 , P2_SUB_1108_U19 , P2_SUB_1108_U20 , P2_SUB_1108_U21 , P2_SUB_1108_U22 , P2_SUB_1108_U23 , P2_SUB_1108_U24 , P2_SUB_1108_U25;
wire P2_SUB_1108_U26 , P2_SUB_1108_U27 , P2_SUB_1108_U28 , P2_SUB_1108_U29 , P2_SUB_1108_U30 , P2_SUB_1108_U31 , P2_SUB_1108_U32 , P2_SUB_1108_U33 , P2_SUB_1108_U34 , P2_SUB_1108_U35;
wire P2_SUB_1108_U36 , P2_SUB_1108_U37 , P2_SUB_1108_U38 , P2_SUB_1108_U39 , P2_SUB_1108_U40 , P2_SUB_1108_U41 , P2_SUB_1108_U42 , P2_SUB_1108_U43 , P2_SUB_1108_U44 , P2_SUB_1108_U45;
wire P2_SUB_1108_U46 , P2_SUB_1108_U47 , P2_SUB_1108_U48 , P2_SUB_1108_U49 , P2_SUB_1108_U50 , P2_SUB_1108_U51 , P2_SUB_1108_U52 , P2_SUB_1108_U53 , P2_SUB_1108_U54 , P2_SUB_1108_U55;
wire P2_SUB_1108_U56 , P2_SUB_1108_U57 , P2_SUB_1108_U58 , P2_SUB_1108_U59 , P2_SUB_1108_U60 , P2_SUB_1108_U61 , P2_SUB_1108_U62 , P2_SUB_1108_U63 , P2_SUB_1108_U64 , P2_SUB_1108_U65;
wire P2_SUB_1108_U66 , P2_SUB_1108_U67 , P2_SUB_1108_U68 , P2_SUB_1108_U69 , P2_SUB_1108_U70 , P2_SUB_1108_U71 , P2_SUB_1108_U72 , P2_SUB_1108_U73 , P2_SUB_1108_U74 , P2_SUB_1108_U75;
wire P2_SUB_1108_U76 , P2_SUB_1108_U77 , P2_SUB_1108_U78 , P2_SUB_1108_U79 , P2_SUB_1108_U80 , P2_SUB_1108_U81 , P2_SUB_1108_U82 , P2_SUB_1108_U83 , P2_SUB_1108_U84 , P2_SUB_1108_U85;
wire P2_SUB_1108_U86 , P2_SUB_1108_U87 , P2_SUB_1108_U88 , P2_SUB_1108_U89 , P2_SUB_1108_U90 , P2_SUB_1108_U91 , P2_SUB_1108_U92 , P2_SUB_1108_U93 , P2_SUB_1108_U94 , P2_SUB_1108_U95;
wire P2_SUB_1108_U96 , P2_SUB_1108_U97 , P2_SUB_1108_U98 , P2_SUB_1108_U99 , P2_SUB_1108_U100 , P2_SUB_1108_U101 , P2_SUB_1108_U102 , P2_SUB_1108_U103 , P2_SUB_1108_U104 , P2_SUB_1108_U105;
wire P2_SUB_1108_U106 , P2_SUB_1108_U107 , P2_SUB_1108_U108 , P2_SUB_1108_U109 , P2_SUB_1108_U110 , P2_SUB_1108_U111 , P2_SUB_1108_U112 , P2_SUB_1108_U113 , P2_SUB_1108_U114 , P2_SUB_1108_U115;
wire P2_SUB_1108_U116 , P2_SUB_1108_U117 , P2_SUB_1108_U118 , P2_SUB_1108_U119 , P2_SUB_1108_U120 , P2_SUB_1108_U121 , P2_SUB_1108_U122 , P2_SUB_1108_U123 , P2_SUB_1108_U124 , P2_SUB_1108_U125;
wire P2_SUB_1108_U126 , P2_SUB_1108_U127 , P2_SUB_1108_U128 , P2_SUB_1108_U129 , P2_SUB_1108_U130 , P2_SUB_1108_U131 , P2_SUB_1108_U132 , P2_SUB_1108_U133 , P2_SUB_1108_U134 , P2_SUB_1108_U135;
wire P2_SUB_1108_U136 , P2_SUB_1108_U137 , P2_SUB_1108_U138 , P2_SUB_1108_U139 , P2_SUB_1108_U140 , P2_SUB_1108_U141 , P2_SUB_1108_U142 , P2_SUB_1108_U143 , P2_SUB_1108_U144 , P2_SUB_1108_U145;
wire P2_SUB_1108_U146 , P2_SUB_1108_U147 , P2_SUB_1108_U148 , P2_SUB_1108_U149 , P2_SUB_1108_U150 , P2_SUB_1108_U151 , P2_SUB_1108_U152 , P2_SUB_1108_U153 , P2_SUB_1108_U154 , P2_SUB_1108_U155;
wire P2_SUB_1108_U156 , P2_SUB_1108_U157 , P2_SUB_1108_U158 , P2_SUB_1108_U159 , P2_SUB_1108_U160 , P2_SUB_1108_U161 , P2_SUB_1108_U162 , P2_SUB_1108_U163 , P2_SUB_1108_U164 , P2_SUB_1108_U165;
wire P2_SUB_1108_U166 , P2_SUB_1108_U167 , P2_SUB_1108_U168 , P2_SUB_1108_U169 , P2_SUB_1108_U170 , P2_SUB_1108_U171 , P2_SUB_1108_U172 , P2_SUB_1108_U173 , P2_SUB_1108_U174 , P2_SUB_1108_U175;
wire P2_SUB_1108_U176 , P2_SUB_1108_U177 , P2_SUB_1108_U178 , P2_SUB_1108_U179 , P2_SUB_1108_U180 , P2_SUB_1108_U181 , P2_SUB_1108_U182 , P2_SUB_1108_U183 , P2_SUB_1108_U184 , P2_SUB_1108_U185;
wire P2_SUB_1108_U186 , P2_SUB_1108_U187 , P2_SUB_1108_U188 , P2_SUB_1108_U189 , P2_SUB_1108_U190 , P2_SUB_1108_U191 , P2_SUB_1108_U192 , P2_SUB_1108_U193 , P2_SUB_1108_U194 , P2_SUB_1108_U195;
wire P2_SUB_1108_U196 , P2_SUB_1108_U197 , P2_SUB_1108_U198 , P2_SUB_1108_U199 , P2_SUB_1108_U200 , P2_SUB_1108_U201 , P2_SUB_1108_U202 , P2_R1299_U6 , P2_R1299_U7 , P2_R1312_U6;
wire P2_R1312_U7 , P2_R1312_U8 , P2_R1312_U9 , P2_R1312_U10 , P2_R1312_U11 , P2_R1312_U12 , P2_R1312_U13 , P2_R1312_U14 , P2_R1312_U15 , P2_R1312_U16;
wire P2_R1312_U17 , P2_R1312_U18 , P2_R1312_U19 , P2_R1312_U20 , P2_R1312_U21 , P2_R1312_U22 , P2_R1312_U23 , P2_R1312_U24 , P2_R1312_U25 , P2_R1312_U26;
wire P2_R1312_U27 , P2_R1312_U28 , P2_R1312_U29 , P2_R1312_U30 , P2_R1312_U31 , P2_R1312_U32 , P2_R1312_U33 , P2_R1312_U34 , P2_R1312_U35 , P2_R1312_U36;
wire P2_R1312_U37 , P2_R1312_U38 , P2_R1312_U39 , P2_R1312_U40 , P2_R1312_U41 , P2_R1312_U42 , P2_R1312_U43 , P2_R1312_U44 , P2_R1312_U45 , P2_R1312_U46;
wire P2_R1312_U47 , P2_R1312_U48 , P2_R1312_U49 , P2_R1312_U50 , P2_R1312_U51 , P2_R1312_U52 , P2_R1312_U53 , P2_R1312_U54 , P2_R1312_U55 , P2_R1312_U56;
wire P2_R1312_U57 , P2_R1312_U58 , P2_R1312_U59 , P2_R1312_U60 , P2_R1312_U61 , P2_R1312_U62 , P2_R1312_U63 , P2_R1312_U64 , P2_R1312_U65 , P2_R1312_U66;
wire P2_R1312_U67 , P2_R1312_U68 , P2_R1312_U69 , P2_R1312_U70 , P2_R1312_U71 , P2_R1312_U72 , P2_R1312_U73 , P2_R1312_U74 , P2_R1312_U75 , P2_R1312_U76;
wire P2_R1312_U77 , P2_R1312_U78 , P2_R1312_U79 , P2_R1312_U80 , P2_R1312_U81 , P2_R1312_U82 , P2_R1312_U83 , P2_R1312_U84 , P2_R1312_U85 , P2_R1312_U86;
wire P2_R1312_U87 , P2_R1312_U88 , P2_R1312_U89 , P2_R1312_U90 , P2_R1312_U91 , P2_R1312_U92 , P2_R1312_U93 , P2_R1312_U94 , P2_R1312_U95 , P2_R1312_U96;
wire P2_R1312_U97 , P2_R1312_U98 , P2_R1312_U99 , P2_R1312_U100 , P2_R1312_U101 , P2_R1312_U102 , P2_R1312_U103 , P2_R1312_U104 , P2_R1312_U105 , P2_R1312_U106;
wire P2_R1312_U107 , P2_R1312_U108 , P2_R1312_U109 , P2_R1312_U110 , P2_R1312_U111 , P2_R1312_U112 , P2_R1312_U113 , P2_R1312_U114 , P2_R1312_U115 , P2_R1312_U116;
wire P2_R1312_U117 , P2_R1312_U118 , P2_R1312_U119 , P2_R1312_U120 , P2_R1312_U121 , P2_R1312_U122 , P2_R1312_U123 , P2_R1312_U124 , P2_R1312_U125 , P2_R1312_U126;
wire P2_R1312_U127 , P2_R1312_U128 , P2_R1312_U129 , P2_R1312_U130 , P2_R1312_U131 , P2_R1312_U132 , P2_R1312_U133 , P2_R1312_U134 , P2_R1312_U135 , P2_R1312_U136;
wire P2_R1312_U137 , P2_R1312_U138 , P2_R1312_U139 , P2_R1312_U140 , P2_R1312_U141 , P2_R1312_U142 , P2_R1312_U143 , P2_R1312_U144 , P2_R1312_U145 , P2_R1312_U146;
wire P2_R1312_U147 , P2_R1312_U148 , P2_R1312_U149 , P2_R1312_U150 , P2_R1312_U151 , P2_R1312_U152 , P2_R1312_U153 , P2_R1312_U154 , P2_R1312_U155 , P2_R1312_U156;
wire P2_R1312_U157 , P2_R1312_U158 , P2_R1312_U159 , P2_R1312_U160 , P2_R1312_U161 , P2_R1312_U162 , P2_R1312_U163 , P2_R1312_U164 , P2_R1312_U165 , P2_R1312_U166;
wire P2_R1312_U167 , P2_R1312_U168 , P2_R1312_U169 , P2_R1312_U170 , P2_R1312_U171 , P2_R1312_U172 , P2_R1312_U173 , P2_R1312_U174 , P2_R1312_U175 , P2_R1312_U176;
wire P2_R1312_U177 , P2_R1312_U178 , P2_R1312_U179 , P2_R1312_U180 , P2_R1312_U181 , P2_R1312_U182 , P2_R1312_U183 , P2_R1312_U184 , P2_R1312_U185 , P2_R1312_U186;
wire P2_R1312_U187 , P2_R1312_U188 , P2_R1312_U189 , P2_R1312_U190 , P2_R1312_U191 , P2_R1312_U192 , P2_R1312_U193 , P2_R1312_U194 , P2_R1312_U195 , P2_R1312_U196;
wire P2_R1312_U197 , P2_R1312_U198 , P2_R1312_U199 , P2_R1312_U200 , P2_R1312_U201 , P2_R1312_U202 , P2_R1312_U203 , P2_R1312_U204 , P2_R1312_U205 , P2_R1312_U206;
wire P2_R1312_U207 , P2_R1312_U208 , P2_R1312_U209 , P2_R1312_U210 , P2_R1312_U211 , P2_R1312_U212 , P2_R1312_U213 , P2_R1312_U214 , P2_R1312_U215 , P2_R1312_U216;
wire P2_R1312_U217 , P2_R1312_U218 , P2_R1312_U219 , P2_R1312_U220 , P2_R1312_U221 , P2_R1312_U222 , P2_R1312_U223 , P2_R1312_U224 , P2_R1312_U225 , P2_R1312_U226;
wire P2_R1312_U227 , P2_R1335_U6 , P2_R1335_U7 , P2_R1335_U8 , P2_R1335_U9 , P2_R1335_U10 , P2_R1209_U4 , P2_R1209_U5 , P2_R1209_U6 , P2_R1209_U7;
wire P2_R1209_U8 , P2_R1209_U9 , P2_R1209_U10 , P2_R1209_U11 , P2_R1209_U12 , P2_R1209_U13 , P2_R1209_U14 , P2_R1209_U15 , P2_R1209_U16 , P2_R1209_U17;
wire P2_R1209_U18 , P2_R1209_U19 , P2_R1209_U20 , P2_R1209_U21 , P2_R1209_U22 , P2_R1209_U23 , P2_R1209_U24 , P2_R1209_U25 , P2_R1209_U26 , P2_R1209_U27;
wire P2_R1209_U28 , P2_R1209_U29 , P2_R1209_U30 , P2_R1209_U31 , P2_R1209_U32 , P2_R1209_U33 , P2_R1209_U34 , P2_R1209_U35 , P2_R1209_U36 , P2_R1209_U37;
wire P2_R1209_U38 , P2_R1209_U39 , P2_R1209_U40 , P2_R1209_U41 , P2_R1209_U42 , P2_R1209_U43 , P2_R1209_U44 , P2_R1209_U45 , P2_R1209_U46 , P2_R1209_U47;
wire P2_R1209_U48 , P2_R1209_U49 , P2_R1209_U50 , P2_R1209_U51 , P2_R1209_U52 , P2_R1209_U53 , P2_R1209_U54 , P2_R1209_U55 , P2_R1209_U56 , P2_R1209_U57;
wire P2_R1209_U58 , P2_R1209_U59 , P2_R1209_U60 , P2_R1209_U61 , P2_R1209_U62 , P2_R1209_U63 , P2_R1209_U64 , P2_R1209_U65 , P2_R1209_U66 , P2_R1209_U67;
wire P2_R1209_U68 , P2_R1209_U69 , P2_R1209_U70 , P2_R1209_U71 , P2_R1209_U72 , P2_R1209_U73 , P2_R1209_U74 , P2_R1209_U75 , P2_R1209_U76 , P2_R1209_U77;
wire P2_R1209_U78 , P2_R1209_U79 , P2_R1209_U80 , P2_R1209_U81 , P2_R1209_U82 , P2_R1209_U83 , P2_R1209_U84 , P2_R1209_U85 , P2_R1209_U86 , P2_R1209_U87;
wire P2_R1209_U88 , P2_R1209_U89 , P2_R1209_U90 , P2_R1209_U91 , P2_R1209_U92 , P2_R1209_U93 , P2_R1209_U94 , P2_R1209_U95 , P2_R1209_U96 , P2_R1209_U97;
wire P2_R1209_U98 , P2_R1209_U99 , P2_R1209_U100 , P2_R1209_U101 , P2_R1209_U102 , P2_R1209_U103 , P2_R1209_U104 , P2_R1209_U105 , P2_R1209_U106 , P2_R1209_U107;
wire P2_R1209_U108 , P2_R1209_U109 , P2_R1209_U110 , P2_R1209_U111 , P2_R1209_U112 , P2_R1209_U113 , P2_R1209_U114 , P2_R1209_U115 , P2_R1209_U116 , P2_R1209_U117;
wire P2_R1209_U118 , P2_R1209_U119 , P2_R1209_U120 , P2_R1209_U121 , P2_R1209_U122 , P2_R1209_U123 , P2_R1209_U124 , P2_R1209_U125 , P2_R1209_U126 , P2_R1209_U127;
wire P2_R1209_U128 , P2_R1209_U129 , P2_R1209_U130 , P2_R1209_U131 , P2_R1209_U132 , P2_R1209_U133 , P2_R1209_U134 , P2_R1209_U135 , P2_R1209_U136 , P2_R1209_U137;
wire P2_R1209_U138 , P2_R1209_U139 , P2_R1209_U140 , P2_R1209_U141 , P2_R1209_U142 , P2_R1209_U143 , P2_R1209_U144 , P2_R1209_U145 , P2_R1209_U146 , P2_R1209_U147;
wire P2_R1209_U148 , P2_R1209_U149 , P2_R1209_U150 , P2_R1209_U151 , P2_R1209_U152 , P2_R1209_U153 , P2_R1209_U154 , P2_R1209_U155 , P2_R1209_U156 , P2_R1209_U157;
wire P2_R1209_U158 , P2_R1209_U159 , P2_R1209_U160 , P2_R1209_U161 , P2_R1209_U162 , P2_R1209_U163 , P2_R1209_U164 , P2_R1209_U165 , P2_R1209_U166 , P2_R1209_U167;
wire P2_R1209_U168 , P2_R1209_U169 , P2_R1209_U170 , P2_R1209_U171 , P2_R1209_U172 , P2_R1209_U173 , P2_R1209_U174 , P2_R1209_U175 , P2_R1209_U176 , P2_R1209_U177;
wire P2_R1209_U178 , P2_R1209_U179 , P2_R1209_U180 , P2_R1209_U181 , P2_R1209_U182 , P2_R1209_U183 , P2_R1209_U184 , P2_R1209_U185 , P2_R1209_U186 , P2_R1209_U187;
wire P2_R1209_U188 , P2_R1209_U189 , P2_R1209_U190 , P2_R1209_U191 , P2_R1209_U192 , P2_R1209_U193 , P2_R1209_U194 , P2_R1209_U195 , P2_R1209_U196 , P2_R1209_U197;
wire P2_R1209_U198 , P2_R1209_U199 , P2_R1209_U200 , P2_R1209_U201 , P2_R1209_U202 , P2_R1209_U203 , P2_R1209_U204 , P2_R1209_U205 , P2_R1209_U206 , P2_R1209_U207;
wire P2_R1209_U208 , P2_R1209_U209 , P2_R1209_U210 , P2_R1209_U211 , P2_R1209_U212 , P2_R1209_U213 , P2_R1209_U214 , P2_R1209_U215 , P2_R1209_U216 , P2_R1209_U217;
wire P2_R1209_U218 , P2_R1209_U219 , P2_R1209_U220 , P2_R1209_U221 , P2_R1209_U222 , P2_R1209_U223 , P2_R1209_U224 , P2_R1209_U225 , P2_R1209_U226 , P2_R1209_U227;
wire P2_R1209_U228 , P2_R1209_U229 , P2_R1209_U230 , P2_R1209_U231 , P2_R1209_U232 , P2_R1209_U233 , P2_R1209_U234 , P2_R1209_U235 , P2_R1209_U236 , P2_R1209_U237;
wire P2_R1209_U238 , P2_R1209_U239 , P2_R1209_U240 , P2_R1209_U241 , P2_R1209_U242 , P2_R1209_U243 , P2_R1209_U244 , P2_R1209_U245 , P2_R1209_U246 , P2_R1209_U247;
wire P2_R1209_U248 , P2_R1209_U249 , P2_R1209_U250 , P2_R1209_U251 , P2_R1209_U252 , P2_R1209_U253 , P2_R1209_U254 , P2_R1209_U255 , P2_R1209_U256 , P2_R1209_U257;
wire P2_R1209_U258 , P2_R1209_U259 , P2_R1209_U260 , P2_R1209_U261 , P2_R1209_U262 , P2_R1209_U263 , P2_R1209_U264 , P2_R1209_U265 , P2_R1209_U266 , P2_R1209_U267;
wire P2_R1209_U268 , P2_R1209_U269 , P2_R1209_U270 , P2_R1209_U271 , P2_R1209_U272 , P2_R1209_U273 , P2_R1209_U274 , P2_R1209_U275 , P2_R1209_U276 , P2_R1209_U277;
wire P2_R1209_U278 , P2_R1209_U279 , P2_R1209_U280 , P2_R1209_U281 , P2_R1209_U282 , P2_R1209_U283 , P2_R1209_U284 , P2_R1209_U285 , P2_R1209_U286 , P2_R1209_U287;
wire P2_R1209_U288 , P2_R1209_U289 , P2_R1209_U290 , P2_R1209_U291 , P2_R1209_U292 , P2_R1209_U293 , P2_R1209_U294 , P2_R1209_U295 , P2_R1209_U296 , P2_R1209_U297;
wire P2_R1209_U298 , P2_R1209_U299 , P2_R1209_U300 , P2_R1209_U301 , P2_R1209_U302 , P2_R1209_U303 , P2_R1209_U304 , P2_R1209_U305 , P2_R1209_U306 , P2_R1209_U307;
wire P2_R1209_U308 , P2_R1170_U4 , P2_R1170_U5 , P2_R1170_U6 , P2_R1170_U7 , P2_R1170_U8 , P2_R1170_U9 , P2_R1170_U10 , P2_R1170_U11 , P2_R1170_U12;
wire P2_R1170_U13 , P2_R1170_U14 , P2_R1170_U15 , P2_R1170_U16 , P2_R1170_U17 , P2_R1170_U18 , P2_R1170_U19 , P2_R1170_U20 , P2_R1170_U21 , P2_R1170_U22;
wire P2_R1170_U23 , P2_R1170_U24 , P2_R1170_U25 , P2_R1170_U26 , P2_R1170_U27 , P2_R1170_U28 , P2_R1170_U29 , P2_R1170_U30 , P2_R1170_U31 , P2_R1170_U32;
wire P2_R1170_U33 , P2_R1170_U34 , P2_R1170_U35 , P2_R1170_U36 , P2_R1170_U37 , P2_R1170_U38 , P2_R1170_U39 , P2_R1170_U40 , P2_R1170_U41 , P2_R1170_U42;
wire P2_R1170_U43 , P2_R1170_U44 , P2_R1170_U45 , P2_R1170_U46 , P2_R1170_U47 , P2_R1170_U48 , P2_R1170_U49 , P2_R1170_U50 , P2_R1170_U51 , P2_R1170_U52;
wire P2_R1170_U53 , P2_R1170_U54 , P2_R1170_U55 , P2_R1170_U56 , P2_R1170_U57 , P2_R1170_U58 , P2_R1170_U59 , P2_R1170_U60 , P2_R1170_U61 , P2_R1170_U62;
wire P2_R1170_U63 , P2_R1170_U64 , P2_R1170_U65 , P2_R1170_U66 , P2_R1170_U67 , P2_R1170_U68 , P2_R1170_U69 , P2_R1170_U70 , P2_R1170_U71 , P2_R1170_U72;
wire P2_R1170_U73 , P2_R1170_U74 , P2_R1170_U75 , P2_R1170_U76 , P2_R1170_U77 , P2_R1170_U78 , P2_R1170_U79 , P2_R1170_U80 , P2_R1170_U81 , P2_R1170_U82;
wire P2_R1170_U83 , P2_R1170_U84 , P2_R1170_U85 , P2_R1170_U86 , P2_R1170_U87 , P2_R1170_U88 , P2_R1170_U89 , P2_R1170_U90 , P2_R1170_U91 , P2_R1170_U92;
wire P2_R1170_U93 , P2_R1170_U94 , P2_R1170_U95 , P2_R1170_U96 , P2_R1170_U97 , P2_R1170_U98 , P2_R1170_U99 , P2_R1170_U100 , P2_R1170_U101 , P2_R1170_U102;
wire P2_R1170_U103 , P2_R1170_U104 , P2_R1170_U105 , P2_R1170_U106 , P2_R1170_U107 , P2_R1170_U108 , P2_R1170_U109 , P2_R1170_U110 , P2_R1170_U111 , P2_R1170_U112;
wire P2_R1170_U113 , P2_R1170_U114 , P2_R1170_U115 , P2_R1170_U116 , P2_R1170_U117 , P2_R1170_U118 , P2_R1170_U119 , P2_R1170_U120 , P2_R1170_U121 , P2_R1170_U122;
wire P2_R1170_U123 , P2_R1170_U124 , P2_R1170_U125 , P2_R1170_U126 , P2_R1170_U127 , P2_R1170_U128 , P2_R1170_U129 , P2_R1170_U130 , P2_R1170_U131 , P2_R1170_U132;
wire P2_R1170_U133 , P2_R1170_U134 , P2_R1170_U135 , P2_R1170_U136 , P2_R1170_U137 , P2_R1170_U138 , P2_R1170_U139 , P2_R1170_U140 , P2_R1170_U141 , P2_R1170_U142;
wire P2_R1170_U143 , P2_R1170_U144 , P2_R1170_U145 , P2_R1170_U146 , P2_R1170_U147 , P2_R1170_U148 , P2_R1170_U149 , P2_R1170_U150 , P2_R1170_U151 , P2_R1170_U152;
wire P2_R1170_U153 , P2_R1170_U154 , P2_R1170_U155 , P2_R1170_U156 , P2_R1170_U157 , P2_R1170_U158 , P2_R1170_U159 , P2_R1170_U160 , P2_R1170_U161 , P2_R1170_U162;
wire P2_R1170_U163 , P2_R1170_U164 , P2_R1170_U165 , P2_R1170_U166 , P2_R1170_U167 , P2_R1170_U168 , P2_R1170_U169 , P2_R1170_U170 , P2_R1170_U171 , P2_R1170_U172;
wire P2_R1170_U173 , P2_R1170_U174 , P2_R1170_U175 , P2_R1170_U176 , P2_R1170_U177 , P2_R1170_U178 , P2_R1170_U179 , P2_R1170_U180 , P2_R1170_U181 , P2_R1170_U182;
wire P2_R1170_U183 , P2_R1170_U184 , P2_R1170_U185 , P2_R1170_U186 , P2_R1170_U187 , P2_R1170_U188 , P2_R1170_U189 , P2_R1170_U190 , P2_R1170_U191 , P2_R1170_U192;
wire P2_R1170_U193 , P2_R1170_U194 , P2_R1170_U195 , P2_R1170_U196 , P2_R1170_U197 , P2_R1170_U198 , P2_R1170_U199 , P2_R1170_U200 , P2_R1170_U201 , P2_R1170_U202;
wire P2_R1170_U203 , P2_R1170_U204 , P2_R1170_U205 , P2_R1170_U206 , P2_R1170_U207 , P2_R1170_U208 , P2_R1170_U209 , P2_R1170_U210 , P2_R1170_U211 , P2_R1170_U212;
wire P2_R1170_U213 , P2_R1170_U214 , P2_R1170_U215 , P2_R1170_U216 , P2_R1170_U217 , P2_R1170_U218 , P2_R1170_U219 , P2_R1170_U220 , P2_R1170_U221 , P2_R1170_U222;
wire P2_R1170_U223 , P2_R1170_U224 , P2_R1170_U225 , P2_R1170_U226 , P2_R1170_U227 , P2_R1170_U228 , P2_R1170_U229 , P2_R1170_U230 , P2_R1170_U231 , P2_R1170_U232;
wire P2_R1170_U233 , P2_R1170_U234 , P2_R1170_U235 , P2_R1170_U236 , P2_R1170_U237 , P2_R1170_U238 , P2_R1170_U239 , P2_R1170_U240 , P2_R1170_U241 , P2_R1170_U242;
wire P2_R1170_U243 , P2_R1170_U244 , P2_R1170_U245 , P2_R1170_U246 , P2_R1170_U247 , P2_R1170_U248 , P2_R1170_U249 , P2_R1170_U250 , P2_R1170_U251 , P2_R1170_U252;
wire P2_R1170_U253 , P2_R1170_U254 , P2_R1170_U255 , P2_R1170_U256 , P2_R1170_U257 , P2_R1170_U258 , P2_R1170_U259 , P2_R1170_U260 , P2_R1170_U261 , P2_R1170_U262;
wire P2_R1170_U263 , P2_R1170_U264 , P2_R1170_U265 , P2_R1170_U266 , P2_R1170_U267 , P2_R1170_U268 , P2_R1170_U269 , P2_R1170_U270 , P2_R1170_U271 , P2_R1170_U272;
wire P2_R1170_U273 , P2_R1170_U274 , P2_R1170_U275 , P2_R1170_U276 , P2_R1170_U277 , P2_R1170_U278 , P2_R1170_U279 , P2_R1170_U280 , P2_R1170_U281 , P2_R1170_U282;
wire P2_R1170_U283 , P2_R1170_U284 , P2_R1170_U285 , P2_R1170_U286 , P2_R1170_U287 , P2_R1170_U288 , P2_R1170_U289 , P2_R1170_U290 , P2_R1170_U291 , P2_R1170_U292;
wire P2_R1170_U293 , P2_R1170_U294 , P2_R1170_U295 , P2_R1170_U296 , P2_R1170_U297 , P2_R1170_U298 , P2_R1170_U299 , P2_R1170_U300 , P2_R1170_U301 , P2_R1170_U302;
wire P2_R1170_U303 , P2_R1170_U304 , P2_R1170_U305 , P2_R1170_U306 , P2_R1170_U307 , P2_R1170_U308 , P2_R1275_U6 , P2_R1275_U7 , P2_R1275_U8 , P2_R1275_U9;
wire P2_R1275_U10 , P2_R1275_U11 , P2_R1275_U12 , P2_R1275_U13 , P2_R1275_U14 , P2_R1275_U15 , P2_R1275_U16 , P2_R1275_U17 , P2_R1275_U18 , P2_R1275_U19;
wire P2_R1275_U20 , P2_R1275_U21 , P2_R1275_U22 , P2_R1275_U23 , P2_R1275_U24 , P2_R1275_U25 , P2_R1275_U26 , P2_R1275_U27 , P2_R1275_U28 , P2_R1275_U29;
wire P2_R1275_U30 , P2_R1275_U31 , P2_R1275_U32 , P2_R1275_U33 , P2_R1275_U34 , P2_R1275_U35 , P2_R1275_U36 , P2_R1275_U37 , P2_R1275_U38 , P2_R1275_U39;
wire P2_R1275_U40 , P2_R1275_U41 , P2_R1275_U42 , P2_R1275_U43 , P2_R1275_U44 , P2_R1275_U45 , P2_R1275_U46 , P2_R1275_U47 , P2_R1275_U48 , P2_R1275_U49;
wire P2_R1275_U50 , P2_R1275_U51 , P2_R1275_U52 , P2_R1275_U53 , P2_R1275_U54 , P2_R1275_U55 , P2_R1275_U56 , P2_R1275_U57 , P2_R1275_U58 , P2_R1275_U59;
wire P2_R1275_U60 , P2_R1275_U61 , P2_R1275_U62 , P2_R1275_U63 , P2_R1275_U64 , P2_R1275_U65 , P2_R1275_U66 , P2_R1275_U67 , P2_R1275_U68 , P2_R1275_U69;
wire P2_R1275_U70 , P2_R1275_U71 , P2_R1275_U72 , P2_R1275_U73 , P2_R1275_U74 , P2_R1275_U75 , P2_R1275_U76 , P2_R1275_U77 , P2_R1275_U78 , P2_R1275_U79;
wire P2_R1275_U80 , P2_R1275_U81 , P2_R1275_U82 , P2_R1275_U83 , P2_R1275_U84 , P2_R1275_U85 , P2_R1275_U86 , P2_R1275_U87 , P2_R1275_U88 , P2_R1275_U89;
wire P2_R1275_U90 , P2_R1275_U91 , P2_R1275_U92 , P2_R1275_U93 , P2_R1275_U94 , P2_R1275_U95 , P2_R1275_U96 , P2_R1275_U97 , P2_R1275_U98 , P2_R1275_U99;
wire P2_R1275_U100 , P2_R1275_U101 , P2_R1275_U102 , P2_R1275_U103 , P2_R1275_U104 , P2_R1275_U105 , P2_R1275_U106 , P2_R1275_U107 , P2_R1275_U108 , P2_R1275_U109;
wire P2_R1275_U110 , P2_R1275_U111 , P2_R1275_U112 , P2_R1275_U113 , P2_R1275_U114 , P2_R1275_U115 , P2_R1275_U116 , P2_R1275_U117 , P2_R1275_U118 , P2_R1275_U119;
wire P2_R1275_U120 , P2_R1275_U121 , P2_R1275_U122 , P2_R1275_U123 , P2_R1275_U124 , P2_R1275_U125 , P2_R1275_U126 , P2_R1275_U127 , P2_R1275_U128 , P2_R1275_U129;
wire P2_R1275_U130 , P2_R1275_U131 , P2_R1275_U132 , P2_R1275_U133 , P2_R1275_U134 , P2_R1275_U135 , P2_R1275_U136 , P2_R1275_U137 , P2_R1275_U138 , P2_R1275_U139;
wire P2_R1275_U140 , P2_R1275_U141 , P2_R1275_U142 , P2_R1275_U143 , P2_R1275_U144 , P2_R1275_U145 , P2_R1275_U146 , P2_R1275_U147 , P2_R1275_U148 , P2_R1275_U149;
wire P2_R1275_U150 , P2_R1275_U151 , P2_R1275_U152 , P2_R1275_U153 , P2_R1275_U154 , P2_R1275_U155 , P2_R1275_U156 , P2_R1275_U157 , P2_R1275_U158 , P2_R1275_U159;
wire P2_R1179_U6 , P2_R1179_U7 , P2_R1179_U8 , P2_R1179_U9 , P2_R1179_U10 , P2_R1179_U11 , P2_R1179_U12 , P2_R1179_U13 , P2_R1179_U14 , P2_R1179_U15;
wire P2_R1179_U16 , P2_R1179_U17 , P2_R1179_U18 , P2_R1179_U19 , P2_R1179_U20 , P2_R1179_U21 , P2_R1179_U22 , P2_R1179_U23 , P2_R1179_U24 , P2_R1179_U25;
wire P2_R1179_U26 , P2_R1179_U27 , P2_R1179_U28 , P2_R1179_U29 , P2_R1179_U30 , P2_R1179_U31 , P2_R1179_U32 , P2_R1179_U33 , P2_R1179_U34 , P2_R1179_U35;
wire P2_R1179_U36 , P2_R1179_U37 , P2_R1179_U38 , P2_R1179_U39 , P2_R1179_U40 , P2_R1179_U41 , P2_R1179_U42 , P2_R1179_U43 , P2_R1179_U44 , P2_R1179_U45;
wire P2_R1179_U46 , P2_R1179_U47 , P2_R1179_U48 , P2_R1179_U49 , P2_R1179_U50 , P2_R1179_U51 , P2_R1179_U52 , P2_R1179_U53 , P2_R1179_U54 , P2_R1179_U55;
wire P2_R1179_U56 , P2_R1179_U57 , P2_R1179_U58 , P2_R1179_U59 , P2_R1179_U60 , P2_R1179_U61 , P2_R1179_U62 , P2_R1179_U63 , P2_R1179_U64 , P2_R1179_U65;
wire P2_R1179_U66 , P2_R1179_U67 , P2_R1179_U68 , P2_R1179_U69 , P2_R1179_U70 , P2_R1179_U71 , P2_R1179_U72 , P2_R1179_U73 , P2_R1179_U74 , P2_R1179_U75;
wire P2_R1179_U76 , P2_R1179_U77 , P2_R1179_U78 , P2_R1179_U79 , P2_R1179_U80 , P2_R1179_U81 , P2_R1179_U82 , P2_R1179_U83 , P2_R1179_U84 , P2_R1179_U85;
wire P2_R1179_U86 , P2_R1179_U87 , P2_R1179_U88 , P2_R1179_U89 , P2_R1179_U90 , P2_R1179_U91 , P2_R1179_U92 , P2_R1179_U93 , P2_R1179_U94 , P2_R1179_U95;
wire P2_R1179_U96 , P2_R1179_U97 , P2_R1179_U98 , P2_R1179_U99 , P2_R1179_U100 , P2_R1179_U101 , P2_R1179_U102 , P2_R1179_U103 , P2_R1179_U104 , P2_R1179_U105;
wire P2_R1179_U106 , P2_R1179_U107 , P2_R1179_U108 , P2_R1179_U109 , P2_R1179_U110 , P2_R1179_U111 , P2_R1179_U112 , P2_R1179_U113 , P2_R1179_U114 , P2_R1179_U115;
wire P2_R1179_U116 , P2_R1179_U117 , P2_R1179_U118 , P2_R1179_U119 , P2_R1179_U120 , P2_R1179_U121 , P2_R1179_U122 , P2_R1179_U123 , P2_R1179_U124 , P2_R1179_U125;
wire P2_R1179_U126 , P2_R1179_U127 , P2_R1179_U128 , P2_R1179_U129 , P2_R1179_U130 , P2_R1179_U131 , P2_R1179_U132 , P2_R1179_U133 , P2_R1179_U134 , P2_R1179_U135;
wire P2_R1179_U136 , P2_R1179_U137 , P2_R1179_U138 , P2_R1179_U139 , P2_R1179_U140 , P2_R1179_U141 , P2_R1179_U142 , P2_R1179_U143 , P2_R1179_U144 , P2_R1179_U145;
wire P2_R1179_U146 , P2_R1179_U147 , P2_R1179_U148 , P2_R1179_U149 , P2_R1179_U150 , P2_R1179_U151 , P2_R1179_U152 , P2_R1179_U153 , P2_R1179_U154 , P2_R1179_U155;
wire P2_R1179_U156 , P2_R1179_U157 , P2_R1179_U158 , P2_R1179_U159 , P2_R1179_U160 , P2_R1179_U161 , P2_R1179_U162 , P2_R1179_U163 , P2_R1179_U164 , P2_R1179_U165;
wire P2_R1179_U166 , P2_R1179_U167 , P2_R1179_U168 , P2_R1179_U169 , P2_R1179_U170 , P2_R1179_U171 , P2_R1179_U172 , P2_R1179_U173 , P2_R1179_U174 , P2_R1179_U175;
wire P2_R1179_U176 , P2_R1179_U177 , P2_R1179_U178 , P2_R1179_U179 , P2_R1179_U180 , P2_R1179_U181 , P2_R1179_U182 , P2_R1179_U183 , P2_R1179_U184 , P2_R1179_U185;
wire P2_R1179_U186 , P2_R1179_U187 , P2_R1179_U188 , P2_R1179_U189 , P2_R1179_U190 , P2_R1179_U191 , P2_R1179_U192 , P2_R1179_U193 , P2_R1179_U194 , P2_R1179_U195;
wire P2_R1179_U196 , P2_R1179_U197 , P2_R1179_U198 , P2_R1179_U199 , P2_R1179_U200 , P2_R1179_U201 , P2_R1179_U202 , P2_R1179_U203 , P2_R1179_U204 , P2_R1179_U205;
wire P2_R1179_U206 , P2_R1179_U207 , P2_R1179_U208 , P2_R1179_U209 , P2_R1179_U210 , P2_R1179_U211 , P2_R1179_U212 , P2_R1179_U213 , P2_R1179_U214 , P2_R1179_U215;
wire P2_R1179_U216 , P2_R1179_U217 , P2_R1179_U218 , P2_R1179_U219 , P2_R1179_U220 , P2_R1179_U221 , P2_R1179_U222 , P2_R1179_U223 , P2_R1179_U224 , P2_R1179_U225;
wire P2_R1179_U226 , P2_R1179_U227 , P2_R1179_U228 , P2_R1179_U229 , P2_R1179_U230 , P2_R1179_U231 , P2_R1179_U232 , P2_R1179_U233 , P2_R1179_U234 , P2_R1179_U235;
wire P2_R1179_U236 , P2_R1179_U237 , P2_R1179_U238 , P2_R1179_U239 , P2_R1179_U240 , P2_R1179_U241 , P2_R1179_U242 , P2_R1179_U243 , P2_R1179_U244 , P2_R1179_U245;
wire P2_R1179_U246 , P2_R1179_U247 , P2_R1179_U248 , P2_R1179_U249 , P2_R1179_U250 , P2_R1179_U251 , P2_R1179_U252 , P2_R1179_U253 , P2_R1179_U254 , P2_R1179_U255;
wire P2_R1179_U256 , P2_R1179_U257 , P2_R1179_U258 , P2_R1179_U259 , P2_R1179_U260 , P2_R1179_U261 , P2_R1179_U262 , P2_R1179_U263 , P2_R1179_U264 , P2_R1179_U265;
wire P2_R1179_U266 , P2_R1179_U267 , P2_R1179_U268 , P2_R1179_U269 , P2_R1179_U270 , P2_R1179_U271 , P2_R1179_U272 , P2_R1179_U273 , P2_R1179_U274 , P2_R1179_U275;
wire P2_R1179_U276 , P2_R1179_U277 , P2_R1179_U278 , P2_R1179_U279 , P2_R1179_U280 , P2_R1179_U281 , P2_R1179_U282 , P2_R1179_U283 , P2_R1179_U284 , P2_R1179_U285;
wire P2_R1179_U286 , P2_R1179_U287 , P2_R1179_U288 , P2_R1179_U289 , P2_R1179_U290 , P2_R1179_U291 , P2_R1179_U292 , P2_R1179_U293 , P2_R1179_U294 , P2_R1179_U295;
wire P2_R1179_U296 , P2_R1179_U297 , P2_R1179_U298 , P2_R1179_U299 , P2_R1179_U300 , P2_R1179_U301 , P2_R1179_U302 , P2_R1179_U303 , P2_R1179_U304 , P2_R1179_U305;
wire P2_R1179_U306 , P2_R1179_U307 , P2_R1179_U308 , P2_R1179_U309 , P2_R1179_U310 , P2_R1179_U311 , P2_R1179_U312 , P2_R1179_U313 , P2_R1179_U314 , P2_R1179_U315;
wire P2_R1179_U316 , P2_R1179_U317 , P2_R1179_U318 , P2_R1179_U319 , P2_R1179_U320 , P2_R1179_U321 , P2_R1179_U322 , P2_R1179_U323 , P2_R1179_U324 , P2_R1179_U325;
wire P2_R1179_U326 , P2_R1179_U327 , P2_R1179_U328 , P2_R1179_U329 , P2_R1179_U330 , P2_R1179_U331 , P2_R1179_U332 , P2_R1179_U333 , P2_R1179_U334 , P2_R1179_U335;
wire P2_R1179_U336 , P2_R1179_U337 , P2_R1179_U338 , P2_R1179_U339 , P2_R1179_U340 , P2_R1179_U341 , P2_R1179_U342 , P2_R1179_U343 , P2_R1179_U344 , P2_R1179_U345;
wire P2_R1179_U346 , P2_R1179_U347 , P2_R1179_U348 , P2_R1179_U349 , P2_R1179_U350 , P2_R1179_U351 , P2_R1179_U352 , P2_R1179_U353 , P2_R1179_U354 , P2_R1179_U355;
wire P2_R1179_U356 , P2_R1179_U357 , P2_R1179_U358 , P2_R1179_U359 , P2_R1179_U360 , P2_R1179_U361 , P2_R1179_U362 , P2_R1179_U363 , P2_R1179_U364 , P2_R1179_U365;
wire P2_R1179_U366 , P2_R1179_U367 , P2_R1179_U368 , P2_R1179_U369 , P2_R1179_U370 , P2_R1179_U371 , P2_R1179_U372 , P2_R1179_U373 , P2_R1179_U374 , P2_R1179_U375;
wire P2_R1179_U376 , P2_R1179_U377 , P2_R1179_U378 , P2_R1179_U379 , P2_R1179_U380 , P2_R1179_U381 , P2_R1179_U382 , P2_R1179_U383 , P2_R1179_U384 , P2_R1179_U385;
wire P2_R1179_U386 , P2_R1179_U387 , P2_R1179_U388 , P2_R1179_U389 , P2_R1179_U390 , P2_R1179_U391 , P2_R1179_U392 , P2_R1179_U393 , P2_R1179_U394 , P2_R1179_U395;
wire P2_R1179_U396 , P2_R1179_U397 , P2_R1179_U398 , P2_R1179_U399 , P2_R1179_U400 , P2_R1179_U401 , P2_R1179_U402 , P2_R1179_U403 , P2_R1179_U404 , P2_R1179_U405;
wire P2_R1179_U406 , P2_R1179_U407 , P2_R1179_U408 , P2_R1179_U409 , P2_R1179_U410 , P2_R1179_U411 , P2_R1179_U412 , P2_R1179_U413 , P2_R1179_U414 , P2_R1179_U415;
wire P2_R1179_U416 , P2_R1179_U417 , P2_R1179_U418 , P2_R1179_U419 , P2_R1179_U420 , P2_R1179_U421 , P2_R1179_U422 , P2_R1179_U423 , P2_R1179_U424 , P2_R1179_U425;
wire P2_R1179_U426 , P2_R1179_U427 , P2_R1179_U428 , P2_R1179_U429 , P2_R1179_U430 , P2_R1179_U431 , P2_R1179_U432 , P2_R1179_U433 , P2_R1179_U434 , P2_R1179_U435;
wire P2_R1179_U436 , P2_R1179_U437 , P2_R1179_U438 , P2_R1179_U439 , P2_R1179_U440 , P2_R1179_U441 , P2_R1179_U442 , P2_R1179_U443 , P2_R1179_U444 , P2_R1179_U445;
wire P2_R1179_U446 , P2_R1179_U447 , P2_R1179_U448 , P2_R1179_U449 , P2_R1179_U450 , P2_R1179_U451 , P2_R1179_U452 , P2_R1179_U453 , P2_R1179_U454 , P2_R1179_U455;
wire P2_R1179_U456 , P2_R1179_U457 , P2_R1179_U458 , P2_R1179_U459 , P2_R1179_U460 , P2_R1179_U461 , P2_R1179_U462 , P2_R1179_U463 , P2_R1179_U464 , P2_R1179_U465;
wire P2_R1179_U466 , P2_R1179_U467 , P2_R1179_U468 , P2_R1179_U469 , P2_R1179_U470 , P2_R1179_U471 , P2_R1179_U472 , P2_R1179_U473 , P2_R1179_U474 , P2_R1179_U475;
wire P2_R1179_U476 , P2_R1179_U477 , P2_R1179_U478 , P2_R1215_U4 , P2_R1215_U5 , P2_R1215_U6 , P2_R1215_U7 , P2_R1215_U8 , P2_R1215_U9 , P2_R1215_U10;
wire P2_R1215_U11 , P2_R1215_U12 , P2_R1215_U13 , P2_R1215_U14 , P2_R1215_U15 , P2_R1215_U16 , P2_R1215_U17 , P2_R1215_U18 , P2_R1215_U19 , P2_R1215_U20;
wire P2_R1215_U21 , P2_R1215_U22 , P2_R1215_U23 , P2_R1215_U24 , P2_R1215_U25 , P2_R1215_U26 , P2_R1215_U27 , P2_R1215_U28 , P2_R1215_U29 , P2_R1215_U30;
wire P2_R1215_U31 , P2_R1215_U32 , P2_R1215_U33 , P2_R1215_U34 , P2_R1215_U35 , P2_R1215_U36 , P2_R1215_U37 , P2_R1215_U38 , P2_R1215_U39 , P2_R1215_U40;
wire P2_R1215_U41 , P2_R1215_U42 , P2_R1215_U43 , P2_R1215_U44 , P2_R1215_U45 , P2_R1215_U46 , P2_R1215_U47 , P2_R1215_U48 , P2_R1215_U49 , P2_R1215_U50;
wire P2_R1215_U51 , P2_R1215_U52 , P2_R1215_U53 , P2_R1215_U54 , P2_R1215_U55 , P2_R1215_U56 , P2_R1215_U57 , P2_R1215_U58 , P2_R1215_U59 , P2_R1215_U60;
wire P2_R1215_U61 , P2_R1215_U62 , P2_R1215_U63 , P2_R1215_U64 , P2_R1215_U65 , P2_R1215_U66 , P2_R1215_U67 , P2_R1215_U68 , P2_R1215_U69 , P2_R1215_U70;
wire P2_R1215_U71 , P2_R1215_U72 , P2_R1215_U73 , P2_R1215_U74 , P2_R1215_U75 , P2_R1215_U76 , P2_R1215_U77 , P2_R1215_U78 , P2_R1215_U79 , P2_R1215_U80;
wire P2_R1215_U81 , P2_R1215_U82 , P2_R1215_U83 , P2_R1215_U84 , P2_R1215_U85 , P2_R1215_U86 , P2_R1215_U87 , P2_R1215_U88 , P2_R1215_U89 , P2_R1215_U90;
wire P2_R1215_U91 , P2_R1215_U92 , P2_R1215_U93 , P2_R1215_U94 , P2_R1215_U95 , P2_R1215_U96 , P2_R1215_U97 , P2_R1215_U98 , P2_R1215_U99 , P2_R1215_U100;
wire P2_R1215_U101 , P2_R1215_U102 , P2_R1215_U103 , P2_R1215_U104 , P2_R1215_U105 , P2_R1215_U106 , P2_R1215_U107 , P2_R1215_U108 , P2_R1215_U109 , P2_R1215_U110;
wire P2_R1215_U111 , P2_R1215_U112 , P2_R1215_U113 , P2_R1215_U114 , P2_R1215_U115 , P2_R1215_U116 , P2_R1215_U117 , P2_R1215_U118 , P2_R1215_U119 , P2_R1215_U120;
wire P2_R1215_U121 , P2_R1215_U122 , P2_R1215_U123 , P2_R1215_U124 , P2_R1215_U125 , P2_R1215_U126 , P2_R1215_U127 , P2_R1215_U128 , P2_R1215_U129 , P2_R1215_U130;
wire P2_R1215_U131 , P2_R1215_U132 , P2_R1215_U133 , P2_R1215_U134 , P2_R1215_U135 , P2_R1215_U136 , P2_R1215_U137 , P2_R1215_U138 , P2_R1215_U139 , P2_R1215_U140;
wire P2_R1215_U141 , P2_R1215_U142 , P2_R1215_U143 , P2_R1215_U144 , P2_R1215_U145 , P2_R1215_U146 , P2_R1215_U147 , P2_R1215_U148 , P2_R1215_U149 , P2_R1215_U150;
wire P2_R1215_U151 , P2_R1215_U152 , P2_R1215_U153 , P2_R1215_U154 , P2_R1215_U155 , P2_R1215_U156 , P2_R1215_U157 , P2_R1215_U158 , P2_R1215_U159 , P2_R1215_U160;
wire P2_R1215_U161 , P2_R1215_U162 , P2_R1215_U163 , P2_R1215_U164 , P2_R1215_U165 , P2_R1215_U166 , P2_R1215_U167 , P2_R1215_U168 , P2_R1215_U169 , P2_R1215_U170;
wire P2_R1215_U171 , P2_R1215_U172 , P2_R1215_U173 , P2_R1215_U174 , P2_R1215_U175 , P2_R1215_U176 , P2_R1215_U177 , P2_R1215_U178 , P2_R1215_U179 , P2_R1215_U180;
wire P2_R1215_U181 , P2_R1215_U182 , P2_R1215_U183 , P2_R1215_U184 , P2_R1215_U185 , P2_R1215_U186 , P2_R1215_U187 , P2_R1215_U188 , P2_R1215_U189 , P2_R1215_U190;
wire P2_R1215_U191 , P2_R1215_U192 , P2_R1215_U193 , P2_R1215_U194 , P2_R1215_U195 , P2_R1215_U196 , P2_R1215_U197 , P2_R1215_U198 , P2_R1215_U199 , P2_R1215_U200;
wire P2_R1215_U201 , P2_R1215_U202 , P2_R1215_U203 , P2_R1215_U204 , P2_R1215_U205 , P2_R1215_U206 , P2_R1215_U207 , P2_R1215_U208 , P2_R1215_U209 , P2_R1215_U210;
wire P2_R1215_U211 , P2_R1215_U212 , P2_R1215_U213 , P2_R1215_U214 , P2_R1215_U215 , P2_R1215_U216 , P2_R1215_U217 , P2_R1215_U218 , P2_R1215_U219 , P2_R1215_U220;
wire P2_R1215_U221 , P2_R1215_U222 , P2_R1215_U223 , P2_R1215_U224 , P2_R1215_U225 , P2_R1215_U226 , P2_R1215_U227 , P2_R1215_U228 , P2_R1215_U229 , P2_R1215_U230;
wire P2_R1215_U231 , P2_R1215_U232 , P2_R1215_U233 , P2_R1215_U234 , P2_R1215_U235 , P2_R1215_U236 , P2_R1215_U237 , P2_R1215_U238 , P2_R1215_U239 , P2_R1215_U240;
wire P2_R1215_U241 , P2_R1215_U242 , P2_R1215_U243 , P2_R1215_U244 , P2_R1215_U245 , P2_R1215_U246 , P2_R1215_U247 , P2_R1215_U248 , P2_R1215_U249 , P2_R1215_U250;
wire P2_R1215_U251 , P2_R1215_U252 , P2_R1215_U253 , P2_R1215_U254 , P2_R1215_U255 , P2_R1215_U256 , P2_R1215_U257 , P2_R1215_U258 , P2_R1215_U259 , P2_R1215_U260;
wire P2_R1215_U261 , P2_R1215_U262 , P2_R1215_U263 , P2_R1215_U264 , P2_R1215_U265 , P2_R1215_U266 , P2_R1215_U267 , P2_R1215_U268 , P2_R1215_U269 , P2_R1215_U270;
wire P2_R1215_U271 , P2_R1215_U272 , P2_R1215_U273 , P2_R1215_U274 , P2_R1215_U275 , P2_R1215_U276 , P2_R1215_U277 , P2_R1215_U278 , P2_R1215_U279 , P2_R1215_U280;
wire P2_R1215_U281 , P2_R1215_U282 , P2_R1215_U283 , P2_R1215_U284 , P2_R1215_U285 , P2_R1215_U286 , P2_R1215_U287 , P2_R1215_U288 , P2_R1215_U289 , P2_R1215_U290;
wire P2_R1215_U291 , P2_R1215_U292 , P2_R1215_U293 , P2_R1215_U294 , P2_R1215_U295 , P2_R1215_U296 , P2_R1215_U297 , P2_R1215_U298 , P2_R1215_U299 , P2_R1215_U300;
wire P2_R1215_U301 , P2_R1215_U302 , P2_R1215_U303 , P2_R1215_U304 , P2_R1215_U305 , P2_R1215_U306 , P2_R1215_U307 , P2_R1215_U308 , P2_R1215_U309 , P2_R1215_U310;
wire P2_R1215_U311 , P2_R1215_U312 , P2_R1215_U313 , P2_R1215_U314 , P2_R1215_U315 , P2_R1215_U316 , P2_R1215_U317 , P2_R1215_U318 , P2_R1215_U319 , P2_R1215_U320;
wire P2_R1215_U321 , P2_R1215_U322 , P2_R1215_U323 , P2_R1215_U324 , P2_R1215_U325 , P2_R1215_U326 , P2_R1215_U327 , P2_R1215_U328 , P2_R1215_U329 , P2_R1215_U330;
wire P2_R1215_U331 , P2_R1215_U332 , P2_R1215_U333 , P2_R1215_U334 , P2_R1215_U335 , P2_R1215_U336 , P2_R1215_U337 , P2_R1215_U338 , P2_R1215_U339 , P2_R1215_U340;
wire P2_R1215_U341 , P2_R1215_U342 , P2_R1215_U343 , P2_R1215_U344 , P2_R1215_U345 , P2_R1215_U346 , P2_R1215_U347 , P2_R1215_U348 , P2_R1215_U349 , P2_R1215_U350;
wire P2_R1215_U351 , P2_R1215_U352 , P2_R1215_U353 , P2_R1215_U354 , P2_R1215_U355 , P2_R1215_U356 , P2_R1215_U357 , P2_R1215_U358 , P2_R1215_U359 , P2_R1215_U360;
wire P2_R1215_U361 , P2_R1215_U362 , P2_R1215_U363 , P2_R1215_U364 , P2_R1215_U365 , P2_R1215_U366 , P2_R1215_U367 , P2_R1215_U368 , P2_R1215_U369 , P2_R1215_U370;
wire P2_R1215_U371 , P2_R1215_U372 , P2_R1215_U373 , P2_R1215_U374 , P2_R1215_U375 , P2_R1215_U376 , P2_R1215_U377 , P2_R1215_U378 , P2_R1215_U379 , P2_R1215_U380;
wire P2_R1215_U381 , P2_R1215_U382 , P2_R1215_U383 , P2_R1215_U384 , P2_R1215_U385 , P2_R1215_U386 , P2_R1215_U387 , P2_R1215_U388 , P2_R1215_U389 , P2_R1215_U390;
wire P2_R1215_U391 , P2_R1215_U392 , P2_R1215_U393 , P2_R1215_U394 , P2_R1215_U395 , P2_R1215_U396 , P2_R1215_U397 , P2_R1215_U398 , P2_R1215_U399 , P2_R1215_U400;
wire P2_R1215_U401 , P2_R1215_U402 , P2_R1215_U403 , P2_R1215_U404 , P2_R1215_U405 , P2_R1215_U406 , P2_R1215_U407 , P2_R1215_U408 , P2_R1215_U409 , P2_R1215_U410;
wire P2_R1215_U411 , P2_R1215_U412 , P2_R1215_U413 , P2_R1215_U414 , P2_R1215_U415 , P2_R1215_U416 , P2_R1215_U417 , P2_R1215_U418 , P2_R1215_U419 , P2_R1215_U420;
wire P2_R1215_U421 , P2_R1215_U422 , P2_R1215_U423 , P2_R1215_U424 , P2_R1215_U425 , P2_R1215_U426 , P2_R1215_U427 , P2_R1215_U428 , P2_R1215_U429 , P2_R1215_U430;
wire P2_R1215_U431 , P2_R1215_U432 , P2_R1215_U433 , P2_R1215_U434 , P2_R1215_U435 , P2_R1215_U436 , P2_R1215_U437 , P2_R1215_U438 , P2_R1215_U439 , P2_R1215_U440;
wire P2_R1215_U441 , P2_R1215_U442 , P2_R1215_U443 , P2_R1215_U444 , P2_R1215_U445 , P2_R1215_U446 , P2_R1215_U447 , P2_R1215_U448 , P2_R1215_U449 , P2_R1215_U450;
wire P2_R1215_U451 , P2_R1215_U452 , P2_R1215_U453 , P2_R1215_U454 , P2_R1215_U455 , P2_R1215_U456 , P2_R1215_U457 , P2_R1215_U458 , P2_R1215_U459 , P2_R1215_U460;
wire P2_R1215_U461 , P2_R1215_U462 , P2_R1215_U463 , P2_R1215_U464 , P2_R1215_U465 , P2_R1215_U466 , P2_R1215_U467 , P2_R1215_U468 , P2_R1215_U469 , P2_R1215_U470;
wire P2_R1215_U471 , P2_R1215_U472 , P2_R1215_U473 , P2_R1215_U474 , P2_R1215_U475 , P2_R1215_U476 , P2_R1215_U477 , P2_R1215_U478 , P2_R1215_U479 , P2_R1215_U480;
wire P2_R1215_U481 , P2_R1215_U482 , P2_R1215_U483 , P2_R1215_U484 , P2_R1215_U485 , P2_R1215_U486 , P2_R1215_U487 , P2_R1215_U488 , P2_R1215_U489 , P2_R1215_U490;
wire P2_R1215_U491 , P2_R1215_U492 , P2_R1215_U493 , P2_R1215_U494 , P2_R1215_U495 , P2_R1215_U496 , P2_R1215_U497 , P2_R1215_U498 , P2_R1215_U499 , P2_R1215_U500;
wire P2_R1215_U501 , P2_R1215_U502 , P2_R1215_U503 , P2_R1215_U504 , P2_R1164_U4 , P2_R1164_U5 , P2_R1164_U6 , P2_R1164_U7 , P2_R1164_U8 , P2_R1164_U9;
wire P2_R1164_U10 , P2_R1164_U11 , P2_R1164_U12 , P2_R1164_U13 , P2_R1164_U14 , P2_R1164_U15 , P2_R1164_U16 , P2_R1164_U17 , P2_R1164_U18 , P2_R1164_U19;
wire P2_R1164_U20 , P2_R1164_U21 , P2_R1164_U22 , P2_R1164_U23 , P2_R1164_U24 , P2_R1164_U25 , P2_R1164_U26 , P2_R1164_U27 , P2_R1164_U28 , P2_R1164_U29;
wire P2_R1164_U30 , P2_R1164_U31 , P2_R1164_U32 , P2_R1164_U33 , P2_R1164_U34 , P2_R1164_U35 , P2_R1164_U36 , P2_R1164_U37 , P2_R1164_U38 , P2_R1164_U39;
wire P2_R1164_U40 , P2_R1164_U41 , P2_R1164_U42 , P2_R1164_U43 , P2_R1164_U44 , P2_R1164_U45 , P2_R1164_U46 , P2_R1164_U47 , P2_R1164_U48 , P2_R1164_U49;
wire P2_R1164_U50 , P2_R1164_U51 , P2_R1164_U52 , P2_R1164_U53 , P2_R1164_U54 , P2_R1164_U55 , P2_R1164_U56 , P2_R1164_U57 , P2_R1164_U58 , P2_R1164_U59;
wire P2_R1164_U60 , P2_R1164_U61 , P2_R1164_U62 , P2_R1164_U63 , P2_R1164_U64 , P2_R1164_U65 , P2_R1164_U66 , P2_R1164_U67 , P2_R1164_U68 , P2_R1164_U69;
wire P2_R1164_U70 , P2_R1164_U71 , P2_R1164_U72 , P2_R1164_U73 , P2_R1164_U74 , P2_R1164_U75 , P2_R1164_U76 , P2_R1164_U77 , P2_R1164_U78 , P2_R1164_U79;
wire P2_R1164_U80 , P2_R1164_U81 , P2_R1164_U82 , P2_R1164_U83 , P2_R1164_U84 , P2_R1164_U85 , P2_R1164_U86 , P2_R1164_U87 , P2_R1164_U88 , P2_R1164_U89;
wire P2_R1164_U90 , P2_R1164_U91 , P2_R1164_U92 , P2_R1164_U93 , P2_R1164_U94 , P2_R1164_U95 , P2_R1164_U96 , P2_R1164_U97 , P2_R1164_U98 , P2_R1164_U99;
wire P2_R1164_U100 , P2_R1164_U101 , P2_R1164_U102 , P2_R1164_U103 , P2_R1164_U104 , P2_R1164_U105 , P2_R1164_U106 , P2_R1164_U107 , P2_R1164_U108 , P2_R1164_U109;
wire P2_R1164_U110 , P2_R1164_U111 , P2_R1164_U112 , P2_R1164_U113 , P2_R1164_U114 , P2_R1164_U115 , P2_R1164_U116 , P2_R1164_U117 , P2_R1164_U118 , P2_R1164_U119;
wire P2_R1164_U120 , P2_R1164_U121 , P2_R1164_U122 , P2_R1164_U123 , P2_R1164_U124 , P2_R1164_U125 , P2_R1164_U126 , P2_R1164_U127 , P2_R1164_U128 , P2_R1164_U129;
wire P2_R1164_U130 , P2_R1164_U131 , P2_R1164_U132 , P2_R1164_U133 , P2_R1164_U134 , P2_R1164_U135 , P2_R1164_U136 , P2_R1164_U137 , P2_R1164_U138 , P2_R1164_U139;
wire P2_R1164_U140 , P2_R1164_U141 , P2_R1164_U142 , P2_R1164_U143 , P2_R1164_U144 , P2_R1164_U145 , P2_R1164_U146 , P2_R1164_U147 , P2_R1164_U148 , P2_R1164_U149;
wire P2_R1164_U150 , P2_R1164_U151 , P2_R1164_U152 , P2_R1164_U153 , P2_R1164_U154 , P2_R1164_U155 , P2_R1164_U156 , P2_R1164_U157 , P2_R1164_U158 , P2_R1164_U159;
wire P2_R1164_U160 , P2_R1164_U161 , P2_R1164_U162 , P2_R1164_U163 , P2_R1164_U164 , P2_R1164_U165 , P2_R1164_U166 , P2_R1164_U167 , P2_R1164_U168 , P2_R1164_U169;
wire P2_R1164_U170 , P2_R1164_U171 , P2_R1164_U172 , P2_R1164_U173 , P2_R1164_U174 , P2_R1164_U175 , P2_R1164_U176 , P2_R1164_U177 , P2_R1164_U178 , P2_R1164_U179;
wire P2_R1164_U180 , P2_R1164_U181 , P2_R1164_U182 , P2_R1164_U183 , P2_R1164_U184 , P2_R1164_U185 , P2_R1164_U186 , P2_R1164_U187 , P2_R1164_U188 , P2_R1164_U189;
wire P2_R1164_U190 , P2_R1164_U191 , P2_R1164_U192 , P2_R1164_U193 , P2_R1164_U194 , P2_R1164_U195 , P2_R1164_U196 , P2_R1164_U197 , P2_R1164_U198 , P2_R1164_U199;
wire P2_R1164_U200 , P2_R1164_U201 , P2_R1164_U202 , P2_R1164_U203 , P2_R1164_U204 , P2_R1164_U205 , P2_R1164_U206 , P2_R1164_U207 , P2_R1164_U208 , P2_R1164_U209;
wire P2_R1164_U210 , P2_R1164_U211 , P2_R1164_U212 , P2_R1164_U213 , P2_R1164_U214 , P2_R1164_U215 , P2_R1164_U216 , P2_R1164_U217 , P2_R1164_U218 , P2_R1164_U219;
wire P2_R1164_U220 , P2_R1164_U221 , P2_R1164_U222 , P2_R1164_U223 , P2_R1164_U224 , P2_R1164_U225 , P2_R1164_U226 , P2_R1164_U227 , P2_R1164_U228 , P2_R1164_U229;
wire P2_R1164_U230 , P2_R1164_U231 , P2_R1164_U232 , P2_R1164_U233 , P2_R1164_U234 , P2_R1164_U235 , P2_R1164_U236 , P2_R1164_U237 , P2_R1164_U238 , P2_R1164_U239;
wire P2_R1164_U240 , P2_R1164_U241 , P2_R1164_U242 , P2_R1164_U243 , P2_R1164_U244 , P2_R1164_U245 , P2_R1164_U246 , P2_R1164_U247 , P2_R1164_U248 , P2_R1164_U249;
wire P2_R1164_U250 , P2_R1164_U251 , P2_R1164_U252 , P2_R1164_U253 , P2_R1164_U254 , P2_R1164_U255 , P2_R1164_U256 , P2_R1164_U257 , P2_R1164_U258 , P2_R1164_U259;
wire P2_R1164_U260 , P2_R1164_U261 , P2_R1164_U262 , P2_R1164_U263 , P2_R1164_U264 , P2_R1164_U265 , P2_R1164_U266 , P2_R1164_U267 , P2_R1164_U268 , P2_R1164_U269;
wire P2_R1164_U270 , P2_R1164_U271 , P2_R1164_U272 , P2_R1164_U273 , P2_R1164_U274 , P2_R1164_U275 , P2_R1164_U276 , P2_R1164_U277 , P2_R1164_U278 , P2_R1164_U279;
wire P2_R1164_U280 , P2_R1164_U281 , P2_R1164_U282 , P2_R1164_U283 , P2_R1164_U284 , P2_R1164_U285 , P2_R1164_U286 , P2_R1164_U287 , P2_R1164_U288 , P2_R1164_U289;
wire P2_R1164_U290 , P2_R1164_U291 , P2_R1164_U292 , P2_R1164_U293 , P2_R1164_U294 , P2_R1164_U295 , P2_R1164_U296 , P2_R1164_U297 , P2_R1164_U298 , P2_R1164_U299;
wire P2_R1164_U300 , P2_R1164_U301 , P2_R1164_U302 , P2_R1164_U303 , P2_R1164_U304 , P2_R1164_U305 , P2_R1164_U306 , P2_R1164_U307 , P2_R1164_U308 , P2_R1164_U309;
wire P2_R1164_U310 , P2_R1164_U311 , P2_R1164_U312 , P2_R1164_U313 , P2_R1164_U314 , P2_R1164_U315 , P2_R1164_U316 , P2_R1164_U317 , P2_R1164_U318 , P2_R1164_U319;
wire P2_R1164_U320 , P2_R1164_U321 , P2_R1164_U322 , P2_R1164_U323 , P2_R1164_U324 , P2_R1164_U325 , P2_R1164_U326 , P2_R1164_U327 , P2_R1164_U328 , P2_R1164_U329;
wire P2_R1164_U330 , P2_R1164_U331 , P2_R1164_U332 , P2_R1164_U333 , P2_R1164_U334 , P2_R1164_U335 , P2_R1164_U336 , P2_R1164_U337 , P2_R1164_U338 , P2_R1164_U339;
wire P2_R1164_U340 , P2_R1164_U341 , P2_R1164_U342 , P2_R1164_U343 , P2_R1164_U344 , P2_R1164_U345 , P2_R1164_U346 , P2_R1164_U347 , P2_R1164_U348 , P2_R1164_U349;
wire P2_R1164_U350 , P2_R1164_U351 , P2_R1164_U352 , P2_R1164_U353 , P2_R1164_U354 , P2_R1164_U355 , P2_R1164_U356 , P2_R1164_U357 , P2_R1164_U358 , P2_R1164_U359;
wire P2_R1164_U360 , P2_R1164_U361 , P2_R1164_U362 , P2_R1164_U363 , P2_R1164_U364 , P2_R1164_U365 , P2_R1164_U366 , P2_R1164_U367 , P2_R1164_U368 , P2_R1164_U369;
wire P2_R1164_U370 , P2_R1164_U371 , P2_R1164_U372 , P2_R1164_U373 , P2_R1164_U374 , P2_R1164_U375 , P2_R1164_U376 , P2_R1164_U377 , P2_R1164_U378 , P2_R1164_U379;
wire P2_R1164_U380 , P2_R1164_U381 , P2_R1164_U382 , P2_R1164_U383 , P2_R1164_U384 , P2_R1164_U385 , P2_R1164_U386 , P2_R1164_U387 , P2_R1164_U388 , P2_R1164_U389;
wire P2_R1164_U390 , P2_R1164_U391 , P2_R1164_U392 , P2_R1164_U393 , P2_R1164_U394 , P2_R1164_U395 , P2_R1164_U396 , P2_R1164_U397 , P2_R1164_U398 , P2_R1164_U399;
wire P2_R1164_U400 , P2_R1164_U401 , P2_R1164_U402 , P2_R1164_U403 , P2_R1164_U404 , P2_R1164_U405 , P2_R1164_U406 , P2_R1164_U407 , P2_R1164_U408 , P2_R1164_U409;
wire P2_R1164_U410 , P2_R1164_U411 , P2_R1164_U412 , P2_R1164_U413 , P2_R1164_U414 , P2_R1164_U415 , P2_R1164_U416 , P2_R1164_U417 , P2_R1164_U418 , P2_R1164_U419;
wire P2_R1164_U420 , P2_R1164_U421 , P2_R1164_U422 , P2_R1164_U423 , P2_R1164_U424 , P2_R1164_U425 , P2_R1164_U426 , P2_R1164_U427 , P2_R1164_U428 , P2_R1164_U429;
wire P2_R1164_U430 , P2_R1164_U431 , P2_R1164_U432 , P2_R1164_U433 , P2_R1164_U434 , P2_R1164_U435 , P2_R1164_U436 , P2_R1164_U437 , P2_R1164_U438 , P2_R1164_U439;
wire P2_R1164_U440 , P2_R1164_U441 , P2_R1164_U442 , P2_R1164_U443 , P2_R1164_U444 , P2_R1164_U445 , P2_R1164_U446 , P2_R1164_U447 , P2_R1164_U448 , P2_R1164_U449;
wire P2_R1164_U450 , P2_R1164_U451 , P2_R1164_U452 , P2_R1164_U453 , P2_R1164_U454 , P2_R1164_U455 , P2_R1164_U456 , P2_R1164_U457 , P2_R1164_U458 , P2_R1164_U459;
wire P2_R1164_U460 , P2_R1164_U461 , P2_R1164_U462 , P2_R1164_U463 , P2_R1164_U464 , P2_R1164_U465 , P2_R1164_U466 , P2_R1164_U467 , P2_R1164_U468 , P2_R1164_U469;
wire P2_R1164_U470 , P2_R1164_U471 , P2_R1164_U472 , P2_R1164_U473 , P2_R1164_U474 , P2_R1164_U475 , P2_R1164_U476 , P2_R1164_U477 , P2_R1164_U478 , P2_R1164_U479;
wire P2_R1164_U480 , P2_R1164_U481 , P2_R1164_U482 , P2_R1164_U483 , P2_R1164_U484 , P2_R1164_U485 , P2_R1164_U486 , P2_R1164_U487 , P2_R1164_U488 , P2_R1164_U489;
wire P2_R1164_U490 , P2_R1164_U491 , P2_R1164_U492 , P2_R1164_U493 , P2_R1164_U494 , P2_R1164_U495 , P2_R1164_U496 , P2_R1164_U497 , P2_R1164_U498 , P2_R1164_U499;
wire P2_R1164_U500 , P2_R1164_U501 , P2_R1164_U502 , P2_R1164_U503 , P2_R1164_U504 , P2_R1233_U4 , P2_R1233_U5 , P2_R1233_U6 , P2_R1233_U7 , P2_R1233_U8;
wire P2_R1233_U9 , P2_R1233_U10 , P2_R1233_U11 , P2_R1233_U12 , P2_R1233_U13 , P2_R1233_U14 , P2_R1233_U15 , P2_R1233_U16 , P2_R1233_U17 , P2_R1233_U18;
wire P2_R1233_U19 , P2_R1233_U20 , P2_R1233_U21 , P2_R1233_U22 , P2_R1233_U23 , P2_R1233_U24 , P2_R1233_U25 , P2_R1233_U26 , P2_R1233_U27 , P2_R1233_U28;
wire P2_R1233_U29 , P2_R1233_U30 , P2_R1233_U31 , P2_R1233_U32 , P2_R1233_U33 , P2_R1233_U34 , P2_R1233_U35 , P2_R1233_U36 , P2_R1233_U37 , P2_R1233_U38;
wire P2_R1233_U39 , P2_R1233_U40 , P2_R1233_U41 , P2_R1233_U42 , P2_R1233_U43 , P2_R1233_U44 , P2_R1233_U45 , P2_R1233_U46 , P2_R1233_U47 , P2_R1233_U48;
wire P2_R1233_U49 , P2_R1233_U50 , P2_R1233_U51 , P2_R1233_U52 , P2_R1233_U53 , P2_R1233_U54 , P2_R1233_U55 , P2_R1233_U56 , P2_R1233_U57 , P2_R1233_U58;
wire P2_R1233_U59 , P2_R1233_U60 , P2_R1233_U61 , P2_R1233_U62 , P2_R1233_U63 , P2_R1233_U64 , P2_R1233_U65 , P2_R1233_U66 , P2_R1233_U67 , P2_R1233_U68;
wire P2_R1233_U69 , P2_R1233_U70 , P2_R1233_U71 , P2_R1233_U72 , P2_R1233_U73 , P2_R1233_U74 , P2_R1233_U75 , P2_R1233_U76 , P2_R1233_U77 , P2_R1233_U78;
wire P2_R1233_U79 , P2_R1233_U80 , P2_R1233_U81 , P2_R1233_U82 , P2_R1233_U83 , P2_R1233_U84 , P2_R1233_U85 , P2_R1233_U86 , P2_R1233_U87 , P2_R1233_U88;
wire P2_R1233_U89 , P2_R1233_U90 , P2_R1233_U91 , P2_R1233_U92 , P2_R1233_U93 , P2_R1233_U94 , P2_R1233_U95 , P2_R1233_U96 , P2_R1233_U97 , P2_R1233_U98;
wire P2_R1233_U99 , P2_R1233_U100 , P2_R1233_U101 , P2_R1233_U102 , P2_R1233_U103 , P2_R1233_U104 , P2_R1233_U105 , P2_R1233_U106 , P2_R1233_U107 , P2_R1233_U108;
wire P2_R1233_U109 , P2_R1233_U110 , P2_R1233_U111 , P2_R1233_U112 , P2_R1233_U113 , P2_R1233_U114 , P2_R1233_U115 , P2_R1233_U116 , P2_R1233_U117 , P2_R1233_U118;
wire P2_R1233_U119 , P2_R1233_U120 , P2_R1233_U121 , P2_R1233_U122 , P2_R1233_U123 , P2_R1233_U124 , P2_R1233_U125 , P2_R1233_U126 , P2_R1233_U127 , P2_R1233_U128;
wire P2_R1233_U129 , P2_R1233_U130 , P2_R1233_U131 , P2_R1233_U132 , P2_R1233_U133 , P2_R1233_U134 , P2_R1233_U135 , P2_R1233_U136 , P2_R1233_U137 , P2_R1233_U138;
wire P2_R1233_U139 , P2_R1233_U140 , P2_R1233_U141 , P2_R1233_U142 , P2_R1233_U143 , P2_R1233_U144 , P2_R1233_U145 , P2_R1233_U146 , P2_R1233_U147 , P2_R1233_U148;
wire P2_R1233_U149 , P2_R1233_U150 , P2_R1233_U151 , P2_R1233_U152 , P2_R1233_U153 , P2_R1233_U154 , P2_R1233_U155 , P2_R1233_U156 , P2_R1233_U157 , P2_R1233_U158;
wire P2_R1233_U159 , P2_R1233_U160 , P2_R1233_U161 , P2_R1233_U162 , P2_R1233_U163 , P2_R1233_U164 , P2_R1233_U165 , P2_R1233_U166 , P2_R1233_U167 , P2_R1233_U168;
wire P2_R1233_U169 , P2_R1233_U170 , P2_R1233_U171 , P2_R1233_U172 , P2_R1233_U173 , P2_R1233_U174 , P2_R1233_U175 , P2_R1233_U176 , P2_R1233_U177 , P2_R1233_U178;
wire P2_R1233_U179 , P2_R1233_U180 , P2_R1233_U181 , P2_R1233_U182 , P2_R1233_U183 , P2_R1233_U184 , P2_R1233_U185 , P2_R1233_U186 , P2_R1233_U187 , P2_R1233_U188;
wire P2_R1233_U189 , P2_R1233_U190 , P2_R1233_U191 , P2_R1233_U192 , P2_R1233_U193 , P2_R1233_U194 , P2_R1233_U195 , P2_R1233_U196 , P2_R1233_U197 , P2_R1233_U198;
wire P2_R1233_U199 , P2_R1233_U200 , P2_R1233_U201 , P2_R1233_U202 , P2_R1233_U203 , P2_R1233_U204 , P2_R1233_U205 , P2_R1233_U206 , P2_R1233_U207 , P2_R1233_U208;
wire P2_R1233_U209 , P2_R1233_U210 , P2_R1233_U211 , P2_R1233_U212 , P2_R1233_U213 , P2_R1233_U214 , P2_R1233_U215 , P2_R1233_U216 , P2_R1233_U217 , P2_R1233_U218;
wire P2_R1233_U219 , P2_R1233_U220 , P2_R1233_U221 , P2_R1233_U222 , P2_R1233_U223 , P2_R1233_U224 , P2_R1233_U225 , P2_R1233_U226 , P2_R1233_U227 , P2_R1233_U228;
wire P2_R1233_U229 , P2_R1233_U230 , P2_R1233_U231 , P2_R1233_U232 , P2_R1233_U233 , P2_R1233_U234 , P2_R1233_U235 , P2_R1233_U236 , P2_R1233_U237 , P2_R1233_U238;
wire P2_R1233_U239 , P2_R1233_U240 , P2_R1233_U241 , P2_R1233_U242 , P2_R1233_U243 , P2_R1233_U244 , P2_R1233_U245 , P2_R1233_U246 , P2_R1233_U247 , P2_R1233_U248;
wire P2_R1233_U249 , P2_R1233_U250 , P2_R1233_U251 , P2_R1233_U252 , P2_R1233_U253 , P2_R1233_U254 , P2_R1233_U255 , P2_R1233_U256 , P2_R1233_U257 , P2_R1233_U258;
wire P2_R1233_U259 , P2_R1233_U260 , P2_R1233_U261 , P2_R1233_U262 , P2_R1233_U263 , P2_R1233_U264 , P2_R1233_U265 , P2_R1233_U266 , P2_R1233_U267 , P2_R1233_U268;
wire P2_R1233_U269 , P2_R1233_U270 , P2_R1233_U271 , P2_R1233_U272 , P2_R1233_U273 , P2_R1233_U274 , P2_R1233_U275 , P2_R1233_U276 , P2_R1233_U277 , P2_R1233_U278;
wire P2_R1233_U279 , P2_R1233_U280 , P2_R1233_U281 , P2_R1233_U282 , P2_R1233_U283 , P2_R1233_U284 , P2_R1233_U285 , P2_R1233_U286 , P2_R1233_U287 , P2_R1233_U288;
wire P2_R1233_U289 , P2_R1233_U290 , P2_R1233_U291 , P2_R1233_U292 , P2_R1233_U293 , P2_R1233_U294 , P2_R1233_U295 , P2_R1233_U296 , P2_R1233_U297 , P2_R1233_U298;
wire P2_R1233_U299 , P2_R1233_U300 , P2_R1233_U301 , P2_R1233_U302 , P2_R1233_U303 , P2_R1233_U304 , P2_R1233_U305 , P2_R1233_U306 , P2_R1233_U307 , P2_R1233_U308;
wire P2_R1233_U309 , P2_R1233_U310 , P2_R1233_U311 , P2_R1233_U312 , P2_R1233_U313 , P2_R1233_U314 , P2_R1233_U315 , P2_R1233_U316 , P2_R1233_U317 , P2_R1233_U318;
wire P2_R1233_U319 , P2_R1233_U320 , P2_R1233_U321 , P2_R1233_U322 , P2_R1233_U323 , P2_R1233_U324 , P2_R1233_U325 , P2_R1233_U326 , P2_R1233_U327 , P2_R1233_U328;
wire P2_R1233_U329 , P2_R1233_U330 , P2_R1233_U331 , P2_R1233_U332 , P2_R1233_U333 , P2_R1233_U334 , P2_R1233_U335 , P2_R1233_U336 , P2_R1233_U337 , P2_R1233_U338;
wire P2_R1233_U339 , P2_R1233_U340 , P2_R1233_U341 , P2_R1233_U342 , P2_R1233_U343 , P2_R1233_U344 , P2_R1233_U345 , P2_R1233_U346 , P2_R1233_U347 , P2_R1233_U348;
wire P2_R1233_U349 , P2_R1233_U350 , P2_R1233_U351 , P2_R1233_U352 , P2_R1233_U353 , P2_R1233_U354 , P2_R1233_U355 , P2_R1233_U356 , P2_R1233_U357 , P2_R1233_U358;
wire P2_R1233_U359 , P2_R1233_U360 , P2_R1233_U361 , P2_R1233_U362 , P2_R1233_U363 , P2_R1233_U364 , P2_R1233_U365 , P2_R1233_U366 , P2_R1233_U367 , P2_R1233_U368;
wire P2_R1233_U369 , P2_R1233_U370 , P2_R1233_U371 , P2_R1233_U372 , P2_R1233_U373 , P2_R1233_U374 , P2_R1233_U375 , P2_R1233_U376 , P2_R1233_U377 , P2_R1233_U378;
wire P2_R1233_U379 , P2_R1233_U380 , P2_R1233_U381 , P2_R1233_U382 , P2_R1233_U383 , P2_R1233_U384 , P2_R1233_U385 , P2_R1233_U386 , P2_R1233_U387 , P2_R1233_U388;
wire P2_R1233_U389 , P2_R1233_U390 , P2_R1233_U391 , P2_R1233_U392 , P2_R1233_U393 , P2_R1233_U394 , P2_R1233_U395 , P2_R1233_U396 , P2_R1233_U397 , P2_R1233_U398;
wire P2_R1233_U399 , P2_R1233_U400 , P2_R1233_U401 , P2_R1233_U402 , P2_R1233_U403 , P2_R1233_U404 , P2_R1233_U405 , P2_R1233_U406 , P2_R1233_U407 , P2_R1233_U408;
wire P2_R1233_U409 , P2_R1233_U410 , P2_R1233_U411 , P2_R1233_U412 , P2_R1233_U413 , P2_R1233_U414 , P2_R1233_U415 , P2_R1233_U416 , P2_R1233_U417 , P2_R1233_U418;
wire P2_R1233_U419 , P2_R1233_U420 , P2_R1233_U421 , P2_R1233_U422 , P2_R1233_U423 , P2_R1233_U424 , P2_R1233_U425 , P2_R1233_U426 , P2_R1233_U427 , P2_R1233_U428;
wire P2_R1233_U429 , P2_R1233_U430 , P2_R1233_U431 , P2_R1233_U432 , P2_R1233_U433 , P2_R1233_U434 , P2_R1233_U435 , P2_R1233_U436 , P2_R1233_U437 , P2_R1233_U438;
wire P2_R1233_U439 , P2_R1233_U440 , P2_R1233_U441 , P2_R1233_U442 , P2_R1233_U443 , P2_R1233_U444 , P2_R1233_U445 , P2_R1233_U446 , P2_R1233_U447 , P2_R1233_U448;
wire P2_R1233_U449 , P2_R1233_U450 , P2_R1233_U451 , P2_R1233_U452 , P2_R1233_U453 , P2_R1233_U454 , P2_R1233_U455 , P2_R1233_U456 , P2_R1233_U457 , P2_R1233_U458;
wire P2_R1233_U459 , P2_R1233_U460 , P2_R1233_U461 , P2_R1233_U462 , P2_R1233_U463 , P2_R1233_U464 , P2_R1233_U465 , P2_R1233_U466 , P2_R1233_U467 , P2_R1233_U468;
wire P2_R1233_U469 , P2_R1233_U470 , P2_R1233_U471 , P2_R1233_U472 , P2_R1233_U473 , P2_R1233_U474 , P2_R1233_U475 , P2_R1233_U476 , P2_R1233_U477 , P2_R1233_U478;
wire P2_R1233_U479 , P2_R1233_U480 , P2_R1233_U481 , P2_R1233_U482 , P2_R1233_U483 , P2_R1233_U484 , P2_R1233_U485 , P2_R1233_U486 , P2_R1233_U487 , P2_R1233_U488;
wire P2_R1233_U489 , P2_R1233_U490 , P2_R1233_U491 , P2_R1233_U492 , P2_R1233_U493 , P2_R1233_U494 , P2_R1233_U495 , P2_R1233_U496 , P2_R1233_U497 , P2_R1233_U498;
wire P2_R1233_U499 , P2_R1233_U500 , P2_R1233_U501 , P2_R1233_U502 , P2_R1233_U503 , P2_R1233_U504 , P2_R1176_U4 , P2_R1176_U5 , P2_R1176_U6 , P2_R1176_U7;
wire P2_R1176_U8 , P2_R1176_U9 , P2_R1176_U10 , P2_R1176_U11 , P2_R1176_U12 , P2_R1176_U13 , P2_R1176_U14 , P2_R1176_U15 , P2_R1176_U16 , P2_R1176_U17;
wire P2_R1176_U18 , P2_R1176_U19 , P2_R1176_U20 , P2_R1176_U21 , P2_R1176_U22 , P2_R1176_U23 , P2_R1176_U24 , P2_R1176_U25 , P2_R1176_U26 , P2_R1176_U27;
wire P2_R1176_U28 , P2_R1176_U29 , P2_R1176_U30 , P2_R1176_U31 , P2_R1176_U32 , P2_R1176_U33 , P2_R1176_U34 , P2_R1176_U35 , P2_R1176_U36 , P2_R1176_U37;
wire P2_R1176_U38 , P2_R1176_U39 , P2_R1176_U40 , P2_R1176_U41 , P2_R1176_U42 , P2_R1176_U43 , P2_R1176_U44 , P2_R1176_U45 , P2_R1176_U46 , P2_R1176_U47;
wire P2_R1176_U48 , P2_R1176_U49 , P2_R1176_U50 , P2_R1176_U51 , P2_R1176_U52 , P2_R1176_U53 , P2_R1176_U54 , P2_R1176_U55 , P2_R1176_U56 , P2_R1176_U57;
wire P2_R1176_U58 , P2_R1176_U59 , P2_R1176_U60 , P2_R1176_U61 , P2_R1176_U62 , P2_R1176_U63 , P2_R1176_U64 , P2_R1176_U65 , P2_R1176_U66 , P2_R1176_U67;
wire P2_R1176_U68 , P2_R1176_U69 , P2_R1176_U70 , P2_R1176_U71 , P2_R1176_U72 , P2_R1176_U73 , P2_R1176_U74 , P2_R1176_U75 , P2_R1176_U76 , P2_R1176_U77;
wire P2_R1176_U78 , P2_R1176_U79 , P2_R1176_U80 , P2_R1176_U81 , P2_R1176_U82 , P2_R1176_U83 , P2_R1176_U84 , P2_R1176_U85 , P2_R1176_U86 , P2_R1176_U87;
wire P2_R1176_U88 , P2_R1176_U89 , P2_R1176_U90 , P2_R1176_U91 , P2_R1176_U92 , P2_R1176_U93 , P2_R1176_U94 , P2_R1176_U95 , P2_R1176_U96 , P2_R1176_U97;
wire P2_R1176_U98 , P2_R1176_U99 , P2_R1176_U100 , P2_R1176_U101 , P2_R1176_U102 , P2_R1176_U103 , P2_R1176_U104 , P2_R1176_U105 , P2_R1176_U106 , P2_R1176_U107;
wire P2_R1176_U108 , P2_R1176_U109 , P2_R1176_U110 , P2_R1176_U111 , P2_R1176_U112 , P2_R1176_U113 , P2_R1176_U114 , P2_R1176_U115 , P2_R1176_U116 , P2_R1176_U117;
wire P2_R1176_U118 , P2_R1176_U119 , P2_R1176_U120 , P2_R1176_U121 , P2_R1176_U122 , P2_R1176_U123 , P2_R1176_U124 , P2_R1176_U125 , P2_R1176_U126 , P2_R1176_U127;
wire P2_R1176_U128 , P2_R1176_U129 , P2_R1176_U130 , P2_R1176_U131 , P2_R1176_U132 , P2_R1176_U133 , P2_R1176_U134 , P2_R1176_U135 , P2_R1176_U136 , P2_R1176_U137;
wire P2_R1176_U138 , P2_R1176_U139 , P2_R1176_U140 , P2_R1176_U141 , P2_R1176_U142 , P2_R1176_U143 , P2_R1176_U144 , P2_R1176_U145 , P2_R1176_U146 , P2_R1176_U147;
wire P2_R1176_U148 , P2_R1176_U149 , P2_R1176_U150 , P2_R1176_U151 , P2_R1176_U152 , P2_R1176_U153 , P2_R1176_U154 , P2_R1176_U155 , P2_R1176_U156 , P2_R1176_U157;
wire P2_R1176_U158 , P2_R1176_U159 , P2_R1176_U160 , P2_R1176_U161 , P2_R1176_U162 , P2_R1176_U163 , P2_R1176_U164 , P2_R1176_U165 , P2_R1176_U166 , P2_R1176_U167;
wire P2_R1176_U168 , P2_R1176_U169 , P2_R1176_U170 , P2_R1176_U171 , P2_R1176_U172 , P2_R1176_U173 , P2_R1176_U174 , P2_R1176_U175 , P2_R1176_U176 , P2_R1176_U177;
wire P2_R1176_U178 , P2_R1176_U179 , P2_R1176_U180 , P2_R1176_U181 , P2_R1176_U182 , P2_R1176_U183 , P2_R1176_U184 , P2_R1176_U185 , P2_R1176_U186 , P2_R1176_U187;
wire P2_R1176_U188 , P2_R1176_U189 , P2_R1176_U190 , P2_R1176_U191 , P2_R1176_U192 , P2_R1176_U193 , P2_R1176_U194 , P2_R1176_U195 , P2_R1176_U196 , P2_R1176_U197;
wire P2_R1176_U198 , P2_R1176_U199 , P2_R1176_U200 , P2_R1176_U201 , P2_R1176_U202 , P2_R1176_U203 , P2_R1176_U204 , P2_R1176_U205 , P2_R1176_U206 , P2_R1176_U207;
wire P2_R1176_U208 , P2_R1176_U209 , P2_R1176_U210 , P2_R1176_U211 , P2_R1176_U212 , P2_R1176_U213 , P2_R1176_U214 , P2_R1176_U215 , P2_R1176_U216 , P2_R1176_U217;
wire P2_R1176_U218 , P2_R1176_U219 , P2_R1176_U220 , P2_R1176_U221 , P2_R1176_U222 , P2_R1176_U223 , P2_R1176_U224 , P2_R1176_U225 , P2_R1176_U226 , P2_R1176_U227;
wire P2_R1176_U228 , P2_R1176_U229 , P2_R1176_U230 , P2_R1176_U231 , P2_R1176_U232 , P2_R1176_U233 , P2_R1176_U234 , P2_R1176_U235 , P2_R1176_U236 , P2_R1176_U237;
wire P2_R1176_U238 , P2_R1176_U239 , P2_R1176_U240 , P2_R1176_U241 , P2_R1176_U242 , P2_R1176_U243 , P2_R1176_U244 , P2_R1176_U245 , P2_R1176_U246 , P2_R1176_U247;
wire P2_R1176_U248 , P2_R1176_U249 , P2_R1176_U250 , P2_R1176_U251 , P2_R1176_U252 , P2_R1176_U253 , P2_R1176_U254 , P2_R1176_U255 , P2_R1176_U256 , P2_R1176_U257;
wire P2_R1176_U258 , P2_R1176_U259 , P2_R1176_U260 , P2_R1176_U261 , P2_R1176_U262 , P2_R1176_U263 , P2_R1176_U264 , P2_R1176_U265 , P2_R1176_U266 , P2_R1176_U267;
wire P2_R1176_U268 , P2_R1176_U269 , P2_R1176_U270 , P2_R1176_U271 , P2_R1176_U272 , P2_R1176_U273 , P2_R1176_U274 , P2_R1176_U275 , P2_R1176_U276 , P2_R1176_U277;
wire P2_R1176_U278 , P2_R1176_U279 , P2_R1176_U280 , P2_R1176_U281 , P2_R1176_U282 , P2_R1176_U283 , P2_R1176_U284 , P2_R1176_U285 , P2_R1176_U286 , P2_R1176_U287;
wire P2_R1176_U288 , P2_R1176_U289 , P2_R1176_U290 , P2_R1176_U291 , P2_R1176_U292 , P2_R1176_U293 , P2_R1176_U294 , P2_R1176_U295 , P2_R1176_U296 , P2_R1176_U297;
wire P2_R1176_U298 , P2_R1176_U299 , P2_R1176_U300 , P2_R1176_U301 , P2_R1176_U302 , P2_R1176_U303 , P2_R1176_U304 , P2_R1176_U305 , P2_R1176_U306 , P2_R1176_U307;
wire P2_R1176_U308 , P2_R1176_U309 , P2_R1176_U310 , P2_R1176_U311 , P2_R1176_U312 , P2_R1176_U313 , P2_R1176_U314 , P2_R1176_U315 , P2_R1176_U316 , P2_R1176_U317;
wire P2_R1176_U318 , P2_R1176_U319 , P2_R1176_U320 , P2_R1176_U321 , P2_R1176_U322 , P2_R1176_U323 , P2_R1176_U324 , P2_R1176_U325 , P2_R1176_U326 , P2_R1176_U327;
wire P2_R1176_U328 , P2_R1176_U329 , P2_R1176_U330 , P2_R1176_U331 , P2_R1176_U332 , P2_R1176_U333 , P2_R1176_U334 , P2_R1176_U335 , P2_R1176_U336 , P2_R1176_U337;
wire P2_R1176_U338 , P2_R1176_U339 , P2_R1176_U340 , P2_R1176_U341 , P2_R1176_U342 , P2_R1176_U343 , P2_R1176_U344 , P2_R1176_U345 , P2_R1176_U346 , P2_R1176_U347;
wire P2_R1176_U348 , P2_R1176_U349 , P2_R1176_U350 , P2_R1176_U351 , P2_R1176_U352 , P2_R1176_U353 , P2_R1176_U354 , P2_R1176_U355 , P2_R1176_U356 , P2_R1176_U357;
wire P2_R1176_U358 , P2_R1176_U359 , P2_R1176_U360 , P2_R1176_U361 , P2_R1176_U362 , P2_R1176_U363 , P2_R1176_U364 , P2_R1176_U365 , P2_R1176_U366 , P2_R1176_U367;
wire P2_R1176_U368 , P2_R1176_U369 , P2_R1176_U370 , P2_R1176_U371 , P2_R1176_U372 , P2_R1176_U373 , P2_R1176_U374 , P2_R1176_U375 , P2_R1176_U376 , P2_R1176_U377;
wire P2_R1176_U378 , P2_R1176_U379 , P2_R1176_U380 , P2_R1176_U381 , P2_R1176_U382 , P2_R1176_U383 , P2_R1176_U384 , P2_R1176_U385 , P2_R1176_U386 , P2_R1176_U387;
wire P2_R1176_U388 , P2_R1176_U389 , P2_R1176_U390 , P2_R1176_U391 , P2_R1176_U392 , P2_R1176_U393 , P2_R1176_U394 , P2_R1176_U395 , P2_R1176_U396 , P2_R1176_U397;
wire P2_R1176_U398 , P2_R1176_U399 , P2_R1176_U400 , P2_R1176_U401 , P2_R1176_U402 , P2_R1176_U403 , P2_R1176_U404 , P2_R1176_U405 , P2_R1176_U406 , P2_R1176_U407;
wire P2_R1176_U408 , P2_R1176_U409 , P2_R1176_U410 , P2_R1176_U411 , P2_R1176_U412 , P2_R1176_U413 , P2_R1176_U414 , P2_R1176_U415 , P2_R1176_U416 , P2_R1176_U417;
wire P2_R1176_U418 , P2_R1176_U419 , P2_R1176_U420 , P2_R1176_U421 , P2_R1176_U422 , P2_R1176_U423 , P2_R1176_U424 , P2_R1176_U425 , P2_R1176_U426 , P2_R1176_U427;
wire P2_R1176_U428 , P2_R1176_U429 , P2_R1176_U430 , P2_R1176_U431 , P2_R1176_U432 , P2_R1176_U433 , P2_R1176_U434 , P2_R1176_U435 , P2_R1176_U436 , P2_R1176_U437;
wire P2_R1176_U438 , P2_R1176_U439 , P2_R1176_U440 , P2_R1176_U441 , P2_R1176_U442 , P2_R1176_U443 , P2_R1176_U444 , P2_R1176_U445 , P2_R1176_U446 , P2_R1176_U447;
wire P2_R1176_U448 , P2_R1176_U449 , P2_R1176_U450 , P2_R1176_U451 , P2_R1176_U452 , P2_R1176_U453 , P2_R1176_U454 , P2_R1176_U455 , P2_R1176_U456 , P2_R1176_U457;
wire P2_R1176_U458 , P2_R1176_U459 , P2_R1176_U460 , P2_R1176_U461 , P2_R1176_U462 , P2_R1176_U463 , P2_R1176_U464 , P2_R1176_U465 , P2_R1176_U466 , P2_R1176_U467;
wire P2_R1176_U468 , P2_R1176_U469 , P2_R1176_U470 , P2_R1176_U471 , P2_R1176_U472 , P2_R1176_U473 , P2_R1176_U474 , P2_R1176_U475 , P2_R1176_U476 , P2_R1176_U477;
wire P2_R1176_U478 , P2_R1176_U479 , P2_R1176_U480 , P2_R1176_U481 , P2_R1176_U482 , P2_R1176_U483 , P2_R1176_U484 , P2_R1176_U485 , P2_R1176_U486 , P2_R1176_U487;
wire P2_R1176_U488 , P2_R1176_U489 , P2_R1176_U490 , P2_R1176_U491 , P2_R1176_U492 , P2_R1176_U493 , P2_R1176_U494 , P2_R1176_U495 , P2_R1176_U496 , P2_R1176_U497;
wire P2_R1176_U498 , P2_R1176_U499 , P2_R1176_U500 , P2_R1176_U501 , P2_R1176_U502 , P2_R1176_U503 , P2_R1176_U504 , P2_R1176_U505 , P2_R1176_U506 , P2_R1176_U507;
wire P2_R1176_U508 , P2_R1176_U509 , P2_R1176_U510 , P2_R1176_U511 , P2_R1176_U512 , P2_R1176_U513 , P2_R1176_U514 , P2_R1176_U515 , P2_R1176_U516 , P2_R1176_U517;
wire P2_R1176_U518 , P2_R1176_U519 , P2_R1176_U520 , P2_R1176_U521 , P2_R1176_U522 , P2_R1176_U523 , P2_R1176_U524 , P2_R1176_U525 , P2_R1176_U526 , P2_R1176_U527;
wire P2_R1176_U528 , P2_R1176_U529 , P2_R1176_U530 , P2_R1176_U531 , P2_R1176_U532 , P2_R1176_U533 , P2_R1176_U534 , P2_R1176_U535 , P2_R1176_U536 , P2_R1176_U537;
wire P2_R1176_U538 , P2_R1176_U539 , P2_R1176_U540 , P2_R1176_U541 , P2_R1176_U542 , P2_R1176_U543 , P2_R1176_U544 , P2_R1176_U545 , P2_R1176_U546 , P2_R1176_U547;
wire P2_R1176_U548 , P2_R1176_U549 , P2_R1176_U550 , P2_R1176_U551 , P2_R1176_U552 , P2_R1176_U553 , P2_R1176_U554 , P2_R1176_U555 , P2_R1176_U556 , P2_R1176_U557;
wire P2_R1176_U558 , P2_R1176_U559 , P2_R1176_U560 , P2_R1176_U561 , P2_R1176_U562 , P2_R1176_U563 , P2_R1176_U564 , P2_R1176_U565 , P2_R1176_U566 , P2_R1176_U567;
wire P2_R1176_U568 , P2_R1176_U569 , P2_R1176_U570 , P2_R1176_U571 , P2_R1176_U572 , P2_R1176_U573 , P2_R1176_U574 , P2_R1176_U575 , P2_R1176_U576 , P2_R1176_U577;
wire P2_R1176_U578 , P2_R1176_U579 , P2_R1176_U580 , P2_R1176_U581 , P2_R1176_U582 , P2_R1176_U583 , P2_R1176_U584 , P2_R1176_U585 , P2_R1176_U586 , P2_R1176_U587;
wire P2_R1176_U588 , P2_R1176_U589 , P2_R1176_U590 , P2_R1176_U591 , P2_R1176_U592 , P2_R1176_U593 , P2_R1176_U594 , P2_R1176_U595 , P2_R1176_U596 , P2_R1176_U597;
wire P2_R1176_U598 , P2_R1176_U599 , P2_R1176_U600 , P2_R1176_U601 , P2_R1176_U602 , P2_R1176_U603 , P2_R1176_U604 , P2_R1176_U605 , P2_R1176_U606 , P2_R1176_U607;
wire P2_R1176_U608 , P2_R1176_U609 , P2_R1176_U610 , P2_R1176_U611 , P2_R1176_U612 , P2_R1176_U613 , P2_R1176_U614 , P2_R1176_U615 , P2_R1176_U616 , P2_R1176_U617;
wire P2_R1176_U618 , P2_R1176_U619 , P2_R1176_U620 , P2_R1176_U621 , P2_R1176_U622 , P2_R1176_U623 , P2_R1131_U4 , P2_R1131_U5 , P2_R1131_U6 , P2_R1131_U7;
wire P2_R1131_U8 , P2_R1131_U9 , P2_R1131_U10 , P2_R1131_U11 , P2_R1131_U12 , P2_R1131_U13 , P2_R1131_U14 , P2_R1131_U15 , P2_R1131_U16 , P2_R1131_U17;
wire P2_R1131_U18 , P2_R1131_U19 , P2_R1131_U20 , P2_R1131_U21 , P2_R1131_U22 , P2_R1131_U23 , P2_R1131_U24 , P2_R1131_U25 , P2_R1131_U26 , P2_R1131_U27;
wire P2_R1131_U28 , P2_R1131_U29 , P2_R1131_U30 , P2_R1131_U31 , P2_R1131_U32 , P2_R1131_U33 , P2_R1131_U34 , P2_R1131_U35 , P2_R1131_U36 , P2_R1131_U37;
wire P2_R1131_U38 , P2_R1131_U39 , P2_R1131_U40 , P2_R1131_U41 , P2_R1131_U42 , P2_R1131_U43 , P2_R1131_U44 , P2_R1131_U45 , P2_R1131_U46 , P2_R1131_U47;
wire P2_R1131_U48 , P2_R1131_U49 , P2_R1131_U50 , P2_R1131_U51 , P2_R1131_U52 , P2_R1131_U53 , P2_R1131_U54 , P2_R1131_U55 , P2_R1131_U56 , P2_R1131_U57;
wire P2_R1131_U58 , P2_R1131_U59 , P2_R1131_U60 , P2_R1131_U61 , P2_R1131_U62 , P2_R1131_U63 , P2_R1131_U64 , P2_R1131_U65 , P2_R1131_U66 , P2_R1131_U67;
wire P2_R1131_U68 , P2_R1131_U69 , P2_R1131_U70 , P2_R1131_U71 , P2_R1131_U72 , P2_R1131_U73 , P2_R1131_U74 , P2_R1131_U75 , P2_R1131_U76 , P2_R1131_U77;
wire P2_R1131_U78 , P2_R1131_U79 , P2_R1131_U80 , P2_R1131_U81 , P2_R1131_U82 , P2_R1131_U83 , P2_R1131_U84 , P2_R1131_U85 , P2_R1131_U86 , P2_R1131_U87;
wire P2_R1131_U88 , P2_R1131_U89 , P2_R1131_U90 , P2_R1131_U91 , P2_R1131_U92 , P2_R1131_U93 , P2_R1131_U94 , P2_R1131_U95 , P2_R1131_U96 , P2_R1131_U97;
wire P2_R1131_U98 , P2_R1131_U99 , P2_R1131_U100 , P2_R1131_U101 , P2_R1131_U102 , P2_R1131_U103 , P2_R1131_U104 , P2_R1131_U105 , P2_R1131_U106 , P2_R1131_U107;
wire P2_R1131_U108 , P2_R1131_U109 , P2_R1131_U110 , P2_R1131_U111 , P2_R1131_U112 , P2_R1131_U113 , P2_R1131_U114 , P2_R1131_U115 , P2_R1131_U116 , P2_R1131_U117;
wire P2_R1131_U118 , P2_R1131_U119 , P2_R1131_U120 , P2_R1131_U121 , P2_R1131_U122 , P2_R1131_U123 , P2_R1131_U124 , P2_R1131_U125 , P2_R1131_U126 , P2_R1131_U127;
wire P2_R1131_U128 , P2_R1131_U129 , P2_R1131_U130 , P2_R1131_U131 , P2_R1131_U132 , P2_R1131_U133 , P2_R1131_U134 , P2_R1131_U135 , P2_R1131_U136 , P2_R1131_U137;
wire P2_R1131_U138 , P2_R1131_U139 , P2_R1131_U140 , P2_R1131_U141 , P2_R1131_U142 , P2_R1131_U143 , P2_R1131_U144 , P2_R1131_U145 , P2_R1131_U146 , P2_R1131_U147;
wire P2_R1131_U148 , P2_R1131_U149 , P2_R1131_U150 , P2_R1131_U151 , P2_R1131_U152 , P2_R1131_U153 , P2_R1131_U154 , P2_R1131_U155 , P2_R1131_U156 , P2_R1131_U157;
wire P2_R1131_U158 , P2_R1131_U159 , P2_R1131_U160 , P2_R1131_U161 , P2_R1131_U162 , P2_R1131_U163 , P2_R1131_U164 , P2_R1131_U165 , P2_R1131_U166 , P2_R1131_U167;
wire P2_R1131_U168 , P2_R1131_U169 , P2_R1131_U170 , P2_R1131_U171 , P2_R1131_U172 , P2_R1131_U173 , P2_R1131_U174 , P2_R1131_U175 , P2_R1131_U176 , P2_R1131_U177;
wire P2_R1131_U178 , P2_R1131_U179 , P2_R1131_U180 , P2_R1131_U181 , P2_R1131_U182 , P2_R1131_U183 , P2_R1131_U184 , P2_R1131_U185 , P2_R1131_U186 , P2_R1131_U187;
wire P2_R1131_U188 , P2_R1131_U189 , P2_R1131_U190 , P2_R1131_U191 , P2_R1131_U192 , P2_R1131_U193 , P2_R1131_U194 , P2_R1131_U195 , P2_R1131_U196 , P2_R1131_U197;
wire P2_R1131_U198 , P2_R1131_U199 , P2_R1131_U200 , P2_R1131_U201 , P2_R1131_U202 , P2_R1131_U203 , P2_R1131_U204 , P2_R1131_U205 , P2_R1131_U206 , P2_R1131_U207;
wire P2_R1131_U208 , P2_R1131_U209 , P2_R1131_U210 , P2_R1131_U211 , P2_R1131_U212 , P2_R1131_U213 , P2_R1131_U214 , P2_R1131_U215 , P2_R1131_U216 , P2_R1131_U217;
wire P2_R1131_U218 , P2_R1131_U219 , P2_R1131_U220 , P2_R1131_U221 , P2_R1131_U222 , P2_R1131_U223 , P2_R1131_U224 , P2_R1131_U225 , P2_R1131_U226 , P2_R1131_U227;
wire P2_R1131_U228 , P2_R1131_U229 , P2_R1131_U230 , P2_R1131_U231 , P2_R1131_U232 , P2_R1131_U233 , P2_R1131_U234 , P2_R1131_U235 , P2_R1131_U236 , P2_R1131_U237;
wire P2_R1131_U238 , P2_R1131_U239 , P2_R1131_U240 , P2_R1131_U241 , P2_R1131_U242 , P2_R1131_U243 , P2_R1131_U244 , P2_R1131_U245 , P2_R1131_U246 , P2_R1131_U247;
wire P2_R1131_U248 , P2_R1131_U249 , P2_R1131_U250 , P2_R1131_U251 , P2_R1131_U252 , P2_R1131_U253 , P2_R1131_U254 , P2_R1131_U255 , P2_R1131_U256 , P2_R1131_U257;
wire P2_R1131_U258 , P2_R1131_U259 , P2_R1131_U260 , P2_R1131_U261 , P2_R1131_U262 , P2_R1131_U263 , P2_R1131_U264 , P2_R1131_U265 , P2_R1131_U266 , P2_R1131_U267;
wire P2_R1131_U268 , P2_R1131_U269 , P2_R1131_U270 , P2_R1131_U271 , P2_R1131_U272 , P2_R1131_U273 , P2_R1131_U274 , P2_R1131_U275 , P2_R1131_U276 , P2_R1131_U277;
wire P2_R1131_U278 , P2_R1131_U279 , P2_R1131_U280 , P2_R1131_U281 , P2_R1131_U282 , P2_R1131_U283 , P2_R1131_U284 , P2_R1131_U285 , P2_R1131_U286 , P2_R1131_U287;
wire P2_R1131_U288 , P2_R1131_U289 , P2_R1131_U290 , P2_R1131_U291 , P2_R1131_U292 , P2_R1131_U293 , P2_R1131_U294 , P2_R1131_U295 , P2_R1131_U296 , P2_R1131_U297;
wire P2_R1131_U298 , P2_R1131_U299 , P2_R1131_U300 , P2_R1131_U301 , P2_R1131_U302 , P2_R1131_U303 , P2_R1131_U304 , P2_R1131_U305 , P2_R1131_U306 , P2_R1131_U307;
wire P2_R1131_U308 , P2_R1131_U309 , P2_R1131_U310 , P2_R1131_U311 , P2_R1131_U312 , P2_R1131_U313 , P2_R1131_U314 , P2_R1131_U315 , P2_R1131_U316 , P2_R1131_U317;
wire P2_R1131_U318 , P2_R1131_U319 , P2_R1131_U320 , P2_R1131_U321 , P2_R1131_U322 , P2_R1131_U323 , P2_R1131_U324 , P2_R1131_U325 , P2_R1131_U326 , P2_R1131_U327;
wire P2_R1131_U328 , P2_R1131_U329 , P2_R1131_U330 , P2_R1131_U331 , P2_R1131_U332 , P2_R1131_U333 , P2_R1131_U334 , P2_R1131_U335 , P2_R1131_U336 , P2_R1131_U337;
wire P2_R1131_U338 , P2_R1131_U339 , P2_R1131_U340 , P2_R1131_U341 , P2_R1131_U342 , P2_R1131_U343 , P2_R1131_U344 , P2_R1131_U345 , P2_R1131_U346 , P2_R1131_U347;
wire P2_R1131_U348 , P2_R1131_U349 , P2_R1131_U350 , P2_R1131_U351 , P2_R1131_U352 , P2_R1131_U353 , P2_R1131_U354 , P2_R1131_U355 , P2_R1131_U356 , P2_R1131_U357;
wire P2_R1131_U358 , P2_R1131_U359 , P2_R1131_U360 , P2_R1131_U361 , P2_R1131_U362 , P2_R1131_U363 , P2_R1131_U364 , P2_R1131_U365 , P2_R1131_U366 , P2_R1131_U367;
wire P2_R1131_U368 , P2_R1131_U369 , P2_R1131_U370 , P2_R1131_U371 , P2_R1131_U372 , P2_R1131_U373 , P2_R1131_U374 , P2_R1131_U375 , P2_R1131_U376 , P2_R1131_U377;
wire P2_R1131_U378 , P2_R1131_U379 , P2_R1131_U380 , P2_R1131_U381 , P2_R1131_U382 , P2_R1131_U383 , P2_R1131_U384 , P2_R1131_U385 , P2_R1131_U386 , P2_R1131_U387;
wire P2_R1131_U388 , P2_R1131_U389 , P2_R1131_U390 , P2_R1131_U391 , P2_R1131_U392 , P2_R1131_U393 , P2_R1131_U394 , P2_R1131_U395 , P2_R1131_U396 , P2_R1131_U397;
wire P2_R1131_U398 , P2_R1131_U399 , P2_R1131_U400 , P2_R1131_U401 , P2_R1131_U402 , P2_R1131_U403 , P2_R1131_U404 , P2_R1131_U405 , P2_R1131_U406 , P2_R1131_U407;
wire P2_R1131_U408 , P2_R1131_U409 , P2_R1131_U410 , P2_R1131_U411 , P2_R1131_U412 , P2_R1131_U413 , P2_R1131_U414 , P2_R1131_U415 , P2_R1131_U416 , P2_R1131_U417;
wire P2_R1131_U418 , P2_R1131_U419 , P2_R1131_U420 , P2_R1131_U421 , P2_R1131_U422 , P2_R1131_U423 , P2_R1131_U424 , P2_R1131_U425 , P2_R1131_U426 , P2_R1131_U427;
wire P2_R1131_U428 , P2_R1131_U429 , P2_R1131_U430 , P2_R1131_U431 , P2_R1131_U432 , P2_R1131_U433 , P2_R1131_U434 , P2_R1131_U435 , P2_R1131_U436 , P2_R1131_U437;
wire P2_R1131_U438 , P2_R1131_U439 , P2_R1131_U440 , P2_R1131_U441 , P2_R1131_U442 , P2_R1131_U443 , P2_R1131_U444 , P2_R1131_U445 , P2_R1131_U446 , P2_R1131_U447;
wire P2_R1131_U448 , P2_R1131_U449 , P2_R1131_U450 , P2_R1131_U451 , P2_R1131_U452 , P2_R1131_U453 , P2_R1131_U454 , P2_R1131_U455 , P2_R1131_U456 , P2_R1131_U457;
wire P2_R1131_U458 , P2_R1131_U459 , P2_R1131_U460 , P2_R1131_U461 , P2_R1131_U462 , P2_R1131_U463 , P2_R1131_U464 , P2_R1131_U465 , P2_R1131_U466 , P2_R1131_U467;
wire P2_R1131_U468 , P2_R1131_U469 , P2_R1131_U470 , P2_R1131_U471 , P2_R1131_U472 , P2_R1131_U473 , P2_R1131_U474 , P2_R1131_U475 , P2_R1131_U476 , P2_R1131_U477;
wire P2_R1131_U478 , P2_R1131_U479 , P2_R1131_U480 , P2_R1131_U481 , P2_R1131_U482 , P2_R1131_U483 , P2_R1131_U484 , P2_R1131_U485 , P2_R1131_U486 , P2_R1131_U487;
wire P2_R1131_U488 , P2_R1131_U489 , P2_R1131_U490 , P2_R1131_U491 , P2_R1131_U492 , P2_R1131_U493 , P2_R1131_U494 , P2_R1131_U495 , P2_R1131_U496 , P2_R1131_U497;
wire P2_R1131_U498 , P2_R1131_U499 , P2_R1131_U500 , P2_R1131_U501 , P2_R1131_U502 , P2_R1131_U503 , P2_R1131_U504 , P2_R1146_U6 , P2_R1146_U7 , P2_R1146_U8;
wire P2_R1146_U9 , P2_R1146_U10 , P2_R1146_U11 , P2_R1146_U12 , P2_R1146_U13 , P2_R1146_U14 , P2_R1146_U15 , P2_R1146_U16 , P2_R1146_U17 , P2_R1146_U18;
wire P2_R1146_U19 , P2_R1146_U20 , P2_R1146_U21 , P2_R1146_U22 , P2_R1146_U23 , P2_R1146_U24 , P2_R1146_U25 , P2_R1146_U26 , P2_R1146_U27 , P2_R1146_U28;
wire P2_R1146_U29 , P2_R1146_U30 , P2_R1146_U31 , P2_R1146_U32 , P2_R1146_U33 , P2_R1146_U34 , P2_R1146_U35 , P2_R1146_U36 , P2_R1146_U37 , P2_R1146_U38;
wire P2_R1146_U39 , P2_R1146_U40 , P2_R1146_U41 , P2_R1146_U42 , P2_R1146_U43 , P2_R1146_U44 , P2_R1146_U45 , P2_R1146_U46 , P2_R1146_U47 , P2_R1146_U48;
wire P2_R1146_U49 , P2_R1146_U50 , P2_R1146_U51 , P2_R1146_U52 , P2_R1146_U53 , P2_R1146_U54 , P2_R1146_U55 , P2_R1146_U56 , P2_R1146_U57 , P2_R1146_U58;
wire P2_R1146_U59 , P2_R1146_U60 , P2_R1146_U61 , P2_R1146_U62 , P2_R1146_U63 , P2_R1146_U64 , P2_R1146_U65 , P2_R1146_U66 , P2_R1146_U67 , P2_R1146_U68;
wire P2_R1146_U69 , P2_R1146_U70 , P2_R1146_U71 , P2_R1146_U72 , P2_R1146_U73 , P2_R1146_U74 , P2_R1146_U75 , P2_R1146_U76 , P2_R1146_U77 , P2_R1146_U78;
wire P2_R1146_U79 , P2_R1146_U80 , P2_R1146_U81 , P2_R1146_U82 , P2_R1146_U83 , P2_R1146_U84 , P2_R1146_U85 , P2_R1146_U86 , P2_R1146_U87 , P2_R1146_U88;
wire P2_R1146_U89 , P2_R1146_U90 , P2_R1146_U91 , P2_R1146_U92 , P2_R1146_U93 , P2_R1146_U94 , P2_R1146_U95 , P2_R1146_U96 , P2_R1146_U97 , P2_R1146_U98;
wire P2_R1146_U99 , P2_R1146_U100 , P2_R1146_U101 , P2_R1146_U102 , P2_R1146_U103 , P2_R1146_U104 , P2_R1146_U105 , P2_R1146_U106 , P2_R1146_U107 , P2_R1146_U108;
wire P2_R1146_U109 , P2_R1146_U110 , P2_R1146_U111 , P2_R1146_U112 , P2_R1146_U113 , P2_R1146_U114 , P2_R1146_U115 , P2_R1146_U116 , P2_R1146_U117 , P2_R1146_U118;
wire P2_R1146_U119 , P2_R1146_U120 , P2_R1146_U121 , P2_R1146_U122 , P2_R1146_U123 , P2_R1146_U124 , P2_R1146_U125 , P2_R1146_U126 , P2_R1146_U127 , P2_R1146_U128;
wire P2_R1146_U129 , P2_R1146_U130 , P2_R1146_U131 , P2_R1146_U132 , P2_R1146_U133 , P2_R1146_U134 , P2_R1146_U135 , P2_R1146_U136 , P2_R1146_U137 , P2_R1146_U138;
wire P2_R1146_U139 , P2_R1146_U140 , P2_R1146_U141 , P2_R1146_U142 , P2_R1146_U143 , P2_R1146_U144 , P2_R1146_U145 , P2_R1146_U146 , P2_R1146_U147 , P2_R1146_U148;
wire P2_R1146_U149 , P2_R1146_U150 , P2_R1146_U151 , P2_R1146_U152 , P2_R1146_U153 , P2_R1146_U154 , P2_R1146_U155 , P2_R1146_U156 , P2_R1146_U157 , P2_R1146_U158;
wire P2_R1146_U159 , P2_R1146_U160 , P2_R1146_U161 , P2_R1146_U162 , P2_R1146_U163 , P2_R1146_U164 , P2_R1146_U165 , P2_R1146_U166 , P2_R1146_U167 , P2_R1146_U168;
wire P2_R1146_U169 , P2_R1146_U170 , P2_R1146_U171 , P2_R1146_U172 , P2_R1146_U173 , P2_R1146_U174 , P2_R1146_U175 , P2_R1146_U176 , P2_R1146_U177 , P2_R1146_U178;
wire P2_R1146_U179 , P2_R1146_U180 , P2_R1146_U181 , P2_R1146_U182 , P2_R1146_U183 , P2_R1146_U184 , P2_R1146_U185 , P2_R1146_U186 , P2_R1146_U187 , P2_R1146_U188;
wire P2_R1146_U189 , P2_R1146_U190 , P2_R1146_U191 , P2_R1146_U192 , P2_R1146_U193 , P2_R1146_U194 , P2_R1146_U195 , P2_R1146_U196 , P2_R1146_U197 , P2_R1146_U198;
wire P2_R1146_U199 , P2_R1146_U200 , P2_R1146_U201 , P2_R1146_U202 , P2_R1146_U203 , P2_R1146_U204 , P2_R1146_U205 , P2_R1146_U206 , P2_R1146_U207 , P2_R1146_U208;
wire P2_R1146_U209 , P2_R1146_U210 , P2_R1146_U211 , P2_R1146_U212 , P2_R1146_U213 , P2_R1146_U214 , P2_R1146_U215 , P2_R1146_U216 , P2_R1146_U217 , P2_R1146_U218;
wire P2_R1146_U219 , P2_R1146_U220 , P2_R1146_U221 , P2_R1146_U222 , P2_R1146_U223 , P2_R1146_U224 , P2_R1146_U225 , P2_R1146_U226 , P2_R1146_U227 , P2_R1146_U228;
wire P2_R1146_U229 , P2_R1146_U230 , P2_R1146_U231 , P2_R1146_U232 , P2_R1146_U233 , P2_R1146_U234 , P2_R1146_U235 , P2_R1146_U236 , P2_R1146_U237 , P2_R1146_U238;
wire P2_R1146_U239 , P2_R1146_U240 , P2_R1146_U241 , P2_R1146_U242 , P2_R1146_U243 , P2_R1146_U244 , P2_R1146_U245 , P2_R1146_U246 , P2_R1146_U247 , P2_R1146_U248;
wire P2_R1146_U249 , P2_R1146_U250 , P2_R1146_U251 , P2_R1146_U252 , P2_R1146_U253 , P2_R1146_U254 , P2_R1146_U255 , P2_R1146_U256 , P2_R1146_U257 , P2_R1146_U258;
wire P2_R1146_U259 , P2_R1146_U260 , P2_R1146_U261 , P2_R1146_U262 , P2_R1146_U263 , P2_R1146_U264 , P2_R1146_U265 , P2_R1146_U266 , P2_R1146_U267 , P2_R1146_U268;
wire P2_R1146_U269 , P2_R1146_U270 , P2_R1146_U271 , P2_R1146_U272 , P2_R1146_U273 , P2_R1146_U274 , P2_R1146_U275 , P2_R1146_U276 , P2_R1146_U277 , P2_R1146_U278;
wire P2_R1146_U279 , P2_R1146_U280 , P2_R1146_U281 , P2_R1146_U282 , P2_R1146_U283 , P2_R1146_U284 , P2_R1146_U285 , P2_R1146_U286 , P2_R1146_U287 , P2_R1146_U288;
wire P2_R1146_U289 , P2_R1146_U290 , P2_R1146_U291 , P2_R1146_U292 , P2_R1146_U293 , P2_R1146_U294 , P2_R1146_U295 , P2_R1146_U296 , P2_R1146_U297 , P2_R1146_U298;
wire P2_R1146_U299 , P2_R1146_U300 , P2_R1146_U301 , P2_R1146_U302 , P2_R1146_U303 , P2_R1146_U304 , P2_R1146_U305 , P2_R1146_U306 , P2_R1146_U307 , P2_R1146_U308;
wire P2_R1146_U309 , P2_R1146_U310 , P2_R1146_U311 , P2_R1146_U312 , P2_R1146_U313 , P2_R1146_U314 , P2_R1146_U315 , P2_R1146_U316 , P2_R1146_U317 , P2_R1146_U318;
wire P2_R1146_U319 , P2_R1146_U320 , P2_R1146_U321 , P2_R1146_U322 , P2_R1146_U323 , P2_R1146_U324 , P2_R1146_U325 , P2_R1146_U326 , P2_R1146_U327 , P2_R1146_U328;
wire P2_R1146_U329 , P2_R1146_U330 , P2_R1146_U331 , P2_R1146_U332 , P2_R1146_U333 , P2_R1146_U334 , P2_R1146_U335 , P2_R1146_U336 , P2_R1146_U337 , P2_R1146_U338;
wire P2_R1146_U339 , P2_R1146_U340 , P2_R1146_U341 , P2_R1146_U342 , P2_R1146_U343 , P2_R1146_U344 , P2_R1146_U345 , P2_R1146_U346 , P2_R1146_U347 , P2_R1146_U348;
wire P2_R1146_U349 , P2_R1146_U350 , P2_R1146_U351 , P2_R1146_U352 , P2_R1146_U353 , P2_R1146_U354 , P2_R1146_U355 , P2_R1146_U356 , P2_R1146_U357 , P2_R1146_U358;
wire P2_R1146_U359 , P2_R1146_U360 , P2_R1146_U361 , P2_R1146_U362 , P2_R1146_U363 , P2_R1146_U364 , P2_R1146_U365 , P2_R1146_U366 , P2_R1146_U367 , P2_R1146_U368;
wire P2_R1146_U369 , P2_R1146_U370 , P2_R1146_U371 , P2_R1146_U372 , P2_R1146_U373 , P2_R1146_U374 , P2_R1146_U375 , P2_R1146_U376 , P2_R1146_U377 , P2_R1146_U378;
wire P2_R1146_U379 , P2_R1146_U380 , P2_R1146_U381 , P2_R1146_U382 , P2_R1146_U383 , P2_R1146_U384 , P2_R1146_U385 , P2_R1146_U386 , P2_R1146_U387 , P2_R1146_U388;
wire P2_R1146_U389 , P2_R1146_U390 , P2_R1146_U391 , P2_R1146_U392 , P2_R1146_U393 , P2_R1146_U394 , P2_R1146_U395 , P2_R1146_U396 , P2_R1146_U397 , P2_R1146_U398;
wire P2_R1146_U399 , P2_R1146_U400 , P2_R1146_U401 , P2_R1146_U402 , P2_R1146_U403 , P2_R1146_U404 , P2_R1146_U405 , P2_R1146_U406 , P2_R1146_U407 , P2_R1146_U408;
wire P2_R1146_U409 , P2_R1146_U410 , P2_R1146_U411 , P2_R1146_U412 , P2_R1146_U413 , P2_R1146_U414 , P2_R1146_U415 , P2_R1146_U416 , P2_R1146_U417 , P2_R1146_U418;
wire P2_R1146_U419 , P2_R1146_U420 , P2_R1146_U421 , P2_R1146_U422 , P2_R1146_U423 , P2_R1146_U424 , P2_R1146_U425 , P2_R1146_U426 , P2_R1146_U427 , P2_R1146_U428;
wire P2_R1146_U429 , P2_R1146_U430 , P2_R1146_U431 , P2_R1146_U432 , P2_R1146_U433 , P2_R1146_U434 , P2_R1146_U435 , P2_R1146_U436 , P2_R1146_U437 , P2_R1146_U438;
wire P2_R1146_U439 , P2_R1146_U440 , P2_R1146_U441 , P2_R1146_U442 , P2_R1146_U443 , P2_R1146_U444 , P2_R1146_U445 , P2_R1146_U446 , P2_R1146_U447 , P2_R1146_U448;
wire P2_R1146_U449 , P2_R1146_U450 , P2_R1146_U451 , P2_R1146_U452 , P2_R1146_U453 , P2_R1146_U454 , P2_R1146_U455 , P2_R1146_U456 , P2_R1146_U457 , P2_R1146_U458;
wire P2_R1146_U459 , P2_R1146_U460 , P2_R1146_U461 , P2_R1146_U462 , P2_R1146_U463 , P2_R1146_U464 , P2_R1146_U465 , P2_R1146_U466 , P2_R1146_U467 , P2_R1146_U468;
wire P2_R1146_U469 , P2_R1146_U470 , P2_R1146_U471 , P2_R1146_U472 , P2_R1146_U473 , P2_R1146_U474 , P2_R1146_U475 , P2_R1146_U476 , P2_R1146_U477 , P2_R1146_U478;
wire P2_R1203_U6 , P2_R1203_U7 , P2_R1203_U8 , P2_R1203_U9 , P2_R1203_U10 , P2_R1203_U11 , P2_R1203_U12 , P2_R1203_U13 , P2_R1203_U14 , P2_R1203_U15;
wire P2_R1203_U16 , P2_R1203_U17 , P2_R1203_U18 , P2_R1203_U19 , P2_R1203_U20 , P2_R1203_U21 , P2_R1203_U22 , P2_R1203_U23 , P2_R1203_U24 , P2_R1203_U25;
wire P2_R1203_U26 , P2_R1203_U27 , P2_R1203_U28 , P2_R1203_U29 , P2_R1203_U30 , P2_R1203_U31 , P2_R1203_U32 , P2_R1203_U33 , P2_R1203_U34 , P2_R1203_U35;
wire P2_R1203_U36 , P2_R1203_U37 , P2_R1203_U38 , P2_R1203_U39 , P2_R1203_U40 , P2_R1203_U41 , P2_R1203_U42 , P2_R1203_U43 , P2_R1203_U44 , P2_R1203_U45;
wire P2_R1203_U46 , P2_R1203_U47 , P2_R1203_U48 , P2_R1203_U49 , P2_R1203_U50 , P2_R1203_U51 , P2_R1203_U52 , P2_R1203_U53 , P2_R1203_U54 , P2_R1203_U55;
wire P2_R1203_U56 , P2_R1203_U57 , P2_R1203_U58 , P2_R1203_U59 , P2_R1203_U60 , P2_R1203_U61 , P2_R1203_U62 , P2_R1203_U63 , P2_R1203_U64 , P2_R1203_U65;
wire P2_R1203_U66 , P2_R1203_U67 , P2_R1203_U68 , P2_R1203_U69 , P2_R1203_U70 , P2_R1203_U71 , P2_R1203_U72 , P2_R1203_U73 , P2_R1203_U74 , P2_R1203_U75;
wire P2_R1203_U76 , P2_R1203_U77 , P2_R1203_U78 , P2_R1203_U79 , P2_R1203_U80 , P2_R1203_U81 , P2_R1203_U82 , P2_R1203_U83 , P2_R1203_U84 , P2_R1203_U85;
wire P2_R1203_U86 , P2_R1203_U87 , P2_R1203_U88 , P2_R1203_U89 , P2_R1203_U90 , P2_R1203_U91 , P2_R1203_U92 , P2_R1203_U93 , P2_R1203_U94 , P2_R1203_U95;
wire P2_R1203_U96 , P2_R1203_U97 , P2_R1203_U98 , P2_R1203_U99 , P2_R1203_U100 , P2_R1203_U101 , P2_R1203_U102 , P2_R1203_U103 , P2_R1203_U104 , P2_R1203_U105;
wire P2_R1203_U106 , P2_R1203_U107 , P2_R1203_U108 , P2_R1203_U109 , P2_R1203_U110 , P2_R1203_U111 , P2_R1203_U112 , P2_R1203_U113 , P2_R1203_U114 , P2_R1203_U115;
wire P2_R1203_U116 , P2_R1203_U117 , P2_R1203_U118 , P2_R1203_U119 , P2_R1203_U120 , P2_R1203_U121 , P2_R1203_U122 , P2_R1203_U123 , P2_R1203_U124 , P2_R1203_U125;
wire P2_R1203_U126 , P2_R1203_U127 , P2_R1203_U128 , P2_R1203_U129 , P2_R1203_U130 , P2_R1203_U131 , P2_R1203_U132 , P2_R1203_U133 , P2_R1203_U134 , P2_R1203_U135;
wire P2_R1203_U136 , P2_R1203_U137 , P2_R1203_U138 , P2_R1203_U139 , P2_R1203_U140 , P2_R1203_U141 , P2_R1203_U142 , P2_R1203_U143 , P2_R1203_U144 , P2_R1203_U145;
wire P2_R1203_U146 , P2_R1203_U147 , P2_R1203_U148 , P2_R1203_U149 , P2_R1203_U150 , P2_R1203_U151 , P2_R1203_U152 , P2_R1203_U153 , P2_R1203_U154 , P2_R1203_U155;
wire P2_R1203_U156 , P2_R1203_U157 , P2_R1203_U158 , P2_R1203_U159 , P2_R1203_U160 , P2_R1203_U161 , P2_R1203_U162 , P2_R1203_U163 , P2_R1203_U164 , P2_R1203_U165;
wire P2_R1203_U166 , P2_R1203_U167 , P2_R1203_U168 , P2_R1203_U169 , P2_R1203_U170 , P2_R1203_U171 , P2_R1203_U172 , P2_R1203_U173 , P2_R1203_U174 , P2_R1203_U175;
wire P2_R1203_U176 , P2_R1203_U177 , P2_R1203_U178 , P2_R1203_U179 , P2_R1203_U180 , P2_R1203_U181 , P2_R1203_U182 , P2_R1203_U183 , P2_R1203_U184 , P2_R1203_U185;
wire P2_R1203_U186 , P2_R1203_U187 , P2_R1203_U188 , P2_R1203_U189 , P2_R1203_U190 , P2_R1203_U191 , P2_R1203_U192 , P2_R1203_U193 , P2_R1203_U194 , P2_R1203_U195;
wire P2_R1203_U196 , P2_R1203_U197 , P2_R1203_U198 , P2_R1203_U199 , P2_R1203_U200 , P2_R1203_U201 , P2_R1203_U202 , P2_R1203_U203 , P2_R1203_U204 , P2_R1203_U205;
wire P2_R1203_U206 , P2_R1203_U207 , P2_R1203_U208 , P2_R1203_U209 , P2_R1203_U210 , P2_R1203_U211 , P2_R1203_U212 , P2_R1203_U213 , P2_R1203_U214 , P2_R1203_U215;
wire P2_R1203_U216 , P2_R1203_U217 , P2_R1203_U218 , P2_R1203_U219 , P2_R1203_U220 , P2_R1203_U221 , P2_R1203_U222 , P2_R1203_U223 , P2_R1203_U224 , P2_R1203_U225;
wire P2_R1203_U226 , P2_R1203_U227 , P2_R1203_U228 , P2_R1203_U229 , P2_R1203_U230 , P2_R1203_U231 , P2_R1203_U232 , P2_R1203_U233 , P2_R1203_U234 , P2_R1203_U235;
wire P2_R1203_U236 , P2_R1203_U237 , P2_R1203_U238 , P2_R1203_U239 , P2_R1203_U240 , P2_R1203_U241 , P2_R1203_U242 , P2_R1203_U243 , P2_R1203_U244 , P2_R1203_U245;
wire P2_R1203_U246 , P2_R1203_U247 , P2_R1203_U248 , P2_R1203_U249 , P2_R1203_U250 , P2_R1203_U251 , P2_R1203_U252 , P2_R1203_U253 , P2_R1203_U254 , P2_R1203_U255;
wire P2_R1203_U256 , P2_R1203_U257 , P2_R1203_U258 , P2_R1203_U259 , P2_R1203_U260 , P2_R1203_U261 , P2_R1203_U262 , P2_R1203_U263 , P2_R1203_U264 , P2_R1203_U265;
wire P2_R1203_U266 , P2_R1203_U267 , P2_R1203_U268 , P2_R1203_U269 , P2_R1203_U270 , P2_R1203_U271 , P2_R1203_U272 , P2_R1203_U273 , P2_R1203_U274 , P2_R1203_U275;
wire P2_R1203_U276 , P2_R1203_U277 , P2_R1203_U278 , P2_R1203_U279 , P2_R1203_U280 , P2_R1203_U281 , P2_R1203_U282 , P2_R1203_U283 , P2_R1203_U284 , P2_R1203_U285;
wire P2_R1203_U286 , P2_R1203_U287 , P2_R1203_U288 , P2_R1203_U289 , P2_R1203_U290 , P2_R1203_U291 , P2_R1203_U292 , P2_R1203_U293 , P2_R1203_U294 , P2_R1203_U295;
wire P2_R1203_U296 , P2_R1203_U297 , P2_R1203_U298 , P2_R1203_U299 , P2_R1203_U300 , P2_R1203_U301 , P2_R1203_U302 , P2_R1203_U303 , P2_R1203_U304 , P2_R1203_U305;
wire P2_R1203_U306 , P2_R1203_U307 , P2_R1203_U308 , P2_R1203_U309 , P2_R1203_U310 , P2_R1203_U311 , P2_R1203_U312 , P2_R1203_U313 , P2_R1203_U314 , P2_R1203_U315;
wire P2_R1203_U316 , P2_R1203_U317 , P2_R1203_U318 , P2_R1203_U319 , P2_R1203_U320 , P2_R1203_U321 , P2_R1203_U322 , P2_R1203_U323 , P2_R1203_U324 , P2_R1203_U325;
wire P2_R1203_U326 , P2_R1203_U327 , P2_R1203_U328 , P2_R1203_U329 , P2_R1203_U330 , P2_R1203_U331 , P2_R1203_U332 , P2_R1203_U333 , P2_R1203_U334 , P2_R1203_U335;
wire P2_R1203_U336 , P2_R1203_U337 , P2_R1203_U338 , P2_R1203_U339 , P2_R1203_U340 , P2_R1203_U341 , P2_R1203_U342 , P2_R1203_U343 , P2_R1203_U344 , P2_R1203_U345;
wire P2_R1203_U346 , P2_R1203_U347 , P2_R1203_U348 , P2_R1203_U349 , P2_R1203_U350 , P2_R1203_U351 , P2_R1203_U352 , P2_R1203_U353 , P2_R1203_U354 , P2_R1203_U355;
wire P2_R1203_U356 , P2_R1203_U357 , P2_R1203_U358 , P2_R1203_U359 , P2_R1203_U360 , P2_R1203_U361 , P2_R1203_U362 , P2_R1203_U363 , P2_R1203_U364 , P2_R1203_U365;
wire P2_R1203_U366 , P2_R1203_U367 , P2_R1203_U368 , P2_R1203_U369 , P2_R1203_U370 , P2_R1203_U371 , P2_R1203_U372 , P2_R1203_U373 , P2_R1203_U374 , P2_R1203_U375;
wire P2_R1203_U376 , P2_R1203_U377 , P2_R1203_U378 , P2_R1203_U379 , P2_R1203_U380 , P2_R1203_U381 , P2_R1203_U382 , P2_R1203_U383 , P2_R1203_U384 , P2_R1203_U385;
wire P2_R1203_U386 , P2_R1203_U387 , P2_R1203_U388 , P2_R1203_U389 , P2_R1203_U390 , P2_R1203_U391 , P2_R1203_U392 , P2_R1203_U393 , P2_R1203_U394 , P2_R1203_U395;
wire P2_R1203_U396 , P2_R1203_U397 , P2_R1203_U398 , P2_R1203_U399 , P2_R1203_U400 , P2_R1203_U401 , P2_R1203_U402 , P2_R1203_U403 , P2_R1203_U404 , P2_R1203_U405;
wire P2_R1203_U406 , P2_R1203_U407 , P2_R1203_U408 , P2_R1203_U409 , P2_R1203_U410 , P2_R1203_U411 , P2_R1203_U412 , P2_R1203_U413 , P2_R1203_U414 , P2_R1203_U415;
wire P2_R1203_U416 , P2_R1203_U417 , P2_R1203_U418 , P2_R1203_U419 , P2_R1203_U420 , P2_R1203_U421 , P2_R1203_U422 , P2_R1203_U423 , P2_R1203_U424 , P2_R1203_U425;
wire P2_R1203_U426 , P2_R1203_U427 , P2_R1203_U428 , P2_R1203_U429 , P2_R1203_U430 , P2_R1203_U431 , P2_R1203_U432 , P2_R1203_U433 , P2_R1203_U434 , P2_R1203_U435;
wire P2_R1203_U436 , P2_R1203_U437 , P2_R1203_U438 , P2_R1203_U439 , P2_R1203_U440 , P2_R1203_U441 , P2_R1203_U442 , P2_R1203_U443 , P2_R1203_U444 , P2_R1203_U445;
wire P2_R1203_U446 , P2_R1203_U447 , P2_R1203_U448 , P2_R1203_U449 , P2_R1203_U450 , P2_R1203_U451 , P2_R1203_U452 , P2_R1203_U453 , P2_R1203_U454 , P2_R1203_U455;
wire P2_R1203_U456 , P2_R1203_U457 , P2_R1203_U458 , P2_R1203_U459 , P2_R1203_U460 , P2_R1203_U461 , P2_R1203_U462 , P2_R1203_U463 , P2_R1203_U464 , P2_R1203_U465;
wire P2_R1203_U466 , P2_R1203_U467 , P2_R1203_U468 , P2_R1203_U469 , P2_R1203_U470 , P2_R1203_U471 , P2_R1203_U472 , P2_R1203_U473 , P2_R1203_U474 , P2_R1203_U475;
wire P2_R1203_U476 , P2_R1203_U477 , P2_R1203_U478 , P2_R1113_U6 , P2_R1113_U7 , P2_R1113_U8 , P2_R1113_U9 , P2_R1113_U10 , P2_R1113_U11 , P2_R1113_U12;
wire P2_R1113_U13 , P2_R1113_U14 , P2_R1113_U15 , P2_R1113_U16 , P2_R1113_U17 , P2_R1113_U18 , P2_R1113_U19 , P2_R1113_U20 , P2_R1113_U21 , P2_R1113_U22;
wire P2_R1113_U23 , P2_R1113_U24 , P2_R1113_U25 , P2_R1113_U26 , P2_R1113_U27 , P2_R1113_U28 , P2_R1113_U29 , P2_R1113_U30 , P2_R1113_U31 , P2_R1113_U32;
wire P2_R1113_U33 , P2_R1113_U34 , P2_R1113_U35 , P2_R1113_U36 , P2_R1113_U37 , P2_R1113_U38 , P2_R1113_U39 , P2_R1113_U40 , P2_R1113_U41 , P2_R1113_U42;
wire P2_R1113_U43 , P2_R1113_U44 , P2_R1113_U45 , P2_R1113_U46 , P2_R1113_U47 , P2_R1113_U48 , P2_R1113_U49 , P2_R1113_U50 , P2_R1113_U51 , P2_R1113_U52;
wire P2_R1113_U53 , P2_R1113_U54 , P2_R1113_U55 , P2_R1113_U56 , P2_R1113_U57 , P2_R1113_U58 , P2_R1113_U59 , P2_R1113_U60 , P2_R1113_U61 , P2_R1113_U62;
wire P2_R1113_U63 , P2_R1113_U64 , P2_R1113_U65 , P2_R1113_U66 , P2_R1113_U67 , P2_R1113_U68 , P2_R1113_U69 , P2_R1113_U70 , P2_R1113_U71 , P2_R1113_U72;
wire P2_R1113_U73 , P2_R1113_U74 , P2_R1113_U75 , P2_R1113_U76 , P2_R1113_U77 , P2_R1113_U78 , P2_R1113_U79 , P2_R1113_U80 , P2_R1113_U81 , P2_R1113_U82;
wire P2_R1113_U83 , P2_R1113_U84 , P2_R1113_U85 , P2_R1113_U86 , P2_R1113_U87 , P2_R1113_U88 , P2_R1113_U89 , P2_R1113_U90 , P2_R1113_U91 , P2_R1113_U92;
wire P2_R1113_U93 , P2_R1113_U94 , P2_R1113_U95 , P2_R1113_U96 , P2_R1113_U97 , P2_R1113_U98 , P2_R1113_U99 , P2_R1113_U100 , P2_R1113_U101 , P2_R1113_U102;
wire P2_R1113_U103 , P2_R1113_U104 , P2_R1113_U105 , P2_R1113_U106 , P2_R1113_U107 , P2_R1113_U108 , P2_R1113_U109 , P2_R1113_U110 , P2_R1113_U111 , P2_R1113_U112;
wire P2_R1113_U113 , P2_R1113_U114 , P2_R1113_U115 , P2_R1113_U116 , P2_R1113_U117 , P2_R1113_U118 , P2_R1113_U119 , P2_R1113_U120 , P2_R1113_U121 , P2_R1113_U122;
wire P2_R1113_U123 , P2_R1113_U124 , P2_R1113_U125 , P2_R1113_U126 , P2_R1113_U127 , P2_R1113_U128 , P2_R1113_U129 , P2_R1113_U130 , P2_R1113_U131 , P2_R1113_U132;
wire P2_R1113_U133 , P2_R1113_U134 , P2_R1113_U135 , P2_R1113_U136 , P2_R1113_U137 , P2_R1113_U138 , P2_R1113_U139 , P2_R1113_U140 , P2_R1113_U141 , P2_R1113_U142;
wire P2_R1113_U143 , P2_R1113_U144 , P2_R1113_U145 , P2_R1113_U146 , P2_R1113_U147 , P2_R1113_U148 , P2_R1113_U149 , P2_R1113_U150 , P2_R1113_U151 , P2_R1113_U152;
wire P2_R1113_U153 , P2_R1113_U154 , P2_R1113_U155 , P2_R1113_U156 , P2_R1113_U157 , P2_R1113_U158 , P2_R1113_U159 , P2_R1113_U160 , P2_R1113_U161 , P2_R1113_U162;
wire P2_R1113_U163 , P2_R1113_U164 , P2_R1113_U165 , P2_R1113_U166 , P2_R1113_U167 , P2_R1113_U168 , P2_R1113_U169 , P2_R1113_U170 , P2_R1113_U171 , P2_R1113_U172;
wire P2_R1113_U173 , P2_R1113_U174 , P2_R1113_U175 , P2_R1113_U176 , P2_R1113_U177 , P2_R1113_U178 , P2_R1113_U179 , P2_R1113_U180 , P2_R1113_U181 , P2_R1113_U182;
wire P2_R1113_U183 , P2_R1113_U184 , P2_R1113_U185 , P2_R1113_U186 , P2_R1113_U187 , P2_R1113_U188 , P2_R1113_U189 , P2_R1113_U190 , P2_R1113_U191 , P2_R1113_U192;
wire P2_R1113_U193 , P2_R1113_U194 , P2_R1113_U195 , P2_R1113_U196 , P2_R1113_U197 , P2_R1113_U198 , P2_R1113_U199 , P2_R1113_U200 , P2_R1113_U201 , P2_R1113_U202;
wire P2_R1113_U203 , P2_R1113_U204 , P2_R1113_U205 , P2_R1113_U206 , P2_R1113_U207 , P2_R1113_U208 , P2_R1113_U209 , P2_R1113_U210 , P2_R1113_U211 , P2_R1113_U212;
wire P2_R1113_U213 , P2_R1113_U214 , P2_R1113_U215 , P2_R1113_U216 , P2_R1113_U217 , P2_R1113_U218 , P2_R1113_U219 , P2_R1113_U220 , P2_R1113_U221 , P2_R1113_U222;
wire P2_R1113_U223 , P2_R1113_U224 , P2_R1113_U225 , P2_R1113_U226 , P2_R1113_U227 , P2_R1113_U228 , P2_R1113_U229 , P2_R1113_U230 , P2_R1113_U231 , P2_R1113_U232;
wire P2_R1113_U233 , P2_R1113_U234 , P2_R1113_U235 , P2_R1113_U236 , P2_R1113_U237 , P2_R1113_U238 , P2_R1113_U239 , P2_R1113_U240 , P2_R1113_U241 , P2_R1113_U242;
wire P2_R1113_U243 , P2_R1113_U244 , P2_R1113_U245 , P2_R1113_U246 , P2_R1113_U247 , P2_R1113_U248 , P2_R1113_U249 , P2_R1113_U250 , P2_R1113_U251 , P2_R1113_U252;
wire P2_R1113_U253 , P2_R1113_U254 , P2_R1113_U255 , P2_R1113_U256 , P2_R1113_U257 , P2_R1113_U258 , P2_R1113_U259 , P2_R1113_U260 , P2_R1113_U261 , P2_R1113_U262;
wire P2_R1113_U263 , P2_R1113_U264 , P2_R1113_U265 , P2_R1113_U266 , P2_R1113_U267 , P2_R1113_U268 , P2_R1113_U269 , P2_R1113_U270 , P2_R1113_U271 , P2_R1113_U272;
wire P2_R1113_U273 , P2_R1113_U274 , P2_R1113_U275 , P2_R1113_U276 , P2_R1113_U277 , P2_R1113_U278 , P2_R1113_U279 , P2_R1113_U280 , P2_R1113_U281 , P2_R1113_U282;
wire P2_R1113_U283 , P2_R1113_U284 , P2_R1113_U285 , P2_R1113_U286 , P2_R1113_U287 , P2_R1113_U288 , P2_R1113_U289 , P2_R1113_U290 , P2_R1113_U291 , P2_R1113_U292;
wire P2_R1113_U293 , P2_R1113_U294 , P2_R1113_U295 , P2_R1113_U296 , P2_R1113_U297 , P2_R1113_U298 , P2_R1113_U299 , P2_R1113_U300 , P2_R1113_U301 , P2_R1113_U302;
wire P2_R1113_U303 , P2_R1113_U304 , P2_R1113_U305 , P2_R1113_U306 , P2_R1113_U307 , P2_R1113_U308 , P2_R1113_U309 , P2_R1113_U310 , P2_R1113_U311 , P2_R1113_U312;
wire P2_R1113_U313 , P2_R1113_U314 , P2_R1113_U315 , P2_R1113_U316 , P2_R1113_U317 , P2_R1113_U318 , P2_R1113_U319 , P2_R1113_U320 , P2_R1113_U321 , P2_R1113_U322;
wire P2_R1113_U323 , P2_R1113_U324 , P2_R1113_U325 , P2_R1113_U326 , P2_R1113_U327 , P2_R1113_U328 , P2_R1113_U329 , P2_R1113_U330 , P2_R1113_U331 , P2_R1113_U332;
wire P2_R1113_U333 , P2_R1113_U334 , P2_R1113_U335 , P2_R1113_U336 , P2_R1113_U337 , P2_R1113_U338 , P2_R1113_U339 , P2_R1113_U340 , P2_R1113_U341 , P2_R1113_U342;
wire P2_R1113_U343 , P2_R1113_U344 , P2_R1113_U345 , P2_R1113_U346 , P2_R1113_U347 , P2_R1113_U348 , P2_R1113_U349 , P2_R1113_U350 , P2_R1113_U351 , P2_R1113_U352;
wire P2_R1113_U353 , P2_R1113_U354 , P2_R1113_U355 , P2_R1113_U356 , P2_R1113_U357 , P2_R1113_U358 , P2_R1113_U359 , P2_R1113_U360 , P2_R1113_U361 , P2_R1113_U362;
wire P2_R1113_U363 , P2_R1113_U364 , P2_R1113_U365 , P2_R1113_U366 , P2_R1113_U367 , P2_R1113_U368 , P2_R1113_U369 , P2_R1113_U370 , P2_R1113_U371 , P2_R1113_U372;
wire P2_R1113_U373 , P2_R1113_U374 , P2_R1113_U375 , P2_R1113_U376 , P2_R1113_U377 , P2_R1113_U378 , P2_R1113_U379 , P2_R1113_U380 , P2_R1113_U381 , P2_R1113_U382;
wire P2_R1113_U383 , P2_R1113_U384 , P2_R1113_U385 , P2_R1113_U386 , P2_R1113_U387 , P2_R1113_U388 , P2_R1113_U389 , P2_R1113_U390 , P2_R1113_U391 , P2_R1113_U392;
wire P2_R1113_U393 , P2_R1113_U394 , P2_R1113_U395 , P2_R1113_U396 , P2_R1113_U397 , P2_R1113_U398 , P2_R1113_U399 , P2_R1113_U400 , P2_R1113_U401 , P2_R1113_U402;
wire P2_R1113_U403 , P2_R1113_U404 , P2_R1113_U405 , P2_R1113_U406 , P2_R1113_U407 , P2_R1113_U408 , P2_R1113_U409 , P2_R1113_U410 , P2_R1113_U411 , P2_R1113_U412;
wire P2_R1113_U413 , P2_R1113_U414 , P2_R1113_U415 , P2_R1113_U416 , P2_R1113_U417 , P2_R1113_U418 , P2_R1113_U419 , P2_R1113_U420 , P2_R1113_U421 , P2_R1113_U422;
wire P2_R1113_U423 , P2_R1113_U424 , P2_R1113_U425 , P2_R1113_U426 , P2_R1113_U427 , P2_R1113_U428 , P2_R1113_U429 , P2_R1113_U430 , P2_R1113_U431 , P2_R1113_U432;
wire P2_R1113_U433 , P2_R1113_U434 , P2_R1113_U435 , P2_R1113_U436 , P2_R1113_U437 , P2_R1113_U438 , P2_R1113_U439 , P2_R1113_U440 , P2_R1113_U441 , P2_R1113_U442;
wire P2_R1113_U443 , P2_R1113_U444 , P2_R1113_U445 , P2_R1113_U446 , P2_R1113_U447 , P2_R1113_U448 , P2_R1113_U449 , P2_R1113_U450 , P2_R1113_U451 , P2_R1113_U452;
wire P2_R1113_U453 , P2_R1113_U454 , P2_R1113_U455 , P2_R1113_U456 , P2_R1113_U457 , P2_R1113_U458 , P2_R1113_U459 , P2_R1113_U460 , P2_R1113_U461 , P2_R1113_U462;
wire P2_R1113_U463 , P2_R1113_U464 , P2_R1113_U465 , P2_R1113_U466 , P2_R1113_U467 , P2_R1113_U468 , P2_R1113_U469 , P2_R1113_U470 , P2_R1113_U471 , P2_R1113_U472;
wire P2_R1113_U473 , P2_R1113_U474 , P2_R1113_U475 , P2_R1113_U476 , P2_R1113_U477 , P2_R1113_U478 , P3_SUB_598_U6 , P3_SUB_598_U7 , P3_SUB_598_U8 , P3_SUB_598_U9;
wire P3_SUB_598_U10 , P3_SUB_598_U11 , P3_SUB_598_U12 , P3_SUB_598_U13 , P3_SUB_598_U14 , P3_SUB_598_U15 , P3_SUB_598_U16 , P3_SUB_598_U17 , P3_SUB_598_U18 , P3_SUB_598_U19;
wire P3_SUB_598_U20 , P3_SUB_598_U21 , P3_SUB_598_U22 , P3_SUB_598_U23 , P3_SUB_598_U24 , P3_SUB_598_U25 , P3_SUB_598_U26 , P3_SUB_598_U27 , P3_SUB_598_U28 , P3_SUB_598_U29;
wire P3_SUB_598_U30 , P3_SUB_598_U31 , P3_SUB_598_U32 , P3_SUB_598_U33 , P3_SUB_598_U34 , P3_SUB_598_U35 , P3_SUB_598_U36 , P3_SUB_598_U37 , P3_SUB_598_U38 , P3_SUB_598_U39;
wire P3_SUB_598_U40 , P3_SUB_598_U41 , P3_SUB_598_U42 , P3_SUB_598_U43 , P3_SUB_598_U44 , P3_SUB_598_U45 , P3_SUB_598_U46 , P3_SUB_598_U47 , P3_SUB_598_U48 , P3_SUB_598_U49;
wire P3_SUB_598_U50 , P3_SUB_598_U51 , P3_SUB_598_U52 , P3_SUB_598_U53 , P3_SUB_598_U54 , P3_SUB_598_U55 , P3_SUB_598_U56 , P3_SUB_598_U57 , P3_SUB_598_U58 , P3_SUB_598_U59;
wire P3_SUB_598_U60 , P3_SUB_598_U61 , P3_SUB_598_U62 , P3_SUB_598_U63 , P3_SUB_598_U64 , P3_SUB_598_U65 , P3_SUB_598_U66 , P3_SUB_598_U67 , P3_SUB_598_U68 , P3_SUB_598_U69;
wire P3_SUB_598_U70 , P3_SUB_598_U71 , P3_SUB_598_U72 , P3_SUB_598_U73 , P3_SUB_598_U74 , P3_SUB_598_U75 , P3_SUB_598_U76 , P3_SUB_598_U77 , P3_SUB_598_U78 , P3_SUB_598_U79;
wire P3_SUB_598_U80 , P3_SUB_598_U81 , P3_SUB_598_U82 , P3_SUB_598_U83 , P3_SUB_598_U84 , P3_SUB_598_U85 , P3_SUB_598_U86 , P3_SUB_598_U87 , P3_SUB_598_U88 , P3_SUB_598_U89;
wire P3_SUB_598_U90 , P3_SUB_598_U91 , P3_SUB_598_U92 , P3_SUB_598_U93 , P3_SUB_598_U94 , P3_SUB_598_U95 , P3_SUB_598_U96 , P3_SUB_598_U97 , P3_SUB_598_U98 , P3_SUB_598_U99;
wire P3_SUB_598_U100 , P3_SUB_598_U101 , P3_SUB_598_U102 , P3_SUB_598_U103 , P3_SUB_598_U104 , P3_SUB_598_U105 , P3_SUB_598_U106 , P3_SUB_598_U107 , P3_SUB_598_U108 , P3_SUB_598_U109;
wire P3_SUB_598_U110 , P3_SUB_598_U111 , P3_SUB_598_U112 , P3_SUB_598_U113 , P3_SUB_598_U114 , P3_SUB_598_U115 , P3_SUB_598_U116 , P3_SUB_598_U117 , P3_SUB_598_U118 , P3_SUB_598_U119;
wire P3_SUB_598_U120 , P3_SUB_598_U121 , P3_SUB_598_U122 , P3_SUB_598_U123 , P3_SUB_598_U124 , P3_SUB_598_U125 , P3_SUB_598_U126 , P3_SUB_598_U127 , P3_SUB_598_U128 , P3_SUB_598_U129;
wire P3_SUB_598_U130 , P3_SUB_598_U131 , P3_SUB_598_U132 , P3_SUB_598_U133 , P3_SUB_598_U134 , P3_SUB_598_U135 , P3_SUB_598_U136 , P3_SUB_598_U137 , P3_SUB_598_U138 , P3_SUB_598_U139;
wire P3_SUB_598_U140 , P3_SUB_598_U141 , P3_SUB_598_U142 , P3_SUB_598_U143 , P3_SUB_598_U144 , P3_SUB_598_U145 , P3_SUB_598_U146 , P3_SUB_598_U147 , P3_SUB_598_U148 , P3_SUB_598_U149;
wire P3_SUB_598_U150 , P3_SUB_598_U151 , P3_SUB_598_U152 , P3_SUB_598_U153 , P3_SUB_598_U154 , P3_SUB_598_U155 , P3_SUB_598_U156 , P3_SUB_598_U157 , P3_SUB_598_U158 , P3_SUB_598_U159;
wire P3_SUB_598_U160 , P3_R693_U6 , P3_R693_U7 , P3_R693_U8 , P3_R693_U9 , P3_R693_U10 , P3_R693_U11 , P3_R693_U12 , P3_R693_U13 , P3_R693_U14;
wire P3_R693_U15 , P3_R693_U16 , P3_R693_U17 , P3_R693_U18 , P3_R693_U19 , P3_R693_U20 , P3_R693_U21 , P3_R693_U22 , P3_R693_U23 , P3_R693_U24;
wire P3_R693_U25 , P3_R693_U26 , P3_R693_U27 , P3_R693_U28 , P3_R693_U29 , P3_R693_U30 , P3_R693_U31 , P3_R693_U32 , P3_R693_U33 , P3_R693_U34;
wire P3_R693_U35 , P3_R693_U36 , P3_R693_U37 , P3_R693_U38 , P3_R693_U39 , P3_R693_U40 , P3_R693_U41 , P3_R693_U42 , P3_R693_U43 , P3_R693_U44;
wire P3_R693_U45 , P3_R693_U46 , P3_R693_U47 , P3_R693_U48 , P3_R693_U49 , P3_R693_U50 , P3_R693_U51 , P3_R693_U52 , P3_R693_U53 , P3_R693_U54;
wire P3_R693_U55 , P3_R693_U56 , P3_R693_U57 , P3_R693_U58 , P3_R693_U59 , P3_R693_U60 , P3_R693_U61 , P3_R693_U62 , P3_R693_U63 , P3_R693_U64;
wire P3_R693_U65 , P3_R693_U66 , P3_R693_U67 , P3_R693_U68 , P3_R693_U69 , P3_R693_U70 , P3_R693_U71 , P3_R693_U72 , P3_R693_U73 , P3_R693_U74;
wire P3_R693_U75 , P3_R693_U76 , P3_R693_U77 , P3_R693_U78 , P3_R693_U79 , P3_R693_U80 , P3_R693_U81 , P3_R693_U82 , P3_R693_U83 , P3_R693_U84;
wire P3_R693_U85 , P3_R693_U86 , P3_R693_U87 , P3_R693_U88 , P3_R693_U89 , P3_R693_U90 , P3_R693_U91 , P3_R693_U92 , P3_R693_U93 , P3_R693_U94;
wire P3_R693_U95 , P3_R693_U96 , P3_R693_U97 , P3_R693_U98 , P3_R693_U99 , P3_R693_U100 , P3_R693_U101 , P3_R693_U102 , P3_R693_U103 , P3_R693_U104;
wire P3_R693_U105 , P3_R693_U106 , P3_R693_U107 , P3_R693_U108 , P3_R693_U109 , P3_R693_U110 , P3_R693_U111 , P3_R693_U112 , P3_R693_U113 , P3_R693_U114;
wire P3_R693_U115 , P3_R693_U116 , P3_R693_U117 , P3_R693_U118 , P3_R693_U119 , P3_R693_U120 , P3_R693_U121 , P3_R693_U122 , P3_R693_U123 , P3_R693_U124;
wire P3_R693_U125 , P3_R693_U126 , P3_R693_U127 , P3_R693_U128 , P3_R693_U129 , P3_R693_U130 , P3_R693_U131 , P3_R693_U132 , P3_R693_U133 , P3_R693_U134;
wire P3_R693_U135 , P3_R693_U136 , P3_R693_U137 , P3_R693_U138 , P3_R693_U139 , P3_R693_U140 , P3_R693_U141 , P3_R693_U142 , P3_R693_U143 , P3_R693_U144;
wire P3_R693_U145 , P3_R693_U146 , P3_R693_U147 , P3_R693_U148 , P3_R693_U149 , P3_R693_U150 , P3_R693_U151 , P3_R693_U152 , P3_R693_U153 , P3_R693_U154;
wire P3_R693_U155 , P3_R693_U156 , P3_R693_U157 , P3_R693_U158 , P3_R693_U159 , P3_R693_U160 , P3_R693_U161 , P3_R693_U162 , P3_R693_U163 , P3_R693_U164;
wire P3_R693_U165 , P3_R693_U166 , P3_R693_U167 , P3_R693_U168 , P3_R693_U169 , P3_R693_U170 , P3_R693_U171 , P3_R693_U172 , P3_R693_U173 , P3_R693_U174;
wire P3_R693_U175 , P3_R693_U176 , P3_R693_U177 , P3_R693_U178 , P3_R693_U179 , P3_R693_U180 , P3_R693_U181 , P3_R693_U182 , P3_R693_U183 , P3_R693_U184;
wire P3_R693_U185 , P3_R693_U186 , P3_R693_U187 , P3_R693_U188 , P3_R693_U189 , P3_R693_U190 , P3_R693_U191 , P3_R693_U192 , P3_R693_U193 , P3_R693_U194;
wire P3_R693_U195 , P3_R693_U196 , P3_SUB_609_U6 , P3_SUB_609_U7 , P3_SUB_609_U8 , P3_SUB_609_U9 , P3_SUB_609_U10 , P3_SUB_609_U11 , P3_SUB_609_U12 , P3_SUB_609_U13;
wire P3_SUB_609_U14 , P3_SUB_609_U15 , P3_SUB_609_U16 , P3_SUB_609_U17 , P3_SUB_609_U18 , P3_SUB_609_U19 , P3_SUB_609_U20 , P3_SUB_609_U21 , P3_SUB_609_U22 , P3_SUB_609_U23;
wire P3_SUB_609_U24 , P3_SUB_609_U25 , P3_SUB_609_U26 , P3_SUB_609_U27 , P3_SUB_609_U28 , P3_SUB_609_U29 , P3_SUB_609_U30 , P3_SUB_609_U31 , P3_SUB_609_U32 , P3_SUB_609_U33;
wire P3_SUB_609_U34 , P3_SUB_609_U35 , P3_SUB_609_U36 , P3_SUB_609_U37 , P3_SUB_609_U38 , P3_SUB_609_U39 , P3_SUB_609_U40 , P3_SUB_609_U41 , P3_SUB_609_U42 , P3_SUB_609_U43;
wire P3_SUB_609_U44 , P3_SUB_609_U45 , P3_SUB_609_U46 , P3_SUB_609_U47 , P3_SUB_609_U48 , P3_SUB_609_U49 , P3_SUB_609_U50 , P3_SUB_609_U51 , P3_SUB_609_U52 , P3_SUB_609_U53;
wire P3_SUB_609_U54 , P3_SUB_609_U55 , P3_SUB_609_U56 , P3_SUB_609_U57 , P3_SUB_609_U58 , P3_SUB_609_U59 , P3_SUB_609_U60 , P3_SUB_609_U61 , P3_SUB_609_U62 , P3_SUB_609_U63;
wire P3_SUB_609_U64 , P3_SUB_609_U65 , P3_SUB_609_U66 , P3_SUB_609_U67 , P3_SUB_609_U68 , P3_SUB_609_U69 , P3_SUB_609_U70 , P3_SUB_609_U71 , P3_SUB_609_U72 , P3_SUB_609_U73;
wire P3_SUB_609_U74 , P3_SUB_609_U75 , P3_SUB_609_U76 , P3_SUB_609_U77 , P3_SUB_609_U78 , P3_SUB_609_U79 , P3_SUB_609_U80 , P3_SUB_609_U81 , P3_SUB_609_U82 , P3_SUB_609_U83;
wire P3_SUB_609_U84 , P3_SUB_609_U85 , P3_SUB_609_U86 , P3_SUB_609_U87 , P3_SUB_609_U88 , P3_SUB_609_U89 , P3_SUB_609_U90 , P3_SUB_609_U91 , P3_SUB_609_U92 , P3_SUB_609_U93;
wire P3_SUB_609_U94 , P3_SUB_609_U95 , P3_SUB_609_U96 , P3_SUB_609_U97 , P3_SUB_609_U98 , P3_SUB_609_U99 , P3_SUB_609_U100 , P3_SUB_609_U101 , P3_SUB_609_U102 , P3_SUB_609_U103;
wire P3_SUB_609_U104 , P3_SUB_609_U105 , P3_SUB_609_U106 , P3_SUB_609_U107 , P3_SUB_609_U108 , P3_SUB_609_U109 , P3_SUB_609_U110 , P3_SUB_609_U111 , P3_SUB_609_U112 , P3_SUB_609_U113;
wire P3_SUB_609_U114 , P3_SUB_609_U115 , P3_R1095_U6 , P3_R1095_U7 , P3_R1095_U8 , P3_R1095_U9 , P3_R1095_U10 , P3_R1095_U11 , P3_R1095_U12 , P3_R1095_U13;
wire P3_R1095_U14 , P3_R1095_U15 , P3_R1095_U16 , P3_R1095_U17 , P3_R1095_U18 , P3_R1095_U19 , P3_R1095_U20 , P3_R1095_U21 , P3_R1095_U22 , P3_R1095_U23;
wire P3_R1095_U24 , P3_R1095_U25 , P3_R1095_U26 , P3_R1095_U27 , P3_R1095_U28 , P3_R1095_U29 , P3_R1095_U30 , P3_R1095_U31 , P3_R1095_U32 , P3_R1095_U33;
wire P3_R1095_U34 , P3_R1095_U35 , P3_R1095_U36 , P3_R1095_U37 , P3_R1095_U38 , P3_R1095_U39 , P3_R1095_U40 , P3_R1095_U41 , P3_R1095_U42 , P3_R1095_U43;
wire P3_R1095_U44 , P3_R1095_U45 , P3_R1095_U46 , P3_R1095_U47 , P3_R1095_U48 , P3_R1095_U49 , P3_R1095_U50 , P3_R1095_U51 , P3_R1095_U52 , P3_R1095_U53;
wire P3_R1095_U54 , P3_R1095_U55 , P3_R1095_U56 , P3_R1095_U57 , P3_R1095_U58 , P3_R1095_U59 , P3_R1095_U60 , P3_R1095_U61 , P3_R1095_U62 , P3_R1095_U63;
wire P3_R1095_U64 , P3_R1095_U65 , P3_R1095_U66 , P3_R1095_U67 , P3_R1095_U68 , P3_R1095_U69 , P3_R1095_U70 , P3_R1095_U71 , P3_R1095_U72 , P3_R1095_U73;
wire P3_R1095_U74 , P3_R1095_U75 , P3_R1095_U76 , P3_R1095_U77 , P3_R1095_U78 , P3_R1095_U79 , P3_R1095_U80 , P3_R1095_U81 , P3_R1095_U82 , P3_R1095_U83;
wire P3_R1095_U84 , P3_R1095_U85 , P3_R1095_U86 , P3_R1095_U87 , P3_R1095_U88 , P3_R1095_U89 , P3_R1095_U90 , P3_R1095_U91 , P3_R1095_U92 , P3_R1095_U93;
wire P3_R1095_U94 , P3_R1095_U95 , P3_R1095_U96 , P3_R1095_U97 , P3_R1095_U98 , P3_R1095_U99 , P3_R1095_U100 , P3_R1095_U101 , P3_R1095_U102 , P3_R1095_U103;
wire P3_R1095_U104 , P3_R1095_U105 , P3_R1095_U106 , P3_R1095_U107 , P3_R1095_U108 , P3_R1095_U109 , P3_R1095_U110 , P3_R1095_U111 , P3_R1095_U112 , P3_R1095_U113;
wire P3_R1095_U114 , P3_R1095_U115 , P3_R1095_U116 , P3_R1095_U117 , P3_R1095_U118 , P3_R1095_U119 , P3_R1095_U120 , P3_R1095_U121 , P3_R1095_U122 , P3_R1095_U123;
wire P3_R1095_U124 , P3_R1095_U125 , P3_R1095_U126 , P3_R1095_U127 , P3_R1095_U128 , P3_R1095_U129 , P3_R1095_U130 , P3_R1095_U131 , P3_R1095_U132 , P3_R1095_U133;
wire P3_R1095_U134 , P3_R1095_U135 , P3_R1095_U136 , P3_R1095_U137 , P3_R1095_U138 , P3_R1095_U139 , P3_R1095_U140 , P3_R1095_U141 , P3_R1095_U142 , P3_R1095_U143;
wire P3_R1095_U144 , P3_R1095_U145 , P3_R1095_U146 , P3_R1095_U147 , P3_R1095_U148 , P3_R1095_U149 , P3_R1095_U150 , P3_R1095_U151 , P3_R1095_U152 , P3_R1095_U153;
wire P3_R1095_U154 , P3_R1095_U155 , P3_R1095_U156 , P3_R1095_U157 , P3_R1095_U158 , P3_R1095_U159 , P3_R1095_U160 , P3_R1095_U161 , P3_R1095_U162 , P3_R1095_U163;
wire P3_R1095_U164 , P3_R1095_U165 , P3_R1095_U166 , P3_R1095_U167 , P3_R1095_U168 , P3_R1095_U169 , P3_R1095_U170 , P3_R1095_U171 , P3_R1095_U172 , P3_R1095_U173;
wire P3_R1095_U174 , P3_R1095_U175 , P3_R1095_U176 , P3_R1095_U177 , P3_R1095_U178 , P3_R1095_U179 , P3_R1095_U180 , P3_R1095_U181 , P3_R1095_U182 , P3_R1095_U183;
wire P3_R1095_U184 , P3_R1095_U185 , P3_R1095_U186 , P3_R1095_U187 , P3_R1095_U188 , P3_R1095_U189 , P3_R1095_U190 , P3_R1095_U191 , P3_R1095_U192 , P3_R1095_U193;
wire P3_R1095_U194 , P3_R1095_U195 , P3_R1095_U196 , P3_R1095_U197 , P3_R1095_U198 , P3_R1095_U199 , P3_R1095_U200 , P3_R1095_U201 , P3_R1095_U202 , P3_R1095_U203;
wire P3_R1095_U204 , P3_R1095_U205 , P3_R1095_U206 , P3_R1095_U207 , P3_R1095_U208 , P3_R1095_U209 , P3_R1095_U210 , P3_R1095_U211 , P3_R1095_U212 , P3_R1095_U213;
wire P3_R1095_U214 , P3_R1095_U215 , P3_R1095_U216 , P3_R1095_U217 , P3_R1095_U218 , P3_R1095_U219 , P3_R1095_U220 , P3_R1095_U221 , P3_R1095_U222 , P3_R1095_U223;
wire P3_R1095_U224 , P3_R1095_U225 , P3_R1095_U226 , P3_R1095_U227 , P3_R1095_U228 , P3_R1095_U229 , P3_R1095_U230 , P3_R1095_U231 , P3_R1095_U232 , P3_R1095_U233;
wire P3_R1095_U234 , P3_R1095_U235 , P3_R1095_U236 , P3_R1095_U237 , P3_R1095_U238 , P3_R1095_U239 , P3_R1095_U240 , P3_R1095_U241 , P3_R1095_U242 , P3_R1095_U243;
wire P3_R1095_U244 , P3_R1095_U245 , P3_R1095_U246 , P3_R1095_U247 , P3_R1095_U248 , P3_R1095_U249 , P3_R1095_U250 , P3_R1095_U251 , P3_R1095_U252 , P3_R1095_U253;
wire P3_R1095_U254 , P3_R1095_U255 , P3_R1095_U256 , P3_R1095_U257 , P3_R1095_U258 , P3_R1095_U259 , P3_R1095_U260 , P3_R1095_U261 , P3_R1095_U262 , P3_R1095_U263;
wire P3_R1095_U264 , P3_R1095_U265 , P3_R1095_U266 , P3_R1095_U267 , P3_R1095_U268 , P3_R1095_U269 , P3_R1095_U270 , P3_R1095_U271 , P3_R1095_U272 , P3_R1095_U273;
wire P3_R1095_U274 , P3_R1095_U275 , P3_R1095_U276 , P3_R1095_U277 , P3_R1095_U278 , P3_R1095_U279 , P3_R1095_U280 , P3_R1095_U281 , P3_R1095_U282 , P3_R1095_U283;
wire P3_R1095_U284 , P3_R1095_U285 , P3_R1095_U286 , P3_R1095_U287 , P3_R1095_U288 , P3_R1095_U289 , P3_R1095_U290 , P3_R1095_U291 , P3_R1095_U292 , P3_R1095_U293;
wire P3_R1095_U294 , P3_R1095_U295 , P3_R1095_U296 , P3_R1095_U297 , P3_R1095_U298 , P3_R1095_U299 , P3_R1095_U300 , P3_R1095_U301 , P3_R1095_U302 , P3_R1095_U303;
wire P3_R1095_U304 , P3_R1095_U305 , P3_R1095_U306 , P3_R1095_U307 , P3_R1095_U308 , P3_R1095_U309 , P3_R1095_U310 , P3_R1095_U311 , P3_R1095_U312 , P3_R1095_U313;
wire P3_R1095_U314 , P3_R1095_U315 , P3_R1095_U316 , P3_R1095_U317 , P3_R1095_U318 , P3_R1095_U319 , P3_R1095_U320 , P3_R1095_U321 , P3_R1095_U322 , P3_R1095_U323;
wire P3_R1095_U324 , P3_R1095_U325 , P3_R1095_U326 , P3_R1095_U327 , P3_R1095_U328 , P3_R1095_U329 , P3_R1095_U330 , P3_R1095_U331 , P3_R1095_U332 , P3_R1095_U333;
wire P3_R1095_U334 , P3_R1095_U335 , P3_R1095_U336 , P3_R1095_U337 , P3_R1095_U338 , P3_R1095_U339 , P3_R1095_U340 , P3_R1095_U341 , P3_R1095_U342 , P3_R1095_U343;
wire P3_R1095_U344 , P3_R1095_U345 , P3_R1095_U346 , P3_R1095_U347 , P3_R1095_U348 , P3_R1095_U349 , P3_R1095_U350 , P3_R1095_U351 , P3_R1095_U352 , P3_R1095_U353;
wire P3_R1095_U354 , P3_R1095_U355 , P3_R1095_U356 , P3_R1095_U357 , P3_R1095_U358 , P3_R1095_U359 , P3_R1095_U360 , P3_R1095_U361 , P3_R1095_U362 , P3_R1095_U363;
wire P3_R1095_U364 , P3_R1095_U365 , P3_R1095_U366 , P3_R1095_U367 , P3_R1095_U368 , P3_R1095_U369 , P3_R1095_U370 , P3_R1095_U371 , P3_R1095_U372 , P3_R1095_U373;
wire P3_R1095_U374 , P3_R1095_U375 , P3_R1095_U376 , P3_R1095_U377 , P3_R1095_U378 , P3_R1095_U379 , P3_R1095_U380 , P3_R1095_U381 , P3_R1095_U382 , P3_R1095_U383;
wire P3_R1095_U384 , P3_R1095_U385 , P3_R1095_U386 , P3_R1095_U387 , P3_R1095_U388 , P3_R1095_U389 , P3_R1095_U390 , P3_R1095_U391 , P3_R1095_U392 , P3_R1095_U393;
wire P3_R1095_U394 , P3_R1095_U395 , P3_R1095_U396 , P3_R1095_U397 , P3_R1095_U398 , P3_R1095_U399 , P3_R1095_U400 , P3_R1095_U401 , P3_R1095_U402 , P3_R1095_U403;
wire P3_R1095_U404 , P3_R1095_U405 , P3_R1095_U406 , P3_R1095_U407 , P3_R1095_U408 , P3_R1095_U409 , P3_R1095_U410 , P3_R1095_U411 , P3_R1095_U412 , P3_R1095_U413;
wire P3_R1095_U414 , P3_R1095_U415 , P3_R1095_U416 , P3_R1095_U417 , P3_R1095_U418 , P3_R1095_U419 , P3_R1095_U420 , P3_R1095_U421 , P3_R1095_U422 , P3_R1095_U423;
wire P3_R1095_U424 , P3_R1095_U425 , P3_R1095_U426 , P3_R1095_U427 , P3_R1095_U428 , P3_R1095_U429 , P3_R1095_U430 , P3_R1095_U431 , P3_R1095_U432 , P3_R1095_U433;
wire P3_R1095_U434 , P3_R1095_U435 , P3_R1095_U436 , P3_R1095_U437 , P3_R1095_U438 , P3_R1095_U439 , P3_R1095_U440 , P3_R1095_U441 , P3_R1095_U442 , P3_R1095_U443;
wire P3_R1095_U444 , P3_R1095_U445 , P3_R1095_U446 , P3_R1095_U447 , P3_R1095_U448 , P3_R1095_U449 , P3_R1095_U450 , P3_R1095_U451 , P3_R1095_U452 , P3_R1095_U453;
wire P3_R1095_U454 , P3_R1095_U455 , P3_R1095_U456 , P3_R1095_U457 , P3_R1095_U458 , P3_R1095_U459 , P3_R1095_U460 , P3_R1095_U461 , P3_R1095_U462 , P3_R1095_U463;
wire P3_R1095_U464 , P3_R1095_U465 , P3_R1095_U466 , P3_R1095_U467 , P3_R1095_U468 , P3_R1095_U469 , P3_R1095_U470 , P3_R1095_U471 , P3_R1095_U472 , P3_R1095_U473;
wire P3_R1095_U474 , P3_R1095_U475 , P3_R1095_U476 , P3_R1095_U477 , P3_R1095_U478 , P3_R1095_U479 , P3_R1095_U480 , P3_R1095_U481 , P3_R1095_U482 , P3_R1095_U483;
wire P3_R1095_U484 , P3_R1095_U485 , P3_R1212_U6 , P3_R1212_U7 , P3_R1212_U8 , P3_R1212_U9 , P3_R1212_U10 , P3_R1212_U11 , P3_R1212_U12 , P3_R1212_U13;
wire P3_R1212_U14 , P3_R1212_U15 , P3_R1212_U16 , P3_R1212_U17 , P3_R1212_U18 , P3_R1212_U19 , P3_R1212_U20 , P3_R1212_U21 , P3_R1212_U22 , P3_R1212_U23;
wire P3_R1212_U24 , P3_R1212_U25 , P3_R1212_U26 , P3_R1212_U27 , P3_R1212_U28 , P3_R1212_U29 , P3_R1212_U30 , P3_R1212_U31 , P3_R1212_U32 , P3_R1212_U33;
wire P3_R1212_U34 , P3_R1212_U35 , P3_R1212_U36 , P3_R1212_U37 , P3_R1212_U38 , P3_R1212_U39 , P3_R1212_U40 , P3_R1212_U41 , P3_R1212_U42 , P3_R1212_U43;
wire P3_R1212_U44 , P3_R1212_U45 , P3_R1212_U46 , P3_R1212_U47 , P3_R1212_U48 , P3_R1212_U49 , P3_R1212_U50 , P3_R1212_U51 , P3_R1212_U52 , P3_R1212_U53;
wire P3_R1212_U54 , P3_R1212_U55 , P3_R1212_U56 , P3_R1212_U57 , P3_R1212_U58 , P3_R1212_U59 , P3_R1212_U60 , P3_R1212_U61 , P3_R1212_U62 , P3_R1212_U63;
wire P3_R1212_U64 , P3_R1212_U65 , P3_R1212_U66 , P3_R1212_U67 , P3_R1212_U68 , P3_R1212_U69 , P3_R1212_U70 , P3_R1212_U71 , P3_R1212_U72 , P3_R1212_U73;
wire P3_R1212_U74 , P3_R1212_U75 , P3_R1212_U76 , P3_R1212_U77 , P3_R1212_U78 , P3_R1212_U79 , P3_R1212_U80 , P3_R1212_U81 , P3_R1212_U82 , P3_R1212_U83;
wire P3_R1212_U84 , P3_R1212_U85 , P3_R1212_U86 , P3_R1212_U87 , P3_R1212_U88 , P3_R1212_U89 , P3_R1212_U90 , P3_R1212_U91 , P3_R1212_U92 , P3_R1212_U93;
wire P3_R1212_U94 , P3_R1212_U95 , P3_R1212_U96 , P3_R1212_U97 , P3_R1212_U98 , P3_R1212_U99 , P3_R1212_U100 , P3_R1212_U101 , P3_R1212_U102 , P3_R1212_U103;
wire P3_R1212_U104 , P3_R1212_U105 , P3_R1212_U106 , P3_R1212_U107 , P3_R1212_U108 , P3_R1212_U109 , P3_R1212_U110 , P3_R1212_U111 , P3_R1212_U112 , P3_R1212_U113;
wire P3_R1212_U114 , P3_R1212_U115 , P3_R1212_U116 , P3_R1212_U117 , P3_R1212_U118 , P3_R1212_U119 , P3_R1212_U120 , P3_R1212_U121 , P3_R1212_U122 , P3_R1212_U123;
wire P3_R1212_U124 , P3_R1212_U125 , P3_R1212_U126 , P3_R1212_U127 , P3_R1212_U128 , P3_R1212_U129 , P3_R1212_U130 , P3_R1212_U131 , P3_R1212_U132 , P3_R1212_U133;
wire P3_R1212_U134 , P3_R1212_U135 , P3_R1212_U136 , P3_R1212_U137 , P3_R1212_U138 , P3_R1212_U139 , P3_R1212_U140 , P3_R1212_U141 , P3_R1212_U142 , P3_R1212_U143;
wire P3_R1212_U144 , P3_R1212_U145 , P3_R1212_U146 , P3_R1212_U147 , P3_R1212_U148 , P3_R1212_U149 , P3_R1212_U150 , P3_R1212_U151 , P3_R1212_U152 , P3_R1212_U153;
wire P3_R1212_U154 , P3_R1212_U155 , P3_R1212_U156 , P3_R1212_U157 , P3_R1212_U158 , P3_R1212_U159 , P3_R1212_U160 , P3_R1212_U161 , P3_R1212_U162 , P3_R1212_U163;
wire P3_R1212_U164 , P3_R1212_U165 , P3_R1212_U166 , P3_R1212_U167 , P3_R1212_U168 , P3_R1212_U169 , P3_R1212_U170 , P3_R1212_U171 , P3_R1212_U172 , P3_R1212_U173;
wire P3_R1212_U174 , P3_R1212_U175 , P3_R1212_U176 , P3_R1212_U177 , P3_R1212_U178 , P3_R1212_U179 , P3_R1212_U180 , P3_R1212_U181 , P3_R1212_U182 , P3_R1212_U183;
wire P3_R1212_U184 , P3_R1212_U185 , P3_R1212_U186 , P3_R1212_U187 , P3_R1212_U188 , P3_R1212_U189 , P3_R1212_U190 , P3_R1212_U191 , P3_R1212_U192 , P3_R1212_U193;
wire P3_R1212_U194 , P3_R1212_U195 , P3_R1212_U196 , P3_R1212_U197 , P3_R1212_U198 , P3_R1212_U199 , P3_R1212_U200 , P3_R1212_U201 , P3_R1212_U202 , P3_R1212_U203;
wire P3_R1212_U204 , P3_R1212_U205 , P3_R1212_U206 , P3_R1212_U207 , P3_R1212_U208 , P3_R1212_U209 , P3_R1212_U210 , P3_R1212_U211 , P3_R1212_U212 , P3_R1212_U213;
wire P3_R1212_U214 , P3_R1212_U215 , P3_R1212_U216 , P3_R1212_U217 , P3_R1212_U218 , P3_R1212_U219 , P3_R1212_U220 , P3_R1212_U221 , P3_R1212_U222 , P3_R1212_U223;
wire P3_R1212_U224 , P3_R1212_U225 , P3_R1212_U226 , P3_R1212_U227 , P3_R1212_U228 , P3_R1212_U229 , P3_R1212_U230 , P3_R1212_U231 , P3_R1212_U232 , P3_R1212_U233;
wire P3_R1212_U234 , P3_R1212_U235 , P3_R1212_U236 , P3_R1212_U237 , P3_R1212_U238 , P3_R1212_U239 , P3_R1212_U240 , P3_R1212_U241 , P3_R1212_U242 , P3_R1212_U243;
wire P3_R1212_U244 , P3_R1212_U245 , P3_R1212_U246 , P3_R1212_U247 , P3_R1212_U248 , P3_R1212_U249 , P3_R1212_U250 , P3_R1212_U251 , P3_R1212_U252 , P3_R1212_U253;
wire P3_R1212_U254 , P3_R1212_U255 , P3_R1212_U256 , P3_R1212_U257 , P3_R1212_U258 , P3_R1212_U259 , P3_R1212_U260 , P3_R1212_U261 , P3_R1212_U262 , P3_R1212_U263;
wire P3_R1212_U264 , P3_R1212_U265 , P3_R1212_U266 , P3_R1212_U267 , P3_R1212_U268 , P3_R1212_U269 , P3_R1212_U270 , P3_R1212_U271 , P3_R1212_U272 , P3_R1212_U273;
wire P3_R1212_U274 , P3_R1212_U275 , P3_R1212_U276 , P3_R1209_U6 , P3_R1209_U7 , P3_R1209_U8 , P3_R1209_U9 , P3_R1209_U10 , P3_R1209_U11 , P3_R1209_U12;
wire P3_R1209_U13 , P3_R1209_U14 , P3_R1209_U15 , P3_R1209_U16 , P3_R1209_U17 , P3_R1209_U18 , P3_R1209_U19 , P3_R1209_U20 , P3_R1209_U21 , P3_R1209_U22;
wire P3_R1209_U23 , P3_R1209_U24 , P3_R1209_U25 , P3_R1209_U26 , P3_R1209_U27 , P3_R1209_U28 , P3_R1209_U29 , P3_R1209_U30 , P3_R1209_U31 , P3_R1209_U32;
wire P3_R1209_U33 , P3_R1209_U34 , P3_R1209_U35 , P3_R1209_U36 , P3_R1209_U37 , P3_R1209_U38 , P3_R1209_U39 , P3_R1209_U40 , P3_R1209_U41 , P3_R1209_U42;
wire P3_R1209_U43 , P3_R1209_U44 , P3_R1209_U45 , P3_R1209_U46 , P3_R1209_U47 , P3_R1209_U48 , P3_R1209_U49 , P3_R1209_U50 , P3_R1209_U51 , P3_R1209_U52;
wire P3_R1209_U53 , P3_R1209_U54 , P3_R1209_U55 , P3_R1209_U56 , P3_R1209_U57 , P3_R1209_U58 , P3_R1209_U59 , P3_R1209_U60 , P3_R1209_U61 , P3_R1209_U62;
wire P3_R1209_U63 , P3_R1209_U64 , P3_R1209_U65 , P3_R1209_U66 , P3_R1209_U67 , P3_R1209_U68 , P3_R1209_U69 , P3_R1209_U70 , P3_R1209_U71 , P3_R1209_U72;
wire P3_R1209_U73 , P3_R1209_U74 , P3_R1209_U75 , P3_R1209_U76 , P3_R1209_U77 , P3_R1209_U78 , P3_R1209_U79 , P3_R1209_U80 , P3_R1209_U81 , P3_R1209_U82;
wire P3_R1209_U83 , P3_R1209_U84 , P3_R1209_U85 , P3_R1209_U86 , P3_R1209_U87 , P3_R1209_U88 , P3_R1209_U89 , P3_R1209_U90 , P3_R1209_U91 , P3_R1209_U92;
wire P3_R1209_U93 , P3_R1209_U94 , P3_R1209_U95 , P3_R1209_U96 , P3_R1209_U97 , P3_R1209_U98 , P3_R1209_U99 , P3_R1209_U100 , P3_R1209_U101 , P3_R1209_U102;
wire P3_R1209_U103 , P3_R1209_U104 , P3_R1209_U105 , P3_R1209_U106 , P3_R1209_U107 , P3_R1209_U108 , P3_R1209_U109 , P3_R1209_U110 , P3_R1209_U111 , P3_R1209_U112;
wire P3_R1209_U113 , P3_R1209_U114 , P3_R1209_U115 , P3_R1209_U116 , P3_R1209_U117 , P3_R1209_U118 , P3_R1209_U119 , P3_R1209_U120 , P3_R1209_U121 , P3_R1209_U122;
wire P3_R1209_U123 , P3_R1209_U124 , P3_R1209_U125 , P3_R1209_U126 , P3_R1209_U127 , P3_R1209_U128 , P3_R1209_U129 , P3_R1209_U130 , P3_R1209_U131 , P3_R1209_U132;
wire P3_R1209_U133 , P3_R1209_U134 , P3_R1209_U135 , P3_R1209_U136 , P3_R1209_U137 , P3_R1209_U138 , P3_R1209_U139 , P3_R1209_U140 , P3_R1209_U141 , P3_R1209_U142;
wire P3_R1209_U143 , P3_R1209_U144 , P3_R1209_U145 , P3_R1209_U146 , P3_R1209_U147 , P3_R1209_U148 , P3_R1209_U149 , P3_R1209_U150 , P3_R1209_U151 , P3_R1209_U152;
wire P3_R1209_U153 , P3_R1209_U154 , P3_R1209_U155 , P3_R1209_U156 , P3_R1209_U157 , P3_R1209_U158 , P3_R1209_U159 , P3_R1209_U160 , P3_R1209_U161 , P3_R1209_U162;
wire P3_R1209_U163 , P3_R1209_U164 , P3_R1209_U165 , P3_R1209_U166 , P3_R1209_U167 , P3_R1209_U168 , P3_R1209_U169 , P3_R1209_U170 , P3_R1209_U171 , P3_R1209_U172;
wire P3_R1209_U173 , P3_R1209_U174 , P3_R1209_U175 , P3_R1209_U176 , P3_R1209_U177 , P3_R1209_U178 , P3_R1209_U179 , P3_R1209_U180 , P3_R1209_U181 , P3_R1209_U182;
wire P3_R1209_U183 , P3_R1209_U184 , P3_R1209_U185 , P3_R1209_U186 , P3_R1209_U187 , P3_R1209_U188 , P3_R1209_U189 , P3_R1209_U190 , P3_R1209_U191 , P3_R1209_U192;
wire P3_R1209_U193 , P3_R1209_U194 , P3_R1209_U195 , P3_R1209_U196 , P3_R1209_U197 , P3_R1209_U198 , P3_R1209_U199 , P3_R1209_U200 , P3_R1209_U201 , P3_R1209_U202;
wire P3_R1209_U203 , P3_R1209_U204 , P3_R1209_U205 , P3_R1209_U206 , P3_R1209_U207 , P3_R1209_U208 , P3_R1209_U209 , P3_R1209_U210 , P3_R1209_U211 , P3_R1209_U212;
wire P3_R1209_U213 , P3_R1209_U214 , P3_R1209_U215 , P3_R1209_U216 , P3_R1209_U217 , P3_R1209_U218 , P3_R1209_U219 , P3_R1209_U220 , P3_R1209_U221 , P3_R1209_U222;
wire P3_R1209_U223 , P3_R1209_U224 , P3_R1209_U225 , P3_R1209_U226 , P3_R1209_U227 , P3_R1209_U228 , P3_R1209_U229 , P3_R1209_U230 , P3_R1209_U231 , P3_R1209_U232;
wire P3_R1209_U233 , P3_R1209_U234 , P3_R1209_U235 , P3_R1209_U236 , P3_R1209_U237 , P3_R1209_U238 , P3_R1209_U239 , P3_R1209_U240 , P3_R1209_U241 , P3_R1209_U242;
wire P3_R1209_U243 , P3_R1209_U244 , P3_R1209_U245 , P3_R1209_U246 , P3_R1209_U247 , P3_R1209_U248 , P3_R1209_U249 , P3_R1209_U250 , P3_R1209_U251 , P3_R1209_U252;
wire P3_R1209_U253 , P3_R1209_U254 , P3_R1209_U255 , P3_R1209_U256 , P3_R1209_U257 , P3_R1209_U258 , P3_R1209_U259 , P3_R1209_U260 , P3_R1209_U261 , P3_R1209_U262;
wire P3_R1209_U263 , P3_R1209_U264 , P3_R1209_U265 , P3_R1209_U266 , P3_R1209_U267 , P3_R1209_U268 , P3_R1209_U269 , P3_R1209_U270 , P3_R1209_U271 , P3_R1209_U272;
wire P3_R1209_U273 , P3_R1209_U274 , P3_R1209_U275 , P3_R1209_U276 , P3_R1300_U6 , P3_R1300_U7 , P3_R1300_U8 , P3_R1300_U9 , P3_R1300_U10 , P3_R1200_U6;
wire P3_R1200_U7 , P3_R1200_U8 , P3_R1200_U9 , P3_R1200_U10 , P3_R1200_U11 , P3_R1200_U12 , P3_R1200_U13 , P3_R1200_U14 , P3_R1200_U15 , P3_R1200_U16;
wire P3_R1200_U17 , P3_R1200_U18 , P3_R1200_U19 , P3_R1200_U20 , P3_R1200_U21 , P3_R1200_U22 , P3_R1200_U23 , P3_R1200_U24 , P3_R1200_U25 , P3_R1200_U26;
wire P3_R1200_U27 , P3_R1200_U28 , P3_R1200_U29 , P3_R1200_U30 , P3_R1200_U31 , P3_R1200_U32 , P3_R1200_U33 , P3_R1200_U34 , P3_R1200_U35 , P3_R1200_U36;
wire P3_R1200_U37 , P3_R1200_U38 , P3_R1200_U39 , P3_R1200_U40 , P3_R1200_U41 , P3_R1200_U42 , P3_R1200_U43 , P3_R1200_U44 , P3_R1200_U45 , P3_R1200_U46;
wire P3_R1200_U47 , P3_R1200_U48 , P3_R1200_U49 , P3_R1200_U50 , P3_R1200_U51 , P3_R1200_U52 , P3_R1200_U53 , P3_R1200_U54 , P3_R1200_U55 , P3_R1200_U56;
wire P3_R1200_U57 , P3_R1200_U58 , P3_R1200_U59 , P3_R1200_U60 , P3_R1200_U61 , P3_R1200_U62 , P3_R1200_U63 , P3_R1200_U64 , P3_R1200_U65 , P3_R1200_U66;
wire P3_R1200_U67 , P3_R1200_U68 , P3_R1200_U69 , P3_R1200_U70 , P3_R1200_U71 , P3_R1200_U72 , P3_R1200_U73 , P3_R1200_U74 , P3_R1200_U75 , P3_R1200_U76;
wire P3_R1200_U77 , P3_R1200_U78 , P3_R1200_U79 , P3_R1200_U80 , P3_R1200_U81 , P3_R1200_U82 , P3_R1200_U83 , P3_R1200_U84 , P3_R1200_U85 , P3_R1200_U86;
wire P3_R1200_U87 , P3_R1200_U88 , P3_R1200_U89 , P3_R1200_U90 , P3_R1200_U91 , P3_R1200_U92 , P3_R1200_U93 , P3_R1200_U94 , P3_R1200_U95 , P3_R1200_U96;
wire P3_R1200_U97 , P3_R1200_U98 , P3_R1200_U99 , P3_R1200_U100 , P3_R1200_U101 , P3_R1200_U102 , P3_R1200_U103 , P3_R1200_U104 , P3_R1200_U105 , P3_R1200_U106;
wire P3_R1200_U107 , P3_R1200_U108 , P3_R1200_U109 , P3_R1200_U110 , P3_R1200_U111 , P3_R1200_U112 , P3_R1200_U113 , P3_R1200_U114 , P3_R1200_U115 , P3_R1200_U116;
wire P3_R1200_U117 , P3_R1200_U118 , P3_R1200_U119 , P3_R1200_U120 , P3_R1200_U121 , P3_R1200_U122 , P3_R1200_U123 , P3_R1200_U124 , P3_R1200_U125 , P3_R1200_U126;
wire P3_R1200_U127 , P3_R1200_U128 , P3_R1200_U129 , P3_R1200_U130 , P3_R1200_U131 , P3_R1200_U132 , P3_R1200_U133 , P3_R1200_U134 , P3_R1200_U135 , P3_R1200_U136;
wire P3_R1200_U137 , P3_R1200_U138 , P3_R1200_U139 , P3_R1200_U140 , P3_R1200_U141 , P3_R1200_U142 , P3_R1200_U143 , P3_R1200_U144 , P3_R1200_U145 , P3_R1200_U146;
wire P3_R1200_U147 , P3_R1200_U148 , P3_R1200_U149 , P3_R1200_U150 , P3_R1200_U151 , P3_R1200_U152 , P3_R1200_U153 , P3_R1200_U154 , P3_R1200_U155 , P3_R1200_U156;
wire P3_R1200_U157 , P3_R1200_U158 , P3_R1200_U159 , P3_R1200_U160 , P3_R1200_U161 , P3_R1200_U162 , P3_R1200_U163 , P3_R1200_U164 , P3_R1200_U165 , P3_R1200_U166;
wire P3_R1200_U167 , P3_R1200_U168 , P3_R1200_U169 , P3_R1200_U170 , P3_R1200_U171 , P3_R1200_U172 , P3_R1200_U173 , P3_R1200_U174 , P3_R1200_U175 , P3_R1200_U176;
wire P3_R1200_U177 , P3_R1200_U178 , P3_R1200_U179 , P3_R1200_U180 , P3_R1200_U181 , P3_R1200_U182 , P3_R1200_U183 , P3_R1200_U184 , P3_R1200_U185 , P3_R1200_U186;
wire P3_R1200_U187 , P3_R1200_U188 , P3_R1200_U189 , P3_R1200_U190 , P3_R1200_U191 , P3_R1200_U192 , P3_R1200_U193 , P3_R1200_U194 , P3_R1200_U195 , P3_R1200_U196;
wire P3_R1200_U197 , P3_R1200_U198 , P3_R1200_U199 , P3_R1200_U200 , P3_R1200_U201 , P3_R1200_U202 , P3_R1200_U203 , P3_R1200_U204 , P3_R1200_U205 , P3_R1200_U206;
wire P3_R1200_U207 , P3_R1200_U208 , P3_R1200_U209 , P3_R1200_U210 , P3_R1200_U211 , P3_R1200_U212 , P3_R1200_U213 , P3_R1200_U214 , P3_R1200_U215 , P3_R1200_U216;
wire P3_R1200_U217 , P3_R1200_U218 , P3_R1200_U219 , P3_R1200_U220 , P3_R1200_U221 , P3_R1200_U222 , P3_R1200_U223 , P3_R1200_U224 , P3_R1200_U225 , P3_R1200_U226;
wire P3_R1200_U227 , P3_R1200_U228 , P3_R1200_U229 , P3_R1200_U230 , P3_R1200_U231 , P3_R1200_U232 , P3_R1200_U233 , P3_R1200_U234 , P3_R1200_U235 , P3_R1200_U236;
wire P3_R1200_U237 , P3_R1200_U238 , P3_R1200_U239 , P3_R1200_U240 , P3_R1200_U241 , P3_R1200_U242 , P3_R1200_U243 , P3_R1200_U244 , P3_R1200_U245 , P3_R1200_U246;
wire P3_R1200_U247 , P3_R1200_U248 , P3_R1200_U249 , P3_R1200_U250 , P3_R1200_U251 , P3_R1200_U252 , P3_R1200_U253 , P3_R1200_U254 , P3_R1200_U255 , P3_R1200_U256;
wire P3_R1200_U257 , P3_R1200_U258 , P3_R1200_U259 , P3_R1200_U260 , P3_R1200_U261 , P3_R1200_U262 , P3_R1200_U263 , P3_R1200_U264 , P3_R1200_U265 , P3_R1200_U266;
wire P3_R1200_U267 , P3_R1200_U268 , P3_R1200_U269 , P3_R1200_U270 , P3_R1200_U271 , P3_R1200_U272 , P3_R1200_U273 , P3_R1200_U274 , P3_R1200_U275 , P3_R1200_U276;
wire P3_R1200_U277 , P3_R1200_U278 , P3_R1200_U279 , P3_R1200_U280 , P3_R1200_U281 , P3_R1200_U282 , P3_R1200_U283 , P3_R1200_U284 , P3_R1200_U285 , P3_R1200_U286;
wire P3_R1200_U287 , P3_R1200_U288 , P3_R1200_U289 , P3_R1200_U290 , P3_R1200_U291 , P3_R1200_U292 , P3_R1200_U293 , P3_R1200_U294 , P3_R1200_U295 , P3_R1200_U296;
wire P3_R1200_U297 , P3_R1200_U298 , P3_R1200_U299 , P3_R1200_U300 , P3_R1200_U301 , P3_R1200_U302 , P3_R1200_U303 , P3_R1200_U304 , P3_R1200_U305 , P3_R1200_U306;
wire P3_R1200_U307 , P3_R1200_U308 , P3_R1200_U309 , P3_R1200_U310 , P3_R1200_U311 , P3_R1200_U312 , P3_R1200_U313 , P3_R1200_U314 , P3_R1200_U315 , P3_R1200_U316;
wire P3_R1200_U317 , P3_R1200_U318 , P3_R1200_U319 , P3_R1200_U320 , P3_R1200_U321 , P3_R1200_U322 , P3_R1200_U323 , P3_R1200_U324 , P3_R1200_U325 , P3_R1200_U326;
wire P3_R1200_U327 , P3_R1200_U328 , P3_R1200_U329 , P3_R1200_U330 , P3_R1200_U331 , P3_R1200_U332 , P3_R1200_U333 , P3_R1200_U334 , P3_R1200_U335 , P3_R1200_U336;
wire P3_R1200_U337 , P3_R1200_U338 , P3_R1200_U339 , P3_R1200_U340 , P3_R1200_U341 , P3_R1200_U342 , P3_R1200_U343 , P3_R1200_U344 , P3_R1200_U345 , P3_R1200_U346;
wire P3_R1200_U347 , P3_R1200_U348 , P3_R1200_U349 , P3_R1200_U350 , P3_R1200_U351 , P3_R1200_U352 , P3_R1200_U353 , P3_R1200_U354 , P3_R1200_U355 , P3_R1200_U356;
wire P3_R1200_U357 , P3_R1200_U358 , P3_R1200_U359 , P3_R1200_U360 , P3_R1200_U361 , P3_R1200_U362 , P3_R1200_U363 , P3_R1200_U364 , P3_R1200_U365 , P3_R1200_U366;
wire P3_R1200_U367 , P3_R1200_U368 , P3_R1200_U369 , P3_R1200_U370 , P3_R1200_U371 , P3_R1200_U372 , P3_R1200_U373 , P3_R1200_U374 , P3_R1200_U375 , P3_R1200_U376;
wire P3_R1200_U377 , P3_R1200_U378 , P3_R1200_U379 , P3_R1200_U380 , P3_R1200_U381 , P3_R1200_U382 , P3_R1200_U383 , P3_R1200_U384 , P3_R1200_U385 , P3_R1200_U386;
wire P3_R1200_U387 , P3_R1200_U388 , P3_R1200_U389 , P3_R1200_U390 , P3_R1200_U391 , P3_R1200_U392 , P3_R1200_U393 , P3_R1200_U394 , P3_R1200_U395 , P3_R1200_U396;
wire P3_R1200_U397 , P3_R1200_U398 , P3_R1200_U399 , P3_R1200_U400 , P3_R1200_U401 , P3_R1200_U402 , P3_R1200_U403 , P3_R1200_U404 , P3_R1200_U405 , P3_R1200_U406;
wire P3_R1200_U407 , P3_R1200_U408 , P3_R1200_U409 , P3_R1200_U410 , P3_R1200_U411 , P3_R1200_U412 , P3_R1200_U413 , P3_R1200_U414 , P3_R1200_U415 , P3_R1200_U416;
wire P3_R1200_U417 , P3_R1200_U418 , P3_R1200_U419 , P3_R1200_U420 , P3_R1200_U421 , P3_R1200_U422 , P3_R1200_U423 , P3_R1200_U424 , P3_R1200_U425 , P3_R1200_U426;
wire P3_R1200_U427 , P3_R1200_U428 , P3_R1200_U429 , P3_R1200_U430 , P3_R1200_U431 , P3_R1200_U432 , P3_R1200_U433 , P3_R1200_U434 , P3_R1200_U435 , P3_R1200_U436;
wire P3_R1200_U437 , P3_R1200_U438 , P3_R1200_U439 , P3_R1200_U440 , P3_R1200_U441 , P3_R1200_U442 , P3_R1200_U443 , P3_R1200_U444 , P3_R1200_U445 , P3_R1200_U446;
wire P3_R1200_U447 , P3_R1200_U448 , P3_R1200_U449 , P3_R1200_U450 , P3_R1200_U451 , P3_R1200_U452 , P3_R1200_U453 , P3_R1200_U454 , P3_R1200_U455 , P3_R1200_U456;
wire P3_R1200_U457 , P3_R1200_U458 , P3_R1200_U459 , P3_R1200_U460 , P3_R1200_U461 , P3_R1200_U462 , P3_R1200_U463 , P3_R1200_U464 , P3_R1200_U465 , P3_R1200_U466;
wire P3_R1200_U467 , P3_R1200_U468 , P3_R1200_U469 , P3_R1200_U470 , P3_R1200_U471 , P3_R1200_U472 , P3_R1200_U473 , P3_R1200_U474 , P3_R1200_U475 , P3_R1200_U476;
wire P3_R1200_U477 , P3_R1200_U478 , P3_R1200_U479 , P3_R1200_U480 , P3_R1200_U481 , P3_R1200_U482 , P3_R1200_U483 , P3_R1200_U484 , P3_R1200_U485 , P3_R1179_U6;
wire P3_R1179_U7 , P3_R1179_U8 , P3_R1179_U9 , P3_R1179_U10 , P3_R1179_U11 , P3_R1179_U12 , P3_R1179_U13 , P3_R1179_U14 , P3_R1179_U15 , P3_R1179_U16;
wire P3_R1179_U17 , P3_R1179_U18 , P3_R1179_U19 , P3_R1179_U20 , P3_R1179_U21 , P3_R1179_U22 , P3_R1179_U23 , P3_R1179_U24 , P3_R1179_U25 , P3_R1179_U26;
wire P3_R1179_U27 , P3_R1179_U28 , P3_R1179_U29 , P3_R1179_U30 , P3_R1179_U31 , P3_R1179_U32 , P3_R1179_U33 , P3_R1179_U34 , P3_R1179_U35 , P3_R1179_U36;
wire P3_R1179_U37 , P3_R1179_U38 , P3_R1179_U39 , P3_R1179_U40 , P3_R1179_U41 , P3_R1179_U42 , P3_R1179_U43 , P3_R1179_U44 , P3_R1179_U45 , P3_R1179_U46;
wire P3_R1179_U47 , P3_R1179_U48 , P3_R1179_U49 , P3_R1179_U50 , P3_R1179_U51 , P3_R1179_U52 , P3_R1179_U53 , P3_R1179_U54 , P3_R1179_U55 , P3_R1179_U56;
wire P3_R1179_U57 , P3_R1179_U58 , P3_R1179_U59 , P3_R1179_U60 , P3_R1179_U61 , P3_R1179_U62 , P3_R1179_U63 , P3_R1179_U64 , P3_R1179_U65 , P3_R1179_U66;
wire P3_R1179_U67 , P3_R1179_U68 , P3_R1179_U69 , P3_R1179_U70 , P3_R1179_U71 , P3_R1179_U72 , P3_R1179_U73 , P3_R1179_U74 , P3_R1179_U75 , P3_R1179_U76;
wire P3_R1179_U77 , P3_R1179_U78 , P3_R1179_U79 , P3_R1179_U80 , P3_R1179_U81 , P3_R1179_U82 , P3_R1179_U83 , P3_R1179_U84 , P3_R1179_U85 , P3_R1179_U86;
wire P3_R1179_U87 , P3_R1179_U88 , P3_R1179_U89 , P3_R1179_U90 , P3_R1179_U91 , P3_R1179_U92 , P3_R1179_U93 , P3_R1179_U94 , P3_R1179_U95 , P3_R1179_U96;
wire P3_R1179_U97 , P3_R1179_U98 , P3_R1179_U99 , P3_R1179_U100 , P3_R1179_U101 , P3_R1179_U102 , P3_R1179_U103 , P3_R1179_U104 , P3_R1179_U105 , P3_R1179_U106;
wire P3_R1179_U107 , P3_R1179_U108 , P3_R1179_U109 , P3_R1179_U110 , P3_R1179_U111 , P3_R1179_U112 , P3_R1179_U113 , P3_R1179_U114 , P3_R1179_U115 , P3_R1179_U116;
wire P3_R1179_U117 , P3_R1179_U118 , P3_R1179_U119 , P3_R1179_U120 , P3_R1179_U121 , P3_R1179_U122 , P3_R1179_U123 , P3_R1179_U124 , P3_R1179_U125 , P3_R1179_U126;
wire P3_R1179_U127 , P3_R1179_U128 , P3_R1179_U129 , P3_R1179_U130 , P3_R1179_U131 , P3_R1179_U132 , P3_R1179_U133 , P3_R1179_U134 , P3_R1179_U135 , P3_R1179_U136;
wire P3_R1179_U137 , P3_R1179_U138 , P3_R1179_U139 , P3_R1179_U140 , P3_R1179_U141 , P3_R1179_U142 , P3_R1179_U143 , P3_R1179_U144 , P3_R1179_U145 , P3_R1179_U146;
wire P3_R1179_U147 , P3_R1179_U148 , P3_R1179_U149 , P3_R1179_U150 , P3_R1179_U151 , P3_R1179_U152 , P3_R1179_U153 , P3_R1179_U154 , P3_R1179_U155 , P3_R1179_U156;
wire P3_R1179_U157 , P3_R1179_U158 , P3_R1179_U159 , P3_R1179_U160 , P3_R1179_U161 , P3_R1179_U162 , P3_R1179_U163 , P3_R1179_U164 , P3_R1179_U165 , P3_R1179_U166;
wire P3_R1179_U167 , P3_R1179_U168 , P3_R1179_U169 , P3_R1179_U170 , P3_R1179_U171 , P3_R1179_U172 , P3_R1179_U173 , P3_R1179_U174 , P3_R1179_U175 , P3_R1179_U176;
wire P3_R1179_U177 , P3_R1179_U178 , P3_R1179_U179 , P3_R1179_U180 , P3_R1179_U181 , P3_R1179_U182 , P3_R1179_U183 , P3_R1179_U184 , P3_R1179_U185 , P3_R1179_U186;
wire P3_R1179_U187 , P3_R1179_U188 , P3_R1179_U189 , P3_R1179_U190 , P3_R1179_U191 , P3_R1179_U192 , P3_R1179_U193 , P3_R1179_U194 , P3_R1179_U195 , P3_R1179_U196;
wire P3_R1179_U197 , P3_R1179_U198 , P3_R1179_U199 , P3_R1179_U200 , P3_R1179_U201 , P3_R1179_U202 , P3_R1179_U203 , P3_R1179_U204 , P3_R1179_U205 , P3_R1179_U206;
wire P3_R1179_U207 , P3_R1179_U208 , P3_R1179_U209 , P3_R1179_U210 , P3_R1179_U211 , P3_R1179_U212 , P3_R1179_U213 , P3_R1179_U214 , P3_R1179_U215 , P3_R1179_U216;
wire P3_R1179_U217 , P3_R1179_U218 , P3_R1179_U219 , P3_R1179_U220 , P3_R1179_U221 , P3_R1179_U222 , P3_R1179_U223 , P3_R1179_U224 , P3_R1179_U225 , P3_R1179_U226;
wire P3_R1179_U227 , P3_R1179_U228 , P3_R1179_U229 , P3_R1179_U230 , P3_R1179_U231 , P3_R1179_U232 , P3_R1179_U233 , P3_R1179_U234 , P3_R1179_U235 , P3_R1179_U236;
wire P3_R1179_U237 , P3_R1179_U238 , P3_R1179_U239 , P3_R1179_U240 , P3_R1179_U241 , P3_R1179_U242 , P3_R1179_U243 , P3_R1179_U244 , P3_R1179_U245 , P3_R1179_U246;
wire P3_R1179_U247 , P3_R1179_U248 , P3_R1179_U249 , P3_R1179_U250 , P3_R1179_U251 , P3_R1179_U252 , P3_R1179_U253 , P3_R1179_U254 , P3_R1179_U255 , P3_R1179_U256;
wire P3_R1179_U257 , P3_R1179_U258 , P3_R1179_U259 , P3_R1179_U260 , P3_R1179_U261 , P3_R1179_U262 , P3_R1179_U263 , P3_R1179_U264 , P3_R1179_U265 , P3_R1179_U266;
wire P3_R1179_U267 , P3_R1179_U268 , P3_R1179_U269 , P3_R1179_U270 , P3_R1179_U271 , P3_R1179_U272 , P3_R1179_U273 , P3_R1179_U274 , P3_R1179_U275 , P3_R1179_U276;
wire P3_R1179_U277 , P3_R1179_U278 , P3_R1179_U279 , P3_R1179_U280 , P3_R1179_U281 , P3_R1179_U282 , P3_R1179_U283 , P3_R1179_U284 , P3_R1179_U285 , P3_R1179_U286;
wire P3_R1179_U287 , P3_R1179_U288 , P3_R1179_U289 , P3_R1179_U290 , P3_R1179_U291 , P3_R1179_U292 , P3_R1179_U293 , P3_R1179_U294 , P3_R1179_U295 , P3_R1179_U296;
wire P3_R1179_U297 , P3_R1179_U298 , P3_R1179_U299 , P3_R1179_U300 , P3_R1179_U301 , P3_R1179_U302 , P3_R1179_U303 , P3_R1179_U304 , P3_R1179_U305 , P3_R1179_U306;
wire P3_R1179_U307 , P3_R1179_U308 , P3_R1179_U309 , P3_R1179_U310 , P3_R1179_U311 , P3_R1179_U312 , P3_R1179_U313 , P3_R1179_U314 , P3_R1179_U315 , P3_R1179_U316;
wire P3_R1179_U317 , P3_R1179_U318 , P3_R1179_U319 , P3_R1179_U320 , P3_R1179_U321 , P3_R1179_U322 , P3_R1179_U323 , P3_R1179_U324 , P3_R1179_U325 , P3_R1179_U326;
wire P3_R1179_U327 , P3_R1179_U328 , P3_R1179_U329 , P3_R1179_U330 , P3_R1179_U331 , P3_R1179_U332 , P3_R1179_U333 , P3_R1179_U334 , P3_R1179_U335 , P3_R1179_U336;
wire P3_R1179_U337 , P3_R1179_U338 , P3_R1179_U339 , P3_R1179_U340 , P3_R1179_U341 , P3_R1179_U342 , P3_R1179_U343 , P3_R1179_U344 , P3_R1179_U345 , P3_R1179_U346;
wire P3_R1179_U347 , P3_R1179_U348 , P3_R1179_U349 , P3_R1179_U350 , P3_R1179_U351 , P3_R1179_U352 , P3_R1179_U353 , P3_R1179_U354 , P3_R1179_U355 , P3_R1179_U356;
wire P3_R1179_U357 , P3_R1179_U358 , P3_R1179_U359 , P3_R1179_U360 , P3_R1179_U361 , P3_R1179_U362 , P3_R1179_U363 , P3_R1179_U364 , P3_R1179_U365 , P3_R1179_U366;
wire P3_R1179_U367 , P3_R1179_U368 , P3_R1179_U369 , P3_R1179_U370 , P3_R1179_U371 , P3_R1179_U372 , P3_R1179_U373 , P3_R1179_U374 , P3_R1179_U375 , P3_R1179_U376;
wire P3_R1179_U377 , P3_R1179_U378 , P3_R1179_U379 , P3_R1179_U380 , P3_R1179_U381 , P3_R1179_U382 , P3_R1179_U383 , P3_R1179_U384 , P3_R1179_U385 , P3_R1179_U386;
wire P3_R1179_U387 , P3_R1179_U388 , P3_R1179_U389 , P3_R1179_U390 , P3_R1179_U391 , P3_R1179_U392 , P3_R1179_U393 , P3_R1179_U394 , P3_R1179_U395 , P3_R1179_U396;
wire P3_R1179_U397 , P3_R1179_U398 , P3_R1179_U399 , P3_R1179_U400 , P3_R1179_U401 , P3_R1179_U402 , P3_R1179_U403 , P3_R1179_U404 , P3_R1179_U405 , P3_R1179_U406;
wire P3_R1179_U407 , P3_R1179_U408 , P3_R1179_U409 , P3_R1179_U410 , P3_R1179_U411 , P3_R1179_U412 , P3_R1179_U413 , P3_R1179_U414 , P3_R1179_U415 , P3_R1179_U416;
wire P3_R1179_U417 , P3_R1179_U418 , P3_R1179_U419 , P3_R1179_U420 , P3_R1179_U421 , P3_R1179_U422 , P3_R1179_U423 , P3_R1179_U424 , P3_R1179_U425 , P3_R1179_U426;
wire P3_R1179_U427 , P3_R1179_U428 , P3_R1179_U429 , P3_R1179_U430 , P3_R1179_U431 , P3_R1179_U432 , P3_R1179_U433 , P3_R1179_U434 , P3_R1179_U435 , P3_R1179_U436;
wire P3_R1179_U437 , P3_R1179_U438 , P3_R1179_U439 , P3_R1179_U440 , P3_R1179_U441 , P3_R1179_U442 , P3_R1179_U443 , P3_R1179_U444 , P3_R1179_U445 , P3_R1179_U446;
wire P3_R1179_U447 , P3_R1179_U448 , P3_R1179_U449 , P3_R1179_U450 , P3_R1179_U451 , P3_R1179_U452 , P3_R1179_U453 , P3_R1179_U454 , P3_R1179_U455 , P3_R1179_U456;
wire P3_R1179_U457 , P3_R1179_U458 , P3_R1179_U459 , P3_R1179_U460 , P3_R1179_U461 , P3_R1179_U462 , P3_R1179_U463 , P3_R1179_U464 , P3_R1179_U465 , P3_R1179_U466;
wire P3_R1179_U467 , P3_R1179_U468 , P3_R1179_U469 , P3_R1179_U470 , P3_R1179_U471 , P3_R1179_U472 , P3_R1179_U473 , P3_R1179_U474 , P3_R1179_U475 , P3_R1179_U476;
wire P3_R1179_U477 , P3_R1179_U478 , P3_R1179_U479 , P3_R1179_U480 , P3_R1179_U481 , P3_R1179_U482 , P3_R1179_U483 , P3_R1179_U484 , P3_R1179_U485 , P3_R1269_U6;
wire P3_R1269_U7 , P3_R1269_U8 , P3_R1269_U9 , P3_R1269_U10 , P3_R1269_U11 , P3_R1269_U12 , P3_R1269_U13 , P3_R1269_U14 , P3_R1269_U15 , P3_R1269_U16;
wire P3_R1269_U17 , P3_R1269_U18 , P3_R1269_U19 , P3_R1269_U20 , P3_R1269_U21 , P3_R1269_U22 , P3_R1269_U23 , P3_R1269_U24 , P3_R1269_U25 , P3_R1269_U26;
wire P3_R1269_U27 , P3_R1269_U28 , P3_R1269_U29 , P3_R1269_U30 , P3_R1269_U31 , P3_R1269_U32 , P3_R1269_U33 , P3_R1269_U34 , P3_R1269_U35 , P3_R1269_U36;
wire P3_R1269_U37 , P3_R1269_U38 , P3_R1269_U39 , P3_R1269_U40 , P3_R1269_U41 , P3_R1269_U42 , P3_R1269_U43 , P3_R1269_U44 , P3_R1269_U45 , P3_R1269_U46;
wire P3_R1269_U47 , P3_R1269_U48 , P3_R1269_U49 , P3_R1269_U50 , P3_R1269_U51 , P3_R1269_U52 , P3_R1269_U53 , P3_R1269_U54 , P3_R1269_U55 , P3_R1269_U56;
wire P3_R1269_U57 , P3_R1269_U58 , P3_R1269_U59 , P3_R1269_U60 , P3_R1269_U61 , P3_R1269_U62 , P3_R1269_U63 , P3_R1269_U64 , P3_R1269_U65 , P3_R1269_U66;
wire P3_R1269_U67 , P3_R1269_U68 , P3_R1269_U69 , P3_R1269_U70 , P3_R1269_U71 , P3_R1269_U72 , P3_R1269_U73 , P3_R1269_U74 , P3_R1269_U75 , P3_R1269_U76;
wire P3_R1269_U77 , P3_R1269_U78 , P3_R1269_U79 , P3_R1269_U80 , P3_R1269_U81 , P3_R1269_U82 , P3_R1269_U83 , P3_R1269_U84 , P3_R1269_U85 , P3_R1269_U86;
wire P3_R1269_U87 , P3_R1269_U88 , P3_R1269_U89 , P3_R1269_U90 , P3_R1269_U91 , P3_R1269_U92 , P3_R1269_U93 , P3_R1269_U94 , P3_R1269_U95 , P3_R1269_U96;
wire P3_R1269_U97 , P3_R1269_U98 , P3_R1269_U99 , P3_R1269_U100 , P3_R1269_U101 , P3_R1269_U102 , P3_R1269_U103 , P3_R1269_U104 , P3_R1269_U105 , P3_R1269_U106;
wire P3_R1269_U107 , P3_R1269_U108 , P3_R1269_U109 , P3_R1269_U110 , P3_R1269_U111 , P3_R1269_U112 , P3_R1269_U113 , P3_R1269_U114 , P3_R1269_U115 , P3_R1269_U116;
wire P3_R1269_U117 , P3_R1269_U118 , P3_R1269_U119 , P3_R1269_U120 , P3_R1269_U121 , P3_R1269_U122 , P3_R1269_U123 , P3_R1269_U124 , P3_R1269_U125 , P3_R1269_U126;
wire P3_R1269_U127 , P3_R1269_U128 , P3_R1269_U129 , P3_R1269_U130 , P3_R1269_U131 , P3_R1269_U132 , P3_R1269_U133 , P3_R1269_U134 , P3_R1269_U135 , P3_R1269_U136;
wire P3_R1269_U137 , P3_R1269_U138 , P3_R1269_U139 , P3_R1269_U140 , P3_R1269_U141 , P3_R1269_U142 , P3_R1269_U143 , P3_R1269_U144 , P3_R1269_U145 , P3_R1269_U146;
wire P3_R1269_U147 , P3_R1269_U148 , P3_R1269_U149 , P3_R1269_U150 , P3_R1269_U151 , P3_R1269_U152 , P3_R1269_U153 , P3_R1269_U154 , P3_R1269_U155 , P3_R1269_U156;
wire P3_R1269_U157 , P3_R1269_U158 , P3_R1269_U159 , P3_R1269_U160 , P3_R1269_U161 , P3_R1269_U162 , P3_R1269_U163 , P3_R1269_U164 , P3_R1269_U165 , P3_R1269_U166;
wire P3_R1269_U167 , P3_R1269_U168 , P3_R1269_U169 , P3_R1269_U170 , P3_R1269_U171 , P3_R1269_U172 , P3_R1269_U173 , P3_R1269_U174 , P3_R1269_U175 , P3_R1269_U176;
wire P3_R1269_U177 , P3_R1269_U178 , P3_R1269_U179 , P3_R1269_U180 , P3_R1269_U181 , P3_R1269_U182 , P3_R1269_U183 , P3_R1269_U184 , P3_R1269_U185 , P3_R1269_U186;
wire P3_R1269_U187 , P3_R1269_U188 , P3_R1269_U189 , P3_R1269_U190 , P3_R1269_U191 , P3_R1269_U192 , P3_R1269_U193 , P3_R1269_U194 , P3_R1269_U195 , P3_R1269_U196;
wire P3_R1269_U197 , P3_R1269_U198 , P3_R1269_U199 , P3_R1269_U200 , P3_R1269_U201 , P3_R1269_U202 , P3_R1110_U4 , P3_R1110_U5 , P3_R1110_U6 , P3_R1110_U7;
wire P3_R1110_U8 , P3_R1110_U9 , P3_R1110_U10 , P3_R1110_U11 , P3_R1110_U12 , P3_R1110_U13 , P3_R1110_U14 , P3_R1110_U15 , P3_R1110_U16 , P3_R1110_U17;
wire P3_R1110_U18 , P3_R1110_U19 , P3_R1110_U20 , P3_R1110_U21 , P3_R1110_U22 , P3_R1110_U23 , P3_R1110_U24 , P3_R1110_U25 , P3_R1110_U26 , P3_R1110_U27;
wire P3_R1110_U28 , P3_R1110_U29 , P3_R1110_U30 , P3_R1110_U31 , P3_R1110_U32 , P3_R1110_U33 , P3_R1110_U34 , P3_R1110_U35 , P3_R1110_U36 , P3_R1110_U37;
wire P3_R1110_U38 , P3_R1110_U39 , P3_R1110_U40 , P3_R1110_U41 , P3_R1110_U42 , P3_R1110_U43 , P3_R1110_U44 , P3_R1110_U45 , P3_R1110_U46 , P3_R1110_U47;
wire P3_R1110_U48 , P3_R1110_U49 , P3_R1110_U50 , P3_R1110_U51 , P3_R1110_U52 , P3_R1110_U53 , P3_R1110_U54 , P3_R1110_U55 , P3_R1110_U56 , P3_R1110_U57;
wire P3_R1110_U58 , P3_R1110_U59 , P3_R1110_U60 , P3_R1110_U61 , P3_R1110_U62 , P3_R1110_U63 , P3_R1110_U64 , P3_R1110_U65 , P3_R1110_U66 , P3_R1110_U67;
wire P3_R1110_U68 , P3_R1110_U69 , P3_R1110_U70 , P3_R1110_U71 , P3_R1110_U72 , P3_R1110_U73 , P3_R1110_U74 , P3_R1110_U75 , P3_R1110_U76 , P3_R1110_U77;
wire P3_R1110_U78 , P3_R1110_U79 , P3_R1110_U80 , P3_R1110_U81 , P3_R1110_U82 , P3_R1110_U83 , P3_R1110_U84 , P3_R1110_U85 , P3_R1110_U86 , P3_R1110_U87;
wire P3_R1110_U88 , P3_R1110_U89 , P3_R1110_U90 , P3_R1110_U91 , P3_R1110_U92 , P3_R1110_U93 , P3_R1110_U94 , P3_R1110_U95 , P3_R1110_U96 , P3_R1110_U97;
wire P3_R1110_U98 , P3_R1110_U99 , P3_R1110_U100 , P3_R1110_U101 , P3_R1110_U102 , P3_R1110_U103 , P3_R1110_U104 , P3_R1110_U105 , P3_R1110_U106 , P3_R1110_U107;
wire P3_R1110_U108 , P3_R1110_U109 , P3_R1110_U110 , P3_R1110_U111 , P3_R1110_U112 , P3_R1110_U113 , P3_R1110_U114 , P3_R1110_U115 , P3_R1110_U116 , P3_R1110_U117;
wire P3_R1110_U118 , P3_R1110_U119 , P3_R1110_U120 , P3_R1110_U121 , P3_R1110_U122 , P3_R1110_U123 , P3_R1110_U124 , P3_R1110_U125 , P3_R1110_U126 , P3_R1110_U127;
wire P3_R1110_U128 , P3_R1110_U129 , P3_R1110_U130 , P3_R1110_U131 , P3_R1110_U132 , P3_R1110_U133 , P3_R1110_U134 , P3_R1110_U135 , P3_R1110_U136 , P3_R1110_U137;
wire P3_R1110_U138 , P3_R1110_U139 , P3_R1110_U140 , P3_R1110_U141 , P3_R1110_U142 , P3_R1110_U143 , P3_R1110_U144 , P3_R1110_U145 , P3_R1110_U146 , P3_R1110_U147;
wire P3_R1110_U148 , P3_R1110_U149 , P3_R1110_U150 , P3_R1110_U151 , P3_R1110_U152 , P3_R1110_U153 , P3_R1110_U154 , P3_R1110_U155 , P3_R1110_U156 , P3_R1110_U157;
wire P3_R1110_U158 , P3_R1110_U159 , P3_R1110_U160 , P3_R1110_U161 , P3_R1110_U162 , P3_R1110_U163 , P3_R1110_U164 , P3_R1110_U165 , P3_R1110_U166 , P3_R1110_U167;
wire P3_R1110_U168 , P3_R1110_U169 , P3_R1110_U170 , P3_R1110_U171 , P3_R1110_U172 , P3_R1110_U173 , P3_R1110_U174 , P3_R1110_U175 , P3_R1110_U176 , P3_R1110_U177;
wire P3_R1110_U178 , P3_R1110_U179 , P3_R1110_U180 , P3_R1110_U181 , P3_R1110_U182 , P3_R1110_U183 , P3_R1110_U184 , P3_R1110_U185 , P3_R1110_U186 , P3_R1110_U187;
wire P3_R1110_U188 , P3_R1110_U189 , P3_R1110_U190 , P3_R1110_U191 , P3_R1110_U192 , P3_R1110_U193 , P3_R1110_U194 , P3_R1110_U195 , P3_R1110_U196 , P3_R1110_U197;
wire P3_R1110_U198 , P3_R1110_U199 , P3_R1110_U200 , P3_R1110_U201 , P3_R1110_U202 , P3_R1110_U203 , P3_R1110_U204 , P3_R1110_U205 , P3_R1110_U206 , P3_R1110_U207;
wire P3_R1110_U208 , P3_R1110_U209 , P3_R1110_U210 , P3_R1110_U211 , P3_R1110_U212 , P3_R1110_U213 , P3_R1110_U214 , P3_R1110_U215 , P3_R1110_U216 , P3_R1110_U217;
wire P3_R1110_U218 , P3_R1110_U219 , P3_R1110_U220 , P3_R1110_U221 , P3_R1110_U222 , P3_R1110_U223 , P3_R1110_U224 , P3_R1110_U225 , P3_R1110_U226 , P3_R1110_U227;
wire P3_R1110_U228 , P3_R1110_U229 , P3_R1110_U230 , P3_R1110_U231 , P3_R1110_U232 , P3_R1110_U233 , P3_R1110_U234 , P3_R1110_U235 , P3_R1110_U236 , P3_R1110_U237;
wire P3_R1110_U238 , P3_R1110_U239 , P3_R1110_U240 , P3_R1110_U241 , P3_R1110_U242 , P3_R1110_U243 , P3_R1110_U244 , P3_R1110_U245 , P3_R1110_U246 , P3_R1110_U247;
wire P3_R1110_U248 , P3_R1110_U249 , P3_R1110_U250 , P3_R1110_U251 , P3_R1110_U252 , P3_R1110_U253 , P3_R1110_U254 , P3_R1110_U255 , P3_R1110_U256 , P3_R1110_U257;
wire P3_R1110_U258 , P3_R1110_U259 , P3_R1110_U260 , P3_R1110_U261 , P3_R1110_U262 , P3_R1110_U263 , P3_R1110_U264 , P3_R1110_U265 , P3_R1110_U266 , P3_R1110_U267;
wire P3_R1110_U268 , P3_R1110_U269 , P3_R1110_U270 , P3_R1110_U271 , P3_R1110_U272 , P3_R1110_U273 , P3_R1110_U274 , P3_R1110_U275 , P3_R1110_U276 , P3_R1110_U277;
wire P3_R1110_U278 , P3_R1110_U279 , P3_R1110_U280 , P3_R1110_U281 , P3_R1110_U282 , P3_R1110_U283 , P3_R1110_U284 , P3_R1110_U285 , P3_R1110_U286 , P3_R1110_U287;
wire P3_R1110_U288 , P3_R1110_U289 , P3_R1110_U290 , P3_R1110_U291 , P3_R1110_U292 , P3_R1110_U293 , P3_R1110_U294 , P3_R1110_U295 , P3_R1110_U296 , P3_R1110_U297;
wire P3_R1110_U298 , P3_R1110_U299 , P3_R1110_U300 , P3_R1110_U301 , P3_R1110_U302 , P3_R1110_U303 , P3_R1110_U304 , P3_R1110_U305 , P3_R1110_U306 , P3_R1110_U307;
wire P3_R1110_U308 , P3_R1110_U309 , P3_R1110_U310 , P3_R1110_U311 , P3_R1110_U312 , P3_R1110_U313 , P3_R1110_U314 , P3_R1110_U315 , P3_R1110_U316 , P3_R1110_U317;
wire P3_R1110_U318 , P3_R1110_U319 , P3_R1110_U320 , P3_R1110_U321 , P3_R1110_U322 , P3_R1110_U323 , P3_R1110_U324 , P3_R1110_U325 , P3_R1110_U326 , P3_R1110_U327;
wire P3_R1110_U328 , P3_R1110_U329 , P3_R1110_U330 , P3_R1110_U331 , P3_R1110_U332 , P3_R1110_U333 , P3_R1110_U334 , P3_R1110_U335 , P3_R1110_U336 , P3_R1110_U337;
wire P3_R1110_U338 , P3_R1110_U339 , P3_R1110_U340 , P3_R1110_U341 , P3_R1110_U342 , P3_R1110_U343 , P3_R1110_U344 , P3_R1110_U345 , P3_R1110_U346 , P3_R1110_U347;
wire P3_R1110_U348 , P3_R1110_U349 , P3_R1110_U350 , P3_R1110_U351 , P3_R1110_U352 , P3_R1110_U353 , P3_R1110_U354 , P3_R1110_U355 , P3_R1110_U356 , P3_R1110_U357;
wire P3_R1110_U358 , P3_R1110_U359 , P3_R1110_U360 , P3_R1110_U361 , P3_R1110_U362 , P3_R1110_U363 , P3_R1110_U364 , P3_R1110_U365 , P3_R1110_U366 , P3_R1110_U367;
wire P3_R1110_U368 , P3_R1110_U369 , P3_R1110_U370 , P3_R1110_U371 , P3_R1110_U372 , P3_R1110_U373 , P3_R1110_U374 , P3_R1110_U375 , P3_R1110_U376 , P3_R1110_U377;
wire P3_R1110_U378 , P3_R1110_U379 , P3_R1110_U380 , P3_R1110_U381 , P3_R1110_U382 , P3_R1110_U383 , P3_R1110_U384 , P3_R1110_U385 , P3_R1110_U386 , P3_R1110_U387;
wire P3_R1110_U388 , P3_R1110_U389 , P3_R1110_U390 , P3_R1110_U391 , P3_R1110_U392 , P3_R1110_U393 , P3_R1110_U394 , P3_R1110_U395 , P3_R1110_U396 , P3_R1110_U397;
wire P3_R1110_U398 , P3_R1110_U399 , P3_R1110_U400 , P3_R1110_U401 , P3_R1110_U402 , P3_R1110_U403 , P3_R1110_U404 , P3_R1110_U405 , P3_R1110_U406 , P3_R1110_U407;
wire P3_R1110_U408 , P3_R1110_U409 , P3_R1110_U410 , P3_R1110_U411 , P3_R1110_U412 , P3_R1110_U413 , P3_R1110_U414 , P3_R1110_U415 , P3_R1110_U416 , P3_R1110_U417;
wire P3_R1110_U418 , P3_R1110_U419 , P3_R1110_U420 , P3_R1110_U421 , P3_R1110_U422 , P3_R1110_U423 , P3_R1110_U424 , P3_R1110_U425 , P3_R1110_U426 , P3_R1110_U427;
wire P3_R1110_U428 , P3_R1110_U429 , P3_R1110_U430 , P3_R1110_U431 , P3_R1110_U432 , P3_R1110_U433 , P3_R1110_U434 , P3_R1110_U435 , P3_R1110_U436 , P3_R1110_U437;
wire P3_R1110_U438 , P3_R1110_U439 , P3_R1110_U440 , P3_R1110_U441 , P3_R1110_U442 , P3_R1110_U443 , P3_R1110_U444 , P3_R1110_U445 , P3_R1110_U446 , P3_R1110_U447;
wire P3_R1110_U448 , P3_R1110_U449 , P3_R1110_U450 , P3_R1110_U451 , P3_R1110_U452 , P3_R1110_U453 , P3_R1110_U454 , P3_R1110_U455 , P3_R1110_U456 , P3_R1110_U457;
wire P3_R1110_U458 , P3_R1110_U459 , P3_R1110_U460 , P3_R1110_U461 , P3_R1110_U462 , P3_R1110_U463 , P3_R1110_U464 , P3_R1110_U465 , P3_R1110_U466 , P3_R1110_U467;
wire P3_R1110_U468 , P3_R1110_U469 , P3_R1110_U470 , P3_R1110_U471 , P3_R1110_U472 , P3_R1110_U473 , P3_R1110_U474 , P3_R1110_U475 , P3_R1110_U476 , P3_R1110_U477;
wire P3_R1110_U478 , P3_R1110_U479 , P3_R1110_U480 , P3_R1110_U481 , P3_R1110_U482 , P3_R1110_U483 , P3_R1110_U484 , P3_R1110_U485 , P3_R1110_U486 , P3_R1110_U487;
wire P3_R1110_U488 , P3_R1110_U489 , P3_R1110_U490 , P3_R1110_U491 , P3_R1110_U492 , P3_R1110_U493 , P3_R1110_U494 , P3_R1110_U495 , P3_R1110_U496 , P3_R1110_U497;
wire P3_R1110_U498 , P3_R1110_U499 , P3_R1110_U500 , P3_R1110_U501 , P3_R1110_U502 , P3_R1110_U503 , P3_R1110_U504 , P3_R1297_U6 , P3_R1297_U7 , P3_R1077_U4;
wire P3_R1077_U5 , P3_R1077_U6 , P3_R1077_U7 , P3_R1077_U8 , P3_R1077_U9 , P3_R1077_U10 , P3_R1077_U11 , P3_R1077_U12 , P3_R1077_U13 , P3_R1077_U14;
wire P3_R1077_U15 , P3_R1077_U16 , P3_R1077_U17 , P3_R1077_U18 , P3_R1077_U19 , P3_R1077_U20 , P3_R1077_U21 , P3_R1077_U22 , P3_R1077_U23 , P3_R1077_U24;
wire P3_R1077_U25 , P3_R1077_U26 , P3_R1077_U27 , P3_R1077_U28 , P3_R1077_U29 , P3_R1077_U30 , P3_R1077_U31 , P3_R1077_U32 , P3_R1077_U33 , P3_R1077_U34;
wire P3_R1077_U35 , P3_R1077_U36 , P3_R1077_U37 , P3_R1077_U38 , P3_R1077_U39 , P3_R1077_U40 , P3_R1077_U41 , P3_R1077_U42 , P3_R1077_U43 , P3_R1077_U44;
wire P3_R1077_U45 , P3_R1077_U46 , P3_R1077_U47 , P3_R1077_U48 , P3_R1077_U49 , P3_R1077_U50 , P3_R1077_U51 , P3_R1077_U52 , P3_R1077_U53 , P3_R1077_U54;
wire P3_R1077_U55 , P3_R1077_U56 , P3_R1077_U57 , P3_R1077_U58 , P3_R1077_U59 , P3_R1077_U60 , P3_R1077_U61 , P3_R1077_U62 , P3_R1077_U63 , P3_R1077_U64;
wire P3_R1077_U65 , P3_R1077_U66 , P3_R1077_U67 , P3_R1077_U68 , P3_R1077_U69 , P3_R1077_U70 , P3_R1077_U71 , P3_R1077_U72 , P3_R1077_U73 , P3_R1077_U74;
wire P3_R1077_U75 , P3_R1077_U76 , P3_R1077_U77 , P3_R1077_U78 , P3_R1077_U79 , P3_R1077_U80 , P3_R1077_U81 , P3_R1077_U82 , P3_R1077_U83 , P3_R1077_U84;
wire P3_R1077_U85 , P3_R1077_U86 , P3_R1077_U87 , P3_R1077_U88 , P3_R1077_U89 , P3_R1077_U90 , P3_R1077_U91 , P3_R1077_U92 , P3_R1077_U93 , P3_R1077_U94;
wire P3_R1077_U95 , P3_R1077_U96 , P3_R1077_U97 , P3_R1077_U98 , P3_R1077_U99 , P3_R1077_U100 , P3_R1077_U101 , P3_R1077_U102 , P3_R1077_U103 , P3_R1077_U104;
wire P3_R1077_U105 , P3_R1077_U106 , P3_R1077_U107 , P3_R1077_U108 , P3_R1077_U109 , P3_R1077_U110 , P3_R1077_U111 , P3_R1077_U112 , P3_R1077_U113 , P3_R1077_U114;
wire P3_R1077_U115 , P3_R1077_U116 , P3_R1077_U117 , P3_R1077_U118 , P3_R1077_U119 , P3_R1077_U120 , P3_R1077_U121 , P3_R1077_U122 , P3_R1077_U123 , P3_R1077_U124;
wire P3_R1077_U125 , P3_R1077_U126 , P3_R1077_U127 , P3_R1077_U128 , P3_R1077_U129 , P3_R1077_U130 , P3_R1077_U131 , P3_R1077_U132 , P3_R1077_U133 , P3_R1077_U134;
wire P3_R1077_U135 , P3_R1077_U136 , P3_R1077_U137 , P3_R1077_U138 , P3_R1077_U139 , P3_R1077_U140 , P3_R1077_U141 , P3_R1077_U142 , P3_R1077_U143 , P3_R1077_U144;
wire P3_R1077_U145 , P3_R1077_U146 , P3_R1077_U147 , P3_R1077_U148 , P3_R1077_U149 , P3_R1077_U150 , P3_R1077_U151 , P3_R1077_U152 , P3_R1077_U153 , P3_R1077_U154;
wire P3_R1077_U155 , P3_R1077_U156 , P3_R1077_U157 , P3_R1077_U158 , P3_R1077_U159 , P3_R1077_U160 , P3_R1077_U161 , P3_R1077_U162 , P3_R1077_U163 , P3_R1077_U164;
wire P3_R1077_U165 , P3_R1077_U166 , P3_R1077_U167 , P3_R1077_U168 , P3_R1077_U169 , P3_R1077_U170 , P3_R1077_U171 , P3_R1077_U172 , P3_R1077_U173 , P3_R1077_U174;
wire P3_R1077_U175 , P3_R1077_U176 , P3_R1077_U177 , P3_R1077_U178 , P3_R1077_U179 , P3_R1077_U180 , P3_R1077_U181 , P3_R1077_U182 , P3_R1077_U183 , P3_R1077_U184;
wire P3_R1077_U185 , P3_R1077_U186 , P3_R1077_U187 , P3_R1077_U188 , P3_R1077_U189 , P3_R1077_U190 , P3_R1077_U191 , P3_R1077_U192 , P3_R1077_U193 , P3_R1077_U194;
wire P3_R1077_U195 , P3_R1077_U196 , P3_R1077_U197 , P3_R1077_U198 , P3_R1077_U199 , P3_R1077_U200 , P3_R1077_U201 , P3_R1077_U202 , P3_R1077_U203 , P3_R1077_U204;
wire P3_R1077_U205 , P3_R1077_U206 , P3_R1077_U207 , P3_R1077_U208 , P3_R1077_U209 , P3_R1077_U210 , P3_R1077_U211 , P3_R1077_U212 , P3_R1077_U213 , P3_R1077_U214;
wire P3_R1077_U215 , P3_R1077_U216 , P3_R1077_U217 , P3_R1077_U218 , P3_R1077_U219 , P3_R1077_U220 , P3_R1077_U221 , P3_R1077_U222 , P3_R1077_U223 , P3_R1077_U224;
wire P3_R1077_U225 , P3_R1077_U226 , P3_R1077_U227 , P3_R1077_U228 , P3_R1077_U229 , P3_R1077_U230 , P3_R1077_U231 , P3_R1077_U232 , P3_R1077_U233 , P3_R1077_U234;
wire P3_R1077_U235 , P3_R1077_U236 , P3_R1077_U237 , P3_R1077_U238 , P3_R1077_U239 , P3_R1077_U240 , P3_R1077_U241 , P3_R1077_U242 , P3_R1077_U243 , P3_R1077_U244;
wire P3_R1077_U245 , P3_R1077_U246 , P3_R1077_U247 , P3_R1077_U248 , P3_R1077_U249 , P3_R1077_U250 , P3_R1077_U251 , P3_R1077_U252 , P3_R1077_U253 , P3_R1077_U254;
wire P3_R1077_U255 , P3_R1077_U256 , P3_R1077_U257 , P3_R1077_U258 , P3_R1077_U259 , P3_R1077_U260 , P3_R1077_U261 , P3_R1077_U262 , P3_R1077_U263 , P3_R1077_U264;
wire P3_R1077_U265 , P3_R1077_U266 , P3_R1077_U267 , P3_R1077_U268 , P3_R1077_U269 , P3_R1077_U270 , P3_R1077_U271 , P3_R1077_U272 , P3_R1077_U273 , P3_R1077_U274;
wire P3_R1077_U275 , P3_R1077_U276 , P3_R1077_U277 , P3_R1077_U278 , P3_R1077_U279 , P3_R1077_U280 , P3_R1077_U281 , P3_R1077_U282 , P3_R1077_U283 , P3_R1077_U284;
wire P3_R1077_U285 , P3_R1077_U286 , P3_R1077_U287 , P3_R1077_U288 , P3_R1077_U289 , P3_R1077_U290 , P3_R1077_U291 , P3_R1077_U292 , P3_R1077_U293 , P3_R1077_U294;
wire P3_R1077_U295 , P3_R1077_U296 , P3_R1077_U297 , P3_R1077_U298 , P3_R1077_U299 , P3_R1077_U300 , P3_R1077_U301 , P3_R1077_U302 , P3_R1077_U303 , P3_R1077_U304;
wire P3_R1077_U305 , P3_R1077_U306 , P3_R1077_U307 , P3_R1077_U308 , P3_R1077_U309 , P3_R1077_U310 , P3_R1077_U311 , P3_R1077_U312 , P3_R1077_U313 , P3_R1077_U314;
wire P3_R1077_U315 , P3_R1077_U316 , P3_R1077_U317 , P3_R1077_U318 , P3_R1077_U319 , P3_R1077_U320 , P3_R1077_U321 , P3_R1077_U322 , P3_R1077_U323 , P3_R1077_U324;
wire P3_R1077_U325 , P3_R1077_U326 , P3_R1077_U327 , P3_R1077_U328 , P3_R1077_U329 , P3_R1077_U330 , P3_R1077_U331 , P3_R1077_U332 , P3_R1077_U333 , P3_R1077_U334;
wire P3_R1077_U335 , P3_R1077_U336 , P3_R1077_U337 , P3_R1077_U338 , P3_R1077_U339 , P3_R1077_U340 , P3_R1077_U341 , P3_R1077_U342 , P3_R1077_U343 , P3_R1077_U344;
wire P3_R1077_U345 , P3_R1077_U346 , P3_R1077_U347 , P3_R1077_U348 , P3_R1077_U349 , P3_R1077_U350 , P3_R1077_U351 , P3_R1077_U352 , P3_R1077_U353 , P3_R1077_U354;
wire P3_R1077_U355 , P3_R1077_U356 , P3_R1077_U357 , P3_R1077_U358 , P3_R1077_U359 , P3_R1077_U360 , P3_R1077_U361 , P3_R1077_U362 , P3_R1077_U363 , P3_R1077_U364;
wire P3_R1077_U365 , P3_R1077_U366 , P3_R1077_U367 , P3_R1077_U368 , P3_R1077_U369 , P3_R1077_U370 , P3_R1077_U371 , P3_R1077_U372 , P3_R1077_U373 , P3_R1077_U374;
wire P3_R1077_U375 , P3_R1077_U376 , P3_R1077_U377 , P3_R1077_U378 , P3_R1077_U379 , P3_R1077_U380 , P3_R1077_U381 , P3_R1077_U382 , P3_R1077_U383 , P3_R1077_U384;
wire P3_R1077_U385 , P3_R1077_U386 , P3_R1077_U387 , P3_R1077_U388 , P3_R1077_U389 , P3_R1077_U390 , P3_R1077_U391 , P3_R1077_U392 , P3_R1077_U393 , P3_R1077_U394;
wire P3_R1077_U395 , P3_R1077_U396 , P3_R1077_U397 , P3_R1077_U398 , P3_R1077_U399 , P3_R1077_U400 , P3_R1077_U401 , P3_R1077_U402 , P3_R1077_U403 , P3_R1077_U404;
wire P3_R1077_U405 , P3_R1077_U406 , P3_R1077_U407 , P3_R1077_U408 , P3_R1077_U409 , P3_R1077_U410 , P3_R1077_U411 , P3_R1077_U412 , P3_R1077_U413 , P3_R1077_U414;
wire P3_R1077_U415 , P3_R1077_U416 , P3_R1077_U417 , P3_R1077_U418 , P3_R1077_U419 , P3_R1077_U420 , P3_R1077_U421 , P3_R1077_U422 , P3_R1077_U423 , P3_R1077_U424;
wire P3_R1077_U425 , P3_R1077_U426 , P3_R1077_U427 , P3_R1077_U428 , P3_R1077_U429 , P3_R1077_U430 , P3_R1077_U431 , P3_R1077_U432 , P3_R1077_U433 , P3_R1077_U434;
wire P3_R1077_U435 , P3_R1077_U436 , P3_R1077_U437 , P3_R1077_U438 , P3_R1077_U439 , P3_R1077_U440 , P3_R1077_U441 , P3_R1077_U442 , P3_R1077_U443 , P3_R1077_U444;
wire P3_R1077_U445 , P3_R1077_U446 , P3_R1077_U447 , P3_R1077_U448 , P3_R1077_U449 , P3_R1077_U450 , P3_R1077_U451 , P3_R1077_U452 , P3_R1077_U453 , P3_R1077_U454;
wire P3_R1077_U455 , P3_R1077_U456 , P3_R1077_U457 , P3_R1077_U458 , P3_R1077_U459 , P3_R1077_U460 , P3_R1077_U461 , P3_R1077_U462 , P3_R1077_U463 , P3_R1077_U464;
wire P3_R1077_U465 , P3_R1077_U466 , P3_R1077_U467 , P3_R1077_U468 , P3_R1077_U469 , P3_R1077_U470 , P3_R1077_U471 , P3_R1077_U472 , P3_R1077_U473 , P3_R1077_U474;
wire P3_R1077_U475 , P3_R1077_U476 , P3_R1077_U477 , P3_R1077_U478 , P3_R1077_U479 , P3_R1077_U480 , P3_R1077_U481 , P3_R1077_U482 , P3_R1077_U483 , P3_R1077_U484;
wire P3_R1077_U485 , P3_R1077_U486 , P3_R1077_U487 , P3_R1077_U488 , P3_R1077_U489 , P3_R1077_U490 , P3_R1077_U491 , P3_R1077_U492 , P3_R1077_U493 , P3_R1077_U494;
wire P3_R1077_U495 , P3_R1077_U496 , P3_R1077_U497 , P3_R1077_U498 , P3_R1077_U499 , P3_R1077_U500 , P3_R1077_U501 , P3_R1077_U502 , P3_R1077_U503 , P3_R1077_U504;
wire P3_R1143_U4 , P3_R1143_U5 , P3_R1143_U6 , P3_R1143_U7 , P3_R1143_U8 , P3_R1143_U9 , P3_R1143_U10 , P3_R1143_U11 , P3_R1143_U12 , P3_R1143_U13;
wire P3_R1143_U14 , P3_R1143_U15 , P3_R1143_U16 , P3_R1143_U17 , P3_R1143_U18 , P3_R1143_U19 , P3_R1143_U20 , P3_R1143_U21 , P3_R1143_U22 , P3_R1143_U23;
wire P3_R1143_U24 , P3_R1143_U25 , P3_R1143_U26 , P3_R1143_U27 , P3_R1143_U28 , P3_R1143_U29 , P3_R1143_U30 , P3_R1143_U31 , P3_R1143_U32 , P3_R1143_U33;
wire P3_R1143_U34 , P3_R1143_U35 , P3_R1143_U36 , P3_R1143_U37 , P3_R1143_U38 , P3_R1143_U39 , P3_R1143_U40 , P3_R1143_U41 , P3_R1143_U42 , P3_R1143_U43;
wire P3_R1143_U44 , P3_R1143_U45 , P3_R1143_U46 , P3_R1143_U47 , P3_R1143_U48 , P3_R1143_U49 , P3_R1143_U50 , P3_R1143_U51 , P3_R1143_U52 , P3_R1143_U53;
wire P3_R1143_U54 , P3_R1143_U55 , P3_R1143_U56 , P3_R1143_U57 , P3_R1143_U58 , P3_R1143_U59 , P3_R1143_U60 , P3_R1143_U61 , P3_R1143_U62 , P3_R1143_U63;
wire P3_R1143_U64 , P3_R1143_U65 , P3_R1143_U66 , P3_R1143_U67 , P3_R1143_U68 , P3_R1143_U69 , P3_R1143_U70 , P3_R1143_U71 , P3_R1143_U72 , P3_R1143_U73;
wire P3_R1143_U74 , P3_R1143_U75 , P3_R1143_U76 , P3_R1143_U77 , P3_R1143_U78 , P3_R1143_U79 , P3_R1143_U80 , P3_R1143_U81 , P3_R1143_U82 , P3_R1143_U83;
wire P3_R1143_U84 , P3_R1143_U85 , P3_R1143_U86 , P3_R1143_U87 , P3_R1143_U88 , P3_R1143_U89 , P3_R1143_U90 , P3_R1143_U91 , P3_R1143_U92 , P3_R1143_U93;
wire P3_R1143_U94 , P3_R1143_U95 , P3_R1143_U96 , P3_R1143_U97 , P3_R1143_U98 , P3_R1143_U99 , P3_R1143_U100 , P3_R1143_U101 , P3_R1143_U102 , P3_R1143_U103;
wire P3_R1143_U104 , P3_R1143_U105 , P3_R1143_U106 , P3_R1143_U107 , P3_R1143_U108 , P3_R1143_U109 , P3_R1143_U110 , P3_R1143_U111 , P3_R1143_U112 , P3_R1143_U113;
wire P3_R1143_U114 , P3_R1143_U115 , P3_R1143_U116 , P3_R1143_U117 , P3_R1143_U118 , P3_R1143_U119 , P3_R1143_U120 , P3_R1143_U121 , P3_R1143_U122 , P3_R1143_U123;
wire P3_R1143_U124 , P3_R1143_U125 , P3_R1143_U126 , P3_R1143_U127 , P3_R1143_U128 , P3_R1143_U129 , P3_R1143_U130 , P3_R1143_U131 , P3_R1143_U132 , P3_R1143_U133;
wire P3_R1143_U134 , P3_R1143_U135 , P3_R1143_U136 , P3_R1143_U137 , P3_R1143_U138 , P3_R1143_U139 , P3_R1143_U140 , P3_R1143_U141 , P3_R1143_U142 , P3_R1143_U143;
wire P3_R1143_U144 , P3_R1143_U145 , P3_R1143_U146 , P3_R1143_U147 , P3_R1143_U148 , P3_R1143_U149 , P3_R1143_U150 , P3_R1143_U151 , P3_R1143_U152 , P3_R1143_U153;
wire P3_R1143_U154 , P3_R1143_U155 , P3_R1143_U156 , P3_R1143_U157 , P3_R1143_U158 , P3_R1143_U159 , P3_R1143_U160 , P3_R1143_U161 , P3_R1143_U162 , P3_R1143_U163;
wire P3_R1143_U164 , P3_R1143_U165 , P3_R1143_U166 , P3_R1143_U167 , P3_R1143_U168 , P3_R1143_U169 , P3_R1143_U170 , P3_R1143_U171 , P3_R1143_U172 , P3_R1143_U173;
wire P3_R1143_U174 , P3_R1143_U175 , P3_R1143_U176 , P3_R1143_U177 , P3_R1143_U178 , P3_R1143_U179 , P3_R1143_U180 , P3_R1143_U181 , P3_R1143_U182 , P3_R1143_U183;
wire P3_R1143_U184 , P3_R1143_U185 , P3_R1143_U186 , P3_R1143_U187 , P3_R1143_U188 , P3_R1143_U189 , P3_R1143_U190 , P3_R1143_U191 , P3_R1143_U192 , P3_R1143_U193;
wire P3_R1143_U194 , P3_R1143_U195 , P3_R1143_U196 , P3_R1143_U197 , P3_R1143_U198 , P3_R1143_U199 , P3_R1143_U200 , P3_R1143_U201 , P3_R1143_U202 , P3_R1143_U203;
wire P3_R1143_U204 , P3_R1143_U205 , P3_R1143_U206 , P3_R1143_U207 , P3_R1143_U208 , P3_R1143_U209 , P3_R1143_U210 , P3_R1143_U211 , P3_R1143_U212 , P3_R1143_U213;
wire P3_R1143_U214 , P3_R1143_U215 , P3_R1143_U216 , P3_R1143_U217 , P3_R1143_U218 , P3_R1143_U219 , P3_R1143_U220 , P3_R1143_U221 , P3_R1143_U222 , P3_R1143_U223;
wire P3_R1143_U224 , P3_R1143_U225 , P3_R1143_U226 , P3_R1143_U227 , P3_R1143_U228 , P3_R1143_U229 , P3_R1143_U230 , P3_R1143_U231 , P3_R1143_U232 , P3_R1143_U233;
wire P3_R1143_U234 , P3_R1143_U235 , P3_R1143_U236 , P3_R1143_U237 , P3_R1143_U238 , P3_R1143_U239 , P3_R1143_U240 , P3_R1143_U241 , P3_R1143_U242 , P3_R1143_U243;
wire P3_R1143_U244 , P3_R1143_U245 , P3_R1143_U246 , P3_R1143_U247 , P3_R1143_U248 , P3_R1143_U249 , P3_R1143_U250 , P3_R1143_U251 , P3_R1143_U252 , P3_R1143_U253;
wire P3_R1143_U254 , P3_R1143_U255 , P3_R1143_U256 , P3_R1143_U257 , P3_R1143_U258 , P3_R1143_U259 , P3_R1143_U260 , P3_R1143_U261 , P3_R1143_U262 , P3_R1143_U263;
wire P3_R1143_U264 , P3_R1143_U265 , P3_R1143_U266 , P3_R1143_U267 , P3_R1143_U268 , P3_R1143_U269 , P3_R1143_U270 , P3_R1143_U271 , P3_R1143_U272 , P3_R1143_U273;
wire P3_R1143_U274 , P3_R1143_U275 , P3_R1143_U276 , P3_R1143_U277 , P3_R1143_U278 , P3_R1143_U279 , P3_R1143_U280 , P3_R1143_U281 , P3_R1143_U282 , P3_R1143_U283;
wire P3_R1143_U284 , P3_R1143_U285 , P3_R1143_U286 , P3_R1143_U287 , P3_R1143_U288 , P3_R1143_U289 , P3_R1143_U290 , P3_R1143_U291 , P3_R1143_U292 , P3_R1143_U293;
wire P3_R1143_U294 , P3_R1143_U295 , P3_R1143_U296 , P3_R1143_U297 , P3_R1143_U298 , P3_R1143_U299 , P3_R1143_U300 , P3_R1143_U301 , P3_R1143_U302 , P3_R1143_U303;
wire P3_R1143_U304 , P3_R1143_U305 , P3_R1143_U306 , P3_R1143_U307 , P3_R1143_U308 , P3_R1143_U309 , P3_R1143_U310 , P3_R1143_U311 , P3_R1143_U312 , P3_R1143_U313;
wire P3_R1143_U314 , P3_R1143_U315 , P3_R1143_U316 , P3_R1143_U317 , P3_R1143_U318 , P3_R1143_U319 , P3_R1143_U320 , P3_R1143_U321 , P3_R1143_U322 , P3_R1143_U323;
wire P3_R1143_U324 , P3_R1143_U325 , P3_R1143_U326 , P3_R1143_U327 , P3_R1143_U328 , P3_R1143_U329 , P3_R1143_U330 , P3_R1143_U331 , P3_R1143_U332 , P3_R1143_U333;
wire P3_R1143_U334 , P3_R1143_U335 , P3_R1143_U336 , P3_R1143_U337 , P3_R1143_U338 , P3_R1143_U339 , P3_R1143_U340 , P3_R1143_U341 , P3_R1143_U342 , P3_R1143_U343;
wire P3_R1143_U344 , P3_R1143_U345 , P3_R1143_U346 , P3_R1143_U347 , P3_R1143_U348 , P3_R1143_U349 , P3_R1143_U350 , P3_R1143_U351 , P3_R1143_U352 , P3_R1143_U353;
wire P3_R1143_U354 , P3_R1143_U355 , P3_R1143_U356 , P3_R1143_U357 , P3_R1143_U358 , P3_R1143_U359 , P3_R1143_U360 , P3_R1143_U361 , P3_R1143_U362 , P3_R1143_U363;
wire P3_R1143_U364 , P3_R1143_U365 , P3_R1143_U366 , P3_R1143_U367 , P3_R1143_U368 , P3_R1143_U369 , P3_R1143_U370 , P3_R1143_U371 , P3_R1143_U372 , P3_R1143_U373;
wire P3_R1143_U374 , P3_R1143_U375 , P3_R1143_U376 , P3_R1143_U377 , P3_R1143_U378 , P3_R1143_U379 , P3_R1143_U380 , P3_R1143_U381 , P3_R1143_U382 , P3_R1143_U383;
wire P3_R1143_U384 , P3_R1143_U385 , P3_R1143_U386 , P3_R1143_U387 , P3_R1143_U388 , P3_R1143_U389 , P3_R1143_U390 , P3_R1143_U391 , P3_R1143_U392 , P3_R1143_U393;
wire P3_R1143_U394 , P3_R1143_U395 , P3_R1143_U396 , P3_R1143_U397 , P3_R1143_U398 , P3_R1143_U399 , P3_R1143_U400 , P3_R1143_U401 , P3_R1143_U402 , P3_R1143_U403;
wire P3_R1143_U404 , P3_R1143_U405 , P3_R1143_U406 , P3_R1143_U407 , P3_R1143_U408 , P3_R1143_U409 , P3_R1143_U410 , P3_R1143_U411 , P3_R1143_U412 , P3_R1143_U413;
wire P3_R1143_U414 , P3_R1143_U415 , P3_R1143_U416 , P3_R1143_U417 , P3_R1143_U418 , P3_R1143_U419 , P3_R1143_U420 , P3_R1143_U421 , P3_R1143_U422 , P3_R1143_U423;
wire P3_R1143_U424 , P3_R1143_U425 , P3_R1143_U426 , P3_R1143_U427 , P3_R1143_U428 , P3_R1143_U429 , P3_R1143_U430 , P3_R1143_U431 , P3_R1143_U432 , P3_R1143_U433;
wire P3_R1143_U434 , P3_R1143_U435 , P3_R1143_U436 , P3_R1143_U437 , P3_R1143_U438 , P3_R1143_U439 , P3_R1143_U440 , P3_R1143_U441 , P3_R1143_U442 , P3_R1143_U443;
wire P3_R1143_U444 , P3_R1143_U445 , P3_R1143_U446 , P3_R1143_U447 , P3_R1143_U448 , P3_R1143_U449 , P3_R1143_U450 , P3_R1143_U451 , P3_R1143_U452 , P3_R1143_U453;
wire P3_R1143_U454 , P3_R1143_U455 , P3_R1143_U456 , P3_R1143_U457 , P3_R1143_U458 , P3_R1143_U459 , P3_R1143_U460 , P3_R1143_U461 , P3_R1143_U462 , P3_R1143_U463;
wire P3_R1143_U464 , P3_R1143_U465 , P3_R1143_U466 , P3_R1143_U467 , P3_R1143_U468 , P3_R1143_U469 , P3_R1143_U470 , P3_R1143_U471 , P3_R1143_U472 , P3_R1143_U473;
wire P3_R1143_U474 , P3_R1143_U475 , P3_R1143_U476 , P3_R1143_U477 , P3_R1143_U478 , P3_R1143_U479 , P3_R1143_U480 , P3_R1143_U481 , P3_R1143_U482 , P3_R1143_U483;
wire P3_R1143_U484 , P3_R1143_U485 , P3_R1143_U486 , P3_R1143_U487 , P3_R1143_U488 , P3_R1143_U489 , P3_R1143_U490 , P3_R1143_U491 , P3_R1143_U492 , P3_R1143_U493;
wire P3_R1143_U494 , P3_R1143_U495 , P3_R1143_U496 , P3_R1143_U497 , P3_R1143_U498 , P3_R1143_U499 , P3_R1143_U500 , P3_R1143_U501 , P3_R1143_U502 , P3_R1143_U503;
wire P3_R1143_U504 , P3_R1158_U4 , P3_R1158_U5 , P3_R1158_U6 , P3_R1158_U7 , P3_R1158_U8 , P3_R1158_U9 , P3_R1158_U10 , P3_R1158_U11 , P3_R1158_U12;
wire P3_R1158_U13 , P3_R1158_U14 , P3_R1158_U15 , P3_R1158_U16 , P3_R1158_U17 , P3_R1158_U18 , P3_R1158_U19 , P3_R1158_U20 , P3_R1158_U21 , P3_R1158_U22;
wire P3_R1158_U23 , P3_R1158_U24 , P3_R1158_U25 , P3_R1158_U26 , P3_R1158_U27 , P3_R1158_U28 , P3_R1158_U29 , P3_R1158_U30 , P3_R1158_U31 , P3_R1158_U32;
wire P3_R1158_U33 , P3_R1158_U34 , P3_R1158_U35 , P3_R1158_U36 , P3_R1158_U37 , P3_R1158_U38 , P3_R1158_U39 , P3_R1158_U40 , P3_R1158_U41 , P3_R1158_U42;
wire P3_R1158_U43 , P3_R1158_U44 , P3_R1158_U45 , P3_R1158_U46 , P3_R1158_U47 , P3_R1158_U48 , P3_R1158_U49 , P3_R1158_U50 , P3_R1158_U51 , P3_R1158_U52;
wire P3_R1158_U53 , P3_R1158_U54 , P3_R1158_U55 , P3_R1158_U56 , P3_R1158_U57 , P3_R1158_U58 , P3_R1158_U59 , P3_R1158_U60 , P3_R1158_U61 , P3_R1158_U62;
wire P3_R1158_U63 , P3_R1158_U64 , P3_R1158_U65 , P3_R1158_U66 , P3_R1158_U67 , P3_R1158_U68 , P3_R1158_U69 , P3_R1158_U70 , P3_R1158_U71 , P3_R1158_U72;
wire P3_R1158_U73 , P3_R1158_U74 , P3_R1158_U75 , P3_R1158_U76 , P3_R1158_U77 , P3_R1158_U78 , P3_R1158_U79 , P3_R1158_U80 , P3_R1158_U81 , P3_R1158_U82;
wire P3_R1158_U83 , P3_R1158_U84 , P3_R1158_U85 , P3_R1158_U86 , P3_R1158_U87 , P3_R1158_U88 , P3_R1158_U89 , P3_R1158_U90 , P3_R1158_U91 , P3_R1158_U92;
wire P3_R1158_U93 , P3_R1158_U94 , P3_R1158_U95 , P3_R1158_U96 , P3_R1158_U97 , P3_R1158_U98 , P3_R1158_U99 , P3_R1158_U100 , P3_R1158_U101 , P3_R1158_U102;
wire P3_R1158_U103 , P3_R1158_U104 , P3_R1158_U105 , P3_R1158_U106 , P3_R1158_U107 , P3_R1158_U108 , P3_R1158_U109 , P3_R1158_U110 , P3_R1158_U111 , P3_R1158_U112;
wire P3_R1158_U113 , P3_R1158_U114 , P3_R1158_U115 , P3_R1158_U116 , P3_R1158_U117 , P3_R1158_U118 , P3_R1158_U119 , P3_R1158_U120 , P3_R1158_U121 , P3_R1158_U122;
wire P3_R1158_U123 , P3_R1158_U124 , P3_R1158_U125 , P3_R1158_U126 , P3_R1158_U127 , P3_R1158_U128 , P3_R1158_U129 , P3_R1158_U130 , P3_R1158_U131 , P3_R1158_U132;
wire P3_R1158_U133 , P3_R1158_U134 , P3_R1158_U135 , P3_R1158_U136 , P3_R1158_U137 , P3_R1158_U138 , P3_R1158_U139 , P3_R1158_U140 , P3_R1158_U141 , P3_R1158_U142;
wire P3_R1158_U143 , P3_R1158_U144 , P3_R1158_U145 , P3_R1158_U146 , P3_R1158_U147 , P3_R1158_U148 , P3_R1158_U149 , P3_R1158_U150 , P3_R1158_U151 , P3_R1158_U152;
wire P3_R1158_U153 , P3_R1158_U154 , P3_R1158_U155 , P3_R1158_U156 , P3_R1158_U157 , P3_R1158_U158 , P3_R1158_U159 , P3_R1158_U160 , P3_R1158_U161 , P3_R1158_U162;
wire P3_R1158_U163 , P3_R1158_U164 , P3_R1158_U165 , P3_R1158_U166 , P3_R1158_U167 , P3_R1158_U168 , P3_R1158_U169 , P3_R1158_U170 , P3_R1158_U171 , P3_R1158_U172;
wire P3_R1158_U173 , P3_R1158_U174 , P3_R1158_U175 , P3_R1158_U176 , P3_R1158_U177 , P3_R1158_U178 , P3_R1158_U179 , P3_R1158_U180 , P3_R1158_U181 , P3_R1158_U182;
wire P3_R1158_U183 , P3_R1158_U184 , P3_R1158_U185 , P3_R1158_U186 , P3_R1158_U187 , P3_R1158_U188 , P3_R1158_U189 , P3_R1158_U190 , P3_R1158_U191 , P3_R1158_U192;
wire P3_R1158_U193 , P3_R1158_U194 , P3_R1158_U195 , P3_R1158_U196 , P3_R1158_U197 , P3_R1158_U198 , P3_R1158_U199 , P3_R1158_U200 , P3_R1158_U201 , P3_R1158_U202;
wire P3_R1158_U203 , P3_R1158_U204 , P3_R1158_U205 , P3_R1158_U206 , P3_R1158_U207 , P3_R1158_U208 , P3_R1158_U209 , P3_R1158_U210 , P3_R1158_U211 , P3_R1158_U212;
wire P3_R1158_U213 , P3_R1158_U214 , P3_R1158_U215 , P3_R1158_U216 , P3_R1158_U217 , P3_R1158_U218 , P3_R1158_U219 , P3_R1158_U220 , P3_R1158_U221 , P3_R1158_U222;
wire P3_R1158_U223 , P3_R1158_U224 , P3_R1158_U225 , P3_R1158_U226 , P3_R1158_U227 , P3_R1158_U228 , P3_R1158_U229 , P3_R1158_U230 , P3_R1158_U231 , P3_R1158_U232;
wire P3_R1158_U233 , P3_R1158_U234 , P3_R1158_U235 , P3_R1158_U236 , P3_R1158_U237 , P3_R1158_U238 , P3_R1158_U239 , P3_R1158_U240 , P3_R1158_U241 , P3_R1158_U242;
wire P3_R1158_U243 , P3_R1158_U244 , P3_R1158_U245 , P3_R1158_U246 , P3_R1158_U247 , P3_R1158_U248 , P3_R1158_U249 , P3_R1158_U250 , P3_R1158_U251 , P3_R1158_U252;
wire P3_R1158_U253 , P3_R1158_U254 , P3_R1158_U255 , P3_R1158_U256 , P3_R1158_U257 , P3_R1158_U258 , P3_R1158_U259 , P3_R1158_U260 , P3_R1158_U261 , P3_R1158_U262;
wire P3_R1158_U263 , P3_R1158_U264 , P3_R1158_U265 , P3_R1158_U266 , P3_R1158_U267 , P3_R1158_U268 , P3_R1158_U269 , P3_R1158_U270 , P3_R1158_U271 , P3_R1158_U272;
wire P3_R1158_U273 , P3_R1158_U274 , P3_R1158_U275 , P3_R1158_U276 , P3_R1158_U277 , P3_R1158_U278 , P3_R1158_U279 , P3_R1158_U280 , P3_R1158_U281 , P3_R1158_U282;
wire P3_R1158_U283 , P3_R1158_U284 , P3_R1158_U285 , P3_R1158_U286 , P3_R1158_U287 , P3_R1158_U288 , P3_R1158_U289 , P3_R1158_U290 , P3_R1158_U291 , P3_R1158_U292;
wire P3_R1158_U293 , P3_R1158_U294 , P3_R1158_U295 , P3_R1158_U296 , P3_R1158_U297 , P3_R1158_U298 , P3_R1158_U299 , P3_R1158_U300 , P3_R1158_U301 , P3_R1158_U302;
wire P3_R1158_U303 , P3_R1158_U304 , P3_R1158_U305 , P3_R1158_U306 , P3_R1158_U307 , P3_R1158_U308 , P3_R1158_U309 , P3_R1158_U310 , P3_R1158_U311 , P3_R1158_U312;
wire P3_R1158_U313 , P3_R1158_U314 , P3_R1158_U315 , P3_R1158_U316 , P3_R1158_U317 , P3_R1158_U318 , P3_R1158_U319 , P3_R1158_U320 , P3_R1158_U321 , P3_R1158_U322;
wire P3_R1158_U323 , P3_R1158_U324 , P3_R1158_U325 , P3_R1158_U326 , P3_R1158_U327 , P3_R1158_U328 , P3_R1158_U329 , P3_R1158_U330 , P3_R1158_U331 , P3_R1158_U332;
wire P3_R1158_U333 , P3_R1158_U334 , P3_R1158_U335 , P3_R1158_U336 , P3_R1158_U337 , P3_R1158_U338 , P3_R1158_U339 , P3_R1158_U340 , P3_R1158_U341 , P3_R1158_U342;
wire P3_R1158_U343 , P3_R1158_U344 , P3_R1158_U345 , P3_R1158_U346 , P3_R1158_U347 , P3_R1158_U348 , P3_R1158_U349 , P3_R1158_U350 , P3_R1158_U351 , P3_R1158_U352;
wire P3_R1158_U353 , P3_R1158_U354 , P3_R1158_U355 , P3_R1158_U356 , P3_R1158_U357 , P3_R1158_U358 , P3_R1158_U359 , P3_R1158_U360 , P3_R1158_U361 , P3_R1158_U362;
wire P3_R1158_U363 , P3_R1158_U364 , P3_R1158_U365 , P3_R1158_U366 , P3_R1158_U367 , P3_R1158_U368 , P3_R1158_U369 , P3_R1158_U370 , P3_R1158_U371 , P3_R1158_U372;
wire P3_R1158_U373 , P3_R1158_U374 , P3_R1158_U375 , P3_R1158_U376 , P3_R1158_U377 , P3_R1158_U378 , P3_R1158_U379 , P3_R1158_U380 , P3_R1158_U381 , P3_R1158_U382;
wire P3_R1158_U383 , P3_R1158_U384 , P3_R1158_U385 , P3_R1158_U386 , P3_R1158_U387 , P3_R1158_U388 , P3_R1158_U389 , P3_R1158_U390 , P3_R1158_U391 , P3_R1158_U392;
wire P3_R1158_U393 , P3_R1158_U394 , P3_R1158_U395 , P3_R1158_U396 , P3_R1158_U397 , P3_R1158_U398 , P3_R1158_U399 , P3_R1158_U400 , P3_R1158_U401 , P3_R1158_U402;
wire P3_R1158_U403 , P3_R1158_U404 , P3_R1158_U405 , P3_R1158_U406 , P3_R1158_U407 , P3_R1158_U408 , P3_R1158_U409 , P3_R1158_U410 , P3_R1158_U411 , P3_R1158_U412;
wire P3_R1158_U413 , P3_R1158_U414 , P3_R1158_U415 , P3_R1158_U416 , P3_R1158_U417 , P3_R1158_U418 , P3_R1158_U419 , P3_R1158_U420 , P3_R1158_U421 , P3_R1158_U422;
wire P3_R1158_U423 , P3_R1158_U424 , P3_R1158_U425 , P3_R1158_U426 , P3_R1158_U427 , P3_R1158_U428 , P3_R1158_U429 , P3_R1158_U430 , P3_R1158_U431 , P3_R1158_U432;
wire P3_R1158_U433 , P3_R1158_U434 , P3_R1158_U435 , P3_R1158_U436 , P3_R1158_U437 , P3_R1158_U438 , P3_R1158_U439 , P3_R1158_U440 , P3_R1158_U441 , P3_R1158_U442;
wire P3_R1158_U443 , P3_R1158_U444 , P3_R1158_U445 , P3_R1158_U446 , P3_R1158_U447 , P3_R1158_U448 , P3_R1158_U449 , P3_R1158_U450 , P3_R1158_U451 , P3_R1158_U452;
wire P3_R1158_U453 , P3_R1158_U454 , P3_R1158_U455 , P3_R1158_U456 , P3_R1158_U457 , P3_R1158_U458 , P3_R1158_U459 , P3_R1158_U460 , P3_R1158_U461 , P3_R1158_U462;
wire P3_R1158_U463 , P3_R1158_U464 , P3_R1158_U465 , P3_R1158_U466 , P3_R1158_U467 , P3_R1158_U468 , P3_R1158_U469 , P3_R1158_U470 , P3_R1158_U471 , P3_R1158_U472;
wire P3_R1158_U473 , P3_R1158_U474 , P3_R1158_U475 , P3_R1158_U476 , P3_R1158_U477 , P3_R1158_U478 , P3_R1158_U479 , P3_R1158_U480 , P3_R1158_U481 , P3_R1158_U482;
wire P3_R1158_U483 , P3_R1158_U484 , P3_R1158_U485 , P3_R1158_U486 , P3_R1158_U487 , P3_R1158_U488 , P3_R1158_U489 , P3_R1158_U490 , P3_R1158_U491 , P3_R1158_U492;
wire P3_R1158_U493 , P3_R1158_U494 , P3_R1158_U495 , P3_R1158_U496 , P3_R1158_U497 , P3_R1158_U498 , P3_R1158_U499 , P3_R1158_U500 , P3_R1158_U501 , P3_R1158_U502;
wire P3_R1158_U503 , P3_R1158_U504 , P3_R1158_U505 , P3_R1158_U506 , P3_R1158_U507 , P3_R1158_U508 , P3_R1158_U509 , P3_R1158_U510 , P3_R1158_U511 , P3_R1158_U512;
wire P3_R1158_U513 , P3_R1158_U514 , P3_R1158_U515 , P3_R1158_U516 , P3_R1158_U517 , P3_R1158_U518 , P3_R1158_U519 , P3_R1158_U520 , P3_R1158_U521 , P3_R1158_U522;
wire P3_R1158_U523 , P3_R1158_U524 , P3_R1158_U525 , P3_R1158_U526 , P3_R1158_U527 , P3_R1158_U528 , P3_R1158_U529 , P3_R1158_U530 , P3_R1158_U531 , P3_R1158_U532;
wire P3_R1158_U533 , P3_R1158_U534 , P3_R1158_U535 , P3_R1158_U536 , P3_R1158_U537 , P3_R1158_U538 , P3_R1158_U539 , P3_R1158_U540 , P3_R1158_U541 , P3_R1158_U542;
wire P3_R1158_U543 , P3_R1158_U544 , P3_R1158_U545 , P3_R1158_U546 , P3_R1158_U547 , P3_R1158_U548 , P3_R1158_U549 , P3_R1158_U550 , P3_R1158_U551 , P3_R1158_U552;
wire P3_R1158_U553 , P3_R1158_U554 , P3_R1158_U555 , P3_R1158_U556 , P3_R1158_U557 , P3_R1158_U558 , P3_R1158_U559 , P3_R1158_U560 , P3_R1158_U561 , P3_R1158_U562;
wire P3_R1158_U563 , P3_R1158_U564 , P3_R1158_U565 , P3_R1158_U566 , P3_R1158_U567 , P3_R1158_U568 , P3_R1158_U569 , P3_R1158_U570 , P3_R1158_U571 , P3_R1158_U572;
wire P3_R1158_U573 , P3_R1158_U574 , P3_R1158_U575 , P3_R1158_U576 , P3_R1158_U577 , P3_R1158_U578 , P3_R1158_U579 , P3_R1158_U580 , P3_R1158_U581 , P3_R1158_U582;
wire P3_R1158_U583 , P3_R1158_U584 , P3_R1158_U585 , P3_R1158_U586 , P3_R1158_U587 , P3_R1158_U588 , P3_R1158_U589 , P3_R1158_U590 , P3_R1158_U591 , P3_R1158_U592;
wire P3_R1158_U593 , P3_R1158_U594 , P3_R1158_U595 , P3_R1158_U596 , P3_R1158_U597 , P3_R1158_U598 , P3_R1158_U599 , P3_R1158_U600 , P3_R1158_U601 , P3_R1158_U602;
wire P3_R1158_U603 , P3_R1158_U604 , P3_R1158_U605 , P3_R1158_U606 , P3_R1158_U607 , P3_R1158_U608 , P3_R1158_U609 , P3_R1158_U610 , P3_R1158_U611 , P3_R1158_U612;
wire P3_R1158_U613 , P3_R1158_U614 , P3_R1158_U615 , P3_R1158_U616 , P3_R1158_U617 , P3_R1158_U618 , P3_R1158_U619 , P3_R1158_U620 , P3_R1158_U621 , P3_R1158_U622;
wire P3_R1158_U623 , P3_R1158_U624 , P3_R1158_U625 , P3_R1158_U626 , P3_R1158_U627 , P3_R1158_U628 , P3_R1158_U629 , P3_R1158_U630 , P3_R1158_U631 , P3_R1158_U632;
wire P3_R1131_U6 , P3_R1131_U7 , P3_R1131_U8 , P3_R1131_U9 , P3_R1131_U10 , P3_R1131_U11 , P3_R1131_U12 , P3_R1131_U13 , P3_R1131_U14 , P3_R1131_U15;
wire P3_R1131_U16 , P3_R1131_U17 , P3_R1131_U18 , P3_R1131_U19 , P3_R1131_U20 , P3_R1131_U21 , P3_R1131_U22 , P3_R1131_U23 , P3_R1131_U24 , P3_R1131_U25;
wire P3_R1131_U26 , P3_R1131_U27 , P3_R1131_U28 , P3_R1131_U29 , P3_R1131_U30 , P3_R1131_U31 , P3_R1131_U32 , P3_R1131_U33 , P3_R1131_U34 , P3_R1131_U35;
wire P3_R1131_U36 , P3_R1131_U37 , P3_R1131_U38 , P3_R1131_U39 , P3_R1131_U40 , P3_R1131_U41 , P3_R1131_U42 , P3_R1131_U43 , P3_R1131_U44 , P3_R1131_U45;
wire P3_R1131_U46 , P3_R1131_U47 , P3_R1131_U48 , P3_R1131_U49 , P3_R1131_U50 , P3_R1131_U51 , P3_R1131_U52 , P3_R1131_U53 , P3_R1131_U54 , P3_R1131_U55;
wire P3_R1131_U56 , P3_R1131_U57 , P3_R1131_U58 , P3_R1131_U59 , P3_R1131_U60 , P3_R1131_U61 , P3_R1131_U62 , P3_R1131_U63 , P3_R1131_U64 , P3_R1131_U65;
wire P3_R1131_U66 , P3_R1131_U67 , P3_R1131_U68 , P3_R1131_U69 , P3_R1131_U70 , P3_R1131_U71 , P3_R1131_U72 , P3_R1131_U73 , P3_R1131_U74 , P3_R1131_U75;
wire P3_R1131_U76 , P3_R1131_U77 , P3_R1131_U78 , P3_R1131_U79 , P3_R1131_U80 , P3_R1131_U81 , P3_R1131_U82 , P3_R1131_U83 , P3_R1131_U84 , P3_R1131_U85;
wire P3_R1131_U86 , P3_R1131_U87 , P3_R1131_U88 , P3_R1131_U89 , P3_R1131_U90 , P3_R1131_U91 , P3_R1131_U92 , P3_R1131_U93 , P3_R1131_U94 , P3_R1131_U95;
wire P3_R1131_U96 , P3_R1131_U97 , P3_R1131_U98 , P3_R1131_U99 , P3_R1131_U100 , P3_R1131_U101 , P3_R1131_U102 , P3_R1131_U103 , P3_R1131_U104 , P3_R1131_U105;
wire P3_R1131_U106 , P3_R1131_U107 , P3_R1131_U108 , P3_R1131_U109 , P3_R1131_U110 , P3_R1131_U111 , P3_R1131_U112 , P3_R1131_U113 , P3_R1131_U114 , P3_R1131_U115;
wire P3_R1131_U116 , P3_R1131_U117 , P3_R1131_U118 , P3_R1131_U119 , P3_R1131_U120 , P3_R1131_U121 , P3_R1131_U122 , P3_R1131_U123 , P3_R1131_U124 , P3_R1131_U125;
wire P3_R1131_U126 , P3_R1131_U127 , P3_R1131_U128 , P3_R1131_U129 , P3_R1131_U130 , P3_R1131_U131 , P3_R1131_U132 , P3_R1131_U133 , P3_R1131_U134 , P3_R1131_U135;
wire P3_R1131_U136 , P3_R1131_U137 , P3_R1131_U138 , P3_R1131_U139 , P3_R1131_U140 , P3_R1131_U141 , P3_R1131_U142 , P3_R1131_U143 , P3_R1131_U144 , P3_R1131_U145;
wire P3_R1131_U146 , P3_R1131_U147 , P3_R1131_U148 , P3_R1131_U149 , P3_R1131_U150 , P3_R1131_U151 , P3_R1131_U152 , P3_R1131_U153 , P3_R1131_U154 , P3_R1131_U155;
wire P3_R1131_U156 , P3_R1131_U157 , P3_R1131_U158 , P3_R1131_U159 , P3_R1131_U160 , P3_R1131_U161 , P3_R1131_U162 , P3_R1131_U163 , P3_R1131_U164 , P3_R1131_U165;
wire P3_R1131_U166 , P3_R1131_U167 , P3_R1131_U168 , P3_R1131_U169 , P3_R1131_U170 , P3_R1131_U171 , P3_R1131_U172 , P3_R1131_U173 , P3_R1131_U174 , P3_R1131_U175;
wire P3_R1131_U176 , P3_R1131_U177 , P3_R1131_U178 , P3_R1131_U179 , P3_R1131_U180 , P3_R1131_U181 , P3_R1131_U182 , P3_R1131_U183 , P3_R1131_U184 , P3_R1131_U185;
wire P3_R1131_U186 , P3_R1131_U187 , P3_R1131_U188 , P3_R1131_U189 , P3_R1131_U190 , P3_R1131_U191 , P3_R1131_U192 , P3_R1131_U193 , P3_R1131_U194 , P3_R1131_U195;
wire P3_R1131_U196 , P3_R1131_U197 , P3_R1131_U198 , P3_R1131_U199 , P3_R1131_U200 , P3_R1131_U201 , P3_R1131_U202 , P3_R1131_U203 , P3_R1131_U204 , P3_R1131_U205;
wire P3_R1131_U206 , P3_R1131_U207 , P3_R1131_U208 , P3_R1131_U209 , P3_R1131_U210 , P3_R1131_U211 , P3_R1131_U212 , P3_R1131_U213 , P3_R1131_U214 , P3_R1131_U215;
wire P3_R1131_U216 , P3_R1131_U217 , P3_R1131_U218 , P3_R1131_U219 , P3_R1131_U220 , P3_R1131_U221 , P3_R1131_U222 , P3_R1131_U223 , P3_R1131_U224 , P3_R1131_U225;
wire P3_R1131_U226 , P3_R1131_U227 , P3_R1131_U228 , P3_R1131_U229 , P3_R1131_U230 , P3_R1131_U231 , P3_R1131_U232 , P3_R1131_U233 , P3_R1131_U234 , P3_R1131_U235;
wire P3_R1131_U236 , P3_R1131_U237 , P3_R1131_U238 , P3_R1131_U239 , P3_R1131_U240 , P3_R1131_U241 , P3_R1131_U242 , P3_R1131_U243 , P3_R1131_U244 , P3_R1131_U245;
wire P3_R1131_U246 , P3_R1131_U247 , P3_R1131_U248 , P3_R1131_U249 , P3_R1131_U250 , P3_R1131_U251 , P3_R1131_U252 , P3_R1131_U253 , P3_R1131_U254 , P3_R1131_U255;
wire P3_R1131_U256 , P3_R1131_U257 , P3_R1131_U258 , P3_R1131_U259 , P3_R1131_U260 , P3_R1131_U261 , P3_R1131_U262 , P3_R1131_U263 , P3_R1131_U264 , P3_R1131_U265;
wire P3_R1131_U266 , P3_R1131_U267 , P3_R1131_U268 , P3_R1131_U269 , P3_R1131_U270 , P3_R1131_U271 , P3_R1131_U272 , P3_R1131_U273 , P3_R1131_U274 , P3_R1131_U275;
wire P3_R1131_U276 , P3_R1131_U277 , P3_R1131_U278 , P3_R1131_U279 , P3_R1131_U280 , P3_R1131_U281 , P3_R1131_U282 , P3_R1131_U283 , P3_R1131_U284 , P3_R1131_U285;
wire P3_R1131_U286 , P3_R1131_U287 , P3_R1131_U288 , P3_R1131_U289 , P3_R1131_U290 , P3_R1131_U291 , P3_R1131_U292 , P3_R1131_U293 , P3_R1131_U294 , P3_R1131_U295;
wire P3_R1131_U296 , P3_R1131_U297 , P3_R1131_U298 , P3_R1131_U299 , P3_R1131_U300 , P3_R1131_U301 , P3_R1131_U302 , P3_R1131_U303 , P3_R1131_U304 , P3_R1131_U305;
wire P3_R1131_U306 , P3_R1131_U307 , P3_R1131_U308 , P3_R1131_U309 , P3_R1131_U310 , P3_R1131_U311 , P3_R1131_U312 , P3_R1131_U313 , P3_R1131_U314 , P3_R1131_U315;
wire P3_R1131_U316 , P3_R1131_U317 , P3_R1131_U318 , P3_R1131_U319 , P3_R1131_U320 , P3_R1131_U321 , P3_R1131_U322 , P3_R1131_U323 , P3_R1131_U324 , P3_R1131_U325;
wire P3_R1131_U326 , P3_R1131_U327 , P3_R1131_U328 , P3_R1131_U329 , P3_R1131_U330 , P3_R1131_U331 , P3_R1131_U332 , P3_R1131_U333 , P3_R1131_U334 , P3_R1131_U335;
wire P3_R1131_U336 , P3_R1131_U337 , P3_R1131_U338 , P3_R1131_U339 , P3_R1131_U340 , P3_R1131_U341 , P3_R1131_U342 , P3_R1131_U343 , P3_R1131_U344 , P3_R1131_U345;
wire P3_R1131_U346 , P3_R1131_U347 , P3_R1131_U348 , P3_R1131_U349 , P3_R1131_U350 , P3_R1131_U351 , P3_R1131_U352 , P3_R1131_U353 , P3_R1131_U354 , P3_R1131_U355;
wire P3_R1131_U356 , P3_R1131_U357 , P3_R1131_U358 , P3_R1131_U359 , P3_R1131_U360 , P3_R1131_U361 , P3_R1131_U362 , P3_R1131_U363 , P3_R1131_U364 , P3_R1131_U365;
wire P3_R1131_U366 , P3_R1131_U367 , P3_R1131_U368 , P3_R1131_U369 , P3_R1131_U370 , P3_R1131_U371 , P3_R1131_U372 , P3_R1131_U373 , P3_R1131_U374 , P3_R1131_U375;
wire P3_R1131_U376 , P3_R1131_U377 , P3_R1131_U378 , P3_R1131_U379 , P3_R1131_U380 , P3_R1131_U381 , P3_R1131_U382 , P3_R1131_U383 , P3_R1131_U384 , P3_R1131_U385;
wire P3_R1131_U386 , P3_R1131_U387 , P3_R1131_U388 , P3_R1131_U389 , P3_R1131_U390 , P3_R1131_U391 , P3_R1131_U392 , P3_R1131_U393 , P3_R1131_U394 , P3_R1131_U395;
wire P3_R1131_U396 , P3_R1131_U397 , P3_R1131_U398 , P3_R1131_U399 , P3_R1131_U400 , P3_R1131_U401 , P3_R1131_U402 , P3_R1131_U403 , P3_R1131_U404 , P3_R1131_U405;
wire P3_R1131_U406 , P3_R1131_U407 , P3_R1131_U408 , P3_R1131_U409 , P3_R1131_U410 , P3_R1131_U411 , P3_R1131_U412 , P3_R1131_U413 , P3_R1131_U414 , P3_R1131_U415;
wire P3_R1131_U416 , P3_R1131_U417 , P3_R1131_U418 , P3_R1131_U419 , P3_R1131_U420 , P3_R1131_U421 , P3_R1131_U422 , P3_R1131_U423 , P3_R1131_U424 , P3_R1131_U425;
wire P3_R1131_U426 , P3_R1131_U427 , P3_R1131_U428 , P3_R1131_U429 , P3_R1131_U430 , P3_R1131_U431 , P3_R1131_U432 , P3_R1131_U433 , P3_R1131_U434 , P3_R1131_U435;
wire P3_R1131_U436 , P3_R1131_U437 , P3_R1131_U438 , P3_R1131_U439 , P3_R1131_U440 , P3_R1131_U441 , P3_R1131_U442 , P3_R1131_U443 , P3_R1131_U444 , P3_R1131_U445;
wire P3_R1131_U446 , P3_R1131_U447 , P3_R1131_U448 , P3_R1131_U449 , P3_R1131_U450 , P3_R1131_U451 , P3_R1131_U452 , P3_R1131_U453 , P3_R1131_U454 , P3_R1131_U455;
wire P3_R1131_U456 , P3_R1131_U457 , P3_R1131_U458 , P3_R1131_U459 , P3_R1131_U460 , P3_R1131_U461 , P3_R1131_U462 , P3_R1131_U463 , P3_R1131_U464 , P3_R1131_U465;
wire P3_R1131_U466 , P3_R1131_U467 , P3_R1131_U468 , P3_R1131_U469 , P3_R1131_U470 , P3_R1131_U471 , P3_R1131_U472 , P3_R1131_U473 , P3_R1131_U474 , P3_R1131_U475;
wire P3_R1131_U476 , P3_R1131_U477 , P3_R1131_U478 , P3_R1131_U479 , P3_R1131_U480 , P3_R1131_U481 , P3_R1131_U482 , P3_R1131_U483 , P3_R1131_U484 , P3_R1131_U485;
wire P3_R1054_U6 , P3_R1054_U7 , P3_R1054_U8 , P3_R1054_U9 , P3_R1054_U10 , P3_R1054_U11 , P3_R1054_U12 , P3_R1054_U13 , P3_R1054_U14 , P3_R1054_U15;
wire P3_R1054_U16 , P3_R1054_U17 , P3_R1054_U18 , P3_R1054_U19 , P3_R1054_U20 , P3_R1054_U21 , P3_R1054_U22 , P3_R1054_U23 , P3_R1054_U24 , P3_R1054_U25;
wire P3_R1054_U26 , P3_R1054_U27 , P3_R1054_U28 , P3_R1054_U29 , P3_R1054_U30 , P3_R1054_U31 , P3_R1054_U32 , P3_R1054_U33 , P3_R1054_U34 , P3_R1054_U35;
wire P3_R1054_U36 , P3_R1054_U37 , P3_R1054_U38 , P3_R1054_U39 , P3_R1054_U40 , P3_R1054_U41 , P3_R1054_U42 , P3_R1054_U43 , P3_R1054_U44 , P3_R1054_U45;
wire P3_R1054_U46 , P3_R1054_U47 , P3_R1054_U48 , P3_R1054_U49 , P3_R1054_U50 , P3_R1054_U51 , P3_R1054_U52 , P3_R1054_U53 , P3_R1054_U54 , P3_R1054_U55;
wire P3_R1054_U56 , P3_R1054_U57 , P3_R1054_U58 , P3_R1054_U59 , P3_R1054_U60 , P3_R1054_U61 , P3_R1054_U62 , P3_R1054_U63 , P3_R1054_U64 , P3_R1054_U65;
wire P3_R1054_U66 , P3_R1054_U67 , P3_R1054_U68 , P3_R1054_U69 , P3_R1054_U70 , P3_R1054_U71 , P3_R1054_U72 , P3_R1054_U73 , P3_R1054_U74 , P3_R1054_U75;
wire P3_R1054_U76 , P3_R1054_U77 , P3_R1054_U78 , P3_R1054_U79 , P3_R1054_U80 , P3_R1054_U81 , P3_R1054_U82 , P3_R1054_U83 , P3_R1054_U84 , P3_R1054_U85;
wire P3_R1054_U86 , P3_R1054_U87 , P3_R1054_U88 , P3_R1054_U89 , P3_R1054_U90 , P3_R1054_U91 , P3_R1054_U92 , P3_R1054_U93 , P3_R1054_U94 , P3_R1054_U95;
wire P3_R1054_U96 , P3_R1054_U97 , P3_R1054_U98 , P3_R1054_U99 , P3_R1054_U100 , P3_R1054_U101 , P3_R1054_U102 , P3_R1054_U103 , P3_R1054_U104 , P3_R1054_U105;
wire P3_R1054_U106 , P3_R1054_U107 , P3_R1054_U108 , P3_R1054_U109 , P3_R1054_U110 , P3_R1054_U111 , P3_R1054_U112 , P3_R1054_U113 , P3_R1054_U114 , P3_R1054_U115;
wire P3_R1054_U116 , P3_R1054_U117 , P3_R1054_U118 , P3_R1054_U119 , P3_R1054_U120 , P3_R1054_U121 , P3_R1054_U122 , P3_R1054_U123 , P3_R1054_U124 , P3_R1054_U125;
wire P3_R1054_U126 , P3_R1054_U127 , P3_R1054_U128 , P3_R1054_U129 , P3_R1054_U130 , P3_R1054_U131 , P3_R1054_U132 , P3_R1054_U133 , P3_R1054_U134 , P3_R1054_U135;
wire P3_R1054_U136 , P3_R1054_U137 , P3_R1054_U138 , P3_R1054_U139 , P3_R1054_U140 , P3_R1054_U141 , P3_R1054_U142 , P3_R1054_U143 , P3_R1054_U144 , P3_R1054_U145;
wire P3_R1054_U146 , P3_R1054_U147 , P3_R1054_U148 , P3_R1054_U149 , P3_R1054_U150 , P3_R1054_U151 , P3_R1054_U152 , P3_R1054_U153 , P3_R1054_U154 , P3_R1054_U155;
wire P3_R1054_U156 , P3_R1054_U157 , P3_R1054_U158 , P3_R1054_U159 , P3_R1054_U160 , P3_R1054_U161 , P3_R1054_U162 , P3_R1054_U163 , P3_R1054_U164 , P3_R1054_U165;
wire P3_R1054_U166 , P3_R1054_U167 , P3_R1054_U168 , P3_R1054_U169 , P3_R1054_U170 , P3_R1054_U171 , P3_R1054_U172 , P3_R1054_U173 , P3_R1054_U174 , P3_R1054_U175;
wire P3_R1054_U176 , P3_R1054_U177 , P3_R1054_U178 , P3_R1054_U179 , P3_R1054_U180 , P3_R1054_U181 , P3_R1054_U182 , P3_R1054_U183 , P3_R1054_U184 , P3_R1054_U185;
wire P3_R1054_U186 , P3_R1054_U187 , P3_R1054_U188 , P3_R1054_U189 , P3_R1054_U190 , P3_R1054_U191 , P3_R1054_U192 , P3_R1054_U193 , P3_R1054_U194 , P3_R1054_U195;
wire P3_R1054_U196 , P3_R1054_U197 , P3_R1054_U198 , P3_R1054_U199 , P3_R1054_U200 , P3_R1054_U201 , P3_R1054_U202 , P3_R1054_U203 , P3_R1054_U204 , P3_R1054_U205;
wire P3_R1054_U206 , P3_R1054_U207 , P3_R1054_U208 , P3_R1054_U209 , P3_R1054_U210 , P3_R1054_U211 , P3_R1054_U212 , P3_R1054_U213 , P3_R1054_U214 , P3_R1054_U215;
wire P3_R1054_U216 , P3_R1054_U217 , P3_R1054_U218 , P3_R1054_U219 , P3_R1054_U220 , P3_R1054_U221 , P3_R1054_U222 , P3_R1054_U223 , P3_R1054_U224 , P3_R1054_U225;
wire P3_R1054_U226 , P3_R1054_U227 , P3_R1054_U228 , P3_R1054_U229 , P3_R1054_U230 , P3_R1054_U231 , P3_R1054_U232 , P3_R1054_U233 , P3_R1054_U234 , P3_R1054_U235;
wire P3_R1054_U236 , P3_R1054_U237 , P3_R1054_U238 , P3_R1054_U239 , P3_R1054_U240 , P3_R1054_U241 , P3_R1054_U242 , P3_R1054_U243 , P3_R1054_U244 , P3_R1054_U245;
wire P3_R1054_U246 , P3_R1054_U247 , P3_R1054_U248 , P3_R1054_U249 , P3_R1054_U250 , P3_R1054_U251 , P3_R1054_U252 , P3_R1054_U253 , P3_R1054_U254 , P3_R1054_U255;
wire P3_R1054_U256 , P3_R1054_U257 , P3_R1054_U258 , P3_R1054_U259 , P3_R1054_U260 , P3_R1054_U261 , P3_R1054_U262 , P3_R1054_U263 , P3_R1054_U264 , P3_R1054_U265;
wire P3_R1054_U266 , P3_R1054_U267 , P3_R1054_U268 , P3_R1054_U269 , P3_R1054_U270 , P3_R1054_U271 , P3_R1054_U272 , P3_R1054_U273 , P3_R1054_U274 , P3_R1054_U275;
wire P3_R1054_U276 , P3_R1054_U277 , P3_R1054_U278 , P3_R1054_U279 , P3_R1054_U280 , P3_R1054_U281 , P3_R1054_U282 , P3_R1054_U283 , P3_R1054_U284 , P3_R1054_U285;
wire P3_R1054_U286 , P3_R1054_U287 , P3_R1054_U288 , P3_R1054_U289 , P3_R1054_U290 , P3_R1054_U291 , P3_R1054_U292 , P3_R1054_U293 , P3_R1054_U294 , P3_R1161_U4;
wire P3_R1161_U5 , P3_R1161_U6 , P3_R1161_U7 , P3_R1161_U8 , P3_R1161_U9 , P3_R1161_U10 , P3_R1161_U11 , P3_R1161_U12 , P3_R1161_U13 , P3_R1161_U14;
wire P3_R1161_U15 , P3_R1161_U16 , P3_R1161_U17 , P3_R1161_U18 , P3_R1161_U19 , P3_R1161_U20 , P3_R1161_U21 , P3_R1161_U22 , P3_R1161_U23 , P3_R1161_U24;
wire P3_R1161_U25 , P3_R1161_U26 , P3_R1161_U27 , P3_R1161_U28 , P3_R1161_U29 , P3_R1161_U30 , P3_R1161_U31 , P3_R1161_U32 , P3_R1161_U33 , P3_R1161_U34;
wire P3_R1161_U35 , P3_R1161_U36 , P3_R1161_U37 , P3_R1161_U38 , P3_R1161_U39 , P3_R1161_U40 , P3_R1161_U41 , P3_R1161_U42 , P3_R1161_U43 , P3_R1161_U44;
wire P3_R1161_U45 , P3_R1161_U46 , P3_R1161_U47 , P3_R1161_U48 , P3_R1161_U49 , P3_R1161_U50 , P3_R1161_U51 , P3_R1161_U52 , P3_R1161_U53 , P3_R1161_U54;
wire P3_R1161_U55 , P3_R1161_U56 , P3_R1161_U57 , P3_R1161_U58 , P3_R1161_U59 , P3_R1161_U60 , P3_R1161_U61 , P3_R1161_U62 , P3_R1161_U63 , P3_R1161_U64;
wire P3_R1161_U65 , P3_R1161_U66 , P3_R1161_U67 , P3_R1161_U68 , P3_R1161_U69 , P3_R1161_U70 , P3_R1161_U71 , P3_R1161_U72 , P3_R1161_U73 , P3_R1161_U74;
wire P3_R1161_U75 , P3_R1161_U76 , P3_R1161_U77 , P3_R1161_U78 , P3_R1161_U79 , P3_R1161_U80 , P3_R1161_U81 , P3_R1161_U82 , P3_R1161_U83 , P3_R1161_U84;
wire P3_R1161_U85 , P3_R1161_U86 , P3_R1161_U87 , P3_R1161_U88 , P3_R1161_U89 , P3_R1161_U90 , P3_R1161_U91 , P3_R1161_U92 , P3_R1161_U93 , P3_R1161_U94;
wire P3_R1161_U95 , P3_R1161_U96 , P3_R1161_U97 , P3_R1161_U98 , P3_R1161_U99 , P3_R1161_U100 , P3_R1161_U101 , P3_R1161_U102 , P3_R1161_U103 , P3_R1161_U104;
wire P3_R1161_U105 , P3_R1161_U106 , P3_R1161_U107 , P3_R1161_U108 , P3_R1161_U109 , P3_R1161_U110 , P3_R1161_U111 , P3_R1161_U112 , P3_R1161_U113 , P3_R1161_U114;
wire P3_R1161_U115 , P3_R1161_U116 , P3_R1161_U117 , P3_R1161_U118 , P3_R1161_U119 , P3_R1161_U120 , P3_R1161_U121 , P3_R1161_U122 , P3_R1161_U123 , P3_R1161_U124;
wire P3_R1161_U125 , P3_R1161_U126 , P3_R1161_U127 , P3_R1161_U128 , P3_R1161_U129 , P3_R1161_U130 , P3_R1161_U131 , P3_R1161_U132 , P3_R1161_U133 , P3_R1161_U134;
wire P3_R1161_U135 , P3_R1161_U136 , P3_R1161_U137 , P3_R1161_U138 , P3_R1161_U139 , P3_R1161_U140 , P3_R1161_U141 , P3_R1161_U142 , P3_R1161_U143 , P3_R1161_U144;
wire P3_R1161_U145 , P3_R1161_U146 , P3_R1161_U147 , P3_R1161_U148 , P3_R1161_U149 , P3_R1161_U150 , P3_R1161_U151 , P3_R1161_U152 , P3_R1161_U153 , P3_R1161_U154;
wire P3_R1161_U155 , P3_R1161_U156 , P3_R1161_U157 , P3_R1161_U158 , P3_R1161_U159 , P3_R1161_U160 , P3_R1161_U161 , P3_R1161_U162 , P3_R1161_U163 , P3_R1161_U164;
wire P3_R1161_U165 , P3_R1161_U166 , P3_R1161_U167 , P3_R1161_U168 , P3_R1161_U169 , P3_R1161_U170 , P3_R1161_U171 , P3_R1161_U172 , P3_R1161_U173 , P3_R1161_U174;
wire P3_R1161_U175 , P3_R1161_U176 , P3_R1161_U177 , P3_R1161_U178 , P3_R1161_U179 , P3_R1161_U180 , P3_R1161_U181 , P3_R1161_U182 , P3_R1161_U183 , P3_R1161_U184;
wire P3_R1161_U185 , P3_R1161_U186 , P3_R1161_U187 , P3_R1161_U188 , P3_R1161_U189 , P3_R1161_U190 , P3_R1161_U191 , P3_R1161_U192 , P3_R1161_U193 , P3_R1161_U194;
wire P3_R1161_U195 , P3_R1161_U196 , P3_R1161_U197 , P3_R1161_U198 , P3_R1161_U199 , P3_R1161_U200 , P3_R1161_U201 , P3_R1161_U202 , P3_R1161_U203 , P3_R1161_U204;
wire P3_R1161_U205 , P3_R1161_U206 , P3_R1161_U207 , P3_R1161_U208 , P3_R1161_U209 , P3_R1161_U210 , P3_R1161_U211 , P3_R1161_U212 , P3_R1161_U213 , P3_R1161_U214;
wire P3_R1161_U215 , P3_R1161_U216 , P3_R1161_U217 , P3_R1161_U218 , P3_R1161_U219 , P3_R1161_U220 , P3_R1161_U221 , P3_R1161_U222 , P3_R1161_U223 , P3_R1161_U224;
wire P3_R1161_U225 , P3_R1161_U226 , P3_R1161_U227 , P3_R1161_U228 , P3_R1161_U229 , P3_R1161_U230 , P3_R1161_U231 , P3_R1161_U232 , P3_R1161_U233 , P3_R1161_U234;
wire P3_R1161_U235 , P3_R1161_U236 , P3_R1161_U237 , P3_R1161_U238 , P3_R1161_U239 , P3_R1161_U240 , P3_R1161_U241 , P3_R1161_U242 , P3_R1161_U243 , P3_R1161_U244;
wire P3_R1161_U245 , P3_R1161_U246 , P3_R1161_U247 , P3_R1161_U248 , P3_R1161_U249 , P3_R1161_U250 , P3_R1161_U251 , P3_R1161_U252 , P3_R1161_U253 , P3_R1161_U254;
wire P3_R1161_U255 , P3_R1161_U256 , P3_R1161_U257 , P3_R1161_U258 , P3_R1161_U259 , P3_R1161_U260 , P3_R1161_U261 , P3_R1161_U262 , P3_R1161_U263 , P3_R1161_U264;
wire P3_R1161_U265 , P3_R1161_U266 , P3_R1161_U267 , P3_R1161_U268 , P3_R1161_U269 , P3_R1161_U270 , P3_R1161_U271 , P3_R1161_U272 , P3_R1161_U273 , P3_R1161_U274;
wire P3_R1161_U275 , P3_R1161_U276 , P3_R1161_U277 , P3_R1161_U278 , P3_R1161_U279 , P3_R1161_U280 , P3_R1161_U281 , P3_R1161_U282 , P3_R1161_U283 , P3_R1161_U284;
wire P3_R1161_U285 , P3_R1161_U286 , P3_R1161_U287 , P3_R1161_U288 , P3_R1161_U289 , P3_R1161_U290 , P3_R1161_U291 , P3_R1161_U292 , P3_R1161_U293 , P3_R1161_U294;
wire P3_R1161_U295 , P3_R1161_U296 , P3_R1161_U297 , P3_R1161_U298 , P3_R1161_U299 , P3_R1161_U300 , P3_R1161_U301 , P3_R1161_U302 , P3_R1161_U303 , P3_R1161_U304;
wire P3_R1161_U305 , P3_R1161_U306 , P3_R1161_U307 , P3_R1161_U308 , P3_R1161_U309 , P3_R1161_U310 , P3_R1161_U311 , P3_R1161_U312 , P3_R1161_U313 , P3_R1161_U314;
wire P3_R1161_U315 , P3_R1161_U316 , P3_R1161_U317 , P3_R1161_U318 , P3_R1161_U319 , P3_R1161_U320 , P3_R1161_U321 , P3_R1161_U322 , P3_R1161_U323 , P3_R1161_U324;
wire P3_R1161_U325 , P3_R1161_U326 , P3_R1161_U327 , P3_R1161_U328 , P3_R1161_U329 , P3_R1161_U330 , P3_R1161_U331 , P3_R1161_U332 , P3_R1161_U333 , P3_R1161_U334;
wire P3_R1161_U335 , P3_R1161_U336 , P3_R1161_U337 , P3_R1161_U338 , P3_R1161_U339 , P3_R1161_U340 , P3_R1161_U341 , P3_R1161_U342 , P3_R1161_U343 , P3_R1161_U344;
wire P3_R1161_U345 , P3_R1161_U346 , P3_R1161_U347 , P3_R1161_U348 , P3_R1161_U349 , P3_R1161_U350 , P3_R1161_U351 , P3_R1161_U352 , P3_R1161_U353 , P3_R1161_U354;
wire P3_R1161_U355 , P3_R1161_U356 , P3_R1161_U357 , P3_R1161_U358 , P3_R1161_U359 , P3_R1161_U360 , P3_R1161_U361 , P3_R1161_U362 , P3_R1161_U363 , P3_R1161_U364;
wire P3_R1161_U365 , P3_R1161_U366 , P3_R1161_U367 , P3_R1161_U368 , P3_R1161_U369 , P3_R1161_U370 , P3_R1161_U371 , P3_R1161_U372 , P3_R1161_U373 , P3_R1161_U374;
wire P3_R1161_U375 , P3_R1161_U376 , P3_R1161_U377 , P3_R1161_U378 , P3_R1161_U379 , P3_R1161_U380 , P3_R1161_U381 , P3_R1161_U382 , P3_R1161_U383 , P3_R1161_U384;
wire P3_R1161_U385 , P3_R1161_U386 , P3_R1161_U387 , P3_R1161_U388 , P3_R1161_U389 , P3_R1161_U390 , P3_R1161_U391 , P3_R1161_U392 , P3_R1161_U393 , P3_R1161_U394;
wire P3_R1161_U395 , P3_R1161_U396 , P3_R1161_U397 , P3_R1161_U398 , P3_R1161_U399 , P3_R1161_U400 , P3_R1161_U401 , P3_R1161_U402 , P3_R1161_U403 , P3_R1161_U404;
wire P3_R1161_U405 , P3_R1161_U406 , P3_R1161_U407 , P3_R1161_U408 , P3_R1161_U409 , P3_R1161_U410 , P3_R1161_U411 , P3_R1161_U412 , P3_R1161_U413 , P3_R1161_U414;
wire P3_R1161_U415 , P3_R1161_U416 , P3_R1161_U417 , P3_R1161_U418 , P3_R1161_U419 , P3_R1161_U420 , P3_R1161_U421 , P3_R1161_U422 , P3_R1161_U423 , P3_R1161_U424;
wire P3_R1161_U425 , P3_R1161_U426 , P3_R1161_U427 , P3_R1161_U428 , P3_R1161_U429;


nand NAND2_1 ( P3_R1161_U504 , P3_U3387 , P3_R1161_U30 );
nand NAND2_2 ( P3_R1161_U503 , P3_U3076 , P3_R1161_U29 );
nand NAND2_3 ( P3_R1161_U502 , P3_U3419 , P3_R1161_U62 );
or OR2_4 ( U28 , P3_WR_REG , U160 );
or OR2_5 ( U29 , P3_RD_REG , U163 );
nand NAND2_6 ( U30 , U173 , U172 );
nand NAND2_7 ( U31 , U175 , U174 );
nand NAND2_8 ( U32 , U177 , U176 );
nand NAND2_9 ( U33 , U179 , U178 );
nand NAND2_10 ( U34 , U181 , U180 );
nand NAND2_11 ( U35 , U183 , U182 );
nand NAND2_12 ( U36 , U185 , U184 );
nand NAND2_13 ( U37 , U187 , U186 );
nand NAND2_14 ( U38 , U189 , U188 );
nand NAND2_15 ( U39 , U191 , U190 );
nand NAND2_16 ( U40 , U193 , U192 );
nand NAND2_17 ( U41 , U195 , U194 );
nand NAND2_18 ( U42 , U197 , U196 );
nand NAND2_19 ( U43 , U199 , U198 );
nand NAND2_20 ( U44 , U201 , U200 );
nand NAND2_21 ( U45 , U203 , U202 );
nand NAND2_22 ( U46 , U205 , U204 );
nand NAND2_23 ( U47 , U207 , U206 );
nand NAND2_24 ( U48 , U209 , U208 );
nand NAND2_25 ( U49 , U211 , U210 );
nand NAND2_26 ( U50 , U213 , U212 );
nand NAND2_27 ( U51 , U215 , U214 );
nand NAND2_28 ( U52 , U217 , U216 );
nand NAND2_29 ( U53 , U219 , U218 );
nand NAND2_30 ( U54 , U221 , U220 );
nand NAND2_31 ( U55 , U223 , U222 );
nand NAND2_32 ( U56 , U225 , U224 );
nand NAND2_33 ( U57 , U227 , U226 );
nand NAND2_34 ( U58 , U229 , U228 );
nand NAND2_35 ( U59 , U231 , U230 );
nand NAND2_36 ( U60 , U233 , U232 );
nand NAND2_37 ( U61 , U235 , U234 );
nand NAND2_38 ( U62 , U237 , U236 );
nand NAND2_39 ( U63 , U239 , U238 );
nand NAND2_40 ( U64 , U241 , U240 );
nand NAND2_41 ( U65 , U243 , U242 );
nand NAND2_42 ( U66 , U245 , U244 );
nand NAND2_43 ( U67 , U247 , U246 );
nand NAND2_44 ( U68 , U249 , U248 );
nand NAND2_45 ( U69 , U251 , U250 );
nand NAND2_46 ( U70 , U253 , U252 );
nand NAND2_47 ( U71 , U255 , U254 );
nand NAND2_48 ( U72 , U257 , U256 );
nand NAND2_49 ( U73 , U259 , U258 );
nand NAND2_50 ( U74 , U261 , U260 );
nand NAND2_51 ( U75 , U263 , U262 );
nand NAND2_52 ( U76 , U265 , U264 );
nand NAND2_53 ( U77 , U267 , U266 );
nand NAND2_54 ( U78 , U269 , U268 );
nand NAND2_55 ( U79 , U271 , U270 );
nand NAND2_56 ( U80 , U273 , U272 );
nand NAND2_57 ( U81 , U275 , U274 );
nand NAND2_58 ( U82 , U277 , U276 );
nand NAND2_59 ( U83 , U279 , U278 );
nand NAND2_60 ( U84 , U281 , U280 );
nand NAND2_61 ( U85 , U283 , U282 );
nand NAND2_62 ( U86 , U285 , U284 );
nand NAND2_63 ( U87 , U287 , U286 );
nand NAND2_64 ( U88 , U289 , U288 );
nand NAND2_65 ( U89 , U291 , U290 );
nand NAND2_66 ( U90 , U293 , U292 );
nand NAND2_67 ( U91 , U295 , U294 );
nand NAND2_68 ( U92 , U297 , U296 );
nand NAND2_69 ( U93 , U299 , U298 );
nand NAND2_70 ( U94 , U301 , U300 );
nand NAND2_71 ( U95 , U303 , U302 );
nand NAND2_72 ( U96 , U305 , U304 );
nand NAND2_73 ( U97 , U307 , U306 );
nand NAND2_74 ( U98 , U309 , U308 );
nand NAND2_75 ( U99 , U311 , U310 );
nand NAND2_76 ( U100 , U313 , U312 );
nand NAND2_77 ( U101 , U315 , U314 );
nand NAND2_78 ( U102 , U317 , U316 );
nand NAND2_79 ( U103 , U319 , U318 );
nand NAND2_80 ( U104 , U321 , U320 );
nand NAND2_81 ( U105 , U323 , U322 );
nand NAND2_82 ( U106 , U325 , U324 );
nand NAND2_83 ( U107 , U327 , U326 );
nand NAND2_84 ( U108 , U329 , U328 );
nand NAND2_85 ( U109 , U331 , U330 );
nand NAND2_86 ( U110 , U333 , U332 );
nand NAND2_87 ( U111 , U335 , U334 );
nand NAND2_88 ( U112 , U337 , U336 );
nand NAND2_89 ( U113 , U339 , U338 );
nand NAND2_90 ( U114 , U341 , U340 );
nand NAND2_91 ( U115 , U343 , U342 );
nand NAND2_92 ( U116 , U345 , U344 );
nand NAND2_93 ( U117 , U347 , U346 );
nand NAND2_94 ( U118 , U349 , U348 );
nand NAND2_95 ( U119 , U351 , U350 );
nand NAND2_96 ( U120 , U353 , U352 );
nand NAND2_97 ( U121 , U355 , U354 );
nand NAND2_98 ( U122 , U357 , U356 );
nand NAND2_99 ( U123 , U359 , U358 );
nand NAND2_100 ( U124 , U361 , U360 );
nand NAND2_101 ( U125 , U363 , U362 );
nand NAND2_102 ( U126 , U365 , U364 );
nand NAND2_103 ( U127 , U367 , U366 );
nand NAND2_104 ( U128 , U369 , U368 );
nand NAND2_105 ( U129 , U371 , U370 );
nand NAND2_106 ( U130 , U373 , U372 );
nand NAND2_107 ( U131 , U375 , U374 );
nand NAND2_108 ( U132 , U377 , U376 );
nand NAND2_109 ( U133 , U379 , U378 );
nand NAND2_110 ( U134 , U381 , U380 );
nand NAND2_111 ( U135 , U383 , U382 );
nand NAND2_112 ( U136 , U385 , U384 );
nand NAND2_113 ( U137 , U387 , U386 );
nand NAND2_114 ( U138 , U389 , U388 );
nand NAND2_115 ( U139 , U391 , U390 );
nand NAND2_116 ( U140 , U393 , U392 );
nand NAND2_117 ( U141 , U395 , U394 );
nand NAND2_118 ( U142 , U397 , U396 );
nand NAND2_119 ( U143 , U399 , U398 );
nand NAND2_120 ( U144 , U401 , U400 );
nand NAND2_121 ( U145 , U403 , U402 );
nand NAND2_122 ( U146 , U405 , U404 );
nand NAND2_123 ( U147 , U407 , U406 );
nand NAND2_124 ( U148 , U409 , U408 );
nand NAND2_125 ( U149 , U411 , U410 );
nand NAND2_126 ( U150 , U413 , U412 );
nand NAND2_127 ( U151 , U415 , U414 );
nand NAND2_128 ( U152 , U417 , U416 );
nand NAND2_129 ( U153 , U419 , U418 );
nand NAND2_130 ( U154 , U421 , U420 );
nand NAND2_131 ( U155 , U423 , U422 );
nand NAND2_132 ( U156 , U425 , U424 );
nand NAND2_133 ( U157 , U427 , U426 );
not NOT1_134 ( U158 , P2_WR_REG );
not NOT1_135 ( U159 , P1_WR_REG );
and AND2_136 ( U160 , U169 , U168 );
not NOT1_137 ( U161 , P2_RD_REG );
not NOT1_138 ( U162 , P1_RD_REG );
and AND2_139 ( U163 , U171 , U170 );
nand NAND2_140 ( U164 , U166 , U165 );
nand NAND4_141 ( U165 , P1_ADDR_REG_19_ , P2_ADDR_REG_19_ , LT_1602_U6 , U161 );
nand NAND4_142 ( U166 , LT_1601_U6 , LT_1601_21_U6 , P3_ADDR_REG_19_ , U162 );
not NOT1_143 ( U167 , U164 );
nand NAND2_144 ( U168 , P2_WR_REG , U159 );
nand NAND2_145 ( U169 , P1_WR_REG , U158 );
nand NAND2_146 ( U170 , P2_RD_REG , U162 );
nand NAND2_147 ( U171 , P1_RD_REG , U161 );
nand NAND2_148 ( U172 , SUB_1605_U79 , U164 );
nand NAND2_149 ( U173 , SI_9_ , U167 );
nand NAND2_150 ( U174 , SUB_1605_U80 , U164 );
nand NAND2_151 ( U175 , SI_8_ , U167 );
nand NAND2_152 ( U176 , SUB_1605_U81 , U164 );
nand NAND2_153 ( U177 , SI_7_ , U167 );
nand NAND2_154 ( U178 , SUB_1605_U82 , U164 );
nand NAND2_155 ( U179 , SI_6_ , U167 );
nand NAND2_156 ( U180 , SUB_1605_U83 , U164 );
nand NAND2_157 ( U181 , SI_5_ , U167 );
nand NAND2_158 ( U182 , SUB_1605_U84 , U164 );
nand NAND2_159 ( U183 , SI_4_ , U167 );
nand NAND2_160 ( U184 , SUB_1605_U85 , U164 );
nand NAND2_161 ( U185 , SI_3_ , U167 );
nand NAND2_162 ( U186 , SUB_1605_U12 , U164 );
nand NAND2_163 ( U187 , SI_31_ , U167 );
nand NAND2_164 ( U188 , SUB_1605_U86 , U164 );
nand NAND2_165 ( U189 , SI_30_ , U167 );
nand NAND2_166 ( U190 , SUB_1605_U87 , U164 );
nand NAND2_167 ( U191 , SI_2_ , U167 );
nand NAND2_168 ( U192 , SUB_1605_U88 , U164 );
nand NAND2_169 ( U193 , SI_29_ , U167 );
nand NAND2_170 ( U194 , SUB_1605_U89 , U164 );
nand NAND2_171 ( U195 , SI_28_ , U167 );
nand NAND2_172 ( U196 , SUB_1605_U90 , U164 );
nand NAND2_173 ( U197 , SI_27_ , U167 );
nand NAND2_174 ( U198 , SUB_1605_U91 , U164 );
nand NAND2_175 ( U199 , SI_26_ , U167 );
nand NAND2_176 ( U200 , SUB_1605_U92 , U164 );
nand NAND2_177 ( U201 , SI_25_ , U167 );
nand NAND2_178 ( U202 , SUB_1605_U93 , U164 );
nand NAND2_179 ( U203 , SI_24_ , U167 );
nand NAND2_180 ( U204 , SUB_1605_U94 , U164 );
nand NAND2_181 ( U205 , SI_23_ , U167 );
nand NAND2_182 ( U206 , SUB_1605_U95 , U164 );
nand NAND2_183 ( U207 , SI_22_ , U167 );
nand NAND2_184 ( U208 , SUB_1605_U96 , U164 );
nand NAND2_185 ( U209 , SI_21_ , U167 );
nand NAND2_186 ( U210 , SUB_1605_U97 , U164 );
nand NAND2_187 ( U211 , SI_20_ , U167 );
nand NAND2_188 ( U212 , SUB_1605_U98 , U164 );
nand NAND2_189 ( U213 , SI_1_ , U167 );
nand NAND2_190 ( U214 , SUB_1605_U99 , U164 );
nand NAND2_191 ( U215 , SI_19_ , U167 );
nand NAND2_192 ( U216 , SUB_1605_U100 , U164 );
nand NAND2_193 ( U217 , SI_18_ , U167 );
nand NAND2_194 ( U218 , SUB_1605_U101 , U164 );
nand NAND2_195 ( U219 , SI_17_ , U167 );
nand NAND2_196 ( U220 , SUB_1605_U102 , U164 );
nand NAND2_197 ( U221 , SI_16_ , U167 );
nand NAND2_198 ( U222 , SUB_1605_U103 , U164 );
nand NAND2_199 ( U223 , SI_15_ , U167 );
nand NAND2_200 ( U224 , SUB_1605_U104 , U164 );
nand NAND2_201 ( U225 , SI_14_ , U167 );
nand NAND2_202 ( U226 , SUB_1605_U105 , U164 );
nand NAND2_203 ( U227 , SI_13_ , U167 );
nand NAND2_204 ( U228 , SUB_1605_U106 , U164 );
nand NAND2_205 ( U229 , SI_12_ , U167 );
nand NAND2_206 ( U230 , SUB_1605_U107 , U164 );
nand NAND2_207 ( U231 , SI_11_ , U167 );
nand NAND2_208 ( U232 , SUB_1605_U108 , U164 );
nand NAND2_209 ( U233 , SI_10_ , U167 );
nand NAND2_210 ( U234 , SUB_1605_U13 , U164 );
nand NAND2_211 ( U235 , SI_0_ , U167 );
nand NAND2_212 ( U236 , P1_DATAO_REG_9_ , U164 );
nand NAND2_213 ( U237 , R152_U85 , U167 );
nand NAND2_214 ( U238 , P1_DATAO_REG_8_ , U164 );
nand NAND2_215 ( U239 , R152_U86 , U167 );
nand NAND2_216 ( U240 , P1_DATAO_REG_7_ , U164 );
nand NAND2_217 ( U241 , R152_U87 , U167 );
nand NAND2_218 ( U242 , P1_DATAO_REG_6_ , U164 );
nand NAND2_219 ( U243 , R152_U88 , U167 );
nand NAND2_220 ( U244 , P1_DATAO_REG_5_ , U164 );
nand NAND2_221 ( U245 , R152_U89 , U167 );
nand NAND2_222 ( U246 , P1_DATAO_REG_4_ , U164 );
nand NAND2_223 ( U247 , R152_U90 , U167 );
nand NAND2_224 ( U248 , P1_DATAO_REG_3_ , U164 );
nand NAND2_225 ( U249 , R152_U91 , U167 );
nand NAND2_226 ( U250 , P1_DATAO_REG_31_ , U164 );
nand NAND2_227 ( U251 , R152_U12 , U167 );
nand NAND2_228 ( U252 , P1_DATAO_REG_30_ , U164 );
nand NAND2_229 ( U253 , R152_U92 , U167 );
nand NAND2_230 ( U254 , P1_DATAO_REG_2_ , U164 );
nand NAND2_231 ( U255 , R152_U93 , U167 );
nand NAND2_232 ( U256 , P1_DATAO_REG_29_ , U164 );
nand NAND2_233 ( U257 , R152_U94 , U167 );
nand NAND2_234 ( U258 , P1_DATAO_REG_28_ , U164 );
nand NAND2_235 ( U259 , R152_U95 , U167 );
nand NAND2_236 ( U260 , P1_DATAO_REG_27_ , U164 );
nand NAND2_237 ( U261 , R152_U96 , U167 );
nand NAND2_238 ( U262 , P1_DATAO_REG_26_ , U164 );
nand NAND2_239 ( U263 , R152_U97 , U167 );
nand NAND2_240 ( U264 , P1_DATAO_REG_25_ , U164 );
nand NAND2_241 ( U265 , R152_U98 , U167 );
nand NAND2_242 ( U266 , P1_DATAO_REG_24_ , U164 );
nand NAND2_243 ( U267 , R152_U99 , U167 );
nand NAND2_244 ( U268 , P1_DATAO_REG_23_ , U164 );
nand NAND2_245 ( U269 , R152_U100 , U167 );
nand NAND2_246 ( U270 , P1_DATAO_REG_22_ , U164 );
nand NAND2_247 ( U271 , R152_U101 , U167 );
nand NAND2_248 ( U272 , P1_DATAO_REG_21_ , U164 );
nand NAND2_249 ( U273 , R152_U102 , U167 );
nand NAND2_250 ( U274 , P1_DATAO_REG_20_ , U164 );
nand NAND2_251 ( U275 , R152_U103 , U167 );
nand NAND2_252 ( U276 , P1_DATAO_REG_1_ , U164 );
nand NAND2_253 ( U277 , R152_U13 , U167 );
nand NAND2_254 ( U278 , P1_DATAO_REG_19_ , U164 );
nand NAND2_255 ( U279 , R152_U104 , U167 );
nand NAND2_256 ( U280 , P1_DATAO_REG_18_ , U164 );
nand NAND2_257 ( U281 , R152_U105 , U167 );
nand NAND2_258 ( U282 , P1_DATAO_REG_17_ , U164 );
nand NAND2_259 ( U283 , R152_U106 , U167 );
nand NAND2_260 ( U284 , P1_DATAO_REG_16_ , U164 );
nand NAND2_261 ( U285 , R152_U107 , U167 );
nand NAND2_262 ( U286 , P1_DATAO_REG_15_ , U164 );
nand NAND2_263 ( U287 , R152_U108 , U167 );
nand NAND2_264 ( U288 , P1_DATAO_REG_14_ , U164 );
nand NAND2_265 ( U289 , R152_U109 , U167 );
nand NAND2_266 ( U290 , P1_DATAO_REG_13_ , U164 );
nand NAND2_267 ( U291 , R152_U110 , U167 );
nand NAND2_268 ( U292 , P1_DATAO_REG_12_ , U164 );
nand NAND2_269 ( U293 , R152_U111 , U167 );
nand NAND2_270 ( U294 , P1_DATAO_REG_11_ , U164 );
nand NAND2_271 ( U295 , R152_U112 , U167 );
nand NAND2_272 ( U296 , P1_DATAO_REG_10_ , U164 );
nand NAND2_273 ( U297 , R152_U113 , U167 );
nand NAND2_274 ( U298 , P1_DATAO_REG_0_ , U164 );
nand NAND2_275 ( U299 , R152_U84 , U167 );
nand NAND2_276 ( U300 , R152_U85 , U164 );
nand NAND2_277 ( U301 , P2_DATAO_REG_9_ , U167 );
nand NAND2_278 ( U302 , R152_U86 , U164 );
nand NAND2_279 ( U303 , P2_DATAO_REG_8_ , U167 );
nand NAND2_280 ( U304 , R152_U87 , U164 );
nand NAND2_281 ( U305 , P2_DATAO_REG_7_ , U167 );
nand NAND2_282 ( U306 , R152_U88 , U164 );
nand NAND2_283 ( U307 , P2_DATAO_REG_6_ , U167 );
nand NAND2_284 ( U308 , R152_U89 , U164 );
nand NAND2_285 ( U309 , P2_DATAO_REG_5_ , U167 );
nand NAND2_286 ( U310 , R152_U90 , U164 );
nand NAND2_287 ( U311 , P2_DATAO_REG_4_ , U167 );
nand NAND2_288 ( U312 , R152_U91 , U164 );
nand NAND2_289 ( U313 , P2_DATAO_REG_3_ , U167 );
nand NAND2_290 ( U314 , R152_U12 , U164 );
nand NAND2_291 ( U315 , P2_DATAO_REG_31_ , U167 );
nand NAND2_292 ( U316 , R152_U92 , U164 );
nand NAND2_293 ( U317 , P2_DATAO_REG_30_ , U167 );
nand NAND2_294 ( U318 , R152_U93 , U164 );
nand NAND2_295 ( U319 , P2_DATAO_REG_2_ , U167 );
nand NAND2_296 ( U320 , R152_U94 , U164 );
nand NAND2_297 ( U321 , P2_DATAO_REG_29_ , U167 );
nand NAND2_298 ( U322 , R152_U95 , U164 );
nand NAND2_299 ( U323 , P2_DATAO_REG_28_ , U167 );
nand NAND2_300 ( U324 , R152_U96 , U164 );
nand NAND2_301 ( U325 , P2_DATAO_REG_27_ , U167 );
nand NAND2_302 ( U326 , R152_U97 , U164 );
nand NAND2_303 ( U327 , P2_DATAO_REG_26_ , U167 );
nand NAND2_304 ( U328 , R152_U98 , U164 );
nand NAND2_305 ( U329 , P2_DATAO_REG_25_ , U167 );
nand NAND2_306 ( U330 , R152_U99 , U164 );
nand NAND2_307 ( U331 , P2_DATAO_REG_24_ , U167 );
nand NAND2_308 ( U332 , R152_U100 , U164 );
nand NAND2_309 ( U333 , P2_DATAO_REG_23_ , U167 );
nand NAND2_310 ( U334 , R152_U101 , U164 );
nand NAND2_311 ( U335 , P2_DATAO_REG_22_ , U167 );
nand NAND2_312 ( U336 , R152_U102 , U164 );
nand NAND2_313 ( U337 , P2_DATAO_REG_21_ , U167 );
nand NAND2_314 ( U338 , R152_U103 , U164 );
nand NAND2_315 ( U339 , P2_DATAO_REG_20_ , U167 );
nand NAND2_316 ( U340 , R152_U13 , U164 );
nand NAND2_317 ( U341 , P2_DATAO_REG_1_ , U167 );
nand NAND2_318 ( U342 , R152_U104 , U164 );
nand NAND2_319 ( U343 , P2_DATAO_REG_19_ , U167 );
nand NAND2_320 ( U344 , R152_U105 , U164 );
nand NAND2_321 ( U345 , P2_DATAO_REG_18_ , U167 );
nand NAND2_322 ( U346 , R152_U106 , U164 );
nand NAND2_323 ( U347 , P2_DATAO_REG_17_ , U167 );
nand NAND2_324 ( U348 , R152_U107 , U164 );
nand NAND2_325 ( U349 , P2_DATAO_REG_16_ , U167 );
nand NAND2_326 ( U350 , R152_U108 , U164 );
nand NAND2_327 ( U351 , P2_DATAO_REG_15_ , U167 );
nand NAND2_328 ( U352 , R152_U109 , U164 );
nand NAND2_329 ( U353 , P2_DATAO_REG_14_ , U167 );
nand NAND2_330 ( U354 , R152_U110 , U164 );
nand NAND2_331 ( U355 , P2_DATAO_REG_13_ , U167 );
nand NAND2_332 ( U356 , R152_U111 , U164 );
nand NAND2_333 ( U357 , P2_DATAO_REG_12_ , U167 );
nand NAND2_334 ( U358 , R152_U112 , U164 );
nand NAND2_335 ( U359 , P2_DATAO_REG_11_ , U167 );
nand NAND2_336 ( U360 , R152_U113 , U164 );
nand NAND2_337 ( U361 , P2_DATAO_REG_10_ , U167 );
nand NAND2_338 ( U362 , R152_U84 , U164 );
nand NAND2_339 ( U363 , P2_DATAO_REG_0_ , U167 );
nand NAND2_340 ( U364 , P2_DATAO_REG_9_ , U164 );
nand NAND2_341 ( U365 , P1_DATAO_REG_9_ , U167 );
nand NAND2_342 ( U366 , P2_DATAO_REG_8_ , U164 );
nand NAND2_343 ( U367 , P1_DATAO_REG_8_ , U167 );
nand NAND2_344 ( U368 , P2_DATAO_REG_7_ , U164 );
nand NAND2_345 ( U369 , P1_DATAO_REG_7_ , U167 );
nand NAND2_346 ( U370 , P2_DATAO_REG_6_ , U164 );
nand NAND2_347 ( U371 , P1_DATAO_REG_6_ , U167 );
nand NAND2_348 ( U372 , P2_DATAO_REG_5_ , U164 );
nand NAND2_349 ( U373 , P1_DATAO_REG_5_ , U167 );
nand NAND2_350 ( U374 , P2_DATAO_REG_4_ , U164 );
nand NAND2_351 ( U375 , P1_DATAO_REG_4_ , U167 );
nand NAND2_352 ( U376 , P2_DATAO_REG_31_ , U164 );
nand NAND2_353 ( U377 , P1_DATAO_REG_31_ , U167 );
nand NAND2_354 ( U378 , P2_DATAO_REG_30_ , U164 );
nand NAND2_355 ( U379 , P1_DATAO_REG_30_ , U167 );
nand NAND2_356 ( U380 , P2_DATAO_REG_3_ , U164 );
nand NAND2_357 ( U381 , P1_DATAO_REG_3_ , U167 );
nand NAND2_358 ( U382 , P2_DATAO_REG_29_ , U164 );
nand NAND2_359 ( U383 , P1_DATAO_REG_29_ , U167 );
nand NAND2_360 ( U384 , P2_DATAO_REG_28_ , U164 );
nand NAND2_361 ( U385 , P1_DATAO_REG_28_ , U167 );
nand NAND2_362 ( U386 , P2_DATAO_REG_27_ , U164 );
nand NAND2_363 ( U387 , P1_DATAO_REG_27_ , U167 );
nand NAND2_364 ( U388 , P2_DATAO_REG_26_ , U164 );
nand NAND2_365 ( U389 , P1_DATAO_REG_26_ , U167 );
nand NAND2_366 ( U390 , P2_DATAO_REG_25_ , U164 );
nand NAND2_367 ( U391 , P1_DATAO_REG_25_ , U167 );
nand NAND2_368 ( U392 , P2_DATAO_REG_24_ , U164 );
nand NAND2_369 ( U393 , P1_DATAO_REG_24_ , U167 );
nand NAND2_370 ( U394 , P2_DATAO_REG_23_ , U164 );
nand NAND2_371 ( U395 , P1_DATAO_REG_23_ , U167 );
nand NAND2_372 ( U396 , P2_DATAO_REG_22_ , U164 );
nand NAND2_373 ( U397 , P1_DATAO_REG_22_ , U167 );
nand NAND2_374 ( U398 , P2_DATAO_REG_21_ , U164 );
nand NAND2_375 ( U399 , P1_DATAO_REG_21_ , U167 );
nand NAND2_376 ( U400 , P2_DATAO_REG_20_ , U164 );
nand NAND2_377 ( U401 , P1_DATAO_REG_20_ , U167 );
nand NAND2_378 ( U402 , P2_DATAO_REG_2_ , U164 );
nand NAND2_379 ( U403 , P1_DATAO_REG_2_ , U167 );
nand NAND2_380 ( U404 , P2_DATAO_REG_19_ , U164 );
nand NAND2_381 ( U405 , P1_DATAO_REG_19_ , U167 );
nand NAND2_382 ( U406 , P2_DATAO_REG_18_ , U164 );
nand NAND2_383 ( U407 , P1_DATAO_REG_18_ , U167 );
nand NAND2_384 ( U408 , P2_DATAO_REG_17_ , U164 );
nand NAND2_385 ( U409 , P1_DATAO_REG_17_ , U167 );
nand NAND2_386 ( U410 , P2_DATAO_REG_16_ , U164 );
nand NAND2_387 ( U411 , P1_DATAO_REG_16_ , U167 );
nand NAND2_388 ( U412 , P2_DATAO_REG_15_ , U164 );
nand NAND2_389 ( U413 , P1_DATAO_REG_15_ , U167 );
nand NAND2_390 ( U414 , P2_DATAO_REG_14_ , U164 );
nand NAND2_391 ( U415 , P1_DATAO_REG_14_ , U167 );
nand NAND2_392 ( U416 , P2_DATAO_REG_13_ , U164 );
nand NAND2_393 ( U417 , P1_DATAO_REG_13_ , U167 );
nand NAND2_394 ( U418 , P2_DATAO_REG_12_ , U164 );
nand NAND2_395 ( U419 , P1_DATAO_REG_12_ , U167 );
nand NAND2_396 ( U420 , P2_DATAO_REG_11_ , U164 );
nand NAND2_397 ( U421 , P1_DATAO_REG_11_ , U167 );
nand NAND2_398 ( U422 , P2_DATAO_REG_10_ , U164 );
nand NAND2_399 ( U423 , P1_DATAO_REG_10_ , U167 );
nand NAND2_400 ( U424 , P2_DATAO_REG_1_ , U164 );
nand NAND2_401 ( U425 , P1_DATAO_REG_1_ , U167 );
nand NAND2_402 ( U426 , P2_DATAO_REG_0_ , U164 );
nand NAND2_403 ( U427 , P1_DATAO_REG_0_ , U167 );
nand NAND2_404 ( P3_R1161_U501 , P3_U3061 , P3_R1161_U61 );
nand NAND2_405 ( P3_R1161_U500 , P3_R1161_U244 , P3_R1161_U498 );
nand NAND2_406 ( P3_R1161_U499 , P3_R1161_U363 , P3_R1161_U167 );
nand NAND2_407 ( P3_R1161_U498 , P3_R1161_U497 , P3_R1161_U496 );
nand NAND2_408 ( P3_R1161_U497 , P3_U3422 , P3_R1161_U67 );
nand NAND2_409 ( P3_R1161_U496 , P3_U3062 , P3_R1161_U66 );
nand NAND2_410 ( P3_R1161_U495 , P3_R1161_U493 , P3_R1161_U338 );
nand NAND2_411 ( P3_R1161_U494 , P3_R1161_U362 , P3_R1161_U93 );
nand NAND2_412 ( P3_R1161_U493 , P3_R1161_U492 , P3_R1161_U491 );
nand NAND2_413 ( P3_R1161_U492 , P3_U3425 , P3_R1161_U65 );
nand NAND2_414 ( P3_R1161_U491 , P3_U3071 , P3_R1161_U64 );
nand NAND2_415 ( P3_R1161_U490 , P3_U3428 , P3_R1161_U70 );
and AND2_416 ( P1_U3014 , P1_U4002 , P1_U3451 );
and AND2_417 ( P1_U3015 , P1_U3455 , P1_U3449 );
and AND2_418 ( P1_U3016 , P1_U3605 , P1_U3600 );
and AND2_419 ( P1_U3017 , P1_U3447 , P1_U3448 );
and AND2_420 ( P1_U3018 , P1_U5808 , P1_U3447 );
and AND2_421 ( P1_U3019 , P1_U5805 , P1_U3448 );
and AND2_422 ( P1_U3020 , P1_U5805 , P1_U5808 );
and AND2_423 ( P1_U3021 , P1_U5412 , P1_U3425 );
and AND2_424 ( P1_U3022 , P1_U3592 , P1_U3425 );
and AND2_425 ( P1_U3023 , P1_U4043 , P1_U3428 );
and AND2_426 ( P1_U3024 , P1_U3048 , P1_U5793 );
and AND2_427 ( P1_U3025 , P1_U4030 , P1_U5811 );
and AND2_428 ( P1_U3026 , P1_U3851 , P1_U4015 );
and AND2_429 ( P1_U3027 , P1_R1352_U6 , P1_U3437 );
and AND2_430 ( P1_U3028 , P1_R1352_U6 , P1_U3440 );
and AND2_431 ( P1_U3029 , P1_U3357 , P1_STATE_REG );
and AND2_432 ( P1_U3030 , P1_U4008 , P1_U4031 );
and AND2_433 ( P1_U3031 , P1_U4031 , P1_U3426 );
and AND2_434 ( P1_U3032 , P1_U4003 , P1_U4031 );
and AND2_435 ( P1_U3033 , P1_U4009 , P1_U4031 );
and AND2_436 ( P1_U3034 , P1_U4030 , P1_U3449 );
and AND2_437 ( P1_U3035 , P1_U4015 , P1_U5811 );
and AND2_438 ( P1_U3036 , P1_U4031 , P1_U3025 );
and AND2_439 ( P1_U3037 , P1_U4015 , P1_U3449 );
and AND2_440 ( P1_U3038 , P1_U5817 , P1_U4923 );
and AND2_441 ( P1_U3039 , P1_U3023 , P1_U5817 );
and AND2_442 ( P1_U3040 , P1_U5811 , P1_U4923 );
and AND2_443 ( P1_U3041 , P1_U3023 , P1_U5811 );
and AND2_444 ( P1_U3042 , P1_U3015 , P1_U4923 );
and AND2_445 ( P1_U3043 , P1_U3023 , P1_U3015 );
and AND2_446 ( P1_U3044 , P1_U3022 , P1_U3428 );
and AND2_447 ( P1_U3045 , P1_U3022 , P1_U5159 );
and AND2_448 ( P1_U3046 , P1_U3606 , P1_U3016 );
and AND2_449 ( P1_U3047 , P1_U3452 , P1_U3453 );
and AND2_450 ( P1_U3048 , P1_U5799 , P1_U3452 );
and AND2_451 ( P1_U3049 , P1_U5802 , P1_U5796 );
and AND2_452 ( P1_U3050 , P1_U3850 , P1_U5148 );
and AND2_453 ( P1_U3051 , P1_U3419 , P1_U3367 );
and AND3_454 ( P1_U3052 , P1_U5541 , P1_U3422 , P1_U3879 );
nand NAND4_455 ( P1_U3053 , P1_U4680 , P1_U4681 , P1_U4679 , P1_U4682 );
nand NAND4_456 ( P1_U3054 , P1_U4699 , P1_U4700 , P1_U4698 , P1_U4701 );
nand NAND4_457 ( P1_U3055 , P1_U4720 , P1_U4719 , P1_U4718 , P1_U4717 );
nand NAND3_458 ( P1_U3056 , P1_U4757 , P1_U4758 , P1_U4756 );
nand NAND4_459 ( P1_U3057 , P1_U4661 , P1_U4662 , P1_U4660 , P1_U4663 );
nand NAND4_460 ( P1_U3058 , P1_U4642 , P1_U4643 , P1_U4641 , P1_U4644 );
nand NAND3_461 ( P1_U3059 , P1_U4737 , P1_U4738 , P1_U4736 );
nand NAND4_462 ( P1_U3060 , P1_U4245 , P1_U4244 , P1_U4243 , P1_U4242 );
nand NAND4_463 ( P1_U3061 , P1_U4585 , P1_U4586 , P1_U4584 , P1_U4587 );
nand NAND4_464 ( P1_U3062 , P1_U4357 , P1_U4358 , P1_U4356 , P1_U4359 );
nand NAND4_465 ( P1_U3063 , P1_U4376 , P1_U4377 , P1_U4375 , P1_U4378 );
nand NAND4_466 ( P1_U3064 , P1_U4226 , P1_U4225 , P1_U4224 , P1_U4223 );
nand NAND4_467 ( P1_U3065 , P1_U4623 , P1_U4624 , P1_U4622 , P1_U4625 );
nand NAND4_468 ( P1_U3066 , P1_U4604 , P1_U4605 , P1_U4603 , P1_U4606 );
nand NAND4_469 ( P1_U3067 , P1_U4264 , P1_U4263 , P1_U4262 , P1_U4261 );
nand NAND4_470 ( P1_U3068 , P1_U4202 , P1_U4201 , P1_U4200 , P1_U4199 );
nand NAND4_471 ( P1_U3069 , P1_U4490 , P1_U4491 , P1_U4489 , P1_U4492 );
nand NAND4_472 ( P1_U3070 , P1_U4302 , P1_U4301 , P1_U4300 , P1_U4299 );
nand NAND4_473 ( P1_U3071 , P1_U4283 , P1_U4282 , P1_U4281 , P1_U4280 );
nand NAND4_474 ( P1_U3072 , P1_U4395 , P1_U4396 , P1_U4394 , P1_U4397 );
nand NAND4_475 ( P1_U3073 , P1_U4471 , P1_U4472 , P1_U4470 , P1_U4473 );
nand NAND4_476 ( P1_U3074 , P1_U4452 , P1_U4453 , P1_U4451 , P1_U4454 );
nand NAND4_477 ( P1_U3075 , P1_U4566 , P1_U4567 , P1_U4565 , P1_U4568 );
nand NAND4_478 ( P1_U3076 , P1_U4547 , P1_U4548 , P1_U4546 , P1_U4549 );
nand NAND4_479 ( P1_U3077 , P1_U4207 , P1_U4206 , P1_U4205 , P1_U4204 );
nand NAND4_480 ( P1_U3078 , P1_U4183 , P1_U4182 , P1_U4181 , P1_U4180 );
nand NAND4_481 ( P1_U3079 , P1_U4433 , P1_U4434 , P1_U4432 , P1_U4435 );
nand NAND4_482 ( P1_U3080 , P1_U4414 , P1_U4415 , P1_U4413 , P1_U4416 );
nand NAND4_483 ( P1_U3081 , P1_U4528 , P1_U4529 , P1_U4527 , P1_U4530 );
nand NAND4_484 ( P1_U3082 , P1_U4509 , P1_U4510 , P1_U4508 , P1_U4511 );
nand NAND4_485 ( P1_U3083 , P1_U4338 , P1_U4339 , P1_U4337 , P1_U4340 );
nand NAND4_486 ( P1_U3084 , P1_U4321 , P1_U4320 , P1_U4319 , P1_U4318 );
nand NAND2_487 ( P1_U3085 , P1_U4930 , P1_STATE_REG );
not NOT1_488 ( P1_U3086 , P1_STATE_REG );
nand NAND3_489 ( P1_U3087 , P1_U5668 , P1_U5666 , P1_U5667 );
nand NAND3_490 ( P1_U3088 , P1_U5671 , P1_U5669 , P1_U5670 );
nand NAND3_491 ( P1_U3089 , P1_U3929 , P1_U5678 , P1_U5679 );
nand NAND3_492 ( P1_U3090 , P1_U5683 , P1_U5682 , P1_U3930 );
nand NAND3_493 ( P1_U3091 , P1_U5687 , P1_U5686 , P1_U3931 );
nand NAND3_494 ( P1_U3092 , P1_U5691 , P1_U5690 , P1_U3932 );
nand NAND3_495 ( P1_U3093 , P1_U5695 , P1_U5694 , P1_U3933 );
nand NAND3_496 ( P1_U3094 , P1_U5699 , P1_U5698 , P1_U3934 );
nand NAND3_497 ( P1_U3095 , P1_U5703 , P1_U5702 , P1_U3935 );
nand NAND3_498 ( P1_U3096 , P1_U5707 , P1_U5706 , P1_U3936 );
nand NAND3_499 ( P1_U3097 , P1_U5711 , P1_U5710 , P1_U3937 );
nand NAND3_500 ( P1_U3098 , P1_U5715 , P1_U5714 , P1_U3938 );
nand NAND3_501 ( P1_U3099 , P1_U5723 , P1_U5722 , P1_U3940 );
nand NAND3_502 ( P1_U3100 , P1_U5727 , P1_U5726 , P1_U3941 );
nand NAND3_503 ( P1_U3101 , P1_U5731 , P1_U5730 , P1_U3942 );
nand NAND3_504 ( P1_U3102 , P1_U5735 , P1_U5734 , P1_U3943 );
nand NAND3_505 ( P1_U3103 , P1_U5739 , P1_U5738 , P1_U3944 );
nand NAND3_506 ( P1_U3104 , P1_U5743 , P1_U5742 , P1_U3945 );
nand NAND3_507 ( P1_U3105 , P1_U5747 , P1_U5746 , P1_U3946 );
nand NAND3_508 ( P1_U3106 , P1_U5751 , P1_U5750 , P1_U3947 );
nand NAND3_509 ( P1_U3107 , P1_U5755 , P1_U5754 , P1_U3948 );
nand NAND3_510 ( P1_U3108 , P1_U5759 , P1_U5758 , P1_U3949 );
nand NAND3_511 ( P1_U3109 , P1_U3922 , P1_U5644 , P1_U5643 );
nand NAND3_512 ( P1_U3110 , P1_U3923 , P1_U5648 , P1_U5647 );
nand NAND3_513 ( P1_U3111 , P1_U5653 , P1_U5652 , P1_U3924 );
nand NAND3_514 ( P1_U3112 , P1_U5657 , P1_U5656 , P1_U3925 );
nand NAND3_515 ( P1_U3113 , P1_U5661 , P1_U5660 , P1_U3926 );
nand NAND3_516 ( P1_U3114 , P1_U5665 , P1_U5664 , P1_U3927 );
nand NAND2_517 ( P1_U3115 , P1_U3928 , P1_U5674 );
nand NAND2_518 ( P1_U3116 , P1_U3939 , P1_U5718 );
nand NAND2_519 ( P1_U3117 , P1_U3950 , P1_U5762 );
nand NAND2_520 ( P1_U3118 , P1_U3951 , P1_U5766 );
nand NAND2_521 ( P1_U3119 , P1_U3892 , P1_U5563 );
nand NAND2_522 ( P1_U3120 , P1_U3893 , P1_U5566 );
nand NAND3_523 ( P1_U3121 , P1_U5572 , P1_U5571 , P1_U3896 );
nand NAND3_524 ( P1_U3122 , P1_U5575 , P1_U5574 , P1_U3897 );
nand NAND3_525 ( P1_U3123 , P1_U5578 , P1_U5577 , P1_U3898 );
nand NAND3_526 ( P1_U3124 , P1_U5581 , P1_U5580 , P1_U3899 );
nand NAND3_527 ( P1_U3125 , P1_U5584 , P1_U5583 , P1_U3900 );
nand NAND3_528 ( P1_U3126 , P1_U5587 , P1_U5586 , P1_U3901 );
nand NAND3_529 ( P1_U3127 , P1_U5590 , P1_U5589 , P1_U3902 );
nand NAND3_530 ( P1_U3128 , P1_U5593 , P1_U5592 , P1_U3903 );
nand NAND3_531 ( P1_U3129 , P1_U5596 , P1_U5595 , P1_U3904 );
nand NAND3_532 ( P1_U3130 , P1_U5599 , P1_U5598 , P1_U3905 );
nand NAND3_533 ( P1_U3131 , P1_U5605 , P1_U5604 , P1_U3908 );
nand NAND3_534 ( P1_U3132 , P1_U5608 , P1_U5607 , P1_U3909 );
nand NAND3_535 ( P1_U3133 , P1_U5611 , P1_U5610 , P1_U3910 );
nand NAND3_536 ( P1_U3134 , P1_U5614 , P1_U5613 , P1_U3911 );
nand NAND3_537 ( P1_U3135 , P1_U5617 , P1_U5616 , P1_U3912 );
nand NAND3_538 ( P1_U3136 , P1_U5620 , P1_U5619 , P1_U3913 );
nand NAND3_539 ( P1_U3137 , P1_U5623 , P1_U5622 , P1_U3914 );
nand NAND3_540 ( P1_U3138 , P1_U5626 , P1_U5625 , P1_U3915 );
nand NAND3_541 ( P1_U3139 , P1_U5629 , P1_U5628 , P1_U3916 );
nand NAND3_542 ( P1_U3140 , P1_U5632 , P1_U5631 , P1_U3917 );
nand NAND2_543 ( P1_U3141 , P1_U5545 , P1_U3880 );
nand NAND2_544 ( P1_U3142 , P1_U5548 , P1_U3882 );
nand NAND2_545 ( P1_U3143 , P1_U5551 , P1_U3884 );
nand NAND2_546 ( P1_U3144 , P1_U5554 , P1_U3886 );
nand NAND2_547 ( P1_U3145 , P1_U5557 , P1_U3888 );
nand NAND2_548 ( P1_U3146 , P1_U5560 , P1_U3890 );
nand NAND2_549 ( P1_U3147 , P1_U5569 , P1_U3894 );
nand NAND2_550 ( P1_U3148 , P1_U5602 , P1_U3906 );
nand NAND2_551 ( P1_U3149 , P1_U5635 , P1_U3918 );
nand NAND2_552 ( P1_U3150 , P1_U5638 , P1_U3920 );
nand NAND2_553 ( P1_U3151 , P1_U3877 , P1_U5537 );
nand NAND2_554 ( P1_U3152 , P1_U3014 , P1_U5786 );
nand NAND2_555 ( P1_U3153 , P1_U5492 , P1_U5491 );
nand NAND2_556 ( P1_U3154 , P1_U5494 , P1_U5493 );
nand NAND2_557 ( P1_U3155 , P1_U5496 , P1_U5495 );
nand NAND2_558 ( P1_U3156 , P1_U5498 , P1_U5497 );
nand NAND2_559 ( P1_U3157 , P1_U5500 , P1_U5499 );
nand NAND2_560 ( P1_U3158 , P1_U5502 , P1_U5501 );
nand NAND2_561 ( P1_U3159 , P1_U5504 , P1_U5503 );
nand NAND2_562 ( P1_U3160 , P1_U5506 , P1_U5505 );
nand NAND2_563 ( P1_U3161 , P1_U5508 , P1_U5507 );
nand NAND2_564 ( P1_U3162 , P1_U5512 , P1_U5511 );
nand NAND2_565 ( P1_U3163 , P1_U5514 , P1_U5513 );
nand NAND2_566 ( P1_U3164 , P1_U5516 , P1_U5515 );
nand NAND2_567 ( P1_U3165 , P1_U5518 , P1_U5517 );
nand NAND2_568 ( P1_U3166 , P1_U5520 , P1_U5519 );
nand NAND2_569 ( P1_U3167 , P1_U5522 , P1_U5521 );
nand NAND2_570 ( P1_U3168 , P1_U5524 , P1_U5523 );
nand NAND2_571 ( P1_U3169 , P1_U5526 , P1_U5525 );
nand NAND2_572 ( P1_U3170 , P1_U5528 , P1_U5527 );
nand NAND2_573 ( P1_U3171 , P1_U5530 , P1_U5529 );
nand NAND2_574 ( P1_U3172 , P1_U5478 , P1_U5477 );
nand NAND2_575 ( P1_U3173 , P1_U5480 , P1_U5479 );
nand NAND2_576 ( P1_U3174 , P1_U5482 , P1_U5481 );
nand NAND2_577 ( P1_U3175 , P1_U5484 , P1_U5483 );
nand NAND2_578 ( P1_U3176 , P1_U5486 , P1_U5485 );
nand NAND2_579 ( P1_U3177 , P1_U5488 , P1_U5487 );
nand NAND2_580 ( P1_U3178 , P1_U5490 , P1_U5489 );
nand NAND2_581 ( P1_U3179 , P1_U5510 , P1_U5509 );
nand NAND2_582 ( P1_U3180 , P1_U5532 , P1_U5531 );
nand NAND2_583 ( P1_U3181 , P1_U3876 , P1_U5534 );
nand NAND2_584 ( P1_U3182 , P1_U5433 , P1_U5432 );
nand NAND2_585 ( P1_U3183 , P1_U5435 , P1_U5434 );
nand NAND2_586 ( P1_U3184 , P1_U5437 , P1_U5436 );
nand NAND2_587 ( P1_U3185 , P1_U5439 , P1_U5438 );
nand NAND2_588 ( P1_U3186 , P1_U5441 , P1_U5440 );
nand NAND2_589 ( P1_U3187 , P1_U5443 , P1_U5442 );
nand NAND2_590 ( P1_U3188 , P1_U5445 , P1_U5444 );
nand NAND2_591 ( P1_U3189 , P1_U5447 , P1_U5446 );
nand NAND2_592 ( P1_U3190 , P1_U5449 , P1_U5448 );
nand NAND2_593 ( P1_U3191 , P1_U5453 , P1_U5452 );
nand NAND2_594 ( P1_U3192 , P1_U5455 , P1_U5454 );
nand NAND2_595 ( P1_U3193 , P1_U5457 , P1_U5456 );
nand NAND2_596 ( P1_U3194 , P1_U5459 , P1_U5458 );
nand NAND2_597 ( P1_U3195 , P1_U5461 , P1_U5460 );
nand NAND2_598 ( P1_U3196 , P1_U5463 , P1_U5462 );
nand NAND2_599 ( P1_U3197 , P1_U5465 , P1_U5464 );
nand NAND2_600 ( P1_U3198 , P1_U5467 , P1_U5466 );
nand NAND2_601 ( P1_U3199 , P1_U5469 , P1_U5468 );
nand NAND2_602 ( P1_U3200 , P1_U5471 , P1_U5470 );
nand NAND2_603 ( P1_U3201 , P1_U5419 , P1_U5418 );
nand NAND2_604 ( P1_U3202 , P1_U5421 , P1_U5420 );
nand NAND2_605 ( P1_U3203 , P1_U5423 , P1_U5422 );
nand NAND2_606 ( P1_U3204 , P1_U5425 , P1_U5424 );
nand NAND2_607 ( P1_U3205 , P1_U5427 , P1_U5426 );
nand NAND2_608 ( P1_U3206 , P1_U5429 , P1_U5428 );
nand NAND2_609 ( P1_U3207 , P1_U5431 , P1_U5430 );
nand NAND2_610 ( P1_U3208 , P1_U5451 , P1_U5450 );
nand NAND2_611 ( P1_U3209 , P1_U5473 , P1_U5472 );
nand NAND2_612 ( P1_U3210 , P1_U3875 , P1_U5474 );
and AND2_613 ( P1_U3211 , P1_U5411 , P1_U3425 );
nand NAND3_614 ( P1_U3212 , P1_U6285 , P1_U6284 , P1_U5409 );
nand NAND4_615 ( P1_U3213 , P1_U5403 , P1_U5402 , P1_U3872 , P1_U5404 );
nand NAND5_616 ( P1_U3214 , P1_U5394 , P1_U5393 , P1_U5397 , P1_U5396 , P1_U5395 );
nand NAND5_617 ( P1_U3215 , P1_U5385 , P1_U5384 , P1_U5388 , P1_U5387 , P1_U5386 );
nand NAND5_618 ( P1_U3216 , P1_U5376 , P1_U5375 , P1_U5379 , P1_U5378 , P1_U5377 );
nand NAND4_619 ( P1_U3217 , P1_U5367 , P1_U5366 , P1_U3871 , P1_U5368 );
nand NAND3_620 ( P1_U3218 , P1_U3869 , P1_U5358 , P1_U3870 );
nand NAND5_621 ( P1_U3219 , P1_U5349 , P1_U5348 , P1_U5352 , P1_U5351 , P1_U5350 );
nand NAND5_622 ( P1_U3220 , P1_U5340 , P1_U5339 , P1_U5343 , P1_U5342 , P1_U5341 );
nand NAND4_623 ( P1_U3221 , P1_U5331 , P1_U5330 , P1_U3868 , P1_U5332 );
nand NAND3_624 ( P1_U3222 , P1_U3866 , P1_U5322 , P1_U3867 );
nand NAND5_625 ( P1_U3223 , P1_U5313 , P1_U5312 , P1_U5316 , P1_U5315 , P1_U5314 );
nand NAND4_626 ( P1_U3224 , P1_U5304 , P1_U5303 , P1_U3865 , P1_U5305 );
nand NAND5_627 ( P1_U3225 , P1_U5295 , P1_U5294 , P1_U5298 , P1_U5297 , P1_U5296 );
nand NAND5_628 ( P1_U3226 , P1_U5286 , P1_U5285 , P1_U5289 , P1_U5288 , P1_U5287 );
nand NAND4_629 ( P1_U3227 , P1_U5277 , P1_U5276 , P1_U5278 , P1_U3864 );
nand NAND5_630 ( P1_U3228 , P1_U5268 , P1_U5267 , P1_U5271 , P1_U5270 , P1_U5269 );
nand NAND5_631 ( P1_U3229 , P1_U5259 , P1_U5258 , P1_U5262 , P1_U5261 , P1_U5260 );
nand NAND3_632 ( P1_U3230 , P1_U3862 , P1_U5250 , P1_U3863 );
nand NAND4_633 ( P1_U3231 , P1_U5241 , P1_U5240 , P1_U3861 , P1_U5242 );
nand NAND2_634 ( P1_U3232 , P1_U5233 , P1_U3859 );
nand NAND5_635 ( P1_U3233 , P1_U5224 , P1_U5223 , P1_U5227 , P1_U5226 , P1_U5225 );
nand NAND4_636 ( P1_U3234 , P1_U5215 , P1_U5214 , P1_U3857 , P1_U5216 );
nand NAND5_637 ( P1_U3235 , P1_U5206 , P1_U5205 , P1_U5209 , P1_U5208 , P1_U5207 );
nand NAND4_638 ( P1_U3236 , P1_U5197 , P1_U5196 , P1_U3856 , P1_U5198 );
nand NAND3_639 ( P1_U3237 , P1_U3854 , P1_U5188 , P1_U3855 );
nand NAND5_640 ( P1_U3238 , P1_U5179 , P1_U5178 , P1_U5182 , P1_U5181 , P1_U5180 );
nand NAND4_641 ( P1_U3239 , P1_U5170 , P1_U5169 , P1_U3853 , P1_U5171 );
nand NAND5_642 ( P1_U3240 , P1_U5161 , P1_U5160 , P1_U5164 , P1_U5163 , P1_U5162 );
nand NAND5_643 ( P1_U3241 , P1_U5150 , P1_U5149 , P1_U5153 , P1_U5152 , P1_U5151 );
nand NAND2_644 ( P1_U3242 , P1_U3846 , P1_U5137 );
nand NAND3_645 ( P1_U3243 , P1_U3830 , P1_U5123 , P1_U3831 );
nand NAND3_646 ( P1_U3244 , P1_U3828 , P1_U5113 , P1_U3829 );
nand NAND3_647 ( P1_U3245 , P1_U5103 , P1_U3825 , P1_U3827 );
nand NAND3_648 ( P1_U3246 , P1_U3823 , P1_U5093 , P1_U3824 );
nand NAND3_649 ( P1_U3247 , P1_U5083 , P1_U3820 , P1_U3822 );
nand NAND3_650 ( P1_U3248 , P1_U3818 , P1_U5073 , P1_U3819 );
nand NAND3_651 ( P1_U3249 , P1_U3816 , P1_U3817 , P1_U5063 );
nand NAND3_652 ( P1_U3250 , P1_U3814 , P1_U3815 , P1_U5053 );
nand NAND3_653 ( P1_U3251 , P1_U3812 , P1_U3813 , P1_U5043 );
nand NAND3_654 ( P1_U3252 , P1_U3810 , P1_U3811 , P1_U5033 );
nand NAND3_655 ( P1_U3253 , P1_U3808 , P1_U3809 , P1_U5023 );
nand NAND3_656 ( P1_U3254 , P1_U3806 , P1_U3807 , P1_U5013 );
nand NAND3_657 ( P1_U3255 , P1_U3804 , P1_U3805 , P1_U5003 );
nand NAND3_658 ( P1_U3256 , P1_U3802 , P1_U3803 , P1_U4993 );
nand NAND3_659 ( P1_U3257 , P1_U3800 , P1_U3801 , P1_U4983 );
nand NAND3_660 ( P1_U3258 , P1_U3798 , P1_U3799 , P1_U4973 );
nand NAND3_661 ( P1_U3259 , P1_U3796 , P1_U3797 , P1_U4963 );
nand NAND3_662 ( P1_U3260 , P1_U3794 , P1_U3795 , P1_U4953 );
nand NAND3_663 ( P1_U3261 , P1_U3792 , P1_U3793 , P1_U4943 );
nand NAND3_664 ( P1_U3262 , P1_U3790 , P1_U3791 , P1_U4933 );
nand NAND3_665 ( P1_U3263 , P1_U3989 , P1_U4921 , P1_U4922 );
nand NAND3_666 ( P1_U3264 , P1_U3988 , P1_U4919 , P1_U4920 );
nand NAND4_667 ( P1_U3265 , P1_U3784 , P1_U3785 , P1_U4912 , P1_U3985 );
nand NAND4_668 ( P1_U3266 , P1_U3782 , P1_U3783 , P1_U4907 , P1_U3984 );
nand NAND4_669 ( P1_U3267 , P1_U3780 , P1_U3781 , P1_U4902 , P1_U3983 );
nand NAND4_670 ( P1_U3268 , P1_U3778 , P1_U3779 , P1_U4897 , P1_U3982 );
nand NAND4_671 ( P1_U3269 , P1_U3776 , P1_U3777 , P1_U4892 , P1_U3981 );
nand NAND4_672 ( P1_U3270 , P1_U3774 , P1_U3775 , P1_U4887 , P1_U3980 );
nand NAND4_673 ( P1_U3271 , P1_U3772 , P1_U3773 , P1_U4882 , P1_U3979 );
nand NAND4_674 ( P1_U3272 , P1_U3770 , P1_U3771 , P1_U4877 , P1_U3978 );
nand NAND4_675 ( P1_U3273 , P1_U3768 , P1_U3769 , P1_U4872 , P1_U3977 );
nand NAND4_676 ( P1_U3274 , P1_U3766 , P1_U3767 , P1_U4867 , P1_U3976 );
nand NAND3_677 ( P1_U3275 , P1_U3765 , P1_U3764 , P1_U3975 );
nand NAND3_678 ( P1_U3276 , P1_U3763 , P1_U3762 , P1_U3974 );
nand NAND4_679 ( P1_U3277 , P1_U3760 , P1_U3761 , P1_U4852 , P1_U3973 );
nand NAND4_680 ( P1_U3278 , P1_U3758 , P1_U3759 , P1_U4847 , P1_U3972 );
nand NAND3_681 ( P1_U3279 , P1_U3757 , P1_U3756 , P1_U3971 );
nand NAND3_682 ( P1_U3280 , P1_U3755 , P1_U3754 , P1_U3970 );
nand NAND3_683 ( P1_U3281 , P1_U3753 , P1_U3752 , P1_U3969 );
nand NAND3_684 ( P1_U3282 , P1_U3751 , P1_U3750 , P1_U3968 );
nand NAND4_685 ( P1_U3283 , P1_U3748 , P1_U3749 , P1_U4822 , P1_U3967 );
nand NAND4_686 ( P1_U3284 , P1_U3746 , P1_U3747 , P1_U4817 , P1_U3966 );
nand NAND3_687 ( P1_U3285 , P1_U3745 , P1_U3744 , P1_U3965 );
nand NAND3_688 ( P1_U3286 , P1_U3743 , P1_U3742 , P1_U3964 );
nand NAND3_689 ( P1_U3287 , P1_U3741 , P1_U3740 , P1_U3963 );
nand NAND3_690 ( P1_U3288 , P1_U3739 , P1_U3738 , P1_U3962 );
nand NAND2_691 ( P1_U3289 , P1_U3737 , P1_U3736 );
nand NAND2_692 ( P1_U3290 , P1_U3735 , P1_U3734 );
nand NAND2_693 ( P1_U3291 , P1_U3733 , P1_U3732 );
nand NAND2_694 ( P1_U3292 , P1_U3731 , P1_U3730 );
nand NAND2_695 ( P1_U3293 , P1_U3729 , P1_U3728 );
and AND2_696 ( P1_U3294 , P1_D_REG_31_ , P1_U3953 );
and AND2_697 ( P1_U3295 , P1_D_REG_30_ , P1_U3953 );
and AND2_698 ( P1_U3296 , P1_D_REG_29_ , P1_U3953 );
and AND2_699 ( P1_U3297 , P1_D_REG_28_ , P1_U3953 );
and AND2_700 ( P1_U3298 , P1_D_REG_27_ , P1_U3953 );
and AND2_701 ( P1_U3299 , P1_D_REG_26_ , P1_U3953 );
and AND2_702 ( P1_U3300 , P1_D_REG_25_ , P1_U3953 );
and AND2_703 ( P1_U3301 , P1_D_REG_24_ , P1_U3953 );
and AND2_704 ( P1_U3302 , P1_D_REG_23_ , P1_U3953 );
and AND2_705 ( P1_U3303 , P1_D_REG_22_ , P1_U3953 );
and AND2_706 ( P1_U3304 , P1_D_REG_21_ , P1_U3953 );
and AND2_707 ( P1_U3305 , P1_D_REG_20_ , P1_U3953 );
and AND2_708 ( P1_U3306 , P1_D_REG_19_ , P1_U3953 );
and AND2_709 ( P1_U3307 , P1_D_REG_18_ , P1_U3953 );
and AND2_710 ( P1_U3308 , P1_D_REG_17_ , P1_U3953 );
and AND2_711 ( P1_U3309 , P1_D_REG_16_ , P1_U3953 );
and AND2_712 ( P1_U3310 , P1_D_REG_15_ , P1_U3953 );
and AND2_713 ( P1_U3311 , P1_D_REG_14_ , P1_U3953 );
and AND2_714 ( P1_U3312 , P1_D_REG_13_ , P1_U3953 );
and AND2_715 ( P1_U3313 , P1_D_REG_12_ , P1_U3953 );
and AND2_716 ( P1_U3314 , P1_D_REG_11_ , P1_U3953 );
and AND2_717 ( P1_U3315 , P1_D_REG_10_ , P1_U3953 );
and AND2_718 ( P1_U3316 , P1_D_REG_9_ , P1_U3953 );
and AND2_719 ( P1_U3317 , P1_D_REG_8_ , P1_U3953 );
and AND2_720 ( P1_U3318 , P1_D_REG_7_ , P1_U3953 );
and AND2_721 ( P1_U3319 , P1_D_REG_6_ , P1_U3953 );
and AND2_722 ( P1_U3320 , P1_D_REG_5_ , P1_U3953 );
and AND2_723 ( P1_U3321 , P1_D_REG_4_ , P1_U3953 );
and AND2_724 ( P1_U3322 , P1_D_REG_3_ , P1_U3953 );
and AND2_725 ( P1_U3323 , P1_D_REG_2_ , P1_U3953 );
nand NAND3_726 ( P1_U3324 , P1_U4142 , P1_U4143 , P1_U4141 );
nand NAND3_727 ( P1_U3325 , P1_U4139 , P1_U4140 , P1_U4138 );
nand NAND3_728 ( P1_U3326 , P1_U4136 , P1_U4137 , P1_U4135 );
nand NAND3_729 ( P1_U3327 , P1_U4133 , P1_U4134 , P1_U4132 );
nand NAND3_730 ( P1_U3328 , P1_U4130 , P1_U4131 , P1_U4129 );
nand NAND3_731 ( P1_U3329 , P1_U4127 , P1_U4128 , P1_U4126 );
nand NAND3_732 ( P1_U3330 , P1_U4124 , P1_U4125 , P1_U4123 );
nand NAND3_733 ( P1_U3331 , P1_U4121 , P1_U4122 , P1_U4120 );
nand NAND3_734 ( P1_U3332 , P1_U4118 , P1_U4119 , P1_U4117 );
nand NAND3_735 ( P1_U3333 , P1_U4115 , P1_U4116 , P1_U4114 );
nand NAND3_736 ( P1_U3334 , P1_U4112 , P1_U4113 , P1_U4111 );
nand NAND3_737 ( P1_U3335 , P1_U4109 , P1_U4110 , P1_U4108 );
nand NAND3_738 ( P1_U3336 , P1_U4106 , P1_U4107 , P1_U4105 );
nand NAND3_739 ( P1_U3337 , P1_U4103 , P1_U4104 , P1_U4102 );
nand NAND3_740 ( P1_U3338 , P1_U4100 , P1_U4101 , P1_U4099 );
nand NAND3_741 ( P1_U3339 , P1_U4097 , P1_U4098 , P1_U4096 );
nand NAND3_742 ( P1_U3340 , P1_U4094 , P1_U4095 , P1_U4093 );
nand NAND3_743 ( P1_U3341 , P1_U4091 , P1_U4092 , P1_U4090 );
nand NAND3_744 ( P1_U3342 , P1_U4088 , P1_U4089 , P1_U4087 );
nand NAND3_745 ( P1_U3343 , P1_U4085 , P1_U4086 , P1_U4084 );
nand NAND3_746 ( P1_U3344 , P1_U4082 , P1_U4083 , P1_U4081 );
nand NAND3_747 ( P1_U3345 , P1_U4079 , P1_U4080 , P1_U4078 );
nand NAND3_748 ( P1_U3346 , P1_U4076 , P1_U4077 , P1_U4075 );
nand NAND3_749 ( P1_U3347 , P1_U4073 , P1_U4074 , P1_U4072 );
nand NAND3_750 ( P1_U3348 , P1_U4070 , P1_U4071 , P1_U4069 );
nand NAND3_751 ( P1_U3349 , P1_U4067 , P1_U4068 , P1_U4066 );
nand NAND3_752 ( P1_U3350 , P1_U4064 , P1_U4065 , P1_U4063 );
nand NAND3_753 ( P1_U3351 , P1_U4061 , P1_U4062 , P1_U4060 );
nand NAND3_754 ( P1_U3352 , P1_U4058 , P1_U4059 , P1_U4057 );
nand NAND3_755 ( P1_U3353 , P1_U4055 , P1_U4056 , P1_U4054 );
nand NAND3_756 ( P1_U3354 , P1_U4052 , P1_U4053 , P1_U4051 );
nand NAND3_757 ( P1_U3355 , P1_U4049 , P1_U4050 , P1_U4048 );
nand NAND5_758 ( P1_U3356 , P1_U4917 , P1_U4915 , P1_U4918 , P1_U4916 , P1_U3986 );
nand NAND2_759 ( P1_U3357 , P1_STATE_REG , P1_U3952 );
nand NAND2_760 ( P1_U3358 , P1_U3443 , P1_U5778 );
not NOT1_761 ( P1_U3359 , P1_B_REG );
nand NAND3_762 ( P1_U3360 , P1_U5783 , P1_U5782 , P1_U3443 );
nand NAND2_763 ( P1_U3361 , P1_U3048 , P1_U3451 );
nand NAND2_764 ( P1_U3362 , P1_U3047 , P1_U3451 );
nand NAND2_765 ( P1_U3363 , P1_U3453 , P1_U5796 );
nand NAND2_766 ( P1_U3364 , P1_U4042 , P1_U3451 );
nand NAND2_767 ( P1_U3365 , P1_U3047 , P1_U3450 );
nand NAND2_768 ( P1_U3366 , P1_U4042 , P1_U3450 );
nand NAND2_769 ( P1_U3367 , P1_U3049 , P1_U3451 );
nand NAND2_770 ( P1_U3368 , P1_U4001 , P1_U5799 );
nand NAND2_771 ( P1_U3369 , P1_U5799 , P1_U5796 );
nand NAND2_772 ( P1_U3370 , P1_U4044 , P1_U3450 );
nand NAND2_773 ( P1_U3371 , P1_U4002 , P1_U5793 );
nand NAND2_774 ( P1_U3372 , P1_U3451 , P1_U3450 );
nand NAND3_775 ( P1_U3373 , P1_U5799 , P1_U5793 , P1_U5802 );
nand NAND2_776 ( P1_U3374 , P1_U3049 , P1_U5793 );
nand NAND2_777 ( P1_U3375 , P1_U5802 , P1_U3452 );
nand NAND5_778 ( P1_U3376 , P1_U4191 , P1_U4190 , P1_U4192 , P1_U3594 , P1_U3593 );
not NOT1_779 ( P1_U3377 , P1_REG2_REG_0_ );
nand NAND4_780 ( P1_U3378 , P1_U4210 , P1_U4209 , P1_U3608 , P1_U3610 );
nand NAND4_781 ( P1_U3379 , P1_U4229 , P1_U4228 , P1_U3612 , P1_U3614 );
nand NAND4_782 ( P1_U3380 , P1_U4248 , P1_U4247 , P1_U3616 , P1_U3618 );
nand NAND4_783 ( P1_U3381 , P1_U4267 , P1_U4266 , P1_U3620 , P1_U3622 );
nand NAND4_784 ( P1_U3382 , P1_U4286 , P1_U4285 , P1_U3624 , P1_U3626 );
nand NAND4_785 ( P1_U3383 , P1_U4305 , P1_U4304 , P1_U3628 , P1_U3630 );
nand NAND4_786 ( P1_U3384 , P1_U4324 , P1_U4323 , P1_U3632 , P1_U3634 );
nand NAND4_787 ( P1_U3385 , P1_U4343 , P1_U4342 , P1_U3636 , P1_U3638 );
nand NAND4_788 ( P1_U3386 , P1_U4362 , P1_U4361 , P1_U3640 , P1_U3642 );
nand NAND4_789 ( P1_U3387 , P1_U4381 , P1_U4380 , P1_U3644 , P1_U3646 );
nand NAND4_790 ( P1_U3388 , P1_U4400 , P1_U4399 , P1_U3648 , P1_U3650 );
nand NAND4_791 ( P1_U3389 , P1_U4419 , P1_U4418 , P1_U3652 , P1_U3654 );
nand NAND4_792 ( P1_U3390 , P1_U4438 , P1_U4437 , P1_U3656 , P1_U3658 );
nand NAND4_793 ( P1_U3391 , P1_U4457 , P1_U4456 , P1_U3660 , P1_U3662 );
nand NAND4_794 ( P1_U3392 , P1_U4476 , P1_U4475 , P1_U3664 , P1_U3666 );
nand NAND4_795 ( P1_U3393 , P1_U4495 , P1_U4494 , P1_U3668 , P1_U3670 );
nand NAND4_796 ( P1_U3394 , P1_U4514 , P1_U4513 , P1_U3672 , P1_U3674 );
nand NAND4_797 ( P1_U3395 , P1_U4533 , P1_U4532 , P1_U3676 , P1_U3678 );
nand NAND4_798 ( P1_U3396 , P1_U4552 , P1_U4551 , P1_U3680 , P1_U3682 );
nand NAND2_799 ( P1_U3397 , U113 , P1_U3954 );
nand NAND4_800 ( P1_U3398 , P1_U4571 , P1_U4570 , P1_U3684 , P1_U3686 );
nand NAND2_801 ( P1_U3399 , U112 , P1_U3954 );
nand NAND4_802 ( P1_U3400 , P1_U4590 , P1_U4589 , P1_U3688 , P1_U3690 );
nand NAND2_803 ( P1_U3401 , U111 , P1_U3954 );
nand NAND4_804 ( P1_U3402 , P1_U4609 , P1_U4608 , P1_U3692 , P1_U3694 );
nand NAND2_805 ( P1_U3403 , U110 , P1_U3954 );
nand NAND4_806 ( P1_U3404 , P1_U4628 , P1_U4627 , P1_U3696 , P1_U3698 );
nand NAND2_807 ( P1_U3405 , U109 , P1_U3954 );
nand NAND4_808 ( P1_U3406 , P1_U4647 , P1_U4646 , P1_U3700 , P1_U3702 );
nand NAND2_809 ( P1_U3407 , U108 , P1_U3954 );
nand NAND4_810 ( P1_U3408 , P1_U4666 , P1_U4665 , P1_U3704 , P1_U3706 );
nand NAND2_811 ( P1_U3409 , U107 , P1_U3954 );
nand NAND4_812 ( P1_U3410 , P1_U4685 , P1_U4684 , P1_U3708 , P1_U3710 );
nand NAND2_813 ( P1_U3411 , U106 , P1_U3954 );
nand NAND4_814 ( P1_U3412 , P1_U4704 , P1_U4703 , P1_U3712 , P1_U3714 );
nand NAND2_815 ( P1_U3413 , U105 , P1_U3954 );
nand NAND4_816 ( P1_U3414 , P1_U4723 , P1_U4722 , P1_U3716 , P1_U3718 );
nand NAND2_817 ( P1_U3415 , U104 , P1_U3954 );
nand NAND2_818 ( P1_U3416 , P1_U3723 , P1_U3721 );
nand NAND2_819 ( P1_U3417 , U102 , P1_U3954 );
nand NAND2_820 ( P1_U3418 , U101 , P1_U3954 );
nand NAND2_821 ( P1_U3419 , P1_U4041 , P1_U5793 );
nand NAND2_822 ( P1_U3420 , P1_U3022 , P1_U4767 );
nand NAND2_823 ( P1_U3421 , P1_U3998 , P1_U5799 );
nand NAND2_824 ( P1_U3422 , P1_U3048 , P1_U3450 );
nand NAND2_825 ( P1_U3423 , P1_U3047 , P1_U5793 );
nand NAND2_826 ( P1_U3424 , P1_U3993 , P1_U5799 );
nand NAND3_827 ( P1_U3425 , P1_U3441 , P1_U3443 , P1_U3442 );
nand NAND2_828 ( P1_U3426 , P1_U4010 , P1_U4768 );
nand NAND2_829 ( P1_U3427 , P1_U3444 , P1_STATE_REG );
nand NAND2_830 ( P1_U3428 , P1_U3429 , P1_U4931 );
nand NAND2_831 ( P1_U3429 , P1_U4145 , P1_U5786 );
nand NAND2_832 ( P1_U3430 , P1_U4045 , P1_STATE_REG );
nand NAND2_833 ( P1_U3431 , P1_U3014 , P1_U3015 );
not NOT1_834 ( P1_U3432 , P1_R1375_U9 );
nand NAND2_835 ( P1_U3433 , P1_U3022 , P1_U3426 );
nand NAND2_836 ( P1_U3434 , P1_U3847 , P1_U3016 );
nand NAND2_837 ( P1_U3435 , P1_U3852 , P1_U5143 );
nand NAND2_838 ( P1_U3436 , P1_U5415 , P1_U5414 );
nand NAND2_839 ( P1_U3437 , P1_U3999 , P1_U3362 );
nand NAND2_840 ( P1_U3438 , P1_U5536 , P1_U3051 );
not NOT1_841 ( P1_U3439 , P1_R1352_U6 );
nand NAND2_842 ( P1_U3440 , P1_U3364 , P1_U3423 );
nand NAND2_843 ( P1_U3441 , P1_U5774 , P1_U5773 );
nand NAND2_844 ( P1_U3442 , P1_U5777 , P1_U5776 );
nand NAND2_845 ( P1_U3443 , P1_U5780 , P1_U5779 );
nand NAND2_846 ( P1_U3444 , P1_U5785 , P1_U5784 );
nand NAND2_847 ( P1_U3445 , P1_U5788 , P1_U5787 );
nand NAND2_848 ( P1_U3446 , P1_U5790 , P1_U5789 );
nand NAND2_849 ( P1_U3447 , P1_U5804 , P1_U5803 );
nand NAND2_850 ( P1_U3448 , P1_U5807 , P1_U5806 );
nand NAND2_851 ( P1_U3449 , P1_U5810 , P1_U5809 );
nand NAND2_852 ( P1_U3450 , P1_U5801 , P1_U5800 );
nand NAND2_853 ( P1_U3451 , P1_U5792 , P1_U5791 );
nand NAND2_854 ( P1_U3452 , P1_U5795 , P1_U5794 );
nand NAND2_855 ( P1_U3453 , P1_U5798 , P1_U5797 );
nand NAND2_856 ( P1_U3454 , P1_U5813 , P1_U5812 );
nand NAND2_857 ( P1_U3455 , P1_U5816 , P1_U5815 );
nand NAND2_858 ( P1_U3456 , P1_U5819 , P1_U5818 );
nand NAND2_859 ( P1_U3457 , P1_U5827 , P1_U5826 );
nand NAND2_860 ( P1_U3458 , P1_U5824 , P1_U5823 );
nand NAND2_861 ( P1_U3459 , P1_U5830 , P1_U5829 );
nand NAND2_862 ( P1_U3460 , P1_U5832 , P1_U5831 );
nand NAND2_863 ( P1_U3461 , P1_U5834 , P1_U5833 );
nand NAND2_864 ( P1_U3462 , P1_U5837 , P1_U5836 );
nand NAND2_865 ( P1_U3463 , P1_U5839 , P1_U5838 );
nand NAND2_866 ( P1_U3464 , P1_U5841 , P1_U5840 );
nand NAND2_867 ( P1_U3465 , P1_U5844 , P1_U5843 );
nand NAND2_868 ( P1_U3466 , P1_U5846 , P1_U5845 );
nand NAND2_869 ( P1_U3467 , P1_U5848 , P1_U5847 );
nand NAND2_870 ( P1_U3468 , P1_U5851 , P1_U5850 );
nand NAND2_871 ( P1_U3469 , P1_U5853 , P1_U5852 );
nand NAND2_872 ( P1_U3470 , P1_U5855 , P1_U5854 );
nand NAND2_873 ( P1_U3471 , P1_U5858 , P1_U5857 );
nand NAND2_874 ( P1_U3472 , P1_U5860 , P1_U5859 );
nand NAND2_875 ( P1_U3473 , P1_U5862 , P1_U5861 );
nand NAND2_876 ( P1_U3474 , P1_U5865 , P1_U5864 );
nand NAND2_877 ( P1_U3475 , P1_U5867 , P1_U5866 );
nand NAND2_878 ( P1_U3476 , P1_U5869 , P1_U5868 );
nand NAND2_879 ( P1_U3477 , P1_U5872 , P1_U5871 );
nand NAND2_880 ( P1_U3478 , P1_U5874 , P1_U5873 );
nand NAND2_881 ( P1_U3479 , P1_U5876 , P1_U5875 );
nand NAND2_882 ( P1_U3480 , P1_U5879 , P1_U5878 );
nand NAND2_883 ( P1_U3481 , P1_U5881 , P1_U5880 );
nand NAND2_884 ( P1_U3482 , P1_U5883 , P1_U5882 );
nand NAND2_885 ( P1_U3483 , P1_U5886 , P1_U5885 );
nand NAND2_886 ( P1_U3484 , P1_U5888 , P1_U5887 );
nand NAND2_887 ( P1_U3485 , P1_U5890 , P1_U5889 );
nand NAND2_888 ( P1_U3486 , P1_U5893 , P1_U5892 );
nand NAND2_889 ( P1_U3487 , P1_U5895 , P1_U5894 );
nand NAND2_890 ( P1_U3488 , P1_U5897 , P1_U5896 );
nand NAND2_891 ( P1_U3489 , P1_U5900 , P1_U5899 );
nand NAND2_892 ( P1_U3490 , P1_U5902 , P1_U5901 );
nand NAND2_893 ( P1_U3491 , P1_U5904 , P1_U5903 );
nand NAND2_894 ( P1_U3492 , P1_U5907 , P1_U5906 );
nand NAND2_895 ( P1_U3493 , P1_U5909 , P1_U5908 );
nand NAND2_896 ( P1_U3494 , P1_U5911 , P1_U5910 );
nand NAND2_897 ( P1_U3495 , P1_U5914 , P1_U5913 );
nand NAND2_898 ( P1_U3496 , P1_U5916 , P1_U5915 );
nand NAND2_899 ( P1_U3497 , P1_U5918 , P1_U5917 );
nand NAND2_900 ( P1_U3498 , P1_U5921 , P1_U5920 );
nand NAND2_901 ( P1_U3499 , P1_U5923 , P1_U5922 );
nand NAND2_902 ( P1_U3500 , P1_U5925 , P1_U5924 );
nand NAND2_903 ( P1_U3501 , P1_U5928 , P1_U5927 );
nand NAND2_904 ( P1_U3502 , P1_U5930 , P1_U5929 );
nand NAND2_905 ( P1_U3503 , P1_U5932 , P1_U5931 );
nand NAND2_906 ( P1_U3504 , P1_U5935 , P1_U5934 );
nand NAND2_907 ( P1_U3505 , P1_U5937 , P1_U5936 );
nand NAND2_908 ( P1_U3506 , P1_U5939 , P1_U5938 );
nand NAND2_909 ( P1_U3507 , P1_U5942 , P1_U5941 );
nand NAND2_910 ( P1_U3508 , P1_U5944 , P1_U5943 );
nand NAND2_911 ( P1_U3509 , P1_U5946 , P1_U5945 );
nand NAND2_912 ( P1_U3510 , P1_U5949 , P1_U5948 );
nand NAND2_913 ( P1_U3511 , P1_U5951 , P1_U5950 );
nand NAND2_914 ( P1_U3512 , P1_U5953 , P1_U5952 );
nand NAND2_915 ( P1_U3513 , P1_U5956 , P1_U5955 );
nand NAND2_916 ( P1_U3514 , P1_U5958 , P1_U5957 );
nand NAND2_917 ( P1_U3515 , P1_U5961 , P1_U5960 );
nand NAND2_918 ( P1_U3516 , P1_U5963 , P1_U5962 );
nand NAND2_919 ( P1_U3517 , P1_U5965 , P1_U5964 );
nand NAND2_920 ( P1_U3518 , P1_U5967 , P1_U5966 );
nand NAND2_921 ( P1_U3519 , P1_U5969 , P1_U5968 );
nand NAND2_922 ( P1_U3520 , P1_U5971 , P1_U5970 );
nand NAND2_923 ( P1_U3521 , P1_U5973 , P1_U5972 );
nand NAND2_924 ( P1_U3522 , P1_U5975 , P1_U5974 );
nand NAND2_925 ( P1_U3523 , P1_U5977 , P1_U5976 );
nand NAND2_926 ( P1_U3524 , P1_U5979 , P1_U5978 );
nand NAND2_927 ( P1_U3525 , P1_U5981 , P1_U5980 );
nand NAND2_928 ( P1_U3526 , P1_U5983 , P1_U5982 );
nand NAND2_929 ( P1_U3527 , P1_U5985 , P1_U5984 );
nand NAND2_930 ( P1_U3528 , P1_U5987 , P1_U5986 );
nand NAND2_931 ( P1_U3529 , P1_U5989 , P1_U5988 );
nand NAND2_932 ( P1_U3530 , P1_U5991 , P1_U5990 );
nand NAND2_933 ( P1_U3531 , P1_U5993 , P1_U5992 );
nand NAND2_934 ( P1_U3532 , P1_U5995 , P1_U5994 );
nand NAND2_935 ( P1_U3533 , P1_U5997 , P1_U5996 );
nand NAND2_936 ( P1_U3534 , P1_U5999 , P1_U5998 );
nand NAND2_937 ( P1_U3535 , P1_U6001 , P1_U6000 );
nand NAND2_938 ( P1_U3536 , P1_U6003 , P1_U6002 );
nand NAND2_939 ( P1_U3537 , P1_U6005 , P1_U6004 );
nand NAND2_940 ( P1_U3538 , P1_U6007 , P1_U6006 );
nand NAND2_941 ( P1_U3539 , P1_U6009 , P1_U6008 );
nand NAND2_942 ( P1_U3540 , P1_U6011 , P1_U6010 );
nand NAND2_943 ( P1_U3541 , P1_U6013 , P1_U6012 );
nand NAND2_944 ( P1_U3542 , P1_U6015 , P1_U6014 );
nand NAND2_945 ( P1_U3543 , P1_U6017 , P1_U6016 );
nand NAND2_946 ( P1_U3544 , P1_U6019 , P1_U6018 );
nand NAND2_947 ( P1_U3545 , P1_U6021 , P1_U6020 );
nand NAND2_948 ( P1_U3546 , P1_U6023 , P1_U6022 );
nand NAND2_949 ( P1_U3547 , P1_U6025 , P1_U6024 );
nand NAND2_950 ( P1_U3548 , P1_U6027 , P1_U6026 );
nand NAND2_951 ( P1_U3549 , P1_U6029 , P1_U6028 );
nand NAND2_952 ( P1_U3550 , P1_U6031 , P1_U6030 );
nand NAND2_953 ( P1_U3551 , P1_U6033 , P1_U6032 );
nand NAND2_954 ( P1_U3552 , P1_U6035 , P1_U6034 );
nand NAND2_955 ( P1_U3553 , P1_U6037 , P1_U6036 );
nand NAND2_956 ( P1_U3554 , P1_U6039 , P1_U6038 );
nand NAND2_957 ( P1_U3555 , P1_U6041 , P1_U6040 );
nand NAND2_958 ( P1_U3556 , P1_U6043 , P1_U6042 );
nand NAND2_959 ( P1_U3557 , P1_U6045 , P1_U6044 );
nand NAND2_960 ( P1_U3558 , P1_U6047 , P1_U6046 );
nand NAND2_961 ( P1_U3559 , P1_U6049 , P1_U6048 );
nand NAND2_962 ( P1_U3560 , P1_U6115 , P1_U6114 );
nand NAND2_963 ( P1_U3561 , P1_U6117 , P1_U6116 );
nand NAND2_964 ( P1_U3562 , P1_U6119 , P1_U6118 );
nand NAND2_965 ( P1_U3563 , P1_U6121 , P1_U6120 );
nand NAND2_966 ( P1_U3564 , P1_U6123 , P1_U6122 );
nand NAND2_967 ( P1_U3565 , P1_U6125 , P1_U6124 );
nand NAND2_968 ( P1_U3566 , P1_U6127 , P1_U6126 );
nand NAND2_969 ( P1_U3567 , P1_U6129 , P1_U6128 );
nand NAND2_970 ( P1_U3568 , P1_U6131 , P1_U6130 );
nand NAND2_971 ( P1_U3569 , P1_U6133 , P1_U6132 );
nand NAND2_972 ( P1_U3570 , P1_U6135 , P1_U6134 );
nand NAND2_973 ( P1_U3571 , P1_U6137 , P1_U6136 );
nand NAND2_974 ( P1_U3572 , P1_U6139 , P1_U6138 );
nand NAND2_975 ( P1_U3573 , P1_U6141 , P1_U6140 );
nand NAND2_976 ( P1_U3574 , P1_U6143 , P1_U6142 );
nand NAND2_977 ( P1_U3575 , P1_U6145 , P1_U6144 );
nand NAND2_978 ( P1_U3576 , P1_U6147 , P1_U6146 );
nand NAND2_979 ( P1_U3577 , P1_U6149 , P1_U6148 );
nand NAND2_980 ( P1_U3578 , P1_U6151 , P1_U6150 );
nand NAND2_981 ( P1_U3579 , P1_U6153 , P1_U6152 );
nand NAND2_982 ( P1_U3580 , P1_U6155 , P1_U6154 );
nand NAND2_983 ( P1_U3581 , P1_U6157 , P1_U6156 );
nand NAND2_984 ( P1_U3582 , P1_U6159 , P1_U6158 );
nand NAND2_985 ( P1_U3583 , P1_U6161 , P1_U6160 );
nand NAND2_986 ( P1_U3584 , P1_U6163 , P1_U6162 );
nand NAND2_987 ( P1_U3585 , P1_U6165 , P1_U6164 );
nand NAND2_988 ( P1_U3586 , P1_U6167 , P1_U6166 );
nand NAND2_989 ( P1_U3587 , P1_U6169 , P1_U6168 );
nand NAND2_990 ( P1_U3588 , P1_U6171 , P1_U6170 );
nand NAND2_991 ( P1_U3589 , P1_U6173 , P1_U6172 );
nand NAND2_992 ( P1_U3590 , P1_U6175 , P1_U6174 );
nand NAND2_993 ( P1_U3591 , P1_U6177 , P1_U6176 );
and AND2_994 ( P1_U3592 , P1_U5786 , P1_STATE_REG );
and AND2_995 ( P1_U3593 , P1_U4187 , P1_U4186 );
and AND2_996 ( P1_U3594 , P1_U4189 , P1_U4188 );
and AND2_997 ( P1_U3595 , P1_U4195 , P1_U4196 );
and AND4_998 ( P1_U3596 , P1_U4151 , P1_U4150 , P1_U4149 , P1_U4148 );
and AND4_999 ( P1_U3597 , P1_U4155 , P1_U4154 , P1_U4153 , P1_U4152 );
and AND4_1000 ( P1_U3598 , P1_U4159 , P1_U4158 , P1_U4157 , P1_U4156 );
and AND3_1001 ( P1_U3599 , P1_U4161 , P1_U4160 , P1_U4162 );
and AND4_1002 ( P1_U3600 , P1_U3599 , P1_U3598 , P1_U3597 , P1_U3596 );
and AND4_1003 ( P1_U3601 , P1_U4166 , P1_U4165 , P1_U4164 , P1_U4163 );
and AND4_1004 ( P1_U3602 , P1_U4170 , P1_U4169 , P1_U4168 , P1_U4167 );
and AND4_1005 ( P1_U3603 , P1_U4174 , P1_U4173 , P1_U4172 , P1_U4171 );
and AND3_1006 ( P1_U3604 , P1_U4176 , P1_U4175 , P1_U4177 );
and AND4_1007 ( P1_U3605 , P1_U3604 , P1_U3603 , P1_U3602 , P1_U3601 );
and AND2_1008 ( P1_U3606 , P1_U5825 , P1_U4179 );
and AND2_1009 ( P1_U3607 , P1_U5828 , P1_U3022 );
and AND2_1010 ( P1_U3608 , P1_U4212 , P1_U4211 );
and AND2_1011 ( P1_U3609 , P1_U4214 , P1_U4213 );
and AND3_1012 ( P1_U3610 , P1_U4216 , P1_U4215 , P1_U3609 );
and AND4_1013 ( P1_U3611 , P1_U4220 , P1_U4218 , P1_U4221 , P1_U4219 );
and AND2_1014 ( P1_U3612 , P1_U4231 , P1_U4230 );
and AND2_1015 ( P1_U3613 , P1_U4233 , P1_U4232 );
and AND3_1016 ( P1_U3614 , P1_U4235 , P1_U4234 , P1_U3613 );
and AND4_1017 ( P1_U3615 , P1_U4239 , P1_U4237 , P1_U4240 , P1_U4238 );
and AND2_1018 ( P1_U3616 , P1_U4250 , P1_U4249 );
and AND2_1019 ( P1_U3617 , P1_U4252 , P1_U4251 );
and AND3_1020 ( P1_U3618 , P1_U4254 , P1_U4253 , P1_U3617 );
and AND4_1021 ( P1_U3619 , P1_U4258 , P1_U4256 , P1_U4259 , P1_U4257 );
and AND2_1022 ( P1_U3620 , P1_U4269 , P1_U4268 );
and AND2_1023 ( P1_U3621 , P1_U4271 , P1_U4270 );
and AND3_1024 ( P1_U3622 , P1_U4273 , P1_U4272 , P1_U3621 );
and AND4_1025 ( P1_U3623 , P1_U4277 , P1_U4275 , P1_U4278 , P1_U4276 );
and AND2_1026 ( P1_U3624 , P1_U4288 , P1_U4287 );
and AND2_1027 ( P1_U3625 , P1_U4290 , P1_U4289 );
and AND3_1028 ( P1_U3626 , P1_U4292 , P1_U4291 , P1_U3625 );
and AND4_1029 ( P1_U3627 , P1_U4296 , P1_U4294 , P1_U4297 , P1_U4295 );
and AND2_1030 ( P1_U3628 , P1_U4307 , P1_U4306 );
and AND2_1031 ( P1_U3629 , P1_U4309 , P1_U4308 );
and AND3_1032 ( P1_U3630 , P1_U4311 , P1_U4310 , P1_U3629 );
and AND4_1033 ( P1_U3631 , P1_U4315 , P1_U4313 , P1_U4316 , P1_U4314 );
and AND2_1034 ( P1_U3632 , P1_U4326 , P1_U4325 );
and AND2_1035 ( P1_U3633 , P1_U4328 , P1_U4327 );
and AND3_1036 ( P1_U3634 , P1_U4330 , P1_U4329 , P1_U3633 );
and AND4_1037 ( P1_U3635 , P1_U4334 , P1_U4332 , P1_U4335 , P1_U4333 );
and AND2_1038 ( P1_U3636 , P1_U4345 , P1_U4344 );
and AND2_1039 ( P1_U3637 , P1_U4347 , P1_U4346 );
and AND3_1040 ( P1_U3638 , P1_U4349 , P1_U4348 , P1_U3637 );
and AND4_1041 ( P1_U3639 , P1_U4353 , P1_U4351 , P1_U4354 , P1_U4352 );
and AND2_1042 ( P1_U3640 , P1_U4364 , P1_U4363 );
and AND2_1043 ( P1_U3641 , P1_U4366 , P1_U4365 );
and AND3_1044 ( P1_U3642 , P1_U4368 , P1_U4367 , P1_U3641 );
and AND4_1045 ( P1_U3643 , P1_U4372 , P1_U4370 , P1_U4373 , P1_U4371 );
and AND2_1046 ( P1_U3644 , P1_U4383 , P1_U4382 );
and AND2_1047 ( P1_U3645 , P1_U4385 , P1_U4384 );
and AND3_1048 ( P1_U3646 , P1_U4387 , P1_U4386 , P1_U3645 );
and AND4_1049 ( P1_U3647 , P1_U4391 , P1_U4389 , P1_U4392 , P1_U4390 );
and AND2_1050 ( P1_U3648 , P1_U4402 , P1_U4401 );
and AND2_1051 ( P1_U3649 , P1_U4404 , P1_U4403 );
and AND3_1052 ( P1_U3650 , P1_U4406 , P1_U4405 , P1_U3649 );
and AND4_1053 ( P1_U3651 , P1_U4411 , P1_U4410 , P1_U4409 , P1_U4408 );
and AND2_1054 ( P1_U3652 , P1_U4421 , P1_U4420 );
and AND2_1055 ( P1_U3653 , P1_U4423 , P1_U4422 );
and AND3_1056 ( P1_U3654 , P1_U4425 , P1_U4424 , P1_U3653 );
and AND4_1057 ( P1_U3655 , P1_U4430 , P1_U4428 , P1_U4429 , P1_U4427 );
and AND2_1058 ( P1_U3656 , P1_U4440 , P1_U4439 );
and AND2_1059 ( P1_U3657 , P1_U4442 , P1_U4441 );
and AND3_1060 ( P1_U3658 , P1_U4444 , P1_U4443 , P1_U3657 );
and AND4_1061 ( P1_U3659 , P1_U4449 , P1_U4448 , P1_U4447 , P1_U4446 );
and AND2_1062 ( P1_U3660 , P1_U4459 , P1_U4458 );
and AND2_1063 ( P1_U3661 , P1_U4461 , P1_U4460 );
and AND3_1064 ( P1_U3662 , P1_U4463 , P1_U4462 , P1_U3661 );
and AND4_1065 ( P1_U3663 , P1_U4468 , P1_U4466 , P1_U4467 , P1_U4465 );
and AND2_1066 ( P1_U3664 , P1_U4478 , P1_U4477 );
and AND2_1067 ( P1_U3665 , P1_U4480 , P1_U4479 );
and AND3_1068 ( P1_U3666 , P1_U4482 , P1_U4481 , P1_U3665 );
and AND4_1069 ( P1_U3667 , P1_U4486 , P1_U4484 , P1_U4487 , P1_U4485 );
and AND2_1070 ( P1_U3668 , P1_U4497 , P1_U4496 );
and AND2_1071 ( P1_U3669 , P1_U4499 , P1_U4498 );
and AND3_1072 ( P1_U3670 , P1_U4501 , P1_U4500 , P1_U3669 );
and AND4_1073 ( P1_U3671 , P1_U4505 , P1_U4503 , P1_U4506 , P1_U4504 );
and AND2_1074 ( P1_U3672 , P1_U4516 , P1_U4515 );
and AND2_1075 ( P1_U3673 , P1_U4518 , P1_U4517 );
and AND3_1076 ( P1_U3674 , P1_U4520 , P1_U4519 , P1_U3673 );
and AND4_1077 ( P1_U3675 , P1_U4525 , P1_U4523 , P1_U4524 , P1_U4522 );
and AND2_1078 ( P1_U3676 , P1_U4535 , P1_U4534 );
and AND2_1079 ( P1_U3677 , P1_U4537 , P1_U4536 );
and AND3_1080 ( P1_U3678 , P1_U4539 , P1_U4538 , P1_U3677 );
and AND4_1081 ( P1_U3679 , P1_U4544 , P1_U4542 , P1_U4543 , P1_U4541 );
and AND2_1082 ( P1_U3680 , P1_U4554 , P1_U4553 );
and AND2_1083 ( P1_U3681 , P1_U4556 , P1_U4555 );
and AND3_1084 ( P1_U3682 , P1_U4558 , P1_U4557 , P1_U3681 );
and AND4_1085 ( P1_U3683 , P1_U4562 , P1_U4560 , P1_U4563 , P1_U4561 );
and AND2_1086 ( P1_U3684 , P1_U4573 , P1_U4572 );
and AND2_1087 ( P1_U3685 , P1_U4575 , P1_U4574 );
and AND3_1088 ( P1_U3686 , P1_U4577 , P1_U4576 , P1_U3685 );
and AND4_1089 ( P1_U3687 , P1_U4581 , P1_U4579 , P1_U4582 , P1_U4580 );
and AND2_1090 ( P1_U3688 , P1_U4592 , P1_U4591 );
and AND2_1091 ( P1_U3689 , P1_U4594 , P1_U4593 );
and AND3_1092 ( P1_U3690 , P1_U4596 , P1_U4595 , P1_U3689 );
and AND4_1093 ( P1_U3691 , P1_U4600 , P1_U4598 , P1_U4601 , P1_U4599 );
and AND2_1094 ( P1_U3692 , P1_U4611 , P1_U4610 );
and AND2_1095 ( P1_U3693 , P1_U4613 , P1_U4612 );
and AND3_1096 ( P1_U3694 , P1_U4615 , P1_U4614 , P1_U3693 );
and AND4_1097 ( P1_U3695 , P1_U4619 , P1_U4617 , P1_U4620 , P1_U4618 );
and AND2_1098 ( P1_U3696 , P1_U4630 , P1_U4629 );
and AND2_1099 ( P1_U3697 , P1_U4632 , P1_U4631 );
and AND3_1100 ( P1_U3698 , P1_U4634 , P1_U4633 , P1_U3697 );
and AND4_1101 ( P1_U3699 , P1_U4638 , P1_U4636 , P1_U4639 , P1_U4637 );
and AND2_1102 ( P1_U3700 , P1_U4649 , P1_U4648 );
and AND2_1103 ( P1_U3701 , P1_U4651 , P1_U4650 );
and AND3_1104 ( P1_U3702 , P1_U4653 , P1_U4652 , P1_U3701 );
and AND4_1105 ( P1_U3703 , P1_U4657 , P1_U4655 , P1_U4658 , P1_U4656 );
and AND2_1106 ( P1_U3704 , P1_U4668 , P1_U4667 );
and AND2_1107 ( P1_U3705 , P1_U4670 , P1_U4669 );
and AND3_1108 ( P1_U3706 , P1_U4672 , P1_U4671 , P1_U3705 );
and AND4_1109 ( P1_U3707 , P1_U4676 , P1_U4674 , P1_U4677 , P1_U4675 );
and AND2_1110 ( P1_U3708 , P1_U4687 , P1_U4686 );
and AND2_1111 ( P1_U3709 , P1_U4689 , P1_U4688 );
and AND3_1112 ( P1_U3710 , P1_U4691 , P1_U4690 , P1_U3709 );
and AND4_1113 ( P1_U3711 , P1_U4695 , P1_U4693 , P1_U4696 , P1_U4694 );
and AND2_1114 ( P1_U3712 , P1_U4706 , P1_U4705 );
and AND2_1115 ( P1_U3713 , P1_U4708 , P1_U4707 );
and AND3_1116 ( P1_U3714 , P1_U4710 , P1_U4709 , P1_U3713 );
and AND4_1117 ( P1_U3715 , P1_U4714 , P1_U4712 , P1_U4715 , P1_U4713 );
and AND2_1118 ( P1_U3716 , P1_U4725 , P1_U4724 );
and AND2_1119 ( P1_U3717 , P1_U4727 , P1_U4726 );
and AND3_1120 ( P1_U3718 , P1_U4729 , P1_U4728 , P1_U3717 );
and AND4_1121 ( P1_U3719 , P1_U4733 , P1_U4731 , P1_U4734 , P1_U4732 );
and AND2_1122 ( P1_U3720 , P1_U4741 , P1_U4030 );
and AND5_1123 ( P1_U3721 , P1_U4743 , P1_U4742 , P1_U4744 , P1_U4745 , P1_U4746 );
and AND2_1124 ( P1_U3722 , P1_U4748 , P1_U4747 );
and AND3_1125 ( P1_U3723 , P1_U4750 , P1_U4749 , P1_U3722 );
and AND3_1126 ( P1_U3724 , P1_U4753 , P1_U4754 , P1_U4752 );
and AND2_1127 ( P1_U3725 , P1_U4030 , P1_U4741 );
and AND2_1128 ( P1_U3726 , P1_U3022 , P1_U3457 );
and AND3_1129 ( P1_U3727 , P1_U5828 , P1_U4012 , P1_U3458 );
and AND3_1130 ( P1_U3728 , P1_U4771 , P1_U4770 , P1_U4772 );
and AND3_1131 ( P1_U3729 , P1_U4774 , P1_U4773 , P1_U3957 );
and AND3_1132 ( P1_U3730 , P1_U4776 , P1_U4775 , P1_U4777 );
and AND3_1133 ( P1_U3731 , P1_U4779 , P1_U4778 , P1_U3958 );
and AND3_1134 ( P1_U3732 , P1_U4781 , P1_U4780 , P1_U4782 );
and AND3_1135 ( P1_U3733 , P1_U4784 , P1_U4783 , P1_U3959 );
and AND3_1136 ( P1_U3734 , P1_U4786 , P1_U4785 , P1_U4787 );
and AND3_1137 ( P1_U3735 , P1_U4789 , P1_U4788 , P1_U3960 );
and AND3_1138 ( P1_U3736 , P1_U4791 , P1_U4790 , P1_U4792 );
and AND3_1139 ( P1_U3737 , P1_U4794 , P1_U4793 , P1_U3961 );
and AND3_1140 ( P1_U3738 , P1_U4796 , P1_U4795 , P1_U4797 );
and AND2_1141 ( P1_U3739 , P1_U4799 , P1_U4798 );
and AND3_1142 ( P1_U3740 , P1_U4801 , P1_U4800 , P1_U4802 );
and AND2_1143 ( P1_U3741 , P1_U4804 , P1_U4803 );
and AND3_1144 ( P1_U3742 , P1_U4806 , P1_U4805 , P1_U4807 );
and AND2_1145 ( P1_U3743 , P1_U4809 , P1_U4808 );
and AND3_1146 ( P1_U3744 , P1_U4811 , P1_U4810 , P1_U4812 );
and AND2_1147 ( P1_U3745 , P1_U4814 , P1_U4813 );
and AND2_1148 ( P1_U3746 , P1_U4816 , P1_U4815 );
and AND2_1149 ( P1_U3747 , P1_U4819 , P1_U4818 );
and AND2_1150 ( P1_U3748 , P1_U4821 , P1_U4820 );
and AND2_1151 ( P1_U3749 , P1_U4824 , P1_U4823 );
and AND3_1152 ( P1_U3750 , P1_U4826 , P1_U4825 , P1_U4827 );
and AND2_1153 ( P1_U3751 , P1_U4829 , P1_U4828 );
and AND3_1154 ( P1_U3752 , P1_U4831 , P1_U4830 , P1_U4832 );
and AND2_1155 ( P1_U3753 , P1_U4834 , P1_U4833 );
and AND3_1156 ( P1_U3754 , P1_U4836 , P1_U4835 , P1_U4837 );
and AND2_1157 ( P1_U3755 , P1_U4839 , P1_U4838 );
and AND3_1158 ( P1_U3756 , P1_U4841 , P1_U4840 , P1_U4842 );
and AND2_1159 ( P1_U3757 , P1_U4844 , P1_U4843 );
and AND2_1160 ( P1_U3758 , P1_U4846 , P1_U4845 );
and AND2_1161 ( P1_U3759 , P1_U4849 , P1_U4848 );
and AND2_1162 ( P1_U3760 , P1_U4851 , P1_U4850 );
and AND2_1163 ( P1_U3761 , P1_U4854 , P1_U4853 );
and AND3_1164 ( P1_U3762 , P1_U4856 , P1_U4855 , P1_U4857 );
and AND2_1165 ( P1_U3763 , P1_U4859 , P1_U4858 );
and AND3_1166 ( P1_U3764 , P1_U4861 , P1_U4860 , P1_U4862 );
and AND2_1167 ( P1_U3765 , P1_U4864 , P1_U4863 );
and AND2_1168 ( P1_U3766 , P1_U4866 , P1_U4865 );
and AND2_1169 ( P1_U3767 , P1_U4869 , P1_U4868 );
and AND2_1170 ( P1_U3768 , P1_U4871 , P1_U4870 );
and AND2_1171 ( P1_U3769 , P1_U4874 , P1_U4873 );
and AND2_1172 ( P1_U3770 , P1_U4876 , P1_U4875 );
and AND2_1173 ( P1_U3771 , P1_U4879 , P1_U4878 );
and AND2_1174 ( P1_U3772 , P1_U4881 , P1_U4880 );
and AND2_1175 ( P1_U3773 , P1_U4884 , P1_U4883 );
and AND2_1176 ( P1_U3774 , P1_U4886 , P1_U4885 );
and AND2_1177 ( P1_U3775 , P1_U4889 , P1_U4888 );
and AND2_1178 ( P1_U3776 , P1_U4891 , P1_U4890 );
and AND2_1179 ( P1_U3777 , P1_U4894 , P1_U4893 );
and AND2_1180 ( P1_U3778 , P1_U4896 , P1_U4895 );
and AND2_1181 ( P1_U3779 , P1_U4899 , P1_U4898 );
and AND2_1182 ( P1_U3780 , P1_U4901 , P1_U4900 );
and AND2_1183 ( P1_U3781 , P1_U4904 , P1_U4903 );
and AND2_1184 ( P1_U3782 , P1_U4906 , P1_U4905 );
and AND2_1185 ( P1_U3783 , P1_U4909 , P1_U4908 );
and AND2_1186 ( P1_U3784 , P1_U4911 , P1_U4910 );
and AND2_1187 ( P1_U3785 , P1_U4914 , P1_U4913 );
and AND3_1188 ( P1_U3786 , P1_U3362 , P1_U3364 , P1_U3370 );
and AND3_1189 ( P1_U3787 , P1_U3366 , P1_U3422 , P1_U3365 );
and AND2_1190 ( P1_U3788 , P1_U3361 , P1_U4006 );
and AND2_1191 ( P1_U3789 , P1_U3788 , P1_U3424 );
and AND2_1192 ( P1_U3790 , P1_U4934 , P1_U4935 );
and AND3_1193 ( P1_U3791 , P1_U4938 , P1_U4936 , P1_U4937 );
and AND2_1194 ( P1_U3792 , P1_U4944 , P1_U4945 );
and AND3_1195 ( P1_U3793 , P1_U4948 , P1_U4946 , P1_U4947 );
and AND2_1196 ( P1_U3794 , P1_U4954 , P1_U4955 );
and AND3_1197 ( P1_U3795 , P1_U4958 , P1_U4956 , P1_U4957 );
and AND2_1198 ( P1_U3796 , P1_U4964 , P1_U4965 );
and AND3_1199 ( P1_U3797 , P1_U4968 , P1_U4966 , P1_U4967 );
and AND2_1200 ( P1_U3798 , P1_U4974 , P1_U4975 );
and AND3_1201 ( P1_U3799 , P1_U4978 , P1_U4976 , P1_U4977 );
and AND2_1202 ( P1_U3800 , P1_U4984 , P1_U4985 );
and AND3_1203 ( P1_U3801 , P1_U4988 , P1_U4986 , P1_U4987 );
and AND2_1204 ( P1_U3802 , P1_U4994 , P1_U4995 );
and AND3_1205 ( P1_U3803 , P1_U4998 , P1_U4996 , P1_U4997 );
and AND2_1206 ( P1_U3804 , P1_U5004 , P1_U5005 );
and AND3_1207 ( P1_U3805 , P1_U5008 , P1_U5006 , P1_U5007 );
and AND2_1208 ( P1_U3806 , P1_U5014 , P1_U5015 );
and AND3_1209 ( P1_U3807 , P1_U5018 , P1_U5016 , P1_U5017 );
and AND2_1210 ( P1_U3808 , P1_U5024 , P1_U5025 );
and AND3_1211 ( P1_U3809 , P1_U5028 , P1_U5026 , P1_U5027 );
and AND2_1212 ( P1_U3810 , P1_U5034 , P1_U5035 );
and AND3_1213 ( P1_U3811 , P1_U5038 , P1_U5036 , P1_U5037 );
and AND2_1214 ( P1_U3812 , P1_U5044 , P1_U5045 );
and AND3_1215 ( P1_U3813 , P1_U5048 , P1_U5046 , P1_U5047 );
and AND2_1216 ( P1_U3814 , P1_U5054 , P1_U5055 );
and AND3_1217 ( P1_U3815 , P1_U5058 , P1_U5056 , P1_U5057 );
and AND2_1218 ( P1_U3816 , P1_U5064 , P1_U5065 );
and AND3_1219 ( P1_U3817 , P1_U5067 , P1_U5066 , P1_U5068 );
and AND2_1220 ( P1_U3818 , P1_U5074 , P1_U5075 );
and AND3_1221 ( P1_U3819 , P1_U5077 , P1_U5076 , P1_U5078 );
and AND2_1222 ( P1_U3820 , P1_U3821 , P1_U5084 );
and AND2_1223 ( P1_U3821 , P1_U5085 , P1_U4040 );
and AND3_1224 ( P1_U3822 , P1_U5087 , P1_U5086 , P1_U5088 );
and AND2_1225 ( P1_U3823 , P1_U5094 , P1_U5095 );
and AND3_1226 ( P1_U3824 , P1_U5097 , P1_U5096 , P1_U5098 );
and AND2_1227 ( P1_U3825 , P1_U3826 , P1_U5104 );
and AND2_1228 ( P1_U3826 , P1_U5105 , P1_U4040 );
and AND3_1229 ( P1_U3827 , P1_U5107 , P1_U5106 , P1_U5108 );
and AND2_1230 ( P1_U3828 , P1_U5114 , P1_U5115 );
and AND3_1231 ( P1_U3829 , P1_U5117 , P1_U5116 , P1_U5118 );
and AND2_1232 ( P1_U3830 , P1_U5124 , P1_U5125 );
and AND3_1233 ( P1_U3831 , P1_U5127 , P1_U5126 , P1_U5128 );
and AND3_1234 ( P1_U3832 , P1_U6218 , P1_U6215 , P1_U6221 );
and AND3_1235 ( P1_U3833 , P1_U3834 , P1_U3832 , P1_U6233 );
and AND3_1236 ( P1_U3834 , P1_U6230 , P1_U6227 , P1_U6224 );
and AND3_1237 ( P1_U3835 , P1_U6242 , P1_U6239 , P1_U6245 );
and AND3_1238 ( P1_U3836 , P1_U6251 , P1_U6248 , P1_U6254 );
and AND3_1239 ( P1_U3837 , P1_U3836 , P1_U3835 , P1_U6236 );
and AND3_1240 ( P1_U3838 , P1_U6188 , P1_U6185 , P1_U6191 );
and AND5_1241 ( P1_U3839 , P1_U6203 , P1_U6200 , P1_U6197 , P1_U6194 , P1_U6206 );
and AND4_1242 ( P1_U3840 , P1_U6269 , P1_U6266 , P1_U6263 , P1_U6260 );
and AND2_1243 ( P1_U3841 , P1_U6275 , P1_U6272 );
and AND2_1244 ( P1_U3842 , P1_U3841 , P1_U3840 );
and AND5_1245 ( P1_U3843 , P1_U3837 , P1_U3833 , P1_U6212 , P1_U6257 , P1_U6209 );
and AND3_1246 ( P1_U3844 , P1_U3839 , P1_U3838 , P1_U6182 );
and AND2_1247 ( P1_U3845 , P1_U3429 , P1_STATE_REG );
and AND2_1248 ( P1_U3846 , P1_U5138 , P1_U5136 );
and AND2_1249 ( P1_U3847 , P1_U3457 , P1_U3458 );
and AND3_1250 ( P1_U3848 , P1_U3997 , P1_U3371 , P1_U3996 );
and AND2_1251 ( P1_U3849 , P1_U3368 , P1_U3424 );
and AND2_1252 ( P1_U3850 , P1_U3427 , P1_U3430 );
and AND2_1253 ( P1_U3851 , P1_U3022 , P1_U5145 );
and AND2_1254 ( P1_U3852 , P1_U3425 , P1_STATE_REG );
and AND2_1255 ( P1_U3853 , P1_U5173 , P1_U5172 );
and AND2_1256 ( P1_U3854 , P1_U5189 , P1_U5187 );
and AND2_1257 ( P1_U3855 , P1_U5191 , P1_U5190 );
and AND2_1258 ( P1_U3856 , P1_U5200 , P1_U5199 );
and AND2_1259 ( P1_U3857 , P1_U5218 , P1_U5217 );
and AND2_1260 ( P1_U3858 , P1_U4037 , P1_U3078 );
and AND3_1261 ( P1_U3859 , P1_U5232 , P1_U5231 , P1_U3860 );
and AND2_1262 ( P1_U3860 , P1_U5235 , P1_U5234 );
and AND2_1263 ( P1_U3861 , P1_U5244 , P1_U5243 );
and AND2_1264 ( P1_U3862 , P1_U5251 , P1_U5249 );
and AND2_1265 ( P1_U3863 , P1_U5253 , P1_U5252 );
and AND2_1266 ( P1_U3864 , P1_U5280 , P1_U5279 );
and AND2_1267 ( P1_U3865 , P1_U5307 , P1_U5306 );
and AND2_1268 ( P1_U3866 , P1_U5323 , P1_U5321 );
and AND2_1269 ( P1_U3867 , P1_U5325 , P1_U5324 );
and AND2_1270 ( P1_U3868 , P1_U5334 , P1_U5333 );
and AND2_1271 ( P1_U3869 , P1_U5359 , P1_U5357 );
and AND2_1272 ( P1_U3870 , P1_U5361 , P1_U5360 );
and AND2_1273 ( P1_U3871 , P1_U5370 , P1_U5369 );
and AND2_1274 ( P1_U3872 , P1_U5406 , P1_U5405 );
and AND2_1275 ( P1_U3873 , P1_U5802 , P1_U5793 );
and AND2_1276 ( P1_U3874 , P1_U3375 , P1_U5410 );
and AND2_1277 ( P1_U3875 , P1_U5475 , P1_U5476 );
and AND2_1278 ( P1_U3876 , P1_U5535 , P1_U5533 );
and AND2_1279 ( P1_U3877 , P1_U3444 , P1_U5538 );
and AND2_1280 ( P1_U3878 , P1_U3374 , P1_U3997 );
and AND2_1281 ( P1_U3879 , P1_U3878 , P1_U3371 );
and AND2_1282 ( P1_U3880 , P1_U3881 , P1_U5546 );
and AND2_1283 ( P1_U3881 , P1_U3444 , P1_U5544 );
and AND2_1284 ( P1_U3882 , P1_U3883 , P1_U5549 );
and AND2_1285 ( P1_U3883 , P1_U3444 , P1_U5547 );
and AND2_1286 ( P1_U3884 , P1_U3885 , P1_U5552 );
and AND2_1287 ( P1_U3885 , P1_U3444 , P1_U5550 );
and AND2_1288 ( P1_U3886 , P1_U3887 , P1_U5555 );
and AND2_1289 ( P1_U3887 , P1_U3444 , P1_U5553 );
and AND2_1290 ( P1_U3888 , P1_U3889 , P1_U5558 );
and AND2_1291 ( P1_U3889 , P1_U3444 , P1_U5556 );
and AND2_1292 ( P1_U3890 , P1_U3891 , P1_U5561 );
and AND2_1293 ( P1_U3891 , P1_U3444 , P1_U5559 );
and AND2_1294 ( P1_U3892 , P1_U5564 , P1_U5562 );
and AND2_1295 ( P1_U3893 , P1_U5567 , P1_U5565 );
and AND2_1296 ( P1_U3894 , P1_U3895 , P1_U5570 );
and AND2_1297 ( P1_U3895 , P1_U3444 , P1_U5568 );
and AND2_1298 ( P1_U3896 , P1_U3444 , P1_U5573 );
and AND2_1299 ( P1_U3897 , P1_U3444 , P1_U5576 );
and AND2_1300 ( P1_U3898 , P1_U3444 , P1_U5579 );
and AND2_1301 ( P1_U3899 , P1_U3444 , P1_U5582 );
and AND2_1302 ( P1_U3900 , P1_U3444 , P1_U5585 );
and AND2_1303 ( P1_U3901 , P1_U3444 , P1_U5588 );
and AND2_1304 ( P1_U3902 , P1_U3444 , P1_U5591 );
and AND2_1305 ( P1_U3903 , P1_U3444 , P1_U5594 );
and AND2_1306 ( P1_U3904 , P1_U3444 , P1_U5597 );
and AND2_1307 ( P1_U3905 , P1_U3444 , P1_U5600 );
and AND2_1308 ( P1_U3906 , P1_U3907 , P1_U5603 );
and AND2_1309 ( P1_U3907 , P1_U3444 , P1_U5601 );
and AND2_1310 ( P1_U3908 , P1_U3444 , P1_U5606 );
and AND2_1311 ( P1_U3909 , P1_U3444 , P1_U5609 );
and AND2_1312 ( P1_U3910 , P1_U3444 , P1_U5612 );
and AND2_1313 ( P1_U3911 , P1_U3444 , P1_U5615 );
and AND2_1314 ( P1_U3912 , P1_U3444 , P1_U5618 );
and AND2_1315 ( P1_U3913 , P1_U3444 , P1_U5621 );
and AND2_1316 ( P1_U3914 , P1_U3444 , P1_U5624 );
and AND2_1317 ( P1_U3915 , P1_U3444 , P1_U5627 );
and AND2_1318 ( P1_U3916 , P1_U3444 , P1_U5630 );
and AND2_1319 ( P1_U3917 , P1_U3444 , P1_U5633 );
and AND2_1320 ( P1_U3918 , P1_U3919 , P1_U5636 );
and AND2_1321 ( P1_U3919 , P1_U3444 , P1_U5634 );
and AND2_1322 ( P1_U3920 , P1_U3921 , P1_U5639 );
and AND2_1323 ( P1_U3921 , P1_U3444 , P1_U5637 );
and AND2_1324 ( P1_U3922 , P1_U5645 , P1_U5642 );
and AND2_1325 ( P1_U3923 , P1_U5649 , P1_U5646 );
and AND2_1326 ( P1_U3924 , P1_U5651 , P1_U5650 );
and AND2_1327 ( P1_U3925 , P1_U5655 , P1_U5654 );
and AND2_1328 ( P1_U3926 , P1_U5659 , P1_U5658 );
and AND2_1329 ( P1_U3927 , P1_U5663 , P1_U5662 );
and AND3_1330 ( P1_U3928 , P1_U5673 , P1_U5672 , P1_U5675 );
and AND2_1331 ( P1_U3929 , P1_U5677 , P1_U5676 );
and AND2_1332 ( P1_U3930 , P1_U5681 , P1_U5680 );
and AND2_1333 ( P1_U3931 , P1_U5685 , P1_U5684 );
and AND2_1334 ( P1_U3932 , P1_U5689 , P1_U5688 );
and AND2_1335 ( P1_U3933 , P1_U5693 , P1_U5692 );
and AND2_1336 ( P1_U3934 , P1_U5697 , P1_U5696 );
and AND2_1337 ( P1_U3935 , P1_U5701 , P1_U5700 );
and AND2_1338 ( P1_U3936 , P1_U5705 , P1_U5704 );
and AND2_1339 ( P1_U3937 , P1_U5709 , P1_U5708 );
and AND2_1340 ( P1_U3938 , P1_U5713 , P1_U5712 );
and AND3_1341 ( P1_U3939 , P1_U5717 , P1_U5716 , P1_U5719 );
and AND2_1342 ( P1_U3940 , P1_U5721 , P1_U5720 );
and AND2_1343 ( P1_U3941 , P1_U5725 , P1_U5724 );
and AND2_1344 ( P1_U3942 , P1_U5729 , P1_U5728 );
and AND2_1345 ( P1_U3943 , P1_U5733 , P1_U5732 );
and AND2_1346 ( P1_U3944 , P1_U5737 , P1_U5736 );
and AND2_1347 ( P1_U3945 , P1_U5741 , P1_U5740 );
and AND2_1348 ( P1_U3946 , P1_U5745 , P1_U5744 );
and AND2_1349 ( P1_U3947 , P1_U5749 , P1_U5748 );
and AND2_1350 ( P1_U3948 , P1_U5753 , P1_U5752 );
and AND2_1351 ( P1_U3949 , P1_U5757 , P1_U5756 );
and AND3_1352 ( P1_U3950 , P1_U5761 , P1_U5760 , P1_U5763 );
and AND2_1353 ( P1_U3951 , P1_U5765 , P1_U5764 );
not NOT1_1354 ( P1_U3952 , P1_IR_REG_31_ );
nand NAND2_1355 ( P1_U3953 , P1_U3022 , P1_U3360 );
nand NAND2_1356 ( P1_U3954 , P1_U5817 , P1_U5811 );
nand NAND2_1357 ( P1_U3955 , P1_U3607 , P1_U3046 );
nand NAND2_1358 ( P1_U3956 , P1_U3726 , P1_U3046 );
and AND2_1359 ( P1_U3957 , P1_U6051 , P1_U6050 );
and AND2_1360 ( P1_U3958 , P1_U6053 , P1_U6052 );
and AND2_1361 ( P1_U3959 , P1_U6055 , P1_U6054 );
and AND2_1362 ( P1_U3960 , P1_U6057 , P1_U6056 );
and AND2_1363 ( P1_U3961 , P1_U6059 , P1_U6058 );
and AND2_1364 ( P1_U3962 , P1_U6061 , P1_U6060 );
and AND2_1365 ( P1_U3963 , P1_U6063 , P1_U6062 );
and AND2_1366 ( P1_U3964 , P1_U6065 , P1_U6064 );
and AND2_1367 ( P1_U3965 , P1_U6067 , P1_U6066 );
and AND2_1368 ( P1_U3966 , P1_U6069 , P1_U6068 );
and AND2_1369 ( P1_U3967 , P1_U6071 , P1_U6070 );
and AND2_1370 ( P1_U3968 , P1_U6073 , P1_U6072 );
and AND2_1371 ( P1_U3969 , P1_U6075 , P1_U6074 );
and AND2_1372 ( P1_U3970 , P1_U6077 , P1_U6076 );
and AND2_1373 ( P1_U3971 , P1_U6079 , P1_U6078 );
and AND2_1374 ( P1_U3972 , P1_U6081 , P1_U6080 );
and AND2_1375 ( P1_U3973 , P1_U6083 , P1_U6082 );
and AND2_1376 ( P1_U3974 , P1_U6085 , P1_U6084 );
and AND2_1377 ( P1_U3975 , P1_U6087 , P1_U6086 );
and AND2_1378 ( P1_U3976 , P1_U6089 , P1_U6088 );
and AND2_1379 ( P1_U3977 , P1_U6091 , P1_U6090 );
and AND2_1380 ( P1_U3978 , P1_U6093 , P1_U6092 );
and AND2_1381 ( P1_U3979 , P1_U6095 , P1_U6094 );
and AND2_1382 ( P1_U3980 , P1_U6097 , P1_U6096 );
and AND2_1383 ( P1_U3981 , P1_U6099 , P1_U6098 );
and AND2_1384 ( P1_U3982 , P1_U6101 , P1_U6100 );
and AND2_1385 ( P1_U3983 , P1_U6103 , P1_U6102 );
and AND2_1386 ( P1_U3984 , P1_U6105 , P1_U6104 );
and AND2_1387 ( P1_U3985 , P1_U6107 , P1_U6106 );
and AND2_1388 ( P1_U3986 , P1_U6109 , P1_U6108 );
nand NAND2_1389 ( P1_U3987 , P1_U3725 , P1_U3056 );
and AND2_1390 ( P1_U3988 , P1_U6111 , P1_U6110 );
and AND2_1391 ( P1_U3989 , P1_U6113 , P1_U6112 );
and AND2_1392 ( P1_U3990 , P1_U6179 , P1_U6178 );
nand NAND3_1393 ( P1_U3991 , P1_U3842 , P1_U3843 , P1_U3844 );
not NOT1_1394 ( P1_U3992 , P1_U3371 );
not NOT1_1395 ( P1_U3993 , P1_U3374 );
not NOT1_1396 ( P1_U3994 , P1_U3364 );
not NOT1_1397 ( P1_U3995 , P1_U3423 );
nand NAND2_1398 ( P1_U3996 , P1_U4003 , P1_U5793 );
nand NAND2_1399 ( P1_U3997 , P1_U4041 , P1_U3451 );
not NOT1_1400 ( P1_U3998 , P1_U3419 );
nand NAND2_1401 ( P1_U3999 , P1_U4042 , P1_U5793 );
not NOT1_1402 ( P1_U4000 , P1_U3362 );
not NOT1_1403 ( P1_U4001 , P1_U3367 );
not NOT1_1404 ( P1_U4002 , P1_U3370 );
not NOT1_1405 ( P1_U4003 , P1_U3422 );
not NOT1_1406 ( P1_U4004 , P1_U3366 );
not NOT1_1407 ( P1_U4005 , P1_U3365 );
nand NAND2_1408 ( P1_U4006 , P1_U4044 , P1_U3451 );
not NOT1_1409 ( P1_U4007 , P1_U3361 );
not NOT1_1410 ( P1_U4008 , P1_U3424 );
not NOT1_1411 ( P1_U4009 , P1_U3421 );
nand NAND2_1412 ( P1_U4010 , P1_U3993 , P1_U3453 );
not NOT1_1413 ( P1_U4011 , P1_U3368 );
nand NAND2_1414 ( P1_U4012 , P1_U4030 , P1_U3369 );
nand NAND2_1415 ( P1_U4013 , P1_U3873 , P1_U3425 );
not NOT1_1416 ( P1_U4014 , P1_U3954 );
not NOT1_1417 ( P1_U4015 , P1_U3434 );
not NOT1_1418 ( P1_U4016 , P1_U3430 );
not NOT1_1419 ( P1_U4017 , P1_U3413 );
not NOT1_1420 ( P1_U4018 , P1_U3411 );
not NOT1_1421 ( P1_U4019 , P1_U3409 );
not NOT1_1422 ( P1_U4020 , P1_U3407 );
not NOT1_1423 ( P1_U4021 , P1_U3405 );
not NOT1_1424 ( P1_U4022 , P1_U3403 );
not NOT1_1425 ( P1_U4023 , P1_U3401 );
not NOT1_1426 ( P1_U4024 , P1_U3399 );
not NOT1_1427 ( P1_U4025 , P1_U3397 );
not NOT1_1428 ( P1_U4026 , P1_U3418 );
not NOT1_1429 ( P1_U4027 , P1_U3417 );
not NOT1_1430 ( P1_U4028 , P1_U3415 );
not NOT1_1431 ( P1_U4029 , P1_U3431 );
not NOT1_1432 ( P1_U4030 , P1_U3372 );
not NOT1_1433 ( P1_U4031 , P1_U3420 );
not NOT1_1434 ( P1_U4032 , P1_U3956 );
not NOT1_1435 ( P1_U4033 , P1_U3955 );
not NOT1_1436 ( P1_U4034 , P1_U3953 );
not NOT1_1437 ( P1_U4035 , P1_U3987 );
not NOT1_1438 ( P1_U4036 , P1_U3373 );
not NOT1_1439 ( P1_U4037 , P1_U3435 );
not NOT1_1440 ( P1_U4038 , P1_U3433 );
nand NAND2_1441 ( P1_U4039 , P1_U4009 , P1_U3022 );
nand NAND2_1442 ( P1_U4040 , P1_U4016 , P1_U3212 );
not NOT1_1443 ( P1_U4041 , P1_U3375 );
not NOT1_1444 ( P1_U4042 , P1_U3363 );
not NOT1_1445 ( P1_U4043 , P1_U3427 );
not NOT1_1446 ( P1_U4044 , P1_U3369 );
not NOT1_1447 ( P1_U4045 , P1_U3429 );
not NOT1_1448 ( P1_U4046 , P1_U3358 );
not NOT1_1449 ( P1_U4047 , P1_U3357 );
nand NAND2_1450 ( P1_U4048 , U125 , P1_U3086 );
nand NAND2_1451 ( P1_U4049 , P1_IR_REG_0_ , P1_U3029 );
nand NAND2_1452 ( P1_U4050 , P1_IR_REG_0_ , P1_U4047 );
nand NAND2_1453 ( P1_U4051 , U114 , P1_U3086 );
nand NAND2_1454 ( P1_U4052 , P1_SUB_88_U40 , P1_U3029 );
nand NAND2_1455 ( P1_U4053 , P1_IR_REG_1_ , P1_U4047 );
nand NAND2_1456 ( P1_U4054 , U103 , P1_U3086 );
nand NAND2_1457 ( P1_U4055 , P1_SUB_88_U21 , P1_U3029 );
nand NAND2_1458 ( P1_U4056 , P1_IR_REG_2_ , P1_U4047 );
nand NAND2_1459 ( P1_U4057 , U100 , P1_U3086 );
nand NAND2_1460 ( P1_U4058 , P1_SUB_88_U22 , P1_U3029 );
nand NAND2_1461 ( P1_U4059 , P1_IR_REG_3_ , P1_U4047 );
nand NAND2_1462 ( P1_U4060 , U99 , P1_U3086 );
nand NAND2_1463 ( P1_U4061 , P1_SUB_88_U23 , P1_U3029 );
nand NAND2_1464 ( P1_U4062 , P1_IR_REG_4_ , P1_U4047 );
nand NAND2_1465 ( P1_U4063 , U98 , P1_U3086 );
nand NAND2_1466 ( P1_U4064 , P1_SUB_88_U162 , P1_U3029 );
nand NAND2_1467 ( P1_U4065 , P1_IR_REG_5_ , P1_U4047 );
nand NAND2_1468 ( P1_U4066 , U97 , P1_U3086 );
nand NAND2_1469 ( P1_U4067 , P1_SUB_88_U24 , P1_U3029 );
nand NAND2_1470 ( P1_U4068 , P1_IR_REG_6_ , P1_U4047 );
nand NAND2_1471 ( P1_U4069 , U96 , P1_U3086 );
nand NAND2_1472 ( P1_U4070 , P1_SUB_88_U25 , P1_U3029 );
nand NAND2_1473 ( P1_U4071 , P1_IR_REG_7_ , P1_U4047 );
nand NAND2_1474 ( P1_U4072 , U95 , P1_U3086 );
nand NAND2_1475 ( P1_U4073 , P1_SUB_88_U26 , P1_U3029 );
nand NAND2_1476 ( P1_U4074 , P1_IR_REG_8_ , P1_U4047 );
nand NAND2_1477 ( P1_U4075 , U94 , P1_U3086 );
nand NAND2_1478 ( P1_U4076 , P1_SUB_88_U160 , P1_U3029 );
nand NAND2_1479 ( P1_U4077 , P1_IR_REG_9_ , P1_U4047 );
nand NAND2_1480 ( P1_U4078 , U124 , P1_U3086 );
nand NAND2_1481 ( P1_U4079 , P1_SUB_88_U6 , P1_U3029 );
nand NAND2_1482 ( P1_U4080 , P1_IR_REG_10_ , P1_U4047 );
nand NAND2_1483 ( P1_U4081 , U123 , P1_U3086 );
nand NAND2_1484 ( P1_U4082 , P1_SUB_88_U7 , P1_U3029 );
nand NAND2_1485 ( P1_U4083 , P1_IR_REG_11_ , P1_U4047 );
nand NAND2_1486 ( P1_U4084 , U122 , P1_U3086 );
nand NAND2_1487 ( P1_U4085 , P1_SUB_88_U8 , P1_U3029 );
nand NAND2_1488 ( P1_U4086 , P1_IR_REG_12_ , P1_U4047 );
nand NAND2_1489 ( P1_U4087 , U121 , P1_U3086 );
nand NAND2_1490 ( P1_U4088 , P1_SUB_88_U179 , P1_U3029 );
nand NAND2_1491 ( P1_U4089 , P1_IR_REG_13_ , P1_U4047 );
nand NAND2_1492 ( P1_U4090 , U120 , P1_U3086 );
nand NAND2_1493 ( P1_U4091 , P1_SUB_88_U9 , P1_U3029 );
nand NAND2_1494 ( P1_U4092 , P1_IR_REG_14_ , P1_U4047 );
nand NAND2_1495 ( P1_U4093 , U119 , P1_U3086 );
nand NAND2_1496 ( P1_U4094 , P1_SUB_88_U10 , P1_U3029 );
nand NAND2_1497 ( P1_U4095 , P1_IR_REG_15_ , P1_U4047 );
nand NAND2_1498 ( P1_U4096 , U118 , P1_U3086 );
nand NAND2_1499 ( P1_U4097 , P1_SUB_88_U11 , P1_U3029 );
nand NAND2_1500 ( P1_U4098 , P1_IR_REG_16_ , P1_U4047 );
nand NAND2_1501 ( P1_U4099 , U117 , P1_U3086 );
nand NAND2_1502 ( P1_U4100 , P1_SUB_88_U177 , P1_U3029 );
nand NAND2_1503 ( P1_U4101 , P1_IR_REG_17_ , P1_U4047 );
nand NAND2_1504 ( P1_U4102 , U116 , P1_U3086 );
nand NAND2_1505 ( P1_U4103 , P1_SUB_88_U12 , P1_U3029 );
nand NAND2_1506 ( P1_U4104 , P1_IR_REG_18_ , P1_U4047 );
nand NAND2_1507 ( P1_U4105 , U115 , P1_U3086 );
nand NAND2_1508 ( P1_U4106 , P1_SUB_88_U13 , P1_U3029 );
nand NAND2_1509 ( P1_U4107 , P1_IR_REG_19_ , P1_U4047 );
nand NAND2_1510 ( P1_U4108 , U113 , P1_U3086 );
nand NAND2_1511 ( P1_U4109 , P1_SUB_88_U14 , P1_U3029 );
nand NAND2_1512 ( P1_U4110 , P1_IR_REG_20_ , P1_U4047 );
nand NAND2_1513 ( P1_U4111 , U112 , P1_U3086 );
nand NAND2_1514 ( P1_U4112 , P1_SUB_88_U173 , P1_U3029 );
nand NAND2_1515 ( P1_U4113 , P1_IR_REG_21_ , P1_U4047 );
nand NAND2_1516 ( P1_U4114 , U111 , P1_U3086 );
nand NAND2_1517 ( P1_U4115 , P1_SUB_88_U15 , P1_U3029 );
nand NAND2_1518 ( P1_U4116 , P1_IR_REG_22_ , P1_U4047 );
nand NAND2_1519 ( P1_U4117 , U110 , P1_U3086 );
nand NAND2_1520 ( P1_U4118 , P1_SUB_88_U16 , P1_U3029 );
nand NAND2_1521 ( P1_U4119 , P1_IR_REG_23_ , P1_U4047 );
nand NAND2_1522 ( P1_U4120 , U109 , P1_U3086 );
nand NAND2_1523 ( P1_U4121 , P1_SUB_88_U17 , P1_U3029 );
nand NAND2_1524 ( P1_U4122 , P1_IR_REG_24_ , P1_U4047 );
nand NAND2_1525 ( P1_U4123 , U108 , P1_U3086 );
nand NAND2_1526 ( P1_U4124 , P1_SUB_88_U170 , P1_U3029 );
nand NAND2_1527 ( P1_U4125 , P1_IR_REG_25_ , P1_U4047 );
nand NAND2_1528 ( P1_U4126 , U107 , P1_U3086 );
nand NAND2_1529 ( P1_U4127 , P1_SUB_88_U18 , P1_U3029 );
nand NAND2_1530 ( P1_U4128 , P1_IR_REG_26_ , P1_U4047 );
nand NAND2_1531 ( P1_U4129 , U106 , P1_U3086 );
nand NAND2_1532 ( P1_U4130 , P1_SUB_88_U42 , P1_U3029 );
nand NAND2_1533 ( P1_U4131 , P1_IR_REG_27_ , P1_U4047 );
nand NAND2_1534 ( P1_U4132 , U105 , P1_U3086 );
nand NAND2_1535 ( P1_U4133 , P1_SUB_88_U19 , P1_U3029 );
nand NAND2_1536 ( P1_U4134 , P1_IR_REG_28_ , P1_U4047 );
nand NAND2_1537 ( P1_U4135 , U104 , P1_U3086 );
nand NAND2_1538 ( P1_U4136 , P1_SUB_88_U20 , P1_U3029 );
nand NAND2_1539 ( P1_U4137 , P1_IR_REG_29_ , P1_U4047 );
nand NAND2_1540 ( P1_U4138 , U102 , P1_U3086 );
nand NAND2_1541 ( P1_U4139 , P1_SUB_88_U165 , P1_U3029 );
nand NAND2_1542 ( P1_U4140 , P1_IR_REG_30_ , P1_U4047 );
nand NAND2_1543 ( P1_U4141 , U101 , P1_U3086 );
nand NAND2_1544 ( P1_U4142 , P1_SUB_88_U41 , P1_U3029 );
nand NAND2_1545 ( P1_U4143 , P1_IR_REG_31_ , P1_U4047 );
not NOT1_1546 ( P1_U4144 , P1_U3360 );
not NOT1_1547 ( P1_U4145 , P1_U3425 );
nand NAND2_1548 ( P1_U4146 , P1_U3358 , P1_U5775 );
nand NAND2_1549 ( P1_U4147 , P1_U3358 , P1_U5778 );
nand NAND2_1550 ( P1_U4148 , P1_U4144 , P1_D_REG_10_ );
nand NAND2_1551 ( P1_U4149 , P1_U4144 , P1_D_REG_11_ );
nand NAND2_1552 ( P1_U4150 , P1_U4144 , P1_D_REG_12_ );
nand NAND2_1553 ( P1_U4151 , P1_U4144 , P1_D_REG_13_ );
nand NAND2_1554 ( P1_U4152 , P1_U4144 , P1_D_REG_14_ );
nand NAND2_1555 ( P1_U4153 , P1_U4144 , P1_D_REG_15_ );
nand NAND2_1556 ( P1_U4154 , P1_U4144 , P1_D_REG_16_ );
nand NAND2_1557 ( P1_U4155 , P1_U4144 , P1_D_REG_17_ );
nand NAND2_1558 ( P1_U4156 , P1_U4144 , P1_D_REG_18_ );
nand NAND2_1559 ( P1_U4157 , P1_U4144 , P1_D_REG_19_ );
nand NAND2_1560 ( P1_U4158 , P1_U4144 , P1_D_REG_20_ );
nand NAND2_1561 ( P1_U4159 , P1_U4144 , P1_D_REG_21_ );
nand NAND2_1562 ( P1_U4160 , P1_U4144 , P1_D_REG_22_ );
nand NAND2_1563 ( P1_U4161 , P1_U4144 , P1_D_REG_23_ );
nand NAND2_1564 ( P1_U4162 , P1_U4144 , P1_D_REG_24_ );
nand NAND2_1565 ( P1_U4163 , P1_U4144 , P1_D_REG_25_ );
nand NAND2_1566 ( P1_U4164 , P1_U4144 , P1_D_REG_26_ );
nand NAND2_1567 ( P1_U4165 , P1_U4144 , P1_D_REG_27_ );
nand NAND2_1568 ( P1_U4166 , P1_U4144 , P1_D_REG_28_ );
nand NAND2_1569 ( P1_U4167 , P1_U4144 , P1_D_REG_29_ );
nand NAND2_1570 ( P1_U4168 , P1_U4144 , P1_D_REG_2_ );
nand NAND2_1571 ( P1_U4169 , P1_U4144 , P1_D_REG_30_ );
nand NAND2_1572 ( P1_U4170 , P1_U4144 , P1_D_REG_31_ );
nand NAND2_1573 ( P1_U4171 , P1_U4144 , P1_D_REG_3_ );
nand NAND2_1574 ( P1_U4172 , P1_U4144 , P1_D_REG_4_ );
nand NAND2_1575 ( P1_U4173 , P1_U4144 , P1_D_REG_5_ );
nand NAND2_1576 ( P1_U4174 , P1_U4144 , P1_D_REG_6_ );
nand NAND2_1577 ( P1_U4175 , P1_U4144 , P1_D_REG_7_ );
nand NAND2_1578 ( P1_U4176 , P1_U4144 , P1_D_REG_8_ );
nand NAND2_1579 ( P1_U4177 , P1_U4144 , P1_D_REG_9_ );
nand NAND2_1580 ( P1_U4178 , P1_U5802 , P1_U5799 );
nand NAND3_1581 ( P1_U4179 , P1_U5822 , P1_U5821 , P1_U3369 );
nand NAND2_1582 ( P1_U4180 , P1_U3018 , P1_REG2_REG_1_ );
nand NAND2_1583 ( P1_U4181 , P1_U3019 , P1_REG1_REG_1_ );
nand NAND2_1584 ( P1_U4182 , P1_U3020 , P1_REG0_REG_1_ );
nand NAND2_1585 ( P1_U4183 , P1_REG3_REG_1_ , P1_U3017 );
not NOT1_1586 ( P1_U4184 , P1_U3078 );
nand NAND2_1587 ( P1_U4185 , P1_U3419 , P1_U4010 );
nand NAND2_1588 ( P1_U4186 , P1_U4007 , P1_R1150_U21 );
nand NAND2_1589 ( P1_U4187 , P1_U4000 , P1_R1117_U21 );
nand NAND2_1590 ( P1_U4188 , P1_U3994 , P1_R1138_U96 );
nand NAND2_1591 ( P1_U4189 , P1_U4005 , P1_R1192_U21 );
nand NAND2_1592 ( P1_U4190 , P1_U4004 , P1_R1207_U21 );
nand NAND2_1593 ( P1_U4191 , P1_U4011 , P1_R1171_U96 );
nand NAND2_1594 ( P1_U4192 , P1_U3992 , P1_R1240_U96 );
not NOT1_1595 ( P1_U4193 , P1_U3376 );
nand NAND2_1596 ( P1_U4194 , P1_U3025 , P1_U3078 );
nand NAND2_1597 ( P1_U4195 , P1_R1222_U96 , P1_U3024 );
nand NAND2_1598 ( P1_U4196 , P1_U3456 , P1_U4036 );
nand NAND2_1599 ( P1_U4197 , P1_U3456 , P1_U4185 );
nand NAND4_1600 ( P1_U4198 , P1_U4197 , P1_U4194 , P1_U3595 , P1_U4193 );
nand NAND2_1601 ( P1_U4199 , P1_REG2_REG_2_ , P1_U3018 );
nand NAND2_1602 ( P1_U4200 , P1_REG1_REG_2_ , P1_U3019 );
nand NAND2_1603 ( P1_U4201 , P1_REG0_REG_2_ , P1_U3020 );
nand NAND2_1604 ( P1_U4202 , P1_REG3_REG_2_ , P1_U3017 );
not NOT1_1605 ( P1_U4203 , P1_U3068 );
nand NAND2_1606 ( P1_U4204 , P1_REG0_REG_0_ , P1_U3020 );
nand NAND2_1607 ( P1_U4205 , P1_REG1_REG_0_ , P1_U3019 );
nand NAND2_1608 ( P1_U4206 , P1_REG2_REG_0_ , P1_U3018 );
nand NAND2_1609 ( P1_U4207 , P1_REG3_REG_0_ , P1_U3017 );
not NOT1_1610 ( P1_U4208 , P1_U3077 );
nand NAND2_1611 ( P1_U4209 , P1_U3034 , P1_U3077 );
nand NAND2_1612 ( P1_U4210 , P1_R1150_U98 , P1_U4007 );
nand NAND2_1613 ( P1_U4211 , P1_R1117_U98 , P1_U4000 );
nand NAND2_1614 ( P1_U4212 , P1_R1138_U95 , P1_U3994 );
nand NAND2_1615 ( P1_U4213 , P1_R1192_U98 , P1_U4005 );
nand NAND2_1616 ( P1_U4214 , P1_R1207_U98 , P1_U4004 );
nand NAND2_1617 ( P1_U4215 , P1_R1171_U95 , P1_U4011 );
nand NAND2_1618 ( P1_U4216 , P1_R1240_U95 , P1_U3992 );
not NOT1_1619 ( P1_U4217 , P1_U3378 );
nand NAND2_1620 ( P1_U4218 , P1_U3025 , P1_U3068 );
nand NAND2_1621 ( P1_U4219 , P1_R1222_U95 , P1_U3024 );
nand NAND2_1622 ( P1_U4220 , P1_R1282_U56 , P1_U4036 );
nand NAND2_1623 ( P1_U4221 , P1_U3461 , P1_U4185 );
nand NAND2_1624 ( P1_U4222 , P1_U3611 , P1_U4217 );
nand NAND2_1625 ( P1_U4223 , P1_REG2_REG_3_ , P1_U3018 );
nand NAND2_1626 ( P1_U4224 , P1_REG1_REG_3_ , P1_U3019 );
nand NAND2_1627 ( P1_U4225 , P1_REG0_REG_3_ , P1_U3020 );
nand NAND2_1628 ( P1_U4226 , P1_ADD_99_U4 , P1_U3017 );
not NOT1_1629 ( P1_U4227 , P1_U3064 );
nand NAND2_1630 ( P1_U4228 , P1_U3034 , P1_U3078 );
nand NAND2_1631 ( P1_U4229 , P1_R1150_U108 , P1_U4007 );
nand NAND2_1632 ( P1_U4230 , P1_R1117_U108 , P1_U4000 );
nand NAND2_1633 ( P1_U4231 , P1_R1138_U17 , P1_U3994 );
nand NAND2_1634 ( P1_U4232 , P1_R1192_U108 , P1_U4005 );
nand NAND2_1635 ( P1_U4233 , P1_R1207_U108 , P1_U4004 );
nand NAND2_1636 ( P1_U4234 , P1_R1171_U17 , P1_U4011 );
nand NAND2_1637 ( P1_U4235 , P1_R1240_U17 , P1_U3992 );
not NOT1_1638 ( P1_U4236 , P1_U3379 );
nand NAND2_1639 ( P1_U4237 , P1_U3025 , P1_U3064 );
nand NAND2_1640 ( P1_U4238 , P1_R1222_U17 , P1_U3024 );
nand NAND2_1641 ( P1_U4239 , P1_R1282_U18 , P1_U4036 );
nand NAND2_1642 ( P1_U4240 , P1_U3464 , P1_U4185 );
nand NAND2_1643 ( P1_U4241 , P1_U3615 , P1_U4236 );
nand NAND2_1644 ( P1_U4242 , P1_REG2_REG_4_ , P1_U3018 );
nand NAND2_1645 ( P1_U4243 , P1_REG1_REG_4_ , P1_U3019 );
nand NAND2_1646 ( P1_U4244 , P1_REG0_REG_4_ , P1_U3020 );
nand NAND2_1647 ( P1_U4245 , P1_ADD_99_U59 , P1_U3017 );
not NOT1_1648 ( P1_U4246 , P1_U3060 );
nand NAND2_1649 ( P1_U4247 , P1_U3034 , P1_U3068 );
nand NAND2_1650 ( P1_U4248 , P1_R1150_U18 , P1_U4007 );
nand NAND2_1651 ( P1_U4249 , P1_R1117_U18 , P1_U4000 );
nand NAND2_1652 ( P1_U4250 , P1_R1138_U101 , P1_U3994 );
nand NAND2_1653 ( P1_U4251 , P1_R1192_U18 , P1_U4005 );
nand NAND2_1654 ( P1_U4252 , P1_R1207_U18 , P1_U4004 );
nand NAND2_1655 ( P1_U4253 , P1_R1171_U101 , P1_U4011 );
nand NAND2_1656 ( P1_U4254 , P1_R1240_U101 , P1_U3992 );
not NOT1_1657 ( P1_U4255 , P1_U3380 );
nand NAND2_1658 ( P1_U4256 , P1_U3025 , P1_U3060 );
nand NAND2_1659 ( P1_U4257 , P1_R1222_U101 , P1_U3024 );
nand NAND2_1660 ( P1_U4258 , P1_R1282_U20 , P1_U4036 );
nand NAND2_1661 ( P1_U4259 , P1_U3467 , P1_U4185 );
nand NAND2_1662 ( P1_U4260 , P1_U3619 , P1_U4255 );
nand NAND2_1663 ( P1_U4261 , P1_REG2_REG_5_ , P1_U3018 );
nand NAND2_1664 ( P1_U4262 , P1_REG1_REG_5_ , P1_U3019 );
nand NAND2_1665 ( P1_U4263 , P1_REG0_REG_5_ , P1_U3020 );
nand NAND2_1666 ( P1_U4264 , P1_ADD_99_U58 , P1_U3017 );
not NOT1_1667 ( P1_U4265 , P1_U3067 );
nand NAND2_1668 ( P1_U4266 , P1_U3034 , P1_U3064 );
nand NAND2_1669 ( P1_U4267 , P1_R1150_U107 , P1_U4007 );
nand NAND2_1670 ( P1_U4268 , P1_R1117_U107 , P1_U4000 );
nand NAND2_1671 ( P1_U4269 , P1_R1138_U100 , P1_U3994 );
nand NAND2_1672 ( P1_U4270 , P1_R1192_U107 , P1_U4005 );
nand NAND2_1673 ( P1_U4271 , P1_R1207_U107 , P1_U4004 );
nand NAND2_1674 ( P1_U4272 , P1_R1171_U100 , P1_U4011 );
nand NAND2_1675 ( P1_U4273 , P1_R1240_U100 , P1_U3992 );
not NOT1_1676 ( P1_U4274 , P1_U3381 );
nand NAND2_1677 ( P1_U4275 , P1_U3025 , P1_U3067 );
nand NAND2_1678 ( P1_U4276 , P1_R1222_U100 , P1_U3024 );
nand NAND2_1679 ( P1_U4277 , P1_R1282_U21 , P1_U4036 );
nand NAND2_1680 ( P1_U4278 , P1_U3470 , P1_U4185 );
nand NAND2_1681 ( P1_U4279 , P1_U3623 , P1_U4274 );
nand NAND2_1682 ( P1_U4280 , P1_REG2_REG_6_ , P1_U3018 );
nand NAND2_1683 ( P1_U4281 , P1_REG1_REG_6_ , P1_U3019 );
nand NAND2_1684 ( P1_U4282 , P1_REG0_REG_6_ , P1_U3020 );
nand NAND2_1685 ( P1_U4283 , P1_ADD_99_U57 , P1_U3017 );
not NOT1_1686 ( P1_U4284 , P1_U3071 );
nand NAND2_1687 ( P1_U4285 , P1_U3034 , P1_U3060 );
nand NAND2_1688 ( P1_U4286 , P1_R1150_U106 , P1_U4007 );
nand NAND2_1689 ( P1_U4287 , P1_R1117_U106 , P1_U4000 );
nand NAND2_1690 ( P1_U4288 , P1_R1138_U18 , P1_U3994 );
nand NAND2_1691 ( P1_U4289 , P1_R1192_U106 , P1_U4005 );
nand NAND2_1692 ( P1_U4290 , P1_R1207_U106 , P1_U4004 );
nand NAND2_1693 ( P1_U4291 , P1_R1171_U18 , P1_U4011 );
nand NAND2_1694 ( P1_U4292 , P1_R1240_U18 , P1_U3992 );
not NOT1_1695 ( P1_U4293 , P1_U3382 );
nand NAND2_1696 ( P1_U4294 , P1_U3025 , P1_U3071 );
nand NAND2_1697 ( P1_U4295 , P1_R1222_U18 , P1_U3024 );
nand NAND2_1698 ( P1_U4296 , P1_R1282_U65 , P1_U4036 );
nand NAND2_1699 ( P1_U4297 , P1_U3473 , P1_U4185 );
nand NAND2_1700 ( P1_U4298 , P1_U3627 , P1_U4293 );
nand NAND2_1701 ( P1_U4299 , P1_REG2_REG_7_ , P1_U3018 );
nand NAND2_1702 ( P1_U4300 , P1_REG1_REG_7_ , P1_U3019 );
nand NAND2_1703 ( P1_U4301 , P1_REG0_REG_7_ , P1_U3020 );
nand NAND2_1704 ( P1_U4302 , P1_ADD_99_U56 , P1_U3017 );
not NOT1_1705 ( P1_U4303 , P1_U3070 );
nand NAND2_1706 ( P1_U4304 , P1_U3034 , P1_U3067 );
nand NAND2_1707 ( P1_U4305 , P1_R1150_U19 , P1_U4007 );
nand NAND2_1708 ( P1_U4306 , P1_R1117_U19 , P1_U4000 );
nand NAND2_1709 ( P1_U4307 , P1_R1138_U99 , P1_U3994 );
nand NAND2_1710 ( P1_U4308 , P1_R1192_U19 , P1_U4005 );
nand NAND2_1711 ( P1_U4309 , P1_R1207_U19 , P1_U4004 );
nand NAND2_1712 ( P1_U4310 , P1_R1171_U99 , P1_U4011 );
nand NAND2_1713 ( P1_U4311 , P1_R1240_U99 , P1_U3992 );
not NOT1_1714 ( P1_U4312 , P1_U3383 );
nand NAND2_1715 ( P1_U4313 , P1_U3025 , P1_U3070 );
nand NAND2_1716 ( P1_U4314 , P1_R1222_U99 , P1_U3024 );
nand NAND2_1717 ( P1_U4315 , P1_R1282_U22 , P1_U4036 );
nand NAND2_1718 ( P1_U4316 , P1_U3476 , P1_U4185 );
nand NAND2_1719 ( P1_U4317 , P1_U3631 , P1_U4312 );
nand NAND2_1720 ( P1_U4318 , P1_REG2_REG_8_ , P1_U3018 );
nand NAND2_1721 ( P1_U4319 , P1_REG1_REG_8_ , P1_U3019 );
nand NAND2_1722 ( P1_U4320 , P1_REG0_REG_8_ , P1_U3020 );
nand NAND2_1723 ( P1_U4321 , P1_ADD_99_U55 , P1_U3017 );
not NOT1_1724 ( P1_U4322 , P1_U3084 );
nand NAND2_1725 ( P1_U4323 , P1_U3034 , P1_U3071 );
nand NAND2_1726 ( P1_U4324 , P1_R1150_U105 , P1_U4007 );
nand NAND2_1727 ( P1_U4325 , P1_R1117_U105 , P1_U4000 );
nand NAND2_1728 ( P1_U4326 , P1_R1138_U19 , P1_U3994 );
nand NAND2_1729 ( P1_U4327 , P1_R1192_U105 , P1_U4005 );
nand NAND2_1730 ( P1_U4328 , P1_R1207_U105 , P1_U4004 );
nand NAND2_1731 ( P1_U4329 , P1_R1171_U19 , P1_U4011 );
nand NAND2_1732 ( P1_U4330 , P1_R1240_U19 , P1_U3992 );
not NOT1_1733 ( P1_U4331 , P1_U3384 );
nand NAND2_1734 ( P1_U4332 , P1_U3025 , P1_U3084 );
nand NAND2_1735 ( P1_U4333 , P1_R1222_U19 , P1_U3024 );
nand NAND2_1736 ( P1_U4334 , P1_R1282_U23 , P1_U4036 );
nand NAND2_1737 ( P1_U4335 , P1_U3479 , P1_U4185 );
nand NAND2_1738 ( P1_U4336 , P1_U3635 , P1_U4331 );
nand NAND2_1739 ( P1_U4337 , P1_REG2_REG_9_ , P1_U3018 );
nand NAND2_1740 ( P1_U4338 , P1_REG1_REG_9_ , P1_U3019 );
nand NAND2_1741 ( P1_U4339 , P1_REG0_REG_9_ , P1_U3020 );
nand NAND2_1742 ( P1_U4340 , P1_ADD_99_U54 , P1_U3017 );
not NOT1_1743 ( P1_U4341 , P1_U3083 );
nand NAND2_1744 ( P1_U4342 , P1_U3034 , P1_U3070 );
nand NAND2_1745 ( P1_U4343 , P1_R1150_U20 , P1_U4007 );
nand NAND2_1746 ( P1_U4344 , P1_R1117_U20 , P1_U4000 );
nand NAND2_1747 ( P1_U4345 , P1_R1138_U98 , P1_U3994 );
nand NAND2_1748 ( P1_U4346 , P1_R1192_U20 , P1_U4005 );
nand NAND2_1749 ( P1_U4347 , P1_R1207_U20 , P1_U4004 );
nand NAND2_1750 ( P1_U4348 , P1_R1171_U98 , P1_U4011 );
nand NAND2_1751 ( P1_U4349 , P1_R1240_U98 , P1_U3992 );
not NOT1_1752 ( P1_U4350 , P1_U3385 );
nand NAND2_1753 ( P1_U4351 , P1_U3025 , P1_U3083 );
nand NAND2_1754 ( P1_U4352 , P1_R1222_U98 , P1_U3024 );
nand NAND2_1755 ( P1_U4353 , P1_R1282_U24 , P1_U4036 );
nand NAND2_1756 ( P1_U4354 , P1_U3482 , P1_U4185 );
nand NAND2_1757 ( P1_U4355 , P1_U3639 , P1_U4350 );
nand NAND2_1758 ( P1_U4356 , P1_REG2_REG_10_ , P1_U3018 );
nand NAND2_1759 ( P1_U4357 , P1_REG1_REG_10_ , P1_U3019 );
nand NAND2_1760 ( P1_U4358 , P1_REG0_REG_10_ , P1_U3020 );
nand NAND2_1761 ( P1_U4359 , P1_ADD_99_U78 , P1_U3017 );
not NOT1_1762 ( P1_U4360 , P1_U3062 );
nand NAND2_1763 ( P1_U4361 , P1_U3034 , P1_U3084 );
nand NAND2_1764 ( P1_U4362 , P1_R1150_U104 , P1_U4007 );
nand NAND2_1765 ( P1_U4363 , P1_R1117_U104 , P1_U4000 );
nand NAND2_1766 ( P1_U4364 , P1_R1138_U97 , P1_U3994 );
nand NAND2_1767 ( P1_U4365 , P1_R1192_U104 , P1_U4005 );
nand NAND2_1768 ( P1_U4366 , P1_R1207_U104 , P1_U4004 );
nand NAND2_1769 ( P1_U4367 , P1_R1171_U97 , P1_U4011 );
nand NAND2_1770 ( P1_U4368 , P1_R1240_U97 , P1_U3992 );
not NOT1_1771 ( P1_U4369 , P1_U3386 );
nand NAND2_1772 ( P1_U4370 , P1_U3025 , P1_U3062 );
nand NAND2_1773 ( P1_U4371 , P1_R1222_U97 , P1_U3024 );
nand NAND2_1774 ( P1_U4372 , P1_R1282_U63 , P1_U4036 );
nand NAND2_1775 ( P1_U4373 , P1_U3485 , P1_U4185 );
nand NAND2_1776 ( P1_U4374 , P1_U3643 , P1_U4369 );
nand NAND2_1777 ( P1_U4375 , P1_REG2_REG_11_ , P1_U3018 );
nand NAND2_1778 ( P1_U4376 , P1_REG1_REG_11_ , P1_U3019 );
nand NAND2_1779 ( P1_U4377 , P1_REG0_REG_11_ , P1_U3020 );
nand NAND2_1780 ( P1_U4378 , P1_ADD_99_U77 , P1_U3017 );
not NOT1_1781 ( P1_U4379 , P1_U3063 );
nand NAND2_1782 ( P1_U4380 , P1_U3034 , P1_U3083 );
nand NAND2_1783 ( P1_U4381 , P1_R1150_U114 , P1_U4007 );
nand NAND2_1784 ( P1_U4382 , P1_R1117_U114 , P1_U4000 );
nand NAND2_1785 ( P1_U4383 , P1_R1138_U11 , P1_U3994 );
nand NAND2_1786 ( P1_U4384 , P1_R1192_U114 , P1_U4005 );
nand NAND2_1787 ( P1_U4385 , P1_R1207_U114 , P1_U4004 );
nand NAND2_1788 ( P1_U4386 , P1_R1171_U11 , P1_U4011 );
nand NAND2_1789 ( P1_U4387 , P1_R1240_U11 , P1_U3992 );
not NOT1_1790 ( P1_U4388 , P1_U3387 );
nand NAND2_1791 ( P1_U4389 , P1_U3025 , P1_U3063 );
nand NAND2_1792 ( P1_U4390 , P1_R1222_U11 , P1_U3024 );
nand NAND2_1793 ( P1_U4391 , P1_R1282_U6 , P1_U4036 );
nand NAND2_1794 ( P1_U4392 , P1_U3488 , P1_U4185 );
nand NAND2_1795 ( P1_U4393 , P1_U3647 , P1_U4388 );
nand NAND2_1796 ( P1_U4394 , P1_REG2_REG_12_ , P1_U3018 );
nand NAND2_1797 ( P1_U4395 , P1_REG1_REG_12_ , P1_U3019 );
nand NAND2_1798 ( P1_U4396 , P1_REG0_REG_12_ , P1_U3020 );
nand NAND2_1799 ( P1_U4397 , P1_ADD_99_U76 , P1_U3017 );
not NOT1_1800 ( P1_U4398 , P1_U3072 );
nand NAND2_1801 ( P1_U4399 , P1_U3034 , P1_U3062 );
nand NAND2_1802 ( P1_U4400 , P1_R1150_U13 , P1_U4007 );
nand NAND2_1803 ( P1_U4401 , P1_R1117_U13 , P1_U4000 );
nand NAND2_1804 ( P1_U4402 , P1_R1138_U115 , P1_U3994 );
nand NAND2_1805 ( P1_U4403 , P1_R1192_U13 , P1_U4005 );
nand NAND2_1806 ( P1_U4404 , P1_R1207_U13 , P1_U4004 );
nand NAND2_1807 ( P1_U4405 , P1_R1171_U115 , P1_U4011 );
nand NAND2_1808 ( P1_U4406 , P1_R1240_U115 , P1_U3992 );
not NOT1_1809 ( P1_U4407 , P1_U3388 );
nand NAND2_1810 ( P1_U4408 , P1_U3025 , P1_U3072 );
nand NAND2_1811 ( P1_U4409 , P1_R1222_U115 , P1_U3024 );
nand NAND2_1812 ( P1_U4410 , P1_R1282_U7 , P1_U4036 );
nand NAND2_1813 ( P1_U4411 , P1_U3491 , P1_U4185 );
nand NAND2_1814 ( P1_U4412 , P1_U3651 , P1_U4407 );
nand NAND2_1815 ( P1_U4413 , P1_REG2_REG_13_ , P1_U3018 );
nand NAND2_1816 ( P1_U4414 , P1_REG1_REG_13_ , P1_U3019 );
nand NAND2_1817 ( P1_U4415 , P1_REG0_REG_13_ , P1_U3020 );
nand NAND2_1818 ( P1_U4416 , P1_ADD_99_U75 , P1_U3017 );
not NOT1_1819 ( P1_U4417 , P1_U3080 );
nand NAND2_1820 ( P1_U4418 , P1_U3034 , P1_U3063 );
nand NAND2_1821 ( P1_U4419 , P1_R1150_U103 , P1_U4007 );
nand NAND2_1822 ( P1_U4420 , P1_R1117_U103 , P1_U4000 );
nand NAND2_1823 ( P1_U4421 , P1_R1138_U114 , P1_U3994 );
nand NAND2_1824 ( P1_U4422 , P1_R1192_U103 , P1_U4005 );
nand NAND2_1825 ( P1_U4423 , P1_R1207_U103 , P1_U4004 );
nand NAND2_1826 ( P1_U4424 , P1_R1171_U114 , P1_U4011 );
nand NAND2_1827 ( P1_U4425 , P1_R1240_U114 , P1_U3992 );
not NOT1_1828 ( P1_U4426 , P1_U3389 );
nand NAND2_1829 ( P1_U4427 , P1_U3025 , P1_U3080 );
nand NAND2_1830 ( P1_U4428 , P1_R1222_U114 , P1_U3024 );
nand NAND2_1831 ( P1_U4429 , P1_R1282_U8 , P1_U4036 );
nand NAND2_1832 ( P1_U4430 , P1_U3494 , P1_U4185 );
nand NAND2_1833 ( P1_U4431 , P1_U3655 , P1_U4426 );
nand NAND2_1834 ( P1_U4432 , P1_REG2_REG_14_ , P1_U3018 );
nand NAND2_1835 ( P1_U4433 , P1_REG1_REG_14_ , P1_U3019 );
nand NAND2_1836 ( P1_U4434 , P1_REG0_REG_14_ , P1_U3020 );
nand NAND2_1837 ( P1_U4435 , P1_ADD_99_U74 , P1_U3017 );
not NOT1_1838 ( P1_U4436 , P1_U3079 );
nand NAND2_1839 ( P1_U4437 , P1_U3034 , P1_U3072 );
nand NAND2_1840 ( P1_U4438 , P1_R1150_U102 , P1_U4007 );
nand NAND2_1841 ( P1_U4439 , P1_R1117_U102 , P1_U4000 );
nand NAND2_1842 ( P1_U4440 , P1_R1138_U12 , P1_U3994 );
nand NAND2_1843 ( P1_U4441 , P1_R1192_U102 , P1_U4005 );
nand NAND2_1844 ( P1_U4442 , P1_R1207_U102 , P1_U4004 );
nand NAND2_1845 ( P1_U4443 , P1_R1171_U12 , P1_U4011 );
nand NAND2_1846 ( P1_U4444 , P1_R1240_U12 , P1_U3992 );
not NOT1_1847 ( P1_U4445 , P1_U3390 );
nand NAND2_1848 ( P1_U4446 , P1_U3025 , P1_U3079 );
nand NAND2_1849 ( P1_U4447 , P1_R1222_U12 , P1_U3024 );
nand NAND2_1850 ( P1_U4448 , P1_R1282_U86 , P1_U4036 );
nand NAND2_1851 ( P1_U4449 , P1_U3497 , P1_U4185 );
nand NAND2_1852 ( P1_U4450 , P1_U3659 , P1_U4445 );
nand NAND2_1853 ( P1_U4451 , P1_REG2_REG_15_ , P1_U3018 );
nand NAND2_1854 ( P1_U4452 , P1_REG1_REG_15_ , P1_U3019 );
nand NAND2_1855 ( P1_U4453 , P1_REG0_REG_15_ , P1_U3020 );
nand NAND2_1856 ( P1_U4454 , P1_ADD_99_U73 , P1_U3017 );
not NOT1_1857 ( P1_U4455 , P1_U3074 );
nand NAND2_1858 ( P1_U4456 , P1_U3034 , P1_U3080 );
nand NAND2_1859 ( P1_U4457 , P1_R1150_U113 , P1_U4007 );
nand NAND2_1860 ( P1_U4458 , P1_R1117_U113 , P1_U4000 );
nand NAND2_1861 ( P1_U4459 , P1_R1138_U113 , P1_U3994 );
nand NAND2_1862 ( P1_U4460 , P1_R1192_U113 , P1_U4005 );
nand NAND2_1863 ( P1_U4461 , P1_R1207_U113 , P1_U4004 );
nand NAND2_1864 ( P1_U4462 , P1_R1171_U113 , P1_U4011 );
nand NAND2_1865 ( P1_U4463 , P1_R1240_U113 , P1_U3992 );
not NOT1_1866 ( P1_U4464 , P1_U3391 );
nand NAND2_1867 ( P1_U4465 , P1_U3025 , P1_U3074 );
nand NAND2_1868 ( P1_U4466 , P1_R1222_U113 , P1_U3024 );
nand NAND2_1869 ( P1_U4467 , P1_R1282_U9 , P1_U4036 );
nand NAND2_1870 ( P1_U4468 , P1_U3500 , P1_U4185 );
nand NAND2_1871 ( P1_U4469 , P1_U3663 , P1_U4464 );
nand NAND2_1872 ( P1_U4470 , P1_REG2_REG_16_ , P1_U3018 );
nand NAND2_1873 ( P1_U4471 , P1_REG1_REG_16_ , P1_U3019 );
nand NAND2_1874 ( P1_U4472 , P1_REG0_REG_16_ , P1_U3020 );
nand NAND2_1875 ( P1_U4473 , P1_ADD_99_U72 , P1_U3017 );
not NOT1_1876 ( P1_U4474 , P1_U3073 );
nand NAND2_1877 ( P1_U4475 , P1_U3034 , P1_U3079 );
nand NAND2_1878 ( P1_U4476 , P1_R1150_U112 , P1_U4007 );
nand NAND2_1879 ( P1_U4477 , P1_R1117_U112 , P1_U4000 );
nand NAND2_1880 ( P1_U4478 , P1_R1138_U112 , P1_U3994 );
nand NAND2_1881 ( P1_U4479 , P1_R1192_U112 , P1_U4005 );
nand NAND2_1882 ( P1_U4480 , P1_R1207_U112 , P1_U4004 );
nand NAND2_1883 ( P1_U4481 , P1_R1171_U112 , P1_U4011 );
nand NAND2_1884 ( P1_U4482 , P1_R1240_U112 , P1_U3992 );
not NOT1_1885 ( P1_U4483 , P1_U3392 );
nand NAND2_1886 ( P1_U4484 , P1_U3025 , P1_U3073 );
nand NAND2_1887 ( P1_U4485 , P1_R1222_U112 , P1_U3024 );
nand NAND2_1888 ( P1_U4486 , P1_R1282_U10 , P1_U4036 );
nand NAND2_1889 ( P1_U4487 , P1_U3503 , P1_U4185 );
nand NAND2_1890 ( P1_U4488 , P1_U3667 , P1_U4483 );
nand NAND2_1891 ( P1_U4489 , P1_REG2_REG_17_ , P1_U3018 );
nand NAND2_1892 ( P1_U4490 , P1_REG1_REG_17_ , P1_U3019 );
nand NAND2_1893 ( P1_U4491 , P1_REG0_REG_17_ , P1_U3020 );
nand NAND2_1894 ( P1_U4492 , P1_ADD_99_U71 , P1_U3017 );
not NOT1_1895 ( P1_U4493 , P1_U3069 );
nand NAND2_1896 ( P1_U4494 , P1_U3034 , P1_U3074 );
nand NAND2_1897 ( P1_U4495 , P1_R1150_U14 , P1_U4007 );
nand NAND2_1898 ( P1_U4496 , P1_R1117_U14 , P1_U4000 );
nand NAND2_1899 ( P1_U4497 , P1_R1138_U111 , P1_U3994 );
nand NAND2_1900 ( P1_U4498 , P1_R1192_U14 , P1_U4005 );
nand NAND2_1901 ( P1_U4499 , P1_R1207_U14 , P1_U4004 );
nand NAND2_1902 ( P1_U4500 , P1_R1171_U111 , P1_U4011 );
nand NAND2_1903 ( P1_U4501 , P1_R1240_U111 , P1_U3992 );
not NOT1_1904 ( P1_U4502 , P1_U3393 );
nand NAND2_1905 ( P1_U4503 , P1_U3025 , P1_U3069 );
nand NAND2_1906 ( P1_U4504 , P1_R1222_U111 , P1_U3024 );
nand NAND2_1907 ( P1_U4505 , P1_R1282_U11 , P1_U4036 );
nand NAND2_1908 ( P1_U4506 , P1_U3506 , P1_U4185 );
nand NAND2_1909 ( P1_U4507 , P1_U3671 , P1_U4502 );
nand NAND2_1910 ( P1_U4508 , P1_REG2_REG_18_ , P1_U3018 );
nand NAND2_1911 ( P1_U4509 , P1_REG1_REG_18_ , P1_U3019 );
nand NAND2_1912 ( P1_U4510 , P1_REG0_REG_18_ , P1_U3020 );
nand NAND2_1913 ( P1_U4511 , P1_ADD_99_U70 , P1_U3017 );
not NOT1_1914 ( P1_U4512 , P1_U3082 );
nand NAND2_1915 ( P1_U4513 , P1_U3034 , P1_U3073 );
nand NAND2_1916 ( P1_U4514 , P1_R1150_U101 , P1_U4007 );
nand NAND2_1917 ( P1_U4515 , P1_R1117_U101 , P1_U4000 );
nand NAND2_1918 ( P1_U4516 , P1_R1138_U13 , P1_U3994 );
nand NAND2_1919 ( P1_U4517 , P1_R1192_U101 , P1_U4005 );
nand NAND2_1920 ( P1_U4518 , P1_R1207_U101 , P1_U4004 );
nand NAND2_1921 ( P1_U4519 , P1_R1171_U13 , P1_U4011 );
nand NAND2_1922 ( P1_U4520 , P1_R1240_U13 , P1_U3992 );
not NOT1_1923 ( P1_U4521 , P1_U3394 );
nand NAND2_1924 ( P1_U4522 , P1_U3025 , P1_U3082 );
nand NAND2_1925 ( P1_U4523 , P1_R1222_U13 , P1_U3024 );
nand NAND2_1926 ( P1_U4524 , P1_R1282_U84 , P1_U4036 );
nand NAND2_1927 ( P1_U4525 , P1_U3509 , P1_U4185 );
nand NAND2_1928 ( P1_U4526 , P1_U3675 , P1_U4521 );
nand NAND2_1929 ( P1_U4527 , P1_REG2_REG_19_ , P1_U3018 );
nand NAND2_1930 ( P1_U4528 , P1_REG1_REG_19_ , P1_U3019 );
nand NAND2_1931 ( P1_U4529 , P1_REG0_REG_19_ , P1_U3020 );
nand NAND2_1932 ( P1_U4530 , P1_ADD_99_U69 , P1_U3017 );
not NOT1_1933 ( P1_U4531 , P1_U3081 );
nand NAND2_1934 ( P1_U4532 , P1_U3034 , P1_U3069 );
nand NAND2_1935 ( P1_U4533 , P1_R1150_U100 , P1_U4007 );
nand NAND2_1936 ( P1_U4534 , P1_R1117_U100 , P1_U4000 );
nand NAND2_1937 ( P1_U4535 , P1_R1138_U110 , P1_U3994 );
nand NAND2_1938 ( P1_U4536 , P1_R1192_U100 , P1_U4005 );
nand NAND2_1939 ( P1_U4537 , P1_R1207_U100 , P1_U4004 );
nand NAND2_1940 ( P1_U4538 , P1_R1171_U110 , P1_U4011 );
nand NAND2_1941 ( P1_U4539 , P1_R1240_U110 , P1_U3992 );
not NOT1_1942 ( P1_U4540 , P1_U3395 );
nand NAND2_1943 ( P1_U4541 , P1_U3025 , P1_U3081 );
nand NAND2_1944 ( P1_U4542 , P1_R1222_U110 , P1_U3024 );
nand NAND2_1945 ( P1_U4543 , P1_R1282_U12 , P1_U4036 );
nand NAND2_1946 ( P1_U4544 , P1_U3512 , P1_U4185 );
nand NAND2_1947 ( P1_U4545 , P1_U3679 , P1_U4540 );
nand NAND2_1948 ( P1_U4546 , P1_REG2_REG_20_ , P1_U3018 );
nand NAND2_1949 ( P1_U4547 , P1_REG1_REG_20_ , P1_U3019 );
nand NAND2_1950 ( P1_U4548 , P1_REG0_REG_20_ , P1_U3020 );
nand NAND2_1951 ( P1_U4549 , P1_ADD_99_U68 , P1_U3017 );
not NOT1_1952 ( P1_U4550 , P1_U3076 );
nand NAND2_1953 ( P1_U4551 , P1_U3034 , P1_U3082 );
nand NAND2_1954 ( P1_U4552 , P1_R1150_U99 , P1_U4007 );
nand NAND2_1955 ( P1_U4553 , P1_R1117_U99 , P1_U4000 );
nand NAND2_1956 ( P1_U4554 , P1_R1138_U109 , P1_U3994 );
nand NAND2_1957 ( P1_U4555 , P1_R1192_U99 , P1_U4005 );
nand NAND2_1958 ( P1_U4556 , P1_R1207_U99 , P1_U4004 );
nand NAND2_1959 ( P1_U4557 , P1_R1171_U109 , P1_U4011 );
nand NAND2_1960 ( P1_U4558 , P1_R1240_U109 , P1_U3992 );
not NOT1_1961 ( P1_U4559 , P1_U3396 );
nand NAND2_1962 ( P1_U4560 , P1_U3025 , P1_U3076 );
nand NAND2_1963 ( P1_U4561 , P1_R1222_U109 , P1_U3024 );
nand NAND2_1964 ( P1_U4562 , P1_R1282_U82 , P1_U4036 );
nand NAND2_1965 ( P1_U4563 , P1_U3514 , P1_U4185 );
nand NAND2_1966 ( P1_U4564 , P1_U3683 , P1_U4559 );
nand NAND2_1967 ( P1_U4565 , P1_REG2_REG_21_ , P1_U3018 );
nand NAND2_1968 ( P1_U4566 , P1_REG1_REG_21_ , P1_U3019 );
nand NAND2_1969 ( P1_U4567 , P1_REG0_REG_21_ , P1_U3020 );
nand NAND2_1970 ( P1_U4568 , P1_ADD_99_U67 , P1_U3017 );
not NOT1_1971 ( P1_U4569 , P1_U3075 );
nand NAND2_1972 ( P1_U4570 , P1_U3034 , P1_U3081 );
nand NAND2_1973 ( P1_U4571 , P1_R1150_U97 , P1_U4007 );
nand NAND2_1974 ( P1_U4572 , P1_R1117_U97 , P1_U4000 );
nand NAND2_1975 ( P1_U4573 , P1_R1138_U14 , P1_U3994 );
nand NAND2_1976 ( P1_U4574 , P1_R1192_U97 , P1_U4005 );
nand NAND2_1977 ( P1_U4575 , P1_R1207_U97 , P1_U4004 );
nand NAND2_1978 ( P1_U4576 , P1_R1171_U14 , P1_U4011 );
nand NAND2_1979 ( P1_U4577 , P1_R1240_U14 , P1_U3992 );
not NOT1_1980 ( P1_U4578 , P1_U3398 );
nand NAND2_1981 ( P1_U4579 , P1_U3025 , P1_U3075 );
nand NAND2_1982 ( P1_U4580 , P1_R1222_U14 , P1_U3024 );
nand NAND2_1983 ( P1_U4581 , P1_R1282_U13 , P1_U4036 );
nand NAND2_1984 ( P1_U4582 , P1_U4025 , P1_U4185 );
nand NAND2_1985 ( P1_U4583 , P1_U3687 , P1_U4578 );
nand NAND2_1986 ( P1_U4584 , P1_REG2_REG_22_ , P1_U3018 );
nand NAND2_1987 ( P1_U4585 , P1_REG1_REG_22_ , P1_U3019 );
nand NAND2_1988 ( P1_U4586 , P1_REG0_REG_22_ , P1_U3020 );
nand NAND2_1989 ( P1_U4587 , P1_ADD_99_U66 , P1_U3017 );
not NOT1_1990 ( P1_U4588 , P1_U3061 );
nand NAND2_1991 ( P1_U4589 , P1_U3034 , P1_U3076 );
nand NAND2_1992 ( P1_U4590 , P1_R1150_U111 , P1_U4007 );
nand NAND2_1993 ( P1_U4591 , P1_R1117_U111 , P1_U4000 );
nand NAND2_1994 ( P1_U4592 , P1_R1138_U15 , P1_U3994 );
nand NAND2_1995 ( P1_U4593 , P1_R1192_U111 , P1_U4005 );
nand NAND2_1996 ( P1_U4594 , P1_R1207_U111 , P1_U4004 );
nand NAND2_1997 ( P1_U4595 , P1_R1171_U15 , P1_U4011 );
nand NAND2_1998 ( P1_U4596 , P1_R1240_U15 , P1_U3992 );
not NOT1_1999 ( P1_U4597 , P1_U3400 );
nand NAND2_2000 ( P1_U4598 , P1_U3025 , P1_U3061 );
nand NAND2_2001 ( P1_U4599 , P1_R1222_U15 , P1_U3024 );
nand NAND2_2002 ( P1_U4600 , P1_R1282_U78 , P1_U4036 );
nand NAND2_2003 ( P1_U4601 , P1_U4024 , P1_U4185 );
nand NAND2_2004 ( P1_U4602 , P1_U3691 , P1_U4597 );
nand NAND2_2005 ( P1_U4603 , P1_REG2_REG_23_ , P1_U3018 );
nand NAND2_2006 ( P1_U4604 , P1_REG1_REG_23_ , P1_U3019 );
nand NAND2_2007 ( P1_U4605 , P1_REG0_REG_23_ , P1_U3020 );
nand NAND2_2008 ( P1_U4606 , P1_ADD_99_U65 , P1_U3017 );
not NOT1_2009 ( P1_U4607 , P1_U3066 );
nand NAND2_2010 ( P1_U4608 , P1_U3034 , P1_U3075 );
nand NAND2_2011 ( P1_U4609 , P1_R1150_U110 , P1_U4007 );
nand NAND2_2012 ( P1_U4610 , P1_R1117_U110 , P1_U4000 );
nand NAND2_2013 ( P1_U4611 , P1_R1138_U108 , P1_U3994 );
nand NAND2_2014 ( P1_U4612 , P1_R1192_U110 , P1_U4005 );
nand NAND2_2015 ( P1_U4613 , P1_R1207_U110 , P1_U4004 );
nand NAND2_2016 ( P1_U4614 , P1_R1171_U108 , P1_U4011 );
nand NAND2_2017 ( P1_U4615 , P1_R1240_U108 , P1_U3992 );
not NOT1_2018 ( P1_U4616 , P1_U3402 );
nand NAND2_2019 ( P1_U4617 , P1_U3025 , P1_U3066 );
nand NAND2_2020 ( P1_U4618 , P1_R1222_U108 , P1_U3024 );
nand NAND2_2021 ( P1_U4619 , P1_R1282_U14 , P1_U4036 );
nand NAND2_2022 ( P1_U4620 , P1_U4023 , P1_U4185 );
nand NAND2_2023 ( P1_U4621 , P1_U3695 , P1_U4616 );
nand NAND2_2024 ( P1_U4622 , P1_REG2_REG_24_ , P1_U3018 );
nand NAND2_2025 ( P1_U4623 , P1_REG1_REG_24_ , P1_U3019 );
nand NAND2_2026 ( P1_U4624 , P1_REG0_REG_24_ , P1_U3020 );
nand NAND2_2027 ( P1_U4625 , P1_ADD_99_U64 , P1_U3017 );
not NOT1_2028 ( P1_U4626 , P1_U3065 );
nand NAND2_2029 ( P1_U4627 , P1_U3034 , P1_U3061 );
nand NAND2_2030 ( P1_U4628 , P1_R1150_U15 , P1_U4007 );
nand NAND2_2031 ( P1_U4629 , P1_R1117_U15 , P1_U4000 );
nand NAND2_2032 ( P1_U4630 , P1_R1138_U107 , P1_U3994 );
nand NAND2_2033 ( P1_U4631 , P1_R1192_U15 , P1_U4005 );
nand NAND2_2034 ( P1_U4632 , P1_R1207_U15 , P1_U4004 );
nand NAND2_2035 ( P1_U4633 , P1_R1171_U107 , P1_U4011 );
nand NAND2_2036 ( P1_U4634 , P1_R1240_U107 , P1_U3992 );
not NOT1_2037 ( P1_U4635 , P1_U3404 );
nand NAND2_2038 ( P1_U4636 , P1_U3025 , P1_U3065 );
nand NAND2_2039 ( P1_U4637 , P1_R1222_U107 , P1_U3024 );
nand NAND2_2040 ( P1_U4638 , P1_R1282_U76 , P1_U4036 );
nand NAND2_2041 ( P1_U4639 , P1_U4022 , P1_U4185 );
nand NAND2_2042 ( P1_U4640 , P1_U3699 , P1_U4635 );
nand NAND2_2043 ( P1_U4641 , P1_REG2_REG_25_ , P1_U3018 );
nand NAND2_2044 ( P1_U4642 , P1_REG1_REG_25_ , P1_U3019 );
nand NAND2_2045 ( P1_U4643 , P1_REG0_REG_25_ , P1_U3020 );
nand NAND2_2046 ( P1_U4644 , P1_ADD_99_U63 , P1_U3017 );
not NOT1_2047 ( P1_U4645 , P1_U3058 );
nand NAND2_2048 ( P1_U4646 , P1_U3034 , P1_U3066 );
nand NAND2_2049 ( P1_U4647 , P1_R1150_U96 , P1_U4007 );
nand NAND2_2050 ( P1_U4648 , P1_R1117_U96 , P1_U4000 );
nand NAND2_2051 ( P1_U4649 , P1_R1138_U106 , P1_U3994 );
nand NAND2_2052 ( P1_U4650 , P1_R1192_U96 , P1_U4005 );
nand NAND2_2053 ( P1_U4651 , P1_R1207_U96 , P1_U4004 );
nand NAND2_2054 ( P1_U4652 , P1_R1171_U106 , P1_U4011 );
nand NAND2_2055 ( P1_U4653 , P1_R1240_U106 , P1_U3992 );
not NOT1_2056 ( P1_U4654 , P1_U3406 );
nand NAND2_2057 ( P1_U4655 , P1_U3025 , P1_U3058 );
nand NAND2_2058 ( P1_U4656 , P1_R1222_U106 , P1_U3024 );
nand NAND2_2059 ( P1_U4657 , P1_R1282_U15 , P1_U4036 );
nand NAND2_2060 ( P1_U4658 , P1_U4021 , P1_U4185 );
nand NAND2_2061 ( P1_U4659 , P1_U3703 , P1_U4654 );
nand NAND2_2062 ( P1_U4660 , P1_REG2_REG_26_ , P1_U3018 );
nand NAND2_2063 ( P1_U4661 , P1_REG1_REG_26_ , P1_U3019 );
nand NAND2_2064 ( P1_U4662 , P1_REG0_REG_26_ , P1_U3020 );
nand NAND2_2065 ( P1_U4663 , P1_ADD_99_U62 , P1_U3017 );
not NOT1_2066 ( P1_U4664 , P1_U3057 );
nand NAND2_2067 ( P1_U4665 , P1_U3034 , P1_U3065 );
nand NAND2_2068 ( P1_U4666 , P1_R1150_U95 , P1_U4007 );
nand NAND2_2069 ( P1_U4667 , P1_R1117_U95 , P1_U4000 );
nand NAND2_2070 ( P1_U4668 , P1_R1138_U105 , P1_U3994 );
nand NAND2_2071 ( P1_U4669 , P1_R1192_U95 , P1_U4005 );
nand NAND2_2072 ( P1_U4670 , P1_R1207_U95 , P1_U4004 );
nand NAND2_2073 ( P1_U4671 , P1_R1171_U105 , P1_U4011 );
nand NAND2_2074 ( P1_U4672 , P1_R1240_U105 , P1_U3992 );
not NOT1_2075 ( P1_U4673 , P1_U3408 );
nand NAND2_2076 ( P1_U4674 , P1_U3025 , P1_U3057 );
nand NAND2_2077 ( P1_U4675 , P1_R1222_U105 , P1_U3024 );
nand NAND2_2078 ( P1_U4676 , P1_R1282_U74 , P1_U4036 );
nand NAND2_2079 ( P1_U4677 , P1_U4020 , P1_U4185 );
nand NAND2_2080 ( P1_U4678 , P1_U3707 , P1_U4673 );
nand NAND2_2081 ( P1_U4679 , P1_REG2_REG_27_ , P1_U3018 );
nand NAND2_2082 ( P1_U4680 , P1_REG1_REG_27_ , P1_U3019 );
nand NAND2_2083 ( P1_U4681 , P1_REG0_REG_27_ , P1_U3020 );
nand NAND2_2084 ( P1_U4682 , P1_ADD_99_U61 , P1_U3017 );
not NOT1_2085 ( P1_U4683 , P1_U3053 );
nand NAND2_2086 ( P1_U4684 , P1_U3034 , P1_U3058 );
nand NAND2_2087 ( P1_U4685 , P1_R1150_U109 , P1_U4007 );
nand NAND2_2088 ( P1_U4686 , P1_R1117_U109 , P1_U4000 );
nand NAND2_2089 ( P1_U4687 , P1_R1138_U16 , P1_U3994 );
nand NAND2_2090 ( P1_U4688 , P1_R1192_U109 , P1_U4005 );
nand NAND2_2091 ( P1_U4689 , P1_R1207_U109 , P1_U4004 );
nand NAND2_2092 ( P1_U4690 , P1_R1171_U16 , P1_U4011 );
nand NAND2_2093 ( P1_U4691 , P1_R1240_U16 , P1_U3992 );
not NOT1_2094 ( P1_U4692 , P1_U3410 );
nand NAND2_2095 ( P1_U4693 , P1_U3025 , P1_U3053 );
nand NAND2_2096 ( P1_U4694 , P1_R1222_U16 , P1_U3024 );
nand NAND2_2097 ( P1_U4695 , P1_R1282_U16 , P1_U4036 );
nand NAND2_2098 ( P1_U4696 , P1_U4019 , P1_U4185 );
nand NAND2_2099 ( P1_U4697 , P1_U3711 , P1_U4692 );
nand NAND2_2100 ( P1_U4698 , P1_REG2_REG_28_ , P1_U3018 );
nand NAND2_2101 ( P1_U4699 , P1_REG1_REG_28_ , P1_U3019 );
nand NAND2_2102 ( P1_U4700 , P1_REG0_REG_28_ , P1_U3020 );
nand NAND2_2103 ( P1_U4701 , P1_ADD_99_U60 , P1_U3017 );
not NOT1_2104 ( P1_U4702 , P1_U3054 );
nand NAND2_2105 ( P1_U4703 , P1_U3034 , P1_U3057 );
nand NAND2_2106 ( P1_U4704 , P1_R1150_U16 , P1_U4007 );
nand NAND2_2107 ( P1_U4705 , P1_R1117_U16 , P1_U4000 );
nand NAND2_2108 ( P1_U4706 , P1_R1138_U104 , P1_U3994 );
nand NAND2_2109 ( P1_U4707 , P1_R1192_U16 , P1_U4005 );
nand NAND2_2110 ( P1_U4708 , P1_R1207_U16 , P1_U4004 );
nand NAND2_2111 ( P1_U4709 , P1_R1171_U104 , P1_U4011 );
nand NAND2_2112 ( P1_U4710 , P1_R1240_U104 , P1_U3992 );
not NOT1_2113 ( P1_U4711 , P1_U3412 );
nand NAND2_2114 ( P1_U4712 , P1_U3025 , P1_U3054 );
nand NAND2_2115 ( P1_U4713 , P1_R1222_U104 , P1_U3024 );
nand NAND2_2116 ( P1_U4714 , P1_R1282_U72 , P1_U4036 );
nand NAND2_2117 ( P1_U4715 , P1_U4018 , P1_U4185 );
nand NAND2_2118 ( P1_U4716 , P1_U3715 , P1_U4711 );
nand NAND2_2119 ( P1_U4717 , P1_ADD_99_U5 , P1_U3017 );
nand NAND2_2120 ( P1_U4718 , P1_REG2_REG_29_ , P1_U3018 );
nand NAND2_2121 ( P1_U4719 , P1_REG1_REG_29_ , P1_U3019 );
nand NAND2_2122 ( P1_U4720 , P1_REG0_REG_29_ , P1_U3020 );
not NOT1_2123 ( P1_U4721 , P1_U3055 );
nand NAND2_2124 ( P1_U4722 , P1_U3034 , P1_U3053 );
nand NAND2_2125 ( P1_U4723 , P1_R1150_U94 , P1_U4007 );
nand NAND2_2126 ( P1_U4724 , P1_R1117_U94 , P1_U4000 );
nand NAND2_2127 ( P1_U4725 , P1_R1138_U103 , P1_U3994 );
nand NAND2_2128 ( P1_U4726 , P1_R1192_U94 , P1_U4005 );
nand NAND2_2129 ( P1_U4727 , P1_R1207_U94 , P1_U4004 );
nand NAND2_2130 ( P1_U4728 , P1_R1171_U103 , P1_U4011 );
nand NAND2_2131 ( P1_U4729 , P1_R1240_U103 , P1_U3992 );
not NOT1_2132 ( P1_U4730 , P1_U3414 );
nand NAND2_2133 ( P1_U4731 , P1_U3025 , P1_U3055 );
nand NAND2_2134 ( P1_U4732 , P1_R1222_U103 , P1_U3024 );
nand NAND2_2135 ( P1_U4733 , P1_R1282_U17 , P1_U4036 );
nand NAND2_2136 ( P1_U4734 , P1_U4017 , P1_U4185 );
nand NAND2_2137 ( P1_U4735 , P1_U3719 , P1_U4730 );
nand NAND2_2138 ( P1_U4736 , P1_REG2_REG_30_ , P1_U3018 );
nand NAND2_2139 ( P1_U4737 , P1_REG1_REG_30_ , P1_U3019 );
nand NAND2_2140 ( P1_U4738 , P1_REG0_REG_30_ , P1_U3020 );
not NOT1_2141 ( P1_U4739 , P1_U3059 );
nand NAND2_2142 ( P1_U4740 , P1_U5811 , P1_U3359 );
nand NAND2_2143 ( P1_U4741 , P1_U3954 , P1_U4740 );
nand NAND2_2144 ( P1_U4742 , P1_U3720 , P1_U3059 );
nand NAND2_2145 ( P1_U4743 , P1_U3034 , P1_U3054 );
nand NAND2_2146 ( P1_U4744 , P1_R1150_U17 , P1_U4007 );
nand NAND2_2147 ( P1_U4745 , P1_R1117_U17 , P1_U4000 );
nand NAND2_2148 ( P1_U4746 , P1_R1138_U102 , P1_U3994 );
nand NAND2_2149 ( P1_U4747 , P1_R1192_U17 , P1_U4005 );
nand NAND2_2150 ( P1_U4748 , P1_R1207_U17 , P1_U4004 );
nand NAND2_2151 ( P1_U4749 , P1_R1171_U102 , P1_U4011 );
nand NAND2_2152 ( P1_U4750 , P1_R1240_U102 , P1_U3992 );
not NOT1_2153 ( P1_U4751 , P1_U3416 );
nand NAND2_2154 ( P1_U4752 , P1_R1222_U102 , P1_U3024 );
nand NAND2_2155 ( P1_U4753 , P1_R1282_U70 , P1_U4036 );
nand NAND2_2156 ( P1_U4754 , P1_U4028 , P1_U4185 );
nand NAND2_2157 ( P1_U4755 , P1_U3724 , P1_U4751 );
nand NAND2_2158 ( P1_U4756 , P1_REG2_REG_31_ , P1_U3018 );
nand NAND2_2159 ( P1_U4757 , P1_REG1_REG_31_ , P1_U3019 );
nand NAND2_2160 ( P1_U4758 , P1_REG0_REG_31_ , P1_U3020 );
not NOT1_2161 ( P1_U4759 , P1_U3056 );
nand NAND2_2162 ( P1_U4760 , P1_R1282_U19 , P1_U4036 );
nand NAND2_2163 ( P1_U4761 , P1_U4027 , P1_U4185 );
nand NAND3_2164 ( P1_U4762 , P1_U4761 , P1_U3987 , P1_U4760 );
nand NAND2_2165 ( P1_U4763 , P1_R1282_U68 , P1_U4036 );
nand NAND2_2166 ( P1_U4764 , P1_U4026 , P1_U4185 );
nand NAND3_2167 ( P1_U4765 , P1_U4764 , P1_U3987 , P1_U4763 );
nand NAND2_2168 ( P1_U4766 , P1_U3727 , P1_U3016 );
nand NAND2_2169 ( P1_U4767 , P1_U3421 , P1_U4766 );
nand NAND2_2170 ( P1_U4768 , P1_U3995 , P1_U5802 );
not NOT1_2171 ( P1_U4769 , P1_U3426 );
nand NAND2_2172 ( P1_U4770 , P1_U3036 , P1_U3078 );
nand NAND2_2173 ( P1_U4771 , P1_U3033 , P1_REG3_REG_0_ );
nand NAND2_2174 ( P1_U4772 , P1_U3032 , P1_R1222_U96 );
nand NAND2_2175 ( P1_U4773 , P1_U3031 , P1_U3456 );
nand NAND2_2176 ( P1_U4774 , P1_U3030 , P1_U3456 );
nand NAND2_2177 ( P1_U4775 , P1_U3036 , P1_U3068 );
nand NAND2_2178 ( P1_U4776 , P1_U3033 , P1_REG3_REG_1_ );
nand NAND2_2179 ( P1_U4777 , P1_U3032 , P1_R1222_U95 );
nand NAND2_2180 ( P1_U4778 , P1_U3031 , P1_U3461 );
nand NAND2_2181 ( P1_U4779 , P1_U3030 , P1_R1282_U56 );
nand NAND2_2182 ( P1_U4780 , P1_U3036 , P1_U3064 );
nand NAND2_2183 ( P1_U4781 , P1_U3033 , P1_REG3_REG_2_ );
nand NAND2_2184 ( P1_U4782 , P1_U3032 , P1_R1222_U17 );
nand NAND2_2185 ( P1_U4783 , P1_U3031 , P1_U3464 );
nand NAND2_2186 ( P1_U4784 , P1_U3030 , P1_R1282_U18 );
nand NAND2_2187 ( P1_U4785 , P1_U3036 , P1_U3060 );
nand NAND2_2188 ( P1_U4786 , P1_U3033 , P1_ADD_99_U4 );
nand NAND2_2189 ( P1_U4787 , P1_U3032 , P1_R1222_U101 );
nand NAND2_2190 ( P1_U4788 , P1_U3031 , P1_U3467 );
nand NAND2_2191 ( P1_U4789 , P1_U3030 , P1_R1282_U20 );
nand NAND2_2192 ( P1_U4790 , P1_U3036 , P1_U3067 );
nand NAND2_2193 ( P1_U4791 , P1_U3033 , P1_ADD_99_U59 );
nand NAND2_2194 ( P1_U4792 , P1_U3032 , P1_R1222_U100 );
nand NAND2_2195 ( P1_U4793 , P1_U3031 , P1_U3470 );
nand NAND2_2196 ( P1_U4794 , P1_U3030 , P1_R1282_U21 );
nand NAND2_2197 ( P1_U4795 , P1_U3036 , P1_U3071 );
nand NAND2_2198 ( P1_U4796 , P1_U3033 , P1_ADD_99_U58 );
nand NAND2_2199 ( P1_U4797 , P1_U3032 , P1_R1222_U18 );
nand NAND2_2200 ( P1_U4798 , P1_U3031 , P1_U3473 );
nand NAND2_2201 ( P1_U4799 , P1_U3030 , P1_R1282_U65 );
nand NAND2_2202 ( P1_U4800 , P1_U3036 , P1_U3070 );
nand NAND2_2203 ( P1_U4801 , P1_U3033 , P1_ADD_99_U57 );
nand NAND2_2204 ( P1_U4802 , P1_U3032 , P1_R1222_U99 );
nand NAND2_2205 ( P1_U4803 , P1_U3031 , P1_U3476 );
nand NAND2_2206 ( P1_U4804 , P1_U3030 , P1_R1282_U22 );
nand NAND2_2207 ( P1_U4805 , P1_U3036 , P1_U3084 );
nand NAND2_2208 ( P1_U4806 , P1_U3033 , P1_ADD_99_U56 );
nand NAND2_2209 ( P1_U4807 , P1_U3032 , P1_R1222_U19 );
nand NAND2_2210 ( P1_U4808 , P1_U3031 , P1_U3479 );
nand NAND2_2211 ( P1_U4809 , P1_U3030 , P1_R1282_U23 );
nand NAND2_2212 ( P1_U4810 , P1_U3036 , P1_U3083 );
nand NAND2_2213 ( P1_U4811 , P1_U3033 , P1_ADD_99_U55 );
nand NAND2_2214 ( P1_U4812 , P1_U3032 , P1_R1222_U98 );
nand NAND2_2215 ( P1_U4813 , P1_U3031 , P1_U3482 );
nand NAND2_2216 ( P1_U4814 , P1_U3030 , P1_R1282_U24 );
nand NAND2_2217 ( P1_U4815 , P1_U3036 , P1_U3062 );
nand NAND2_2218 ( P1_U4816 , P1_U3033 , P1_ADD_99_U54 );
nand NAND2_2219 ( P1_U4817 , P1_U3032 , P1_R1222_U97 );
nand NAND2_2220 ( P1_U4818 , P1_U3031 , P1_U3485 );
nand NAND2_2221 ( P1_U4819 , P1_U3030 , P1_R1282_U63 );
nand NAND2_2222 ( P1_U4820 , P1_U3036 , P1_U3063 );
nand NAND2_2223 ( P1_U4821 , P1_U3033 , P1_ADD_99_U78 );
nand NAND2_2224 ( P1_U4822 , P1_U3032 , P1_R1222_U11 );
nand NAND2_2225 ( P1_U4823 , P1_U3031 , P1_U3488 );
nand NAND2_2226 ( P1_U4824 , P1_U3030 , P1_R1282_U6 );
nand NAND2_2227 ( P1_U4825 , P1_U3036 , P1_U3072 );
nand NAND2_2228 ( P1_U4826 , P1_U3033 , P1_ADD_99_U77 );
nand NAND2_2229 ( P1_U4827 , P1_U3032 , P1_R1222_U115 );
nand NAND2_2230 ( P1_U4828 , P1_U3031 , P1_U3491 );
nand NAND2_2231 ( P1_U4829 , P1_U3030 , P1_R1282_U7 );
nand NAND2_2232 ( P1_U4830 , P1_U3036 , P1_U3080 );
nand NAND2_2233 ( P1_U4831 , P1_U3033 , P1_ADD_99_U76 );
nand NAND2_2234 ( P1_U4832 , P1_U3032 , P1_R1222_U114 );
nand NAND2_2235 ( P1_U4833 , P1_U3031 , P1_U3494 );
nand NAND2_2236 ( P1_U4834 , P1_U3030 , P1_R1282_U8 );
nand NAND2_2237 ( P1_U4835 , P1_U3036 , P1_U3079 );
nand NAND2_2238 ( P1_U4836 , P1_U3033 , P1_ADD_99_U75 );
nand NAND2_2239 ( P1_U4837 , P1_U3032 , P1_R1222_U12 );
nand NAND2_2240 ( P1_U4838 , P1_U3031 , P1_U3497 );
nand NAND2_2241 ( P1_U4839 , P1_U3030 , P1_R1282_U86 );
nand NAND2_2242 ( P1_U4840 , P1_U3036 , P1_U3074 );
nand NAND2_2243 ( P1_U4841 , P1_U3033 , P1_ADD_99_U74 );
nand NAND2_2244 ( P1_U4842 , P1_U3032 , P1_R1222_U113 );
nand NAND2_2245 ( P1_U4843 , P1_U3031 , P1_U3500 );
nand NAND2_2246 ( P1_U4844 , P1_U3030 , P1_R1282_U9 );
nand NAND2_2247 ( P1_U4845 , P1_U3036 , P1_U3073 );
nand NAND2_2248 ( P1_U4846 , P1_U3033 , P1_ADD_99_U73 );
nand NAND2_2249 ( P1_U4847 , P1_U3032 , P1_R1222_U112 );
nand NAND2_2250 ( P1_U4848 , P1_U3031 , P1_U3503 );
nand NAND2_2251 ( P1_U4849 , P1_U3030 , P1_R1282_U10 );
nand NAND2_2252 ( P1_U4850 , P1_U3036 , P1_U3069 );
nand NAND2_2253 ( P1_U4851 , P1_U3033 , P1_ADD_99_U72 );
nand NAND2_2254 ( P1_U4852 , P1_U3032 , P1_R1222_U111 );
nand NAND2_2255 ( P1_U4853 , P1_U3031 , P1_U3506 );
nand NAND2_2256 ( P1_U4854 , P1_U3030 , P1_R1282_U11 );
nand NAND2_2257 ( P1_U4855 , P1_U3036 , P1_U3082 );
nand NAND2_2258 ( P1_U4856 , P1_U3033 , P1_ADD_99_U71 );
nand NAND2_2259 ( P1_U4857 , P1_U3032 , P1_R1222_U13 );
nand NAND2_2260 ( P1_U4858 , P1_U3031 , P1_U3509 );
nand NAND2_2261 ( P1_U4859 , P1_U3030 , P1_R1282_U84 );
nand NAND2_2262 ( P1_U4860 , P1_U3036 , P1_U3081 );
nand NAND2_2263 ( P1_U4861 , P1_U3033 , P1_ADD_99_U70 );
nand NAND2_2264 ( P1_U4862 , P1_U3032 , P1_R1222_U110 );
nand NAND2_2265 ( P1_U4863 , P1_U3031 , P1_U3512 );
nand NAND2_2266 ( P1_U4864 , P1_U3030 , P1_R1282_U12 );
nand NAND2_2267 ( P1_U4865 , P1_U3036 , P1_U3076 );
nand NAND2_2268 ( P1_U4866 , P1_U3033 , P1_ADD_99_U69 );
nand NAND2_2269 ( P1_U4867 , P1_U3032 , P1_R1222_U109 );
nand NAND2_2270 ( P1_U4868 , P1_U3031 , P1_U3514 );
nand NAND2_2271 ( P1_U4869 , P1_U3030 , P1_R1282_U82 );
nand NAND2_2272 ( P1_U4870 , P1_U3036 , P1_U3075 );
nand NAND2_2273 ( P1_U4871 , P1_U3033 , P1_ADD_99_U68 );
nand NAND2_2274 ( P1_U4872 , P1_U3032 , P1_R1222_U14 );
nand NAND2_2275 ( P1_U4873 , P1_U3031 , P1_U4025 );
nand NAND2_2276 ( P1_U4874 , P1_U3030 , P1_R1282_U13 );
nand NAND2_2277 ( P1_U4875 , P1_U3036 , P1_U3061 );
nand NAND2_2278 ( P1_U4876 , P1_U3033 , P1_ADD_99_U67 );
nand NAND2_2279 ( P1_U4877 , P1_U3032 , P1_R1222_U15 );
nand NAND2_2280 ( P1_U4878 , P1_U3031 , P1_U4024 );
nand NAND2_2281 ( P1_U4879 , P1_U3030 , P1_R1282_U78 );
nand NAND2_2282 ( P1_U4880 , P1_U3036 , P1_U3066 );
nand NAND2_2283 ( P1_U4881 , P1_U3033 , P1_ADD_99_U66 );
nand NAND2_2284 ( P1_U4882 , P1_U3032 , P1_R1222_U108 );
nand NAND2_2285 ( P1_U4883 , P1_U3031 , P1_U4023 );
nand NAND2_2286 ( P1_U4884 , P1_U3030 , P1_R1282_U14 );
nand NAND2_2287 ( P1_U4885 , P1_U3036 , P1_U3065 );
nand NAND2_2288 ( P1_U4886 , P1_U3033 , P1_ADD_99_U65 );
nand NAND2_2289 ( P1_U4887 , P1_U3032 , P1_R1222_U107 );
nand NAND2_2290 ( P1_U4888 , P1_U3031 , P1_U4022 );
nand NAND2_2291 ( P1_U4889 , P1_U3030 , P1_R1282_U76 );
nand NAND2_2292 ( P1_U4890 , P1_U3036 , P1_U3058 );
nand NAND2_2293 ( P1_U4891 , P1_U3033 , P1_ADD_99_U64 );
nand NAND2_2294 ( P1_U4892 , P1_U3032 , P1_R1222_U106 );
nand NAND2_2295 ( P1_U4893 , P1_U3031 , P1_U4021 );
nand NAND2_2296 ( P1_U4894 , P1_U3030 , P1_R1282_U15 );
nand NAND2_2297 ( P1_U4895 , P1_U3036 , P1_U3057 );
nand NAND2_2298 ( P1_U4896 , P1_U3033 , P1_ADD_99_U63 );
nand NAND2_2299 ( P1_U4897 , P1_U3032 , P1_R1222_U105 );
nand NAND2_2300 ( P1_U4898 , P1_U3031 , P1_U4020 );
nand NAND2_2301 ( P1_U4899 , P1_U3030 , P1_R1282_U74 );
nand NAND2_2302 ( P1_U4900 , P1_U3036 , P1_U3053 );
nand NAND2_2303 ( P1_U4901 , P1_U3033 , P1_ADD_99_U62 );
nand NAND2_2304 ( P1_U4902 , P1_U3032 , P1_R1222_U16 );
nand NAND2_2305 ( P1_U4903 , P1_U3031 , P1_U4019 );
nand NAND2_2306 ( P1_U4904 , P1_U3030 , P1_R1282_U16 );
nand NAND2_2307 ( P1_U4905 , P1_U3036 , P1_U3054 );
nand NAND2_2308 ( P1_U4906 , P1_U3033 , P1_ADD_99_U61 );
nand NAND2_2309 ( P1_U4907 , P1_U3032 , P1_R1222_U104 );
nand NAND2_2310 ( P1_U4908 , P1_U3031 , P1_U4018 );
nand NAND2_2311 ( P1_U4909 , P1_U3030 , P1_R1282_U72 );
nand NAND2_2312 ( P1_U4910 , P1_U3036 , P1_U3055 );
nand NAND2_2313 ( P1_U4911 , P1_U3033 , P1_ADD_99_U60 );
nand NAND2_2314 ( P1_U4912 , P1_U3032 , P1_R1222_U103 );
nand NAND2_2315 ( P1_U4913 , P1_U3031 , P1_U4017 );
nand NAND2_2316 ( P1_U4914 , P1_U3030 , P1_R1282_U17 );
nand NAND2_2317 ( P1_U4915 , P1_U3033 , P1_ADD_99_U5 );
nand NAND2_2318 ( P1_U4916 , P1_U3032 , P1_R1222_U102 );
nand NAND2_2319 ( P1_U4917 , P1_U3031 , P1_U4028 );
nand NAND2_2320 ( P1_U4918 , P1_U3030 , P1_R1282_U70 );
nand NAND2_2321 ( P1_U4919 , P1_U3031 , P1_U4027 );
nand NAND2_2322 ( P1_U4920 , P1_U3030 , P1_R1282_U19 );
nand NAND2_2323 ( P1_U4921 , P1_U3031 , P1_U4026 );
nand NAND2_2324 ( P1_U4922 , P1_U3030 , P1_R1282_U68 );
nand NAND5_2325 ( P1_U4923 , P1_U3787 , P1_U3786 , P1_U3789 , P1_U4769 , P1_U3421 );
nand NAND2_2326 ( P1_U4924 , P1_R1105_U13 , P1_U3042 );
nand NAND2_2327 ( P1_U4925 , P1_U3040 , P1_U3452 );
nand NAND2_2328 ( P1_U4926 , P1_R1162_U13 , P1_U3038 );
nand NAND3_2329 ( P1_U4927 , P1_U4925 , P1_U4924 , P1_U4926 );
nand NAND2_2330 ( P1_U4928 , P1_U3425 , P1_U3372 );
nand NAND2_2331 ( P1_U4929 , P1_U5786 , P1_U4928 );
nand NAND2_2332 ( P1_U4930 , P1_U4929 , P1_U3954 );
not NOT1_2333 ( P1_U4931 , P1_U3085 );
not NOT1_2334 ( P1_U4932 , P1_U3428 );
nand NAND2_2335 ( P1_U4933 , P1_U3044 , P1_U4927 );
nand NAND2_2336 ( P1_U4934 , P1_U3043 , P1_R1105_U13 );
nand NAND2_2337 ( P1_U4935 , P1_REG3_REG_19_ , P1_U3086 );
nand NAND2_2338 ( P1_U4936 , P1_U3041 , P1_U3452 );
nand NAND2_2339 ( P1_U4937 , P1_U3039 , P1_R1162_U13 );
nand NAND2_2340 ( P1_U4938 , P1_ADDR_REG_19_ , P1_U4932 );
nand NAND2_2341 ( P1_U4939 , P1_R1105_U75 , P1_U3042 );
nand NAND2_2342 ( P1_U4940 , P1_U3040 , P1_U3511 );
nand NAND2_2343 ( P1_U4941 , P1_R1162_U75 , P1_U3038 );
nand NAND3_2344 ( P1_U4942 , P1_U4940 , P1_U4939 , P1_U4941 );
nand NAND2_2345 ( P1_U4943 , P1_U3044 , P1_U4942 );
nand NAND2_2346 ( P1_U4944 , P1_R1105_U75 , P1_U3043 );
nand NAND2_2347 ( P1_U4945 , P1_REG3_REG_18_ , P1_U3086 );
nand NAND2_2348 ( P1_U4946 , P1_U3041 , P1_U3511 );
nand NAND2_2349 ( P1_U4947 , P1_R1162_U75 , P1_U3039 );
nand NAND2_2350 ( P1_U4948 , P1_ADDR_REG_18_ , P1_U4932 );
nand NAND2_2351 ( P1_U4949 , P1_R1105_U12 , P1_U3042 );
nand NAND2_2352 ( P1_U4950 , P1_U3040 , P1_U3508 );
nand NAND2_2353 ( P1_U4951 , P1_R1162_U12 , P1_U3038 );
nand NAND3_2354 ( P1_U4952 , P1_U4950 , P1_U4949 , P1_U4951 );
nand NAND2_2355 ( P1_U4953 , P1_U3044 , P1_U4952 );
nand NAND2_2356 ( P1_U4954 , P1_R1105_U12 , P1_U3043 );
nand NAND2_2357 ( P1_U4955 , P1_REG3_REG_17_ , P1_U3086 );
nand NAND2_2358 ( P1_U4956 , P1_U3041 , P1_U3508 );
nand NAND2_2359 ( P1_U4957 , P1_R1162_U12 , P1_U3039 );
nand NAND2_2360 ( P1_U4958 , P1_ADDR_REG_17_ , P1_U4932 );
nand NAND2_2361 ( P1_U4959 , P1_R1105_U76 , P1_U3042 );
nand NAND2_2362 ( P1_U4960 , P1_U3040 , P1_U3505 );
nand NAND2_2363 ( P1_U4961 , P1_R1162_U76 , P1_U3038 );
nand NAND3_2364 ( P1_U4962 , P1_U4960 , P1_U4959 , P1_U4961 );
nand NAND2_2365 ( P1_U4963 , P1_U3044 , P1_U4962 );
nand NAND2_2366 ( P1_U4964 , P1_R1105_U76 , P1_U3043 );
nand NAND2_2367 ( P1_U4965 , P1_REG3_REG_16_ , P1_U3086 );
nand NAND2_2368 ( P1_U4966 , P1_U3041 , P1_U3505 );
nand NAND2_2369 ( P1_U4967 , P1_R1162_U76 , P1_U3039 );
nand NAND2_2370 ( P1_U4968 , P1_ADDR_REG_16_ , P1_U4932 );
nand NAND2_2371 ( P1_U4969 , P1_R1105_U77 , P1_U3042 );
nand NAND2_2372 ( P1_U4970 , P1_U3040 , P1_U3502 );
nand NAND2_2373 ( P1_U4971 , P1_R1162_U77 , P1_U3038 );
nand NAND3_2374 ( P1_U4972 , P1_U4970 , P1_U4969 , P1_U4971 );
nand NAND2_2375 ( P1_U4973 , P1_U3044 , P1_U4972 );
nand NAND2_2376 ( P1_U4974 , P1_R1105_U77 , P1_U3043 );
nand NAND2_2377 ( P1_U4975 , P1_REG3_REG_15_ , P1_U3086 );
nand NAND2_2378 ( P1_U4976 , P1_U3041 , P1_U3502 );
nand NAND2_2379 ( P1_U4977 , P1_R1162_U77 , P1_U3039 );
nand NAND2_2380 ( P1_U4978 , P1_ADDR_REG_15_ , P1_U4932 );
nand NAND2_2381 ( P1_U4979 , P1_R1105_U78 , P1_U3042 );
nand NAND2_2382 ( P1_U4980 , P1_U3040 , P1_U3499 );
nand NAND2_2383 ( P1_U4981 , P1_R1162_U78 , P1_U3038 );
nand NAND3_2384 ( P1_U4982 , P1_U4980 , P1_U4979 , P1_U4981 );
nand NAND2_2385 ( P1_U4983 , P1_U3044 , P1_U4982 );
nand NAND2_2386 ( P1_U4984 , P1_R1105_U78 , P1_U3043 );
nand NAND2_2387 ( P1_U4985 , P1_REG3_REG_14_ , P1_U3086 );
nand NAND2_2388 ( P1_U4986 , P1_U3041 , P1_U3499 );
nand NAND2_2389 ( P1_U4987 , P1_R1162_U78 , P1_U3039 );
nand NAND2_2390 ( P1_U4988 , P1_ADDR_REG_14_ , P1_U4932 );
nand NAND2_2391 ( P1_U4989 , P1_R1105_U11 , P1_U3042 );
nand NAND2_2392 ( P1_U4990 , P1_U3040 , P1_U3496 );
nand NAND2_2393 ( P1_U4991 , P1_R1162_U11 , P1_U3038 );
nand NAND3_2394 ( P1_U4992 , P1_U4990 , P1_U4989 , P1_U4991 );
nand NAND2_2395 ( P1_U4993 , P1_U3044 , P1_U4992 );
nand NAND2_2396 ( P1_U4994 , P1_R1105_U11 , P1_U3043 );
nand NAND2_2397 ( P1_U4995 , P1_REG3_REG_13_ , P1_U3086 );
nand NAND2_2398 ( P1_U4996 , P1_U3041 , P1_U3496 );
nand NAND2_2399 ( P1_U4997 , P1_R1162_U11 , P1_U3039 );
nand NAND2_2400 ( P1_U4998 , P1_ADDR_REG_13_ , P1_U4932 );
nand NAND2_2401 ( P1_U4999 , P1_R1105_U79 , P1_U3042 );
nand NAND2_2402 ( P1_U5000 , P1_U3040 , P1_U3493 );
nand NAND2_2403 ( P1_U5001 , P1_R1162_U79 , P1_U3038 );
nand NAND3_2404 ( P1_U5002 , P1_U5000 , P1_U4999 , P1_U5001 );
nand NAND2_2405 ( P1_U5003 , P1_U3044 , P1_U5002 );
nand NAND2_2406 ( P1_U5004 , P1_R1105_U79 , P1_U3043 );
nand NAND2_2407 ( P1_U5005 , P1_REG3_REG_12_ , P1_U3086 );
nand NAND2_2408 ( P1_U5006 , P1_U3041 , P1_U3493 );
nand NAND2_2409 ( P1_U5007 , P1_R1162_U79 , P1_U3039 );
nand NAND2_2410 ( P1_U5008 , P1_ADDR_REG_12_ , P1_U4932 );
nand NAND2_2411 ( P1_U5009 , P1_R1105_U80 , P1_U3042 );
nand NAND2_2412 ( P1_U5010 , P1_U3040 , P1_U3490 );
nand NAND2_2413 ( P1_U5011 , P1_R1162_U80 , P1_U3038 );
nand NAND3_2414 ( P1_U5012 , P1_U5010 , P1_U5009 , P1_U5011 );
nand NAND2_2415 ( P1_U5013 , P1_U3044 , P1_U5012 );
nand NAND2_2416 ( P1_U5014 , P1_R1105_U80 , P1_U3043 );
nand NAND2_2417 ( P1_U5015 , P1_REG3_REG_11_ , P1_U3086 );
nand NAND2_2418 ( P1_U5016 , P1_U3041 , P1_U3490 );
nand NAND2_2419 ( P1_U5017 , P1_R1162_U80 , P1_U3039 );
nand NAND2_2420 ( P1_U5018 , P1_ADDR_REG_11_ , P1_U4932 );
nand NAND2_2421 ( P1_U5019 , P1_R1105_U10 , P1_U3042 );
nand NAND2_2422 ( P1_U5020 , P1_U3040 , P1_U3487 );
nand NAND2_2423 ( P1_U5021 , P1_R1162_U10 , P1_U3038 );
nand NAND3_2424 ( P1_U5022 , P1_U5020 , P1_U5019 , P1_U5021 );
nand NAND2_2425 ( P1_U5023 , P1_U3044 , P1_U5022 );
nand NAND2_2426 ( P1_U5024 , P1_R1105_U10 , P1_U3043 );
nand NAND2_2427 ( P1_U5025 , P1_REG3_REG_10_ , P1_U3086 );
nand NAND2_2428 ( P1_U5026 , P1_U3041 , P1_U3487 );
nand NAND2_2429 ( P1_U5027 , P1_R1162_U10 , P1_U3039 );
nand NAND2_2430 ( P1_U5028 , P1_ADDR_REG_10_ , P1_U4932 );
nand NAND2_2431 ( P1_U5029 , P1_R1105_U70 , P1_U3042 );
nand NAND2_2432 ( P1_U5030 , P1_U3040 , P1_U3484 );
nand NAND2_2433 ( P1_U5031 , P1_R1162_U70 , P1_U3038 );
nand NAND3_2434 ( P1_U5032 , P1_U5030 , P1_U5029 , P1_U5031 );
nand NAND2_2435 ( P1_U5033 , P1_U3044 , P1_U5032 );
nand NAND2_2436 ( P1_U5034 , P1_R1105_U70 , P1_U3043 );
nand NAND2_2437 ( P1_U5035 , P1_REG3_REG_9_ , P1_U3086 );
nand NAND2_2438 ( P1_U5036 , P1_U3041 , P1_U3484 );
nand NAND2_2439 ( P1_U5037 , P1_R1162_U70 , P1_U3039 );
nand NAND2_2440 ( P1_U5038 , P1_ADDR_REG_9_ , P1_U4932 );
nand NAND2_2441 ( P1_U5039 , P1_R1105_U71 , P1_U3042 );
nand NAND2_2442 ( P1_U5040 , P1_U3040 , P1_U3481 );
nand NAND2_2443 ( P1_U5041 , P1_R1162_U71 , P1_U3038 );
nand NAND3_2444 ( P1_U5042 , P1_U5040 , P1_U5039 , P1_U5041 );
nand NAND2_2445 ( P1_U5043 , P1_U3044 , P1_U5042 );
nand NAND2_2446 ( P1_U5044 , P1_R1105_U71 , P1_U3043 );
nand NAND2_2447 ( P1_U5045 , P1_REG3_REG_8_ , P1_U3086 );
nand NAND2_2448 ( P1_U5046 , P1_U3041 , P1_U3481 );
nand NAND2_2449 ( P1_U5047 , P1_R1162_U71 , P1_U3039 );
nand NAND2_2450 ( P1_U5048 , P1_ADDR_REG_8_ , P1_U4932 );
nand NAND2_2451 ( P1_U5049 , P1_R1105_U16 , P1_U3042 );
nand NAND2_2452 ( P1_U5050 , P1_U3040 , P1_U3478 );
nand NAND2_2453 ( P1_U5051 , P1_R1162_U16 , P1_U3038 );
nand NAND3_2454 ( P1_U5052 , P1_U5050 , P1_U5049 , P1_U5051 );
nand NAND2_2455 ( P1_U5053 , P1_U3044 , P1_U5052 );
nand NAND2_2456 ( P1_U5054 , P1_R1105_U16 , P1_U3043 );
nand NAND2_2457 ( P1_U5055 , P1_REG3_REG_7_ , P1_U3086 );
nand NAND2_2458 ( P1_U5056 , P1_U3041 , P1_U3478 );
nand NAND2_2459 ( P1_U5057 , P1_R1162_U16 , P1_U3039 );
nand NAND2_2460 ( P1_U5058 , P1_ADDR_REG_7_ , P1_U4932 );
nand NAND2_2461 ( P1_U5059 , P1_R1105_U72 , P1_U3042 );
nand NAND2_2462 ( P1_U5060 , P1_U3040 , P1_U3475 );
nand NAND2_2463 ( P1_U5061 , P1_R1162_U72 , P1_U3038 );
nand NAND3_2464 ( P1_U5062 , P1_U5060 , P1_U5059 , P1_U5061 );
nand NAND2_2465 ( P1_U5063 , P1_U3044 , P1_U5062 );
nand NAND2_2466 ( P1_U5064 , P1_R1105_U72 , P1_U3043 );
nand NAND2_2467 ( P1_U5065 , P1_REG3_REG_6_ , P1_U3086 );
nand NAND2_2468 ( P1_U5066 , P1_U3041 , P1_U3475 );
nand NAND2_2469 ( P1_U5067 , P1_R1162_U72 , P1_U3039 );
nand NAND2_2470 ( P1_U5068 , P1_ADDR_REG_6_ , P1_U4932 );
nand NAND2_2471 ( P1_U5069 , P1_R1105_U15 , P1_U3042 );
nand NAND2_2472 ( P1_U5070 , P1_U3040 , P1_U3472 );
nand NAND2_2473 ( P1_U5071 , P1_R1162_U15 , P1_U3038 );
nand NAND3_2474 ( P1_U5072 , P1_U5070 , P1_U5069 , P1_U5071 );
nand NAND2_2475 ( P1_U5073 , P1_U3044 , P1_U5072 );
nand NAND2_2476 ( P1_U5074 , P1_R1105_U15 , P1_U3043 );
nand NAND2_2477 ( P1_U5075 , P1_REG3_REG_5_ , P1_U3086 );
nand NAND2_2478 ( P1_U5076 , P1_U3041 , P1_U3472 );
nand NAND2_2479 ( P1_U5077 , P1_R1162_U15 , P1_U3039 );
nand NAND2_2480 ( P1_U5078 , P1_ADDR_REG_5_ , P1_U4932 );
nand NAND2_2481 ( P1_U5079 , P1_R1105_U73 , P1_U3042 );
nand NAND2_2482 ( P1_U5080 , P1_U3040 , P1_U3469 );
nand NAND2_2483 ( P1_U5081 , P1_R1162_U73 , P1_U3038 );
nand NAND3_2484 ( P1_U5082 , P1_U5080 , P1_U5079 , P1_U5081 );
nand NAND2_2485 ( P1_U5083 , P1_U3044 , P1_U5082 );
nand NAND2_2486 ( P1_U5084 , P1_R1105_U73 , P1_U3043 );
nand NAND2_2487 ( P1_U5085 , P1_REG3_REG_4_ , P1_U3086 );
nand NAND2_2488 ( P1_U5086 , P1_U3041 , P1_U3469 );
nand NAND2_2489 ( P1_U5087 , P1_R1162_U73 , P1_U3039 );
nand NAND2_2490 ( P1_U5088 , P1_ADDR_REG_4_ , P1_U4932 );
nand NAND2_2491 ( P1_U5089 , P1_R1105_U74 , P1_U3042 );
nand NAND2_2492 ( P1_U5090 , P1_U3040 , P1_U3466 );
nand NAND2_2493 ( P1_U5091 , P1_R1162_U74 , P1_U3038 );
nand NAND3_2494 ( P1_U5092 , P1_U5090 , P1_U5089 , P1_U5091 );
nand NAND2_2495 ( P1_U5093 , P1_U3044 , P1_U5092 );
nand NAND2_2496 ( P1_U5094 , P1_R1105_U74 , P1_U3043 );
nand NAND2_2497 ( P1_U5095 , P1_REG3_REG_3_ , P1_U3086 );
nand NAND2_2498 ( P1_U5096 , P1_U3041 , P1_U3466 );
nand NAND2_2499 ( P1_U5097 , P1_R1162_U74 , P1_U3039 );
nand NAND2_2500 ( P1_U5098 , P1_ADDR_REG_3_ , P1_U4932 );
nand NAND2_2501 ( P1_U5099 , P1_R1105_U14 , P1_U3042 );
nand NAND2_2502 ( P1_U5100 , P1_U3040 , P1_U3463 );
nand NAND2_2503 ( P1_U5101 , P1_R1162_U14 , P1_U3038 );
nand NAND3_2504 ( P1_U5102 , P1_U5100 , P1_U5099 , P1_U5101 );
nand NAND2_2505 ( P1_U5103 , P1_U3044 , P1_U5102 );
nand NAND2_2506 ( P1_U5104 , P1_R1105_U14 , P1_U3043 );
nand NAND2_2507 ( P1_U5105 , P1_REG3_REG_2_ , P1_U3086 );
nand NAND2_2508 ( P1_U5106 , P1_U3041 , P1_U3463 );
nand NAND2_2509 ( P1_U5107 , P1_R1162_U14 , P1_U3039 );
nand NAND2_2510 ( P1_U5108 , P1_ADDR_REG_2_ , P1_U4932 );
nand NAND2_2511 ( P1_U5109 , P1_R1105_U68 , P1_U3042 );
nand NAND2_2512 ( P1_U5110 , P1_U3040 , P1_U3460 );
nand NAND2_2513 ( P1_U5111 , P1_R1162_U68 , P1_U3038 );
nand NAND3_2514 ( P1_U5112 , P1_U5110 , P1_U5109 , P1_U5111 );
nand NAND2_2515 ( P1_U5113 , P1_U3044 , P1_U5112 );
nand NAND2_2516 ( P1_U5114 , P1_R1105_U68 , P1_U3043 );
nand NAND2_2517 ( P1_U5115 , P1_REG3_REG_1_ , P1_U3086 );
nand NAND2_2518 ( P1_U5116 , P1_U3041 , P1_U3460 );
nand NAND2_2519 ( P1_U5117 , P1_R1162_U68 , P1_U3039 );
nand NAND2_2520 ( P1_U5118 , P1_ADDR_REG_1_ , P1_U4932 );
nand NAND2_2521 ( P1_U5119 , P1_R1105_U69 , P1_U3042 );
nand NAND2_2522 ( P1_U5120 , P1_U3040 , P1_U3454 );
nand NAND2_2523 ( P1_U5121 , P1_R1162_U69 , P1_U3038 );
nand NAND3_2524 ( P1_U5122 , P1_U5120 , P1_U5119 , P1_U5121 );
nand NAND2_2525 ( P1_U5123 , P1_U3044 , P1_U5122 );
nand NAND2_2526 ( P1_U5124 , P1_R1105_U69 , P1_U3043 );
nand NAND2_2527 ( P1_U5125 , P1_REG3_REG_0_ , P1_U3086 );
nand NAND2_2528 ( P1_U5126 , P1_U3041 , P1_U3454 );
nand NAND2_2529 ( P1_U5127 , P1_R1162_U69 , P1_U3039 );
nand NAND2_2530 ( P1_U5128 , P1_ADDR_REG_0_ , P1_U4932 );
not NOT1_2531 ( P1_U5129 , P1_U3991 );
nand NAND3_2532 ( P1_U5130 , P1_U6277 , P1_U6276 , P1_U3990 );
nand NAND2_2533 ( P1_U5131 , P1_U3370 , P1_U3373 );
nand NAND2_2534 ( P1_U5132 , P1_U5802 , P1_U3451 );
nand NAND2_2535 ( P1_U5133 , P1_U3422 , P1_U5132 );
nand NAND3_2536 ( P1_U5134 , P1_U6279 , P1_U6278 , P1_U5772 );
nand NAND3_2537 ( P1_U5135 , P1_U6281 , P1_U6280 , P1_U3845 );
nand NAND3_2538 ( P1_U5136 , P1_U3022 , P1_U4029 , P1_U3432 );
nand NAND2_2539 ( P1_U5137 , P1_U4043 , P1_U5134 );
nand NAND2_2540 ( P1_U5138 , P1_B_REG , P1_U5135 );
nand NAND2_2541 ( P1_U5139 , P1_U3037 , P1_U3079 );
nand NAND2_2542 ( P1_U5140 , P1_U3035 , P1_U3073 );
nand NAND2_2543 ( P1_U5141 , P1_ADD_99_U73 , P1_U3434 );
nand NAND3_2544 ( P1_U5142 , P1_U5141 , P1_U5139 , P1_U5140 );
not NOT1_2545 ( P1_U5143 , P1_U3152 );
nand NAND2_2546 ( P1_U5144 , P1_U3423 , P1_U3999 );
nand NAND4_2547 ( P1_U5145 , P1_U6283 , P1_U6282 , P1_U3849 , P1_U3848 );
nand NAND2_2548 ( P1_U5146 , P1_U5145 , P1_U3434 );
nand NAND2_2549 ( P1_U5147 , P1_U4012 , P1_U5146 );
nand NAND2_2550 ( P1_U5148 , P1_U3022 , P1_U5147 );
nand NAND2_2551 ( P1_U5149 , P1_U3503 , P1_U5770 );
nand NAND2_2552 ( P1_U5150 , P1_ADD_99_U73 , P1_U5769 );
nand NAND2_2553 ( P1_U5151 , P1_R1165_U105 , P1_U3026 );
nand NAND2_2554 ( P1_U5152 , P1_U4037 , P1_U5142 );
nand NAND2_2555 ( P1_U5153 , P1_REG3_REG_15_ , P1_U3086 );
nand NAND2_2556 ( P1_U5154 , P1_U3037 , P1_U3058 );
nand NAND2_2557 ( P1_U5155 , P1_U3035 , P1_U3053 );
nand NAND2_2558 ( P1_U5156 , P1_ADD_99_U62 , P1_U3434 );
nand NAND3_2559 ( P1_U5157 , P1_U5156 , P1_U5154 , P1_U5155 );
nand NAND2_2560 ( P1_U5158 , P1_U4015 , P1_U3426 );
nand NAND2_2561 ( P1_U5159 , P1_U3421 , P1_U5158 );
nand NAND2_2562 ( P1_U5160 , P1_U3045 , P1_U4019 );
nand NAND2_2563 ( P1_U5161 , P1_ADD_99_U62 , P1_U5769 );
nand NAND2_2564 ( P1_U5162 , P1_R1165_U12 , P1_U3026 );
nand NAND2_2565 ( P1_U5163 , P1_U4037 , P1_U5157 );
nand NAND2_2566 ( P1_U5164 , P1_REG3_REG_26_ , P1_U3086 );
nand NAND2_2567 ( P1_U5165 , P1_U3037 , P1_U3067 );
nand NAND2_2568 ( P1_U5166 , P1_U3035 , P1_U3070 );
nand NAND2_2569 ( P1_U5167 , P1_ADD_99_U57 , P1_U3434 );
nand NAND3_2570 ( P1_U5168 , P1_U5166 , P1_U5165 , P1_U5167 );
nand NAND2_2571 ( P1_U5169 , P1_U3476 , P1_U5770 );
nand NAND2_2572 ( P1_U5170 , P1_ADD_99_U57 , P1_U5769 );
nand NAND2_2573 ( P1_U5171 , P1_R1165_U90 , P1_U3026 );
nand NAND2_2574 ( P1_U5172 , P1_U4037 , P1_U5168 );
nand NAND2_2575 ( P1_U5173 , P1_REG3_REG_6_ , P1_U3086 );
nand NAND2_2576 ( P1_U5174 , P1_U3037 , P1_U3069 );
nand NAND2_2577 ( P1_U5175 , P1_U3035 , P1_U3081 );
nand NAND2_2578 ( P1_U5176 , P1_ADD_99_U70 , P1_U3434 );
nand NAND3_2579 ( P1_U5177 , P1_U5176 , P1_U5174 , P1_U5175 );
nand NAND2_2580 ( P1_U5178 , P1_U3512 , P1_U5770 );
nand NAND2_2581 ( P1_U5179 , P1_ADD_99_U70 , P1_U5769 );
nand NAND2_2582 ( P1_U5180 , P1_R1165_U103 , P1_U3026 );
nand NAND2_2583 ( P1_U5181 , P1_U4037 , P1_U5177 );
nand NAND2_2584 ( P1_U5182 , P1_REG3_REG_18_ , P1_U3086 );
nand NAND2_2585 ( P1_U5183 , P1_U3037 , P1_U3078 );
nand NAND2_2586 ( P1_U5184 , P1_U3035 , P1_U3064 );
nand NAND2_2587 ( P1_U5185 , P1_REG3_REG_2_ , P1_U3434 );
nand NAND3_2588 ( P1_U5186 , P1_U5184 , P1_U5183 , P1_U5185 );
nand NAND2_2589 ( P1_U5187 , P1_U3464 , P1_U5770 );
nand NAND2_2590 ( P1_U5188 , P1_REG3_REG_2_ , P1_U5769 );
nand NAND2_2591 ( P1_U5189 , P1_R1165_U93 , P1_U3026 );
nand NAND2_2592 ( P1_U5190 , P1_U4037 , P1_U5186 );
nand NAND2_2593 ( P1_U5191 , P1_REG3_REG_2_ , P1_U3086 );
nand NAND2_2594 ( P1_U5192 , P1_U3037 , P1_U3062 );
nand NAND2_2595 ( P1_U5193 , P1_U3035 , P1_U3072 );
nand NAND2_2596 ( P1_U5194 , P1_ADD_99_U77 , P1_U3434 );
nand NAND3_2597 ( P1_U5195 , P1_U5193 , P1_U5192 , P1_U5194 );
nand NAND2_2598 ( P1_U5196 , P1_U3491 , P1_U5770 );
nand NAND2_2599 ( P1_U5197 , P1_ADD_99_U77 , P1_U5769 );
nand NAND2_2600 ( P1_U5198 , P1_R1165_U108 , P1_U3026 );
nand NAND2_2601 ( P1_U5199 , P1_U4037 , P1_U5195 );
nand NAND2_2602 ( P1_U5200 , P1_REG3_REG_11_ , P1_U3086 );
nand NAND2_2603 ( P1_U5201 , P1_U3037 , P1_U3075 );
nand NAND2_2604 ( P1_U5202 , P1_U3035 , P1_U3066 );
nand NAND2_2605 ( P1_U5203 , P1_ADD_99_U66 , P1_U3434 );
nand NAND3_2606 ( P1_U5204 , P1_U5203 , P1_U5201 , P1_U5202 );
nand NAND2_2607 ( P1_U5205 , P1_U3045 , P1_U4023 );
nand NAND2_2608 ( P1_U5206 , P1_ADD_99_U66 , P1_U5769 );
nand NAND2_2609 ( P1_U5207 , P1_R1165_U99 , P1_U3026 );
nand NAND2_2610 ( P1_U5208 , P1_U4037 , P1_U5204 );
nand NAND2_2611 ( P1_U5209 , P1_REG3_REG_22_ , P1_U3086 );
nand NAND2_2612 ( P1_U5210 , P1_U3037 , P1_U3072 );
nand NAND2_2613 ( P1_U5211 , P1_U3035 , P1_U3079 );
nand NAND2_2614 ( P1_U5212 , P1_ADD_99_U75 , P1_U3434 );
nand NAND3_2615 ( P1_U5213 , P1_U5212 , P1_U5210 , P1_U5211 );
nand NAND2_2616 ( P1_U5214 , P1_U3497 , P1_U5770 );
nand NAND2_2617 ( P1_U5215 , P1_ADD_99_U75 , P1_U5769 );
nand NAND2_2618 ( P1_U5216 , P1_R1165_U9 , P1_U3026 );
nand NAND2_2619 ( P1_U5217 , P1_U4037 , P1_U5213 );
nand NAND2_2620 ( P1_U5218 , P1_REG3_REG_13_ , P1_U3086 );
nand NAND2_2621 ( P1_U5219 , P1_U3037 , P1_U3081 );
nand NAND2_2622 ( P1_U5220 , P1_U3035 , P1_U3075 );
nand NAND2_2623 ( P1_U5221 , P1_ADD_99_U68 , P1_U3434 );
nand NAND3_2624 ( P1_U5222 , P1_U5221 , P1_U5219 , P1_U5220 );
nand NAND2_2625 ( P1_U5223 , P1_U3045 , P1_U4025 );
nand NAND2_2626 ( P1_U5224 , P1_ADD_99_U68 , P1_U5769 );
nand NAND2_2627 ( P1_U5225 , P1_R1165_U100 , P1_U3026 );
nand NAND2_2628 ( P1_U5226 , P1_U4037 , P1_U5222 );
nand NAND2_2629 ( P1_U5227 , P1_REG3_REG_20_ , P1_U3086 );
nand NAND2_2630 ( P1_U5228 , P1_U3435 , P1_U3433 );
nand NAND2_2631 ( P1_U5229 , P1_U5228 , P1_U3434 );
nand NAND2_2632 ( P1_U5230 , P1_U3050 , P1_U5229 );
nand NAND2_2633 ( P1_U5231 , P1_U3858 , P1_U3035 );
nand NAND2_2634 ( P1_U5232 , P1_U3456 , P1_U5770 );
nand NAND2_2635 ( P1_U5233 , P1_REG3_REG_0_ , P1_U5230 );
nand NAND2_2636 ( P1_U5234 , P1_R1165_U87 , P1_U3026 );
nand NAND2_2637 ( P1_U5235 , P1_REG3_REG_0_ , P1_U3086 );
nand NAND2_2638 ( P1_U5236 , P1_U3037 , P1_U3084 );
nand NAND2_2639 ( P1_U5237 , P1_U3035 , P1_U3062 );
nand NAND2_2640 ( P1_U5238 , P1_ADD_99_U54 , P1_U3434 );
nand NAND3_2641 ( P1_U5239 , P1_U5237 , P1_U5236 , P1_U5238 );
nand NAND2_2642 ( P1_U5240 , P1_U3485 , P1_U5770 );
nand NAND2_2643 ( P1_U5241 , P1_ADD_99_U54 , P1_U5769 );
nand NAND2_2644 ( P1_U5242 , P1_R1165_U88 , P1_U3026 );
nand NAND2_2645 ( P1_U5243 , P1_U4037 , P1_U5239 );
nand NAND2_2646 ( P1_U5244 , P1_REG3_REG_9_ , P1_U3086 );
nand NAND2_2647 ( P1_U5245 , P1_U3037 , P1_U3064 );
nand NAND2_2648 ( P1_U5246 , P1_U3035 , P1_U3067 );
nand NAND2_2649 ( P1_U5247 , P1_ADD_99_U59 , P1_U3434 );
nand NAND3_2650 ( P1_U5248 , P1_U5246 , P1_U5245 , P1_U5247 );
nand NAND2_2651 ( P1_U5249 , P1_U3470 , P1_U5770 );
nand NAND2_2652 ( P1_U5250 , P1_ADD_99_U59 , P1_U5769 );
nand NAND2_2653 ( P1_U5251 , P1_R1165_U92 , P1_U3026 );
nand NAND2_2654 ( P1_U5252 , P1_U4037 , P1_U5248 );
nand NAND2_2655 ( P1_U5253 , P1_REG3_REG_4_ , P1_U3086 );
nand NAND2_2656 ( P1_U5254 , P1_U3037 , P1_U3066 );
nand NAND2_2657 ( P1_U5255 , P1_U3035 , P1_U3058 );
nand NAND2_2658 ( P1_U5256 , P1_ADD_99_U64 , P1_U3434 );
nand NAND3_2659 ( P1_U5257 , P1_U5256 , P1_U5254 , P1_U5255 );
nand NAND2_2660 ( P1_U5258 , P1_U3045 , P1_U4021 );
nand NAND2_2661 ( P1_U5259 , P1_ADD_99_U64 , P1_U5769 );
nand NAND2_2662 ( P1_U5260 , P1_R1165_U97 , P1_U3026 );
nand NAND2_2663 ( P1_U5261 , P1_U4037 , P1_U5257 );
nand NAND2_2664 ( P1_U5262 , P1_REG3_REG_24_ , P1_U3086 );
nand NAND2_2665 ( P1_U5263 , P1_U3037 , P1_U3073 );
nand NAND2_2666 ( P1_U5264 , P1_U3035 , P1_U3082 );
nand NAND2_2667 ( P1_U5265 , P1_ADD_99_U71 , P1_U3434 );
nand NAND3_2668 ( P1_U5266 , P1_U5265 , P1_U5263 , P1_U5264 );
nand NAND2_2669 ( P1_U5267 , P1_U3509 , P1_U5770 );
nand NAND2_2670 ( P1_U5268 , P1_ADD_99_U71 , P1_U5769 );
nand NAND2_2671 ( P1_U5269 , P1_R1165_U10 , P1_U3026 );
nand NAND2_2672 ( P1_U5270 , P1_U4037 , P1_U5266 );
nand NAND2_2673 ( P1_U5271 , P1_REG3_REG_17_ , P1_U3086 );
nand NAND2_2674 ( P1_U5272 , P1_U3037 , P1_U3060 );
nand NAND2_2675 ( P1_U5273 , P1_U3035 , P1_U3071 );
nand NAND2_2676 ( P1_U5274 , P1_ADD_99_U58 , P1_U3434 );
nand NAND3_2677 ( P1_U5275 , P1_U5273 , P1_U5272 , P1_U5274 );
nand NAND2_2678 ( P1_U5276 , P1_U3473 , P1_U5770 );
nand NAND2_2679 ( P1_U5277 , P1_ADD_99_U58 , P1_U5769 );
nand NAND2_2680 ( P1_U5278 , P1_R1165_U91 , P1_U3026 );
nand NAND2_2681 ( P1_U5279 , P1_U4037 , P1_U5275 );
nand NAND2_2682 ( P1_U5280 , P1_REG3_REG_5_ , P1_U3086 );
nand NAND2_2683 ( P1_U5281 , P1_U3037 , P1_U3074 );
nand NAND2_2684 ( P1_U5282 , P1_U3035 , P1_U3069 );
nand NAND2_2685 ( P1_U5283 , P1_ADD_99_U72 , P1_U3434 );
nand NAND3_2686 ( P1_U5284 , P1_U5283 , P1_U5281 , P1_U5282 );
nand NAND2_2687 ( P1_U5285 , P1_U3506 , P1_U5770 );
nand NAND2_2688 ( P1_U5286 , P1_ADD_99_U72 , P1_U5769 );
nand NAND2_2689 ( P1_U5287 , P1_R1165_U104 , P1_U3026 );
nand NAND2_2690 ( P1_U5288 , P1_U4037 , P1_U5284 );
nand NAND2_2691 ( P1_U5289 , P1_REG3_REG_16_ , P1_U3086 );
nand NAND2_2692 ( P1_U5290 , P1_U3037 , P1_U3065 );
nand NAND2_2693 ( P1_U5291 , P1_U3035 , P1_U3057 );
nand NAND2_2694 ( P1_U5292 , P1_ADD_99_U63 , P1_U3434 );
nand NAND3_2695 ( P1_U5293 , P1_U5292 , P1_U5290 , P1_U5291 );
nand NAND2_2696 ( P1_U5294 , P1_U3045 , P1_U4020 );
nand NAND2_2697 ( P1_U5295 , P1_ADD_99_U63 , P1_U5769 );
nand NAND2_2698 ( P1_U5296 , P1_R1165_U96 , P1_U3026 );
nand NAND2_2699 ( P1_U5297 , P1_U4037 , P1_U5293 );
nand NAND2_2700 ( P1_U5298 , P1_REG3_REG_25_ , P1_U3086 );
nand NAND2_2701 ( P1_U5299 , P1_U3037 , P1_U3063 );
nand NAND2_2702 ( P1_U5300 , P1_U3035 , P1_U3080 );
nand NAND2_2703 ( P1_U5301 , P1_ADD_99_U76 , P1_U3434 );
nand NAND3_2704 ( P1_U5302 , P1_U5301 , P1_U5299 , P1_U5300 );
nand NAND2_2705 ( P1_U5303 , P1_U3494 , P1_U5770 );
nand NAND2_2706 ( P1_U5304 , P1_ADD_99_U76 , P1_U5769 );
nand NAND2_2707 ( P1_U5305 , P1_R1165_U107 , P1_U3026 );
nand NAND2_2708 ( P1_U5306 , P1_U4037 , P1_U5302 );
nand NAND2_2709 ( P1_U5307 , P1_REG3_REG_12_ , P1_U3086 );
nand NAND2_2710 ( P1_U5308 , P1_U3037 , P1_U3076 );
nand NAND2_2711 ( P1_U5309 , P1_U3035 , P1_U3061 );
nand NAND2_2712 ( P1_U5310 , P1_ADD_99_U67 , P1_U3434 );
nand NAND3_2713 ( P1_U5311 , P1_U5310 , P1_U5308 , P1_U5309 );
nand NAND2_2714 ( P1_U5312 , P1_U3045 , P1_U4024 );
nand NAND2_2715 ( P1_U5313 , P1_ADD_99_U67 , P1_U5769 );
nand NAND2_2716 ( P1_U5314 , P1_R1165_U11 , P1_U3026 );
nand NAND2_2717 ( P1_U5315 , P1_U4037 , P1_U5311 );
nand NAND2_2718 ( P1_U5316 , P1_REG3_REG_21_ , P1_U3086 );
nand NAND2_2719 ( P1_U5317 , P1_U3037 , P1_U3077 );
nand NAND2_2720 ( P1_U5318 , P1_U3035 , P1_U3068 );
nand NAND2_2721 ( P1_U5319 , P1_REG3_REG_1_ , P1_U3434 );
nand NAND3_2722 ( P1_U5320 , P1_U5318 , P1_U5317 , P1_U5319 );
nand NAND2_2723 ( P1_U5321 , P1_U3461 , P1_U5770 );
nand NAND2_2724 ( P1_U5322 , P1_REG3_REG_1_ , P1_U5769 );
nand NAND2_2725 ( P1_U5323 , P1_R1165_U101 , P1_U3026 );
nand NAND2_2726 ( P1_U5324 , P1_U4037 , P1_U5320 );
nand NAND2_2727 ( P1_U5325 , P1_REG3_REG_1_ , P1_U3086 );
nand NAND2_2728 ( P1_U5326 , P1_U3037 , P1_U3070 );
nand NAND2_2729 ( P1_U5327 , P1_U3035 , P1_U3083 );
nand NAND2_2730 ( P1_U5328 , P1_ADD_99_U55 , P1_U3434 );
nand NAND3_2731 ( P1_U5329 , P1_U5327 , P1_U5326 , P1_U5328 );
nand NAND2_2732 ( P1_U5330 , P1_U3482 , P1_U5770 );
nand NAND2_2733 ( P1_U5331 , P1_ADD_99_U55 , P1_U5769 );
nand NAND2_2734 ( P1_U5332 , P1_R1165_U89 , P1_U3026 );
nand NAND2_2735 ( P1_U5333 , P1_U4037 , P1_U5329 );
nand NAND2_2736 ( P1_U5334 , P1_REG3_REG_8_ , P1_U3086 );
nand NAND2_2737 ( P1_U5335 , P1_U3037 , P1_U3053 );
nand NAND2_2738 ( P1_U5336 , P1_U3035 , P1_U3055 );
nand NAND2_2739 ( P1_U5337 , P1_ADD_99_U60 , P1_U3434 );
nand NAND3_2740 ( P1_U5338 , P1_U5336 , P1_U5335 , P1_U5337 );
nand NAND2_2741 ( P1_U5339 , P1_U3045 , P1_U4017 );
nand NAND2_2742 ( P1_U5340 , P1_ADD_99_U60 , P1_U5769 );
nand NAND2_2743 ( P1_U5341 , P1_R1165_U94 , P1_U3026 );
nand NAND2_2744 ( P1_U5342 , P1_U4037 , P1_U5338 );
nand NAND2_2745 ( P1_U5343 , P1_REG3_REG_28_ , P1_U3086 );
nand NAND2_2746 ( P1_U5344 , P1_U3037 , P1_U3082 );
nand NAND2_2747 ( P1_U5345 , P1_U3035 , P1_U3076 );
nand NAND2_2748 ( P1_U5346 , P1_ADD_99_U69 , P1_U3434 );
nand NAND3_2749 ( P1_U5347 , P1_U5346 , P1_U5344 , P1_U5345 );
nand NAND2_2750 ( P1_U5348 , P1_U3514 , P1_U5770 );
nand NAND2_2751 ( P1_U5349 , P1_ADD_99_U69 , P1_U5769 );
nand NAND2_2752 ( P1_U5350 , P1_R1165_U102 , P1_U3026 );
nand NAND2_2753 ( P1_U5351 , P1_U4037 , P1_U5347 );
nand NAND2_2754 ( P1_U5352 , P1_REG3_REG_19_ , P1_U3086 );
nand NAND2_2755 ( P1_U5353 , P1_U3037 , P1_U3068 );
nand NAND2_2756 ( P1_U5354 , P1_U3035 , P1_U3060 );
nand NAND2_2757 ( P1_U5355 , P1_ADD_99_U4 , P1_U3434 );
nand NAND3_2758 ( P1_U5356 , P1_U5354 , P1_U5353 , P1_U5355 );
nand NAND2_2759 ( P1_U5357 , P1_U3467 , P1_U5770 );
nand NAND2_2760 ( P1_U5358 , P1_ADD_99_U4 , P1_U5769 );
nand NAND2_2761 ( P1_U5359 , P1_R1165_U13 , P1_U3026 );
nand NAND2_2762 ( P1_U5360 , P1_U4037 , P1_U5356 );
nand NAND2_2763 ( P1_U5361 , P1_REG3_REG_3_ , P1_U3086 );
nand NAND2_2764 ( P1_U5362 , P1_U3037 , P1_U3083 );
nand NAND2_2765 ( P1_U5363 , P1_U3035 , P1_U3063 );
nand NAND2_2766 ( P1_U5364 , P1_ADD_99_U78 , P1_U3434 );
nand NAND3_2767 ( P1_U5365 , P1_U5363 , P1_U5362 , P1_U5364 );
nand NAND2_2768 ( P1_U5366 , P1_U3488 , P1_U5770 );
nand NAND2_2769 ( P1_U5367 , P1_ADD_99_U78 , P1_U5769 );
nand NAND2_2770 ( P1_U5368 , P1_R1165_U109 , P1_U3026 );
nand NAND2_2771 ( P1_U5369 , P1_U4037 , P1_U5365 );
nand NAND2_2772 ( P1_U5370 , P1_REG3_REG_10_ , P1_U3086 );
nand NAND2_2773 ( P1_U5371 , P1_U3037 , P1_U3061 );
nand NAND2_2774 ( P1_U5372 , P1_U3035 , P1_U3065 );
nand NAND2_2775 ( P1_U5373 , P1_ADD_99_U65 , P1_U3434 );
nand NAND3_2776 ( P1_U5374 , P1_U5373 , P1_U5371 , P1_U5372 );
nand NAND2_2777 ( P1_U5375 , P1_U3045 , P1_U4022 );
nand NAND2_2778 ( P1_U5376 , P1_ADD_99_U65 , P1_U5769 );
nand NAND2_2779 ( P1_U5377 , P1_R1165_U98 , P1_U3026 );
nand NAND2_2780 ( P1_U5378 , P1_U4037 , P1_U5374 );
nand NAND2_2781 ( P1_U5379 , P1_REG3_REG_23_ , P1_U3086 );
nand NAND2_2782 ( P1_U5380 , P1_U3037 , P1_U3080 );
nand NAND2_2783 ( P1_U5381 , P1_U3035 , P1_U3074 );
nand NAND2_2784 ( P1_U5382 , P1_ADD_99_U74 , P1_U3434 );
nand NAND3_2785 ( P1_U5383 , P1_U5382 , P1_U5380 , P1_U5381 );
nand NAND2_2786 ( P1_U5384 , P1_U3500 , P1_U5770 );
nand NAND2_2787 ( P1_U5385 , P1_ADD_99_U74 , P1_U5769 );
nand NAND2_2788 ( P1_U5386 , P1_R1165_U106 , P1_U3026 );
nand NAND2_2789 ( P1_U5387 , P1_U4037 , P1_U5383 );
nand NAND2_2790 ( P1_U5388 , P1_REG3_REG_14_ , P1_U3086 );
nand NAND2_2791 ( P1_U5389 , P1_U3037 , P1_U3057 );
nand NAND2_2792 ( P1_U5390 , P1_U3035 , P1_U3054 );
nand NAND2_2793 ( P1_U5391 , P1_ADD_99_U61 , P1_U3434 );
nand NAND3_2794 ( P1_U5392 , P1_U5391 , P1_U5389 , P1_U5390 );
nand NAND2_2795 ( P1_U5393 , P1_U3045 , P1_U4018 );
nand NAND2_2796 ( P1_U5394 , P1_ADD_99_U61 , P1_U5769 );
nand NAND2_2797 ( P1_U5395 , P1_R1165_U95 , P1_U3026 );
nand NAND2_2798 ( P1_U5396 , P1_U4037 , P1_U5392 );
nand NAND2_2799 ( P1_U5397 , P1_REG3_REG_27_ , P1_U3086 );
nand NAND2_2800 ( P1_U5398 , P1_U3037 , P1_U3071 );
nand NAND2_2801 ( P1_U5399 , P1_U3035 , P1_U3084 );
nand NAND2_2802 ( P1_U5400 , P1_ADD_99_U56 , P1_U3434 );
nand NAND3_2803 ( P1_U5401 , P1_U5399 , P1_U5398 , P1_U5400 );
nand NAND2_2804 ( P1_U5402 , P1_U3479 , P1_U5770 );
nand NAND2_2805 ( P1_U5403 , P1_ADD_99_U56 , P1_U5769 );
nand NAND2_2806 ( P1_U5404 , P1_R1165_U14 , P1_U3026 );
nand NAND2_2807 ( P1_U5405 , P1_U4037 , P1_U5401 );
nand NAND2_2808 ( P1_U5406 , P1_REG3_REG_7_ , P1_U3086 );
nand NAND2_2809 ( P1_U5407 , P1_U3455 , P1_U3377 );
nand NAND2_2810 ( P1_U5408 , P1_U3449 , P1_U5407 );
nand NAND3_2811 ( P1_U5409 , P1_U5817 , P1_U3449 , P1_R1165_U87 );
nand NAND2_2812 ( P1_U5410 , P1_U3450 , P1_U3453 );
nand NAND2_2813 ( P1_U5411 , P1_U3874 , P1_U4013 );
nand NAND2_2814 ( P1_U5412 , P1_U3370 , P1_U3422 );
nand NAND3_2815 ( P1_U5413 , P1_U4006 , P1_U3363 , P1_U3365 );
nand NAND2_2816 ( P1_U5414 , P1_U4041 , P1_U3425 );
nand NAND2_2817 ( P1_U5415 , P1_U5413 , P1_U3425 );
not NOT1_2818 ( P1_U5416 , P1_U3436 );
nand NAND2_2819 ( P1_U5417 , P1_U5416 , P1_U4013 );
nand NAND2_2820 ( P1_U5418 , P1_U3485 , P1_U5417 );
nand NAND2_2821 ( P1_U5419 , P1_U3021 , P1_U3083 );
nand NAND2_2822 ( P1_U5420 , P1_U3482 , P1_U5417 );
nand NAND2_2823 ( P1_U5421 , P1_U3021 , P1_U3084 );
nand NAND2_2824 ( P1_U5422 , P1_U3479 , P1_U5417 );
nand NAND2_2825 ( P1_U5423 , P1_U3021 , P1_U3070 );
nand NAND2_2826 ( P1_U5424 , P1_U3476 , P1_U5417 );
nand NAND2_2827 ( P1_U5425 , P1_U3021 , P1_U3071 );
nand NAND2_2828 ( P1_U5426 , P1_U3473 , P1_U5417 );
nand NAND2_2829 ( P1_U5427 , P1_U3021 , P1_U3067 );
nand NAND2_2830 ( P1_U5428 , P1_U3470 , P1_U5417 );
nand NAND2_2831 ( P1_U5429 , P1_U3021 , P1_U3060 );
nand NAND2_2832 ( P1_U5430 , P1_U3467 , P1_U5417 );
nand NAND2_2833 ( P1_U5431 , P1_U3021 , P1_U3064 );
nand NAND2_2834 ( P1_U5432 , P1_U4017 , P1_U5417 );
nand NAND2_2835 ( P1_U5433 , P1_U3021 , P1_U3054 );
nand NAND2_2836 ( P1_U5434 , P1_U4018 , P1_U5417 );
nand NAND2_2837 ( P1_U5435 , P1_U3021 , P1_U3053 );
nand NAND2_2838 ( P1_U5436 , P1_U4019 , P1_U5417 );
nand NAND2_2839 ( P1_U5437 , P1_U3021 , P1_U3057 );
nand NAND2_2840 ( P1_U5438 , P1_U4020 , P1_U5417 );
nand NAND2_2841 ( P1_U5439 , P1_U3021 , P1_U3058 );
nand NAND2_2842 ( P1_U5440 , P1_U4021 , P1_U5417 );
nand NAND2_2843 ( P1_U5441 , P1_U3021 , P1_U3065 );
nand NAND2_2844 ( P1_U5442 , P1_U4022 , P1_U5417 );
nand NAND2_2845 ( P1_U5443 , P1_U3021 , P1_U3066 );
nand NAND2_2846 ( P1_U5444 , P1_U4023 , P1_U5417 );
nand NAND2_2847 ( P1_U5445 , P1_U3021 , P1_U3061 );
nand NAND2_2848 ( P1_U5446 , P1_U4024 , P1_U5417 );
nand NAND2_2849 ( P1_U5447 , P1_U3021 , P1_U3075 );
nand NAND2_2850 ( P1_U5448 , P1_U4025 , P1_U5417 );
nand NAND2_2851 ( P1_U5449 , P1_U3021 , P1_U3076 );
nand NAND2_2852 ( P1_U5450 , P1_U3464 , P1_U5417 );
nand NAND2_2853 ( P1_U5451 , P1_U3021 , P1_U3068 );
nand NAND2_2854 ( P1_U5452 , P1_U3514 , P1_U5417 );
nand NAND2_2855 ( P1_U5453 , P1_U3021 , P1_U3081 );
nand NAND2_2856 ( P1_U5454 , P1_U3512 , P1_U5417 );
nand NAND2_2857 ( P1_U5455 , P1_U3021 , P1_U3082 );
nand NAND2_2858 ( P1_U5456 , P1_U3509 , P1_U5417 );
nand NAND2_2859 ( P1_U5457 , P1_U3021 , P1_U3069 );
nand NAND2_2860 ( P1_U5458 , P1_U3506 , P1_U5417 );
nand NAND2_2861 ( P1_U5459 , P1_U3021 , P1_U3073 );
nand NAND2_2862 ( P1_U5460 , P1_U3503 , P1_U5417 );
nand NAND2_2863 ( P1_U5461 , P1_U3021 , P1_U3074 );
nand NAND2_2864 ( P1_U5462 , P1_U3500 , P1_U5417 );
nand NAND2_2865 ( P1_U5463 , P1_U3021 , P1_U3079 );
nand NAND2_2866 ( P1_U5464 , P1_U3497 , P1_U5417 );
nand NAND2_2867 ( P1_U5465 , P1_U3021 , P1_U3080 );
nand NAND2_2868 ( P1_U5466 , P1_U3494 , P1_U5417 );
nand NAND2_2869 ( P1_U5467 , P1_U3021 , P1_U3072 );
nand NAND2_2870 ( P1_U5468 , P1_U3491 , P1_U5417 );
nand NAND2_2871 ( P1_U5469 , P1_U3021 , P1_U3063 );
nand NAND2_2872 ( P1_U5470 , P1_U3488 , P1_U5417 );
nand NAND2_2873 ( P1_U5471 , P1_U3021 , P1_U3062 );
nand NAND2_2874 ( P1_U5472 , P1_U3461 , P1_U5417 );
nand NAND2_2875 ( P1_U5473 , P1_U3021 , P1_U3078 );
nand NAND2_2876 ( P1_U5474 , P1_U3456 , P1_U5417 );
nand NAND2_2877 ( P1_U5475 , P1_U3021 , P1_U3077 );
nand NAND2_2878 ( P1_U5476 , P1_U4145 , P1_REG1_REG_0_ );
nand NAND2_2879 ( P1_U5477 , P1_U3021 , P1_U3485 );
nand NAND2_2880 ( P1_U5478 , P1_U3436 , P1_U3083 );
nand NAND2_2881 ( P1_U5479 , P1_U3021 , P1_U3482 );
nand NAND2_2882 ( P1_U5480 , P1_U3436 , P1_U3084 );
nand NAND2_2883 ( P1_U5481 , P1_U3021 , P1_U3479 );
nand NAND2_2884 ( P1_U5482 , P1_U3436 , P1_U3070 );
nand NAND2_2885 ( P1_U5483 , P1_U3021 , P1_U3476 );
nand NAND2_2886 ( P1_U5484 , P1_U3436 , P1_U3071 );
nand NAND2_2887 ( P1_U5485 , P1_U3021 , P1_U3473 );
nand NAND2_2888 ( P1_U5486 , P1_U3436 , P1_U3067 );
nand NAND2_2889 ( P1_U5487 , P1_U3021 , P1_U3470 );
nand NAND2_2890 ( P1_U5488 , P1_U3436 , P1_U3060 );
nand NAND2_2891 ( P1_U5489 , P1_U3021 , P1_U3467 );
nand NAND2_2892 ( P1_U5490 , P1_U3436 , P1_U3064 );
nand NAND2_2893 ( P1_U5491 , P1_U3021 , P1_U4017 );
nand NAND2_2894 ( P1_U5492 , P1_U3436 , P1_U3054 );
nand NAND2_2895 ( P1_U5493 , P1_U3021 , P1_U4018 );
nand NAND2_2896 ( P1_U5494 , P1_U3436 , P1_U3053 );
nand NAND2_2897 ( P1_U5495 , P1_U3021 , P1_U4019 );
nand NAND2_2898 ( P1_U5496 , P1_U3436 , P1_U3057 );
nand NAND2_2899 ( P1_U5497 , P1_U3021 , P1_U4020 );
nand NAND2_2900 ( P1_U5498 , P1_U3436 , P1_U3058 );
nand NAND2_2901 ( P1_U5499 , P1_U3021 , P1_U4021 );
nand NAND2_2902 ( P1_U5500 , P1_U3436 , P1_U3065 );
nand NAND2_2903 ( P1_U5501 , P1_U3021 , P1_U4022 );
nand NAND2_2904 ( P1_U5502 , P1_U3436 , P1_U3066 );
nand NAND2_2905 ( P1_U5503 , P1_U3021 , P1_U4023 );
nand NAND2_2906 ( P1_U5504 , P1_U3436 , P1_U3061 );
nand NAND2_2907 ( P1_U5505 , P1_U3021 , P1_U4024 );
nand NAND2_2908 ( P1_U5506 , P1_U3436 , P1_U3075 );
nand NAND2_2909 ( P1_U5507 , P1_U3021 , P1_U4025 );
nand NAND2_2910 ( P1_U5508 , P1_U3436 , P1_U3076 );
nand NAND2_2911 ( P1_U5509 , P1_U3021 , P1_U3464 );
nand NAND2_2912 ( P1_U5510 , P1_U3436 , P1_U3068 );
nand NAND2_2913 ( P1_U5511 , P1_U3021 , P1_U3514 );
nand NAND2_2914 ( P1_U5512 , P1_U3436 , P1_U3081 );
nand NAND2_2915 ( P1_U5513 , P1_U3021 , P1_U3512 );
nand NAND2_2916 ( P1_U5514 , P1_U3436 , P1_U3082 );
nand NAND2_2917 ( P1_U5515 , P1_U3021 , P1_U3509 );
nand NAND2_2918 ( P1_U5516 , P1_U3436 , P1_U3069 );
nand NAND2_2919 ( P1_U5517 , P1_U3021 , P1_U3506 );
nand NAND2_2920 ( P1_U5518 , P1_U3436 , P1_U3073 );
nand NAND2_2921 ( P1_U5519 , P1_U3021 , P1_U3503 );
nand NAND2_2922 ( P1_U5520 , P1_U3436 , P1_U3074 );
nand NAND2_2923 ( P1_U5521 , P1_U3021 , P1_U3500 );
nand NAND2_2924 ( P1_U5522 , P1_U3436 , P1_U3079 );
nand NAND2_2925 ( P1_U5523 , P1_U3021 , P1_U3497 );
nand NAND2_2926 ( P1_U5524 , P1_U3436 , P1_U3080 );
nand NAND2_2927 ( P1_U5525 , P1_U3021 , P1_U3494 );
nand NAND2_2928 ( P1_U5526 , P1_U3436 , P1_U3072 );
nand NAND2_2929 ( P1_U5527 , P1_U3021 , P1_U3491 );
nand NAND2_2930 ( P1_U5528 , P1_U3436 , P1_U3063 );
nand NAND2_2931 ( P1_U5529 , P1_U3021 , P1_U3488 );
nand NAND2_2932 ( P1_U5530 , P1_U3436 , P1_U3062 );
nand NAND2_2933 ( P1_U5531 , P1_U3021 , P1_U3461 );
nand NAND2_2934 ( P1_U5532 , P1_U3436 , P1_U3078 );
nand NAND2_2935 ( P1_U5533 , P1_U3021 , P1_U3456 );
nand NAND2_2936 ( P1_U5534 , P1_U3436 , P1_U3077 );
nand NAND2_2937 ( P1_U5535 , P1_U4145 , P1_U3454 );
not NOT1_2938 ( P1_U5536 , P1_U3437 );
not NOT1_2939 ( P1_U5537 , P1_U3438 );
nand NAND2_2940 ( P1_U5538 , P1_U5799 , P1_U3450 );
nand NAND2_2941 ( P1_U5539 , P1_U3437 , P1_U3439 );
nand NAND2_2942 ( P1_U5540 , P1_U3051 , P1_U5539 );
nand NAND2_2943 ( P1_U5541 , P1_U3014 , P1_U3444 );
not NOT1_2944 ( P1_U5542 , P1_U3440 );
nand NAND2_2945 ( P1_U5543 , P1_U3052 , P1_U5542 );
nand NAND2_2946 ( P1_U5544 , P1_U3083 , P1_U3027 );
nand NAND2_2947 ( P1_U5545 , P1_U3485 , P1_U5543 );
nand NAND2_2948 ( P1_U5546 , P1_U5540 , P1_U3083 );
nand NAND2_2949 ( P1_U5547 , P1_U3084 , P1_U3027 );
nand NAND2_2950 ( P1_U5548 , P1_U3482 , P1_U5543 );
nand NAND2_2951 ( P1_U5549 , P1_U5540 , P1_U3084 );
nand NAND2_2952 ( P1_U5550 , P1_U3070 , P1_U3027 );
nand NAND2_2953 ( P1_U5551 , P1_U3479 , P1_U5543 );
nand NAND2_2954 ( P1_U5552 , P1_U5540 , P1_U3070 );
nand NAND2_2955 ( P1_U5553 , P1_U3071 , P1_U3027 );
nand NAND2_2956 ( P1_U5554 , P1_U3476 , P1_U5543 );
nand NAND2_2957 ( P1_U5555 , P1_U5540 , P1_U3071 );
nand NAND2_2958 ( P1_U5556 , P1_U3067 , P1_U3027 );
nand NAND2_2959 ( P1_U5557 , P1_U3473 , P1_U5543 );
nand NAND2_2960 ( P1_U5558 , P1_U5540 , P1_U3067 );
nand NAND2_2961 ( P1_U5559 , P1_U3060 , P1_U3027 );
nand NAND2_2962 ( P1_U5560 , P1_U3470 , P1_U5543 );
nand NAND2_2963 ( P1_U5561 , P1_U5540 , P1_U3060 );
nand NAND2_2964 ( P1_U5562 , P1_R1309_U8 , P1_U3027 );
nand NAND2_2965 ( P1_U5563 , P1_U4026 , P1_U5543 );
nand NAND2_2966 ( P1_U5564 , P1_U5540 , P1_U3056 );
nand NAND2_2967 ( P1_U5565 , P1_R1309_U6 , P1_U3027 );
nand NAND2_2968 ( P1_U5566 , P1_U4027 , P1_U5543 );
nand NAND2_2969 ( P1_U5567 , P1_U5540 , P1_U3059 );
nand NAND2_2970 ( P1_U5568 , P1_U3064 , P1_U3027 );
nand NAND2_2971 ( P1_U5569 , P1_U3467 , P1_U5543 );
nand NAND2_2972 ( P1_U5570 , P1_U5540 , P1_U3064 );
nand NAND2_2973 ( P1_U5571 , P1_U3055 , P1_U3027 );
nand NAND2_2974 ( P1_U5572 , P1_U4028 , P1_U5543 );
nand NAND2_2975 ( P1_U5573 , P1_U5540 , P1_U3055 );
nand NAND2_2976 ( P1_U5574 , P1_U3054 , P1_U3027 );
nand NAND2_2977 ( P1_U5575 , P1_U4017 , P1_U5543 );
nand NAND2_2978 ( P1_U5576 , P1_U5540 , P1_U3054 );
nand NAND2_2979 ( P1_U5577 , P1_U3053 , P1_U3027 );
nand NAND2_2980 ( P1_U5578 , P1_U4018 , P1_U5543 );
nand NAND2_2981 ( P1_U5579 , P1_U5540 , P1_U3053 );
nand NAND2_2982 ( P1_U5580 , P1_U3057 , P1_U3027 );
nand NAND2_2983 ( P1_U5581 , P1_U4019 , P1_U5543 );
nand NAND2_2984 ( P1_U5582 , P1_U5540 , P1_U3057 );
nand NAND2_2985 ( P1_U5583 , P1_U3058 , P1_U3027 );
nand NAND2_2986 ( P1_U5584 , P1_U4020 , P1_U5543 );
nand NAND2_2987 ( P1_U5585 , P1_U5540 , P1_U3058 );
nand NAND2_2988 ( P1_U5586 , P1_U3065 , P1_U3027 );
nand NAND2_2989 ( P1_U5587 , P1_U4021 , P1_U5543 );
nand NAND2_2990 ( P1_U5588 , P1_U5540 , P1_U3065 );
nand NAND2_2991 ( P1_U5589 , P1_U3066 , P1_U3027 );
nand NAND2_2992 ( P1_U5590 , P1_U4022 , P1_U5543 );
nand NAND2_2993 ( P1_U5591 , P1_U5540 , P1_U3066 );
nand NAND2_2994 ( P1_U5592 , P1_U3061 , P1_U3027 );
nand NAND2_2995 ( P1_U5593 , P1_U4023 , P1_U5543 );
nand NAND2_2996 ( P1_U5594 , P1_U5540 , P1_U3061 );
nand NAND2_2997 ( P1_U5595 , P1_U3075 , P1_U3027 );
nand NAND2_2998 ( P1_U5596 , P1_U4024 , P1_U5543 );
nand NAND2_2999 ( P1_U5597 , P1_U5540 , P1_U3075 );
nand NAND2_3000 ( P1_U5598 , P1_U3076 , P1_U3027 );
nand NAND2_3001 ( P1_U5599 , P1_U4025 , P1_U5543 );
nand NAND2_3002 ( P1_U5600 , P1_U5540 , P1_U3076 );
nand NAND2_3003 ( P1_U5601 , P1_U3068 , P1_U3027 );
nand NAND2_3004 ( P1_U5602 , P1_U3464 , P1_U5543 );
nand NAND2_3005 ( P1_U5603 , P1_U5540 , P1_U3068 );
nand NAND2_3006 ( P1_U5604 , P1_U3081 , P1_U3027 );
nand NAND2_3007 ( P1_U5605 , P1_U3514 , P1_U5543 );
nand NAND2_3008 ( P1_U5606 , P1_U5540 , P1_U3081 );
nand NAND2_3009 ( P1_U5607 , P1_U3082 , P1_U3027 );
nand NAND2_3010 ( P1_U5608 , P1_U3512 , P1_U5543 );
nand NAND2_3011 ( P1_U5609 , P1_U5540 , P1_U3082 );
nand NAND2_3012 ( P1_U5610 , P1_U3069 , P1_U3027 );
nand NAND2_3013 ( P1_U5611 , P1_U3509 , P1_U5543 );
nand NAND2_3014 ( P1_U5612 , P1_U5540 , P1_U3069 );
nand NAND2_3015 ( P1_U5613 , P1_U3073 , P1_U3027 );
nand NAND2_3016 ( P1_U5614 , P1_U3506 , P1_U5543 );
nand NAND2_3017 ( P1_U5615 , P1_U5540 , P1_U3073 );
nand NAND2_3018 ( P1_U5616 , P1_U3074 , P1_U3027 );
nand NAND2_3019 ( P1_U5617 , P1_U3503 , P1_U5543 );
nand NAND2_3020 ( P1_U5618 , P1_U5540 , P1_U3074 );
nand NAND2_3021 ( P1_U5619 , P1_U3079 , P1_U3027 );
nand NAND2_3022 ( P1_U5620 , P1_U3500 , P1_U5543 );
nand NAND2_3023 ( P1_U5621 , P1_U5540 , P1_U3079 );
nand NAND2_3024 ( P1_U5622 , P1_U3080 , P1_U3027 );
nand NAND2_3025 ( P1_U5623 , P1_U3497 , P1_U5543 );
nand NAND2_3026 ( P1_U5624 , P1_U5540 , P1_U3080 );
nand NAND2_3027 ( P1_U5625 , P1_U3072 , P1_U3027 );
nand NAND2_3028 ( P1_U5626 , P1_U3494 , P1_U5543 );
nand NAND2_3029 ( P1_U5627 , P1_U5540 , P1_U3072 );
nand NAND2_3030 ( P1_U5628 , P1_U3063 , P1_U3027 );
nand NAND2_3031 ( P1_U5629 , P1_U3491 , P1_U5543 );
nand NAND2_3032 ( P1_U5630 , P1_U5540 , P1_U3063 );
nand NAND2_3033 ( P1_U5631 , P1_U3062 , P1_U3027 );
nand NAND2_3034 ( P1_U5632 , P1_U3488 , P1_U5543 );
nand NAND2_3035 ( P1_U5633 , P1_U5540 , P1_U3062 );
nand NAND2_3036 ( P1_U5634 , P1_U3078 , P1_U3027 );
nand NAND2_3037 ( P1_U5635 , P1_U3461 , P1_U5543 );
nand NAND2_3038 ( P1_U5636 , P1_U5540 , P1_U3078 );
nand NAND2_3039 ( P1_U5637 , P1_U3077 , P1_U3027 );
nand NAND2_3040 ( P1_U5638 , P1_U3456 , P1_U5543 );
nand NAND2_3041 ( P1_U5639 , P1_U5540 , P1_U3077 );
nand NAND2_3042 ( P1_U5640 , P1_U3440 , P1_U3439 );
nand NAND2_3043 ( P1_U5641 , P1_U3052 , P1_U5640 );
nand NAND2_3044 ( P1_U5642 , P1_U3028 , P1_U3083 );
nand NAND2_3045 ( P1_U5643 , P1_U3485 , P1_U3438 );
nand NAND2_3046 ( P1_U5644 , P1_U5641 , P1_U3083 );
nand NAND2_3047 ( P1_U5645 , P1_U5786 , P1_U3084 );
nand NAND2_3048 ( P1_U5646 , P1_U3028 , P1_U3084 );
nand NAND2_3049 ( P1_U5647 , P1_U3482 , P1_U3438 );
nand NAND2_3050 ( P1_U5648 , P1_U5641 , P1_U3084 );
nand NAND2_3051 ( P1_U5649 , P1_U5786 , P1_U3070 );
nand NAND2_3052 ( P1_U5650 , P1_U3028 , P1_U3070 );
nand NAND2_3053 ( P1_U5651 , P1_U3479 , P1_U3438 );
nand NAND2_3054 ( P1_U5652 , P1_U5641 , P1_U3070 );
nand NAND2_3055 ( P1_U5653 , P1_U5786 , P1_U3071 );
nand NAND2_3056 ( P1_U5654 , P1_U3028 , P1_U3071 );
nand NAND2_3057 ( P1_U5655 , P1_U3476 , P1_U3438 );
nand NAND2_3058 ( P1_U5656 , P1_U5641 , P1_U3071 );
nand NAND2_3059 ( P1_U5657 , P1_U5786 , P1_U3067 );
nand NAND2_3060 ( P1_U5658 , P1_U3028 , P1_U3067 );
nand NAND2_3061 ( P1_U5659 , P1_U3473 , P1_U3438 );
nand NAND2_3062 ( P1_U5660 , P1_U5641 , P1_U3067 );
nand NAND2_3063 ( P1_U5661 , P1_U5786 , P1_U3060 );
nand NAND2_3064 ( P1_U5662 , P1_U3028 , P1_U3060 );
nand NAND2_3065 ( P1_U5663 , P1_U3470 , P1_U3438 );
nand NAND2_3066 ( P1_U5664 , P1_U5641 , P1_U3060 );
nand NAND2_3067 ( P1_U5665 , P1_U5786 , P1_U3064 );
nand NAND2_3068 ( P1_U5666 , P1_U3028 , P1_R1309_U8 );
nand NAND2_3069 ( P1_U5667 , P1_U4026 , P1_U3438 );
nand NAND2_3070 ( P1_U5668 , P1_U5641 , P1_U3056 );
nand NAND2_3071 ( P1_U5669 , P1_U3028 , P1_R1309_U6 );
nand NAND2_3072 ( P1_U5670 , P1_U4027 , P1_U3438 );
nand NAND2_3073 ( P1_U5671 , P1_U5641 , P1_U3059 );
nand NAND2_3074 ( P1_U5672 , P1_U3028 , P1_U3064 );
nand NAND2_3075 ( P1_U5673 , P1_U3467 , P1_U3438 );
nand NAND2_3076 ( P1_U5674 , P1_U5641 , P1_U3064 );
nand NAND2_3077 ( P1_U5675 , P1_U5786 , P1_U3068 );
nand NAND2_3078 ( P1_U5676 , P1_U3028 , P1_U3055 );
nand NAND2_3079 ( P1_U5677 , P1_U4028 , P1_U3438 );
nand NAND2_3080 ( P1_U5678 , P1_U5641 , P1_U3055 );
nand NAND2_3081 ( P1_U5679 , P1_U5786 , P1_U3054 );
nand NAND2_3082 ( P1_U5680 , P1_U3028 , P1_U3054 );
nand NAND2_3083 ( P1_U5681 , P1_U4017 , P1_U3438 );
nand NAND2_3084 ( P1_U5682 , P1_U5641 , P1_U3054 );
nand NAND2_3085 ( P1_U5683 , P1_U5786 , P1_U3053 );
nand NAND2_3086 ( P1_U5684 , P1_U3028 , P1_U3053 );
nand NAND2_3087 ( P1_U5685 , P1_U4018 , P1_U3438 );
nand NAND2_3088 ( P1_U5686 , P1_U5641 , P1_U3053 );
nand NAND2_3089 ( P1_U5687 , P1_U5786 , P1_U3057 );
nand NAND2_3090 ( P1_U5688 , P1_U3028 , P1_U3057 );
nand NAND2_3091 ( P1_U5689 , P1_U4019 , P1_U3438 );
nand NAND2_3092 ( P1_U5690 , P1_U5641 , P1_U3057 );
nand NAND2_3093 ( P1_U5691 , P1_U5786 , P1_U3058 );
nand NAND2_3094 ( P1_U5692 , P1_U3028 , P1_U3058 );
nand NAND2_3095 ( P1_U5693 , P1_U4020 , P1_U3438 );
nand NAND2_3096 ( P1_U5694 , P1_U5641 , P1_U3058 );
nand NAND2_3097 ( P1_U5695 , P1_U5786 , P1_U3065 );
nand NAND2_3098 ( P1_U5696 , P1_U3028 , P1_U3065 );
nand NAND2_3099 ( P1_U5697 , P1_U4021 , P1_U3438 );
nand NAND2_3100 ( P1_U5698 , P1_U5641 , P1_U3065 );
nand NAND2_3101 ( P1_U5699 , P1_U5786 , P1_U3066 );
nand NAND2_3102 ( P1_U5700 , P1_U3028 , P1_U3066 );
nand NAND2_3103 ( P1_U5701 , P1_U4022 , P1_U3438 );
nand NAND2_3104 ( P1_U5702 , P1_U5641 , P1_U3066 );
nand NAND2_3105 ( P1_U5703 , P1_U5786 , P1_U3061 );
nand NAND2_3106 ( P1_U5704 , P1_U3028 , P1_U3061 );
nand NAND2_3107 ( P1_U5705 , P1_U4023 , P1_U3438 );
nand NAND2_3108 ( P1_U5706 , P1_U5641 , P1_U3061 );
nand NAND2_3109 ( P1_U5707 , P1_U5786 , P1_U3075 );
nand NAND2_3110 ( P1_U5708 , P1_U3028 , P1_U3075 );
nand NAND2_3111 ( P1_U5709 , P1_U4024 , P1_U3438 );
nand NAND2_3112 ( P1_U5710 , P1_U5641 , P1_U3075 );
nand NAND2_3113 ( P1_U5711 , P1_U5786 , P1_U3076 );
nand NAND2_3114 ( P1_U5712 , P1_U3028 , P1_U3076 );
nand NAND2_3115 ( P1_U5713 , P1_U4025 , P1_U3438 );
nand NAND2_3116 ( P1_U5714 , P1_U5641 , P1_U3076 );
nand NAND2_3117 ( P1_U5715 , P1_U5786 , P1_U3081 );
nand NAND2_3118 ( P1_U5716 , P1_U3028 , P1_U3068 );
nand NAND2_3119 ( P1_U5717 , P1_U3464 , P1_U3438 );
nand NAND2_3120 ( P1_U5718 , P1_U5641 , P1_U3068 );
nand NAND2_3121 ( P1_U5719 , P1_U5786 , P1_U3078 );
nand NAND2_3122 ( P1_U5720 , P1_U3028 , P1_U3081 );
nand NAND2_3123 ( P1_U5721 , P1_U3514 , P1_U3438 );
nand NAND2_3124 ( P1_U5722 , P1_U5641 , P1_U3081 );
nand NAND2_3125 ( P1_U5723 , P1_U5786 , P1_U3082 );
nand NAND2_3126 ( P1_U5724 , P1_U3028 , P1_U3082 );
nand NAND2_3127 ( P1_U5725 , P1_U3512 , P1_U3438 );
nand NAND2_3128 ( P1_U5726 , P1_U5641 , P1_U3082 );
nand NAND2_3129 ( P1_U5727 , P1_U5786 , P1_U3069 );
nand NAND2_3130 ( P1_U5728 , P1_U3028 , P1_U3069 );
nand NAND2_3131 ( P1_U5729 , P1_U3509 , P1_U3438 );
nand NAND2_3132 ( P1_U5730 , P1_U5641 , P1_U3069 );
nand NAND2_3133 ( P1_U5731 , P1_U5786 , P1_U3073 );
nand NAND2_3134 ( P1_U5732 , P1_U3028 , P1_U3073 );
nand NAND2_3135 ( P1_U5733 , P1_U3506 , P1_U3438 );
nand NAND2_3136 ( P1_U5734 , P1_U5641 , P1_U3073 );
nand NAND2_3137 ( P1_U5735 , P1_U5786 , P1_U3074 );
nand NAND2_3138 ( P1_U5736 , P1_U3028 , P1_U3074 );
nand NAND2_3139 ( P1_U5737 , P1_U3503 , P1_U3438 );
nand NAND2_3140 ( P1_U5738 , P1_U5641 , P1_U3074 );
nand NAND2_3141 ( P1_U5739 , P1_U5786 , P1_U3079 );
nand NAND2_3142 ( P1_U5740 , P1_U3028 , P1_U3079 );
nand NAND2_3143 ( P1_U5741 , P1_U3500 , P1_U3438 );
nand NAND2_3144 ( P1_U5742 , P1_U5641 , P1_U3079 );
nand NAND2_3145 ( P1_U5743 , P1_U5786 , P1_U3080 );
nand NAND2_3146 ( P1_U5744 , P1_U3028 , P1_U3080 );
nand NAND2_3147 ( P1_U5745 , P1_U3497 , P1_U3438 );
nand NAND2_3148 ( P1_U5746 , P1_U5641 , P1_U3080 );
nand NAND2_3149 ( P1_U5747 , P1_U5786 , P1_U3072 );
nand NAND2_3150 ( P1_U5748 , P1_U3028 , P1_U3072 );
nand NAND2_3151 ( P1_U5749 , P1_U3494 , P1_U3438 );
nand NAND2_3152 ( P1_U5750 , P1_U5641 , P1_U3072 );
nand NAND2_3153 ( P1_U5751 , P1_U5786 , P1_U3063 );
nand NAND2_3154 ( P1_U5752 , P1_U3028 , P1_U3063 );
nand NAND2_3155 ( P1_U5753 , P1_U3491 , P1_U3438 );
nand NAND2_3156 ( P1_U5754 , P1_U5641 , P1_U3063 );
nand NAND2_3157 ( P1_U5755 , P1_U5786 , P1_U3062 );
nand NAND2_3158 ( P1_U5756 , P1_U3028 , P1_U3062 );
nand NAND2_3159 ( P1_U5757 , P1_U3488 , P1_U3438 );
nand NAND2_3160 ( P1_U5758 , P1_U5641 , P1_U3062 );
nand NAND2_3161 ( P1_U5759 , P1_U5786 , P1_U3083 );
nand NAND2_3162 ( P1_U5760 , P1_U3028 , P1_U3078 );
nand NAND2_3163 ( P1_U5761 , P1_U3461 , P1_U3438 );
nand NAND2_3164 ( P1_U5762 , P1_U5641 , P1_U3078 );
nand NAND2_3165 ( P1_U5763 , P1_U5786 , P1_U3077 );
nand NAND2_3166 ( P1_U5764 , P1_U3028 , P1_U3077 );
nand NAND2_3167 ( P1_U5765 , P1_U3456 , P1_U3438 );
nand NAND2_3168 ( P1_U5766 , P1_U5641 , P1_U3077 );
nand NAND2_3169 ( P1_U5767 , P1_U4038 , P1_U3434 );
nand NAND2_3170 ( P1_U5768 , P1_U4015 , P1_U4038 );
nand NAND2_3171 ( P1_U5769 , P1_U3050 , P1_U5767 );
nand NAND2_3172 ( P1_U5770 , P1_U5768 , P1_U4039 );
nand NAND2_3173 ( P1_U5771 , P1_U5775 , P1_U5781 );
nand NAND2_3174 ( P1_U5772 , P1_R1375_U9 , P1_U5131 );
nand NAND2_3175 ( P1_U5773 , P1_IR_REG_24_ , P1_U3952 );
nand NAND2_3176 ( P1_U5774 , P1_IR_REG_31_ , P1_SUB_88_U17 );
not NOT1_3177 ( P1_U5775 , P1_U3441 );
nand NAND2_3178 ( P1_U5776 , P1_IR_REG_25_ , P1_U3952 );
nand NAND2_3179 ( P1_U5777 , P1_IR_REG_31_ , P1_SUB_88_U170 );
not NOT1_3180 ( P1_U5778 , P1_U3442 );
nand NAND2_3181 ( P1_U5779 , P1_IR_REG_26_ , P1_U3952 );
nand NAND2_3182 ( P1_U5780 , P1_IR_REG_31_ , P1_SUB_88_U18 );
not NOT1_3183 ( P1_U5781 , P1_U3443 );
nand NAND2_3184 ( P1_U5782 , P1_U3441 , P1_U3359 );
nand NAND3_3185 ( P1_U5783 , P1_U4046 , P1_U5775 , P1_B_REG );
nand NAND2_3186 ( P1_U5784 , P1_IR_REG_23_ , P1_U3952 );
nand NAND2_3187 ( P1_U5785 , P1_IR_REG_31_ , P1_SUB_88_U16 );
not NOT1_3188 ( P1_U5786 , P1_U3444 );
nand NAND2_3189 ( P1_U5787 , P1_D_REG_0_ , P1_U3953 );
nand NAND2_3190 ( P1_U5788 , P1_U4034 , P1_U4146 );
nand NAND2_3191 ( P1_U5789 , P1_D_REG_1_ , P1_U3953 );
nand NAND2_3192 ( P1_U5790 , P1_U4034 , P1_U4147 );
nand NAND2_3193 ( P1_U5791 , P1_IR_REG_22_ , P1_U3952 );
nand NAND2_3194 ( P1_U5792 , P1_IR_REG_31_ , P1_SUB_88_U15 );
not NOT1_3195 ( P1_U5793 , P1_U3451 );
nand NAND2_3196 ( P1_U5794 , P1_IR_REG_19_ , P1_U3952 );
nand NAND2_3197 ( P1_U5795 , P1_IR_REG_31_ , P1_SUB_88_U13 );
not NOT1_3198 ( P1_U5796 , P1_U3452 );
nand NAND2_3199 ( P1_U5797 , P1_IR_REG_20_ , P1_U3952 );
nand NAND2_3200 ( P1_U5798 , P1_IR_REG_31_ , P1_SUB_88_U14 );
not NOT1_3201 ( P1_U5799 , P1_U3453 );
nand NAND2_3202 ( P1_U5800 , P1_IR_REG_21_ , P1_U3952 );
nand NAND2_3203 ( P1_U5801 , P1_IR_REG_31_ , P1_SUB_88_U173 );
not NOT1_3204 ( P1_U5802 , P1_U3450 );
nand NAND2_3205 ( P1_U5803 , P1_IR_REG_30_ , P1_U3952 );
nand NAND2_3206 ( P1_U5804 , P1_IR_REG_31_ , P1_SUB_88_U165 );
not NOT1_3207 ( P1_U5805 , P1_U3447 );
nand NAND2_3208 ( P1_U5806 , P1_IR_REG_29_ , P1_U3952 );
nand NAND2_3209 ( P1_U5807 , P1_IR_REG_31_ , P1_SUB_88_U20 );
not NOT1_3210 ( P1_U5808 , P1_U3448 );
nand NAND2_3211 ( P1_U5809 , P1_IR_REG_28_ , P1_U3952 );
nand NAND2_3212 ( P1_U5810 , P1_IR_REG_31_ , P1_SUB_88_U19 );
not NOT1_3213 ( P1_U5811 , P1_U3449 );
nand NAND2_3214 ( P1_U5812 , P1_IR_REG_0_ , P1_U3952 );
nand NAND2_3215 ( P1_U5813 , P1_IR_REG_31_ , P1_IR_REG_0_ );
not NOT1_3216 ( P1_U5814 , P1_U3454 );
nand NAND2_3217 ( P1_U5815 , P1_IR_REG_27_ , P1_U3952 );
nand NAND2_3218 ( P1_U5816 , P1_IR_REG_31_ , P1_SUB_88_U42 );
not NOT1_3219 ( P1_U5817 , P1_U3455 );
nand NAND2_3220 ( P1_U5818 , U125 , P1_U3954 );
nand NAND2_3221 ( P1_U5819 , P1_U4014 , P1_U3454 );
not NOT1_3222 ( P1_U5820 , P1_U3456 );
nand NAND2_3223 ( P1_U5821 , P1_U3451 , P1_U5802 );
nand NAND2_3224 ( P1_U5822 , P1_U5793 , P1_U4178 );
nand NAND2_3225 ( P1_U5823 , P1_D_REG_1_ , P1_U4144 );
nand NAND2_3226 ( P1_U5824 , P1_U4147 , P1_U3360 );
not NOT1_3227 ( P1_U5825 , P1_U3458 );
nand NAND2_3228 ( P1_U5826 , P1_U5771 , P1_U3360 );
nand NAND2_3229 ( P1_U5827 , P1_D_REG_0_ , P1_U4144 );
not NOT1_3230 ( P1_U5828 , P1_U3457 );
nand NAND2_3231 ( P1_U5829 , P1_REG0_REG_0_ , P1_U3955 );
nand NAND2_3232 ( P1_U5830 , P1_U4033 , P1_U4198 );
nand NAND2_3233 ( P1_U5831 , P1_IR_REG_1_ , P1_U3952 );
nand NAND2_3234 ( P1_U5832 , P1_IR_REG_31_ , P1_SUB_88_U40 );
nand NAND2_3235 ( P1_U5833 , U114 , P1_U3954 );
nand NAND2_3236 ( P1_U5834 , P1_U3460 , P1_U4014 );
not NOT1_3237 ( P1_U5835 , P1_U3461 );
nand NAND2_3238 ( P1_U5836 , P1_REG0_REG_1_ , P1_U3955 );
nand NAND2_3239 ( P1_U5837 , P1_U4033 , P1_U4222 );
nand NAND2_3240 ( P1_U5838 , P1_IR_REG_2_ , P1_U3952 );
nand NAND2_3241 ( P1_U5839 , P1_IR_REG_31_ , P1_SUB_88_U21 );
nand NAND2_3242 ( P1_U5840 , U103 , P1_U3954 );
nand NAND2_3243 ( P1_U5841 , P1_U3463 , P1_U4014 );
not NOT1_3244 ( P1_U5842 , P1_U3464 );
nand NAND2_3245 ( P1_U5843 , P1_REG0_REG_2_ , P1_U3955 );
nand NAND2_3246 ( P1_U5844 , P1_U4033 , P1_U4241 );
nand NAND2_3247 ( P1_U5845 , P1_IR_REG_3_ , P1_U3952 );
nand NAND2_3248 ( P1_U5846 , P1_IR_REG_31_ , P1_SUB_88_U22 );
nand NAND2_3249 ( P1_U5847 , U100 , P1_U3954 );
nand NAND2_3250 ( P1_U5848 , P1_U3466 , P1_U4014 );
not NOT1_3251 ( P1_U5849 , P1_U3467 );
nand NAND2_3252 ( P1_U5850 , P1_REG0_REG_3_ , P1_U3955 );
nand NAND2_3253 ( P1_U5851 , P1_U4033 , P1_U4260 );
nand NAND2_3254 ( P1_U5852 , P1_IR_REG_4_ , P1_U3952 );
nand NAND2_3255 ( P1_U5853 , P1_IR_REG_31_ , P1_SUB_88_U23 );
nand NAND2_3256 ( P1_U5854 , U99 , P1_U3954 );
nand NAND2_3257 ( P1_U5855 , P1_U3469 , P1_U4014 );
not NOT1_3258 ( P1_U5856 , P1_U3470 );
nand NAND2_3259 ( P1_U5857 , P1_REG0_REG_4_ , P1_U3955 );
nand NAND2_3260 ( P1_U5858 , P1_U4033 , P1_U4279 );
nand NAND2_3261 ( P1_U5859 , P1_IR_REG_5_ , P1_U3952 );
nand NAND2_3262 ( P1_U5860 , P1_IR_REG_31_ , P1_SUB_88_U162 );
nand NAND2_3263 ( P1_U5861 , U98 , P1_U3954 );
nand NAND2_3264 ( P1_U5862 , P1_U3472 , P1_U4014 );
not NOT1_3265 ( P1_U5863 , P1_U3473 );
nand NAND2_3266 ( P1_U5864 , P1_REG0_REG_5_ , P1_U3955 );
nand NAND2_3267 ( P1_U5865 , P1_U4033 , P1_U4298 );
nand NAND2_3268 ( P1_U5866 , P1_IR_REG_6_ , P1_U3952 );
nand NAND2_3269 ( P1_U5867 , P1_IR_REG_31_ , P1_SUB_88_U24 );
nand NAND2_3270 ( P1_U5868 , U97 , P1_U3954 );
nand NAND2_3271 ( P1_U5869 , P1_U3475 , P1_U4014 );
not NOT1_3272 ( P1_U5870 , P1_U3476 );
nand NAND2_3273 ( P1_U5871 , P1_REG0_REG_6_ , P1_U3955 );
nand NAND2_3274 ( P1_U5872 , P1_U4033 , P1_U4317 );
nand NAND2_3275 ( P1_U5873 , P1_IR_REG_7_ , P1_U3952 );
nand NAND2_3276 ( P1_U5874 , P1_IR_REG_31_ , P1_SUB_88_U25 );
nand NAND2_3277 ( P1_U5875 , U96 , P1_U3954 );
nand NAND2_3278 ( P1_U5876 , P1_U3478 , P1_U4014 );
not NOT1_3279 ( P1_U5877 , P1_U3479 );
nand NAND2_3280 ( P1_U5878 , P1_REG0_REG_7_ , P1_U3955 );
nand NAND2_3281 ( P1_U5879 , P1_U4033 , P1_U4336 );
nand NAND2_3282 ( P1_U5880 , P1_IR_REG_8_ , P1_U3952 );
nand NAND2_3283 ( P1_U5881 , P1_IR_REG_31_ , P1_SUB_88_U26 );
nand NAND2_3284 ( P1_U5882 , U95 , P1_U3954 );
nand NAND2_3285 ( P1_U5883 , P1_U3481 , P1_U4014 );
not NOT1_3286 ( P1_U5884 , P1_U3482 );
nand NAND2_3287 ( P1_U5885 , P1_REG0_REG_8_ , P1_U3955 );
nand NAND2_3288 ( P1_U5886 , P1_U4033 , P1_U4355 );
nand NAND2_3289 ( P1_U5887 , P1_IR_REG_9_ , P1_U3952 );
nand NAND2_3290 ( P1_U5888 , P1_IR_REG_31_ , P1_SUB_88_U160 );
nand NAND2_3291 ( P1_U5889 , U94 , P1_U3954 );
nand NAND2_3292 ( P1_U5890 , P1_U3484 , P1_U4014 );
not NOT1_3293 ( P1_U5891 , P1_U3485 );
nand NAND2_3294 ( P1_U5892 , P1_REG0_REG_9_ , P1_U3955 );
nand NAND2_3295 ( P1_U5893 , P1_U4033 , P1_U4374 );
nand NAND2_3296 ( P1_U5894 , P1_IR_REG_10_ , P1_U3952 );
nand NAND2_3297 ( P1_U5895 , P1_IR_REG_31_ , P1_SUB_88_U6 );
nand NAND2_3298 ( P1_U5896 , U124 , P1_U3954 );
nand NAND2_3299 ( P1_U5897 , P1_U3487 , P1_U4014 );
not NOT1_3300 ( P1_U5898 , P1_U3488 );
nand NAND2_3301 ( P1_U5899 , P1_REG0_REG_10_ , P1_U3955 );
nand NAND2_3302 ( P1_U5900 , P1_U4033 , P1_U4393 );
nand NAND2_3303 ( P1_U5901 , P1_IR_REG_11_ , P1_U3952 );
nand NAND2_3304 ( P1_U5902 , P1_IR_REG_31_ , P1_SUB_88_U7 );
nand NAND2_3305 ( P1_U5903 , U123 , P1_U3954 );
nand NAND2_3306 ( P1_U5904 , P1_U3490 , P1_U4014 );
not NOT1_3307 ( P1_U5905 , P1_U3491 );
nand NAND2_3308 ( P1_U5906 , P1_REG0_REG_11_ , P1_U3955 );
nand NAND2_3309 ( P1_U5907 , P1_U4033 , P1_U4412 );
nand NAND2_3310 ( P1_U5908 , P1_IR_REG_12_ , P1_U3952 );
nand NAND2_3311 ( P1_U5909 , P1_IR_REG_31_ , P1_SUB_88_U8 );
nand NAND2_3312 ( P1_U5910 , U122 , P1_U3954 );
nand NAND2_3313 ( P1_U5911 , P1_U3493 , P1_U4014 );
not NOT1_3314 ( P1_U5912 , P1_U3494 );
nand NAND2_3315 ( P1_U5913 , P1_REG0_REG_12_ , P1_U3955 );
nand NAND2_3316 ( P1_U5914 , P1_U4033 , P1_U4431 );
nand NAND2_3317 ( P1_U5915 , P1_IR_REG_13_ , P1_U3952 );
nand NAND2_3318 ( P1_U5916 , P1_IR_REG_31_ , P1_SUB_88_U179 );
nand NAND2_3319 ( P1_U5917 , U121 , P1_U3954 );
nand NAND2_3320 ( P1_U5918 , P1_U3496 , P1_U4014 );
not NOT1_3321 ( P1_U5919 , P1_U3497 );
nand NAND2_3322 ( P1_U5920 , P1_REG0_REG_13_ , P1_U3955 );
nand NAND2_3323 ( P1_U5921 , P1_U4033 , P1_U4450 );
nand NAND2_3324 ( P1_U5922 , P1_IR_REG_14_ , P1_U3952 );
nand NAND2_3325 ( P1_U5923 , P1_IR_REG_31_ , P1_SUB_88_U9 );
nand NAND2_3326 ( P1_U5924 , U120 , P1_U3954 );
nand NAND2_3327 ( P1_U5925 , P1_U3499 , P1_U4014 );
not NOT1_3328 ( P1_U5926 , P1_U3500 );
nand NAND2_3329 ( P1_U5927 , P1_REG0_REG_14_ , P1_U3955 );
nand NAND2_3330 ( P1_U5928 , P1_U4033 , P1_U4469 );
nand NAND2_3331 ( P1_U5929 , P1_IR_REG_15_ , P1_U3952 );
nand NAND2_3332 ( P1_U5930 , P1_IR_REG_31_ , P1_SUB_88_U10 );
nand NAND2_3333 ( P1_U5931 , U119 , P1_U3954 );
nand NAND2_3334 ( P1_U5932 , P1_U3502 , P1_U4014 );
not NOT1_3335 ( P1_U5933 , P1_U3503 );
nand NAND2_3336 ( P1_U5934 , P1_REG0_REG_15_ , P1_U3955 );
nand NAND2_3337 ( P1_U5935 , P1_U4033 , P1_U4488 );
nand NAND2_3338 ( P1_U5936 , P1_IR_REG_16_ , P1_U3952 );
nand NAND2_3339 ( P1_U5937 , P1_IR_REG_31_ , P1_SUB_88_U11 );
nand NAND2_3340 ( P1_U5938 , U118 , P1_U3954 );
nand NAND2_3341 ( P1_U5939 , P1_U3505 , P1_U4014 );
not NOT1_3342 ( P1_U5940 , P1_U3506 );
nand NAND2_3343 ( P1_U5941 , P1_REG0_REG_16_ , P1_U3955 );
nand NAND2_3344 ( P1_U5942 , P1_U4033 , P1_U4507 );
nand NAND2_3345 ( P1_U5943 , P1_IR_REG_17_ , P1_U3952 );
nand NAND2_3346 ( P1_U5944 , P1_IR_REG_31_ , P1_SUB_88_U177 );
nand NAND2_3347 ( P1_U5945 , U117 , P1_U3954 );
nand NAND2_3348 ( P1_U5946 , P1_U3508 , P1_U4014 );
not NOT1_3349 ( P1_U5947 , P1_U3509 );
nand NAND2_3350 ( P1_U5948 , P1_REG0_REG_17_ , P1_U3955 );
nand NAND2_3351 ( P1_U5949 , P1_U4033 , P1_U4526 );
nand NAND2_3352 ( P1_U5950 , P1_IR_REG_18_ , P1_U3952 );
nand NAND2_3353 ( P1_U5951 , P1_IR_REG_31_ , P1_SUB_88_U12 );
nand NAND2_3354 ( P1_U5952 , U116 , P1_U3954 );
nand NAND2_3355 ( P1_U5953 , P1_U3511 , P1_U4014 );
not NOT1_3356 ( P1_U5954 , P1_U3512 );
nand NAND2_3357 ( P1_U5955 , P1_REG0_REG_18_ , P1_U3955 );
nand NAND2_3358 ( P1_U5956 , P1_U4033 , P1_U4545 );
nand NAND2_3359 ( P1_U5957 , U115 , P1_U3954 );
nand NAND2_3360 ( P1_U5958 , P1_U4014 , P1_U3452 );
not NOT1_3361 ( P1_U5959 , P1_U3514 );
nand NAND2_3362 ( P1_U5960 , P1_REG0_REG_19_ , P1_U3955 );
nand NAND2_3363 ( P1_U5961 , P1_U4033 , P1_U4564 );
nand NAND2_3364 ( P1_U5962 , P1_REG0_REG_20_ , P1_U3955 );
nand NAND2_3365 ( P1_U5963 , P1_U4033 , P1_U4583 );
nand NAND2_3366 ( P1_U5964 , P1_REG0_REG_21_ , P1_U3955 );
nand NAND2_3367 ( P1_U5965 , P1_U4033 , P1_U4602 );
nand NAND2_3368 ( P1_U5966 , P1_REG0_REG_22_ , P1_U3955 );
nand NAND2_3369 ( P1_U5967 , P1_U4033 , P1_U4621 );
nand NAND2_3370 ( P1_U5968 , P1_REG0_REG_23_ , P1_U3955 );
nand NAND2_3371 ( P1_U5969 , P1_U4033 , P1_U4640 );
nand NAND2_3372 ( P1_U5970 , P1_REG0_REG_24_ , P1_U3955 );
nand NAND2_3373 ( P1_U5971 , P1_U4033 , P1_U4659 );
nand NAND2_3374 ( P1_U5972 , P1_REG0_REG_25_ , P1_U3955 );
nand NAND2_3375 ( P1_U5973 , P1_U4033 , P1_U4678 );
nand NAND2_3376 ( P1_U5974 , P1_REG0_REG_26_ , P1_U3955 );
nand NAND2_3377 ( P1_U5975 , P1_U4033 , P1_U4697 );
nand NAND2_3378 ( P1_U5976 , P1_REG0_REG_27_ , P1_U3955 );
nand NAND2_3379 ( P1_U5977 , P1_U4033 , P1_U4716 );
nand NAND2_3380 ( P1_U5978 , P1_REG0_REG_28_ , P1_U3955 );
nand NAND2_3381 ( P1_U5979 , P1_U4033 , P1_U4735 );
nand NAND2_3382 ( P1_U5980 , P1_REG0_REG_29_ , P1_U3955 );
nand NAND2_3383 ( P1_U5981 , P1_U4033 , P1_U4755 );
nand NAND2_3384 ( P1_U5982 , P1_REG0_REG_30_ , P1_U3955 );
nand NAND2_3385 ( P1_U5983 , P1_U4033 , P1_U4762 );
nand NAND2_3386 ( P1_U5984 , P1_REG0_REG_31_ , P1_U3955 );
nand NAND2_3387 ( P1_U5985 , P1_U4033 , P1_U4765 );
nand NAND2_3388 ( P1_U5986 , P1_REG1_REG_0_ , P1_U3956 );
nand NAND2_3389 ( P1_U5987 , P1_U4032 , P1_U4198 );
nand NAND2_3390 ( P1_U5988 , P1_REG1_REG_1_ , P1_U3956 );
nand NAND2_3391 ( P1_U5989 , P1_U4032 , P1_U4222 );
nand NAND2_3392 ( P1_U5990 , P1_REG1_REG_2_ , P1_U3956 );
nand NAND2_3393 ( P1_U5991 , P1_U4032 , P1_U4241 );
nand NAND2_3394 ( P1_U5992 , P1_REG1_REG_3_ , P1_U3956 );
nand NAND2_3395 ( P1_U5993 , P1_U4032 , P1_U4260 );
nand NAND2_3396 ( P1_U5994 , P1_REG1_REG_4_ , P1_U3956 );
nand NAND2_3397 ( P1_U5995 , P1_U4032 , P1_U4279 );
nand NAND2_3398 ( P1_U5996 , P1_REG1_REG_5_ , P1_U3956 );
nand NAND2_3399 ( P1_U5997 , P1_U4032 , P1_U4298 );
nand NAND2_3400 ( P1_U5998 , P1_REG1_REG_6_ , P1_U3956 );
nand NAND2_3401 ( P1_U5999 , P1_U4032 , P1_U4317 );
nand NAND2_3402 ( P1_U6000 , P1_REG1_REG_7_ , P1_U3956 );
nand NAND2_3403 ( P1_U6001 , P1_U4032 , P1_U4336 );
nand NAND2_3404 ( P1_U6002 , P1_REG1_REG_8_ , P1_U3956 );
nand NAND2_3405 ( P1_U6003 , P1_U4032 , P1_U4355 );
nand NAND2_3406 ( P1_U6004 , P1_REG1_REG_9_ , P1_U3956 );
nand NAND2_3407 ( P1_U6005 , P1_U4032 , P1_U4374 );
nand NAND2_3408 ( P1_U6006 , P1_REG1_REG_10_ , P1_U3956 );
nand NAND2_3409 ( P1_U6007 , P1_U4032 , P1_U4393 );
nand NAND2_3410 ( P1_U6008 , P1_REG1_REG_11_ , P1_U3956 );
nand NAND2_3411 ( P1_U6009 , P1_U4032 , P1_U4412 );
nand NAND2_3412 ( P1_U6010 , P1_REG1_REG_12_ , P1_U3956 );
nand NAND2_3413 ( P1_U6011 , P1_U4032 , P1_U4431 );
nand NAND2_3414 ( P1_U6012 , P1_REG1_REG_13_ , P1_U3956 );
nand NAND2_3415 ( P1_U6013 , P1_U4032 , P1_U4450 );
nand NAND2_3416 ( P1_U6014 , P1_REG1_REG_14_ , P1_U3956 );
nand NAND2_3417 ( P1_U6015 , P1_U4032 , P1_U4469 );
nand NAND2_3418 ( P1_U6016 , P1_REG1_REG_15_ , P1_U3956 );
nand NAND2_3419 ( P1_U6017 , P1_U4032 , P1_U4488 );
nand NAND2_3420 ( P1_U6018 , P1_REG1_REG_16_ , P1_U3956 );
nand NAND2_3421 ( P1_U6019 , P1_U4032 , P1_U4507 );
nand NAND2_3422 ( P1_U6020 , P1_REG1_REG_17_ , P1_U3956 );
nand NAND2_3423 ( P1_U6021 , P1_U4032 , P1_U4526 );
nand NAND2_3424 ( P1_U6022 , P1_REG1_REG_18_ , P1_U3956 );
nand NAND2_3425 ( P1_U6023 , P1_U4032 , P1_U4545 );
nand NAND2_3426 ( P1_U6024 , P1_REG1_REG_19_ , P1_U3956 );
nand NAND2_3427 ( P1_U6025 , P1_U4032 , P1_U4564 );
nand NAND2_3428 ( P1_U6026 , P1_REG1_REG_20_ , P1_U3956 );
nand NAND2_3429 ( P1_U6027 , P1_U4032 , P1_U4583 );
nand NAND2_3430 ( P1_U6028 , P1_REG1_REG_21_ , P1_U3956 );
nand NAND2_3431 ( P1_U6029 , P1_U4032 , P1_U4602 );
nand NAND2_3432 ( P1_U6030 , P1_REG1_REG_22_ , P1_U3956 );
nand NAND2_3433 ( P1_U6031 , P1_U4032 , P1_U4621 );
nand NAND2_3434 ( P1_U6032 , P1_REG1_REG_23_ , P1_U3956 );
nand NAND2_3435 ( P1_U6033 , P1_U4032 , P1_U4640 );
nand NAND2_3436 ( P1_U6034 , P1_REG1_REG_24_ , P1_U3956 );
nand NAND2_3437 ( P1_U6035 , P1_U4032 , P1_U4659 );
nand NAND2_3438 ( P1_U6036 , P1_REG1_REG_25_ , P1_U3956 );
nand NAND2_3439 ( P1_U6037 , P1_U4032 , P1_U4678 );
nand NAND2_3440 ( P1_U6038 , P1_REG1_REG_26_ , P1_U3956 );
nand NAND2_3441 ( P1_U6039 , P1_U4032 , P1_U4697 );
nand NAND2_3442 ( P1_U6040 , P1_REG1_REG_27_ , P1_U3956 );
nand NAND2_3443 ( P1_U6041 , P1_U4032 , P1_U4716 );
nand NAND2_3444 ( P1_U6042 , P1_REG1_REG_28_ , P1_U3956 );
nand NAND2_3445 ( P1_U6043 , P1_U4032 , P1_U4735 );
nand NAND2_3446 ( P1_U6044 , P1_REG1_REG_29_ , P1_U3956 );
nand NAND2_3447 ( P1_U6045 , P1_U4032 , P1_U4755 );
nand NAND2_3448 ( P1_U6046 , P1_REG1_REG_30_ , P1_U3956 );
nand NAND2_3449 ( P1_U6047 , P1_U4032 , P1_U4762 );
nand NAND2_3450 ( P1_U6048 , P1_REG1_REG_31_ , P1_U3956 );
nand NAND2_3451 ( P1_U6049 , P1_U4032 , P1_U4765 );
nand NAND2_3452 ( P1_U6050 , P1_REG2_REG_0_ , P1_U3420 );
nand NAND2_3453 ( P1_U6051 , P1_U4031 , P1_U3376 );
nand NAND2_3454 ( P1_U6052 , P1_REG2_REG_1_ , P1_U3420 );
nand NAND2_3455 ( P1_U6053 , P1_U4031 , P1_U3378 );
nand NAND2_3456 ( P1_U6054 , P1_REG2_REG_2_ , P1_U3420 );
nand NAND2_3457 ( P1_U6055 , P1_U4031 , P1_U3379 );
nand NAND2_3458 ( P1_U6056 , P1_REG2_REG_3_ , P1_U3420 );
nand NAND2_3459 ( P1_U6057 , P1_U4031 , P1_U3380 );
nand NAND2_3460 ( P1_U6058 , P1_REG2_REG_4_ , P1_U3420 );
nand NAND2_3461 ( P1_U6059 , P1_U4031 , P1_U3381 );
nand NAND2_3462 ( P1_U6060 , P1_REG2_REG_5_ , P1_U3420 );
nand NAND2_3463 ( P1_U6061 , P1_U4031 , P1_U3382 );
nand NAND2_3464 ( P1_U6062 , P1_REG2_REG_6_ , P1_U3420 );
nand NAND2_3465 ( P1_U6063 , P1_U4031 , P1_U3383 );
nand NAND2_3466 ( P1_U6064 , P1_REG2_REG_7_ , P1_U3420 );
nand NAND2_3467 ( P1_U6065 , P1_U4031 , P1_U3384 );
nand NAND2_3468 ( P1_U6066 , P1_REG2_REG_8_ , P1_U3420 );
nand NAND2_3469 ( P1_U6067 , P1_U4031 , P1_U3385 );
nand NAND2_3470 ( P1_U6068 , P1_REG2_REG_9_ , P1_U3420 );
nand NAND2_3471 ( P1_U6069 , P1_U4031 , P1_U3386 );
nand NAND2_3472 ( P1_U6070 , P1_REG2_REG_10_ , P1_U3420 );
nand NAND2_3473 ( P1_U6071 , P1_U4031 , P1_U3387 );
nand NAND2_3474 ( P1_U6072 , P1_REG2_REG_11_ , P1_U3420 );
nand NAND2_3475 ( P1_U6073 , P1_U4031 , P1_U3388 );
nand NAND2_3476 ( P1_U6074 , P1_REG2_REG_12_ , P1_U3420 );
nand NAND2_3477 ( P1_U6075 , P1_U4031 , P1_U3389 );
nand NAND2_3478 ( P1_U6076 , P1_REG2_REG_13_ , P1_U3420 );
nand NAND2_3479 ( P1_U6077 , P1_U4031 , P1_U3390 );
nand NAND2_3480 ( P1_U6078 , P1_REG2_REG_14_ , P1_U3420 );
nand NAND2_3481 ( P1_U6079 , P1_U4031 , P1_U3391 );
nand NAND2_3482 ( P1_U6080 , P1_REG2_REG_15_ , P1_U3420 );
nand NAND2_3483 ( P1_U6081 , P1_U4031 , P1_U3392 );
nand NAND2_3484 ( P1_U6082 , P1_REG2_REG_16_ , P1_U3420 );
nand NAND2_3485 ( P1_U6083 , P1_U4031 , P1_U3393 );
nand NAND2_3486 ( P1_U6084 , P1_REG2_REG_17_ , P1_U3420 );
nand NAND2_3487 ( P1_U6085 , P1_U4031 , P1_U3394 );
nand NAND2_3488 ( P1_U6086 , P1_REG2_REG_18_ , P1_U3420 );
nand NAND2_3489 ( P1_U6087 , P1_U4031 , P1_U3395 );
nand NAND2_3490 ( P1_U6088 , P1_REG2_REG_19_ , P1_U3420 );
nand NAND2_3491 ( P1_U6089 , P1_U4031 , P1_U3396 );
nand NAND2_3492 ( P1_U6090 , P1_REG2_REG_20_ , P1_U3420 );
nand NAND2_3493 ( P1_U6091 , P1_U4031 , P1_U3398 );
nand NAND2_3494 ( P1_U6092 , P1_REG2_REG_21_ , P1_U3420 );
nand NAND2_3495 ( P1_U6093 , P1_U4031 , P1_U3400 );
nand NAND2_3496 ( P1_U6094 , P1_REG2_REG_22_ , P1_U3420 );
nand NAND2_3497 ( P1_U6095 , P1_U4031 , P1_U3402 );
nand NAND2_3498 ( P1_U6096 , P1_REG2_REG_23_ , P1_U3420 );
nand NAND2_3499 ( P1_U6097 , P1_U4031 , P1_U3404 );
nand NAND2_3500 ( P1_U6098 , P1_REG2_REG_24_ , P1_U3420 );
nand NAND2_3501 ( P1_U6099 , P1_U4031 , P1_U3406 );
nand NAND2_3502 ( P1_U6100 , P1_REG2_REG_25_ , P1_U3420 );
nand NAND2_3503 ( P1_U6101 , P1_U4031 , P1_U3408 );
nand NAND2_3504 ( P1_U6102 , P1_REG2_REG_26_ , P1_U3420 );
nand NAND2_3505 ( P1_U6103 , P1_U4031 , P1_U3410 );
nand NAND2_3506 ( P1_U6104 , P1_REG2_REG_27_ , P1_U3420 );
nand NAND2_3507 ( P1_U6105 , P1_U4031 , P1_U3412 );
nand NAND2_3508 ( P1_U6106 , P1_REG2_REG_28_ , P1_U3420 );
nand NAND2_3509 ( P1_U6107 , P1_U4031 , P1_U3414 );
nand NAND2_3510 ( P1_U6108 , P1_REG2_REG_29_ , P1_U3420 );
nand NAND2_3511 ( P1_U6109 , P1_U4031 , P1_U3416 );
nand NAND2_3512 ( P1_U6110 , P1_REG2_REG_30_ , P1_U3420 );
nand NAND2_3513 ( P1_U6111 , P1_U4035 , P1_U4031 );
nand NAND2_3514 ( P1_U6112 , P1_REG2_REG_31_ , P1_U3420 );
nand NAND2_3515 ( P1_U6113 , P1_U4035 , P1_U4031 );
nand NAND2_3516 ( P1_U6114 , P1_DATAO_REG_0_ , P1_U3430 );
nand NAND2_3517 ( P1_U6115 , P1_U4016 , P1_U3077 );
nand NAND2_3518 ( P1_U6116 , P1_DATAO_REG_1_ , P1_U3430 );
nand NAND2_3519 ( P1_U6117 , P1_U4016 , P1_U3078 );
nand NAND2_3520 ( P1_U6118 , P1_DATAO_REG_2_ , P1_U3430 );
nand NAND2_3521 ( P1_U6119 , P1_U4016 , P1_U3068 );
nand NAND2_3522 ( P1_U6120 , P1_DATAO_REG_3_ , P1_U3430 );
nand NAND2_3523 ( P1_U6121 , P1_U4016 , P1_U3064 );
nand NAND2_3524 ( P1_U6122 , P1_DATAO_REG_4_ , P1_U3430 );
nand NAND2_3525 ( P1_U6123 , P1_U4016 , P1_U3060 );
nand NAND2_3526 ( P1_U6124 , P1_DATAO_REG_5_ , P1_U3430 );
nand NAND2_3527 ( P1_U6125 , P1_U4016 , P1_U3067 );
nand NAND2_3528 ( P1_U6126 , P1_DATAO_REG_6_ , P1_U3430 );
nand NAND2_3529 ( P1_U6127 , P1_U4016 , P1_U3071 );
nand NAND2_3530 ( P1_U6128 , P1_DATAO_REG_7_ , P1_U3430 );
nand NAND2_3531 ( P1_U6129 , P1_U4016 , P1_U3070 );
nand NAND2_3532 ( P1_U6130 , P1_DATAO_REG_8_ , P1_U3430 );
nand NAND2_3533 ( P1_U6131 , P1_U4016 , P1_U3084 );
nand NAND2_3534 ( P1_U6132 , P1_DATAO_REG_9_ , P1_U3430 );
nand NAND2_3535 ( P1_U6133 , P1_U4016 , P1_U3083 );
nand NAND2_3536 ( P1_U6134 , P1_DATAO_REG_10_ , P1_U3430 );
nand NAND2_3537 ( P1_U6135 , P1_U4016 , P1_U3062 );
nand NAND2_3538 ( P1_U6136 , P1_DATAO_REG_11_ , P1_U3430 );
nand NAND2_3539 ( P1_U6137 , P1_U4016 , P1_U3063 );
nand NAND2_3540 ( P1_U6138 , P1_DATAO_REG_12_ , P1_U3430 );
nand NAND2_3541 ( P1_U6139 , P1_U4016 , P1_U3072 );
nand NAND2_3542 ( P1_U6140 , P1_DATAO_REG_13_ , P1_U3430 );
nand NAND2_3543 ( P1_U6141 , P1_U4016 , P1_U3080 );
nand NAND2_3544 ( P1_U6142 , P1_DATAO_REG_14_ , P1_U3430 );
nand NAND2_3545 ( P1_U6143 , P1_U4016 , P1_U3079 );
nand NAND2_3546 ( P1_U6144 , P1_DATAO_REG_15_ , P1_U3430 );
nand NAND2_3547 ( P1_U6145 , P1_U4016 , P1_U3074 );
nand NAND2_3548 ( P1_U6146 , P1_DATAO_REG_16_ , P1_U3430 );
nand NAND2_3549 ( P1_U6147 , P1_U4016 , P1_U3073 );
nand NAND2_3550 ( P1_U6148 , P1_DATAO_REG_17_ , P1_U3430 );
nand NAND2_3551 ( P1_U6149 , P1_U4016 , P1_U3069 );
nand NAND2_3552 ( P1_U6150 , P1_DATAO_REG_18_ , P1_U3430 );
nand NAND2_3553 ( P1_U6151 , P1_U4016 , P1_U3082 );
nand NAND2_3554 ( P1_U6152 , P1_DATAO_REG_19_ , P1_U3430 );
nand NAND2_3555 ( P1_U6153 , P1_U4016 , P1_U3081 );
nand NAND2_3556 ( P1_U6154 , P1_DATAO_REG_20_ , P1_U3430 );
nand NAND2_3557 ( P1_U6155 , P1_U4016 , P1_U3076 );
nand NAND2_3558 ( P1_U6156 , P1_DATAO_REG_21_ , P1_U3430 );
nand NAND2_3559 ( P1_U6157 , P1_U4016 , P1_U3075 );
nand NAND2_3560 ( P1_U6158 , P1_DATAO_REG_22_ , P1_U3430 );
nand NAND2_3561 ( P1_U6159 , P1_U4016 , P1_U3061 );
nand NAND2_3562 ( P1_U6160 , P1_DATAO_REG_23_ , P1_U3430 );
nand NAND2_3563 ( P1_U6161 , P1_U4016 , P1_U3066 );
nand NAND2_3564 ( P1_U6162 , P1_DATAO_REG_24_ , P1_U3430 );
nand NAND2_3565 ( P1_U6163 , P1_U4016 , P1_U3065 );
nand NAND2_3566 ( P1_U6164 , P1_DATAO_REG_25_ , P1_U3430 );
nand NAND2_3567 ( P1_U6165 , P1_U4016 , P1_U3058 );
nand NAND2_3568 ( P1_U6166 , P1_DATAO_REG_26_ , P1_U3430 );
nand NAND2_3569 ( P1_U6167 , P1_U4016 , P1_U3057 );
nand NAND2_3570 ( P1_U6168 , P1_DATAO_REG_27_ , P1_U3430 );
nand NAND2_3571 ( P1_U6169 , P1_U4016 , P1_U3053 );
nand NAND2_3572 ( P1_U6170 , P1_DATAO_REG_28_ , P1_U3430 );
nand NAND2_3573 ( P1_U6171 , P1_U4016 , P1_U3054 );
nand NAND2_3574 ( P1_U6172 , P1_DATAO_REG_29_ , P1_U3430 );
nand NAND2_3575 ( P1_U6173 , P1_U4016 , P1_U3055 );
nand NAND2_3576 ( P1_U6174 , P1_DATAO_REG_30_ , P1_U3430 );
nand NAND2_3577 ( P1_U6175 , P1_U4016 , P1_U3059 );
nand NAND2_3578 ( P1_U6176 , P1_DATAO_REG_31_ , P1_U3430 );
nand NAND2_3579 ( P1_U6177 , P1_U4016 , P1_U3056 );
nand NAND3_3580 ( P1_U6178 , P1_U3450 , P1_U5793 , P1_U3432 );
nand NAND2_3581 ( P1_U6179 , P1_R1375_U9 , P1_U4030 );
nand NAND2_3582 ( P1_U6180 , P1_U4017 , P1_U3054 );
nand NAND2_3583 ( P1_U6181 , P1_U3413 , P1_U4702 );
nand NAND2_3584 ( P1_U6182 , P1_U6181 , P1_U6180 );
nand NAND2_3585 ( P1_U6183 , P1_U4026 , P1_U3056 );
nand NAND2_3586 ( P1_U6184 , P1_U3418 , P1_U4759 );
nand NAND2_3587 ( P1_U6185 , P1_U6184 , P1_U6183 );
nand NAND2_3588 ( P1_U6186 , P1_U4025 , P1_U3076 );
nand NAND2_3589 ( P1_U6187 , P1_U3397 , P1_U4550 );
nand NAND2_3590 ( P1_U6188 , P1_U6187 , P1_U6186 );
nand NAND2_3591 ( P1_U6189 , P1_U4027 , P1_U3059 );
nand NAND2_3592 ( P1_U6190 , P1_U3417 , P1_U4739 );
nand NAND2_3593 ( P1_U6191 , P1_U6190 , P1_U6189 );
nand NAND2_3594 ( P1_U6192 , P1_U5959 , P1_U4531 );
nand NAND2_3595 ( P1_U6193 , P1_U3514 , P1_U3081 );
nand NAND2_3596 ( P1_U6194 , P1_U6193 , P1_U6192 );
nand NAND2_3597 ( P1_U6195 , P1_U5905 , P1_U4379 );
nand NAND2_3598 ( P1_U6196 , P1_U3491 , P1_U3063 );
nand NAND2_3599 ( P1_U6197 , P1_U6196 , P1_U6195 );
nand NAND2_3600 ( P1_U6198 , P1_U5856 , P1_U4246 );
nand NAND2_3601 ( P1_U6199 , P1_U3470 , P1_U3060 );
nand NAND2_3602 ( P1_U6200 , P1_U6199 , P1_U6198 );
nand NAND2_3603 ( P1_U6201 , P1_U5898 , P1_U4360 );
nand NAND2_3604 ( P1_U6202 , P1_U3488 , P1_U3062 );
nand NAND2_3605 ( P1_U6203 , P1_U6202 , P1_U6201 );
nand NAND2_3606 ( P1_U6204 , P1_U4028 , P1_U3055 );
nand NAND2_3607 ( P1_U6205 , P1_U3415 , P1_U4721 );
nand NAND2_3608 ( P1_U6206 , P1_U6205 , P1_U6204 );
nand NAND2_3609 ( P1_U6207 , P1_U4018 , P1_U3053 );
nand NAND2_3610 ( P1_U6208 , P1_U3411 , P1_U4683 );
nand NAND2_3611 ( P1_U6209 , P1_U6208 , P1_U6207 );
nand NAND2_3612 ( P1_U6210 , P1_U5947 , P1_U4493 );
nand NAND2_3613 ( P1_U6211 , P1_U3509 , P1_U3069 );
nand NAND2_3614 ( P1_U6212 , P1_U6211 , P1_U6210 );
nand NAND2_3615 ( P1_U6213 , P1_U5884 , P1_U4322 );
nand NAND2_3616 ( P1_U6214 , P1_U3482 , P1_U3084 );
nand NAND2_3617 ( P1_U6215 , P1_U6214 , P1_U6213 );
nand NAND2_3618 ( P1_U6216 , P1_U5891 , P1_U4341 );
nand NAND2_3619 ( P1_U6217 , P1_U3485 , P1_U3083 );
nand NAND2_3620 ( P1_U6218 , P1_U6217 , P1_U6216 );
nand NAND2_3621 ( P1_U6219 , P1_U5919 , P1_U4417 );
nand NAND2_3622 ( P1_U6220 , P1_U3497 , P1_U3080 );
nand NAND2_3623 ( P1_U6221 , P1_U6220 , P1_U6219 );
nand NAND2_3624 ( P1_U6222 , P1_U5926 , P1_U4436 );
nand NAND2_3625 ( P1_U6223 , P1_U3500 , P1_U3079 );
nand NAND2_3626 ( P1_U6224 , P1_U6223 , P1_U6222 );
nand NAND2_3627 ( P1_U6225 , P1_U5820 , P1_U4208 );
nand NAND2_3628 ( P1_U6226 , P1_U3456 , P1_U3077 );
nand NAND2_3629 ( P1_U6227 , P1_U6226 , P1_U6225 );
nand NAND2_3630 ( P1_U6228 , P1_U5835 , P1_U4184 );
nand NAND2_3631 ( P1_U6229 , P1_U3461 , P1_U3078 );
nand NAND2_3632 ( P1_U6230 , P1_U6229 , P1_U6228 );
nand NAND2_3633 ( P1_U6231 , P1_U5933 , P1_U4455 );
nand NAND2_3634 ( P1_U6232 , P1_U3503 , P1_U3074 );
nand NAND2_3635 ( P1_U6233 , P1_U6232 , P1_U6231 );
nand NAND2_3636 ( P1_U6234 , P1_U5940 , P1_U4474 );
nand NAND2_3637 ( P1_U6235 , P1_U3506 , P1_U3073 );
nand NAND2_3638 ( P1_U6236 , P1_U6235 , P1_U6234 );
nand NAND2_3639 ( P1_U6237 , P1_U5870 , P1_U4284 );
nand NAND2_3640 ( P1_U6238 , P1_U3476 , P1_U3071 );
nand NAND2_3641 ( P1_U6239 , P1_U6238 , P1_U6237 );
nand NAND2_3642 ( P1_U6240 , P1_U5877 , P1_U4303 );
nand NAND2_3643 ( P1_U6241 , P1_U3479 , P1_U3070 );
nand NAND2_3644 ( P1_U6242 , P1_U6241 , P1_U6240 );
nand NAND2_3645 ( P1_U6243 , P1_U5912 , P1_U4398 );
nand NAND2_3646 ( P1_U6244 , P1_U3494 , P1_U3072 );
nand NAND2_3647 ( P1_U6245 , P1_U6244 , P1_U6243 );
nand NAND2_3648 ( P1_U6246 , P1_U5842 , P1_U4203 );
nand NAND2_3649 ( P1_U6247 , P1_U3464 , P1_U3068 );
nand NAND2_3650 ( P1_U6248 , P1_U6247 , P1_U6246 );
nand NAND2_3651 ( P1_U6249 , P1_U5849 , P1_U4227 );
nand NAND2_3652 ( P1_U6250 , P1_U3467 , P1_U3064 );
nand NAND2_3653 ( P1_U6251 , P1_U6250 , P1_U6249 );
nand NAND2_3654 ( P1_U6252 , P1_U5863 , P1_U4265 );
nand NAND2_3655 ( P1_U6253 , P1_U3473 , P1_U3067 );
nand NAND2_3656 ( P1_U6254 , P1_U6253 , P1_U6252 );
nand NAND2_3657 ( P1_U6255 , P1_U5954 , P1_U4512 );
nand NAND2_3658 ( P1_U6256 , P1_U3512 , P1_U3082 );
nand NAND2_3659 ( P1_U6257 , P1_U6256 , P1_U6255 );
nand NAND2_3660 ( P1_U6258 , P1_U4021 , P1_U3065 );
nand NAND2_3661 ( P1_U6259 , P1_U3405 , P1_U4626 );
nand NAND2_3662 ( P1_U6260 , P1_U6259 , P1_U6258 );
nand NAND2_3663 ( P1_U6261 , P1_U4022 , P1_U3066 );
nand NAND2_3664 ( P1_U6262 , P1_U3403 , P1_U4607 );
nand NAND2_3665 ( P1_U6263 , P1_U6262 , P1_U6261 );
nand NAND2_3666 ( P1_U6264 , P1_U4024 , P1_U3075 );
nand NAND2_3667 ( P1_U6265 , P1_U3399 , P1_U4569 );
nand NAND2_3668 ( P1_U6266 , P1_U6265 , P1_U6264 );
nand NAND2_3669 ( P1_U6267 , P1_U4023 , P1_U3061 );
nand NAND2_3670 ( P1_U6268 , P1_U3401 , P1_U4588 );
nand NAND2_3671 ( P1_U6269 , P1_U6268 , P1_U6267 );
nand NAND2_3672 ( P1_U6270 , P1_U4020 , P1_U3058 );
nand NAND2_3673 ( P1_U6271 , P1_U3407 , P1_U4645 );
nand NAND2_3674 ( P1_U6272 , P1_U6271 , P1_U6270 );
nand NAND2_3675 ( P1_U6273 , P1_U4019 , P1_U3057 );
nand NAND2_3676 ( P1_U6274 , P1_U3409 , P1_U4664 );
nand NAND2_3677 ( P1_U6275 , P1_U6274 , P1_U6273 );
nand NAND2_3678 ( P1_U6276 , P1_U4041 , P1_U3991 );
nand NAND2_3679 ( P1_U6277 , P1_U5129 , P1_U3049 );
nand NAND3_3680 ( P1_U6278 , P1_U5133 , P1_U3432 , P1_U5799 );
nand NAND2_3681 ( P1_U6279 , P1_U3453 , P1_U5130 );
nand NAND2_3682 ( P1_U6280 , P1_U5786 , P1_U3431 );
nand NAND2_3683 ( P1_U6281 , P1_U3451 , P1_U3444 );
nand NAND2_3684 ( P1_U6282 , P1_U3450 , P1_U5144 );
nand NAND2_3685 ( P1_U6283 , P1_U5802 , P1_U3994 );
nand NAND2_3686 ( P1_U6284 , P1_U3454 , P1_U5408 );
nand NAND3_3687 ( P1_U6285 , P1_U3015 , P1_REG2_REG_0_ , P1_U5814 );
nand NAND2_3688 ( P3_R1161_U489 , P3_U3079 , P3_R1161_U69 );
nand NAND2_3689 ( P3_R1161_U488 , P3_R1161_U254 , P3_R1161_U486 );
nand NAND2_3690 ( P3_R1161_U487 , P3_R1161_U165 , P3_R1161_U166 );
nand NAND2_3691 ( P3_R1161_U486 , P3_R1161_U485 , P3_R1161_U484 );
nand NAND2_3692 ( P3_R1161_U485 , P3_U3431 , P3_R1161_U72 );
nand NAND2_3693 ( P3_R1161_U484 , P3_U3078 , P3_R1161_U71 );
nand NAND2_3694 ( P3_R1161_U483 , P3_U3431 , P3_R1161_U72 );
nand NAND2_3695 ( P3_R1161_U482 , P3_U3078 , P3_R1161_U71 );
nand NAND2_3696 ( P3_R1161_U481 , P3_R1161_U258 , P3_R1161_U479 );
nand NAND2_3697 ( P3_R1161_U480 , P3_R1161_U163 , P3_R1161_U164 );
nand NAND2_3698 ( P3_R1161_U479 , P3_R1161_U478 , P3_R1161_U477 );
nand NAND2_3699 ( P3_R1161_U478 , P3_U3434 , P3_R1161_U74 );
nand NAND2_3700 ( P3_R1161_U477 , P3_U3073 , P3_R1161_U73 );
nand NAND2_3701 ( P3_R1161_U476 , P3_U3434 , P3_R1161_U74 );
nand NAND2_3702 ( P3_R1161_U475 , P3_U3073 , P3_R1161_U73 );
nand NAND2_3703 ( P3_R1161_U474 , P3_R1161_U472 , P3_R1161_U262 );
nand NAND2_3704 ( P3_R1161_U473 , P3_R1161_U361 , P3_R1161_U92 );
nand NAND2_3705 ( P3_R1161_U472 , P3_R1161_U471 , P3_R1161_U470 );
nand NAND2_3706 ( P3_R1161_U471 , P3_U3437 , P3_R1161_U57 );
nand NAND2_3707 ( P3_R1161_U470 , P3_U3072 , P3_R1161_U56 );
nand NAND2_3708 ( P3_R1161_U469 , P3_U3440 , P3_R1161_U58 );
and AND2_3709 ( P2_U3014 , P2_U3924 , P2_U5671 );
and AND2_3710 ( P2_U3015 , P2_U3937 , P2_U3419 );
and AND2_3711 ( P2_U3016 , P2_U3575 , P2_U3570 );
and AND2_3712 ( P2_U3017 , P2_U5688 , P2_U3423 );
and AND2_3713 ( P2_U3018 , P2_U3426 , P2_U3423 );
and AND2_3714 ( P2_U3019 , P2_U3421 , P2_U3422 );
and AND2_3715 ( P2_U3020 , P2_U5680 , P2_U3421 );
and AND2_3716 ( P2_U3021 , P2_U5677 , P2_U3422 );
and AND2_3717 ( P2_U3022 , P2_U5677 , P2_U5680 );
and AND2_3718 ( P2_U3023 , P2_U3048 , P2_STATE_REG );
and AND2_3719 ( P2_U3024 , P2_U3757 , P2_U3401 );
and AND2_3720 ( P2_U3025 , P2_U3976 , P2_U5671 );
and AND2_3721 ( P2_U3026 , P2_U3963 , P2_U5683 );
and AND2_3722 ( P2_U3027 , P2_U3944 , P2_U5671 );
and AND2_3723 ( P2_U3028 , P2_U3803 , P2_U3946 );
and AND2_3724 ( P2_U3029 , P2_R1299_U6 , P2_U3411 );
and AND2_3725 ( P2_U3030 , P2_U3329 , P2_STATE_REG );
and AND2_3726 ( P2_U3031 , P2_U3932 , P2_U3964 );
and AND2_3727 ( P2_U3032 , P2_U3964 , P2_U3398 );
and AND2_3728 ( P2_U3033 , P2_U3933 , P2_U3964 );
and AND2_3729 ( P2_U3034 , P2_U3938 , P2_U3964 );
and AND2_3730 ( P2_U3035 , P2_U3963 , P2_U3423 );
and AND2_3731 ( P2_U3036 , P2_U3946 , P2_U5683 );
and AND2_3732 ( P2_U3037 , P2_U3964 , P2_U3026 );
and AND2_3733 ( P2_U3038 , P2_U3946 , P2_U3423 );
and AND2_3734 ( P2_U3039 , P2_U5688 , P2_U4854 );
and AND2_3735 ( P2_U3040 , P2_U3024 , P2_U5688 );
and AND2_3736 ( P2_U3041 , P2_U5683 , P2_U4854 );
and AND2_3737 ( P2_U3042 , P2_U3024 , P2_U5683 );
and AND2_3738 ( P2_U3043 , P2_U3018 , P2_U4854 );
and AND2_3739 ( P2_U3044 , P2_U3024 , P2_U3018 );
and AND2_3740 ( P2_U3045 , P2_U3023 , P2_U3401 );
and AND2_3741 ( P2_U3046 , P2_U5184 , P2_STATE_REG );
and AND2_3742 ( P2_U3047 , P2_U3023 , P2_U5186 );
and AND2_3743 ( P2_U3048 , P2_U5658 , P2_U3396 );
and AND2_3744 ( P2_U3049 , P2_U3418 , P2_U5668 );
and AND2_3745 ( P2_U3050 , P2_U3576 , P2_U3016 );
and AND5_3746 ( P2_U3051 , P2_U3341 , P2_U3402 , P2_U3392 , P2_U3338 , P2_U3337 );
and AND2_3747 ( P2_U3052 , P2_U3399 , P2_STATE_REG );
and AND3_3748 ( P2_U3053 , P2_U3820 , P2_U5439 , P2_U3819 );
and AND2_3749 ( P2_U3054 , P2_U5461 , P2_U5460 );
nand NAND4_3750 ( P2_U3055 , P2_U4611 , P2_U4612 , P2_U4610 , P2_U4613 );
nand NAND4_3751 ( P2_U3056 , P2_U4630 , P2_U4631 , P2_U4629 , P2_U4632 );
nand NAND4_3752 ( P2_U3057 , P2_U4651 , P2_U4650 , P2_U4649 , P2_U4648 );
nand NAND3_3753 ( P2_U3058 , P2_U4688 , P2_U4689 , P2_U4687 );
nand NAND4_3754 ( P2_U3059 , P2_U4592 , P2_U4593 , P2_U4591 , P2_U4594 );
nand NAND4_3755 ( P2_U3060 , P2_U4573 , P2_U4574 , P2_U4572 , P2_U4575 );
nand NAND3_3756 ( P2_U3061 , P2_U4668 , P2_U4669 , P2_U4667 );
nand NAND4_3757 ( P2_U3062 , P2_U4176 , P2_U4175 , P2_U4174 , P2_U4173 );
nand NAND4_3758 ( P2_U3063 , P2_U4516 , P2_U4517 , P2_U4515 , P2_U4518 );
nand NAND4_3759 ( P2_U3064 , P2_U4290 , P2_U4289 , P2_U4288 , P2_U4287 );
nand NAND4_3760 ( P2_U3065 , P2_U4309 , P2_U4308 , P2_U4307 , P2_U4306 );
nand NAND4_3761 ( P2_U3066 , P2_U4157 , P2_U4156 , P2_U4155 , P2_U4154 );
nand NAND4_3762 ( P2_U3067 , P2_U4554 , P2_U4555 , P2_U4553 , P2_U4556 );
nand NAND4_3763 ( P2_U3068 , P2_U4535 , P2_U4536 , P2_U4534 , P2_U4537 );
nand NAND4_3764 ( P2_U3069 , P2_U4195 , P2_U4194 , P2_U4193 , P2_U4192 );
nand NAND4_3765 ( P2_U3070 , P2_U4133 , P2_U4132 , P2_U4131 , P2_U4130 );
nand NAND4_3766 ( P2_U3071 , P2_U4421 , P2_U4422 , P2_U4420 , P2_U4423 );
nand NAND4_3767 ( P2_U3072 , P2_U4233 , P2_U4232 , P2_U4231 , P2_U4230 );
nand NAND4_3768 ( P2_U3073 , P2_U4214 , P2_U4213 , P2_U4212 , P2_U4211 );
nand NAND4_3769 ( P2_U3074 , P2_U4328 , P2_U4327 , P2_U4326 , P2_U4325 );
nand NAND4_3770 ( P2_U3075 , P2_U4404 , P2_U4403 , P2_U4402 , P2_U4401 );
nand NAND4_3771 ( P2_U3076 , P2_U4385 , P2_U4384 , P2_U4383 , P2_U4382 );
nand NAND4_3772 ( P2_U3077 , P2_U4497 , P2_U4498 , P2_U4496 , P2_U4499 );
nand NAND4_3773 ( P2_U3078 , P2_U4478 , P2_U4479 , P2_U4477 , P2_U4480 );
nand NAND4_3774 ( P2_U3079 , P2_U4138 , P2_U4137 , P2_U4136 , P2_U4135 );
nand NAND4_3775 ( P2_U3080 , P2_U4114 , P2_U4113 , P2_U4112 , P2_U4111 );
nand NAND4_3776 ( P2_U3081 , P2_U4366 , P2_U4365 , P2_U4364 , P2_U4363 );
nand NAND4_3777 ( P2_U3082 , P2_U4347 , P2_U4346 , P2_U4345 , P2_U4344 );
nand NAND4_3778 ( P2_U3083 , P2_U4459 , P2_U4460 , P2_U4458 , P2_U4461 );
nand NAND4_3779 ( P2_U3084 , P2_U4440 , P2_U4441 , P2_U4439 , P2_U4442 );
nand NAND4_3780 ( P2_U3085 , P2_U4271 , P2_U4270 , P2_U4269 , P2_U4268 );
nand NAND4_3781 ( P2_U3086 , P2_U4252 , P2_U4251 , P2_U4250 , P2_U4249 );
nand NAND2_3782 ( P2_U3087 , P2_U3815 , P2_U5434 );
not NOT1_3783 ( P2_U3088 , P2_STATE_REG );
nand NAND2_3784 ( P2_U3089 , P2_U5557 , P2_U5556 );
nand NAND2_3785 ( P2_U3090 , P2_U5559 , P2_U5558 );
nand NAND2_3786 ( P2_U3091 , P2_U3859 , P2_U5563 );
nand NAND2_3787 ( P2_U3092 , P2_U3860 , P2_U5566 );
nand NAND2_3788 ( P2_U3093 , P2_U3861 , P2_U5569 );
nand NAND2_3789 ( P2_U3094 , P2_U3862 , P2_U5572 );
nand NAND2_3790 ( P2_U3095 , P2_U3863 , P2_U5575 );
nand NAND2_3791 ( P2_U3096 , P2_U3864 , P2_U5578 );
nand NAND2_3792 ( P2_U3097 , P2_U3865 , P2_U5581 );
nand NAND2_3793 ( P2_U3098 , P2_U3866 , P2_U5584 );
nand NAND2_3794 ( P2_U3099 , P2_U3867 , P2_U5587 );
nand NAND2_3795 ( P2_U3100 , P2_U3868 , P2_U5590 );
nand NAND2_3796 ( P2_U3101 , P2_U3869 , P2_U5596 );
nand NAND2_3797 ( P2_U3102 , P2_U3870 , P2_U5599 );
nand NAND2_3798 ( P2_U3103 , P2_U3871 , P2_U5602 );
nand NAND2_3799 ( P2_U3104 , P2_U3872 , P2_U5605 );
nand NAND2_3800 ( P2_U3105 , P2_U3873 , P2_U5608 );
nand NAND2_3801 ( P2_U3106 , P2_U3874 , P2_U5611 );
nand NAND2_3802 ( P2_U3107 , P2_U3875 , P2_U5614 );
nand NAND2_3803 ( P2_U3108 , P2_U3876 , P2_U5617 );
nand NAND2_3804 ( P2_U3109 , P2_U3877 , P2_U5620 );
nand NAND2_3805 ( P2_U3110 , P2_U3878 , P2_U5623 );
nand NAND2_3806 ( P2_U3111 , P2_U3857 , P2_U5538 );
nand NAND2_3807 ( P2_U3112 , P2_U3858 , P2_U5541 );
nand NAND3_3808 ( P2_U3113 , P2_U5545 , P2_U5544 , P2_U5546 );
nand NAND3_3809 ( P2_U3114 , P2_U5548 , P2_U5547 , P2_U5549 );
nand NAND3_3810 ( P2_U3115 , P2_U5551 , P2_U5550 , P2_U5552 );
nand NAND3_3811 ( P2_U3116 , P2_U5554 , P2_U5553 , P2_U5555 );
nand NAND3_3812 ( P2_U3117 , P2_U5561 , P2_U5560 , P2_U5562 );
nand NAND3_3813 ( P2_U3118 , P2_U5594 , P2_U5593 , P2_U5595 );
nand NAND3_3814 ( P2_U3119 , P2_U5627 , P2_U5626 , P2_U5628 );
nand NAND2_3815 ( P2_U3120 , P2_U5630 , P2_U5629 );
and AND3_3816 ( P2_U3121 , P2_U5637 , P2_U5632 , P2_U5638 );
nand NAND3_3817 ( P2_U3122 , P2_U5463 , P2_U5462 , P2_U5464 );
nand NAND3_3818 ( P2_U3123 , P2_U5469 , P2_U3831 , P2_U5470 );
nand NAND3_3819 ( P2_U3124 , P2_U5472 , P2_U3832 , P2_U5473 );
nand NAND3_3820 ( P2_U3125 , P2_U5475 , P2_U3833 , P2_U5476 );
nand NAND3_3821 ( P2_U3126 , P2_U5478 , P2_U3834 , P2_U5479 );
nand NAND3_3822 ( P2_U3127 , P2_U5481 , P2_U3835 , P2_U5482 );
nand NAND3_3823 ( P2_U3128 , P2_U5484 , P2_U3836 , P2_U5485 );
nand NAND3_3824 ( P2_U3129 , P2_U5487 , P2_U3837 , P2_U5488 );
nand NAND3_3825 ( P2_U3130 , P2_U5490 , P2_U3838 , P2_U5491 );
nand NAND3_3826 ( P2_U3131 , P2_U5493 , P2_U3839 , P2_U5494 );
nand NAND3_3827 ( P2_U3132 , P2_U5496 , P2_U3840 , P2_U5497 );
nand NAND3_3828 ( P2_U3133 , P2_U5502 , P2_U3843 , P2_U5503 );
nand NAND3_3829 ( P2_U3134 , P2_U5505 , P2_U3844 , P2_U5506 );
nand NAND3_3830 ( P2_U3135 , P2_U5508 , P2_U3845 , P2_U5509 );
nand NAND3_3831 ( P2_U3136 , P2_U5511 , P2_U3846 , P2_U5512 );
nand NAND3_3832 ( P2_U3137 , P2_U5514 , P2_U3847 , P2_U5515 );
nand NAND3_3833 ( P2_U3138 , P2_U5517 , P2_U3848 , P2_U5518 );
nand NAND3_3834 ( P2_U3139 , P2_U5520 , P2_U3849 , P2_U5521 );
nand NAND3_3835 ( P2_U3140 , P2_U5523 , P2_U3850 , P2_U5524 );
nand NAND3_3836 ( P2_U3141 , P2_U5526 , P2_U5525 , P2_U3851 );
nand NAND3_3837 ( P2_U3142 , P2_U5529 , P2_U5528 , P2_U3852 );
nand NAND3_3838 ( P2_U3143 , P2_U5443 , P2_U5442 , P2_U3821 );
nand NAND3_3839 ( P2_U3144 , P2_U5446 , P2_U5445 , P2_U3822 );
nand NAND3_3840 ( P2_U3145 , P2_U5449 , P2_U5448 , P2_U3823 );
nand NAND3_3841 ( P2_U3146 , P2_U5452 , P2_U5451 , P2_U3824 );
nand NAND3_3842 ( P2_U3147 , P2_U5455 , P2_U5454 , P2_U3825 );
nand NAND2_3843 ( P2_U3148 , P2_U5458 , P2_U3826 );
nand NAND2_3844 ( P2_U3149 , P2_U5466 , P2_U3829 );
nand NAND2_3845 ( P2_U3150 , P2_U5499 , P2_U3841 );
nand NAND2_3846 ( P2_U3151 , P2_U5532 , P2_U3853 );
nand NAND2_3847 ( P2_U3152 , P2_U5535 , P2_U3855 );
nand NAND3_3848 ( P2_U3153 , P2_U3817 , P2_U3345 , P2_U3415 );
nand NAND2_3849 ( P2_U3154 , P2_U3015 , P2_U5658 );
and AND2_3850 ( P2_U3155 , P2_U5437 , P2_U3056 );
and AND2_3851 ( P2_U3156 , P2_U5437 , P2_U3055 );
and AND2_3852 ( P2_U3157 , P2_U5437 , P2_U3059 );
and AND2_3853 ( P2_U3158 , P2_U5437 , P2_U3060 );
and AND2_3854 ( P2_U3159 , P2_U5437 , P2_U3067 );
and AND2_3855 ( P2_U3160 , P2_U5437 , P2_U3068 );
and AND2_3856 ( P2_U3161 , P2_U5437 , P2_U3063 );
and AND2_3857 ( P2_U3162 , P2_U5437 , P2_U3077 );
and AND2_3858 ( P2_U3163 , P2_U5437 , P2_U3078 );
and AND2_3859 ( P2_U3164 , P2_U5437 , P2_U3083 );
and AND2_3860 ( P2_U3165 , P2_U5437 , P2_U3084 );
and AND2_3861 ( P2_U3166 , P2_U5437 , P2_U3071 );
and AND2_3862 ( P2_U3167 , P2_U5437 , P2_U3075 );
and AND2_3863 ( P2_U3168 , P2_U5437 , P2_U3076 );
and AND2_3864 ( P2_U3169 , P2_U5437 , P2_U3081 );
and AND2_3865 ( P2_U3170 , P2_U5437 , P2_U3082 );
and AND2_3866 ( P2_U3171 , P2_U5437 , P2_U3074 );
and AND2_3867 ( P2_U3172 , P2_U5437 , P2_U3065 );
and AND2_3868 ( P2_U3173 , P2_U5437 , P2_U3064 );
and AND2_3869 ( P2_U3174 , P2_U5437 , P2_U3085 );
and AND2_3870 ( P2_U3175 , P2_U5437 , P2_U3086 );
and AND2_3871 ( P2_U3176 , P2_U5437 , P2_U3072 );
and AND2_3872 ( P2_U3177 , P2_U5437 , P2_U3073 );
and AND2_3873 ( P2_U3178 , P2_U5437 , P2_U3069 );
and AND2_3874 ( P2_U3179 , P2_U5437 , P2_U3062 );
and AND2_3875 ( P2_U3180 , P2_U5437 , P2_U3066 );
and AND2_3876 ( P2_U3181 , P2_U5437 , P2_U3070 );
and AND2_3877 ( P2_U3182 , P2_U5437 , P2_U3080 );
and AND2_3878 ( P2_U3183 , P2_U5437 , P2_U3079 );
nand NAND3_3879 ( P2_U3184 , P2_U3404 , P2_U5436 , P2_U3343 );
nand NAND4_3880 ( P2_U3185 , P2_U5433 , P2_U5432 , P2_U3814 , P2_U5430 );
nand NAND5_3881 ( P2_U3186 , P2_U5424 , P2_U5423 , P2_U5421 , P2_U5420 , P2_U5422 );
nand NAND5_3882 ( P2_U3187 , P2_U5412 , P2_U5411 , P2_U5415 , P2_U5414 , P2_U5413 );
nand NAND5_3883 ( P2_U3188 , P2_U5406 , P2_U5405 , P2_U5403 , P2_U5402 , P2_U5404 );
nand NAND5_3884 ( P2_U3189 , P2_U5394 , P2_U5393 , P2_U5395 , P2_U5397 , P2_U5396 );
nand NAND4_3885 ( P2_U3190 , P2_U5388 , P2_U5387 , P2_U3813 , P2_U5385 );
nand NAND5_3886 ( P2_U3191 , P2_U5376 , P2_U5375 , P2_U5379 , P2_U5378 , P2_U5377 );
nand NAND5_3887 ( P2_U3192 , P2_U5370 , P2_U5369 , P2_U5367 , P2_U5366 , P2_U5368 );
nand NAND4_3888 ( P2_U3193 , P2_U5361 , P2_U5360 , P2_U3812 , P2_U5358 );
nand NAND4_3889 ( P2_U3194 , P2_U5352 , P2_U5351 , P2_U3811 , P2_U5349 );
nand NAND5_3890 ( P2_U3195 , P2_U5340 , P2_U5339 , P2_U5343 , P2_U5342 , P2_U5341 );
nand NAND5_3891 ( P2_U3196 , P2_U5331 , P2_U5330 , P2_U5334 , P2_U5333 , P2_U5332 );
nand NAND5_3892 ( P2_U3197 , P2_U5325 , P2_U5324 , P2_U5322 , P2_U5321 , P2_U5323 );
nand NAND5_3893 ( P2_U3198 , P2_U5313 , P2_U5312 , P2_U5316 , P2_U5315 , P2_U5314 );
nand NAND4_3894 ( P2_U3199 , P2_U5307 , P2_U5306 , P2_U3810 , P2_U5304 );
nand NAND5_3895 ( P2_U3200 , P2_U5295 , P2_U5294 , P2_U5298 , P2_U5297 , P2_U5296 );
nand NAND5_3896 ( P2_U3201 , P2_U5289 , P2_U5288 , P2_U5286 , P2_U5285 , P2_U5287 );
nand NAND4_3897 ( P2_U3202 , P2_U5280 , P2_U5279 , P2_U3809 , P2_U5277 );
nand NAND5_3898 ( P2_U3203 , P2_U5268 , P2_U5267 , P2_U5269 , P2_U5271 , P2_U5270 );
nand NAND3_3899 ( P2_U3204 , P2_U3808 , P2_U5260 , P2_U3807 );
nand NAND5_3900 ( P2_U3205 , P2_U5251 , P2_U5250 , P2_U5254 , P2_U5253 , P2_U5252 );
nand NAND5_3901 ( P2_U3206 , P2_U5242 , P2_U5241 , P2_U5245 , P2_U5244 , P2_U5243 );
nand NAND5_3902 ( P2_U3207 , P2_U5236 , P2_U5235 , P2_U5233 , P2_U5232 , P2_U5234 );
nand NAND5_3903 ( P2_U3208 , P2_U5224 , P2_U5223 , P2_U5225 , P2_U5227 , P2_U5226 );
nand NAND4_3904 ( P2_U3209 , P2_U5218 , P2_U5217 , P2_U3805 , P2_U5215 );
nand NAND5_3905 ( P2_U3210 , P2_U5206 , P2_U5205 , P2_U5209 , P2_U5208 , P2_U5207 );
nand NAND4_3906 ( P2_U3211 , P2_U5200 , P2_U5199 , P2_U3804 , P2_U5197 );
nand NAND5_3907 ( P2_U3212 , P2_U5191 , P2_U5190 , P2_U5188 , P2_U5187 , P2_U5189 );
nand NAND5_3908 ( P2_U3213 , P2_U5175 , P2_U5174 , P2_U5178 , P2_U5177 , P2_U5176 );
nand NAND4_3909 ( P2_U3214 , P2_U5150 , P2_U5149 , P2_U3785 , P2_U3786 );
nand NAND4_3910 ( P2_U3215 , P2_U5135 , P2_U5134 , P2_U3783 , P2_U3784 );
nand NAND4_3911 ( P2_U3216 , P2_U5120 , P2_U5119 , P2_U3781 , P2_U3782 );
nand NAND4_3912 ( P2_U3217 , P2_U5105 , P2_U5104 , P2_U3779 , P2_U3780 );
nand NAND4_3913 ( P2_U3218 , P2_U5090 , P2_U5089 , P2_U3777 , P2_U3778 );
nand NAND4_3914 ( P2_U3219 , P2_U5075 , P2_U5074 , P2_U3775 , P2_U3776 );
nand NAND4_3915 ( P2_U3220 , P2_U5060 , P2_U5059 , P2_U3773 , P2_U3774 );
nand NAND4_3916 ( P2_U3221 , P2_U5045 , P2_U5044 , P2_U3771 , P2_U3772 );
nand NAND4_3917 ( P2_U3222 , P2_U5030 , P2_U5029 , P2_U3769 , P2_U3770 );
nand NAND3_3918 ( P2_U3223 , P2_U5015 , P2_U5014 , P2_U3768 );
nand NAND3_3919 ( P2_U3224 , P2_U5000 , P2_U4999 , P2_U3767 );
nand NAND3_3920 ( P2_U3225 , P2_U4985 , P2_U4984 , P2_U3766 );
nand NAND3_3921 ( P2_U3226 , P2_U4970 , P2_U4969 , P2_U3765 );
nand NAND3_3922 ( P2_U3227 , P2_U4955 , P2_U4954 , P2_U3764 );
nand NAND3_3923 ( P2_U3228 , P2_U4940 , P2_U4939 , P2_U3763 );
nand NAND3_3924 ( P2_U3229 , P2_U4925 , P2_U4924 , P2_U3762 );
nand NAND3_3925 ( P2_U3230 , P2_U4910 , P2_U4909 , P2_U3761 );
nand NAND3_3926 ( P2_U3231 , P2_U4895 , P2_U4894 , P2_U3760 );
nand NAND3_3927 ( P2_U3232 , P2_U4880 , P2_U4879 , P2_U3759 );
nand NAND3_3928 ( P2_U3233 , P2_U4865 , P2_U4864 , P2_U3758 );
nand NAND3_3929 ( P2_U3234 , P2_U3915 , P2_U4852 , P2_U4853 );
nand NAND3_3930 ( P2_U3235 , P2_U3914 , P2_U4850 , P2_U4851 );
nand NAND5_3931 ( P2_U3236 , P2_U4847 , P2_U4848 , P2_U4849 , P2_U4846 , P2_U3912 );
nand NAND4_3932 ( P2_U3237 , P2_U3753 , P2_U3754 , P2_U4842 , P2_U3911 );
nand NAND4_3933 ( P2_U3238 , P2_U3751 , P2_U3752 , P2_U4837 , P2_U3910 );
nand NAND4_3934 ( P2_U3239 , P2_U3749 , P2_U3750 , P2_U4832 , P2_U3909 );
nand NAND4_3935 ( P2_U3240 , P2_U3747 , P2_U3748 , P2_U4827 , P2_U3908 );
nand NAND4_3936 ( P2_U3241 , P2_U3745 , P2_U3746 , P2_U4822 , P2_U3907 );
nand NAND4_3937 ( P2_U3242 , P2_U3743 , P2_U3744 , P2_U4817 , P2_U3906 );
nand NAND4_3938 ( P2_U3243 , P2_U3741 , P2_U3742 , P2_U4812 , P2_U3905 );
nand NAND4_3939 ( P2_U3244 , P2_U3739 , P2_U3740 , P2_U4807 , P2_U3904 );
nand NAND4_3940 ( P2_U3245 , P2_U3737 , P2_U3738 , P2_U4802 , P2_U3903 );
nand NAND4_3941 ( P2_U3246 , P2_U3735 , P2_U3736 , P2_U4797 , P2_U3902 );
nand NAND4_3942 ( P2_U3247 , P2_U3733 , P2_U3734 , P2_U4792 , P2_U3901 );
nand NAND4_3943 ( P2_U3248 , P2_U3731 , P2_U3732 , P2_U4787 , P2_U3900 );
nand NAND4_3944 ( P2_U3249 , P2_U3729 , P2_U3730 , P2_U4782 , P2_U3899 );
nand NAND3_3945 ( P2_U3250 , P2_U3728 , P2_U3727 , P2_U3898 );
nand NAND3_3946 ( P2_U3251 , P2_U3726 , P2_U3725 , P2_U3897 );
nand NAND3_3947 ( P2_U3252 , P2_U3724 , P2_U3723 , P2_U3896 );
nand NAND3_3948 ( P2_U3253 , P2_U3722 , P2_U3721 , P2_U3895 );
nand NAND3_3949 ( P2_U3254 , P2_U3720 , P2_U3719 , P2_U3894 );
nand NAND3_3950 ( P2_U3255 , P2_U3718 , P2_U3717 , P2_U3893 );
nand NAND2_3951 ( P2_U3256 , P2_U3716 , P2_U3715 );
nand NAND2_3952 ( P2_U3257 , P2_U3714 , P2_U3713 );
nand NAND2_3953 ( P2_U3258 , P2_U3712 , P2_U3711 );
nand NAND2_3954 ( P2_U3259 , P2_U3710 , P2_U3709 );
nand NAND2_3955 ( P2_U3260 , P2_U3708 , P2_U3707 );
nand NAND2_3956 ( P2_U3261 , P2_U3706 , P2_U3705 );
nand NAND2_3957 ( P2_U3262 , P2_U3704 , P2_U3703 );
nand NAND2_3958 ( P2_U3263 , P2_U3702 , P2_U3701 );
nand NAND2_3959 ( P2_U3264 , P2_U3700 , P2_U3699 );
nand NAND2_3960 ( P2_U3265 , P2_U3698 , P2_U3697 );
and AND2_3961 ( P2_U3266 , P2_D_REG_31_ , P2_U3880 );
and AND2_3962 ( P2_U3267 , P2_D_REG_30_ , P2_U3880 );
and AND2_3963 ( P2_U3268 , P2_D_REG_29_ , P2_U3880 );
and AND2_3964 ( P2_U3269 , P2_D_REG_28_ , P2_U3880 );
and AND2_3965 ( P2_U3270 , P2_D_REG_27_ , P2_U3880 );
and AND2_3966 ( P2_U3271 , P2_D_REG_26_ , P2_U3880 );
and AND2_3967 ( P2_U3272 , P2_D_REG_25_ , P2_U3880 );
and AND2_3968 ( P2_U3273 , P2_D_REG_24_ , P2_U3880 );
and AND2_3969 ( P2_U3274 , P2_D_REG_23_ , P2_U3880 );
and AND2_3970 ( P2_U3275 , P2_D_REG_22_ , P2_U3880 );
and AND2_3971 ( P2_U3276 , P2_D_REG_21_ , P2_U3880 );
and AND2_3972 ( P2_U3277 , P2_D_REG_20_ , P2_U3880 );
and AND2_3973 ( P2_U3278 , P2_D_REG_19_ , P2_U3880 );
and AND2_3974 ( P2_U3279 , P2_D_REG_18_ , P2_U3880 );
and AND2_3975 ( P2_U3280 , P2_D_REG_17_ , P2_U3880 );
and AND2_3976 ( P2_U3281 , P2_D_REG_16_ , P2_U3880 );
and AND2_3977 ( P2_U3282 , P2_D_REG_15_ , P2_U3880 );
and AND2_3978 ( P2_U3283 , P2_D_REG_14_ , P2_U3880 );
and AND2_3979 ( P2_U3284 , P2_D_REG_13_ , P2_U3880 );
and AND2_3980 ( P2_U3285 , P2_D_REG_12_ , P2_U3880 );
and AND2_3981 ( P2_U3286 , P2_D_REG_11_ , P2_U3880 );
and AND2_3982 ( P2_U3287 , P2_D_REG_10_ , P2_U3880 );
and AND2_3983 ( P2_U3288 , P2_D_REG_9_ , P2_U3880 );
and AND2_3984 ( P2_U3289 , P2_D_REG_8_ , P2_U3880 );
and AND2_3985 ( P2_U3290 , P2_D_REG_7_ , P2_U3880 );
and AND2_3986 ( P2_U3291 , P2_D_REG_6_ , P2_U3880 );
and AND2_3987 ( P2_U3292 , P2_D_REG_5_ , P2_U3880 );
and AND2_3988 ( P2_U3293 , P2_D_REG_4_ , P2_U3880 );
and AND2_3989 ( P2_U3294 , P2_D_REG_3_ , P2_U3880 );
and AND2_3990 ( P2_U3295 , P2_D_REG_2_ , P2_U3880 );
nand NAND3_3991 ( P2_U3296 , P2_U4073 , P2_U4074 , P2_U4072 );
nand NAND3_3992 ( P2_U3297 , P2_U4070 , P2_U4071 , P2_U4069 );
nand NAND3_3993 ( P2_U3298 , P2_U4067 , P2_U4068 , P2_U4066 );
nand NAND3_3994 ( P2_U3299 , P2_U4064 , P2_U4065 , P2_U4063 );
nand NAND3_3995 ( P2_U3300 , P2_U4061 , P2_U4062 , P2_U4060 );
nand NAND3_3996 ( P2_U3301 , P2_U4058 , P2_U4059 , P2_U4057 );
nand NAND3_3997 ( P2_U3302 , P2_U4055 , P2_U4056 , P2_U4054 );
nand NAND3_3998 ( P2_U3303 , P2_U4052 , P2_U4053 , P2_U4051 );
nand NAND3_3999 ( P2_U3304 , P2_U4049 , P2_U4050 , P2_U4048 );
nand NAND3_4000 ( P2_U3305 , P2_U4046 , P2_U4047 , P2_U4045 );
nand NAND3_4001 ( P2_U3306 , P2_U4043 , P2_U4044 , P2_U4042 );
nand NAND3_4002 ( P2_U3307 , P2_U4040 , P2_U4041 , P2_U4039 );
nand NAND3_4003 ( P2_U3308 , P2_U4037 , P2_U4038 , P2_U4036 );
nand NAND3_4004 ( P2_U3309 , P2_U4034 , P2_U4035 , P2_U4033 );
nand NAND3_4005 ( P2_U3310 , P2_U4031 , P2_U4032 , P2_U4030 );
nand NAND3_4006 ( P2_U3311 , P2_U4028 , P2_U4029 , P2_U4027 );
nand NAND3_4007 ( P2_U3312 , P2_U4025 , P2_U4026 , P2_U4024 );
nand NAND3_4008 ( P2_U3313 , P2_U4022 , P2_U4023 , P2_U4021 );
nand NAND3_4009 ( P2_U3314 , P2_U4019 , P2_U4020 , P2_U4018 );
nand NAND3_4010 ( P2_U3315 , P2_U4016 , P2_U4017 , P2_U4015 );
nand NAND3_4011 ( P2_U3316 , P2_U4013 , P2_U4014 , P2_U4012 );
nand NAND3_4012 ( P2_U3317 , P2_U4010 , P2_U4011 , P2_U4009 );
nand NAND3_4013 ( P2_U3318 , P2_U4007 , P2_U4008 , P2_U4006 );
nand NAND3_4014 ( P2_U3319 , P2_U4004 , P2_U4005 , P2_U4003 );
nand NAND3_4015 ( P2_U3320 , P2_U4001 , P2_U4002 , P2_U4000 );
nand NAND3_4016 ( P2_U3321 , P2_U3998 , P2_U3999 , P2_U3997 );
nand NAND3_4017 ( P2_U3322 , P2_U3995 , P2_U3996 , P2_U3994 );
nand NAND3_4018 ( P2_U3323 , P2_U3992 , P2_U3993 , P2_U3991 );
nand NAND3_4019 ( P2_U3324 , P2_U3989 , P2_U3990 , P2_U3988 );
nand NAND3_4020 ( P2_U3325 , P2_U3986 , P2_U3987 , P2_U3985 );
nand NAND3_4021 ( P2_U3326 , P2_U3983 , P2_U3984 , P2_U3982 );
nand NAND3_4022 ( P2_U3327 , P2_U3980 , P2_U3981 , P2_U3979 );
and AND2_4023 ( P2_U3328 , P2_U3797 , P2_U5641 );
nand NAND2_4024 ( P2_U3329 , P2_STATE_REG , P2_U3879 );
not NOT1_4025 ( P2_U3330 , U69 );
not NOT1_4026 ( P2_U3331 , P2_B_REG );
nand NAND2_4027 ( P2_U3332 , P2_U3414 , P2_U5649 );
nand NAND2_4028 ( P2_U3333 , P2_U3414 , P2_U4075 );
nand NAND3_4029 ( P2_U3334 , P2_U5671 , P2_U3424 , P2_U3420 );
nand NAND3_4030 ( P2_U3335 , P2_U3418 , P2_U3424 , P2_U3420 );
nand NAND2_4031 ( P2_U3336 , P2_U3049 , P2_U3420 );
nand NAND3_4032 ( P2_U3337 , P2_U3418 , P2_U3424 , P2_U3419 );
nand NAND2_4033 ( P2_U3338 , P2_U3049 , P2_U3419 );
nand NAND3_4034 ( P2_U3339 , P2_U5668 , P2_U5674 , P2_U3420 );
nand NAND2_4035 ( P2_U3340 , P2_U5671 , P2_U5668 );
nand NAND2_4036 ( P2_U3341 , P2_U3974 , P2_U3419 );
nand NAND2_4037 ( P2_U3342 , P2_U3939 , P2_U5665 );
nand NAND2_4038 ( P2_U3343 , P2_U5665 , P2_U5674 );
nand NAND2_4039 ( P2_U3344 , P2_U3420 , P2_U3419 );
nand NAND2_4040 ( P2_U3345 , P2_U5665 , P2_U3424 );
nand NAND2_4041 ( P2_U3346 , P2_U3049 , P2_U5665 );
nand NAND2_4042 ( P2_U3347 , P2_U5688 , P2_U5683 );
nand NAND3_4043 ( P2_U3348 , P2_U3564 , P2_U4123 , P2_U3563 );
nand NAND4_4044 ( P2_U3349 , P2_U4141 , P2_U4140 , P2_U3578 , P2_U3580 );
nand NAND4_4045 ( P2_U3350 , P2_U4160 , P2_U4159 , P2_U3582 , P2_U3584 );
nand NAND4_4046 ( P2_U3351 , P2_U4179 , P2_U4178 , P2_U3586 , P2_U3588 );
nand NAND4_4047 ( P2_U3352 , P2_U4198 , P2_U4197 , P2_U3590 , P2_U3592 );
nand NAND4_4048 ( P2_U3353 , P2_U4217 , P2_U4216 , P2_U3594 , P2_U3596 );
nand NAND4_4049 ( P2_U3354 , P2_U4236 , P2_U4235 , P2_U3598 , P2_U3600 );
nand NAND4_4050 ( P2_U3355 , P2_U4255 , P2_U4254 , P2_U3602 , P2_U3604 );
nand NAND4_4051 ( P2_U3356 , P2_U4274 , P2_U4273 , P2_U3606 , P2_U3608 );
nand NAND4_4052 ( P2_U3357 , P2_U4293 , P2_U4292 , P2_U3610 , P2_U3612 );
nand NAND4_4053 ( P2_U3358 , P2_U4312 , P2_U4311 , P2_U3614 , P2_U3616 );
nand NAND4_4054 ( P2_U3359 , P2_U4331 , P2_U4330 , P2_U3618 , P2_U3620 );
nand NAND4_4055 ( P2_U3360 , P2_U4350 , P2_U4349 , P2_U3622 , P2_U3624 );
nand NAND4_4056 ( P2_U3361 , P2_U4369 , P2_U4368 , P2_U3626 , P2_U3628 );
nand NAND4_4057 ( P2_U3362 , P2_U4388 , P2_U4387 , P2_U3630 , P2_U3632 );
nand NAND4_4058 ( P2_U3363 , P2_U4407 , P2_U4406 , P2_U3634 , P2_U3636 );
nand NAND4_4059 ( P2_U3364 , P2_U4426 , P2_U4425 , P2_U3638 , P2_U3640 );
nand NAND4_4060 ( P2_U3365 , P2_U4445 , P2_U4444 , P2_U3642 , P2_U3644 );
nand NAND4_4061 ( P2_U3366 , P2_U4464 , P2_U4463 , P2_U3646 , P2_U3648 );
nand NAND4_4062 ( P2_U3367 , P2_U4483 , P2_U4482 , P2_U3650 , P2_U3652 );
nand NAND2_4063 ( P2_U3368 , U81 , P2_U3347 );
nand NAND4_4064 ( P2_U3369 , P2_U4502 , P2_U4501 , P2_U3654 , P2_U3656 );
nand NAND2_4065 ( P2_U3370 , U80 , P2_U3347 );
nand NAND4_4066 ( P2_U3371 , P2_U4521 , P2_U4520 , P2_U3658 , P2_U3660 );
nand NAND2_4067 ( P2_U3372 , U79 , P2_U3347 );
nand NAND4_4068 ( P2_U3373 , P2_U4540 , P2_U4539 , P2_U3662 , P2_U3664 );
nand NAND2_4069 ( P2_U3374 , U78 , P2_U3347 );
nand NAND4_4070 ( P2_U3375 , P2_U4559 , P2_U4558 , P2_U3666 , P2_U3668 );
nand NAND2_4071 ( P2_U3376 , U77 , P2_U3347 );
nand NAND4_4072 ( P2_U3377 , P2_U4578 , P2_U4577 , P2_U3670 , P2_U3672 );
nand NAND2_4073 ( P2_U3378 , U76 , P2_U3347 );
nand NAND4_4074 ( P2_U3379 , P2_U4597 , P2_U4596 , P2_U3674 , P2_U3676 );
nand NAND2_4075 ( P2_U3380 , U75 , P2_U3347 );
nand NAND4_4076 ( P2_U3381 , P2_U4616 , P2_U4615 , P2_U3678 , P2_U3680 );
nand NAND2_4077 ( P2_U3382 , U74 , P2_U3347 );
nand NAND4_4078 ( P2_U3383 , P2_U4635 , P2_U4634 , P2_U3682 , P2_U3684 );
nand NAND2_4079 ( P2_U3384 , U73 , P2_U3347 );
nand NAND5_4080 ( P2_U3385 , P2_U4654 , P2_U4653 , P2_U4655 , P2_U4656 , P2_U3687 );
nand NAND2_4081 ( P2_U3386 , U72 , P2_U3347 );
nand NAND5_4082 ( P2_U3387 , P2_U4674 , P2_U4673 , P2_U4675 , P2_U3690 , P2_U3692 );
nand NAND2_4083 ( P2_U3388 , U70 , P2_U3347 );
nand NAND2_4084 ( P2_U3389 , U69 , P2_U3347 );
nand NAND2_4085 ( P2_U3390 , P2_U3944 , P2_U3424 );
nand NAND2_4086 ( P2_U3391 , P2_U3023 , P2_U4698 );
nand NAND3_4087 ( P2_U3392 , P2_U5671 , P2_U3424 , P2_U3419 );
nand NAND2_4088 ( P2_U3393 , P2_U3921 , P2_U5671 );
nand NAND2_4089 ( P2_U3394 , P2_U3944 , P2_U5668 );
nand NAND2_4090 ( P2_U3395 , P2_U3927 , P2_U5671 );
nand NAND3_4091 ( P2_U3396 , P2_U3413 , P2_U3412 , P2_U3414 );
nand NAND2_4092 ( P2_U3397 , P2_U3344 , P2_U3347 );
nand NAND2_4093 ( P2_U3398 , P2_U3934 , P2_U4699 );
nand NAND2_4094 ( P2_U3399 , P2_U3962 , P2_U5658 );
nand NAND2_4095 ( P2_U3400 , P2_U3977 , P2_STATE_REG );
nand NAND2_4096 ( P2_U3401 , P2_U3756 , P2_U3052 );
nand NAND2_4097 ( P2_U3402 , P2_U3974 , P2_U3420 );
nand NAND2_4098 ( P2_U3403 , P2_U3015 , P2_U3018 );
nand NAND2_4099 ( P2_U3404 , P2_U5674 , P2_U3424 );
nand NAND2_4100 ( P2_U3405 , P2_U3023 , P2_U3398 );
nand NAND2_4101 ( P2_U3406 , P2_U3798 , P2_U3016 );
nand NAND3_4102 ( P2_U3407 , P2_U5168 , P2_STATE_REG , P2_U3396 );
nand NAND2_4103 ( P2_U3408 , P2_U3802 , P2_U5172 );
not NOT1_4104 ( P2_U3409 , P2_R1299_U6 );
nand NAND2_4105 ( P2_U3410 , P2_U3938 , P2_U5665 );
nand NAND4_4106 ( P2_U3411 , P2_U3335 , P2_U3336 , P2_U3346 , P2_U3923 );
nand NAND2_4107 ( P2_U3412 , P2_U5645 , P2_U5644 );
nand NAND2_4108 ( P2_U3413 , P2_U5648 , P2_U5647 );
nand NAND2_4109 ( P2_U3414 , P2_U5651 , P2_U5650 );
nand NAND2_4110 ( P2_U3415 , P2_U5657 , P2_U5656 );
nand NAND2_4111 ( P2_U3416 , P2_U5660 , P2_U5659 );
nand NAND2_4112 ( P2_U3417 , P2_U5662 , P2_U5661 );
nand NAND2_4113 ( P2_U3418 , P2_U5670 , P2_U5669 );
nand NAND2_4114 ( P2_U3419 , P2_U5673 , P2_U5672 );
nand NAND2_4115 ( P2_U3420 , P2_U5664 , P2_U5663 );
nand NAND2_4116 ( P2_U3421 , P2_U5676 , P2_U5675 );
nand NAND2_4117 ( P2_U3422 , P2_U5679 , P2_U5678 );
nand NAND2_4118 ( P2_U3423 , P2_U5682 , P2_U5681 );
nand NAND2_4119 ( P2_U3424 , P2_U5667 , P2_U5666 );
nand NAND2_4120 ( P2_U3425 , P2_U5685 , P2_U5684 );
nand NAND2_4121 ( P2_U3426 , P2_U5687 , P2_U5686 );
nand NAND2_4122 ( P2_U3427 , P2_U5690 , P2_U5689 );
nand NAND2_4123 ( P2_U3428 , P2_U5698 , P2_U5697 );
nand NAND2_4124 ( P2_U3429 , P2_U5695 , P2_U5694 );
nand NAND2_4125 ( P2_U3430 , P2_U5701 , P2_U5700 );
nand NAND2_4126 ( P2_U3431 , P2_U5703 , P2_U5702 );
nand NAND2_4127 ( P2_U3432 , P2_U5705 , P2_U5704 );
nand NAND2_4128 ( P2_U3433 , P2_U5708 , P2_U5707 );
nand NAND2_4129 ( P2_U3434 , P2_U5710 , P2_U5709 );
nand NAND2_4130 ( P2_U3435 , P2_U5712 , P2_U5711 );
nand NAND2_4131 ( P2_U3436 , P2_U5715 , P2_U5714 );
nand NAND2_4132 ( P2_U3437 , P2_U5717 , P2_U5716 );
nand NAND2_4133 ( P2_U3438 , P2_U5719 , P2_U5718 );
nand NAND2_4134 ( P2_U3439 , P2_U5722 , P2_U5721 );
nand NAND2_4135 ( P2_U3440 , P2_U5724 , P2_U5723 );
nand NAND2_4136 ( P2_U3441 , P2_U5726 , P2_U5725 );
nand NAND2_4137 ( P2_U3442 , P2_U5729 , P2_U5728 );
nand NAND2_4138 ( P2_U3443 , P2_U5731 , P2_U5730 );
nand NAND2_4139 ( P2_U3444 , P2_U5733 , P2_U5732 );
nand NAND2_4140 ( P2_U3445 , P2_U5736 , P2_U5735 );
nand NAND2_4141 ( P2_U3446 , P2_U5738 , P2_U5737 );
nand NAND2_4142 ( P2_U3447 , P2_U5740 , P2_U5739 );
nand NAND2_4143 ( P2_U3448 , P2_U5743 , P2_U5742 );
nand NAND2_4144 ( P2_U3449 , P2_U5745 , P2_U5744 );
nand NAND2_4145 ( P2_U3450 , P2_U5747 , P2_U5746 );
nand NAND2_4146 ( P2_U3451 , P2_U5750 , P2_U5749 );
nand NAND2_4147 ( P2_U3452 , P2_U5752 , P2_U5751 );
nand NAND2_4148 ( P2_U3453 , P2_U5754 , P2_U5753 );
nand NAND2_4149 ( P2_U3454 , P2_U5757 , P2_U5756 );
nand NAND2_4150 ( P2_U3455 , P2_U5759 , P2_U5758 );
nand NAND2_4151 ( P2_U3456 , P2_U5761 , P2_U5760 );
nand NAND2_4152 ( P2_U3457 , P2_U5764 , P2_U5763 );
nand NAND2_4153 ( P2_U3458 , P2_U5766 , P2_U5765 );
nand NAND2_4154 ( P2_U3459 , P2_U5768 , P2_U5767 );
nand NAND2_4155 ( P2_U3460 , P2_U5771 , P2_U5770 );
nand NAND2_4156 ( P2_U3461 , P2_U5773 , P2_U5772 );
nand NAND2_4157 ( P2_U3462 , P2_U5775 , P2_U5774 );
nand NAND2_4158 ( P2_U3463 , P2_U5778 , P2_U5777 );
nand NAND2_4159 ( P2_U3464 , P2_U5780 , P2_U5779 );
nand NAND2_4160 ( P2_U3465 , P2_U5782 , P2_U5781 );
nand NAND2_4161 ( P2_U3466 , P2_U5785 , P2_U5784 );
nand NAND2_4162 ( P2_U3467 , P2_U5787 , P2_U5786 );
nand NAND2_4163 ( P2_U3468 , P2_U5789 , P2_U5788 );
nand NAND2_4164 ( P2_U3469 , P2_U5792 , P2_U5791 );
nand NAND2_4165 ( P2_U3470 , P2_U5794 , P2_U5793 );
nand NAND2_4166 ( P2_U3471 , P2_U5796 , P2_U5795 );
nand NAND2_4167 ( P2_U3472 , P2_U5799 , P2_U5798 );
nand NAND2_4168 ( P2_U3473 , P2_U5801 , P2_U5800 );
nand NAND2_4169 ( P2_U3474 , P2_U5803 , P2_U5802 );
nand NAND2_4170 ( P2_U3475 , P2_U5806 , P2_U5805 );
nand NAND2_4171 ( P2_U3476 , P2_U5808 , P2_U5807 );
nand NAND2_4172 ( P2_U3477 , P2_U5810 , P2_U5809 );
nand NAND2_4173 ( P2_U3478 , P2_U5813 , P2_U5812 );
nand NAND2_4174 ( P2_U3479 , P2_U5815 , P2_U5814 );
nand NAND2_4175 ( P2_U3480 , P2_U5817 , P2_U5816 );
nand NAND2_4176 ( P2_U3481 , P2_U5820 , P2_U5819 );
nand NAND2_4177 ( P2_U3482 , P2_U5822 , P2_U5821 );
nand NAND2_4178 ( P2_U3483 , P2_U5824 , P2_U5823 );
nand NAND2_4179 ( P2_U3484 , P2_U5827 , P2_U5826 );
nand NAND2_4180 ( P2_U3485 , P2_U5829 , P2_U5828 );
nand NAND2_4181 ( P2_U3486 , P2_U5832 , P2_U5831 );
nand NAND2_4182 ( P2_U3487 , P2_U5834 , P2_U5833 );
nand NAND2_4183 ( P2_U3488 , P2_U5836 , P2_U5835 );
nand NAND2_4184 ( P2_U3489 , P2_U5838 , P2_U5837 );
nand NAND2_4185 ( P2_U3490 , P2_U5840 , P2_U5839 );
nand NAND2_4186 ( P2_U3491 , P2_U5842 , P2_U5841 );
nand NAND2_4187 ( P2_U3492 , P2_U5844 , P2_U5843 );
nand NAND2_4188 ( P2_U3493 , P2_U5846 , P2_U5845 );
nand NAND2_4189 ( P2_U3494 , P2_U5848 , P2_U5847 );
nand NAND2_4190 ( P2_U3495 , P2_U5850 , P2_U5849 );
nand NAND2_4191 ( P2_U3496 , P2_U5852 , P2_U5851 );
nand NAND2_4192 ( P2_U3497 , P2_U5854 , P2_U5853 );
nand NAND2_4193 ( P2_U3498 , P2_U5856 , P2_U5855 );
nand NAND2_4194 ( P2_U3499 , P2_U5858 , P2_U5857 );
nand NAND2_4195 ( P2_U3500 , P2_U5860 , P2_U5859 );
nand NAND2_4196 ( P2_U3501 , P2_U5862 , P2_U5861 );
nand NAND2_4197 ( P2_U3502 , P2_U5864 , P2_U5863 );
nand NAND2_4198 ( P2_U3503 , P2_U5866 , P2_U5865 );
nand NAND2_4199 ( P2_U3504 , P2_U5868 , P2_U5867 );
nand NAND2_4200 ( P2_U3505 , P2_U5870 , P2_U5869 );
nand NAND2_4201 ( P2_U3506 , P2_U5872 , P2_U5871 );
nand NAND2_4202 ( P2_U3507 , P2_U5874 , P2_U5873 );
nand NAND2_4203 ( P2_U3508 , P2_U5876 , P2_U5875 );
nand NAND2_4204 ( P2_U3509 , P2_U5878 , P2_U5877 );
nand NAND2_4205 ( P2_U3510 , P2_U5880 , P2_U5879 );
nand NAND2_4206 ( P2_U3511 , P2_U5882 , P2_U5881 );
nand NAND2_4207 ( P2_U3512 , P2_U5884 , P2_U5883 );
nand NAND2_4208 ( P2_U3513 , P2_U5886 , P2_U5885 );
nand NAND2_4209 ( P2_U3514 , P2_U5888 , P2_U5887 );
nand NAND2_4210 ( P2_U3515 , P2_U5890 , P2_U5889 );
nand NAND2_4211 ( P2_U3516 , P2_U5892 , P2_U5891 );
nand NAND2_4212 ( P2_U3517 , P2_U5894 , P2_U5893 );
nand NAND2_4213 ( P2_U3518 , P2_U5896 , P2_U5895 );
nand NAND2_4214 ( P2_U3519 , P2_U5898 , P2_U5897 );
nand NAND2_4215 ( P2_U3520 , P2_U5900 , P2_U5899 );
nand NAND2_4216 ( P2_U3521 , P2_U5902 , P2_U5901 );
nand NAND2_4217 ( P2_U3522 , P2_U5904 , P2_U5903 );
nand NAND2_4218 ( P2_U3523 , P2_U5906 , P2_U5905 );
nand NAND2_4219 ( P2_U3524 , P2_U5908 , P2_U5907 );
nand NAND2_4220 ( P2_U3525 , P2_U5910 , P2_U5909 );
nand NAND2_4221 ( P2_U3526 , P2_U5912 , P2_U5911 );
nand NAND2_4222 ( P2_U3527 , P2_U5914 , P2_U5913 );
nand NAND2_4223 ( P2_U3528 , P2_U5916 , P2_U5915 );
nand NAND2_4224 ( P2_U3529 , P2_U5918 , P2_U5917 );
nand NAND2_4225 ( P2_U3530 , P2_U5920 , P2_U5919 );
nand NAND2_4226 ( P2_U3531 , P2_U5986 , P2_U5985 );
nand NAND2_4227 ( P2_U3532 , P2_U5988 , P2_U5987 );
nand NAND2_4228 ( P2_U3533 , P2_U5990 , P2_U5989 );
nand NAND2_4229 ( P2_U3534 , P2_U5992 , P2_U5991 );
nand NAND2_4230 ( P2_U3535 , P2_U5994 , P2_U5993 );
nand NAND2_4231 ( P2_U3536 , P2_U5996 , P2_U5995 );
nand NAND2_4232 ( P2_U3537 , P2_U5998 , P2_U5997 );
nand NAND2_4233 ( P2_U3538 , P2_U6000 , P2_U5999 );
nand NAND2_4234 ( P2_U3539 , P2_U6002 , P2_U6001 );
nand NAND2_4235 ( P2_U3540 , P2_U6004 , P2_U6003 );
nand NAND2_4236 ( P2_U3541 , P2_U6006 , P2_U6005 );
nand NAND2_4237 ( P2_U3542 , P2_U6008 , P2_U6007 );
nand NAND2_4238 ( P2_U3543 , P2_U6010 , P2_U6009 );
nand NAND2_4239 ( P2_U3544 , P2_U6012 , P2_U6011 );
nand NAND2_4240 ( P2_U3545 , P2_U6014 , P2_U6013 );
nand NAND2_4241 ( P2_U3546 , P2_U6016 , P2_U6015 );
nand NAND2_4242 ( P2_U3547 , P2_U6018 , P2_U6017 );
nand NAND2_4243 ( P2_U3548 , P2_U6020 , P2_U6019 );
nand NAND2_4244 ( P2_U3549 , P2_U6022 , P2_U6021 );
nand NAND2_4245 ( P2_U3550 , P2_U6024 , P2_U6023 );
nand NAND2_4246 ( P2_U3551 , P2_U6026 , P2_U6025 );
nand NAND2_4247 ( P2_U3552 , P2_U6028 , P2_U6027 );
nand NAND2_4248 ( P2_U3553 , P2_U6030 , P2_U6029 );
nand NAND2_4249 ( P2_U3554 , P2_U6032 , P2_U6031 );
nand NAND2_4250 ( P2_U3555 , P2_U6034 , P2_U6033 );
nand NAND2_4251 ( P2_U3556 , P2_U6036 , P2_U6035 );
nand NAND2_4252 ( P2_U3557 , P2_U6038 , P2_U6037 );
nand NAND2_4253 ( P2_U3558 , P2_U6040 , P2_U6039 );
nand NAND2_4254 ( P2_U3559 , P2_U6042 , P2_U6041 );
nand NAND2_4255 ( P2_U3560 , P2_U6044 , P2_U6043 );
nand NAND2_4256 ( P2_U3561 , P2_U6046 , P2_U6045 );
nand NAND2_4257 ( P2_U3562 , P2_U6048 , P2_U6047 );
and AND4_4258 ( P2_U3563 , P2_U4120 , P2_U4119 , P2_U4118 , P2_U4117 );
and AND2_4259 ( P2_U3564 , P2_U4122 , P2_U4121 );
and AND2_4260 ( P2_U3565 , P2_U4127 , P2_U4125 );
and AND4_4261 ( P2_U3566 , P2_U4082 , P2_U4081 , P2_U4080 , P2_U4079 );
and AND4_4262 ( P2_U3567 , P2_U4086 , P2_U4085 , P2_U4084 , P2_U4083 );
and AND4_4263 ( P2_U3568 , P2_U4090 , P2_U4089 , P2_U4088 , P2_U4087 );
and AND3_4264 ( P2_U3569 , P2_U4092 , P2_U4091 , P2_U4093 );
and AND4_4265 ( P2_U3570 , P2_U3569 , P2_U3568 , P2_U3567 , P2_U3566 );
and AND4_4266 ( P2_U3571 , P2_U4097 , P2_U4096 , P2_U4095 , P2_U4094 );
and AND4_4267 ( P2_U3572 , P2_U4101 , P2_U4100 , P2_U4099 , P2_U4098 );
and AND4_4268 ( P2_U3573 , P2_U4105 , P2_U4104 , P2_U4103 , P2_U4102 );
and AND3_4269 ( P2_U3574 , P2_U4107 , P2_U4106 , P2_U4108 );
and AND4_4270 ( P2_U3575 , P2_U3574 , P2_U3573 , P2_U3572 , P2_U3571 );
and AND2_4271 ( P2_U3576 , P2_U5696 , P2_U4110 );
and AND2_4272 ( P2_U3577 , P2_U5699 , P2_U3023 );
and AND2_4273 ( P2_U3578 , P2_U4143 , P2_U4142 );
and AND2_4274 ( P2_U3579 , P2_U4145 , P2_U4144 );
and AND3_4275 ( P2_U3580 , P2_U4147 , P2_U4146 , P2_U3579 );
and AND4_4276 ( P2_U3581 , P2_U4150 , P2_U4149 , P2_U4152 , P2_U4151 );
and AND2_4277 ( P2_U3582 , P2_U4162 , P2_U4161 );
and AND2_4278 ( P2_U3583 , P2_U4164 , P2_U4163 );
and AND3_4279 ( P2_U3584 , P2_U4166 , P2_U4165 , P2_U3583 );
and AND4_4280 ( P2_U3585 , P2_U4169 , P2_U4168 , P2_U4171 , P2_U4170 );
and AND2_4281 ( P2_U3586 , P2_U4181 , P2_U4180 );
and AND2_4282 ( P2_U3587 , P2_U4183 , P2_U4182 );
and AND3_4283 ( P2_U3588 , P2_U4185 , P2_U4184 , P2_U3587 );
and AND4_4284 ( P2_U3589 , P2_U4188 , P2_U4187 , P2_U4190 , P2_U4189 );
and AND2_4285 ( P2_U3590 , P2_U4200 , P2_U4199 );
and AND2_4286 ( P2_U3591 , P2_U4202 , P2_U4201 );
and AND3_4287 ( P2_U3592 , P2_U4204 , P2_U4203 , P2_U3591 );
and AND4_4288 ( P2_U3593 , P2_U4207 , P2_U4206 , P2_U4209 , P2_U4208 );
and AND2_4289 ( P2_U3594 , P2_U4219 , P2_U4218 );
and AND2_4290 ( P2_U3595 , P2_U4221 , P2_U4220 );
and AND3_4291 ( P2_U3596 , P2_U4223 , P2_U4222 , P2_U3595 );
and AND4_4292 ( P2_U3597 , P2_U4226 , P2_U4225 , P2_U4228 , P2_U4227 );
and AND2_4293 ( P2_U3598 , P2_U4238 , P2_U4237 );
and AND2_4294 ( P2_U3599 , P2_U4240 , P2_U4239 );
and AND3_4295 ( P2_U3600 , P2_U4242 , P2_U4241 , P2_U3599 );
and AND4_4296 ( P2_U3601 , P2_U4245 , P2_U4244 , P2_U4247 , P2_U4246 );
and AND2_4297 ( P2_U3602 , P2_U4257 , P2_U4256 );
and AND2_4298 ( P2_U3603 , P2_U4259 , P2_U4258 );
and AND3_4299 ( P2_U3604 , P2_U4261 , P2_U4260 , P2_U3603 );
and AND4_4300 ( P2_U3605 , P2_U4264 , P2_U4263 , P2_U4266 , P2_U4265 );
and AND2_4301 ( P2_U3606 , P2_U4276 , P2_U4275 );
and AND2_4302 ( P2_U3607 , P2_U4278 , P2_U4277 );
and AND3_4303 ( P2_U3608 , P2_U4280 , P2_U4279 , P2_U3607 );
and AND4_4304 ( P2_U3609 , P2_U4283 , P2_U4282 , P2_U4285 , P2_U4284 );
and AND2_4305 ( P2_U3610 , P2_U4295 , P2_U4294 );
and AND2_4306 ( P2_U3611 , P2_U4297 , P2_U4296 );
and AND3_4307 ( P2_U3612 , P2_U4299 , P2_U4298 , P2_U3611 );
and AND4_4308 ( P2_U3613 , P2_U4302 , P2_U4301 , P2_U4304 , P2_U4303 );
and AND2_4309 ( P2_U3614 , P2_U4314 , P2_U4313 );
and AND2_4310 ( P2_U3615 , P2_U4316 , P2_U4315 );
and AND3_4311 ( P2_U3616 , P2_U4318 , P2_U4317 , P2_U3615 );
and AND4_4312 ( P2_U3617 , P2_U4321 , P2_U4320 , P2_U4323 , P2_U4322 );
and AND2_4313 ( P2_U3618 , P2_U4333 , P2_U4332 );
and AND2_4314 ( P2_U3619 , P2_U4335 , P2_U4334 );
and AND3_4315 ( P2_U3620 , P2_U4337 , P2_U4336 , P2_U3619 );
and AND4_4316 ( P2_U3621 , P2_U4340 , P2_U4339 , P2_U4342 , P2_U4341 );
and AND2_4317 ( P2_U3622 , P2_U4352 , P2_U4351 );
and AND2_4318 ( P2_U3623 , P2_U4354 , P2_U4353 );
and AND3_4319 ( P2_U3624 , P2_U4356 , P2_U4355 , P2_U3623 );
and AND4_4320 ( P2_U3625 , P2_U4359 , P2_U4358 , P2_U4361 , P2_U4360 );
and AND2_4321 ( P2_U3626 , P2_U4371 , P2_U4370 );
and AND2_4322 ( P2_U3627 , P2_U4373 , P2_U4372 );
and AND3_4323 ( P2_U3628 , P2_U4375 , P2_U4374 , P2_U3627 );
and AND4_4324 ( P2_U3629 , P2_U4378 , P2_U4377 , P2_U4380 , P2_U4379 );
and AND2_4325 ( P2_U3630 , P2_U4390 , P2_U4389 );
and AND2_4326 ( P2_U3631 , P2_U4392 , P2_U4391 );
and AND3_4327 ( P2_U3632 , P2_U4394 , P2_U4393 , P2_U3631 );
and AND4_4328 ( P2_U3633 , P2_U4397 , P2_U4396 , P2_U4399 , P2_U4398 );
and AND2_4329 ( P2_U3634 , P2_U4409 , P2_U4408 );
and AND2_4330 ( P2_U3635 , P2_U4411 , P2_U4410 );
and AND3_4331 ( P2_U3636 , P2_U4413 , P2_U4412 , P2_U3635 );
and AND4_4332 ( P2_U3637 , P2_U4416 , P2_U4415 , P2_U4418 , P2_U4417 );
and AND2_4333 ( P2_U3638 , P2_U4428 , P2_U4427 );
and AND2_4334 ( P2_U3639 , P2_U4430 , P2_U4429 );
and AND3_4335 ( P2_U3640 , P2_U4432 , P2_U4431 , P2_U3639 );
and AND4_4336 ( P2_U3641 , P2_U4435 , P2_U4434 , P2_U4437 , P2_U4436 );
and AND2_4337 ( P2_U3642 , P2_U4447 , P2_U4446 );
and AND2_4338 ( P2_U3643 , P2_U4449 , P2_U4448 );
and AND3_4339 ( P2_U3644 , P2_U4451 , P2_U4450 , P2_U3643 );
and AND4_4340 ( P2_U3645 , P2_U4454 , P2_U4453 , P2_U4456 , P2_U4455 );
and AND2_4341 ( P2_U3646 , P2_U4466 , P2_U4465 );
and AND2_4342 ( P2_U3647 , P2_U4468 , P2_U4467 );
and AND3_4343 ( P2_U3648 , P2_U4470 , P2_U4469 , P2_U3647 );
and AND4_4344 ( P2_U3649 , P2_U4473 , P2_U4472 , P2_U4475 , P2_U4474 );
and AND2_4345 ( P2_U3650 , P2_U4485 , P2_U4484 );
and AND2_4346 ( P2_U3651 , P2_U4487 , P2_U4486 );
and AND3_4347 ( P2_U3652 , P2_U4489 , P2_U4488 , P2_U3651 );
and AND4_4348 ( P2_U3653 , P2_U4492 , P2_U4491 , P2_U4494 , P2_U4493 );
and AND2_4349 ( P2_U3654 , P2_U4504 , P2_U4503 );
and AND2_4350 ( P2_U3655 , P2_U4506 , P2_U4505 );
and AND3_4351 ( P2_U3656 , P2_U4508 , P2_U4507 , P2_U3655 );
and AND4_4352 ( P2_U3657 , P2_U4511 , P2_U4510 , P2_U4513 , P2_U4512 );
and AND2_4353 ( P2_U3658 , P2_U4523 , P2_U4522 );
and AND2_4354 ( P2_U3659 , P2_U4525 , P2_U4524 );
and AND3_4355 ( P2_U3660 , P2_U4527 , P2_U4526 , P2_U3659 );
and AND4_4356 ( P2_U3661 , P2_U4530 , P2_U4529 , P2_U4532 , P2_U4531 );
and AND2_4357 ( P2_U3662 , P2_U4542 , P2_U4541 );
and AND2_4358 ( P2_U3663 , P2_U4544 , P2_U4543 );
and AND3_4359 ( P2_U3664 , P2_U4546 , P2_U4545 , P2_U3663 );
and AND4_4360 ( P2_U3665 , P2_U4549 , P2_U4548 , P2_U4551 , P2_U4550 );
and AND2_4361 ( P2_U3666 , P2_U4561 , P2_U4560 );
and AND2_4362 ( P2_U3667 , P2_U4563 , P2_U4562 );
and AND3_4363 ( P2_U3668 , P2_U4565 , P2_U4564 , P2_U3667 );
and AND4_4364 ( P2_U3669 , P2_U4568 , P2_U4567 , P2_U4570 , P2_U4569 );
and AND2_4365 ( P2_U3670 , P2_U4580 , P2_U4579 );
and AND2_4366 ( P2_U3671 , P2_U4582 , P2_U4581 );
and AND3_4367 ( P2_U3672 , P2_U4584 , P2_U4583 , P2_U3671 );
and AND4_4368 ( P2_U3673 , P2_U4587 , P2_U4586 , P2_U4589 , P2_U4588 );
and AND2_4369 ( P2_U3674 , P2_U4599 , P2_U4598 );
and AND2_4370 ( P2_U3675 , P2_U4601 , P2_U4600 );
and AND3_4371 ( P2_U3676 , P2_U4603 , P2_U4602 , P2_U3675 );
and AND4_4372 ( P2_U3677 , P2_U4606 , P2_U4605 , P2_U4608 , P2_U4607 );
and AND2_4373 ( P2_U3678 , P2_U4618 , P2_U4617 );
and AND2_4374 ( P2_U3679 , P2_U4620 , P2_U4619 );
and AND3_4375 ( P2_U3680 , P2_U4622 , P2_U4621 , P2_U3679 );
and AND4_4376 ( P2_U3681 , P2_U4625 , P2_U4624 , P2_U4627 , P2_U4626 );
and AND2_4377 ( P2_U3682 , P2_U4637 , P2_U4636 );
and AND2_4378 ( P2_U3683 , P2_U4639 , P2_U4638 );
and AND3_4379 ( P2_U3684 , P2_U4641 , P2_U4640 , P2_U3683 );
and AND4_4380 ( P2_U3685 , P2_U4644 , P2_U4643 , P2_U4646 , P2_U4645 );
and AND2_4381 ( P2_U3686 , P2_U4658 , P2_U4657 );
and AND3_4382 ( P2_U3687 , P2_U4660 , P2_U4659 , P2_U3686 );
and AND4_4383 ( P2_U3688 , P2_U4663 , P2_U4662 , P2_U4665 , P2_U4664 );
and AND2_4384 ( P2_U3689 , P2_U4672 , P2_U3963 );
and AND2_4385 ( P2_U3690 , P2_U4677 , P2_U4676 );
and AND2_4386 ( P2_U3691 , P2_U4679 , P2_U4678 );
and AND3_4387 ( P2_U3692 , P2_U4681 , P2_U4680 , P2_U3691 );
and AND3_4388 ( P2_U3693 , P2_U4685 , P2_U4683 , P2_U4684 );
and AND2_4389 ( P2_U3694 , P2_U3963 , P2_U4672 );
and AND2_4390 ( P2_U3695 , P2_U3023 , P2_U3428 );
and AND3_4391 ( P2_U3696 , P2_U5699 , P2_U3935 , P2_U3429 );
and AND3_4392 ( P2_U3697 , P2_U4702 , P2_U4701 , P2_U4703 );
and AND3_4393 ( P2_U3698 , P2_U4705 , P2_U4704 , P2_U3883 );
and AND3_4394 ( P2_U3699 , P2_U4707 , P2_U4706 , P2_U4708 );
and AND3_4395 ( P2_U3700 , P2_U4710 , P2_U4709 , P2_U3884 );
and AND3_4396 ( P2_U3701 , P2_U4712 , P2_U4711 , P2_U4713 );
and AND3_4397 ( P2_U3702 , P2_U4715 , P2_U4714 , P2_U3885 );
and AND3_4398 ( P2_U3703 , P2_U4717 , P2_U4716 , P2_U4718 );
and AND3_4399 ( P2_U3704 , P2_U4720 , P2_U4719 , P2_U3886 );
and AND3_4400 ( P2_U3705 , P2_U4722 , P2_U4721 , P2_U4723 );
and AND3_4401 ( P2_U3706 , P2_U4725 , P2_U4724 , P2_U3887 );
and AND3_4402 ( P2_U3707 , P2_U4727 , P2_U4726 , P2_U4728 );
and AND3_4403 ( P2_U3708 , P2_U4730 , P2_U4729 , P2_U3888 );
and AND3_4404 ( P2_U3709 , P2_U4732 , P2_U4731 , P2_U4733 );
and AND3_4405 ( P2_U3710 , P2_U4735 , P2_U4734 , P2_U3889 );
and AND3_4406 ( P2_U3711 , P2_U4737 , P2_U4736 , P2_U4738 );
and AND3_4407 ( P2_U3712 , P2_U4740 , P2_U4739 , P2_U3890 );
and AND3_4408 ( P2_U3713 , P2_U4742 , P2_U4741 , P2_U4743 );
and AND3_4409 ( P2_U3714 , P2_U4745 , P2_U4744 , P2_U3891 );
and AND3_4410 ( P2_U3715 , P2_U4747 , P2_U4746 , P2_U4748 );
and AND3_4411 ( P2_U3716 , P2_U4750 , P2_U4749 , P2_U3892 );
and AND3_4412 ( P2_U3717 , P2_U4752 , P2_U4751 , P2_U4753 );
and AND2_4413 ( P2_U3718 , P2_U4755 , P2_U4754 );
and AND3_4414 ( P2_U3719 , P2_U4757 , P2_U4756 , P2_U4758 );
and AND2_4415 ( P2_U3720 , P2_U4760 , P2_U4759 );
and AND3_4416 ( P2_U3721 , P2_U4762 , P2_U4761 , P2_U4763 );
and AND2_4417 ( P2_U3722 , P2_U4765 , P2_U4764 );
and AND3_4418 ( P2_U3723 , P2_U4768 , P2_U4766 , P2_U4767 );
and AND2_4419 ( P2_U3724 , P2_U4770 , P2_U4769 );
and AND3_4420 ( P2_U3725 , P2_U4772 , P2_U4771 , P2_U4773 );
and AND2_4421 ( P2_U3726 , P2_U4775 , P2_U4774 );
and AND3_4422 ( P2_U3727 , P2_U4778 , P2_U4776 , P2_U4777 );
and AND2_4423 ( P2_U3728 , P2_U4780 , P2_U4779 );
and AND2_4424 ( P2_U3729 , P2_U4783 , P2_U4781 );
and AND2_4425 ( P2_U3730 , P2_U4785 , P2_U4784 );
and AND2_4426 ( P2_U3731 , P2_U4788 , P2_U4786 );
and AND2_4427 ( P2_U3732 , P2_U4790 , P2_U4789 );
and AND2_4428 ( P2_U3733 , P2_U4793 , P2_U4791 );
and AND2_4429 ( P2_U3734 , P2_U4795 , P2_U4794 );
and AND2_4430 ( P2_U3735 , P2_U4798 , P2_U4796 );
and AND2_4431 ( P2_U3736 , P2_U4800 , P2_U4799 );
and AND2_4432 ( P2_U3737 , P2_U4803 , P2_U4801 );
and AND2_4433 ( P2_U3738 , P2_U4805 , P2_U4804 );
and AND2_4434 ( P2_U3739 , P2_U4808 , P2_U4806 );
and AND2_4435 ( P2_U3740 , P2_U4810 , P2_U4809 );
and AND2_4436 ( P2_U3741 , P2_U4813 , P2_U4811 );
and AND2_4437 ( P2_U3742 , P2_U4815 , P2_U4814 );
and AND2_4438 ( P2_U3743 , P2_U4818 , P2_U4816 );
and AND2_4439 ( P2_U3744 , P2_U4820 , P2_U4819 );
and AND2_4440 ( P2_U3745 , P2_U4823 , P2_U4821 );
and AND2_4441 ( P2_U3746 , P2_U4825 , P2_U4824 );
and AND2_4442 ( P2_U3747 , P2_U4828 , P2_U4826 );
and AND2_4443 ( P2_U3748 , P2_U4830 , P2_U4829 );
and AND2_4444 ( P2_U3749 , P2_U4833 , P2_U4831 );
and AND2_4445 ( P2_U3750 , P2_U4835 , P2_U4834 );
and AND2_4446 ( P2_U3751 , P2_U4838 , P2_U4836 );
and AND2_4447 ( P2_U3752 , P2_U4840 , P2_U4839 );
and AND2_4448 ( P2_U3753 , P2_U4843 , P2_U4841 );
and AND2_4449 ( P2_U3754 , P2_U4845 , P2_U4844 );
and AND3_4450 ( P2_U3755 , P2_U3335 , P2_U3336 , P2_U3334 );
and AND2_4451 ( P2_U3756 , P2_U5643 , P2_U3397 );
and AND2_4452 ( P2_U3757 , P2_U3415 , P2_STATE_REG );
and AND5_4453 ( P2_U3758 , P2_U4870 , P2_U4868 , P2_U4869 , P2_U4867 , P2_U4866 );
and AND5_4454 ( P2_U3759 , P2_U4885 , P2_U4883 , P2_U4884 , P2_U4882 , P2_U4881 );
and AND5_4455 ( P2_U3760 , P2_U4900 , P2_U4898 , P2_U4899 , P2_U4897 , P2_U4896 );
and AND5_4456 ( P2_U3761 , P2_U4915 , P2_U4913 , P2_U4914 , P2_U4912 , P2_U4911 );
and AND5_4457 ( P2_U3762 , P2_U4930 , P2_U4928 , P2_U4929 , P2_U4927 , P2_U4926 );
and AND5_4458 ( P2_U3763 , P2_U4945 , P2_U4943 , P2_U4944 , P2_U4942 , P2_U4941 );
and AND5_4459 ( P2_U3764 , P2_U4960 , P2_U4958 , P2_U4959 , P2_U4957 , P2_U4956 );
and AND5_4460 ( P2_U3765 , P2_U4975 , P2_U4973 , P2_U4974 , P2_U4972 , P2_U4971 );
and AND5_4461 ( P2_U3766 , P2_U4989 , P2_U4988 , P2_U4990 , P2_U4987 , P2_U4986 );
and AND5_4462 ( P2_U3767 , P2_U5005 , P2_U5003 , P2_U5004 , P2_U5002 , P2_U5001 );
and AND5_4463 ( P2_U3768 , P2_U5019 , P2_U5018 , P2_U5020 , P2_U5017 , P2_U5016 );
and AND2_4464 ( P2_U3769 , P2_U5032 , P2_U5031 );
and AND3_4465 ( P2_U3770 , P2_U5034 , P2_U5033 , P2_U5035 );
and AND2_4466 ( P2_U3771 , P2_U5047 , P2_U5046 );
and AND3_4467 ( P2_U3772 , P2_U5049 , P2_U5048 , P2_U5050 );
and AND2_4468 ( P2_U3773 , P2_U5062 , P2_U5061 );
and AND3_4469 ( P2_U3774 , P2_U5064 , P2_U5063 , P2_U5065 );
and AND2_4470 ( P2_U3775 , P2_U5077 , P2_U5076 );
and AND3_4471 ( P2_U3776 , P2_U5079 , P2_U5078 , P2_U5080 );
and AND2_4472 ( P2_U3777 , P2_U5092 , P2_U5091 );
and AND3_4473 ( P2_U3778 , P2_U5094 , P2_U5093 , P2_U5095 );
and AND2_4474 ( P2_U3779 , P2_U5107 , P2_U5106 );
and AND3_4475 ( P2_U3780 , P2_U5109 , P2_U5108 , P2_U5110 );
and AND2_4476 ( P2_U3781 , P2_U5122 , P2_U5121 );
and AND3_4477 ( P2_U3782 , P2_U5124 , P2_U5123 , P2_U5125 );
and AND2_4478 ( P2_U3783 , P2_U5137 , P2_U5136 );
and AND3_4479 ( P2_U3784 , P2_U5139 , P2_U5138 , P2_U5140 );
and AND2_4480 ( P2_U3785 , P2_U5152 , P2_U5151 );
and AND3_4481 ( P2_U3786 , P2_U5154 , P2_U5153 , P2_U5155 );
and AND2_4482 ( P2_U3787 , P2_U5639 , P2_U5658 );
and AND3_4483 ( P2_U3788 , P2_U6103 , P2_U6100 , P2_U6106 );
and AND4_4484 ( P2_U3789 , P2_U6097 , P2_U6094 , P2_U6091 , P2_U6088 );
and AND4_4485 ( P2_U3790 , P2_U6121 , P2_U6118 , P2_U6115 , P2_U6112 );
and AND4_4486 ( P2_U3791 , P2_U6127 , P2_U6124 , P2_U6130 , P2_U6133 );
and AND5_4487 ( P2_U3792 , P2_U3788 , P2_U3789 , P2_U6109 , P2_U3791 , P2_U3790 );
and AND5_4488 ( P2_U3793 , P2_U3796 , P2_U3795 , P2_U6061 , P2_U6058 , P2_U6055 );
and AND5_4489 ( P2_U3794 , P2_U6145 , P2_U6142 , P2_U6139 , P2_U6136 , P2_U6148 );
and AND4_4490 ( P2_U3795 , P2_U6073 , P2_U6070 , P2_U6067 , P2_U6064 );
and AND2_4491 ( P2_U3796 , P2_U6079 , P2_U6076 );
and AND2_4492 ( P2_U3797 , P2_U5640 , P2_U5631 );
and AND2_4493 ( P2_U3798 , P2_U3428 , P2_U3429 );
and AND2_4494 ( P2_U3799 , P2_U3339 , P2_U3928 );
and AND2_4495 ( P2_U3800 , P2_U3799 , P2_U3342 );
and AND2_4496 ( P2_U3801 , P2_U3395 , P2_U3410 );
and AND3_4497 ( P2_U3802 , P2_U5658 , P2_U3935 , P2_U3399 );
and AND2_4498 ( P2_U3803 , P2_U3023 , P2_U5171 );
and AND2_4499 ( P2_U3804 , P2_U5198 , P2_U5196 );
and AND2_4500 ( P2_U3805 , P2_U5216 , P2_U5214 );
and AND2_4501 ( P2_U3806 , P2_U3969 , P2_U3080 );
and AND2_4502 ( P2_U3807 , P2_U5259 , P2_U5258 );
and AND2_4503 ( P2_U3808 , P2_U5262 , P2_U5261 );
and AND2_4504 ( P2_U3809 , P2_U5278 , P2_U5276 );
and AND2_4505 ( P2_U3810 , P2_U5305 , P2_U5303 );
and AND2_4506 ( P2_U3811 , P2_U5350 , P2_U5348 );
and AND2_4507 ( P2_U3812 , P2_U5359 , P2_U5357 );
and AND2_4508 ( P2_U3813 , P2_U5386 , P2_U5384 );
and AND2_4509 ( P2_U3814 , P2_U5431 , P2_U5429 );
and AND2_4510 ( P2_U3815 , P2_U5435 , P2_STATE_REG );
and AND3_4511 ( P2_U3816 , P2_U3919 , P2_U3936 , P2_U3920 );
and AND2_4512 ( P2_U3817 , P2_U5671 , P2_U3419 );
and AND2_4513 ( P2_U3818 , P2_U3394 , P2_U3339 );
and AND3_4514 ( P2_U3819 , P2_U3342 , P2_U3390 , P2_U3818 );
and AND2_4515 ( P2_U3820 , P2_U3334 , P2_U3928 );
and AND2_4516 ( P2_U3821 , P2_U3415 , P2_U5444 );
and AND2_4517 ( P2_U3822 , P2_U3415 , P2_U5447 );
and AND2_4518 ( P2_U3823 , P2_U3415 , P2_U5450 );
and AND2_4519 ( P2_U3824 , P2_U3415 , P2_U5453 );
and AND2_4520 ( P2_U3825 , P2_U3415 , P2_U5456 );
and AND2_4521 ( P2_U3826 , P2_U3827 , P2_U5457 );
and AND2_4522 ( P2_U3827 , P2_U3415 , P2_U5459 );
and AND2_4523 ( P2_U3828 , P2_U5460 , P2_U3410 );
and AND2_4524 ( P2_U3829 , P2_U3830 , P2_U5465 );
and AND2_4525 ( P2_U3830 , P2_U3415 , P2_U5467 );
and AND2_4526 ( P2_U3831 , P2_U3415 , P2_U5468 );
and AND2_4527 ( P2_U3832 , P2_U3415 , P2_U5471 );
and AND2_4528 ( P2_U3833 , P2_U3415 , P2_U5474 );
and AND2_4529 ( P2_U3834 , P2_U3415 , P2_U5477 );
and AND2_4530 ( P2_U3835 , P2_U3415 , P2_U5480 );
and AND2_4531 ( P2_U3836 , P2_U3415 , P2_U5483 );
and AND2_4532 ( P2_U3837 , P2_U3415 , P2_U5486 );
and AND2_4533 ( P2_U3838 , P2_U3415 , P2_U5489 );
and AND2_4534 ( P2_U3839 , P2_U3415 , P2_U5492 );
and AND2_4535 ( P2_U3840 , P2_U3415 , P2_U5495 );
and AND2_4536 ( P2_U3841 , P2_U3842 , P2_U5498 );
and AND2_4537 ( P2_U3842 , P2_U3415 , P2_U5500 );
and AND2_4538 ( P2_U3843 , P2_U3415 , P2_U5501 );
and AND2_4539 ( P2_U3844 , P2_U3415 , P2_U5504 );
and AND2_4540 ( P2_U3845 , P2_U3415 , P2_U5507 );
and AND2_4541 ( P2_U3846 , P2_U3415 , P2_U5510 );
and AND2_4542 ( P2_U3847 , P2_U3415 , P2_U5513 );
and AND2_4543 ( P2_U3848 , P2_U3415 , P2_U5516 );
and AND2_4544 ( P2_U3849 , P2_U3415 , P2_U5519 );
and AND2_4545 ( P2_U3850 , P2_U3415 , P2_U5522 );
and AND2_4546 ( P2_U3851 , P2_U3415 , P2_U5527 );
and AND2_4547 ( P2_U3852 , P2_U3415 , P2_U5530 );
and AND2_4548 ( P2_U3853 , P2_U3854 , P2_U5531 );
and AND2_4549 ( P2_U3854 , P2_U3415 , P2_U5533 );
and AND2_4550 ( P2_U3855 , P2_U3856 , P2_U5534 );
and AND2_4551 ( P2_U3856 , P2_U3415 , P2_U5536 );
and AND2_4552 ( P2_U3857 , P2_U5539 , P2_U5540 );
and AND2_4553 ( P2_U3858 , P2_U5542 , P2_U5543 );
and AND2_4554 ( P2_U3859 , P2_U5564 , P2_U5565 );
and AND2_4555 ( P2_U3860 , P2_U5567 , P2_U5568 );
and AND2_4556 ( P2_U3861 , P2_U5570 , P2_U5571 );
and AND2_4557 ( P2_U3862 , P2_U5573 , P2_U5574 );
and AND2_4558 ( P2_U3863 , P2_U5576 , P2_U5577 );
and AND2_4559 ( P2_U3864 , P2_U5579 , P2_U5580 );
and AND2_4560 ( P2_U3865 , P2_U5582 , P2_U5583 );
and AND2_4561 ( P2_U3866 , P2_U5585 , P2_U5586 );
and AND2_4562 ( P2_U3867 , P2_U5588 , P2_U5589 );
and AND2_4563 ( P2_U3868 , P2_U5591 , P2_U5592 );
and AND2_4564 ( P2_U3869 , P2_U5597 , P2_U5598 );
and AND2_4565 ( P2_U3870 , P2_U5600 , P2_U5601 );
and AND2_4566 ( P2_U3871 , P2_U5603 , P2_U5604 );
and AND2_4567 ( P2_U3872 , P2_U5606 , P2_U5607 );
and AND2_4568 ( P2_U3873 , P2_U5609 , P2_U5610 );
and AND2_4569 ( P2_U3874 , P2_U5612 , P2_U5613 );
and AND2_4570 ( P2_U3875 , P2_U5615 , P2_U5616 );
and AND2_4571 ( P2_U3876 , P2_U5618 , P2_U5619 );
and AND2_4572 ( P2_U3877 , P2_U5621 , P2_U5622 );
and AND2_4573 ( P2_U3878 , P2_U5624 , P2_U5625 );
not NOT1_4574 ( P2_U3879 , P2_IR_REG_31_ );
nand NAND2_4575 ( P2_U3880 , P2_U3023 , P2_U3333 );
nand NAND2_4576 ( P2_U3881 , P2_U3577 , P2_U3050 );
nand NAND2_4577 ( P2_U3882 , P2_U3695 , P2_U3050 );
and AND2_4578 ( P2_U3883 , P2_U5922 , P2_U5921 );
and AND2_4579 ( P2_U3884 , P2_U5924 , P2_U5923 );
and AND2_4580 ( P2_U3885 , P2_U5926 , P2_U5925 );
and AND2_4581 ( P2_U3886 , P2_U5928 , P2_U5927 );
and AND2_4582 ( P2_U3887 , P2_U5930 , P2_U5929 );
and AND2_4583 ( P2_U3888 , P2_U5932 , P2_U5931 );
and AND2_4584 ( P2_U3889 , P2_U5934 , P2_U5933 );
and AND2_4585 ( P2_U3890 , P2_U5936 , P2_U5935 );
and AND2_4586 ( P2_U3891 , P2_U5938 , P2_U5937 );
and AND2_4587 ( P2_U3892 , P2_U5940 , P2_U5939 );
and AND2_4588 ( P2_U3893 , P2_U5942 , P2_U5941 );
and AND2_4589 ( P2_U3894 , P2_U5944 , P2_U5943 );
and AND2_4590 ( P2_U3895 , P2_U5946 , P2_U5945 );
and AND2_4591 ( P2_U3896 , P2_U5948 , P2_U5947 );
and AND2_4592 ( P2_U3897 , P2_U5950 , P2_U5949 );
and AND2_4593 ( P2_U3898 , P2_U5952 , P2_U5951 );
and AND2_4594 ( P2_U3899 , P2_U5954 , P2_U5953 );
and AND2_4595 ( P2_U3900 , P2_U5956 , P2_U5955 );
and AND2_4596 ( P2_U3901 , P2_U5958 , P2_U5957 );
and AND2_4597 ( P2_U3902 , P2_U5960 , P2_U5959 );
and AND2_4598 ( P2_U3903 , P2_U5962 , P2_U5961 );
and AND2_4599 ( P2_U3904 , P2_U5964 , P2_U5963 );
and AND2_4600 ( P2_U3905 , P2_U5966 , P2_U5965 );
and AND2_4601 ( P2_U3906 , P2_U5968 , P2_U5967 );
and AND2_4602 ( P2_U3907 , P2_U5970 , P2_U5969 );
and AND2_4603 ( P2_U3908 , P2_U5972 , P2_U5971 );
and AND2_4604 ( P2_U3909 , P2_U5974 , P2_U5973 );
and AND2_4605 ( P2_U3910 , P2_U5976 , P2_U5975 );
and AND2_4606 ( P2_U3911 , P2_U5978 , P2_U5977 );
and AND2_4607 ( P2_U3912 , P2_U5980 , P2_U5979 );
nand NAND2_4608 ( P2_U3913 , P2_U3694 , P2_U3058 );
and AND2_4609 ( P2_U3914 , P2_U5982 , P2_U5981 );
and AND2_4610 ( P2_U3915 , P2_U5984 , P2_U5983 );
not NOT1_4611 ( P2_U3916 , P2_R1312_U18 );
and AND2_4612 ( P2_U3917 , P2_U6050 , P2_U6049 );
nand NAND5_4613 ( P2_U3918 , P2_U3794 , P2_U3792 , P2_U6085 , P2_U6082 , P2_U3793 );
nand NAND2_4614 ( P2_U3919 , P2_U3049 , P2_U5674 );
nand NAND2_4615 ( P2_U3920 , P2_U3973 , P2_U3418 );
not NOT1_4616 ( P2_U3921 , P2_U3390 );
not NOT1_4617 ( P2_U3922 , P2_U3342 );
nand NAND2_4618 ( P2_U3923 , P2_U3976 , P2_U3418 );
not NOT1_4619 ( P2_U3924 , P2_U3339 );
not NOT1_4620 ( P2_U3925 , P2_U3346 );
not NOT1_4621 ( P2_U3926 , P2_U3336 );
not NOT1_4622 ( P2_U3927 , P2_U3394 );
nand NAND2_4623 ( P2_U3928 , P2_U3973 , P2_U3420 );
not NOT1_4624 ( P2_U3929 , P2_U3410 );
not NOT1_4625 ( P2_U3930 , P2_U3335 );
not NOT1_4626 ( P2_U3931 , P2_U3334 );
not NOT1_4627 ( P2_U3932 , P2_U3395 );
not NOT1_4628 ( P2_U3933 , P2_U3393 );
nand NAND2_4629 ( P2_U3934 , P2_U3925 , P2_U5674 );
nand NAND2_4630 ( P2_U3935 , P2_U3963 , P2_U3340 );
nand NAND2_4631 ( P2_U3936 , P2_U3973 , P2_U5671 );
not NOT1_4632 ( P2_U3937 , P2_U3402 );
not NOT1_4633 ( P2_U3938 , P2_U3392 );
not NOT1_4634 ( P2_U3939 , P2_U3341 );
not NOT1_4635 ( P2_U3940 , P2_U3919 );
not NOT1_4636 ( P2_U3941 , P2_U3337 );
not NOT1_4637 ( P2_U3942 , P2_U3920 );
not NOT1_4638 ( P2_U3943 , P2_U3338 );
not NOT1_4639 ( P2_U3944 , P2_U3343 );
not NOT1_4640 ( P2_U3945 , P2_U3347 );
not NOT1_4641 ( P2_U3946 , P2_U3406 );
not NOT1_4642 ( P2_U3947 , P2_U3400 );
not NOT1_4643 ( P2_U3948 , P2_U3397 );
not NOT1_4644 ( P2_U3949 , P2_U3384 );
not NOT1_4645 ( P2_U3950 , P2_U3382 );
not NOT1_4646 ( P2_U3951 , P2_U3380 );
not NOT1_4647 ( P2_U3952 , P2_U3378 );
not NOT1_4648 ( P2_U3953 , P2_U3376 );
not NOT1_4649 ( P2_U3954 , P2_U3374 );
not NOT1_4650 ( P2_U3955 , P2_U3372 );
not NOT1_4651 ( P2_U3956 , P2_U3370 );
not NOT1_4652 ( P2_U3957 , P2_U3368 );
not NOT1_4653 ( P2_U3958 , P2_U3389 );
not NOT1_4654 ( P2_U3959 , P2_U3388 );
not NOT1_4655 ( P2_U3960 , P2_U3386 );
not NOT1_4656 ( P2_U3961 , P2_U3403 );
not NOT1_4657 ( P2_U3962 , P2_U3396 );
not NOT1_4658 ( P2_U3963 , P2_U3344 );
not NOT1_4659 ( P2_U3964 , P2_U3391 );
not NOT1_4660 ( P2_U3965 , P2_U3882 );
not NOT1_4661 ( P2_U3966 , P2_U3881 );
not NOT1_4662 ( P2_U3967 , P2_U3880 );
not NOT1_4663 ( P2_U3968 , P2_U3913 );
not NOT1_4664 ( P2_U3969 , P2_U3407 );
nand NAND2_4665 ( P2_U3970 , P2_U3408 , P2_STATE_REG );
nand NAND2_4666 ( P2_U3971 , P2_U3933 , P2_U3023 );
not NOT1_4667 ( P2_U3972 , P2_U3405 );
not NOT1_4668 ( P2_U3973 , P2_U3404 );
not NOT1_4669 ( P2_U3974 , P2_U3340 );
not NOT1_4670 ( P2_U3975 , P2_U3332 );
not NOT1_4671 ( P2_U3976 , P2_U3345 );
not NOT1_4672 ( P2_U3977 , P2_U3399 );
not NOT1_4673 ( P2_U3978 , P2_U3329 );
nand NAND2_4674 ( P2_U3979 , U93 , P2_U3088 );
nand NAND2_4675 ( P2_U3980 , P2_IR_REG_0_ , P2_U3030 );
nand NAND2_4676 ( P2_U3981 , P2_IR_REG_0_ , P2_U3978 );
nand NAND2_4677 ( P2_U3982 , U82 , P2_U3088 );
nand NAND2_4678 ( P2_U3983 , P2_SUB_1108_U42 , P2_U3030 );
nand NAND2_4679 ( P2_U3984 , P2_IR_REG_1_ , P2_U3978 );
nand NAND2_4680 ( P2_U3985 , U71 , P2_U3088 );
nand NAND2_4681 ( P2_U3986 , P2_SUB_1108_U17 , P2_U3030 );
nand NAND2_4682 ( P2_U3987 , P2_IR_REG_2_ , P2_U3978 );
nand NAND2_4683 ( P2_U3988 , U68 , P2_U3088 );
nand NAND2_4684 ( P2_U3989 , P2_SUB_1108_U18 , P2_U3030 );
nand NAND2_4685 ( P2_U3990 , P2_IR_REG_3_ , P2_U3978 );
nand NAND2_4686 ( P2_U3991 , U67 , P2_U3088 );
nand NAND2_4687 ( P2_U3992 , P2_SUB_1108_U19 , P2_U3030 );
nand NAND2_4688 ( P2_U3993 , P2_IR_REG_4_ , P2_U3978 );
nand NAND2_4689 ( P2_U3994 , U66 , P2_U3088 );
nand NAND2_4690 ( P2_U3995 , P2_SUB_1108_U101 , P2_U3030 );
nand NAND2_4691 ( P2_U3996 , P2_IR_REG_5_ , P2_U3978 );
nand NAND2_4692 ( P2_U3997 , U65 , P2_U3088 );
nand NAND2_4693 ( P2_U3998 , P2_SUB_1108_U20 , P2_U3030 );
nand NAND2_4694 ( P2_U3999 , P2_IR_REG_6_ , P2_U3978 );
nand NAND2_4695 ( P2_U4000 , U64 , P2_U3088 );
nand NAND2_4696 ( P2_U4001 , P2_SUB_1108_U21 , P2_U3030 );
nand NAND2_4697 ( P2_U4002 , P2_IR_REG_7_ , P2_U3978 );
nand NAND2_4698 ( P2_U4003 , U63 , P2_U3088 );
nand NAND2_4699 ( P2_U4004 , P2_SUB_1108_U22 , P2_U3030 );
nand NAND2_4700 ( P2_U4005 , P2_IR_REG_8_ , P2_U3978 );
nand NAND2_4701 ( P2_U4006 , U62 , P2_U3088 );
nand NAND2_4702 ( P2_U4007 , P2_SUB_1108_U99 , P2_U3030 );
nand NAND2_4703 ( P2_U4008 , P2_IR_REG_9_ , P2_U3978 );
nand NAND2_4704 ( P2_U4009 , U92 , P2_U3088 );
nand NAND2_4705 ( P2_U4010 , P2_SUB_1108_U6 , P2_U3030 );
nand NAND2_4706 ( P2_U4011 , P2_IR_REG_10_ , P2_U3978 );
nand NAND2_4707 ( P2_U4012 , U91 , P2_U3088 );
nand NAND2_4708 ( P2_U4013 , P2_SUB_1108_U7 , P2_U3030 );
nand NAND2_4709 ( P2_U4014 , P2_IR_REG_11_ , P2_U3978 );
nand NAND2_4710 ( P2_U4015 , U90 , P2_U3088 );
nand NAND2_4711 ( P2_U4016 , P2_SUB_1108_U8 , P2_U3030 );
nand NAND2_4712 ( P2_U4017 , P2_IR_REG_12_ , P2_U3978 );
nand NAND2_4713 ( P2_U4018 , U89 , P2_U3088 );
nand NAND2_4714 ( P2_U4019 , P2_SUB_1108_U127 , P2_U3030 );
nand NAND2_4715 ( P2_U4020 , P2_IR_REG_13_ , P2_U3978 );
nand NAND2_4716 ( P2_U4021 , U88 , P2_U3088 );
nand NAND2_4717 ( P2_U4022 , P2_SUB_1108_U9 , P2_U3030 );
nand NAND2_4718 ( P2_U4023 , P2_IR_REG_14_ , P2_U3978 );
nand NAND2_4719 ( P2_U4024 , U87 , P2_U3088 );
nand NAND2_4720 ( P2_U4025 , P2_SUB_1108_U10 , P2_U3030 );
nand NAND2_4721 ( P2_U4026 , P2_IR_REG_15_ , P2_U3978 );
nand NAND2_4722 ( P2_U4027 , U86 , P2_U3088 );
nand NAND2_4723 ( P2_U4028 , P2_SUB_1108_U11 , P2_U3030 );
nand NAND2_4724 ( P2_U4029 , P2_IR_REG_16_ , P2_U3978 );
nand NAND2_4725 ( P2_U4030 , U85 , P2_U3088 );
nand NAND2_4726 ( P2_U4031 , P2_SUB_1108_U125 , P2_U3030 );
nand NAND2_4727 ( P2_U4032 , P2_IR_REG_17_ , P2_U3978 );
nand NAND2_4728 ( P2_U4033 , U84 , P2_U3088 );
nand NAND2_4729 ( P2_U4034 , P2_SUB_1108_U12 , P2_U3030 );
nand NAND2_4730 ( P2_U4035 , P2_IR_REG_18_ , P2_U3978 );
nand NAND2_4731 ( P2_U4036 , U83 , P2_U3088 );
nand NAND2_4732 ( P2_U4037 , P2_SUB_1108_U123 , P2_U3030 );
nand NAND2_4733 ( P2_U4038 , P2_IR_REG_19_ , P2_U3978 );
nand NAND2_4734 ( P2_U4039 , U81 , P2_U3088 );
nand NAND2_4735 ( P2_U4040 , P2_SUB_1108_U119 , P2_U3030 );
nand NAND2_4736 ( P2_U4041 , P2_IR_REG_20_ , P2_U3978 );
nand NAND2_4737 ( P2_U4042 , U80 , P2_U3088 );
nand NAND2_4738 ( P2_U4043 , P2_SUB_1108_U116 , P2_U3030 );
nand NAND2_4739 ( P2_U4044 , P2_IR_REG_21_ , P2_U3978 );
nand NAND2_4740 ( P2_U4045 , U79 , P2_U3088 );
nand NAND2_4741 ( P2_U4046 , P2_SUB_1108_U114 , P2_U3030 );
nand NAND2_4742 ( P2_U4047 , P2_IR_REG_22_ , P2_U3978 );
nand NAND2_4743 ( P2_U4048 , U78 , P2_U3088 );
nand NAND2_4744 ( P2_U4049 , P2_SUB_1108_U13 , P2_U3030 );
nand NAND2_4745 ( P2_U4050 , P2_IR_REG_23_ , P2_U3978 );
nand NAND2_4746 ( P2_U4051 , U77 , P2_U3088 );
nand NAND2_4747 ( P2_U4052 , P2_SUB_1108_U14 , P2_U3030 );
nand NAND2_4748 ( P2_U4053 , P2_IR_REG_24_ , P2_U3978 );
nand NAND2_4749 ( P2_U4054 , U76 , P2_U3088 );
nand NAND2_4750 ( P2_U4055 , P2_SUB_1108_U112 , P2_U3030 );
nand NAND2_4751 ( P2_U4056 , P2_IR_REG_25_ , P2_U3978 );
nand NAND2_4752 ( P2_U4057 , U75 , P2_U3088 );
nand NAND2_4753 ( P2_U4058 , P2_SUB_1108_U15 , P2_U3030 );
nand NAND2_4754 ( P2_U4059 , P2_IR_REG_26_ , P2_U3978 );
nand NAND2_4755 ( P2_U4060 , U74 , P2_U3088 );
nand NAND2_4756 ( P2_U4061 , P2_SUB_1108_U110 , P2_U3030 );
nand NAND2_4757 ( P2_U4062 , P2_IR_REG_27_ , P2_U3978 );
nand NAND2_4758 ( P2_U4063 , U73 , P2_U3088 );
nand NAND2_4759 ( P2_U4064 , P2_SUB_1108_U107 , P2_U3030 );
nand NAND2_4760 ( P2_U4065 , P2_IR_REG_28_ , P2_U3978 );
nand NAND2_4761 ( P2_U4066 , U72 , P2_U3088 );
nand NAND2_4762 ( P2_U4067 , P2_SUB_1108_U16 , P2_U3030 );
nand NAND2_4763 ( P2_U4068 , P2_IR_REG_29_ , P2_U3978 );
nand NAND2_4764 ( P2_U4069 , U70 , P2_U3088 );
nand NAND2_4765 ( P2_U4070 , P2_SUB_1108_U104 , P2_U3030 );
nand NAND2_4766 ( P2_U4071 , P2_IR_REG_30_ , P2_U3978 );
nand NAND2_4767 ( P2_U4072 , U69 , P2_U3088 );
nand NAND2_4768 ( P2_U4073 , P2_SUB_1108_U43 , P2_U3030 );
nand NAND2_4769 ( P2_U4074 , P2_IR_REG_31_ , P2_U3978 );
nand NAND2_4770 ( P2_U4075 , P2_U3975 , P2_U5655 );
not NOT1_4771 ( P2_U4076 , P2_U3333 );
nand NAND2_4772 ( P2_U4077 , P2_U3332 , P2_U5646 );
nand NAND2_4773 ( P2_U4078 , P2_U3332 , P2_U5649 );
nand NAND2_4774 ( P2_U4079 , P2_U4076 , P2_D_REG_10_ );
nand NAND2_4775 ( P2_U4080 , P2_U4076 , P2_D_REG_11_ );
nand NAND2_4776 ( P2_U4081 , P2_U4076 , P2_D_REG_12_ );
nand NAND2_4777 ( P2_U4082 , P2_U4076 , P2_D_REG_13_ );
nand NAND2_4778 ( P2_U4083 , P2_U4076 , P2_D_REG_14_ );
nand NAND2_4779 ( P2_U4084 , P2_U4076 , P2_D_REG_15_ );
nand NAND2_4780 ( P2_U4085 , P2_U4076 , P2_D_REG_16_ );
nand NAND2_4781 ( P2_U4086 , P2_U4076 , P2_D_REG_17_ );
nand NAND2_4782 ( P2_U4087 , P2_U4076 , P2_D_REG_18_ );
nand NAND2_4783 ( P2_U4088 , P2_U4076 , P2_D_REG_19_ );
nand NAND2_4784 ( P2_U4089 , P2_U4076 , P2_D_REG_20_ );
nand NAND2_4785 ( P2_U4090 , P2_U4076 , P2_D_REG_21_ );
nand NAND2_4786 ( P2_U4091 , P2_U4076 , P2_D_REG_22_ );
nand NAND2_4787 ( P2_U4092 , P2_U4076 , P2_D_REG_23_ );
nand NAND2_4788 ( P2_U4093 , P2_U4076 , P2_D_REG_24_ );
nand NAND2_4789 ( P2_U4094 , P2_U4076 , P2_D_REG_25_ );
nand NAND2_4790 ( P2_U4095 , P2_U4076 , P2_D_REG_26_ );
nand NAND2_4791 ( P2_U4096 , P2_U4076 , P2_D_REG_27_ );
nand NAND2_4792 ( P2_U4097 , P2_U4076 , P2_D_REG_28_ );
nand NAND2_4793 ( P2_U4098 , P2_U4076 , P2_D_REG_29_ );
nand NAND2_4794 ( P2_U4099 , P2_U4076 , P2_D_REG_2_ );
nand NAND2_4795 ( P2_U4100 , P2_U4076 , P2_D_REG_30_ );
nand NAND2_4796 ( P2_U4101 , P2_U4076 , P2_D_REG_31_ );
nand NAND2_4797 ( P2_U4102 , P2_U4076 , P2_D_REG_3_ );
nand NAND2_4798 ( P2_U4103 , P2_U4076 , P2_D_REG_4_ );
nand NAND2_4799 ( P2_U4104 , P2_U4076 , P2_D_REG_5_ );
nand NAND2_4800 ( P2_U4105 , P2_U4076 , P2_D_REG_6_ );
nand NAND2_4801 ( P2_U4106 , P2_U4076 , P2_D_REG_7_ );
nand NAND2_4802 ( P2_U4107 , P2_U4076 , P2_D_REG_8_ );
nand NAND2_4803 ( P2_U4108 , P2_U4076 , P2_D_REG_9_ );
nand NAND2_4804 ( P2_U4109 , P2_U5674 , P2_U5671 );
nand NAND3_4805 ( P2_U4110 , P2_U5693 , P2_U5692 , P2_U3340 );
nand NAND2_4806 ( P2_U4111 , P2_U3020 , P2_REG2_REG_1_ );
nand NAND2_4807 ( P2_U4112 , P2_U3021 , P2_REG1_REG_1_ );
nand NAND2_4808 ( P2_U4113 , P2_U3022 , P2_REG0_REG_1_ );
nand NAND2_4809 ( P2_U4114 , P2_REG3_REG_1_ , P2_U3019 );
not NOT1_4810 ( P2_U4115 , P2_U3080 );
nand NAND2_4811 ( P2_U4116 , P2_U3390 , P2_U3934 );
nand NAND2_4812 ( P2_U4117 , P2_U3931 , P2_R1146_U20 );
nand NAND2_4813 ( P2_U4118 , P2_U3930 , P2_R1113_U20 );
nand NAND2_4814 ( P2_U4119 , P2_U3926 , P2_R1131_U95 );
nand NAND2_4815 ( P2_U4120 , P2_U3941 , P2_R1179_U20 );
nand NAND2_4816 ( P2_U4121 , P2_U3943 , P2_R1203_U20 );
nand NAND2_4817 ( P2_U4122 , P2_U3014 , P2_R1164_U95 );
nand NAND2_4818 ( P2_U4123 , P2_U3922 , P2_R1233_U95 );
not NOT1_4819 ( P2_U4124 , P2_U3348 );
nand NAND2_4820 ( P2_U4125 , P2_U3427 , P2_U3027 );
nand NAND2_4821 ( P2_U4126 , P2_U3026 , P2_U3080 );
nand NAND2_4822 ( P2_U4127 , P2_R1215_U96 , P2_U3025 );
nand NAND2_4823 ( P2_U4128 , P2_U3427 , P2_U4116 );
nand NAND4_4824 ( P2_U4129 , P2_U4128 , P2_U4126 , P2_U3565 , P2_U4124 );
nand NAND2_4825 ( P2_U4130 , P2_REG2_REG_2_ , P2_U3020 );
nand NAND2_4826 ( P2_U4131 , P2_REG1_REG_2_ , P2_U3021 );
nand NAND2_4827 ( P2_U4132 , P2_REG0_REG_2_ , P2_U3022 );
nand NAND2_4828 ( P2_U4133 , P2_REG3_REG_2_ , P2_U3019 );
not NOT1_4829 ( P2_U4134 , P2_U3070 );
nand NAND2_4830 ( P2_U4135 , P2_REG2_REG_0_ , P2_U3020 );
nand NAND2_4831 ( P2_U4136 , P2_REG1_REG_0_ , P2_U3021 );
nand NAND2_4832 ( P2_U4137 , P2_REG0_REG_0_ , P2_U3022 );
nand NAND2_4833 ( P2_U4138 , P2_REG3_REG_0_ , P2_U3019 );
not NOT1_4834 ( P2_U4139 , P2_U3079 );
nand NAND2_4835 ( P2_U4140 , P2_U3035 , P2_U3079 );
nand NAND2_4836 ( P2_U4141 , P2_R1146_U97 , P2_U3931 );
nand NAND2_4837 ( P2_U4142 , P2_R1113_U97 , P2_U3930 );
nand NAND2_4838 ( P2_U4143 , P2_R1131_U94 , P2_U3926 );
nand NAND2_4839 ( P2_U4144 , P2_R1179_U97 , P2_U3941 );
nand NAND2_4840 ( P2_U4145 , P2_R1203_U97 , P2_U3943 );
nand NAND2_4841 ( P2_U4146 , P2_R1164_U94 , P2_U3014 );
nand NAND2_4842 ( P2_U4147 , P2_R1233_U94 , P2_U3922 );
not NOT1_4843 ( P2_U4148 , P2_U3349 );
nand NAND2_4844 ( P2_U4149 , P2_R1275_U55 , P2_U3027 );
nand NAND2_4845 ( P2_U4150 , P2_U3026 , P2_U3070 );
nand NAND2_4846 ( P2_U4151 , P2_R1215_U95 , P2_U3025 );
nand NAND2_4847 ( P2_U4152 , P2_U3432 , P2_U4116 );
nand NAND2_4848 ( P2_U4153 , P2_U3581 , P2_U4148 );
nand NAND2_4849 ( P2_U4154 , P2_REG2_REG_3_ , P2_U3020 );
nand NAND2_4850 ( P2_U4155 , P2_REG1_REG_3_ , P2_U3021 );
nand NAND2_4851 ( P2_U4156 , P2_REG0_REG_3_ , P2_U3022 );
nand NAND2_4852 ( P2_U4157 , P2_ADD_1119_U4 , P2_U3019 );
not NOT1_4853 ( P2_U4158 , P2_U3066 );
nand NAND2_4854 ( P2_U4159 , P2_U3035 , P2_U3080 );
nand NAND2_4855 ( P2_U4160 , P2_R1146_U107 , P2_U3931 );
nand NAND2_4856 ( P2_U4161 , P2_R1113_U107 , P2_U3930 );
nand NAND2_4857 ( P2_U4162 , P2_R1131_U16 , P2_U3926 );
nand NAND2_4858 ( P2_U4163 , P2_R1179_U107 , P2_U3941 );
nand NAND2_4859 ( P2_U4164 , P2_R1203_U107 , P2_U3943 );
nand NAND2_4860 ( P2_U4165 , P2_R1164_U16 , P2_U3014 );
nand NAND2_4861 ( P2_U4166 , P2_R1233_U16 , P2_U3922 );
not NOT1_4862 ( P2_U4167 , P2_U3350 );
nand NAND2_4863 ( P2_U4168 , P2_R1275_U18 , P2_U3027 );
nand NAND2_4864 ( P2_U4169 , P2_U3026 , P2_U3066 );
nand NAND2_4865 ( P2_U4170 , P2_R1215_U17 , P2_U3025 );
nand NAND2_4866 ( P2_U4171 , P2_U3435 , P2_U4116 );
nand NAND2_4867 ( P2_U4172 , P2_U3585 , P2_U4167 );
nand NAND2_4868 ( P2_U4173 , P2_REG2_REG_4_ , P2_U3020 );
nand NAND2_4869 ( P2_U4174 , P2_REG1_REG_4_ , P2_U3021 );
nand NAND2_4870 ( P2_U4175 , P2_REG0_REG_4_ , P2_U3022 );
nand NAND2_4871 ( P2_U4176 , P2_ADD_1119_U55 , P2_U3019 );
not NOT1_4872 ( P2_U4177 , P2_U3062 );
nand NAND2_4873 ( P2_U4178 , P2_U3035 , P2_U3070 );
nand NAND2_4874 ( P2_U4179 , P2_R1146_U17 , P2_U3931 );
nand NAND2_4875 ( P2_U4180 , P2_R1113_U17 , P2_U3930 );
nand NAND2_4876 ( P2_U4181 , P2_R1131_U100 , P2_U3926 );
nand NAND2_4877 ( P2_U4182 , P2_R1179_U17 , P2_U3941 );
nand NAND2_4878 ( P2_U4183 , P2_R1203_U17 , P2_U3943 );
nand NAND2_4879 ( P2_U4184 , P2_R1164_U100 , P2_U3014 );
nand NAND2_4880 ( P2_U4185 , P2_R1233_U100 , P2_U3922 );
not NOT1_4881 ( P2_U4186 , P2_U3351 );
nand NAND2_4882 ( P2_U4187 , P2_R1275_U20 , P2_U3027 );
nand NAND2_4883 ( P2_U4188 , P2_U3026 , P2_U3062 );
nand NAND2_4884 ( P2_U4189 , P2_R1215_U101 , P2_U3025 );
nand NAND2_4885 ( P2_U4190 , P2_U3438 , P2_U4116 );
nand NAND2_4886 ( P2_U4191 , P2_U3589 , P2_U4186 );
nand NAND2_4887 ( P2_U4192 , P2_REG2_REG_5_ , P2_U3020 );
nand NAND2_4888 ( P2_U4193 , P2_REG1_REG_5_ , P2_U3021 );
nand NAND2_4889 ( P2_U4194 , P2_REG0_REG_5_ , P2_U3022 );
nand NAND2_4890 ( P2_U4195 , P2_ADD_1119_U54 , P2_U3019 );
not NOT1_4891 ( P2_U4196 , P2_U3069 );
nand NAND2_4892 ( P2_U4197 , P2_U3035 , P2_U3066 );
nand NAND2_4893 ( P2_U4198 , P2_R1146_U106 , P2_U3931 );
nand NAND2_4894 ( P2_U4199 , P2_R1113_U106 , P2_U3930 );
nand NAND2_4895 ( P2_U4200 , P2_R1131_U99 , P2_U3926 );
nand NAND2_4896 ( P2_U4201 , P2_R1179_U106 , P2_U3941 );
nand NAND2_4897 ( P2_U4202 , P2_R1203_U106 , P2_U3943 );
nand NAND2_4898 ( P2_U4203 , P2_R1164_U99 , P2_U3014 );
nand NAND2_4899 ( P2_U4204 , P2_R1233_U99 , P2_U3922 );
not NOT1_4900 ( P2_U4205 , P2_U3352 );
nand NAND2_4901 ( P2_U4206 , P2_R1275_U21 , P2_U3027 );
nand NAND2_4902 ( P2_U4207 , P2_U3026 , P2_U3069 );
nand NAND2_4903 ( P2_U4208 , P2_R1215_U100 , P2_U3025 );
nand NAND2_4904 ( P2_U4209 , P2_U3441 , P2_U4116 );
nand NAND2_4905 ( P2_U4210 , P2_U3593 , P2_U4205 );
nand NAND2_4906 ( P2_U4211 , P2_REG2_REG_6_ , P2_U3020 );
nand NAND2_4907 ( P2_U4212 , P2_REG1_REG_6_ , P2_U3021 );
nand NAND2_4908 ( P2_U4213 , P2_REG0_REG_6_ , P2_U3022 );
nand NAND2_4909 ( P2_U4214 , P2_ADD_1119_U53 , P2_U3019 );
not NOT1_4910 ( P2_U4215 , P2_U3073 );
nand NAND2_4911 ( P2_U4216 , P2_U3035 , P2_U3062 );
nand NAND2_4912 ( P2_U4217 , P2_R1146_U105 , P2_U3931 );
nand NAND2_4913 ( P2_U4218 , P2_R1113_U105 , P2_U3930 );
nand NAND2_4914 ( P2_U4219 , P2_R1131_U17 , P2_U3926 );
nand NAND2_4915 ( P2_U4220 , P2_R1179_U105 , P2_U3941 );
nand NAND2_4916 ( P2_U4221 , P2_R1203_U105 , P2_U3943 );
nand NAND2_4917 ( P2_U4222 , P2_R1164_U17 , P2_U3014 );
nand NAND2_4918 ( P2_U4223 , P2_R1233_U17 , P2_U3922 );
not NOT1_4919 ( P2_U4224 , P2_U3353 );
nand NAND2_4920 ( P2_U4225 , P2_R1275_U65 , P2_U3027 );
nand NAND2_4921 ( P2_U4226 , P2_U3026 , P2_U3073 );
nand NAND2_4922 ( P2_U4227 , P2_R1215_U18 , P2_U3025 );
nand NAND2_4923 ( P2_U4228 , P2_U3444 , P2_U4116 );
nand NAND2_4924 ( P2_U4229 , P2_U3597 , P2_U4224 );
nand NAND2_4925 ( P2_U4230 , P2_REG2_REG_7_ , P2_U3020 );
nand NAND2_4926 ( P2_U4231 , P2_REG1_REG_7_ , P2_U3021 );
nand NAND2_4927 ( P2_U4232 , P2_REG0_REG_7_ , P2_U3022 );
nand NAND2_4928 ( P2_U4233 , P2_ADD_1119_U52 , P2_U3019 );
not NOT1_4929 ( P2_U4234 , P2_U3072 );
nand NAND2_4930 ( P2_U4235 , P2_U3035 , P2_U3069 );
nand NAND2_4931 ( P2_U4236 , P2_R1146_U18 , P2_U3931 );
nand NAND2_4932 ( P2_U4237 , P2_R1113_U18 , P2_U3930 );
nand NAND2_4933 ( P2_U4238 , P2_R1131_U98 , P2_U3926 );
nand NAND2_4934 ( P2_U4239 , P2_R1179_U18 , P2_U3941 );
nand NAND2_4935 ( P2_U4240 , P2_R1203_U18 , P2_U3943 );
nand NAND2_4936 ( P2_U4241 , P2_R1164_U98 , P2_U3014 );
nand NAND2_4937 ( P2_U4242 , P2_R1233_U98 , P2_U3922 );
not NOT1_4938 ( P2_U4243 , P2_U3354 );
nand NAND2_4939 ( P2_U4244 , P2_R1275_U22 , P2_U3027 );
nand NAND2_4940 ( P2_U4245 , P2_U3026 , P2_U3072 );
nand NAND2_4941 ( P2_U4246 , P2_R1215_U99 , P2_U3025 );
nand NAND2_4942 ( P2_U4247 , P2_U3447 , P2_U4116 );
nand NAND2_4943 ( P2_U4248 , P2_U3601 , P2_U4243 );
nand NAND2_4944 ( P2_U4249 , P2_REG2_REG_8_ , P2_U3020 );
nand NAND2_4945 ( P2_U4250 , P2_REG1_REG_8_ , P2_U3021 );
nand NAND2_4946 ( P2_U4251 , P2_REG0_REG_8_ , P2_U3022 );
nand NAND2_4947 ( P2_U4252 , P2_ADD_1119_U51 , P2_U3019 );
not NOT1_4948 ( P2_U4253 , P2_U3086 );
nand NAND2_4949 ( P2_U4254 , P2_U3035 , P2_U3073 );
nand NAND2_4950 ( P2_U4255 , P2_R1146_U104 , P2_U3931 );
nand NAND2_4951 ( P2_U4256 , P2_R1113_U104 , P2_U3930 );
nand NAND2_4952 ( P2_U4257 , P2_R1131_U18 , P2_U3926 );
nand NAND2_4953 ( P2_U4258 , P2_R1179_U104 , P2_U3941 );
nand NAND2_4954 ( P2_U4259 , P2_R1203_U104 , P2_U3943 );
nand NAND2_4955 ( P2_U4260 , P2_R1164_U18 , P2_U3014 );
nand NAND2_4956 ( P2_U4261 , P2_R1233_U18 , P2_U3922 );
not NOT1_4957 ( P2_U4262 , P2_U3355 );
nand NAND2_4958 ( P2_U4263 , P2_R1275_U23 , P2_U3027 );
nand NAND2_4959 ( P2_U4264 , P2_U3026 , P2_U3086 );
nand NAND2_4960 ( P2_U4265 , P2_R1215_U19 , P2_U3025 );
nand NAND2_4961 ( P2_U4266 , P2_U3450 , P2_U4116 );
nand NAND2_4962 ( P2_U4267 , P2_U3605 , P2_U4262 );
nand NAND2_4963 ( P2_U4268 , P2_REG2_REG_9_ , P2_U3020 );
nand NAND2_4964 ( P2_U4269 , P2_REG1_REG_9_ , P2_U3021 );
nand NAND2_4965 ( P2_U4270 , P2_REG0_REG_9_ , P2_U3022 );
nand NAND2_4966 ( P2_U4271 , P2_ADD_1119_U50 , P2_U3019 );
not NOT1_4967 ( P2_U4272 , P2_U3085 );
nand NAND2_4968 ( P2_U4273 , P2_U3035 , P2_U3072 );
nand NAND2_4969 ( P2_U4274 , P2_R1146_U19 , P2_U3931 );
nand NAND2_4970 ( P2_U4275 , P2_R1113_U19 , P2_U3930 );
nand NAND2_4971 ( P2_U4276 , P2_R1131_U97 , P2_U3926 );
nand NAND2_4972 ( P2_U4277 , P2_R1179_U19 , P2_U3941 );
nand NAND2_4973 ( P2_U4278 , P2_R1203_U19 , P2_U3943 );
nand NAND2_4974 ( P2_U4279 , P2_R1164_U97 , P2_U3014 );
nand NAND2_4975 ( P2_U4280 , P2_R1233_U97 , P2_U3922 );
not NOT1_4976 ( P2_U4281 , P2_U3356 );
nand NAND2_4977 ( P2_U4282 , P2_R1275_U24 , P2_U3027 );
nand NAND2_4978 ( P2_U4283 , P2_U3026 , P2_U3085 );
nand NAND2_4979 ( P2_U4284 , P2_R1215_U98 , P2_U3025 );
nand NAND2_4980 ( P2_U4285 , P2_U3453 , P2_U4116 );
nand NAND2_4981 ( P2_U4286 , P2_U3609 , P2_U4281 );
nand NAND2_4982 ( P2_U4287 , P2_REG2_REG_10_ , P2_U3020 );
nand NAND2_4983 ( P2_U4288 , P2_REG1_REG_10_ , P2_U3021 );
nand NAND2_4984 ( P2_U4289 , P2_REG0_REG_10_ , P2_U3022 );
nand NAND2_4985 ( P2_U4290 , P2_ADD_1119_U74 , P2_U3019 );
not NOT1_4986 ( P2_U4291 , P2_U3064 );
nand NAND2_4987 ( P2_U4292 , P2_U3035 , P2_U3086 );
nand NAND2_4988 ( P2_U4293 , P2_R1146_U103 , P2_U3931 );
nand NAND2_4989 ( P2_U4294 , P2_R1113_U103 , P2_U3930 );
nand NAND2_4990 ( P2_U4295 , P2_R1131_U96 , P2_U3926 );
nand NAND2_4991 ( P2_U4296 , P2_R1179_U103 , P2_U3941 );
nand NAND2_4992 ( P2_U4297 , P2_R1203_U103 , P2_U3943 );
nand NAND2_4993 ( P2_U4298 , P2_R1164_U96 , P2_U3014 );
nand NAND2_4994 ( P2_U4299 , P2_R1233_U96 , P2_U3922 );
not NOT1_4995 ( P2_U4300 , P2_U3357 );
nand NAND2_4996 ( P2_U4301 , P2_R1275_U63 , P2_U3027 );
nand NAND2_4997 ( P2_U4302 , P2_U3026 , P2_U3064 );
nand NAND2_4998 ( P2_U4303 , P2_R1215_U97 , P2_U3025 );
nand NAND2_4999 ( P2_U4304 , P2_U3456 , P2_U4116 );
nand NAND2_5000 ( P2_U4305 , P2_U3613 , P2_U4300 );
nand NAND2_5001 ( P2_U4306 , P2_REG2_REG_11_ , P2_U3020 );
nand NAND2_5002 ( P2_U4307 , P2_REG1_REG_11_ , P2_U3021 );
nand NAND2_5003 ( P2_U4308 , P2_REG0_REG_11_ , P2_U3022 );
nand NAND2_5004 ( P2_U4309 , P2_ADD_1119_U73 , P2_U3019 );
not NOT1_5005 ( P2_U4310 , P2_U3065 );
nand NAND2_5006 ( P2_U4311 , P2_U3035 , P2_U3085 );
nand NAND2_5007 ( P2_U4312 , P2_R1146_U113 , P2_U3931 );
nand NAND2_5008 ( P2_U4313 , P2_R1113_U113 , P2_U3930 );
nand NAND2_5009 ( P2_U4314 , P2_R1131_U10 , P2_U3926 );
nand NAND2_5010 ( P2_U4315 , P2_R1179_U113 , P2_U3941 );
nand NAND2_5011 ( P2_U4316 , P2_R1203_U113 , P2_U3943 );
nand NAND2_5012 ( P2_U4317 , P2_R1164_U10 , P2_U3014 );
nand NAND2_5013 ( P2_U4318 , P2_R1233_U10 , P2_U3922 );
not NOT1_5014 ( P2_U4319 , P2_U3358 );
nand NAND2_5015 ( P2_U4320 , P2_R1275_U6 , P2_U3027 );
nand NAND2_5016 ( P2_U4321 , P2_U3026 , P2_U3065 );
nand NAND2_5017 ( P2_U4322 , P2_R1215_U11 , P2_U3025 );
nand NAND2_5018 ( P2_U4323 , P2_U3459 , P2_U4116 );
nand NAND2_5019 ( P2_U4324 , P2_U3617 , P2_U4319 );
nand NAND2_5020 ( P2_U4325 , P2_REG2_REG_12_ , P2_U3020 );
nand NAND2_5021 ( P2_U4326 , P2_REG1_REG_12_ , P2_U3021 );
nand NAND2_5022 ( P2_U4327 , P2_REG0_REG_12_ , P2_U3022 );
nand NAND2_5023 ( P2_U4328 , P2_ADD_1119_U72 , P2_U3019 );
not NOT1_5024 ( P2_U4329 , P2_U3074 );
nand NAND2_5025 ( P2_U4330 , P2_U3035 , P2_U3064 );
nand NAND2_5026 ( P2_U4331 , P2_R1146_U12 , P2_U3931 );
nand NAND2_5027 ( P2_U4332 , P2_R1113_U12 , P2_U3930 );
nand NAND2_5028 ( P2_U4333 , P2_R1131_U114 , P2_U3926 );
nand NAND2_5029 ( P2_U4334 , P2_R1179_U12 , P2_U3941 );
nand NAND2_5030 ( P2_U4335 , P2_R1203_U12 , P2_U3943 );
nand NAND2_5031 ( P2_U4336 , P2_R1164_U114 , P2_U3014 );
nand NAND2_5032 ( P2_U4337 , P2_R1233_U114 , P2_U3922 );
not NOT1_5033 ( P2_U4338 , P2_U3359 );
nand NAND2_5034 ( P2_U4339 , P2_R1275_U7 , P2_U3027 );
nand NAND2_5035 ( P2_U4340 , P2_U3026 , P2_U3074 );
nand NAND2_5036 ( P2_U4341 , P2_R1215_U115 , P2_U3025 );
nand NAND2_5037 ( P2_U4342 , P2_U3462 , P2_U4116 );
nand NAND2_5038 ( P2_U4343 , P2_U3621 , P2_U4338 );
nand NAND2_5039 ( P2_U4344 , P2_REG2_REG_13_ , P2_U3020 );
nand NAND2_5040 ( P2_U4345 , P2_REG1_REG_13_ , P2_U3021 );
nand NAND2_5041 ( P2_U4346 , P2_REG0_REG_13_ , P2_U3022 );
nand NAND2_5042 ( P2_U4347 , P2_ADD_1119_U71 , P2_U3019 );
not NOT1_5043 ( P2_U4348 , P2_U3082 );
nand NAND2_5044 ( P2_U4349 , P2_U3035 , P2_U3065 );
nand NAND2_5045 ( P2_U4350 , P2_R1146_U102 , P2_U3931 );
nand NAND2_5046 ( P2_U4351 , P2_R1113_U102 , P2_U3930 );
nand NAND2_5047 ( P2_U4352 , P2_R1131_U113 , P2_U3926 );
nand NAND2_5048 ( P2_U4353 , P2_R1179_U102 , P2_U3941 );
nand NAND2_5049 ( P2_U4354 , P2_R1203_U102 , P2_U3943 );
nand NAND2_5050 ( P2_U4355 , P2_R1164_U113 , P2_U3014 );
nand NAND2_5051 ( P2_U4356 , P2_R1233_U113 , P2_U3922 );
not NOT1_5052 ( P2_U4357 , P2_U3360 );
nand NAND2_5053 ( P2_U4358 , P2_R1275_U8 , P2_U3027 );
nand NAND2_5054 ( P2_U4359 , P2_U3026 , P2_U3082 );
nand NAND2_5055 ( P2_U4360 , P2_R1215_U114 , P2_U3025 );
nand NAND2_5056 ( P2_U4361 , P2_U3465 , P2_U4116 );
nand NAND2_5057 ( P2_U4362 , P2_U3625 , P2_U4357 );
nand NAND2_5058 ( P2_U4363 , P2_REG2_REG_14_ , P2_U3020 );
nand NAND2_5059 ( P2_U4364 , P2_REG1_REG_14_ , P2_U3021 );
nand NAND2_5060 ( P2_U4365 , P2_REG0_REG_14_ , P2_U3022 );
nand NAND2_5061 ( P2_U4366 , P2_ADD_1119_U70 , P2_U3019 );
not NOT1_5062 ( P2_U4367 , P2_U3081 );
nand NAND2_5063 ( P2_U4368 , P2_U3035 , P2_U3074 );
nand NAND2_5064 ( P2_U4369 , P2_R1146_U101 , P2_U3931 );
nand NAND2_5065 ( P2_U4370 , P2_R1113_U101 , P2_U3930 );
nand NAND2_5066 ( P2_U4371 , P2_R1131_U11 , P2_U3926 );
nand NAND2_5067 ( P2_U4372 , P2_R1179_U101 , P2_U3941 );
nand NAND2_5068 ( P2_U4373 , P2_R1203_U101 , P2_U3943 );
nand NAND2_5069 ( P2_U4374 , P2_R1164_U11 , P2_U3014 );
nand NAND2_5070 ( P2_U4375 , P2_R1233_U11 , P2_U3922 );
not NOT1_5071 ( P2_U4376 , P2_U3361 );
nand NAND2_5072 ( P2_U4377 , P2_R1275_U86 , P2_U3027 );
nand NAND2_5073 ( P2_U4378 , P2_U3026 , P2_U3081 );
nand NAND2_5074 ( P2_U4379 , P2_R1215_U12 , P2_U3025 );
nand NAND2_5075 ( P2_U4380 , P2_U3468 , P2_U4116 );
nand NAND2_5076 ( P2_U4381 , P2_U3629 , P2_U4376 );
nand NAND2_5077 ( P2_U4382 , P2_REG2_REG_15_ , P2_U3020 );
nand NAND2_5078 ( P2_U4383 , P2_REG1_REG_15_ , P2_U3021 );
nand NAND2_5079 ( P2_U4384 , P2_REG0_REG_15_ , P2_U3022 );
nand NAND2_5080 ( P2_U4385 , P2_ADD_1119_U69 , P2_U3019 );
not NOT1_5081 ( P2_U4386 , P2_U3076 );
nand NAND2_5082 ( P2_U4387 , P2_U3035 , P2_U3082 );
nand NAND2_5083 ( P2_U4388 , P2_R1146_U112 , P2_U3931 );
nand NAND2_5084 ( P2_U4389 , P2_R1113_U112 , P2_U3930 );
nand NAND2_5085 ( P2_U4390 , P2_R1131_U112 , P2_U3926 );
nand NAND2_5086 ( P2_U4391 , P2_R1179_U112 , P2_U3941 );
nand NAND2_5087 ( P2_U4392 , P2_R1203_U112 , P2_U3943 );
nand NAND2_5088 ( P2_U4393 , P2_R1164_U112 , P2_U3014 );
nand NAND2_5089 ( P2_U4394 , P2_R1233_U112 , P2_U3922 );
not NOT1_5090 ( P2_U4395 , P2_U3362 );
nand NAND2_5091 ( P2_U4396 , P2_R1275_U9 , P2_U3027 );
nand NAND2_5092 ( P2_U4397 , P2_U3026 , P2_U3076 );
nand NAND2_5093 ( P2_U4398 , P2_R1215_U113 , P2_U3025 );
nand NAND2_5094 ( P2_U4399 , P2_U3471 , P2_U4116 );
nand NAND2_5095 ( P2_U4400 , P2_U3633 , P2_U4395 );
nand NAND2_5096 ( P2_U4401 , P2_REG2_REG_16_ , P2_U3020 );
nand NAND2_5097 ( P2_U4402 , P2_REG1_REG_16_ , P2_U3021 );
nand NAND2_5098 ( P2_U4403 , P2_REG0_REG_16_ , P2_U3022 );
nand NAND2_5099 ( P2_U4404 , P2_ADD_1119_U68 , P2_U3019 );
not NOT1_5100 ( P2_U4405 , P2_U3075 );
nand NAND2_5101 ( P2_U4406 , P2_U3035 , P2_U3081 );
nand NAND2_5102 ( P2_U4407 , P2_R1146_U111 , P2_U3931 );
nand NAND2_5103 ( P2_U4408 , P2_R1113_U111 , P2_U3930 );
nand NAND2_5104 ( P2_U4409 , P2_R1131_U111 , P2_U3926 );
nand NAND2_5105 ( P2_U4410 , P2_R1179_U111 , P2_U3941 );
nand NAND2_5106 ( P2_U4411 , P2_R1203_U111 , P2_U3943 );
nand NAND2_5107 ( P2_U4412 , P2_R1164_U111 , P2_U3014 );
nand NAND2_5108 ( P2_U4413 , P2_R1233_U111 , P2_U3922 );
not NOT1_5109 ( P2_U4414 , P2_U3363 );
nand NAND2_5110 ( P2_U4415 , P2_R1275_U10 , P2_U3027 );
nand NAND2_5111 ( P2_U4416 , P2_U3026 , P2_U3075 );
nand NAND2_5112 ( P2_U4417 , P2_R1215_U112 , P2_U3025 );
nand NAND2_5113 ( P2_U4418 , P2_U3474 , P2_U4116 );
nand NAND2_5114 ( P2_U4419 , P2_U3637 , P2_U4414 );
nand NAND2_5115 ( P2_U4420 , P2_REG2_REG_17_ , P2_U3020 );
nand NAND2_5116 ( P2_U4421 , P2_REG1_REG_17_ , P2_U3021 );
nand NAND2_5117 ( P2_U4422 , P2_REG0_REG_17_ , P2_U3022 );
nand NAND2_5118 ( P2_U4423 , P2_ADD_1119_U67 , P2_U3019 );
not NOT1_5119 ( P2_U4424 , P2_U3071 );
nand NAND2_5120 ( P2_U4425 , P2_U3035 , P2_U3076 );
nand NAND2_5121 ( P2_U4426 , P2_R1146_U13 , P2_U3931 );
nand NAND2_5122 ( P2_U4427 , P2_R1113_U13 , P2_U3930 );
nand NAND2_5123 ( P2_U4428 , P2_R1131_U110 , P2_U3926 );
nand NAND2_5124 ( P2_U4429 , P2_R1179_U13 , P2_U3941 );
nand NAND2_5125 ( P2_U4430 , P2_R1203_U13 , P2_U3943 );
nand NAND2_5126 ( P2_U4431 , P2_R1164_U110 , P2_U3014 );
nand NAND2_5127 ( P2_U4432 , P2_R1233_U110 , P2_U3922 );
not NOT1_5128 ( P2_U4433 , P2_U3364 );
nand NAND2_5129 ( P2_U4434 , P2_R1275_U11 , P2_U3027 );
nand NAND2_5130 ( P2_U4435 , P2_U3026 , P2_U3071 );
nand NAND2_5131 ( P2_U4436 , P2_R1215_U111 , P2_U3025 );
nand NAND2_5132 ( P2_U4437 , P2_U3477 , P2_U4116 );
nand NAND2_5133 ( P2_U4438 , P2_U3641 , P2_U4433 );
nand NAND2_5134 ( P2_U4439 , P2_REG2_REG_18_ , P2_U3020 );
nand NAND2_5135 ( P2_U4440 , P2_REG1_REG_18_ , P2_U3021 );
nand NAND2_5136 ( P2_U4441 , P2_REG0_REG_18_ , P2_U3022 );
nand NAND2_5137 ( P2_U4442 , P2_ADD_1119_U66 , P2_U3019 );
not NOT1_5138 ( P2_U4443 , P2_U3084 );
nand NAND2_5139 ( P2_U4444 , P2_U3035 , P2_U3075 );
nand NAND2_5140 ( P2_U4445 , P2_R1146_U100 , P2_U3931 );
nand NAND2_5141 ( P2_U4446 , P2_R1113_U100 , P2_U3930 );
nand NAND2_5142 ( P2_U4447 , P2_R1131_U12 , P2_U3926 );
nand NAND2_5143 ( P2_U4448 , P2_R1179_U100 , P2_U3941 );
nand NAND2_5144 ( P2_U4449 , P2_R1203_U100 , P2_U3943 );
nand NAND2_5145 ( P2_U4450 , P2_R1164_U12 , P2_U3014 );
nand NAND2_5146 ( P2_U4451 , P2_R1233_U12 , P2_U3922 );
not NOT1_5147 ( P2_U4452 , P2_U3365 );
nand NAND2_5148 ( P2_U4453 , P2_R1275_U84 , P2_U3027 );
nand NAND2_5149 ( P2_U4454 , P2_U3026 , P2_U3084 );
nand NAND2_5150 ( P2_U4455 , P2_R1215_U13 , P2_U3025 );
nand NAND2_5151 ( P2_U4456 , P2_U3480 , P2_U4116 );
nand NAND2_5152 ( P2_U4457 , P2_U3645 , P2_U4452 );
nand NAND2_5153 ( P2_U4458 , P2_REG2_REG_19_ , P2_U3020 );
nand NAND2_5154 ( P2_U4459 , P2_REG1_REG_19_ , P2_U3021 );
nand NAND2_5155 ( P2_U4460 , P2_REG0_REG_19_ , P2_U3022 );
nand NAND2_5156 ( P2_U4461 , P2_ADD_1119_U65 , P2_U3019 );
not NOT1_5157 ( P2_U4462 , P2_U3083 );
nand NAND2_5158 ( P2_U4463 , P2_U3035 , P2_U3071 );
nand NAND2_5159 ( P2_U4464 , P2_R1146_U99 , P2_U3931 );
nand NAND2_5160 ( P2_U4465 , P2_R1113_U99 , P2_U3930 );
nand NAND2_5161 ( P2_U4466 , P2_R1131_U109 , P2_U3926 );
nand NAND2_5162 ( P2_U4467 , P2_R1179_U99 , P2_U3941 );
nand NAND2_5163 ( P2_U4468 , P2_R1203_U99 , P2_U3943 );
nand NAND2_5164 ( P2_U4469 , P2_R1164_U109 , P2_U3014 );
nand NAND2_5165 ( P2_U4470 , P2_R1233_U109 , P2_U3922 );
not NOT1_5166 ( P2_U4471 , P2_U3366 );
nand NAND2_5167 ( P2_U4472 , P2_R1275_U12 , P2_U3027 );
nand NAND2_5168 ( P2_U4473 , P2_U3026 , P2_U3083 );
nand NAND2_5169 ( P2_U4474 , P2_R1215_U110 , P2_U3025 );
nand NAND2_5170 ( P2_U4475 , P2_U3483 , P2_U4116 );
nand NAND2_5171 ( P2_U4476 , P2_U3649 , P2_U4471 );
nand NAND2_5172 ( P2_U4477 , P2_REG2_REG_20_ , P2_U3020 );
nand NAND2_5173 ( P2_U4478 , P2_REG1_REG_20_ , P2_U3021 );
nand NAND2_5174 ( P2_U4479 , P2_REG0_REG_20_ , P2_U3022 );
nand NAND2_5175 ( P2_U4480 , P2_ADD_1119_U64 , P2_U3019 );
not NOT1_5176 ( P2_U4481 , P2_U3078 );
nand NAND2_5177 ( P2_U4482 , P2_U3035 , P2_U3084 );
nand NAND2_5178 ( P2_U4483 , P2_R1146_U98 , P2_U3931 );
nand NAND2_5179 ( P2_U4484 , P2_R1113_U98 , P2_U3930 );
nand NAND2_5180 ( P2_U4485 , P2_R1131_U108 , P2_U3926 );
nand NAND2_5181 ( P2_U4486 , P2_R1179_U98 , P2_U3941 );
nand NAND2_5182 ( P2_U4487 , P2_R1203_U98 , P2_U3943 );
nand NAND2_5183 ( P2_U4488 , P2_R1164_U108 , P2_U3014 );
nand NAND2_5184 ( P2_U4489 , P2_R1233_U108 , P2_U3922 );
not NOT1_5185 ( P2_U4490 , P2_U3367 );
nand NAND2_5186 ( P2_U4491 , P2_R1275_U82 , P2_U3027 );
nand NAND2_5187 ( P2_U4492 , P2_U3026 , P2_U3078 );
nand NAND2_5188 ( P2_U4493 , P2_R1215_U109 , P2_U3025 );
nand NAND2_5189 ( P2_U4494 , P2_U3485 , P2_U4116 );
nand NAND2_5190 ( P2_U4495 , P2_U3653 , P2_U4490 );
nand NAND2_5191 ( P2_U4496 , P2_REG2_REG_21_ , P2_U3020 );
nand NAND2_5192 ( P2_U4497 , P2_REG1_REG_21_ , P2_U3021 );
nand NAND2_5193 ( P2_U4498 , P2_REG0_REG_21_ , P2_U3022 );
nand NAND2_5194 ( P2_U4499 , P2_ADD_1119_U63 , P2_U3019 );
not NOT1_5195 ( P2_U4500 , P2_U3077 );
nand NAND2_5196 ( P2_U4501 , P2_U3035 , P2_U3083 );
nand NAND2_5197 ( P2_U4502 , P2_R1146_U96 , P2_U3931 );
nand NAND2_5198 ( P2_U4503 , P2_R1113_U96 , P2_U3930 );
nand NAND2_5199 ( P2_U4504 , P2_R1131_U13 , P2_U3926 );
nand NAND2_5200 ( P2_U4505 , P2_R1179_U96 , P2_U3941 );
nand NAND2_5201 ( P2_U4506 , P2_R1203_U96 , P2_U3943 );
nand NAND2_5202 ( P2_U4507 , P2_R1164_U13 , P2_U3014 );
nand NAND2_5203 ( P2_U4508 , P2_R1233_U13 , P2_U3922 );
not NOT1_5204 ( P2_U4509 , P2_U3369 );
nand NAND2_5205 ( P2_U4510 , P2_R1275_U13 , P2_U3027 );
nand NAND2_5206 ( P2_U4511 , P2_U3026 , P2_U3077 );
nand NAND2_5207 ( P2_U4512 , P2_R1215_U14 , P2_U3025 );
nand NAND2_5208 ( P2_U4513 , P2_U3957 , P2_U4116 );
nand NAND2_5209 ( P2_U4514 , P2_U3657 , P2_U4509 );
nand NAND2_5210 ( P2_U4515 , P2_REG2_REG_22_ , P2_U3020 );
nand NAND2_5211 ( P2_U4516 , P2_REG1_REG_22_ , P2_U3021 );
nand NAND2_5212 ( P2_U4517 , P2_REG0_REG_22_ , P2_U3022 );
nand NAND2_5213 ( P2_U4518 , P2_ADD_1119_U62 , P2_U3019 );
not NOT1_5214 ( P2_U4519 , P2_U3063 );
nand NAND2_5215 ( P2_U4520 , P2_U3035 , P2_U3078 );
nand NAND2_5216 ( P2_U4521 , P2_R1146_U110 , P2_U3931 );
nand NAND2_5217 ( P2_U4522 , P2_R1113_U110 , P2_U3930 );
nand NAND2_5218 ( P2_U4523 , P2_R1131_U14 , P2_U3926 );
nand NAND2_5219 ( P2_U4524 , P2_R1179_U110 , P2_U3941 );
nand NAND2_5220 ( P2_U4525 , P2_R1203_U110 , P2_U3943 );
nand NAND2_5221 ( P2_U4526 , P2_R1164_U14 , P2_U3014 );
nand NAND2_5222 ( P2_U4527 , P2_R1233_U14 , P2_U3922 );
not NOT1_5223 ( P2_U4528 , P2_U3371 );
nand NAND2_5224 ( P2_U4529 , P2_R1275_U78 , P2_U3027 );
nand NAND2_5225 ( P2_U4530 , P2_U3026 , P2_U3063 );
nand NAND2_5226 ( P2_U4531 , P2_R1215_U15 , P2_U3025 );
nand NAND2_5227 ( P2_U4532 , P2_U3956 , P2_U4116 );
nand NAND2_5228 ( P2_U4533 , P2_U3661 , P2_U4528 );
nand NAND2_5229 ( P2_U4534 , P2_REG2_REG_23_ , P2_U3020 );
nand NAND2_5230 ( P2_U4535 , P2_REG1_REG_23_ , P2_U3021 );
nand NAND2_5231 ( P2_U4536 , P2_REG0_REG_23_ , P2_U3022 );
nand NAND2_5232 ( P2_U4537 , P2_ADD_1119_U61 , P2_U3019 );
not NOT1_5233 ( P2_U4538 , P2_U3068 );
nand NAND2_5234 ( P2_U4539 , P2_U3035 , P2_U3077 );
nand NAND2_5235 ( P2_U4540 , P2_R1146_U109 , P2_U3931 );
nand NAND2_5236 ( P2_U4541 , P2_R1113_U109 , P2_U3930 );
nand NAND2_5237 ( P2_U4542 , P2_R1131_U107 , P2_U3926 );
nand NAND2_5238 ( P2_U4543 , P2_R1179_U109 , P2_U3941 );
nand NAND2_5239 ( P2_U4544 , P2_R1203_U109 , P2_U3943 );
nand NAND2_5240 ( P2_U4545 , P2_R1164_U107 , P2_U3014 );
nand NAND2_5241 ( P2_U4546 , P2_R1233_U107 , P2_U3922 );
not NOT1_5242 ( P2_U4547 , P2_U3373 );
nand NAND2_5243 ( P2_U4548 , P2_R1275_U14 , P2_U3027 );
nand NAND2_5244 ( P2_U4549 , P2_U3026 , P2_U3068 );
nand NAND2_5245 ( P2_U4550 , P2_R1215_U108 , P2_U3025 );
nand NAND2_5246 ( P2_U4551 , P2_U3955 , P2_U4116 );
nand NAND2_5247 ( P2_U4552 , P2_U3665 , P2_U4547 );
nand NAND2_5248 ( P2_U4553 , P2_REG2_REG_24_ , P2_U3020 );
nand NAND2_5249 ( P2_U4554 , P2_REG1_REG_24_ , P2_U3021 );
nand NAND2_5250 ( P2_U4555 , P2_REG0_REG_24_ , P2_U3022 );
nand NAND2_5251 ( P2_U4556 , P2_ADD_1119_U60 , P2_U3019 );
not NOT1_5252 ( P2_U4557 , P2_U3067 );
nand NAND2_5253 ( P2_U4558 , P2_U3035 , P2_U3063 );
nand NAND2_5254 ( P2_U4559 , P2_R1146_U14 , P2_U3931 );
nand NAND2_5255 ( P2_U4560 , P2_R1113_U14 , P2_U3930 );
nand NAND2_5256 ( P2_U4561 , P2_R1131_U106 , P2_U3926 );
nand NAND2_5257 ( P2_U4562 , P2_R1179_U14 , P2_U3941 );
nand NAND2_5258 ( P2_U4563 , P2_R1203_U14 , P2_U3943 );
nand NAND2_5259 ( P2_U4564 , P2_R1164_U106 , P2_U3014 );
nand NAND2_5260 ( P2_U4565 , P2_R1233_U106 , P2_U3922 );
not NOT1_5261 ( P2_U4566 , P2_U3375 );
nand NAND2_5262 ( P2_U4567 , P2_R1275_U76 , P2_U3027 );
nand NAND2_5263 ( P2_U4568 , P2_U3026 , P2_U3067 );
nand NAND2_5264 ( P2_U4569 , P2_R1215_U107 , P2_U3025 );
nand NAND2_5265 ( P2_U4570 , P2_U3954 , P2_U4116 );
nand NAND2_5266 ( P2_U4571 , P2_U3669 , P2_U4566 );
nand NAND2_5267 ( P2_U4572 , P2_REG2_REG_25_ , P2_U3020 );
nand NAND2_5268 ( P2_U4573 , P2_REG1_REG_25_ , P2_U3021 );
nand NAND2_5269 ( P2_U4574 , P2_REG0_REG_25_ , P2_U3022 );
nand NAND2_5270 ( P2_U4575 , P2_ADD_1119_U59 , P2_U3019 );
not NOT1_5271 ( P2_U4576 , P2_U3060 );
nand NAND2_5272 ( P2_U4577 , P2_U3035 , P2_U3068 );
nand NAND2_5273 ( P2_U4578 , P2_R1146_U95 , P2_U3931 );
nand NAND2_5274 ( P2_U4579 , P2_R1113_U95 , P2_U3930 );
nand NAND2_5275 ( P2_U4580 , P2_R1131_U105 , P2_U3926 );
nand NAND2_5276 ( P2_U4581 , P2_R1179_U95 , P2_U3941 );
nand NAND2_5277 ( P2_U4582 , P2_R1203_U95 , P2_U3943 );
nand NAND2_5278 ( P2_U4583 , P2_R1164_U105 , P2_U3014 );
nand NAND2_5279 ( P2_U4584 , P2_R1233_U105 , P2_U3922 );
not NOT1_5280 ( P2_U4585 , P2_U3377 );
nand NAND2_5281 ( P2_U4586 , P2_R1275_U15 , P2_U3027 );
nand NAND2_5282 ( P2_U4587 , P2_U3026 , P2_U3060 );
nand NAND2_5283 ( P2_U4588 , P2_R1215_U106 , P2_U3025 );
nand NAND2_5284 ( P2_U4589 , P2_U3953 , P2_U4116 );
nand NAND2_5285 ( P2_U4590 , P2_U3673 , P2_U4585 );
nand NAND2_5286 ( P2_U4591 , P2_REG2_REG_26_ , P2_U3020 );
nand NAND2_5287 ( P2_U4592 , P2_REG1_REG_26_ , P2_U3021 );
nand NAND2_5288 ( P2_U4593 , P2_REG0_REG_26_ , P2_U3022 );
nand NAND2_5289 ( P2_U4594 , P2_ADD_1119_U58 , P2_U3019 );
not NOT1_5290 ( P2_U4595 , P2_U3059 );
nand NAND2_5291 ( P2_U4596 , P2_U3035 , P2_U3067 );
nand NAND2_5292 ( P2_U4597 , P2_R1146_U94 , P2_U3931 );
nand NAND2_5293 ( P2_U4598 , P2_R1113_U94 , P2_U3930 );
nand NAND2_5294 ( P2_U4599 , P2_R1131_U104 , P2_U3926 );
nand NAND2_5295 ( P2_U4600 , P2_R1179_U94 , P2_U3941 );
nand NAND2_5296 ( P2_U4601 , P2_R1203_U94 , P2_U3943 );
nand NAND2_5297 ( P2_U4602 , P2_R1164_U104 , P2_U3014 );
nand NAND2_5298 ( P2_U4603 , P2_R1233_U104 , P2_U3922 );
not NOT1_5299 ( P2_U4604 , P2_U3379 );
nand NAND2_5300 ( P2_U4605 , P2_R1275_U74 , P2_U3027 );
nand NAND2_5301 ( P2_U4606 , P2_U3026 , P2_U3059 );
nand NAND2_5302 ( P2_U4607 , P2_R1215_U105 , P2_U3025 );
nand NAND2_5303 ( P2_U4608 , P2_U3952 , P2_U4116 );
nand NAND2_5304 ( P2_U4609 , P2_U3677 , P2_U4604 );
nand NAND2_5305 ( P2_U4610 , P2_REG2_REG_27_ , P2_U3020 );
nand NAND2_5306 ( P2_U4611 , P2_REG1_REG_27_ , P2_U3021 );
nand NAND2_5307 ( P2_U4612 , P2_REG0_REG_27_ , P2_U3022 );
nand NAND2_5308 ( P2_U4613 , P2_ADD_1119_U57 , P2_U3019 );
not NOT1_5309 ( P2_U4614 , P2_U3055 );
nand NAND2_5310 ( P2_U4615 , P2_U3035 , P2_U3060 );
nand NAND2_5311 ( P2_U4616 , P2_R1146_U108 , P2_U3931 );
nand NAND2_5312 ( P2_U4617 , P2_R1113_U108 , P2_U3930 );
nand NAND2_5313 ( P2_U4618 , P2_R1131_U15 , P2_U3926 );
nand NAND2_5314 ( P2_U4619 , P2_R1179_U108 , P2_U3941 );
nand NAND2_5315 ( P2_U4620 , P2_R1203_U108 , P2_U3943 );
nand NAND2_5316 ( P2_U4621 , P2_R1164_U15 , P2_U3014 );
nand NAND2_5317 ( P2_U4622 , P2_R1233_U15 , P2_U3922 );
not NOT1_5318 ( P2_U4623 , P2_U3381 );
nand NAND2_5319 ( P2_U4624 , P2_R1275_U16 , P2_U3027 );
nand NAND2_5320 ( P2_U4625 , P2_U3026 , P2_U3055 );
nand NAND2_5321 ( P2_U4626 , P2_R1215_U16 , P2_U3025 );
nand NAND2_5322 ( P2_U4627 , P2_U3951 , P2_U4116 );
nand NAND2_5323 ( P2_U4628 , P2_U3681 , P2_U4623 );
nand NAND2_5324 ( P2_U4629 , P2_REG2_REG_28_ , P2_U3020 );
nand NAND2_5325 ( P2_U4630 , P2_REG1_REG_28_ , P2_U3021 );
nand NAND2_5326 ( P2_U4631 , P2_REG0_REG_28_ , P2_U3022 );
nand NAND2_5327 ( P2_U4632 , P2_ADD_1119_U56 , P2_U3019 );
not NOT1_5328 ( P2_U4633 , P2_U3056 );
nand NAND2_5329 ( P2_U4634 , P2_U3035 , P2_U3059 );
nand NAND2_5330 ( P2_U4635 , P2_R1146_U15 , P2_U3931 );
nand NAND2_5331 ( P2_U4636 , P2_R1113_U15 , P2_U3930 );
nand NAND2_5332 ( P2_U4637 , P2_R1131_U103 , P2_U3926 );
nand NAND2_5333 ( P2_U4638 , P2_R1179_U15 , P2_U3941 );
nand NAND2_5334 ( P2_U4639 , P2_R1203_U15 , P2_U3943 );
nand NAND2_5335 ( P2_U4640 , P2_R1164_U103 , P2_U3014 );
nand NAND2_5336 ( P2_U4641 , P2_R1233_U103 , P2_U3922 );
not NOT1_5337 ( P2_U4642 , P2_U3383 );
nand NAND2_5338 ( P2_U4643 , P2_R1275_U72 , P2_U3027 );
nand NAND2_5339 ( P2_U4644 , P2_U3026 , P2_U3056 );
nand NAND2_5340 ( P2_U4645 , P2_R1215_U104 , P2_U3025 );
nand NAND2_5341 ( P2_U4646 , P2_U3950 , P2_U4116 );
nand NAND2_5342 ( P2_U4647 , P2_U3685 , P2_U4642 );
nand NAND2_5343 ( P2_U4648 , P2_ADD_1119_U5 , P2_U3019 );
nand NAND2_5344 ( P2_U4649 , P2_REG2_REG_29_ , P2_U3020 );
nand NAND2_5345 ( P2_U4650 , P2_REG1_REG_29_ , P2_U3021 );
nand NAND2_5346 ( P2_U4651 , P2_REG0_REG_29_ , P2_U3022 );
not NOT1_5347 ( P2_U4652 , P2_U3057 );
nand NAND2_5348 ( P2_U4653 , P2_U3035 , P2_U3055 );
nand NAND2_5349 ( P2_U4654 , P2_R1146_U93 , P2_U3931 );
nand NAND2_5350 ( P2_U4655 , P2_R1113_U93 , P2_U3930 );
nand NAND2_5351 ( P2_U4656 , P2_R1131_U102 , P2_U3926 );
nand NAND2_5352 ( P2_U4657 , P2_R1179_U93 , P2_U3941 );
nand NAND2_5353 ( P2_U4658 , P2_R1203_U93 , P2_U3943 );
nand NAND2_5354 ( P2_U4659 , P2_R1164_U102 , P2_U3014 );
nand NAND2_5355 ( P2_U4660 , P2_R1233_U102 , P2_U3922 );
not NOT1_5356 ( P2_U4661 , P2_U3385 );
nand NAND2_5357 ( P2_U4662 , P2_R1275_U17 , P2_U3027 );
nand NAND2_5358 ( P2_U4663 , P2_U3026 , P2_U3057 );
nand NAND2_5359 ( P2_U4664 , P2_R1215_U103 , P2_U3025 );
nand NAND2_5360 ( P2_U4665 , P2_U3949 , P2_U4116 );
nand NAND2_5361 ( P2_U4666 , P2_U3688 , P2_U4661 );
nand NAND2_5362 ( P2_U4667 , P2_REG2_REG_30_ , P2_U3020 );
nand NAND2_5363 ( P2_U4668 , P2_REG1_REG_30_ , P2_U3021 );
nand NAND2_5364 ( P2_U4669 , P2_REG0_REG_30_ , P2_U3022 );
not NOT1_5365 ( P2_U4670 , P2_U3061 );
nand NAND2_5366 ( P2_U4671 , P2_U5683 , P2_U3331 );
nand NAND2_5367 ( P2_U4672 , P2_U3347 , P2_U4671 );
nand NAND2_5368 ( P2_U4673 , P2_U3689 , P2_U3061 );
nand NAND2_5369 ( P2_U4674 , P2_U3035 , P2_U3056 );
nand NAND2_5370 ( P2_U4675 , P2_R1146_U16 , P2_U3931 );
nand NAND2_5371 ( P2_U4676 , P2_R1113_U16 , P2_U3930 );
nand NAND2_5372 ( P2_U4677 , P2_R1131_U101 , P2_U3926 );
nand NAND2_5373 ( P2_U4678 , P2_R1179_U16 , P2_U3941 );
nand NAND2_5374 ( P2_U4679 , P2_R1203_U16 , P2_U3943 );
nand NAND2_5375 ( P2_U4680 , P2_R1164_U101 , P2_U3014 );
nand NAND2_5376 ( P2_U4681 , P2_R1233_U101 , P2_U3922 );
not NOT1_5377 ( P2_U4682 , P2_U3387 );
nand NAND2_5378 ( P2_U4683 , P2_R1275_U70 , P2_U3027 );
nand NAND2_5379 ( P2_U4684 , P2_R1215_U102 , P2_U3025 );
nand NAND2_5380 ( P2_U4685 , P2_U3960 , P2_U4116 );
nand NAND2_5381 ( P2_U4686 , P2_U3693 , P2_U4682 );
nand NAND2_5382 ( P2_U4687 , P2_REG2_REG_31_ , P2_U3020 );
nand NAND2_5383 ( P2_U4688 , P2_REG1_REG_31_ , P2_U3021 );
nand NAND2_5384 ( P2_U4689 , P2_REG0_REG_31_ , P2_U3022 );
not NOT1_5385 ( P2_U4690 , P2_U3058 );
nand NAND2_5386 ( P2_U4691 , P2_R1275_U19 , P2_U3027 );
nand NAND2_5387 ( P2_U4692 , P2_U3959 , P2_U4116 );
nand NAND3_5388 ( P2_U4693 , P2_U4692 , P2_U3913 , P2_U4691 );
nand NAND2_5389 ( P2_U4694 , P2_R1275_U68 , P2_U3027 );
nand NAND2_5390 ( P2_U4695 , P2_U3958 , P2_U4116 );
nand NAND3_5391 ( P2_U4696 , P2_U4695 , P2_U3913 , P2_U4694 );
nand NAND2_5392 ( P2_U4697 , P2_U3696 , P2_U3016 );
nand NAND2_5393 ( P2_U4698 , P2_U3393 , P2_U4697 );
nand NAND2_5394 ( P2_U4699 , P2_U3921 , P2_U3418 );
not NOT1_5395 ( P2_U4700 , P2_U3398 );
nand NAND2_5396 ( P2_U4701 , P2_U3037 , P2_U3080 );
nand NAND2_5397 ( P2_U4702 , P2_U3034 , P2_R1215_U96 );
nand NAND2_5398 ( P2_U4703 , P2_U3033 , P2_REG3_REG_0_ );
nand NAND2_5399 ( P2_U4704 , P2_U3032 , P2_U3427 );
nand NAND2_5400 ( P2_U4705 , P2_U3031 , P2_U3427 );
nand NAND2_5401 ( P2_U4706 , P2_U3037 , P2_U3070 );
nand NAND2_5402 ( P2_U4707 , P2_U3034 , P2_R1215_U95 );
nand NAND2_5403 ( P2_U4708 , P2_U3033 , P2_REG3_REG_1_ );
nand NAND2_5404 ( P2_U4709 , P2_U3032 , P2_U3432 );
nand NAND2_5405 ( P2_U4710 , P2_U3031 , P2_R1275_U55 );
nand NAND2_5406 ( P2_U4711 , P2_U3037 , P2_U3066 );
nand NAND2_5407 ( P2_U4712 , P2_U3034 , P2_R1215_U17 );
nand NAND2_5408 ( P2_U4713 , P2_U3033 , P2_REG3_REG_2_ );
nand NAND2_5409 ( P2_U4714 , P2_U3032 , P2_U3435 );
nand NAND2_5410 ( P2_U4715 , P2_U3031 , P2_R1275_U18 );
nand NAND2_5411 ( P2_U4716 , P2_U3037 , P2_U3062 );
nand NAND2_5412 ( P2_U4717 , P2_U3034 , P2_R1215_U101 );
nand NAND2_5413 ( P2_U4718 , P2_U3033 , P2_ADD_1119_U4 );
nand NAND2_5414 ( P2_U4719 , P2_U3032 , P2_U3438 );
nand NAND2_5415 ( P2_U4720 , P2_U3031 , P2_R1275_U20 );
nand NAND2_5416 ( P2_U4721 , P2_U3037 , P2_U3069 );
nand NAND2_5417 ( P2_U4722 , P2_U3034 , P2_R1215_U100 );
nand NAND2_5418 ( P2_U4723 , P2_U3033 , P2_ADD_1119_U55 );
nand NAND2_5419 ( P2_U4724 , P2_U3032 , P2_U3441 );
nand NAND2_5420 ( P2_U4725 , P2_U3031 , P2_R1275_U21 );
nand NAND2_5421 ( P2_U4726 , P2_U3037 , P2_U3073 );
nand NAND2_5422 ( P2_U4727 , P2_U3034 , P2_R1215_U18 );
nand NAND2_5423 ( P2_U4728 , P2_U3033 , P2_ADD_1119_U54 );
nand NAND2_5424 ( P2_U4729 , P2_U3032 , P2_U3444 );
nand NAND2_5425 ( P2_U4730 , P2_U3031 , P2_R1275_U65 );
nand NAND2_5426 ( P2_U4731 , P2_U3037 , P2_U3072 );
nand NAND2_5427 ( P2_U4732 , P2_U3034 , P2_R1215_U99 );
nand NAND2_5428 ( P2_U4733 , P2_U3033 , P2_ADD_1119_U53 );
nand NAND2_5429 ( P2_U4734 , P2_U3032 , P2_U3447 );
nand NAND2_5430 ( P2_U4735 , P2_U3031 , P2_R1275_U22 );
nand NAND2_5431 ( P2_U4736 , P2_U3037 , P2_U3086 );
nand NAND2_5432 ( P2_U4737 , P2_U3034 , P2_R1215_U19 );
nand NAND2_5433 ( P2_U4738 , P2_U3033 , P2_ADD_1119_U52 );
nand NAND2_5434 ( P2_U4739 , P2_U3032 , P2_U3450 );
nand NAND2_5435 ( P2_U4740 , P2_U3031 , P2_R1275_U23 );
nand NAND2_5436 ( P2_U4741 , P2_U3037 , P2_U3085 );
nand NAND2_5437 ( P2_U4742 , P2_U3034 , P2_R1215_U98 );
nand NAND2_5438 ( P2_U4743 , P2_U3033 , P2_ADD_1119_U51 );
nand NAND2_5439 ( P2_U4744 , P2_U3032 , P2_U3453 );
nand NAND2_5440 ( P2_U4745 , P2_U3031 , P2_R1275_U24 );
nand NAND2_5441 ( P2_U4746 , P2_U3037 , P2_U3064 );
nand NAND2_5442 ( P2_U4747 , P2_U3034 , P2_R1215_U97 );
nand NAND2_5443 ( P2_U4748 , P2_U3033 , P2_ADD_1119_U50 );
nand NAND2_5444 ( P2_U4749 , P2_U3032 , P2_U3456 );
nand NAND2_5445 ( P2_U4750 , P2_U3031 , P2_R1275_U63 );
nand NAND2_5446 ( P2_U4751 , P2_U3037 , P2_U3065 );
nand NAND2_5447 ( P2_U4752 , P2_U3034 , P2_R1215_U11 );
nand NAND2_5448 ( P2_U4753 , P2_U3033 , P2_ADD_1119_U74 );
nand NAND2_5449 ( P2_U4754 , P2_U3032 , P2_U3459 );
nand NAND2_5450 ( P2_U4755 , P2_U3031 , P2_R1275_U6 );
nand NAND2_5451 ( P2_U4756 , P2_U3037 , P2_U3074 );
nand NAND2_5452 ( P2_U4757 , P2_U3034 , P2_R1215_U115 );
nand NAND2_5453 ( P2_U4758 , P2_U3033 , P2_ADD_1119_U73 );
nand NAND2_5454 ( P2_U4759 , P2_U3032 , P2_U3462 );
nand NAND2_5455 ( P2_U4760 , P2_U3031 , P2_R1275_U7 );
nand NAND2_5456 ( P2_U4761 , P2_U3037 , P2_U3082 );
nand NAND2_5457 ( P2_U4762 , P2_U3034 , P2_R1215_U114 );
nand NAND2_5458 ( P2_U4763 , P2_U3033 , P2_ADD_1119_U72 );
nand NAND2_5459 ( P2_U4764 , P2_U3032 , P2_U3465 );
nand NAND2_5460 ( P2_U4765 , P2_U3031 , P2_R1275_U8 );
nand NAND2_5461 ( P2_U4766 , P2_U3037 , P2_U3081 );
nand NAND2_5462 ( P2_U4767 , P2_U3034 , P2_R1215_U12 );
nand NAND2_5463 ( P2_U4768 , P2_U3033 , P2_ADD_1119_U71 );
nand NAND2_5464 ( P2_U4769 , P2_U3032 , P2_U3468 );
nand NAND2_5465 ( P2_U4770 , P2_U3031 , P2_R1275_U86 );
nand NAND2_5466 ( P2_U4771 , P2_U3037 , P2_U3076 );
nand NAND2_5467 ( P2_U4772 , P2_U3034 , P2_R1215_U113 );
nand NAND2_5468 ( P2_U4773 , P2_U3033 , P2_ADD_1119_U70 );
nand NAND2_5469 ( P2_U4774 , P2_U3032 , P2_U3471 );
nand NAND2_5470 ( P2_U4775 , P2_U3031 , P2_R1275_U9 );
nand NAND2_5471 ( P2_U4776 , P2_U3037 , P2_U3075 );
nand NAND2_5472 ( P2_U4777 , P2_U3034 , P2_R1215_U112 );
nand NAND2_5473 ( P2_U4778 , P2_U3033 , P2_ADD_1119_U69 );
nand NAND2_5474 ( P2_U4779 , P2_U3032 , P2_U3474 );
nand NAND2_5475 ( P2_U4780 , P2_U3031 , P2_R1275_U10 );
nand NAND2_5476 ( P2_U4781 , P2_U3037 , P2_U3071 );
nand NAND2_5477 ( P2_U4782 , P2_U3034 , P2_R1215_U111 );
nand NAND2_5478 ( P2_U4783 , P2_U3033 , P2_ADD_1119_U68 );
nand NAND2_5479 ( P2_U4784 , P2_U3032 , P2_U3477 );
nand NAND2_5480 ( P2_U4785 , P2_U3031 , P2_R1275_U11 );
nand NAND2_5481 ( P2_U4786 , P2_U3037 , P2_U3084 );
nand NAND2_5482 ( P2_U4787 , P2_U3034 , P2_R1215_U13 );
nand NAND2_5483 ( P2_U4788 , P2_U3033 , P2_ADD_1119_U67 );
nand NAND2_5484 ( P2_U4789 , P2_U3032 , P2_U3480 );
nand NAND2_5485 ( P2_U4790 , P2_U3031 , P2_R1275_U84 );
nand NAND2_5486 ( P2_U4791 , P2_U3037 , P2_U3083 );
nand NAND2_5487 ( P2_U4792 , P2_U3034 , P2_R1215_U110 );
nand NAND2_5488 ( P2_U4793 , P2_U3033 , P2_ADD_1119_U66 );
nand NAND2_5489 ( P2_U4794 , P2_U3032 , P2_U3483 );
nand NAND2_5490 ( P2_U4795 , P2_U3031 , P2_R1275_U12 );
nand NAND2_5491 ( P2_U4796 , P2_U3037 , P2_U3078 );
nand NAND2_5492 ( P2_U4797 , P2_U3034 , P2_R1215_U109 );
nand NAND2_5493 ( P2_U4798 , P2_U3033 , P2_ADD_1119_U65 );
nand NAND2_5494 ( P2_U4799 , P2_U3032 , P2_U3485 );
nand NAND2_5495 ( P2_U4800 , P2_U3031 , P2_R1275_U82 );
nand NAND2_5496 ( P2_U4801 , P2_U3037 , P2_U3077 );
nand NAND2_5497 ( P2_U4802 , P2_U3034 , P2_R1215_U14 );
nand NAND2_5498 ( P2_U4803 , P2_U3033 , P2_ADD_1119_U64 );
nand NAND2_5499 ( P2_U4804 , P2_U3032 , P2_U3957 );
nand NAND2_5500 ( P2_U4805 , P2_U3031 , P2_R1275_U13 );
nand NAND2_5501 ( P2_U4806 , P2_U3037 , P2_U3063 );
nand NAND2_5502 ( P2_U4807 , P2_U3034 , P2_R1215_U15 );
nand NAND2_5503 ( P2_U4808 , P2_U3033 , P2_ADD_1119_U63 );
nand NAND2_5504 ( P2_U4809 , P2_U3032 , P2_U3956 );
nand NAND2_5505 ( P2_U4810 , P2_U3031 , P2_R1275_U78 );
nand NAND2_5506 ( P2_U4811 , P2_U3037 , P2_U3068 );
nand NAND2_5507 ( P2_U4812 , P2_U3034 , P2_R1215_U108 );
nand NAND2_5508 ( P2_U4813 , P2_U3033 , P2_ADD_1119_U62 );
nand NAND2_5509 ( P2_U4814 , P2_U3032 , P2_U3955 );
nand NAND2_5510 ( P2_U4815 , P2_U3031 , P2_R1275_U14 );
nand NAND2_5511 ( P2_U4816 , P2_U3037 , P2_U3067 );
nand NAND2_5512 ( P2_U4817 , P2_U3034 , P2_R1215_U107 );
nand NAND2_5513 ( P2_U4818 , P2_U3033 , P2_ADD_1119_U61 );
nand NAND2_5514 ( P2_U4819 , P2_U3032 , P2_U3954 );
nand NAND2_5515 ( P2_U4820 , P2_U3031 , P2_R1275_U76 );
nand NAND2_5516 ( P2_U4821 , P2_U3037 , P2_U3060 );
nand NAND2_5517 ( P2_U4822 , P2_U3034 , P2_R1215_U106 );
nand NAND2_5518 ( P2_U4823 , P2_U3033 , P2_ADD_1119_U60 );
nand NAND2_5519 ( P2_U4824 , P2_U3032 , P2_U3953 );
nand NAND2_5520 ( P2_U4825 , P2_U3031 , P2_R1275_U15 );
nand NAND2_5521 ( P2_U4826 , P2_U3037 , P2_U3059 );
nand NAND2_5522 ( P2_U4827 , P2_U3034 , P2_R1215_U105 );
nand NAND2_5523 ( P2_U4828 , P2_U3033 , P2_ADD_1119_U59 );
nand NAND2_5524 ( P2_U4829 , P2_U3032 , P2_U3952 );
nand NAND2_5525 ( P2_U4830 , P2_U3031 , P2_R1275_U74 );
nand NAND2_5526 ( P2_U4831 , P2_U3037 , P2_U3055 );
nand NAND2_5527 ( P2_U4832 , P2_U3034 , P2_R1215_U16 );
nand NAND2_5528 ( P2_U4833 , P2_U3033 , P2_ADD_1119_U58 );
nand NAND2_5529 ( P2_U4834 , P2_U3032 , P2_U3951 );
nand NAND2_5530 ( P2_U4835 , P2_U3031 , P2_R1275_U16 );
nand NAND2_5531 ( P2_U4836 , P2_U3037 , P2_U3056 );
nand NAND2_5532 ( P2_U4837 , P2_U3034 , P2_R1215_U104 );
nand NAND2_5533 ( P2_U4838 , P2_U3033 , P2_ADD_1119_U57 );
nand NAND2_5534 ( P2_U4839 , P2_U3032 , P2_U3950 );
nand NAND2_5535 ( P2_U4840 , P2_U3031 , P2_R1275_U72 );
nand NAND2_5536 ( P2_U4841 , P2_U3037 , P2_U3057 );
nand NAND2_5537 ( P2_U4842 , P2_U3034 , P2_R1215_U103 );
nand NAND2_5538 ( P2_U4843 , P2_U3033 , P2_ADD_1119_U56 );
nand NAND2_5539 ( P2_U4844 , P2_U3032 , P2_U3949 );
nand NAND2_5540 ( P2_U4845 , P2_U3031 , P2_R1275_U17 );
nand NAND2_5541 ( P2_U4846 , P2_U3034 , P2_R1215_U102 );
nand NAND2_5542 ( P2_U4847 , P2_U3033 , P2_ADD_1119_U5 );
nand NAND2_5543 ( P2_U4848 , P2_U3032 , P2_U3960 );
nand NAND2_5544 ( P2_U4849 , P2_U3031 , P2_R1275_U70 );
nand NAND2_5545 ( P2_U4850 , P2_U3032 , P2_U3959 );
nand NAND2_5546 ( P2_U4851 , P2_U3031 , P2_R1275_U19 );
nand NAND2_5547 ( P2_U4852 , P2_U3032 , P2_U3958 );
nand NAND2_5548 ( P2_U4853 , P2_U3031 , P2_R1275_U68 );
nand NAND5_5549 ( P2_U4854 , P2_U3755 , P2_U3395 , P2_U3051 , P2_U4700 , P2_U3393 );
nand NAND2_5550 ( P2_U4855 , P2_R1170_U13 , P2_U3043 );
nand NAND2_5551 ( P2_U4856 , P2_U3041 , P2_U3424 );
nand NAND2_5552 ( P2_U4857 , P2_R1209_U13 , P2_U3039 );
nand NAND3_5553 ( P2_U4858 , P2_U4856 , P2_U4855 , P2_U4857 );
nand NAND2_5554 ( P2_U4859 , P2_R1170_U13 , P2_U3018 );
nand NAND2_5555 ( P2_U4860 , P2_U3017 , P2_R1209_U13 );
nand NAND2_5556 ( P2_U4861 , P2_U5683 , P2_U3424 );
nand NAND3_5557 ( P2_U4862 , P2_U4860 , P2_U4859 , P2_U4861 );
not NOT1_5558 ( P2_U4863 , P2_U3401 );
nand NAND2_5559 ( P2_U4864 , P2_U3045 , P2_U4858 );
nand NAND2_5560 ( P2_U4865 , P2_U3947 , P2_U4862 );
nand NAND2_5561 ( P2_U4866 , P2_U3044 , P2_R1170_U13 );
nand NAND2_5562 ( P2_U4867 , P2_REG3_REG_19_ , P2_U3088 );
nand NAND2_5563 ( P2_U4868 , P2_U3042 , P2_U3424 );
nand NAND2_5564 ( P2_U4869 , P2_U3040 , P2_R1209_U13 );
nand NAND2_5565 ( P2_U4870 , P2_ADDR_REG_19_ , P2_U4863 );
nand NAND2_5566 ( P2_U4871 , P2_R1170_U75 , P2_U3043 );
nand NAND2_5567 ( P2_U4872 , P2_U3041 , P2_U3482 );
nand NAND2_5568 ( P2_U4873 , P2_R1209_U75 , P2_U3039 );
nand NAND3_5569 ( P2_U4874 , P2_U4872 , P2_U4871 , P2_U4873 );
nand NAND2_5570 ( P2_U4875 , P2_R1170_U75 , P2_U3018 );
nand NAND2_5571 ( P2_U4876 , P2_R1209_U75 , P2_U3017 );
nand NAND2_5572 ( P2_U4877 , P2_U5683 , P2_U3482 );
nand NAND3_5573 ( P2_U4878 , P2_U4876 , P2_U4875 , P2_U4877 );
nand NAND2_5574 ( P2_U4879 , P2_U3045 , P2_U4874 );
nand NAND2_5575 ( P2_U4880 , P2_U3947 , P2_U4878 );
nand NAND2_5576 ( P2_U4881 , P2_R1170_U75 , P2_U3044 );
nand NAND2_5577 ( P2_U4882 , P2_REG3_REG_18_ , P2_U3088 );
nand NAND2_5578 ( P2_U4883 , P2_U3042 , P2_U3482 );
nand NAND2_5579 ( P2_U4884 , P2_R1209_U75 , P2_U3040 );
nand NAND2_5580 ( P2_U4885 , P2_ADDR_REG_18_ , P2_U4863 );
nand NAND2_5581 ( P2_U4886 , P2_R1170_U12 , P2_U3043 );
nand NAND2_5582 ( P2_U4887 , P2_U3041 , P2_U3479 );
nand NAND2_5583 ( P2_U4888 , P2_R1209_U12 , P2_U3039 );
nand NAND3_5584 ( P2_U4889 , P2_U4887 , P2_U4886 , P2_U4888 );
nand NAND2_5585 ( P2_U4890 , P2_R1170_U12 , P2_U3018 );
nand NAND2_5586 ( P2_U4891 , P2_R1209_U12 , P2_U3017 );
nand NAND2_5587 ( P2_U4892 , P2_U5683 , P2_U3479 );
nand NAND3_5588 ( P2_U4893 , P2_U4891 , P2_U4890 , P2_U4892 );
nand NAND2_5589 ( P2_U4894 , P2_U3045 , P2_U4889 );
nand NAND2_5590 ( P2_U4895 , P2_U3947 , P2_U4893 );
nand NAND2_5591 ( P2_U4896 , P2_R1170_U12 , P2_U3044 );
nand NAND2_5592 ( P2_U4897 , P2_REG3_REG_17_ , P2_U3088 );
nand NAND2_5593 ( P2_U4898 , P2_U3042 , P2_U3479 );
nand NAND2_5594 ( P2_U4899 , P2_R1209_U12 , P2_U3040 );
nand NAND2_5595 ( P2_U4900 , P2_ADDR_REG_17_ , P2_U4863 );
nand NAND2_5596 ( P2_U4901 , P2_R1170_U76 , P2_U3043 );
nand NAND2_5597 ( P2_U4902 , P2_U3041 , P2_U3476 );
nand NAND2_5598 ( P2_U4903 , P2_R1209_U76 , P2_U3039 );
nand NAND3_5599 ( P2_U4904 , P2_U4902 , P2_U4901 , P2_U4903 );
nand NAND2_5600 ( P2_U4905 , P2_R1170_U76 , P2_U3018 );
nand NAND2_5601 ( P2_U4906 , P2_R1209_U76 , P2_U3017 );
nand NAND2_5602 ( P2_U4907 , P2_U5683 , P2_U3476 );
nand NAND3_5603 ( P2_U4908 , P2_U4906 , P2_U4905 , P2_U4907 );
nand NAND2_5604 ( P2_U4909 , P2_U3045 , P2_U4904 );
nand NAND2_5605 ( P2_U4910 , P2_U3947 , P2_U4908 );
nand NAND2_5606 ( P2_U4911 , P2_R1170_U76 , P2_U3044 );
nand NAND2_5607 ( P2_U4912 , P2_REG3_REG_16_ , P2_U3088 );
nand NAND2_5608 ( P2_U4913 , P2_U3042 , P2_U3476 );
nand NAND2_5609 ( P2_U4914 , P2_R1209_U76 , P2_U3040 );
nand NAND2_5610 ( P2_U4915 , P2_ADDR_REG_16_ , P2_U4863 );
nand NAND2_5611 ( P2_U4916 , P2_R1170_U77 , P2_U3043 );
nand NAND2_5612 ( P2_U4917 , P2_U3041 , P2_U3473 );
nand NAND2_5613 ( P2_U4918 , P2_R1209_U77 , P2_U3039 );
nand NAND3_5614 ( P2_U4919 , P2_U4917 , P2_U4916 , P2_U4918 );
nand NAND2_5615 ( P2_U4920 , P2_R1170_U77 , P2_U3018 );
nand NAND2_5616 ( P2_U4921 , P2_R1209_U77 , P2_U3017 );
nand NAND2_5617 ( P2_U4922 , P2_U5683 , P2_U3473 );
nand NAND3_5618 ( P2_U4923 , P2_U4921 , P2_U4920 , P2_U4922 );
nand NAND2_5619 ( P2_U4924 , P2_U3045 , P2_U4919 );
nand NAND2_5620 ( P2_U4925 , P2_U3947 , P2_U4923 );
nand NAND2_5621 ( P2_U4926 , P2_R1170_U77 , P2_U3044 );
nand NAND2_5622 ( P2_U4927 , P2_REG3_REG_15_ , P2_U3088 );
nand NAND2_5623 ( P2_U4928 , P2_U3042 , P2_U3473 );
nand NAND2_5624 ( P2_U4929 , P2_R1209_U77 , P2_U3040 );
nand NAND2_5625 ( P2_U4930 , P2_ADDR_REG_15_ , P2_U4863 );
nand NAND2_5626 ( P2_U4931 , P2_R1170_U78 , P2_U3043 );
nand NAND2_5627 ( P2_U4932 , P2_U3041 , P2_U3470 );
nand NAND2_5628 ( P2_U4933 , P2_R1209_U78 , P2_U3039 );
nand NAND3_5629 ( P2_U4934 , P2_U4932 , P2_U4931 , P2_U4933 );
nand NAND2_5630 ( P2_U4935 , P2_R1170_U78 , P2_U3018 );
nand NAND2_5631 ( P2_U4936 , P2_R1209_U78 , P2_U3017 );
nand NAND2_5632 ( P2_U4937 , P2_U5683 , P2_U3470 );
nand NAND3_5633 ( P2_U4938 , P2_U4936 , P2_U4935 , P2_U4937 );
nand NAND2_5634 ( P2_U4939 , P2_U3045 , P2_U4934 );
nand NAND2_5635 ( P2_U4940 , P2_U3947 , P2_U4938 );
nand NAND2_5636 ( P2_U4941 , P2_R1170_U78 , P2_U3044 );
nand NAND2_5637 ( P2_U4942 , P2_REG3_REG_14_ , P2_U3088 );
nand NAND2_5638 ( P2_U4943 , P2_U3042 , P2_U3470 );
nand NAND2_5639 ( P2_U4944 , P2_R1209_U78 , P2_U3040 );
nand NAND2_5640 ( P2_U4945 , P2_ADDR_REG_14_ , P2_U4863 );
nand NAND2_5641 ( P2_U4946 , P2_R1170_U11 , P2_U3043 );
nand NAND2_5642 ( P2_U4947 , P2_U3041 , P2_U3467 );
nand NAND2_5643 ( P2_U4948 , P2_R1209_U11 , P2_U3039 );
nand NAND3_5644 ( P2_U4949 , P2_U4947 , P2_U4946 , P2_U4948 );
nand NAND2_5645 ( P2_U4950 , P2_R1170_U11 , P2_U3018 );
nand NAND2_5646 ( P2_U4951 , P2_R1209_U11 , P2_U3017 );
nand NAND2_5647 ( P2_U4952 , P2_U5683 , P2_U3467 );
nand NAND3_5648 ( P2_U4953 , P2_U4951 , P2_U4950 , P2_U4952 );
nand NAND2_5649 ( P2_U4954 , P2_U3045 , P2_U4949 );
nand NAND2_5650 ( P2_U4955 , P2_U3947 , P2_U4953 );
nand NAND2_5651 ( P2_U4956 , P2_R1170_U11 , P2_U3044 );
nand NAND2_5652 ( P2_U4957 , P2_REG3_REG_13_ , P2_U3088 );
nand NAND2_5653 ( P2_U4958 , P2_U3042 , P2_U3467 );
nand NAND2_5654 ( P2_U4959 , P2_R1209_U11 , P2_U3040 );
nand NAND2_5655 ( P2_U4960 , P2_ADDR_REG_13_ , P2_U4863 );
nand NAND2_5656 ( P2_U4961 , P2_R1170_U79 , P2_U3043 );
nand NAND2_5657 ( P2_U4962 , P2_U3041 , P2_U3464 );
nand NAND2_5658 ( P2_U4963 , P2_R1209_U79 , P2_U3039 );
nand NAND3_5659 ( P2_U4964 , P2_U4962 , P2_U4961 , P2_U4963 );
nand NAND2_5660 ( P2_U4965 , P2_R1170_U79 , P2_U3018 );
nand NAND2_5661 ( P2_U4966 , P2_R1209_U79 , P2_U3017 );
nand NAND2_5662 ( P2_U4967 , P2_U5683 , P2_U3464 );
nand NAND3_5663 ( P2_U4968 , P2_U4966 , P2_U4965 , P2_U4967 );
nand NAND2_5664 ( P2_U4969 , P2_U3045 , P2_U4964 );
nand NAND2_5665 ( P2_U4970 , P2_U3947 , P2_U4968 );
nand NAND2_5666 ( P2_U4971 , P2_R1170_U79 , P2_U3044 );
nand NAND2_5667 ( P2_U4972 , P2_REG3_REG_12_ , P2_U3088 );
nand NAND2_5668 ( P2_U4973 , P2_U3042 , P2_U3464 );
nand NAND2_5669 ( P2_U4974 , P2_R1209_U79 , P2_U3040 );
nand NAND2_5670 ( P2_U4975 , P2_ADDR_REG_12_ , P2_U4863 );
nand NAND2_5671 ( P2_U4976 , P2_R1170_U80 , P2_U3043 );
nand NAND2_5672 ( P2_U4977 , P2_U3041 , P2_U3461 );
nand NAND2_5673 ( P2_U4978 , P2_R1209_U80 , P2_U3039 );
nand NAND3_5674 ( P2_U4979 , P2_U4977 , P2_U4976 , P2_U4978 );
nand NAND2_5675 ( P2_U4980 , P2_R1170_U80 , P2_U3018 );
nand NAND2_5676 ( P2_U4981 , P2_R1209_U80 , P2_U3017 );
nand NAND2_5677 ( P2_U4982 , P2_U5683 , P2_U3461 );
nand NAND3_5678 ( P2_U4983 , P2_U4981 , P2_U4980 , P2_U4982 );
nand NAND2_5679 ( P2_U4984 , P2_U3045 , P2_U4979 );
nand NAND2_5680 ( P2_U4985 , P2_U3947 , P2_U4983 );
nand NAND2_5681 ( P2_U4986 , P2_R1170_U80 , P2_U3044 );
nand NAND2_5682 ( P2_U4987 , P2_REG3_REG_11_ , P2_U3088 );
nand NAND2_5683 ( P2_U4988 , P2_U3042 , P2_U3461 );
nand NAND2_5684 ( P2_U4989 , P2_R1209_U80 , P2_U3040 );
nand NAND2_5685 ( P2_U4990 , P2_ADDR_REG_11_ , P2_U4863 );
nand NAND2_5686 ( P2_U4991 , P2_R1170_U10 , P2_U3043 );
nand NAND2_5687 ( P2_U4992 , P2_U3041 , P2_U3458 );
nand NAND2_5688 ( P2_U4993 , P2_R1209_U10 , P2_U3039 );
nand NAND3_5689 ( P2_U4994 , P2_U4992 , P2_U4991 , P2_U4993 );
nand NAND2_5690 ( P2_U4995 , P2_R1170_U10 , P2_U3018 );
nand NAND2_5691 ( P2_U4996 , P2_R1209_U10 , P2_U3017 );
nand NAND2_5692 ( P2_U4997 , P2_U5683 , P2_U3458 );
nand NAND3_5693 ( P2_U4998 , P2_U4996 , P2_U4995 , P2_U4997 );
nand NAND2_5694 ( P2_U4999 , P2_U3045 , P2_U4994 );
nand NAND2_5695 ( P2_U5000 , P2_U3947 , P2_U4998 );
nand NAND2_5696 ( P2_U5001 , P2_R1170_U10 , P2_U3044 );
nand NAND2_5697 ( P2_U5002 , P2_REG3_REG_10_ , P2_U3088 );
nand NAND2_5698 ( P2_U5003 , P2_U3042 , P2_U3458 );
nand NAND2_5699 ( P2_U5004 , P2_R1209_U10 , P2_U3040 );
nand NAND2_5700 ( P2_U5005 , P2_ADDR_REG_10_ , P2_U4863 );
nand NAND2_5701 ( P2_U5006 , P2_R1170_U70 , P2_U3043 );
nand NAND2_5702 ( P2_U5007 , P2_U3041 , P2_U3455 );
nand NAND2_5703 ( P2_U5008 , P2_R1209_U70 , P2_U3039 );
nand NAND3_5704 ( P2_U5009 , P2_U5007 , P2_U5006 , P2_U5008 );
nand NAND2_5705 ( P2_U5010 , P2_R1170_U70 , P2_U3018 );
nand NAND2_5706 ( P2_U5011 , P2_R1209_U70 , P2_U3017 );
nand NAND2_5707 ( P2_U5012 , P2_U5683 , P2_U3455 );
nand NAND3_5708 ( P2_U5013 , P2_U5011 , P2_U5010 , P2_U5012 );
nand NAND2_5709 ( P2_U5014 , P2_U3045 , P2_U5009 );
nand NAND2_5710 ( P2_U5015 , P2_U3947 , P2_U5013 );
nand NAND2_5711 ( P2_U5016 , P2_R1170_U70 , P2_U3044 );
nand NAND2_5712 ( P2_U5017 , P2_REG3_REG_9_ , P2_U3088 );
nand NAND2_5713 ( P2_U5018 , P2_U3042 , P2_U3455 );
nand NAND2_5714 ( P2_U5019 , P2_R1209_U70 , P2_U3040 );
nand NAND2_5715 ( P2_U5020 , P2_ADDR_REG_9_ , P2_U4863 );
nand NAND2_5716 ( P2_U5021 , P2_R1170_U71 , P2_U3043 );
nand NAND2_5717 ( P2_U5022 , P2_U3041 , P2_U3452 );
nand NAND2_5718 ( P2_U5023 , P2_R1209_U71 , P2_U3039 );
nand NAND3_5719 ( P2_U5024 , P2_U5022 , P2_U5021 , P2_U5023 );
nand NAND2_5720 ( P2_U5025 , P2_R1170_U71 , P2_U3018 );
nand NAND2_5721 ( P2_U5026 , P2_R1209_U71 , P2_U3017 );
nand NAND2_5722 ( P2_U5027 , P2_U5683 , P2_U3452 );
nand NAND3_5723 ( P2_U5028 , P2_U5026 , P2_U5025 , P2_U5027 );
nand NAND2_5724 ( P2_U5029 , P2_U3045 , P2_U5024 );
nand NAND2_5725 ( P2_U5030 , P2_U3947 , P2_U5028 );
nand NAND2_5726 ( P2_U5031 , P2_R1170_U71 , P2_U3044 );
nand NAND2_5727 ( P2_U5032 , P2_REG3_REG_8_ , P2_U3088 );
nand NAND2_5728 ( P2_U5033 , P2_U3042 , P2_U3452 );
nand NAND2_5729 ( P2_U5034 , P2_R1209_U71 , P2_U3040 );
nand NAND2_5730 ( P2_U5035 , P2_ADDR_REG_8_ , P2_U4863 );
nand NAND2_5731 ( P2_U5036 , P2_R1170_U16 , P2_U3043 );
nand NAND2_5732 ( P2_U5037 , P2_U3041 , P2_U3449 );
nand NAND2_5733 ( P2_U5038 , P2_R1209_U16 , P2_U3039 );
nand NAND3_5734 ( P2_U5039 , P2_U5037 , P2_U5036 , P2_U5038 );
nand NAND2_5735 ( P2_U5040 , P2_R1170_U16 , P2_U3018 );
nand NAND2_5736 ( P2_U5041 , P2_R1209_U16 , P2_U3017 );
nand NAND2_5737 ( P2_U5042 , P2_U5683 , P2_U3449 );
nand NAND3_5738 ( P2_U5043 , P2_U5041 , P2_U5040 , P2_U5042 );
nand NAND2_5739 ( P2_U5044 , P2_U3045 , P2_U5039 );
nand NAND2_5740 ( P2_U5045 , P2_U3947 , P2_U5043 );
nand NAND2_5741 ( P2_U5046 , P2_R1170_U16 , P2_U3044 );
nand NAND2_5742 ( P2_U5047 , P2_REG3_REG_7_ , P2_U3088 );
nand NAND2_5743 ( P2_U5048 , P2_U3042 , P2_U3449 );
nand NAND2_5744 ( P2_U5049 , P2_R1209_U16 , P2_U3040 );
nand NAND2_5745 ( P2_U5050 , P2_ADDR_REG_7_ , P2_U4863 );
nand NAND2_5746 ( P2_U5051 , P2_R1170_U72 , P2_U3043 );
nand NAND2_5747 ( P2_U5052 , P2_U3041 , P2_U3446 );
nand NAND2_5748 ( P2_U5053 , P2_R1209_U72 , P2_U3039 );
nand NAND3_5749 ( P2_U5054 , P2_U5052 , P2_U5051 , P2_U5053 );
nand NAND2_5750 ( P2_U5055 , P2_R1170_U72 , P2_U3018 );
nand NAND2_5751 ( P2_U5056 , P2_R1209_U72 , P2_U3017 );
nand NAND2_5752 ( P2_U5057 , P2_U5683 , P2_U3446 );
nand NAND3_5753 ( P2_U5058 , P2_U5056 , P2_U5055 , P2_U5057 );
nand NAND2_5754 ( P2_U5059 , P2_U3045 , P2_U5054 );
nand NAND2_5755 ( P2_U5060 , P2_U3947 , P2_U5058 );
nand NAND2_5756 ( P2_U5061 , P2_R1170_U72 , P2_U3044 );
nand NAND2_5757 ( P2_U5062 , P2_REG3_REG_6_ , P2_U3088 );
nand NAND2_5758 ( P2_U5063 , P2_U3042 , P2_U3446 );
nand NAND2_5759 ( P2_U5064 , P2_R1209_U72 , P2_U3040 );
nand NAND2_5760 ( P2_U5065 , P2_ADDR_REG_6_ , P2_U4863 );
nand NAND2_5761 ( P2_U5066 , P2_R1170_U15 , P2_U3043 );
nand NAND2_5762 ( P2_U5067 , P2_U3041 , P2_U3443 );
nand NAND2_5763 ( P2_U5068 , P2_R1209_U15 , P2_U3039 );
nand NAND3_5764 ( P2_U5069 , P2_U5067 , P2_U5066 , P2_U5068 );
nand NAND2_5765 ( P2_U5070 , P2_R1170_U15 , P2_U3018 );
nand NAND2_5766 ( P2_U5071 , P2_R1209_U15 , P2_U3017 );
nand NAND2_5767 ( P2_U5072 , P2_U5683 , P2_U3443 );
nand NAND3_5768 ( P2_U5073 , P2_U5071 , P2_U5070 , P2_U5072 );
nand NAND2_5769 ( P2_U5074 , P2_U3045 , P2_U5069 );
nand NAND2_5770 ( P2_U5075 , P2_U3947 , P2_U5073 );
nand NAND2_5771 ( P2_U5076 , P2_R1170_U15 , P2_U3044 );
nand NAND2_5772 ( P2_U5077 , P2_REG3_REG_5_ , P2_U3088 );
nand NAND2_5773 ( P2_U5078 , P2_U3042 , P2_U3443 );
nand NAND2_5774 ( P2_U5079 , P2_R1209_U15 , P2_U3040 );
nand NAND2_5775 ( P2_U5080 , P2_ADDR_REG_5_ , P2_U4863 );
nand NAND2_5776 ( P2_U5081 , P2_R1170_U73 , P2_U3043 );
nand NAND2_5777 ( P2_U5082 , P2_U3041 , P2_U3440 );
nand NAND2_5778 ( P2_U5083 , P2_R1209_U73 , P2_U3039 );
nand NAND3_5779 ( P2_U5084 , P2_U5082 , P2_U5081 , P2_U5083 );
nand NAND2_5780 ( P2_U5085 , P2_R1170_U73 , P2_U3018 );
nand NAND2_5781 ( P2_U5086 , P2_R1209_U73 , P2_U3017 );
nand NAND2_5782 ( P2_U5087 , P2_U5683 , P2_U3440 );
nand NAND3_5783 ( P2_U5088 , P2_U5086 , P2_U5085 , P2_U5087 );
nand NAND2_5784 ( P2_U5089 , P2_U3045 , P2_U5084 );
nand NAND2_5785 ( P2_U5090 , P2_U3947 , P2_U5088 );
nand NAND2_5786 ( P2_U5091 , P2_R1170_U73 , P2_U3044 );
nand NAND2_5787 ( P2_U5092 , P2_REG3_REG_4_ , P2_U3088 );
nand NAND2_5788 ( P2_U5093 , P2_U3042 , P2_U3440 );
nand NAND2_5789 ( P2_U5094 , P2_R1209_U73 , P2_U3040 );
nand NAND2_5790 ( P2_U5095 , P2_ADDR_REG_4_ , P2_U4863 );
nand NAND2_5791 ( P2_U5096 , P2_R1170_U74 , P2_U3043 );
nand NAND2_5792 ( P2_U5097 , P2_U3041 , P2_U3437 );
nand NAND2_5793 ( P2_U5098 , P2_R1209_U74 , P2_U3039 );
nand NAND3_5794 ( P2_U5099 , P2_U5097 , P2_U5096 , P2_U5098 );
nand NAND2_5795 ( P2_U5100 , P2_R1170_U74 , P2_U3018 );
nand NAND2_5796 ( P2_U5101 , P2_R1209_U74 , P2_U3017 );
nand NAND2_5797 ( P2_U5102 , P2_U5683 , P2_U3437 );
nand NAND3_5798 ( P2_U5103 , P2_U5101 , P2_U5100 , P2_U5102 );
nand NAND2_5799 ( P2_U5104 , P2_U3045 , P2_U5099 );
nand NAND2_5800 ( P2_U5105 , P2_U3947 , P2_U5103 );
nand NAND2_5801 ( P2_U5106 , P2_R1170_U74 , P2_U3044 );
nand NAND2_5802 ( P2_U5107 , P2_REG3_REG_3_ , P2_U3088 );
nand NAND2_5803 ( P2_U5108 , P2_U3042 , P2_U3437 );
nand NAND2_5804 ( P2_U5109 , P2_R1209_U74 , P2_U3040 );
nand NAND2_5805 ( P2_U5110 , P2_ADDR_REG_3_ , P2_U4863 );
nand NAND2_5806 ( P2_U5111 , P2_R1170_U14 , P2_U3043 );
nand NAND2_5807 ( P2_U5112 , P2_U3041 , P2_U3434 );
nand NAND2_5808 ( P2_U5113 , P2_R1209_U14 , P2_U3039 );
nand NAND3_5809 ( P2_U5114 , P2_U5112 , P2_U5111 , P2_U5113 );
nand NAND2_5810 ( P2_U5115 , P2_R1170_U14 , P2_U3018 );
nand NAND2_5811 ( P2_U5116 , P2_R1209_U14 , P2_U3017 );
nand NAND2_5812 ( P2_U5117 , P2_U5683 , P2_U3434 );
nand NAND3_5813 ( P2_U5118 , P2_U5116 , P2_U5115 , P2_U5117 );
nand NAND2_5814 ( P2_U5119 , P2_U3045 , P2_U5114 );
nand NAND2_5815 ( P2_U5120 , P2_U3947 , P2_U5118 );
nand NAND2_5816 ( P2_U5121 , P2_R1170_U14 , P2_U3044 );
nand NAND2_5817 ( P2_U5122 , P2_REG3_REG_2_ , P2_U3088 );
nand NAND2_5818 ( P2_U5123 , P2_U3042 , P2_U3434 );
nand NAND2_5819 ( P2_U5124 , P2_R1209_U14 , P2_U3040 );
nand NAND2_5820 ( P2_U5125 , P2_ADDR_REG_2_ , P2_U4863 );
nand NAND2_5821 ( P2_U5126 , P2_R1170_U68 , P2_U3043 );
nand NAND2_5822 ( P2_U5127 , P2_U3041 , P2_U3431 );
nand NAND2_5823 ( P2_U5128 , P2_R1209_U68 , P2_U3039 );
nand NAND3_5824 ( P2_U5129 , P2_U5127 , P2_U5126 , P2_U5128 );
nand NAND2_5825 ( P2_U5130 , P2_R1170_U68 , P2_U3018 );
nand NAND2_5826 ( P2_U5131 , P2_R1209_U68 , P2_U3017 );
nand NAND2_5827 ( P2_U5132 , P2_U5683 , P2_U3431 );
nand NAND3_5828 ( P2_U5133 , P2_U5131 , P2_U5130 , P2_U5132 );
nand NAND2_5829 ( P2_U5134 , P2_U3045 , P2_U5129 );
nand NAND2_5830 ( P2_U5135 , P2_U3947 , P2_U5133 );
nand NAND2_5831 ( P2_U5136 , P2_R1170_U68 , P2_U3044 );
nand NAND2_5832 ( P2_U5137 , P2_REG3_REG_1_ , P2_U3088 );
nand NAND2_5833 ( P2_U5138 , P2_U3042 , P2_U3431 );
nand NAND2_5834 ( P2_U5139 , P2_R1209_U68 , P2_U3040 );
nand NAND2_5835 ( P2_U5140 , P2_ADDR_REG_1_ , P2_U4863 );
nand NAND2_5836 ( P2_U5141 , P2_R1170_U69 , P2_U3043 );
nand NAND2_5837 ( P2_U5142 , P2_U3041 , P2_U3425 );
nand NAND2_5838 ( P2_U5143 , P2_R1209_U69 , P2_U3039 );
nand NAND3_5839 ( P2_U5144 , P2_U5142 , P2_U5141 , P2_U5143 );
nand NAND2_5840 ( P2_U5145 , P2_R1170_U69 , P2_U3018 );
nand NAND2_5841 ( P2_U5146 , P2_R1209_U69 , P2_U3017 );
nand NAND2_5842 ( P2_U5147 , P2_U5683 , P2_U3425 );
nand NAND3_5843 ( P2_U5148 , P2_U5146 , P2_U5145 , P2_U5147 );
nand NAND2_5844 ( P2_U5149 , P2_U3045 , P2_U5144 );
nand NAND2_5845 ( P2_U5150 , P2_U3947 , P2_U5148 );
nand NAND2_5846 ( P2_U5151 , P2_R1170_U69 , P2_U3044 );
nand NAND2_5847 ( P2_U5152 , P2_REG3_REG_0_ , P2_U3088 );
nand NAND2_5848 ( P2_U5153 , P2_U3042 , P2_U3425 );
nand NAND2_5849 ( P2_U5154 , P2_R1209_U69 , P2_U3040 );
nand NAND2_5850 ( P2_U5155 , P2_ADDR_REG_0_ , P2_U4863 );
not NOT1_5851 ( P2_U5156 , P2_U3918 );
nand NAND3_5852 ( P2_U5157 , P2_U3936 , P2_U3334 , P2_U3337 );
nand NAND2_5853 ( P2_U5158 , P2_U5665 , P2_U5671 );
nand NAND2_5854 ( P2_U5159 , P2_U3424 , P2_U5158 );
nand NAND2_5855 ( P2_U5160 , P2_U3419 , P2_U5159 );
nand NAND2_5856 ( P2_U5161 , P2_U3340 , P2_U5160 );
nand NAND3_5857 ( P2_U5162 , P2_U6052 , P2_U6051 , P2_U3052 );
nand NAND2_5858 ( P2_U5163 , P2_B_REG , P2_U5162 );
nand NAND2_5859 ( P2_U5164 , P2_U3038 , P2_U3081 );
nand NAND2_5860 ( P2_U5165 , P2_U3036 , P2_U3075 );
nand NAND2_5861 ( P2_U5166 , P2_ADD_1119_U69 , P2_U3406 );
nand NAND3_5862 ( P2_U5167 , P2_U5165 , P2_U5164 , P2_U5166 );
not NOT1_5863 ( P2_U5168 , P2_U3154 );
nand NAND2_5864 ( P2_U5169 , P2_U3923 , P2_U3346 );
nand NAND2_5865 ( P2_U5170 , P2_U3419 , P2_U5169 );
nand NAND3_5866 ( P2_U5171 , P2_U3800 , P2_U5170 , P2_U3801 );
nand NAND2_5867 ( P2_U5172 , P2_U5171 , P2_U3406 );
not NOT1_5868 ( P2_U5173 , P2_U3408 );
nand NAND2_5869 ( P2_U5174 , P2_U3474 , P2_U5636 );
nand NAND2_5870 ( P2_U5175 , P2_ADD_1119_U69 , P2_U5635 );
nand NAND2_5871 ( P2_U5176 , P2_R1176_U111 , P2_U3028 );
nand NAND2_5872 ( P2_U5177 , P2_U3969 , P2_U5167 );
nand NAND2_5873 ( P2_U5178 , P2_REG3_REG_15_ , P2_U3088 );
nand NAND2_5874 ( P2_U5179 , P2_U3038 , P2_U3060 );
nand NAND2_5875 ( P2_U5180 , P2_U3036 , P2_U3055 );
nand NAND2_5876 ( P2_U5181 , P2_ADD_1119_U58 , P2_U3406 );
nand NAND3_5877 ( P2_U5182 , P2_U5181 , P2_U5179 , P2_U5180 );
nand NAND2_5878 ( P2_U5183 , P2_U3398 , P2_U3406 );
nand NAND2_5879 ( P2_U5184 , P2_U5173 , P2_U5183 );
nand NAND2_5880 ( P2_U5185 , P2_U3946 , P2_U3398 );
nand NAND2_5881 ( P2_U5186 , P2_U3393 , P2_U5185 );
nand NAND2_5882 ( P2_U5187 , P2_U3047 , P2_U3951 );
nand NAND2_5883 ( P2_U5188 , P2_U3046 , P2_ADD_1119_U58 );
nand NAND2_5884 ( P2_U5189 , P2_R1176_U16 , P2_U3028 );
nand NAND2_5885 ( P2_U5190 , P2_U3969 , P2_U5182 );
nand NAND2_5886 ( P2_U5191 , P2_REG3_REG_26_ , P2_U3088 );
nand NAND2_5887 ( P2_U5192 , P2_U3038 , P2_U3069 );
nand NAND2_5888 ( P2_U5193 , P2_U3036 , P2_U3072 );
nand NAND2_5889 ( P2_U5194 , P2_ADD_1119_U53 , P2_U3406 );
nand NAND3_5890 ( P2_U5195 , P2_U5193 , P2_U5192 , P2_U5194 );
nand NAND2_5891 ( P2_U5196 , P2_U3447 , P2_U5636 );
nand NAND2_5892 ( P2_U5197 , P2_ADD_1119_U53 , P2_U5635 );
nand NAND2_5893 ( P2_U5198 , P2_R1176_U96 , P2_U3028 );
nand NAND2_5894 ( P2_U5199 , P2_U3969 , P2_U5195 );
nand NAND2_5895 ( P2_U5200 , P2_REG3_REG_6_ , P2_U3088 );
nand NAND2_5896 ( P2_U5201 , P2_U3038 , P2_U3071 );
nand NAND2_5897 ( P2_U5202 , P2_U3036 , P2_U3083 );
nand NAND2_5898 ( P2_U5203 , P2_ADD_1119_U66 , P2_U3406 );
nand NAND3_5899 ( P2_U5204 , P2_U5202 , P2_U5201 , P2_U5203 );
nand NAND2_5900 ( P2_U5205 , P2_U3483 , P2_U5636 );
nand NAND2_5901 ( P2_U5206 , P2_ADD_1119_U66 , P2_U5635 );
nand NAND2_5902 ( P2_U5207 , P2_R1176_U109 , P2_U3028 );
nand NAND2_5903 ( P2_U5208 , P2_U3969 , P2_U5204 );
nand NAND2_5904 ( P2_U5209 , P2_REG3_REG_18_ , P2_U3088 );
nand NAND2_5905 ( P2_U5210 , P2_U3038 , P2_U3080 );
nand NAND2_5906 ( P2_U5211 , P2_U3036 , P2_U3066 );
nand NAND2_5907 ( P2_U5212 , P2_REG3_REG_2_ , P2_U3406 );
nand NAND3_5908 ( P2_U5213 , P2_U5211 , P2_U5210 , P2_U5212 );
nand NAND2_5909 ( P2_U5214 , P2_U3435 , P2_U5636 );
nand NAND2_5910 ( P2_U5215 , P2_REG3_REG_2_ , P2_U5635 );
nand NAND2_5911 ( P2_U5216 , P2_R1176_U99 , P2_U3028 );
nand NAND2_5912 ( P2_U5217 , P2_U3969 , P2_U5213 );
nand NAND2_5913 ( P2_U5218 , P2_REG3_REG_2_ , P2_U3088 );
nand NAND2_5914 ( P2_U5219 , P2_U3038 , P2_U3064 );
nand NAND2_5915 ( P2_U5220 , P2_U3036 , P2_U3074 );
nand NAND2_5916 ( P2_U5221 , P2_ADD_1119_U73 , P2_U3406 );
nand NAND3_5917 ( P2_U5222 , P2_U5220 , P2_U5219 , P2_U5221 );
nand NAND2_5918 ( P2_U5223 , P2_U3462 , P2_U5636 );
nand NAND2_5919 ( P2_U5224 , P2_ADD_1119_U73 , P2_U5635 );
nand NAND2_5920 ( P2_U5225 , P2_R1176_U114 , P2_U3028 );
nand NAND2_5921 ( P2_U5226 , P2_U3969 , P2_U5222 );
nand NAND2_5922 ( P2_U5227 , P2_REG3_REG_11_ , P2_U3088 );
nand NAND2_5923 ( P2_U5228 , P2_U3038 , P2_U3077 );
nand NAND2_5924 ( P2_U5229 , P2_U3036 , P2_U3068 );
nand NAND2_5925 ( P2_U5230 , P2_ADD_1119_U62 , P2_U3406 );
nand NAND3_5926 ( P2_U5231 , P2_U5229 , P2_U5228 , P2_U5230 );
nand NAND2_5927 ( P2_U5232 , P2_U3047 , P2_U3955 );
nand NAND2_5928 ( P2_U5233 , P2_U3046 , P2_ADD_1119_U62 );
nand NAND2_5929 ( P2_U5234 , P2_R1176_U105 , P2_U3028 );
nand NAND2_5930 ( P2_U5235 , P2_U3969 , P2_U5231 );
nand NAND2_5931 ( P2_U5236 , P2_REG3_REG_22_ , P2_U3088 );
nand NAND2_5932 ( P2_U5237 , P2_U3038 , P2_U3074 );
nand NAND2_5933 ( P2_U5238 , P2_U3036 , P2_U3081 );
nand NAND2_5934 ( P2_U5239 , P2_ADD_1119_U71 , P2_U3406 );
nand NAND3_5935 ( P2_U5240 , P2_U5238 , P2_U5237 , P2_U5239 );
nand NAND2_5936 ( P2_U5241 , P2_U3468 , P2_U5636 );
nand NAND2_5937 ( P2_U5242 , P2_ADD_1119_U71 , P2_U5635 );
nand NAND2_5938 ( P2_U5243 , P2_R1176_U13 , P2_U3028 );
nand NAND2_5939 ( P2_U5244 , P2_U3969 , P2_U5240 );
nand NAND2_5940 ( P2_U5245 , P2_REG3_REG_13_ , P2_U3088 );
nand NAND2_5941 ( P2_U5246 , P2_U3038 , P2_U3083 );
nand NAND2_5942 ( P2_U5247 , P2_U3036 , P2_U3077 );
nand NAND2_5943 ( P2_U5248 , P2_ADD_1119_U64 , P2_U3406 );
nand NAND3_5944 ( P2_U5249 , P2_U5247 , P2_U5246 , P2_U5248 );
nand NAND2_5945 ( P2_U5250 , P2_U3047 , P2_U3957 );
nand NAND2_5946 ( P2_U5251 , P2_U3046 , P2_ADD_1119_U64 );
nand NAND2_5947 ( P2_U5252 , P2_R1176_U106 , P2_U3028 );
nand NAND2_5948 ( P2_U5253 , P2_U3969 , P2_U5249 );
nand NAND2_5949 ( P2_U5254 , P2_REG3_REG_20_ , P2_U3088 );
nand NAND2_5950 ( P2_U5255 , P2_U3407 , P2_U3405 );
nand NAND2_5951 ( P2_U5256 , P2_U5255 , P2_U3406 );
nand NAND2_5952 ( P2_U5257 , P2_U3970 , P2_U5256 );
nand NAND2_5953 ( P2_U5258 , P2_U3806 , P2_U3036 );
nand NAND2_5954 ( P2_U5259 , P2_U3427 , P2_U5636 );
nand NAND2_5955 ( P2_U5260 , P2_REG3_REG_0_ , P2_U5257 );
nand NAND2_5956 ( P2_U5261 , P2_R1176_U93 , P2_U3028 );
nand NAND2_5957 ( P2_U5262 , P2_REG3_REG_0_ , P2_U3088 );
nand NAND2_5958 ( P2_U5263 , P2_U3038 , P2_U3086 );
nand NAND2_5959 ( P2_U5264 , P2_U3036 , P2_U3064 );
nand NAND2_5960 ( P2_U5265 , P2_ADD_1119_U50 , P2_U3406 );
nand NAND3_5961 ( P2_U5266 , P2_U5264 , P2_U5263 , P2_U5265 );
nand NAND2_5962 ( P2_U5267 , P2_U3456 , P2_U5636 );
nand NAND2_5963 ( P2_U5268 , P2_ADD_1119_U50 , P2_U5635 );
nand NAND2_5964 ( P2_U5269 , P2_R1176_U94 , P2_U3028 );
nand NAND2_5965 ( P2_U5270 , P2_U3969 , P2_U5266 );
nand NAND2_5966 ( P2_U5271 , P2_REG3_REG_9_ , P2_U3088 );
nand NAND2_5967 ( P2_U5272 , P2_U3038 , P2_U3066 );
nand NAND2_5968 ( P2_U5273 , P2_U3036 , P2_U3069 );
nand NAND2_5969 ( P2_U5274 , P2_ADD_1119_U55 , P2_U3406 );
nand NAND3_5970 ( P2_U5275 , P2_U5273 , P2_U5272 , P2_U5274 );
nand NAND2_5971 ( P2_U5276 , P2_U3441 , P2_U5636 );
nand NAND2_5972 ( P2_U5277 , P2_ADD_1119_U55 , P2_U5635 );
nand NAND2_5973 ( P2_U5278 , P2_R1176_U98 , P2_U3028 );
nand NAND2_5974 ( P2_U5279 , P2_U3969 , P2_U5275 );
nand NAND2_5975 ( P2_U5280 , P2_REG3_REG_4_ , P2_U3088 );
nand NAND2_5976 ( P2_U5281 , P2_U3038 , P2_U3068 );
nand NAND2_5977 ( P2_U5282 , P2_U3036 , P2_U3060 );
nand NAND2_5978 ( P2_U5283 , P2_ADD_1119_U60 , P2_U3406 );
nand NAND3_5979 ( P2_U5284 , P2_U5282 , P2_U5281 , P2_U5283 );
nand NAND2_5980 ( P2_U5285 , P2_U3047 , P2_U3953 );
nand NAND2_5981 ( P2_U5286 , P2_U3046 , P2_ADD_1119_U60 );
nand NAND2_5982 ( P2_U5287 , P2_R1176_U103 , P2_U3028 );
nand NAND2_5983 ( P2_U5288 , P2_U3969 , P2_U5284 );
nand NAND2_5984 ( P2_U5289 , P2_REG3_REG_24_ , P2_U3088 );
nand NAND2_5985 ( P2_U5290 , P2_U3038 , P2_U3075 );
nand NAND2_5986 ( P2_U5291 , P2_U3036 , P2_U3084 );
nand NAND2_5987 ( P2_U5292 , P2_ADD_1119_U67 , P2_U3406 );
nand NAND3_5988 ( P2_U5293 , P2_U5291 , P2_U5290 , P2_U5292 );
nand NAND2_5989 ( P2_U5294 , P2_U3480 , P2_U5636 );
nand NAND2_5990 ( P2_U5295 , P2_ADD_1119_U67 , P2_U5635 );
nand NAND2_5991 ( P2_U5296 , P2_R1176_U14 , P2_U3028 );
nand NAND2_5992 ( P2_U5297 , P2_U3969 , P2_U5293 );
nand NAND2_5993 ( P2_U5298 , P2_REG3_REG_17_ , P2_U3088 );
nand NAND2_5994 ( P2_U5299 , P2_U3038 , P2_U3062 );
nand NAND2_5995 ( P2_U5300 , P2_U3036 , P2_U3073 );
nand NAND2_5996 ( P2_U5301 , P2_ADD_1119_U54 , P2_U3406 );
nand NAND3_5997 ( P2_U5302 , P2_U5300 , P2_U5299 , P2_U5301 );
nand NAND2_5998 ( P2_U5303 , P2_U3444 , P2_U5636 );
nand NAND2_5999 ( P2_U5304 , P2_ADD_1119_U54 , P2_U5635 );
nand NAND2_6000 ( P2_U5305 , P2_R1176_U97 , P2_U3028 );
nand NAND2_6001 ( P2_U5306 , P2_U3969 , P2_U5302 );
nand NAND2_6002 ( P2_U5307 , P2_REG3_REG_5_ , P2_U3088 );
nand NAND2_6003 ( P2_U5308 , P2_U3038 , P2_U3076 );
nand NAND2_6004 ( P2_U5309 , P2_U3036 , P2_U3071 );
nand NAND2_6005 ( P2_U5310 , P2_ADD_1119_U68 , P2_U3406 );
nand NAND3_6006 ( P2_U5311 , P2_U5309 , P2_U5308 , P2_U5310 );
nand NAND2_6007 ( P2_U5312 , P2_U3477 , P2_U5636 );
nand NAND2_6008 ( P2_U5313 , P2_ADD_1119_U68 , P2_U5635 );
nand NAND2_6009 ( P2_U5314 , P2_R1176_U110 , P2_U3028 );
nand NAND2_6010 ( P2_U5315 , P2_U3969 , P2_U5311 );
nand NAND2_6011 ( P2_U5316 , P2_REG3_REG_16_ , P2_U3088 );
nand NAND2_6012 ( P2_U5317 , P2_U3038 , P2_U3067 );
nand NAND2_6013 ( P2_U5318 , P2_U3036 , P2_U3059 );
nand NAND2_6014 ( P2_U5319 , P2_ADD_1119_U59 , P2_U3406 );
nand NAND3_6015 ( P2_U5320 , P2_U5318 , P2_U5317 , P2_U5319 );
nand NAND2_6016 ( P2_U5321 , P2_U3047 , P2_U3952 );
nand NAND2_6017 ( P2_U5322 , P2_U3046 , P2_ADD_1119_U59 );
nand NAND2_6018 ( P2_U5323 , P2_R1176_U102 , P2_U3028 );
nand NAND2_6019 ( P2_U5324 , P2_U3969 , P2_U5320 );
nand NAND2_6020 ( P2_U5325 , P2_REG3_REG_25_ , P2_U3088 );
nand NAND2_6021 ( P2_U5326 , P2_U3038 , P2_U3065 );
nand NAND2_6022 ( P2_U5327 , P2_U3036 , P2_U3082 );
nand NAND2_6023 ( P2_U5328 , P2_ADD_1119_U72 , P2_U3406 );
nand NAND3_6024 ( P2_U5329 , P2_U5327 , P2_U5326 , P2_U5328 );
nand NAND2_6025 ( P2_U5330 , P2_U3465 , P2_U5636 );
nand NAND2_6026 ( P2_U5331 , P2_ADD_1119_U72 , P2_U5635 );
nand NAND2_6027 ( P2_U5332 , P2_R1176_U113 , P2_U3028 );
nand NAND2_6028 ( P2_U5333 , P2_U3969 , P2_U5329 );
nand NAND2_6029 ( P2_U5334 , P2_REG3_REG_12_ , P2_U3088 );
nand NAND2_6030 ( P2_U5335 , P2_U3038 , P2_U3078 );
nand NAND2_6031 ( P2_U5336 , P2_U3036 , P2_U3063 );
nand NAND2_6032 ( P2_U5337 , P2_ADD_1119_U63 , P2_U3406 );
nand NAND3_6033 ( P2_U5338 , P2_U5336 , P2_U5335 , P2_U5337 );
nand NAND2_6034 ( P2_U5339 , P2_U3047 , P2_U3956 );
nand NAND2_6035 ( P2_U5340 , P2_U3046 , P2_ADD_1119_U63 );
nand NAND2_6036 ( P2_U5341 , P2_R1176_U15 , P2_U3028 );
nand NAND2_6037 ( P2_U5342 , P2_U3969 , P2_U5338 );
nand NAND2_6038 ( P2_U5343 , P2_REG3_REG_21_ , P2_U3088 );
nand NAND2_6039 ( P2_U5344 , P2_U3038 , P2_U3079 );
nand NAND2_6040 ( P2_U5345 , P2_U3036 , P2_U3070 );
nand NAND2_6041 ( P2_U5346 , P2_REG3_REG_1_ , P2_U3406 );
nand NAND3_6042 ( P2_U5347 , P2_U5345 , P2_U5344 , P2_U5346 );
nand NAND2_6043 ( P2_U5348 , P2_U3432 , P2_U5636 );
nand NAND2_6044 ( P2_U5349 , P2_REG3_REG_1_ , P2_U5635 );
nand NAND2_6045 ( P2_U5350 , P2_R1176_U107 , P2_U3028 );
nand NAND2_6046 ( P2_U5351 , P2_U3969 , P2_U5347 );
nand NAND2_6047 ( P2_U5352 , P2_REG3_REG_1_ , P2_U3088 );
nand NAND2_6048 ( P2_U5353 , P2_U3038 , P2_U3072 );
nand NAND2_6049 ( P2_U5354 , P2_U3036 , P2_U3085 );
nand NAND2_6050 ( P2_U5355 , P2_ADD_1119_U51 , P2_U3406 );
nand NAND3_6051 ( P2_U5356 , P2_U5354 , P2_U5353 , P2_U5355 );
nand NAND2_6052 ( P2_U5357 , P2_U3453 , P2_U5636 );
nand NAND2_6053 ( P2_U5358 , P2_ADD_1119_U51 , P2_U5635 );
nand NAND2_6054 ( P2_U5359 , P2_R1176_U95 , P2_U3028 );
nand NAND2_6055 ( P2_U5360 , P2_U3969 , P2_U5356 );
nand NAND2_6056 ( P2_U5361 , P2_REG3_REG_8_ , P2_U3088 );
nand NAND2_6057 ( P2_U5362 , P2_U3038 , P2_U3055 );
nand NAND2_6058 ( P2_U5363 , P2_U3036 , P2_U3057 );
nand NAND2_6059 ( P2_U5364 , P2_ADD_1119_U56 , P2_U3406 );
nand NAND3_6060 ( P2_U5365 , P2_U5363 , P2_U5364 , P2_U5362 );
nand NAND2_6061 ( P2_U5366 , P2_U3047 , P2_U3949 );
nand NAND2_6062 ( P2_U5367 , P2_U3046 , P2_ADD_1119_U56 );
nand NAND2_6063 ( P2_U5368 , P2_R1176_U100 , P2_U3028 );
nand NAND2_6064 ( P2_U5369 , P2_U3969 , P2_U5365 );
nand NAND2_6065 ( P2_U5370 , P2_REG3_REG_28_ , P2_U3088 );
nand NAND2_6066 ( P2_U5371 , P2_U3038 , P2_U3084 );
nand NAND2_6067 ( P2_U5372 , P2_U3036 , P2_U3078 );
nand NAND2_6068 ( P2_U5373 , P2_ADD_1119_U65 , P2_U3406 );
nand NAND3_6069 ( P2_U5374 , P2_U5372 , P2_U5371 , P2_U5373 );
nand NAND2_6070 ( P2_U5375 , P2_U3485 , P2_U5636 );
nand NAND2_6071 ( P2_U5376 , P2_ADD_1119_U65 , P2_U5635 );
nand NAND2_6072 ( P2_U5377 , P2_R1176_U108 , P2_U3028 );
nand NAND2_6073 ( P2_U5378 , P2_U3969 , P2_U5374 );
nand NAND2_6074 ( P2_U5379 , P2_REG3_REG_19_ , P2_U3088 );
nand NAND2_6075 ( P2_U5380 , P2_U3038 , P2_U3070 );
nand NAND2_6076 ( P2_U5381 , P2_U3036 , P2_U3062 );
nand NAND2_6077 ( P2_U5382 , P2_ADD_1119_U4 , P2_U3406 );
nand NAND3_6078 ( P2_U5383 , P2_U5381 , P2_U5380 , P2_U5382 );
nand NAND2_6079 ( P2_U5384 , P2_U3438 , P2_U5636 );
nand NAND2_6080 ( P2_U5385 , P2_ADD_1119_U4 , P2_U5635 );
nand NAND2_6081 ( P2_U5386 , P2_R1176_U17 , P2_U3028 );
nand NAND2_6082 ( P2_U5387 , P2_U3969 , P2_U5383 );
nand NAND2_6083 ( P2_U5388 , P2_REG3_REG_3_ , P2_U3088 );
nand NAND2_6084 ( P2_U5389 , P2_U3038 , P2_U3085 );
nand NAND2_6085 ( P2_U5390 , P2_U3036 , P2_U3065 );
nand NAND2_6086 ( P2_U5391 , P2_ADD_1119_U74 , P2_U3406 );
nand NAND3_6087 ( P2_U5392 , P2_U5390 , P2_U5389 , P2_U5391 );
nand NAND2_6088 ( P2_U5393 , P2_U3459 , P2_U5636 );
nand NAND2_6089 ( P2_U5394 , P2_ADD_1119_U74 , P2_U5635 );
nand NAND2_6090 ( P2_U5395 , P2_R1176_U115 , P2_U3028 );
nand NAND2_6091 ( P2_U5396 , P2_U3969 , P2_U5392 );
nand NAND2_6092 ( P2_U5397 , P2_REG3_REG_10_ , P2_U3088 );
nand NAND2_6093 ( P2_U5398 , P2_U3038 , P2_U3063 );
nand NAND2_6094 ( P2_U5399 , P2_U3036 , P2_U3067 );
nand NAND2_6095 ( P2_U5400 , P2_ADD_1119_U61 , P2_U3406 );
nand NAND3_6096 ( P2_U5401 , P2_U5399 , P2_U5398 , P2_U5400 );
nand NAND2_6097 ( P2_U5402 , P2_U3047 , P2_U3954 );
nand NAND2_6098 ( P2_U5403 , P2_U3046 , P2_ADD_1119_U61 );
nand NAND2_6099 ( P2_U5404 , P2_R1176_U104 , P2_U3028 );
nand NAND2_6100 ( P2_U5405 , P2_U3969 , P2_U5401 );
nand NAND2_6101 ( P2_U5406 , P2_REG3_REG_23_ , P2_U3088 );
nand NAND2_6102 ( P2_U5407 , P2_U3038 , P2_U3082 );
nand NAND2_6103 ( P2_U5408 , P2_U3036 , P2_U3076 );
nand NAND2_6104 ( P2_U5409 , P2_ADD_1119_U70 , P2_U3406 );
nand NAND3_6105 ( P2_U5410 , P2_U5408 , P2_U5407 , P2_U5409 );
nand NAND2_6106 ( P2_U5411 , P2_U3471 , P2_U5636 );
nand NAND2_6107 ( P2_U5412 , P2_ADD_1119_U70 , P2_U5635 );
nand NAND2_6108 ( P2_U5413 , P2_R1176_U112 , P2_U3028 );
nand NAND2_6109 ( P2_U5414 , P2_U3969 , P2_U5410 );
nand NAND2_6110 ( P2_U5415 , P2_REG3_REG_14_ , P2_U3088 );
nand NAND2_6111 ( P2_U5416 , P2_U3038 , P2_U3059 );
nand NAND2_6112 ( P2_U5417 , P2_U3036 , P2_U3056 );
nand NAND2_6113 ( P2_U5418 , P2_ADD_1119_U57 , P2_U3406 );
nand NAND3_6114 ( P2_U5419 , P2_U5418 , P2_U5416 , P2_U5417 );
nand NAND2_6115 ( P2_U5420 , P2_U3047 , P2_U3950 );
nand NAND2_6116 ( P2_U5421 , P2_U3046 , P2_ADD_1119_U57 );
nand NAND2_6117 ( P2_U5422 , P2_R1176_U101 , P2_U3028 );
nand NAND2_6118 ( P2_U5423 , P2_U3969 , P2_U5419 );
nand NAND2_6119 ( P2_U5424 , P2_REG3_REG_27_ , P2_U3088 );
nand NAND2_6120 ( P2_U5425 , P2_U3038 , P2_U3073 );
nand NAND2_6121 ( P2_U5426 , P2_U3036 , P2_U3086 );
nand NAND2_6122 ( P2_U5427 , P2_ADD_1119_U52 , P2_U3406 );
nand NAND3_6123 ( P2_U5428 , P2_U5426 , P2_U5425 , P2_U5427 );
nand NAND2_6124 ( P2_U5429 , P2_U3450 , P2_U5636 );
nand NAND2_6125 ( P2_U5430 , P2_ADD_1119_U52 , P2_U5635 );
nand NAND2_6126 ( P2_U5431 , P2_R1176_U18 , P2_U3028 );
nand NAND2_6127 ( P2_U5432 , P2_U3969 , P2_U5428 );
nand NAND2_6128 ( P2_U5433 , P2_REG3_REG_7_ , P2_U3088 );
nand NAND2_6129 ( P2_U5434 , P2_U3948 , P2_U3048 );
nand NAND2_6130 ( P2_U5435 , P2_U3415 , P2_U3347 );
nand NAND2_6131 ( P2_U5436 , P2_U3419 , P2_U3418 );
nand NAND2_6132 ( P2_U5437 , P2_U3816 , P2_U3051 );
not NOT1_6133 ( P2_U5438 , P2_U3411 );
nand NAND2_6134 ( P2_U5439 , P2_U3015 , P2_U3415 );
nand NAND2_6135 ( P2_U5440 , P2_U3411 , P2_U3409 );
nand NAND2_6136 ( P2_U5441 , P2_U3053 , P2_U5440 );
nand NAND2_6137 ( P2_U5442 , P2_U3085 , P2_U3029 );
nand NAND2_6138 ( P2_U5443 , P2_U5441 , P2_U3085 );
nand NAND2_6139 ( P2_U5444 , P2_U3929 , P2_U3456 );
nand NAND2_6140 ( P2_U5445 , P2_U3086 , P2_U3029 );
nand NAND2_6141 ( P2_U5446 , P2_U5441 , P2_U3086 );
nand NAND2_6142 ( P2_U5447 , P2_U3929 , P2_U3453 );
nand NAND2_6143 ( P2_U5448 , P2_U3072 , P2_U3029 );
nand NAND2_6144 ( P2_U5449 , P2_U5441 , P2_U3072 );
nand NAND2_6145 ( P2_U5450 , P2_U3929 , P2_U3450 );
nand NAND2_6146 ( P2_U5451 , P2_U3073 , P2_U3029 );
nand NAND2_6147 ( P2_U5452 , P2_U5441 , P2_U3073 );
nand NAND2_6148 ( P2_U5453 , P2_U3929 , P2_U3447 );
nand NAND2_6149 ( P2_U5454 , P2_U3069 , P2_U3029 );
nand NAND2_6150 ( P2_U5455 , P2_U5441 , P2_U3069 );
nand NAND2_6151 ( P2_U5456 , P2_U3929 , P2_U3444 );
nand NAND2_6152 ( P2_U5457 , P2_U3062 , P2_U3029 );
nand NAND2_6153 ( P2_U5458 , P2_U5441 , P2_U3062 );
nand NAND2_6154 ( P2_U5459 , P2_U3929 , P2_U3441 );
nand NAND2_6155 ( P2_U5460 , P2_R1335_U8 , P2_U3029 );
nand NAND2_6156 ( P2_U5461 , P2_U5441 , P2_U3058 );
nand NAND2_6157 ( P2_U5462 , P2_R1335_U6 , P2_U3029 );
nand NAND2_6158 ( P2_U5463 , P2_U5441 , P2_U3061 );
nand NAND3_6159 ( P2_U5464 , P2_U3929 , P2_U3347 , U70 );
nand NAND2_6160 ( P2_U5465 , P2_U3066 , P2_U3029 );
nand NAND2_6161 ( P2_U5466 , P2_U5441 , P2_U3066 );
nand NAND2_6162 ( P2_U5467 , P2_U3929 , P2_U3438 );
nand NAND2_6163 ( P2_U5468 , P2_U3057 , P2_U3029 );
nand NAND2_6164 ( P2_U5469 , P2_U5441 , P2_U3057 );
nand NAND2_6165 ( P2_U5470 , P2_U3929 , P2_U3960 );
nand NAND2_6166 ( P2_U5471 , P2_U3056 , P2_U3029 );
nand NAND2_6167 ( P2_U5472 , P2_U5441 , P2_U3056 );
nand NAND2_6168 ( P2_U5473 , P2_U3929 , P2_U3949 );
nand NAND2_6169 ( P2_U5474 , P2_U3055 , P2_U3029 );
nand NAND2_6170 ( P2_U5475 , P2_U5441 , P2_U3055 );
nand NAND2_6171 ( P2_U5476 , P2_U3929 , P2_U3950 );
nand NAND2_6172 ( P2_U5477 , P2_U3059 , P2_U3029 );
nand NAND2_6173 ( P2_U5478 , P2_U5441 , P2_U3059 );
nand NAND2_6174 ( P2_U5479 , P2_U3929 , P2_U3951 );
nand NAND2_6175 ( P2_U5480 , P2_U3060 , P2_U3029 );
nand NAND2_6176 ( P2_U5481 , P2_U5441 , P2_U3060 );
nand NAND2_6177 ( P2_U5482 , P2_U3929 , P2_U3952 );
nand NAND2_6178 ( P2_U5483 , P2_U3067 , P2_U3029 );
nand NAND2_6179 ( P2_U5484 , P2_U5441 , P2_U3067 );
nand NAND2_6180 ( P2_U5485 , P2_U3929 , P2_U3953 );
nand NAND2_6181 ( P2_U5486 , P2_U3068 , P2_U3029 );
nand NAND2_6182 ( P2_U5487 , P2_U5441 , P2_U3068 );
nand NAND2_6183 ( P2_U5488 , P2_U3929 , P2_U3954 );
nand NAND2_6184 ( P2_U5489 , P2_U3063 , P2_U3029 );
nand NAND2_6185 ( P2_U5490 , P2_U5441 , P2_U3063 );
nand NAND2_6186 ( P2_U5491 , P2_U3929 , P2_U3955 );
nand NAND2_6187 ( P2_U5492 , P2_U3077 , P2_U3029 );
nand NAND2_6188 ( P2_U5493 , P2_U5441 , P2_U3077 );
nand NAND2_6189 ( P2_U5494 , P2_U3929 , P2_U3956 );
nand NAND2_6190 ( P2_U5495 , P2_U3078 , P2_U3029 );
nand NAND2_6191 ( P2_U5496 , P2_U5441 , P2_U3078 );
nand NAND2_6192 ( P2_U5497 , P2_U3929 , P2_U3957 );
nand NAND2_6193 ( P2_U5498 , P2_U3070 , P2_U3029 );
nand NAND2_6194 ( P2_U5499 , P2_U5441 , P2_U3070 );
nand NAND2_6195 ( P2_U5500 , P2_U3929 , P2_U3435 );
nand NAND2_6196 ( P2_U5501 , P2_U3083 , P2_U3029 );
nand NAND2_6197 ( P2_U5502 , P2_U5441 , P2_U3083 );
nand NAND2_6198 ( P2_U5503 , P2_U3929 , P2_U3485 );
nand NAND2_6199 ( P2_U5504 , P2_U3084 , P2_U3029 );
nand NAND2_6200 ( P2_U5505 , P2_U5441 , P2_U3084 );
nand NAND2_6201 ( P2_U5506 , P2_U3929 , P2_U3483 );
nand NAND2_6202 ( P2_U5507 , P2_U3071 , P2_U3029 );
nand NAND2_6203 ( P2_U5508 , P2_U5441 , P2_U3071 );
nand NAND2_6204 ( P2_U5509 , P2_U3929 , P2_U3480 );
nand NAND2_6205 ( P2_U5510 , P2_U3075 , P2_U3029 );
nand NAND2_6206 ( P2_U5511 , P2_U5441 , P2_U3075 );
nand NAND2_6207 ( P2_U5512 , P2_U3929 , P2_U3477 );
nand NAND2_6208 ( P2_U5513 , P2_U3076 , P2_U3029 );
nand NAND2_6209 ( P2_U5514 , P2_U5441 , P2_U3076 );
nand NAND2_6210 ( P2_U5515 , P2_U3929 , P2_U3474 );
nand NAND2_6211 ( P2_U5516 , P2_U3081 , P2_U3029 );
nand NAND2_6212 ( P2_U5517 , P2_U5441 , P2_U3081 );
nand NAND2_6213 ( P2_U5518 , P2_U3929 , P2_U3471 );
nand NAND2_6214 ( P2_U5519 , P2_U3082 , P2_U3029 );
nand NAND2_6215 ( P2_U5520 , P2_U5441 , P2_U3082 );
nand NAND2_6216 ( P2_U5521 , P2_U3929 , P2_U3468 );
nand NAND2_6217 ( P2_U5522 , P2_U3074 , P2_U3029 );
nand NAND2_6218 ( P2_U5523 , P2_U5441 , P2_U3074 );
nand NAND2_6219 ( P2_U5524 , P2_U3929 , P2_U3465 );
nand NAND2_6220 ( P2_U5525 , P2_U3065 , P2_U3029 );
nand NAND2_6221 ( P2_U5526 , P2_U5441 , P2_U3065 );
nand NAND2_6222 ( P2_U5527 , P2_U3929 , P2_U3462 );
nand NAND2_6223 ( P2_U5528 , P2_U3064 , P2_U3029 );
nand NAND2_6224 ( P2_U5529 , P2_U5441 , P2_U3064 );
nand NAND2_6225 ( P2_U5530 , P2_U3929 , P2_U3459 );
nand NAND2_6226 ( P2_U5531 , P2_U3080 , P2_U3029 );
nand NAND2_6227 ( P2_U5532 , P2_U5441 , P2_U3080 );
nand NAND2_6228 ( P2_U5533 , P2_U3929 , P2_U3432 );
nand NAND2_6229 ( P2_U5534 , P2_U3079 , P2_U3029 );
nand NAND2_6230 ( P2_U5535 , P2_U5441 , P2_U3079 );
nand NAND2_6231 ( P2_U5536 , P2_U3929 , P2_U3427 );
nand NAND2_6232 ( P2_U5537 , P2_U5438 , P2_U3053 );
nand NAND2_6233 ( P2_U5538 , P2_U3456 , P2_U5537 );
nand NAND2_6234 ( P2_U5539 , P2_U3929 , P2_U3085 );
nand NAND2_6235 ( P2_U5540 , P2_U5658 , P2_U3086 );
nand NAND2_6236 ( P2_U5541 , P2_U3453 , P2_U5537 );
nand NAND2_6237 ( P2_U5542 , P2_U3929 , P2_U3086 );
nand NAND2_6238 ( P2_U5543 , P2_U5658 , P2_U3072 );
nand NAND2_6239 ( P2_U5544 , P2_U3450 , P2_U5537 );
nand NAND2_6240 ( P2_U5545 , P2_U3929 , P2_U3072 );
nand NAND2_6241 ( P2_U5546 , P2_U5658 , P2_U3073 );
nand NAND2_6242 ( P2_U5547 , P2_U3447 , P2_U5537 );
nand NAND2_6243 ( P2_U5548 , P2_U3929 , P2_U3073 );
nand NAND2_6244 ( P2_U5549 , P2_U5658 , P2_U3069 );
nand NAND2_6245 ( P2_U5550 , P2_U3444 , P2_U5537 );
nand NAND2_6246 ( P2_U5551 , P2_U3929 , P2_U3069 );
nand NAND2_6247 ( P2_U5552 , P2_U5658 , P2_U3062 );
nand NAND2_6248 ( P2_U5553 , P2_U3441 , P2_U5537 );
nand NAND2_6249 ( P2_U5554 , P2_U3929 , P2_U3062 );
nand NAND2_6250 ( P2_U5555 , P2_U5658 , P2_U3066 );
nand NAND3_6251 ( P2_U5556 , P2_U5537 , P2_U3347 , U69 );
nand NAND2_6252 ( P2_U5557 , P2_U3929 , P2_U3058 );
nand NAND2_6253 ( P2_U5558 , P2_U3959 , P2_U5537 );
nand NAND2_6254 ( P2_U5559 , P2_U3929 , P2_U3061 );
nand NAND2_6255 ( P2_U5560 , P2_U3438 , P2_U5537 );
nand NAND2_6256 ( P2_U5561 , P2_U3929 , P2_U3066 );
nand NAND2_6257 ( P2_U5562 , P2_U5658 , P2_U3070 );
nand NAND2_6258 ( P2_U5563 , P2_U3960 , P2_U5537 );
nand NAND2_6259 ( P2_U5564 , P2_U3929 , P2_U3057 );
nand NAND2_6260 ( P2_U5565 , P2_U5658 , P2_U3056 );
nand NAND2_6261 ( P2_U5566 , P2_U3949 , P2_U5537 );
nand NAND2_6262 ( P2_U5567 , P2_U3929 , P2_U3056 );
nand NAND2_6263 ( P2_U5568 , P2_U5658 , P2_U3055 );
nand NAND2_6264 ( P2_U5569 , P2_U3950 , P2_U5537 );
nand NAND2_6265 ( P2_U5570 , P2_U3929 , P2_U3055 );
nand NAND2_6266 ( P2_U5571 , P2_U5658 , P2_U3059 );
nand NAND2_6267 ( P2_U5572 , P2_U3951 , P2_U5537 );
nand NAND2_6268 ( P2_U5573 , P2_U3929 , P2_U3059 );
nand NAND2_6269 ( P2_U5574 , P2_U5658 , P2_U3060 );
nand NAND2_6270 ( P2_U5575 , P2_U3952 , P2_U5537 );
nand NAND2_6271 ( P2_U5576 , P2_U3929 , P2_U3060 );
nand NAND2_6272 ( P2_U5577 , P2_U5658 , P2_U3067 );
nand NAND2_6273 ( P2_U5578 , P2_U3953 , P2_U5537 );
nand NAND2_6274 ( P2_U5579 , P2_U3929 , P2_U3067 );
nand NAND2_6275 ( P2_U5580 , P2_U5658 , P2_U3068 );
nand NAND2_6276 ( P2_U5581 , P2_U3954 , P2_U5537 );
nand NAND2_6277 ( P2_U5582 , P2_U3929 , P2_U3068 );
nand NAND2_6278 ( P2_U5583 , P2_U5658 , P2_U3063 );
nand NAND2_6279 ( P2_U5584 , P2_U3955 , P2_U5537 );
nand NAND2_6280 ( P2_U5585 , P2_U3929 , P2_U3063 );
nand NAND2_6281 ( P2_U5586 , P2_U5658 , P2_U3077 );
nand NAND2_6282 ( P2_U5587 , P2_U3956 , P2_U5537 );
nand NAND2_6283 ( P2_U5588 , P2_U3929 , P2_U3077 );
nand NAND2_6284 ( P2_U5589 , P2_U5658 , P2_U3078 );
nand NAND2_6285 ( P2_U5590 , P2_U3957 , P2_U5537 );
nand NAND2_6286 ( P2_U5591 , P2_U3929 , P2_U3078 );
nand NAND2_6287 ( P2_U5592 , P2_U5658 , P2_U3083 );
nand NAND2_6288 ( P2_U5593 , P2_U3435 , P2_U5537 );
nand NAND2_6289 ( P2_U5594 , P2_U3929 , P2_U3070 );
nand NAND2_6290 ( P2_U5595 , P2_U5658 , P2_U3080 );
nand NAND2_6291 ( P2_U5596 , P2_U3485 , P2_U5537 );
nand NAND2_6292 ( P2_U5597 , P2_U3929 , P2_U3083 );
nand NAND2_6293 ( P2_U5598 , P2_U5658 , P2_U3084 );
nand NAND2_6294 ( P2_U5599 , P2_U3483 , P2_U5537 );
nand NAND2_6295 ( P2_U5600 , P2_U3929 , P2_U3084 );
nand NAND2_6296 ( P2_U5601 , P2_U5658 , P2_U3071 );
nand NAND2_6297 ( P2_U5602 , P2_U3480 , P2_U5537 );
nand NAND2_6298 ( P2_U5603 , P2_U3929 , P2_U3071 );
nand NAND2_6299 ( P2_U5604 , P2_U5658 , P2_U3075 );
nand NAND2_6300 ( P2_U5605 , P2_U3477 , P2_U5537 );
nand NAND2_6301 ( P2_U5606 , P2_U3929 , P2_U3075 );
nand NAND2_6302 ( P2_U5607 , P2_U5658 , P2_U3076 );
nand NAND2_6303 ( P2_U5608 , P2_U3474 , P2_U5537 );
nand NAND2_6304 ( P2_U5609 , P2_U3929 , P2_U3076 );
nand NAND2_6305 ( P2_U5610 , P2_U5658 , P2_U3081 );
nand NAND2_6306 ( P2_U5611 , P2_U3471 , P2_U5537 );
nand NAND2_6307 ( P2_U5612 , P2_U3929 , P2_U3081 );
nand NAND2_6308 ( P2_U5613 , P2_U5658 , P2_U3082 );
nand NAND2_6309 ( P2_U5614 , P2_U3468 , P2_U5537 );
nand NAND2_6310 ( P2_U5615 , P2_U3929 , P2_U3082 );
nand NAND2_6311 ( P2_U5616 , P2_U5658 , P2_U3074 );
nand NAND2_6312 ( P2_U5617 , P2_U3465 , P2_U5537 );
nand NAND2_6313 ( P2_U5618 , P2_U3929 , P2_U3074 );
nand NAND2_6314 ( P2_U5619 , P2_U5658 , P2_U3065 );
nand NAND2_6315 ( P2_U5620 , P2_U3462 , P2_U5537 );
nand NAND2_6316 ( P2_U5621 , P2_U3929 , P2_U3065 );
nand NAND2_6317 ( P2_U5622 , P2_U5658 , P2_U3064 );
nand NAND2_6318 ( P2_U5623 , P2_U3459 , P2_U5537 );
nand NAND2_6319 ( P2_U5624 , P2_U3929 , P2_U3064 );
nand NAND2_6320 ( P2_U5625 , P2_U5658 , P2_U3085 );
nand NAND2_6321 ( P2_U5626 , P2_U3432 , P2_U5537 );
nand NAND2_6322 ( P2_U5627 , P2_U3929 , P2_U3080 );
nand NAND2_6323 ( P2_U5628 , P2_U5658 , P2_U3079 );
nand NAND2_6324 ( P2_U5629 , P2_U3427 , P2_U5537 );
nand NAND2_6325 ( P2_U5630 , P2_U3929 , P2_U3079 );
nand NAND2_6326 ( P2_U5631 , P2_U5163 , P2_U3088 );
nand NAND2_6327 ( P2_U5632 , P2_U3828 , P2_U5461 );
nand NAND2_6328 ( P2_U5633 , P2_U3972 , P2_U3406 );
nand NAND2_6329 ( P2_U5634 , P2_U3946 , P2_U3972 );
nand NAND2_6330 ( P2_U5635 , P2_U5633 , P2_U3970 );
nand NAND2_6331 ( P2_U5636 , P2_U5634 , P2_U3971 );
nand NAND2_6332 ( P2_U5637 , P2_U3054 , P2_U3945 );
nand NAND2_6333 ( P2_U5638 , P2_U3054 , P2_U3330 );
nand NAND2_6334 ( P2_U5639 , P2_U3961 , P2_U3023 );
nand NAND2_6335 ( P2_U5640 , P2_U3787 , P2_U5163 );
nand NAND4_6336 ( P2_U5641 , P2_U6150 , P2_U6149 , P2_U5163 , P2_U3917 );
nand NAND2_6337 ( P2_U5642 , P2_U5652 , P2_U5646 );
nand NAND2_6338 ( P2_U5643 , P2_U3415 , P2_U3347 );
nand NAND2_6339 ( P2_U5644 , P2_IR_REG_24_ , P2_U3879 );
nand NAND2_6340 ( P2_U5645 , P2_IR_REG_31_ , P2_SUB_1108_U14 );
not NOT1_6341 ( P2_U5646 , P2_U3412 );
nand NAND2_6342 ( P2_U5647 , P2_IR_REG_25_ , P2_U3879 );
nand NAND2_6343 ( P2_U5648 , P2_IR_REG_31_ , P2_SUB_1108_U112 );
not NOT1_6344 ( P2_U5649 , P2_U3413 );
nand NAND2_6345 ( P2_U5650 , P2_IR_REG_26_ , P2_U3879 );
nand NAND2_6346 ( P2_U5651 , P2_IR_REG_31_ , P2_SUB_1108_U15 );
not NOT1_6347 ( P2_U5652 , P2_U3414 );
nand NAND2_6348 ( P2_U5653 , P2_U5646 , P2_B_REG );
nand NAND2_6349 ( P2_U5654 , P2_U3412 , P2_U3331 );
nand NAND2_6350 ( P2_U5655 , P2_U5654 , P2_U5653 );
nand NAND2_6351 ( P2_U5656 , P2_IR_REG_23_ , P2_U3879 );
nand NAND2_6352 ( P2_U5657 , P2_IR_REG_31_ , P2_SUB_1108_U13 );
not NOT1_6353 ( P2_U5658 , P2_U3415 );
nand NAND2_6354 ( P2_U5659 , P2_D_REG_0_ , P2_U3880 );
nand NAND2_6355 ( P2_U5660 , P2_U3967 , P2_U4077 );
nand NAND2_6356 ( P2_U5661 , P2_D_REG_1_ , P2_U3880 );
nand NAND2_6357 ( P2_U5662 , P2_U3967 , P2_U4078 );
nand NAND2_6358 ( P2_U5663 , P2_IR_REG_22_ , P2_U3879 );
nand NAND2_6359 ( P2_U5664 , P2_IR_REG_31_ , P2_SUB_1108_U114 );
not NOT1_6360 ( P2_U5665 , P2_U3420 );
nand NAND2_6361 ( P2_U5666 , P2_IR_REG_19_ , P2_U3879 );
nand NAND2_6362 ( P2_U5667 , P2_IR_REG_31_ , P2_SUB_1108_U123 );
not NOT1_6363 ( P2_U5668 , P2_U3424 );
nand NAND2_6364 ( P2_U5669 , P2_IR_REG_20_ , P2_U3879 );
nand NAND2_6365 ( P2_U5670 , P2_IR_REG_31_ , P2_SUB_1108_U119 );
not NOT1_6366 ( P2_U5671 , P2_U3418 );
nand NAND2_6367 ( P2_U5672 , P2_IR_REG_21_ , P2_U3879 );
nand NAND2_6368 ( P2_U5673 , P2_IR_REG_31_ , P2_SUB_1108_U116 );
not NOT1_6369 ( P2_U5674 , P2_U3419 );
nand NAND2_6370 ( P2_U5675 , P2_IR_REG_30_ , P2_U3879 );
nand NAND2_6371 ( P2_U5676 , P2_IR_REG_31_ , P2_SUB_1108_U104 );
not NOT1_6372 ( P2_U5677 , P2_U3421 );
nand NAND2_6373 ( P2_U5678 , P2_IR_REG_29_ , P2_U3879 );
nand NAND2_6374 ( P2_U5679 , P2_IR_REG_31_ , P2_SUB_1108_U16 );
not NOT1_6375 ( P2_U5680 , P2_U3422 );
nand NAND2_6376 ( P2_U5681 , P2_IR_REG_28_ , P2_U3879 );
nand NAND2_6377 ( P2_U5682 , P2_IR_REG_31_ , P2_SUB_1108_U107 );
not NOT1_6378 ( P2_U5683 , P2_U3423 );
nand NAND2_6379 ( P2_U5684 , P2_IR_REG_0_ , P2_U3879 );
nand NAND2_6380 ( P2_U5685 , P2_IR_REG_31_ , P2_IR_REG_0_ );
nand NAND2_6381 ( P2_U5686 , P2_IR_REG_27_ , P2_U3879 );
nand NAND2_6382 ( P2_U5687 , P2_IR_REG_31_ , P2_SUB_1108_U110 );
not NOT1_6383 ( P2_U5688 , P2_U3426 );
nand NAND2_6384 ( P2_U5689 , U93 , P2_U3347 );
nand NAND2_6385 ( P2_U5690 , P2_U3425 , P2_U3945 );
not NOT1_6386 ( P2_U5691 , P2_U3427 );
nand NAND2_6387 ( P2_U5692 , P2_U3420 , P2_U5674 );
nand NAND2_6388 ( P2_U5693 , P2_U5665 , P2_U4109 );
nand NAND2_6389 ( P2_U5694 , P2_D_REG_1_ , P2_U4076 );
nand NAND2_6390 ( P2_U5695 , P2_U4078 , P2_U3333 );
not NOT1_6391 ( P2_U5696 , P2_U3429 );
nand NAND2_6392 ( P2_U5697 , P2_U5642 , P2_U3333 );
nand NAND2_6393 ( P2_U5698 , P2_D_REG_0_ , P2_U4076 );
not NOT1_6394 ( P2_U5699 , P2_U3428 );
nand NAND2_6395 ( P2_U5700 , P2_REG0_REG_0_ , P2_U3881 );
nand NAND2_6396 ( P2_U5701 , P2_U3966 , P2_U4129 );
nand NAND2_6397 ( P2_U5702 , P2_IR_REG_1_ , P2_U3879 );
nand NAND2_6398 ( P2_U5703 , P2_IR_REG_31_ , P2_SUB_1108_U42 );
nand NAND2_6399 ( P2_U5704 , U82 , P2_U3347 );
nand NAND2_6400 ( P2_U5705 , P2_U3431 , P2_U3945 );
not NOT1_6401 ( P2_U5706 , P2_U3432 );
nand NAND2_6402 ( P2_U5707 , P2_REG0_REG_1_ , P2_U3881 );
nand NAND2_6403 ( P2_U5708 , P2_U3966 , P2_U4153 );
nand NAND2_6404 ( P2_U5709 , P2_IR_REG_2_ , P2_U3879 );
nand NAND2_6405 ( P2_U5710 , P2_IR_REG_31_ , P2_SUB_1108_U17 );
nand NAND2_6406 ( P2_U5711 , U71 , P2_U3347 );
nand NAND2_6407 ( P2_U5712 , P2_U3434 , P2_U3945 );
not NOT1_6408 ( P2_U5713 , P2_U3435 );
nand NAND2_6409 ( P2_U5714 , P2_REG0_REG_2_ , P2_U3881 );
nand NAND2_6410 ( P2_U5715 , P2_U3966 , P2_U4172 );
nand NAND2_6411 ( P2_U5716 , P2_IR_REG_3_ , P2_U3879 );
nand NAND2_6412 ( P2_U5717 , P2_IR_REG_31_ , P2_SUB_1108_U18 );
nand NAND2_6413 ( P2_U5718 , U68 , P2_U3347 );
nand NAND2_6414 ( P2_U5719 , P2_U3437 , P2_U3945 );
not NOT1_6415 ( P2_U5720 , P2_U3438 );
nand NAND2_6416 ( P2_U5721 , P2_REG0_REG_3_ , P2_U3881 );
nand NAND2_6417 ( P2_U5722 , P2_U3966 , P2_U4191 );
nand NAND2_6418 ( P2_U5723 , P2_IR_REG_4_ , P2_U3879 );
nand NAND2_6419 ( P2_U5724 , P2_IR_REG_31_ , P2_SUB_1108_U19 );
nand NAND2_6420 ( P2_U5725 , U67 , P2_U3347 );
nand NAND2_6421 ( P2_U5726 , P2_U3440 , P2_U3945 );
not NOT1_6422 ( P2_U5727 , P2_U3441 );
nand NAND2_6423 ( P2_U5728 , P2_REG0_REG_4_ , P2_U3881 );
nand NAND2_6424 ( P2_U5729 , P2_U3966 , P2_U4210 );
nand NAND2_6425 ( P2_U5730 , P2_IR_REG_5_ , P2_U3879 );
nand NAND2_6426 ( P2_U5731 , P2_IR_REG_31_ , P2_SUB_1108_U101 );
nand NAND2_6427 ( P2_U5732 , U66 , P2_U3347 );
nand NAND2_6428 ( P2_U5733 , P2_U3443 , P2_U3945 );
not NOT1_6429 ( P2_U5734 , P2_U3444 );
nand NAND2_6430 ( P2_U5735 , P2_REG0_REG_5_ , P2_U3881 );
nand NAND2_6431 ( P2_U5736 , P2_U3966 , P2_U4229 );
nand NAND2_6432 ( P2_U5737 , P2_IR_REG_6_ , P2_U3879 );
nand NAND2_6433 ( P2_U5738 , P2_IR_REG_31_ , P2_SUB_1108_U20 );
nand NAND2_6434 ( P2_U5739 , U65 , P2_U3347 );
nand NAND2_6435 ( P2_U5740 , P2_U3446 , P2_U3945 );
not NOT1_6436 ( P2_U5741 , P2_U3447 );
nand NAND2_6437 ( P2_U5742 , P2_REG0_REG_6_ , P2_U3881 );
nand NAND2_6438 ( P2_U5743 , P2_U3966 , P2_U4248 );
nand NAND2_6439 ( P2_U5744 , P2_IR_REG_7_ , P2_U3879 );
nand NAND2_6440 ( P2_U5745 , P2_IR_REG_31_ , P2_SUB_1108_U21 );
nand NAND2_6441 ( P2_U5746 , U64 , P2_U3347 );
nand NAND2_6442 ( P2_U5747 , P2_U3449 , P2_U3945 );
not NOT1_6443 ( P2_U5748 , P2_U3450 );
nand NAND2_6444 ( P2_U5749 , P2_REG0_REG_7_ , P2_U3881 );
nand NAND2_6445 ( P2_U5750 , P2_U3966 , P2_U4267 );
nand NAND2_6446 ( P2_U5751 , P2_IR_REG_8_ , P2_U3879 );
nand NAND2_6447 ( P2_U5752 , P2_IR_REG_31_ , P2_SUB_1108_U22 );
nand NAND2_6448 ( P2_U5753 , U63 , P2_U3347 );
nand NAND2_6449 ( P2_U5754 , P2_U3452 , P2_U3945 );
not NOT1_6450 ( P2_U5755 , P2_U3453 );
nand NAND2_6451 ( P2_U5756 , P2_REG0_REG_8_ , P2_U3881 );
nand NAND2_6452 ( P2_U5757 , P2_U3966 , P2_U4286 );
nand NAND2_6453 ( P2_U5758 , P2_IR_REG_9_ , P2_U3879 );
nand NAND2_6454 ( P2_U5759 , P2_IR_REG_31_ , P2_SUB_1108_U99 );
nand NAND2_6455 ( P2_U5760 , U62 , P2_U3347 );
nand NAND2_6456 ( P2_U5761 , P2_U3455 , P2_U3945 );
not NOT1_6457 ( P2_U5762 , P2_U3456 );
nand NAND2_6458 ( P2_U5763 , P2_REG0_REG_9_ , P2_U3881 );
nand NAND2_6459 ( P2_U5764 , P2_U3966 , P2_U4305 );
nand NAND2_6460 ( P2_U5765 , P2_IR_REG_10_ , P2_U3879 );
nand NAND2_6461 ( P2_U5766 , P2_IR_REG_31_ , P2_SUB_1108_U6 );
nand NAND2_6462 ( P2_U5767 , U92 , P2_U3347 );
nand NAND2_6463 ( P2_U5768 , P2_U3458 , P2_U3945 );
not NOT1_6464 ( P2_U5769 , P2_U3459 );
nand NAND2_6465 ( P2_U5770 , P2_REG0_REG_10_ , P2_U3881 );
nand NAND2_6466 ( P2_U5771 , P2_U3966 , P2_U4324 );
nand NAND2_6467 ( P2_U5772 , P2_IR_REG_11_ , P2_U3879 );
nand NAND2_6468 ( P2_U5773 , P2_IR_REG_31_ , P2_SUB_1108_U7 );
nand NAND2_6469 ( P2_U5774 , U91 , P2_U3347 );
nand NAND2_6470 ( P2_U5775 , P2_U3461 , P2_U3945 );
not NOT1_6471 ( P2_U5776 , P2_U3462 );
nand NAND2_6472 ( P2_U5777 , P2_REG0_REG_11_ , P2_U3881 );
nand NAND2_6473 ( P2_U5778 , P2_U3966 , P2_U4343 );
nand NAND2_6474 ( P2_U5779 , P2_IR_REG_12_ , P2_U3879 );
nand NAND2_6475 ( P2_U5780 , P2_IR_REG_31_ , P2_SUB_1108_U8 );
nand NAND2_6476 ( P2_U5781 , U90 , P2_U3347 );
nand NAND2_6477 ( P2_U5782 , P2_U3464 , P2_U3945 );
not NOT1_6478 ( P2_U5783 , P2_U3465 );
nand NAND2_6479 ( P2_U5784 , P2_REG0_REG_12_ , P2_U3881 );
nand NAND2_6480 ( P2_U5785 , P2_U3966 , P2_U4362 );
nand NAND2_6481 ( P2_U5786 , P2_IR_REG_13_ , P2_U3879 );
nand NAND2_6482 ( P2_U5787 , P2_IR_REG_31_ , P2_SUB_1108_U127 );
nand NAND2_6483 ( P2_U5788 , U89 , P2_U3347 );
nand NAND2_6484 ( P2_U5789 , P2_U3467 , P2_U3945 );
not NOT1_6485 ( P2_U5790 , P2_U3468 );
nand NAND2_6486 ( P2_U5791 , P2_REG0_REG_13_ , P2_U3881 );
nand NAND2_6487 ( P2_U5792 , P2_U3966 , P2_U4381 );
nand NAND2_6488 ( P2_U5793 , P2_IR_REG_14_ , P2_U3879 );
nand NAND2_6489 ( P2_U5794 , P2_IR_REG_31_ , P2_SUB_1108_U9 );
nand NAND2_6490 ( P2_U5795 , U88 , P2_U3347 );
nand NAND2_6491 ( P2_U5796 , P2_U3470 , P2_U3945 );
not NOT1_6492 ( P2_U5797 , P2_U3471 );
nand NAND2_6493 ( P2_U5798 , P2_REG0_REG_14_ , P2_U3881 );
nand NAND2_6494 ( P2_U5799 , P2_U3966 , P2_U4400 );
nand NAND2_6495 ( P2_U5800 , P2_IR_REG_15_ , P2_U3879 );
nand NAND2_6496 ( P2_U5801 , P2_IR_REG_31_ , P2_SUB_1108_U10 );
nand NAND2_6497 ( P2_U5802 , U87 , P2_U3347 );
nand NAND2_6498 ( P2_U5803 , P2_U3473 , P2_U3945 );
not NOT1_6499 ( P2_U5804 , P2_U3474 );
nand NAND2_6500 ( P2_U5805 , P2_REG0_REG_15_ , P2_U3881 );
nand NAND2_6501 ( P2_U5806 , P2_U3966 , P2_U4419 );
nand NAND2_6502 ( P2_U5807 , P2_IR_REG_16_ , P2_U3879 );
nand NAND2_6503 ( P2_U5808 , P2_IR_REG_31_ , P2_SUB_1108_U11 );
nand NAND2_6504 ( P2_U5809 , U86 , P2_U3347 );
nand NAND2_6505 ( P2_U5810 , P2_U3476 , P2_U3945 );
not NOT1_6506 ( P2_U5811 , P2_U3477 );
nand NAND2_6507 ( P2_U5812 , P2_REG0_REG_16_ , P2_U3881 );
nand NAND2_6508 ( P2_U5813 , P2_U3966 , P2_U4438 );
nand NAND2_6509 ( P2_U5814 , P2_IR_REG_17_ , P2_U3879 );
nand NAND2_6510 ( P2_U5815 , P2_IR_REG_31_ , P2_SUB_1108_U125 );
nand NAND2_6511 ( P2_U5816 , U85 , P2_U3347 );
nand NAND2_6512 ( P2_U5817 , P2_U3479 , P2_U3945 );
not NOT1_6513 ( P2_U5818 , P2_U3480 );
nand NAND2_6514 ( P2_U5819 , P2_REG0_REG_17_ , P2_U3881 );
nand NAND2_6515 ( P2_U5820 , P2_U3966 , P2_U4457 );
nand NAND2_6516 ( P2_U5821 , P2_IR_REG_18_ , P2_U3879 );
nand NAND2_6517 ( P2_U5822 , P2_IR_REG_31_ , P2_SUB_1108_U12 );
nand NAND2_6518 ( P2_U5823 , U84 , P2_U3347 );
nand NAND2_6519 ( P2_U5824 , P2_U3482 , P2_U3945 );
not NOT1_6520 ( P2_U5825 , P2_U3483 );
nand NAND2_6521 ( P2_U5826 , P2_REG0_REG_18_ , P2_U3881 );
nand NAND2_6522 ( P2_U5827 , P2_U3966 , P2_U4476 );
nand NAND2_6523 ( P2_U5828 , U83 , P2_U3347 );
nand NAND2_6524 ( P2_U5829 , P2_U3424 , P2_U3945 );
not NOT1_6525 ( P2_U5830 , P2_U3485 );
nand NAND2_6526 ( P2_U5831 , P2_REG0_REG_19_ , P2_U3881 );
nand NAND2_6527 ( P2_U5832 , P2_U3966 , P2_U4495 );
nand NAND2_6528 ( P2_U5833 , P2_REG0_REG_20_ , P2_U3881 );
nand NAND2_6529 ( P2_U5834 , P2_U3966 , P2_U4514 );
nand NAND2_6530 ( P2_U5835 , P2_REG0_REG_21_ , P2_U3881 );
nand NAND2_6531 ( P2_U5836 , P2_U3966 , P2_U4533 );
nand NAND2_6532 ( P2_U5837 , P2_REG0_REG_22_ , P2_U3881 );
nand NAND2_6533 ( P2_U5838 , P2_U3966 , P2_U4552 );
nand NAND2_6534 ( P2_U5839 , P2_REG0_REG_23_ , P2_U3881 );
nand NAND2_6535 ( P2_U5840 , P2_U3966 , P2_U4571 );
nand NAND2_6536 ( P2_U5841 , P2_REG0_REG_24_ , P2_U3881 );
nand NAND2_6537 ( P2_U5842 , P2_U3966 , P2_U4590 );
nand NAND2_6538 ( P2_U5843 , P2_REG0_REG_25_ , P2_U3881 );
nand NAND2_6539 ( P2_U5844 , P2_U3966 , P2_U4609 );
nand NAND2_6540 ( P2_U5845 , P2_REG0_REG_26_ , P2_U3881 );
nand NAND2_6541 ( P2_U5846 , P2_U3966 , P2_U4628 );
nand NAND2_6542 ( P2_U5847 , P2_REG0_REG_27_ , P2_U3881 );
nand NAND2_6543 ( P2_U5848 , P2_U3966 , P2_U4647 );
nand NAND2_6544 ( P2_U5849 , P2_REG0_REG_28_ , P2_U3881 );
nand NAND2_6545 ( P2_U5850 , P2_U3966 , P2_U4666 );
nand NAND2_6546 ( P2_U5851 , P2_REG0_REG_29_ , P2_U3881 );
nand NAND2_6547 ( P2_U5852 , P2_U3966 , P2_U4686 );
nand NAND2_6548 ( P2_U5853 , P2_REG0_REG_30_ , P2_U3881 );
nand NAND2_6549 ( P2_U5854 , P2_U3966 , P2_U4693 );
nand NAND2_6550 ( P2_U5855 , P2_REG0_REG_31_ , P2_U3881 );
nand NAND2_6551 ( P2_U5856 , P2_U3966 , P2_U4696 );
nand NAND2_6552 ( P2_U5857 , P2_REG1_REG_0_ , P2_U3882 );
nand NAND2_6553 ( P2_U5858 , P2_U3965 , P2_U4129 );
nand NAND2_6554 ( P2_U5859 , P2_REG1_REG_1_ , P2_U3882 );
nand NAND2_6555 ( P2_U5860 , P2_U3965 , P2_U4153 );
nand NAND2_6556 ( P2_U5861 , P2_REG1_REG_2_ , P2_U3882 );
nand NAND2_6557 ( P2_U5862 , P2_U3965 , P2_U4172 );
nand NAND2_6558 ( P2_U5863 , P2_REG1_REG_3_ , P2_U3882 );
nand NAND2_6559 ( P2_U5864 , P2_U3965 , P2_U4191 );
nand NAND2_6560 ( P2_U5865 , P2_REG1_REG_4_ , P2_U3882 );
nand NAND2_6561 ( P2_U5866 , P2_U3965 , P2_U4210 );
nand NAND2_6562 ( P2_U5867 , P2_REG1_REG_5_ , P2_U3882 );
nand NAND2_6563 ( P2_U5868 , P2_U3965 , P2_U4229 );
nand NAND2_6564 ( P2_U5869 , P2_REG1_REG_6_ , P2_U3882 );
nand NAND2_6565 ( P2_U5870 , P2_U3965 , P2_U4248 );
nand NAND2_6566 ( P2_U5871 , P2_REG1_REG_7_ , P2_U3882 );
nand NAND2_6567 ( P2_U5872 , P2_U3965 , P2_U4267 );
nand NAND2_6568 ( P2_U5873 , P2_REG1_REG_8_ , P2_U3882 );
nand NAND2_6569 ( P2_U5874 , P2_U3965 , P2_U4286 );
nand NAND2_6570 ( P2_U5875 , P2_REG1_REG_9_ , P2_U3882 );
nand NAND2_6571 ( P2_U5876 , P2_U3965 , P2_U4305 );
nand NAND2_6572 ( P2_U5877 , P2_REG1_REG_10_ , P2_U3882 );
nand NAND2_6573 ( P2_U5878 , P2_U3965 , P2_U4324 );
nand NAND2_6574 ( P2_U5879 , P2_REG1_REG_11_ , P2_U3882 );
nand NAND2_6575 ( P2_U5880 , P2_U3965 , P2_U4343 );
nand NAND2_6576 ( P2_U5881 , P2_REG1_REG_12_ , P2_U3882 );
nand NAND2_6577 ( P2_U5882 , P2_U3965 , P2_U4362 );
nand NAND2_6578 ( P2_U5883 , P2_REG1_REG_13_ , P2_U3882 );
nand NAND2_6579 ( P2_U5884 , P2_U3965 , P2_U4381 );
nand NAND2_6580 ( P2_U5885 , P2_REG1_REG_14_ , P2_U3882 );
nand NAND2_6581 ( P2_U5886 , P2_U3965 , P2_U4400 );
nand NAND2_6582 ( P2_U5887 , P2_REG1_REG_15_ , P2_U3882 );
nand NAND2_6583 ( P2_U5888 , P2_U3965 , P2_U4419 );
nand NAND2_6584 ( P2_U5889 , P2_REG1_REG_16_ , P2_U3882 );
nand NAND2_6585 ( P2_U5890 , P2_U3965 , P2_U4438 );
nand NAND2_6586 ( P2_U5891 , P2_REG1_REG_17_ , P2_U3882 );
nand NAND2_6587 ( P2_U5892 , P2_U3965 , P2_U4457 );
nand NAND2_6588 ( P2_U5893 , P2_REG1_REG_18_ , P2_U3882 );
nand NAND2_6589 ( P2_U5894 , P2_U3965 , P2_U4476 );
nand NAND2_6590 ( P2_U5895 , P2_REG1_REG_19_ , P2_U3882 );
nand NAND2_6591 ( P2_U5896 , P2_U3965 , P2_U4495 );
nand NAND2_6592 ( P2_U5897 , P2_REG1_REG_20_ , P2_U3882 );
nand NAND2_6593 ( P2_U5898 , P2_U3965 , P2_U4514 );
nand NAND2_6594 ( P2_U5899 , P2_REG1_REG_21_ , P2_U3882 );
nand NAND2_6595 ( P2_U5900 , P2_U3965 , P2_U4533 );
nand NAND2_6596 ( P2_U5901 , P2_REG1_REG_22_ , P2_U3882 );
nand NAND2_6597 ( P2_U5902 , P2_U3965 , P2_U4552 );
nand NAND2_6598 ( P2_U5903 , P2_REG1_REG_23_ , P2_U3882 );
nand NAND2_6599 ( P2_U5904 , P2_U3965 , P2_U4571 );
nand NAND2_6600 ( P2_U5905 , P2_REG1_REG_24_ , P2_U3882 );
nand NAND2_6601 ( P2_U5906 , P2_U3965 , P2_U4590 );
nand NAND2_6602 ( P2_U5907 , P2_REG1_REG_25_ , P2_U3882 );
nand NAND2_6603 ( P2_U5908 , P2_U3965 , P2_U4609 );
nand NAND2_6604 ( P2_U5909 , P2_REG1_REG_26_ , P2_U3882 );
nand NAND2_6605 ( P2_U5910 , P2_U3965 , P2_U4628 );
nand NAND2_6606 ( P2_U5911 , P2_REG1_REG_27_ , P2_U3882 );
nand NAND2_6607 ( P2_U5912 , P2_U3965 , P2_U4647 );
nand NAND2_6608 ( P2_U5913 , P2_REG1_REG_28_ , P2_U3882 );
nand NAND2_6609 ( P2_U5914 , P2_U3965 , P2_U4666 );
nand NAND2_6610 ( P2_U5915 , P2_REG1_REG_29_ , P2_U3882 );
nand NAND2_6611 ( P2_U5916 , P2_U3965 , P2_U4686 );
nand NAND2_6612 ( P2_U5917 , P2_REG1_REG_30_ , P2_U3882 );
nand NAND2_6613 ( P2_U5918 , P2_U3965 , P2_U4693 );
nand NAND2_6614 ( P2_U5919 , P2_REG1_REG_31_ , P2_U3882 );
nand NAND2_6615 ( P2_U5920 , P2_U3965 , P2_U4696 );
nand NAND2_6616 ( P2_U5921 , P2_REG2_REG_0_ , P2_U3391 );
nand NAND2_6617 ( P2_U5922 , P2_U3964 , P2_U3348 );
nand NAND2_6618 ( P2_U5923 , P2_REG2_REG_1_ , P2_U3391 );
nand NAND2_6619 ( P2_U5924 , P2_U3964 , P2_U3349 );
nand NAND2_6620 ( P2_U5925 , P2_REG2_REG_2_ , P2_U3391 );
nand NAND2_6621 ( P2_U5926 , P2_U3964 , P2_U3350 );
nand NAND2_6622 ( P2_U5927 , P2_REG2_REG_3_ , P2_U3391 );
nand NAND2_6623 ( P2_U5928 , P2_U3964 , P2_U3351 );
nand NAND2_6624 ( P2_U5929 , P2_REG2_REG_4_ , P2_U3391 );
nand NAND2_6625 ( P2_U5930 , P2_U3964 , P2_U3352 );
nand NAND2_6626 ( P2_U5931 , P2_REG2_REG_5_ , P2_U3391 );
nand NAND2_6627 ( P2_U5932 , P2_U3964 , P2_U3353 );
nand NAND2_6628 ( P2_U5933 , P2_REG2_REG_6_ , P2_U3391 );
nand NAND2_6629 ( P2_U5934 , P2_U3964 , P2_U3354 );
nand NAND2_6630 ( P2_U5935 , P2_REG2_REG_7_ , P2_U3391 );
nand NAND2_6631 ( P2_U5936 , P2_U3964 , P2_U3355 );
nand NAND2_6632 ( P2_U5937 , P2_REG2_REG_8_ , P2_U3391 );
nand NAND2_6633 ( P2_U5938 , P2_U3964 , P2_U3356 );
nand NAND2_6634 ( P2_U5939 , P2_REG2_REG_9_ , P2_U3391 );
nand NAND2_6635 ( P2_U5940 , P2_U3964 , P2_U3357 );
nand NAND2_6636 ( P2_U5941 , P2_REG2_REG_10_ , P2_U3391 );
nand NAND2_6637 ( P2_U5942 , P2_U3964 , P2_U3358 );
nand NAND2_6638 ( P2_U5943 , P2_REG2_REG_11_ , P2_U3391 );
nand NAND2_6639 ( P2_U5944 , P2_U3964 , P2_U3359 );
nand NAND2_6640 ( P2_U5945 , P2_REG2_REG_12_ , P2_U3391 );
nand NAND2_6641 ( P2_U5946 , P2_U3964 , P2_U3360 );
nand NAND2_6642 ( P2_U5947 , P2_REG2_REG_13_ , P2_U3391 );
nand NAND2_6643 ( P2_U5948 , P2_U3964 , P2_U3361 );
nand NAND2_6644 ( P2_U5949 , P2_REG2_REG_14_ , P2_U3391 );
nand NAND2_6645 ( P2_U5950 , P2_U3964 , P2_U3362 );
nand NAND2_6646 ( P2_U5951 , P2_REG2_REG_15_ , P2_U3391 );
nand NAND2_6647 ( P2_U5952 , P2_U3964 , P2_U3363 );
nand NAND2_6648 ( P2_U5953 , P2_REG2_REG_16_ , P2_U3391 );
nand NAND2_6649 ( P2_U5954 , P2_U3964 , P2_U3364 );
nand NAND2_6650 ( P2_U5955 , P2_REG2_REG_17_ , P2_U3391 );
nand NAND2_6651 ( P2_U5956 , P2_U3964 , P2_U3365 );
nand NAND2_6652 ( P2_U5957 , P2_REG2_REG_18_ , P2_U3391 );
nand NAND2_6653 ( P2_U5958 , P2_U3964 , P2_U3366 );
nand NAND2_6654 ( P2_U5959 , P2_REG2_REG_19_ , P2_U3391 );
nand NAND2_6655 ( P2_U5960 , P2_U3964 , P2_U3367 );
nand NAND2_6656 ( P2_U5961 , P2_REG2_REG_20_ , P2_U3391 );
nand NAND2_6657 ( P2_U5962 , P2_U3964 , P2_U3369 );
nand NAND2_6658 ( P2_U5963 , P2_REG2_REG_21_ , P2_U3391 );
nand NAND2_6659 ( P2_U5964 , P2_U3964 , P2_U3371 );
nand NAND2_6660 ( P2_U5965 , P2_REG2_REG_22_ , P2_U3391 );
nand NAND2_6661 ( P2_U5966 , P2_U3964 , P2_U3373 );
nand NAND2_6662 ( P2_U5967 , P2_REG2_REG_23_ , P2_U3391 );
nand NAND2_6663 ( P2_U5968 , P2_U3964 , P2_U3375 );
nand NAND2_6664 ( P2_U5969 , P2_REG2_REG_24_ , P2_U3391 );
nand NAND2_6665 ( P2_U5970 , P2_U3964 , P2_U3377 );
nand NAND2_6666 ( P2_U5971 , P2_REG2_REG_25_ , P2_U3391 );
nand NAND2_6667 ( P2_U5972 , P2_U3964 , P2_U3379 );
nand NAND2_6668 ( P2_U5973 , P2_REG2_REG_26_ , P2_U3391 );
nand NAND2_6669 ( P2_U5974 , P2_U3964 , P2_U3381 );
nand NAND2_6670 ( P2_U5975 , P2_REG2_REG_27_ , P2_U3391 );
nand NAND2_6671 ( P2_U5976 , P2_U3964 , P2_U3383 );
nand NAND2_6672 ( P2_U5977 , P2_REG2_REG_28_ , P2_U3391 );
nand NAND2_6673 ( P2_U5978 , P2_U3964 , P2_U3385 );
nand NAND2_6674 ( P2_U5979 , P2_REG2_REG_29_ , P2_U3391 );
nand NAND2_6675 ( P2_U5980 , P2_U3964 , P2_U3387 );
nand NAND2_6676 ( P2_U5981 , P2_REG2_REG_30_ , P2_U3391 );
nand NAND2_6677 ( P2_U5982 , P2_U3968 , P2_U3964 );
nand NAND2_6678 ( P2_U5983 , P2_REG2_REG_31_ , P2_U3391 );
nand NAND2_6679 ( P2_U5984 , P2_U3968 , P2_U3964 );
nand NAND2_6680 ( P2_U5985 , P2_DATAO_REG_0_ , P2_U3400 );
nand NAND2_6681 ( P2_U5986 , P2_U3947 , P2_U3079 );
nand NAND2_6682 ( P2_U5987 , P2_DATAO_REG_1_ , P2_U3400 );
nand NAND2_6683 ( P2_U5988 , P2_U3947 , P2_U3080 );
nand NAND2_6684 ( P2_U5989 , P2_DATAO_REG_2_ , P2_U3400 );
nand NAND2_6685 ( P2_U5990 , P2_U3947 , P2_U3070 );
nand NAND2_6686 ( P2_U5991 , P2_DATAO_REG_3_ , P2_U3400 );
nand NAND2_6687 ( P2_U5992 , P2_U3947 , P2_U3066 );
nand NAND2_6688 ( P2_U5993 , P2_DATAO_REG_4_ , P2_U3400 );
nand NAND2_6689 ( P2_U5994 , P2_U3947 , P2_U3062 );
nand NAND2_6690 ( P2_U5995 , P2_DATAO_REG_5_ , P2_U3400 );
nand NAND2_6691 ( P2_U5996 , P2_U3947 , P2_U3069 );
nand NAND2_6692 ( P2_U5997 , P2_DATAO_REG_6_ , P2_U3400 );
nand NAND2_6693 ( P2_U5998 , P2_U3947 , P2_U3073 );
nand NAND2_6694 ( P2_U5999 , P2_DATAO_REG_7_ , P2_U3400 );
nand NAND2_6695 ( P2_U6000 , P2_U3947 , P2_U3072 );
nand NAND2_6696 ( P2_U6001 , P2_DATAO_REG_8_ , P2_U3400 );
nand NAND2_6697 ( P2_U6002 , P2_U3947 , P2_U3086 );
nand NAND2_6698 ( P2_U6003 , P2_DATAO_REG_9_ , P2_U3400 );
nand NAND2_6699 ( P2_U6004 , P2_U3947 , P2_U3085 );
nand NAND2_6700 ( P2_U6005 , P2_DATAO_REG_10_ , P2_U3400 );
nand NAND2_6701 ( P2_U6006 , P2_U3947 , P2_U3064 );
nand NAND2_6702 ( P2_U6007 , P2_DATAO_REG_11_ , P2_U3400 );
nand NAND2_6703 ( P2_U6008 , P2_U3947 , P2_U3065 );
nand NAND2_6704 ( P2_U6009 , P2_DATAO_REG_12_ , P2_U3400 );
nand NAND2_6705 ( P2_U6010 , P2_U3947 , P2_U3074 );
nand NAND2_6706 ( P2_U6011 , P2_DATAO_REG_13_ , P2_U3400 );
nand NAND2_6707 ( P2_U6012 , P2_U3947 , P2_U3082 );
nand NAND2_6708 ( P2_U6013 , P2_DATAO_REG_14_ , P2_U3400 );
nand NAND2_6709 ( P2_U6014 , P2_U3947 , P2_U3081 );
nand NAND2_6710 ( P2_U6015 , P2_DATAO_REG_15_ , P2_U3400 );
nand NAND2_6711 ( P2_U6016 , P2_U3947 , P2_U3076 );
nand NAND2_6712 ( P2_U6017 , P2_DATAO_REG_16_ , P2_U3400 );
nand NAND2_6713 ( P2_U6018 , P2_U3947 , P2_U3075 );
nand NAND2_6714 ( P2_U6019 , P2_DATAO_REG_17_ , P2_U3400 );
nand NAND2_6715 ( P2_U6020 , P2_U3947 , P2_U3071 );
nand NAND2_6716 ( P2_U6021 , P2_DATAO_REG_18_ , P2_U3400 );
nand NAND2_6717 ( P2_U6022 , P2_U3947 , P2_U3084 );
nand NAND2_6718 ( P2_U6023 , P2_DATAO_REG_19_ , P2_U3400 );
nand NAND2_6719 ( P2_U6024 , P2_U3947 , P2_U3083 );
nand NAND2_6720 ( P2_U6025 , P2_DATAO_REG_20_ , P2_U3400 );
nand NAND2_6721 ( P2_U6026 , P2_U3947 , P2_U3078 );
nand NAND2_6722 ( P2_U6027 , P2_DATAO_REG_21_ , P2_U3400 );
nand NAND2_6723 ( P2_U6028 , P2_U3947 , P2_U3077 );
nand NAND2_6724 ( P2_U6029 , P2_DATAO_REG_22_ , P2_U3400 );
nand NAND2_6725 ( P2_U6030 , P2_U3947 , P2_U3063 );
nand NAND2_6726 ( P2_U6031 , P2_DATAO_REG_23_ , P2_U3400 );
nand NAND2_6727 ( P2_U6032 , P2_U3947 , P2_U3068 );
nand NAND2_6728 ( P2_U6033 , P2_DATAO_REG_24_ , P2_U3400 );
nand NAND2_6729 ( P2_U6034 , P2_U3947 , P2_U3067 );
nand NAND2_6730 ( P2_U6035 , P2_DATAO_REG_25_ , P2_U3400 );
nand NAND2_6731 ( P2_U6036 , P2_U3947 , P2_U3060 );
nand NAND2_6732 ( P2_U6037 , P2_DATAO_REG_26_ , P2_U3400 );
nand NAND2_6733 ( P2_U6038 , P2_U3947 , P2_U3059 );
nand NAND2_6734 ( P2_U6039 , P2_DATAO_REG_27_ , P2_U3400 );
nand NAND2_6735 ( P2_U6040 , P2_U3947 , P2_U3055 );
nand NAND2_6736 ( P2_U6041 , P2_DATAO_REG_28_ , P2_U3400 );
nand NAND2_6737 ( P2_U6042 , P2_U3947 , P2_U3056 );
nand NAND2_6738 ( P2_U6043 , P2_DATAO_REG_29_ , P2_U3400 );
nand NAND2_6739 ( P2_U6044 , P2_U3947 , P2_U3057 );
nand NAND2_6740 ( P2_U6045 , P2_DATAO_REG_30_ , P2_U3400 );
nand NAND2_6741 ( P2_U6046 , P2_U3947 , P2_U3061 );
nand NAND2_6742 ( P2_U6047 , P2_DATAO_REG_31_ , P2_U3400 );
nand NAND2_6743 ( P2_U6048 , P2_U3947 , P2_U3058 );
nand NAND2_6744 ( P2_U6049 , P2_R1312_U18 , P2_U5157 );
nand NAND2_6745 ( P2_U6050 , P2_U5161 , P2_U3916 );
nand NAND2_6746 ( P2_U6051 , P2_U5658 , P2_U3403 );
nand NAND2_6747 ( P2_U6052 , P2_U3420 , P2_U3415 );
nand NAND2_6748 ( P2_U6053 , P2_U3960 , P2_U3057 );
nand NAND2_6749 ( P2_U6054 , P2_U3386 , P2_U4652 );
nand NAND2_6750 ( P2_U6055 , P2_U6054 , P2_U6053 );
nand NAND2_6751 ( P2_U6056 , P2_U3949 , P2_U3056 );
nand NAND2_6752 ( P2_U6057 , P2_U3384 , P2_U4633 );
nand NAND2_6753 ( P2_U6058 , P2_U6057 , P2_U6056 );
nand NAND2_6754 ( P2_U6059 , P2_U3950 , P2_U3055 );
nand NAND2_6755 ( P2_U6060 , P2_U3382 , P2_U4614 );
nand NAND2_6756 ( P2_U6061 , P2_U6060 , P2_U6059 );
nand NAND2_6757 ( P2_U6062 , P2_U3953 , P2_U3067 );
nand NAND2_6758 ( P2_U6063 , P2_U3376 , P2_U4557 );
nand NAND2_6759 ( P2_U6064 , P2_U6063 , P2_U6062 );
nand NAND2_6760 ( P2_U6065 , P2_U3954 , P2_U3068 );
nand NAND2_6761 ( P2_U6066 , P2_U3374 , P2_U4538 );
nand NAND2_6762 ( P2_U6067 , P2_U6066 , P2_U6065 );
nand NAND2_6763 ( P2_U6068 , P2_U3956 , P2_U3077 );
nand NAND2_6764 ( P2_U6069 , P2_U3370 , P2_U4500 );
nand NAND2_6765 ( P2_U6070 , P2_U6069 , P2_U6068 );
nand NAND2_6766 ( P2_U6071 , P2_U3955 , P2_U3063 );
nand NAND2_6767 ( P2_U6072 , P2_U3372 , P2_U4519 );
nand NAND2_6768 ( P2_U6073 , P2_U6072 , P2_U6071 );
nand NAND2_6769 ( P2_U6074 , P2_U3952 , P2_U3060 );
nand NAND2_6770 ( P2_U6075 , P2_U3378 , P2_U4576 );
nand NAND2_6771 ( P2_U6076 , P2_U6075 , P2_U6074 );
nand NAND2_6772 ( P2_U6077 , P2_U3951 , P2_U3059 );
nand NAND2_6773 ( P2_U6078 , P2_U3380 , P2_U4595 );
nand NAND2_6774 ( P2_U6079 , P2_U6078 , P2_U6077 );
nand NAND2_6775 ( P2_U6080 , P2_U3959 , P2_U3061 );
nand NAND2_6776 ( P2_U6081 , P2_U3388 , P2_U4670 );
nand NAND2_6777 ( P2_U6082 , P2_U6081 , P2_U6080 );
nand NAND2_6778 ( P2_U6083 , P2_U3958 , P2_U3058 );
nand NAND2_6779 ( P2_U6084 , P2_U3389 , P2_U4690 );
nand NAND2_6780 ( P2_U6085 , P2_U6084 , P2_U6083 );
nand NAND2_6781 ( P2_U6086 , P2_U5797 , P2_U4367 );
nand NAND2_6782 ( P2_U6087 , P2_U3471 , P2_U3081 );
nand NAND2_6783 ( P2_U6088 , P2_U6087 , P2_U6086 );
nand NAND2_6784 ( P2_U6089 , P2_U5706 , P2_U4115 );
nand NAND2_6785 ( P2_U6090 , P2_U3432 , P2_U3080 );
nand NAND2_6786 ( P2_U6091 , P2_U6090 , P2_U6089 );
nand NAND2_6787 ( P2_U6092 , P2_U5691 , P2_U4139 );
nand NAND2_6788 ( P2_U6093 , P2_U3427 , P2_U3079 );
nand NAND2_6789 ( P2_U6094 , P2_U6093 , P2_U6092 );
nand NAND2_6790 ( P2_U6095 , P2_U5804 , P2_U4386 );
nand NAND2_6791 ( P2_U6096 , P2_U3474 , P2_U3076 );
nand NAND2_6792 ( P2_U6097 , P2_U6096 , P2_U6095 );
nand NAND2_6793 ( P2_U6098 , P2_U5755 , P2_U4253 );
nand NAND2_6794 ( P2_U6099 , P2_U3453 , P2_U3086 );
nand NAND2_6795 ( P2_U6100 , P2_U6099 , P2_U6098 );
nand NAND2_6796 ( P2_U6101 , P2_U5762 , P2_U4272 );
nand NAND2_6797 ( P2_U6102 , P2_U3456 , P2_U3085 );
nand NAND2_6798 ( P2_U6103 , P2_U6102 , P2_U6101 );
nand NAND2_6799 ( P2_U6104 , P2_U5790 , P2_U4348 );
nand NAND2_6800 ( P2_U6105 , P2_U3468 , P2_U3082 );
nand NAND2_6801 ( P2_U6106 , P2_U6105 , P2_U6104 );
nand NAND2_6802 ( P2_U6107 , P2_U5825 , P2_U4443 );
nand NAND2_6803 ( P2_U6108 , P2_U3483 , P2_U3084 );
nand NAND2_6804 ( P2_U6109 , P2_U6108 , P2_U6107 );
nand NAND2_6805 ( P2_U6110 , P2_U5811 , P2_U4405 );
nand NAND2_6806 ( P2_U6111 , P2_U3477 , P2_U3075 );
nand NAND2_6807 ( P2_U6112 , P2_U6111 , P2_U6110 );
nand NAND2_6808 ( P2_U6113 , P2_U5783 , P2_U4329 );
nand NAND2_6809 ( P2_U6114 , P2_U3465 , P2_U3074 );
nand NAND2_6810 ( P2_U6115 , P2_U6114 , P2_U6113 );
nand NAND2_6811 ( P2_U6116 , P2_U5741 , P2_U4215 );
nand NAND2_6812 ( P2_U6117 , P2_U3447 , P2_U3073 );
nand NAND2_6813 ( P2_U6118 , P2_U6117 , P2_U6116 );
nand NAND2_6814 ( P2_U6119 , P2_U5748 , P2_U4234 );
nand NAND2_6815 ( P2_U6120 , P2_U3450 , P2_U3072 );
nand NAND2_6816 ( P2_U6121 , P2_U6120 , P2_U6119 );
nand NAND2_6817 ( P2_U6122 , P2_U5734 , P2_U4196 );
nand NAND2_6818 ( P2_U6123 , P2_U3444 , P2_U3069 );
nand NAND2_6819 ( P2_U6124 , P2_U6123 , P2_U6122 );
nand NAND2_6820 ( P2_U6125 , P2_U5720 , P2_U4158 );
nand NAND2_6821 ( P2_U6126 , P2_U3438 , P2_U3066 );
nand NAND2_6822 ( P2_U6127 , P2_U6126 , P2_U6125 );
nand NAND2_6823 ( P2_U6128 , P2_U5713 , P2_U4134 );
nand NAND2_6824 ( P2_U6129 , P2_U3435 , P2_U3070 );
nand NAND2_6825 ( P2_U6130 , P2_U6129 , P2_U6128 );
nand NAND2_6826 ( P2_U6131 , P2_U5818 , P2_U4424 );
nand NAND2_6827 ( P2_U6132 , P2_U3480 , P2_U3071 );
nand NAND2_6828 ( P2_U6133 , P2_U6132 , P2_U6131 );
nand NAND2_6829 ( P2_U6134 , P2_U5830 , P2_U4462 );
nand NAND2_6830 ( P2_U6135 , P2_U3485 , P2_U3083 );
nand NAND2_6831 ( P2_U6136 , P2_U6135 , P2_U6134 );
nand NAND2_6832 ( P2_U6137 , P2_U5727 , P2_U4177 );
nand NAND2_6833 ( P2_U6138 , P2_U3441 , P2_U3062 );
nand NAND2_6834 ( P2_U6139 , P2_U6138 , P2_U6137 );
nand NAND2_6835 ( P2_U6140 , P2_U5776 , P2_U4310 );
nand NAND2_6836 ( P2_U6141 , P2_U3462 , P2_U3065 );
nand NAND2_6837 ( P2_U6142 , P2_U6141 , P2_U6140 );
nand NAND2_6838 ( P2_U6143 , P2_U5769 , P2_U4291 );
nand NAND2_6839 ( P2_U6144 , P2_U3459 , P2_U3064 );
nand NAND2_6840 ( P2_U6145 , P2_U6144 , P2_U6143 );
nand NAND2_6841 ( P2_U6146 , P2_U3957 , P2_U3078 );
nand NAND2_6842 ( P2_U6147 , P2_U3368 , P2_U4481 );
nand NAND2_6843 ( P2_U6148 , P2_U6147 , P2_U6146 );
nand NAND2_6844 ( P2_U6149 , P2_U3940 , P2_U5156 );
nand NAND2_6845 ( P2_U6150 , P2_U3942 , P2_U3918 );
nand NAND2_6846 ( P3_R1161_U468 , P3_U3068 , P3_R1161_U60 );
nand NAND2_6847 ( P3_R1161_U467 , P3_R1161_U270 , P3_R1161_U465 );
nand NAND2_6848 ( P3_R1161_U466 , P3_R1161_U360 , P3_R1161_U162 );
nand NAND2_6849 ( P3_R1161_U465 , P3_R1161_U464 , P3_R1161_U463 );
nand NAND2_6850 ( P3_R1161_U464 , P3_U3443 , P3_R1161_U76 );
nand NAND2_6851 ( P3_R1161_U463 , P3_U3081 , P3_R1161_U75 );
nand NAND2_6852 ( P3_R1161_U462 , P3_R1161_U460 , P3_R1161_U316 );
nand NAND2_6853 ( P3_R1161_U461 , P3_R1161_U359 , P3_R1161_U91 );
nand NAND2_6854 ( P3_R1161_U460 , P3_R1161_U459 , P3_R1161_U458 );
nand NAND2_6855 ( P3_R1161_U459 , P3_U3445 , P3_R1161_U79 );
nand NAND2_6856 ( P3_R1161_U458 , P3_U3080 , P3_R1161_U78 );
nand NAND2_6857 ( P3_R1161_U457 , P3_R1161_U328 , P3_R1161_U31 );
nand NAND2_6858 ( P3_R1161_U456 , P3_R1161_U182 , P3_R1161_U161 );
nand NAND2_6859 ( P3_R1161_U455 , P3_U3907 , P3_R1161_U90 );
nand NAND2_6860 ( P3_R1161_U454 , P3_U3075 , P3_R1161_U81 );
nand NAND2_6861 ( P3_R1161_U453 , P3_R1161_U452 , P3_R1161_U451 );
nand NAND2_6862 ( P3_R1161_U452 , P3_U3906 , P3_R1161_U55 );
nand NAND2_6863 ( P3_R1161_U451 , P3_U3074 , P3_R1161_U54 );
nand NAND2_6864 ( P3_R1161_U450 , P3_U3906 , P3_R1161_U55 );
nand NAND2_6865 ( P3_R1161_U449 , P3_U3074 , P3_R1161_U54 );
and AND2_6866 ( P3_U3013 , P3_U3380 , P3_U5450 );
and AND2_6867 ( P3_U3014 , P3_U3380 , P3_U3379 );
and AND2_6868 ( P3_U3015 , P3_U5453 , P3_U3379 );
and AND2_6869 ( P3_U3016 , P3_U5453 , P3_U5450 );
and AND2_6870 ( P3_U3017 , P3_U3874 , P3_U5447 );
and AND2_6871 ( P3_U3018 , P3_U3587 , P3_U3582 );
and AND2_6872 ( P3_U3019 , P3_U3381 , P3_U3382 );
and AND2_6873 ( P3_U3020 , P3_U5462 , P3_U3381 );
and AND2_6874 ( P3_U3021 , P3_U5459 , P3_U3382 );
and AND2_6875 ( P3_U3022 , P3_U5462 , P3_U5459 );
and AND2_6876 ( P3_U3023 , P3_U3046 , P3_STATE_REG );
and AND2_6877 ( P3_U3024 , P3_U3696 , P3_U3366 );
and AND2_6878 ( P3_U3025 , P3_U3911 , P3_U4073 );
and AND2_6879 ( P3_U3026 , P3_U3015 , P3_U5447 );
and AND2_6880 ( P3_U3027 , P3_U3297 , P3_STATE_REG );
and AND2_6881 ( P3_U3028 , P3_U3886 , P3_U3912 );
and AND2_6882 ( P3_U3029 , P3_U3912 , P3_U3365 );
and AND2_6883 ( P3_U3030 , P3_U3693 , P3_U3912 );
and AND2_6884 ( P3_U3031 , P3_U3890 , P3_U3023 );
and AND2_6885 ( P3_U3032 , P3_U3895 , P3_U4073 );
and AND2_6886 ( P3_U3033 , P3_U3911 , P3_U4089 );
and AND2_6887 ( P3_U3034 , P3_U3912 , P3_U3025 );
and AND2_6888 ( P3_U3035 , P3_U3023 , P3_U4989 );
and AND2_6889 ( P3_U3036 , P3_U3895 , P3_U4089 );
and AND2_6890 ( P3_U3037 , P3_U5468 , P3_U4754 );
and AND2_6891 ( P3_U3038 , P3_U3024 , P3_U5468 );
and AND2_6892 ( P3_U3039 , P3_U5465 , P3_U4754 );
and AND2_6893 ( P3_U3040 , P3_U3892 , P3_U4754 );
and AND2_6894 ( P3_U3041 , P3_U3024 , P3_U3892 );
and AND2_6895 ( P3_U3042 , P3_U3023 , P3_U3366 );
and AND2_6896 ( P3_U3043 , P3_U3023 , P3_U3365 );
and AND2_6897 ( P3_U3044 , P3_U5004 , P3_STATE_REG );
and AND2_6898 ( P3_U3045 , P3_U3023 , P3_U5006 );
and AND2_6899 ( P3_U3046 , P3_U5440 , P3_U3362 );
and AND2_6900 ( P3_U3047 , P3_U3692 , P3_U3018 );
and AND2_6901 ( P3_U3048 , P3_U3691 , P3_U3018 );
and AND2_6902 ( P3_U3049 , P3_U4749 , P3_U4748 );
and AND2_6903 ( P3_U3050 , P3_U4759 , P3_STATE_REG );
and AND2_6904 ( P3_U3051 , P3_U3897 , P3_U4761 );
nand NAND4_6905 ( P3_U3052 , P3_U4536 , P3_U4537 , P3_U4535 , P3_U4538 );
nand NAND4_6906 ( P3_U3053 , P3_U4556 , P3_U4555 , P3_U4554 , P3_U4553 );
nand NAND4_6907 ( P3_U3054 , P3_U4574 , P3_U4573 , P3_U4572 , P3_U4571 );
nand NAND4_6908 ( P3_U3055 , P3_U4612 , P3_U4611 , P3_U4610 , P3_U4609 );
nand NAND4_6909 ( P3_U3056 , P3_U4520 , P3_U4519 , P3_U4518 , P3_U4517 );
nand NAND4_6910 ( P3_U3057 , P3_U4502 , P3_U4501 , P3_U4500 , P3_U4499 );
nand NAND4_6911 ( P3_U3058 , P3_U4592 , P3_U4591 , P3_U4590 , P3_U4589 );
nand NAND4_6912 ( P3_U3059 , P3_U4124 , P3_U4123 , P3_U4122 , P3_U4121 );
nand NAND4_6913 ( P3_U3060 , P3_U4448 , P3_U4447 , P3_U4446 , P3_U4445 );
nand NAND4_6914 ( P3_U3061 , P3_U4232 , P3_U4231 , P3_U4230 , P3_U4229 );
nand NAND4_6915 ( P3_U3062 , P3_U4250 , P3_U4249 , P3_U4248 , P3_U4247 );
nand NAND4_6916 ( P3_U3063 , P3_U4106 , P3_U4105 , P3_U4104 , P3_U4103 );
nand NAND4_6917 ( P3_U3064 , P3_U4484 , P3_U4483 , P3_U4482 , P3_U4481 );
nand NAND4_6918 ( P3_U3065 , P3_U4466 , P3_U4465 , P3_U4464 , P3_U4463 );
nand NAND4_6919 ( P3_U3066 , P3_U4142 , P3_U4141 , P3_U4140 , P3_U4139 );
nand NAND4_6920 ( P3_U3067 , P3_U4081 , P3_U4080 , P3_U4079 , P3_U4078 );
nand NAND4_6921 ( P3_U3068 , P3_U4358 , P3_U4357 , P3_U4356 , P3_U4355 );
nand NAND4_6922 ( P3_U3069 , P3_U4178 , P3_U4177 , P3_U4176 , P3_U4175 );
nand NAND4_6923 ( P3_U3070 , P3_U4160 , P3_U4159 , P3_U4158 , P3_U4157 );
nand NAND4_6924 ( P3_U3071 , P3_U4268 , P3_U4267 , P3_U4266 , P3_U4265 );
nand NAND4_6925 ( P3_U3072 , P3_U4340 , P3_U4339 , P3_U4338 , P3_U4337 );
nand NAND4_6926 ( P3_U3073 , P3_U4322 , P3_U4321 , P3_U4320 , P3_U4319 );
nand NAND4_6927 ( P3_U3074 , P3_U4430 , P3_U4429 , P3_U4428 , P3_U4427 );
nand NAND4_6928 ( P3_U3075 , P3_U4412 , P3_U4411 , P3_U4410 , P3_U4409 );
nand NAND4_6929 ( P3_U3076 , P3_U4086 , P3_U4085 , P3_U4084 , P3_U4083 );
nand NAND4_6930 ( P3_U3077 , P3_U4062 , P3_U4061 , P3_U4060 , P3_U4059 );
nand NAND4_6931 ( P3_U3078 , P3_U4304 , P3_U4303 , P3_U4302 , P3_U4301 );
nand NAND4_6932 ( P3_U3079 , P3_U4286 , P3_U4285 , P3_U4284 , P3_U4283 );
nand NAND4_6933 ( P3_U3080 , P3_U4394 , P3_U4393 , P3_U4392 , P3_U4391 );
nand NAND4_6934 ( P3_U3081 , P3_U4376 , P3_U4375 , P3_U4374 , P3_U4373 );
nand NAND4_6935 ( P3_U3082 , P3_U4214 , P3_U4213 , P3_U4212 , P3_U4211 );
nand NAND4_6936 ( P3_U3083 , P3_U4196 , P3_U4195 , P3_U4194 , P3_U4193 );
nand NAND2_6937 ( P3_U3084 , P3_U5341 , P3_U5340 );
nand NAND2_6938 ( P3_U3085 , P3_U5343 , P3_U5342 );
nand NAND3_6939 ( P3_U3086 , P3_U5349 , P3_U5347 , P3_U5348 );
nand NAND3_6940 ( P3_U3087 , P3_U5352 , P3_U5350 , P3_U5351 );
nand NAND3_6941 ( P3_U3088 , P3_U5355 , P3_U5353 , P3_U5354 );
nand NAND3_6942 ( P3_U3089 , P3_U5358 , P3_U5356 , P3_U5357 );
nand NAND3_6943 ( P3_U3090 , P3_U5361 , P3_U5359 , P3_U5360 );
nand NAND3_6944 ( P3_U3091 , P3_U5364 , P3_U5362 , P3_U5363 );
nand NAND3_6945 ( P3_U3092 , P3_U5367 , P3_U5365 , P3_U5366 );
nand NAND3_6946 ( P3_U3093 , P3_U5370 , P3_U5368 , P3_U5369 );
nand NAND3_6947 ( P3_U3094 , P3_U5373 , P3_U5371 , P3_U5372 );
nand NAND3_6948 ( P3_U3095 , P3_U5376 , P3_U5374 , P3_U5375 );
nand NAND3_6949 ( P3_U3096 , P3_U5381 , P3_U5382 , P3_U5380 );
nand NAND3_6950 ( P3_U3097 , P3_U5384 , P3_U5385 , P3_U5383 );
nand NAND3_6951 ( P3_U3098 , P3_U5387 , P3_U5388 , P3_U5386 );
nand NAND3_6952 ( P3_U3099 , P3_U5390 , P3_U5391 , P3_U5389 );
nand NAND3_6953 ( P3_U3100 , P3_U5393 , P3_U5394 , P3_U5392 );
nand NAND3_6954 ( P3_U3101 , P3_U5396 , P3_U5397 , P3_U5395 );
nand NAND3_6955 ( P3_U3102 , P3_U5399 , P3_U5398 , P3_U5400 );
nand NAND3_6956 ( P3_U3103 , P3_U5402 , P3_U5401 , P3_U5403 );
nand NAND3_6957 ( P3_U3104 , P3_U5405 , P3_U5404 , P3_U5406 );
nand NAND3_6958 ( P3_U3105 , P3_U5408 , P3_U5407 , P3_U5409 );
nand NAND3_6959 ( P3_U3106 , P3_U5323 , P3_U5322 , P3_U5324 );
nand NAND3_6960 ( P3_U3107 , P3_U5326 , P3_U5325 , P3_U5327 );
nand NAND3_6961 ( P3_U3108 , P3_U5329 , P3_U5328 , P3_U5330 );
nand NAND3_6962 ( P3_U3109 , P3_U5332 , P3_U5331 , P3_U5333 );
nand NAND3_6963 ( P3_U3110 , P3_U5335 , P3_U5334 , P3_U5336 );
nand NAND3_6964 ( P3_U3111 , P3_U5338 , P3_U5337 , P3_U5339 );
nand NAND3_6965 ( P3_U3112 , P3_U5345 , P3_U5344 , P3_U5346 );
nand NAND3_6966 ( P3_U3113 , P3_U5378 , P3_U5377 , P3_U5379 );
nand NAND3_6967 ( P3_U3114 , P3_U5411 , P3_U5410 , P3_U5412 );
nand NAND2_6968 ( P3_U3115 , P3_U5414 , P3_U5413 );
nand NAND2_6969 ( P3_U3116 , P3_U5271 , P3_U5270 );
nand NAND2_6970 ( P3_U3117 , P3_U5273 , P3_U5272 );
nand NAND3_6971 ( P3_U3118 , P3_U5277 , P3_U3375 , P3_U5276 );
nand NAND3_6972 ( P3_U3119 , P3_U5279 , P3_U3375 , P3_U5278 );
nand NAND3_6973 ( P3_U3120 , P3_U5281 , P3_U3375 , P3_U5280 );
nand NAND3_6974 ( P3_U3121 , P3_U5283 , P3_U3375 , P3_U5282 );
nand NAND3_6975 ( P3_U3122 , P3_U5285 , P3_U3375 , P3_U5284 );
nand NAND3_6976 ( P3_U3123 , P3_U5287 , P3_U3375 , P3_U5286 );
nand NAND3_6977 ( P3_U3124 , P3_U5289 , P3_U3375 , P3_U5288 );
nand NAND3_6978 ( P3_U3125 , P3_U5291 , P3_U3375 , P3_U5290 );
nand NAND3_6979 ( P3_U3126 , P3_U5293 , P3_U3375 , P3_U5292 );
nand NAND3_6980 ( P3_U3127 , P3_U5295 , P3_U3375 , P3_U5294 );
nand NAND3_6981 ( P3_U3128 , P3_U5299 , P3_U3375 , P3_U5298 );
nand NAND3_6982 ( P3_U3129 , P3_U5301 , P3_U3375 , P3_U5300 );
nand NAND3_6983 ( P3_U3130 , P3_U5303 , P3_U3375 , P3_U5302 );
nand NAND3_6984 ( P3_U3131 , P3_U5305 , P3_U3375 , P3_U5304 );
nand NAND3_6985 ( P3_U3132 , P3_U5307 , P3_U3375 , P3_U5306 );
nand NAND3_6986 ( P3_U3133 , P3_U5309 , P3_U3375 , P3_U5308 );
nand NAND2_6987 ( P3_U3134 , P3_U3825 , P3_U5311 );
nand NAND2_6988 ( P3_U3135 , P3_U3826 , P3_U5313 );
nand NAND2_6989 ( P3_U3136 , P3_U3827 , P3_U5315 );
nand NAND2_6990 ( P3_U3137 , P3_U3828 , P3_U5317 );
nand NAND2_6991 ( P3_U3138 , P3_U3817 , P3_U5259 );
nand NAND2_6992 ( P3_U3139 , P3_U3818 , P3_U5261 );
nand NAND2_6993 ( P3_U3140 , P3_U3819 , P3_U5263 );
nand NAND2_6994 ( P3_U3141 , P3_U3820 , P3_U5265 );
nand NAND2_6995 ( P3_U3142 , P3_U3821 , P3_U5267 );
nand NAND2_6996 ( P3_U3143 , P3_U3822 , P3_U5269 );
nand NAND2_6997 ( P3_U3144 , P3_U3823 , P3_U5275 );
nand NAND2_6998 ( P3_U3145 , P3_U3824 , P3_U5297 );
nand NAND2_6999 ( P3_U3146 , P3_U3829 , P3_U5319 );
nand NAND2_7000 ( P3_U3147 , P3_U3830 , P3_U5321 );
nand NAND3_7001 ( P3_U3148 , P3_U3385 , P3_U5453 , P3_U3375 );
nand NAND2_7002 ( P3_U3149 , P3_U3813 , P3_U3013 );
nand NAND2_7003 ( P3_U3150 , P3_U3812 , P3_U5253 );
not NOT1_7004 ( P3_U3151 , P3_STATE_REG );
nand NAND3_7005 ( P3_U3152 , P3_U5944 , P3_U5943 , P3_U3359 );
nand NAND4_7006 ( P3_U3153 , P3_U5249 , P3_U5248 , P3_U3811 , P3_U5250 );
nand NAND4_7007 ( P3_U3154 , P3_U5240 , P3_U3810 , P3_U5239 , P3_U5241 );
nand NAND4_7008 ( P3_U3155 , P3_U5231 , P3_U5230 , P3_U3809 , P3_U5232 );
nand NAND4_7009 ( P3_U3156 , P3_U5222 , P3_U3808 , P3_U5221 , P3_U5223 );
nand NAND4_7010 ( P3_U3157 , P3_U5213 , P3_U5212 , P3_U3807 , P3_U5214 );
nand NAND3_7011 ( P3_U3158 , P3_U3805 , P3_U5204 , P3_U3806 );
nand NAND4_7012 ( P3_U3159 , P3_U5195 , P3_U3804 , P3_U5194 , P3_U5196 );
nand NAND4_7013 ( P3_U3160 , P3_U5186 , P3_U3803 , P3_U5185 , P3_U5187 );
nand NAND4_7014 ( P3_U3161 , P3_U5177 , P3_U5176 , P3_U3802 , P3_U5178 );
nand NAND3_7015 ( P3_U3162 , P3_U3800 , P3_U5168 , P3_U3801 );
nand NAND4_7016 ( P3_U3163 , P3_U5159 , P3_U3799 , P3_U5158 , P3_U5160 );
nand NAND4_7017 ( P3_U3164 , P3_U5150 , P3_U5149 , P3_U3798 , P3_U5151 );
nand NAND4_7018 ( P3_U3165 , P3_U5141 , P3_U3797 , P3_U5140 , P3_U5142 );
nand NAND4_7019 ( P3_U3166 , P3_U5132 , P3_U5131 , P3_U3796 , P3_U5133 );
nand NAND4_7020 ( P3_U3167 , P3_U5123 , P3_U5122 , P3_U3795 , P3_U5124 );
nand NAND4_7021 ( P3_U3168 , P3_U5114 , P3_U5113 , P3_U3794 , P3_U5115 );
nand NAND4_7022 ( P3_U3169 , P3_U5105 , P3_U3793 , P3_U5104 , P3_U5106 );
nand NAND3_7023 ( P3_U3170 , P3_U3791 , P3_U5096 , P3_U3792 );
nand NAND4_7024 ( P3_U3171 , P3_U5087 , P3_U5086 , P3_U3790 , P3_U5088 );
nand NAND2_7025 ( P3_U3172 , P3_U5079 , P3_U3789 );
nand NAND4_7026 ( P3_U3173 , P3_U5071 , P3_U3786 , P3_U5070 , P3_U5072 );
nand NAND4_7027 ( P3_U3174 , P3_U5062 , P3_U5061 , P3_U3785 , P3_U5063 );
nand NAND4_7028 ( P3_U3175 , P3_U5053 , P3_U3784 , P3_U5052 , P3_U5054 );
nand NAND4_7029 ( P3_U3176 , P3_U5044 , P3_U5043 , P3_U3783 , P3_U5045 );
nand NAND3_7030 ( P3_U3177 , P3_U3781 , P3_U5035 , P3_U3782 );
nand NAND4_7031 ( P3_U3178 , P3_U5026 , P3_U5025 , P3_U3780 , P3_U5027 );
nand NAND4_7032 ( P3_U3179 , P3_U5017 , P3_U5016 , P3_U3779 , P3_U5018 );
nand NAND4_7033 ( P3_U3180 , P3_U5008 , P3_U3778 , P3_U5007 , P3_U5009 );
nand NAND4_7034 ( P3_U3181 , P3_U4995 , P3_U4994 , P3_U3777 , P3_U4996 );
nand NAND2_7035 ( P3_U3182 , P3_U4973 , P3_U3756 );
nand NAND2_7036 ( P3_U3183 , P3_U4962 , P3_U3753 );
nand NAND2_7037 ( P3_U3184 , P3_U4951 , P3_U3750 );
nand NAND3_7038 ( P3_U3185 , P3_U4941 , P3_U4940 , P3_U3747 );
nand NAND3_7039 ( P3_U3186 , P3_U4930 , P3_U4929 , P3_U3744 );
nand NAND4_7040 ( P3_U3187 , P3_U4918 , P3_U3741 , P3_U3743 , P3_U4916 );
nand NAND3_7041 ( P3_U3188 , P3_U4907 , P3_U3738 , P3_U4905 );
nand NAND2_7042 ( P3_U3189 , P3_U4896 , P3_U3735 );
nand NAND2_7043 ( P3_U3190 , P3_U4885 , P3_U3732 );
nand NAND2_7044 ( P3_U3191 , P3_U4874 , P3_U3729 );
nand NAND2_7045 ( P3_U3192 , P3_U4863 , P3_U3726 );
nand NAND2_7046 ( P3_U3193 , P3_U4852 , P3_U3723 );
nand NAND2_7047 ( P3_U3194 , P3_U4841 , P3_U3720 );
nand NAND2_7048 ( P3_U3195 , P3_U4830 , P3_U3717 );
nand NAND2_7049 ( P3_U3196 , P3_U4819 , P3_U3714 );
nand NAND2_7050 ( P3_U3197 , P3_U4808 , P3_U3711 );
nand NAND2_7051 ( P3_U3198 , P3_U4797 , P3_U3708 );
nand NAND2_7052 ( P3_U3199 , P3_U4786 , P3_U3705 );
nand NAND2_7053 ( P3_U3200 , P3_U4775 , P3_U3702 );
nand NAND2_7054 ( P3_U3201 , P3_U4764 , P3_U3699 );
nand NAND3_7055 ( P3_U3202 , P3_U4753 , P3_U3049 , P3_U4752 );
nand NAND3_7056 ( P3_U3203 , P3_U4751 , P3_U3049 , P3_U4750 );
nand NAND4_7057 ( P3_U3204 , P3_U4746 , P3_U4747 , P3_U4745 , P3_U3866 );
nand NAND5_7058 ( P3_U3205 , P3_U4743 , P3_U4741 , P3_U4744 , P3_U4742 , P3_U3865 );
nand NAND5_7059 ( P3_U3206 , P3_U4739 , P3_U4737 , P3_U4740 , P3_U4738 , P3_U3864 );
nand NAND5_7060 ( P3_U3207 , P3_U4735 , P3_U4733 , P3_U4736 , P3_U4734 , P3_U3863 );
nand NAND5_7061 ( P3_U3208 , P3_U4731 , P3_U4729 , P3_U4732 , P3_U4730 , P3_U3862 );
nand NAND5_7062 ( P3_U3209 , P3_U4727 , P3_U4725 , P3_U4728 , P3_U4726 , P3_U3861 );
nand NAND5_7063 ( P3_U3210 , P3_U4723 , P3_U4721 , P3_U4724 , P3_U4722 , P3_U3860 );
nand NAND5_7064 ( P3_U3211 , P3_U4719 , P3_U4717 , P3_U4720 , P3_U4718 , P3_U3859 );
nand NAND5_7065 ( P3_U3212 , P3_U4715 , P3_U4713 , P3_U4716 , P3_U4714 , P3_U3858 );
nand NAND5_7066 ( P3_U3213 , P3_U4711 , P3_U4709 , P3_U4712 , P3_U4710 , P3_U3857 );
nand NAND5_7067 ( P3_U3214 , P3_U4707 , P3_U4705 , P3_U4708 , P3_U4706 , P3_U3856 );
nand NAND5_7068 ( P3_U3215 , P3_U4703 , P3_U4701 , P3_U4704 , P3_U4702 , P3_U3855 );
nand NAND5_7069 ( P3_U3216 , P3_U4699 , P3_U4697 , P3_U4700 , P3_U4698 , P3_U3854 );
nand NAND5_7070 ( P3_U3217 , P3_U4695 , P3_U4693 , P3_U4696 , P3_U4694 , P3_U3853 );
nand NAND5_7071 ( P3_U3218 , P3_U4691 , P3_U4689 , P3_U4692 , P3_U4690 , P3_U3852 );
nand NAND5_7072 ( P3_U3219 , P3_U4687 , P3_U4685 , P3_U4688 , P3_U4686 , P3_U3851 );
nand NAND5_7073 ( P3_U3220 , P3_U4684 , P3_U4682 , P3_U4683 , P3_U4681 , P3_U3850 );
nand NAND5_7074 ( P3_U3221 , P3_U4680 , P3_U4679 , P3_U4678 , P3_U4677 , P3_U3849 );
nand NAND5_7075 ( P3_U3222 , P3_U4676 , P3_U4674 , P3_U4675 , P3_U4673 , P3_U3848 );
nand NAND5_7076 ( P3_U3223 , P3_U4672 , P3_U4671 , P3_U4670 , P3_U4669 , P3_U3847 );
nand NAND5_7077 ( P3_U3224 , P3_U4666 , P3_U4665 , P3_U4667 , P3_U3846 , P3_U4668 );
nand NAND5_7078 ( P3_U3225 , P3_U4662 , P3_U4661 , P3_U4663 , P3_U3845 , P3_U4664 );
nand NAND5_7079 ( P3_U3226 , P3_U4658 , P3_U4657 , P3_U4659 , P3_U3844 , P3_U4660 );
nand NAND5_7080 ( P3_U3227 , P3_U4654 , P3_U4653 , P3_U4655 , P3_U3843 , P3_U4656 );
nand NAND5_7081 ( P3_U3228 , P3_U4650 , P3_U4649 , P3_U4651 , P3_U3842 , P3_U4652 );
nand NAND5_7082 ( P3_U3229 , P3_U4646 , P3_U4645 , P3_U4647 , P3_U3841 , P3_U4648 );
nand NAND5_7083 ( P3_U3230 , P3_U4642 , P3_U4641 , P3_U4643 , P3_U3840 , P3_U4644 );
nand NAND5_7084 ( P3_U3231 , P3_U4638 , P3_U4637 , P3_U4639 , P3_U3839 , P3_U4640 );
nand NAND5_7085 ( P3_U3232 , P3_U4634 , P3_U4633 , P3_U4635 , P3_U3838 , P3_U4636 );
nand NAND5_7086 ( P3_U3233 , P3_U4630 , P3_U4629 , P3_U4631 , P3_U3837 , P3_U4632 );
and AND2_7087 ( P3_U3234 , P3_D_REG_31_ , P3_U3832 );
and AND2_7088 ( P3_U3235 , P3_D_REG_30_ , P3_U3832 );
and AND2_7089 ( P3_U3236 , P3_D_REG_29_ , P3_U3832 );
and AND2_7090 ( P3_U3237 , P3_D_REG_28_ , P3_U3832 );
and AND2_7091 ( P3_U3238 , P3_D_REG_27_ , P3_U3832 );
and AND2_7092 ( P3_U3239 , P3_D_REG_26_ , P3_U3832 );
and AND2_7093 ( P3_U3240 , P3_D_REG_25_ , P3_U3832 );
and AND2_7094 ( P3_U3241 , P3_D_REG_24_ , P3_U3832 );
and AND2_7095 ( P3_U3242 , P3_D_REG_23_ , P3_U3832 );
and AND2_7096 ( P3_U3243 , P3_D_REG_22_ , P3_U3832 );
and AND2_7097 ( P3_U3244 , P3_D_REG_21_ , P3_U3832 );
and AND2_7098 ( P3_U3245 , P3_D_REG_20_ , P3_U3832 );
and AND2_7099 ( P3_U3246 , P3_D_REG_19_ , P3_U3832 );
and AND2_7100 ( P3_U3247 , P3_D_REG_18_ , P3_U3832 );
and AND2_7101 ( P3_U3248 , P3_D_REG_17_ , P3_U3832 );
and AND2_7102 ( P3_U3249 , P3_D_REG_16_ , P3_U3832 );
and AND2_7103 ( P3_U3250 , P3_D_REG_15_ , P3_U3832 );
and AND2_7104 ( P3_U3251 , P3_D_REG_14_ , P3_U3832 );
and AND2_7105 ( P3_U3252 , P3_D_REG_13_ , P3_U3832 );
and AND2_7106 ( P3_U3253 , P3_D_REG_12_ , P3_U3832 );
and AND2_7107 ( P3_U3254 , P3_D_REG_11_ , P3_U3832 );
and AND2_7108 ( P3_U3255 , P3_D_REG_10_ , P3_U3832 );
and AND2_7109 ( P3_U3256 , P3_D_REG_9_ , P3_U3832 );
and AND2_7110 ( P3_U3257 , P3_D_REG_8_ , P3_U3832 );
and AND2_7111 ( P3_U3258 , P3_D_REG_7_ , P3_U3832 );
and AND2_7112 ( P3_U3259 , P3_D_REG_6_ , P3_U3832 );
and AND2_7113 ( P3_U3260 , P3_D_REG_5_ , P3_U3832 );
and AND2_7114 ( P3_U3261 , P3_D_REG_4_ , P3_U3832 );
and AND2_7115 ( P3_U3262 , P3_D_REG_3_ , P3_U3832 );
and AND2_7116 ( P3_U3263 , P3_D_REG_2_ , P3_U3832 );
nand NAND3_7117 ( P3_U3264 , P3_U4016 , P3_U4017 , P3_U4015 );
nand NAND3_7118 ( P3_U3265 , P3_U4013 , P3_U4014 , P3_U4012 );
nand NAND3_7119 ( P3_U3266 , P3_U4010 , P3_U4011 , P3_U4009 );
nand NAND3_7120 ( P3_U3267 , P3_U4007 , P3_U4008 , P3_U4006 );
nand NAND3_7121 ( P3_U3268 , P3_U4004 , P3_U4005 , P3_U4003 );
nand NAND3_7122 ( P3_U3269 , P3_U4001 , P3_U4002 , P3_U4000 );
nand NAND3_7123 ( P3_U3270 , P3_U3998 , P3_U3999 , P3_U3997 );
nand NAND3_7124 ( P3_U3271 , P3_U3995 , P3_U3996 , P3_U3994 );
nand NAND3_7125 ( P3_U3272 , P3_U3992 , P3_U3993 , P3_U3991 );
nand NAND3_7126 ( P3_U3273 , P3_U3989 , P3_U3990 , P3_U3988 );
nand NAND3_7127 ( P3_U3274 , P3_U3986 , P3_U3987 , P3_U3985 );
nand NAND3_7128 ( P3_U3275 , P3_U3983 , P3_U3984 , P3_U3982 );
nand NAND3_7129 ( P3_U3276 , P3_U3980 , P3_U3981 , P3_U3979 );
nand NAND3_7130 ( P3_U3277 , P3_U3977 , P3_U3978 , P3_U3976 );
nand NAND3_7131 ( P3_U3278 , P3_U3974 , P3_U3975 , P3_U3973 );
nand NAND3_7132 ( P3_U3279 , P3_U3971 , P3_U3972 , P3_U3970 );
nand NAND3_7133 ( P3_U3280 , P3_U3968 , P3_U3969 , P3_U3967 );
nand NAND3_7134 ( P3_U3281 , P3_U3965 , P3_U3966 , P3_U3964 );
nand NAND3_7135 ( P3_U3282 , P3_U3962 , P3_U3963 , P3_U3961 );
nand NAND3_7136 ( P3_U3283 , P3_U3959 , P3_U3960 , P3_U3958 );
nand NAND3_7137 ( P3_U3284 , P3_U3956 , P3_U3957 , P3_U3955 );
nand NAND3_7138 ( P3_U3285 , P3_U3953 , P3_U3954 , P3_U3952 );
nand NAND3_7139 ( P3_U3286 , P3_U3950 , P3_U3951 , P3_U3949 );
nand NAND3_7140 ( P3_U3287 , P3_U3947 , P3_U3948 , P3_U3946 );
nand NAND3_7141 ( P3_U3288 , P3_U3944 , P3_U3945 , P3_U3943 );
nand NAND3_7142 ( P3_U3289 , P3_U3941 , P3_U3942 , P3_U3940 );
nand NAND3_7143 ( P3_U3290 , P3_U3938 , P3_U3939 , P3_U3937 );
nand NAND3_7144 ( P3_U3291 , P3_U3935 , P3_U3936 , P3_U3934 );
nand NAND3_7145 ( P3_U3292 , P3_U3932 , P3_U3933 , P3_U3931 );
nand NAND3_7146 ( P3_U3293 , P3_U3929 , P3_U3930 , P3_U3928 );
nand NAND3_7147 ( P3_U3294 , P3_U3926 , P3_U3927 , P3_U3925 );
nand NAND3_7148 ( P3_U3295 , P3_U3923 , P3_U3924 , P3_U3922 );
and AND2_7149 ( P3_U3296 , P3_U3775 , P3_U5421 );
nand NAND2_7150 ( P3_U3297 , P3_STATE_REG , P3_U3831 );
not NOT1_7151 ( P3_U3298 , P3_B_REG );
nand NAND2_7152 ( P3_U3299 , P3_U3374 , P3_U5431 );
nand NAND2_7153 ( P3_U3300 , P3_U3374 , P3_U4018 );
nand NAND2_7154 ( P3_U3301 , P3_U3013 , P3_U5447 );
nand NAND2_7155 ( P3_U3302 , P3_U3014 , P3_U5456 );
nand NAND2_7156 ( P3_U3303 , P3_U3588 , P3_U3018 );
nand NAND2_7157 ( P3_U3304 , P3_U3589 , P3_U3018 );
nand NAND2_7158 ( P3_U3305 , P3_U3014 , P3_U5447 );
nand NAND2_7159 ( P3_U3306 , P3_U3014 , P3_U3378 );
nand NAND2_7160 ( P3_U3307 , P3_U3013 , P3_U3378 );
nand NAND3_7161 ( P3_U3308 , P3_U3385 , P3_U3379 , P3_U3378 );
nand NAND3_7162 ( P3_U3309 , P3_U5450 , P3_U3385 , P3_U3378 );
nand NAND2_7163 ( P3_U3310 , P3_U5456 , P3_U3013 );
nand NAND2_7164 ( P3_U3311 , P3_U3878 , P3_U5447 );
nand NAND2_7165 ( P3_U3312 , P3_U3016 , P3_U3385 );
nand NAND2_7166 ( P3_U3313 , P3_U3385 , P3_U3380 );
nand NAND5_7167 ( P3_U3314 , P3_U4070 , P3_U4069 , P3_U4071 , P3_U3576 , P3_U3575 );
nand NAND4_7168 ( P3_U3315 , P3_U4091 , P3_U4090 , P3_U3590 , P3_U3592 );
nand NAND4_7169 ( P3_U3316 , P3_U4109 , P3_U4108 , P3_U3594 , P3_U3596 );
nand NAND4_7170 ( P3_U3317 , P3_U4127 , P3_U4126 , P3_U3598 , P3_U3600 );
nand NAND5_7171 ( P3_U3318 , P3_U4145 , P3_U4144 , P3_U4146 , P3_U4147 , P3_U3603 );
nand NAND5_7172 ( P3_U3319 , P3_U4163 , P3_U4162 , P3_U4164 , P3_U4165 , P3_U3606 );
nand NAND5_7173 ( P3_U3320 , P3_U4181 , P3_U4180 , P3_U4182 , P3_U4183 , P3_U3609 );
nand NAND5_7174 ( P3_U3321 , P3_U4199 , P3_U4198 , P3_U4200 , P3_U4201 , P3_U3612 );
nand NAND5_7175 ( P3_U3322 , P3_U4217 , P3_U4216 , P3_U4218 , P3_U4219 , P3_U3615 );
nand NAND4_7176 ( P3_U3323 , P3_U4235 , P3_U4234 , P3_U3617 , P3_U3619 );
nand NAND4_7177 ( P3_U3324 , P3_U4253 , P3_U4252 , P3_U3621 , P3_U3623 );
nand NAND5_7178 ( P3_U3325 , P3_U4271 , P3_U4270 , P3_U4272 , P3_U4273 , P3_U3626 );
nand NAND4_7179 ( P3_U3326 , P3_U4289 , P3_U4288 , P3_U3628 , P3_U3630 );
nand NAND4_7180 ( P3_U3327 , P3_U4307 , P3_U4306 , P3_U3632 , P3_U3634 );
nand NAND5_7181 ( P3_U3328 , P3_U4325 , P3_U4324 , P3_U4326 , P3_U4327 , P3_U3637 );
nand NAND5_7182 ( P3_U3329 , P3_U4343 , P3_U4342 , P3_U4344 , P3_U4345 , P3_U3640 );
nand NAND5_7183 ( P3_U3330 , P3_U4361 , P3_U4360 , P3_U4362 , P3_U4363 , P3_U3643 );
nand NAND4_7184 ( P3_U3331 , P3_U4379 , P3_U4378 , P3_U3645 , P3_U3647 );
nand NAND5_7185 ( P3_U3332 , P3_U4397 , P3_U4396 , P3_U4398 , P3_U4399 , P3_U3650 );
nand NAND5_7186 ( P3_U3333 , P3_U4415 , P3_U4414 , P3_U4416 , P3_U4417 , P3_U3653 );
nand NAND2_7187 ( P3_U3334 , U49 , P3_U3833 );
nand NAND5_7188 ( P3_U3335 , P3_U4433 , P3_U4432 , P3_U4434 , P3_U4435 , P3_U3656 );
nand NAND2_7189 ( P3_U3336 , U48 , P3_U3833 );
nand NAND5_7190 ( P3_U3337 , P3_U4451 , P3_U4450 , P3_U4452 , P3_U4453 , P3_U3659 );
nand NAND2_7191 ( P3_U3338 , U47 , P3_U3833 );
nand NAND5_7192 ( P3_U3339 , P3_U4469 , P3_U4468 , P3_U4470 , P3_U4471 , P3_U3662 );
nand NAND2_7193 ( P3_U3340 , U46 , P3_U3833 );
nand NAND5_7194 ( P3_U3341 , P3_U4487 , P3_U4486 , P3_U4488 , P3_U4489 , P3_U3665 );
nand NAND2_7195 ( P3_U3342 , U45 , P3_U3833 );
nand NAND4_7196 ( P3_U3343 , P3_U4505 , P3_U4504 , P3_U3667 , P3_U3669 );
nand NAND2_7197 ( P3_U3344 , U44 , P3_U3833 );
nand NAND4_7198 ( P3_U3345 , P3_U4523 , P3_U4522 , P3_U3671 , P3_U3673 );
nand NAND2_7199 ( P3_U3346 , U43 , P3_U3833 );
nand NAND4_7200 ( P3_U3347 , P3_U4541 , P3_U4540 , P3_U3675 , P3_U3677 );
nand NAND2_7201 ( P3_U3348 , U42 , P3_U3833 );
nand NAND4_7202 ( P3_U3349 , P3_U4559 , P3_U4558 , P3_U3679 , P3_U3681 );
nand NAND2_7203 ( P3_U3350 , U41 , P3_U3833 );
nand NAND4_7204 ( P3_U3351 , P3_U4577 , P3_U4576 , P3_U3683 , P3_U3685 );
nand NAND2_7205 ( P3_U3352 , P3_U3383 , P3_U3384 );
nand NAND2_7206 ( P3_U3353 , U40 , P3_U3833 );
nand NAND5_7207 ( P3_U3354 , P3_U4597 , P3_U4596 , P3_U4598 , P3_U3687 , P3_U3689 );
nand NAND2_7208 ( P3_U3355 , U38 , P3_U3833 );
nand NAND2_7209 ( P3_U3356 , U37 , P3_U3833 );
nand NAND2_7210 ( P3_U3357 , P3_U3015 , P3_U5456 );
nand NAND2_7211 ( P3_U3358 , P3_U3023 , P3_U4627 );
nand NAND2_7212 ( P3_U3359 , P3_U5447 , P3_U3385 );
nand NAND2_7213 ( P3_U3360 , P3_U3879 , P3_U5447 );
nand NAND3_7214 ( P3_U3361 , P3_U3911 , P3_U4595 , P3_U3055 );
nand NAND3_7215 ( P3_U3362 , P3_U3373 , P3_U3374 , P3_U3372 );
nand NAND2_7216 ( P3_U3363 , P3_U3694 , P3_U3910 );
nand NAND2_7217 ( P3_U3364 , P3_U3313 , P3_U3833 );
nand NAND2_7218 ( P3_U3365 , P3_U3877 , P3_U5423 );
nand NAND2_7219 ( P3_U3366 , P3_U3695 , P3_U3050 );
nand NAND2_7220 ( P3_U3367 , P3_U3882 , P3_U3385 );
nand NAND2_7221 ( P3_U3368 , P3_U3759 , P3_U3890 );
nand NAND2_7222 ( P3_U3369 , P3_U3876 , P3_U3378 );
nand NAND3_7223 ( P3_U3370 , P3_U4992 , P3_U4991 , P3_U3776 );
nand NAND2_7224 ( P3_U3371 , P3_U5417 , P3_U3917 );
nand NAND2_7225 ( P3_U3372 , P3_U5427 , P3_U5426 );
nand NAND2_7226 ( P3_U3373 , P3_U5430 , P3_U5429 );
nand NAND2_7227 ( P3_U3374 , P3_U5433 , P3_U5432 );
nand NAND2_7228 ( P3_U3375 , P3_U5439 , P3_U5438 );
nand NAND2_7229 ( P3_U3376 , P3_U5442 , P3_U5441 );
nand NAND2_7230 ( P3_U3377 , P3_U5444 , P3_U5443 );
nand NAND2_7231 ( P3_U3378 , P3_U5446 , P3_U5445 );
nand NAND2_7232 ( P3_U3379 , P3_U5449 , P3_U5448 );
nand NAND2_7233 ( P3_U3380 , P3_U5452 , P3_U5451 );
nand NAND2_7234 ( P3_U3381 , P3_U5458 , P3_U5457 );
nand NAND2_7235 ( P3_U3382 , P3_U5461 , P3_U5460 );
nand NAND2_7236 ( P3_U3383 , P3_U5464 , P3_U5463 );
nand NAND2_7237 ( P3_U3384 , P3_U5467 , P3_U5466 );
nand NAND2_7238 ( P3_U3385 , P3_U5455 , P3_U5454 );
nand NAND2_7239 ( P3_U3386 , P3_U5470 , P3_U5469 );
nand NAND2_7240 ( P3_U3387 , P3_U5472 , P3_U5471 );
nand NAND2_7241 ( P3_U3388 , P3_U5475 , P3_U5474 );
nand NAND2_7242 ( P3_U3389 , P3_U5478 , P3_U5477 );
nand NAND2_7243 ( P3_U3390 , P3_U5484 , P3_U5483 );
nand NAND2_7244 ( P3_U3391 , P3_U5486 , P3_U5485 );
nand NAND2_7245 ( P3_U3392 , P3_U5488 , P3_U5487 );
nand NAND2_7246 ( P3_U3393 , P3_U5491 , P3_U5490 );
nand NAND2_7247 ( P3_U3394 , P3_U5493 , P3_U5492 );
nand NAND2_7248 ( P3_U3395 , P3_U5495 , P3_U5494 );
nand NAND2_7249 ( P3_U3396 , P3_U5498 , P3_U5497 );
nand NAND2_7250 ( P3_U3397 , P3_U5500 , P3_U5499 );
nand NAND2_7251 ( P3_U3398 , P3_U5502 , P3_U5501 );
nand NAND2_7252 ( P3_U3399 , P3_U5505 , P3_U5504 );
nand NAND2_7253 ( P3_U3400 , P3_U5507 , P3_U5506 );
nand NAND2_7254 ( P3_U3401 , P3_U5509 , P3_U5508 );
nand NAND2_7255 ( P3_U3402 , P3_U5512 , P3_U5511 );
nand NAND2_7256 ( P3_U3403 , P3_U5514 , P3_U5513 );
nand NAND2_7257 ( P3_U3404 , P3_U5516 , P3_U5515 );
nand NAND2_7258 ( P3_U3405 , P3_U5519 , P3_U5518 );
nand NAND2_7259 ( P3_U3406 , P3_U5521 , P3_U5520 );
nand NAND2_7260 ( P3_U3407 , P3_U5523 , P3_U5522 );
nand NAND2_7261 ( P3_U3408 , P3_U5526 , P3_U5525 );
nand NAND2_7262 ( P3_U3409 , P3_U5528 , P3_U5527 );
nand NAND2_7263 ( P3_U3410 , P3_U5530 , P3_U5529 );
nand NAND2_7264 ( P3_U3411 , P3_U5533 , P3_U5532 );
nand NAND2_7265 ( P3_U3412 , P3_U5535 , P3_U5534 );
nand NAND2_7266 ( P3_U3413 , P3_U5537 , P3_U5536 );
nand NAND2_7267 ( P3_U3414 , P3_U5540 , P3_U5539 );
nand NAND2_7268 ( P3_U3415 , P3_U5542 , P3_U5541 );
nand NAND2_7269 ( P3_U3416 , P3_U5544 , P3_U5543 );
nand NAND2_7270 ( P3_U3417 , P3_U5547 , P3_U5546 );
nand NAND2_7271 ( P3_U3418 , P3_U5549 , P3_U5548 );
nand NAND2_7272 ( P3_U3419 , P3_U5551 , P3_U5550 );
nand NAND2_7273 ( P3_U3420 , P3_U5554 , P3_U5553 );
nand NAND2_7274 ( P3_U3421 , P3_U5556 , P3_U5555 );
nand NAND2_7275 ( P3_U3422 , P3_U5558 , P3_U5557 );
nand NAND2_7276 ( P3_U3423 , P3_U5561 , P3_U5560 );
nand NAND2_7277 ( P3_U3424 , P3_U5563 , P3_U5562 );
nand NAND2_7278 ( P3_U3425 , P3_U5565 , P3_U5564 );
nand NAND2_7279 ( P3_U3426 , P3_U5568 , P3_U5567 );
nand NAND2_7280 ( P3_U3427 , P3_U5570 , P3_U5569 );
nand NAND2_7281 ( P3_U3428 , P3_U5572 , P3_U5571 );
nand NAND2_7282 ( P3_U3429 , P3_U5575 , P3_U5574 );
nand NAND2_7283 ( P3_U3430 , P3_U5577 , P3_U5576 );
nand NAND2_7284 ( P3_U3431 , P3_U5579 , P3_U5578 );
nand NAND2_7285 ( P3_U3432 , P3_U5582 , P3_U5581 );
nand NAND2_7286 ( P3_U3433 , P3_U5584 , P3_U5583 );
nand NAND2_7287 ( P3_U3434 , P3_U5586 , P3_U5585 );
nand NAND2_7288 ( P3_U3435 , P3_U5589 , P3_U5588 );
nand NAND2_7289 ( P3_U3436 , P3_U5591 , P3_U5590 );
nand NAND2_7290 ( P3_U3437 , P3_U5593 , P3_U5592 );
nand NAND2_7291 ( P3_U3438 , P3_U5596 , P3_U5595 );
nand NAND2_7292 ( P3_U3439 , P3_U5598 , P3_U5597 );
nand NAND2_7293 ( P3_U3440 , P3_U5600 , P3_U5599 );
nand NAND2_7294 ( P3_U3441 , P3_U5603 , P3_U5602 );
nand NAND2_7295 ( P3_U3442 , P3_U5605 , P3_U5604 );
nand NAND2_7296 ( P3_U3443 , P3_U5607 , P3_U5606 );
nand NAND2_7297 ( P3_U3444 , P3_U5610 , P3_U5609 );
nand NAND2_7298 ( P3_U3445 , P3_U5612 , P3_U5611 );
nand NAND2_7299 ( P3_U3446 , P3_U5615 , P3_U5614 );
nand NAND2_7300 ( P3_U3447 , P3_U5617 , P3_U5616 );
nand NAND2_7301 ( P3_U3448 , P3_U5619 , P3_U5618 );
nand NAND2_7302 ( P3_U3449 , P3_U5621 , P3_U5620 );
nand NAND2_7303 ( P3_U3450 , P3_U5623 , P3_U5622 );
nand NAND2_7304 ( P3_U3451 , P3_U5625 , P3_U5624 );
nand NAND2_7305 ( P3_U3452 , P3_U5627 , P3_U5626 );
nand NAND2_7306 ( P3_U3453 , P3_U5629 , P3_U5628 );
nand NAND2_7307 ( P3_U3454 , P3_U5631 , P3_U5630 );
nand NAND2_7308 ( P3_U3455 , P3_U5633 , P3_U5632 );
nand NAND2_7309 ( P3_U3456 , P3_U5635 , P3_U5634 );
nand NAND2_7310 ( P3_U3457 , P3_U5637 , P3_U5636 );
nand NAND2_7311 ( P3_U3458 , P3_U5639 , P3_U5638 );
nand NAND2_7312 ( P3_U3459 , P3_U5643 , P3_U5642 );
nand NAND2_7313 ( P3_U3460 , P3_U5645 , P3_U5644 );
nand NAND2_7314 ( P3_U3461 , P3_U5647 , P3_U5646 );
nand NAND2_7315 ( P3_U3462 , P3_U5649 , P3_U5648 );
nand NAND2_7316 ( P3_U3463 , P3_U5651 , P3_U5650 );
nand NAND2_7317 ( P3_U3464 , P3_U5653 , P3_U5652 );
nand NAND2_7318 ( P3_U3465 , P3_U5655 , P3_U5654 );
nand NAND2_7319 ( P3_U3466 , P3_U5657 , P3_U5656 );
nand NAND2_7320 ( P3_U3467 , P3_U5659 , P3_U5658 );
nand NAND2_7321 ( P3_U3468 , P3_U5661 , P3_U5660 );
nand NAND2_7322 ( P3_U3469 , P3_U5663 , P3_U5662 );
nand NAND2_7323 ( P3_U3470 , P3_U5665 , P3_U5664 );
nand NAND2_7324 ( P3_U3471 , P3_U5667 , P3_U5666 );
nand NAND2_7325 ( P3_U3472 , P3_U5669 , P3_U5668 );
nand NAND2_7326 ( P3_U3473 , P3_U5671 , P3_U5670 );
nand NAND2_7327 ( P3_U3474 , P3_U5673 , P3_U5672 );
nand NAND2_7328 ( P3_U3475 , P3_U5675 , P3_U5674 );
nand NAND2_7329 ( P3_U3476 , P3_U5677 , P3_U5676 );
nand NAND2_7330 ( P3_U3477 , P3_U5679 , P3_U5678 );
nand NAND2_7331 ( P3_U3478 , P3_U5681 , P3_U5680 );
nand NAND2_7332 ( P3_U3479 , P3_U5683 , P3_U5682 );
nand NAND2_7333 ( P3_U3480 , P3_U5685 , P3_U5684 );
nand NAND2_7334 ( P3_U3481 , P3_U5687 , P3_U5686 );
nand NAND2_7335 ( P3_U3482 , P3_U5689 , P3_U5688 );
nand NAND2_7336 ( P3_U3483 , P3_U5691 , P3_U5690 );
nand NAND2_7337 ( P3_U3484 , P3_U5693 , P3_U5692 );
nand NAND2_7338 ( P3_U3485 , P3_U5695 , P3_U5694 );
nand NAND2_7339 ( P3_U3486 , P3_U5697 , P3_U5696 );
nand NAND2_7340 ( P3_U3487 , P3_U5699 , P3_U5698 );
nand NAND2_7341 ( P3_U3488 , P3_U5701 , P3_U5700 );
nand NAND2_7342 ( P3_U3489 , P3_U5703 , P3_U5702 );
nand NAND2_7343 ( P3_U3490 , P3_U5705 , P3_U5704 );
nand NAND2_7344 ( P3_U3491 , P3_U5770 , P3_U5769 );
nand NAND2_7345 ( P3_U3492 , P3_U5772 , P3_U5771 );
nand NAND2_7346 ( P3_U3493 , P3_U5774 , P3_U5773 );
nand NAND2_7347 ( P3_U3494 , P3_U5776 , P3_U5775 );
nand NAND2_7348 ( P3_U3495 , P3_U5778 , P3_U5777 );
nand NAND2_7349 ( P3_U3496 , P3_U5780 , P3_U5779 );
nand NAND2_7350 ( P3_U3497 , P3_U5782 , P3_U5781 );
nand NAND2_7351 ( P3_U3498 , P3_U5784 , P3_U5783 );
nand NAND2_7352 ( P3_U3499 , P3_U5786 , P3_U5785 );
nand NAND2_7353 ( P3_U3500 , P3_U5788 , P3_U5787 );
nand NAND2_7354 ( P3_U3501 , P3_U5790 , P3_U5789 );
nand NAND2_7355 ( P3_U3502 , P3_U5792 , P3_U5791 );
nand NAND2_7356 ( P3_U3503 , P3_U5794 , P3_U5793 );
nand NAND2_7357 ( P3_U3504 , P3_U5796 , P3_U5795 );
nand NAND2_7358 ( P3_U3505 , P3_U5798 , P3_U5797 );
nand NAND2_7359 ( P3_U3506 , P3_U5800 , P3_U5799 );
nand NAND2_7360 ( P3_U3507 , P3_U5802 , P3_U5801 );
nand NAND2_7361 ( P3_U3508 , P3_U5804 , P3_U5803 );
nand NAND2_7362 ( P3_U3509 , P3_U5806 , P3_U5805 );
nand NAND2_7363 ( P3_U3510 , P3_U5808 , P3_U5807 );
nand NAND2_7364 ( P3_U3511 , P3_U5810 , P3_U5809 );
nand NAND2_7365 ( P3_U3512 , P3_U5812 , P3_U5811 );
nand NAND2_7366 ( P3_U3513 , P3_U5814 , P3_U5813 );
nand NAND2_7367 ( P3_U3514 , P3_U5816 , P3_U5815 );
nand NAND2_7368 ( P3_U3515 , P3_U5818 , P3_U5817 );
nand NAND2_7369 ( P3_U3516 , P3_U5820 , P3_U5819 );
nand NAND2_7370 ( P3_U3517 , P3_U5822 , P3_U5821 );
nand NAND2_7371 ( P3_U3518 , P3_U5824 , P3_U5823 );
nand NAND2_7372 ( P3_U3519 , P3_U5826 , P3_U5825 );
nand NAND2_7373 ( P3_U3520 , P3_U5828 , P3_U5827 );
nand NAND2_7374 ( P3_U3521 , P3_U5830 , P3_U5829 );
nand NAND2_7375 ( P3_U3522 , P3_U5832 , P3_U5831 );
nand NAND2_7376 ( P3_U3523 , P3_U5946 , P3_U5945 );
nand NAND2_7377 ( P3_U3524 , P3_U5948 , P3_U5947 );
nand NAND2_7378 ( P3_U3525 , P3_U5950 , P3_U5949 );
nand NAND2_7379 ( P3_U3526 , P3_U5952 , P3_U5951 );
nand NAND2_7380 ( P3_U3527 , P3_U5954 , P3_U5953 );
nand NAND2_7381 ( P3_U3528 , P3_U5956 , P3_U5955 );
nand NAND2_7382 ( P3_U3529 , P3_U5958 , P3_U5957 );
nand NAND2_7383 ( P3_U3530 , P3_U5960 , P3_U5959 );
nand NAND2_7384 ( P3_U3531 , P3_U5962 , P3_U5961 );
nand NAND2_7385 ( P3_U3532 , P3_U5964 , P3_U5963 );
nand NAND2_7386 ( P3_U3533 , P3_U5966 , P3_U5965 );
nand NAND2_7387 ( P3_U3534 , P3_U5968 , P3_U5967 );
nand NAND2_7388 ( P3_U3535 , P3_U5970 , P3_U5969 );
nand NAND2_7389 ( P3_U3536 , P3_U5972 , P3_U5971 );
nand NAND2_7390 ( P3_U3537 , P3_U5974 , P3_U5973 );
nand NAND2_7391 ( P3_U3538 , P3_U5976 , P3_U5975 );
nand NAND2_7392 ( P3_U3539 , P3_U5978 , P3_U5977 );
nand NAND2_7393 ( P3_U3540 , P3_U5980 , P3_U5979 );
nand NAND2_7394 ( P3_U3541 , P3_U5982 , P3_U5981 );
nand NAND2_7395 ( P3_U3542 , P3_U5984 , P3_U5983 );
nand NAND2_7396 ( P3_U3543 , P3_U5986 , P3_U5985 );
nand NAND2_7397 ( P3_U3544 , P3_U5988 , P3_U5987 );
nand NAND2_7398 ( P3_U3545 , P3_U5990 , P3_U5989 );
nand NAND2_7399 ( P3_U3546 , P3_U5992 , P3_U5991 );
nand NAND2_7400 ( P3_U3547 , P3_U5994 , P3_U5993 );
nand NAND2_7401 ( P3_U3548 , P3_U5996 , P3_U5995 );
nand NAND2_7402 ( P3_U3549 , P3_U5998 , P3_U5997 );
nand NAND2_7403 ( P3_U3550 , P3_U6000 , P3_U5999 );
nand NAND2_7404 ( P3_U3551 , P3_U6002 , P3_U6001 );
nand NAND2_7405 ( P3_U3552 , P3_U6004 , P3_U6003 );
nand NAND2_7406 ( P3_U3553 , P3_U6006 , P3_U6005 );
nand NAND2_7407 ( P3_U3554 , P3_U6008 , P3_U6007 );
nand NAND2_7408 ( P3_U3555 , P3_U6010 , P3_U6009 );
nand NAND2_7409 ( P3_U3556 , P3_U6012 , P3_U6011 );
nand NAND2_7410 ( P3_U3557 , P3_U6014 , P3_U6013 );
nand NAND2_7411 ( P3_U3558 , P3_U6016 , P3_U6015 );
nand NAND2_7412 ( P3_U3559 , P3_U6018 , P3_U6017 );
nand NAND2_7413 ( P3_U3560 , P3_U6020 , P3_U6019 );
nand NAND2_7414 ( P3_U3561 , P3_U6022 , P3_U6021 );
nand NAND2_7415 ( P3_U3562 , P3_U6024 , P3_U6023 );
nand NAND2_7416 ( P3_U3563 , P3_U6026 , P3_U6025 );
nand NAND2_7417 ( P3_U3564 , P3_U6028 , P3_U6027 );
nand NAND2_7418 ( P3_U3565 , P3_U6030 , P3_U6029 );
nand NAND2_7419 ( P3_U3566 , P3_U6032 , P3_U6031 );
nand NAND2_7420 ( P3_U3567 , P3_U6034 , P3_U6033 );
nand NAND2_7421 ( P3_U3568 , P3_U6036 , P3_U6035 );
nand NAND2_7422 ( P3_U3569 , P3_U6038 , P3_U6037 );
nand NAND2_7423 ( P3_U3570 , P3_U6040 , P3_U6039 );
nand NAND2_7424 ( P3_U3571 , P3_U6042 , P3_U6041 );
nand NAND2_7425 ( P3_U3572 , P3_U6044 , P3_U6043 );
nand NAND2_7426 ( P3_U3573 , P3_U6046 , P3_U6045 );
nand NAND2_7427 ( P3_U3574 , P3_U6048 , P3_U6047 );
and AND2_7428 ( P3_U3575 , P3_U4066 , P3_U4065 );
and AND2_7429 ( P3_U3576 , P3_U4068 , P3_U4067 );
and AND3_7430 ( P3_U3577 , P3_U4076 , P3_U4074 , P3_U4075 );
and AND4_7431 ( P3_U3578 , P3_U4025 , P3_U4024 , P3_U4023 , P3_U4022 );
and AND4_7432 ( P3_U3579 , P3_U4029 , P3_U4028 , P3_U4027 , P3_U4026 );
and AND4_7433 ( P3_U3580 , P3_U4033 , P3_U4032 , P3_U4031 , P3_U4030 );
and AND3_7434 ( P3_U3581 , P3_U4035 , P3_U4034 , P3_U4036 );
and AND4_7435 ( P3_U3582 , P3_U3581 , P3_U3580 , P3_U3579 , P3_U3578 );
and AND4_7436 ( P3_U3583 , P3_U4040 , P3_U4039 , P3_U4038 , P3_U4037 );
and AND4_7437 ( P3_U3584 , P3_U4044 , P3_U4043 , P3_U4042 , P3_U4041 );
and AND4_7438 ( P3_U3585 , P3_U4048 , P3_U4047 , P3_U4046 , P3_U4045 );
and AND3_7439 ( P3_U3586 , P3_U4050 , P3_U4049 , P3_U4051 );
and AND4_7440 ( P3_U3587 , P3_U3586 , P3_U3585 , P3_U3584 , P3_U3583 );
and AND2_7441 ( P3_U3588 , P3_U3389 , P3_U3388 );
and AND2_7442 ( P3_U3589 , P3_U5479 , P3_U5476 );
and AND2_7443 ( P3_U3590 , P3_U4093 , P3_U4092 );
and AND2_7444 ( P3_U3591 , P3_U4095 , P3_U4094 );
and AND3_7445 ( P3_U3592 , P3_U4097 , P3_U4096 , P3_U3591 );
and AND3_7446 ( P3_U3593 , P3_U4100 , P3_U4101 , P3_U4099 );
and AND2_7447 ( P3_U3594 , P3_U4111 , P3_U4110 );
and AND2_7448 ( P3_U3595 , P3_U4113 , P3_U4112 );
and AND3_7449 ( P3_U3596 , P3_U4115 , P3_U4114 , P3_U3595 );
and AND3_7450 ( P3_U3597 , P3_U4118 , P3_U4119 , P3_U4117 );
and AND2_7451 ( P3_U3598 , P3_U4129 , P3_U4128 );
and AND2_7452 ( P3_U3599 , P3_U4131 , P3_U4130 );
and AND3_7453 ( P3_U3600 , P3_U4133 , P3_U4132 , P3_U3599 );
and AND3_7454 ( P3_U3601 , P3_U4136 , P3_U4137 , P3_U4135 );
and AND2_7455 ( P3_U3602 , P3_U4149 , P3_U4148 );
and AND3_7456 ( P3_U3603 , P3_U4151 , P3_U4150 , P3_U3602 );
and AND3_7457 ( P3_U3604 , P3_U4154 , P3_U4155 , P3_U4153 );
and AND2_7458 ( P3_U3605 , P3_U4167 , P3_U4166 );
and AND3_7459 ( P3_U3606 , P3_U4169 , P3_U4168 , P3_U3605 );
and AND3_7460 ( P3_U3607 , P3_U4172 , P3_U4173 , P3_U4171 );
and AND2_7461 ( P3_U3608 , P3_U4185 , P3_U4184 );
and AND3_7462 ( P3_U3609 , P3_U4187 , P3_U4186 , P3_U3608 );
and AND3_7463 ( P3_U3610 , P3_U4190 , P3_U4191 , P3_U4189 );
and AND2_7464 ( P3_U3611 , P3_U4203 , P3_U4202 );
and AND3_7465 ( P3_U3612 , P3_U4205 , P3_U4204 , P3_U3611 );
and AND3_7466 ( P3_U3613 , P3_U4208 , P3_U4209 , P3_U4207 );
and AND2_7467 ( P3_U3614 , P3_U4221 , P3_U4220 );
and AND3_7468 ( P3_U3615 , P3_U4223 , P3_U4222 , P3_U3614 );
and AND3_7469 ( P3_U3616 , P3_U4226 , P3_U4227 , P3_U4225 );
and AND2_7470 ( P3_U3617 , P3_U4237 , P3_U4236 );
and AND2_7471 ( P3_U3618 , P3_U4239 , P3_U4238 );
and AND3_7472 ( P3_U3619 , P3_U4241 , P3_U4240 , P3_U3618 );
and AND3_7473 ( P3_U3620 , P3_U4244 , P3_U4245 , P3_U4243 );
and AND2_7474 ( P3_U3621 , P3_U4255 , P3_U4254 );
and AND2_7475 ( P3_U3622 , P3_U4257 , P3_U4256 );
and AND3_7476 ( P3_U3623 , P3_U4259 , P3_U4258 , P3_U3622 );
and AND3_7477 ( P3_U3624 , P3_U4262 , P3_U4263 , P3_U4261 );
and AND2_7478 ( P3_U3625 , P3_U4275 , P3_U4274 );
and AND3_7479 ( P3_U3626 , P3_U4277 , P3_U4276 , P3_U3625 );
and AND3_7480 ( P3_U3627 , P3_U4280 , P3_U4281 , P3_U4279 );
and AND2_7481 ( P3_U3628 , P3_U4291 , P3_U4290 );
and AND2_7482 ( P3_U3629 , P3_U4293 , P3_U4292 );
and AND3_7483 ( P3_U3630 , P3_U4295 , P3_U4294 , P3_U3629 );
and AND3_7484 ( P3_U3631 , P3_U4298 , P3_U4299 , P3_U4297 );
and AND2_7485 ( P3_U3632 , P3_U4309 , P3_U4308 );
and AND2_7486 ( P3_U3633 , P3_U4311 , P3_U4310 );
and AND3_7487 ( P3_U3634 , P3_U4313 , P3_U4312 , P3_U3633 );
and AND3_7488 ( P3_U3635 , P3_U4316 , P3_U4317 , P3_U4315 );
and AND2_7489 ( P3_U3636 , P3_U4329 , P3_U4328 );
and AND3_7490 ( P3_U3637 , P3_U4331 , P3_U4330 , P3_U3636 );
and AND3_7491 ( P3_U3638 , P3_U4334 , P3_U4335 , P3_U4333 );
and AND2_7492 ( P3_U3639 , P3_U4347 , P3_U4346 );
and AND3_7493 ( P3_U3640 , P3_U4349 , P3_U4348 , P3_U3639 );
and AND3_7494 ( P3_U3641 , P3_U4352 , P3_U4353 , P3_U4351 );
and AND2_7495 ( P3_U3642 , P3_U4365 , P3_U4364 );
and AND3_7496 ( P3_U3643 , P3_U4367 , P3_U4366 , P3_U3642 );
and AND3_7497 ( P3_U3644 , P3_U4370 , P3_U4371 , P3_U4369 );
and AND2_7498 ( P3_U3645 , P3_U4381 , P3_U4380 );
and AND2_7499 ( P3_U3646 , P3_U4383 , P3_U4382 );
and AND3_7500 ( P3_U3647 , P3_U4385 , P3_U4384 , P3_U3646 );
and AND3_7501 ( P3_U3648 , P3_U4388 , P3_U4389 , P3_U4387 );
and AND2_7502 ( P3_U3649 , P3_U4401 , P3_U4400 );
and AND3_7503 ( P3_U3650 , P3_U4403 , P3_U4402 , P3_U3649 );
and AND3_7504 ( P3_U3651 , P3_U4406 , P3_U4407 , P3_U4405 );
and AND2_7505 ( P3_U3652 , P3_U4419 , P3_U4418 );
and AND3_7506 ( P3_U3653 , P3_U4421 , P3_U4420 , P3_U3652 );
and AND3_7507 ( P3_U3654 , P3_U4424 , P3_U4425 , P3_U4423 );
and AND2_7508 ( P3_U3655 , P3_U4437 , P3_U4436 );
and AND3_7509 ( P3_U3656 , P3_U4439 , P3_U4438 , P3_U3655 );
and AND3_7510 ( P3_U3657 , P3_U4442 , P3_U4443 , P3_U4441 );
and AND2_7511 ( P3_U3658 , P3_U4455 , P3_U4454 );
and AND3_7512 ( P3_U3659 , P3_U4457 , P3_U4456 , P3_U3658 );
and AND3_7513 ( P3_U3660 , P3_U4460 , P3_U4461 , P3_U4459 );
and AND2_7514 ( P3_U3661 , P3_U4473 , P3_U4472 );
and AND3_7515 ( P3_U3662 , P3_U4475 , P3_U4474 , P3_U3661 );
and AND3_7516 ( P3_U3663 , P3_U4478 , P3_U4479 , P3_U4477 );
and AND2_7517 ( P3_U3664 , P3_U4491 , P3_U4490 );
and AND3_7518 ( P3_U3665 , P3_U4493 , P3_U4492 , P3_U3664 );
and AND3_7519 ( P3_U3666 , P3_U4496 , P3_U4497 , P3_U4495 );
and AND2_7520 ( P3_U3667 , P3_U4507 , P3_U4506 );
and AND2_7521 ( P3_U3668 , P3_U4509 , P3_U4508 );
and AND3_7522 ( P3_U3669 , P3_U4511 , P3_U4510 , P3_U3668 );
and AND3_7523 ( P3_U3670 , P3_U4514 , P3_U4515 , P3_U4513 );
and AND2_7524 ( P3_U3671 , P3_U4525 , P3_U4524 );
and AND2_7525 ( P3_U3672 , P3_U4527 , P3_U4526 );
and AND3_7526 ( P3_U3673 , P3_U4529 , P3_U4528 , P3_U3672 );
and AND3_7527 ( P3_U3674 , P3_U4532 , P3_U4533 , P3_U4531 );
and AND2_7528 ( P3_U3675 , P3_U4543 , P3_U4542 );
and AND2_7529 ( P3_U3676 , P3_U4545 , P3_U4544 );
and AND3_7530 ( P3_U3677 , P3_U4547 , P3_U4546 , P3_U3676 );
and AND3_7531 ( P3_U3678 , P3_U4550 , P3_U4551 , P3_U4549 );
and AND2_7532 ( P3_U3679 , P3_U4561 , P3_U4560 );
and AND2_7533 ( P3_U3680 , P3_U4563 , P3_U4562 );
and AND3_7534 ( P3_U3681 , P3_U4565 , P3_U4564 , P3_U3680 );
and AND3_7535 ( P3_U3682 , P3_U4568 , P3_U4569 , P3_U4567 );
and AND2_7536 ( P3_U3683 , P3_U4579 , P3_U4578 );
and AND2_7537 ( P3_U3684 , P3_U4581 , P3_U4580 );
and AND3_7538 ( P3_U3685 , P3_U4583 , P3_U4582 , P3_U3684 );
and AND3_7539 ( P3_U3686 , P3_U4586 , P3_U4587 , P3_U4585 );
and AND2_7540 ( P3_U3687 , P3_U4600 , P3_U4599 );
and AND2_7541 ( P3_U3688 , P3_U4602 , P3_U4601 );
and AND3_7542 ( P3_U3689 , P3_U4604 , P3_U4603 , P3_U3688 );
and AND2_7543 ( P3_U3690 , P3_U4607 , P3_U4606 );
and AND2_7544 ( P3_U3691 , P3_U5476 , P3_U3389 );
and AND2_7545 ( P3_U3692 , P3_U5479 , P3_U3388 );
and AND2_7546 ( P3_U3693 , P3_U3920 , P3_U3379 );
and AND2_7547 ( P3_U3694 , P3_U5440 , P3_STATE_REG );
and AND2_7548 ( P3_U3695 , P3_U5424 , P3_U3364 );
and AND2_7549 ( P3_U3696 , P3_U3375 , P3_STATE_REG );
and AND5_7550 ( P3_U3697 , P3_U3301 , P3_U3308 , P3_U3305 , P3_U3306 , P3_U3307 );
and AND2_7551 ( P3_U3698 , P3_U3309 , P3_U3360 );
and AND4_7552 ( P3_U3699 , P3_U4763 , P3_U4762 , P3_U4765 , P3_U3701 );
and AND2_7553 ( P3_U3700 , P3_U4768 , P3_U4766 );
and AND2_7554 ( P3_U3701 , P3_U3700 , P3_U4767 );
and AND4_7555 ( P3_U3702 , P3_U4774 , P3_U4773 , P3_U4776 , P3_U3704 );
and AND2_7556 ( P3_U3703 , P3_U4779 , P3_U4777 );
and AND2_7557 ( P3_U3704 , P3_U3703 , P3_U4778 );
and AND4_7558 ( P3_U3705 , P3_U4785 , P3_U4784 , P3_U4787 , P3_U3707 );
and AND2_7559 ( P3_U3706 , P3_U4790 , P3_U4788 );
and AND2_7560 ( P3_U3707 , P3_U3706 , P3_U4789 );
and AND4_7561 ( P3_U3708 , P3_U4796 , P3_U4795 , P3_U4798 , P3_U3710 );
and AND2_7562 ( P3_U3709 , P3_U4801 , P3_U4799 );
and AND2_7563 ( P3_U3710 , P3_U3709 , P3_U4800 );
and AND4_7564 ( P3_U3711 , P3_U4807 , P3_U4806 , P3_U4809 , P3_U3713 );
and AND2_7565 ( P3_U3712 , P3_U4812 , P3_U4810 );
and AND2_7566 ( P3_U3713 , P3_U3712 , P3_U4811 );
and AND4_7567 ( P3_U3714 , P3_U4818 , P3_U4817 , P3_U4820 , P3_U3716 );
and AND2_7568 ( P3_U3715 , P3_U4823 , P3_U4821 );
and AND2_7569 ( P3_U3716 , P3_U3715 , P3_U4822 );
and AND4_7570 ( P3_U3717 , P3_U4829 , P3_U4828 , P3_U4831 , P3_U3719 );
and AND2_7571 ( P3_U3718 , P3_U4834 , P3_U4832 );
and AND2_7572 ( P3_U3719 , P3_U3718 , P3_U4833 );
and AND4_7573 ( P3_U3720 , P3_U4840 , P3_U4839 , P3_U4842 , P3_U3722 );
and AND2_7574 ( P3_U3721 , P3_U4845 , P3_U4843 );
and AND2_7575 ( P3_U3722 , P3_U3721 , P3_U4844 );
and AND4_7576 ( P3_U3723 , P3_U4851 , P3_U4850 , P3_U4853 , P3_U3725 );
and AND2_7577 ( P3_U3724 , P3_U4856 , P3_U4854 );
and AND2_7578 ( P3_U3725 , P3_U3724 , P3_U4855 );
and AND4_7579 ( P3_U3726 , P3_U4862 , P3_U4861 , P3_U4864 , P3_U3728 );
and AND2_7580 ( P3_U3727 , P3_U4867 , P3_U4865 );
and AND2_7581 ( P3_U3728 , P3_U3727 , P3_U4866 );
and AND4_7582 ( P3_U3729 , P3_U4873 , P3_U4872 , P3_U4875 , P3_U3731 );
and AND2_7583 ( P3_U3730 , P3_U4878 , P3_U4876 );
and AND2_7584 ( P3_U3731 , P3_U3730 , P3_U4877 );
and AND4_7585 ( P3_U3732 , P3_U4884 , P3_U4886 , P3_U4883 , P3_U3734 );
and AND2_7586 ( P3_U3733 , P3_U4889 , P3_U4887 );
and AND2_7587 ( P3_U3734 , P3_U3733 , P3_U4888 );
and AND4_7588 ( P3_U3735 , P3_U4895 , P3_U4897 , P3_U4894 , P3_U3737 );
and AND2_7589 ( P3_U3736 , P3_U4900 , P3_U4898 );
and AND2_7590 ( P3_U3737 , P3_U3736 , P3_U4899 );
and AND3_7591 ( P3_U3738 , P3_U4908 , P3_U4906 , P3_U3740 );
and AND2_7592 ( P3_U3739 , P3_U4911 , P3_U4909 );
and AND2_7593 ( P3_U3740 , P3_U3739 , P3_U4910 );
and AND2_7594 ( P3_U3741 , P3_U4919 , P3_U4917 );
and AND2_7595 ( P3_U3742 , P3_U4922 , P3_U4920 );
and AND2_7596 ( P3_U3743 , P3_U3742 , P3_U4921 );
and AND3_7597 ( P3_U3744 , P3_U4928 , P3_U3746 , P3_U4927 );
and AND2_7598 ( P3_U3745 , P3_U4933 , P3_U4931 );
and AND2_7599 ( P3_U3746 , P3_U3745 , P3_U4932 );
and AND3_7600 ( P3_U3747 , P3_U4939 , P3_U3749 , P3_U4938 );
and AND2_7601 ( P3_U3748 , P3_U4944 , P3_U4942 );
and AND2_7602 ( P3_U3749 , P3_U3748 , P3_U4943 );
and AND4_7603 ( P3_U3750 , P3_U4950 , P3_U4952 , P3_U4949 , P3_U3752 );
and AND2_7604 ( P3_U3751 , P3_U4955 , P3_U4953 );
and AND2_7605 ( P3_U3752 , P3_U3751 , P3_U4954 );
and AND4_7606 ( P3_U3753 , P3_U4961 , P3_U4960 , P3_U4963 , P3_U3755 );
and AND2_7607 ( P3_U3754 , P3_U4966 , P3_U4964 );
and AND2_7608 ( P3_U3755 , P3_U3754 , P3_U4965 );
and AND4_7609 ( P3_U3756 , P3_U4972 , P3_U4971 , P3_U4974 , P3_U3758 );
and AND2_7610 ( P3_U3757 , P3_U4977 , P3_U4975 );
and AND2_7611 ( P3_U3758 , P3_U3757 , P3_U4976 );
and AND2_7612 ( P3_U3759 , P3_U5468 , P3_U3383 );
nand NAND2_7613 ( P3_U3760 , P3_U5834 , P3_U5833 );
and AND2_7614 ( P3_U3761 , P3_U5915 , P3_U5912 );
and AND4_7615 ( P3_U3762 , P3_U3764 , P3_U3763 , P3_U3761 , P3_U5897 );
and AND2_7616 ( P3_U3763 , P3_U5903 , P3_U5900 );
and AND2_7617 ( P3_U3764 , P3_U5909 , P3_U5906 );
and AND3_7618 ( P3_U3765 , P3_U5885 , P3_U5882 , P3_U5879 );
and AND3_7619 ( P3_U3766 , P3_U5894 , P3_U5891 , P3_U5888 );
and AND4_7620 ( P3_U3767 , P3_U3766 , P3_U3765 , P3_U5876 , P3_U5873 );
and AND4_7621 ( P3_U3768 , P3_U5867 , P3_U5864 , P3_U5861 , P3_U5858 );
and AND2_7622 ( P3_U3769 , P3_U5855 , P3_U5852 );
and AND4_7623 ( P3_U3770 , P3_U5930 , P3_U5927 , P3_U5924 , P3_U5921 );
and AND3_7624 ( P3_U3771 , P3_U5843 , P3_U5840 , P3_U5846 );
and AND5_7625 ( P3_U3772 , P3_U3768 , P3_U3769 , P3_U5870 , P3_U5849 , P3_U3771 );
and AND5_7626 ( P3_U3773 , P3_U3762 , P3_U3767 , P3_U5918 , P3_U3770 , P3_U5933 );
and AND3_7627 ( P3_U3774 , P3_U4981 , P3_U3870 , P3_U4980 );
and AND2_7628 ( P3_U3775 , P3_U5416 , P3_U5415 );
and AND4_7629 ( P3_U3776 , P3_U5440 , P3_U3362 , P3_U4990 , P3_U3880 );
and AND2_7630 ( P3_U3777 , P3_U4998 , P3_U4997 );
and AND2_7631 ( P3_U3778 , P3_U5011 , P3_U5010 );
and AND2_7632 ( P3_U3779 , P3_U5020 , P3_U5019 );
and AND2_7633 ( P3_U3780 , P3_U5029 , P3_U5028 );
and AND2_7634 ( P3_U3781 , P3_U5036 , P3_U5034 );
and AND2_7635 ( P3_U3782 , P3_U5038 , P3_U5037 );
and AND2_7636 ( P3_U3783 , P3_U5047 , P3_U5046 );
and AND2_7637 ( P3_U3784 , P3_U5056 , P3_U5055 );
and AND2_7638 ( P3_U3785 , P3_U5065 , P3_U5064 );
and AND2_7639 ( P3_U3786 , P3_U5074 , P3_U5073 );
and AND2_7640 ( P3_U3787 , P3_U3031 , P3_U3077 );
and AND2_7641 ( P3_U3788 , P3_U5078 , P3_U5077 );
and AND3_7642 ( P3_U3789 , P3_U5081 , P3_U5080 , P3_U3788 );
and AND2_7643 ( P3_U3790 , P3_U5090 , P3_U5089 );
and AND2_7644 ( P3_U3791 , P3_U5097 , P3_U5095 );
and AND2_7645 ( P3_U3792 , P3_U5099 , P3_U5098 );
and AND2_7646 ( P3_U3793 , P3_U5108 , P3_U5107 );
and AND2_7647 ( P3_U3794 , P3_U5117 , P3_U5116 );
and AND2_7648 ( P3_U3795 , P3_U5126 , P3_U5125 );
and AND2_7649 ( P3_U3796 , P3_U5135 , P3_U5134 );
and AND2_7650 ( P3_U3797 , P3_U5144 , P3_U5143 );
and AND2_7651 ( P3_U3798 , P3_U5153 , P3_U5152 );
and AND2_7652 ( P3_U3799 , P3_U5162 , P3_U5161 );
and AND2_7653 ( P3_U3800 , P3_U5169 , P3_U5167 );
and AND2_7654 ( P3_U3801 , P3_U5171 , P3_U5170 );
and AND2_7655 ( P3_U3802 , P3_U5180 , P3_U5179 );
and AND2_7656 ( P3_U3803 , P3_U5189 , P3_U5188 );
and AND2_7657 ( P3_U3804 , P3_U5198 , P3_U5197 );
and AND2_7658 ( P3_U3805 , P3_U5205 , P3_U5203 );
and AND2_7659 ( P3_U3806 , P3_U5207 , P3_U5206 );
and AND2_7660 ( P3_U3807 , P3_U5216 , P3_U5215 );
and AND2_7661 ( P3_U3808 , P3_U5225 , P3_U5224 );
and AND2_7662 ( P3_U3809 , P3_U5234 , P3_U5233 );
and AND2_7663 ( P3_U3810 , P3_U5243 , P3_U5242 );
and AND2_7664 ( P3_U3811 , P3_U5252 , P3_U5251 );
and AND2_7665 ( P3_U3812 , P3_U5254 , P3_STATE_REG );
and AND2_7666 ( P3_U3813 , P3_U5440 , P3_U3385 );
and AND2_7667 ( P3_U3814 , P3_U3385 , P3_U3375 );
and AND3_7668 ( P3_U3815 , P3_U3875 , P3_U3312 , P3_U3302 );
and AND3_7669 ( P3_U3816 , P3_U3357 , P3_U3877 , P3_U3310 );
and AND2_7670 ( P3_U3817 , P3_U3375 , P3_U5258 );
and AND2_7671 ( P3_U3818 , P3_U3375 , P3_U5260 );
and AND2_7672 ( P3_U3819 , P3_U3375 , P3_U5262 );
and AND2_7673 ( P3_U3820 , P3_U3375 , P3_U5264 );
and AND2_7674 ( P3_U3821 , P3_U3375 , P3_U5266 );
and AND2_7675 ( P3_U3822 , P3_U3375 , P3_U5268 );
and AND2_7676 ( P3_U3823 , P3_U3375 , P3_U5274 );
and AND2_7677 ( P3_U3824 , P3_U3375 , P3_U5296 );
and AND2_7678 ( P3_U3825 , P3_U3375 , P3_U5310 );
and AND2_7679 ( P3_U3826 , P3_U3375 , P3_U5312 );
and AND2_7680 ( P3_U3827 , P3_U3375 , P3_U5314 );
and AND2_7681 ( P3_U3828 , P3_U3375 , P3_U5316 );
and AND2_7682 ( P3_U3829 , P3_U3375 , P3_U5318 );
and AND2_7683 ( P3_U3830 , P3_U3375 , P3_U5320 );
not NOT1_7684 ( P3_U3831 , P3_IR_REG_31_ );
nand NAND2_7685 ( P3_U3832 , P3_U3023 , P3_U3300 );
nand NAND2_7686 ( P3_U3833 , P3_U5468 , P3_U5465 );
nand NAND2_7687 ( P3_U3834 , P3_U5456 , P3_U5447 );
nand NAND2_7688 ( P3_U3835 , P3_U3023 , P3_U4058 );
nand NAND2_7689 ( P3_U3836 , P3_U3023 , P3_U4622 );
and AND2_7690 ( P3_U3837 , P3_U5707 , P3_U5706 );
and AND2_7691 ( P3_U3838 , P3_U5709 , P3_U5708 );
and AND2_7692 ( P3_U3839 , P3_U5711 , P3_U5710 );
and AND2_7693 ( P3_U3840 , P3_U5713 , P3_U5712 );
and AND2_7694 ( P3_U3841 , P3_U5715 , P3_U5714 );
and AND2_7695 ( P3_U3842 , P3_U5717 , P3_U5716 );
and AND2_7696 ( P3_U3843 , P3_U5719 , P3_U5718 );
and AND2_7697 ( P3_U3844 , P3_U5721 , P3_U5720 );
and AND2_7698 ( P3_U3845 , P3_U5723 , P3_U5722 );
and AND2_7699 ( P3_U3846 , P3_U5725 , P3_U5724 );
and AND2_7700 ( P3_U3847 , P3_U5727 , P3_U5726 );
and AND2_7701 ( P3_U3848 , P3_U5729 , P3_U5728 );
and AND2_7702 ( P3_U3849 , P3_U5731 , P3_U5730 );
and AND2_7703 ( P3_U3850 , P3_U5733 , P3_U5732 );
and AND2_7704 ( P3_U3851 , P3_U5735 , P3_U5734 );
and AND2_7705 ( P3_U3852 , P3_U5737 , P3_U5736 );
and AND2_7706 ( P3_U3853 , P3_U5739 , P3_U5738 );
and AND2_7707 ( P3_U3854 , P3_U5741 , P3_U5740 );
and AND2_7708 ( P3_U3855 , P3_U5743 , P3_U5742 );
and AND2_7709 ( P3_U3856 , P3_U5745 , P3_U5744 );
and AND2_7710 ( P3_U3857 , P3_U5747 , P3_U5746 );
and AND2_7711 ( P3_U3858 , P3_U5749 , P3_U5748 );
and AND2_7712 ( P3_U3859 , P3_U5751 , P3_U5750 );
and AND2_7713 ( P3_U3860 , P3_U5753 , P3_U5752 );
and AND2_7714 ( P3_U3861 , P3_U5755 , P3_U5754 );
and AND2_7715 ( P3_U3862 , P3_U5757 , P3_U5756 );
and AND2_7716 ( P3_U3863 , P3_U5759 , P3_U5758 );
and AND2_7717 ( P3_U3864 , P3_U5761 , P3_U5760 );
and AND2_7718 ( P3_U3865 , P3_U5763 , P3_U5762 );
and AND2_7719 ( P3_U3866 , P3_U5765 , P3_U5764 );
not NOT1_7720 ( P3_U3867 , P3_R1269_U11 );
nand NAND2_7721 ( P3_U3868 , P3_U3773 , P3_U3772 );
not NOT1_7722 ( P3_U3869 , P3_R693_U14 );
and AND2_7723 ( P3_U3870 , P3_U5940 , P3_U5939 );
not NOT1_7724 ( P3_U3871 , P3_R1297_U6 );
not NOT1_7725 ( P3_U3872 , P3_U3356 );
not NOT1_7726 ( P3_U3873 , P3_U3355 );
not NOT1_7727 ( P3_U3874 , P3_U3312 );
nand NAND2_7728 ( P3_U3875 , P3_U3015 , P3_U3385 );
not NOT1_7729 ( P3_U3876 , P3_U3302 );
nand NAND2_7730 ( P3_U3877 , P3_U3016 , P3_U5456 );
not NOT1_7731 ( P3_U3878 , P3_U3310 );
not NOT1_7732 ( P3_U3879 , P3_U3357 );
nand NAND2_7733 ( P3_U3880 , P3_U3014 , P3_U3385 );
not NOT1_7734 ( P3_U3881 , P3_U3308 );
not NOT1_7735 ( P3_U3882 , P3_U3301 );
not NOT1_7736 ( P3_U3883 , P3_U3305 );
not NOT1_7737 ( P3_U3884 , P3_U3307 );
not NOT1_7738 ( P3_U3885 , P3_U3306 );
not NOT1_7739 ( P3_U3886 , P3_U3360 );
not NOT1_7740 ( P3_U3887 , P3_U3311 );
nand NAND2_7741 ( P3_U3888 , P3_U3878 , P3_U3378 );
not NOT1_7742 ( P3_U3889 , P3_U3369 );
not NOT1_7743 ( P3_U3890 , P3_U3367 );
not NOT1_7744 ( P3_U3891 , P3_U3309 );
not NOT1_7745 ( P3_U3892 , P3_U3352 );
not NOT1_7746 ( P3_U3893 , P3_U3833 );
not NOT1_7747 ( P3_U3894 , P3_U3303 );
not NOT1_7748 ( P3_U3895 , P3_U3304 );
nand NAND2_7749 ( P3_U3896 , P3_U5465 , P3_U3384 );
not NOT1_7750 ( P3_U3897 , P3_U3363 );
not NOT1_7751 ( P3_U3898 , P3_U3364 );
not NOT1_7752 ( P3_U3899 , P3_U3350 );
not NOT1_7753 ( P3_U3900 , P3_U3348 );
not NOT1_7754 ( P3_U3901 , P3_U3346 );
not NOT1_7755 ( P3_U3902 , P3_U3344 );
not NOT1_7756 ( P3_U3903 , P3_U3342 );
not NOT1_7757 ( P3_U3904 , P3_U3340 );
not NOT1_7758 ( P3_U3905 , P3_U3338 );
not NOT1_7759 ( P3_U3906 , P3_U3336 );
not NOT1_7760 ( P3_U3907 , P3_U3334 );
not NOT1_7761 ( P3_U3908 , P3_U3353 );
not NOT1_7762 ( P3_U3909 , P3_U3368 );
not NOT1_7763 ( P3_U3910 , P3_U3362 );
not NOT1_7764 ( P3_U3911 , P3_U3313 );
not NOT1_7765 ( P3_U3912 , P3_U3358 );
not NOT1_7766 ( P3_U3913 , P3_U3836 );
not NOT1_7767 ( P3_U3914 , P3_U3835 );
not NOT1_7768 ( P3_U3915 , P3_U3832 );
not NOT1_7769 ( P3_U3916 , P3_U3361 );
nand NAND2_7770 ( P3_U3917 , P3_U3370 , P3_STATE_REG );
nand NAND2_7771 ( P3_U3918 , P3_U3886 , P3_U3023 );
not NOT1_7772 ( P3_U3919 , P3_U3299 );
not NOT1_7773 ( P3_U3920 , P3_U3359 );
not NOT1_7774 ( P3_U3921 , P3_U3297 );
nand NAND2_7775 ( P3_U3922 , U61 , P3_U3151 );
nand NAND2_7776 ( P3_U3923 , P3_IR_REG_0_ , P3_U3027 );
nand NAND2_7777 ( P3_U3924 , P3_IR_REG_0_ , P3_U3921 );
nand NAND2_7778 ( P3_U3925 , U50 , P3_U3151 );
nand NAND2_7779 ( P3_U3926 , P3_SUB_598_U51 , P3_U3027 );
nand NAND2_7780 ( P3_U3927 , P3_IR_REG_1_ , P3_U3921 );
nand NAND2_7781 ( P3_U3928 , U39 , P3_U3151 );
nand NAND2_7782 ( P3_U3929 , P3_SUB_598_U22 , P3_U3027 );
nand NAND2_7783 ( P3_U3930 , P3_IR_REG_2_ , P3_U3921 );
nand NAND2_7784 ( P3_U3931 , U36 , P3_U3151 );
nand NAND2_7785 ( P3_U3932 , P3_SUB_598_U23 , P3_U3027 );
nand NAND2_7786 ( P3_U3933 , P3_IR_REG_3_ , P3_U3921 );
nand NAND2_7787 ( P3_U3934 , U35 , P3_U3151 );
nand NAND2_7788 ( P3_U3935 , P3_SUB_598_U24 , P3_U3027 );
nand NAND2_7789 ( P3_U3936 , P3_IR_REG_4_ , P3_U3921 );
nand NAND2_7790 ( P3_U3937 , U34 , P3_U3151 );
nand NAND2_7791 ( P3_U3938 , P3_SUB_598_U74 , P3_U3027 );
nand NAND2_7792 ( P3_U3939 , P3_IR_REG_5_ , P3_U3921 );
nand NAND2_7793 ( P3_U3940 , U33 , P3_U3151 );
nand NAND2_7794 ( P3_U3941 , P3_SUB_598_U25 , P3_U3027 );
nand NAND2_7795 ( P3_U3942 , P3_IR_REG_6_ , P3_U3921 );
nand NAND2_7796 ( P3_U3943 , U32 , P3_U3151 );
nand NAND2_7797 ( P3_U3944 , P3_SUB_598_U26 , P3_U3027 );
nand NAND2_7798 ( P3_U3945 , P3_IR_REG_7_ , P3_U3921 );
nand NAND2_7799 ( P3_U3946 , U31 , P3_U3151 );
nand NAND2_7800 ( P3_U3947 , P3_SUB_598_U27 , P3_U3027 );
nand NAND2_7801 ( P3_U3948 , P3_IR_REG_8_ , P3_U3921 );
nand NAND2_7802 ( P3_U3949 , U30 , P3_U3151 );
nand NAND2_7803 ( P3_U3950 , P3_SUB_598_U72 , P3_U3027 );
nand NAND2_7804 ( P3_U3951 , P3_IR_REG_9_ , P3_U3921 );
nand NAND2_7805 ( P3_U3952 , U60 , P3_U3151 );
nand NAND2_7806 ( P3_U3953 , P3_SUB_598_U7 , P3_U3027 );
nand NAND2_7807 ( P3_U3954 , P3_IR_REG_10_ , P3_U3921 );
nand NAND2_7808 ( P3_U3955 , U59 , P3_U3151 );
nand NAND2_7809 ( P3_U3956 , P3_SUB_598_U8 , P3_U3027 );
nand NAND2_7810 ( P3_U3957 , P3_IR_REG_11_ , P3_U3921 );
nand NAND2_7811 ( P3_U3958 , U58 , P3_U3151 );
nand NAND2_7812 ( P3_U3959 , P3_SUB_598_U9 , P3_U3027 );
nand NAND2_7813 ( P3_U3960 , P3_IR_REG_12_ , P3_U3921 );
nand NAND2_7814 ( P3_U3961 , U57 , P3_U3151 );
nand NAND2_7815 ( P3_U3962 , P3_SUB_598_U89 , P3_U3027 );
nand NAND2_7816 ( P3_U3963 , P3_IR_REG_13_ , P3_U3921 );
nand NAND2_7817 ( P3_U3964 , U56 , P3_U3151 );
nand NAND2_7818 ( P3_U3965 , P3_SUB_598_U10 , P3_U3027 );
nand NAND2_7819 ( P3_U3966 , P3_IR_REG_14_ , P3_U3921 );
nand NAND2_7820 ( P3_U3967 , U55 , P3_U3151 );
nand NAND2_7821 ( P3_U3968 , P3_SUB_598_U11 , P3_U3027 );
nand NAND2_7822 ( P3_U3969 , P3_IR_REG_15_ , P3_U3921 );
nand NAND2_7823 ( P3_U3970 , U54 , P3_U3151 );
nand NAND2_7824 ( P3_U3971 , P3_SUB_598_U12 , P3_U3027 );
nand NAND2_7825 ( P3_U3972 , P3_IR_REG_16_ , P3_U3921 );
nand NAND2_7826 ( P3_U3973 , U53 , P3_U3151 );
nand NAND2_7827 ( P3_U3974 , P3_SUB_598_U87 , P3_U3027 );
nand NAND2_7828 ( P3_U3975 , P3_IR_REG_17_ , P3_U3921 );
nand NAND2_7829 ( P3_U3976 , U52 , P3_U3151 );
nand NAND2_7830 ( P3_U3977 , P3_SUB_598_U13 , P3_U3027 );
nand NAND2_7831 ( P3_U3978 , P3_IR_REG_18_ , P3_U3921 );
nand NAND2_7832 ( P3_U3979 , U51 , P3_U3151 );
nand NAND2_7833 ( P3_U3980 , P3_SUB_598_U14 , P3_U3027 );
nand NAND2_7834 ( P3_U3981 , P3_IR_REG_19_ , P3_U3921 );
nand NAND2_7835 ( P3_U3982 , U49 , P3_U3151 );
nand NAND2_7836 ( P3_U3983 , P3_SUB_598_U15 , P3_U3027 );
nand NAND2_7837 ( P3_U3984 , P3_IR_REG_20_ , P3_U3921 );
nand NAND2_7838 ( P3_U3985 , U48 , P3_U3151 );
nand NAND2_7839 ( P3_U3986 , P3_SUB_598_U83 , P3_U3027 );
nand NAND2_7840 ( P3_U3987 , P3_IR_REG_21_ , P3_U3921 );
nand NAND2_7841 ( P3_U3988 , U47 , P3_U3151 );
nand NAND2_7842 ( P3_U3989 , P3_SUB_598_U16 , P3_U3027 );
nand NAND2_7843 ( P3_U3990 , P3_IR_REG_22_ , P3_U3921 );
nand NAND2_7844 ( P3_U3991 , U46 , P3_U3151 );
nand NAND2_7845 ( P3_U3992 , P3_SUB_598_U17 , P3_U3027 );
nand NAND2_7846 ( P3_U3993 , P3_IR_REG_23_ , P3_U3921 );
nand NAND2_7847 ( P3_U3994 , U45 , P3_U3151 );
nand NAND2_7848 ( P3_U3995 , P3_SUB_598_U18 , P3_U3027 );
nand NAND2_7849 ( P3_U3996 , P3_IR_REG_24_ , P3_U3921 );
nand NAND2_7850 ( P3_U3997 , U44 , P3_U3151 );
nand NAND2_7851 ( P3_U3998 , P3_SUB_598_U81 , P3_U3027 );
nand NAND2_7852 ( P3_U3999 , P3_IR_REG_25_ , P3_U3921 );
nand NAND2_7853 ( P3_U4000 , U43 , P3_U3151 );
nand NAND2_7854 ( P3_U4001 , P3_SUB_598_U19 , P3_U3027 );
nand NAND2_7855 ( P3_U4002 , P3_IR_REG_26_ , P3_U3921 );
nand NAND2_7856 ( P3_U4003 , U42 , P3_U3151 );
nand NAND2_7857 ( P3_U4004 , P3_SUB_598_U79 , P3_U3027 );
nand NAND2_7858 ( P3_U4005 , P3_IR_REG_27_ , P3_U3921 );
nand NAND2_7859 ( P3_U4006 , U41 , P3_U3151 );
nand NAND2_7860 ( P3_U4007 , P3_SUB_598_U20 , P3_U3027 );
nand NAND2_7861 ( P3_U4008 , P3_IR_REG_28_ , P3_U3921 );
nand NAND2_7862 ( P3_U4009 , U40 , P3_U3151 );
nand NAND2_7863 ( P3_U4010 , P3_SUB_598_U21 , P3_U3027 );
nand NAND2_7864 ( P3_U4011 , P3_IR_REG_29_ , P3_U3921 );
nand NAND2_7865 ( P3_U4012 , U38 , P3_U3151 );
nand NAND2_7866 ( P3_U4013 , P3_SUB_598_U77 , P3_U3027 );
nand NAND2_7867 ( P3_U4014 , P3_IR_REG_30_ , P3_U3921 );
nand NAND2_7868 ( P3_U4015 , U37 , P3_U3151 );
nand NAND2_7869 ( P3_U4016 , P3_SUB_598_U52 , P3_U3027 );
nand NAND2_7870 ( P3_U4017 , P3_IR_REG_31_ , P3_U3921 );
nand NAND2_7871 ( P3_U4018 , P3_U3919 , P3_U5437 );
not NOT1_7872 ( P3_U4019 , P3_U3300 );
nand NAND2_7873 ( P3_U4020 , P3_U3299 , P3_U5428 );
nand NAND2_7874 ( P3_U4021 , P3_U3299 , P3_U5431 );
nand NAND2_7875 ( P3_U4022 , P3_U4019 , P3_D_REG_10_ );
nand NAND2_7876 ( P3_U4023 , P3_U4019 , P3_D_REG_11_ );
nand NAND2_7877 ( P3_U4024 , P3_U4019 , P3_D_REG_12_ );
nand NAND2_7878 ( P3_U4025 , P3_U4019 , P3_D_REG_13_ );
nand NAND2_7879 ( P3_U4026 , P3_U4019 , P3_D_REG_14_ );
nand NAND2_7880 ( P3_U4027 , P3_U4019 , P3_D_REG_15_ );
nand NAND2_7881 ( P3_U4028 , P3_U4019 , P3_D_REG_16_ );
nand NAND2_7882 ( P3_U4029 , P3_U4019 , P3_D_REG_17_ );
nand NAND2_7883 ( P3_U4030 , P3_U4019 , P3_D_REG_18_ );
nand NAND2_7884 ( P3_U4031 , P3_U4019 , P3_D_REG_19_ );
nand NAND2_7885 ( P3_U4032 , P3_U4019 , P3_D_REG_20_ );
nand NAND2_7886 ( P3_U4033 , P3_U4019 , P3_D_REG_21_ );
nand NAND2_7887 ( P3_U4034 , P3_U4019 , P3_D_REG_22_ );
nand NAND2_7888 ( P3_U4035 , P3_U4019 , P3_D_REG_23_ );
nand NAND2_7889 ( P3_U4036 , P3_U4019 , P3_D_REG_24_ );
nand NAND2_7890 ( P3_U4037 , P3_U4019 , P3_D_REG_25_ );
nand NAND2_7891 ( P3_U4038 , P3_U4019 , P3_D_REG_26_ );
nand NAND2_7892 ( P3_U4039 , P3_U4019 , P3_D_REG_27_ );
nand NAND2_7893 ( P3_U4040 , P3_U4019 , P3_D_REG_28_ );
nand NAND2_7894 ( P3_U4041 , P3_U4019 , P3_D_REG_29_ );
nand NAND2_7895 ( P3_U4042 , P3_U4019 , P3_D_REG_2_ );
nand NAND2_7896 ( P3_U4043 , P3_U4019 , P3_D_REG_30_ );
nand NAND2_7897 ( P3_U4044 , P3_U4019 , P3_D_REG_31_ );
nand NAND2_7898 ( P3_U4045 , P3_U4019 , P3_D_REG_3_ );
nand NAND2_7899 ( P3_U4046 , P3_U4019 , P3_D_REG_4_ );
nand NAND2_7900 ( P3_U4047 , P3_U4019 , P3_D_REG_5_ );
nand NAND2_7901 ( P3_U4048 , P3_U4019 , P3_D_REG_6_ );
nand NAND2_7902 ( P3_U4049 , P3_U4019 , P3_D_REG_7_ );
nand NAND2_7903 ( P3_U4050 , P3_U4019 , P3_D_REG_8_ );
nand NAND2_7904 ( P3_U4051 , P3_U4019 , P3_D_REG_9_ );
not NOT1_7905 ( P3_U4052 , P3_U3834 );
nand NAND2_7906 ( P3_U4053 , P3_U5456 , P3_U5450 );
nand NAND2_7907 ( P3_U4054 , P3_U5482 , P3_U4053 );
nand NAND2_7908 ( P3_U4055 , P3_U3369 , P3_U3367 );
nand NAND2_7909 ( P3_U4056 , P3_U3894 , P3_U4055 );
nand NAND2_7910 ( P3_U4057 , P3_U3895 , P3_U4054 );
nand NAND2_7911 ( P3_U4058 , P3_U4057 , P3_U4056 );
nand NAND2_7912 ( P3_U4059 , P3_U3022 , P3_REG0_REG_1_ );
nand NAND2_7913 ( P3_U4060 , P3_REG1_REG_1_ , P3_U3021 );
nand NAND2_7914 ( P3_U4061 , P3_REG2_REG_1_ , P3_U3020 );
nand NAND2_7915 ( P3_U4062 , P3_REG3_REG_1_ , P3_U3019 );
not NOT1_7916 ( P3_U4063 , P3_U3077 );
nand NAND2_7917 ( P3_U4064 , P3_U3877 , P3_U3357 );
nand NAND2_7918 ( P3_U4065 , P3_U3883 , P3_R1110_U95 );
nand NAND2_7919 ( P3_U4066 , P3_U3885 , P3_R1077_U95 );
nand NAND2_7920 ( P3_U4067 , P3_U3884 , P3_R1095_U24 );
nand NAND2_7921 ( P3_U4068 , P3_U3881 , P3_R1143_U95 );
nand NAND2_7922 ( P3_U4069 , P3_U3891 , P3_R1161_U95 );
nand NAND2_7923 ( P3_U4070 , P3_U3887 , P3_R1131_U24 );
nand NAND2_7924 ( P3_U4071 , P3_U3017 , P3_R1200_U24 );
not NOT1_7925 ( P3_U4072 , P3_U3314 );
nand NAND2_7926 ( P3_U4073 , P3_U3352 , P3_U3833 );
nand NAND2_7927 ( P3_U4074 , P3_R1179_U24 , P3_U3026 );
nand NAND2_7928 ( P3_U4075 , P3_U3025 , P3_U3077 );
nand NAND2_7929 ( P3_U4076 , P3_U3387 , P3_U4064 );
nand NAND2_7930 ( P3_U4077 , P3_U3577 , P3_U4072 );
nand NAND2_7931 ( P3_U4078 , P3_REG0_REG_2_ , P3_U3022 );
nand NAND2_7932 ( P3_U4079 , P3_REG1_REG_2_ , P3_U3021 );
nand NAND2_7933 ( P3_U4080 , P3_REG2_REG_2_ , P3_U3020 );
nand NAND2_7934 ( P3_U4081 , P3_REG3_REG_2_ , P3_U3019 );
not NOT1_7935 ( P3_U4082 , P3_U3067 );
nand NAND2_7936 ( P3_U4083 , P3_REG0_REG_0_ , P3_U3022 );
nand NAND2_7937 ( P3_U4084 , P3_REG1_REG_0_ , P3_U3021 );
nand NAND2_7938 ( P3_U4085 , P3_REG2_REG_0_ , P3_U3020 );
nand NAND2_7939 ( P3_U4086 , P3_REG3_REG_0_ , P3_U3019 );
not NOT1_7940 ( P3_U4087 , P3_U3076 );
nand NAND2_7941 ( P3_U4088 , P3_U5468 , P3_U3383 );
nand NAND2_7942 ( P3_U4089 , P3_U3896 , P3_U4088 );
nand NAND2_7943 ( P3_U4090 , P3_U3033 , P3_U3076 );
nand NAND2_7944 ( P3_U4091 , P3_R1110_U94 , P3_U3883 );
nand NAND2_7945 ( P3_U4092 , P3_R1077_U94 , P3_U3885 );
nand NAND2_7946 ( P3_U4093 , P3_R1095_U100 , P3_U3884 );
nand NAND2_7947 ( P3_U4094 , P3_R1143_U94 , P3_U3881 );
nand NAND2_7948 ( P3_U4095 , P3_R1161_U94 , P3_U3891 );
nand NAND2_7949 ( P3_U4096 , P3_R1131_U100 , P3_U3887 );
nand NAND2_7950 ( P3_U4097 , P3_R1200_U100 , P3_U3017 );
not NOT1_7951 ( P3_U4098 , P3_U3315 );
nand NAND2_7952 ( P3_U4099 , P3_R1179_U100 , P3_U3026 );
nand NAND2_7953 ( P3_U4100 , P3_U3025 , P3_U3067 );
nand NAND2_7954 ( P3_U4101 , P3_U3392 , P3_U4064 );
nand NAND2_7955 ( P3_U4102 , P3_U3593 , P3_U4098 );
nand NAND2_7956 ( P3_U4103 , P3_REG0_REG_3_ , P3_U3022 );
nand NAND2_7957 ( P3_U4104 , P3_REG1_REG_3_ , P3_U3021 );
nand NAND2_7958 ( P3_U4105 , P3_REG2_REG_3_ , P3_U3020 );
nand NAND2_7959 ( P3_U4106 , P3_SUB_609_U25 , P3_U3019 );
not NOT1_7960 ( P3_U4107 , P3_U3063 );
nand NAND2_7961 ( P3_U4108 , P3_U3033 , P3_U3077 );
nand NAND2_7962 ( P3_U4109 , P3_R1110_U16 , P3_U3883 );
nand NAND2_7963 ( P3_U4110 , P3_R1077_U16 , P3_U3885 );
nand NAND2_7964 ( P3_U4111 , P3_R1095_U110 , P3_U3884 );
nand NAND2_7965 ( P3_U4112 , P3_R1143_U16 , P3_U3881 );
nand NAND2_7966 ( P3_U4113 , P3_R1161_U16 , P3_U3891 );
nand NAND2_7967 ( P3_U4114 , P3_R1131_U110 , P3_U3887 );
nand NAND2_7968 ( P3_U4115 , P3_R1200_U110 , P3_U3017 );
not NOT1_7969 ( P3_U4116 , P3_U3316 );
nand NAND2_7970 ( P3_U4117 , P3_R1179_U110 , P3_U3026 );
nand NAND2_7971 ( P3_U4118 , P3_U3025 , P3_U3063 );
nand NAND2_7972 ( P3_U4119 , P3_U3395 , P3_U4064 );
nand NAND2_7973 ( P3_U4120 , P3_U3597 , P3_U4116 );
nand NAND2_7974 ( P3_U4121 , P3_REG0_REG_4_ , P3_U3022 );
nand NAND2_7975 ( P3_U4122 , P3_REG1_REG_4_ , P3_U3021 );
nand NAND2_7976 ( P3_U4123 , P3_REG2_REG_4_ , P3_U3020 );
nand NAND2_7977 ( P3_U4124 , P3_SUB_609_U29 , P3_U3019 );
not NOT1_7978 ( P3_U4125 , P3_U3059 );
nand NAND2_7979 ( P3_U4126 , P3_U3033 , P3_U3067 );
nand NAND2_7980 ( P3_U4127 , P3_R1110_U100 , P3_U3883 );
nand NAND2_7981 ( P3_U4128 , P3_R1077_U100 , P3_U3885 );
nand NAND2_7982 ( P3_U4129 , P3_R1095_U21 , P3_U3884 );
nand NAND2_7983 ( P3_U4130 , P3_R1143_U100 , P3_U3881 );
nand NAND2_7984 ( P3_U4131 , P3_R1161_U100 , P3_U3891 );
nand NAND2_7985 ( P3_U4132 , P3_R1131_U21 , P3_U3887 );
nand NAND2_7986 ( P3_U4133 , P3_R1200_U21 , P3_U3017 );
not NOT1_7987 ( P3_U4134 , P3_U3317 );
nand NAND2_7988 ( P3_U4135 , P3_R1179_U21 , P3_U3026 );
nand NAND2_7989 ( P3_U4136 , P3_U3025 , P3_U3059 );
nand NAND2_7990 ( P3_U4137 , P3_U3398 , P3_U4064 );
nand NAND2_7991 ( P3_U4138 , P3_U3601 , P3_U4134 );
nand NAND2_7992 ( P3_U4139 , P3_REG0_REG_5_ , P3_U3022 );
nand NAND2_7993 ( P3_U4140 , P3_REG1_REG_5_ , P3_U3021 );
nand NAND2_7994 ( P3_U4141 , P3_REG2_REG_5_ , P3_U3020 );
nand NAND2_7995 ( P3_U4142 , P3_SUB_609_U53 , P3_U3019 );
not NOT1_7996 ( P3_U4143 , P3_U3066 );
nand NAND2_7997 ( P3_U4144 , P3_U3033 , P3_U3063 );
nand NAND2_7998 ( P3_U4145 , P3_R1110_U99 , P3_U3883 );
nand NAND2_7999 ( P3_U4146 , P3_R1077_U99 , P3_U3885 );
nand NAND2_8000 ( P3_U4147 , P3_R1095_U109 , P3_U3884 );
nand NAND2_8001 ( P3_U4148 , P3_R1143_U99 , P3_U3881 );
nand NAND2_8002 ( P3_U4149 , P3_R1161_U99 , P3_U3891 );
nand NAND2_8003 ( P3_U4150 , P3_R1131_U109 , P3_U3887 );
nand NAND2_8004 ( P3_U4151 , P3_R1200_U109 , P3_U3017 );
not NOT1_8005 ( P3_U4152 , P3_U3318 );
nand NAND2_8006 ( P3_U4153 , P3_R1179_U109 , P3_U3026 );
nand NAND2_8007 ( P3_U4154 , P3_U3025 , P3_U3066 );
nand NAND2_8008 ( P3_U4155 , P3_U3401 , P3_U4064 );
nand NAND2_8009 ( P3_U4156 , P3_U3604 , P3_U4152 );
nand NAND2_8010 ( P3_U4157 , P3_REG0_REG_6_ , P3_U3022 );
nand NAND2_8011 ( P3_U4158 , P3_REG1_REG_6_ , P3_U3021 );
nand NAND2_8012 ( P3_U4159 , P3_REG2_REG_6_ , P3_U3020 );
nand NAND2_8013 ( P3_U4160 , P3_SUB_609_U8 , P3_U3019 );
not NOT1_8014 ( P3_U4161 , P3_U3070 );
nand NAND2_8015 ( P3_U4162 , P3_U3033 , P3_U3059 );
nand NAND2_8016 ( P3_U4163 , P3_R1110_U17 , P3_U3883 );
nand NAND2_8017 ( P3_U4164 , P3_R1077_U17 , P3_U3885 );
nand NAND2_8018 ( P3_U4165 , P3_R1095_U108 , P3_U3884 );
nand NAND2_8019 ( P3_U4166 , P3_R1143_U17 , P3_U3881 );
nand NAND2_8020 ( P3_U4167 , P3_R1161_U17 , P3_U3891 );
nand NAND2_8021 ( P3_U4168 , P3_R1131_U108 , P3_U3887 );
nand NAND2_8022 ( P3_U4169 , P3_R1200_U108 , P3_U3017 );
not NOT1_8023 ( P3_U4170 , P3_U3319 );
nand NAND2_8024 ( P3_U4171 , P3_R1179_U108 , P3_U3026 );
nand NAND2_8025 ( P3_U4172 , P3_U3025 , P3_U3070 );
nand NAND2_8026 ( P3_U4173 , P3_U3404 , P3_U4064 );
nand NAND2_8027 ( P3_U4174 , P3_U3607 , P3_U4170 );
nand NAND2_8028 ( P3_U4175 , P3_REG0_REG_7_ , P3_U3022 );
nand NAND2_8029 ( P3_U4176 , P3_REG1_REG_7_ , P3_U3021 );
nand NAND2_8030 ( P3_U4177 , P3_REG2_REG_7_ , P3_U3020 );
nand NAND2_8031 ( P3_U4178 , P3_SUB_609_U18 , P3_U3019 );
not NOT1_8032 ( P3_U4179 , P3_U3069 );
nand NAND2_8033 ( P3_U4180 , P3_U3033 , P3_U3066 );
nand NAND2_8034 ( P3_U4181 , P3_R1110_U98 , P3_U3883 );
nand NAND2_8035 ( P3_U4182 , P3_R1077_U98 , P3_U3885 );
nand NAND2_8036 ( P3_U4183 , P3_R1095_U22 , P3_U3884 );
nand NAND2_8037 ( P3_U4184 , P3_R1143_U98 , P3_U3881 );
nand NAND2_8038 ( P3_U4185 , P3_R1161_U98 , P3_U3891 );
nand NAND2_8039 ( P3_U4186 , P3_R1131_U22 , P3_U3887 );
nand NAND2_8040 ( P3_U4187 , P3_R1200_U22 , P3_U3017 );
not NOT1_8041 ( P3_U4188 , P3_U3320 );
nand NAND2_8042 ( P3_U4189 , P3_R1179_U22 , P3_U3026 );
nand NAND2_8043 ( P3_U4190 , P3_U3025 , P3_U3069 );
nand NAND2_8044 ( P3_U4191 , P3_U3407 , P3_U4064 );
nand NAND2_8045 ( P3_U4192 , P3_U3610 , P3_U4188 );
nand NAND2_8046 ( P3_U4193 , P3_REG0_REG_8_ , P3_U3022 );
nand NAND2_8047 ( P3_U4194 , P3_REG1_REG_8_ , P3_U3021 );
nand NAND2_8048 ( P3_U4195 , P3_REG2_REG_8_ , P3_U3020 );
nand NAND2_8049 ( P3_U4196 , P3_SUB_609_U12 , P3_U3019 );
not NOT1_8050 ( P3_U4197 , P3_U3083 );
nand NAND2_8051 ( P3_U4198 , P3_U3033 , P3_U3070 );
nand NAND2_8052 ( P3_U4199 , P3_R1110_U18 , P3_U3883 );
nand NAND2_8053 ( P3_U4200 , P3_R1077_U18 , P3_U3885 );
nand NAND2_8054 ( P3_U4201 , P3_R1095_U107 , P3_U3884 );
nand NAND2_8055 ( P3_U4202 , P3_R1143_U18 , P3_U3881 );
nand NAND2_8056 ( P3_U4203 , P3_R1161_U18 , P3_U3891 );
nand NAND2_8057 ( P3_U4204 , P3_R1131_U107 , P3_U3887 );
nand NAND2_8058 ( P3_U4205 , P3_R1200_U107 , P3_U3017 );
not NOT1_8059 ( P3_U4206 , P3_U3321 );
nand NAND2_8060 ( P3_U4207 , P3_R1179_U107 , P3_U3026 );
nand NAND2_8061 ( P3_U4208 , P3_U3025 , P3_U3083 );
nand NAND2_8062 ( P3_U4209 , P3_U3410 , P3_U4064 );
nand NAND2_8063 ( P3_U4210 , P3_U3613 , P3_U4206 );
nand NAND2_8064 ( P3_U4211 , P3_REG0_REG_9_ , P3_U3022 );
nand NAND2_8065 ( P3_U4212 , P3_REG1_REG_9_ , P3_U3021 );
nand NAND2_8066 ( P3_U4213 , P3_REG2_REG_9_ , P3_U3020 );
nand NAND2_8067 ( P3_U4214 , P3_SUB_609_U14 , P3_U3019 );
not NOT1_8068 ( P3_U4215 , P3_U3082 );
nand NAND2_8069 ( P3_U4216 , P3_U3033 , P3_U3069 );
nand NAND2_8070 ( P3_U4217 , P3_R1110_U97 , P3_U3883 );
nand NAND2_8071 ( P3_U4218 , P3_R1077_U97 , P3_U3885 );
nand NAND2_8072 ( P3_U4219 , P3_R1095_U23 , P3_U3884 );
nand NAND2_8073 ( P3_U4220 , P3_R1143_U97 , P3_U3881 );
nand NAND2_8074 ( P3_U4221 , P3_R1161_U97 , P3_U3891 );
nand NAND2_8075 ( P3_U4222 , P3_R1131_U23 , P3_U3887 );
nand NAND2_8076 ( P3_U4223 , P3_R1200_U23 , P3_U3017 );
not NOT1_8077 ( P3_U4224 , P3_U3322 );
nand NAND2_8078 ( P3_U4225 , P3_R1179_U23 , P3_U3026 );
nand NAND2_8079 ( P3_U4226 , P3_U3025 , P3_U3082 );
nand NAND2_8080 ( P3_U4227 , P3_U3413 , P3_U4064 );
nand NAND2_8081 ( P3_U4228 , P3_U3616 , P3_U4224 );
nand NAND2_8082 ( P3_U4229 , P3_REG0_REG_10_ , P3_U3022 );
nand NAND2_8083 ( P3_U4230 , P3_REG1_REG_10_ , P3_U3021 );
nand NAND2_8084 ( P3_U4231 , P3_REG2_REG_10_ , P3_U3020 );
nand NAND2_8085 ( P3_U4232 , P3_SUB_609_U13 , P3_U3019 );
not NOT1_8086 ( P3_U4233 , P3_U3061 );
nand NAND2_8087 ( P3_U4234 , P3_U3033 , P3_U3083 );
nand NAND2_8088 ( P3_U4235 , P3_R1110_U96 , P3_U3883 );
nand NAND2_8089 ( P3_U4236 , P3_R1077_U96 , P3_U3885 );
nand NAND2_8090 ( P3_U4237 , P3_R1095_U106 , P3_U3884 );
nand NAND2_8091 ( P3_U4238 , P3_R1143_U96 , P3_U3881 );
nand NAND2_8092 ( P3_U4239 , P3_R1161_U96 , P3_U3891 );
nand NAND2_8093 ( P3_U4240 , P3_R1131_U106 , P3_U3887 );
nand NAND2_8094 ( P3_U4241 , P3_R1200_U106 , P3_U3017 );
not NOT1_8095 ( P3_U4242 , P3_U3323 );
nand NAND2_8096 ( P3_U4243 , P3_R1179_U106 , P3_U3026 );
nand NAND2_8097 ( P3_U4244 , P3_U3025 , P3_U3061 );
nand NAND2_8098 ( P3_U4245 , P3_U3416 , P3_U4064 );
nand NAND2_8099 ( P3_U4246 , P3_U3620 , P3_U4242 );
nand NAND2_8100 ( P3_U4247 , P3_REG0_REG_11_ , P3_U3022 );
nand NAND2_8101 ( P3_U4248 , P3_REG1_REG_11_ , P3_U3021 );
nand NAND2_8102 ( P3_U4249 , P3_REG2_REG_11_ , P3_U3020 );
nand NAND2_8103 ( P3_U4250 , P3_SUB_609_U9 , P3_U3019 );
not NOT1_8104 ( P3_U4251 , P3_U3062 );
nand NAND2_8105 ( P3_U4252 , P3_U3033 , P3_U3082 );
nand NAND2_8106 ( P3_U4253 , P3_R1110_U10 , P3_U3883 );
nand NAND2_8107 ( P3_U4254 , P3_R1077_U10 , P3_U3885 );
nand NAND2_8108 ( P3_U4255 , P3_R1095_U116 , P3_U3884 );
nand NAND2_8109 ( P3_U4256 , P3_R1143_U10 , P3_U3881 );
nand NAND2_8110 ( P3_U4257 , P3_R1161_U10 , P3_U3891 );
nand NAND2_8111 ( P3_U4258 , P3_R1131_U116 , P3_U3887 );
nand NAND2_8112 ( P3_U4259 , P3_R1200_U116 , P3_U3017 );
not NOT1_8113 ( P3_U4260 , P3_U3324 );
nand NAND2_8114 ( P3_U4261 , P3_R1179_U116 , P3_U3026 );
nand NAND2_8115 ( P3_U4262 , P3_U3025 , P3_U3062 );
nand NAND2_8116 ( P3_U4263 , P3_U3419 , P3_U4064 );
nand NAND2_8117 ( P3_U4264 , P3_U3624 , P3_U4260 );
nand NAND2_8118 ( P3_U4265 , P3_REG0_REG_12_ , P3_U3022 );
nand NAND2_8119 ( P3_U4266 , P3_REG1_REG_12_ , P3_U3021 );
nand NAND2_8120 ( P3_U4267 , P3_REG2_REG_12_ , P3_U3020 );
nand NAND2_8121 ( P3_U4268 , P3_SUB_609_U23 , P3_U3019 );
not NOT1_8122 ( P3_U4269 , P3_U3071 );
nand NAND2_8123 ( P3_U4270 , P3_U3033 , P3_U3061 );
nand NAND2_8124 ( P3_U4271 , P3_R1110_U114 , P3_U3883 );
nand NAND2_8125 ( P3_U4272 , P3_R1077_U114 , P3_U3885 );
nand NAND2_8126 ( P3_U4273 , P3_R1095_U16 , P3_U3884 );
nand NAND2_8127 ( P3_U4274 , P3_R1143_U114 , P3_U3881 );
nand NAND2_8128 ( P3_U4275 , P3_R1161_U114 , P3_U3891 );
nand NAND2_8129 ( P3_U4276 , P3_R1131_U16 , P3_U3887 );
nand NAND2_8130 ( P3_U4277 , P3_R1200_U16 , P3_U3017 );
not NOT1_8131 ( P3_U4278 , P3_U3325 );
nand NAND2_8132 ( P3_U4279 , P3_R1179_U16 , P3_U3026 );
nand NAND2_8133 ( P3_U4280 , P3_U3025 , P3_U3071 );
nand NAND2_8134 ( P3_U4281 , P3_U3422 , P3_U4064 );
nand NAND2_8135 ( P3_U4282 , P3_U3627 , P3_U4278 );
nand NAND2_8136 ( P3_U4283 , P3_REG0_REG_13_ , P3_U3022 );
nand NAND2_8137 ( P3_U4284 , P3_REG1_REG_13_ , P3_U3021 );
nand NAND2_8138 ( P3_U4285 , P3_REG2_REG_13_ , P3_U3020 );
nand NAND2_8139 ( P3_U4286 , P3_SUB_609_U24 , P3_U3019 );
not NOT1_8140 ( P3_U4287 , P3_U3079 );
nand NAND2_8141 ( P3_U4288 , P3_U3033 , P3_U3062 );
nand NAND2_8142 ( P3_U4289 , P3_R1110_U113 , P3_U3883 );
nand NAND2_8143 ( P3_U4290 , P3_R1077_U113 , P3_U3885 );
nand NAND2_8144 ( P3_U4291 , P3_R1095_U105 , P3_U3884 );
nand NAND2_8145 ( P3_U4292 , P3_R1143_U113 , P3_U3881 );
nand NAND2_8146 ( P3_U4293 , P3_R1161_U113 , P3_U3891 );
nand NAND2_8147 ( P3_U4294 , P3_R1131_U105 , P3_U3887 );
nand NAND2_8148 ( P3_U4295 , P3_R1200_U105 , P3_U3017 );
not NOT1_8149 ( P3_U4296 , P3_U3326 );
nand NAND2_8150 ( P3_U4297 , P3_R1179_U105 , P3_U3026 );
nand NAND2_8151 ( P3_U4298 , P3_U3025 , P3_U3079 );
nand NAND2_8152 ( P3_U4299 , P3_U3425 , P3_U4064 );
nand NAND2_8153 ( P3_U4300 , P3_U3631 , P3_U4296 );
nand NAND2_8154 ( P3_U4301 , P3_REG0_REG_14_ , P3_U3022 );
nand NAND2_8155 ( P3_U4302 , P3_REG1_REG_14_ , P3_U3021 );
nand NAND2_8156 ( P3_U4303 , P3_REG2_REG_14_ , P3_U3020 );
nand NAND2_8157 ( P3_U4304 , P3_SUB_609_U30 , P3_U3019 );
not NOT1_8158 ( P3_U4305 , P3_U3078 );
nand NAND2_8159 ( P3_U4306 , P3_U3033 , P3_U3071 );
nand NAND2_8160 ( P3_U4307 , P3_R1110_U11 , P3_U3883 );
nand NAND2_8161 ( P3_U4308 , P3_R1077_U11 , P3_U3885 );
nand NAND2_8162 ( P3_U4309 , P3_R1095_U104 , P3_U3884 );
nand NAND2_8163 ( P3_U4310 , P3_R1143_U11 , P3_U3881 );
nand NAND2_8164 ( P3_U4311 , P3_R1161_U11 , P3_U3891 );
nand NAND2_8165 ( P3_U4312 , P3_R1131_U104 , P3_U3887 );
nand NAND2_8166 ( P3_U4313 , P3_R1200_U104 , P3_U3017 );
not NOT1_8167 ( P3_U4314 , P3_U3327 );
nand NAND2_8168 ( P3_U4315 , P3_R1179_U104 , P3_U3026 );
nand NAND2_8169 ( P3_U4316 , P3_U3025 , P3_U3078 );
nand NAND2_8170 ( P3_U4317 , P3_U3428 , P3_U4064 );
nand NAND2_8171 ( P3_U4318 , P3_U3635 , P3_U4314 );
nand NAND2_8172 ( P3_U4319 , P3_REG0_REG_15_ , P3_U3022 );
nand NAND2_8173 ( P3_U4320 , P3_REG1_REG_15_ , P3_U3021 );
nand NAND2_8174 ( P3_U4321 , P3_REG2_REG_15_ , P3_U3020 );
nand NAND2_8175 ( P3_U4322 , P3_SUB_609_U21 , P3_U3019 );
not NOT1_8176 ( P3_U4323 , P3_U3073 );
nand NAND2_8177 ( P3_U4324 , P3_U3033 , P3_U3079 );
nand NAND2_8178 ( P3_U4325 , P3_R1110_U112 , P3_U3883 );
nand NAND2_8179 ( P3_U4326 , P3_R1077_U112 , P3_U3885 );
nand NAND2_8180 ( P3_U4327 , P3_R1095_U115 , P3_U3884 );
nand NAND2_8181 ( P3_U4328 , P3_R1143_U112 , P3_U3881 );
nand NAND2_8182 ( P3_U4329 , P3_R1161_U112 , P3_U3891 );
nand NAND2_8183 ( P3_U4330 , P3_R1131_U115 , P3_U3887 );
nand NAND2_8184 ( P3_U4331 , P3_R1200_U115 , P3_U3017 );
not NOT1_8185 ( P3_U4332 , P3_U3328 );
nand NAND2_8186 ( P3_U4333 , P3_R1179_U115 , P3_U3026 );
nand NAND2_8187 ( P3_U4334 , P3_U3025 , P3_U3073 );
nand NAND2_8188 ( P3_U4335 , P3_U3431 , P3_U4064 );
nand NAND2_8189 ( P3_U4336 , P3_U3638 , P3_U4332 );
nand NAND2_8190 ( P3_U4337 , P3_REG0_REG_16_ , P3_U3022 );
nand NAND2_8191 ( P3_U4338 , P3_REG1_REG_16_ , P3_U3021 );
nand NAND2_8192 ( P3_U4339 , P3_REG2_REG_16_ , P3_U3020 );
nand NAND2_8193 ( P3_U4340 , P3_SUB_609_U7 , P3_U3019 );
not NOT1_8194 ( P3_U4341 , P3_U3072 );
nand NAND2_8195 ( P3_U4342 , P3_U3033 , P3_U3078 );
nand NAND2_8196 ( P3_U4343 , P3_R1110_U111 , P3_U3883 );
nand NAND2_8197 ( P3_U4344 , P3_R1077_U111 , P3_U3885 );
nand NAND2_8198 ( P3_U4345 , P3_R1095_U114 , P3_U3884 );
nand NAND2_8199 ( P3_U4346 , P3_R1143_U111 , P3_U3881 );
nand NAND2_8200 ( P3_U4347 , P3_R1161_U111 , P3_U3891 );
nand NAND2_8201 ( P3_U4348 , P3_R1131_U114 , P3_U3887 );
nand NAND2_8202 ( P3_U4349 , P3_R1200_U114 , P3_U3017 );
not NOT1_8203 ( P3_U4350 , P3_U3329 );
nand NAND2_8204 ( P3_U4351 , P3_R1179_U114 , P3_U3026 );
nand NAND2_8205 ( P3_U4352 , P3_U3025 , P3_U3072 );
nand NAND2_8206 ( P3_U4353 , P3_U3434 , P3_U4064 );
nand NAND2_8207 ( P3_U4354 , P3_U3641 , P3_U4350 );
nand NAND2_8208 ( P3_U4355 , P3_REG0_REG_17_ , P3_U3022 );
nand NAND2_8209 ( P3_U4356 , P3_REG1_REG_17_ , P3_U3021 );
nand NAND2_8210 ( P3_U4357 , P3_REG2_REG_17_ , P3_U3020 );
nand NAND2_8211 ( P3_U4358 , P3_SUB_609_U19 , P3_U3019 );
not NOT1_8212 ( P3_U4359 , P3_U3068 );
nand NAND2_8213 ( P3_U4360 , P3_U3033 , P3_U3073 );
nand NAND2_8214 ( P3_U4361 , P3_R1110_U110 , P3_U3883 );
nand NAND2_8215 ( P3_U4362 , P3_R1077_U110 , P3_U3885 );
nand NAND2_8216 ( P3_U4363 , P3_R1095_U17 , P3_U3884 );
nand NAND2_8217 ( P3_U4364 , P3_R1143_U110 , P3_U3881 );
nand NAND2_8218 ( P3_U4365 , P3_R1161_U110 , P3_U3891 );
nand NAND2_8219 ( P3_U4366 , P3_R1131_U17 , P3_U3887 );
nand NAND2_8220 ( P3_U4367 , P3_R1200_U17 , P3_U3017 );
not NOT1_8221 ( P3_U4368 , P3_U3330 );
nand NAND2_8222 ( P3_U4369 , P3_R1179_U17 , P3_U3026 );
nand NAND2_8223 ( P3_U4370 , P3_U3025 , P3_U3068 );
nand NAND2_8224 ( P3_U4371 , P3_U3437 , P3_U4064 );
nand NAND2_8225 ( P3_U4372 , P3_U3644 , P3_U4368 );
nand NAND2_8226 ( P3_U4373 , P3_REG0_REG_18_ , P3_U3022 );
nand NAND2_8227 ( P3_U4374 , P3_REG1_REG_18_ , P3_U3021 );
nand NAND2_8228 ( P3_U4375 , P3_REG2_REG_18_ , P3_U3020 );
nand NAND2_8229 ( P3_U4376 , P3_SUB_609_U11 , P3_U3019 );
not NOT1_8230 ( P3_U4377 , P3_U3081 );
nand NAND2_8231 ( P3_U4378 , P3_U3033 , P3_U3072 );
nand NAND2_8232 ( P3_U4379 , P3_R1110_U12 , P3_U3883 );
nand NAND2_8233 ( P3_U4380 , P3_R1077_U12 , P3_U3885 );
nand NAND2_8234 ( P3_U4381 , P3_R1095_U103 , P3_U3884 );
nand NAND2_8235 ( P3_U4382 , P3_R1143_U12 , P3_U3881 );
nand NAND2_8236 ( P3_U4383 , P3_R1161_U12 , P3_U3891 );
nand NAND2_8237 ( P3_U4384 , P3_R1131_U103 , P3_U3887 );
nand NAND2_8238 ( P3_U4385 , P3_R1200_U103 , P3_U3017 );
not NOT1_8239 ( P3_U4386 , P3_U3331 );
nand NAND2_8240 ( P3_U4387 , P3_R1179_U103 , P3_U3026 );
nand NAND2_8241 ( P3_U4388 , P3_U3025 , P3_U3081 );
nand NAND2_8242 ( P3_U4389 , P3_U3440 , P3_U4064 );
nand NAND2_8243 ( P3_U4390 , P3_U3648 , P3_U4386 );
nand NAND2_8244 ( P3_U4391 , P3_REG0_REG_19_ , P3_U3022 );
nand NAND2_8245 ( P3_U4392 , P3_REG1_REG_19_ , P3_U3021 );
nand NAND2_8246 ( P3_U4393 , P3_REG2_REG_19_ , P3_U3020 );
nand NAND2_8247 ( P3_U4394 , P3_SUB_609_U15 , P3_U3019 );
not NOT1_8248 ( P3_U4395 , P3_U3080 );
nand NAND2_8249 ( P3_U4396 , P3_U3033 , P3_U3068 );
nand NAND2_8250 ( P3_U4397 , P3_R1110_U109 , P3_U3883 );
nand NAND2_8251 ( P3_U4398 , P3_R1077_U109 , P3_U3885 );
nand NAND2_8252 ( P3_U4399 , P3_R1095_U102 , P3_U3884 );
nand NAND2_8253 ( P3_U4400 , P3_R1143_U109 , P3_U3881 );
nand NAND2_8254 ( P3_U4401 , P3_R1161_U109 , P3_U3891 );
nand NAND2_8255 ( P3_U4402 , P3_R1131_U102 , P3_U3887 );
nand NAND2_8256 ( P3_U4403 , P3_R1200_U102 , P3_U3017 );
not NOT1_8257 ( P3_U4404 , P3_U3332 );
nand NAND2_8258 ( P3_U4405 , P3_R1179_U102 , P3_U3026 );
nand NAND2_8259 ( P3_U4406 , P3_U3025 , P3_U3080 );
nand NAND2_8260 ( P3_U4407 , P3_U3443 , P3_U4064 );
nand NAND2_8261 ( P3_U4408 , P3_U3651 , P3_U4404 );
nand NAND2_8262 ( P3_U4409 , P3_REG2_REG_20_ , P3_U3020 );
nand NAND2_8263 ( P3_U4410 , P3_REG1_REG_20_ , P3_U3021 );
nand NAND2_8264 ( P3_U4411 , P3_REG0_REG_20_ , P3_U3022 );
nand NAND2_8265 ( P3_U4412 , P3_SUB_609_U20 , P3_U3019 );
not NOT1_8266 ( P3_U4413 , P3_U3075 );
nand NAND2_8267 ( P3_U4414 , P3_U3033 , P3_U3081 );
nand NAND2_8268 ( P3_U4415 , P3_R1110_U108 , P3_U3883 );
nand NAND2_8269 ( P3_U4416 , P3_R1077_U108 , P3_U3885 );
nand NAND2_8270 ( P3_U4417 , P3_R1095_U101 , P3_U3884 );
nand NAND2_8271 ( P3_U4418 , P3_R1143_U108 , P3_U3881 );
nand NAND2_8272 ( P3_U4419 , P3_R1161_U108 , P3_U3891 );
nand NAND2_8273 ( P3_U4420 , P3_R1131_U101 , P3_U3887 );
nand NAND2_8274 ( P3_U4421 , P3_R1200_U101 , P3_U3017 );
not NOT1_8275 ( P3_U4422 , P3_U3333 );
nand NAND2_8276 ( P3_U4423 , P3_R1179_U101 , P3_U3026 );
nand NAND2_8277 ( P3_U4424 , P3_U3025 , P3_U3075 );
nand NAND2_8278 ( P3_U4425 , P3_U3445 , P3_U4064 );
nand NAND2_8279 ( P3_U4426 , P3_U3654 , P3_U4422 );
nand NAND2_8280 ( P3_U4427 , P3_REG2_REG_21_ , P3_U3020 );
nand NAND2_8281 ( P3_U4428 , P3_REG1_REG_21_ , P3_U3021 );
nand NAND2_8282 ( P3_U4429 , P3_REG0_REG_21_ , P3_U3022 );
nand NAND2_8283 ( P3_U4430 , P3_SUB_609_U27 , P3_U3019 );
not NOT1_8284 ( P3_U4431 , P3_U3074 );
nand NAND2_8285 ( P3_U4432 , P3_U3033 , P3_U3080 );
nand NAND2_8286 ( P3_U4433 , P3_R1110_U13 , P3_U3883 );
nand NAND2_8287 ( P3_U4434 , P3_R1077_U13 , P3_U3885 );
nand NAND2_8288 ( P3_U4435 , P3_R1095_U99 , P3_U3884 );
nand NAND2_8289 ( P3_U4436 , P3_R1143_U13 , P3_U3881 );
nand NAND2_8290 ( P3_U4437 , P3_R1161_U13 , P3_U3891 );
nand NAND2_8291 ( P3_U4438 , P3_R1131_U99 , P3_U3887 );
nand NAND2_8292 ( P3_U4439 , P3_R1200_U99 , P3_U3017 );
not NOT1_8293 ( P3_U4440 , P3_U3335 );
nand NAND2_8294 ( P3_U4441 , P3_R1179_U99 , P3_U3026 );
nand NAND2_8295 ( P3_U4442 , P3_U3025 , P3_U3074 );
nand NAND2_8296 ( P3_U4443 , P3_U3907 , P3_U4064 );
nand NAND2_8297 ( P3_U4444 , P3_U3657 , P3_U4440 );
nand NAND2_8298 ( P3_U4445 , P3_REG2_REG_22_ , P3_U3020 );
nand NAND2_8299 ( P3_U4446 , P3_REG1_REG_22_ , P3_U3021 );
nand NAND2_8300 ( P3_U4447 , P3_REG0_REG_22_ , P3_U3022 );
nand NAND2_8301 ( P3_U4448 , P3_SUB_609_U17 , P3_U3019 );
not NOT1_8302 ( P3_U4449 , P3_U3060 );
nand NAND2_8303 ( P3_U4450 , P3_U3033 , P3_U3075 );
nand NAND2_8304 ( P3_U4451 , P3_R1110_U14 , P3_U3883 );
nand NAND2_8305 ( P3_U4452 , P3_R1077_U14 , P3_U3885 );
nand NAND2_8306 ( P3_U4453 , P3_R1095_U113 , P3_U3884 );
nand NAND2_8307 ( P3_U4454 , P3_R1143_U14 , P3_U3881 );
nand NAND2_8308 ( P3_U4455 , P3_R1161_U14 , P3_U3891 );
nand NAND2_8309 ( P3_U4456 , P3_R1131_U113 , P3_U3887 );
nand NAND2_8310 ( P3_U4457 , P3_R1200_U113 , P3_U3017 );
not NOT1_8311 ( P3_U4458 , P3_U3337 );
nand NAND2_8312 ( P3_U4459 , P3_R1179_U113 , P3_U3026 );
nand NAND2_8313 ( P3_U4460 , P3_U3025 , P3_U3060 );
nand NAND2_8314 ( P3_U4461 , P3_U3906 , P3_U4064 );
nand NAND2_8315 ( P3_U4462 , P3_U3660 , P3_U4458 );
nand NAND2_8316 ( P3_U4463 , P3_REG2_REG_23_ , P3_U3020 );
nand NAND2_8317 ( P3_U4464 , P3_REG1_REG_23_ , P3_U3021 );
nand NAND2_8318 ( P3_U4465 , P3_REG0_REG_23_ , P3_U3022 );
nand NAND2_8319 ( P3_U4466 , P3_SUB_609_U6 , P3_U3019 );
not NOT1_8320 ( P3_U4467 , P3_U3065 );
nand NAND2_8321 ( P3_U4468 , P3_U3033 , P3_U3074 );
nand NAND2_8322 ( P3_U4469 , P3_R1110_U107 , P3_U3883 );
nand NAND2_8323 ( P3_U4470 , P3_R1077_U107 , P3_U3885 );
nand NAND2_8324 ( P3_U4471 , P3_R1095_U112 , P3_U3884 );
nand NAND2_8325 ( P3_U4472 , P3_R1143_U107 , P3_U3881 );
nand NAND2_8326 ( P3_U4473 , P3_R1161_U107 , P3_U3891 );
nand NAND2_8327 ( P3_U4474 , P3_R1131_U112 , P3_U3887 );
nand NAND2_8328 ( P3_U4475 , P3_R1200_U112 , P3_U3017 );
not NOT1_8329 ( P3_U4476 , P3_U3339 );
nand NAND2_8330 ( P3_U4477 , P3_R1179_U112 , P3_U3026 );
nand NAND2_8331 ( P3_U4478 , P3_U3025 , P3_U3065 );
nand NAND2_8332 ( P3_U4479 , P3_U3905 , P3_U4064 );
nand NAND2_8333 ( P3_U4480 , P3_U3663 , P3_U4476 );
nand NAND2_8334 ( P3_U4481 , P3_REG2_REG_24_ , P3_U3020 );
nand NAND2_8335 ( P3_U4482 , P3_REG1_REG_24_ , P3_U3021 );
nand NAND2_8336 ( P3_U4483 , P3_REG0_REG_24_ , P3_U3022 );
nand NAND2_8337 ( P3_U4484 , P3_SUB_609_U10 , P3_U3019 );
not NOT1_8338 ( P3_U4485 , P3_U3064 );
nand NAND2_8339 ( P3_U4486 , P3_U3033 , P3_U3060 );
nand NAND2_8340 ( P3_U4487 , P3_R1110_U106 , P3_U3883 );
nand NAND2_8341 ( P3_U4488 , P3_R1077_U106 , P3_U3885 );
nand NAND2_8342 ( P3_U4489 , P3_R1095_U18 , P3_U3884 );
nand NAND2_8343 ( P3_U4490 , P3_R1143_U106 , P3_U3881 );
nand NAND2_8344 ( P3_U4491 , P3_R1161_U106 , P3_U3891 );
nand NAND2_8345 ( P3_U4492 , P3_R1131_U18 , P3_U3887 );
nand NAND2_8346 ( P3_U4493 , P3_R1200_U18 , P3_U3017 );
not NOT1_8347 ( P3_U4494 , P3_U3341 );
nand NAND2_8348 ( P3_U4495 , P3_R1179_U18 , P3_U3026 );
nand NAND2_8349 ( P3_U4496 , P3_U3025 , P3_U3064 );
nand NAND2_8350 ( P3_U4497 , P3_U3904 , P3_U4064 );
nand NAND2_8351 ( P3_U4498 , P3_U3666 , P3_U4494 );
nand NAND2_8352 ( P3_U4499 , P3_REG2_REG_25_ , P3_U3020 );
nand NAND2_8353 ( P3_U4500 , P3_REG1_REG_25_ , P3_U3021 );
nand NAND2_8354 ( P3_U4501 , P3_REG0_REG_25_ , P3_U3022 );
nand NAND2_8355 ( P3_U4502 , P3_SUB_609_U16 , P3_U3019 );
not NOT1_8356 ( P3_U4503 , P3_U3057 );
nand NAND2_8357 ( P3_U4504 , P3_U3033 , P3_U3065 );
nand NAND2_8358 ( P3_U4505 , P3_R1110_U105 , P3_U3883 );
nand NAND2_8359 ( P3_U4506 , P3_R1077_U105 , P3_U3885 );
nand NAND2_8360 ( P3_U4507 , P3_R1095_U98 , P3_U3884 );
nand NAND2_8361 ( P3_U4508 , P3_R1143_U105 , P3_U3881 );
nand NAND2_8362 ( P3_U4509 , P3_R1161_U105 , P3_U3891 );
nand NAND2_8363 ( P3_U4510 , P3_R1131_U98 , P3_U3887 );
nand NAND2_8364 ( P3_U4511 , P3_R1200_U98 , P3_U3017 );
not NOT1_8365 ( P3_U4512 , P3_U3343 );
nand NAND2_8366 ( P3_U4513 , P3_R1179_U98 , P3_U3026 );
nand NAND2_8367 ( P3_U4514 , P3_U3025 , P3_U3057 );
nand NAND2_8368 ( P3_U4515 , P3_U3903 , P3_U4064 );
nand NAND2_8369 ( P3_U4516 , P3_U3670 , P3_U4512 );
nand NAND2_8370 ( P3_U4517 , P3_REG2_REG_26_ , P3_U3020 );
nand NAND2_8371 ( P3_U4518 , P3_REG1_REG_26_ , P3_U3021 );
nand NAND2_8372 ( P3_U4519 , P3_REG0_REG_26_ , P3_U3022 );
nand NAND2_8373 ( P3_U4520 , P3_SUB_609_U26 , P3_U3019 );
not NOT1_8374 ( P3_U4521 , P3_U3056 );
nand NAND2_8375 ( P3_U4522 , P3_U3033 , P3_U3064 );
nand NAND2_8376 ( P3_U4523 , P3_R1110_U104 , P3_U3883 );
nand NAND2_8377 ( P3_U4524 , P3_R1077_U104 , P3_U3885 );
nand NAND2_8378 ( P3_U4525 , P3_R1095_U97 , P3_U3884 );
nand NAND2_8379 ( P3_U4526 , P3_R1143_U104 , P3_U3881 );
nand NAND2_8380 ( P3_U4527 , P3_R1161_U104 , P3_U3891 );
nand NAND2_8381 ( P3_U4528 , P3_R1131_U97 , P3_U3887 );
nand NAND2_8382 ( P3_U4529 , P3_R1200_U97 , P3_U3017 );
not NOT1_8383 ( P3_U4530 , P3_U3345 );
nand NAND2_8384 ( P3_U4531 , P3_R1179_U97 , P3_U3026 );
nand NAND2_8385 ( P3_U4532 , P3_U3025 , P3_U3056 );
nand NAND2_8386 ( P3_U4533 , P3_U3902 , P3_U4064 );
nand NAND2_8387 ( P3_U4534 , P3_U3674 , P3_U4530 );
nand NAND2_8388 ( P3_U4535 , P3_REG2_REG_27_ , P3_U3020 );
nand NAND2_8389 ( P3_U4536 , P3_REG1_REG_27_ , P3_U3021 );
nand NAND2_8390 ( P3_U4537 , P3_REG0_REG_27_ , P3_U3022 );
nand NAND2_8391 ( P3_U4538 , P3_SUB_609_U22 , P3_U3019 );
not NOT1_8392 ( P3_U4539 , P3_U3052 );
nand NAND2_8393 ( P3_U4540 , P3_U3033 , P3_U3057 );
nand NAND2_8394 ( P3_U4541 , P3_R1110_U15 , P3_U3883 );
nand NAND2_8395 ( P3_U4542 , P3_R1077_U15 , P3_U3885 );
nand NAND2_8396 ( P3_U4543 , P3_R1095_U111 , P3_U3884 );
nand NAND2_8397 ( P3_U4544 , P3_R1143_U15 , P3_U3881 );
nand NAND2_8398 ( P3_U4545 , P3_R1161_U15 , P3_U3891 );
nand NAND2_8399 ( P3_U4546 , P3_R1131_U111 , P3_U3887 );
nand NAND2_8400 ( P3_U4547 , P3_R1200_U111 , P3_U3017 );
not NOT1_8401 ( P3_U4548 , P3_U3347 );
nand NAND2_8402 ( P3_U4549 , P3_R1179_U111 , P3_U3026 );
nand NAND2_8403 ( P3_U4550 , P3_U3025 , P3_U3052 );
nand NAND2_8404 ( P3_U4551 , P3_U3901 , P3_U4064 );
nand NAND2_8405 ( P3_U4552 , P3_U3678 , P3_U4548 );
nand NAND2_8406 ( P3_U4553 , P3_REG2_REG_28_ , P3_U3020 );
nand NAND2_8407 ( P3_U4554 , P3_REG1_REG_28_ , P3_U3021 );
nand NAND2_8408 ( P3_U4555 , P3_REG0_REG_28_ , P3_U3022 );
nand NAND2_8409 ( P3_U4556 , P3_SUB_609_U28 , P3_U3019 );
not NOT1_8410 ( P3_U4557 , P3_U3053 );
nand NAND2_8411 ( P3_U4558 , P3_U3033 , P3_U3056 );
nand NAND2_8412 ( P3_U4559 , P3_R1110_U103 , P3_U3883 );
nand NAND2_8413 ( P3_U4560 , P3_R1077_U103 , P3_U3885 );
nand NAND2_8414 ( P3_U4561 , P3_R1095_U19 , P3_U3884 );
nand NAND2_8415 ( P3_U4562 , P3_R1143_U103 , P3_U3881 );
nand NAND2_8416 ( P3_U4563 , P3_R1161_U103 , P3_U3891 );
nand NAND2_8417 ( P3_U4564 , P3_R1131_U19 , P3_U3887 );
nand NAND2_8418 ( P3_U4565 , P3_R1200_U19 , P3_U3017 );
not NOT1_8419 ( P3_U4566 , P3_U3349 );
nand NAND2_8420 ( P3_U4567 , P3_R1179_U19 , P3_U3026 );
nand NAND2_8421 ( P3_U4568 , P3_U3025 , P3_U3053 );
nand NAND2_8422 ( P3_U4569 , P3_U3900 , P3_U4064 );
nand NAND2_8423 ( P3_U4570 , P3_U3682 , P3_U4566 );
nand NAND2_8424 ( P3_U4571 , P3_SUB_609_U92 , P3_U3019 );
nand NAND2_8425 ( P3_U4572 , P3_REG2_REG_29_ , P3_U3020 );
nand NAND2_8426 ( P3_U4573 , P3_REG1_REG_29_ , P3_U3021 );
nand NAND2_8427 ( P3_U4574 , P3_REG0_REG_29_ , P3_U3022 );
not NOT1_8428 ( P3_U4575 , P3_U3054 );
nand NAND2_8429 ( P3_U4576 , P3_U3033 , P3_U3052 );
nand NAND2_8430 ( P3_U4577 , P3_R1110_U102 , P3_U3883 );
nand NAND2_8431 ( P3_U4578 , P3_R1077_U102 , P3_U3885 );
nand NAND2_8432 ( P3_U4579 , P3_R1095_U96 , P3_U3884 );
nand NAND2_8433 ( P3_U4580 , P3_R1143_U102 , P3_U3881 );
nand NAND2_8434 ( P3_U4581 , P3_R1161_U102 , P3_U3891 );
nand NAND2_8435 ( P3_U4582 , P3_R1131_U96 , P3_U3887 );
nand NAND2_8436 ( P3_U4583 , P3_R1200_U96 , P3_U3017 );
not NOT1_8437 ( P3_U4584 , P3_U3351 );
nand NAND2_8438 ( P3_U4585 , P3_R1179_U96 , P3_U3026 );
nand NAND2_8439 ( P3_U4586 , P3_U3025 , P3_U3054 );
nand NAND2_8440 ( P3_U4587 , P3_U3899 , P3_U4064 );
nand NAND2_8441 ( P3_U4588 , P3_U3686 , P3_U4584 );
nand NAND2_8442 ( P3_U4589 , P3_REG2_REG_30_ , P3_U3020 );
nand NAND2_8443 ( P3_U4590 , P3_REG1_REG_30_ , P3_U3021 );
nand NAND2_8444 ( P3_U4591 , P3_REG0_REG_30_ , P3_U3022 );
nand NAND2_8445 ( P3_U4592 , P3_SUB_609_U92 , P3_U3019 );
not NOT1_8446 ( P3_U4593 , P3_U3058 );
nand NAND2_8447 ( P3_U4594 , P3_U3892 , P3_U3298 );
nand NAND2_8448 ( P3_U4595 , P3_U3833 , P3_U4594 );
nand NAND3_8449 ( P3_U4596 , P3_U4595 , P3_U3911 , P3_U3058 );
nand NAND2_8450 ( P3_U4597 , P3_U3033 , P3_U3053 );
nand NAND2_8451 ( P3_U4598 , P3_R1110_U101 , P3_U3883 );
nand NAND2_8452 ( P3_U4599 , P3_R1077_U101 , P3_U3885 );
nand NAND2_8453 ( P3_U4600 , P3_R1095_U20 , P3_U3884 );
nand NAND2_8454 ( P3_U4601 , P3_R1143_U101 , P3_U3881 );
nand NAND2_8455 ( P3_U4602 , P3_R1161_U101 , P3_U3891 );
nand NAND2_8456 ( P3_U4603 , P3_R1131_U20 , P3_U3887 );
nand NAND2_8457 ( P3_U4604 , P3_R1200_U20 , P3_U3017 );
not NOT1_8458 ( P3_U4605 , P3_U3354 );
nand NAND2_8459 ( P3_U4606 , P3_R1179_U20 , P3_U3026 );
nand NAND2_8460 ( P3_U4607 , P3_U3908 , P3_U4064 );
nand NAND2_8461 ( P3_U4608 , P3_U3690 , P3_U4605 );
nand NAND2_8462 ( P3_U4609 , P3_SUB_609_U92 , P3_U3019 );
nand NAND2_8463 ( P3_U4610 , P3_REG2_REG_31_ , P3_U3020 );
nand NAND2_8464 ( P3_U4611 , P3_REG1_REG_31_ , P3_U3021 );
nand NAND2_8465 ( P3_U4612 , P3_REG0_REG_31_ , P3_U3022 );
not NOT1_8466 ( P3_U4613 , P3_U3055 );
nand NAND2_8467 ( P3_U4614 , P3_U3873 , P3_U4064 );
nand NAND2_8468 ( P3_U4615 , P3_U3361 , P3_U4614 );
nand NAND2_8469 ( P3_U4616 , P3_U3872 , P3_U4064 );
nand NAND2_8470 ( P3_U4617 , P3_U3361 , P3_U4616 );
nand NAND3_8471 ( P3_U4618 , P3_U5641 , P3_U5640 , P3_U3302 );
nand NAND2_8472 ( P3_U4619 , P3_U3888 , P3_U3367 );
nand NAND2_8473 ( P3_U4620 , P3_U3048 , P3_U4619 );
nand NAND2_8474 ( P3_U4621 , P3_U3047 , P3_U4618 );
nand NAND2_8475 ( P3_U4622 , P3_U4621 , P3_U4620 );
nand NAND2_8476 ( P3_U4623 , P3_U5456 , P3_U3379 );
nand NAND3_8477 ( P3_U4624 , P3_U4623 , P3_U3380 , P3_U3834 );
nand NAND2_8478 ( P3_U4625 , P3_U3048 , P3_U4624 );
nand NAND2_8479 ( P3_U4626 , P3_U3047 , P3_U4619 );
nand NAND3_8480 ( P3_U4627 , P3_U4625 , P3_U3360 , P3_U4626 );
not NOT1_8481 ( P3_U4628 , P3_U3365 );
nand NAND2_8482 ( P3_U4629 , P3_U3034 , P3_U3077 );
nand NAND2_8483 ( P3_U4630 , P3_U3030 , P3_R1179_U24 );
nand NAND2_8484 ( P3_U4631 , P3_U3029 , P3_U3387 );
nand NAND2_8485 ( P3_U4632 , P3_U3028 , P3_REG3_REG_0_ );
nand NAND2_8486 ( P3_U4633 , P3_U3034 , P3_U3067 );
nand NAND2_8487 ( P3_U4634 , P3_U3030 , P3_R1179_U100 );
nand NAND2_8488 ( P3_U4635 , P3_U3029 , P3_U3392 );
nand NAND2_8489 ( P3_U4636 , P3_U3028 , P3_REG3_REG_1_ );
nand NAND2_8490 ( P3_U4637 , P3_U3034 , P3_U3063 );
nand NAND2_8491 ( P3_U4638 , P3_U3030 , P3_R1179_U110 );
nand NAND2_8492 ( P3_U4639 , P3_U3029 , P3_U3395 );
nand NAND2_8493 ( P3_U4640 , P3_U3028 , P3_REG3_REG_2_ );
nand NAND2_8494 ( P3_U4641 , P3_U3034 , P3_U3059 );
nand NAND2_8495 ( P3_U4642 , P3_U3030 , P3_R1179_U21 );
nand NAND2_8496 ( P3_U4643 , P3_U3029 , P3_U3398 );
nand NAND2_8497 ( P3_U4644 , P3_U3028 , P3_SUB_609_U25 );
nand NAND2_8498 ( P3_U4645 , P3_U3034 , P3_U3066 );
nand NAND2_8499 ( P3_U4646 , P3_U3030 , P3_R1179_U109 );
nand NAND2_8500 ( P3_U4647 , P3_U3029 , P3_U3401 );
nand NAND2_8501 ( P3_U4648 , P3_U3028 , P3_SUB_609_U29 );
nand NAND2_8502 ( P3_U4649 , P3_U3034 , P3_U3070 );
nand NAND2_8503 ( P3_U4650 , P3_U3030 , P3_R1179_U108 );
nand NAND2_8504 ( P3_U4651 , P3_U3029 , P3_U3404 );
nand NAND2_8505 ( P3_U4652 , P3_U3028 , P3_SUB_609_U53 );
nand NAND2_8506 ( P3_U4653 , P3_U3034 , P3_U3069 );
nand NAND2_8507 ( P3_U4654 , P3_U3030 , P3_R1179_U22 );
nand NAND2_8508 ( P3_U4655 , P3_U3029 , P3_U3407 );
nand NAND2_8509 ( P3_U4656 , P3_U3028 , P3_SUB_609_U8 );
nand NAND2_8510 ( P3_U4657 , P3_U3034 , P3_U3083 );
nand NAND2_8511 ( P3_U4658 , P3_U3030 , P3_R1179_U107 );
nand NAND2_8512 ( P3_U4659 , P3_U3029 , P3_U3410 );
nand NAND2_8513 ( P3_U4660 , P3_U3028 , P3_SUB_609_U18 );
nand NAND2_8514 ( P3_U4661 , P3_U3034 , P3_U3082 );
nand NAND2_8515 ( P3_U4662 , P3_U3030 , P3_R1179_U23 );
nand NAND2_8516 ( P3_U4663 , P3_U3029 , P3_U3413 );
nand NAND2_8517 ( P3_U4664 , P3_U3028 , P3_SUB_609_U12 );
nand NAND2_8518 ( P3_U4665 , P3_U3034 , P3_U3061 );
nand NAND2_8519 ( P3_U4666 , P3_U3030 , P3_R1179_U106 );
nand NAND2_8520 ( P3_U4667 , P3_U3029 , P3_U3416 );
nand NAND2_8521 ( P3_U4668 , P3_U3028 , P3_SUB_609_U14 );
nand NAND2_8522 ( P3_U4669 , P3_U3034 , P3_U3062 );
nand NAND2_8523 ( P3_U4670 , P3_U3030 , P3_R1179_U116 );
nand NAND2_8524 ( P3_U4671 , P3_U3029 , P3_U3419 );
nand NAND2_8525 ( P3_U4672 , P3_U3028 , P3_SUB_609_U13 );
nand NAND2_8526 ( P3_U4673 , P3_U3034 , P3_U3071 );
nand NAND2_8527 ( P3_U4674 , P3_U3030 , P3_R1179_U16 );
nand NAND2_8528 ( P3_U4675 , P3_U3029 , P3_U3422 );
nand NAND2_8529 ( P3_U4676 , P3_U3028 , P3_SUB_609_U9 );
nand NAND2_8530 ( P3_U4677 , P3_U3034 , P3_U3079 );
nand NAND2_8531 ( P3_U4678 , P3_U3030 , P3_R1179_U105 );
nand NAND2_8532 ( P3_U4679 , P3_U3029 , P3_U3425 );
nand NAND2_8533 ( P3_U4680 , P3_U3028 , P3_SUB_609_U23 );
nand NAND2_8534 ( P3_U4681 , P3_U3034 , P3_U3078 );
nand NAND2_8535 ( P3_U4682 , P3_U3030 , P3_R1179_U104 );
nand NAND2_8536 ( P3_U4683 , P3_U3029 , P3_U3428 );
nand NAND2_8537 ( P3_U4684 , P3_U3028 , P3_SUB_609_U24 );
nand NAND2_8538 ( P3_U4685 , P3_U3034 , P3_U3073 );
nand NAND2_8539 ( P3_U4686 , P3_U3030 , P3_R1179_U115 );
nand NAND2_8540 ( P3_U4687 , P3_U3029 , P3_U3431 );
nand NAND2_8541 ( P3_U4688 , P3_U3028 , P3_SUB_609_U30 );
nand NAND2_8542 ( P3_U4689 , P3_U3034 , P3_U3072 );
nand NAND2_8543 ( P3_U4690 , P3_U3030 , P3_R1179_U114 );
nand NAND2_8544 ( P3_U4691 , P3_U3029 , P3_U3434 );
nand NAND2_8545 ( P3_U4692 , P3_U3028 , P3_SUB_609_U21 );
nand NAND2_8546 ( P3_U4693 , P3_U3034 , P3_U3068 );
nand NAND2_8547 ( P3_U4694 , P3_U3030 , P3_R1179_U17 );
nand NAND2_8548 ( P3_U4695 , P3_U3029 , P3_U3437 );
nand NAND2_8549 ( P3_U4696 , P3_U3028 , P3_SUB_609_U7 );
nand NAND2_8550 ( P3_U4697 , P3_U3034 , P3_U3081 );
nand NAND2_8551 ( P3_U4698 , P3_U3030 , P3_R1179_U103 );
nand NAND2_8552 ( P3_U4699 , P3_U3029 , P3_U3440 );
nand NAND2_8553 ( P3_U4700 , P3_U3028 , P3_SUB_609_U19 );
nand NAND2_8554 ( P3_U4701 , P3_U3034 , P3_U3080 );
nand NAND2_8555 ( P3_U4702 , P3_U3030 , P3_R1179_U102 );
nand NAND2_8556 ( P3_U4703 , P3_U3029 , P3_U3443 );
nand NAND2_8557 ( P3_U4704 , P3_U3028 , P3_SUB_609_U11 );
nand NAND2_8558 ( P3_U4705 , P3_U3034 , P3_U3075 );
nand NAND2_8559 ( P3_U4706 , P3_U3030 , P3_R1179_U101 );
nand NAND2_8560 ( P3_U4707 , P3_U3029 , P3_U3445 );
nand NAND2_8561 ( P3_U4708 , P3_U3028 , P3_SUB_609_U15 );
nand NAND2_8562 ( P3_U4709 , P3_U3034 , P3_U3074 );
nand NAND2_8563 ( P3_U4710 , P3_U3030 , P3_R1179_U99 );
nand NAND2_8564 ( P3_U4711 , P3_U3029 , P3_U3907 );
nand NAND2_8565 ( P3_U4712 , P3_U3028 , P3_SUB_609_U20 );
nand NAND2_8566 ( P3_U4713 , P3_U3034 , P3_U3060 );
nand NAND2_8567 ( P3_U4714 , P3_U3030 , P3_R1179_U113 );
nand NAND2_8568 ( P3_U4715 , P3_U3029 , P3_U3906 );
nand NAND2_8569 ( P3_U4716 , P3_U3028 , P3_SUB_609_U27 );
nand NAND2_8570 ( P3_U4717 , P3_U3034 , P3_U3065 );
nand NAND2_8571 ( P3_U4718 , P3_U3030 , P3_R1179_U112 );
nand NAND2_8572 ( P3_U4719 , P3_U3029 , P3_U3905 );
nand NAND2_8573 ( P3_U4720 , P3_U3028 , P3_SUB_609_U17 );
nand NAND2_8574 ( P3_U4721 , P3_U3034 , P3_U3064 );
nand NAND2_8575 ( P3_U4722 , P3_U3030 , P3_R1179_U18 );
nand NAND2_8576 ( P3_U4723 , P3_U3029 , P3_U3904 );
nand NAND2_8577 ( P3_U4724 , P3_U3028 , P3_SUB_609_U6 );
nand NAND2_8578 ( P3_U4725 , P3_U3034 , P3_U3057 );
nand NAND2_8579 ( P3_U4726 , P3_U3030 , P3_R1179_U98 );
nand NAND2_8580 ( P3_U4727 , P3_U3029 , P3_U3903 );
nand NAND2_8581 ( P3_U4728 , P3_U3028 , P3_SUB_609_U10 );
nand NAND2_8582 ( P3_U4729 , P3_U3034 , P3_U3056 );
nand NAND2_8583 ( P3_U4730 , P3_U3030 , P3_R1179_U97 );
nand NAND2_8584 ( P3_U4731 , P3_U3029 , P3_U3902 );
nand NAND2_8585 ( P3_U4732 , P3_U3028 , P3_SUB_609_U16 );
nand NAND2_8586 ( P3_U4733 , P3_U3034 , P3_U3052 );
nand NAND2_8587 ( P3_U4734 , P3_U3030 , P3_R1179_U111 );
nand NAND2_8588 ( P3_U4735 , P3_U3029 , P3_U3901 );
nand NAND2_8589 ( P3_U4736 , P3_U3028 , P3_SUB_609_U26 );
nand NAND2_8590 ( P3_U4737 , P3_U3034 , P3_U3053 );
nand NAND2_8591 ( P3_U4738 , P3_U3030 , P3_R1179_U19 );
nand NAND2_8592 ( P3_U4739 , P3_U3029 , P3_U3900 );
nand NAND2_8593 ( P3_U4740 , P3_U3028 , P3_SUB_609_U22 );
nand NAND2_8594 ( P3_U4741 , P3_U3034 , P3_U3054 );
nand NAND2_8595 ( P3_U4742 , P3_U3030 , P3_R1179_U96 );
nand NAND2_8596 ( P3_U4743 , P3_U3029 , P3_U3899 );
nand NAND2_8597 ( P3_U4744 , P3_U3028 , P3_SUB_609_U28 );
nand NAND2_8598 ( P3_U4745 , P3_U3030 , P3_R1179_U20 );
nand NAND2_8599 ( P3_U4746 , P3_U3029 , P3_U3908 );
nand NAND2_8600 ( P3_U4747 , P3_U3028 , P3_SUB_609_U92 );
nand NAND2_8601 ( P3_U4748 , P3_U3028 , P3_SUB_609_U92 );
nand NAND2_8602 ( P3_U4749 , P3_U3916 , P3_U3912 );
nand NAND2_8603 ( P3_U4750 , P3_U3029 , P3_U3873 );
nand NAND2_8604 ( P3_U4751 , P3_REG2_REG_30_ , P3_U3358 );
nand NAND2_8605 ( P3_U4752 , P3_U3029 , P3_U3872 );
nand NAND2_8606 ( P3_U4753 , P3_REG2_REG_31_ , P3_U3358 );
nand NAND4_8607 ( P3_U4754 , P3_U4628 , P3_U3359 , P3_U3698 , P3_U3697 );
nand NAND2_8608 ( P3_U4755 , P3_R1212_U6 , P3_U3040 );
nand NAND2_8609 ( P3_U4756 , P3_U3039 , P3_U3379 );
nand NAND2_8610 ( P3_U4757 , P3_R1209_U6 , P3_U3037 );
nand NAND3_8611 ( P3_U4758 , P3_U4756 , P3_U4755 , P3_U4757 );
nand NAND2_8612 ( P3_U4759 , P3_U3910 , P3_U5440 );
not NOT1_8613 ( P3_U4760 , P3_U3366 );
nand NAND2_8614 ( P3_U4761 , P3_U3833 , P3_U3896 );
nand NAND2_8615 ( P3_U4762 , P3_R1054_U67 , P3_U3051 );
nand NAND2_8616 ( P3_U4763 , P3_U5768 , P3_U3379 );
nand NAND2_8617 ( P3_U4764 , P3_U3042 , P3_U4758 );
nand NAND2_8618 ( P3_U4765 , P3_U3041 , P3_R1212_U6 );
nand NAND2_8619 ( P3_U4766 , P3_REG3_REG_19_ , P3_U3151 );
nand NAND2_8620 ( P3_U4767 , P3_U3038 , P3_R1209_U6 );
nand NAND2_8621 ( P3_U4768 , P3_ADDR_REG_19_ , P3_U4760 );
nand NAND2_8622 ( P3_U4769 , P3_R1212_U58 , P3_U3040 );
nand NAND2_8623 ( P3_U4770 , P3_U3039 , P3_U3442 );
nand NAND2_8624 ( P3_U4771 , P3_R1209_U58 , P3_U3037 );
nand NAND3_8625 ( P3_U4772 , P3_U4770 , P3_U4769 , P3_U4771 );
nand NAND2_8626 ( P3_U4773 , P3_R1054_U68 , P3_U3051 );
nand NAND2_8627 ( P3_U4774 , P3_U5768 , P3_U3442 );
nand NAND2_8628 ( P3_U4775 , P3_U3042 , P3_U4772 );
nand NAND2_8629 ( P3_U4776 , P3_R1212_U58 , P3_U3041 );
nand NAND2_8630 ( P3_U4777 , P3_REG3_REG_18_ , P3_U3151 );
nand NAND2_8631 ( P3_U4778 , P3_R1209_U58 , P3_U3038 );
nand NAND2_8632 ( P3_U4779 , P3_ADDR_REG_18_ , P3_U4760 );
nand NAND2_8633 ( P3_U4780 , P3_R1212_U59 , P3_U3040 );
nand NAND2_8634 ( P3_U4781 , P3_U3039 , P3_U3439 );
nand NAND2_8635 ( P3_U4782 , P3_R1209_U59 , P3_U3037 );
nand NAND3_8636 ( P3_U4783 , P3_U4781 , P3_U4780 , P3_U4782 );
nand NAND2_8637 ( P3_U4784 , P3_R1054_U69 , P3_U3051 );
nand NAND2_8638 ( P3_U4785 , P3_U5768 , P3_U3439 );
nand NAND2_8639 ( P3_U4786 , P3_U3042 , P3_U4783 );
nand NAND2_8640 ( P3_U4787 , P3_R1212_U59 , P3_U3041 );
nand NAND2_8641 ( P3_U4788 , P3_REG3_REG_17_ , P3_U3151 );
nand NAND2_8642 ( P3_U4789 , P3_R1209_U59 , P3_U3038 );
nand NAND2_8643 ( P3_U4790 , P3_ADDR_REG_17_ , P3_U4760 );
nand NAND2_8644 ( P3_U4791 , P3_R1212_U60 , P3_U3040 );
nand NAND2_8645 ( P3_U4792 , P3_U3039 , P3_U3436 );
nand NAND2_8646 ( P3_U4793 , P3_R1209_U60 , P3_U3037 );
nand NAND3_8647 ( P3_U4794 , P3_U4792 , P3_U4791 , P3_U4793 );
nand NAND2_8648 ( P3_U4795 , P3_R1054_U13 , P3_U3051 );
nand NAND2_8649 ( P3_U4796 , P3_U5768 , P3_U3436 );
nand NAND2_8650 ( P3_U4797 , P3_U3042 , P3_U4794 );
nand NAND2_8651 ( P3_U4798 , P3_R1212_U60 , P3_U3041 );
nand NAND2_8652 ( P3_U4799 , P3_REG3_REG_16_ , P3_U3151 );
nand NAND2_8653 ( P3_U4800 , P3_R1209_U60 , P3_U3038 );
nand NAND2_8654 ( P3_U4801 , P3_ADDR_REG_16_ , P3_U4760 );
nand NAND2_8655 ( P3_U4802 , P3_R1212_U61 , P3_U3040 );
nand NAND2_8656 ( P3_U4803 , P3_U3039 , P3_U3433 );
nand NAND2_8657 ( P3_U4804 , P3_R1209_U61 , P3_U3037 );
nand NAND3_8658 ( P3_U4805 , P3_U4803 , P3_U4802 , P3_U4804 );
nand NAND2_8659 ( P3_U4806 , P3_R1054_U77 , P3_U3051 );
nand NAND2_8660 ( P3_U4807 , P3_U5768 , P3_U3433 );
nand NAND2_8661 ( P3_U4808 , P3_U3042 , P3_U4805 );
nand NAND2_8662 ( P3_U4809 , P3_R1212_U61 , P3_U3041 );
nand NAND2_8663 ( P3_U4810 , P3_REG3_REG_15_ , P3_U3151 );
nand NAND2_8664 ( P3_U4811 , P3_R1209_U61 , P3_U3038 );
nand NAND2_8665 ( P3_U4812 , P3_ADDR_REG_15_ , P3_U4760 );
nand NAND2_8666 ( P3_U4813 , P3_R1212_U62 , P3_U3040 );
nand NAND2_8667 ( P3_U4814 , P3_U3039 , P3_U3430 );
nand NAND2_8668 ( P3_U4815 , P3_R1209_U62 , P3_U3037 );
nand NAND3_8669 ( P3_U4816 , P3_U4814 , P3_U4813 , P3_U4815 );
nand NAND2_8670 ( P3_U4817 , P3_R1054_U78 , P3_U3051 );
nand NAND2_8671 ( P3_U4818 , P3_U5768 , P3_U3430 );
nand NAND2_8672 ( P3_U4819 , P3_U3042 , P3_U4816 );
nand NAND2_8673 ( P3_U4820 , P3_R1212_U62 , P3_U3041 );
nand NAND2_8674 ( P3_U4821 , P3_REG3_REG_14_ , P3_U3151 );
nand NAND2_8675 ( P3_U4822 , P3_R1209_U62 , P3_U3038 );
nand NAND2_8676 ( P3_U4823 , P3_ADDR_REG_14_ , P3_U4760 );
nand NAND2_8677 ( P3_U4824 , P3_R1212_U63 , P3_U3040 );
nand NAND2_8678 ( P3_U4825 , P3_U3039 , P3_U3427 );
nand NAND2_8679 ( P3_U4826 , P3_R1209_U63 , P3_U3037 );
nand NAND3_8680 ( P3_U4827 , P3_U4825 , P3_U4824 , P3_U4826 );
nand NAND2_8681 ( P3_U4828 , P3_R1054_U70 , P3_U3051 );
nand NAND2_8682 ( P3_U4829 , P3_U5768 , P3_U3427 );
nand NAND2_8683 ( P3_U4830 , P3_U3042 , P3_U4827 );
nand NAND2_8684 ( P3_U4831 , P3_R1212_U63 , P3_U3041 );
nand NAND2_8685 ( P3_U4832 , P3_REG3_REG_13_ , P3_U3151 );
nand NAND2_8686 ( P3_U4833 , P3_R1209_U63 , P3_U3038 );
nand NAND2_8687 ( P3_U4834 , P3_ADDR_REG_13_ , P3_U4760 );
nand NAND2_8688 ( P3_U4835 , P3_R1212_U64 , P3_U3040 );
nand NAND2_8689 ( P3_U4836 , P3_U3039 , P3_U3424 );
nand NAND2_8690 ( P3_U4837 , P3_R1209_U64 , P3_U3037 );
nand NAND3_8691 ( P3_U4838 , P3_U4836 , P3_U4835 , P3_U4837 );
nand NAND2_8692 ( P3_U4839 , P3_R1054_U71 , P3_U3051 );
nand NAND2_8693 ( P3_U4840 , P3_U5768 , P3_U3424 );
nand NAND2_8694 ( P3_U4841 , P3_U3042 , P3_U4838 );
nand NAND2_8695 ( P3_U4842 , P3_R1212_U64 , P3_U3041 );
nand NAND2_8696 ( P3_U4843 , P3_REG3_REG_12_ , P3_U3151 );
nand NAND2_8697 ( P3_U4844 , P3_R1209_U64 , P3_U3038 );
nand NAND2_8698 ( P3_U4845 , P3_ADDR_REG_12_ , P3_U4760 );
nand NAND2_8699 ( P3_U4846 , P3_R1212_U65 , P3_U3040 );
nand NAND2_8700 ( P3_U4847 , P3_U3039 , P3_U3421 );
nand NAND2_8701 ( P3_U4848 , P3_R1209_U65 , P3_U3037 );
nand NAND3_8702 ( P3_U4849 , P3_U4847 , P3_U4846 , P3_U4848 );
nand NAND2_8703 ( P3_U4850 , P3_R1054_U12 , P3_U3051 );
nand NAND2_8704 ( P3_U4851 , P3_U5768 , P3_U3421 );
nand NAND2_8705 ( P3_U4852 , P3_U3042 , P3_U4849 );
nand NAND2_8706 ( P3_U4853 , P3_R1212_U65 , P3_U3041 );
nand NAND2_8707 ( P3_U4854 , P3_REG3_REG_11_ , P3_U3151 );
nand NAND2_8708 ( P3_U4855 , P3_R1209_U65 , P3_U3038 );
nand NAND2_8709 ( P3_U4856 , P3_ADDR_REG_11_ , P3_U4760 );
nand NAND2_8710 ( P3_U4857 , P3_R1212_U66 , P3_U3040 );
nand NAND2_8711 ( P3_U4858 , P3_U3039 , P3_U3418 );
nand NAND2_8712 ( P3_U4859 , P3_R1209_U66 , P3_U3037 );
nand NAND3_8713 ( P3_U4860 , P3_U4858 , P3_U4857 , P3_U4859 );
nand NAND2_8714 ( P3_U4861 , P3_R1054_U79 , P3_U3051 );
nand NAND2_8715 ( P3_U4862 , P3_U5768 , P3_U3418 );
nand NAND2_8716 ( P3_U4863 , P3_U3042 , P3_U4860 );
nand NAND2_8717 ( P3_U4864 , P3_R1212_U66 , P3_U3041 );
nand NAND2_8718 ( P3_U4865 , P3_REG3_REG_10_ , P3_U3151 );
nand NAND2_8719 ( P3_U4866 , P3_R1209_U66 , P3_U3038 );
nand NAND2_8720 ( P3_U4867 , P3_ADDR_REG_10_ , P3_U4760 );
nand NAND2_8721 ( P3_U4868 , P3_R1212_U49 , P3_U3040 );
nand NAND2_8722 ( P3_U4869 , P3_U3039 , P3_U3415 );
nand NAND2_8723 ( P3_U4870 , P3_R1209_U49 , P3_U3037 );
nand NAND3_8724 ( P3_U4871 , P3_U4869 , P3_U4868 , P3_U4870 );
nand NAND2_8725 ( P3_U4872 , P3_R1054_U72 , P3_U3051 );
nand NAND2_8726 ( P3_U4873 , P3_U5768 , P3_U3415 );
nand NAND2_8727 ( P3_U4874 , P3_U3042 , P3_U4871 );
nand NAND2_8728 ( P3_U4875 , P3_R1212_U49 , P3_U3041 );
nand NAND2_8729 ( P3_U4876 , P3_REG3_REG_9_ , P3_U3151 );
nand NAND2_8730 ( P3_U4877 , P3_R1209_U49 , P3_U3038 );
nand NAND2_8731 ( P3_U4878 , P3_ADDR_REG_9_ , P3_U4760 );
nand NAND2_8732 ( P3_U4879 , P3_R1212_U50 , P3_U3040 );
nand NAND2_8733 ( P3_U4880 , P3_U3039 , P3_U3412 );
nand NAND2_8734 ( P3_U4881 , P3_R1209_U50 , P3_U3037 );
nand NAND3_8735 ( P3_U4882 , P3_U4880 , P3_U4879 , P3_U4881 );
nand NAND2_8736 ( P3_U4883 , P3_R1054_U16 , P3_U3051 );
nand NAND2_8737 ( P3_U4884 , P3_U5768 , P3_U3412 );
nand NAND2_8738 ( P3_U4885 , P3_U3042 , P3_U4882 );
nand NAND2_8739 ( P3_U4886 , P3_R1212_U50 , P3_U3041 );
nand NAND2_8740 ( P3_U4887 , P3_REG3_REG_8_ , P3_U3151 );
nand NAND2_8741 ( P3_U4888 , P3_R1209_U50 , P3_U3038 );
nand NAND2_8742 ( P3_U4889 , P3_ADDR_REG_8_ , P3_U4760 );
nand NAND2_8743 ( P3_U4890 , P3_R1212_U51 , P3_U3040 );
nand NAND2_8744 ( P3_U4891 , P3_U3039 , P3_U3409 );
nand NAND2_8745 ( P3_U4892 , P3_R1209_U51 , P3_U3037 );
nand NAND3_8746 ( P3_U4893 , P3_U4891 , P3_U4890 , P3_U4892 );
nand NAND2_8747 ( P3_U4894 , P3_R1054_U73 , P3_U3051 );
nand NAND2_8748 ( P3_U4895 , P3_U5768 , P3_U3409 );
nand NAND2_8749 ( P3_U4896 , P3_U3042 , P3_U4893 );
nand NAND2_8750 ( P3_U4897 , P3_R1212_U51 , P3_U3041 );
nand NAND2_8751 ( P3_U4898 , P3_REG3_REG_7_ , P3_U3151 );
nand NAND2_8752 ( P3_U4899 , P3_R1209_U51 , P3_U3038 );
nand NAND2_8753 ( P3_U4900 , P3_ADDR_REG_7_ , P3_U4760 );
nand NAND2_8754 ( P3_U4901 , P3_R1212_U52 , P3_U3040 );
nand NAND2_8755 ( P3_U4902 , P3_U3039 , P3_U3406 );
nand NAND2_8756 ( P3_U4903 , P3_R1209_U52 , P3_U3037 );
nand NAND3_8757 ( P3_U4904 , P3_U4902 , P3_U4901 , P3_U4903 );
nand NAND2_8758 ( P3_U4905 , P3_R1054_U15 , P3_U3051 );
nand NAND2_8759 ( P3_U4906 , P3_U5768 , P3_U3406 );
nand NAND2_8760 ( P3_U4907 , P3_U3042 , P3_U4904 );
nand NAND2_8761 ( P3_U4908 , P3_R1212_U52 , P3_U3041 );
nand NAND2_8762 ( P3_U4909 , P3_REG3_REG_6_ , P3_U3151 );
nand NAND2_8763 ( P3_U4910 , P3_R1209_U52 , P3_U3038 );
nand NAND2_8764 ( P3_U4911 , P3_ADDR_REG_6_ , P3_U4760 );
nand NAND2_8765 ( P3_U4912 , P3_R1212_U53 , P3_U3040 );
nand NAND2_8766 ( P3_U4913 , P3_U3039 , P3_U3403 );
nand NAND2_8767 ( P3_U4914 , P3_R1209_U53 , P3_U3037 );
nand NAND3_8768 ( P3_U4915 , P3_U4913 , P3_U4912 , P3_U4914 );
nand NAND2_8769 ( P3_U4916 , P3_R1054_U74 , P3_U3051 );
nand NAND2_8770 ( P3_U4917 , P3_U5768 , P3_U3403 );
nand NAND2_8771 ( P3_U4918 , P3_U3042 , P3_U4915 );
nand NAND2_8772 ( P3_U4919 , P3_R1212_U53 , P3_U3041 );
nand NAND2_8773 ( P3_U4920 , P3_REG3_REG_5_ , P3_U3151 );
nand NAND2_8774 ( P3_U4921 , P3_R1209_U53 , P3_U3038 );
nand NAND2_8775 ( P3_U4922 , P3_ADDR_REG_5_ , P3_U4760 );
nand NAND2_8776 ( P3_U4923 , P3_R1212_U54 , P3_U3040 );
nand NAND2_8777 ( P3_U4924 , P3_U3039 , P3_U3400 );
nand NAND2_8778 ( P3_U4925 , P3_R1209_U54 , P3_U3037 );
nand NAND3_8779 ( P3_U4926 , P3_U4924 , P3_U4923 , P3_U4925 );
nand NAND2_8780 ( P3_U4927 , P3_R1054_U75 , P3_U3051 );
nand NAND2_8781 ( P3_U4928 , P3_U5768 , P3_U3400 );
nand NAND2_8782 ( P3_U4929 , P3_U3042 , P3_U4926 );
nand NAND2_8783 ( P3_U4930 , P3_R1212_U54 , P3_U3041 );
nand NAND2_8784 ( P3_U4931 , P3_REG3_REG_4_ , P3_U3151 );
nand NAND2_8785 ( P3_U4932 , P3_R1209_U54 , P3_U3038 );
nand NAND2_8786 ( P3_U4933 , P3_ADDR_REG_4_ , P3_U4760 );
nand NAND2_8787 ( P3_U4934 , P3_R1212_U55 , P3_U3040 );
nand NAND2_8788 ( P3_U4935 , P3_U3039 , P3_U3397 );
nand NAND2_8789 ( P3_U4936 , P3_R1209_U55 , P3_U3037 );
nand NAND3_8790 ( P3_U4937 , P3_U4935 , P3_U4934 , P3_U4936 );
nand NAND2_8791 ( P3_U4938 , P3_R1054_U14 , P3_U3051 );
nand NAND2_8792 ( P3_U4939 , P3_U5768 , P3_U3397 );
nand NAND2_8793 ( P3_U4940 , P3_U3042 , P3_U4937 );
nand NAND2_8794 ( P3_U4941 , P3_R1212_U55 , P3_U3041 );
nand NAND2_8795 ( P3_U4942 , P3_REG3_REG_3_ , P3_U3151 );
nand NAND2_8796 ( P3_U4943 , P3_R1209_U55 , P3_U3038 );
nand NAND2_8797 ( P3_U4944 , P3_ADDR_REG_3_ , P3_U4760 );
nand NAND2_8798 ( P3_U4945 , P3_R1212_U56 , P3_U3040 );
nand NAND2_8799 ( P3_U4946 , P3_U3039 , P3_U3394 );
nand NAND2_8800 ( P3_U4947 , P3_R1209_U56 , P3_U3037 );
nand NAND3_8801 ( P3_U4948 , P3_U4946 , P3_U4945 , P3_U4947 );
nand NAND2_8802 ( P3_U4949 , P3_R1054_U76 , P3_U3051 );
nand NAND2_8803 ( P3_U4950 , P3_U5768 , P3_U3394 );
nand NAND2_8804 ( P3_U4951 , P3_U3042 , P3_U4948 );
nand NAND2_8805 ( P3_U4952 , P3_R1212_U56 , P3_U3041 );
nand NAND2_8806 ( P3_U4953 , P3_REG3_REG_2_ , P3_U3151 );
nand NAND2_8807 ( P3_U4954 , P3_R1209_U56 , P3_U3038 );
nand NAND2_8808 ( P3_U4955 , P3_ADDR_REG_2_ , P3_U4760 );
nand NAND2_8809 ( P3_U4956 , P3_R1212_U57 , P3_U3040 );
nand NAND2_8810 ( P3_U4957 , P3_U3039 , P3_U3391 );
nand NAND2_8811 ( P3_U4958 , P3_R1209_U57 , P3_U3037 );
nand NAND3_8812 ( P3_U4959 , P3_U4957 , P3_U4956 , P3_U4958 );
nand NAND2_8813 ( P3_U4960 , P3_R1054_U66 , P3_U3051 );
nand NAND2_8814 ( P3_U4961 , P3_U5768 , P3_U3391 );
nand NAND2_8815 ( P3_U4962 , P3_U3042 , P3_U4959 );
nand NAND2_8816 ( P3_U4963 , P3_R1212_U57 , P3_U3041 );
nand NAND2_8817 ( P3_U4964 , P3_REG3_REG_1_ , P3_U3151 );
nand NAND2_8818 ( P3_U4965 , P3_R1209_U57 , P3_U3038 );
nand NAND2_8819 ( P3_U4966 , P3_ADDR_REG_1_ , P3_U4760 );
nand NAND2_8820 ( P3_U4967 , P3_R1212_U7 , P3_U3040 );
nand NAND2_8821 ( P3_U4968 , P3_U3039 , P3_U3386 );
nand NAND2_8822 ( P3_U4969 , P3_R1209_U7 , P3_U3037 );
nand NAND3_8823 ( P3_U4970 , P3_U4968 , P3_U4967 , P3_U4969 );
nand NAND2_8824 ( P3_U4971 , P3_R1054_U17 , P3_U3051 );
nand NAND2_8825 ( P3_U4972 , P3_U5768 , P3_U3386 );
nand NAND2_8826 ( P3_U4973 , P3_U3042 , P3_U4970 );
nand NAND2_8827 ( P3_U4974 , P3_R1212_U7 , P3_U3041 );
nand NAND2_8828 ( P3_U4975 , P3_REG3_REG_0_ , P3_U3151 );
nand NAND2_8829 ( P3_U4976 , P3_R1209_U7 , P3_U3038 );
nand NAND2_8830 ( P3_U4977 , P3_ADDR_REG_0_ , P3_U4760 );
not NOT1_8831 ( P3_U4978 , P3_U3868 );
nand NAND3_8832 ( P3_U4979 , P3_U5942 , P3_U5941 , P3_U3050 );
nand NAND3_8833 ( P3_U4980 , P3_U3023 , P3_U3909 , P3_U3867 );
nand NAND2_8834 ( P3_U4981 , P3_B_REG , P3_U4979 );
nand NAND2_8835 ( P3_U4982 , P3_U3036 , P3_U3078 );
nand NAND2_8836 ( P3_U4983 , P3_U3032 , P3_U3072 );
nand NAND2_8837 ( P3_U4984 , P3_SUB_609_U21 , P3_U3304 );
nand NAND3_8838 ( P3_U4985 , P3_U4983 , P3_U4982 , P3_U4984 );
nand NAND5_8839 ( P3_U4986 , P3_U3311 , P3_U3875 , P3_U3888 , P3_U5425 , P3_U3312 );
nand NAND2_8840 ( P3_U4987 , P3_U3894 , P3_U4986 );
nand NAND2_8841 ( P3_U4988 , P3_U3889 , P3_U3895 );
nand NAND2_8842 ( P3_U4989 , P3_U4988 , P3_U4987 );
nand NAND2_8843 ( P3_U4990 , P3_U3911 , P3_U3378 );
nand NAND2_8844 ( P3_U4991 , P3_U3889 , P3_U3304 );
nand NAND2_8845 ( P3_U4992 , P3_U4986 , P3_U3303 );
not NOT1_8846 ( P3_U4993 , P3_U3370 );
nand NAND2_8847 ( P3_U4994 , P3_U3434 , P3_U5420 );
nand NAND2_8848 ( P3_U4995 , P3_SUB_609_U21 , P3_U3371 );
nand NAND2_8849 ( P3_U4996 , P3_R1158_U114 , P3_U3035 );
nand NAND2_8850 ( P3_U4997 , P3_U3031 , P3_U4985 );
nand NAND2_8851 ( P3_U4998 , P3_REG3_REG_15_ , P3_U3151 );
nand NAND2_8852 ( P3_U4999 , P3_U3036 , P3_U3057 );
nand NAND2_8853 ( P3_U5000 , P3_U3032 , P3_U3052 );
nand NAND2_8854 ( P3_U5001 , P3_SUB_609_U26 , P3_U3304 );
nand NAND3_8855 ( P3_U5002 , P3_U5000 , P3_U4999 , P3_U5001 );
nand NAND2_8856 ( P3_U5003 , P3_U3365 , P3_U3303 );
nand NAND2_8857 ( P3_U5004 , P3_U4993 , P3_U5003 );
nand NAND2_8858 ( P3_U5005 , P3_U3894 , P3_U3365 );
nand NAND2_8859 ( P3_U5006 , P3_U3360 , P3_U5005 );
nand NAND2_8860 ( P3_U5007 , P3_U3045 , P3_U3901 );
nand NAND2_8861 ( P3_U5008 , P3_U3044 , P3_SUB_609_U26 );
nand NAND2_8862 ( P3_U5009 , P3_R1158_U16 , P3_U3035 );
nand NAND2_8863 ( P3_U5010 , P3_U3031 , P3_U5002 );
nand NAND2_8864 ( P3_U5011 , P3_REG3_REG_26_ , P3_U3151 );
nand NAND2_8865 ( P3_U5012 , P3_U3036 , P3_U3066 );
nand NAND2_8866 ( P3_U5013 , P3_U3032 , P3_U3069 );
nand NAND2_8867 ( P3_U5014 , P3_SUB_609_U8 , P3_U3304 );
nand NAND3_8868 ( P3_U5015 , P3_U5013 , P3_U5012 , P3_U5014 );
nand NAND2_8869 ( P3_U5016 , P3_U3407 , P3_U5420 );
nand NAND2_8870 ( P3_U5017 , P3_SUB_609_U8 , P3_U3371 );
nand NAND2_8871 ( P3_U5018 , P3_R1158_U97 , P3_U3035 );
nand NAND2_8872 ( P3_U5019 , P3_U3031 , P3_U5015 );
nand NAND2_8873 ( P3_U5020 , P3_REG3_REG_6_ , P3_U3151 );
nand NAND2_8874 ( P3_U5021 , P3_U3036 , P3_U3068 );
nand NAND2_8875 ( P3_U5022 , P3_U3032 , P3_U3080 );
nand NAND2_8876 ( P3_U5023 , P3_SUB_609_U11 , P3_U3304 );
nand NAND3_8877 ( P3_U5024 , P3_U5022 , P3_U5021 , P3_U5023 );
nand NAND2_8878 ( P3_U5025 , P3_U3443 , P3_U5420 );
nand NAND2_8879 ( P3_U5026 , P3_SUB_609_U11 , P3_U3371 );
nand NAND2_8880 ( P3_U5027 , P3_R1158_U112 , P3_U3035 );
nand NAND2_8881 ( P3_U5028 , P3_U3031 , P3_U5024 );
nand NAND2_8882 ( P3_U5029 , P3_REG3_REG_18_ , P3_U3151 );
nand NAND2_8883 ( P3_U5030 , P3_U3036 , P3_U3077 );
nand NAND2_8884 ( P3_U5031 , P3_U3032 , P3_U3063 );
nand NAND2_8885 ( P3_U5032 , P3_REG3_REG_2_ , P3_U3304 );
nand NAND3_8886 ( P3_U5033 , P3_U5031 , P3_U5030 , P3_U5032 );
nand NAND2_8887 ( P3_U5034 , P3_U3395 , P3_U5420 );
nand NAND2_8888 ( P3_U5035 , P3_REG3_REG_2_ , P3_U3371 );
nand NAND2_8889 ( P3_U5036 , P3_R1158_U100 , P3_U3035 );
nand NAND2_8890 ( P3_U5037 , P3_U3031 , P3_U5033 );
nand NAND2_8891 ( P3_U5038 , P3_REG3_REG_2_ , P3_U3151 );
nand NAND2_8892 ( P3_U5039 , P3_U3036 , P3_U3061 );
nand NAND2_8893 ( P3_U5040 , P3_U3032 , P3_U3071 );
nand NAND2_8894 ( P3_U5041 , P3_SUB_609_U9 , P3_U3304 );
nand NAND3_8895 ( P3_U5042 , P3_U5040 , P3_U5039 , P3_U5041 );
nand NAND2_8896 ( P3_U5043 , P3_U3422 , P3_U5420 );
nand NAND2_8897 ( P3_U5044 , P3_SUB_609_U9 , P3_U3371 );
nand NAND2_8898 ( P3_U5045 , P3_R1158_U117 , P3_U3035 );
nand NAND2_8899 ( P3_U5046 , P3_U3031 , P3_U5042 );
nand NAND2_8900 ( P3_U5047 , P3_REG3_REG_11_ , P3_U3151 );
nand NAND2_8901 ( P3_U5048 , P3_U3036 , P3_U3074 );
nand NAND2_8902 ( P3_U5049 , P3_U3032 , P3_U3065 );
nand NAND2_8903 ( P3_U5050 , P3_SUB_609_U17 , P3_U3304 );
nand NAND3_8904 ( P3_U5051 , P3_U5049 , P3_U5048 , P3_U5050 );
nand NAND2_8905 ( P3_U5052 , P3_U3045 , P3_U3905 );
nand NAND2_8906 ( P3_U5053 , P3_U3044 , P3_SUB_609_U17 );
nand NAND2_8907 ( P3_U5054 , P3_R1158_U108 , P3_U3035 );
nand NAND2_8908 ( P3_U5055 , P3_U3031 , P3_U5051 );
nand NAND2_8909 ( P3_U5056 , P3_REG3_REG_22_ , P3_U3151 );
nand NAND2_8910 ( P3_U5057 , P3_U3036 , P3_U3071 );
nand NAND2_8911 ( P3_U5058 , P3_U3032 , P3_U3078 );
nand NAND2_8912 ( P3_U5059 , P3_SUB_609_U24 , P3_U3304 );
nand NAND3_8913 ( P3_U5060 , P3_U5058 , P3_U5057 , P3_U5059 );
nand NAND2_8914 ( P3_U5061 , P3_U3428 , P3_U5420 );
nand NAND2_8915 ( P3_U5062 , P3_SUB_609_U24 , P3_U3371 );
nand NAND2_8916 ( P3_U5063 , P3_R1158_U13 , P3_U3035 );
nand NAND2_8917 ( P3_U5064 , P3_U3031 , P3_U5060 );
nand NAND2_8918 ( P3_U5065 , P3_REG3_REG_13_ , P3_U3151 );
nand NAND2_8919 ( P3_U5066 , P3_U3036 , P3_U3080 );
nand NAND2_8920 ( P3_U5067 , P3_U3032 , P3_U3074 );
nand NAND2_8921 ( P3_U5068 , P3_SUB_609_U20 , P3_U3304 );
nand NAND3_8922 ( P3_U5069 , P3_U5067 , P3_U5066 , P3_U5068 );
nand NAND2_8923 ( P3_U5070 , P3_U3045 , P3_U3907 );
nand NAND2_8924 ( P3_U5071 , P3_U3044 , P3_SUB_609_U20 );
nand NAND2_8925 ( P3_U5072 , P3_R1158_U109 , P3_U3035 );
nand NAND2_8926 ( P3_U5073 , P3_U3031 , P3_U5069 );
nand NAND2_8927 ( P3_U5074 , P3_REG3_REG_20_ , P3_U3151 );
nand NAND2_8928 ( P3_U5075 , P3_U3031 , P3_U3304 );
nand NAND2_8929 ( P3_U5076 , P3_U5419 , P3_U5075 );
nand NAND2_8930 ( P3_U5077 , P3_U3787 , P3_U3032 );
nand NAND2_8931 ( P3_U5078 , P3_U3387 , P3_U5420 );
nand NAND2_8932 ( P3_U5079 , P3_REG3_REG_0_ , P3_U5076 );
nand NAND2_8933 ( P3_U5080 , P3_R1158_U94 , P3_U3035 );
nand NAND2_8934 ( P3_U5081 , P3_REG3_REG_0_ , P3_U3151 );
nand NAND2_8935 ( P3_U5082 , P3_U3036 , P3_U3083 );
nand NAND2_8936 ( P3_U5083 , P3_U3032 , P3_U3061 );
nand NAND2_8937 ( P3_U5084 , P3_SUB_609_U14 , P3_U3304 );
nand NAND3_8938 ( P3_U5085 , P3_U5083 , P3_U5082 , P3_U5084 );
nand NAND2_8939 ( P3_U5086 , P3_U3416 , P3_U5420 );
nand NAND2_8940 ( P3_U5087 , P3_SUB_609_U14 , P3_U3371 );
nand NAND2_8941 ( P3_U5088 , P3_R1158_U95 , P3_U3035 );
nand NAND2_8942 ( P3_U5089 , P3_U3031 , P3_U5085 );
nand NAND2_8943 ( P3_U5090 , P3_REG3_REG_9_ , P3_U3151 );
nand NAND2_8944 ( P3_U5091 , P3_U3036 , P3_U3063 );
nand NAND2_8945 ( P3_U5092 , P3_U3032 , P3_U3066 );
nand NAND2_8946 ( P3_U5093 , P3_SUB_609_U29 , P3_U3304 );
nand NAND3_8947 ( P3_U5094 , P3_U5092 , P3_U5091 , P3_U5093 );
nand NAND2_8948 ( P3_U5095 , P3_U3401 , P3_U5420 );
nand NAND2_8949 ( P3_U5096 , P3_SUB_609_U29 , P3_U3371 );
nand NAND2_8950 ( P3_U5097 , P3_R1158_U99 , P3_U3035 );
nand NAND2_8951 ( P3_U5098 , P3_U3031 , P3_U5094 );
nand NAND2_8952 ( P3_U5099 , P3_REG3_REG_4_ , P3_U3151 );
nand NAND2_8953 ( P3_U5100 , P3_U3036 , P3_U3065 );
nand NAND2_8954 ( P3_U5101 , P3_U3032 , P3_U3057 );
nand NAND2_8955 ( P3_U5102 , P3_SUB_609_U10 , P3_U3304 );
nand NAND3_8956 ( P3_U5103 , P3_U5101 , P3_U5100 , P3_U5102 );
nand NAND2_8957 ( P3_U5104 , P3_U3045 , P3_U3903 );
nand NAND2_8958 ( P3_U5105 , P3_U3044 , P3_SUB_609_U10 );
nand NAND2_8959 ( P3_U5106 , P3_R1158_U106 , P3_U3035 );
nand NAND2_8960 ( P3_U5107 , P3_U3031 , P3_U5103 );
nand NAND2_8961 ( P3_U5108 , P3_REG3_REG_24_ , P3_U3151 );
nand NAND2_8962 ( P3_U5109 , P3_U3036 , P3_U3072 );
nand NAND2_8963 ( P3_U5110 , P3_U3032 , P3_U3081 );
nand NAND2_8964 ( P3_U5111 , P3_SUB_609_U19 , P3_U3304 );
nand NAND3_8965 ( P3_U5112 , P3_U5110 , P3_U5109 , P3_U5111 );
nand NAND2_8966 ( P3_U5113 , P3_U3440 , P3_U5420 );
nand NAND2_8967 ( P3_U5114 , P3_SUB_609_U19 , P3_U3371 );
nand NAND2_8968 ( P3_U5115 , P3_R1158_U14 , P3_U3035 );
nand NAND2_8969 ( P3_U5116 , P3_U3031 , P3_U5112 );
nand NAND2_8970 ( P3_U5117 , P3_REG3_REG_17_ , P3_U3151 );
nand NAND2_8971 ( P3_U5118 , P3_U3036 , P3_U3059 );
nand NAND2_8972 ( P3_U5119 , P3_U3032 , P3_U3070 );
nand NAND2_8973 ( P3_U5120 , P3_SUB_609_U53 , P3_U3304 );
nand NAND3_8974 ( P3_U5121 , P3_U5119 , P3_U5118 , P3_U5120 );
nand NAND2_8975 ( P3_U5122 , P3_U3404 , P3_U5420 );
nand NAND2_8976 ( P3_U5123 , P3_SUB_609_U53 , P3_U3371 );
nand NAND2_8977 ( P3_U5124 , P3_R1158_U98 , P3_U3035 );
nand NAND2_8978 ( P3_U5125 , P3_U3031 , P3_U5121 );
nand NAND2_8979 ( P3_U5126 , P3_REG3_REG_5_ , P3_U3151 );
nand NAND2_8980 ( P3_U5127 , P3_U3036 , P3_U3073 );
nand NAND2_8981 ( P3_U5128 , P3_U3032 , P3_U3068 );
nand NAND2_8982 ( P3_U5129 , P3_SUB_609_U7 , P3_U3304 );
nand NAND3_8983 ( P3_U5130 , P3_U5128 , P3_U5127 , P3_U5129 );
nand NAND2_8984 ( P3_U5131 , P3_U3437 , P3_U5420 );
nand NAND2_8985 ( P3_U5132 , P3_SUB_609_U7 , P3_U3371 );
nand NAND2_8986 ( P3_U5133 , P3_R1158_U113 , P3_U3035 );
nand NAND2_8987 ( P3_U5134 , P3_U3031 , P3_U5130 );
nand NAND2_8988 ( P3_U5135 , P3_REG3_REG_16_ , P3_U3151 );
nand NAND2_8989 ( P3_U5136 , P3_U3036 , P3_U3064 );
nand NAND2_8990 ( P3_U5137 , P3_U3032 , P3_U3056 );
nand NAND2_8991 ( P3_U5138 , P3_SUB_609_U16 , P3_U3304 );
nand NAND3_8992 ( P3_U5139 , P3_U5137 , P3_U5136 , P3_U5138 );
nand NAND2_8993 ( P3_U5140 , P3_U3045 , P3_U3902 );
nand NAND2_8994 ( P3_U5141 , P3_U3044 , P3_SUB_609_U16 );
nand NAND2_8995 ( P3_U5142 , P3_R1158_U105 , P3_U3035 );
nand NAND2_8996 ( P3_U5143 , P3_U3031 , P3_U5139 );
nand NAND2_8997 ( P3_U5144 , P3_REG3_REG_25_ , P3_U3151 );
nand NAND2_8998 ( P3_U5145 , P3_U3036 , P3_U3062 );
nand NAND2_8999 ( P3_U5146 , P3_U3032 , P3_U3079 );
nand NAND2_9000 ( P3_U5147 , P3_SUB_609_U23 , P3_U3304 );
nand NAND3_9001 ( P3_U5148 , P3_U5146 , P3_U5145 , P3_U5147 );
nand NAND2_9002 ( P3_U5149 , P3_U3425 , P3_U5420 );
nand NAND2_9003 ( P3_U5150 , P3_SUB_609_U23 , P3_U3371 );
nand NAND2_9004 ( P3_U5151 , P3_R1158_U116 , P3_U3035 );
nand NAND2_9005 ( P3_U5152 , P3_U3031 , P3_U5148 );
nand NAND2_9006 ( P3_U5153 , P3_REG3_REG_12_ , P3_U3151 );
nand NAND2_9007 ( P3_U5154 , P3_U3036 , P3_U3075 );
nand NAND2_9008 ( P3_U5155 , P3_U3032 , P3_U3060 );
nand NAND2_9009 ( P3_U5156 , P3_SUB_609_U27 , P3_U3304 );
nand NAND3_9010 ( P3_U5157 , P3_U5155 , P3_U5154 , P3_U5156 );
nand NAND2_9011 ( P3_U5158 , P3_U3045 , P3_U3906 );
nand NAND2_9012 ( P3_U5159 , P3_U3044 , P3_SUB_609_U27 );
nand NAND2_9013 ( P3_U5160 , P3_R1158_U15 , P3_U3035 );
nand NAND2_9014 ( P3_U5161 , P3_U3031 , P3_U5157 );
nand NAND2_9015 ( P3_U5162 , P3_REG3_REG_21_ , P3_U3151 );
nand NAND2_9016 ( P3_U5163 , P3_U3036 , P3_U3076 );
nand NAND2_9017 ( P3_U5164 , P3_U3032 , P3_U3067 );
nand NAND2_9018 ( P3_U5165 , P3_REG3_REG_1_ , P3_U3304 );
nand NAND3_9019 ( P3_U5166 , P3_U5164 , P3_U5163 , P3_U5165 );
nand NAND2_9020 ( P3_U5167 , P3_U3392 , P3_U5420 );
nand NAND2_9021 ( P3_U5168 , P3_REG3_REG_1_ , P3_U3371 );
nand NAND2_9022 ( P3_U5169 , P3_R1158_U110 , P3_U3035 );
nand NAND2_9023 ( P3_U5170 , P3_U3031 , P3_U5166 );
nand NAND2_9024 ( P3_U5171 , P3_REG3_REG_1_ , P3_U3151 );
nand NAND2_9025 ( P3_U5172 , P3_U3036 , P3_U3069 );
nand NAND2_9026 ( P3_U5173 , P3_U3032 , P3_U3082 );
nand NAND2_9027 ( P3_U5174 , P3_SUB_609_U12 , P3_U3304 );
nand NAND3_9028 ( P3_U5175 , P3_U5173 , P3_U5172 , P3_U5174 );
nand NAND2_9029 ( P3_U5176 , P3_U3413 , P3_U5420 );
nand NAND2_9030 ( P3_U5177 , P3_SUB_609_U12 , P3_U3371 );
nand NAND2_9031 ( P3_U5178 , P3_R1158_U96 , P3_U3035 );
nand NAND2_9032 ( P3_U5179 , P3_U3031 , P3_U5175 );
nand NAND2_9033 ( P3_U5180 , P3_REG3_REG_8_ , P3_U3151 );
nand NAND2_9034 ( P3_U5181 , P3_U3036 , P3_U3052 );
nand NAND2_9035 ( P3_U5182 , P3_U3032 , P3_U3054 );
nand NAND2_9036 ( P3_U5183 , P3_SUB_609_U28 , P3_U3304 );
nand NAND3_9037 ( P3_U5184 , P3_U5182 , P3_U5181 , P3_U5183 );
nand NAND2_9038 ( P3_U5185 , P3_U3045 , P3_U3899 );
nand NAND2_9039 ( P3_U5186 , P3_U3044 , P3_SUB_609_U28 );
nand NAND2_9040 ( P3_U5187 , P3_R1158_U101 , P3_U3035 );
nand NAND2_9041 ( P3_U5188 , P3_U3031 , P3_U5184 );
nand NAND2_9042 ( P3_U5189 , P3_REG3_REG_28_ , P3_U3151 );
nand NAND2_9043 ( P3_U5190 , P3_U3036 , P3_U3081 );
nand NAND2_9044 ( P3_U5191 , P3_U3032 , P3_U3075 );
nand NAND2_9045 ( P3_U5192 , P3_SUB_609_U15 , P3_U3304 );
nand NAND3_9046 ( P3_U5193 , P3_U5191 , P3_U5190 , P3_U5192 );
nand NAND2_9047 ( P3_U5194 , P3_U3445 , P3_U5420 );
nand NAND2_9048 ( P3_U5195 , P3_SUB_609_U15 , P3_U3371 );
nand NAND2_9049 ( P3_U5196 , P3_R1158_U111 , P3_U3035 );
nand NAND2_9050 ( P3_U5197 , P3_U3031 , P3_U5193 );
nand NAND2_9051 ( P3_U5198 , P3_REG3_REG_19_ , P3_U3151 );
nand NAND2_9052 ( P3_U5199 , P3_U3036 , P3_U3067 );
nand NAND2_9053 ( P3_U5200 , P3_U3032 , P3_U3059 );
nand NAND2_9054 ( P3_U5201 , P3_SUB_609_U25 , P3_U3304 );
nand NAND3_9055 ( P3_U5202 , P3_U5200 , P3_U5199 , P3_U5201 );
nand NAND2_9056 ( P3_U5203 , P3_U3398 , P3_U5420 );
nand NAND2_9057 ( P3_U5204 , P3_SUB_609_U25 , P3_U3371 );
nand NAND2_9058 ( P3_U5205 , P3_R1158_U17 , P3_U3035 );
nand NAND2_9059 ( P3_U5206 , P3_U3031 , P3_U5202 );
nand NAND2_9060 ( P3_U5207 , P3_REG3_REG_3_ , P3_U3151 );
nand NAND2_9061 ( P3_U5208 , P3_U3036 , P3_U3082 );
nand NAND2_9062 ( P3_U5209 , P3_U3032 , P3_U3062 );
nand NAND2_9063 ( P3_U5210 , P3_SUB_609_U13 , P3_U3304 );
nand NAND3_9064 ( P3_U5211 , P3_U5209 , P3_U5208 , P3_U5210 );
nand NAND2_9065 ( P3_U5212 , P3_U3419 , P3_U5420 );
nand NAND2_9066 ( P3_U5213 , P3_SUB_609_U13 , P3_U3371 );
nand NAND2_9067 ( P3_U5214 , P3_R1158_U118 , P3_U3035 );
nand NAND2_9068 ( P3_U5215 , P3_U3031 , P3_U5211 );
nand NAND2_9069 ( P3_U5216 , P3_REG3_REG_10_ , P3_U3151 );
nand NAND2_9070 ( P3_U5217 , P3_U3036 , P3_U3060 );
nand NAND2_9071 ( P3_U5218 , P3_U3032 , P3_U3064 );
nand NAND2_9072 ( P3_U5219 , P3_SUB_609_U6 , P3_U3304 );
nand NAND3_9073 ( P3_U5220 , P3_U5218 , P3_U5217 , P3_U5219 );
nand NAND2_9074 ( P3_U5221 , P3_U3045 , P3_U3904 );
nand NAND2_9075 ( P3_U5222 , P3_U3044 , P3_SUB_609_U6 );
nand NAND2_9076 ( P3_U5223 , P3_R1158_U107 , P3_U3035 );
nand NAND2_9077 ( P3_U5224 , P3_U3031 , P3_U5220 );
nand NAND2_9078 ( P3_U5225 , P3_REG3_REG_23_ , P3_U3151 );
nand NAND2_9079 ( P3_U5226 , P3_U3036 , P3_U3079 );
nand NAND2_9080 ( P3_U5227 , P3_U3032 , P3_U3073 );
nand NAND2_9081 ( P3_U5228 , P3_SUB_609_U30 , P3_U3304 );
nand NAND3_9082 ( P3_U5229 , P3_U5227 , P3_U5226 , P3_U5228 );
nand NAND2_9083 ( P3_U5230 , P3_U3431 , P3_U5420 );
nand NAND2_9084 ( P3_U5231 , P3_SUB_609_U30 , P3_U3371 );
nand NAND2_9085 ( P3_U5232 , P3_R1158_U115 , P3_U3035 );
nand NAND2_9086 ( P3_U5233 , P3_U3031 , P3_U5229 );
nand NAND2_9087 ( P3_U5234 , P3_REG3_REG_14_ , P3_U3151 );
nand NAND2_9088 ( P3_U5235 , P3_U3036 , P3_U3056 );
nand NAND2_9089 ( P3_U5236 , P3_U3032 , P3_U3053 );
nand NAND2_9090 ( P3_U5237 , P3_SUB_609_U22 , P3_U3304 );
nand NAND3_9091 ( P3_U5238 , P3_U5236 , P3_U5235 , P3_U5237 );
nand NAND2_9092 ( P3_U5239 , P3_U3045 , P3_U3900 );
nand NAND2_9093 ( P3_U5240 , P3_U3044 , P3_SUB_609_U22 );
nand NAND2_9094 ( P3_U5241 , P3_R1158_U102 , P3_U3035 );
nand NAND2_9095 ( P3_U5242 , P3_U3031 , P3_U5238 );
nand NAND2_9096 ( P3_U5243 , P3_REG3_REG_27_ , P3_U3151 );
nand NAND2_9097 ( P3_U5244 , P3_U3036 , P3_U3070 );
nand NAND2_9098 ( P3_U5245 , P3_U3032 , P3_U3083 );
nand NAND2_9099 ( P3_U5246 , P3_SUB_609_U18 , P3_U3304 );
nand NAND3_9100 ( P3_U5247 , P3_U5245 , P3_U5244 , P3_U5246 );
nand NAND2_9101 ( P3_U5248 , P3_U3410 , P3_U5420 );
nand NAND2_9102 ( P3_U5249 , P3_SUB_609_U18 , P3_U3371 );
nand NAND2_9103 ( P3_U5250 , P3_R1158_U18 , P3_U3035 );
nand NAND2_9104 ( P3_U5251 , P3_U3031 , P3_U5247 );
nand NAND2_9105 ( P3_U5252 , P3_REG3_REG_7_ , P3_U3151 );
nand NAND2_9106 ( P3_U5253 , P3_U3898 , P3_U3046 );
nand NAND2_9107 ( P3_U5254 , P3_U3375 , P3_U3833 );
nand NAND2_9108 ( P3_U5255 , P3_U3816 , P3_U3815 );
nand NAND2_9109 ( P3_U5256 , P3_U3814 , P3_U3013 );
nand NAND2_9110 ( P3_U5257 , P3_U3880 , P3_U5256 );
nand NAND2_9111 ( P3_U5258 , P3_U3416 , P3_U5257 );
nand NAND2_9112 ( P3_U5259 , P3_U5255 , P3_U3082 );
nand NAND2_9113 ( P3_U5260 , P3_U3413 , P3_U5257 );
nand NAND2_9114 ( P3_U5261 , P3_U5255 , P3_U3083 );
nand NAND2_9115 ( P3_U5262 , P3_U3410 , P3_U5257 );
nand NAND2_9116 ( P3_U5263 , P3_U5255 , P3_U3069 );
nand NAND2_9117 ( P3_U5264 , P3_U3407 , P3_U5257 );
nand NAND2_9118 ( P3_U5265 , P3_U5255 , P3_U3070 );
nand NAND2_9119 ( P3_U5266 , P3_U3404 , P3_U5257 );
nand NAND2_9120 ( P3_U5267 , P3_U5255 , P3_U3066 );
nand NAND2_9121 ( P3_U5268 , P3_U3401 , P3_U5257 );
nand NAND2_9122 ( P3_U5269 , P3_U5255 , P3_U3059 );
nand NAND2_9123 ( P3_U5270 , P3_U3872 , P3_U5257 );
nand NAND2_9124 ( P3_U5271 , P3_U5255 , P3_U3055 );
nand NAND2_9125 ( P3_U5272 , P3_U3873 , P3_U5257 );
nand NAND2_9126 ( P3_U5273 , P3_U5255 , P3_U3058 );
nand NAND2_9127 ( P3_U5274 , P3_U3398 , P3_U5257 );
nand NAND2_9128 ( P3_U5275 , P3_U5255 , P3_U3063 );
nand NAND2_9129 ( P3_U5276 , P3_U3908 , P3_U5257 );
nand NAND2_9130 ( P3_U5277 , P3_U5255 , P3_U3054 );
nand NAND2_9131 ( P3_U5278 , P3_U3899 , P3_U5257 );
nand NAND2_9132 ( P3_U5279 , P3_U5255 , P3_U3053 );
nand NAND2_9133 ( P3_U5280 , P3_U3900 , P3_U5257 );
nand NAND2_9134 ( P3_U5281 , P3_U5255 , P3_U3052 );
nand NAND2_9135 ( P3_U5282 , P3_U3901 , P3_U5257 );
nand NAND2_9136 ( P3_U5283 , P3_U5255 , P3_U3056 );
nand NAND2_9137 ( P3_U5284 , P3_U3902 , P3_U5257 );
nand NAND2_9138 ( P3_U5285 , P3_U5255 , P3_U3057 );
nand NAND2_9139 ( P3_U5286 , P3_U3903 , P3_U5257 );
nand NAND2_9140 ( P3_U5287 , P3_U5255 , P3_U3064 );
nand NAND2_9141 ( P3_U5288 , P3_U3904 , P3_U5257 );
nand NAND2_9142 ( P3_U5289 , P3_U5255 , P3_U3065 );
nand NAND2_9143 ( P3_U5290 , P3_U3905 , P3_U5257 );
nand NAND2_9144 ( P3_U5291 , P3_U5255 , P3_U3060 );
nand NAND2_9145 ( P3_U5292 , P3_U3906 , P3_U5257 );
nand NAND2_9146 ( P3_U5293 , P3_U5255 , P3_U3074 );
nand NAND2_9147 ( P3_U5294 , P3_U3907 , P3_U5257 );
nand NAND2_9148 ( P3_U5295 , P3_U5255 , P3_U3075 );
nand NAND2_9149 ( P3_U5296 , P3_U3395 , P3_U5257 );
nand NAND2_9150 ( P3_U5297 , P3_U5255 , P3_U3067 );
nand NAND2_9151 ( P3_U5298 , P3_U3445 , P3_U5257 );
nand NAND2_9152 ( P3_U5299 , P3_U5255 , P3_U3080 );
nand NAND2_9153 ( P3_U5300 , P3_U3443 , P3_U5257 );
nand NAND2_9154 ( P3_U5301 , P3_U5255 , P3_U3081 );
nand NAND2_9155 ( P3_U5302 , P3_U3440 , P3_U5257 );
nand NAND2_9156 ( P3_U5303 , P3_U5255 , P3_U3068 );
nand NAND2_9157 ( P3_U5304 , P3_U3437 , P3_U5257 );
nand NAND2_9158 ( P3_U5305 , P3_U5255 , P3_U3072 );
nand NAND2_9159 ( P3_U5306 , P3_U3434 , P3_U5257 );
nand NAND2_9160 ( P3_U5307 , P3_U5255 , P3_U3073 );
nand NAND2_9161 ( P3_U5308 , P3_U3431 , P3_U5257 );
nand NAND2_9162 ( P3_U5309 , P3_U5255 , P3_U3078 );
nand NAND2_9163 ( P3_U5310 , P3_U3428 , P3_U5257 );
nand NAND2_9164 ( P3_U5311 , P3_U5255 , P3_U3079 );
nand NAND2_9165 ( P3_U5312 , P3_U3425 , P3_U5257 );
nand NAND2_9166 ( P3_U5313 , P3_U5255 , P3_U3071 );
nand NAND2_9167 ( P3_U5314 , P3_U3422 , P3_U5257 );
nand NAND2_9168 ( P3_U5315 , P3_U5255 , P3_U3062 );
nand NAND2_9169 ( P3_U5316 , P3_U3419 , P3_U5257 );
nand NAND2_9170 ( P3_U5317 , P3_U5255 , P3_U3061 );
nand NAND2_9171 ( P3_U5318 , P3_U3392 , P3_U5257 );
nand NAND2_9172 ( P3_U5319 , P3_U5255 , P3_U3077 );
nand NAND2_9173 ( P3_U5320 , P3_U3387 , P3_U5257 );
nand NAND2_9174 ( P3_U5321 , P3_U5255 , P3_U3076 );
nand NAND2_9175 ( P3_U5322 , P3_U3416 , P3_U5255 );
nand NAND2_9176 ( P3_U5323 , P3_U5257 , P3_U3082 );
nand NAND2_9177 ( P3_U5324 , P3_U5440 , P3_U3083 );
nand NAND2_9178 ( P3_U5325 , P3_U3413 , P3_U5255 );
nand NAND2_9179 ( P3_U5326 , P3_U5257 , P3_U3083 );
nand NAND2_9180 ( P3_U5327 , P3_U5440 , P3_U3069 );
nand NAND2_9181 ( P3_U5328 , P3_U3410 , P3_U5255 );
nand NAND2_9182 ( P3_U5329 , P3_U5257 , P3_U3069 );
nand NAND2_9183 ( P3_U5330 , P3_U5440 , P3_U3070 );
nand NAND2_9184 ( P3_U5331 , P3_U3407 , P3_U5255 );
nand NAND2_9185 ( P3_U5332 , P3_U5257 , P3_U3070 );
nand NAND2_9186 ( P3_U5333 , P3_U5440 , P3_U3066 );
nand NAND2_9187 ( P3_U5334 , P3_U3404 , P3_U5255 );
nand NAND2_9188 ( P3_U5335 , P3_U5257 , P3_U3066 );
nand NAND2_9189 ( P3_U5336 , P3_U5440 , P3_U3059 );
nand NAND2_9190 ( P3_U5337 , P3_U3401 , P3_U5255 );
nand NAND2_9191 ( P3_U5338 , P3_U5257 , P3_U3059 );
nand NAND2_9192 ( P3_U5339 , P3_U5440 , P3_U3063 );
nand NAND2_9193 ( P3_U5340 , P3_U5257 , P3_U3055 );
nand NAND2_9194 ( P3_U5341 , P3_U3872 , P3_U5255 );
nand NAND2_9195 ( P3_U5342 , P3_U5257 , P3_U3058 );
nand NAND2_9196 ( P3_U5343 , P3_U3873 , P3_U5255 );
nand NAND2_9197 ( P3_U5344 , P3_U3398 , P3_U5255 );
nand NAND2_9198 ( P3_U5345 , P3_U5257 , P3_U3063 );
nand NAND2_9199 ( P3_U5346 , P3_U5440 , P3_U3067 );
nand NAND2_9200 ( P3_U5347 , P3_U5257 , P3_U3054 );
nand NAND2_9201 ( P3_U5348 , P3_U3908 , P3_U5255 );
nand NAND2_9202 ( P3_U5349 , P3_U5440 , P3_U3053 );
nand NAND2_9203 ( P3_U5350 , P3_U5257 , P3_U3053 );
nand NAND2_9204 ( P3_U5351 , P3_U3899 , P3_U5255 );
nand NAND2_9205 ( P3_U5352 , P3_U5440 , P3_U3052 );
nand NAND2_9206 ( P3_U5353 , P3_U5257 , P3_U3052 );
nand NAND2_9207 ( P3_U5354 , P3_U3900 , P3_U5255 );
nand NAND2_9208 ( P3_U5355 , P3_U5440 , P3_U3056 );
nand NAND2_9209 ( P3_U5356 , P3_U5257 , P3_U3056 );
nand NAND2_9210 ( P3_U5357 , P3_U3901 , P3_U5255 );
nand NAND2_9211 ( P3_U5358 , P3_U5440 , P3_U3057 );
nand NAND2_9212 ( P3_U5359 , P3_U5257 , P3_U3057 );
nand NAND2_9213 ( P3_U5360 , P3_U3902 , P3_U5255 );
nand NAND2_9214 ( P3_U5361 , P3_U5440 , P3_U3064 );
nand NAND2_9215 ( P3_U5362 , P3_U5257 , P3_U3064 );
nand NAND2_9216 ( P3_U5363 , P3_U3903 , P3_U5255 );
nand NAND2_9217 ( P3_U5364 , P3_U5440 , P3_U3065 );
nand NAND2_9218 ( P3_U5365 , P3_U5257 , P3_U3065 );
nand NAND2_9219 ( P3_U5366 , P3_U3904 , P3_U5255 );
nand NAND2_9220 ( P3_U5367 , P3_U5440 , P3_U3060 );
nand NAND2_9221 ( P3_U5368 , P3_U5257 , P3_U3060 );
nand NAND2_9222 ( P3_U5369 , P3_U3905 , P3_U5255 );
nand NAND2_9223 ( P3_U5370 , P3_U5440 , P3_U3074 );
nand NAND2_9224 ( P3_U5371 , P3_U5257 , P3_U3074 );
nand NAND2_9225 ( P3_U5372 , P3_U3906 , P3_U5255 );
nand NAND2_9226 ( P3_U5373 , P3_U5440 , P3_U3075 );
nand NAND2_9227 ( P3_U5374 , P3_U5257 , P3_U3075 );
nand NAND2_9228 ( P3_U5375 , P3_U3907 , P3_U5255 );
nand NAND2_9229 ( P3_U5376 , P3_U5440 , P3_U3080 );
nand NAND2_9230 ( P3_U5377 , P3_U3395 , P3_U5255 );
nand NAND2_9231 ( P3_U5378 , P3_U5257 , P3_U3067 );
nand NAND2_9232 ( P3_U5379 , P3_U5440 , P3_U3077 );
nand NAND2_9233 ( P3_U5380 , P3_U3445 , P3_U5255 );
nand NAND2_9234 ( P3_U5381 , P3_U5257 , P3_U3080 );
nand NAND2_9235 ( P3_U5382 , P3_U5440 , P3_U3081 );
nand NAND2_9236 ( P3_U5383 , P3_U3443 , P3_U5255 );
nand NAND2_9237 ( P3_U5384 , P3_U5257 , P3_U3081 );
nand NAND2_9238 ( P3_U5385 , P3_U5440 , P3_U3068 );
nand NAND2_9239 ( P3_U5386 , P3_U3440 , P3_U5255 );
nand NAND2_9240 ( P3_U5387 , P3_U5257 , P3_U3068 );
nand NAND2_9241 ( P3_U5388 , P3_U5440 , P3_U3072 );
nand NAND2_9242 ( P3_U5389 , P3_U3437 , P3_U5255 );
nand NAND2_9243 ( P3_U5390 , P3_U5257 , P3_U3072 );
nand NAND2_9244 ( P3_U5391 , P3_U5440 , P3_U3073 );
nand NAND2_9245 ( P3_U5392 , P3_U3434 , P3_U5255 );
nand NAND2_9246 ( P3_U5393 , P3_U5257 , P3_U3073 );
nand NAND2_9247 ( P3_U5394 , P3_U5440 , P3_U3078 );
nand NAND2_9248 ( P3_U5395 , P3_U3431 , P3_U5255 );
nand NAND2_9249 ( P3_U5396 , P3_U5257 , P3_U3078 );
nand NAND2_9250 ( P3_U5397 , P3_U5440 , P3_U3079 );
nand NAND2_9251 ( P3_U5398 , P3_U3428 , P3_U5255 );
nand NAND2_9252 ( P3_U5399 , P3_U5257 , P3_U3079 );
nand NAND2_9253 ( P3_U5400 , P3_U5440 , P3_U3071 );
nand NAND2_9254 ( P3_U5401 , P3_U3425 , P3_U5255 );
nand NAND2_9255 ( P3_U5402 , P3_U5257 , P3_U3071 );
nand NAND2_9256 ( P3_U5403 , P3_U5440 , P3_U3062 );
nand NAND2_9257 ( P3_U5404 , P3_U3422 , P3_U5255 );
nand NAND2_9258 ( P3_U5405 , P3_U5257 , P3_U3062 );
nand NAND2_9259 ( P3_U5406 , P3_U5440 , P3_U3061 );
nand NAND2_9260 ( P3_U5407 , P3_U3419 , P3_U5255 );
nand NAND2_9261 ( P3_U5408 , P3_U5257 , P3_U3061 );
nand NAND2_9262 ( P3_U5409 , P3_U5440 , P3_U3082 );
nand NAND2_9263 ( P3_U5410 , P3_U3392 , P3_U5255 );
nand NAND2_9264 ( P3_U5411 , P3_U5257 , P3_U3077 );
nand NAND2_9265 ( P3_U5412 , P3_U5440 , P3_U3076 );
nand NAND2_9266 ( P3_U5413 , P3_U3387 , P3_U5255 );
nand NAND2_9267 ( P3_U5414 , P3_U5257 , P3_U3076 );
nand NAND2_9268 ( P3_U5415 , P3_U4981 , P3_U3151 );
nand NAND3_9269 ( P3_U5416 , P3_U4981 , P3_U5440 , P3_U4980 );
nand NAND2_9270 ( P3_U5417 , P3_U3043 , P3_U3303 );
nand NAND2_9271 ( P3_U5418 , P3_U3043 , P3_U3894 );
not NOT1_9272 ( P3_U5419 , P3_U3371 );
nand NAND2_9273 ( P3_U5420 , P3_U5418 , P3_U3918 );
nand NAND3_9274 ( P3_U5421 , P3_U5938 , P3_U5937 , P3_U3774 );
nand NAND2_9275 ( P3_U5422 , P3_U5434 , P3_U5428 );
nand NAND2_9276 ( P3_U5423 , P3_U3879 , P3_U3378 );
nand NAND2_9277 ( P3_U5424 , P3_U3375 , P3_U3833 );
nand NAND2_9278 ( P3_U5425 , P3_U3876 , P3_U5447 );
nand NAND2_9279 ( P3_U5426 , P3_IR_REG_24_ , P3_U3831 );
nand NAND2_9280 ( P3_U5427 , P3_IR_REG_31_ , P3_SUB_598_U18 );
not NOT1_9281 ( P3_U5428 , P3_U3372 );
nand NAND2_9282 ( P3_U5429 , P3_IR_REG_25_ , P3_U3831 );
nand NAND2_9283 ( P3_U5430 , P3_IR_REG_31_ , P3_SUB_598_U81 );
not NOT1_9284 ( P3_U5431 , P3_U3373 );
nand NAND2_9285 ( P3_U5432 , P3_IR_REG_26_ , P3_U3831 );
nand NAND2_9286 ( P3_U5433 , P3_IR_REG_31_ , P3_SUB_598_U19 );
not NOT1_9287 ( P3_U5434 , P3_U3374 );
nand NAND2_9288 ( P3_U5435 , P3_U5428 , P3_B_REG );
nand NAND2_9289 ( P3_U5436 , P3_U3372 , P3_U3298 );
nand NAND2_9290 ( P3_U5437 , P3_U5436 , P3_U5435 );
nand NAND2_9291 ( P3_U5438 , P3_IR_REG_23_ , P3_U3831 );
nand NAND2_9292 ( P3_U5439 , P3_IR_REG_31_ , P3_SUB_598_U17 );
not NOT1_9293 ( P3_U5440 , P3_U3375 );
nand NAND2_9294 ( P3_U5441 , P3_D_REG_0_ , P3_U3832 );
nand NAND2_9295 ( P3_U5442 , P3_U3915 , P3_U4020 );
nand NAND2_9296 ( P3_U5443 , P3_D_REG_1_ , P3_U3832 );
nand NAND2_9297 ( P3_U5444 , P3_U3915 , P3_U4021 );
nand NAND2_9298 ( P3_U5445 , P3_IR_REG_20_ , P3_U3831 );
nand NAND2_9299 ( P3_U5446 , P3_IR_REG_31_ , P3_SUB_598_U15 );
not NOT1_9300 ( P3_U5447 , P3_U3378 );
nand NAND2_9301 ( P3_U5448 , P3_IR_REG_19_ , P3_U3831 );
nand NAND2_9302 ( P3_U5449 , P3_IR_REG_31_ , P3_SUB_598_U14 );
not NOT1_9303 ( P3_U5450 , P3_U3379 );
nand NAND2_9304 ( P3_U5451 , P3_IR_REG_22_ , P3_U3831 );
nand NAND2_9305 ( P3_U5452 , P3_IR_REG_31_ , P3_SUB_598_U16 );
not NOT1_9306 ( P3_U5453 , P3_U3380 );
nand NAND2_9307 ( P3_U5454 , P3_IR_REG_21_ , P3_U3831 );
nand NAND2_9308 ( P3_U5455 , P3_IR_REG_31_ , P3_SUB_598_U83 );
not NOT1_9309 ( P3_U5456 , P3_U3385 );
nand NAND2_9310 ( P3_U5457 , P3_IR_REG_30_ , P3_U3831 );
nand NAND2_9311 ( P3_U5458 , P3_IR_REG_31_ , P3_SUB_598_U77 );
not NOT1_9312 ( P3_U5459 , P3_U3381 );
nand NAND2_9313 ( P3_U5460 , P3_IR_REG_29_ , P3_U3831 );
nand NAND2_9314 ( P3_U5461 , P3_IR_REG_31_ , P3_SUB_598_U21 );
not NOT1_9315 ( P3_U5462 , P3_U3382 );
nand NAND2_9316 ( P3_U5463 , P3_IR_REG_28_ , P3_U3831 );
nand NAND2_9317 ( P3_U5464 , P3_IR_REG_31_ , P3_SUB_598_U20 );
not NOT1_9318 ( P3_U5465 , P3_U3383 );
nand NAND2_9319 ( P3_U5466 , P3_IR_REG_27_ , P3_U3831 );
nand NAND2_9320 ( P3_U5467 , P3_IR_REG_31_ , P3_SUB_598_U79 );
not NOT1_9321 ( P3_U5468 , P3_U3384 );
nand NAND2_9322 ( P3_U5469 , P3_IR_REG_0_ , P3_U3831 );
nand NAND2_9323 ( P3_U5470 , P3_IR_REG_31_ , P3_IR_REG_0_ );
nand NAND2_9324 ( P3_U5471 , U61 , P3_U3833 );
nand NAND2_9325 ( P3_U5472 , P3_U3893 , P3_U3386 );
not NOT1_9326 ( P3_U5473 , P3_U3387 );
nand NAND2_9327 ( P3_U5474 , P3_U5422 , P3_U3300 );
nand NAND2_9328 ( P3_U5475 , P3_D_REG_0_ , P3_U4019 );
not NOT1_9329 ( P3_U5476 , P3_U3388 );
nand NAND2_9330 ( P3_U5477 , P3_D_REG_1_ , P3_U4019 );
nand NAND2_9331 ( P3_U5478 , P3_U4021 , P3_U3300 );
not NOT1_9332 ( P3_U5479 , P3_U3389 );
nand NAND2_9333 ( P3_U5480 , P3_U4052 , P3_U5453 );
nand NAND2_9334 ( P3_U5481 , P3_U3380 , P3_U3834 );
nand NAND2_9335 ( P3_U5482 , P3_U5481 , P3_U5480 );
nand NAND2_9336 ( P3_U5483 , P3_REG0_REG_0_ , P3_U3835 );
nand NAND2_9337 ( P3_U5484 , P3_U3914 , P3_U4077 );
nand NAND2_9338 ( P3_U5485 , P3_IR_REG_1_ , P3_U3831 );
nand NAND2_9339 ( P3_U5486 , P3_IR_REG_31_ , P3_SUB_598_U51 );
nand NAND2_9340 ( P3_U5487 , U50 , P3_U3833 );
nand NAND2_9341 ( P3_U5488 , P3_U3391 , P3_U3893 );
not NOT1_9342 ( P3_U5489 , P3_U3392 );
nand NAND2_9343 ( P3_U5490 , P3_REG0_REG_1_ , P3_U3835 );
nand NAND2_9344 ( P3_U5491 , P3_U3914 , P3_U4102 );
nand NAND2_9345 ( P3_U5492 , P3_IR_REG_2_ , P3_U3831 );
nand NAND2_9346 ( P3_U5493 , P3_IR_REG_31_ , P3_SUB_598_U22 );
nand NAND2_9347 ( P3_U5494 , U39 , P3_U3833 );
nand NAND2_9348 ( P3_U5495 , P3_U3394 , P3_U3893 );
not NOT1_9349 ( P3_U5496 , P3_U3395 );
nand NAND2_9350 ( P3_U5497 , P3_REG0_REG_2_ , P3_U3835 );
nand NAND2_9351 ( P3_U5498 , P3_U3914 , P3_U4120 );
nand NAND2_9352 ( P3_U5499 , P3_IR_REG_3_ , P3_U3831 );
nand NAND2_9353 ( P3_U5500 , P3_IR_REG_31_ , P3_SUB_598_U23 );
nand NAND2_9354 ( P3_U5501 , U36 , P3_U3833 );
nand NAND2_9355 ( P3_U5502 , P3_U3397 , P3_U3893 );
not NOT1_9356 ( P3_U5503 , P3_U3398 );
nand NAND2_9357 ( P3_U5504 , P3_REG0_REG_3_ , P3_U3835 );
nand NAND2_9358 ( P3_U5505 , P3_U3914 , P3_U4138 );
nand NAND2_9359 ( P3_U5506 , P3_IR_REG_4_ , P3_U3831 );
nand NAND2_9360 ( P3_U5507 , P3_IR_REG_31_ , P3_SUB_598_U24 );
nand NAND2_9361 ( P3_U5508 , U35 , P3_U3833 );
nand NAND2_9362 ( P3_U5509 , P3_U3400 , P3_U3893 );
not NOT1_9363 ( P3_U5510 , P3_U3401 );
nand NAND2_9364 ( P3_U5511 , P3_REG0_REG_4_ , P3_U3835 );
nand NAND2_9365 ( P3_U5512 , P3_U3914 , P3_U4156 );
nand NAND2_9366 ( P3_U5513 , P3_IR_REG_5_ , P3_U3831 );
nand NAND2_9367 ( P3_U5514 , P3_IR_REG_31_ , P3_SUB_598_U74 );
nand NAND2_9368 ( P3_U5515 , U34 , P3_U3833 );
nand NAND2_9369 ( P3_U5516 , P3_U3403 , P3_U3893 );
not NOT1_9370 ( P3_U5517 , P3_U3404 );
nand NAND2_9371 ( P3_U5518 , P3_REG0_REG_5_ , P3_U3835 );
nand NAND2_9372 ( P3_U5519 , P3_U3914 , P3_U4174 );
nand NAND2_9373 ( P3_U5520 , P3_IR_REG_6_ , P3_U3831 );
nand NAND2_9374 ( P3_U5521 , P3_IR_REG_31_ , P3_SUB_598_U25 );
nand NAND2_9375 ( P3_U5522 , U33 , P3_U3833 );
nand NAND2_9376 ( P3_U5523 , P3_U3406 , P3_U3893 );
not NOT1_9377 ( P3_U5524 , P3_U3407 );
nand NAND2_9378 ( P3_U5525 , P3_REG0_REG_6_ , P3_U3835 );
nand NAND2_9379 ( P3_U5526 , P3_U3914 , P3_U4192 );
nand NAND2_9380 ( P3_U5527 , P3_IR_REG_7_ , P3_U3831 );
nand NAND2_9381 ( P3_U5528 , P3_IR_REG_31_ , P3_SUB_598_U26 );
nand NAND2_9382 ( P3_U5529 , U32 , P3_U3833 );
nand NAND2_9383 ( P3_U5530 , P3_U3409 , P3_U3893 );
not NOT1_9384 ( P3_U5531 , P3_U3410 );
nand NAND2_9385 ( P3_U5532 , P3_REG0_REG_7_ , P3_U3835 );
nand NAND2_9386 ( P3_U5533 , P3_U3914 , P3_U4210 );
nand NAND2_9387 ( P3_U5534 , P3_IR_REG_8_ , P3_U3831 );
nand NAND2_9388 ( P3_U5535 , P3_IR_REG_31_ , P3_SUB_598_U27 );
nand NAND2_9389 ( P3_U5536 , U31 , P3_U3833 );
nand NAND2_9390 ( P3_U5537 , P3_U3412 , P3_U3893 );
not NOT1_9391 ( P3_U5538 , P3_U3413 );
nand NAND2_9392 ( P3_U5539 , P3_REG0_REG_8_ , P3_U3835 );
nand NAND2_9393 ( P3_U5540 , P3_U3914 , P3_U4228 );
nand NAND2_9394 ( P3_U5541 , P3_IR_REG_9_ , P3_U3831 );
nand NAND2_9395 ( P3_U5542 , P3_IR_REG_31_ , P3_SUB_598_U72 );
nand NAND2_9396 ( P3_U5543 , U30 , P3_U3833 );
nand NAND2_9397 ( P3_U5544 , P3_U3415 , P3_U3893 );
not NOT1_9398 ( P3_U5545 , P3_U3416 );
nand NAND2_9399 ( P3_U5546 , P3_REG0_REG_9_ , P3_U3835 );
nand NAND2_9400 ( P3_U5547 , P3_U3914 , P3_U4246 );
nand NAND2_9401 ( P3_U5548 , P3_IR_REG_10_ , P3_U3831 );
nand NAND2_9402 ( P3_U5549 , P3_IR_REG_31_ , P3_SUB_598_U7 );
nand NAND2_9403 ( P3_U5550 , U60 , P3_U3833 );
nand NAND2_9404 ( P3_U5551 , P3_U3418 , P3_U3893 );
not NOT1_9405 ( P3_U5552 , P3_U3419 );
nand NAND2_9406 ( P3_U5553 , P3_REG0_REG_10_ , P3_U3835 );
nand NAND2_9407 ( P3_U5554 , P3_U3914 , P3_U4264 );
nand NAND2_9408 ( P3_U5555 , P3_IR_REG_11_ , P3_U3831 );
nand NAND2_9409 ( P3_U5556 , P3_IR_REG_31_ , P3_SUB_598_U8 );
nand NAND2_9410 ( P3_U5557 , U59 , P3_U3833 );
nand NAND2_9411 ( P3_U5558 , P3_U3421 , P3_U3893 );
not NOT1_9412 ( P3_U5559 , P3_U3422 );
nand NAND2_9413 ( P3_U5560 , P3_REG0_REG_11_ , P3_U3835 );
nand NAND2_9414 ( P3_U5561 , P3_U3914 , P3_U4282 );
nand NAND2_9415 ( P3_U5562 , P3_IR_REG_12_ , P3_U3831 );
nand NAND2_9416 ( P3_U5563 , P3_IR_REG_31_ , P3_SUB_598_U9 );
nand NAND2_9417 ( P3_U5564 , U58 , P3_U3833 );
nand NAND2_9418 ( P3_U5565 , P3_U3424 , P3_U3893 );
not NOT1_9419 ( P3_U5566 , P3_U3425 );
nand NAND2_9420 ( P3_U5567 , P3_REG0_REG_12_ , P3_U3835 );
nand NAND2_9421 ( P3_U5568 , P3_U3914 , P3_U4300 );
nand NAND2_9422 ( P3_U5569 , P3_IR_REG_13_ , P3_U3831 );
nand NAND2_9423 ( P3_U5570 , P3_IR_REG_31_ , P3_SUB_598_U89 );
nand NAND2_9424 ( P3_U5571 , U57 , P3_U3833 );
nand NAND2_9425 ( P3_U5572 , P3_U3427 , P3_U3893 );
not NOT1_9426 ( P3_U5573 , P3_U3428 );
nand NAND2_9427 ( P3_U5574 , P3_REG0_REG_13_ , P3_U3835 );
nand NAND2_9428 ( P3_U5575 , P3_U3914 , P3_U4318 );
nand NAND2_9429 ( P3_U5576 , P3_IR_REG_14_ , P3_U3831 );
nand NAND2_9430 ( P3_U5577 , P3_IR_REG_31_ , P3_SUB_598_U10 );
nand NAND2_9431 ( P3_U5578 , U56 , P3_U3833 );
nand NAND2_9432 ( P3_U5579 , P3_U3430 , P3_U3893 );
not NOT1_9433 ( P3_U5580 , P3_U3431 );
nand NAND2_9434 ( P3_U5581 , P3_REG0_REG_14_ , P3_U3835 );
nand NAND2_9435 ( P3_U5582 , P3_U3914 , P3_U4336 );
nand NAND2_9436 ( P3_U5583 , P3_IR_REG_15_ , P3_U3831 );
nand NAND2_9437 ( P3_U5584 , P3_IR_REG_31_ , P3_SUB_598_U11 );
nand NAND2_9438 ( P3_U5585 , U55 , P3_U3833 );
nand NAND2_9439 ( P3_U5586 , P3_U3433 , P3_U3893 );
not NOT1_9440 ( P3_U5587 , P3_U3434 );
nand NAND2_9441 ( P3_U5588 , P3_REG0_REG_15_ , P3_U3835 );
nand NAND2_9442 ( P3_U5589 , P3_U3914 , P3_U4354 );
nand NAND2_9443 ( P3_U5590 , P3_IR_REG_16_ , P3_U3831 );
nand NAND2_9444 ( P3_U5591 , P3_IR_REG_31_ , P3_SUB_598_U12 );
nand NAND2_9445 ( P3_U5592 , U54 , P3_U3833 );
nand NAND2_9446 ( P3_U5593 , P3_U3436 , P3_U3893 );
not NOT1_9447 ( P3_U5594 , P3_U3437 );
nand NAND2_9448 ( P3_U5595 , P3_REG0_REG_16_ , P3_U3835 );
nand NAND2_9449 ( P3_U5596 , P3_U3914 , P3_U4372 );
nand NAND2_9450 ( P3_U5597 , P3_IR_REG_17_ , P3_U3831 );
nand NAND2_9451 ( P3_U5598 , P3_IR_REG_31_ , P3_SUB_598_U87 );
nand NAND2_9452 ( P3_U5599 , U53 , P3_U3833 );
nand NAND2_9453 ( P3_U5600 , P3_U3439 , P3_U3893 );
not NOT1_9454 ( P3_U5601 , P3_U3440 );
nand NAND2_9455 ( P3_U5602 , P3_REG0_REG_17_ , P3_U3835 );
nand NAND2_9456 ( P3_U5603 , P3_U3914 , P3_U4390 );
nand NAND2_9457 ( P3_U5604 , P3_IR_REG_18_ , P3_U3831 );
nand NAND2_9458 ( P3_U5605 , P3_IR_REG_31_ , P3_SUB_598_U13 );
nand NAND2_9459 ( P3_U5606 , U52 , P3_U3833 );
nand NAND2_9460 ( P3_U5607 , P3_U3442 , P3_U3893 );
not NOT1_9461 ( P3_U5608 , P3_U3443 );
nand NAND2_9462 ( P3_U5609 , P3_REG0_REG_18_ , P3_U3835 );
nand NAND2_9463 ( P3_U5610 , P3_U3914 , P3_U4408 );
nand NAND2_9464 ( P3_U5611 , U51 , P3_U3833 );
nand NAND2_9465 ( P3_U5612 , P3_U3893 , P3_U3379 );
not NOT1_9466 ( P3_U5613 , P3_U3445 );
nand NAND2_9467 ( P3_U5614 , P3_REG0_REG_19_ , P3_U3835 );
nand NAND2_9468 ( P3_U5615 , P3_U3914 , P3_U4426 );
nand NAND2_9469 ( P3_U5616 , P3_REG0_REG_20_ , P3_U3835 );
nand NAND2_9470 ( P3_U5617 , P3_U3914 , P3_U4444 );
nand NAND2_9471 ( P3_U5618 , P3_REG0_REG_21_ , P3_U3835 );
nand NAND2_9472 ( P3_U5619 , P3_U3914 , P3_U4462 );
nand NAND2_9473 ( P3_U5620 , P3_REG0_REG_22_ , P3_U3835 );
nand NAND2_9474 ( P3_U5621 , P3_U3914 , P3_U4480 );
nand NAND2_9475 ( P3_U5622 , P3_REG0_REG_23_ , P3_U3835 );
nand NAND2_9476 ( P3_U5623 , P3_U3914 , P3_U4498 );
nand NAND2_9477 ( P3_U5624 , P3_REG0_REG_24_ , P3_U3835 );
nand NAND2_9478 ( P3_U5625 , P3_U3914 , P3_U4516 );
nand NAND2_9479 ( P3_U5626 , P3_REG0_REG_25_ , P3_U3835 );
nand NAND2_9480 ( P3_U5627 , P3_U3914 , P3_U4534 );
nand NAND2_9481 ( P3_U5628 , P3_REG0_REG_26_ , P3_U3835 );
nand NAND2_9482 ( P3_U5629 , P3_U3914 , P3_U4552 );
nand NAND2_9483 ( P3_U5630 , P3_REG0_REG_27_ , P3_U3835 );
nand NAND2_9484 ( P3_U5631 , P3_U3914 , P3_U4570 );
nand NAND2_9485 ( P3_U5632 , P3_REG0_REG_28_ , P3_U3835 );
nand NAND2_9486 ( P3_U5633 , P3_U3914 , P3_U4588 );
nand NAND2_9487 ( P3_U5634 , P3_REG0_REG_29_ , P3_U3835 );
nand NAND2_9488 ( P3_U5635 , P3_U3914 , P3_U4608 );
nand NAND2_9489 ( P3_U5636 , P3_REG0_REG_30_ , P3_U3835 );
nand NAND2_9490 ( P3_U5637 , P3_U3914 , P3_U4615 );
nand NAND2_9491 ( P3_U5638 , P3_REG0_REG_31_ , P3_U3835 );
nand NAND2_9492 ( P3_U5639 , P3_U3914 , P3_U4617 );
nand NAND2_9493 ( P3_U5640 , P3_U5453 , P3_U3834 );
nand NAND2_9494 ( P3_U5641 , P3_U4052 , P3_U5450 );
nand NAND2_9495 ( P3_U5642 , P3_REG1_REG_0_ , P3_U3836 );
nand NAND2_9496 ( P3_U5643 , P3_U3913 , P3_U4077 );
nand NAND2_9497 ( P3_U5644 , P3_REG1_REG_1_ , P3_U3836 );
nand NAND2_9498 ( P3_U5645 , P3_U3913 , P3_U4102 );
nand NAND2_9499 ( P3_U5646 , P3_REG1_REG_2_ , P3_U3836 );
nand NAND2_9500 ( P3_U5647 , P3_U3913 , P3_U4120 );
nand NAND2_9501 ( P3_U5648 , P3_REG1_REG_3_ , P3_U3836 );
nand NAND2_9502 ( P3_U5649 , P3_U3913 , P3_U4138 );
nand NAND2_9503 ( P3_U5650 , P3_REG1_REG_4_ , P3_U3836 );
nand NAND2_9504 ( P3_U5651 , P3_U3913 , P3_U4156 );
nand NAND2_9505 ( P3_U5652 , P3_REG1_REG_5_ , P3_U3836 );
nand NAND2_9506 ( P3_U5653 , P3_U3913 , P3_U4174 );
nand NAND2_9507 ( P3_U5654 , P3_REG1_REG_6_ , P3_U3836 );
nand NAND2_9508 ( P3_U5655 , P3_U3913 , P3_U4192 );
nand NAND2_9509 ( P3_U5656 , P3_REG1_REG_7_ , P3_U3836 );
nand NAND2_9510 ( P3_U5657 , P3_U3913 , P3_U4210 );
nand NAND2_9511 ( P3_U5658 , P3_REG1_REG_8_ , P3_U3836 );
nand NAND2_9512 ( P3_U5659 , P3_U3913 , P3_U4228 );
nand NAND2_9513 ( P3_U5660 , P3_REG1_REG_9_ , P3_U3836 );
nand NAND2_9514 ( P3_U5661 , P3_U3913 , P3_U4246 );
nand NAND2_9515 ( P3_U5662 , P3_REG1_REG_10_ , P3_U3836 );
nand NAND2_9516 ( P3_U5663 , P3_U3913 , P3_U4264 );
nand NAND2_9517 ( P3_U5664 , P3_REG1_REG_11_ , P3_U3836 );
nand NAND2_9518 ( P3_U5665 , P3_U3913 , P3_U4282 );
nand NAND2_9519 ( P3_U5666 , P3_REG1_REG_12_ , P3_U3836 );
nand NAND2_9520 ( P3_U5667 , P3_U3913 , P3_U4300 );
nand NAND2_9521 ( P3_U5668 , P3_REG1_REG_13_ , P3_U3836 );
nand NAND2_9522 ( P3_U5669 , P3_U3913 , P3_U4318 );
nand NAND2_9523 ( P3_U5670 , P3_REG1_REG_14_ , P3_U3836 );
nand NAND2_9524 ( P3_U5671 , P3_U3913 , P3_U4336 );
nand NAND2_9525 ( P3_U5672 , P3_REG1_REG_15_ , P3_U3836 );
nand NAND2_9526 ( P3_U5673 , P3_U3913 , P3_U4354 );
nand NAND2_9527 ( P3_U5674 , P3_REG1_REG_16_ , P3_U3836 );
nand NAND2_9528 ( P3_U5675 , P3_U3913 , P3_U4372 );
nand NAND2_9529 ( P3_U5676 , P3_REG1_REG_17_ , P3_U3836 );
nand NAND2_9530 ( P3_U5677 , P3_U3913 , P3_U4390 );
nand NAND2_9531 ( P3_U5678 , P3_REG1_REG_18_ , P3_U3836 );
nand NAND2_9532 ( P3_U5679 , P3_U3913 , P3_U4408 );
nand NAND2_9533 ( P3_U5680 , P3_REG1_REG_19_ , P3_U3836 );
nand NAND2_9534 ( P3_U5681 , P3_U3913 , P3_U4426 );
nand NAND2_9535 ( P3_U5682 , P3_REG1_REG_20_ , P3_U3836 );
nand NAND2_9536 ( P3_U5683 , P3_U3913 , P3_U4444 );
nand NAND2_9537 ( P3_U5684 , P3_REG1_REG_21_ , P3_U3836 );
nand NAND2_9538 ( P3_U5685 , P3_U3913 , P3_U4462 );
nand NAND2_9539 ( P3_U5686 , P3_REG1_REG_22_ , P3_U3836 );
nand NAND2_9540 ( P3_U5687 , P3_U3913 , P3_U4480 );
nand NAND2_9541 ( P3_U5688 , P3_REG1_REG_23_ , P3_U3836 );
nand NAND2_9542 ( P3_U5689 , P3_U3913 , P3_U4498 );
nand NAND2_9543 ( P3_U5690 , P3_REG1_REG_24_ , P3_U3836 );
nand NAND2_9544 ( P3_U5691 , P3_U3913 , P3_U4516 );
nand NAND2_9545 ( P3_U5692 , P3_REG1_REG_25_ , P3_U3836 );
nand NAND2_9546 ( P3_U5693 , P3_U3913 , P3_U4534 );
nand NAND2_9547 ( P3_U5694 , P3_REG1_REG_26_ , P3_U3836 );
nand NAND2_9548 ( P3_U5695 , P3_U3913 , P3_U4552 );
nand NAND2_9549 ( P3_U5696 , P3_REG1_REG_27_ , P3_U3836 );
nand NAND2_9550 ( P3_U5697 , P3_U3913 , P3_U4570 );
nand NAND2_9551 ( P3_U5698 , P3_REG1_REG_28_ , P3_U3836 );
nand NAND2_9552 ( P3_U5699 , P3_U3913 , P3_U4588 );
nand NAND2_9553 ( P3_U5700 , P3_REG1_REG_29_ , P3_U3836 );
nand NAND2_9554 ( P3_U5701 , P3_U3913 , P3_U4608 );
nand NAND2_9555 ( P3_U5702 , P3_REG1_REG_30_ , P3_U3836 );
nand NAND2_9556 ( P3_U5703 , P3_U3913 , P3_U4615 );
nand NAND2_9557 ( P3_U5704 , P3_REG1_REG_31_ , P3_U3836 );
nand NAND2_9558 ( P3_U5705 , P3_U3913 , P3_U4617 );
nand NAND2_9559 ( P3_U5706 , P3_REG2_REG_0_ , P3_U3358 );
nand NAND2_9560 ( P3_U5707 , P3_U3912 , P3_U3314 );
nand NAND2_9561 ( P3_U5708 , P3_REG2_REG_1_ , P3_U3358 );
nand NAND2_9562 ( P3_U5709 , P3_U3912 , P3_U3315 );
nand NAND2_9563 ( P3_U5710 , P3_REG2_REG_2_ , P3_U3358 );
nand NAND2_9564 ( P3_U5711 , P3_U3912 , P3_U3316 );
nand NAND2_9565 ( P3_U5712 , P3_REG2_REG_3_ , P3_U3358 );
nand NAND2_9566 ( P3_U5713 , P3_U3912 , P3_U3317 );
nand NAND2_9567 ( P3_U5714 , P3_REG2_REG_4_ , P3_U3358 );
nand NAND2_9568 ( P3_U5715 , P3_U3912 , P3_U3318 );
nand NAND2_9569 ( P3_U5716 , P3_REG2_REG_5_ , P3_U3358 );
nand NAND2_9570 ( P3_U5717 , P3_U3912 , P3_U3319 );
nand NAND2_9571 ( P3_U5718 , P3_REG2_REG_6_ , P3_U3358 );
nand NAND2_9572 ( P3_U5719 , P3_U3912 , P3_U3320 );
nand NAND2_9573 ( P3_U5720 , P3_REG2_REG_7_ , P3_U3358 );
nand NAND2_9574 ( P3_U5721 , P3_U3912 , P3_U3321 );
nand NAND2_9575 ( P3_U5722 , P3_REG2_REG_8_ , P3_U3358 );
nand NAND2_9576 ( P3_U5723 , P3_U3912 , P3_U3322 );
nand NAND2_9577 ( P3_U5724 , P3_REG2_REG_9_ , P3_U3358 );
nand NAND2_9578 ( P3_U5725 , P3_U3912 , P3_U3323 );
nand NAND2_9579 ( P3_U5726 , P3_REG2_REG_10_ , P3_U3358 );
nand NAND2_9580 ( P3_U5727 , P3_U3912 , P3_U3324 );
nand NAND2_9581 ( P3_U5728 , P3_REG2_REG_11_ , P3_U3358 );
nand NAND2_9582 ( P3_U5729 , P3_U3912 , P3_U3325 );
nand NAND2_9583 ( P3_U5730 , P3_REG2_REG_12_ , P3_U3358 );
nand NAND2_9584 ( P3_U5731 , P3_U3912 , P3_U3326 );
nand NAND2_9585 ( P3_U5732 , P3_REG2_REG_13_ , P3_U3358 );
nand NAND2_9586 ( P3_U5733 , P3_U3912 , P3_U3327 );
nand NAND2_9587 ( P3_U5734 , P3_REG2_REG_14_ , P3_U3358 );
nand NAND2_9588 ( P3_U5735 , P3_U3912 , P3_U3328 );
nand NAND2_9589 ( P3_U5736 , P3_REG2_REG_15_ , P3_U3358 );
nand NAND2_9590 ( P3_U5737 , P3_U3912 , P3_U3329 );
nand NAND2_9591 ( P3_U5738 , P3_REG2_REG_16_ , P3_U3358 );
nand NAND2_9592 ( P3_U5739 , P3_U3912 , P3_U3330 );
nand NAND2_9593 ( P3_U5740 , P3_REG2_REG_17_ , P3_U3358 );
nand NAND2_9594 ( P3_U5741 , P3_U3912 , P3_U3331 );
nand NAND2_9595 ( P3_U5742 , P3_REG2_REG_18_ , P3_U3358 );
nand NAND2_9596 ( P3_U5743 , P3_U3912 , P3_U3332 );
nand NAND2_9597 ( P3_U5744 , P3_REG2_REG_19_ , P3_U3358 );
nand NAND2_9598 ( P3_U5745 , P3_U3912 , P3_U3333 );
nand NAND2_9599 ( P3_U5746 , P3_REG2_REG_20_ , P3_U3358 );
nand NAND2_9600 ( P3_U5747 , P3_U3912 , P3_U3335 );
nand NAND2_9601 ( P3_U5748 , P3_REG2_REG_21_ , P3_U3358 );
nand NAND2_9602 ( P3_U5749 , P3_U3912 , P3_U3337 );
nand NAND2_9603 ( P3_U5750 , P3_REG2_REG_22_ , P3_U3358 );
nand NAND2_9604 ( P3_U5751 , P3_U3912 , P3_U3339 );
nand NAND2_9605 ( P3_U5752 , P3_REG2_REG_23_ , P3_U3358 );
nand NAND2_9606 ( P3_U5753 , P3_U3912 , P3_U3341 );
nand NAND2_9607 ( P3_U5754 , P3_REG2_REG_24_ , P3_U3358 );
nand NAND2_9608 ( P3_U5755 , P3_U3912 , P3_U3343 );
nand NAND2_9609 ( P3_U5756 , P3_REG2_REG_25_ , P3_U3358 );
nand NAND2_9610 ( P3_U5757 , P3_U3912 , P3_U3345 );
nand NAND2_9611 ( P3_U5758 , P3_REG2_REG_26_ , P3_U3358 );
nand NAND2_9612 ( P3_U5759 , P3_U3912 , P3_U3347 );
nand NAND2_9613 ( P3_U5760 , P3_REG2_REG_27_ , P3_U3358 );
nand NAND2_9614 ( P3_U5761 , P3_U3912 , P3_U3349 );
nand NAND2_9615 ( P3_U5762 , P3_REG2_REG_28_ , P3_U3358 );
nand NAND2_9616 ( P3_U5763 , P3_U3912 , P3_U3351 );
nand NAND2_9617 ( P3_U5764 , P3_REG2_REG_29_ , P3_U3358 );
nand NAND2_9618 ( P3_U5765 , P3_U3912 , P3_U3354 );
nand NAND2_9619 ( P3_U5766 , P3_U5465 , P3_U3024 );
nand NAND2_9620 ( P3_U5767 , P3_U3383 , P3_U3897 );
nand NAND2_9621 ( P3_U5768 , P3_U5767 , P3_U5766 );
nand NAND2_9622 ( P3_U5769 , P3_DATAO_REG_0_ , P3_U3363 );
nand NAND2_9623 ( P3_U5770 , P3_U3897 , P3_U3076 );
nand NAND2_9624 ( P3_U5771 , P3_DATAO_REG_1_ , P3_U3363 );
nand NAND2_9625 ( P3_U5772 , P3_U3897 , P3_U3077 );
nand NAND2_9626 ( P3_U5773 , P3_DATAO_REG_2_ , P3_U3363 );
nand NAND2_9627 ( P3_U5774 , P3_U3897 , P3_U3067 );
nand NAND2_9628 ( P3_U5775 , P3_DATAO_REG_3_ , P3_U3363 );
nand NAND2_9629 ( P3_U5776 , P3_U3897 , P3_U3063 );
nand NAND2_9630 ( P3_U5777 , P3_DATAO_REG_4_ , P3_U3363 );
nand NAND2_9631 ( P3_U5778 , P3_U3897 , P3_U3059 );
nand NAND2_9632 ( P3_U5779 , P3_DATAO_REG_5_ , P3_U3363 );
nand NAND2_9633 ( P3_U5780 , P3_U3897 , P3_U3066 );
nand NAND2_9634 ( P3_U5781 , P3_DATAO_REG_6_ , P3_U3363 );
nand NAND2_9635 ( P3_U5782 , P3_U3897 , P3_U3070 );
nand NAND2_9636 ( P3_U5783 , P3_DATAO_REG_7_ , P3_U3363 );
nand NAND2_9637 ( P3_U5784 , P3_U3897 , P3_U3069 );
nand NAND2_9638 ( P3_U5785 , P3_DATAO_REG_8_ , P3_U3363 );
nand NAND2_9639 ( P3_U5786 , P3_U3897 , P3_U3083 );
nand NAND2_9640 ( P3_U5787 , P3_DATAO_REG_9_ , P3_U3363 );
nand NAND2_9641 ( P3_U5788 , P3_U3897 , P3_U3082 );
nand NAND2_9642 ( P3_U5789 , P3_DATAO_REG_10_ , P3_U3363 );
nand NAND2_9643 ( P3_U5790 , P3_U3897 , P3_U3061 );
nand NAND2_9644 ( P3_U5791 , P3_DATAO_REG_11_ , P3_U3363 );
nand NAND2_9645 ( P3_U5792 , P3_U3897 , P3_U3062 );
nand NAND2_9646 ( P3_U5793 , P3_DATAO_REG_12_ , P3_U3363 );
nand NAND2_9647 ( P3_U5794 , P3_U3897 , P3_U3071 );
nand NAND2_9648 ( P3_U5795 , P3_DATAO_REG_13_ , P3_U3363 );
nand NAND2_9649 ( P3_U5796 , P3_U3897 , P3_U3079 );
nand NAND2_9650 ( P3_U5797 , P3_DATAO_REG_14_ , P3_U3363 );
nand NAND2_9651 ( P3_U5798 , P3_U3897 , P3_U3078 );
nand NAND2_9652 ( P3_U5799 , P3_DATAO_REG_15_ , P3_U3363 );
nand NAND2_9653 ( P3_U5800 , P3_U3897 , P3_U3073 );
nand NAND2_9654 ( P3_U5801 , P3_DATAO_REG_16_ , P3_U3363 );
nand NAND2_9655 ( P3_U5802 , P3_U3897 , P3_U3072 );
nand NAND2_9656 ( P3_U5803 , P3_DATAO_REG_17_ , P3_U3363 );
nand NAND2_9657 ( P3_U5804 , P3_U3897 , P3_U3068 );
nand NAND2_9658 ( P3_U5805 , P3_DATAO_REG_18_ , P3_U3363 );
nand NAND2_9659 ( P3_U5806 , P3_U3897 , P3_U3081 );
nand NAND2_9660 ( P3_U5807 , P3_DATAO_REG_19_ , P3_U3363 );
nand NAND2_9661 ( P3_U5808 , P3_U3897 , P3_U3080 );
nand NAND2_9662 ( P3_U5809 , P3_DATAO_REG_20_ , P3_U3363 );
nand NAND2_9663 ( P3_U5810 , P3_U3897 , P3_U3075 );
nand NAND2_9664 ( P3_U5811 , P3_DATAO_REG_21_ , P3_U3363 );
nand NAND2_9665 ( P3_U5812 , P3_U3897 , P3_U3074 );
nand NAND2_9666 ( P3_U5813 , P3_DATAO_REG_22_ , P3_U3363 );
nand NAND2_9667 ( P3_U5814 , P3_U3897 , P3_U3060 );
nand NAND2_9668 ( P3_U5815 , P3_DATAO_REG_23_ , P3_U3363 );
nand NAND2_9669 ( P3_U5816 , P3_U3897 , P3_U3065 );
nand NAND2_9670 ( P3_U5817 , P3_DATAO_REG_24_ , P3_U3363 );
nand NAND2_9671 ( P3_U5818 , P3_U3897 , P3_U3064 );
nand NAND2_9672 ( P3_U5819 , P3_DATAO_REG_25_ , P3_U3363 );
nand NAND2_9673 ( P3_U5820 , P3_U3897 , P3_U3057 );
nand NAND2_9674 ( P3_U5821 , P3_DATAO_REG_26_ , P3_U3363 );
nand NAND2_9675 ( P3_U5822 , P3_U3897 , P3_U3056 );
nand NAND2_9676 ( P3_U5823 , P3_DATAO_REG_27_ , P3_U3363 );
nand NAND2_9677 ( P3_U5824 , P3_U3897 , P3_U3052 );
nand NAND2_9678 ( P3_U5825 , P3_DATAO_REG_28_ , P3_U3363 );
nand NAND2_9679 ( P3_U5826 , P3_U3897 , P3_U3053 );
nand NAND2_9680 ( P3_U5827 , P3_DATAO_REG_29_ , P3_U3363 );
nand NAND2_9681 ( P3_U5828 , P3_U3897 , P3_U3054 );
nand NAND2_9682 ( P3_U5829 , P3_DATAO_REG_30_ , P3_U3363 );
nand NAND2_9683 ( P3_U5830 , P3_U3897 , P3_U3058 );
nand NAND2_9684 ( P3_U5831 , P3_DATAO_REG_31_ , P3_U3363 );
nand NAND2_9685 ( P3_U5832 , P3_U3897 , P3_U3055 );
nand NAND2_9686 ( P3_U5833 , P3_U3379 , P3_U3313 );
nand NAND2_9687 ( P3_U5834 , P3_U5450 , P3_U3911 );
not NOT1_9688 ( P3_U5835 , P3_U3760 );
nand NAND2_9689 ( P3_U5836 , P3_R1269_U11 , P3_U5835 );
nand NAND2_9690 ( P3_U5837 , P3_U3760 , P3_U3867 );
nand NAND2_9691 ( P3_U5838 , P3_U3900 , P3_U3052 );
nand NAND2_9692 ( P3_U5839 , P3_U3348 , P3_U4539 );
nand NAND2_9693 ( P3_U5840 , P3_U5839 , P3_U5838 );
nand NAND2_9694 ( P3_U5841 , P3_U3899 , P3_U3053 );
nand NAND2_9695 ( P3_U5842 , P3_U3350 , P3_U4557 );
nand NAND2_9696 ( P3_U5843 , P3_U5842 , P3_U5841 );
nand NAND2_9697 ( P3_U5844 , P3_U3872 , P3_U3055 );
nand NAND2_9698 ( P3_U5845 , P3_U3356 , P3_U4613 );
nand NAND2_9699 ( P3_U5846 , P3_U5845 , P3_U5844 );
nand NAND2_9700 ( P3_U5847 , P3_U3908 , P3_U3054 );
nand NAND2_9701 ( P3_U5848 , P3_U3353 , P3_U4575 );
nand NAND2_9702 ( P3_U5849 , P3_U5848 , P3_U5847 );
nand NAND2_9703 ( P3_U5850 , P3_U3906 , P3_U3074 );
nand NAND2_9704 ( P3_U5851 , P3_U3336 , P3_U4431 );
nand NAND2_9705 ( P3_U5852 , P3_U5851 , P3_U5850 );
nand NAND2_9706 ( P3_U5853 , P3_U3907 , P3_U3075 );
nand NAND2_9707 ( P3_U5854 , P3_U3334 , P3_U4413 );
nand NAND2_9708 ( P3_U5855 , P3_U5854 , P3_U5853 );
nand NAND2_9709 ( P3_U5856 , P3_U5503 , P3_U4107 );
nand NAND2_9710 ( P3_U5857 , P3_U3398 , P3_U3063 );
nand NAND2_9711 ( P3_U5858 , P3_U5857 , P3_U5856 );
nand NAND2_9712 ( P3_U5859 , P3_U5559 , P3_U4251 );
nand NAND2_9713 ( P3_U5860 , P3_U3422 , P3_U3062 );
nand NAND2_9714 ( P3_U5861 , P3_U5860 , P3_U5859 );
nand NAND2_9715 ( P3_U5862 , P3_U5552 , P3_U4233 );
nand NAND2_9716 ( P3_U5863 , P3_U3419 , P3_U3061 );
nand NAND2_9717 ( P3_U5864 , P3_U5863 , P3_U5862 );
nand NAND2_9718 ( P3_U5865 , P3_U5510 , P3_U4125 );
nand NAND2_9719 ( P3_U5866 , P3_U3401 , P3_U3059 );
nand NAND2_9720 ( P3_U5867 , P3_U5866 , P3_U5865 );
nand NAND2_9721 ( P3_U5868 , P3_U3905 , P3_U3060 );
nand NAND2_9722 ( P3_U5869 , P3_U3338 , P3_U4449 );
nand NAND2_9723 ( P3_U5870 , P3_U5869 , P3_U5868 );
nand NAND2_9724 ( P3_U5871 , P3_U5601 , P3_U4359 );
nand NAND2_9725 ( P3_U5872 , P3_U3440 , P3_U3068 );
nand NAND2_9726 ( P3_U5873 , P3_U5872 , P3_U5871 );
nand NAND2_9727 ( P3_U5874 , P3_U5594 , P3_U4341 );
nand NAND2_9728 ( P3_U5875 , P3_U3437 , P3_U3072 );
nand NAND2_9729 ( P3_U5876 , P3_U5875 , P3_U5874 );
nand NAND2_9730 ( P3_U5877 , P3_U5587 , P3_U4323 );
nand NAND2_9731 ( P3_U5878 , P3_U3434 , P3_U3073 );
nand NAND2_9732 ( P3_U5879 , P3_U5878 , P3_U5877 );
nand NAND2_9733 ( P3_U5880 , P3_U5566 , P3_U4269 );
nand NAND2_9734 ( P3_U5881 , P3_U3425 , P3_U3071 );
nand NAND2_9735 ( P3_U5882 , P3_U5881 , P3_U5880 );
nand NAND2_9736 ( P3_U5883 , P3_U5524 , P3_U4161 );
nand NAND2_9737 ( P3_U5884 , P3_U3407 , P3_U3070 );
nand NAND2_9738 ( P3_U5885 , P3_U5884 , P3_U5883 );
nand NAND2_9739 ( P3_U5886 , P3_U5531 , P3_U4179 );
nand NAND2_9740 ( P3_U5887 , P3_U3410 , P3_U3069 );
nand NAND2_9741 ( P3_U5888 , P3_U5887 , P3_U5886 );
nand NAND2_9742 ( P3_U5889 , P3_U5496 , P3_U4082 );
nand NAND2_9743 ( P3_U5890 , P3_U3395 , P3_U3067 );
nand NAND2_9744 ( P3_U5891 , P3_U5890 , P3_U5889 );
nand NAND2_9745 ( P3_U5892 , P3_U5517 , P3_U4143 );
nand NAND2_9746 ( P3_U5893 , P3_U3404 , P3_U3066 );
nand NAND2_9747 ( P3_U5894 , P3_U5893 , P3_U5892 );
nand NAND2_9748 ( P3_U5895 , P3_U5608 , P3_U4377 );
nand NAND2_9749 ( P3_U5896 , P3_U3443 , P3_U3081 );
nand NAND2_9750 ( P3_U5897 , P3_U5896 , P3_U5895 );
nand NAND2_9751 ( P3_U5898 , P3_U5573 , P3_U4287 );
nand NAND2_9752 ( P3_U5899 , P3_U3428 , P3_U3079 );
nand NAND2_9753 ( P3_U5900 , P3_U5899 , P3_U5898 );
nand NAND2_9754 ( P3_U5901 , P3_U5580 , P3_U4305 );
nand NAND2_9755 ( P3_U5902 , P3_U3431 , P3_U3078 );
nand NAND2_9756 ( P3_U5903 , P3_U5902 , P3_U5901 );
nand NAND2_9757 ( P3_U5904 , P3_U5489 , P3_U4063 );
nand NAND2_9758 ( P3_U5905 , P3_U3392 , P3_U3077 );
nand NAND2_9759 ( P3_U5906 , P3_U5905 , P3_U5904 );
nand NAND2_9760 ( P3_U5907 , P3_U5473 , P3_U4087 );
nand NAND2_9761 ( P3_U5908 , P3_U3387 , P3_U3076 );
nand NAND2_9762 ( P3_U5909 , P3_U5908 , P3_U5907 );
nand NAND2_9763 ( P3_U5910 , P3_U5538 , P3_U4197 );
nand NAND2_9764 ( P3_U5911 , P3_U3413 , P3_U3083 );
nand NAND2_9765 ( P3_U5912 , P3_U5911 , P3_U5910 );
nand NAND2_9766 ( P3_U5913 , P3_U5545 , P3_U4215 );
nand NAND2_9767 ( P3_U5914 , P3_U3416 , P3_U3082 );
nand NAND2_9768 ( P3_U5915 , P3_U5914 , P3_U5913 );
nand NAND2_9769 ( P3_U5916 , P3_U5613 , P3_U4395 );
nand NAND2_9770 ( P3_U5917 , P3_U3445 , P3_U3080 );
nand NAND2_9771 ( P3_U5918 , P3_U5917 , P3_U5916 );
nand NAND2_9772 ( P3_U5919 , P3_U3901 , P3_U3056 );
nand NAND2_9773 ( P3_U5920 , P3_U3346 , P3_U4521 );
nand NAND2_9774 ( P3_U5921 , P3_U5920 , P3_U5919 );
nand NAND2_9775 ( P3_U5922 , P3_U3902 , P3_U3057 );
nand NAND2_9776 ( P3_U5923 , P3_U3344 , P3_U4503 );
nand NAND2_9777 ( P3_U5924 , P3_U5923 , P3_U5922 );
nand NAND2_9778 ( P3_U5925 , P3_U3904 , P3_U3065 );
nand NAND2_9779 ( P3_U5926 , P3_U3340 , P3_U4467 );
nand NAND2_9780 ( P3_U5927 , P3_U5926 , P3_U5925 );
nand NAND2_9781 ( P3_U5928 , P3_U3903 , P3_U3064 );
nand NAND2_9782 ( P3_U5929 , P3_U3342 , P3_U4485 );
nand NAND2_9783 ( P3_U5930 , P3_U5929 , P3_U5928 );
nand NAND2_9784 ( P3_U5931 , P3_U3873 , P3_U3058 );
nand NAND2_9785 ( P3_U5932 , P3_U3355 , P3_U4593 );
nand NAND2_9786 ( P3_U5933 , P3_U5932 , P3_U5931 );
nand NAND2_9787 ( P3_U5934 , P3_U4978 , P3_U5450 );
nand NAND2_9788 ( P3_U5935 , P3_U3379 , P3_U3868 );
nand NAND2_9789 ( P3_U5936 , P3_U5935 , P3_U5934 );
nand NAND3_9790 ( P3_U5937 , P3_U5837 , P3_U5836 , P3_U5447 );
nand NAND3_9791 ( P3_U5938 , P3_U5456 , P3_U5936 , P3_U3378 );
nand NAND2_9792 ( P3_U5939 , P3_U3881 , P3_U3869 );
nand NAND2_9793 ( P3_U5940 , P3_R693_U14 , P3_U3891 );
nand NAND2_9794 ( P3_U5941 , P3_U5440 , P3_U3368 );
nand NAND2_9795 ( P3_U5942 , P3_U3380 , P3_U3375 );
nand NAND2_9796 ( P3_U5943 , P3_U5450 , P3_U5447 );
nand NAND3_9797 ( P3_U5944 , P3_U3388 , P3_U5456 , P3_U3378 );
nand NAND2_9798 ( P3_U5945 , P3_U3082 , P3_R1297_U6 );
nand NAND2_9799 ( P3_U5946 , P3_U3082 , P3_U3871 );
nand NAND2_9800 ( P3_U5947 , P3_U3083 , P3_R1297_U6 );
nand NAND2_9801 ( P3_U5948 , P3_U3083 , P3_U3871 );
nand NAND2_9802 ( P3_U5949 , P3_U3069 , P3_R1297_U6 );
nand NAND2_9803 ( P3_U5950 , P3_U3069 , P3_U3871 );
nand NAND2_9804 ( P3_U5951 , P3_U3070 , P3_R1297_U6 );
nand NAND2_9805 ( P3_U5952 , P3_U3070 , P3_U3871 );
nand NAND2_9806 ( P3_U5953 , P3_U3066 , P3_R1297_U6 );
nand NAND2_9807 ( P3_U5954 , P3_U3066 , P3_U3871 );
nand NAND2_9808 ( P3_U5955 , P3_U3059 , P3_R1297_U6 );
nand NAND2_9809 ( P3_U5956 , P3_U3059 , P3_U3871 );
nand NAND2_9810 ( P3_U5957 , P3_R1300_U8 , P3_R1297_U6 );
nand NAND2_9811 ( P3_U5958 , P3_U3055 , P3_U3871 );
nand NAND2_9812 ( P3_U5959 , P3_R1300_U6 , P3_R1297_U6 );
nand NAND2_9813 ( P3_U5960 , P3_U3058 , P3_U3871 );
nand NAND2_9814 ( P3_U5961 , P3_U3063 , P3_R1297_U6 );
nand NAND2_9815 ( P3_U5962 , P3_U3063 , P3_U3871 );
nand NAND2_9816 ( P3_U5963 , P3_U3054 , P3_R1297_U6 );
nand NAND2_9817 ( P3_U5964 , P3_U3054 , P3_U3871 );
nand NAND2_9818 ( P3_U5965 , P3_U3053 , P3_R1297_U6 );
nand NAND2_9819 ( P3_U5966 , P3_U3053 , P3_U3871 );
nand NAND2_9820 ( P3_U5967 , P3_U3052 , P3_R1297_U6 );
nand NAND2_9821 ( P3_U5968 , P3_U3052 , P3_U3871 );
nand NAND2_9822 ( P3_U5969 , P3_U3056 , P3_R1297_U6 );
nand NAND2_9823 ( P3_U5970 , P3_U3056 , P3_U3871 );
nand NAND2_9824 ( P3_U5971 , P3_U3057 , P3_R1297_U6 );
nand NAND2_9825 ( P3_U5972 , P3_U3057 , P3_U3871 );
nand NAND2_9826 ( P3_U5973 , P3_U3064 , P3_R1297_U6 );
nand NAND2_9827 ( P3_U5974 , P3_U3064 , P3_U3871 );
nand NAND2_9828 ( P3_U5975 , P3_U3065 , P3_R1297_U6 );
nand NAND2_9829 ( P3_U5976 , P3_U3065 , P3_U3871 );
nand NAND2_9830 ( P3_U5977 , P3_U3060 , P3_R1297_U6 );
nand NAND2_9831 ( P3_U5978 , P3_U3060 , P3_U3871 );
nand NAND2_9832 ( P3_U5979 , P3_U3074 , P3_R1297_U6 );
nand NAND2_9833 ( P3_U5980 , P3_U3074 , P3_U3871 );
nand NAND2_9834 ( P3_U5981 , P3_U3075 , P3_R1297_U6 );
nand NAND2_9835 ( P3_U5982 , P3_U3075 , P3_U3871 );
nand NAND2_9836 ( P3_U5983 , P3_U3067 , P3_R1297_U6 );
nand NAND2_9837 ( P3_U5984 , P3_U3067 , P3_U3871 );
nand NAND2_9838 ( P3_U5985 , P3_U3080 , P3_R1297_U6 );
nand NAND2_9839 ( P3_U5986 , P3_U3080 , P3_U3871 );
nand NAND2_9840 ( P3_U5987 , P3_U3081 , P3_R1297_U6 );
nand NAND2_9841 ( P3_U5988 , P3_U3081 , P3_U3871 );
nand NAND2_9842 ( P3_U5989 , P3_U3068 , P3_R1297_U6 );
nand NAND2_9843 ( P3_U5990 , P3_U3068 , P3_U3871 );
nand NAND2_9844 ( P3_U5991 , P3_U3072 , P3_R1297_U6 );
nand NAND2_9845 ( P3_U5992 , P3_U3072 , P3_U3871 );
nand NAND2_9846 ( P3_U5993 , P3_U3073 , P3_R1297_U6 );
nand NAND2_9847 ( P3_U5994 , P3_U3073 , P3_U3871 );
nand NAND2_9848 ( P3_U5995 , P3_U3078 , P3_R1297_U6 );
nand NAND2_9849 ( P3_U5996 , P3_U3078 , P3_U3871 );
nand NAND2_9850 ( P3_U5997 , P3_U3079 , P3_R1297_U6 );
nand NAND2_9851 ( P3_U5998 , P3_U3079 , P3_U3871 );
nand NAND2_9852 ( P3_U5999 , P3_U3071 , P3_R1297_U6 );
nand NAND2_9853 ( P3_U6000 , P3_U3071 , P3_U3871 );
nand NAND2_9854 ( P3_U6001 , P3_U3062 , P3_R1297_U6 );
nand NAND2_9855 ( P3_U6002 , P3_U3062 , P3_U3871 );
nand NAND2_9856 ( P3_U6003 , P3_U3061 , P3_R1297_U6 );
nand NAND2_9857 ( P3_U6004 , P3_U3061 , P3_U3871 );
nand NAND2_9858 ( P3_U6005 , P3_U3077 , P3_R1297_U6 );
nand NAND2_9859 ( P3_U6006 , P3_U3077 , P3_U3871 );
nand NAND2_9860 ( P3_U6007 , P3_U3076 , P3_R1297_U6 );
nand NAND2_9861 ( P3_U6008 , P3_U3076 , P3_U3871 );
nand NAND2_9862 ( P3_U6009 , P3_U5468 , P3_REG1_REG_9_ );
nand NAND2_9863 ( P3_U6010 , P3_U3384 , P3_REG2_REG_9_ );
nand NAND2_9864 ( P3_U6011 , P3_U5468 , P3_REG1_REG_8_ );
nand NAND2_9865 ( P3_U6012 , P3_U3384 , P3_REG2_REG_8_ );
nand NAND2_9866 ( P3_U6013 , P3_U5468 , P3_REG1_REG_7_ );
nand NAND2_9867 ( P3_U6014 , P3_U3384 , P3_REG2_REG_7_ );
nand NAND2_9868 ( P3_U6015 , P3_U5468 , P3_REG1_REG_6_ );
nand NAND2_9869 ( P3_U6016 , P3_U3384 , P3_REG2_REG_6_ );
nand NAND2_9870 ( P3_U6017 , P3_U5468 , P3_REG1_REG_5_ );
nand NAND2_9871 ( P3_U6018 , P3_U3384 , P3_REG2_REG_5_ );
nand NAND2_9872 ( P3_U6019 , P3_U5468 , P3_REG1_REG_4_ );
nand NAND2_9873 ( P3_U6020 , P3_U3384 , P3_REG2_REG_4_ );
nand NAND2_9874 ( P3_U6021 , P3_U5468 , P3_REG1_REG_3_ );
nand NAND2_9875 ( P3_U6022 , P3_U3384 , P3_REG2_REG_3_ );
nand NAND2_9876 ( P3_U6023 , P3_U5468 , P3_REG1_REG_2_ );
nand NAND2_9877 ( P3_U6024 , P3_U3384 , P3_REG2_REG_2_ );
nand NAND2_9878 ( P3_U6025 , P3_U5468 , P3_REG1_REG_19_ );
nand NAND2_9879 ( P3_U6026 , P3_U3384 , P3_REG2_REG_19_ );
nand NAND2_9880 ( P3_U6027 , P3_U5468 , P3_REG1_REG_18_ );
nand NAND2_9881 ( P3_U6028 , P3_U3384 , P3_REG2_REG_18_ );
nand NAND2_9882 ( P3_U6029 , P3_U5468 , P3_REG1_REG_17_ );
nand NAND2_9883 ( P3_U6030 , P3_U3384 , P3_REG2_REG_17_ );
nand NAND2_9884 ( P3_U6031 , P3_U5468 , P3_REG1_REG_16_ );
nand NAND2_9885 ( P3_U6032 , P3_U3384 , P3_REG2_REG_16_ );
nand NAND2_9886 ( P3_U6033 , P3_U5468 , P3_REG1_REG_15_ );
nand NAND2_9887 ( P3_U6034 , P3_U3384 , P3_REG2_REG_15_ );
nand NAND2_9888 ( P3_U6035 , P3_U5468 , P3_REG1_REG_14_ );
nand NAND2_9889 ( P3_U6036 , P3_U3384 , P3_REG2_REG_14_ );
nand NAND2_9890 ( P3_U6037 , P3_U5468 , P3_REG1_REG_13_ );
nand NAND2_9891 ( P3_U6038 , P3_U3384 , P3_REG2_REG_13_ );
nand NAND2_9892 ( P3_U6039 , P3_U5468 , P3_REG1_REG_12_ );
nand NAND2_9893 ( P3_U6040 , P3_U3384 , P3_REG2_REG_12_ );
nand NAND2_9894 ( P3_U6041 , P3_U5468 , P3_REG1_REG_11_ );
nand NAND2_9895 ( P3_U6042 , P3_U3384 , P3_REG2_REG_11_ );
nand NAND2_9896 ( P3_U6043 , P3_U5468 , P3_REG1_REG_10_ );
nand NAND2_9897 ( P3_U6044 , P3_U3384 , P3_REG2_REG_10_ );
nand NAND2_9898 ( P3_U6045 , P3_U5468 , P3_REG1_REG_1_ );
nand NAND2_9899 ( P3_U6046 , P3_U3384 , P3_REG2_REG_1_ );
nand NAND2_9900 ( P3_U6047 , P3_U5468 , P3_REG1_REG_0_ );
nand NAND2_9901 ( P3_U6048 , P3_U3384 , P3_REG2_REG_0_ );
nand NAND2_9902 ( P3_R1161_U448 , P3_R1161_U286 , P3_R1161_U446 );
nand NAND2_9903 ( P3_R1161_U447 , P3_R1161_U158 , P3_R1161_U159 );
nand NAND2_9904 ( P3_R1161_U446 , P3_R1161_U445 , P3_R1161_U444 );
nand NAND2_9905 ( P3_R1161_U445 , P3_U3905 , P3_R1161_U83 );
nand NAND2_9906 ( P3_R1161_U444 , P3_U3060 , P3_R1161_U82 );
nand NAND2_9907 ( P3_R1161_U443 , P3_U3905 , P3_R1161_U83 );
nand NAND2_9908 ( P3_R1161_U442 , P3_U3060 , P3_R1161_U82 );
nand NAND2_9909 ( P3_R1161_U441 , P3_R1161_U290 , P3_R1161_U439 );
nand NAND2_9910 ( P3_R1161_U440 , P3_R1161_U156 , P3_R1161_U157 );
nand NAND2_9911 ( P3_R1161_U439 , P3_R1161_U438 , P3_R1161_U437 );
nand NAND2_9912 ( P3_R1161_U438 , P3_U3904 , P3_R1161_U85 );
nand NAND2_9913 ( P3_R1161_U437 , P3_U3065 , P3_R1161_U84 );
nand NAND2_9914 ( P3_R1161_U436 , P3_U3904 , P3_R1161_U85 );
nand NAND2_9915 ( P3_R1161_U435 , P3_U3065 , P3_R1161_U84 );
nand NAND2_9916 ( P3_R1161_U434 , P3_R1161_U294 , P3_R1161_U432 );
nand NAND2_9917 ( P3_R1161_U433 , P3_R1161_U358 , P3_R1161_U155 );
nand NAND2_9918 ( P3_R1161_U432 , P3_R1161_U431 , P3_R1161_U430 );
nand NAND2_9919 ( P3_R1161_U431 , P3_U3903 , P3_R1161_U53 );
nand NAND2_9920 ( P3_R1161_U430 , P3_U3064 , P3_R1161_U52 );
and AND2_9921 ( SUB_1605_U6 , SUB_1605_U194 , SUB_1605_U190 );
and AND2_9922 ( SUB_1605_U7 , SUB_1605_U202 , SUB_1605_U200 );
and AND2_9923 ( SUB_1605_U8 , SUB_1605_U7 , SUB_1605_U204 );
and AND2_9924 ( SUB_1605_U9 , SUB_1605_U212 , SUB_1605_U208 );
and AND2_9925 ( SUB_1605_U10 , SUB_1605_U9 , SUB_1605_U215 );
and AND2_9926 ( SUB_1605_U11 , SUB_1605_U363 , SUB_1605_U362 );
nand NAND2_9927 ( SUB_1605_U12 , SUB_1605_U128 , SUB_1605_U323 );
nand NAND2_9928 ( SUB_1605_U13 , SUB_1605_U175 , SUB_1605_U291 );
not NOT1_9929 ( SUB_1605_U14 , P1_DATAO_REG_8_ );
not NOT1_9930 ( SUB_1605_U15 , P2_DATAO_REG_8_ );
not NOT1_9931 ( SUB_1605_U16 , P2_DATAO_REG_7_ );
not NOT1_9932 ( SUB_1605_U17 , P1_DATAO_REG_6_ );
not NOT1_9933 ( SUB_1605_U18 , P1_DATAO_REG_7_ );
not NOT1_9934 ( SUB_1605_U19 , P2_DATAO_REG_6_ );
not NOT1_9935 ( SUB_1605_U20 , P1_DATAO_REG_5_ );
nand NAND2_9936 ( SUB_1605_U21 , SUB_1605_U303 , SUB_1605_U204 );
not NOT1_9937 ( SUB_1605_U22 , P1_DATAO_REG_4_ );
not NOT1_9938 ( SUB_1605_U23 , P2_DATAO_REG_0_ );
not NOT1_9939 ( SUB_1605_U24 , P1_DATAO_REG_1_ );
not NOT1_9940 ( SUB_1605_U25 , P2_DATAO_REG_4_ );
not NOT1_9941 ( SUB_1605_U26 , P2_DATAO_REG_2_ );
not NOT1_9942 ( SUB_1605_U27 , P2_DATAO_REG_3_ );
not NOT1_9943 ( SUB_1605_U28 , P1_DATAO_REG_2_ );
not NOT1_9944 ( SUB_1605_U29 , P1_DATAO_REG_3_ );
not NOT1_9945 ( SUB_1605_U30 , P2_DATAO_REG_5_ );
not NOT1_9946 ( SUB_1605_U31 , P2_DATAO_REG_9_ );
not NOT1_9947 ( SUB_1605_U32 , P1_DATAO_REG_9_ );
not NOT1_9948 ( SUB_1605_U33 , P1_DATAO_REG_12_ );
not NOT1_9949 ( SUB_1605_U34 , P2_DATAO_REG_12_ );
not NOT1_9950 ( SUB_1605_U35 , P2_DATAO_REG_11_ );
not NOT1_9951 ( SUB_1605_U36 , P2_DATAO_REG_10_ );
not NOT1_9952 ( SUB_1605_U37 , P1_DATAO_REG_11_ );
not NOT1_9953 ( SUB_1605_U38 , P1_DATAO_REG_10_ );
nand NAND2_9954 ( SUB_1605_U39 , P1_DATAO_REG_9_ , SUB_1605_U31 );
not NOT1_9955 ( SUB_1605_U40 , P2_DATAO_REG_13_ );
not NOT1_9956 ( SUB_1605_U41 , P1_DATAO_REG_13_ );
not NOT1_9957 ( SUB_1605_U42 , P2_DATAO_REG_14_ );
not NOT1_9958 ( SUB_1605_U43 , P1_DATAO_REG_14_ );
not NOT1_9959 ( SUB_1605_U44 , P2_DATAO_REG_15_ );
not NOT1_9960 ( SUB_1605_U45 , P1_DATAO_REG_15_ );
not NOT1_9961 ( SUB_1605_U46 , P2_DATAO_REG_16_ );
not NOT1_9962 ( SUB_1605_U47 , P1_DATAO_REG_16_ );
not NOT1_9963 ( SUB_1605_U48 , P2_DATAO_REG_17_ );
not NOT1_9964 ( SUB_1605_U49 , P1_DATAO_REG_17_ );
not NOT1_9965 ( SUB_1605_U50 , P2_DATAO_REG_18_ );
not NOT1_9966 ( SUB_1605_U51 , P1_DATAO_REG_18_ );
not NOT1_9967 ( SUB_1605_U52 , P2_DATAO_REG_19_ );
not NOT1_9968 ( SUB_1605_U53 , P1_DATAO_REG_19_ );
not NOT1_9969 ( SUB_1605_U54 , P2_DATAO_REG_20_ );
not NOT1_9970 ( SUB_1605_U55 , P1_DATAO_REG_20_ );
not NOT1_9971 ( SUB_1605_U56 , P2_DATAO_REG_21_ );
not NOT1_9972 ( SUB_1605_U57 , P1_DATAO_REG_21_ );
not NOT1_9973 ( SUB_1605_U58 , P2_DATAO_REG_22_ );
not NOT1_9974 ( SUB_1605_U59 , P1_DATAO_REG_22_ );
not NOT1_9975 ( SUB_1605_U60 , P2_DATAO_REG_23_ );
not NOT1_9976 ( SUB_1605_U61 , P1_DATAO_REG_23_ );
not NOT1_9977 ( SUB_1605_U62 , P2_DATAO_REG_24_ );
not NOT1_9978 ( SUB_1605_U63 , P1_DATAO_REG_24_ );
not NOT1_9979 ( SUB_1605_U64 , P2_DATAO_REG_25_ );
not NOT1_9980 ( SUB_1605_U65 , P1_DATAO_REG_25_ );
not NOT1_9981 ( SUB_1605_U66 , P2_DATAO_REG_26_ );
not NOT1_9982 ( SUB_1605_U67 , P1_DATAO_REG_26_ );
not NOT1_9983 ( SUB_1605_U68 , P2_DATAO_REG_27_ );
not NOT1_9984 ( SUB_1605_U69 , P1_DATAO_REG_27_ );
not NOT1_9985 ( SUB_1605_U70 , P2_DATAO_REG_28_ );
not NOT1_9986 ( SUB_1605_U71 , P1_DATAO_REG_28_ );
not NOT1_9987 ( SUB_1605_U72 , P2_DATAO_REG_29_ );
not NOT1_9988 ( SUB_1605_U73 , P1_DATAO_REG_29_ );
not NOT1_9989 ( SUB_1605_U74 , P1_DATAO_REG_30_ );
not NOT1_9990 ( SUB_1605_U75 , P2_DATAO_REG_30_ );
nand NAND2_9991 ( SUB_1605_U76 , SUB_1605_U308 , SUB_1605_U216 );
nand NAND2_9992 ( SUB_1605_U77 , SUB_1605_U305 , SUB_1605_U213 );
not NOT1_9993 ( SUB_1605_U78 , P1_DATAO_REG_0_ );
nand NAND2_9994 ( SUB_1605_U79 , SUB_1605_U328 , SUB_1605_U327 );
nand NAND2_9995 ( SUB_1605_U80 , SUB_1605_U333 , SUB_1605_U332 );
nand NAND2_9996 ( SUB_1605_U81 , SUB_1605_U338 , SUB_1605_U337 );
nand NAND2_9997 ( SUB_1605_U82 , SUB_1605_U343 , SUB_1605_U342 );
nand NAND2_9998 ( SUB_1605_U83 , SUB_1605_U348 , SUB_1605_U347 );
nand NAND2_9999 ( SUB_1605_U84 , SUB_1605_U353 , SUB_1605_U352 );
nand NAND2_10000 ( SUB_1605_U85 , SUB_1605_U358 , SUB_1605_U357 );
nand NAND2_10001 ( SUB_1605_U86 , SUB_1605_U370 , SUB_1605_U369 );
nand NAND2_10002 ( SUB_1605_U87 , SUB_1605_U375 , SUB_1605_U374 );
nand NAND2_10003 ( SUB_1605_U88 , SUB_1605_U380 , SUB_1605_U379 );
nand NAND2_10004 ( SUB_1605_U89 , SUB_1605_U385 , SUB_1605_U384 );
nand NAND2_10005 ( SUB_1605_U90 , SUB_1605_U390 , SUB_1605_U389 );
nand NAND2_10006 ( SUB_1605_U91 , SUB_1605_U395 , SUB_1605_U394 );
nand NAND2_10007 ( SUB_1605_U92 , SUB_1605_U400 , SUB_1605_U399 );
nand NAND2_10008 ( SUB_1605_U93 , SUB_1605_U405 , SUB_1605_U404 );
nand NAND2_10009 ( SUB_1605_U94 , SUB_1605_U410 , SUB_1605_U409 );
nand NAND2_10010 ( SUB_1605_U95 , SUB_1605_U415 , SUB_1605_U414 );
nand NAND2_10011 ( SUB_1605_U96 , SUB_1605_U420 , SUB_1605_U419 );
nand NAND2_10012 ( SUB_1605_U97 , SUB_1605_U425 , SUB_1605_U424 );
nand NAND2_10013 ( SUB_1605_U98 , SUB_1605_U430 , SUB_1605_U429 );
nand NAND2_10014 ( SUB_1605_U99 , SUB_1605_U435 , SUB_1605_U434 );
nand NAND2_10015 ( SUB_1605_U100 , SUB_1605_U440 , SUB_1605_U439 );
nand NAND2_10016 ( SUB_1605_U101 , SUB_1605_U445 , SUB_1605_U444 );
nand NAND2_10017 ( SUB_1605_U102 , SUB_1605_U450 , SUB_1605_U449 );
nand NAND2_10018 ( SUB_1605_U103 , SUB_1605_U455 , SUB_1605_U454 );
nand NAND2_10019 ( SUB_1605_U104 , SUB_1605_U460 , SUB_1605_U459 );
nand NAND2_10020 ( SUB_1605_U105 , SUB_1605_U465 , SUB_1605_U464 );
nand NAND2_10021 ( SUB_1605_U106 , SUB_1605_U470 , SUB_1605_U469 );
nand NAND2_10022 ( SUB_1605_U107 , SUB_1605_U475 , SUB_1605_U474 );
nand NAND2_10023 ( SUB_1605_U108 , SUB_1605_U480 , SUB_1605_U479 );
and AND2_10024 ( SUB_1605_U109 , P1_DATAO_REG_5_ , SUB_1605_U30 );
and AND2_10025 ( SUB_1605_U110 , SUB_1605_U205 , SUB_1605_U203 );
and AND2_10026 ( SUB_1605_U111 , SUB_1605_U197 , SUB_1605_U6 );
and AND2_10027 ( SUB_1605_U112 , SUB_1605_U299 , SUB_1605_U197 );
and AND2_10028 ( SUB_1605_U113 , SUB_1605_U298 , SUB_1605_U198 );
and AND2_10029 ( SUB_1605_U114 , SUB_1605_U206 , SUB_1605_U8 );
and AND2_10030 ( SUB_1605_U115 , SUB_1605_U302 , SUB_1605_U207 );
nand NAND2_10031 ( SUB_1605_U116 , SUB_1605_U325 , SUB_1605_U324 );
nand NAND2_10032 ( SUB_1605_U117 , SUB_1605_U330 , SUB_1605_U329 );
and AND2_10033 ( SUB_1605_U118 , SUB_1605_U300 , SUB_1605_U203 );
nand NAND2_10034 ( SUB_1605_U119 , SUB_1605_U335 , SUB_1605_U334 );
nand NAND2_10035 ( SUB_1605_U120 , SUB_1605_U340 , SUB_1605_U339 );
nand NAND2_10036 ( SUB_1605_U121 , SUB_1605_U345 , SUB_1605_U344 );
nand NAND2_10037 ( SUB_1605_U122 , SUB_1605_U350 , SUB_1605_U349 );
nand NAND2_10038 ( SUB_1605_U123 , SUB_1605_U355 , SUB_1605_U354 );
and AND2_10039 ( SUB_1605_U124 , SUB_1605_U10 , SUB_1605_U218 );
and AND2_10040 ( SUB_1605_U125 , SUB_1605_U311 , SUB_1605_U219 );
and AND3_10041 ( SUB_1605_U126 , SUB_1605_U11 , SUB_1605_U290 , SUB_1605_U287 );
and AND2_10042 ( SUB_1605_U127 , SUB_1605_U289 , SUB_1605_U361 );
and AND2_10043 ( SUB_1605_U128 , SUB_1605_U161 , SUB_1605_U293 );
nand NAND2_10044 ( SUB_1605_U129 , SUB_1605_U367 , SUB_1605_U366 );
nand NAND2_10045 ( SUB_1605_U130 , SUB_1605_U372 , SUB_1605_U371 );
nand NAND2_10046 ( SUB_1605_U131 , SUB_1605_U377 , SUB_1605_U376 );
nand NAND2_10047 ( SUB_1605_U132 , SUB_1605_U382 , SUB_1605_U381 );
nand NAND2_10048 ( SUB_1605_U133 , SUB_1605_U387 , SUB_1605_U386 );
nand NAND2_10049 ( SUB_1605_U134 , SUB_1605_U392 , SUB_1605_U391 );
nand NAND2_10050 ( SUB_1605_U135 , SUB_1605_U397 , SUB_1605_U396 );
nand NAND2_10051 ( SUB_1605_U136 , SUB_1605_U402 , SUB_1605_U401 );
nand NAND2_10052 ( SUB_1605_U137 , SUB_1605_U407 , SUB_1605_U406 );
nand NAND2_10053 ( SUB_1605_U138 , SUB_1605_U412 , SUB_1605_U411 );
nand NAND2_10054 ( SUB_1605_U139 , SUB_1605_U417 , SUB_1605_U416 );
nand NAND2_10055 ( SUB_1605_U140 , SUB_1605_U422 , SUB_1605_U421 );
nand NAND2_10056 ( SUB_1605_U141 , SUB_1605_U427 , SUB_1605_U426 );
nand NAND2_10057 ( SUB_1605_U142 , SUB_1605_U432 , SUB_1605_U431 );
nand NAND2_10058 ( SUB_1605_U143 , SUB_1605_U437 , SUB_1605_U436 );
nand NAND2_10059 ( SUB_1605_U144 , SUB_1605_U442 , SUB_1605_U441 );
nand NAND2_10060 ( SUB_1605_U145 , SUB_1605_U447 , SUB_1605_U446 );
nand NAND2_10061 ( SUB_1605_U146 , SUB_1605_U452 , SUB_1605_U451 );
nand NAND2_10062 ( SUB_1605_U147 , SUB_1605_U457 , SUB_1605_U456 );
nand NAND2_10063 ( SUB_1605_U148 , SUB_1605_U462 , SUB_1605_U461 );
nand NAND2_10064 ( SUB_1605_U149 , SUB_1605_U467 , SUB_1605_U466 );
nand NAND2_10065 ( SUB_1605_U150 , SUB_1605_U472 , SUB_1605_U471 );
nand NAND2_10066 ( SUB_1605_U151 , SUB_1605_U477 , SUB_1605_U476 );
nand NAND2_10067 ( SUB_1605_U152 , SUB_1605_U115 , SUB_1605_U321 );
nand NAND2_10068 ( SUB_1605_U153 , SUB_1605_U319 , SUB_1605_U21 );
nand NAND2_10069 ( SUB_1605_U154 , SUB_1605_U118 , SUB_1605_U317 );
nand NAND2_10070 ( SUB_1605_U155 , SUB_1605_U315 , SUB_1605_U201 );
nand NAND2_10071 ( SUB_1605_U156 , SUB_1605_U113 , SUB_1605_U297 );
nand NAND2_10072 ( SUB_1605_U157 , SUB_1605_U296 , SUB_1605_U294 );
nand NAND2_10073 ( SUB_1605_U158 , SUB_1605_U192 , SUB_1605_U191 );
not NOT1_10074 ( SUB_1605_U159 , P2_DATAO_REG_31_ );
not NOT1_10075 ( SUB_1605_U160 , P1_DATAO_REG_31_ );
and AND2_10076 ( SUB_1605_U161 , SUB_1605_U365 , SUB_1605_U364 );
nand NAND2_10077 ( SUB_1605_U162 , SUB_1605_U287 , SUB_1605_U286 );
nand NAND3_10078 ( SUB_1605_U163 , SUB_1605_U188 , SUB_1605_U186 , SUB_1605_U292 );
nand NAND2_10079 ( SUB_1605_U164 , SUB_1605_U283 , SUB_1605_U282 );
nand NAND2_10080 ( SUB_1605_U165 , SUB_1605_U279 , SUB_1605_U278 );
nand NAND2_10081 ( SUB_1605_U166 , SUB_1605_U275 , SUB_1605_U274 );
nand NAND2_10082 ( SUB_1605_U167 , SUB_1605_U271 , SUB_1605_U270 );
nand NAND2_10083 ( SUB_1605_U168 , SUB_1605_U267 , SUB_1605_U266 );
nand NAND2_10084 ( SUB_1605_U169 , SUB_1605_U263 , SUB_1605_U262 );
nand NAND2_10085 ( SUB_1605_U170 , SUB_1605_U259 , SUB_1605_U258 );
nand NAND2_10086 ( SUB_1605_U171 , SUB_1605_U255 , SUB_1605_U254 );
nand NAND2_10087 ( SUB_1605_U172 , SUB_1605_U251 , SUB_1605_U250 );
nand NAND2_10088 ( SUB_1605_U173 , SUB_1605_U247 , SUB_1605_U246 );
not NOT1_10089 ( SUB_1605_U174 , P2_DATAO_REG_1_ );
nand NAND2_10090 ( SUB_1605_U175 , P2_DATAO_REG_0_ , SUB_1605_U78 );
nand NAND2_10091 ( SUB_1605_U176 , SUB_1605_U243 , SUB_1605_U242 );
nand NAND2_10092 ( SUB_1605_U177 , SUB_1605_U239 , SUB_1605_U238 );
nand NAND2_10093 ( SUB_1605_U178 , SUB_1605_U235 , SUB_1605_U234 );
nand NAND2_10094 ( SUB_1605_U179 , SUB_1605_U231 , SUB_1605_U230 );
nand NAND2_10095 ( SUB_1605_U180 , SUB_1605_U227 , SUB_1605_U226 );
nand NAND2_10096 ( SUB_1605_U181 , SUB_1605_U223 , SUB_1605_U222 );
nand NAND2_10097 ( SUB_1605_U182 , SUB_1605_U125 , SUB_1605_U310 );
nand NAND2_10098 ( SUB_1605_U183 , SUB_1605_U309 , SUB_1605_U307 );
nand NAND2_10099 ( SUB_1605_U184 , SUB_1605_U306 , SUB_1605_U304 );
nand NAND2_10100 ( SUB_1605_U185 , SUB_1605_U39 , SUB_1605_U209 );
nand NAND2_10101 ( SUB_1605_U186 , SUB_1605_U175 , SUB_1605_U174 );
not NOT1_10102 ( SUB_1605_U187 , SUB_1605_U175 );
nand NAND2_10103 ( SUB_1605_U188 , P1_DATAO_REG_1_ , SUB_1605_U175 );
not NOT1_10104 ( SUB_1605_U189 , SUB_1605_U163 );
nand NAND2_10105 ( SUB_1605_U190 , P2_DATAO_REG_2_ , SUB_1605_U28 );
nand NAND2_10106 ( SUB_1605_U191 , SUB_1605_U190 , SUB_1605_U312 );
nand NAND2_10107 ( SUB_1605_U192 , P1_DATAO_REG_2_ , SUB_1605_U26 );
not NOT1_10108 ( SUB_1605_U193 , SUB_1605_U158 );
nand NAND2_10109 ( SUB_1605_U194 , P2_DATAO_REG_3_ , SUB_1605_U29 );
nand NAND2_10110 ( SUB_1605_U195 , P1_DATAO_REG_3_ , SUB_1605_U27 );
not NOT1_10111 ( SUB_1605_U196 , SUB_1605_U157 );
nand NAND2_10112 ( SUB_1605_U197 , P2_DATAO_REG_4_ , SUB_1605_U22 );
nand NAND2_10113 ( SUB_1605_U198 , P1_DATAO_REG_4_ , SUB_1605_U25 );
not NOT1_10114 ( SUB_1605_U199 , SUB_1605_U156 );
nand NAND2_10115 ( SUB_1605_U200 , P2_DATAO_REG_5_ , SUB_1605_U20 );
nand NAND2_10116 ( SUB_1605_U201 , P1_DATAO_REG_5_ , SUB_1605_U30 );
nand NAND2_10117 ( SUB_1605_U202 , P2_DATAO_REG_6_ , SUB_1605_U17 );
nand NAND2_10118 ( SUB_1605_U203 , P1_DATAO_REG_6_ , SUB_1605_U19 );
nand NAND2_10119 ( SUB_1605_U204 , P2_DATAO_REG_7_ , SUB_1605_U18 );
nand NAND2_10120 ( SUB_1605_U205 , P1_DATAO_REG_7_ , SUB_1605_U16 );
nand NAND2_10121 ( SUB_1605_U206 , P2_DATAO_REG_8_ , SUB_1605_U14 );
nand NAND2_10122 ( SUB_1605_U207 , P1_DATAO_REG_8_ , SUB_1605_U15 );
nand NAND2_10123 ( SUB_1605_U208 , P2_DATAO_REG_9_ , SUB_1605_U32 );
nand NAND2_10124 ( SUB_1605_U209 , SUB_1605_U208 , SUB_1605_U152 );
not NOT1_10125 ( SUB_1605_U210 , SUB_1605_U39 );
not NOT1_10126 ( SUB_1605_U211 , SUB_1605_U185 );
nand NAND2_10127 ( SUB_1605_U212 , P2_DATAO_REG_10_ , SUB_1605_U38 );
nand NAND2_10128 ( SUB_1605_U213 , P1_DATAO_REG_10_ , SUB_1605_U36 );
not NOT1_10129 ( SUB_1605_U214 , SUB_1605_U184 );
nand NAND2_10130 ( SUB_1605_U215 , P2_DATAO_REG_11_ , SUB_1605_U37 );
nand NAND2_10131 ( SUB_1605_U216 , P1_DATAO_REG_11_ , SUB_1605_U35 );
not NOT1_10132 ( SUB_1605_U217 , SUB_1605_U183 );
nand NAND2_10133 ( SUB_1605_U218 , P2_DATAO_REG_12_ , SUB_1605_U33 );
nand NAND2_10134 ( SUB_1605_U219 , P1_DATAO_REG_12_ , SUB_1605_U34 );
not NOT1_10135 ( SUB_1605_U220 , SUB_1605_U182 );
nand NAND2_10136 ( SUB_1605_U221 , P2_DATAO_REG_13_ , SUB_1605_U41 );
nand NAND2_10137 ( SUB_1605_U222 , SUB_1605_U221 , SUB_1605_U182 );
nand NAND2_10138 ( SUB_1605_U223 , P1_DATAO_REG_13_ , SUB_1605_U40 );
not NOT1_10139 ( SUB_1605_U224 , SUB_1605_U181 );
nand NAND2_10140 ( SUB_1605_U225 , P2_DATAO_REG_14_ , SUB_1605_U43 );
nand NAND2_10141 ( SUB_1605_U226 , SUB_1605_U225 , SUB_1605_U181 );
nand NAND2_10142 ( SUB_1605_U227 , P1_DATAO_REG_14_ , SUB_1605_U42 );
not NOT1_10143 ( SUB_1605_U228 , SUB_1605_U180 );
nand NAND2_10144 ( SUB_1605_U229 , P2_DATAO_REG_15_ , SUB_1605_U45 );
nand NAND2_10145 ( SUB_1605_U230 , SUB_1605_U229 , SUB_1605_U180 );
nand NAND2_10146 ( SUB_1605_U231 , P1_DATAO_REG_15_ , SUB_1605_U44 );
not NOT1_10147 ( SUB_1605_U232 , SUB_1605_U179 );
nand NAND2_10148 ( SUB_1605_U233 , P2_DATAO_REG_16_ , SUB_1605_U47 );
nand NAND2_10149 ( SUB_1605_U234 , SUB_1605_U233 , SUB_1605_U179 );
nand NAND2_10150 ( SUB_1605_U235 , P1_DATAO_REG_16_ , SUB_1605_U46 );
not NOT1_10151 ( SUB_1605_U236 , SUB_1605_U178 );
nand NAND2_10152 ( SUB_1605_U237 , P2_DATAO_REG_17_ , SUB_1605_U49 );
nand NAND2_10153 ( SUB_1605_U238 , SUB_1605_U237 , SUB_1605_U178 );
nand NAND2_10154 ( SUB_1605_U239 , P1_DATAO_REG_17_ , SUB_1605_U48 );
not NOT1_10155 ( SUB_1605_U240 , SUB_1605_U177 );
nand NAND2_10156 ( SUB_1605_U241 , P2_DATAO_REG_18_ , SUB_1605_U51 );
nand NAND2_10157 ( SUB_1605_U242 , SUB_1605_U241 , SUB_1605_U177 );
nand NAND2_10158 ( SUB_1605_U243 , P1_DATAO_REG_18_ , SUB_1605_U50 );
not NOT1_10159 ( SUB_1605_U244 , SUB_1605_U176 );
nand NAND2_10160 ( SUB_1605_U245 , P2_DATAO_REG_19_ , SUB_1605_U53 );
nand NAND2_10161 ( SUB_1605_U246 , SUB_1605_U245 , SUB_1605_U176 );
nand NAND2_10162 ( SUB_1605_U247 , P1_DATAO_REG_19_ , SUB_1605_U52 );
not NOT1_10163 ( SUB_1605_U248 , SUB_1605_U173 );
nand NAND2_10164 ( SUB_1605_U249 , P2_DATAO_REG_20_ , SUB_1605_U55 );
nand NAND2_10165 ( SUB_1605_U250 , SUB_1605_U249 , SUB_1605_U173 );
nand NAND2_10166 ( SUB_1605_U251 , P1_DATAO_REG_20_ , SUB_1605_U54 );
not NOT1_10167 ( SUB_1605_U252 , SUB_1605_U172 );
nand NAND2_10168 ( SUB_1605_U253 , P2_DATAO_REG_21_ , SUB_1605_U57 );
nand NAND2_10169 ( SUB_1605_U254 , SUB_1605_U253 , SUB_1605_U172 );
nand NAND2_10170 ( SUB_1605_U255 , P1_DATAO_REG_21_ , SUB_1605_U56 );
not NOT1_10171 ( SUB_1605_U256 , SUB_1605_U171 );
nand NAND2_10172 ( SUB_1605_U257 , P2_DATAO_REG_22_ , SUB_1605_U59 );
nand NAND2_10173 ( SUB_1605_U258 , SUB_1605_U257 , SUB_1605_U171 );
nand NAND2_10174 ( SUB_1605_U259 , P1_DATAO_REG_22_ , SUB_1605_U58 );
not NOT1_10175 ( SUB_1605_U260 , SUB_1605_U170 );
nand NAND2_10176 ( SUB_1605_U261 , P2_DATAO_REG_23_ , SUB_1605_U61 );
nand NAND2_10177 ( SUB_1605_U262 , SUB_1605_U261 , SUB_1605_U170 );
nand NAND2_10178 ( SUB_1605_U263 , P1_DATAO_REG_23_ , SUB_1605_U60 );
not NOT1_10179 ( SUB_1605_U264 , SUB_1605_U169 );
nand NAND2_10180 ( SUB_1605_U265 , P2_DATAO_REG_24_ , SUB_1605_U63 );
nand NAND2_10181 ( SUB_1605_U266 , SUB_1605_U265 , SUB_1605_U169 );
nand NAND2_10182 ( SUB_1605_U267 , P1_DATAO_REG_24_ , SUB_1605_U62 );
not NOT1_10183 ( SUB_1605_U268 , SUB_1605_U168 );
nand NAND2_10184 ( SUB_1605_U269 , P2_DATAO_REG_25_ , SUB_1605_U65 );
nand NAND2_10185 ( SUB_1605_U270 , SUB_1605_U269 , SUB_1605_U168 );
nand NAND2_10186 ( SUB_1605_U271 , P1_DATAO_REG_25_ , SUB_1605_U64 );
not NOT1_10187 ( SUB_1605_U272 , SUB_1605_U167 );
nand NAND2_10188 ( SUB_1605_U273 , P2_DATAO_REG_26_ , SUB_1605_U67 );
nand NAND2_10189 ( SUB_1605_U274 , SUB_1605_U273 , SUB_1605_U167 );
nand NAND2_10190 ( SUB_1605_U275 , P1_DATAO_REG_26_ , SUB_1605_U66 );
not NOT1_10191 ( SUB_1605_U276 , SUB_1605_U166 );
nand NAND2_10192 ( SUB_1605_U277 , P2_DATAO_REG_27_ , SUB_1605_U69 );
nand NAND2_10193 ( SUB_1605_U278 , SUB_1605_U277 , SUB_1605_U166 );
nand NAND2_10194 ( SUB_1605_U279 , P1_DATAO_REG_27_ , SUB_1605_U68 );
not NOT1_10195 ( SUB_1605_U280 , SUB_1605_U165 );
nand NAND2_10196 ( SUB_1605_U281 , P2_DATAO_REG_28_ , SUB_1605_U71 );
nand NAND2_10197 ( SUB_1605_U282 , SUB_1605_U281 , SUB_1605_U165 );
nand NAND2_10198 ( SUB_1605_U283 , P1_DATAO_REG_28_ , SUB_1605_U70 );
not NOT1_10199 ( SUB_1605_U284 , SUB_1605_U164 );
nand NAND2_10200 ( SUB_1605_U285 , P2_DATAO_REG_29_ , SUB_1605_U73 );
nand NAND2_10201 ( SUB_1605_U286 , SUB_1605_U285 , SUB_1605_U164 );
nand NAND2_10202 ( SUB_1605_U287 , P1_DATAO_REG_29_ , SUB_1605_U72 );
not NOT1_10203 ( SUB_1605_U288 , SUB_1605_U162 );
nand NAND2_10204 ( SUB_1605_U289 , P2_DATAO_REG_30_ , SUB_1605_U74 );
nand NAND2_10205 ( SUB_1605_U290 , P1_DATAO_REG_30_ , SUB_1605_U75 );
nand NAND2_10206 ( SUB_1605_U291 , P1_DATAO_REG_0_ , SUB_1605_U23 );
nand NAND2_10207 ( SUB_1605_U292 , P1_DATAO_REG_1_ , SUB_1605_U174 );
nand NAND2_10208 ( SUB_1605_U293 , SUB_1605_U286 , SUB_1605_U126 );
nand NAND2_10209 ( SUB_1605_U294 , SUB_1605_U6 , SUB_1605_U163 );
nand NAND2_10210 ( SUB_1605_U295 , SUB_1605_U195 , SUB_1605_U192 );
nand NAND2_10211 ( SUB_1605_U296 , SUB_1605_U295 , SUB_1605_U299 );
nand NAND2_10212 ( SUB_1605_U297 , SUB_1605_U111 , SUB_1605_U163 );
nand NAND2_10213 ( SUB_1605_U298 , SUB_1605_U112 , SUB_1605_U295 );
nand NAND2_10214 ( SUB_1605_U299 , P2_DATAO_REG_3_ , SUB_1605_U29 );
nand NAND2_10215 ( SUB_1605_U300 , SUB_1605_U109 , SUB_1605_U202 );
not NOT1_10216 ( SUB_1605_U301 , SUB_1605_U21 );
nand NAND2_10217 ( SUB_1605_U302 , SUB_1605_U301 , SUB_1605_U206 );
nand NAND2_10218 ( SUB_1605_U303 , SUB_1605_U110 , SUB_1605_U300 );
nand NAND2_10219 ( SUB_1605_U304 , SUB_1605_U9 , SUB_1605_U152 );
nand NAND2_10220 ( SUB_1605_U305 , SUB_1605_U210 , SUB_1605_U212 );
not NOT1_10221 ( SUB_1605_U306 , SUB_1605_U77 );
nand NAND2_10222 ( SUB_1605_U307 , SUB_1605_U10 , SUB_1605_U152 );
nand NAND2_10223 ( SUB_1605_U308 , SUB_1605_U77 , SUB_1605_U215 );
not NOT1_10224 ( SUB_1605_U309 , SUB_1605_U76 );
nand NAND2_10225 ( SUB_1605_U310 , SUB_1605_U124 , SUB_1605_U152 );
nand NAND2_10226 ( SUB_1605_U311 , SUB_1605_U76 , SUB_1605_U218 );
nand NAND3_10227 ( SUB_1605_U312 , SUB_1605_U313 , SUB_1605_U292 , SUB_1605_U314 );
nand NAND2_10228 ( SUB_1605_U313 , P1_DATAO_REG_1_ , SUB_1605_U175 );
nand NAND2_10229 ( SUB_1605_U314 , SUB_1605_U175 , SUB_1605_U174 );
nand NAND2_10230 ( SUB_1605_U315 , SUB_1605_U200 , SUB_1605_U156 );
not NOT1_10231 ( SUB_1605_U316 , SUB_1605_U155 );
nand NAND2_10232 ( SUB_1605_U317 , SUB_1605_U7 , SUB_1605_U156 );
not NOT1_10233 ( SUB_1605_U318 , SUB_1605_U154 );
nand NAND2_10234 ( SUB_1605_U319 , SUB_1605_U8 , SUB_1605_U156 );
not NOT1_10235 ( SUB_1605_U320 , SUB_1605_U153 );
nand NAND2_10236 ( SUB_1605_U321 , SUB_1605_U114 , SUB_1605_U156 );
not NOT1_10237 ( SUB_1605_U322 , SUB_1605_U152 );
nand NAND2_10238 ( SUB_1605_U323 , SUB_1605_U127 , SUB_1605_U162 );
nand NAND2_10239 ( SUB_1605_U324 , P2_DATAO_REG_9_ , SUB_1605_U32 );
nand NAND2_10240 ( SUB_1605_U325 , P1_DATAO_REG_9_ , SUB_1605_U31 );
not NOT1_10241 ( SUB_1605_U326 , SUB_1605_U116 );
nand NAND2_10242 ( SUB_1605_U327 , SUB_1605_U322 , SUB_1605_U326 );
nand NAND2_10243 ( SUB_1605_U328 , SUB_1605_U116 , SUB_1605_U152 );
nand NAND2_10244 ( SUB_1605_U329 , P2_DATAO_REG_8_ , SUB_1605_U14 );
nand NAND2_10245 ( SUB_1605_U330 , P1_DATAO_REG_8_ , SUB_1605_U15 );
not NOT1_10246 ( SUB_1605_U331 , SUB_1605_U117 );
nand NAND2_10247 ( SUB_1605_U332 , SUB_1605_U320 , SUB_1605_U331 );
nand NAND2_10248 ( SUB_1605_U333 , SUB_1605_U117 , SUB_1605_U153 );
nand NAND2_10249 ( SUB_1605_U334 , P2_DATAO_REG_7_ , SUB_1605_U18 );
nand NAND2_10250 ( SUB_1605_U335 , P1_DATAO_REG_7_ , SUB_1605_U16 );
not NOT1_10251 ( SUB_1605_U336 , SUB_1605_U119 );
nand NAND2_10252 ( SUB_1605_U337 , SUB_1605_U318 , SUB_1605_U336 );
nand NAND2_10253 ( SUB_1605_U338 , SUB_1605_U119 , SUB_1605_U154 );
nand NAND2_10254 ( SUB_1605_U339 , P2_DATAO_REG_6_ , SUB_1605_U17 );
nand NAND2_10255 ( SUB_1605_U340 , P1_DATAO_REG_6_ , SUB_1605_U19 );
not NOT1_10256 ( SUB_1605_U341 , SUB_1605_U120 );
nand NAND2_10257 ( SUB_1605_U342 , SUB_1605_U316 , SUB_1605_U341 );
nand NAND2_10258 ( SUB_1605_U343 , SUB_1605_U120 , SUB_1605_U155 );
nand NAND2_10259 ( SUB_1605_U344 , P2_DATAO_REG_5_ , SUB_1605_U20 );
nand NAND2_10260 ( SUB_1605_U345 , P1_DATAO_REG_5_ , SUB_1605_U30 );
not NOT1_10261 ( SUB_1605_U346 , SUB_1605_U121 );
nand NAND2_10262 ( SUB_1605_U347 , SUB_1605_U199 , SUB_1605_U346 );
nand NAND2_10263 ( SUB_1605_U348 , SUB_1605_U121 , SUB_1605_U156 );
nand NAND2_10264 ( SUB_1605_U349 , P2_DATAO_REG_4_ , SUB_1605_U22 );
nand NAND2_10265 ( SUB_1605_U350 , P1_DATAO_REG_4_ , SUB_1605_U25 );
not NOT1_10266 ( SUB_1605_U351 , SUB_1605_U122 );
nand NAND2_10267 ( SUB_1605_U352 , SUB_1605_U196 , SUB_1605_U351 );
nand NAND2_10268 ( SUB_1605_U353 , SUB_1605_U122 , SUB_1605_U157 );
nand NAND2_10269 ( SUB_1605_U354 , P2_DATAO_REG_3_ , SUB_1605_U29 );
nand NAND2_10270 ( SUB_1605_U355 , P1_DATAO_REG_3_ , SUB_1605_U27 );
not NOT1_10271 ( SUB_1605_U356 , SUB_1605_U123 );
nand NAND2_10272 ( SUB_1605_U357 , SUB_1605_U193 , SUB_1605_U356 );
nand NAND2_10273 ( SUB_1605_U358 , SUB_1605_U123 , SUB_1605_U158 );
nand NAND2_10274 ( SUB_1605_U359 , P2_DATAO_REG_31_ , SUB_1605_U160 );
nand NAND2_10275 ( SUB_1605_U360 , P1_DATAO_REG_31_ , SUB_1605_U159 );
nand NAND2_10276 ( SUB_1605_U361 , SUB_1605_U360 , SUB_1605_U359 );
nand NAND2_10277 ( SUB_1605_U362 , P2_DATAO_REG_31_ , SUB_1605_U160 );
nand NAND2_10278 ( SUB_1605_U363 , P1_DATAO_REG_31_ , SUB_1605_U159 );
nand NAND3_10279 ( SUB_1605_U364 , P1_DATAO_REG_30_ , SUB_1605_U361 , SUB_1605_U75 );
nand NAND3_10280 ( SUB_1605_U365 , SUB_1605_U11 , SUB_1605_U74 , P2_DATAO_REG_30_ );
nand NAND2_10281 ( SUB_1605_U366 , P2_DATAO_REG_30_ , SUB_1605_U74 );
nand NAND2_10282 ( SUB_1605_U367 , P1_DATAO_REG_30_ , SUB_1605_U75 );
not NOT1_10283 ( SUB_1605_U368 , SUB_1605_U129 );
nand NAND2_10284 ( SUB_1605_U369 , SUB_1605_U288 , SUB_1605_U368 );
nand NAND2_10285 ( SUB_1605_U370 , SUB_1605_U129 , SUB_1605_U162 );
nand NAND2_10286 ( SUB_1605_U371 , P2_DATAO_REG_2_ , SUB_1605_U28 );
nand NAND2_10287 ( SUB_1605_U372 , P1_DATAO_REG_2_ , SUB_1605_U26 );
not NOT1_10288 ( SUB_1605_U373 , SUB_1605_U130 );
nand NAND2_10289 ( SUB_1605_U374 , SUB_1605_U189 , SUB_1605_U373 );
nand NAND2_10290 ( SUB_1605_U375 , SUB_1605_U130 , SUB_1605_U163 );
nand NAND2_10291 ( SUB_1605_U376 , P2_DATAO_REG_29_ , SUB_1605_U73 );
nand NAND2_10292 ( SUB_1605_U377 , P1_DATAO_REG_29_ , SUB_1605_U72 );
not NOT1_10293 ( SUB_1605_U378 , SUB_1605_U131 );
nand NAND2_10294 ( SUB_1605_U379 , SUB_1605_U284 , SUB_1605_U378 );
nand NAND2_10295 ( SUB_1605_U380 , SUB_1605_U131 , SUB_1605_U164 );
nand NAND2_10296 ( SUB_1605_U381 , P2_DATAO_REG_28_ , SUB_1605_U71 );
nand NAND2_10297 ( SUB_1605_U382 , P1_DATAO_REG_28_ , SUB_1605_U70 );
not NOT1_10298 ( SUB_1605_U383 , SUB_1605_U132 );
nand NAND2_10299 ( SUB_1605_U384 , SUB_1605_U280 , SUB_1605_U383 );
nand NAND2_10300 ( SUB_1605_U385 , SUB_1605_U132 , SUB_1605_U165 );
nand NAND2_10301 ( SUB_1605_U386 , P2_DATAO_REG_27_ , SUB_1605_U69 );
nand NAND2_10302 ( SUB_1605_U387 , P1_DATAO_REG_27_ , SUB_1605_U68 );
not NOT1_10303 ( SUB_1605_U388 , SUB_1605_U133 );
nand NAND2_10304 ( SUB_1605_U389 , SUB_1605_U276 , SUB_1605_U388 );
nand NAND2_10305 ( SUB_1605_U390 , SUB_1605_U133 , SUB_1605_U166 );
nand NAND2_10306 ( SUB_1605_U391 , P2_DATAO_REG_26_ , SUB_1605_U67 );
nand NAND2_10307 ( SUB_1605_U392 , P1_DATAO_REG_26_ , SUB_1605_U66 );
not NOT1_10308 ( SUB_1605_U393 , SUB_1605_U134 );
nand NAND2_10309 ( SUB_1605_U394 , SUB_1605_U272 , SUB_1605_U393 );
nand NAND2_10310 ( SUB_1605_U395 , SUB_1605_U134 , SUB_1605_U167 );
nand NAND2_10311 ( SUB_1605_U396 , P2_DATAO_REG_25_ , SUB_1605_U65 );
nand NAND2_10312 ( SUB_1605_U397 , P1_DATAO_REG_25_ , SUB_1605_U64 );
not NOT1_10313 ( SUB_1605_U398 , SUB_1605_U135 );
nand NAND2_10314 ( SUB_1605_U399 , SUB_1605_U268 , SUB_1605_U398 );
nand NAND2_10315 ( SUB_1605_U400 , SUB_1605_U135 , SUB_1605_U168 );
nand NAND2_10316 ( SUB_1605_U401 , P2_DATAO_REG_24_ , SUB_1605_U63 );
nand NAND2_10317 ( SUB_1605_U402 , P1_DATAO_REG_24_ , SUB_1605_U62 );
not NOT1_10318 ( SUB_1605_U403 , SUB_1605_U136 );
nand NAND2_10319 ( SUB_1605_U404 , SUB_1605_U264 , SUB_1605_U403 );
nand NAND2_10320 ( SUB_1605_U405 , SUB_1605_U136 , SUB_1605_U169 );
nand NAND2_10321 ( SUB_1605_U406 , P2_DATAO_REG_23_ , SUB_1605_U61 );
nand NAND2_10322 ( SUB_1605_U407 , P1_DATAO_REG_23_ , SUB_1605_U60 );
not NOT1_10323 ( SUB_1605_U408 , SUB_1605_U137 );
nand NAND2_10324 ( SUB_1605_U409 , SUB_1605_U260 , SUB_1605_U408 );
nand NAND2_10325 ( SUB_1605_U410 , SUB_1605_U137 , SUB_1605_U170 );
nand NAND2_10326 ( SUB_1605_U411 , P2_DATAO_REG_22_ , SUB_1605_U59 );
nand NAND2_10327 ( SUB_1605_U412 , P1_DATAO_REG_22_ , SUB_1605_U58 );
not NOT1_10328 ( SUB_1605_U413 , SUB_1605_U138 );
nand NAND2_10329 ( SUB_1605_U414 , SUB_1605_U256 , SUB_1605_U413 );
nand NAND2_10330 ( SUB_1605_U415 , SUB_1605_U138 , SUB_1605_U171 );
nand NAND2_10331 ( SUB_1605_U416 , P2_DATAO_REG_21_ , SUB_1605_U57 );
nand NAND2_10332 ( SUB_1605_U417 , P1_DATAO_REG_21_ , SUB_1605_U56 );
not NOT1_10333 ( SUB_1605_U418 , SUB_1605_U139 );
nand NAND2_10334 ( SUB_1605_U419 , SUB_1605_U252 , SUB_1605_U418 );
nand NAND2_10335 ( SUB_1605_U420 , SUB_1605_U139 , SUB_1605_U172 );
nand NAND2_10336 ( SUB_1605_U421 , P2_DATAO_REG_20_ , SUB_1605_U55 );
nand NAND2_10337 ( SUB_1605_U422 , P1_DATAO_REG_20_ , SUB_1605_U54 );
not NOT1_10338 ( SUB_1605_U423 , SUB_1605_U140 );
nand NAND2_10339 ( SUB_1605_U424 , SUB_1605_U248 , SUB_1605_U423 );
nand NAND2_10340 ( SUB_1605_U425 , SUB_1605_U140 , SUB_1605_U173 );
nand NAND2_10341 ( SUB_1605_U426 , P2_DATAO_REG_1_ , SUB_1605_U24 );
nand NAND2_10342 ( SUB_1605_U427 , P1_DATAO_REG_1_ , SUB_1605_U174 );
not NOT1_10343 ( SUB_1605_U428 , SUB_1605_U141 );
nand NAND2_10344 ( SUB_1605_U429 , SUB_1605_U187 , SUB_1605_U428 );
nand NAND2_10345 ( SUB_1605_U430 , SUB_1605_U141 , SUB_1605_U175 );
nand NAND2_10346 ( SUB_1605_U431 , P2_DATAO_REG_19_ , SUB_1605_U53 );
nand NAND2_10347 ( SUB_1605_U432 , P1_DATAO_REG_19_ , SUB_1605_U52 );
not NOT1_10348 ( SUB_1605_U433 , SUB_1605_U142 );
nand NAND2_10349 ( SUB_1605_U434 , SUB_1605_U244 , SUB_1605_U433 );
nand NAND2_10350 ( SUB_1605_U435 , SUB_1605_U142 , SUB_1605_U176 );
nand NAND2_10351 ( SUB_1605_U436 , P2_DATAO_REG_18_ , SUB_1605_U51 );
nand NAND2_10352 ( SUB_1605_U437 , P1_DATAO_REG_18_ , SUB_1605_U50 );
not NOT1_10353 ( SUB_1605_U438 , SUB_1605_U143 );
nand NAND2_10354 ( SUB_1605_U439 , SUB_1605_U240 , SUB_1605_U438 );
nand NAND2_10355 ( SUB_1605_U440 , SUB_1605_U143 , SUB_1605_U177 );
nand NAND2_10356 ( SUB_1605_U441 , P2_DATAO_REG_17_ , SUB_1605_U49 );
nand NAND2_10357 ( SUB_1605_U442 , P1_DATAO_REG_17_ , SUB_1605_U48 );
not NOT1_10358 ( SUB_1605_U443 , SUB_1605_U144 );
nand NAND2_10359 ( SUB_1605_U444 , SUB_1605_U236 , SUB_1605_U443 );
nand NAND2_10360 ( SUB_1605_U445 , SUB_1605_U144 , SUB_1605_U178 );
nand NAND2_10361 ( SUB_1605_U446 , P2_DATAO_REG_16_ , SUB_1605_U47 );
nand NAND2_10362 ( SUB_1605_U447 , P1_DATAO_REG_16_ , SUB_1605_U46 );
not NOT1_10363 ( SUB_1605_U448 , SUB_1605_U145 );
nand NAND2_10364 ( SUB_1605_U449 , SUB_1605_U232 , SUB_1605_U448 );
nand NAND2_10365 ( SUB_1605_U450 , SUB_1605_U145 , SUB_1605_U179 );
nand NAND2_10366 ( SUB_1605_U451 , P2_DATAO_REG_15_ , SUB_1605_U45 );
nand NAND2_10367 ( SUB_1605_U452 , P1_DATAO_REG_15_ , SUB_1605_U44 );
not NOT1_10368 ( SUB_1605_U453 , SUB_1605_U146 );
nand NAND2_10369 ( SUB_1605_U454 , SUB_1605_U228 , SUB_1605_U453 );
nand NAND2_10370 ( SUB_1605_U455 , SUB_1605_U146 , SUB_1605_U180 );
nand NAND2_10371 ( SUB_1605_U456 , P2_DATAO_REG_14_ , SUB_1605_U43 );
nand NAND2_10372 ( SUB_1605_U457 , P1_DATAO_REG_14_ , SUB_1605_U42 );
not NOT1_10373 ( SUB_1605_U458 , SUB_1605_U147 );
nand NAND2_10374 ( SUB_1605_U459 , SUB_1605_U224 , SUB_1605_U458 );
nand NAND2_10375 ( SUB_1605_U460 , SUB_1605_U147 , SUB_1605_U181 );
nand NAND2_10376 ( SUB_1605_U461 , P2_DATAO_REG_13_ , SUB_1605_U41 );
nand NAND2_10377 ( SUB_1605_U462 , P1_DATAO_REG_13_ , SUB_1605_U40 );
not NOT1_10378 ( SUB_1605_U463 , SUB_1605_U148 );
nand NAND2_10379 ( SUB_1605_U464 , SUB_1605_U220 , SUB_1605_U463 );
nand NAND2_10380 ( SUB_1605_U465 , SUB_1605_U148 , SUB_1605_U182 );
nand NAND2_10381 ( SUB_1605_U466 , P2_DATAO_REG_12_ , SUB_1605_U33 );
nand NAND2_10382 ( SUB_1605_U467 , P1_DATAO_REG_12_ , SUB_1605_U34 );
not NOT1_10383 ( SUB_1605_U468 , SUB_1605_U149 );
nand NAND2_10384 ( SUB_1605_U469 , SUB_1605_U217 , SUB_1605_U468 );
nand NAND2_10385 ( SUB_1605_U470 , SUB_1605_U149 , SUB_1605_U183 );
nand NAND2_10386 ( SUB_1605_U471 , P2_DATAO_REG_11_ , SUB_1605_U37 );
nand NAND2_10387 ( SUB_1605_U472 , P1_DATAO_REG_11_ , SUB_1605_U35 );
not NOT1_10388 ( SUB_1605_U473 , SUB_1605_U150 );
nand NAND2_10389 ( SUB_1605_U474 , SUB_1605_U214 , SUB_1605_U473 );
nand NAND2_10390 ( SUB_1605_U475 , SUB_1605_U150 , SUB_1605_U184 );
nand NAND2_10391 ( SUB_1605_U476 , P2_DATAO_REG_10_ , SUB_1605_U38 );
nand NAND2_10392 ( SUB_1605_U477 , P1_DATAO_REG_10_ , SUB_1605_U36 );
not NOT1_10393 ( SUB_1605_U478 , SUB_1605_U151 );
nand NAND2_10394 ( SUB_1605_U479 , SUB_1605_U211 , SUB_1605_U478 );
nand NAND2_10395 ( SUB_1605_U480 , SUB_1605_U151 , SUB_1605_U185 );
and AND2_10396 ( R152_U4 , R152_U206 , R152_U202 );
and AND2_10397 ( R152_U5 , R152_U214 , R152_U212 );
and AND2_10398 ( R152_U6 , R152_U5 , R152_U216 );
and AND2_10399 ( R152_U7 , R152_U222 , R152_U220 );
and AND2_10400 ( R152_U8 , R152_U7 , R152_U224 );
and AND2_10401 ( R152_U9 , R152_U8 , R152_U226 );
and AND2_10402 ( R152_U10 , R152_U199 , R152_U196 );
and AND2_10403 ( R152_U11 , R152_U391 , R152_U390 );
and AND2_10404 ( R152_U12 , R152_U128 , R152_U193 );
nand NAND2_10405 ( R152_U13 , R152_U172 , R152_U337 );
not NOT1_10406 ( R152_U14 , SI_8_ );
not NOT1_10407 ( R152_U15 , U127 );
not NOT1_10408 ( R152_U16 , SI_7_ );
not NOT1_10409 ( R152_U17 , U128 );
nand NAND2_10410 ( R152_U18 , U128 , SI_7_ );
not NOT1_10411 ( R152_U19 , SI_6_ );
not NOT1_10412 ( R152_U20 , U129 );
not NOT1_10413 ( R152_U21 , SI_3_ );
not NOT1_10414 ( R152_U22 , U134 );
not NOT1_10415 ( R152_U23 , SI_1_ );
not NOT1_10416 ( R152_U24 , SI_0_ );
not NOT1_10417 ( R152_U25 , U157 );
not NOT1_10418 ( R152_U26 , U156 );
not NOT1_10419 ( R152_U27 , SI_2_ );
not NOT1_10420 ( R152_U28 , U145 );
nand NAND2_10421 ( R152_U29 , U145 , SI_2_ );
not NOT1_10422 ( R152_U30 , SI_5_ );
not NOT1_10423 ( R152_U31 , U130 );
not NOT1_10424 ( R152_U32 , SI_4_ );
not NOT1_10425 ( R152_U33 , U131 );
nand NAND2_10426 ( R152_U34 , U131 , SI_4_ );
not NOT1_10427 ( R152_U35 , U126 );
not NOT1_10428 ( R152_U36 , SI_9_ );
nand NAND2_10429 ( R152_U37 , R152_U294 , R152_U207 );
not NOT1_10430 ( R152_U38 , SI_15_ );
not NOT1_10431 ( R152_U39 , U150 );
not NOT1_10432 ( R152_U40 , SI_14_ );
not NOT1_10433 ( R152_U41 , U151 );
not NOT1_10434 ( R152_U42 , SI_13_ );
not NOT1_10435 ( R152_U43 , U152 );
not NOT1_10436 ( R152_U44 , SI_12_ );
not NOT1_10437 ( R152_U45 , U153 );
not NOT1_10438 ( R152_U46 , SI_11_ );
not NOT1_10439 ( R152_U47 , U154 );
nand NAND2_10440 ( R152_U48 , U154 , SI_11_ );
not NOT1_10441 ( R152_U49 , SI_10_ );
not NOT1_10442 ( R152_U50 , U155 );
not NOT1_10443 ( R152_U51 , SI_16_ );
not NOT1_10444 ( R152_U52 , U149 );
not NOT1_10445 ( R152_U53 , SI_17_ );
not NOT1_10446 ( R152_U54 , U148 );
not NOT1_10447 ( R152_U55 , SI_18_ );
not NOT1_10448 ( R152_U56 , U147 );
not NOT1_10449 ( R152_U57 , SI_19_ );
not NOT1_10450 ( R152_U58 , U146 );
not NOT1_10451 ( R152_U59 , SI_20_ );
not NOT1_10452 ( R152_U60 , U144 );
not NOT1_10453 ( R152_U61 , SI_21_ );
not NOT1_10454 ( R152_U62 , U143 );
not NOT1_10455 ( R152_U63 , SI_22_ );
not NOT1_10456 ( R152_U64 , U142 );
not NOT1_10457 ( R152_U65 , SI_23_ );
not NOT1_10458 ( R152_U66 , U141 );
not NOT1_10459 ( R152_U67 , SI_24_ );
not NOT1_10460 ( R152_U68 , U140 );
not NOT1_10461 ( R152_U69 , SI_25_ );
not NOT1_10462 ( R152_U70 , U139 );
not NOT1_10463 ( R152_U71 , SI_26_ );
not NOT1_10464 ( R152_U72 , U138 );
not NOT1_10465 ( R152_U73 , SI_27_ );
not NOT1_10466 ( R152_U74 , U137 );
not NOT1_10467 ( R152_U75 , SI_28_ );
not NOT1_10468 ( R152_U76 , U136 );
not NOT1_10469 ( R152_U77 , SI_29_ );
not NOT1_10470 ( R152_U78 , U135 );
not NOT1_10471 ( R152_U79 , SI_30_ );
not NOT1_10472 ( R152_U80 , U133 );
nand NAND2_10473 ( R152_U81 , R152_U307 , R152_U227 );
nand NAND2_10474 ( R152_U82 , R152_U305 , R152_U225 );
nand NAND2_10475 ( R152_U83 , R152_U300 , R152_U217 );
nand NAND2_10476 ( R152_U84 , R152_U554 , R152_U553 );
nand NAND2_10477 ( R152_U85 , R152_U344 , R152_U343 );
nand NAND2_10478 ( R152_U86 , R152_U351 , R152_U350 );
nand NAND2_10479 ( R152_U87 , R152_U358 , R152_U357 );
nand NAND2_10480 ( R152_U88 , R152_U365 , R152_U364 );
nand NAND2_10481 ( R152_U89 , R152_U372 , R152_U371 );
nand NAND2_10482 ( R152_U90 , R152_U379 , R152_U378 );
nand NAND2_10483 ( R152_U91 , R152_U386 , R152_U385 );
nand NAND2_10484 ( R152_U92 , R152_U400 , R152_U399 );
nand NAND2_10485 ( R152_U93 , R152_U407 , R152_U406 );
nand NAND2_10486 ( R152_U94 , R152_U414 , R152_U413 );
nand NAND2_10487 ( R152_U95 , R152_U421 , R152_U420 );
nand NAND2_10488 ( R152_U96 , R152_U428 , R152_U427 );
nand NAND2_10489 ( R152_U97 , R152_U435 , R152_U434 );
nand NAND2_10490 ( R152_U98 , R152_U442 , R152_U441 );
nand NAND2_10491 ( R152_U99 , R152_U449 , R152_U448 );
nand NAND2_10492 ( R152_U100 , R152_U456 , R152_U455 );
nand NAND2_10493 ( R152_U101 , R152_U463 , R152_U462 );
nand NAND2_10494 ( R152_U102 , R152_U470 , R152_U469 );
nand NAND2_10495 ( R152_U103 , R152_U477 , R152_U476 );
nand NAND2_10496 ( R152_U104 , R152_U489 , R152_U488 );
nand NAND2_10497 ( R152_U105 , R152_U496 , R152_U495 );
nand NAND2_10498 ( R152_U106 , R152_U503 , R152_U502 );
nand NAND2_10499 ( R152_U107 , R152_U510 , R152_U509 );
nand NAND2_10500 ( R152_U108 , R152_U517 , R152_U516 );
nand NAND2_10501 ( R152_U109 , R152_U524 , R152_U523 );
nand NAND2_10502 ( R152_U110 , R152_U531 , R152_U530 );
nand NAND2_10503 ( R152_U111 , R152_U538 , R152_U537 );
nand NAND2_10504 ( R152_U112 , R152_U545 , R152_U544 );
nand NAND2_10505 ( R152_U113 , R152_U552 , R152_U551 );
and AND2_10506 ( R152_U114 , R152_U292 , R152_U200 );
and AND2_10507 ( R152_U115 , R152_U209 , R152_U4 );
and AND2_10508 ( R152_U116 , R152_U297 , R152_U210 );
and AND2_10509 ( R152_U117 , R152_U298 , R152_U215 );
and AND2_10510 ( R152_U118 , R152_U292 , R152_U200 );
and AND2_10511 ( R152_U119 , U156 , U157 );
and AND2_10512 ( R152_U120 , U157 , SI_0_ );
and AND2_10513 ( R152_U121 , SI_1_ , U156 );
and AND2_10514 ( R152_U122 , R152_U218 , R152_U6 );
and AND2_10515 ( R152_U123 , R152_U302 , R152_U219 );
and AND2_10516 ( R152_U124 , R152_U9 , R152_U228 );
and AND2_10517 ( R152_U125 , R152_U309 , R152_U229 );
and AND2_10518 ( R152_U126 , R152_U287 , R152_U389 );
and AND3_10519 ( R152_U127 , R152_U11 , R152_U286 , R152_U284 );
and AND2_10520 ( R152_U128 , R152_U288 , R152_U146 );
and AND2_10521 ( R152_U129 , R152_U303 , R152_U223 );
and AND2_10522 ( R152_U130 , R152_U339 , R152_U338 );
nand NAND2_10523 ( R152_U131 , R152_U117 , R152_U331 );
and AND2_10524 ( R152_U132 , R152_U346 , R152_U345 );
nand NAND2_10525 ( R152_U133 , R152_U329 , R152_U18 );
and AND2_10526 ( R152_U134 , R152_U353 , R152_U352 );
nand NAND2_10527 ( R152_U135 , R152_U116 , R152_U296 );
and AND2_10528 ( R152_U136 , R152_U360 , R152_U359 );
nand NAND2_10529 ( R152_U137 , R152_U295 , R152_U293 );
and AND2_10530 ( R152_U138 , R152_U367 , R152_U366 );
nand NAND2_10531 ( R152_U139 , R152_U34 , R152_U203 );
and AND2_10532 ( R152_U140 , R152_U374 , R152_U373 );
nand NAND2_10533 ( R152_U141 , R152_U118 , R152_U315 );
and AND2_10534 ( R152_U142 , R152_U381 , R152_U380 );
nand NAND4_10535 ( R152_U143 , R152_U312 , R152_U311 , R152_U310 , R152_U29 );
not NOT1_10536 ( R152_U144 , U132 );
not NOT1_10537 ( R152_U145 , SI_31_ );
and AND2_10538 ( R152_U146 , R152_U393 , R152_U392 );
and AND2_10539 ( R152_U147 , R152_U395 , R152_U394 );
nand NAND2_10540 ( R152_U148 , R152_U284 , R152_U283 );
nand NAND3_10541 ( R152_U149 , R152_U290 , R152_U171 , R152_U289 );
and AND2_10542 ( R152_U150 , R152_U409 , R152_U408 );
nand NAND2_10543 ( R152_U151 , R152_U280 , R152_U279 );
and AND2_10544 ( R152_U152 , R152_U416 , R152_U415 );
nand NAND2_10545 ( R152_U153 , R152_U276 , R152_U275 );
and AND2_10546 ( R152_U154 , R152_U423 , R152_U422 );
nand NAND2_10547 ( R152_U155 , R152_U272 , R152_U271 );
and AND2_10548 ( R152_U156 , R152_U430 , R152_U429 );
nand NAND2_10549 ( R152_U157 , R152_U268 , R152_U267 );
and AND2_10550 ( R152_U158 , R152_U437 , R152_U436 );
nand NAND2_10551 ( R152_U159 , R152_U264 , R152_U263 );
and AND2_10552 ( R152_U160 , R152_U444 , R152_U443 );
nand NAND2_10553 ( R152_U161 , R152_U260 , R152_U259 );
and AND2_10554 ( R152_U162 , R152_U451 , R152_U450 );
nand NAND2_10555 ( R152_U163 , R152_U256 , R152_U255 );
and AND2_10556 ( R152_U164 , R152_U458 , R152_U457 );
nand NAND2_10557 ( R152_U165 , R152_U252 , R152_U251 );
and AND2_10558 ( R152_U166 , R152_U465 , R152_U464 );
nand NAND2_10559 ( R152_U167 , R152_U248 , R152_U247 );
and AND2_10560 ( R152_U168 , R152_U472 , R152_U471 );
nand NAND2_10561 ( R152_U169 , R152_U244 , R152_U243 );
nand NAND2_10562 ( R152_U170 , U157 , SI_0_ );
nand NAND3_10563 ( R152_U171 , SI_0_ , SI_1_ , U157 );
and AND2_10564 ( R152_U172 , R152_U482 , R152_U481 );
and AND2_10565 ( R152_U173 , R152_U484 , R152_U483 );
nand NAND2_10566 ( R152_U174 , R152_U240 , R152_U239 );
and AND2_10567 ( R152_U175 , R152_U491 , R152_U490 );
nand NAND2_10568 ( R152_U176 , R152_U236 , R152_U235 );
and AND2_10569 ( R152_U177 , R152_U498 , R152_U497 );
nand NAND2_10570 ( R152_U178 , R152_U232 , R152_U231 );
and AND2_10571 ( R152_U179 , R152_U505 , R152_U504 );
nand NAND2_10572 ( R152_U180 , R152_U125 , R152_U327 );
and AND2_10573 ( R152_U181 , R152_U512 , R152_U511 );
nand NAND2_10574 ( R152_U182 , R152_U308 , R152_U325 );
and AND2_10575 ( R152_U183 , R152_U519 , R152_U518 );
nand NAND2_10576 ( R152_U184 , R152_U306 , R152_U323 );
and AND2_10577 ( R152_U185 , R152_U526 , R152_U525 );
nand NAND2_10578 ( R152_U186 , R152_U129 , R152_U321 );
and AND2_10579 ( R152_U187 , R152_U533 , R152_U532 );
nand NAND2_10580 ( R152_U188 , R152_U319 , R152_U48 );
and AND2_10581 ( R152_U189 , R152_U540 , R152_U539 );
nand NAND2_10582 ( R152_U190 , R152_U123 , R152_U335 );
and AND2_10583 ( R152_U191 , R152_U547 , R152_U546 );
nand NAND2_10584 ( R152_U192 , R152_U301 , R152_U333 );
nand NAND2_10585 ( R152_U193 , R152_U126 , R152_U148 );
not NOT1_10586 ( R152_U194 , R152_U171 );
not NOT1_10587 ( R152_U195 , R152_U149 );
or OR2_10588 ( R152_U196 , SI_2_ , U145 );
not NOT1_10589 ( R152_U197 , R152_U29 );
not NOT1_10590 ( R152_U198 , R152_U143 );
or OR2_10591 ( R152_U199 , SI_3_ , U134 );
nand NAND2_10592 ( R152_U200 , U134 , SI_3_ );
nand NAND2_10593 ( R152_U201 , R152_U114 , R152_U291 );
or OR2_10594 ( R152_U202 , SI_4_ , U131 );
nand NAND2_10595 ( R152_U203 , R152_U202 , R152_U201 );
not NOT1_10596 ( R152_U204 , R152_U34 );
not NOT1_10597 ( R152_U205 , R152_U139 );
or OR2_10598 ( R152_U206 , SI_5_ , U130 );
nand NAND2_10599 ( R152_U207 , U130 , SI_5_ );
not NOT1_10600 ( R152_U208 , R152_U137 );
or OR2_10601 ( R152_U209 , SI_6_ , U129 );
nand NAND2_10602 ( R152_U210 , U129 , SI_6_ );
not NOT1_10603 ( R152_U211 , R152_U135 );
or OR2_10604 ( R152_U212 , SI_7_ , U128 );
not NOT1_10605 ( R152_U213 , R152_U18 );
or OR2_10606 ( R152_U214 , SI_8_ , U127 );
nand NAND2_10607 ( R152_U215 , U127 , SI_8_ );
or OR2_10608 ( R152_U216 , SI_9_ , U126 );
nand NAND2_10609 ( R152_U217 , SI_9_ , U126 );
or OR2_10610 ( R152_U218 , SI_10_ , U155 );
nand NAND2_10611 ( R152_U219 , U155 , SI_10_ );
or OR2_10612 ( R152_U220 , SI_11_ , U154 );
not NOT1_10613 ( R152_U221 , R152_U48 );
or OR2_10614 ( R152_U222 , SI_12_ , U153 );
nand NAND2_10615 ( R152_U223 , U153 , SI_12_ );
or OR2_10616 ( R152_U224 , SI_13_ , U152 );
nand NAND2_10617 ( R152_U225 , U152 , SI_13_ );
or OR2_10618 ( R152_U226 , SI_14_ , U151 );
nand NAND2_10619 ( R152_U227 , U151 , SI_14_ );
or OR2_10620 ( R152_U228 , SI_15_ , U150 );
nand NAND2_10621 ( R152_U229 , U150 , SI_15_ );
or OR2_10622 ( R152_U230 , SI_16_ , U149 );
nand NAND2_10623 ( R152_U231 , R152_U230 , R152_U180 );
nand NAND2_10624 ( R152_U232 , U149 , SI_16_ );
not NOT1_10625 ( R152_U233 , R152_U178 );
or OR2_10626 ( R152_U234 , SI_17_ , U148 );
nand NAND2_10627 ( R152_U235 , R152_U234 , R152_U178 );
nand NAND2_10628 ( R152_U236 , U148 , SI_17_ );
not NOT1_10629 ( R152_U237 , R152_U176 );
or OR2_10630 ( R152_U238 , SI_18_ , U147 );
nand NAND2_10631 ( R152_U239 , R152_U238 , R152_U176 );
nand NAND2_10632 ( R152_U240 , U147 , SI_18_ );
not NOT1_10633 ( R152_U241 , R152_U174 );
or OR2_10634 ( R152_U242 , SI_19_ , U146 );
nand NAND2_10635 ( R152_U243 , R152_U242 , R152_U174 );
nand NAND2_10636 ( R152_U244 , U146 , SI_19_ );
not NOT1_10637 ( R152_U245 , R152_U169 );
or OR2_10638 ( R152_U246 , SI_20_ , U144 );
nand NAND2_10639 ( R152_U247 , R152_U246 , R152_U169 );
nand NAND2_10640 ( R152_U248 , U144 , SI_20_ );
not NOT1_10641 ( R152_U249 , R152_U167 );
or OR2_10642 ( R152_U250 , SI_21_ , U143 );
nand NAND2_10643 ( R152_U251 , R152_U250 , R152_U167 );
nand NAND2_10644 ( R152_U252 , U143 , SI_21_ );
not NOT1_10645 ( R152_U253 , R152_U165 );
or OR2_10646 ( R152_U254 , SI_22_ , U142 );
nand NAND2_10647 ( R152_U255 , R152_U254 , R152_U165 );
nand NAND2_10648 ( R152_U256 , U142 , SI_22_ );
not NOT1_10649 ( R152_U257 , R152_U163 );
or OR2_10650 ( R152_U258 , SI_23_ , U141 );
nand NAND2_10651 ( R152_U259 , R152_U258 , R152_U163 );
nand NAND2_10652 ( R152_U260 , U141 , SI_23_ );
not NOT1_10653 ( R152_U261 , R152_U161 );
or OR2_10654 ( R152_U262 , SI_24_ , U140 );
nand NAND2_10655 ( R152_U263 , R152_U262 , R152_U161 );
nand NAND2_10656 ( R152_U264 , U140 , SI_24_ );
not NOT1_10657 ( R152_U265 , R152_U159 );
or OR2_10658 ( R152_U266 , SI_25_ , U139 );
nand NAND2_10659 ( R152_U267 , R152_U266 , R152_U159 );
nand NAND2_10660 ( R152_U268 , U139 , SI_25_ );
not NOT1_10661 ( R152_U269 , R152_U157 );
or OR2_10662 ( R152_U270 , SI_26_ , U138 );
nand NAND2_10663 ( R152_U271 , R152_U270 , R152_U157 );
nand NAND2_10664 ( R152_U272 , U138 , SI_26_ );
not NOT1_10665 ( R152_U273 , R152_U155 );
or OR2_10666 ( R152_U274 , SI_27_ , U137 );
nand NAND2_10667 ( R152_U275 , R152_U274 , R152_U155 );
nand NAND2_10668 ( R152_U276 , U137 , SI_27_ );
not NOT1_10669 ( R152_U277 , R152_U153 );
or OR2_10670 ( R152_U278 , SI_28_ , U136 );
nand NAND2_10671 ( R152_U279 , R152_U278 , R152_U153 );
nand NAND2_10672 ( R152_U280 , U136 , SI_28_ );
not NOT1_10673 ( R152_U281 , R152_U151 );
or OR2_10674 ( R152_U282 , SI_29_ , U135 );
nand NAND2_10675 ( R152_U283 , R152_U282 , R152_U151 );
nand NAND2_10676 ( R152_U284 , U135 , SI_29_ );
not NOT1_10677 ( R152_U285 , R152_U148 );
nand NAND2_10678 ( R152_U286 , U133 , SI_30_ );
or OR2_10679 ( R152_U287 , U133 , SI_30_ );
nand NAND2_10680 ( R152_U288 , R152_U283 , R152_U127 );
nand NAND3_10681 ( R152_U289 , U157 , SI_0_ , U156 );
nand NAND2_10682 ( R152_U290 , U156 , SI_1_ );
nand NAND2_10683 ( R152_U291 , R152_U10 , R152_U313 );
nand NAND2_10684 ( R152_U292 , R152_U197 , R152_U199 );
nand NAND2_10685 ( R152_U293 , R152_U4 , R152_U201 );
nand NAND2_10686 ( R152_U294 , R152_U204 , R152_U206 );
not NOT1_10687 ( R152_U295 , R152_U37 );
nand NAND2_10688 ( R152_U296 , R152_U115 , R152_U201 );
nand NAND2_10689 ( R152_U297 , R152_U37 , R152_U209 );
nand NAND2_10690 ( R152_U298 , R152_U213 , R152_U214 );
nand NAND2_10691 ( R152_U299 , R152_U298 , R152_U215 );
nand NAND2_10692 ( R152_U300 , R152_U299 , R152_U216 );
not NOT1_10693 ( R152_U301 , R152_U83 );
nand NAND2_10694 ( R152_U302 , R152_U83 , R152_U218 );
nand NAND2_10695 ( R152_U303 , R152_U221 , R152_U222 );
nand NAND2_10696 ( R152_U304 , R152_U303 , R152_U223 );
nand NAND2_10697 ( R152_U305 , R152_U304 , R152_U224 );
not NOT1_10698 ( R152_U306 , R152_U82 );
nand NAND2_10699 ( R152_U307 , R152_U82 , R152_U226 );
not NOT1_10700 ( R152_U308 , R152_U81 );
nand NAND2_10701 ( R152_U309 , R152_U81 , R152_U228 );
nand NAND3_10702 ( R152_U310 , SI_0_ , R152_U196 , R152_U119 );
nand NAND3_10703 ( R152_U311 , SI_1_ , R152_U196 , R152_U120 );
nand NAND2_10704 ( R152_U312 , R152_U121 , R152_U196 );
nand NAND3_10705 ( R152_U313 , R152_U290 , R152_U171 , R152_U289 );
not NOT1_10706 ( R152_U314 , R152_U141 );
nand NAND2_10707 ( R152_U315 , R152_U10 , R152_U316 );
nand NAND3_10708 ( R152_U316 , R152_U318 , R152_U290 , R152_U317 );
nand NAND3_10709 ( R152_U317 , U157 , SI_0_ , U156 );
nand NAND3_10710 ( R152_U318 , SI_0_ , SI_1_ , U157 );
nand NAND2_10711 ( R152_U319 , R152_U220 , R152_U190 );
not NOT1_10712 ( R152_U320 , R152_U188 );
nand NAND2_10713 ( R152_U321 , R152_U7 , R152_U190 );
not NOT1_10714 ( R152_U322 , R152_U186 );
nand NAND2_10715 ( R152_U323 , R152_U8 , R152_U190 );
not NOT1_10716 ( R152_U324 , R152_U184 );
nand NAND2_10717 ( R152_U325 , R152_U9 , R152_U190 );
not NOT1_10718 ( R152_U326 , R152_U182 );
nand NAND2_10719 ( R152_U327 , R152_U124 , R152_U190 );
not NOT1_10720 ( R152_U328 , R152_U180 );
nand NAND2_10721 ( R152_U329 , R152_U212 , R152_U135 );
not NOT1_10722 ( R152_U330 , R152_U133 );
nand NAND2_10723 ( R152_U331 , R152_U5 , R152_U135 );
not NOT1_10724 ( R152_U332 , R152_U131 );
nand NAND2_10725 ( R152_U333 , R152_U6 , R152_U135 );
not NOT1_10726 ( R152_U334 , R152_U192 );
nand NAND2_10727 ( R152_U335 , R152_U122 , R152_U135 );
not NOT1_10728 ( R152_U336 , R152_U190 );
nand NAND2_10729 ( R152_U337 , R152_U480 , R152_U23 );
nand NAND2_10730 ( R152_U338 , U126 , R152_U36 );
nand NAND2_10731 ( R152_U339 , SI_9_ , R152_U35 );
nand NAND2_10732 ( R152_U340 , U126 , R152_U36 );
nand NAND2_10733 ( R152_U341 , SI_9_ , R152_U35 );
nand NAND2_10734 ( R152_U342 , R152_U341 , R152_U340 );
nand NAND2_10735 ( R152_U343 , R152_U130 , R152_U131 );
nand NAND2_10736 ( R152_U344 , R152_U332 , R152_U342 );
nand NAND2_10737 ( R152_U345 , U127 , R152_U14 );
nand NAND2_10738 ( R152_U346 , SI_8_ , R152_U15 );
nand NAND2_10739 ( R152_U347 , U127 , R152_U14 );
nand NAND2_10740 ( R152_U348 , SI_8_ , R152_U15 );
nand NAND2_10741 ( R152_U349 , R152_U348 , R152_U347 );
nand NAND2_10742 ( R152_U350 , R152_U132 , R152_U133 );
nand NAND2_10743 ( R152_U351 , R152_U330 , R152_U349 );
nand NAND2_10744 ( R152_U352 , U128 , R152_U16 );
nand NAND2_10745 ( R152_U353 , SI_7_ , R152_U17 );
nand NAND2_10746 ( R152_U354 , U128 , R152_U16 );
nand NAND2_10747 ( R152_U355 , SI_7_ , R152_U17 );
nand NAND2_10748 ( R152_U356 , R152_U355 , R152_U354 );
nand NAND2_10749 ( R152_U357 , R152_U134 , R152_U135 );
nand NAND2_10750 ( R152_U358 , R152_U211 , R152_U356 );
nand NAND2_10751 ( R152_U359 , U129 , R152_U19 );
nand NAND2_10752 ( R152_U360 , SI_6_ , R152_U20 );
nand NAND2_10753 ( R152_U361 , U129 , R152_U19 );
nand NAND2_10754 ( R152_U362 , SI_6_ , R152_U20 );
nand NAND2_10755 ( R152_U363 , R152_U362 , R152_U361 );
nand NAND2_10756 ( R152_U364 , R152_U136 , R152_U137 );
nand NAND2_10757 ( R152_U365 , R152_U208 , R152_U363 );
nand NAND2_10758 ( R152_U366 , U130 , R152_U30 );
nand NAND2_10759 ( R152_U367 , SI_5_ , R152_U31 );
nand NAND2_10760 ( R152_U368 , U130 , R152_U30 );
nand NAND2_10761 ( R152_U369 , SI_5_ , R152_U31 );
nand NAND2_10762 ( R152_U370 , R152_U369 , R152_U368 );
nand NAND2_10763 ( R152_U371 , R152_U138 , R152_U139 );
nand NAND2_10764 ( R152_U372 , R152_U205 , R152_U370 );
nand NAND2_10765 ( R152_U373 , U131 , R152_U32 );
nand NAND2_10766 ( R152_U374 , SI_4_ , R152_U33 );
nand NAND2_10767 ( R152_U375 , U131 , R152_U32 );
nand NAND2_10768 ( R152_U376 , SI_4_ , R152_U33 );
nand NAND2_10769 ( R152_U377 , R152_U376 , R152_U375 );
nand NAND2_10770 ( R152_U378 , R152_U140 , R152_U141 );
nand NAND2_10771 ( R152_U379 , R152_U314 , R152_U377 );
nand NAND2_10772 ( R152_U380 , U134 , R152_U21 );
nand NAND2_10773 ( R152_U381 , SI_3_ , R152_U22 );
nand NAND2_10774 ( R152_U382 , U134 , R152_U21 );
nand NAND2_10775 ( R152_U383 , SI_3_ , R152_U22 );
nand NAND2_10776 ( R152_U384 , R152_U383 , R152_U382 );
nand NAND2_10777 ( R152_U385 , R152_U142 , R152_U143 );
nand NAND2_10778 ( R152_U386 , R152_U198 , R152_U384 );
nand NAND2_10779 ( R152_U387 , U132 , R152_U145 );
nand NAND2_10780 ( R152_U388 , SI_31_ , R152_U144 );
nand NAND2_10781 ( R152_U389 , R152_U388 , R152_U387 );
nand NAND2_10782 ( R152_U390 , U132 , R152_U145 );
nand NAND2_10783 ( R152_U391 , SI_31_ , R152_U144 );
nand NAND3_10784 ( R152_U392 , R152_U11 , R152_U79 , R152_U80 );
nand NAND3_10785 ( R152_U393 , SI_30_ , R152_U389 , U133 );
nand NAND2_10786 ( R152_U394 , U133 , R152_U79 );
nand NAND2_10787 ( R152_U395 , SI_30_ , R152_U80 );
nand NAND2_10788 ( R152_U396 , U133 , R152_U79 );
nand NAND2_10789 ( R152_U397 , SI_30_ , R152_U80 );
nand NAND2_10790 ( R152_U398 , R152_U397 , R152_U396 );
nand NAND2_10791 ( R152_U399 , R152_U147 , R152_U148 );
nand NAND2_10792 ( R152_U400 , R152_U285 , R152_U398 );
nand NAND2_10793 ( R152_U401 , U145 , R152_U27 );
nand NAND2_10794 ( R152_U402 , SI_2_ , R152_U28 );
nand NAND2_10795 ( R152_U403 , U145 , R152_U27 );
nand NAND2_10796 ( R152_U404 , SI_2_ , R152_U28 );
nand NAND2_10797 ( R152_U405 , R152_U404 , R152_U403 );
nand NAND3_10798 ( R152_U406 , R152_U402 , R152_U401 , R152_U149 );
nand NAND2_10799 ( R152_U407 , R152_U195 , R152_U405 );
nand NAND2_10800 ( R152_U408 , U135 , R152_U77 );
nand NAND2_10801 ( R152_U409 , SI_29_ , R152_U78 );
nand NAND2_10802 ( R152_U410 , U135 , R152_U77 );
nand NAND2_10803 ( R152_U411 , SI_29_ , R152_U78 );
nand NAND2_10804 ( R152_U412 , R152_U411 , R152_U410 );
nand NAND2_10805 ( R152_U413 , R152_U150 , R152_U151 );
nand NAND2_10806 ( R152_U414 , R152_U281 , R152_U412 );
nand NAND2_10807 ( R152_U415 , U136 , R152_U75 );
nand NAND2_10808 ( R152_U416 , SI_28_ , R152_U76 );
nand NAND2_10809 ( R152_U417 , U136 , R152_U75 );
nand NAND2_10810 ( R152_U418 , SI_28_ , R152_U76 );
nand NAND2_10811 ( R152_U419 , R152_U418 , R152_U417 );
nand NAND2_10812 ( R152_U420 , R152_U152 , R152_U153 );
nand NAND2_10813 ( R152_U421 , R152_U277 , R152_U419 );
nand NAND2_10814 ( R152_U422 , U137 , R152_U73 );
nand NAND2_10815 ( R152_U423 , SI_27_ , R152_U74 );
nand NAND2_10816 ( R152_U424 , U137 , R152_U73 );
nand NAND2_10817 ( R152_U425 , SI_27_ , R152_U74 );
nand NAND2_10818 ( R152_U426 , R152_U425 , R152_U424 );
nand NAND2_10819 ( R152_U427 , R152_U154 , R152_U155 );
nand NAND2_10820 ( R152_U428 , R152_U273 , R152_U426 );
nand NAND2_10821 ( R152_U429 , U138 , R152_U71 );
nand NAND2_10822 ( R152_U430 , SI_26_ , R152_U72 );
nand NAND2_10823 ( R152_U431 , U138 , R152_U71 );
nand NAND2_10824 ( R152_U432 , SI_26_ , R152_U72 );
nand NAND2_10825 ( R152_U433 , R152_U432 , R152_U431 );
nand NAND2_10826 ( R152_U434 , R152_U156 , R152_U157 );
nand NAND2_10827 ( R152_U435 , R152_U269 , R152_U433 );
nand NAND2_10828 ( R152_U436 , U139 , R152_U69 );
nand NAND2_10829 ( R152_U437 , SI_25_ , R152_U70 );
nand NAND2_10830 ( R152_U438 , U139 , R152_U69 );
nand NAND2_10831 ( R152_U439 , SI_25_ , R152_U70 );
nand NAND2_10832 ( R152_U440 , R152_U439 , R152_U438 );
nand NAND2_10833 ( R152_U441 , R152_U158 , R152_U159 );
nand NAND2_10834 ( R152_U442 , R152_U265 , R152_U440 );
nand NAND2_10835 ( R152_U443 , U140 , R152_U67 );
nand NAND2_10836 ( R152_U444 , SI_24_ , R152_U68 );
nand NAND2_10837 ( R152_U445 , U140 , R152_U67 );
nand NAND2_10838 ( R152_U446 , SI_24_ , R152_U68 );
nand NAND2_10839 ( R152_U447 , R152_U446 , R152_U445 );
nand NAND2_10840 ( R152_U448 , R152_U160 , R152_U161 );
nand NAND2_10841 ( R152_U449 , R152_U261 , R152_U447 );
nand NAND2_10842 ( R152_U450 , U141 , R152_U65 );
nand NAND2_10843 ( R152_U451 , SI_23_ , R152_U66 );
nand NAND2_10844 ( R152_U452 , U141 , R152_U65 );
nand NAND2_10845 ( R152_U453 , SI_23_ , R152_U66 );
nand NAND2_10846 ( R152_U454 , R152_U453 , R152_U452 );
nand NAND2_10847 ( R152_U455 , R152_U162 , R152_U163 );
nand NAND2_10848 ( R152_U456 , R152_U257 , R152_U454 );
nand NAND2_10849 ( R152_U457 , U142 , R152_U63 );
nand NAND2_10850 ( R152_U458 , SI_22_ , R152_U64 );
nand NAND2_10851 ( R152_U459 , U142 , R152_U63 );
nand NAND2_10852 ( R152_U460 , SI_22_ , R152_U64 );
nand NAND2_10853 ( R152_U461 , R152_U460 , R152_U459 );
nand NAND2_10854 ( R152_U462 , R152_U164 , R152_U165 );
nand NAND2_10855 ( R152_U463 , R152_U253 , R152_U461 );
nand NAND2_10856 ( R152_U464 , U143 , R152_U61 );
nand NAND2_10857 ( R152_U465 , SI_21_ , R152_U62 );
nand NAND2_10858 ( R152_U466 , U143 , R152_U61 );
nand NAND2_10859 ( R152_U467 , SI_21_ , R152_U62 );
nand NAND2_10860 ( R152_U468 , R152_U467 , R152_U466 );
nand NAND2_10861 ( R152_U469 , R152_U166 , R152_U167 );
nand NAND2_10862 ( R152_U470 , R152_U249 , R152_U468 );
nand NAND2_10863 ( R152_U471 , U144 , R152_U59 );
nand NAND2_10864 ( R152_U472 , SI_20_ , R152_U60 );
nand NAND2_10865 ( R152_U473 , U144 , R152_U59 );
nand NAND2_10866 ( R152_U474 , SI_20_ , R152_U60 );
nand NAND2_10867 ( R152_U475 , R152_U474 , R152_U473 );
nand NAND2_10868 ( R152_U476 , R152_U168 , R152_U169 );
nand NAND2_10869 ( R152_U477 , R152_U245 , R152_U475 );
nand NAND2_10870 ( R152_U478 , U156 , R152_U170 );
nand NAND2_10871 ( R152_U479 , R152_U120 , R152_U26 );
nand NAND2_10872 ( R152_U480 , R152_U479 , R152_U478 );
nand NAND3_10873 ( R152_U481 , SI_1_ , R152_U170 , R152_U26 );
nand NAND2_10874 ( R152_U482 , R152_U194 , U156 );
nand NAND2_10875 ( R152_U483 , U146 , R152_U57 );
nand NAND2_10876 ( R152_U484 , SI_19_ , R152_U58 );
nand NAND2_10877 ( R152_U485 , U146 , R152_U57 );
nand NAND2_10878 ( R152_U486 , SI_19_ , R152_U58 );
nand NAND2_10879 ( R152_U487 , R152_U486 , R152_U485 );
nand NAND2_10880 ( R152_U488 , R152_U173 , R152_U174 );
nand NAND2_10881 ( R152_U489 , R152_U241 , R152_U487 );
nand NAND2_10882 ( R152_U490 , U147 , R152_U55 );
nand NAND2_10883 ( R152_U491 , SI_18_ , R152_U56 );
nand NAND2_10884 ( R152_U492 , U147 , R152_U55 );
nand NAND2_10885 ( R152_U493 , SI_18_ , R152_U56 );
nand NAND2_10886 ( R152_U494 , R152_U493 , R152_U492 );
nand NAND2_10887 ( R152_U495 , R152_U175 , R152_U176 );
nand NAND2_10888 ( R152_U496 , R152_U237 , R152_U494 );
nand NAND2_10889 ( R152_U497 , U148 , R152_U53 );
nand NAND2_10890 ( R152_U498 , SI_17_ , R152_U54 );
nand NAND2_10891 ( R152_U499 , U148 , R152_U53 );
nand NAND2_10892 ( R152_U500 , SI_17_ , R152_U54 );
nand NAND2_10893 ( R152_U501 , R152_U500 , R152_U499 );
nand NAND2_10894 ( R152_U502 , R152_U177 , R152_U178 );
nand NAND2_10895 ( R152_U503 , R152_U233 , R152_U501 );
nand NAND2_10896 ( R152_U504 , U149 , R152_U51 );
nand NAND2_10897 ( R152_U505 , SI_16_ , R152_U52 );
nand NAND2_10898 ( R152_U506 , U149 , R152_U51 );
nand NAND2_10899 ( R152_U507 , SI_16_ , R152_U52 );
nand NAND2_10900 ( R152_U508 , R152_U507 , R152_U506 );
nand NAND2_10901 ( R152_U509 , R152_U179 , R152_U180 );
nand NAND2_10902 ( R152_U510 , R152_U328 , R152_U508 );
nand NAND2_10903 ( R152_U511 , U150 , R152_U38 );
nand NAND2_10904 ( R152_U512 , SI_15_ , R152_U39 );
nand NAND2_10905 ( R152_U513 , U150 , R152_U38 );
nand NAND2_10906 ( R152_U514 , SI_15_ , R152_U39 );
nand NAND2_10907 ( R152_U515 , R152_U514 , R152_U513 );
nand NAND2_10908 ( R152_U516 , R152_U181 , R152_U182 );
nand NAND2_10909 ( R152_U517 , R152_U326 , R152_U515 );
nand NAND2_10910 ( R152_U518 , U151 , R152_U40 );
nand NAND2_10911 ( R152_U519 , SI_14_ , R152_U41 );
nand NAND2_10912 ( R152_U520 , U151 , R152_U40 );
nand NAND2_10913 ( R152_U521 , SI_14_ , R152_U41 );
nand NAND2_10914 ( R152_U522 , R152_U521 , R152_U520 );
nand NAND2_10915 ( R152_U523 , R152_U183 , R152_U184 );
nand NAND2_10916 ( R152_U524 , R152_U324 , R152_U522 );
nand NAND2_10917 ( R152_U525 , U152 , R152_U42 );
nand NAND2_10918 ( R152_U526 , SI_13_ , R152_U43 );
nand NAND2_10919 ( R152_U527 , U152 , R152_U42 );
nand NAND2_10920 ( R152_U528 , SI_13_ , R152_U43 );
nand NAND2_10921 ( R152_U529 , R152_U528 , R152_U527 );
nand NAND2_10922 ( R152_U530 , R152_U185 , R152_U186 );
nand NAND2_10923 ( R152_U531 , R152_U322 , R152_U529 );
nand NAND2_10924 ( R152_U532 , U153 , R152_U44 );
nand NAND2_10925 ( R152_U533 , SI_12_ , R152_U45 );
nand NAND2_10926 ( R152_U534 , U153 , R152_U44 );
nand NAND2_10927 ( R152_U535 , SI_12_ , R152_U45 );
nand NAND2_10928 ( R152_U536 , R152_U535 , R152_U534 );
nand NAND2_10929 ( R152_U537 , R152_U187 , R152_U188 );
nand NAND2_10930 ( R152_U538 , R152_U320 , R152_U536 );
nand NAND2_10931 ( R152_U539 , U154 , R152_U46 );
nand NAND2_10932 ( R152_U540 , SI_11_ , R152_U47 );
nand NAND2_10933 ( R152_U541 , U154 , R152_U46 );
nand NAND2_10934 ( R152_U542 , SI_11_ , R152_U47 );
nand NAND2_10935 ( R152_U543 , R152_U542 , R152_U541 );
nand NAND2_10936 ( R152_U544 , R152_U189 , R152_U190 );
nand NAND2_10937 ( R152_U545 , R152_U336 , R152_U543 );
nand NAND2_10938 ( R152_U546 , U155 , R152_U49 );
nand NAND2_10939 ( R152_U547 , SI_10_ , R152_U50 );
nand NAND2_10940 ( R152_U548 , U155 , R152_U49 );
nand NAND2_10941 ( R152_U549 , SI_10_ , R152_U50 );
nand NAND2_10942 ( R152_U550 , R152_U549 , R152_U548 );
nand NAND2_10943 ( R152_U551 , R152_U191 , R152_U192 );
nand NAND2_10944 ( R152_U552 , R152_U334 , R152_U550 );
nand NAND2_10945 ( R152_U553 , U157 , R152_U24 );
nand NAND2_10946 ( R152_U554 , SI_0_ , R152_U25 );
not NOT1_10947 ( LT_1602_U6 , P3_ADDR_REG_19_ );
not NOT1_10948 ( LT_1601_U6 , P1_ADDR_REG_19_ );
and AND2_10949 ( SUB_1596_U4 , SUB_1596_U159 , SUB_1596_U155 );
nand NAND3_10950 ( SUB_1596_U5 , SUB_1596_U221 , SUB_1596_U220 , SUB_1596_U160 );
not NOT1_10951 ( SUB_1596_U6 , ADD_1596_U7 );
not NOT1_10952 ( SUB_1596_U7 , P2_ADDR_REG_0_ );
not NOT1_10953 ( SUB_1596_U8 , P2_ADDR_REG_1_ );
nand NAND2_10954 ( SUB_1596_U9 , P2_ADDR_REG_0_ , ADD_1596_U7 );
not NOT1_10955 ( SUB_1596_U10 , ADD_1596_U55 );
not NOT1_10956 ( SUB_1596_U11 , ADD_1596_U54 );
not NOT1_10957 ( SUB_1596_U12 , P2_ADDR_REG_2_ );
nand NAND2_10958 ( SUB_1596_U13 , SUB_1596_U90 , SUB_1596_U89 );
not NOT1_10959 ( SUB_1596_U14 , ADD_1596_U53 );
not NOT1_10960 ( SUB_1596_U15 , P2_ADDR_REG_3_ );
not NOT1_10961 ( SUB_1596_U16 , ADD_1596_U52 );
not NOT1_10962 ( SUB_1596_U17 , P2_ADDR_REG_4_ );
nand NAND2_10963 ( SUB_1596_U18 , SUB_1596_U98 , SUB_1596_U97 );
not NOT1_10964 ( SUB_1596_U19 , ADD_1596_U51 );
not NOT1_10965 ( SUB_1596_U20 , P2_ADDR_REG_5_ );
not NOT1_10966 ( SUB_1596_U21 , ADD_1596_U50 );
not NOT1_10967 ( SUB_1596_U22 , P2_ADDR_REG_6_ );
not NOT1_10968 ( SUB_1596_U23 , ADD_1596_U49 );
not NOT1_10969 ( SUB_1596_U24 , P2_ADDR_REG_7_ );
nand NAND2_10970 ( SUB_1596_U25 , SUB_1596_U110 , SUB_1596_U109 );
not NOT1_10971 ( SUB_1596_U26 , ADD_1596_U48 );
not NOT1_10972 ( SUB_1596_U27 , P2_ADDR_REG_8_ );
not NOT1_10973 ( SUB_1596_U28 , P2_ADDR_REG_9_ );
not NOT1_10974 ( SUB_1596_U29 , ADD_1596_U47 );
nand NAND2_10975 ( SUB_1596_U30 , SUB_1596_U118 , SUB_1596_U117 );
not NOT1_10976 ( SUB_1596_U31 , ADD_1596_U64 );
not NOT1_10977 ( SUB_1596_U32 , P2_ADDR_REG_10_ );
not NOT1_10978 ( SUB_1596_U33 , ADD_1596_U63 );
not NOT1_10979 ( SUB_1596_U34 , P2_ADDR_REG_11_ );
not NOT1_10980 ( SUB_1596_U35 , ADD_1596_U62 );
not NOT1_10981 ( SUB_1596_U36 , P2_ADDR_REG_12_ );
nand NAND2_10982 ( SUB_1596_U37 , SUB_1596_U130 , SUB_1596_U129 );
not NOT1_10983 ( SUB_1596_U38 , ADD_1596_U61 );
not NOT1_10984 ( SUB_1596_U39 , P2_ADDR_REG_13_ );
nand NAND2_10985 ( SUB_1596_U40 , SUB_1596_U134 , SUB_1596_U133 );
not NOT1_10986 ( SUB_1596_U41 , ADD_1596_U60 );
not NOT1_10987 ( SUB_1596_U42 , P2_ADDR_REG_14_ );
nand NAND2_10988 ( SUB_1596_U43 , SUB_1596_U138 , SUB_1596_U137 );
not NOT1_10989 ( SUB_1596_U44 , ADD_1596_U59 );
not NOT1_10990 ( SUB_1596_U45 , P2_ADDR_REG_15_ );
not NOT1_10991 ( SUB_1596_U46 , ADD_1596_U58 );
not NOT1_10992 ( SUB_1596_U47 , P2_ADDR_REG_16_ );
not NOT1_10993 ( SUB_1596_U48 , ADD_1596_U57 );
not NOT1_10994 ( SUB_1596_U49 , P2_ADDR_REG_17_ );
nand NAND2_10995 ( SUB_1596_U50 , SUB_1596_U150 , SUB_1596_U149 );
not NOT1_10996 ( SUB_1596_U51 , ADD_1596_U56 );
not NOT1_10997 ( SUB_1596_U52 , P2_ADDR_REG_18_ );
nand NAND2_10998 ( SUB_1596_U53 , SUB_1596_U291 , SUB_1596_U290 );
nand NAND2_10999 ( SUB_1596_U54 , SUB_1596_U167 , SUB_1596_U166 );
nand NAND2_11000 ( SUB_1596_U55 , SUB_1596_U174 , SUB_1596_U173 );
nand NAND2_11001 ( SUB_1596_U56 , SUB_1596_U181 , SUB_1596_U180 );
nand NAND2_11002 ( SUB_1596_U57 , SUB_1596_U188 , SUB_1596_U187 );
nand NAND2_11003 ( SUB_1596_U58 , SUB_1596_U195 , SUB_1596_U194 );
nand NAND2_11004 ( SUB_1596_U59 , SUB_1596_U202 , SUB_1596_U201 );
nand NAND2_11005 ( SUB_1596_U60 , SUB_1596_U209 , SUB_1596_U208 );
nand NAND2_11006 ( SUB_1596_U61 , SUB_1596_U216 , SUB_1596_U215 );
nand NAND2_11007 ( SUB_1596_U62 , SUB_1596_U233 , SUB_1596_U232 );
nand NAND2_11008 ( SUB_1596_U63 , SUB_1596_U240 , SUB_1596_U239 );
nand NAND2_11009 ( SUB_1596_U64 , SUB_1596_U247 , SUB_1596_U246 );
nand NAND2_11010 ( SUB_1596_U65 , SUB_1596_U254 , SUB_1596_U253 );
nand NAND2_11011 ( SUB_1596_U66 , SUB_1596_U261 , SUB_1596_U260 );
nand NAND2_11012 ( SUB_1596_U67 , SUB_1596_U268 , SUB_1596_U267 );
nand NAND2_11013 ( SUB_1596_U68 , SUB_1596_U275 , SUB_1596_U274 );
nand NAND2_11014 ( SUB_1596_U69 , SUB_1596_U282 , SUB_1596_U281 );
nand NAND2_11015 ( SUB_1596_U70 , SUB_1596_U289 , SUB_1596_U288 );
nand NAND2_11016 ( SUB_1596_U71 , SUB_1596_U114 , SUB_1596_U113 );
nand NAND2_11017 ( SUB_1596_U72 , SUB_1596_U106 , SUB_1596_U105 );
nand NAND2_11018 ( SUB_1596_U73 , SUB_1596_U102 , SUB_1596_U101 );
nand NAND2_11019 ( SUB_1596_U74 , SUB_1596_U94 , SUB_1596_U93 );
nand NAND2_11020 ( SUB_1596_U75 , SUB_1596_U76 , SUB_1596_U86 );
nand NAND2_11021 ( SUB_1596_U76 , ADD_1596_U55 , SUB_1596_U84 );
not NOT1_11022 ( SUB_1596_U77 , P2_ADDR_REG_19_ );
not NOT1_11023 ( SUB_1596_U78 , ADD_1596_U6 );
nand NAND2_11024 ( SUB_1596_U79 , SUB_1596_U146 , SUB_1596_U145 );
nand NAND2_11025 ( SUB_1596_U80 , SUB_1596_U142 , SUB_1596_U141 );
nand NAND2_11026 ( SUB_1596_U81 , SUB_1596_U126 , SUB_1596_U125 );
nand NAND2_11027 ( SUB_1596_U82 , SUB_1596_U122 , SUB_1596_U121 );
not NOT1_11028 ( SUB_1596_U83 , SUB_1596_U76 );
not NOT1_11029 ( SUB_1596_U84 , SUB_1596_U9 );
nand NAND2_11030 ( SUB_1596_U85 , SUB_1596_U10 , SUB_1596_U9 );
nand NAND2_11031 ( SUB_1596_U86 , P2_ADDR_REG_1_ , SUB_1596_U85 );
not NOT1_11032 ( SUB_1596_U87 , SUB_1596_U75 );
or OR2_11033 ( SUB_1596_U88 , ADD_1596_U54 , P2_ADDR_REG_2_ );
nand NAND2_11034 ( SUB_1596_U89 , SUB_1596_U88 , SUB_1596_U75 );
nand NAND2_11035 ( SUB_1596_U90 , P2_ADDR_REG_2_ , ADD_1596_U54 );
not NOT1_11036 ( SUB_1596_U91 , SUB_1596_U13 );
nand NAND2_11037 ( SUB_1596_U92 , SUB_1596_U91 , SUB_1596_U15 );
nand NAND2_11038 ( SUB_1596_U93 , ADD_1596_U53 , SUB_1596_U92 );
nand NAND2_11039 ( SUB_1596_U94 , P2_ADDR_REG_3_ , SUB_1596_U13 );
not NOT1_11040 ( SUB_1596_U95 , SUB_1596_U74 );
or OR2_11041 ( SUB_1596_U96 , ADD_1596_U52 , P2_ADDR_REG_4_ );
nand NAND2_11042 ( SUB_1596_U97 , SUB_1596_U96 , SUB_1596_U74 );
nand NAND2_11043 ( SUB_1596_U98 , P2_ADDR_REG_4_ , ADD_1596_U52 );
not NOT1_11044 ( SUB_1596_U99 , SUB_1596_U18 );
nand NAND2_11045 ( SUB_1596_U100 , SUB_1596_U99 , SUB_1596_U20 );
nand NAND2_11046 ( SUB_1596_U101 , ADD_1596_U51 , SUB_1596_U100 );
nand NAND2_11047 ( SUB_1596_U102 , P2_ADDR_REG_5_ , SUB_1596_U18 );
not NOT1_11048 ( SUB_1596_U103 , SUB_1596_U73 );
or OR2_11049 ( SUB_1596_U104 , ADD_1596_U50 , P2_ADDR_REG_6_ );
nand NAND2_11050 ( SUB_1596_U105 , SUB_1596_U104 , SUB_1596_U73 );
nand NAND2_11051 ( SUB_1596_U106 , P2_ADDR_REG_6_ , ADD_1596_U50 );
not NOT1_11052 ( SUB_1596_U107 , SUB_1596_U72 );
or OR2_11053 ( SUB_1596_U108 , ADD_1596_U49 , P2_ADDR_REG_7_ );
nand NAND2_11054 ( SUB_1596_U109 , SUB_1596_U108 , SUB_1596_U72 );
nand NAND2_11055 ( SUB_1596_U110 , P2_ADDR_REG_7_ , ADD_1596_U49 );
not NOT1_11056 ( SUB_1596_U111 , SUB_1596_U25 );
nand NAND2_11057 ( SUB_1596_U112 , SUB_1596_U111 , SUB_1596_U27 );
nand NAND2_11058 ( SUB_1596_U113 , ADD_1596_U48 , SUB_1596_U112 );
nand NAND2_11059 ( SUB_1596_U114 , P2_ADDR_REG_8_ , SUB_1596_U25 );
not NOT1_11060 ( SUB_1596_U115 , SUB_1596_U71 );
or OR2_11061 ( SUB_1596_U116 , ADD_1596_U47 , P2_ADDR_REG_9_ );
nand NAND2_11062 ( SUB_1596_U117 , SUB_1596_U116 , SUB_1596_U71 );
nand NAND2_11063 ( SUB_1596_U118 , ADD_1596_U47 , P2_ADDR_REG_9_ );
not NOT1_11064 ( SUB_1596_U119 , SUB_1596_U30 );
nand NAND2_11065 ( SUB_1596_U120 , SUB_1596_U119 , SUB_1596_U32 );
nand NAND2_11066 ( SUB_1596_U121 , ADD_1596_U64 , SUB_1596_U120 );
nand NAND2_11067 ( SUB_1596_U122 , P2_ADDR_REG_10_ , SUB_1596_U30 );
not NOT1_11068 ( SUB_1596_U123 , SUB_1596_U82 );
or OR2_11069 ( SUB_1596_U124 , ADD_1596_U63 , P2_ADDR_REG_11_ );
nand NAND2_11070 ( SUB_1596_U125 , SUB_1596_U124 , SUB_1596_U82 );
nand NAND2_11071 ( SUB_1596_U126 , P2_ADDR_REG_11_ , ADD_1596_U63 );
not NOT1_11072 ( SUB_1596_U127 , SUB_1596_U81 );
or OR2_11073 ( SUB_1596_U128 , ADD_1596_U62 , P2_ADDR_REG_12_ );
nand NAND2_11074 ( SUB_1596_U129 , SUB_1596_U128 , SUB_1596_U81 );
nand NAND2_11075 ( SUB_1596_U130 , P2_ADDR_REG_12_ , ADD_1596_U62 );
not NOT1_11076 ( SUB_1596_U131 , SUB_1596_U37 );
nand NAND2_11077 ( SUB_1596_U132 , SUB_1596_U131 , SUB_1596_U39 );
nand NAND2_11078 ( SUB_1596_U133 , ADD_1596_U61 , SUB_1596_U132 );
nand NAND2_11079 ( SUB_1596_U134 , P2_ADDR_REG_13_ , SUB_1596_U37 );
not NOT1_11080 ( SUB_1596_U135 , SUB_1596_U40 );
nand NAND2_11081 ( SUB_1596_U136 , SUB_1596_U135 , SUB_1596_U42 );
nand NAND2_11082 ( SUB_1596_U137 , ADD_1596_U60 , SUB_1596_U136 );
nand NAND2_11083 ( SUB_1596_U138 , P2_ADDR_REG_14_ , SUB_1596_U40 );
not NOT1_11084 ( SUB_1596_U139 , SUB_1596_U43 );
nand NAND2_11085 ( SUB_1596_U140 , SUB_1596_U139 , SUB_1596_U45 );
nand NAND2_11086 ( SUB_1596_U141 , ADD_1596_U59 , SUB_1596_U140 );
nand NAND2_11087 ( SUB_1596_U142 , P2_ADDR_REG_15_ , SUB_1596_U43 );
not NOT1_11088 ( SUB_1596_U143 , SUB_1596_U80 );
or OR2_11089 ( SUB_1596_U144 , ADD_1596_U58 , P2_ADDR_REG_16_ );
nand NAND2_11090 ( SUB_1596_U145 , SUB_1596_U144 , SUB_1596_U80 );
nand NAND2_11091 ( SUB_1596_U146 , P2_ADDR_REG_16_ , ADD_1596_U58 );
not NOT1_11092 ( SUB_1596_U147 , SUB_1596_U79 );
or OR2_11093 ( SUB_1596_U148 , ADD_1596_U57 , P2_ADDR_REG_17_ );
nand NAND2_11094 ( SUB_1596_U149 , SUB_1596_U148 , SUB_1596_U79 );
nand NAND2_11095 ( SUB_1596_U150 , P2_ADDR_REG_17_ , ADD_1596_U57 );
not NOT1_11096 ( SUB_1596_U151 , SUB_1596_U50 );
nand NAND2_11097 ( SUB_1596_U152 , SUB_1596_U151 , SUB_1596_U52 );
nand NAND2_11098 ( SUB_1596_U153 , ADD_1596_U56 , SUB_1596_U152 );
nand NAND2_11099 ( SUB_1596_U154 , P2_ADDR_REG_18_ , SUB_1596_U50 );
nand NAND4_11100 ( SUB_1596_U155 , SUB_1596_U154 , SUB_1596_U153 , SUB_1596_U223 , SUB_1596_U222 );
nand NAND2_11101 ( SUB_1596_U156 , P2_ADDR_REG_18_ , SUB_1596_U50 );
nand NAND2_11102 ( SUB_1596_U157 , SUB_1596_U156 , SUB_1596_U51 );
nand NAND2_11103 ( SUB_1596_U158 , SUB_1596_U151 , SUB_1596_U52 );
nand NAND3_11104 ( SUB_1596_U159 , SUB_1596_U158 , SUB_1596_U157 , SUB_1596_U226 );
nand NAND2_11105 ( SUB_1596_U160 , SUB_1596_U219 , SUB_1596_U10 );
nand NAND2_11106 ( SUB_1596_U161 , P2_ADDR_REG_9_ , SUB_1596_U29 );
nand NAND2_11107 ( SUB_1596_U162 , ADD_1596_U47 , SUB_1596_U28 );
nand NAND2_11108 ( SUB_1596_U163 , P2_ADDR_REG_9_ , SUB_1596_U29 );
nand NAND2_11109 ( SUB_1596_U164 , ADD_1596_U47 , SUB_1596_U28 );
nand NAND2_11110 ( SUB_1596_U165 , SUB_1596_U164 , SUB_1596_U163 );
nand NAND3_11111 ( SUB_1596_U166 , SUB_1596_U162 , SUB_1596_U161 , SUB_1596_U71 );
nand NAND2_11112 ( SUB_1596_U167 , SUB_1596_U115 , SUB_1596_U165 );
nand NAND2_11113 ( SUB_1596_U168 , P2_ADDR_REG_8_ , SUB_1596_U25 );
nand NAND2_11114 ( SUB_1596_U169 , SUB_1596_U111 , SUB_1596_U27 );
nand NAND2_11115 ( SUB_1596_U170 , P2_ADDR_REG_8_ , SUB_1596_U25 );
nand NAND2_11116 ( SUB_1596_U171 , SUB_1596_U111 , SUB_1596_U27 );
nand NAND2_11117 ( SUB_1596_U172 , SUB_1596_U171 , SUB_1596_U170 );
nand NAND3_11118 ( SUB_1596_U173 , SUB_1596_U169 , SUB_1596_U168 , SUB_1596_U26 );
nand NAND2_11119 ( SUB_1596_U174 , SUB_1596_U172 , ADD_1596_U48 );
nand NAND2_11120 ( SUB_1596_U175 , P2_ADDR_REG_7_ , SUB_1596_U23 );
nand NAND2_11121 ( SUB_1596_U176 , ADD_1596_U49 , SUB_1596_U24 );
nand NAND2_11122 ( SUB_1596_U177 , P2_ADDR_REG_7_ , SUB_1596_U23 );
nand NAND2_11123 ( SUB_1596_U178 , ADD_1596_U49 , SUB_1596_U24 );
nand NAND2_11124 ( SUB_1596_U179 , SUB_1596_U178 , SUB_1596_U177 );
nand NAND3_11125 ( SUB_1596_U180 , SUB_1596_U176 , SUB_1596_U175 , SUB_1596_U72 );
nand NAND2_11126 ( SUB_1596_U181 , SUB_1596_U107 , SUB_1596_U179 );
nand NAND2_11127 ( SUB_1596_U182 , P2_ADDR_REG_6_ , SUB_1596_U21 );
nand NAND2_11128 ( SUB_1596_U183 , ADD_1596_U50 , SUB_1596_U22 );
nand NAND2_11129 ( SUB_1596_U184 , P2_ADDR_REG_6_ , SUB_1596_U21 );
nand NAND2_11130 ( SUB_1596_U185 , ADD_1596_U50 , SUB_1596_U22 );
nand NAND2_11131 ( SUB_1596_U186 , SUB_1596_U185 , SUB_1596_U184 );
nand NAND3_11132 ( SUB_1596_U187 , SUB_1596_U183 , SUB_1596_U182 , SUB_1596_U73 );
nand NAND2_11133 ( SUB_1596_U188 , SUB_1596_U103 , SUB_1596_U186 );
nand NAND2_11134 ( SUB_1596_U189 , P2_ADDR_REG_5_ , SUB_1596_U18 );
nand NAND2_11135 ( SUB_1596_U190 , SUB_1596_U99 , SUB_1596_U20 );
nand NAND2_11136 ( SUB_1596_U191 , P2_ADDR_REG_5_ , SUB_1596_U18 );
nand NAND2_11137 ( SUB_1596_U192 , SUB_1596_U99 , SUB_1596_U20 );
nand NAND2_11138 ( SUB_1596_U193 , SUB_1596_U192 , SUB_1596_U191 );
nand NAND3_11139 ( SUB_1596_U194 , SUB_1596_U190 , SUB_1596_U189 , SUB_1596_U19 );
nand NAND2_11140 ( SUB_1596_U195 , SUB_1596_U193 , ADD_1596_U51 );
nand NAND2_11141 ( SUB_1596_U196 , P2_ADDR_REG_4_ , SUB_1596_U16 );
nand NAND2_11142 ( SUB_1596_U197 , ADD_1596_U52 , SUB_1596_U17 );
nand NAND2_11143 ( SUB_1596_U198 , P2_ADDR_REG_4_ , SUB_1596_U16 );
nand NAND2_11144 ( SUB_1596_U199 , ADD_1596_U52 , SUB_1596_U17 );
nand NAND2_11145 ( SUB_1596_U200 , SUB_1596_U199 , SUB_1596_U198 );
nand NAND3_11146 ( SUB_1596_U201 , SUB_1596_U197 , SUB_1596_U196 , SUB_1596_U74 );
nand NAND2_11147 ( SUB_1596_U202 , SUB_1596_U95 , SUB_1596_U200 );
nand NAND2_11148 ( SUB_1596_U203 , P2_ADDR_REG_3_ , SUB_1596_U13 );
nand NAND2_11149 ( SUB_1596_U204 , SUB_1596_U91 , SUB_1596_U15 );
nand NAND2_11150 ( SUB_1596_U205 , P2_ADDR_REG_3_ , SUB_1596_U13 );
nand NAND2_11151 ( SUB_1596_U206 , SUB_1596_U91 , SUB_1596_U15 );
nand NAND2_11152 ( SUB_1596_U207 , SUB_1596_U206 , SUB_1596_U205 );
nand NAND3_11153 ( SUB_1596_U208 , SUB_1596_U204 , SUB_1596_U203 , SUB_1596_U14 );
nand NAND2_11154 ( SUB_1596_U209 , SUB_1596_U207 , ADD_1596_U53 );
nand NAND2_11155 ( SUB_1596_U210 , P2_ADDR_REG_2_ , SUB_1596_U11 );
nand NAND2_11156 ( SUB_1596_U211 , ADD_1596_U54 , SUB_1596_U12 );
nand NAND2_11157 ( SUB_1596_U212 , P2_ADDR_REG_2_ , SUB_1596_U11 );
nand NAND2_11158 ( SUB_1596_U213 , ADD_1596_U54 , SUB_1596_U12 );
nand NAND2_11159 ( SUB_1596_U214 , SUB_1596_U213 , SUB_1596_U212 );
nand NAND3_11160 ( SUB_1596_U215 , SUB_1596_U211 , SUB_1596_U210 , SUB_1596_U75 );
nand NAND2_11161 ( SUB_1596_U216 , SUB_1596_U87 , SUB_1596_U214 );
nand NAND2_11162 ( SUB_1596_U217 , P2_ADDR_REG_1_ , SUB_1596_U9 );
nand NAND2_11163 ( SUB_1596_U218 , SUB_1596_U84 , SUB_1596_U8 );
nand NAND2_11164 ( SUB_1596_U219 , SUB_1596_U218 , SUB_1596_U217 );
nand NAND3_11165 ( SUB_1596_U220 , ADD_1596_U55 , SUB_1596_U9 , SUB_1596_U8 );
nand NAND2_11166 ( SUB_1596_U221 , SUB_1596_U83 , P2_ADDR_REG_1_ );
nand NAND2_11167 ( SUB_1596_U222 , P2_ADDR_REG_19_ , SUB_1596_U78 );
nand NAND2_11168 ( SUB_1596_U223 , ADD_1596_U6 , SUB_1596_U77 );
nand NAND2_11169 ( SUB_1596_U224 , P2_ADDR_REG_19_ , SUB_1596_U78 );
nand NAND2_11170 ( SUB_1596_U225 , ADD_1596_U6 , SUB_1596_U77 );
nand NAND2_11171 ( SUB_1596_U226 , SUB_1596_U225 , SUB_1596_U224 );
nand NAND2_11172 ( SUB_1596_U227 , P2_ADDR_REG_18_ , SUB_1596_U50 );
nand NAND2_11173 ( SUB_1596_U228 , SUB_1596_U151 , SUB_1596_U52 );
nand NAND2_11174 ( SUB_1596_U229 , P2_ADDR_REG_18_ , SUB_1596_U50 );
nand NAND2_11175 ( SUB_1596_U230 , SUB_1596_U151 , SUB_1596_U52 );
nand NAND2_11176 ( SUB_1596_U231 , SUB_1596_U230 , SUB_1596_U229 );
nand NAND3_11177 ( SUB_1596_U232 , SUB_1596_U228 , SUB_1596_U227 , SUB_1596_U51 );
nand NAND2_11178 ( SUB_1596_U233 , SUB_1596_U231 , ADD_1596_U56 );
nand NAND2_11179 ( SUB_1596_U234 , P2_ADDR_REG_17_ , SUB_1596_U48 );
nand NAND2_11180 ( SUB_1596_U235 , ADD_1596_U57 , SUB_1596_U49 );
nand NAND2_11181 ( SUB_1596_U236 , P2_ADDR_REG_17_ , SUB_1596_U48 );
nand NAND2_11182 ( SUB_1596_U237 , ADD_1596_U57 , SUB_1596_U49 );
nand NAND2_11183 ( SUB_1596_U238 , SUB_1596_U237 , SUB_1596_U236 );
nand NAND3_11184 ( SUB_1596_U239 , SUB_1596_U235 , SUB_1596_U234 , SUB_1596_U79 );
nand NAND2_11185 ( SUB_1596_U240 , SUB_1596_U147 , SUB_1596_U238 );
nand NAND2_11186 ( SUB_1596_U241 , P2_ADDR_REG_16_ , SUB_1596_U46 );
nand NAND2_11187 ( SUB_1596_U242 , ADD_1596_U58 , SUB_1596_U47 );
nand NAND2_11188 ( SUB_1596_U243 , P2_ADDR_REG_16_ , SUB_1596_U46 );
nand NAND2_11189 ( SUB_1596_U244 , ADD_1596_U58 , SUB_1596_U47 );
nand NAND2_11190 ( SUB_1596_U245 , SUB_1596_U244 , SUB_1596_U243 );
nand NAND3_11191 ( SUB_1596_U246 , SUB_1596_U242 , SUB_1596_U241 , SUB_1596_U80 );
nand NAND2_11192 ( SUB_1596_U247 , SUB_1596_U143 , SUB_1596_U245 );
nand NAND2_11193 ( SUB_1596_U248 , P2_ADDR_REG_15_ , SUB_1596_U43 );
nand NAND2_11194 ( SUB_1596_U249 , SUB_1596_U139 , SUB_1596_U45 );
nand NAND2_11195 ( SUB_1596_U250 , P2_ADDR_REG_15_ , SUB_1596_U43 );
nand NAND2_11196 ( SUB_1596_U251 , SUB_1596_U139 , SUB_1596_U45 );
nand NAND2_11197 ( SUB_1596_U252 , SUB_1596_U251 , SUB_1596_U250 );
nand NAND3_11198 ( SUB_1596_U253 , SUB_1596_U249 , SUB_1596_U248 , SUB_1596_U44 );
nand NAND2_11199 ( SUB_1596_U254 , SUB_1596_U252 , ADD_1596_U59 );
nand NAND2_11200 ( SUB_1596_U255 , P2_ADDR_REG_14_ , SUB_1596_U40 );
nand NAND2_11201 ( SUB_1596_U256 , SUB_1596_U135 , SUB_1596_U42 );
nand NAND2_11202 ( SUB_1596_U257 , P2_ADDR_REG_14_ , SUB_1596_U40 );
nand NAND2_11203 ( SUB_1596_U258 , SUB_1596_U135 , SUB_1596_U42 );
nand NAND2_11204 ( SUB_1596_U259 , SUB_1596_U258 , SUB_1596_U257 );
nand NAND3_11205 ( SUB_1596_U260 , SUB_1596_U256 , SUB_1596_U255 , SUB_1596_U41 );
nand NAND2_11206 ( SUB_1596_U261 , SUB_1596_U259 , ADD_1596_U60 );
nand NAND2_11207 ( SUB_1596_U262 , P2_ADDR_REG_13_ , SUB_1596_U37 );
nand NAND2_11208 ( SUB_1596_U263 , SUB_1596_U131 , SUB_1596_U39 );
nand NAND2_11209 ( SUB_1596_U264 , P2_ADDR_REG_13_ , SUB_1596_U37 );
nand NAND2_11210 ( SUB_1596_U265 , SUB_1596_U131 , SUB_1596_U39 );
nand NAND2_11211 ( SUB_1596_U266 , SUB_1596_U265 , SUB_1596_U264 );
nand NAND3_11212 ( SUB_1596_U267 , SUB_1596_U263 , SUB_1596_U262 , SUB_1596_U38 );
nand NAND2_11213 ( SUB_1596_U268 , SUB_1596_U266 , ADD_1596_U61 );
nand NAND2_11214 ( SUB_1596_U269 , P2_ADDR_REG_12_ , SUB_1596_U35 );
nand NAND2_11215 ( SUB_1596_U270 , ADD_1596_U62 , SUB_1596_U36 );
nand NAND2_11216 ( SUB_1596_U271 , P2_ADDR_REG_12_ , SUB_1596_U35 );
nand NAND2_11217 ( SUB_1596_U272 , ADD_1596_U62 , SUB_1596_U36 );
nand NAND2_11218 ( SUB_1596_U273 , SUB_1596_U272 , SUB_1596_U271 );
nand NAND3_11219 ( SUB_1596_U274 , SUB_1596_U270 , SUB_1596_U269 , SUB_1596_U81 );
nand NAND2_11220 ( SUB_1596_U275 , SUB_1596_U127 , SUB_1596_U273 );
nand NAND2_11221 ( SUB_1596_U276 , P2_ADDR_REG_11_ , SUB_1596_U33 );
nand NAND2_11222 ( SUB_1596_U277 , ADD_1596_U63 , SUB_1596_U34 );
nand NAND2_11223 ( SUB_1596_U278 , P2_ADDR_REG_11_ , SUB_1596_U33 );
nand NAND2_11224 ( SUB_1596_U279 , ADD_1596_U63 , SUB_1596_U34 );
nand NAND2_11225 ( SUB_1596_U280 , SUB_1596_U279 , SUB_1596_U278 );
nand NAND3_11226 ( SUB_1596_U281 , SUB_1596_U277 , SUB_1596_U276 , SUB_1596_U82 );
nand NAND2_11227 ( SUB_1596_U282 , SUB_1596_U123 , SUB_1596_U280 );
nand NAND2_11228 ( SUB_1596_U283 , P2_ADDR_REG_10_ , SUB_1596_U30 );
nand NAND2_11229 ( SUB_1596_U284 , SUB_1596_U119 , SUB_1596_U32 );
nand NAND2_11230 ( SUB_1596_U285 , P2_ADDR_REG_10_ , SUB_1596_U30 );
nand NAND2_11231 ( SUB_1596_U286 , SUB_1596_U119 , SUB_1596_U32 );
nand NAND2_11232 ( SUB_1596_U287 , SUB_1596_U286 , SUB_1596_U285 );
nand NAND3_11233 ( SUB_1596_U288 , SUB_1596_U284 , SUB_1596_U283 , SUB_1596_U31 );
nand NAND2_11234 ( SUB_1596_U289 , SUB_1596_U287 , ADD_1596_U64 );
nand NAND2_11235 ( SUB_1596_U290 , P2_ADDR_REG_0_ , SUB_1596_U6 );
nand NAND2_11236 ( SUB_1596_U291 , ADD_1596_U7 , SUB_1596_U7 );
nand NAND2_11237 ( ADD_1596_U6 , ADD_1596_U174 , ADD_1596_U178 );
nand NAND2_11238 ( ADD_1596_U7 , ADD_1596_U9 , ADD_1596_U179 );
not NOT1_11239 ( ADD_1596_U8 , P3_ADDR_REG_0_ );
nand NAND2_11240 ( ADD_1596_U9 , P3_ADDR_REG_0_ , ADD_1596_U46 );
not NOT1_11241 ( ADD_1596_U10 , P1_ADDR_REG_1_ );
not NOT1_11242 ( ADD_1596_U11 , P3_ADDR_REG_2_ );
not NOT1_11243 ( ADD_1596_U12 , P1_ADDR_REG_2_ );
not NOT1_11244 ( ADD_1596_U13 , P3_ADDR_REG_3_ );
not NOT1_11245 ( ADD_1596_U14 , P1_ADDR_REG_3_ );
not NOT1_11246 ( ADD_1596_U15 , P3_ADDR_REG_4_ );
not NOT1_11247 ( ADD_1596_U16 , P1_ADDR_REG_4_ );
not NOT1_11248 ( ADD_1596_U17 , P3_ADDR_REG_5_ );
not NOT1_11249 ( ADD_1596_U18 , P1_ADDR_REG_5_ );
not NOT1_11250 ( ADD_1596_U19 , P3_ADDR_REG_6_ );
not NOT1_11251 ( ADD_1596_U20 , P1_ADDR_REG_6_ );
not NOT1_11252 ( ADD_1596_U21 , P3_ADDR_REG_7_ );
not NOT1_11253 ( ADD_1596_U22 , P1_ADDR_REG_7_ );
not NOT1_11254 ( ADD_1596_U23 , P3_ADDR_REG_8_ );
not NOT1_11255 ( ADD_1596_U24 , P1_ADDR_REG_8_ );
not NOT1_11256 ( ADD_1596_U25 , P3_ADDR_REG_9_ );
not NOT1_11257 ( ADD_1596_U26 , P1_ADDR_REG_9_ );
not NOT1_11258 ( ADD_1596_U27 , P3_ADDR_REG_10_ );
not NOT1_11259 ( ADD_1596_U28 , P1_ADDR_REG_10_ );
not NOT1_11260 ( ADD_1596_U29 , P3_ADDR_REG_11_ );
not NOT1_11261 ( ADD_1596_U30 , P1_ADDR_REG_11_ );
not NOT1_11262 ( ADD_1596_U31 , P3_ADDR_REG_12_ );
not NOT1_11263 ( ADD_1596_U32 , P1_ADDR_REG_12_ );
not NOT1_11264 ( ADD_1596_U33 , P3_ADDR_REG_13_ );
not NOT1_11265 ( ADD_1596_U34 , P1_ADDR_REG_13_ );
not NOT1_11266 ( ADD_1596_U35 , P3_ADDR_REG_14_ );
not NOT1_11267 ( ADD_1596_U36 , P1_ADDR_REG_14_ );
not NOT1_11268 ( ADD_1596_U37 , P3_ADDR_REG_15_ );
not NOT1_11269 ( ADD_1596_U38 , P1_ADDR_REG_15_ );
not NOT1_11270 ( ADD_1596_U39 , P3_ADDR_REG_16_ );
not NOT1_11271 ( ADD_1596_U40 , P1_ADDR_REG_16_ );
not NOT1_11272 ( ADD_1596_U41 , P3_ADDR_REG_17_ );
not NOT1_11273 ( ADD_1596_U42 , P1_ADDR_REG_17_ );
not NOT1_11274 ( ADD_1596_U43 , P3_ADDR_REG_18_ );
not NOT1_11275 ( ADD_1596_U44 , P1_ADDR_REG_18_ );
nand NAND2_11276 ( ADD_1596_U45 , ADD_1596_U169 , ADD_1596_U168 );
not NOT1_11277 ( ADD_1596_U46 , P1_ADDR_REG_0_ );
nand NAND2_11278 ( ADD_1596_U47 , ADD_1596_U184 , ADD_1596_U183 );
nand NAND2_11279 ( ADD_1596_U48 , ADD_1596_U189 , ADD_1596_U188 );
nand NAND2_11280 ( ADD_1596_U49 , ADD_1596_U194 , ADD_1596_U193 );
nand NAND2_11281 ( ADD_1596_U50 , ADD_1596_U199 , ADD_1596_U198 );
nand NAND2_11282 ( ADD_1596_U51 , ADD_1596_U204 , ADD_1596_U203 );
nand NAND2_11283 ( ADD_1596_U52 , ADD_1596_U209 , ADD_1596_U208 );
nand NAND2_11284 ( ADD_1596_U53 , ADD_1596_U214 , ADD_1596_U213 );
nand NAND2_11285 ( ADD_1596_U54 , ADD_1596_U219 , ADD_1596_U218 );
nand NAND2_11286 ( ADD_1596_U55 , ADD_1596_U224 , ADD_1596_U223 );
nand NAND2_11287 ( ADD_1596_U56 , ADD_1596_U234 , ADD_1596_U233 );
nand NAND2_11288 ( ADD_1596_U57 , ADD_1596_U239 , ADD_1596_U238 );
nand NAND2_11289 ( ADD_1596_U58 , ADD_1596_U244 , ADD_1596_U243 );
nand NAND2_11290 ( ADD_1596_U59 , ADD_1596_U249 , ADD_1596_U248 );
nand NAND2_11291 ( ADD_1596_U60 , ADD_1596_U254 , ADD_1596_U253 );
nand NAND2_11292 ( ADD_1596_U61 , ADD_1596_U259 , ADD_1596_U258 );
nand NAND2_11293 ( ADD_1596_U62 , ADD_1596_U264 , ADD_1596_U263 );
nand NAND2_11294 ( ADD_1596_U63 , ADD_1596_U269 , ADD_1596_U268 );
nand NAND2_11295 ( ADD_1596_U64 , ADD_1596_U274 , ADD_1596_U273 );
nand NAND2_11296 ( ADD_1596_U65 , ADD_1596_U181 , ADD_1596_U180 );
nand NAND2_11297 ( ADD_1596_U66 , ADD_1596_U186 , ADD_1596_U185 );
nand NAND2_11298 ( ADD_1596_U67 , ADD_1596_U191 , ADD_1596_U190 );
nand NAND2_11299 ( ADD_1596_U68 , ADD_1596_U196 , ADD_1596_U195 );
nand NAND2_11300 ( ADD_1596_U69 , ADD_1596_U201 , ADD_1596_U200 );
nand NAND2_11301 ( ADD_1596_U70 , ADD_1596_U206 , ADD_1596_U205 );
nand NAND2_11302 ( ADD_1596_U71 , ADD_1596_U211 , ADD_1596_U210 );
nand NAND2_11303 ( ADD_1596_U72 , ADD_1596_U216 , ADD_1596_U215 );
nand NAND2_11304 ( ADD_1596_U73 , ADD_1596_U221 , ADD_1596_U220 );
nand NAND2_11305 ( ADD_1596_U74 , ADD_1596_U231 , ADD_1596_U230 );
nand NAND2_11306 ( ADD_1596_U75 , ADD_1596_U236 , ADD_1596_U235 );
nand NAND2_11307 ( ADD_1596_U76 , ADD_1596_U241 , ADD_1596_U240 );
nand NAND2_11308 ( ADD_1596_U77 , ADD_1596_U246 , ADD_1596_U245 );
nand NAND2_11309 ( ADD_1596_U78 , ADD_1596_U251 , ADD_1596_U250 );
nand NAND2_11310 ( ADD_1596_U79 , ADD_1596_U256 , ADD_1596_U255 );
nand NAND2_11311 ( ADD_1596_U80 , ADD_1596_U261 , ADD_1596_U260 );
nand NAND2_11312 ( ADD_1596_U81 , ADD_1596_U266 , ADD_1596_U265 );
nand NAND2_11313 ( ADD_1596_U82 , ADD_1596_U271 , ADD_1596_U270 );
nand NAND2_11314 ( ADD_1596_U83 , ADD_1596_U133 , ADD_1596_U132 );
nand NAND2_11315 ( ADD_1596_U84 , ADD_1596_U129 , ADD_1596_U128 );
nand NAND2_11316 ( ADD_1596_U85 , ADD_1596_U125 , ADD_1596_U124 );
nand NAND2_11317 ( ADD_1596_U86 , ADD_1596_U121 , ADD_1596_U120 );
nand NAND2_11318 ( ADD_1596_U87 , ADD_1596_U117 , ADD_1596_U116 );
nand NAND2_11319 ( ADD_1596_U88 , ADD_1596_U113 , ADD_1596_U112 );
nand NAND2_11320 ( ADD_1596_U89 , ADD_1596_U109 , ADD_1596_U108 );
nand NAND2_11321 ( ADD_1596_U90 , ADD_1596_U105 , ADD_1596_U104 );
not NOT1_11322 ( ADD_1596_U91 , P3_ADDR_REG_1_ );
not NOT1_11323 ( ADD_1596_U92 , P3_ADDR_REG_19_ );
not NOT1_11324 ( ADD_1596_U93 , P1_ADDR_REG_19_ );
nand NAND2_11325 ( ADD_1596_U94 , ADD_1596_U165 , ADD_1596_U164 );
nand NAND2_11326 ( ADD_1596_U95 , ADD_1596_U161 , ADD_1596_U160 );
nand NAND2_11327 ( ADD_1596_U96 , ADD_1596_U157 , ADD_1596_U156 );
nand NAND2_11328 ( ADD_1596_U97 , ADD_1596_U153 , ADD_1596_U152 );
nand NAND2_11329 ( ADD_1596_U98 , ADD_1596_U149 , ADD_1596_U148 );
nand NAND2_11330 ( ADD_1596_U99 , ADD_1596_U145 , ADD_1596_U144 );
nand NAND2_11331 ( ADD_1596_U100 , ADD_1596_U141 , ADD_1596_U140 );
nand NAND2_11332 ( ADD_1596_U101 , ADD_1596_U137 , ADD_1596_U136 );
not NOT1_11333 ( ADD_1596_U102 , ADD_1596_U9 );
nand NAND2_11334 ( ADD_1596_U103 , ADD_1596_U102 , ADD_1596_U10 );
nand NAND2_11335 ( ADD_1596_U104 , ADD_1596_U103 , ADD_1596_U91 );
nand NAND2_11336 ( ADD_1596_U105 , P1_ADDR_REG_1_ , ADD_1596_U9 );
not NOT1_11337 ( ADD_1596_U106 , ADD_1596_U90 );
nand NAND2_11338 ( ADD_1596_U107 , P3_ADDR_REG_2_ , ADD_1596_U12 );
nand NAND2_11339 ( ADD_1596_U108 , ADD_1596_U107 , ADD_1596_U90 );
nand NAND2_11340 ( ADD_1596_U109 , P1_ADDR_REG_2_ , ADD_1596_U11 );
not NOT1_11341 ( ADD_1596_U110 , ADD_1596_U89 );
nand NAND2_11342 ( ADD_1596_U111 , P3_ADDR_REG_3_ , ADD_1596_U14 );
nand NAND2_11343 ( ADD_1596_U112 , ADD_1596_U111 , ADD_1596_U89 );
nand NAND2_11344 ( ADD_1596_U113 , P1_ADDR_REG_3_ , ADD_1596_U13 );
not NOT1_11345 ( ADD_1596_U114 , ADD_1596_U88 );
nand NAND2_11346 ( ADD_1596_U115 , P3_ADDR_REG_4_ , ADD_1596_U16 );
nand NAND2_11347 ( ADD_1596_U116 , ADD_1596_U115 , ADD_1596_U88 );
nand NAND2_11348 ( ADD_1596_U117 , P1_ADDR_REG_4_ , ADD_1596_U15 );
not NOT1_11349 ( ADD_1596_U118 , ADD_1596_U87 );
nand NAND2_11350 ( ADD_1596_U119 , P3_ADDR_REG_5_ , ADD_1596_U18 );
nand NAND2_11351 ( ADD_1596_U120 , ADD_1596_U119 , ADD_1596_U87 );
nand NAND2_11352 ( ADD_1596_U121 , P1_ADDR_REG_5_ , ADD_1596_U17 );
not NOT1_11353 ( ADD_1596_U122 , ADD_1596_U86 );
nand NAND2_11354 ( ADD_1596_U123 , P3_ADDR_REG_6_ , ADD_1596_U20 );
nand NAND2_11355 ( ADD_1596_U124 , ADD_1596_U123 , ADD_1596_U86 );
nand NAND2_11356 ( ADD_1596_U125 , P1_ADDR_REG_6_ , ADD_1596_U19 );
not NOT1_11357 ( ADD_1596_U126 , ADD_1596_U85 );
nand NAND2_11358 ( ADD_1596_U127 , P3_ADDR_REG_7_ , ADD_1596_U22 );
nand NAND2_11359 ( ADD_1596_U128 , ADD_1596_U127 , ADD_1596_U85 );
nand NAND2_11360 ( ADD_1596_U129 , P1_ADDR_REG_7_ , ADD_1596_U21 );
not NOT1_11361 ( ADD_1596_U130 , ADD_1596_U84 );
nand NAND2_11362 ( ADD_1596_U131 , P3_ADDR_REG_8_ , ADD_1596_U24 );
nand NAND2_11363 ( ADD_1596_U132 , ADD_1596_U131 , ADD_1596_U84 );
nand NAND2_11364 ( ADD_1596_U133 , P1_ADDR_REG_8_ , ADD_1596_U23 );
not NOT1_11365 ( ADD_1596_U134 , ADD_1596_U83 );
nand NAND2_11366 ( ADD_1596_U135 , P3_ADDR_REG_9_ , ADD_1596_U26 );
nand NAND2_11367 ( ADD_1596_U136 , ADD_1596_U135 , ADD_1596_U83 );
nand NAND2_11368 ( ADD_1596_U137 , P1_ADDR_REG_9_ , ADD_1596_U25 );
not NOT1_11369 ( ADD_1596_U138 , ADD_1596_U101 );
nand NAND2_11370 ( ADD_1596_U139 , P3_ADDR_REG_10_ , ADD_1596_U28 );
nand NAND2_11371 ( ADD_1596_U140 , ADD_1596_U139 , ADD_1596_U101 );
nand NAND2_11372 ( ADD_1596_U141 , P1_ADDR_REG_10_ , ADD_1596_U27 );
not NOT1_11373 ( ADD_1596_U142 , ADD_1596_U100 );
nand NAND2_11374 ( ADD_1596_U143 , P3_ADDR_REG_11_ , ADD_1596_U30 );
nand NAND2_11375 ( ADD_1596_U144 , ADD_1596_U143 , ADD_1596_U100 );
nand NAND2_11376 ( ADD_1596_U145 , P1_ADDR_REG_11_ , ADD_1596_U29 );
not NOT1_11377 ( ADD_1596_U146 , ADD_1596_U99 );
nand NAND2_11378 ( ADD_1596_U147 , P3_ADDR_REG_12_ , ADD_1596_U32 );
nand NAND2_11379 ( ADD_1596_U148 , ADD_1596_U147 , ADD_1596_U99 );
nand NAND2_11380 ( ADD_1596_U149 , P1_ADDR_REG_12_ , ADD_1596_U31 );
not NOT1_11381 ( ADD_1596_U150 , ADD_1596_U98 );
nand NAND2_11382 ( ADD_1596_U151 , P3_ADDR_REG_13_ , ADD_1596_U34 );
nand NAND2_11383 ( ADD_1596_U152 , ADD_1596_U151 , ADD_1596_U98 );
nand NAND2_11384 ( ADD_1596_U153 , P1_ADDR_REG_13_ , ADD_1596_U33 );
not NOT1_11385 ( ADD_1596_U154 , ADD_1596_U97 );
nand NAND2_11386 ( ADD_1596_U155 , P3_ADDR_REG_14_ , ADD_1596_U36 );
nand NAND2_11387 ( ADD_1596_U156 , ADD_1596_U155 , ADD_1596_U97 );
nand NAND2_11388 ( ADD_1596_U157 , P1_ADDR_REG_14_ , ADD_1596_U35 );
not NOT1_11389 ( ADD_1596_U158 , ADD_1596_U96 );
nand NAND2_11390 ( ADD_1596_U159 , P3_ADDR_REG_15_ , ADD_1596_U38 );
nand NAND2_11391 ( ADD_1596_U160 , ADD_1596_U159 , ADD_1596_U96 );
nand NAND2_11392 ( ADD_1596_U161 , P1_ADDR_REG_15_ , ADD_1596_U37 );
not NOT1_11393 ( ADD_1596_U162 , ADD_1596_U95 );
nand NAND2_11394 ( ADD_1596_U163 , P3_ADDR_REG_16_ , ADD_1596_U40 );
nand NAND2_11395 ( ADD_1596_U164 , ADD_1596_U163 , ADD_1596_U95 );
nand NAND2_11396 ( ADD_1596_U165 , P1_ADDR_REG_16_ , ADD_1596_U39 );
not NOT1_11397 ( ADD_1596_U166 , ADD_1596_U94 );
nand NAND2_11398 ( ADD_1596_U167 , P3_ADDR_REG_17_ , ADD_1596_U42 );
nand NAND2_11399 ( ADD_1596_U168 , ADD_1596_U167 , ADD_1596_U94 );
nand NAND2_11400 ( ADD_1596_U169 , P1_ADDR_REG_17_ , ADD_1596_U41 );
not NOT1_11401 ( ADD_1596_U170 , ADD_1596_U45 );
nand NAND2_11402 ( ADD_1596_U171 , P1_ADDR_REG_18_ , ADD_1596_U43 );
nand NAND2_11403 ( ADD_1596_U172 , ADD_1596_U170 , ADD_1596_U171 );
nand NAND2_11404 ( ADD_1596_U173 , P3_ADDR_REG_18_ , ADD_1596_U44 );
nand NAND3_11405 ( ADD_1596_U174 , ADD_1596_U173 , ADD_1596_U229 , ADD_1596_U172 );
nand NAND2_11406 ( ADD_1596_U175 , P3_ADDR_REG_18_ , ADD_1596_U44 );
nand NAND2_11407 ( ADD_1596_U176 , ADD_1596_U175 , ADD_1596_U45 );
nand NAND2_11408 ( ADD_1596_U177 , P1_ADDR_REG_18_ , ADD_1596_U43 );
nand NAND4_11409 ( ADD_1596_U178 , ADD_1596_U226 , ADD_1596_U225 , ADD_1596_U177 , ADD_1596_U176 );
nand NAND2_11410 ( ADD_1596_U179 , P1_ADDR_REG_0_ , ADD_1596_U8 );
nand NAND2_11411 ( ADD_1596_U180 , P3_ADDR_REG_9_ , ADD_1596_U26 );
nand NAND2_11412 ( ADD_1596_U181 , P1_ADDR_REG_9_ , ADD_1596_U25 );
not NOT1_11413 ( ADD_1596_U182 , ADD_1596_U65 );
nand NAND2_11414 ( ADD_1596_U183 , ADD_1596_U134 , ADD_1596_U182 );
nand NAND2_11415 ( ADD_1596_U184 , ADD_1596_U65 , ADD_1596_U83 );
nand NAND2_11416 ( ADD_1596_U185 , P3_ADDR_REG_8_ , ADD_1596_U24 );
nand NAND2_11417 ( ADD_1596_U186 , P1_ADDR_REG_8_ , ADD_1596_U23 );
not NOT1_11418 ( ADD_1596_U187 , ADD_1596_U66 );
nand NAND2_11419 ( ADD_1596_U188 , ADD_1596_U130 , ADD_1596_U187 );
nand NAND2_11420 ( ADD_1596_U189 , ADD_1596_U66 , ADD_1596_U84 );
nand NAND2_11421 ( ADD_1596_U190 , P3_ADDR_REG_7_ , ADD_1596_U22 );
nand NAND2_11422 ( ADD_1596_U191 , P1_ADDR_REG_7_ , ADD_1596_U21 );
not NOT1_11423 ( ADD_1596_U192 , ADD_1596_U67 );
nand NAND2_11424 ( ADD_1596_U193 , ADD_1596_U126 , ADD_1596_U192 );
nand NAND2_11425 ( ADD_1596_U194 , ADD_1596_U67 , ADD_1596_U85 );
nand NAND2_11426 ( ADD_1596_U195 , P3_ADDR_REG_6_ , ADD_1596_U20 );
nand NAND2_11427 ( ADD_1596_U196 , P1_ADDR_REG_6_ , ADD_1596_U19 );
not NOT1_11428 ( ADD_1596_U197 , ADD_1596_U68 );
nand NAND2_11429 ( ADD_1596_U198 , ADD_1596_U122 , ADD_1596_U197 );
nand NAND2_11430 ( ADD_1596_U199 , ADD_1596_U68 , ADD_1596_U86 );
nand NAND2_11431 ( ADD_1596_U200 , P3_ADDR_REG_5_ , ADD_1596_U18 );
nand NAND2_11432 ( ADD_1596_U201 , P1_ADDR_REG_5_ , ADD_1596_U17 );
not NOT1_11433 ( ADD_1596_U202 , ADD_1596_U69 );
nand NAND2_11434 ( ADD_1596_U203 , ADD_1596_U118 , ADD_1596_U202 );
nand NAND2_11435 ( ADD_1596_U204 , ADD_1596_U69 , ADD_1596_U87 );
nand NAND2_11436 ( ADD_1596_U205 , P3_ADDR_REG_4_ , ADD_1596_U16 );
nand NAND2_11437 ( ADD_1596_U206 , P1_ADDR_REG_4_ , ADD_1596_U15 );
not NOT1_11438 ( ADD_1596_U207 , ADD_1596_U70 );
nand NAND2_11439 ( ADD_1596_U208 , ADD_1596_U114 , ADD_1596_U207 );
nand NAND2_11440 ( ADD_1596_U209 , ADD_1596_U70 , ADD_1596_U88 );
nand NAND2_11441 ( ADD_1596_U210 , P3_ADDR_REG_3_ , ADD_1596_U14 );
nand NAND2_11442 ( ADD_1596_U211 , P1_ADDR_REG_3_ , ADD_1596_U13 );
not NOT1_11443 ( ADD_1596_U212 , ADD_1596_U71 );
nand NAND2_11444 ( ADD_1596_U213 , ADD_1596_U110 , ADD_1596_U212 );
nand NAND2_11445 ( ADD_1596_U214 , ADD_1596_U71 , ADD_1596_U89 );
nand NAND2_11446 ( ADD_1596_U215 , P3_ADDR_REG_2_ , ADD_1596_U12 );
nand NAND2_11447 ( ADD_1596_U216 , P1_ADDR_REG_2_ , ADD_1596_U11 );
not NOT1_11448 ( ADD_1596_U217 , ADD_1596_U72 );
nand NAND2_11449 ( ADD_1596_U218 , ADD_1596_U106 , ADD_1596_U217 );
nand NAND2_11450 ( ADD_1596_U219 , ADD_1596_U72 , ADD_1596_U90 );
nand NAND2_11451 ( ADD_1596_U220 , P3_ADDR_REG_1_ , ADD_1596_U10 );
nand NAND2_11452 ( ADD_1596_U221 , P1_ADDR_REG_1_ , ADD_1596_U91 );
not NOT1_11453 ( ADD_1596_U222 , ADD_1596_U73 );
nand NAND2_11454 ( ADD_1596_U223 , ADD_1596_U222 , ADD_1596_U102 );
nand NAND2_11455 ( ADD_1596_U224 , ADD_1596_U73 , ADD_1596_U9 );
nand NAND2_11456 ( ADD_1596_U225 , P3_ADDR_REG_19_ , ADD_1596_U93 );
nand NAND2_11457 ( ADD_1596_U226 , P1_ADDR_REG_19_ , ADD_1596_U92 );
nand NAND2_11458 ( ADD_1596_U227 , P3_ADDR_REG_19_ , ADD_1596_U93 );
nand NAND2_11459 ( ADD_1596_U228 , P1_ADDR_REG_19_ , ADD_1596_U92 );
nand NAND2_11460 ( ADD_1596_U229 , ADD_1596_U228 , ADD_1596_U227 );
nand NAND2_11461 ( ADD_1596_U230 , P3_ADDR_REG_18_ , ADD_1596_U44 );
nand NAND2_11462 ( ADD_1596_U231 , P1_ADDR_REG_18_ , ADD_1596_U43 );
not NOT1_11463 ( ADD_1596_U232 , ADD_1596_U74 );
nand NAND2_11464 ( ADD_1596_U233 , ADD_1596_U232 , ADD_1596_U170 );
nand NAND2_11465 ( ADD_1596_U234 , ADD_1596_U74 , ADD_1596_U45 );
nand NAND2_11466 ( ADD_1596_U235 , P3_ADDR_REG_17_ , ADD_1596_U42 );
nand NAND2_11467 ( ADD_1596_U236 , P1_ADDR_REG_17_ , ADD_1596_U41 );
not NOT1_11468 ( ADD_1596_U237 , ADD_1596_U75 );
nand NAND2_11469 ( ADD_1596_U238 , ADD_1596_U166 , ADD_1596_U237 );
nand NAND2_11470 ( ADD_1596_U239 , ADD_1596_U75 , ADD_1596_U94 );
nand NAND2_11471 ( ADD_1596_U240 , P3_ADDR_REG_16_ , ADD_1596_U40 );
nand NAND2_11472 ( ADD_1596_U241 , P1_ADDR_REG_16_ , ADD_1596_U39 );
not NOT1_11473 ( ADD_1596_U242 , ADD_1596_U76 );
nand NAND2_11474 ( ADD_1596_U243 , ADD_1596_U162 , ADD_1596_U242 );
nand NAND2_11475 ( ADD_1596_U244 , ADD_1596_U76 , ADD_1596_U95 );
nand NAND2_11476 ( ADD_1596_U245 , P3_ADDR_REG_15_ , ADD_1596_U38 );
nand NAND2_11477 ( ADD_1596_U246 , P1_ADDR_REG_15_ , ADD_1596_U37 );
not NOT1_11478 ( ADD_1596_U247 , ADD_1596_U77 );
nand NAND2_11479 ( ADD_1596_U248 , ADD_1596_U158 , ADD_1596_U247 );
nand NAND2_11480 ( ADD_1596_U249 , ADD_1596_U77 , ADD_1596_U96 );
nand NAND2_11481 ( ADD_1596_U250 , P3_ADDR_REG_14_ , ADD_1596_U36 );
nand NAND2_11482 ( ADD_1596_U251 , P1_ADDR_REG_14_ , ADD_1596_U35 );
not NOT1_11483 ( ADD_1596_U252 , ADD_1596_U78 );
nand NAND2_11484 ( ADD_1596_U253 , ADD_1596_U154 , ADD_1596_U252 );
nand NAND2_11485 ( ADD_1596_U254 , ADD_1596_U78 , ADD_1596_U97 );
nand NAND2_11486 ( ADD_1596_U255 , P3_ADDR_REG_13_ , ADD_1596_U34 );
nand NAND2_11487 ( ADD_1596_U256 , P1_ADDR_REG_13_ , ADD_1596_U33 );
not NOT1_11488 ( ADD_1596_U257 , ADD_1596_U79 );
nand NAND2_11489 ( ADD_1596_U258 , ADD_1596_U150 , ADD_1596_U257 );
nand NAND2_11490 ( ADD_1596_U259 , ADD_1596_U79 , ADD_1596_U98 );
nand NAND2_11491 ( ADD_1596_U260 , P3_ADDR_REG_12_ , ADD_1596_U32 );
nand NAND2_11492 ( ADD_1596_U261 , P1_ADDR_REG_12_ , ADD_1596_U31 );
not NOT1_11493 ( ADD_1596_U262 , ADD_1596_U80 );
nand NAND2_11494 ( ADD_1596_U263 , ADD_1596_U146 , ADD_1596_U262 );
nand NAND2_11495 ( ADD_1596_U264 , ADD_1596_U80 , ADD_1596_U99 );
nand NAND2_11496 ( ADD_1596_U265 , P3_ADDR_REG_11_ , ADD_1596_U30 );
nand NAND2_11497 ( ADD_1596_U266 , P1_ADDR_REG_11_ , ADD_1596_U29 );
not NOT1_11498 ( ADD_1596_U267 , ADD_1596_U81 );
nand NAND2_11499 ( ADD_1596_U268 , ADD_1596_U142 , ADD_1596_U267 );
nand NAND2_11500 ( ADD_1596_U269 , ADD_1596_U81 , ADD_1596_U100 );
nand NAND2_11501 ( ADD_1596_U270 , P3_ADDR_REG_10_ , ADD_1596_U28 );
nand NAND2_11502 ( ADD_1596_U271 , P1_ADDR_REG_10_ , ADD_1596_U27 );
not NOT1_11503 ( ADD_1596_U272 , ADD_1596_U82 );
nand NAND2_11504 ( ADD_1596_U273 , ADD_1596_U138 , ADD_1596_U272 );
nand NAND2_11505 ( ADD_1596_U274 , ADD_1596_U82 , ADD_1596_U101 );
not NOT1_11506 ( LT_1601_21_U6 , P2_ADDR_REG_19_ );
not NOT1_11507 ( P1_ADD_99_U4 , P1_REG3_REG_3_ );
and AND3_11508 ( P1_ADD_99_U5 , P1_REG3_REG_28_ , P1_REG3_REG_27_ , P1_ADD_99_U102 );
not NOT1_11509 ( P1_ADD_99_U6 , P1_REG3_REG_4_ );
nand NAND2_11510 ( P1_ADD_99_U7 , P1_REG3_REG_4_ , P1_REG3_REG_3_ );
not NOT1_11511 ( P1_ADD_99_U8 , P1_REG3_REG_5_ );
nand NAND2_11512 ( P1_ADD_99_U9 , P1_REG3_REG_5_ , P1_ADD_99_U80 );
not NOT1_11513 ( P1_ADD_99_U10 , P1_REG3_REG_6_ );
nand NAND2_11514 ( P1_ADD_99_U11 , P1_REG3_REG_6_ , P1_ADD_99_U81 );
not NOT1_11515 ( P1_ADD_99_U12 , P1_REG3_REG_7_ );
nand NAND2_11516 ( P1_ADD_99_U13 , P1_REG3_REG_7_ , P1_ADD_99_U82 );
not NOT1_11517 ( P1_ADD_99_U14 , P1_REG3_REG_8_ );
not NOT1_11518 ( P1_ADD_99_U15 , P1_REG3_REG_9_ );
nand NAND2_11519 ( P1_ADD_99_U16 , P1_REG3_REG_8_ , P1_ADD_99_U83 );
nand NAND2_11520 ( P1_ADD_99_U17 , P1_ADD_99_U84 , P1_REG3_REG_9_ );
not NOT1_11521 ( P1_ADD_99_U18 , P1_REG3_REG_10_ );
nand NAND2_11522 ( P1_ADD_99_U19 , P1_REG3_REG_10_ , P1_ADD_99_U85 );
not NOT1_11523 ( P1_ADD_99_U20 , P1_REG3_REG_11_ );
nand NAND2_11524 ( P1_ADD_99_U21 , P1_REG3_REG_11_ , P1_ADD_99_U86 );
not NOT1_11525 ( P1_ADD_99_U22 , P1_REG3_REG_12_ );
nand NAND2_11526 ( P1_ADD_99_U23 , P1_REG3_REG_12_ , P1_ADD_99_U87 );
not NOT1_11527 ( P1_ADD_99_U24 , P1_REG3_REG_13_ );
nand NAND2_11528 ( P1_ADD_99_U25 , P1_REG3_REG_13_ , P1_ADD_99_U88 );
not NOT1_11529 ( P1_ADD_99_U26 , P1_REG3_REG_14_ );
nand NAND2_11530 ( P1_ADD_99_U27 , P1_REG3_REG_14_ , P1_ADD_99_U89 );
not NOT1_11531 ( P1_ADD_99_U28 , P1_REG3_REG_15_ );
nand NAND2_11532 ( P1_ADD_99_U29 , P1_REG3_REG_15_ , P1_ADD_99_U90 );
not NOT1_11533 ( P1_ADD_99_U30 , P1_REG3_REG_16_ );
nand NAND2_11534 ( P1_ADD_99_U31 , P1_REG3_REG_16_ , P1_ADD_99_U91 );
not NOT1_11535 ( P1_ADD_99_U32 , P1_REG3_REG_17_ );
nand NAND2_11536 ( P1_ADD_99_U33 , P1_REG3_REG_17_ , P1_ADD_99_U92 );
not NOT1_11537 ( P1_ADD_99_U34 , P1_REG3_REG_18_ );
nand NAND2_11538 ( P1_ADD_99_U35 , P1_REG3_REG_18_ , P1_ADD_99_U93 );
not NOT1_11539 ( P1_ADD_99_U36 , P1_REG3_REG_19_ );
nand NAND2_11540 ( P1_ADD_99_U37 , P1_REG3_REG_19_ , P1_ADD_99_U94 );
not NOT1_11541 ( P1_ADD_99_U38 , P1_REG3_REG_20_ );
nand NAND2_11542 ( P1_ADD_99_U39 , P1_REG3_REG_20_ , P1_ADD_99_U95 );
not NOT1_11543 ( P1_ADD_99_U40 , P1_REG3_REG_21_ );
nand NAND2_11544 ( P1_ADD_99_U41 , P1_REG3_REG_21_ , P1_ADD_99_U96 );
not NOT1_11545 ( P1_ADD_99_U42 , P1_REG3_REG_22_ );
nand NAND2_11546 ( P1_ADD_99_U43 , P1_REG3_REG_22_ , P1_ADD_99_U97 );
not NOT1_11547 ( P1_ADD_99_U44 , P1_REG3_REG_23_ );
nand NAND2_11548 ( P1_ADD_99_U45 , P1_REG3_REG_23_ , P1_ADD_99_U98 );
not NOT1_11549 ( P1_ADD_99_U46 , P1_REG3_REG_24_ );
nand NAND2_11550 ( P1_ADD_99_U47 , P1_REG3_REG_24_ , P1_ADD_99_U99 );
not NOT1_11551 ( P1_ADD_99_U48 , P1_REG3_REG_25_ );
nand NAND2_11552 ( P1_ADD_99_U49 , P1_REG3_REG_25_ , P1_ADD_99_U100 );
not NOT1_11553 ( P1_ADD_99_U50 , P1_REG3_REG_26_ );
nand NAND2_11554 ( P1_ADD_99_U51 , P1_REG3_REG_26_ , P1_ADD_99_U101 );
not NOT1_11555 ( P1_ADD_99_U52 , P1_REG3_REG_28_ );
not NOT1_11556 ( P1_ADD_99_U53 , P1_REG3_REG_27_ );
nand NAND2_11557 ( P1_ADD_99_U54 , P1_ADD_99_U105 , P1_ADD_99_U104 );
nand NAND2_11558 ( P1_ADD_99_U55 , P1_ADD_99_U107 , P1_ADD_99_U106 );
nand NAND2_11559 ( P1_ADD_99_U56 , P1_ADD_99_U109 , P1_ADD_99_U108 );
nand NAND2_11560 ( P1_ADD_99_U57 , P1_ADD_99_U111 , P1_ADD_99_U110 );
nand NAND2_11561 ( P1_ADD_99_U58 , P1_ADD_99_U113 , P1_ADD_99_U112 );
nand NAND2_11562 ( P1_ADD_99_U59 , P1_ADD_99_U115 , P1_ADD_99_U114 );
nand NAND2_11563 ( P1_ADD_99_U60 , P1_ADD_99_U117 , P1_ADD_99_U116 );
nand NAND2_11564 ( P1_ADD_99_U61 , P1_ADD_99_U119 , P1_ADD_99_U118 );
nand NAND2_11565 ( P1_ADD_99_U62 , P1_ADD_99_U121 , P1_ADD_99_U120 );
nand NAND2_11566 ( P1_ADD_99_U63 , P1_ADD_99_U123 , P1_ADD_99_U122 );
nand NAND2_11567 ( P1_ADD_99_U64 , P1_ADD_99_U125 , P1_ADD_99_U124 );
nand NAND2_11568 ( P1_ADD_99_U65 , P1_ADD_99_U127 , P1_ADD_99_U126 );
nand NAND2_11569 ( P1_ADD_99_U66 , P1_ADD_99_U129 , P1_ADD_99_U128 );
nand NAND2_11570 ( P1_ADD_99_U67 , P1_ADD_99_U131 , P1_ADD_99_U130 );
nand NAND2_11571 ( P1_ADD_99_U68 , P1_ADD_99_U133 , P1_ADD_99_U132 );
nand NAND2_11572 ( P1_ADD_99_U69 , P1_ADD_99_U135 , P1_ADD_99_U134 );
nand NAND2_11573 ( P1_ADD_99_U70 , P1_ADD_99_U137 , P1_ADD_99_U136 );
nand NAND2_11574 ( P1_ADD_99_U71 , P1_ADD_99_U139 , P1_ADD_99_U138 );
nand NAND2_11575 ( P1_ADD_99_U72 , P1_ADD_99_U141 , P1_ADD_99_U140 );
nand NAND2_11576 ( P1_ADD_99_U73 , P1_ADD_99_U143 , P1_ADD_99_U142 );
nand NAND2_11577 ( P1_ADD_99_U74 , P1_ADD_99_U145 , P1_ADD_99_U144 );
nand NAND2_11578 ( P1_ADD_99_U75 , P1_ADD_99_U147 , P1_ADD_99_U146 );
nand NAND2_11579 ( P1_ADD_99_U76 , P1_ADD_99_U149 , P1_ADD_99_U148 );
nand NAND2_11580 ( P1_ADD_99_U77 , P1_ADD_99_U151 , P1_ADD_99_U150 );
nand NAND2_11581 ( P1_ADD_99_U78 , P1_ADD_99_U153 , P1_ADD_99_U152 );
nand NAND2_11582 ( P1_ADD_99_U79 , P1_REG3_REG_27_ , P1_ADD_99_U102 );
not NOT1_11583 ( P1_ADD_99_U80 , P1_ADD_99_U7 );
not NOT1_11584 ( P1_ADD_99_U81 , P1_ADD_99_U9 );
not NOT1_11585 ( P1_ADD_99_U82 , P1_ADD_99_U11 );
not NOT1_11586 ( P1_ADD_99_U83 , P1_ADD_99_U13 );
not NOT1_11587 ( P1_ADD_99_U84 , P1_ADD_99_U16 );
not NOT1_11588 ( P1_ADD_99_U85 , P1_ADD_99_U17 );
not NOT1_11589 ( P1_ADD_99_U86 , P1_ADD_99_U19 );
not NOT1_11590 ( P1_ADD_99_U87 , P1_ADD_99_U21 );
not NOT1_11591 ( P1_ADD_99_U88 , P1_ADD_99_U23 );
not NOT1_11592 ( P1_ADD_99_U89 , P1_ADD_99_U25 );
not NOT1_11593 ( P1_ADD_99_U90 , P1_ADD_99_U27 );
not NOT1_11594 ( P1_ADD_99_U91 , P1_ADD_99_U29 );
not NOT1_11595 ( P1_ADD_99_U92 , P1_ADD_99_U31 );
not NOT1_11596 ( P1_ADD_99_U93 , P1_ADD_99_U33 );
not NOT1_11597 ( P1_ADD_99_U94 , P1_ADD_99_U35 );
not NOT1_11598 ( P1_ADD_99_U95 , P1_ADD_99_U37 );
not NOT1_11599 ( P1_ADD_99_U96 , P1_ADD_99_U39 );
not NOT1_11600 ( P1_ADD_99_U97 , P1_ADD_99_U41 );
not NOT1_11601 ( P1_ADD_99_U98 , P1_ADD_99_U43 );
not NOT1_11602 ( P1_ADD_99_U99 , P1_ADD_99_U45 );
not NOT1_11603 ( P1_ADD_99_U100 , P1_ADD_99_U47 );
not NOT1_11604 ( P1_ADD_99_U101 , P1_ADD_99_U49 );
not NOT1_11605 ( P1_ADD_99_U102 , P1_ADD_99_U51 );
not NOT1_11606 ( P1_ADD_99_U103 , P1_ADD_99_U79 );
nand NAND2_11607 ( P1_ADD_99_U104 , P1_REG3_REG_9_ , P1_ADD_99_U16 );
nand NAND2_11608 ( P1_ADD_99_U105 , P1_ADD_99_U84 , P1_ADD_99_U15 );
nand NAND2_11609 ( P1_ADD_99_U106 , P1_REG3_REG_8_ , P1_ADD_99_U13 );
nand NAND2_11610 ( P1_ADD_99_U107 , P1_ADD_99_U83 , P1_ADD_99_U14 );
nand NAND2_11611 ( P1_ADD_99_U108 , P1_REG3_REG_7_ , P1_ADD_99_U11 );
nand NAND2_11612 ( P1_ADD_99_U109 , P1_ADD_99_U82 , P1_ADD_99_U12 );
nand NAND2_11613 ( P1_ADD_99_U110 , P1_REG3_REG_6_ , P1_ADD_99_U9 );
nand NAND2_11614 ( P1_ADD_99_U111 , P1_ADD_99_U81 , P1_ADD_99_U10 );
nand NAND2_11615 ( P1_ADD_99_U112 , P1_REG3_REG_5_ , P1_ADD_99_U7 );
nand NAND2_11616 ( P1_ADD_99_U113 , P1_ADD_99_U80 , P1_ADD_99_U8 );
nand NAND2_11617 ( P1_ADD_99_U114 , P1_REG3_REG_4_ , P1_ADD_99_U4 );
nand NAND2_11618 ( P1_ADD_99_U115 , P1_REG3_REG_3_ , P1_ADD_99_U6 );
nand NAND2_11619 ( P1_ADD_99_U116 , P1_REG3_REG_28_ , P1_ADD_99_U79 );
nand NAND2_11620 ( P1_ADD_99_U117 , P1_ADD_99_U103 , P1_ADD_99_U52 );
nand NAND2_11621 ( P1_ADD_99_U118 , P1_REG3_REG_27_ , P1_ADD_99_U51 );
nand NAND2_11622 ( P1_ADD_99_U119 , P1_ADD_99_U102 , P1_ADD_99_U53 );
nand NAND2_11623 ( P1_ADD_99_U120 , P1_REG3_REG_26_ , P1_ADD_99_U49 );
nand NAND2_11624 ( P1_ADD_99_U121 , P1_ADD_99_U101 , P1_ADD_99_U50 );
nand NAND2_11625 ( P1_ADD_99_U122 , P1_REG3_REG_25_ , P1_ADD_99_U47 );
nand NAND2_11626 ( P1_ADD_99_U123 , P1_ADD_99_U100 , P1_ADD_99_U48 );
nand NAND2_11627 ( P1_ADD_99_U124 , P1_REG3_REG_24_ , P1_ADD_99_U45 );
nand NAND2_11628 ( P1_ADD_99_U125 , P1_ADD_99_U99 , P1_ADD_99_U46 );
nand NAND2_11629 ( P1_ADD_99_U126 , P1_REG3_REG_23_ , P1_ADD_99_U43 );
nand NAND2_11630 ( P1_ADD_99_U127 , P1_ADD_99_U98 , P1_ADD_99_U44 );
nand NAND2_11631 ( P1_ADD_99_U128 , P1_REG3_REG_22_ , P1_ADD_99_U41 );
nand NAND2_11632 ( P1_ADD_99_U129 , P1_ADD_99_U97 , P1_ADD_99_U42 );
nand NAND2_11633 ( P1_ADD_99_U130 , P1_REG3_REG_21_ , P1_ADD_99_U39 );
nand NAND2_11634 ( P1_ADD_99_U131 , P1_ADD_99_U96 , P1_ADD_99_U40 );
nand NAND2_11635 ( P1_ADD_99_U132 , P1_REG3_REG_20_ , P1_ADD_99_U37 );
nand NAND2_11636 ( P1_ADD_99_U133 , P1_ADD_99_U95 , P1_ADD_99_U38 );
nand NAND2_11637 ( P1_ADD_99_U134 , P1_REG3_REG_19_ , P1_ADD_99_U35 );
nand NAND2_11638 ( P1_ADD_99_U135 , P1_ADD_99_U94 , P1_ADD_99_U36 );
nand NAND2_11639 ( P1_ADD_99_U136 , P1_REG3_REG_18_ , P1_ADD_99_U33 );
nand NAND2_11640 ( P1_ADD_99_U137 , P1_ADD_99_U93 , P1_ADD_99_U34 );
nand NAND2_11641 ( P1_ADD_99_U138 , P1_REG3_REG_17_ , P1_ADD_99_U31 );
nand NAND2_11642 ( P1_ADD_99_U139 , P1_ADD_99_U92 , P1_ADD_99_U32 );
nand NAND2_11643 ( P1_ADD_99_U140 , P1_REG3_REG_16_ , P1_ADD_99_U29 );
nand NAND2_11644 ( P1_ADD_99_U141 , P1_ADD_99_U91 , P1_ADD_99_U30 );
nand NAND2_11645 ( P1_ADD_99_U142 , P1_REG3_REG_15_ , P1_ADD_99_U27 );
nand NAND2_11646 ( P1_ADD_99_U143 , P1_ADD_99_U90 , P1_ADD_99_U28 );
nand NAND2_11647 ( P1_ADD_99_U144 , P1_REG3_REG_14_ , P1_ADD_99_U25 );
nand NAND2_11648 ( P1_ADD_99_U145 , P1_ADD_99_U89 , P1_ADD_99_U26 );
nand NAND2_11649 ( P1_ADD_99_U146 , P1_REG3_REG_13_ , P1_ADD_99_U23 );
nand NAND2_11650 ( P1_ADD_99_U147 , P1_ADD_99_U88 , P1_ADD_99_U24 );
nand NAND2_11651 ( P1_ADD_99_U148 , P1_REG3_REG_12_ , P1_ADD_99_U21 );
nand NAND2_11652 ( P1_ADD_99_U149 , P1_ADD_99_U87 , P1_ADD_99_U22 );
nand NAND2_11653 ( P1_ADD_99_U150 , P1_REG3_REG_11_ , P1_ADD_99_U19 );
nand NAND2_11654 ( P1_ADD_99_U151 , P1_ADD_99_U86 , P1_ADD_99_U20 );
nand NAND2_11655 ( P1_ADD_99_U152 , P1_REG3_REG_10_ , P1_ADD_99_U17 );
nand NAND2_11656 ( P1_ADD_99_U153 , P1_ADD_99_U85 , P1_ADD_99_U18 );
and AND2_11657 ( P1_R1105_U4 , P1_R1105_U95 , P1_R1105_U94 );
and AND2_11658 ( P1_R1105_U5 , P1_R1105_U96 , P1_R1105_U97 );
and AND2_11659 ( P1_R1105_U6 , P1_R1105_U113 , P1_R1105_U112 );
and AND2_11660 ( P1_R1105_U7 , P1_R1105_U155 , P1_R1105_U154 );
and AND2_11661 ( P1_R1105_U8 , P1_R1105_U164 , P1_R1105_U163 );
and AND2_11662 ( P1_R1105_U9 , P1_R1105_U182 , P1_R1105_U181 );
and AND2_11663 ( P1_R1105_U10 , P1_R1105_U218 , P1_R1105_U215 );
and AND2_11664 ( P1_R1105_U11 , P1_R1105_U211 , P1_R1105_U208 );
and AND2_11665 ( P1_R1105_U12 , P1_R1105_U202 , P1_R1105_U199 );
and AND2_11666 ( P1_R1105_U13 , P1_R1105_U196 , P1_R1105_U192 );
and AND2_11667 ( P1_R1105_U14 , P1_R1105_U151 , P1_R1105_U148 );
and AND2_11668 ( P1_R1105_U15 , P1_R1105_U143 , P1_R1105_U140 );
and AND2_11669 ( P1_R1105_U16 , P1_R1105_U129 , P1_R1105_U126 );
not NOT1_11670 ( P1_R1105_U17 , P1_REG2_REG_6_ );
not NOT1_11671 ( P1_R1105_U18 , P1_U3475 );
not NOT1_11672 ( P1_R1105_U19 , P1_U3478 );
nand NAND2_11673 ( P1_R1105_U20 , P1_U3475 , P1_REG2_REG_6_ );
not NOT1_11674 ( P1_R1105_U21 , P1_REG2_REG_7_ );
not NOT1_11675 ( P1_R1105_U22 , P1_REG2_REG_4_ );
not NOT1_11676 ( P1_R1105_U23 , P1_U3469 );
not NOT1_11677 ( P1_R1105_U24 , P1_U3472 );
not NOT1_11678 ( P1_R1105_U25 , P1_REG2_REG_2_ );
not NOT1_11679 ( P1_R1105_U26 , P1_U3463 );
not NOT1_11680 ( P1_R1105_U27 , P1_REG2_REG_0_ );
not NOT1_11681 ( P1_R1105_U28 , P1_U3454 );
nand NAND2_11682 ( P1_R1105_U29 , P1_U3454 , P1_REG2_REG_0_ );
not NOT1_11683 ( P1_R1105_U30 , P1_REG2_REG_3_ );
not NOT1_11684 ( P1_R1105_U31 , P1_U3466 );
nand NAND2_11685 ( P1_R1105_U32 , P1_U3469 , P1_REG2_REG_4_ );
not NOT1_11686 ( P1_R1105_U33 , P1_REG2_REG_5_ );
not NOT1_11687 ( P1_R1105_U34 , P1_REG2_REG_8_ );
not NOT1_11688 ( P1_R1105_U35 , P1_U3481 );
not NOT1_11689 ( P1_R1105_U36 , P1_U3484 );
not NOT1_11690 ( P1_R1105_U37 , P1_REG2_REG_9_ );
nand NAND2_11691 ( P1_R1105_U38 , P1_R1105_U49 , P1_R1105_U121 );
nand NAND3_11692 ( P1_R1105_U39 , P1_R1105_U110 , P1_R1105_U108 , P1_R1105_U109 );
nand NAND2_11693 ( P1_R1105_U40 , P1_R1105_U98 , P1_R1105_U99 );
nand NAND2_11694 ( P1_R1105_U41 , P1_REG2_REG_1_ , P1_U3460 );
nand NAND3_11695 ( P1_R1105_U42 , P1_R1105_U136 , P1_R1105_U134 , P1_R1105_U135 );
nand NAND2_11696 ( P1_R1105_U43 , P1_R1105_U132 , P1_R1105_U131 );
not NOT1_11697 ( P1_R1105_U44 , P1_REG2_REG_16_ );
not NOT1_11698 ( P1_R1105_U45 , P1_U3505 );
not NOT1_11699 ( P1_R1105_U46 , P1_U3508 );
nand NAND2_11700 ( P1_R1105_U47 , P1_U3505 , P1_REG2_REG_16_ );
not NOT1_11701 ( P1_R1105_U48 , P1_REG2_REG_17_ );
nand NAND2_11702 ( P1_R1105_U49 , P1_U3481 , P1_REG2_REG_8_ );
not NOT1_11703 ( P1_R1105_U50 , P1_REG2_REG_10_ );
not NOT1_11704 ( P1_R1105_U51 , P1_U3487 );
not NOT1_11705 ( P1_R1105_U52 , P1_REG2_REG_12_ );
not NOT1_11706 ( P1_R1105_U53 , P1_U3493 );
not NOT1_11707 ( P1_R1105_U54 , P1_REG2_REG_11_ );
not NOT1_11708 ( P1_R1105_U55 , P1_U3490 );
nand NAND2_11709 ( P1_R1105_U56 , P1_U3490 , P1_REG2_REG_11_ );
not NOT1_11710 ( P1_R1105_U57 , P1_REG2_REG_13_ );
not NOT1_11711 ( P1_R1105_U58 , P1_U3496 );
not NOT1_11712 ( P1_R1105_U59 , P1_REG2_REG_14_ );
not NOT1_11713 ( P1_R1105_U60 , P1_U3499 );
not NOT1_11714 ( P1_R1105_U61 , P1_REG2_REG_15_ );
not NOT1_11715 ( P1_R1105_U62 , P1_U3502 );
not NOT1_11716 ( P1_R1105_U63 , P1_REG2_REG_18_ );
not NOT1_11717 ( P1_R1105_U64 , P1_U3511 );
nand NAND3_11718 ( P1_R1105_U65 , P1_R1105_U186 , P1_R1105_U185 , P1_R1105_U187 );
nand NAND2_11719 ( P1_R1105_U66 , P1_R1105_U179 , P1_R1105_U178 );
nand NAND2_11720 ( P1_R1105_U67 , P1_R1105_U56 , P1_R1105_U204 );
nand NAND2_11721 ( P1_R1105_U68 , P1_R1105_U259 , P1_R1105_U258 );
nand NAND2_11722 ( P1_R1105_U69 , P1_R1105_U308 , P1_R1105_U307 );
nand NAND2_11723 ( P1_R1105_U70 , P1_R1105_U231 , P1_R1105_U230 );
nand NAND2_11724 ( P1_R1105_U71 , P1_R1105_U236 , P1_R1105_U235 );
nand NAND2_11725 ( P1_R1105_U72 , P1_R1105_U243 , P1_R1105_U242 );
nand NAND2_11726 ( P1_R1105_U73 , P1_R1105_U250 , P1_R1105_U249 );
nand NAND2_11727 ( P1_R1105_U74 , P1_R1105_U255 , P1_R1105_U254 );
nand NAND2_11728 ( P1_R1105_U75 , P1_R1105_U271 , P1_R1105_U270 );
nand NAND2_11729 ( P1_R1105_U76 , P1_R1105_U278 , P1_R1105_U277 );
nand NAND2_11730 ( P1_R1105_U77 , P1_R1105_U285 , P1_R1105_U284 );
nand NAND2_11731 ( P1_R1105_U78 , P1_R1105_U292 , P1_R1105_U291 );
nand NAND2_11732 ( P1_R1105_U79 , P1_R1105_U299 , P1_R1105_U298 );
nand NAND2_11733 ( P1_R1105_U80 , P1_R1105_U304 , P1_R1105_U303 );
nand NAND3_11734 ( P1_R1105_U81 , P1_R1105_U117 , P1_R1105_U116 , P1_R1105_U118 );
nand NAND2_11735 ( P1_R1105_U82 , P1_R1105_U133 , P1_R1105_U145 );
nand NAND2_11736 ( P1_R1105_U83 , P1_R1105_U41 , P1_R1105_U152 );
not NOT1_11737 ( P1_R1105_U84 , P1_U3452 );
not NOT1_11738 ( P1_R1105_U85 , P1_REG2_REG_19_ );
nand NAND2_11739 ( P1_R1105_U86 , P1_R1105_U175 , P1_R1105_U174 );
nand NAND2_11740 ( P1_R1105_U87 , P1_R1105_U171 , P1_R1105_U170 );
nand NAND2_11741 ( P1_R1105_U88 , P1_R1105_U161 , P1_R1105_U160 );
not NOT1_11742 ( P1_R1105_U89 , P1_R1105_U32 );
nand NAND2_11743 ( P1_R1105_U90 , P1_REG2_REG_9_ , P1_U3484 );
nand NAND2_11744 ( P1_R1105_U91 , P1_U3493 , P1_REG2_REG_12_ );
not NOT1_11745 ( P1_R1105_U92 , P1_R1105_U56 );
not NOT1_11746 ( P1_R1105_U93 , P1_R1105_U49 );
or OR2_11747 ( P1_R1105_U94 , P1_U3472 , P1_REG2_REG_5_ );
or OR2_11748 ( P1_R1105_U95 , P1_U3469 , P1_REG2_REG_4_ );
or OR2_11749 ( P1_R1105_U96 , P1_REG2_REG_3_ , P1_U3466 );
or OR2_11750 ( P1_R1105_U97 , P1_REG2_REG_2_ , P1_U3463 );
not NOT1_11751 ( P1_R1105_U98 , P1_R1105_U29 );
or OR2_11752 ( P1_R1105_U99 , P1_REG2_REG_1_ , P1_U3460 );
not NOT1_11753 ( P1_R1105_U100 , P1_R1105_U40 );
not NOT1_11754 ( P1_R1105_U101 , P1_R1105_U41 );
nand NAND2_11755 ( P1_R1105_U102 , P1_R1105_U40 , P1_R1105_U41 );
nand NAND3_11756 ( P1_R1105_U103 , P1_REG2_REG_2_ , P1_U3463 , P1_R1105_U96 );
nand NAND2_11757 ( P1_R1105_U104 , P1_R1105_U5 , P1_R1105_U102 );
nand NAND2_11758 ( P1_R1105_U105 , P1_U3466 , P1_REG2_REG_3_ );
nand NAND3_11759 ( P1_R1105_U106 , P1_R1105_U105 , P1_R1105_U103 , P1_R1105_U104 );
nand NAND2_11760 ( P1_R1105_U107 , P1_R1105_U33 , P1_R1105_U32 );
nand NAND2_11761 ( P1_R1105_U108 , P1_U3472 , P1_R1105_U107 );
nand NAND2_11762 ( P1_R1105_U109 , P1_R1105_U4 , P1_R1105_U106 );
nand NAND2_11763 ( P1_R1105_U110 , P1_REG2_REG_5_ , P1_R1105_U89 );
not NOT1_11764 ( P1_R1105_U111 , P1_R1105_U39 );
or OR2_11765 ( P1_R1105_U112 , P1_U3478 , P1_REG2_REG_7_ );
or OR2_11766 ( P1_R1105_U113 , P1_U3475 , P1_REG2_REG_6_ );
not NOT1_11767 ( P1_R1105_U114 , P1_R1105_U20 );
nand NAND2_11768 ( P1_R1105_U115 , P1_R1105_U21 , P1_R1105_U20 );
nand NAND2_11769 ( P1_R1105_U116 , P1_U3478 , P1_R1105_U115 );
nand NAND2_11770 ( P1_R1105_U117 , P1_REG2_REG_7_ , P1_R1105_U114 );
nand NAND2_11771 ( P1_R1105_U118 , P1_R1105_U6 , P1_R1105_U39 );
not NOT1_11772 ( P1_R1105_U119 , P1_R1105_U81 );
or OR2_11773 ( P1_R1105_U120 , P1_REG2_REG_8_ , P1_U3481 );
nand NAND2_11774 ( P1_R1105_U121 , P1_R1105_U120 , P1_R1105_U81 );
not NOT1_11775 ( P1_R1105_U122 , P1_R1105_U38 );
or OR2_11776 ( P1_R1105_U123 , P1_U3484 , P1_REG2_REG_9_ );
or OR2_11777 ( P1_R1105_U124 , P1_REG2_REG_6_ , P1_U3475 );
nand NAND2_11778 ( P1_R1105_U125 , P1_R1105_U124 , P1_R1105_U39 );
nand NAND4_11779 ( P1_R1105_U126 , P1_R1105_U238 , P1_R1105_U237 , P1_R1105_U20 , P1_R1105_U125 );
nand NAND2_11780 ( P1_R1105_U127 , P1_R1105_U111 , P1_R1105_U20 );
nand NAND2_11781 ( P1_R1105_U128 , P1_REG2_REG_7_ , P1_U3478 );
nand NAND3_11782 ( P1_R1105_U129 , P1_R1105_U128 , P1_R1105_U6 , P1_R1105_U127 );
or OR2_11783 ( P1_R1105_U130 , P1_U3475 , P1_REG2_REG_6_ );
nand NAND2_11784 ( P1_R1105_U131 , P1_R1105_U101 , P1_R1105_U97 );
nand NAND2_11785 ( P1_R1105_U132 , P1_U3463 , P1_REG2_REG_2_ );
not NOT1_11786 ( P1_R1105_U133 , P1_R1105_U43 );
nand NAND2_11787 ( P1_R1105_U134 , P1_R1105_U100 , P1_R1105_U5 );
nand NAND2_11788 ( P1_R1105_U135 , P1_R1105_U43 , P1_R1105_U96 );
nand NAND2_11789 ( P1_R1105_U136 , P1_U3466 , P1_REG2_REG_3_ );
not NOT1_11790 ( P1_R1105_U137 , P1_R1105_U42 );
or OR2_11791 ( P1_R1105_U138 , P1_REG2_REG_4_ , P1_U3469 );
nand NAND2_11792 ( P1_R1105_U139 , P1_R1105_U138 , P1_R1105_U42 );
nand NAND4_11793 ( P1_R1105_U140 , P1_R1105_U245 , P1_R1105_U244 , P1_R1105_U32 , P1_R1105_U139 );
nand NAND2_11794 ( P1_R1105_U141 , P1_R1105_U137 , P1_R1105_U32 );
nand NAND2_11795 ( P1_R1105_U142 , P1_REG2_REG_5_ , P1_U3472 );
nand NAND3_11796 ( P1_R1105_U143 , P1_R1105_U142 , P1_R1105_U4 , P1_R1105_U141 );
or OR2_11797 ( P1_R1105_U144 , P1_U3469 , P1_REG2_REG_4_ );
nand NAND2_11798 ( P1_R1105_U145 , P1_R1105_U100 , P1_R1105_U97 );
not NOT1_11799 ( P1_R1105_U146 , P1_R1105_U82 );
nand NAND2_11800 ( P1_R1105_U147 , P1_U3466 , P1_REG2_REG_3_ );
nand NAND4_11801 ( P1_R1105_U148 , P1_R1105_U41 , P1_R1105_U40 , P1_R1105_U257 , P1_R1105_U256 );
nand NAND2_11802 ( P1_R1105_U149 , P1_R1105_U41 , P1_R1105_U40 );
nand NAND2_11803 ( P1_R1105_U150 , P1_U3463 , P1_REG2_REG_2_ );
nand NAND3_11804 ( P1_R1105_U151 , P1_R1105_U150 , P1_R1105_U97 , P1_R1105_U149 );
or OR2_11805 ( P1_R1105_U152 , P1_REG2_REG_1_ , P1_U3460 );
not NOT1_11806 ( P1_R1105_U153 , P1_R1105_U83 );
or OR2_11807 ( P1_R1105_U154 , P1_U3484 , P1_REG2_REG_9_ );
or OR2_11808 ( P1_R1105_U155 , P1_U3487 , P1_REG2_REG_10_ );
nand NAND2_11809 ( P1_R1105_U156 , P1_R1105_U93 , P1_R1105_U7 );
nand NAND2_11810 ( P1_R1105_U157 , P1_U3487 , P1_REG2_REG_10_ );
nand NAND3_11811 ( P1_R1105_U158 , P1_R1105_U157 , P1_R1105_U90 , P1_R1105_U156 );
or OR2_11812 ( P1_R1105_U159 , P1_REG2_REG_10_ , P1_U3487 );
nand NAND3_11813 ( P1_R1105_U160 , P1_R1105_U120 , P1_R1105_U7 , P1_R1105_U81 );
nand NAND2_11814 ( P1_R1105_U161 , P1_R1105_U159 , P1_R1105_U158 );
not NOT1_11815 ( P1_R1105_U162 , P1_R1105_U88 );
or OR2_11816 ( P1_R1105_U163 , P1_U3496 , P1_REG2_REG_13_ );
or OR2_11817 ( P1_R1105_U164 , P1_U3493 , P1_REG2_REG_12_ );
nand NAND2_11818 ( P1_R1105_U165 , P1_R1105_U92 , P1_R1105_U8 );
nand NAND2_11819 ( P1_R1105_U166 , P1_U3496 , P1_REG2_REG_13_ );
nand NAND3_11820 ( P1_R1105_U167 , P1_R1105_U166 , P1_R1105_U91 , P1_R1105_U165 );
or OR2_11821 ( P1_R1105_U168 , P1_REG2_REG_11_ , P1_U3490 );
or OR2_11822 ( P1_R1105_U169 , P1_REG2_REG_13_ , P1_U3496 );
nand NAND3_11823 ( P1_R1105_U170 , P1_R1105_U168 , P1_R1105_U8 , P1_R1105_U88 );
nand NAND2_11824 ( P1_R1105_U171 , P1_R1105_U169 , P1_R1105_U167 );
not NOT1_11825 ( P1_R1105_U172 , P1_R1105_U87 );
or OR2_11826 ( P1_R1105_U173 , P1_REG2_REG_14_ , P1_U3499 );
nand NAND2_11827 ( P1_R1105_U174 , P1_R1105_U173 , P1_R1105_U87 );
nand NAND2_11828 ( P1_R1105_U175 , P1_U3499 , P1_REG2_REG_14_ );
not NOT1_11829 ( P1_R1105_U176 , P1_R1105_U86 );
or OR2_11830 ( P1_R1105_U177 , P1_REG2_REG_15_ , P1_U3502 );
nand NAND2_11831 ( P1_R1105_U178 , P1_R1105_U177 , P1_R1105_U86 );
nand NAND2_11832 ( P1_R1105_U179 , P1_U3502 , P1_REG2_REG_15_ );
not NOT1_11833 ( P1_R1105_U180 , P1_R1105_U66 );
or OR2_11834 ( P1_R1105_U181 , P1_U3508 , P1_REG2_REG_17_ );
or OR2_11835 ( P1_R1105_U182 , P1_U3505 , P1_REG2_REG_16_ );
not NOT1_11836 ( P1_R1105_U183 , P1_R1105_U47 );
nand NAND2_11837 ( P1_R1105_U184 , P1_R1105_U48 , P1_R1105_U47 );
nand NAND2_11838 ( P1_R1105_U185 , P1_U3508 , P1_R1105_U184 );
nand NAND2_11839 ( P1_R1105_U186 , P1_REG2_REG_17_ , P1_R1105_U183 );
nand NAND2_11840 ( P1_R1105_U187 , P1_R1105_U9 , P1_R1105_U66 );
not NOT1_11841 ( P1_R1105_U188 , P1_R1105_U65 );
or OR2_11842 ( P1_R1105_U189 , P1_REG2_REG_18_ , P1_U3511 );
nand NAND2_11843 ( P1_R1105_U190 , P1_R1105_U189 , P1_R1105_U65 );
nand NAND2_11844 ( P1_R1105_U191 , P1_U3511 , P1_REG2_REG_18_ );
nand NAND4_11845 ( P1_R1105_U192 , P1_R1105_U261 , P1_R1105_U260 , P1_R1105_U191 , P1_R1105_U190 );
nand NAND2_11846 ( P1_R1105_U193 , P1_U3511 , P1_REG2_REG_18_ );
nand NAND2_11847 ( P1_R1105_U194 , P1_R1105_U188 , P1_R1105_U193 );
or OR2_11848 ( P1_R1105_U195 , P1_U3511 , P1_REG2_REG_18_ );
nand NAND3_11849 ( P1_R1105_U196 , P1_R1105_U195 , P1_R1105_U264 , P1_R1105_U194 );
or OR2_11850 ( P1_R1105_U197 , P1_REG2_REG_16_ , P1_U3505 );
nand NAND2_11851 ( P1_R1105_U198 , P1_R1105_U197 , P1_R1105_U66 );
nand NAND4_11852 ( P1_R1105_U199 , P1_R1105_U273 , P1_R1105_U272 , P1_R1105_U47 , P1_R1105_U198 );
nand NAND2_11853 ( P1_R1105_U200 , P1_R1105_U180 , P1_R1105_U47 );
nand NAND2_11854 ( P1_R1105_U201 , P1_REG2_REG_17_ , P1_U3508 );
nand NAND3_11855 ( P1_R1105_U202 , P1_R1105_U201 , P1_R1105_U9 , P1_R1105_U200 );
or OR2_11856 ( P1_R1105_U203 , P1_U3505 , P1_REG2_REG_16_ );
nand NAND2_11857 ( P1_R1105_U204 , P1_R1105_U168 , P1_R1105_U88 );
not NOT1_11858 ( P1_R1105_U205 , P1_R1105_U67 );
or OR2_11859 ( P1_R1105_U206 , P1_REG2_REG_12_ , P1_U3493 );
nand NAND2_11860 ( P1_R1105_U207 , P1_R1105_U206 , P1_R1105_U67 );
nand NAND4_11861 ( P1_R1105_U208 , P1_R1105_U294 , P1_R1105_U293 , P1_R1105_U91 , P1_R1105_U207 );
nand NAND2_11862 ( P1_R1105_U209 , P1_R1105_U205 , P1_R1105_U91 );
nand NAND2_11863 ( P1_R1105_U210 , P1_U3496 , P1_REG2_REG_13_ );
nand NAND3_11864 ( P1_R1105_U211 , P1_R1105_U210 , P1_R1105_U8 , P1_R1105_U209 );
or OR2_11865 ( P1_R1105_U212 , P1_U3493 , P1_REG2_REG_12_ );
or OR2_11866 ( P1_R1105_U213 , P1_REG2_REG_9_ , P1_U3484 );
nand NAND2_11867 ( P1_R1105_U214 , P1_R1105_U213 , P1_R1105_U38 );
nand NAND4_11868 ( P1_R1105_U215 , P1_R1105_U306 , P1_R1105_U305 , P1_R1105_U90 , P1_R1105_U214 );
nand NAND2_11869 ( P1_R1105_U216 , P1_R1105_U122 , P1_R1105_U90 );
nand NAND2_11870 ( P1_R1105_U217 , P1_U3487 , P1_REG2_REG_10_ );
nand NAND3_11871 ( P1_R1105_U218 , P1_R1105_U217 , P1_R1105_U7 , P1_R1105_U216 );
nand NAND2_11872 ( P1_R1105_U219 , P1_R1105_U123 , P1_R1105_U90 );
nand NAND2_11873 ( P1_R1105_U220 , P1_R1105_U120 , P1_R1105_U49 );
nand NAND2_11874 ( P1_R1105_U221 , P1_R1105_U130 , P1_R1105_U20 );
nand NAND2_11875 ( P1_R1105_U222 , P1_R1105_U144 , P1_R1105_U32 );
nand NAND2_11876 ( P1_R1105_U223 , P1_R1105_U147 , P1_R1105_U96 );
nand NAND2_11877 ( P1_R1105_U224 , P1_R1105_U203 , P1_R1105_U47 );
nand NAND2_11878 ( P1_R1105_U225 , P1_R1105_U212 , P1_R1105_U91 );
nand NAND2_11879 ( P1_R1105_U226 , P1_R1105_U168 , P1_R1105_U56 );
nand NAND2_11880 ( P1_R1105_U227 , P1_U3484 , P1_R1105_U37 );
nand NAND2_11881 ( P1_R1105_U228 , P1_REG2_REG_9_ , P1_R1105_U36 );
nand NAND2_11882 ( P1_R1105_U229 , P1_R1105_U228 , P1_R1105_U227 );
nand NAND2_11883 ( P1_R1105_U230 , P1_R1105_U219 , P1_R1105_U38 );
nand NAND2_11884 ( P1_R1105_U231 , P1_R1105_U229 , P1_R1105_U122 );
nand NAND2_11885 ( P1_R1105_U232 , P1_U3481 , P1_R1105_U34 );
nand NAND2_11886 ( P1_R1105_U233 , P1_REG2_REG_8_ , P1_R1105_U35 );
nand NAND2_11887 ( P1_R1105_U234 , P1_R1105_U233 , P1_R1105_U232 );
nand NAND2_11888 ( P1_R1105_U235 , P1_R1105_U220 , P1_R1105_U81 );
nand NAND2_11889 ( P1_R1105_U236 , P1_R1105_U119 , P1_R1105_U234 );
nand NAND2_11890 ( P1_R1105_U237 , P1_U3478 , P1_R1105_U21 );
nand NAND2_11891 ( P1_R1105_U238 , P1_REG2_REG_7_ , P1_R1105_U19 );
nand NAND2_11892 ( P1_R1105_U239 , P1_U3475 , P1_R1105_U17 );
nand NAND2_11893 ( P1_R1105_U240 , P1_REG2_REG_6_ , P1_R1105_U18 );
nand NAND2_11894 ( P1_R1105_U241 , P1_R1105_U240 , P1_R1105_U239 );
nand NAND2_11895 ( P1_R1105_U242 , P1_R1105_U221 , P1_R1105_U39 );
nand NAND2_11896 ( P1_R1105_U243 , P1_R1105_U241 , P1_R1105_U111 );
nand NAND2_11897 ( P1_R1105_U244 , P1_U3472 , P1_R1105_U33 );
nand NAND2_11898 ( P1_R1105_U245 , P1_REG2_REG_5_ , P1_R1105_U24 );
nand NAND2_11899 ( P1_R1105_U246 , P1_U3469 , P1_R1105_U22 );
nand NAND2_11900 ( P1_R1105_U247 , P1_REG2_REG_4_ , P1_R1105_U23 );
nand NAND2_11901 ( P1_R1105_U248 , P1_R1105_U247 , P1_R1105_U246 );
nand NAND2_11902 ( P1_R1105_U249 , P1_R1105_U222 , P1_R1105_U42 );
nand NAND2_11903 ( P1_R1105_U250 , P1_R1105_U248 , P1_R1105_U137 );
nand NAND2_11904 ( P1_R1105_U251 , P1_U3466 , P1_R1105_U30 );
nand NAND2_11905 ( P1_R1105_U252 , P1_REG2_REG_3_ , P1_R1105_U31 );
nand NAND2_11906 ( P1_R1105_U253 , P1_R1105_U252 , P1_R1105_U251 );
nand NAND2_11907 ( P1_R1105_U254 , P1_R1105_U223 , P1_R1105_U82 );
nand NAND2_11908 ( P1_R1105_U255 , P1_R1105_U146 , P1_R1105_U253 );
nand NAND2_11909 ( P1_R1105_U256 , P1_U3463 , P1_R1105_U25 );
nand NAND2_11910 ( P1_R1105_U257 , P1_REG2_REG_2_ , P1_R1105_U26 );
nand NAND2_11911 ( P1_R1105_U258 , P1_R1105_U98 , P1_R1105_U83 );
nand NAND2_11912 ( P1_R1105_U259 , P1_R1105_U153 , P1_R1105_U29 );
nand NAND2_11913 ( P1_R1105_U260 , P1_U3452 , P1_R1105_U85 );
nand NAND2_11914 ( P1_R1105_U261 , P1_REG2_REG_19_ , P1_R1105_U84 );
nand NAND2_11915 ( P1_R1105_U262 , P1_U3452 , P1_R1105_U85 );
nand NAND2_11916 ( P1_R1105_U263 , P1_REG2_REG_19_ , P1_R1105_U84 );
nand NAND2_11917 ( P1_R1105_U264 , P1_R1105_U263 , P1_R1105_U262 );
nand NAND2_11918 ( P1_R1105_U265 , P1_U3511 , P1_R1105_U63 );
nand NAND2_11919 ( P1_R1105_U266 , P1_REG2_REG_18_ , P1_R1105_U64 );
nand NAND2_11920 ( P1_R1105_U267 , P1_U3511 , P1_R1105_U63 );
nand NAND2_11921 ( P1_R1105_U268 , P1_REG2_REG_18_ , P1_R1105_U64 );
nand NAND2_11922 ( P1_R1105_U269 , P1_R1105_U268 , P1_R1105_U267 );
nand NAND3_11923 ( P1_R1105_U270 , P1_R1105_U266 , P1_R1105_U265 , P1_R1105_U65 );
nand NAND2_11924 ( P1_R1105_U271 , P1_R1105_U269 , P1_R1105_U188 );
nand NAND2_11925 ( P1_R1105_U272 , P1_U3508 , P1_R1105_U48 );
nand NAND2_11926 ( P1_R1105_U273 , P1_REG2_REG_17_ , P1_R1105_U46 );
nand NAND2_11927 ( P1_R1105_U274 , P1_U3505 , P1_R1105_U44 );
nand NAND2_11928 ( P1_R1105_U275 , P1_REG2_REG_16_ , P1_R1105_U45 );
nand NAND2_11929 ( P1_R1105_U276 , P1_R1105_U275 , P1_R1105_U274 );
nand NAND2_11930 ( P1_R1105_U277 , P1_R1105_U224 , P1_R1105_U66 );
nand NAND2_11931 ( P1_R1105_U278 , P1_R1105_U276 , P1_R1105_U180 );
nand NAND2_11932 ( P1_R1105_U279 , P1_U3502 , P1_R1105_U61 );
nand NAND2_11933 ( P1_R1105_U280 , P1_REG2_REG_15_ , P1_R1105_U62 );
nand NAND2_11934 ( P1_R1105_U281 , P1_U3502 , P1_R1105_U61 );
nand NAND2_11935 ( P1_R1105_U282 , P1_REG2_REG_15_ , P1_R1105_U62 );
nand NAND2_11936 ( P1_R1105_U283 , P1_R1105_U282 , P1_R1105_U281 );
nand NAND3_11937 ( P1_R1105_U284 , P1_R1105_U280 , P1_R1105_U279 , P1_R1105_U86 );
nand NAND2_11938 ( P1_R1105_U285 , P1_R1105_U176 , P1_R1105_U283 );
nand NAND2_11939 ( P1_R1105_U286 , P1_U3499 , P1_R1105_U59 );
nand NAND2_11940 ( P1_R1105_U287 , P1_REG2_REG_14_ , P1_R1105_U60 );
nand NAND2_11941 ( P1_R1105_U288 , P1_U3499 , P1_R1105_U59 );
nand NAND2_11942 ( P1_R1105_U289 , P1_REG2_REG_14_ , P1_R1105_U60 );
nand NAND2_11943 ( P1_R1105_U290 , P1_R1105_U289 , P1_R1105_U288 );
nand NAND3_11944 ( P1_R1105_U291 , P1_R1105_U287 , P1_R1105_U286 , P1_R1105_U87 );
nand NAND2_11945 ( P1_R1105_U292 , P1_R1105_U172 , P1_R1105_U290 );
nand NAND2_11946 ( P1_R1105_U293 , P1_U3496 , P1_R1105_U57 );
nand NAND2_11947 ( P1_R1105_U294 , P1_REG2_REG_13_ , P1_R1105_U58 );
nand NAND2_11948 ( P1_R1105_U295 , P1_U3493 , P1_R1105_U52 );
nand NAND2_11949 ( P1_R1105_U296 , P1_REG2_REG_12_ , P1_R1105_U53 );
nand NAND2_11950 ( P1_R1105_U297 , P1_R1105_U296 , P1_R1105_U295 );
nand NAND2_11951 ( P1_R1105_U298 , P1_R1105_U225 , P1_R1105_U67 );
nand NAND2_11952 ( P1_R1105_U299 , P1_R1105_U297 , P1_R1105_U205 );
nand NAND2_11953 ( P1_R1105_U300 , P1_U3490 , P1_R1105_U54 );
nand NAND2_11954 ( P1_R1105_U301 , P1_REG2_REG_11_ , P1_R1105_U55 );
nand NAND2_11955 ( P1_R1105_U302 , P1_R1105_U301 , P1_R1105_U300 );
nand NAND2_11956 ( P1_R1105_U303 , P1_R1105_U226 , P1_R1105_U88 );
nand NAND2_11957 ( P1_R1105_U304 , P1_R1105_U162 , P1_R1105_U302 );
nand NAND2_11958 ( P1_R1105_U305 , P1_U3487 , P1_R1105_U50 );
nand NAND2_11959 ( P1_R1105_U306 , P1_REG2_REG_10_ , P1_R1105_U51 );
nand NAND2_11960 ( P1_R1105_U307 , P1_U3454 , P1_R1105_U27 );
nand NAND2_11961 ( P1_R1105_U308 , P1_REG2_REG_0_ , P1_R1105_U28 );
and AND2_11962 ( P1_SUB_88_U6 , P1_SUB_88_U227 , P1_SUB_88_U38 );
and AND2_11963 ( P1_SUB_88_U7 , P1_SUB_88_U225 , P1_SUB_88_U192 );
and AND2_11964 ( P1_SUB_88_U8 , P1_SUB_88_U224 , P1_SUB_88_U35 );
and AND2_11965 ( P1_SUB_88_U9 , P1_SUB_88_U223 , P1_SUB_88_U36 );
and AND2_11966 ( P1_SUB_88_U10 , P1_SUB_88_U221 , P1_SUB_88_U195 );
and AND2_11967 ( P1_SUB_88_U11 , P1_SUB_88_U220 , P1_SUB_88_U34 );
and AND2_11968 ( P1_SUB_88_U12 , P1_SUB_88_U219 , P1_SUB_88_U197 );
and AND2_11969 ( P1_SUB_88_U13 , P1_SUB_88_U217 , P1_SUB_88_U198 );
and AND2_11970 ( P1_SUB_88_U14 , P1_SUB_88_U216 , P1_SUB_88_U172 );
and AND2_11971 ( P1_SUB_88_U15 , P1_SUB_88_U215 , P1_SUB_88_U200 );
and AND2_11972 ( P1_SUB_88_U16 , P1_SUB_88_U213 , P1_SUB_88_U201 );
and AND2_11973 ( P1_SUB_88_U17 , P1_SUB_88_U212 , P1_SUB_88_U169 );
and AND2_11974 ( P1_SUB_88_U18 , P1_SUB_88_U211 , P1_SUB_88_U167 );
and AND2_11975 ( P1_SUB_88_U19 , P1_SUB_88_U209 , P1_SUB_88_U204 );
and AND2_11976 ( P1_SUB_88_U20 , P1_SUB_88_U208 , P1_SUB_88_U33 );
and AND2_11977 ( P1_SUB_88_U21 , P1_SUB_88_U207 , P1_SUB_88_U27 );
and AND2_11978 ( P1_SUB_88_U22 , P1_SUB_88_U190 , P1_SUB_88_U180 );
and AND2_11979 ( P1_SUB_88_U23 , P1_SUB_88_U189 , P1_SUB_88_U29 );
and AND2_11980 ( P1_SUB_88_U24 , P1_SUB_88_U188 , P1_SUB_88_U30 );
and AND2_11981 ( P1_SUB_88_U25 , P1_SUB_88_U186 , P1_SUB_88_U183 );
and AND2_11982 ( P1_SUB_88_U26 , P1_SUB_88_U185 , P1_SUB_88_U28 );
or OR3_11983 ( P1_SUB_88_U27 , P1_IR_REG_1_ , P1_IR_REG_0_ , P1_IR_REG_2_ );
nand NAND3_11984 ( P1_SUB_88_U28 , P1_SUB_88_U44 , P1_SUB_88_U230 , P1_SUB_88_U43 );
nand NAND2_11985 ( P1_SUB_88_U29 , P1_SUB_88_U45 , P1_SUB_88_U230 );
nand NAND2_11986 ( P1_SUB_88_U30 , P1_SUB_88_U46 , P1_SUB_88_U181 );
not NOT1_11987 ( P1_SUB_88_U31 , P1_IR_REG_7_ );
not NOT1_11988 ( P1_SUB_88_U32 , P1_IR_REG_3_ );
nand NAND2_11989 ( P1_SUB_88_U33 , P1_SUB_88_U56 , P1_SUB_88_U51 );
nand NAND4_11990 ( P1_SUB_88_U34 , P1_SUB_88_U130 , P1_SUB_88_U129 , P1_SUB_88_U128 , P1_SUB_88_U127 );
nand NAND2_11991 ( P1_SUB_88_U35 , P1_SUB_88_U156 , P1_SUB_88_U184 );
nand NAND2_11992 ( P1_SUB_88_U36 , P1_SUB_88_U157 , P1_SUB_88_U193 );
not NOT1_11993 ( P1_SUB_88_U37 , P1_IR_REG_15_ );
nand NAND2_11994 ( P1_SUB_88_U38 , P1_SUB_88_U158 , P1_SUB_88_U184 );
not NOT1_11995 ( P1_SUB_88_U39 , P1_IR_REG_11_ );
nand NAND2_11996 ( P1_SUB_88_U40 , P1_SUB_88_U247 , P1_SUB_88_U246 );
nand NAND2_11997 ( P1_SUB_88_U41 , P1_SUB_88_U237 , P1_SUB_88_U236 );
nand NAND2_11998 ( P1_SUB_88_U42 , P1_SUB_88_U241 , P1_SUB_88_U240 );
nor nor_11999 ( P1_SUB_88_U43 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_12000 ( P1_SUB_88_U44 , P1_IR_REG_7_ , P1_IR_REG_8_ );
nor nor_12001 ( P1_SUB_88_U45 , P1_IR_REG_3_ , P1_IR_REG_4_ );
nor nor_12002 ( P1_SUB_88_U46 , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_12003 ( P1_SUB_88_U47 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_12004 ( P1_SUB_88_U48 , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_12005 ( P1_SUB_88_U49 , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_12006 ( P1_SUB_88_U50 , P1_IR_REG_22_ , P1_IR_REG_20_ , P1_IR_REG_21_ );
and AND4_12007 ( P1_SUB_88_U51 , P1_SUB_88_U50 , P1_SUB_88_U49 , P1_SUB_88_U48 , P1_SUB_88_U47 );
nor nor_12008 ( P1_SUB_88_U52 , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ );
nor nor_12009 ( P1_SUB_88_U53 , P1_IR_REG_27_ , P1_IR_REG_28_ , P1_IR_REG_29_ , P1_IR_REG_2_ );
nor nor_12010 ( P1_SUB_88_U54 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_12011 ( P1_SUB_88_U55 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_12012 ( P1_SUB_88_U56 , P1_SUB_88_U55 , P1_SUB_88_U54 , P1_SUB_88_U53 , P1_SUB_88_U52 );
nor nor_12013 ( P1_SUB_88_U57 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_12014 ( P1_SUB_88_U58 , P1_IR_REG_14_ , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_12015 ( P1_SUB_88_U59 , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_12016 ( P1_SUB_88_U60 , P1_IR_REG_22_ , P1_IR_REG_20_ , P1_IR_REG_21_ );
and AND4_12017 ( P1_SUB_88_U61 , P1_SUB_88_U60 , P1_SUB_88_U59 , P1_SUB_88_U58 , P1_SUB_88_U57 );
nor nor_12018 ( P1_SUB_88_U62 , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ , P1_IR_REG_26_ );
nor nor_12019 ( P1_SUB_88_U63 , P1_IR_REG_2_ , P1_IR_REG_27_ , P1_IR_REG_28_ );
nor nor_12020 ( P1_SUB_88_U64 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_12021 ( P1_SUB_88_U65 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_12022 ( P1_SUB_88_U66 , P1_SUB_88_U65 , P1_SUB_88_U64 , P1_SUB_88_U63 , P1_SUB_88_U62 );
nor nor_12023 ( P1_SUB_88_U67 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_12024 ( P1_SUB_88_U68 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_12025 ( P1_SUB_88_U69 , P1_IR_REG_17_ , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
nor nor_12026 ( P1_SUB_88_U70 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
and AND4_12027 ( P1_SUB_88_U71 , P1_SUB_88_U70 , P1_SUB_88_U69 , P1_SUB_88_U68 , P1_SUB_88_U67 );
nor nor_12028 ( P1_SUB_88_U72 , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ );
nor nor_12029 ( P1_SUB_88_U73 , P1_IR_REG_2_ , P1_IR_REG_26_ , P1_IR_REG_27_ );
nor nor_12030 ( P1_SUB_88_U74 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_12031 ( P1_SUB_88_U75 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_12032 ( P1_SUB_88_U76 , P1_SUB_88_U75 , P1_SUB_88_U74 , P1_SUB_88_U73 , P1_SUB_88_U72 );
nor nor_12033 ( P1_SUB_88_U77 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_12034 ( P1_SUB_88_U78 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_12035 ( P1_SUB_88_U79 , P1_IR_REG_17_ , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
nor nor_12036 ( P1_SUB_88_U80 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
and AND4_12037 ( P1_SUB_88_U81 , P1_SUB_88_U80 , P1_SUB_88_U79 , P1_SUB_88_U78 , P1_SUB_88_U77 );
nor nor_12038 ( P1_SUB_88_U82 , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ );
nor nor_12039 ( P1_SUB_88_U83 , P1_IR_REG_3_ , P1_IR_REG_26_ , P1_IR_REG_2_ );
nor nor_12040 ( P1_SUB_88_U84 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_12041 ( P1_SUB_88_U85 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_12042 ( P1_SUB_88_U86 , P1_SUB_88_U85 , P1_SUB_88_U84 , P1_SUB_88_U83 , P1_SUB_88_U82 );
nor nor_12043 ( P1_SUB_88_U87 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_12044 ( P1_SUB_88_U88 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_12045 ( P1_SUB_88_U89 , P1_IR_REG_17_ , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
nor nor_12046 ( P1_SUB_88_U90 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
and AND4_12047 ( P1_SUB_88_U91 , P1_SUB_88_U90 , P1_SUB_88_U89 , P1_SUB_88_U88 , P1_SUB_88_U87 );
nor nor_12048 ( P1_SUB_88_U92 , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ , P1_IR_REG_25_ );
nor nor_12049 ( P1_SUB_88_U93 , P1_IR_REG_3_ , P1_IR_REG_26_ , P1_IR_REG_2_ );
nor nor_12050 ( P1_SUB_88_U94 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_12051 ( P1_SUB_88_U95 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_12052 ( P1_SUB_88_U96 , P1_SUB_88_U95 , P1_SUB_88_U94 , P1_SUB_88_U93 , P1_SUB_88_U92 );
nor nor_12053 ( P1_SUB_88_U97 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_12054 ( P1_SUB_88_U98 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_12055 ( P1_SUB_88_U99 , P1_IR_REG_19_ , P1_IR_REG_17_ , P1_IR_REG_18_ );
nor nor_12056 ( P1_SUB_88_U100 , P1_IR_REG_20_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
and AND4_12057 ( P1_SUB_88_U101 , P1_SUB_88_U100 , P1_SUB_88_U99 , P1_SUB_88_U98 , P1_SUB_88_U97 );
nor nor_12058 ( P1_SUB_88_U102 , P1_IR_REG_21_ , P1_IR_REG_22_ , P1_IR_REG_23_ , P1_IR_REG_24_ );
nor nor_12059 ( P1_SUB_88_U103 , P1_IR_REG_3_ , P1_IR_REG_25_ , P1_IR_REG_2_ );
nor nor_12060 ( P1_SUB_88_U104 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_12061 ( P1_SUB_88_U105 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_12062 ( P1_SUB_88_U106 , P1_SUB_88_U105 , P1_SUB_88_U104 , P1_SUB_88_U103 , P1_SUB_88_U102 );
nor nor_12063 ( P1_SUB_88_U107 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_13_ );
nor nor_12064 ( P1_SUB_88_U108 , P1_IR_REG_16_ , P1_IR_REG_14_ , P1_IR_REG_15_ );
nor nor_12065 ( P1_SUB_88_U109 , P1_IR_REG_19_ , P1_IR_REG_17_ , P1_IR_REG_18_ );
nor nor_12066 ( P1_SUB_88_U110 , P1_IR_REG_20_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
and AND4_12067 ( P1_SUB_88_U111 , P1_SUB_88_U110 , P1_SUB_88_U109 , P1_SUB_88_U108 , P1_SUB_88_U107 );
nor nor_12068 ( P1_SUB_88_U112 , P1_IR_REG_23_ , P1_IR_REG_21_ , P1_IR_REG_22_ );
nor nor_12069 ( P1_SUB_88_U113 , P1_IR_REG_3_ , P1_IR_REG_24_ , P1_IR_REG_2_ );
nor nor_12070 ( P1_SUB_88_U114 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_12071 ( P1_SUB_88_U115 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_12072 ( P1_SUB_88_U116 , P1_SUB_88_U115 , P1_SUB_88_U114 , P1_SUB_88_U113 , P1_SUB_88_U112 );
nor nor_12073 ( P1_SUB_88_U117 , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_12074 ( P1_SUB_88_U118 , P1_IR_REG_15_ , P1_IR_REG_13_ , P1_IR_REG_14_ );
nor nor_12075 ( P1_SUB_88_U119 , P1_IR_REG_18_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_12076 ( P1_SUB_88_U120 , P1_IR_REG_0_ , P1_IR_REG_19_ , P1_IR_REG_1_ );
and AND4_12077 ( P1_SUB_88_U121 , P1_SUB_88_U120 , P1_SUB_88_U119 , P1_SUB_88_U118 , P1_SUB_88_U117 );
nor nor_12078 ( P1_SUB_88_U122 , P1_IR_REG_22_ , P1_IR_REG_20_ , P1_IR_REG_21_ );
nor nor_12079 ( P1_SUB_88_U123 , P1_IR_REG_3_ , P1_IR_REG_23_ , P1_IR_REG_2_ );
nor nor_12080 ( P1_SUB_88_U124 , P1_IR_REG_6_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_12081 ( P1_SUB_88_U125 , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_8_ );
and AND4_12082 ( P1_SUB_88_U126 , P1_SUB_88_U125 , P1_SUB_88_U124 , P1_SUB_88_U123 , P1_SUB_88_U122 );
nor nor_12083 ( P1_SUB_88_U127 , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_12084 ( P1_SUB_88_U128 , P1_IR_REG_15_ , P1_IR_REG_16_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_12085 ( P1_SUB_88_U129 , P1_IR_REG_2_ , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_5_ );
nor nor_12086 ( P1_SUB_88_U130 , P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ );
nor nor_12087 ( P1_SUB_88_U131 , P1_IR_REG_17_ , P1_IR_REG_18_ );
nor nor_12088 ( P1_SUB_88_U132 , P1_IR_REG_19_ , P1_IR_REG_20_ );
nor nor_12089 ( P1_SUB_88_U133 , P1_IR_REG_21_ , P1_IR_REG_22_ );
and AND3_12090 ( P1_SUB_88_U134 , P1_SUB_88_U132 , P1_SUB_88_U131 , P1_SUB_88_U133 );
nor nor_12091 ( P1_SUB_88_U135 , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_12092 ( P1_SUB_88_U136 , P1_IR_REG_15_ , P1_IR_REG_13_ , P1_IR_REG_14_ );
and AND2_12093 ( P1_SUB_88_U137 , P1_SUB_88_U136 , P1_SUB_88_U135 );
nor nor_12094 ( P1_SUB_88_U138 , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_18_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_12095 ( P1_SUB_88_U139 , P1_IR_REG_21_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
nor nor_12096 ( P1_SUB_88_U140 , P1_IR_REG_4_ , P1_IR_REG_2_ , P1_IR_REG_3_ );
and AND2_12097 ( P1_SUB_88_U141 , P1_SUB_88_U140 , P1_SUB_88_U139 );
nor nor_12098 ( P1_SUB_88_U142 , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_12099 ( P1_SUB_88_U143 , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_12100 ( P1_SUB_88_U144 , P1_IR_REG_15_ , P1_IR_REG_13_ , P1_IR_REG_14_ );
nor nor_12101 ( P1_SUB_88_U145 , P1_IR_REG_19_ , P1_IR_REG_1_ , P1_IR_REG_18_ , P1_IR_REG_16_ , P1_IR_REG_17_ );
nor nor_12102 ( P1_SUB_88_U146 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_2_ , P1_IR_REG_0_ , P1_IR_REG_20_ );
nor nor_12103 ( P1_SUB_88_U147 , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_12104 ( P1_SUB_88_U148 , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_12105 ( P1_SUB_88_U149 , P1_IR_REG_18_ , P1_IR_REG_19_ , P1_IR_REG_17_ , P1_IR_REG_15_ , P1_IR_REG_16_ );
nor nor_12106 ( P1_SUB_88_U150 , P1_IR_REG_3_ , P1_IR_REG_4_ , P1_IR_REG_2_ , P1_IR_REG_1_ , P1_IR_REG_0_ );
nor nor_12107 ( P1_SUB_88_U151 , P1_IR_REG_8_ , P1_IR_REG_9_ , P1_IR_REG_7_ , P1_IR_REG_5_ , P1_IR_REG_6_ );
nor nor_12108 ( P1_SUB_88_U152 , P1_IR_REG_13_ , P1_IR_REG_14_ , P1_IR_REG_12_ , P1_IR_REG_10_ , P1_IR_REG_11_ );
nor nor_12109 ( P1_SUB_88_U153 , P1_IR_REG_18_ , P1_IR_REG_1_ , P1_IR_REG_17_ , P1_IR_REG_15_ , P1_IR_REG_16_ );
nor nor_12110 ( P1_SUB_88_U154 , P1_IR_REG_4_ , P1_IR_REG_5_ , P1_IR_REG_3_ , P1_IR_REG_0_ , P1_IR_REG_2_ );
nor nor_12111 ( P1_SUB_88_U155 , P1_IR_REG_6_ , P1_IR_REG_7_ , P1_IR_REG_8_ , P1_IR_REG_9_ );
nor nor_12112 ( P1_SUB_88_U156 , P1_IR_REG_10_ , P1_IR_REG_11_ , P1_IR_REG_12_ , P1_IR_REG_9_ );
nor nor_12113 ( P1_SUB_88_U157 , P1_IR_REG_13_ , P1_IR_REG_14_ );
nor nor_12114 ( P1_SUB_88_U158 , P1_IR_REG_10_ , P1_IR_REG_9_ );
not NOT1_12115 ( P1_SUB_88_U159 , P1_IR_REG_9_ );
and AND2_12116 ( P1_SUB_88_U160 , P1_SUB_88_U233 , P1_SUB_88_U232 );
not NOT1_12117 ( P1_SUB_88_U161 , P1_IR_REG_5_ );
and AND2_12118 ( P1_SUB_88_U162 , P1_SUB_88_U235 , P1_SUB_88_U234 );
not NOT1_12119 ( P1_SUB_88_U163 , P1_IR_REG_31_ );
not NOT1_12120 ( P1_SUB_88_U164 , P1_IR_REG_30_ );
and AND2_12121 ( P1_SUB_88_U165 , P1_SUB_88_U239 , P1_SUB_88_U238 );
not NOT1_12122 ( P1_SUB_88_U166 , P1_IR_REG_27_ );
nand NAND2_12123 ( P1_SUB_88_U167 , P1_SUB_88_U96 , P1_SUB_88_U91 );
not NOT1_12124 ( P1_SUB_88_U168 , P1_IR_REG_25_ );
nand NAND2_12125 ( P1_SUB_88_U169 , P1_SUB_88_U116 , P1_SUB_88_U111 );
and AND2_12126 ( P1_SUB_88_U170 , P1_SUB_88_U243 , P1_SUB_88_U242 );
not NOT1_12127 ( P1_SUB_88_U171 , P1_IR_REG_21_ );
nand NAND5_12128 ( P1_SUB_88_U172 , P1_SUB_88_U144 , P1_SUB_88_U143 , P1_SUB_88_U145 , P1_SUB_88_U147 , P1_SUB_88_U146 );
and AND2_12129 ( P1_SUB_88_U173 , P1_SUB_88_U245 , P1_SUB_88_U244 );
not NOT1_12130 ( P1_SUB_88_U174 , P1_IR_REG_1_ );
not NOT1_12131 ( P1_SUB_88_U175 , P1_IR_REG_0_ );
not NOT1_12132 ( P1_SUB_88_U176 , P1_IR_REG_17_ );
and AND2_12133 ( P1_SUB_88_U177 , P1_SUB_88_U249 , P1_SUB_88_U248 );
not NOT1_12134 ( P1_SUB_88_U178 , P1_IR_REG_13_ );
and AND2_12135 ( P1_SUB_88_U179 , P1_SUB_88_U251 , P1_SUB_88_U250 );
nand NAND2_12136 ( P1_SUB_88_U180 , P1_SUB_88_U230 , P1_SUB_88_U32 );
not NOT1_12137 ( P1_SUB_88_U181 , P1_SUB_88_U29 );
not NOT1_12138 ( P1_SUB_88_U182 , P1_SUB_88_U30 );
nand NAND2_12139 ( P1_SUB_88_U183 , P1_SUB_88_U182 , P1_SUB_88_U31 );
not NOT1_12140 ( P1_SUB_88_U184 , P1_SUB_88_U28 );
nand NAND2_12141 ( P1_SUB_88_U185 , P1_IR_REG_8_ , P1_SUB_88_U183 );
nand NAND2_12142 ( P1_SUB_88_U186 , P1_IR_REG_7_ , P1_SUB_88_U30 );
nand NAND2_12143 ( P1_SUB_88_U187 , P1_SUB_88_U181 , P1_SUB_88_U161 );
nand NAND2_12144 ( P1_SUB_88_U188 , P1_IR_REG_6_ , P1_SUB_88_U187 );
nand NAND2_12145 ( P1_SUB_88_U189 , P1_IR_REG_4_ , P1_SUB_88_U180 );
nand NAND2_12146 ( P1_SUB_88_U190 , P1_IR_REG_3_ , P1_SUB_88_U27 );
not NOT1_12147 ( P1_SUB_88_U191 , P1_SUB_88_U38 );
nand NAND2_12148 ( P1_SUB_88_U192 , P1_SUB_88_U191 , P1_SUB_88_U39 );
not NOT1_12149 ( P1_SUB_88_U193 , P1_SUB_88_U35 );
not NOT1_12150 ( P1_SUB_88_U194 , P1_SUB_88_U36 );
nand NAND2_12151 ( P1_SUB_88_U195 , P1_SUB_88_U194 , P1_SUB_88_U37 );
not NOT1_12152 ( P1_SUB_88_U196 , P1_SUB_88_U34 );
nand NAND4_12153 ( P1_SUB_88_U197 , P1_SUB_88_U155 , P1_SUB_88_U154 , P1_SUB_88_U153 , P1_SUB_88_U152 );
nand NAND4_12154 ( P1_SUB_88_U198 , P1_SUB_88_U151 , P1_SUB_88_U150 , P1_SUB_88_U149 , P1_SUB_88_U148 );
not NOT1_12155 ( P1_SUB_88_U199 , P1_SUB_88_U172 );
nand NAND2_12156 ( P1_SUB_88_U200 , P1_SUB_88_U134 , P1_SUB_88_U196 );
nand NAND2_12157 ( P1_SUB_88_U201 , P1_SUB_88_U126 , P1_SUB_88_U121 );
not NOT1_12158 ( P1_SUB_88_U202 , P1_SUB_88_U169 );
not NOT1_12159 ( P1_SUB_88_U203 , P1_SUB_88_U167 );
nand NAND2_12160 ( P1_SUB_88_U204 , P1_SUB_88_U66 , P1_SUB_88_U61 );
not NOT1_12161 ( P1_SUB_88_U205 , P1_SUB_88_U33 );
or OR2_12162 ( P1_SUB_88_U206 , P1_IR_REG_1_ , P1_IR_REG_0_ );
nand NAND2_12163 ( P1_SUB_88_U207 , P1_IR_REG_2_ , P1_SUB_88_U206 );
nand NAND2_12164 ( P1_SUB_88_U208 , P1_IR_REG_29_ , P1_SUB_88_U204 );
nand NAND2_12165 ( P1_SUB_88_U209 , P1_IR_REG_28_ , P1_SUB_88_U229 );
nand NAND2_12166 ( P1_SUB_88_U210 , P1_SUB_88_U106 , P1_SUB_88_U101 );
nand NAND2_12167 ( P1_SUB_88_U211 , P1_IR_REG_26_ , P1_SUB_88_U210 );
nand NAND2_12168 ( P1_SUB_88_U212 , P1_IR_REG_24_ , P1_SUB_88_U201 );
nand NAND2_12169 ( P1_SUB_88_U213 , P1_IR_REG_23_ , P1_SUB_88_U200 );
nand NAND4_12170 ( P1_SUB_88_U214 , P1_SUB_88_U142 , P1_SUB_88_U141 , P1_SUB_88_U138 , P1_SUB_88_U137 );
nand NAND2_12171 ( P1_SUB_88_U215 , P1_IR_REG_22_ , P1_SUB_88_U214 );
nand NAND2_12172 ( P1_SUB_88_U216 , P1_IR_REG_20_ , P1_SUB_88_U198 );
nand NAND2_12173 ( P1_SUB_88_U217 , P1_IR_REG_19_ , P1_SUB_88_U197 );
nand NAND2_12174 ( P1_SUB_88_U218 , P1_SUB_88_U196 , P1_SUB_88_U176 );
nand NAND2_12175 ( P1_SUB_88_U219 , P1_IR_REG_18_ , P1_SUB_88_U218 );
nand NAND2_12176 ( P1_SUB_88_U220 , P1_IR_REG_16_ , P1_SUB_88_U195 );
nand NAND2_12177 ( P1_SUB_88_U221 , P1_IR_REG_15_ , P1_SUB_88_U36 );
nand NAND2_12178 ( P1_SUB_88_U222 , P1_SUB_88_U193 , P1_SUB_88_U178 );
nand NAND2_12179 ( P1_SUB_88_U223 , P1_IR_REG_14_ , P1_SUB_88_U222 );
nand NAND2_12180 ( P1_SUB_88_U224 , P1_IR_REG_12_ , P1_SUB_88_U192 );
nand NAND2_12181 ( P1_SUB_88_U225 , P1_IR_REG_11_ , P1_SUB_88_U38 );
nand NAND2_12182 ( P1_SUB_88_U226 , P1_SUB_88_U184 , P1_SUB_88_U159 );
nand NAND2_12183 ( P1_SUB_88_U227 , P1_IR_REG_10_ , P1_SUB_88_U226 );
nand NAND2_12184 ( P1_SUB_88_U228 , P1_SUB_88_U205 , P1_SUB_88_U164 );
nand NAND2_12185 ( P1_SUB_88_U229 , P1_SUB_88_U76 , P1_SUB_88_U71 );
not NOT1_12186 ( P1_SUB_88_U230 , P1_SUB_88_U27 );
nand NAND2_12187 ( P1_SUB_88_U231 , P1_SUB_88_U86 , P1_SUB_88_U81 );
nand NAND2_12188 ( P1_SUB_88_U232 , P1_IR_REG_9_ , P1_SUB_88_U28 );
nand NAND2_12189 ( P1_SUB_88_U233 , P1_SUB_88_U184 , P1_SUB_88_U159 );
nand NAND2_12190 ( P1_SUB_88_U234 , P1_IR_REG_5_ , P1_SUB_88_U29 );
nand NAND2_12191 ( P1_SUB_88_U235 , P1_SUB_88_U181 , P1_SUB_88_U161 );
nand NAND2_12192 ( P1_SUB_88_U236 , P1_SUB_88_U228 , P1_SUB_88_U163 );
nand NAND3_12193 ( P1_SUB_88_U237 , P1_SUB_88_U205 , P1_SUB_88_U164 , P1_IR_REG_31_ );
nand NAND2_12194 ( P1_SUB_88_U238 , P1_IR_REG_30_ , P1_SUB_88_U33 );
nand NAND2_12195 ( P1_SUB_88_U239 , P1_SUB_88_U205 , P1_SUB_88_U164 );
nand NAND2_12196 ( P1_SUB_88_U240 , P1_SUB_88_U203 , P1_IR_REG_27_ );
nand NAND2_12197 ( P1_SUB_88_U241 , P1_SUB_88_U231 , P1_SUB_88_U166 );
nand NAND2_12198 ( P1_SUB_88_U242 , P1_IR_REG_25_ , P1_SUB_88_U169 );
nand NAND2_12199 ( P1_SUB_88_U243 , P1_SUB_88_U202 , P1_SUB_88_U168 );
nand NAND2_12200 ( P1_SUB_88_U244 , P1_IR_REG_21_ , P1_SUB_88_U172 );
nand NAND2_12201 ( P1_SUB_88_U245 , P1_SUB_88_U199 , P1_SUB_88_U171 );
nand NAND2_12202 ( P1_SUB_88_U246 , P1_IR_REG_1_ , P1_SUB_88_U175 );
nand NAND2_12203 ( P1_SUB_88_U247 , P1_IR_REG_0_ , P1_SUB_88_U174 );
nand NAND2_12204 ( P1_SUB_88_U248 , P1_IR_REG_17_ , P1_SUB_88_U34 );
nand NAND2_12205 ( P1_SUB_88_U249 , P1_SUB_88_U196 , P1_SUB_88_U176 );
nand NAND2_12206 ( P1_SUB_88_U250 , P1_IR_REG_13_ , P1_SUB_88_U35 );
nand NAND2_12207 ( P1_SUB_88_U251 , P1_SUB_88_U193 , P1_SUB_88_U178 );
not NOT1_12208 ( P1_R1309_U6 , P1_U3059 );
not NOT1_12209 ( P1_R1309_U7 , P1_U3056 );
and AND2_12210 ( P1_R1309_U8 , P1_R1309_U10 , P1_R1309_U9 );
nand NAND2_12211 ( P1_R1309_U9 , P1_U3056 , P1_R1309_U6 );
nand NAND2_12212 ( P1_R1309_U10 , P1_U3059 , P1_R1309_U7 );
and AND2_12213 ( P1_R1282_U6 , P1_R1282_U135 , P1_R1282_U35 );
and AND2_12214 ( P1_R1282_U7 , P1_R1282_U133 , P1_R1282_U36 );
and AND2_12215 ( P1_R1282_U8 , P1_R1282_U132 , P1_R1282_U37 );
and AND2_12216 ( P1_R1282_U9 , P1_R1282_U131 , P1_R1282_U38 );
and AND2_12217 ( P1_R1282_U10 , P1_R1282_U129 , P1_R1282_U39 );
and AND2_12218 ( P1_R1282_U11 , P1_R1282_U128 , P1_R1282_U40 );
and AND2_12219 ( P1_R1282_U12 , P1_R1282_U127 , P1_R1282_U41 );
and AND2_12220 ( P1_R1282_U13 , P1_R1282_U125 , P1_R1282_U42 );
and AND2_12221 ( P1_R1282_U14 , P1_R1282_U123 , P1_R1282_U43 );
and AND2_12222 ( P1_R1282_U15 , P1_R1282_U121 , P1_R1282_U44 );
and AND2_12223 ( P1_R1282_U16 , P1_R1282_U119 , P1_R1282_U45 );
and AND2_12224 ( P1_R1282_U17 , P1_R1282_U117 , P1_R1282_U46 );
and AND2_12225 ( P1_R1282_U18 , P1_R1282_U115 , P1_R1282_U25 );
and AND2_12226 ( P1_R1282_U19 , P1_R1282_U113 , P1_R1282_U67 );
and AND2_12227 ( P1_R1282_U20 , P1_R1282_U98 , P1_R1282_U26 );
and AND2_12228 ( P1_R1282_U21 , P1_R1282_U97 , P1_R1282_U27 );
and AND2_12229 ( P1_R1282_U22 , P1_R1282_U96 , P1_R1282_U28 );
and AND2_12230 ( P1_R1282_U23 , P1_R1282_U94 , P1_R1282_U29 );
and AND2_12231 ( P1_R1282_U24 , P1_R1282_U93 , P1_R1282_U30 );
or OR3_12232 ( P1_R1282_U25 , P1_U3461 , P1_U3456 , P1_U3464 );
nand NAND2_12233 ( P1_R1282_U26 , P1_R1282_U87 , P1_R1282_U34 );
nand NAND2_12234 ( P1_R1282_U27 , P1_R1282_U88 , P1_R1282_U33 );
nand NAND2_12235 ( P1_R1282_U28 , P1_R1282_U57 , P1_R1282_U89 );
nand NAND2_12236 ( P1_R1282_U29 , P1_R1282_U90 , P1_R1282_U32 );
nand NAND2_12237 ( P1_R1282_U30 , P1_R1282_U91 , P1_R1282_U31 );
not NOT1_12238 ( P1_R1282_U31 , P1_U3482 );
not NOT1_12239 ( P1_R1282_U32 , P1_U3479 );
not NOT1_12240 ( P1_R1282_U33 , P1_U3470 );
not NOT1_12241 ( P1_R1282_U34 , P1_U3467 );
nand NAND2_12242 ( P1_R1282_U35 , P1_R1282_U58 , P1_R1282_U92 );
nand NAND2_12243 ( P1_R1282_U36 , P1_R1282_U99 , P1_R1282_U55 );
nand NAND2_12244 ( P1_R1282_U37 , P1_R1282_U100 , P1_R1282_U54 );
nand NAND2_12245 ( P1_R1282_U38 , P1_R1282_U59 , P1_R1282_U101 );
nand NAND2_12246 ( P1_R1282_U39 , P1_R1282_U102 , P1_R1282_U53 );
nand NAND2_12247 ( P1_R1282_U40 , P1_R1282_U103 , P1_R1282_U52 );
nand NAND2_12248 ( P1_R1282_U41 , P1_R1282_U60 , P1_R1282_U104 );
nand NAND2_12249 ( P1_R1282_U42 , P1_R1282_U61 , P1_R1282_U105 );
nand NAND3_12250 ( P1_R1282_U43 , P1_R1282_U106 , P1_R1282_U77 , P1_R1282_U51 );
nand NAND3_12251 ( P1_R1282_U44 , P1_R1282_U107 , P1_R1282_U75 , P1_R1282_U50 );
nand NAND3_12252 ( P1_R1282_U45 , P1_R1282_U108 , P1_R1282_U73 , P1_R1282_U49 );
nand NAND3_12253 ( P1_R1282_U46 , P1_R1282_U109 , P1_R1282_U71 , P1_R1282_U48 );
not NOT1_12254 ( P1_R1282_U47 , P1_U4027 );
not NOT1_12255 ( P1_R1282_U48 , P1_U4017 );
not NOT1_12256 ( P1_R1282_U49 , P1_U4019 );
not NOT1_12257 ( P1_R1282_U50 , P1_U4021 );
not NOT1_12258 ( P1_R1282_U51 , P1_U4023 );
not NOT1_12259 ( P1_R1282_U52 , P1_U3506 );
not NOT1_12260 ( P1_R1282_U53 , P1_U3503 );
not NOT1_12261 ( P1_R1282_U54 , P1_U3494 );
not NOT1_12262 ( P1_R1282_U55 , P1_U3491 );
nand NAND2_12263 ( P1_R1282_U56 , P1_R1282_U153 , P1_R1282_U152 );
nor nor_12264 ( P1_R1282_U57 , P1_U3473 , P1_U3476 );
nor nor_12265 ( P1_R1282_U58 , P1_U3488 , P1_U3485 );
nor nor_12266 ( P1_R1282_U59 , P1_U3497 , P1_U3500 );
nor nor_12267 ( P1_R1282_U60 , P1_U3509 , P1_U3512 );
nor nor_12268 ( P1_R1282_U61 , P1_U3514 , P1_U4025 );
not NOT1_12269 ( P1_R1282_U62 , P1_U3485 );
and AND2_12270 ( P1_R1282_U63 , P1_R1282_U137 , P1_R1282_U136 );
not NOT1_12271 ( P1_R1282_U64 , P1_U3473 );
and AND2_12272 ( P1_R1282_U65 , P1_R1282_U139 , P1_R1282_U138 );
not NOT1_12273 ( P1_R1282_U66 , P1_U4026 );
nand NAND3_12274 ( P1_R1282_U67 , P1_R1282_U110 , P1_R1282_U69 , P1_R1282_U47 );
and AND2_12275 ( P1_R1282_U68 , P1_R1282_U141 , P1_R1282_U140 );
not NOT1_12276 ( P1_R1282_U69 , P1_U4028 );
and AND2_12277 ( P1_R1282_U70 , P1_R1282_U143 , P1_R1282_U142 );
not NOT1_12278 ( P1_R1282_U71 , P1_U4018 );
and AND2_12279 ( P1_R1282_U72 , P1_R1282_U145 , P1_R1282_U144 );
not NOT1_12280 ( P1_R1282_U73 , P1_U4020 );
and AND2_12281 ( P1_R1282_U74 , P1_R1282_U147 , P1_R1282_U146 );
not NOT1_12282 ( P1_R1282_U75 , P1_U4022 );
and AND2_12283 ( P1_R1282_U76 , P1_R1282_U149 , P1_R1282_U148 );
not NOT1_12284 ( P1_R1282_U77 , P1_U4024 );
and AND2_12285 ( P1_R1282_U78 , P1_R1282_U151 , P1_R1282_U150 );
not NOT1_12286 ( P1_R1282_U79 , P1_U3461 );
not NOT1_12287 ( P1_R1282_U80 , P1_U3456 );
not NOT1_12288 ( P1_R1282_U81 , P1_U3514 );
and AND2_12289 ( P1_R1282_U82 , P1_R1282_U155 , P1_R1282_U154 );
not NOT1_12290 ( P1_R1282_U83 , P1_U3509 );
and AND2_12291 ( P1_R1282_U84 , P1_R1282_U157 , P1_R1282_U156 );
not NOT1_12292 ( P1_R1282_U85 , P1_U3497 );
and AND2_12293 ( P1_R1282_U86 , P1_R1282_U159 , P1_R1282_U158 );
not NOT1_12294 ( P1_R1282_U87 , P1_R1282_U25 );
not NOT1_12295 ( P1_R1282_U88 , P1_R1282_U26 );
not NOT1_12296 ( P1_R1282_U89 , P1_R1282_U27 );
not NOT1_12297 ( P1_R1282_U90 , P1_R1282_U28 );
not NOT1_12298 ( P1_R1282_U91 , P1_R1282_U29 );
not NOT1_12299 ( P1_R1282_U92 , P1_R1282_U30 );
nand NAND2_12300 ( P1_R1282_U93 , P1_U3482 , P1_R1282_U29 );
nand NAND2_12301 ( P1_R1282_U94 , P1_U3479 , P1_R1282_U28 );
nand NAND2_12302 ( P1_R1282_U95 , P1_R1282_U89 , P1_R1282_U64 );
nand NAND2_12303 ( P1_R1282_U96 , P1_U3476 , P1_R1282_U95 );
nand NAND2_12304 ( P1_R1282_U97 , P1_U3470 , P1_R1282_U26 );
nand NAND2_12305 ( P1_R1282_U98 , P1_U3467 , P1_R1282_U25 );
not NOT1_12306 ( P1_R1282_U99 , P1_R1282_U35 );
not NOT1_12307 ( P1_R1282_U100 , P1_R1282_U36 );
not NOT1_12308 ( P1_R1282_U101 , P1_R1282_U37 );
not NOT1_12309 ( P1_R1282_U102 , P1_R1282_U38 );
not NOT1_12310 ( P1_R1282_U103 , P1_R1282_U39 );
not NOT1_12311 ( P1_R1282_U104 , P1_R1282_U40 );
not NOT1_12312 ( P1_R1282_U105 , P1_R1282_U41 );
not NOT1_12313 ( P1_R1282_U106 , P1_R1282_U42 );
not NOT1_12314 ( P1_R1282_U107 , P1_R1282_U43 );
not NOT1_12315 ( P1_R1282_U108 , P1_R1282_U44 );
not NOT1_12316 ( P1_R1282_U109 , P1_R1282_U45 );
not NOT1_12317 ( P1_R1282_U110 , P1_R1282_U46 );
not NOT1_12318 ( P1_R1282_U111 , P1_R1282_U67 );
nand NAND2_12319 ( P1_R1282_U112 , P1_R1282_U110 , P1_R1282_U69 );
nand NAND2_12320 ( P1_R1282_U113 , P1_U4027 , P1_R1282_U112 );
or OR2_12321 ( P1_R1282_U114 , P1_U3461 , P1_U3456 );
nand NAND2_12322 ( P1_R1282_U115 , P1_U3464 , P1_R1282_U114 );
nand NAND2_12323 ( P1_R1282_U116 , P1_R1282_U109 , P1_R1282_U71 );
nand NAND2_12324 ( P1_R1282_U117 , P1_U4017 , P1_R1282_U116 );
nand NAND2_12325 ( P1_R1282_U118 , P1_R1282_U108 , P1_R1282_U73 );
nand NAND2_12326 ( P1_R1282_U119 , P1_U4019 , P1_R1282_U118 );
nand NAND2_12327 ( P1_R1282_U120 , P1_R1282_U107 , P1_R1282_U75 );
nand NAND2_12328 ( P1_R1282_U121 , P1_U4021 , P1_R1282_U120 );
nand NAND2_12329 ( P1_R1282_U122 , P1_R1282_U106 , P1_R1282_U77 );
nand NAND2_12330 ( P1_R1282_U123 , P1_U4023 , P1_R1282_U122 );
nand NAND2_12331 ( P1_R1282_U124 , P1_R1282_U105 , P1_R1282_U81 );
nand NAND2_12332 ( P1_R1282_U125 , P1_U4025 , P1_R1282_U124 );
nand NAND2_12333 ( P1_R1282_U126 , P1_R1282_U104 , P1_R1282_U83 );
nand NAND2_12334 ( P1_R1282_U127 , P1_U3512 , P1_R1282_U126 );
nand NAND2_12335 ( P1_R1282_U128 , P1_U3506 , P1_R1282_U39 );
nand NAND2_12336 ( P1_R1282_U129 , P1_U3503 , P1_R1282_U38 );
nand NAND2_12337 ( P1_R1282_U130 , P1_R1282_U101 , P1_R1282_U85 );
nand NAND2_12338 ( P1_R1282_U131 , P1_U3500 , P1_R1282_U130 );
nand NAND2_12339 ( P1_R1282_U132 , P1_U3494 , P1_R1282_U36 );
nand NAND2_12340 ( P1_R1282_U133 , P1_U3491 , P1_R1282_U35 );
nand NAND2_12341 ( P1_R1282_U134 , P1_R1282_U92 , P1_R1282_U62 );
nand NAND2_12342 ( P1_R1282_U135 , P1_U3488 , P1_R1282_U134 );
nand NAND2_12343 ( P1_R1282_U136 , P1_U3485 , P1_R1282_U30 );
nand NAND2_12344 ( P1_R1282_U137 , P1_R1282_U92 , P1_R1282_U62 );
nand NAND2_12345 ( P1_R1282_U138 , P1_U3473 , P1_R1282_U27 );
nand NAND2_12346 ( P1_R1282_U139 , P1_R1282_U89 , P1_R1282_U64 );
nand NAND2_12347 ( P1_R1282_U140 , P1_U4026 , P1_R1282_U67 );
nand NAND2_12348 ( P1_R1282_U141 , P1_R1282_U111 , P1_R1282_U66 );
nand NAND2_12349 ( P1_R1282_U142 , P1_U4028 , P1_R1282_U46 );
nand NAND2_12350 ( P1_R1282_U143 , P1_R1282_U110 , P1_R1282_U69 );
nand NAND2_12351 ( P1_R1282_U144 , P1_U4018 , P1_R1282_U45 );
nand NAND2_12352 ( P1_R1282_U145 , P1_R1282_U109 , P1_R1282_U71 );
nand NAND2_12353 ( P1_R1282_U146 , P1_U4020 , P1_R1282_U44 );
nand NAND2_12354 ( P1_R1282_U147 , P1_R1282_U108 , P1_R1282_U73 );
nand NAND2_12355 ( P1_R1282_U148 , P1_U4022 , P1_R1282_U43 );
nand NAND2_12356 ( P1_R1282_U149 , P1_R1282_U107 , P1_R1282_U75 );
nand NAND2_12357 ( P1_R1282_U150 , P1_U4024 , P1_R1282_U42 );
nand NAND2_12358 ( P1_R1282_U151 , P1_R1282_U106 , P1_R1282_U77 );
nand NAND2_12359 ( P1_R1282_U152 , P1_U3461 , P1_R1282_U80 );
nand NAND2_12360 ( P1_R1282_U153 , P1_U3456 , P1_R1282_U79 );
nand NAND2_12361 ( P1_R1282_U154 , P1_U3514 , P1_R1282_U41 );
nand NAND2_12362 ( P1_R1282_U155 , P1_R1282_U105 , P1_R1282_U81 );
nand NAND2_12363 ( P1_R1282_U156 , P1_U3509 , P1_R1282_U40 );
nand NAND2_12364 ( P1_R1282_U157 , P1_R1282_U104 , P1_R1282_U83 );
nand NAND2_12365 ( P1_R1282_U158 , P1_U3497 , P1_R1282_U37 );
nand NAND2_12366 ( P1_R1282_U159 , P1_R1282_U101 , P1_R1282_U85 );
and AND2_12367 ( P1_R1240_U4 , P1_R1240_U176 , P1_R1240_U175 );
and AND2_12368 ( P1_R1240_U5 , P1_R1240_U177 , P1_R1240_U178 );
and AND2_12369 ( P1_R1240_U6 , P1_R1240_U194 , P1_R1240_U193 );
and AND2_12370 ( P1_R1240_U7 , P1_R1240_U234 , P1_R1240_U233 );
and AND2_12371 ( P1_R1240_U8 , P1_R1240_U243 , P1_R1240_U242 );
and AND2_12372 ( P1_R1240_U9 , P1_R1240_U261 , P1_R1240_U260 );
and AND2_12373 ( P1_R1240_U10 , P1_R1240_U269 , P1_R1240_U268 );
and AND2_12374 ( P1_R1240_U11 , P1_R1240_U348 , P1_R1240_U345 );
and AND2_12375 ( P1_R1240_U12 , P1_R1240_U341 , P1_R1240_U338 );
and AND2_12376 ( P1_R1240_U13 , P1_R1240_U332 , P1_R1240_U329 );
and AND2_12377 ( P1_R1240_U14 , P1_R1240_U323 , P1_R1240_U320 );
and AND2_12378 ( P1_R1240_U15 , P1_R1240_U317 , P1_R1240_U315 );
and AND2_12379 ( P1_R1240_U16 , P1_R1240_U310 , P1_R1240_U307 );
and AND2_12380 ( P1_R1240_U17 , P1_R1240_U232 , P1_R1240_U229 );
and AND2_12381 ( P1_R1240_U18 , P1_R1240_U224 , P1_R1240_U221 );
and AND2_12382 ( P1_R1240_U19 , P1_R1240_U210 , P1_R1240_U207 );
not NOT1_12383 ( P1_R1240_U20 , P1_U3476 );
not NOT1_12384 ( P1_R1240_U21 , P1_U3071 );
not NOT1_12385 ( P1_R1240_U22 , P1_U3070 );
nand NAND2_12386 ( P1_R1240_U23 , P1_U3071 , P1_U3476 );
not NOT1_12387 ( P1_R1240_U24 , P1_U3479 );
not NOT1_12388 ( P1_R1240_U25 , P1_U3470 );
not NOT1_12389 ( P1_R1240_U26 , P1_U3060 );
not NOT1_12390 ( P1_R1240_U27 , P1_U3067 );
not NOT1_12391 ( P1_R1240_U28 , P1_U3464 );
not NOT1_12392 ( P1_R1240_U29 , P1_U3068 );
not NOT1_12393 ( P1_R1240_U30 , P1_U3456 );
not NOT1_12394 ( P1_R1240_U31 , P1_U3077 );
nand NAND2_12395 ( P1_R1240_U32 , P1_U3077 , P1_U3456 );
not NOT1_12396 ( P1_R1240_U33 , P1_U3467 );
not NOT1_12397 ( P1_R1240_U34 , P1_U3064 );
nand NAND2_12398 ( P1_R1240_U35 , P1_U3060 , P1_U3470 );
not NOT1_12399 ( P1_R1240_U36 , P1_U3473 );
not NOT1_12400 ( P1_R1240_U37 , P1_U3482 );
not NOT1_12401 ( P1_R1240_U38 , P1_U3084 );
not NOT1_12402 ( P1_R1240_U39 , P1_U3083 );
not NOT1_12403 ( P1_R1240_U40 , P1_U3485 );
nand NAND2_12404 ( P1_R1240_U41 , P1_R1240_U62 , P1_R1240_U202 );
nand NAND2_12405 ( P1_R1240_U42 , P1_R1240_U118 , P1_R1240_U190 );
nand NAND2_12406 ( P1_R1240_U43 , P1_R1240_U179 , P1_R1240_U180 );
nand NAND2_12407 ( P1_R1240_U44 , P1_U3461 , P1_U3078 );
nand NAND2_12408 ( P1_R1240_U45 , P1_R1240_U122 , P1_R1240_U216 );
nand NAND2_12409 ( P1_R1240_U46 , P1_R1240_U213 , P1_R1240_U212 );
not NOT1_12410 ( P1_R1240_U47 , P1_U4018 );
not NOT1_12411 ( P1_R1240_U48 , P1_U3053 );
not NOT1_12412 ( P1_R1240_U49 , P1_U3057 );
not NOT1_12413 ( P1_R1240_U50 , P1_U4019 );
not NOT1_12414 ( P1_R1240_U51 , P1_U4020 );
not NOT1_12415 ( P1_R1240_U52 , P1_U3058 );
not NOT1_12416 ( P1_R1240_U53 , P1_U4021 );
not NOT1_12417 ( P1_R1240_U54 , P1_U3065 );
not NOT1_12418 ( P1_R1240_U55 , P1_U4024 );
not NOT1_12419 ( P1_R1240_U56 , P1_U3075 );
not NOT1_12420 ( P1_R1240_U57 , P1_U3506 );
not NOT1_12421 ( P1_R1240_U58 , P1_U3073 );
not NOT1_12422 ( P1_R1240_U59 , P1_U3069 );
nand NAND2_12423 ( P1_R1240_U60 , P1_U3073 , P1_U3506 );
not NOT1_12424 ( P1_R1240_U61 , P1_U3509 );
nand NAND2_12425 ( P1_R1240_U62 , P1_U3084 , P1_U3482 );
not NOT1_12426 ( P1_R1240_U63 , P1_U3488 );
not NOT1_12427 ( P1_R1240_U64 , P1_U3062 );
not NOT1_12428 ( P1_R1240_U65 , P1_U3494 );
not NOT1_12429 ( P1_R1240_U66 , P1_U3072 );
not NOT1_12430 ( P1_R1240_U67 , P1_U3491 );
not NOT1_12431 ( P1_R1240_U68 , P1_U3063 );
nand NAND2_12432 ( P1_R1240_U69 , P1_U3063 , P1_U3491 );
not NOT1_12433 ( P1_R1240_U70 , P1_U3497 );
not NOT1_12434 ( P1_R1240_U71 , P1_U3080 );
not NOT1_12435 ( P1_R1240_U72 , P1_U3500 );
not NOT1_12436 ( P1_R1240_U73 , P1_U3079 );
not NOT1_12437 ( P1_R1240_U74 , P1_U3503 );
not NOT1_12438 ( P1_R1240_U75 , P1_U3074 );
not NOT1_12439 ( P1_R1240_U76 , P1_U3512 );
not NOT1_12440 ( P1_R1240_U77 , P1_U3082 );
nand NAND2_12441 ( P1_R1240_U78 , P1_U3082 , P1_U3512 );
not NOT1_12442 ( P1_R1240_U79 , P1_U3514 );
not NOT1_12443 ( P1_R1240_U80 , P1_U3081 );
nand NAND2_12444 ( P1_R1240_U81 , P1_U3081 , P1_U3514 );
not NOT1_12445 ( P1_R1240_U82 , P1_U4025 );
not NOT1_12446 ( P1_R1240_U83 , P1_U4023 );
not NOT1_12447 ( P1_R1240_U84 , P1_U3061 );
not NOT1_12448 ( P1_R1240_U85 , P1_U4022 );
not NOT1_12449 ( P1_R1240_U86 , P1_U3066 );
nand NAND2_12450 ( P1_R1240_U87 , P1_U4019 , P1_U3057 );
not NOT1_12451 ( P1_R1240_U88 , P1_U3054 );
not NOT1_12452 ( P1_R1240_U89 , P1_U4017 );
nand NAND2_12453 ( P1_R1240_U90 , P1_R1240_U303 , P1_R1240_U173 );
not NOT1_12454 ( P1_R1240_U91 , P1_U3076 );
nand NAND2_12455 ( P1_R1240_U92 , P1_R1240_U78 , P1_R1240_U312 );
nand NAND2_12456 ( P1_R1240_U93 , P1_R1240_U258 , P1_R1240_U257 );
nand NAND2_12457 ( P1_R1240_U94 , P1_R1240_U69 , P1_R1240_U334 );
nand NAND2_12458 ( P1_R1240_U95 , P1_R1240_U454 , P1_R1240_U453 );
nand NAND2_12459 ( P1_R1240_U96 , P1_R1240_U501 , P1_R1240_U500 );
nand NAND2_12460 ( P1_R1240_U97 , P1_R1240_U372 , P1_R1240_U371 );
nand NAND2_12461 ( P1_R1240_U98 , P1_R1240_U377 , P1_R1240_U376 );
nand NAND2_12462 ( P1_R1240_U99 , P1_R1240_U384 , P1_R1240_U383 );
nand NAND2_12463 ( P1_R1240_U100 , P1_R1240_U391 , P1_R1240_U390 );
nand NAND2_12464 ( P1_R1240_U101 , P1_R1240_U396 , P1_R1240_U395 );
nand NAND2_12465 ( P1_R1240_U102 , P1_R1240_U405 , P1_R1240_U404 );
nand NAND2_12466 ( P1_R1240_U103 , P1_R1240_U412 , P1_R1240_U411 );
nand NAND2_12467 ( P1_R1240_U104 , P1_R1240_U419 , P1_R1240_U418 );
nand NAND2_12468 ( P1_R1240_U105 , P1_R1240_U426 , P1_R1240_U425 );
nand NAND2_12469 ( P1_R1240_U106 , P1_R1240_U431 , P1_R1240_U430 );
nand NAND2_12470 ( P1_R1240_U107 , P1_R1240_U438 , P1_R1240_U437 );
nand NAND2_12471 ( P1_R1240_U108 , P1_R1240_U445 , P1_R1240_U444 );
nand NAND2_12472 ( P1_R1240_U109 , P1_R1240_U459 , P1_R1240_U458 );
nand NAND2_12473 ( P1_R1240_U110 , P1_R1240_U464 , P1_R1240_U463 );
nand NAND2_12474 ( P1_R1240_U111 , P1_R1240_U471 , P1_R1240_U470 );
nand NAND2_12475 ( P1_R1240_U112 , P1_R1240_U478 , P1_R1240_U477 );
nand NAND2_12476 ( P1_R1240_U113 , P1_R1240_U485 , P1_R1240_U484 );
nand NAND2_12477 ( P1_R1240_U114 , P1_R1240_U492 , P1_R1240_U491 );
nand NAND2_12478 ( P1_R1240_U115 , P1_R1240_U497 , P1_R1240_U496 );
and AND2_12479 ( P1_R1240_U116 , P1_U3464 , P1_U3068 );
and AND2_12480 ( P1_R1240_U117 , P1_R1240_U186 , P1_R1240_U184 );
and AND2_12481 ( P1_R1240_U118 , P1_R1240_U191 , P1_R1240_U189 );
and AND2_12482 ( P1_R1240_U119 , P1_R1240_U198 , P1_R1240_U197 );
and AND3_12483 ( P1_R1240_U120 , P1_R1240_U379 , P1_R1240_U378 , P1_R1240_U23 );
and AND2_12484 ( P1_R1240_U121 , P1_R1240_U209 , P1_R1240_U6 );
and AND2_12485 ( P1_R1240_U122 , P1_R1240_U217 , P1_R1240_U215 );
and AND3_12486 ( P1_R1240_U123 , P1_R1240_U386 , P1_R1240_U385 , P1_R1240_U35 );
and AND2_12487 ( P1_R1240_U124 , P1_R1240_U223 , P1_R1240_U4 );
and AND2_12488 ( P1_R1240_U125 , P1_R1240_U231 , P1_R1240_U178 );
and AND2_12489 ( P1_R1240_U126 , P1_R1240_U201 , P1_R1240_U7 );
and AND2_12490 ( P1_R1240_U127 , P1_R1240_U236 , P1_R1240_U168 );
and AND2_12491 ( P1_R1240_U128 , P1_R1240_U245 , P1_R1240_U169 );
and AND2_12492 ( P1_R1240_U129 , P1_R1240_U265 , P1_R1240_U264 );
and AND2_12493 ( P1_R1240_U130 , P1_R1240_U10 , P1_R1240_U279 );
and AND2_12494 ( P1_R1240_U131 , P1_R1240_U282 , P1_R1240_U277 );
and AND2_12495 ( P1_R1240_U132 , P1_R1240_U298 , P1_R1240_U295 );
and AND2_12496 ( P1_R1240_U133 , P1_R1240_U365 , P1_R1240_U299 );
and AND2_12497 ( P1_R1240_U134 , P1_R1240_U156 , P1_R1240_U275 );
and AND3_12498 ( P1_R1240_U135 , P1_R1240_U466 , P1_R1240_U465 , P1_R1240_U60 );
and AND3_12499 ( P1_R1240_U136 , P1_R1240_U487 , P1_R1240_U486 , P1_R1240_U169 );
and AND2_12500 ( P1_R1240_U137 , P1_R1240_U340 , P1_R1240_U8 );
and AND3_12501 ( P1_R1240_U138 , P1_R1240_U499 , P1_R1240_U498 , P1_R1240_U168 );
and AND2_12502 ( P1_R1240_U139 , P1_R1240_U347 , P1_R1240_U7 );
nand NAND2_12503 ( P1_R1240_U140 , P1_R1240_U119 , P1_R1240_U199 );
nand NAND2_12504 ( P1_R1240_U141 , P1_R1240_U214 , P1_R1240_U226 );
not NOT1_12505 ( P1_R1240_U142 , P1_U3055 );
not NOT1_12506 ( P1_R1240_U143 , P1_U4028 );
and AND2_12507 ( P1_R1240_U144 , P1_R1240_U400 , P1_R1240_U399 );
nand NAND3_12508 ( P1_R1240_U145 , P1_R1240_U301 , P1_R1240_U166 , P1_R1240_U361 );
and AND2_12509 ( P1_R1240_U146 , P1_R1240_U407 , P1_R1240_U406 );
nand NAND3_12510 ( P1_R1240_U147 , P1_R1240_U367 , P1_R1240_U366 , P1_R1240_U133 );
and AND2_12511 ( P1_R1240_U148 , P1_R1240_U414 , P1_R1240_U413 );
nand NAND3_12512 ( P1_R1240_U149 , P1_R1240_U362 , P1_R1240_U296 , P1_R1240_U87 );
and AND2_12513 ( P1_R1240_U150 , P1_R1240_U421 , P1_R1240_U420 );
nand NAND2_12514 ( P1_R1240_U151 , P1_R1240_U290 , P1_R1240_U289 );
and AND2_12515 ( P1_R1240_U152 , P1_R1240_U433 , P1_R1240_U432 );
nand NAND2_12516 ( P1_R1240_U153 , P1_R1240_U286 , P1_R1240_U285 );
and AND2_12517 ( P1_R1240_U154 , P1_R1240_U440 , P1_R1240_U439 );
nand NAND2_12518 ( P1_R1240_U155 , P1_R1240_U131 , P1_R1240_U281 );
and AND2_12519 ( P1_R1240_U156 , P1_R1240_U447 , P1_R1240_U446 );
and AND2_12520 ( P1_R1240_U157 , P1_R1240_U452 , P1_R1240_U451 );
nand NAND2_12521 ( P1_R1240_U158 , P1_R1240_U44 , P1_R1240_U324 );
nand NAND2_12522 ( P1_R1240_U159 , P1_R1240_U129 , P1_R1240_U266 );
and AND2_12523 ( P1_R1240_U160 , P1_R1240_U473 , P1_R1240_U472 );
nand NAND2_12524 ( P1_R1240_U161 , P1_R1240_U254 , P1_R1240_U253 );
and AND2_12525 ( P1_R1240_U162 , P1_R1240_U480 , P1_R1240_U479 );
nand NAND2_12526 ( P1_R1240_U163 , P1_R1240_U250 , P1_R1240_U249 );
nand NAND2_12527 ( P1_R1240_U164 , P1_R1240_U240 , P1_R1240_U239 );
nand NAND2_12528 ( P1_R1240_U165 , P1_R1240_U364 , P1_R1240_U363 );
nand NAND2_12529 ( P1_R1240_U166 , P1_U3054 , P1_R1240_U147 );
not NOT1_12530 ( P1_R1240_U167 , P1_R1240_U35 );
nand NAND2_12531 ( P1_R1240_U168 , P1_U3485 , P1_U3083 );
nand NAND2_12532 ( P1_R1240_U169 , P1_U3072 , P1_U3494 );
nand NAND2_12533 ( P1_R1240_U170 , P1_U3058 , P1_U4020 );
not NOT1_12534 ( P1_R1240_U171 , P1_R1240_U69 );
not NOT1_12535 ( P1_R1240_U172 , P1_R1240_U78 );
nand NAND2_12536 ( P1_R1240_U173 , P1_U3065 , P1_U4021 );
not NOT1_12537 ( P1_R1240_U174 , P1_R1240_U62 );
or OR2_12538 ( P1_R1240_U175 , P1_U3067 , P1_U3473 );
or OR2_12539 ( P1_R1240_U176 , P1_U3060 , P1_U3470 );
or OR2_12540 ( P1_R1240_U177 , P1_U3467 , P1_U3064 );
or OR2_12541 ( P1_R1240_U178 , P1_U3464 , P1_U3068 );
not NOT1_12542 ( P1_R1240_U179 , P1_R1240_U32 );
or OR2_12543 ( P1_R1240_U180 , P1_U3461 , P1_U3078 );
not NOT1_12544 ( P1_R1240_U181 , P1_R1240_U43 );
not NOT1_12545 ( P1_R1240_U182 , P1_R1240_U44 );
nand NAND2_12546 ( P1_R1240_U183 , P1_R1240_U43 , P1_R1240_U44 );
nand NAND2_12547 ( P1_R1240_U184 , P1_R1240_U116 , P1_R1240_U177 );
nand NAND2_12548 ( P1_R1240_U185 , P1_R1240_U5 , P1_R1240_U183 );
nand NAND2_12549 ( P1_R1240_U186 , P1_U3064 , P1_U3467 );
nand NAND2_12550 ( P1_R1240_U187 , P1_R1240_U117 , P1_R1240_U185 );
nand NAND2_12551 ( P1_R1240_U188 , P1_R1240_U36 , P1_R1240_U35 );
nand NAND2_12552 ( P1_R1240_U189 , P1_U3067 , P1_R1240_U188 );
nand NAND2_12553 ( P1_R1240_U190 , P1_R1240_U4 , P1_R1240_U187 );
nand NAND2_12554 ( P1_R1240_U191 , P1_U3473 , P1_R1240_U167 );
not NOT1_12555 ( P1_R1240_U192 , P1_R1240_U42 );
or OR2_12556 ( P1_R1240_U193 , P1_U3070 , P1_U3479 );
or OR2_12557 ( P1_R1240_U194 , P1_U3071 , P1_U3476 );
not NOT1_12558 ( P1_R1240_U195 , P1_R1240_U23 );
nand NAND2_12559 ( P1_R1240_U196 , P1_R1240_U24 , P1_R1240_U23 );
nand NAND2_12560 ( P1_R1240_U197 , P1_U3070 , P1_R1240_U196 );
nand NAND2_12561 ( P1_R1240_U198 , P1_U3479 , P1_R1240_U195 );
nand NAND2_12562 ( P1_R1240_U199 , P1_R1240_U6 , P1_R1240_U42 );
not NOT1_12563 ( P1_R1240_U200 , P1_R1240_U140 );
or OR2_12564 ( P1_R1240_U201 , P1_U3482 , P1_U3084 );
nand NAND2_12565 ( P1_R1240_U202 , P1_R1240_U201 , P1_R1240_U140 );
not NOT1_12566 ( P1_R1240_U203 , P1_R1240_U41 );
or OR2_12567 ( P1_R1240_U204 , P1_U3083 , P1_U3485 );
or OR2_12568 ( P1_R1240_U205 , P1_U3476 , P1_U3071 );
nand NAND2_12569 ( P1_R1240_U206 , P1_R1240_U205 , P1_R1240_U42 );
nand NAND2_12570 ( P1_R1240_U207 , P1_R1240_U120 , P1_R1240_U206 );
nand NAND2_12571 ( P1_R1240_U208 , P1_R1240_U192 , P1_R1240_U23 );
nand NAND2_12572 ( P1_R1240_U209 , P1_U3479 , P1_U3070 );
nand NAND2_12573 ( P1_R1240_U210 , P1_R1240_U121 , P1_R1240_U208 );
or OR2_12574 ( P1_R1240_U211 , P1_U3071 , P1_U3476 );
nand NAND2_12575 ( P1_R1240_U212 , P1_R1240_U182 , P1_R1240_U178 );
nand NAND2_12576 ( P1_R1240_U213 , P1_U3068 , P1_U3464 );
not NOT1_12577 ( P1_R1240_U214 , P1_R1240_U46 );
nand NAND2_12578 ( P1_R1240_U215 , P1_R1240_U181 , P1_R1240_U5 );
nand NAND2_12579 ( P1_R1240_U216 , P1_R1240_U46 , P1_R1240_U177 );
nand NAND2_12580 ( P1_R1240_U217 , P1_U3064 , P1_U3467 );
not NOT1_12581 ( P1_R1240_U218 , P1_R1240_U45 );
or OR2_12582 ( P1_R1240_U219 , P1_U3470 , P1_U3060 );
nand NAND2_12583 ( P1_R1240_U220 , P1_R1240_U219 , P1_R1240_U45 );
nand NAND2_12584 ( P1_R1240_U221 , P1_R1240_U123 , P1_R1240_U220 );
nand NAND2_12585 ( P1_R1240_U222 , P1_R1240_U218 , P1_R1240_U35 );
nand NAND2_12586 ( P1_R1240_U223 , P1_U3473 , P1_U3067 );
nand NAND2_12587 ( P1_R1240_U224 , P1_R1240_U124 , P1_R1240_U222 );
or OR2_12588 ( P1_R1240_U225 , P1_U3060 , P1_U3470 );
nand NAND2_12589 ( P1_R1240_U226 , P1_R1240_U181 , P1_R1240_U178 );
not NOT1_12590 ( P1_R1240_U227 , P1_R1240_U141 );
nand NAND2_12591 ( P1_R1240_U228 , P1_U3064 , P1_U3467 );
nand NAND4_12592 ( P1_R1240_U229 , P1_R1240_U398 , P1_R1240_U397 , P1_R1240_U44 , P1_R1240_U43 );
nand NAND2_12593 ( P1_R1240_U230 , P1_R1240_U44 , P1_R1240_U43 );
nand NAND2_12594 ( P1_R1240_U231 , P1_U3068 , P1_U3464 );
nand NAND2_12595 ( P1_R1240_U232 , P1_R1240_U125 , P1_R1240_U230 );
or OR2_12596 ( P1_R1240_U233 , P1_U3083 , P1_U3485 );
or OR2_12597 ( P1_R1240_U234 , P1_U3062 , P1_U3488 );
nand NAND2_12598 ( P1_R1240_U235 , P1_R1240_U174 , P1_R1240_U7 );
nand NAND2_12599 ( P1_R1240_U236 , P1_U3062 , P1_U3488 );
nand NAND2_12600 ( P1_R1240_U237 , P1_R1240_U127 , P1_R1240_U235 );
or OR2_12601 ( P1_R1240_U238 , P1_U3488 , P1_U3062 );
nand NAND2_12602 ( P1_R1240_U239 , P1_R1240_U126 , P1_R1240_U140 );
nand NAND2_12603 ( P1_R1240_U240 , P1_R1240_U238 , P1_R1240_U237 );
not NOT1_12604 ( P1_R1240_U241 , P1_R1240_U164 );
or OR2_12605 ( P1_R1240_U242 , P1_U3080 , P1_U3497 );
or OR2_12606 ( P1_R1240_U243 , P1_U3072 , P1_U3494 );
nand NAND2_12607 ( P1_R1240_U244 , P1_R1240_U171 , P1_R1240_U8 );
nand NAND2_12608 ( P1_R1240_U245 , P1_U3080 , P1_U3497 );
nand NAND2_12609 ( P1_R1240_U246 , P1_R1240_U128 , P1_R1240_U244 );
or OR2_12610 ( P1_R1240_U247 , P1_U3491 , P1_U3063 );
or OR2_12611 ( P1_R1240_U248 , P1_U3497 , P1_U3080 );
nand NAND3_12612 ( P1_R1240_U249 , P1_R1240_U247 , P1_R1240_U164 , P1_R1240_U8 );
nand NAND2_12613 ( P1_R1240_U250 , P1_R1240_U248 , P1_R1240_U246 );
not NOT1_12614 ( P1_R1240_U251 , P1_R1240_U163 );
or OR2_12615 ( P1_R1240_U252 , P1_U3500 , P1_U3079 );
nand NAND2_12616 ( P1_R1240_U253 , P1_R1240_U252 , P1_R1240_U163 );
nand NAND2_12617 ( P1_R1240_U254 , P1_U3079 , P1_U3500 );
not NOT1_12618 ( P1_R1240_U255 , P1_R1240_U161 );
or OR2_12619 ( P1_R1240_U256 , P1_U3503 , P1_U3074 );
nand NAND2_12620 ( P1_R1240_U257 , P1_R1240_U256 , P1_R1240_U161 );
nand NAND2_12621 ( P1_R1240_U258 , P1_U3074 , P1_U3503 );
not NOT1_12622 ( P1_R1240_U259 , P1_R1240_U93 );
or OR2_12623 ( P1_R1240_U260 , P1_U3069 , P1_U3509 );
or OR2_12624 ( P1_R1240_U261 , P1_U3073 , P1_U3506 );
not NOT1_12625 ( P1_R1240_U262 , P1_R1240_U60 );
nand NAND2_12626 ( P1_R1240_U263 , P1_R1240_U61 , P1_R1240_U60 );
nand NAND2_12627 ( P1_R1240_U264 , P1_U3069 , P1_R1240_U263 );
nand NAND2_12628 ( P1_R1240_U265 , P1_U3509 , P1_R1240_U262 );
nand NAND2_12629 ( P1_R1240_U266 , P1_R1240_U9 , P1_R1240_U93 );
not NOT1_12630 ( P1_R1240_U267 , P1_R1240_U159 );
or OR2_12631 ( P1_R1240_U268 , P1_U3076 , P1_U4025 );
or OR2_12632 ( P1_R1240_U269 , P1_U3081 , P1_U3514 );
or OR2_12633 ( P1_R1240_U270 , P1_U3075 , P1_U4024 );
not NOT1_12634 ( P1_R1240_U271 , P1_R1240_U81 );
nand NAND2_12635 ( P1_R1240_U272 , P1_U4025 , P1_R1240_U271 );
nand NAND2_12636 ( P1_R1240_U273 , P1_R1240_U272 , P1_R1240_U91 );
nand NAND2_12637 ( P1_R1240_U274 , P1_R1240_U81 , P1_R1240_U82 );
nand NAND2_12638 ( P1_R1240_U275 , P1_R1240_U274 , P1_R1240_U273 );
nand NAND2_12639 ( P1_R1240_U276 , P1_R1240_U172 , P1_R1240_U10 );
nand NAND2_12640 ( P1_R1240_U277 , P1_U3075 , P1_U4024 );
nand NAND2_12641 ( P1_R1240_U278 , P1_R1240_U275 , P1_R1240_U276 );
or OR2_12642 ( P1_R1240_U279 , P1_U3512 , P1_U3082 );
or OR2_12643 ( P1_R1240_U280 , P1_U4024 , P1_U3075 );
nand NAND3_12644 ( P1_R1240_U281 , P1_R1240_U270 , P1_R1240_U159 , P1_R1240_U130 );
nand NAND2_12645 ( P1_R1240_U282 , P1_R1240_U280 , P1_R1240_U278 );
not NOT1_12646 ( P1_R1240_U283 , P1_R1240_U155 );
or OR2_12647 ( P1_R1240_U284 , P1_U4023 , P1_U3061 );
nand NAND2_12648 ( P1_R1240_U285 , P1_R1240_U284 , P1_R1240_U155 );
nand NAND2_12649 ( P1_R1240_U286 , P1_U3061 , P1_U4023 );
not NOT1_12650 ( P1_R1240_U287 , P1_R1240_U153 );
or OR2_12651 ( P1_R1240_U288 , P1_U4022 , P1_U3066 );
nand NAND2_12652 ( P1_R1240_U289 , P1_R1240_U288 , P1_R1240_U153 );
nand NAND2_12653 ( P1_R1240_U290 , P1_U3066 , P1_U4022 );
not NOT1_12654 ( P1_R1240_U291 , P1_R1240_U151 );
or OR2_12655 ( P1_R1240_U292 , P1_U3058 , P1_U4020 );
nand NAND2_12656 ( P1_R1240_U293 , P1_R1240_U173 , P1_R1240_U170 );
not NOT1_12657 ( P1_R1240_U294 , P1_R1240_U87 );
or OR2_12658 ( P1_R1240_U295 , P1_U4021 , P1_U3065 );
nand NAND3_12659 ( P1_R1240_U296 , P1_R1240_U151 , P1_R1240_U295 , P1_R1240_U165 );
not NOT1_12660 ( P1_R1240_U297 , P1_R1240_U149 );
or OR2_12661 ( P1_R1240_U298 , P1_U4018 , P1_U3053 );
nand NAND2_12662 ( P1_R1240_U299 , P1_U3053 , P1_U4018 );
not NOT1_12663 ( P1_R1240_U300 , P1_R1240_U147 );
nand NAND2_12664 ( P1_R1240_U301 , P1_U4017 , P1_R1240_U147 );
not NOT1_12665 ( P1_R1240_U302 , P1_R1240_U145 );
nand NAND2_12666 ( P1_R1240_U303 , P1_R1240_U295 , P1_R1240_U151 );
not NOT1_12667 ( P1_R1240_U304 , P1_R1240_U90 );
or OR2_12668 ( P1_R1240_U305 , P1_U4020 , P1_U3058 );
nand NAND2_12669 ( P1_R1240_U306 , P1_R1240_U305 , P1_R1240_U90 );
nand NAND3_12670 ( P1_R1240_U307 , P1_R1240_U306 , P1_R1240_U170 , P1_R1240_U150 );
nand NAND2_12671 ( P1_R1240_U308 , P1_R1240_U304 , P1_R1240_U170 );
nand NAND2_12672 ( P1_R1240_U309 , P1_U4019 , P1_U3057 );
nand NAND3_12673 ( P1_R1240_U310 , P1_R1240_U308 , P1_R1240_U309 , P1_R1240_U165 );
or OR2_12674 ( P1_R1240_U311 , P1_U3058 , P1_U4020 );
nand NAND2_12675 ( P1_R1240_U312 , P1_R1240_U279 , P1_R1240_U159 );
not NOT1_12676 ( P1_R1240_U313 , P1_R1240_U92 );
nand NAND2_12677 ( P1_R1240_U314 , P1_R1240_U10 , P1_R1240_U92 );
nand NAND2_12678 ( P1_R1240_U315 , P1_R1240_U134 , P1_R1240_U314 );
nand NAND2_12679 ( P1_R1240_U316 , P1_R1240_U314 , P1_R1240_U275 );
nand NAND2_12680 ( P1_R1240_U317 , P1_R1240_U450 , P1_R1240_U316 );
or OR2_12681 ( P1_R1240_U318 , P1_U3514 , P1_U3081 );
nand NAND2_12682 ( P1_R1240_U319 , P1_R1240_U318 , P1_R1240_U92 );
nand NAND3_12683 ( P1_R1240_U320 , P1_R1240_U319 , P1_R1240_U81 , P1_R1240_U157 );
nand NAND2_12684 ( P1_R1240_U321 , P1_R1240_U313 , P1_R1240_U81 );
nand NAND2_12685 ( P1_R1240_U322 , P1_U3076 , P1_U4025 );
nand NAND3_12686 ( P1_R1240_U323 , P1_R1240_U322 , P1_R1240_U321 , P1_R1240_U10 );
or OR2_12687 ( P1_R1240_U324 , P1_U3461 , P1_U3078 );
not NOT1_12688 ( P1_R1240_U325 , P1_R1240_U158 );
or OR2_12689 ( P1_R1240_U326 , P1_U3081 , P1_U3514 );
or OR2_12690 ( P1_R1240_U327 , P1_U3506 , P1_U3073 );
nand NAND2_12691 ( P1_R1240_U328 , P1_R1240_U327 , P1_R1240_U93 );
nand NAND2_12692 ( P1_R1240_U329 , P1_R1240_U135 , P1_R1240_U328 );
nand NAND2_12693 ( P1_R1240_U330 , P1_R1240_U259 , P1_R1240_U60 );
nand NAND2_12694 ( P1_R1240_U331 , P1_U3509 , P1_U3069 );
nand NAND3_12695 ( P1_R1240_U332 , P1_R1240_U331 , P1_R1240_U330 , P1_R1240_U9 );
or OR2_12696 ( P1_R1240_U333 , P1_U3073 , P1_U3506 );
nand NAND2_12697 ( P1_R1240_U334 , P1_R1240_U247 , P1_R1240_U164 );
not NOT1_12698 ( P1_R1240_U335 , P1_R1240_U94 );
or OR2_12699 ( P1_R1240_U336 , P1_U3494 , P1_U3072 );
nand NAND2_12700 ( P1_R1240_U337 , P1_R1240_U336 , P1_R1240_U94 );
nand NAND2_12701 ( P1_R1240_U338 , P1_R1240_U136 , P1_R1240_U337 );
nand NAND2_12702 ( P1_R1240_U339 , P1_R1240_U335 , P1_R1240_U169 );
nand NAND2_12703 ( P1_R1240_U340 , P1_U3080 , P1_U3497 );
nand NAND2_12704 ( P1_R1240_U341 , P1_R1240_U137 , P1_R1240_U339 );
or OR2_12705 ( P1_R1240_U342 , P1_U3072 , P1_U3494 );
or OR2_12706 ( P1_R1240_U343 , P1_U3485 , P1_U3083 );
nand NAND2_12707 ( P1_R1240_U344 , P1_R1240_U343 , P1_R1240_U41 );
nand NAND2_12708 ( P1_R1240_U345 , P1_R1240_U138 , P1_R1240_U344 );
nand NAND2_12709 ( P1_R1240_U346 , P1_R1240_U203 , P1_R1240_U168 );
nand NAND2_12710 ( P1_R1240_U347 , P1_U3062 , P1_U3488 );
nand NAND2_12711 ( P1_R1240_U348 , P1_R1240_U139 , P1_R1240_U346 );
nand NAND2_12712 ( P1_R1240_U349 , P1_R1240_U204 , P1_R1240_U168 );
nand NAND2_12713 ( P1_R1240_U350 , P1_R1240_U201 , P1_R1240_U62 );
nand NAND2_12714 ( P1_R1240_U351 , P1_R1240_U211 , P1_R1240_U23 );
nand NAND2_12715 ( P1_R1240_U352 , P1_R1240_U225 , P1_R1240_U35 );
nand NAND2_12716 ( P1_R1240_U353 , P1_R1240_U228 , P1_R1240_U177 );
nand NAND2_12717 ( P1_R1240_U354 , P1_R1240_U311 , P1_R1240_U170 );
nand NAND2_12718 ( P1_R1240_U355 , P1_R1240_U295 , P1_R1240_U173 );
nand NAND2_12719 ( P1_R1240_U356 , P1_R1240_U326 , P1_R1240_U81 );
nand NAND2_12720 ( P1_R1240_U357 , P1_R1240_U279 , P1_R1240_U78 );
nand NAND2_12721 ( P1_R1240_U358 , P1_R1240_U333 , P1_R1240_U60 );
nand NAND2_12722 ( P1_R1240_U359 , P1_R1240_U342 , P1_R1240_U169 );
nand NAND2_12723 ( P1_R1240_U360 , P1_R1240_U247 , P1_R1240_U69 );
nand NAND2_12724 ( P1_R1240_U361 , P1_U4017 , P1_U3054 );
nand NAND2_12725 ( P1_R1240_U362 , P1_R1240_U293 , P1_R1240_U165 );
nand NAND2_12726 ( P1_R1240_U363 , P1_U3057 , P1_R1240_U292 );
nand NAND2_12727 ( P1_R1240_U364 , P1_U4019 , P1_R1240_U292 );
nand NAND3_12728 ( P1_R1240_U365 , P1_R1240_U293 , P1_R1240_U165 , P1_R1240_U298 );
nand NAND3_12729 ( P1_R1240_U366 , P1_R1240_U151 , P1_R1240_U165 , P1_R1240_U132 );
nand NAND2_12730 ( P1_R1240_U367 , P1_R1240_U294 , P1_R1240_U298 );
nand NAND2_12731 ( P1_R1240_U368 , P1_U3083 , P1_R1240_U40 );
nand NAND2_12732 ( P1_R1240_U369 , P1_U3485 , P1_R1240_U39 );
nand NAND2_12733 ( P1_R1240_U370 , P1_R1240_U369 , P1_R1240_U368 );
nand NAND2_12734 ( P1_R1240_U371 , P1_R1240_U349 , P1_R1240_U41 );
nand NAND2_12735 ( P1_R1240_U372 , P1_R1240_U370 , P1_R1240_U203 );
nand NAND2_12736 ( P1_R1240_U373 , P1_U3084 , P1_R1240_U37 );
nand NAND2_12737 ( P1_R1240_U374 , P1_U3482 , P1_R1240_U38 );
nand NAND2_12738 ( P1_R1240_U375 , P1_R1240_U374 , P1_R1240_U373 );
nand NAND2_12739 ( P1_R1240_U376 , P1_R1240_U350 , P1_R1240_U140 );
nand NAND2_12740 ( P1_R1240_U377 , P1_R1240_U200 , P1_R1240_U375 );
nand NAND2_12741 ( P1_R1240_U378 , P1_U3070 , P1_R1240_U24 );
nand NAND2_12742 ( P1_R1240_U379 , P1_U3479 , P1_R1240_U22 );
nand NAND2_12743 ( P1_R1240_U380 , P1_U3071 , P1_R1240_U20 );
nand NAND2_12744 ( P1_R1240_U381 , P1_U3476 , P1_R1240_U21 );
nand NAND2_12745 ( P1_R1240_U382 , P1_R1240_U381 , P1_R1240_U380 );
nand NAND2_12746 ( P1_R1240_U383 , P1_R1240_U351 , P1_R1240_U42 );
nand NAND2_12747 ( P1_R1240_U384 , P1_R1240_U382 , P1_R1240_U192 );
nand NAND2_12748 ( P1_R1240_U385 , P1_U3067 , P1_R1240_U36 );
nand NAND2_12749 ( P1_R1240_U386 , P1_U3473 , P1_R1240_U27 );
nand NAND2_12750 ( P1_R1240_U387 , P1_U3060 , P1_R1240_U25 );
nand NAND2_12751 ( P1_R1240_U388 , P1_U3470 , P1_R1240_U26 );
nand NAND2_12752 ( P1_R1240_U389 , P1_R1240_U388 , P1_R1240_U387 );
nand NAND2_12753 ( P1_R1240_U390 , P1_R1240_U352 , P1_R1240_U45 );
nand NAND2_12754 ( P1_R1240_U391 , P1_R1240_U389 , P1_R1240_U218 );
nand NAND2_12755 ( P1_R1240_U392 , P1_U3064 , P1_R1240_U33 );
nand NAND2_12756 ( P1_R1240_U393 , P1_U3467 , P1_R1240_U34 );
nand NAND2_12757 ( P1_R1240_U394 , P1_R1240_U393 , P1_R1240_U392 );
nand NAND2_12758 ( P1_R1240_U395 , P1_R1240_U353 , P1_R1240_U141 );
nand NAND2_12759 ( P1_R1240_U396 , P1_R1240_U227 , P1_R1240_U394 );
nand NAND2_12760 ( P1_R1240_U397 , P1_U3068 , P1_R1240_U28 );
nand NAND2_12761 ( P1_R1240_U398 , P1_U3464 , P1_R1240_U29 );
nand NAND2_12762 ( P1_R1240_U399 , P1_U3055 , P1_R1240_U143 );
nand NAND2_12763 ( P1_R1240_U400 , P1_U4028 , P1_R1240_U142 );
nand NAND2_12764 ( P1_R1240_U401 , P1_U3055 , P1_R1240_U143 );
nand NAND2_12765 ( P1_R1240_U402 , P1_U4028 , P1_R1240_U142 );
nand NAND2_12766 ( P1_R1240_U403 , P1_R1240_U402 , P1_R1240_U401 );
nand NAND2_12767 ( P1_R1240_U404 , P1_R1240_U144 , P1_R1240_U145 );
nand NAND2_12768 ( P1_R1240_U405 , P1_R1240_U302 , P1_R1240_U403 );
nand NAND2_12769 ( P1_R1240_U406 , P1_U3054 , P1_R1240_U89 );
nand NAND2_12770 ( P1_R1240_U407 , P1_U4017 , P1_R1240_U88 );
nand NAND2_12771 ( P1_R1240_U408 , P1_U3054 , P1_R1240_U89 );
nand NAND2_12772 ( P1_R1240_U409 , P1_U4017 , P1_R1240_U88 );
nand NAND2_12773 ( P1_R1240_U410 , P1_R1240_U409 , P1_R1240_U408 );
nand NAND2_12774 ( P1_R1240_U411 , P1_R1240_U146 , P1_R1240_U147 );
nand NAND2_12775 ( P1_R1240_U412 , P1_R1240_U300 , P1_R1240_U410 );
nand NAND2_12776 ( P1_R1240_U413 , P1_U3053 , P1_R1240_U47 );
nand NAND2_12777 ( P1_R1240_U414 , P1_U4018 , P1_R1240_U48 );
nand NAND2_12778 ( P1_R1240_U415 , P1_U3053 , P1_R1240_U47 );
nand NAND2_12779 ( P1_R1240_U416 , P1_U4018 , P1_R1240_U48 );
nand NAND2_12780 ( P1_R1240_U417 , P1_R1240_U416 , P1_R1240_U415 );
nand NAND2_12781 ( P1_R1240_U418 , P1_R1240_U148 , P1_R1240_U149 );
nand NAND2_12782 ( P1_R1240_U419 , P1_R1240_U297 , P1_R1240_U417 );
nand NAND2_12783 ( P1_R1240_U420 , P1_U3057 , P1_R1240_U50 );
nand NAND2_12784 ( P1_R1240_U421 , P1_U4019 , P1_R1240_U49 );
nand NAND2_12785 ( P1_R1240_U422 , P1_U3058 , P1_R1240_U51 );
nand NAND2_12786 ( P1_R1240_U423 , P1_U4020 , P1_R1240_U52 );
nand NAND2_12787 ( P1_R1240_U424 , P1_R1240_U423 , P1_R1240_U422 );
nand NAND2_12788 ( P1_R1240_U425 , P1_R1240_U354 , P1_R1240_U90 );
nand NAND2_12789 ( P1_R1240_U426 , P1_R1240_U424 , P1_R1240_U304 );
nand NAND2_12790 ( P1_R1240_U427 , P1_U3065 , P1_R1240_U53 );
nand NAND2_12791 ( P1_R1240_U428 , P1_U4021 , P1_R1240_U54 );
nand NAND2_12792 ( P1_R1240_U429 , P1_R1240_U428 , P1_R1240_U427 );
nand NAND2_12793 ( P1_R1240_U430 , P1_R1240_U355 , P1_R1240_U151 );
nand NAND2_12794 ( P1_R1240_U431 , P1_R1240_U291 , P1_R1240_U429 );
nand NAND2_12795 ( P1_R1240_U432 , P1_U3066 , P1_R1240_U85 );
nand NAND2_12796 ( P1_R1240_U433 , P1_U4022 , P1_R1240_U86 );
nand NAND2_12797 ( P1_R1240_U434 , P1_U3066 , P1_R1240_U85 );
nand NAND2_12798 ( P1_R1240_U435 , P1_U4022 , P1_R1240_U86 );
nand NAND2_12799 ( P1_R1240_U436 , P1_R1240_U435 , P1_R1240_U434 );
nand NAND2_12800 ( P1_R1240_U437 , P1_R1240_U152 , P1_R1240_U153 );
nand NAND2_12801 ( P1_R1240_U438 , P1_R1240_U287 , P1_R1240_U436 );
nand NAND2_12802 ( P1_R1240_U439 , P1_U3061 , P1_R1240_U83 );
nand NAND2_12803 ( P1_R1240_U440 , P1_U4023 , P1_R1240_U84 );
nand NAND2_12804 ( P1_R1240_U441 , P1_U3061 , P1_R1240_U83 );
nand NAND2_12805 ( P1_R1240_U442 , P1_U4023 , P1_R1240_U84 );
nand NAND2_12806 ( P1_R1240_U443 , P1_R1240_U442 , P1_R1240_U441 );
nand NAND2_12807 ( P1_R1240_U444 , P1_R1240_U154 , P1_R1240_U155 );
nand NAND2_12808 ( P1_R1240_U445 , P1_R1240_U283 , P1_R1240_U443 );
nand NAND2_12809 ( P1_R1240_U446 , P1_U3075 , P1_R1240_U55 );
nand NAND2_12810 ( P1_R1240_U447 , P1_U4024 , P1_R1240_U56 );
nand NAND2_12811 ( P1_R1240_U448 , P1_U3075 , P1_R1240_U55 );
nand NAND2_12812 ( P1_R1240_U449 , P1_U4024 , P1_R1240_U56 );
nand NAND2_12813 ( P1_R1240_U450 , P1_R1240_U449 , P1_R1240_U448 );
nand NAND2_12814 ( P1_R1240_U451 , P1_U3076 , P1_R1240_U82 );
nand NAND2_12815 ( P1_R1240_U452 , P1_U4025 , P1_R1240_U91 );
nand NAND2_12816 ( P1_R1240_U453 , P1_R1240_U179 , P1_R1240_U158 );
nand NAND2_12817 ( P1_R1240_U454 , P1_R1240_U325 , P1_R1240_U32 );
nand NAND2_12818 ( P1_R1240_U455 , P1_U3081 , P1_R1240_U79 );
nand NAND2_12819 ( P1_R1240_U456 , P1_U3514 , P1_R1240_U80 );
nand NAND2_12820 ( P1_R1240_U457 , P1_R1240_U456 , P1_R1240_U455 );
nand NAND2_12821 ( P1_R1240_U458 , P1_R1240_U356 , P1_R1240_U92 );
nand NAND2_12822 ( P1_R1240_U459 , P1_R1240_U457 , P1_R1240_U313 );
nand NAND2_12823 ( P1_R1240_U460 , P1_U3082 , P1_R1240_U76 );
nand NAND2_12824 ( P1_R1240_U461 , P1_U3512 , P1_R1240_U77 );
nand NAND2_12825 ( P1_R1240_U462 , P1_R1240_U461 , P1_R1240_U460 );
nand NAND2_12826 ( P1_R1240_U463 , P1_R1240_U357 , P1_R1240_U159 );
nand NAND2_12827 ( P1_R1240_U464 , P1_R1240_U267 , P1_R1240_U462 );
nand NAND2_12828 ( P1_R1240_U465 , P1_U3069 , P1_R1240_U61 );
nand NAND2_12829 ( P1_R1240_U466 , P1_U3509 , P1_R1240_U59 );
nand NAND2_12830 ( P1_R1240_U467 , P1_U3073 , P1_R1240_U57 );
nand NAND2_12831 ( P1_R1240_U468 , P1_U3506 , P1_R1240_U58 );
nand NAND2_12832 ( P1_R1240_U469 , P1_R1240_U468 , P1_R1240_U467 );
nand NAND2_12833 ( P1_R1240_U470 , P1_R1240_U358 , P1_R1240_U93 );
nand NAND2_12834 ( P1_R1240_U471 , P1_R1240_U469 , P1_R1240_U259 );
nand NAND2_12835 ( P1_R1240_U472 , P1_U3074 , P1_R1240_U74 );
nand NAND2_12836 ( P1_R1240_U473 , P1_U3503 , P1_R1240_U75 );
nand NAND2_12837 ( P1_R1240_U474 , P1_U3074 , P1_R1240_U74 );
nand NAND2_12838 ( P1_R1240_U475 , P1_U3503 , P1_R1240_U75 );
nand NAND2_12839 ( P1_R1240_U476 , P1_R1240_U475 , P1_R1240_U474 );
nand NAND2_12840 ( P1_R1240_U477 , P1_R1240_U160 , P1_R1240_U161 );
nand NAND2_12841 ( P1_R1240_U478 , P1_R1240_U255 , P1_R1240_U476 );
nand NAND2_12842 ( P1_R1240_U479 , P1_U3079 , P1_R1240_U72 );
nand NAND2_12843 ( P1_R1240_U480 , P1_U3500 , P1_R1240_U73 );
nand NAND2_12844 ( P1_R1240_U481 , P1_U3079 , P1_R1240_U72 );
nand NAND2_12845 ( P1_R1240_U482 , P1_U3500 , P1_R1240_U73 );
nand NAND2_12846 ( P1_R1240_U483 , P1_R1240_U482 , P1_R1240_U481 );
nand NAND2_12847 ( P1_R1240_U484 , P1_R1240_U162 , P1_R1240_U163 );
nand NAND2_12848 ( P1_R1240_U485 , P1_R1240_U251 , P1_R1240_U483 );
nand NAND2_12849 ( P1_R1240_U486 , P1_U3080 , P1_R1240_U70 );
nand NAND2_12850 ( P1_R1240_U487 , P1_U3497 , P1_R1240_U71 );
nand NAND2_12851 ( P1_R1240_U488 , P1_U3072 , P1_R1240_U65 );
nand NAND2_12852 ( P1_R1240_U489 , P1_U3494 , P1_R1240_U66 );
nand NAND2_12853 ( P1_R1240_U490 , P1_R1240_U489 , P1_R1240_U488 );
nand NAND2_12854 ( P1_R1240_U491 , P1_R1240_U359 , P1_R1240_U94 );
nand NAND2_12855 ( P1_R1240_U492 , P1_R1240_U490 , P1_R1240_U335 );
nand NAND2_12856 ( P1_R1240_U493 , P1_U3063 , P1_R1240_U67 );
nand NAND2_12857 ( P1_R1240_U494 , P1_U3491 , P1_R1240_U68 );
nand NAND2_12858 ( P1_R1240_U495 , P1_R1240_U494 , P1_R1240_U493 );
nand NAND2_12859 ( P1_R1240_U496 , P1_R1240_U360 , P1_R1240_U164 );
nand NAND2_12860 ( P1_R1240_U497 , P1_R1240_U241 , P1_R1240_U495 );
nand NAND2_12861 ( P1_R1240_U498 , P1_U3062 , P1_R1240_U63 );
nand NAND2_12862 ( P1_R1240_U499 , P1_U3488 , P1_R1240_U64 );
nand NAND2_12863 ( P1_R1240_U500 , P1_U3077 , P1_R1240_U30 );
nand NAND2_12864 ( P1_R1240_U501 , P1_U3456 , P1_R1240_U31 );
and AND2_12865 ( P1_R1162_U4 , P1_R1162_U95 , P1_R1162_U94 );
and AND2_12866 ( P1_R1162_U5 , P1_R1162_U96 , P1_R1162_U97 );
and AND2_12867 ( P1_R1162_U6 , P1_R1162_U113 , P1_R1162_U112 );
and AND2_12868 ( P1_R1162_U7 , P1_R1162_U155 , P1_R1162_U154 );
and AND2_12869 ( P1_R1162_U8 , P1_R1162_U164 , P1_R1162_U163 );
and AND2_12870 ( P1_R1162_U9 , P1_R1162_U182 , P1_R1162_U181 );
and AND2_12871 ( P1_R1162_U10 , P1_R1162_U218 , P1_R1162_U215 );
and AND2_12872 ( P1_R1162_U11 , P1_R1162_U211 , P1_R1162_U208 );
and AND2_12873 ( P1_R1162_U12 , P1_R1162_U202 , P1_R1162_U199 );
and AND2_12874 ( P1_R1162_U13 , P1_R1162_U196 , P1_R1162_U192 );
and AND2_12875 ( P1_R1162_U14 , P1_R1162_U151 , P1_R1162_U148 );
and AND2_12876 ( P1_R1162_U15 , P1_R1162_U143 , P1_R1162_U140 );
and AND2_12877 ( P1_R1162_U16 , P1_R1162_U129 , P1_R1162_U126 );
not NOT1_12878 ( P1_R1162_U17 , P1_REG1_REG_6_ );
not NOT1_12879 ( P1_R1162_U18 , P1_U3475 );
not NOT1_12880 ( P1_R1162_U19 , P1_U3478 );
nand NAND2_12881 ( P1_R1162_U20 , P1_U3475 , P1_REG1_REG_6_ );
not NOT1_12882 ( P1_R1162_U21 , P1_REG1_REG_7_ );
not NOT1_12883 ( P1_R1162_U22 , P1_REG1_REG_4_ );
not NOT1_12884 ( P1_R1162_U23 , P1_U3469 );
not NOT1_12885 ( P1_R1162_U24 , P1_U3472 );
not NOT1_12886 ( P1_R1162_U25 , P1_REG1_REG_2_ );
not NOT1_12887 ( P1_R1162_U26 , P1_U3463 );
not NOT1_12888 ( P1_R1162_U27 , P1_REG1_REG_0_ );
not NOT1_12889 ( P1_R1162_U28 , P1_U3454 );
nand NAND2_12890 ( P1_R1162_U29 , P1_U3454 , P1_REG1_REG_0_ );
not NOT1_12891 ( P1_R1162_U30 , P1_REG1_REG_3_ );
not NOT1_12892 ( P1_R1162_U31 , P1_U3466 );
nand NAND2_12893 ( P1_R1162_U32 , P1_U3469 , P1_REG1_REG_4_ );
not NOT1_12894 ( P1_R1162_U33 , P1_REG1_REG_5_ );
not NOT1_12895 ( P1_R1162_U34 , P1_REG1_REG_8_ );
not NOT1_12896 ( P1_R1162_U35 , P1_U3481 );
not NOT1_12897 ( P1_R1162_U36 , P1_U3484 );
not NOT1_12898 ( P1_R1162_U37 , P1_REG1_REG_9_ );
nand NAND2_12899 ( P1_R1162_U38 , P1_R1162_U49 , P1_R1162_U121 );
nand NAND3_12900 ( P1_R1162_U39 , P1_R1162_U110 , P1_R1162_U108 , P1_R1162_U109 );
nand NAND2_12901 ( P1_R1162_U40 , P1_R1162_U98 , P1_R1162_U99 );
nand NAND2_12902 ( P1_R1162_U41 , P1_REG1_REG_1_ , P1_U3460 );
nand NAND3_12903 ( P1_R1162_U42 , P1_R1162_U136 , P1_R1162_U134 , P1_R1162_U135 );
nand NAND2_12904 ( P1_R1162_U43 , P1_R1162_U132 , P1_R1162_U131 );
not NOT1_12905 ( P1_R1162_U44 , P1_REG1_REG_16_ );
not NOT1_12906 ( P1_R1162_U45 , P1_U3505 );
not NOT1_12907 ( P1_R1162_U46 , P1_U3508 );
nand NAND2_12908 ( P1_R1162_U47 , P1_U3505 , P1_REG1_REG_16_ );
not NOT1_12909 ( P1_R1162_U48 , P1_REG1_REG_17_ );
nand NAND2_12910 ( P1_R1162_U49 , P1_U3481 , P1_REG1_REG_8_ );
not NOT1_12911 ( P1_R1162_U50 , P1_REG1_REG_10_ );
not NOT1_12912 ( P1_R1162_U51 , P1_U3487 );
not NOT1_12913 ( P1_R1162_U52 , P1_REG1_REG_12_ );
not NOT1_12914 ( P1_R1162_U53 , P1_U3493 );
not NOT1_12915 ( P1_R1162_U54 , P1_REG1_REG_11_ );
not NOT1_12916 ( P1_R1162_U55 , P1_U3490 );
nand NAND2_12917 ( P1_R1162_U56 , P1_U3490 , P1_REG1_REG_11_ );
not NOT1_12918 ( P1_R1162_U57 , P1_REG1_REG_13_ );
not NOT1_12919 ( P1_R1162_U58 , P1_U3496 );
not NOT1_12920 ( P1_R1162_U59 , P1_REG1_REG_14_ );
not NOT1_12921 ( P1_R1162_U60 , P1_U3499 );
not NOT1_12922 ( P1_R1162_U61 , P1_REG1_REG_15_ );
not NOT1_12923 ( P1_R1162_U62 , P1_U3502 );
not NOT1_12924 ( P1_R1162_U63 , P1_REG1_REG_18_ );
not NOT1_12925 ( P1_R1162_U64 , P1_U3511 );
nand NAND3_12926 ( P1_R1162_U65 , P1_R1162_U186 , P1_R1162_U185 , P1_R1162_U187 );
nand NAND2_12927 ( P1_R1162_U66 , P1_R1162_U179 , P1_R1162_U178 );
nand NAND2_12928 ( P1_R1162_U67 , P1_R1162_U56 , P1_R1162_U204 );
nand NAND2_12929 ( P1_R1162_U68 , P1_R1162_U259 , P1_R1162_U258 );
nand NAND2_12930 ( P1_R1162_U69 , P1_R1162_U308 , P1_R1162_U307 );
nand NAND2_12931 ( P1_R1162_U70 , P1_R1162_U231 , P1_R1162_U230 );
nand NAND2_12932 ( P1_R1162_U71 , P1_R1162_U236 , P1_R1162_U235 );
nand NAND2_12933 ( P1_R1162_U72 , P1_R1162_U243 , P1_R1162_U242 );
nand NAND2_12934 ( P1_R1162_U73 , P1_R1162_U250 , P1_R1162_U249 );
nand NAND2_12935 ( P1_R1162_U74 , P1_R1162_U255 , P1_R1162_U254 );
nand NAND2_12936 ( P1_R1162_U75 , P1_R1162_U271 , P1_R1162_U270 );
nand NAND2_12937 ( P1_R1162_U76 , P1_R1162_U278 , P1_R1162_U277 );
nand NAND2_12938 ( P1_R1162_U77 , P1_R1162_U285 , P1_R1162_U284 );
nand NAND2_12939 ( P1_R1162_U78 , P1_R1162_U292 , P1_R1162_U291 );
nand NAND2_12940 ( P1_R1162_U79 , P1_R1162_U299 , P1_R1162_U298 );
nand NAND2_12941 ( P1_R1162_U80 , P1_R1162_U304 , P1_R1162_U303 );
nand NAND3_12942 ( P1_R1162_U81 , P1_R1162_U117 , P1_R1162_U116 , P1_R1162_U118 );
nand NAND2_12943 ( P1_R1162_U82 , P1_R1162_U133 , P1_R1162_U145 );
nand NAND2_12944 ( P1_R1162_U83 , P1_R1162_U41 , P1_R1162_U152 );
not NOT1_12945 ( P1_R1162_U84 , P1_U3452 );
not NOT1_12946 ( P1_R1162_U85 , P1_REG1_REG_19_ );
nand NAND2_12947 ( P1_R1162_U86 , P1_R1162_U175 , P1_R1162_U174 );
nand NAND2_12948 ( P1_R1162_U87 , P1_R1162_U171 , P1_R1162_U170 );
nand NAND2_12949 ( P1_R1162_U88 , P1_R1162_U161 , P1_R1162_U160 );
not NOT1_12950 ( P1_R1162_U89 , P1_R1162_U32 );
nand NAND2_12951 ( P1_R1162_U90 , P1_REG1_REG_9_ , P1_U3484 );
nand NAND2_12952 ( P1_R1162_U91 , P1_U3493 , P1_REG1_REG_12_ );
not NOT1_12953 ( P1_R1162_U92 , P1_R1162_U56 );
not NOT1_12954 ( P1_R1162_U93 , P1_R1162_U49 );
or OR2_12955 ( P1_R1162_U94 , P1_U3472 , P1_REG1_REG_5_ );
or OR2_12956 ( P1_R1162_U95 , P1_U3469 , P1_REG1_REG_4_ );
or OR2_12957 ( P1_R1162_U96 , P1_REG1_REG_3_ , P1_U3466 );
or OR2_12958 ( P1_R1162_U97 , P1_REG1_REG_2_ , P1_U3463 );
not NOT1_12959 ( P1_R1162_U98 , P1_R1162_U29 );
or OR2_12960 ( P1_R1162_U99 , P1_REG1_REG_1_ , P1_U3460 );
not NOT1_12961 ( P1_R1162_U100 , P1_R1162_U40 );
not NOT1_12962 ( P1_R1162_U101 , P1_R1162_U41 );
nand NAND2_12963 ( P1_R1162_U102 , P1_R1162_U40 , P1_R1162_U41 );
nand NAND3_12964 ( P1_R1162_U103 , P1_REG1_REG_2_ , P1_U3463 , P1_R1162_U96 );
nand NAND2_12965 ( P1_R1162_U104 , P1_R1162_U5 , P1_R1162_U102 );
nand NAND2_12966 ( P1_R1162_U105 , P1_U3466 , P1_REG1_REG_3_ );
nand NAND3_12967 ( P1_R1162_U106 , P1_R1162_U105 , P1_R1162_U103 , P1_R1162_U104 );
nand NAND2_12968 ( P1_R1162_U107 , P1_R1162_U33 , P1_R1162_U32 );
nand NAND2_12969 ( P1_R1162_U108 , P1_U3472 , P1_R1162_U107 );
nand NAND2_12970 ( P1_R1162_U109 , P1_R1162_U4 , P1_R1162_U106 );
nand NAND2_12971 ( P1_R1162_U110 , P1_REG1_REG_5_ , P1_R1162_U89 );
not NOT1_12972 ( P1_R1162_U111 , P1_R1162_U39 );
or OR2_12973 ( P1_R1162_U112 , P1_U3478 , P1_REG1_REG_7_ );
or OR2_12974 ( P1_R1162_U113 , P1_U3475 , P1_REG1_REG_6_ );
not NOT1_12975 ( P1_R1162_U114 , P1_R1162_U20 );
nand NAND2_12976 ( P1_R1162_U115 , P1_R1162_U21 , P1_R1162_U20 );
nand NAND2_12977 ( P1_R1162_U116 , P1_U3478 , P1_R1162_U115 );
nand NAND2_12978 ( P1_R1162_U117 , P1_REG1_REG_7_ , P1_R1162_U114 );
nand NAND2_12979 ( P1_R1162_U118 , P1_R1162_U6 , P1_R1162_U39 );
not NOT1_12980 ( P1_R1162_U119 , P1_R1162_U81 );
or OR2_12981 ( P1_R1162_U120 , P1_REG1_REG_8_ , P1_U3481 );
nand NAND2_12982 ( P1_R1162_U121 , P1_R1162_U120 , P1_R1162_U81 );
not NOT1_12983 ( P1_R1162_U122 , P1_R1162_U38 );
or OR2_12984 ( P1_R1162_U123 , P1_U3484 , P1_REG1_REG_9_ );
or OR2_12985 ( P1_R1162_U124 , P1_REG1_REG_6_ , P1_U3475 );
nand NAND2_12986 ( P1_R1162_U125 , P1_R1162_U124 , P1_R1162_U39 );
nand NAND4_12987 ( P1_R1162_U126 , P1_R1162_U238 , P1_R1162_U237 , P1_R1162_U20 , P1_R1162_U125 );
nand NAND2_12988 ( P1_R1162_U127 , P1_R1162_U111 , P1_R1162_U20 );
nand NAND2_12989 ( P1_R1162_U128 , P1_REG1_REG_7_ , P1_U3478 );
nand NAND3_12990 ( P1_R1162_U129 , P1_R1162_U128 , P1_R1162_U6 , P1_R1162_U127 );
or OR2_12991 ( P1_R1162_U130 , P1_U3475 , P1_REG1_REG_6_ );
nand NAND2_12992 ( P1_R1162_U131 , P1_R1162_U101 , P1_R1162_U97 );
nand NAND2_12993 ( P1_R1162_U132 , P1_U3463 , P1_REG1_REG_2_ );
not NOT1_12994 ( P1_R1162_U133 , P1_R1162_U43 );
nand NAND2_12995 ( P1_R1162_U134 , P1_R1162_U100 , P1_R1162_U5 );
nand NAND2_12996 ( P1_R1162_U135 , P1_R1162_U43 , P1_R1162_U96 );
nand NAND2_12997 ( P1_R1162_U136 , P1_U3466 , P1_REG1_REG_3_ );
not NOT1_12998 ( P1_R1162_U137 , P1_R1162_U42 );
or OR2_12999 ( P1_R1162_U138 , P1_REG1_REG_4_ , P1_U3469 );
nand NAND2_13000 ( P1_R1162_U139 , P1_R1162_U138 , P1_R1162_U42 );
nand NAND4_13001 ( P1_R1162_U140 , P1_R1162_U245 , P1_R1162_U244 , P1_R1162_U32 , P1_R1162_U139 );
nand NAND2_13002 ( P1_R1162_U141 , P1_R1162_U137 , P1_R1162_U32 );
nand NAND2_13003 ( P1_R1162_U142 , P1_REG1_REG_5_ , P1_U3472 );
nand NAND3_13004 ( P1_R1162_U143 , P1_R1162_U142 , P1_R1162_U4 , P1_R1162_U141 );
or OR2_13005 ( P1_R1162_U144 , P1_U3469 , P1_REG1_REG_4_ );
nand NAND2_13006 ( P1_R1162_U145 , P1_R1162_U100 , P1_R1162_U97 );
not NOT1_13007 ( P1_R1162_U146 , P1_R1162_U82 );
nand NAND2_13008 ( P1_R1162_U147 , P1_U3466 , P1_REG1_REG_3_ );
nand NAND4_13009 ( P1_R1162_U148 , P1_R1162_U257 , P1_R1162_U256 , P1_R1162_U41 , P1_R1162_U40 );
nand NAND2_13010 ( P1_R1162_U149 , P1_R1162_U41 , P1_R1162_U40 );
nand NAND2_13011 ( P1_R1162_U150 , P1_U3463 , P1_REG1_REG_2_ );
nand NAND3_13012 ( P1_R1162_U151 , P1_R1162_U150 , P1_R1162_U97 , P1_R1162_U149 );
or OR2_13013 ( P1_R1162_U152 , P1_REG1_REG_1_ , P1_U3460 );
not NOT1_13014 ( P1_R1162_U153 , P1_R1162_U83 );
or OR2_13015 ( P1_R1162_U154 , P1_U3484 , P1_REG1_REG_9_ );
or OR2_13016 ( P1_R1162_U155 , P1_U3487 , P1_REG1_REG_10_ );
nand NAND2_13017 ( P1_R1162_U156 , P1_R1162_U93 , P1_R1162_U7 );
nand NAND2_13018 ( P1_R1162_U157 , P1_U3487 , P1_REG1_REG_10_ );
nand NAND3_13019 ( P1_R1162_U158 , P1_R1162_U157 , P1_R1162_U90 , P1_R1162_U156 );
or OR2_13020 ( P1_R1162_U159 , P1_REG1_REG_10_ , P1_U3487 );
nand NAND3_13021 ( P1_R1162_U160 , P1_R1162_U120 , P1_R1162_U7 , P1_R1162_U81 );
nand NAND2_13022 ( P1_R1162_U161 , P1_R1162_U159 , P1_R1162_U158 );
not NOT1_13023 ( P1_R1162_U162 , P1_R1162_U88 );
or OR2_13024 ( P1_R1162_U163 , P1_U3496 , P1_REG1_REG_13_ );
or OR2_13025 ( P1_R1162_U164 , P1_U3493 , P1_REG1_REG_12_ );
nand NAND2_13026 ( P1_R1162_U165 , P1_R1162_U92 , P1_R1162_U8 );
nand NAND2_13027 ( P1_R1162_U166 , P1_U3496 , P1_REG1_REG_13_ );
nand NAND3_13028 ( P1_R1162_U167 , P1_R1162_U166 , P1_R1162_U91 , P1_R1162_U165 );
or OR2_13029 ( P1_R1162_U168 , P1_REG1_REG_11_ , P1_U3490 );
or OR2_13030 ( P1_R1162_U169 , P1_REG1_REG_13_ , P1_U3496 );
nand NAND3_13031 ( P1_R1162_U170 , P1_R1162_U168 , P1_R1162_U8 , P1_R1162_U88 );
nand NAND2_13032 ( P1_R1162_U171 , P1_R1162_U169 , P1_R1162_U167 );
not NOT1_13033 ( P1_R1162_U172 , P1_R1162_U87 );
or OR2_13034 ( P1_R1162_U173 , P1_REG1_REG_14_ , P1_U3499 );
nand NAND2_13035 ( P1_R1162_U174 , P1_R1162_U173 , P1_R1162_U87 );
nand NAND2_13036 ( P1_R1162_U175 , P1_U3499 , P1_REG1_REG_14_ );
not NOT1_13037 ( P1_R1162_U176 , P1_R1162_U86 );
or OR2_13038 ( P1_R1162_U177 , P1_REG1_REG_15_ , P1_U3502 );
nand NAND2_13039 ( P1_R1162_U178 , P1_R1162_U177 , P1_R1162_U86 );
nand NAND2_13040 ( P1_R1162_U179 , P1_U3502 , P1_REG1_REG_15_ );
not NOT1_13041 ( P1_R1162_U180 , P1_R1162_U66 );
or OR2_13042 ( P1_R1162_U181 , P1_U3508 , P1_REG1_REG_17_ );
or OR2_13043 ( P1_R1162_U182 , P1_U3505 , P1_REG1_REG_16_ );
not NOT1_13044 ( P1_R1162_U183 , P1_R1162_U47 );
nand NAND2_13045 ( P1_R1162_U184 , P1_R1162_U48 , P1_R1162_U47 );
nand NAND2_13046 ( P1_R1162_U185 , P1_U3508 , P1_R1162_U184 );
nand NAND2_13047 ( P1_R1162_U186 , P1_REG1_REG_17_ , P1_R1162_U183 );
nand NAND2_13048 ( P1_R1162_U187 , P1_R1162_U9 , P1_R1162_U66 );
not NOT1_13049 ( P1_R1162_U188 , P1_R1162_U65 );
or OR2_13050 ( P1_R1162_U189 , P1_REG1_REG_18_ , P1_U3511 );
nand NAND2_13051 ( P1_R1162_U190 , P1_R1162_U189 , P1_R1162_U65 );
nand NAND2_13052 ( P1_R1162_U191 , P1_U3511 , P1_REG1_REG_18_ );
nand NAND4_13053 ( P1_R1162_U192 , P1_R1162_U261 , P1_R1162_U260 , P1_R1162_U191 , P1_R1162_U190 );
nand NAND2_13054 ( P1_R1162_U193 , P1_U3511 , P1_REG1_REG_18_ );
nand NAND2_13055 ( P1_R1162_U194 , P1_R1162_U188 , P1_R1162_U193 );
or OR2_13056 ( P1_R1162_U195 , P1_U3511 , P1_REG1_REG_18_ );
nand NAND3_13057 ( P1_R1162_U196 , P1_R1162_U195 , P1_R1162_U264 , P1_R1162_U194 );
or OR2_13058 ( P1_R1162_U197 , P1_REG1_REG_16_ , P1_U3505 );
nand NAND2_13059 ( P1_R1162_U198 , P1_R1162_U197 , P1_R1162_U66 );
nand NAND4_13060 ( P1_R1162_U199 , P1_R1162_U273 , P1_R1162_U272 , P1_R1162_U47 , P1_R1162_U198 );
nand NAND2_13061 ( P1_R1162_U200 , P1_R1162_U180 , P1_R1162_U47 );
nand NAND2_13062 ( P1_R1162_U201 , P1_REG1_REG_17_ , P1_U3508 );
nand NAND3_13063 ( P1_R1162_U202 , P1_R1162_U201 , P1_R1162_U9 , P1_R1162_U200 );
or OR2_13064 ( P1_R1162_U203 , P1_U3505 , P1_REG1_REG_16_ );
nand NAND2_13065 ( P1_R1162_U204 , P1_R1162_U168 , P1_R1162_U88 );
not NOT1_13066 ( P1_R1162_U205 , P1_R1162_U67 );
or OR2_13067 ( P1_R1162_U206 , P1_REG1_REG_12_ , P1_U3493 );
nand NAND2_13068 ( P1_R1162_U207 , P1_R1162_U206 , P1_R1162_U67 );
nand NAND4_13069 ( P1_R1162_U208 , P1_R1162_U294 , P1_R1162_U293 , P1_R1162_U91 , P1_R1162_U207 );
nand NAND2_13070 ( P1_R1162_U209 , P1_R1162_U205 , P1_R1162_U91 );
nand NAND2_13071 ( P1_R1162_U210 , P1_U3496 , P1_REG1_REG_13_ );
nand NAND3_13072 ( P1_R1162_U211 , P1_R1162_U210 , P1_R1162_U8 , P1_R1162_U209 );
or OR2_13073 ( P1_R1162_U212 , P1_U3493 , P1_REG1_REG_12_ );
or OR2_13074 ( P1_R1162_U213 , P1_REG1_REG_9_ , P1_U3484 );
nand NAND2_13075 ( P1_R1162_U214 , P1_R1162_U213 , P1_R1162_U38 );
nand NAND4_13076 ( P1_R1162_U215 , P1_R1162_U306 , P1_R1162_U305 , P1_R1162_U90 , P1_R1162_U214 );
nand NAND2_13077 ( P1_R1162_U216 , P1_R1162_U122 , P1_R1162_U90 );
nand NAND2_13078 ( P1_R1162_U217 , P1_U3487 , P1_REG1_REG_10_ );
nand NAND3_13079 ( P1_R1162_U218 , P1_R1162_U217 , P1_R1162_U7 , P1_R1162_U216 );
nand NAND2_13080 ( P1_R1162_U219 , P1_R1162_U123 , P1_R1162_U90 );
nand NAND2_13081 ( P1_R1162_U220 , P1_R1162_U120 , P1_R1162_U49 );
nand NAND2_13082 ( P1_R1162_U221 , P1_R1162_U130 , P1_R1162_U20 );
nand NAND2_13083 ( P1_R1162_U222 , P1_R1162_U144 , P1_R1162_U32 );
nand NAND2_13084 ( P1_R1162_U223 , P1_R1162_U147 , P1_R1162_U96 );
nand NAND2_13085 ( P1_R1162_U224 , P1_R1162_U203 , P1_R1162_U47 );
nand NAND2_13086 ( P1_R1162_U225 , P1_R1162_U212 , P1_R1162_U91 );
nand NAND2_13087 ( P1_R1162_U226 , P1_R1162_U168 , P1_R1162_U56 );
nand NAND2_13088 ( P1_R1162_U227 , P1_U3484 , P1_R1162_U37 );
nand NAND2_13089 ( P1_R1162_U228 , P1_REG1_REG_9_ , P1_R1162_U36 );
nand NAND2_13090 ( P1_R1162_U229 , P1_R1162_U228 , P1_R1162_U227 );
nand NAND2_13091 ( P1_R1162_U230 , P1_R1162_U219 , P1_R1162_U38 );
nand NAND2_13092 ( P1_R1162_U231 , P1_R1162_U229 , P1_R1162_U122 );
nand NAND2_13093 ( P1_R1162_U232 , P1_U3481 , P1_R1162_U34 );
nand NAND2_13094 ( P1_R1162_U233 , P1_REG1_REG_8_ , P1_R1162_U35 );
nand NAND2_13095 ( P1_R1162_U234 , P1_R1162_U233 , P1_R1162_U232 );
nand NAND2_13096 ( P1_R1162_U235 , P1_R1162_U220 , P1_R1162_U81 );
nand NAND2_13097 ( P1_R1162_U236 , P1_R1162_U119 , P1_R1162_U234 );
nand NAND2_13098 ( P1_R1162_U237 , P1_U3478 , P1_R1162_U21 );
nand NAND2_13099 ( P1_R1162_U238 , P1_REG1_REG_7_ , P1_R1162_U19 );
nand NAND2_13100 ( P1_R1162_U239 , P1_U3475 , P1_R1162_U17 );
nand NAND2_13101 ( P1_R1162_U240 , P1_REG1_REG_6_ , P1_R1162_U18 );
nand NAND2_13102 ( P1_R1162_U241 , P1_R1162_U240 , P1_R1162_U239 );
nand NAND2_13103 ( P1_R1162_U242 , P1_R1162_U221 , P1_R1162_U39 );
nand NAND2_13104 ( P1_R1162_U243 , P1_R1162_U241 , P1_R1162_U111 );
nand NAND2_13105 ( P1_R1162_U244 , P1_U3472 , P1_R1162_U33 );
nand NAND2_13106 ( P1_R1162_U245 , P1_REG1_REG_5_ , P1_R1162_U24 );
nand NAND2_13107 ( P1_R1162_U246 , P1_U3469 , P1_R1162_U22 );
nand NAND2_13108 ( P1_R1162_U247 , P1_REG1_REG_4_ , P1_R1162_U23 );
nand NAND2_13109 ( P1_R1162_U248 , P1_R1162_U247 , P1_R1162_U246 );
nand NAND2_13110 ( P1_R1162_U249 , P1_R1162_U222 , P1_R1162_U42 );
nand NAND2_13111 ( P1_R1162_U250 , P1_R1162_U248 , P1_R1162_U137 );
nand NAND2_13112 ( P1_R1162_U251 , P1_U3466 , P1_R1162_U30 );
nand NAND2_13113 ( P1_R1162_U252 , P1_REG1_REG_3_ , P1_R1162_U31 );
nand NAND2_13114 ( P1_R1162_U253 , P1_R1162_U252 , P1_R1162_U251 );
nand NAND2_13115 ( P1_R1162_U254 , P1_R1162_U223 , P1_R1162_U82 );
nand NAND2_13116 ( P1_R1162_U255 , P1_R1162_U146 , P1_R1162_U253 );
nand NAND2_13117 ( P1_R1162_U256 , P1_U3463 , P1_R1162_U25 );
nand NAND2_13118 ( P1_R1162_U257 , P1_REG1_REG_2_ , P1_R1162_U26 );
nand NAND2_13119 ( P1_R1162_U258 , P1_R1162_U98 , P1_R1162_U83 );
nand NAND2_13120 ( P1_R1162_U259 , P1_R1162_U153 , P1_R1162_U29 );
nand NAND2_13121 ( P1_R1162_U260 , P1_U3452 , P1_R1162_U85 );
nand NAND2_13122 ( P1_R1162_U261 , P1_REG1_REG_19_ , P1_R1162_U84 );
nand NAND2_13123 ( P1_R1162_U262 , P1_U3452 , P1_R1162_U85 );
nand NAND2_13124 ( P1_R1162_U263 , P1_REG1_REG_19_ , P1_R1162_U84 );
nand NAND2_13125 ( P1_R1162_U264 , P1_R1162_U263 , P1_R1162_U262 );
nand NAND2_13126 ( P1_R1162_U265 , P1_U3511 , P1_R1162_U63 );
nand NAND2_13127 ( P1_R1162_U266 , P1_REG1_REG_18_ , P1_R1162_U64 );
nand NAND2_13128 ( P1_R1162_U267 , P1_U3511 , P1_R1162_U63 );
nand NAND2_13129 ( P1_R1162_U268 , P1_REG1_REG_18_ , P1_R1162_U64 );
nand NAND2_13130 ( P1_R1162_U269 , P1_R1162_U268 , P1_R1162_U267 );
nand NAND3_13131 ( P1_R1162_U270 , P1_R1162_U266 , P1_R1162_U265 , P1_R1162_U65 );
nand NAND2_13132 ( P1_R1162_U271 , P1_R1162_U269 , P1_R1162_U188 );
nand NAND2_13133 ( P1_R1162_U272 , P1_U3508 , P1_R1162_U48 );
nand NAND2_13134 ( P1_R1162_U273 , P1_REG1_REG_17_ , P1_R1162_U46 );
nand NAND2_13135 ( P1_R1162_U274 , P1_U3505 , P1_R1162_U44 );
nand NAND2_13136 ( P1_R1162_U275 , P1_REG1_REG_16_ , P1_R1162_U45 );
nand NAND2_13137 ( P1_R1162_U276 , P1_R1162_U275 , P1_R1162_U274 );
nand NAND2_13138 ( P1_R1162_U277 , P1_R1162_U224 , P1_R1162_U66 );
nand NAND2_13139 ( P1_R1162_U278 , P1_R1162_U276 , P1_R1162_U180 );
nand NAND2_13140 ( P1_R1162_U279 , P1_U3502 , P1_R1162_U61 );
nand NAND2_13141 ( P1_R1162_U280 , P1_REG1_REG_15_ , P1_R1162_U62 );
nand NAND2_13142 ( P1_R1162_U281 , P1_U3502 , P1_R1162_U61 );
nand NAND2_13143 ( P1_R1162_U282 , P1_REG1_REG_15_ , P1_R1162_U62 );
nand NAND2_13144 ( P1_R1162_U283 , P1_R1162_U282 , P1_R1162_U281 );
nand NAND3_13145 ( P1_R1162_U284 , P1_R1162_U280 , P1_R1162_U279 , P1_R1162_U86 );
nand NAND2_13146 ( P1_R1162_U285 , P1_R1162_U176 , P1_R1162_U283 );
nand NAND2_13147 ( P1_R1162_U286 , P1_U3499 , P1_R1162_U59 );
nand NAND2_13148 ( P1_R1162_U287 , P1_REG1_REG_14_ , P1_R1162_U60 );
nand NAND2_13149 ( P1_R1162_U288 , P1_U3499 , P1_R1162_U59 );
nand NAND2_13150 ( P1_R1162_U289 , P1_REG1_REG_14_ , P1_R1162_U60 );
nand NAND2_13151 ( P1_R1162_U290 , P1_R1162_U289 , P1_R1162_U288 );
nand NAND3_13152 ( P1_R1162_U291 , P1_R1162_U287 , P1_R1162_U286 , P1_R1162_U87 );
nand NAND2_13153 ( P1_R1162_U292 , P1_R1162_U172 , P1_R1162_U290 );
nand NAND2_13154 ( P1_R1162_U293 , P1_U3496 , P1_R1162_U57 );
nand NAND2_13155 ( P1_R1162_U294 , P1_REG1_REG_13_ , P1_R1162_U58 );
nand NAND2_13156 ( P1_R1162_U295 , P1_U3493 , P1_R1162_U52 );
nand NAND2_13157 ( P1_R1162_U296 , P1_REG1_REG_12_ , P1_R1162_U53 );
nand NAND2_13158 ( P1_R1162_U297 , P1_R1162_U296 , P1_R1162_U295 );
nand NAND2_13159 ( P1_R1162_U298 , P1_R1162_U225 , P1_R1162_U67 );
nand NAND2_13160 ( P1_R1162_U299 , P1_R1162_U297 , P1_R1162_U205 );
nand NAND2_13161 ( P1_R1162_U300 , P1_U3490 , P1_R1162_U54 );
nand NAND2_13162 ( P1_R1162_U301 , P1_REG1_REG_11_ , P1_R1162_U55 );
nand NAND2_13163 ( P1_R1162_U302 , P1_R1162_U301 , P1_R1162_U300 );
nand NAND2_13164 ( P1_R1162_U303 , P1_R1162_U226 , P1_R1162_U88 );
nand NAND2_13165 ( P1_R1162_U304 , P1_R1162_U162 , P1_R1162_U302 );
nand NAND2_13166 ( P1_R1162_U305 , P1_U3487 , P1_R1162_U50 );
nand NAND2_13167 ( P1_R1162_U306 , P1_REG1_REG_10_ , P1_R1162_U51 );
nand NAND2_13168 ( P1_R1162_U307 , P1_U3454 , P1_R1162_U27 );
nand NAND2_13169 ( P1_R1162_U308 , P1_REG1_REG_0_ , P1_R1162_U28 );
and AND2_13170 ( P1_R1117_U6 , P1_R1117_U184 , P1_R1117_U201 );
and AND2_13171 ( P1_R1117_U7 , P1_R1117_U203 , P1_R1117_U202 );
and AND2_13172 ( P1_R1117_U8 , P1_R1117_U179 , P1_R1117_U240 );
and AND2_13173 ( P1_R1117_U9 , P1_R1117_U242 , P1_R1117_U241 );
and AND2_13174 ( P1_R1117_U10 , P1_R1117_U259 , P1_R1117_U258 );
and AND2_13175 ( P1_R1117_U11 , P1_R1117_U285 , P1_R1117_U284 );
and AND2_13176 ( P1_R1117_U12 , P1_R1117_U383 , P1_R1117_U382 );
nand NAND2_13177 ( P1_R1117_U13 , P1_R1117_U340 , P1_R1117_U343 );
nand NAND2_13178 ( P1_R1117_U14 , P1_R1117_U329 , P1_R1117_U332 );
nand NAND2_13179 ( P1_R1117_U15 , P1_R1117_U318 , P1_R1117_U321 );
nand NAND2_13180 ( P1_R1117_U16 , P1_R1117_U310 , P1_R1117_U312 );
nand NAND3_13181 ( P1_R1117_U17 , P1_R1117_U156 , P1_R1117_U175 , P1_R1117_U348 );
nand NAND2_13182 ( P1_R1117_U18 , P1_R1117_U236 , P1_R1117_U238 );
nand NAND2_13183 ( P1_R1117_U19 , P1_R1117_U228 , P1_R1117_U231 );
nand NAND2_13184 ( P1_R1117_U20 , P1_R1117_U220 , P1_R1117_U222 );
nand NAND2_13185 ( P1_R1117_U21 , P1_R1117_U25 , P1_R1117_U346 );
not NOT1_13186 ( P1_R1117_U22 , P1_U3479 );
not NOT1_13187 ( P1_R1117_U23 , P1_U3464 );
not NOT1_13188 ( P1_R1117_U24 , P1_U3456 );
nand NAND2_13189 ( P1_R1117_U25 , P1_U3456 , P1_R1117_U93 );
not NOT1_13190 ( P1_R1117_U26 , P1_U3078 );
not NOT1_13191 ( P1_R1117_U27 , P1_U3467 );
not NOT1_13192 ( P1_R1117_U28 , P1_U3068 );
nand NAND2_13193 ( P1_R1117_U29 , P1_U3068 , P1_R1117_U23 );
not NOT1_13194 ( P1_R1117_U30 , P1_U3064 );
not NOT1_13195 ( P1_R1117_U31 , P1_U3476 );
not NOT1_13196 ( P1_R1117_U32 , P1_U3473 );
not NOT1_13197 ( P1_R1117_U33 , P1_U3470 );
not NOT1_13198 ( P1_R1117_U34 , P1_U3071 );
not NOT1_13199 ( P1_R1117_U35 , P1_U3067 );
not NOT1_13200 ( P1_R1117_U36 , P1_U3060 );
nand NAND2_13201 ( P1_R1117_U37 , P1_U3060 , P1_R1117_U33 );
not NOT1_13202 ( P1_R1117_U38 , P1_U3482 );
not NOT1_13203 ( P1_R1117_U39 , P1_U3070 );
nand NAND2_13204 ( P1_R1117_U40 , P1_U3070 , P1_R1117_U22 );
not NOT1_13205 ( P1_R1117_U41 , P1_U3084 );
not NOT1_13206 ( P1_R1117_U42 , P1_U3485 );
not NOT1_13207 ( P1_R1117_U43 , P1_U3083 );
nand NAND2_13208 ( P1_R1117_U44 , P1_R1117_U209 , P1_R1117_U208 );
nand NAND2_13209 ( P1_R1117_U45 , P1_R1117_U37 , P1_R1117_U224 );
nand NAND2_13210 ( P1_R1117_U46 , P1_R1117_U193 , P1_R1117_U192 );
not NOT1_13211 ( P1_R1117_U47 , P1_U4019 );
not NOT1_13212 ( P1_R1117_U48 , P1_U4023 );
not NOT1_13213 ( P1_R1117_U49 , P1_U3503 );
not NOT1_13214 ( P1_R1117_U50 , P1_U3491 );
not NOT1_13215 ( P1_R1117_U51 , P1_U3488 );
not NOT1_13216 ( P1_R1117_U52 , P1_U3063 );
not NOT1_13217 ( P1_R1117_U53 , P1_U3062 );
nand NAND2_13218 ( P1_R1117_U54 , P1_U3083 , P1_R1117_U42 );
not NOT1_13219 ( P1_R1117_U55 , P1_U3494 );
not NOT1_13220 ( P1_R1117_U56 , P1_U3072 );
not NOT1_13221 ( P1_R1117_U57 , P1_U3497 );
not NOT1_13222 ( P1_R1117_U58 , P1_U3080 );
not NOT1_13223 ( P1_R1117_U59 , P1_U3506 );
not NOT1_13224 ( P1_R1117_U60 , P1_U3500 );
not NOT1_13225 ( P1_R1117_U61 , P1_U3073 );
not NOT1_13226 ( P1_R1117_U62 , P1_U3074 );
not NOT1_13227 ( P1_R1117_U63 , P1_U3079 );
nand NAND2_13228 ( P1_R1117_U64 , P1_U3079 , P1_R1117_U60 );
not NOT1_13229 ( P1_R1117_U65 , P1_U3509 );
not NOT1_13230 ( P1_R1117_U66 , P1_U3069 );
nand NAND2_13231 ( P1_R1117_U67 , P1_R1117_U269 , P1_R1117_U268 );
not NOT1_13232 ( P1_R1117_U68 , P1_U3082 );
not NOT1_13233 ( P1_R1117_U69 , P1_U3514 );
not NOT1_13234 ( P1_R1117_U70 , P1_U3081 );
not NOT1_13235 ( P1_R1117_U71 , P1_U4025 );
not NOT1_13236 ( P1_R1117_U72 , P1_U3076 );
not NOT1_13237 ( P1_R1117_U73 , P1_U4022 );
not NOT1_13238 ( P1_R1117_U74 , P1_U4024 );
not NOT1_13239 ( P1_R1117_U75 , P1_U3066 );
not NOT1_13240 ( P1_R1117_U76 , P1_U3061 );
not NOT1_13241 ( P1_R1117_U77 , P1_U3075 );
nand NAND2_13242 ( P1_R1117_U78 , P1_U3075 , P1_R1117_U74 );
not NOT1_13243 ( P1_R1117_U79 , P1_U4021 );
not NOT1_13244 ( P1_R1117_U80 , P1_U3065 );
not NOT1_13245 ( P1_R1117_U81 , P1_U4020 );
not NOT1_13246 ( P1_R1117_U82 , P1_U3058 );
not NOT1_13247 ( P1_R1117_U83 , P1_U4018 );
not NOT1_13248 ( P1_R1117_U84 , P1_U3057 );
nand NAND2_13249 ( P1_R1117_U85 , P1_U3057 , P1_R1117_U47 );
not NOT1_13250 ( P1_R1117_U86 , P1_U3053 );
not NOT1_13251 ( P1_R1117_U87 , P1_U4017 );
not NOT1_13252 ( P1_R1117_U88 , P1_U3054 );
nand NAND2_13253 ( P1_R1117_U89 , P1_R1117_U299 , P1_R1117_U298 );
nand NAND2_13254 ( P1_R1117_U90 , P1_R1117_U78 , P1_R1117_U314 );
nand NAND2_13255 ( P1_R1117_U91 , P1_R1117_U64 , P1_R1117_U325 );
nand NAND2_13256 ( P1_R1117_U92 , P1_R1117_U54 , P1_R1117_U336 );
not NOT1_13257 ( P1_R1117_U93 , P1_U3077 );
nand NAND2_13258 ( P1_R1117_U94 , P1_R1117_U393 , P1_R1117_U392 );
nand NAND2_13259 ( P1_R1117_U95 , P1_R1117_U407 , P1_R1117_U406 );
nand NAND2_13260 ( P1_R1117_U96 , P1_R1117_U412 , P1_R1117_U411 );
nand NAND2_13261 ( P1_R1117_U97 , P1_R1117_U428 , P1_R1117_U427 );
nand NAND2_13262 ( P1_R1117_U98 , P1_R1117_U433 , P1_R1117_U432 );
nand NAND2_13263 ( P1_R1117_U99 , P1_R1117_U438 , P1_R1117_U437 );
nand NAND2_13264 ( P1_R1117_U100 , P1_R1117_U443 , P1_R1117_U442 );
nand NAND2_13265 ( P1_R1117_U101 , P1_R1117_U448 , P1_R1117_U447 );
nand NAND2_13266 ( P1_R1117_U102 , P1_R1117_U464 , P1_R1117_U463 );
nand NAND2_13267 ( P1_R1117_U103 , P1_R1117_U469 , P1_R1117_U468 );
nand NAND2_13268 ( P1_R1117_U104 , P1_R1117_U352 , P1_R1117_U351 );
nand NAND2_13269 ( P1_R1117_U105 , P1_R1117_U361 , P1_R1117_U360 );
nand NAND2_13270 ( P1_R1117_U106 , P1_R1117_U368 , P1_R1117_U367 );
nand NAND2_13271 ( P1_R1117_U107 , P1_R1117_U372 , P1_R1117_U371 );
nand NAND2_13272 ( P1_R1117_U108 , P1_R1117_U381 , P1_R1117_U380 );
nand NAND2_13273 ( P1_R1117_U109 , P1_R1117_U402 , P1_R1117_U401 );
nand NAND2_13274 ( P1_R1117_U110 , P1_R1117_U419 , P1_R1117_U418 );
nand NAND2_13275 ( P1_R1117_U111 , P1_R1117_U423 , P1_R1117_U422 );
nand NAND2_13276 ( P1_R1117_U112 , P1_R1117_U455 , P1_R1117_U454 );
nand NAND2_13277 ( P1_R1117_U113 , P1_R1117_U459 , P1_R1117_U458 );
nand NAND2_13278 ( P1_R1117_U114 , P1_R1117_U476 , P1_R1117_U475 );
and AND2_13279 ( P1_R1117_U115 , P1_R1117_U195 , P1_R1117_U183 );
and AND2_13280 ( P1_R1117_U116 , P1_R1117_U198 , P1_R1117_U199 );
and AND2_13281 ( P1_R1117_U117 , P1_R1117_U211 , P1_R1117_U185 );
and AND2_13282 ( P1_R1117_U118 , P1_R1117_U214 , P1_R1117_U215 );
and AND3_13283 ( P1_R1117_U119 , P1_R1117_U354 , P1_R1117_U353 , P1_R1117_U40 );
and AND2_13284 ( P1_R1117_U120 , P1_R1117_U357 , P1_R1117_U185 );
and AND2_13285 ( P1_R1117_U121 , P1_R1117_U230 , P1_R1117_U7 );
and AND2_13286 ( P1_R1117_U122 , P1_R1117_U364 , P1_R1117_U184 );
and AND3_13287 ( P1_R1117_U123 , P1_R1117_U374 , P1_R1117_U373 , P1_R1117_U29 );
and AND2_13288 ( P1_R1117_U124 , P1_R1117_U377 , P1_R1117_U183 );
and AND2_13289 ( P1_R1117_U125 , P1_R1117_U217 , P1_R1117_U8 );
and AND2_13290 ( P1_R1117_U126 , P1_R1117_U262 , P1_R1117_U180 );
and AND2_13291 ( P1_R1117_U127 , P1_R1117_U288 , P1_R1117_U181 );
and AND2_13292 ( P1_R1117_U128 , P1_R1117_U304 , P1_R1117_U305 );
and AND2_13293 ( P1_R1117_U129 , P1_R1117_U307 , P1_R1117_U386 );
and AND3_13294 ( P1_R1117_U130 , P1_R1117_U305 , P1_R1117_U304 , P1_R1117_U308 );
nand NAND2_13295 ( P1_R1117_U131 , P1_R1117_U390 , P1_R1117_U389 );
and AND3_13296 ( P1_R1117_U132 , P1_R1117_U395 , P1_R1117_U394 , P1_R1117_U85 );
and AND2_13297 ( P1_R1117_U133 , P1_R1117_U398 , P1_R1117_U182 );
nand NAND2_13298 ( P1_R1117_U134 , P1_R1117_U404 , P1_R1117_U403 );
nand NAND2_13299 ( P1_R1117_U135 , P1_R1117_U409 , P1_R1117_U408 );
and AND2_13300 ( P1_R1117_U136 , P1_R1117_U415 , P1_R1117_U181 );
nand NAND2_13301 ( P1_R1117_U137 , P1_R1117_U425 , P1_R1117_U424 );
nand NAND2_13302 ( P1_R1117_U138 , P1_R1117_U430 , P1_R1117_U429 );
nand NAND2_13303 ( P1_R1117_U139 , P1_R1117_U435 , P1_R1117_U434 );
nand NAND2_13304 ( P1_R1117_U140 , P1_R1117_U440 , P1_R1117_U439 );
nand NAND2_13305 ( P1_R1117_U141 , P1_R1117_U445 , P1_R1117_U444 );
and AND2_13306 ( P1_R1117_U142 , P1_R1117_U451 , P1_R1117_U180 );
nand NAND2_13307 ( P1_R1117_U143 , P1_R1117_U461 , P1_R1117_U460 );
nand NAND2_13308 ( P1_R1117_U144 , P1_R1117_U466 , P1_R1117_U465 );
and AND2_13309 ( P1_R1117_U145 , P1_R1117_U342 , P1_R1117_U9 );
and AND2_13310 ( P1_R1117_U146 , P1_R1117_U472 , P1_R1117_U179 );
and AND2_13311 ( P1_R1117_U147 , P1_R1117_U350 , P1_R1117_U349 );
nand NAND2_13312 ( P1_R1117_U148 , P1_R1117_U118 , P1_R1117_U212 );
and AND2_13313 ( P1_R1117_U149 , P1_R1117_U359 , P1_R1117_U358 );
and AND2_13314 ( P1_R1117_U150 , P1_R1117_U366 , P1_R1117_U365 );
and AND2_13315 ( P1_R1117_U151 , P1_R1117_U370 , P1_R1117_U369 );
nand NAND2_13316 ( P1_R1117_U152 , P1_R1117_U116 , P1_R1117_U196 );
and AND2_13317 ( P1_R1117_U153 , P1_R1117_U379 , P1_R1117_U378 );
not NOT1_13318 ( P1_R1117_U154 , P1_U4028 );
not NOT1_13319 ( P1_R1117_U155 , P1_U3055 );
and AND2_13320 ( P1_R1117_U156 , P1_R1117_U388 , P1_R1117_U387 );
nand NAND2_13321 ( P1_R1117_U157 , P1_R1117_U128 , P1_R1117_U302 );
and AND2_13322 ( P1_R1117_U158 , P1_R1117_U400 , P1_R1117_U399 );
nand NAND2_13323 ( P1_R1117_U159 , P1_R1117_U295 , P1_R1117_U294 );
nand NAND2_13324 ( P1_R1117_U160 , P1_R1117_U291 , P1_R1117_U290 );
and AND2_13325 ( P1_R1117_U161 , P1_R1117_U417 , P1_R1117_U416 );
and AND2_13326 ( P1_R1117_U162 , P1_R1117_U421 , P1_R1117_U420 );
nand NAND2_13327 ( P1_R1117_U163 , P1_R1117_U281 , P1_R1117_U280 );
nand NAND2_13328 ( P1_R1117_U164 , P1_R1117_U277 , P1_R1117_U276 );
not NOT1_13329 ( P1_R1117_U165 , P1_U3461 );
nand NAND2_13330 ( P1_R1117_U166 , P1_R1117_U273 , P1_R1117_U272 );
not NOT1_13331 ( P1_R1117_U167 , P1_U3512 );
nand NAND2_13332 ( P1_R1117_U168 , P1_R1117_U265 , P1_R1117_U264 );
and AND2_13333 ( P1_R1117_U169 , P1_R1117_U453 , P1_R1117_U452 );
and AND2_13334 ( P1_R1117_U170 , P1_R1117_U457 , P1_R1117_U456 );
nand NAND2_13335 ( P1_R1117_U171 , P1_R1117_U255 , P1_R1117_U254 );
nand NAND2_13336 ( P1_R1117_U172 , P1_R1117_U251 , P1_R1117_U250 );
nand NAND2_13337 ( P1_R1117_U173 , P1_R1117_U247 , P1_R1117_U246 );
and AND2_13338 ( P1_R1117_U174 , P1_R1117_U474 , P1_R1117_U473 );
nand NAND2_13339 ( P1_R1117_U175 , P1_R1117_U129 , P1_R1117_U157 );
not NOT1_13340 ( P1_R1117_U176 , P1_R1117_U85 );
not NOT1_13341 ( P1_R1117_U177 , P1_R1117_U29 );
not NOT1_13342 ( P1_R1117_U178 , P1_R1117_U40 );
nand NAND2_13343 ( P1_R1117_U179 , P1_U3488 , P1_R1117_U53 );
nand NAND2_13344 ( P1_R1117_U180 , P1_U3503 , P1_R1117_U62 );
nand NAND2_13345 ( P1_R1117_U181 , P1_U4023 , P1_R1117_U76 );
nand NAND2_13346 ( P1_R1117_U182 , P1_U4019 , P1_R1117_U84 );
nand NAND2_13347 ( P1_R1117_U183 , P1_U3464 , P1_R1117_U28 );
nand NAND2_13348 ( P1_R1117_U184 , P1_U3473 , P1_R1117_U35 );
nand NAND2_13349 ( P1_R1117_U185 , P1_U3479 , P1_R1117_U39 );
not NOT1_13350 ( P1_R1117_U186 , P1_R1117_U64 );
not NOT1_13351 ( P1_R1117_U187 , P1_R1117_U78 );
not NOT1_13352 ( P1_R1117_U188 , P1_R1117_U37 );
not NOT1_13353 ( P1_R1117_U189 , P1_R1117_U54 );
not NOT1_13354 ( P1_R1117_U190 , P1_R1117_U25 );
nand NAND2_13355 ( P1_R1117_U191 , P1_R1117_U190 , P1_R1117_U26 );
nand NAND2_13356 ( P1_R1117_U192 , P1_R1117_U191 , P1_R1117_U165 );
nand NAND2_13357 ( P1_R1117_U193 , P1_U3078 , P1_R1117_U25 );
not NOT1_13358 ( P1_R1117_U194 , P1_R1117_U46 );
nand NAND2_13359 ( P1_R1117_U195 , P1_U3467 , P1_R1117_U30 );
nand NAND2_13360 ( P1_R1117_U196 , P1_R1117_U115 , P1_R1117_U46 );
nand NAND2_13361 ( P1_R1117_U197 , P1_R1117_U30 , P1_R1117_U29 );
nand NAND2_13362 ( P1_R1117_U198 , P1_R1117_U197 , P1_R1117_U27 );
nand NAND2_13363 ( P1_R1117_U199 , P1_U3064 , P1_R1117_U177 );
not NOT1_13364 ( P1_R1117_U200 , P1_R1117_U152 );
nand NAND2_13365 ( P1_R1117_U201 , P1_U3476 , P1_R1117_U34 );
nand NAND2_13366 ( P1_R1117_U202 , P1_U3071 , P1_R1117_U31 );
nand NAND2_13367 ( P1_R1117_U203 , P1_U3067 , P1_R1117_U32 );
nand NAND2_13368 ( P1_R1117_U204 , P1_R1117_U188 , P1_R1117_U6 );
nand NAND2_13369 ( P1_R1117_U205 , P1_R1117_U7 , P1_R1117_U204 );
nand NAND2_13370 ( P1_R1117_U206 , P1_U3470 , P1_R1117_U36 );
nand NAND2_13371 ( P1_R1117_U207 , P1_U3476 , P1_R1117_U34 );
nand NAND3_13372 ( P1_R1117_U208 , P1_R1117_U206 , P1_R1117_U152 , P1_R1117_U6 );
nand NAND2_13373 ( P1_R1117_U209 , P1_R1117_U207 , P1_R1117_U205 );
not NOT1_13374 ( P1_R1117_U210 , P1_R1117_U44 );
nand NAND2_13375 ( P1_R1117_U211 , P1_U3482 , P1_R1117_U41 );
nand NAND2_13376 ( P1_R1117_U212 , P1_R1117_U117 , P1_R1117_U44 );
nand NAND2_13377 ( P1_R1117_U213 , P1_R1117_U41 , P1_R1117_U40 );
nand NAND2_13378 ( P1_R1117_U214 , P1_R1117_U213 , P1_R1117_U38 );
nand NAND2_13379 ( P1_R1117_U215 , P1_U3084 , P1_R1117_U178 );
not NOT1_13380 ( P1_R1117_U216 , P1_R1117_U148 );
nand NAND2_13381 ( P1_R1117_U217 , P1_U3485 , P1_R1117_U43 );
nand NAND2_13382 ( P1_R1117_U218 , P1_R1117_U217 , P1_R1117_U54 );
nand NAND2_13383 ( P1_R1117_U219 , P1_R1117_U210 , P1_R1117_U40 );
nand NAND2_13384 ( P1_R1117_U220 , P1_R1117_U120 , P1_R1117_U219 );
nand NAND2_13385 ( P1_R1117_U221 , P1_R1117_U44 , P1_R1117_U185 );
nand NAND2_13386 ( P1_R1117_U222 , P1_R1117_U119 , P1_R1117_U221 );
nand NAND2_13387 ( P1_R1117_U223 , P1_R1117_U40 , P1_R1117_U185 );
nand NAND2_13388 ( P1_R1117_U224 , P1_R1117_U206 , P1_R1117_U152 );
not NOT1_13389 ( P1_R1117_U225 , P1_R1117_U45 );
nand NAND2_13390 ( P1_R1117_U226 , P1_U3067 , P1_R1117_U32 );
nand NAND2_13391 ( P1_R1117_U227 , P1_R1117_U225 , P1_R1117_U226 );
nand NAND2_13392 ( P1_R1117_U228 , P1_R1117_U122 , P1_R1117_U227 );
nand NAND2_13393 ( P1_R1117_U229 , P1_R1117_U45 , P1_R1117_U184 );
nand NAND2_13394 ( P1_R1117_U230 , P1_U3476 , P1_R1117_U34 );
nand NAND2_13395 ( P1_R1117_U231 , P1_R1117_U121 , P1_R1117_U229 );
nand NAND2_13396 ( P1_R1117_U232 , P1_U3067 , P1_R1117_U32 );
nand NAND2_13397 ( P1_R1117_U233 , P1_R1117_U184 , P1_R1117_U232 );
nand NAND2_13398 ( P1_R1117_U234 , P1_R1117_U206 , P1_R1117_U37 );
nand NAND2_13399 ( P1_R1117_U235 , P1_R1117_U194 , P1_R1117_U29 );
nand NAND2_13400 ( P1_R1117_U236 , P1_R1117_U124 , P1_R1117_U235 );
nand NAND2_13401 ( P1_R1117_U237 , P1_R1117_U46 , P1_R1117_U183 );
nand NAND2_13402 ( P1_R1117_U238 , P1_R1117_U123 , P1_R1117_U237 );
nand NAND2_13403 ( P1_R1117_U239 , P1_R1117_U29 , P1_R1117_U183 );
nand NAND2_13404 ( P1_R1117_U240 , P1_U3491 , P1_R1117_U52 );
nand NAND2_13405 ( P1_R1117_U241 , P1_U3063 , P1_R1117_U50 );
nand NAND2_13406 ( P1_R1117_U242 , P1_U3062 , P1_R1117_U51 );
nand NAND2_13407 ( P1_R1117_U243 , P1_R1117_U189 , P1_R1117_U8 );
nand NAND2_13408 ( P1_R1117_U244 , P1_R1117_U9 , P1_R1117_U243 );
nand NAND2_13409 ( P1_R1117_U245 , P1_U3491 , P1_R1117_U52 );
nand NAND2_13410 ( P1_R1117_U246 , P1_R1117_U125 , P1_R1117_U148 );
nand NAND2_13411 ( P1_R1117_U247 , P1_R1117_U245 , P1_R1117_U244 );
not NOT1_13412 ( P1_R1117_U248 , P1_R1117_U173 );
nand NAND2_13413 ( P1_R1117_U249 , P1_U3494 , P1_R1117_U56 );
nand NAND2_13414 ( P1_R1117_U250 , P1_R1117_U249 , P1_R1117_U173 );
nand NAND2_13415 ( P1_R1117_U251 , P1_U3072 , P1_R1117_U55 );
not NOT1_13416 ( P1_R1117_U252 , P1_R1117_U172 );
nand NAND2_13417 ( P1_R1117_U253 , P1_U3497 , P1_R1117_U58 );
nand NAND2_13418 ( P1_R1117_U254 , P1_R1117_U253 , P1_R1117_U172 );
nand NAND2_13419 ( P1_R1117_U255 , P1_U3080 , P1_R1117_U57 );
not NOT1_13420 ( P1_R1117_U256 , P1_R1117_U171 );
nand NAND2_13421 ( P1_R1117_U257 , P1_U3506 , P1_R1117_U61 );
nand NAND2_13422 ( P1_R1117_U258 , P1_U3073 , P1_R1117_U59 );
nand NAND2_13423 ( P1_R1117_U259 , P1_U3074 , P1_R1117_U49 );
nand NAND2_13424 ( P1_R1117_U260 , P1_R1117_U186 , P1_R1117_U180 );
nand NAND2_13425 ( P1_R1117_U261 , P1_R1117_U10 , P1_R1117_U260 );
nand NAND2_13426 ( P1_R1117_U262 , P1_U3500 , P1_R1117_U63 );
nand NAND2_13427 ( P1_R1117_U263 , P1_U3506 , P1_R1117_U61 );
nand NAND3_13428 ( P1_R1117_U264 , P1_R1117_U171 , P1_R1117_U126 , P1_R1117_U257 );
nand NAND2_13429 ( P1_R1117_U265 , P1_R1117_U263 , P1_R1117_U261 );
not NOT1_13430 ( P1_R1117_U266 , P1_R1117_U168 );
nand NAND2_13431 ( P1_R1117_U267 , P1_U3509 , P1_R1117_U66 );
nand NAND2_13432 ( P1_R1117_U268 , P1_R1117_U267 , P1_R1117_U168 );
nand NAND2_13433 ( P1_R1117_U269 , P1_U3069 , P1_R1117_U65 );
not NOT1_13434 ( P1_R1117_U270 , P1_R1117_U67 );
nand NAND2_13435 ( P1_R1117_U271 , P1_R1117_U270 , P1_R1117_U68 );
nand NAND2_13436 ( P1_R1117_U272 , P1_R1117_U271 , P1_R1117_U167 );
nand NAND2_13437 ( P1_R1117_U273 , P1_U3082 , P1_R1117_U67 );
not NOT1_13438 ( P1_R1117_U274 , P1_R1117_U166 );
nand NAND2_13439 ( P1_R1117_U275 , P1_U3514 , P1_R1117_U70 );
nand NAND2_13440 ( P1_R1117_U276 , P1_R1117_U275 , P1_R1117_U166 );
nand NAND2_13441 ( P1_R1117_U277 , P1_U3081 , P1_R1117_U69 );
not NOT1_13442 ( P1_R1117_U278 , P1_R1117_U164 );
nand NAND2_13443 ( P1_R1117_U279 , P1_U4025 , P1_R1117_U72 );
nand NAND2_13444 ( P1_R1117_U280 , P1_R1117_U279 , P1_R1117_U164 );
nand NAND2_13445 ( P1_R1117_U281 , P1_U3076 , P1_R1117_U71 );
not NOT1_13446 ( P1_R1117_U282 , P1_R1117_U163 );
nand NAND2_13447 ( P1_R1117_U283 , P1_U4022 , P1_R1117_U75 );
nand NAND2_13448 ( P1_R1117_U284 , P1_U3066 , P1_R1117_U73 );
nand NAND2_13449 ( P1_R1117_U285 , P1_U3061 , P1_R1117_U48 );
nand NAND2_13450 ( P1_R1117_U286 , P1_R1117_U187 , P1_R1117_U181 );
nand NAND2_13451 ( P1_R1117_U287 , P1_R1117_U11 , P1_R1117_U286 );
nand NAND2_13452 ( P1_R1117_U288 , P1_U4024 , P1_R1117_U77 );
nand NAND2_13453 ( P1_R1117_U289 , P1_U4022 , P1_R1117_U75 );
nand NAND3_13454 ( P1_R1117_U290 , P1_R1117_U163 , P1_R1117_U127 , P1_R1117_U283 );
nand NAND2_13455 ( P1_R1117_U291 , P1_R1117_U289 , P1_R1117_U287 );
not NOT1_13456 ( P1_R1117_U292 , P1_R1117_U160 );
nand NAND2_13457 ( P1_R1117_U293 , P1_U4021 , P1_R1117_U80 );
nand NAND2_13458 ( P1_R1117_U294 , P1_R1117_U293 , P1_R1117_U160 );
nand NAND2_13459 ( P1_R1117_U295 , P1_U3065 , P1_R1117_U79 );
not NOT1_13460 ( P1_R1117_U296 , P1_R1117_U159 );
nand NAND2_13461 ( P1_R1117_U297 , P1_U4020 , P1_R1117_U82 );
nand NAND2_13462 ( P1_R1117_U298 , P1_R1117_U297 , P1_R1117_U159 );
nand NAND2_13463 ( P1_R1117_U299 , P1_U3058 , P1_R1117_U81 );
not NOT1_13464 ( P1_R1117_U300 , P1_R1117_U89 );
nand NAND2_13465 ( P1_R1117_U301 , P1_U4018 , P1_R1117_U86 );
nand NAND3_13466 ( P1_R1117_U302 , P1_R1117_U89 , P1_R1117_U182 , P1_R1117_U301 );
nand NAND2_13467 ( P1_R1117_U303 , P1_R1117_U86 , P1_R1117_U85 );
nand NAND2_13468 ( P1_R1117_U304 , P1_R1117_U303 , P1_R1117_U83 );
nand NAND2_13469 ( P1_R1117_U305 , P1_U3053 , P1_R1117_U176 );
not NOT1_13470 ( P1_R1117_U306 , P1_R1117_U157 );
nand NAND2_13471 ( P1_R1117_U307 , P1_U4017 , P1_R1117_U88 );
nand NAND2_13472 ( P1_R1117_U308 , P1_U3054 , P1_R1117_U87 );
nand NAND2_13473 ( P1_R1117_U309 , P1_R1117_U300 , P1_R1117_U85 );
nand NAND2_13474 ( P1_R1117_U310 , P1_R1117_U133 , P1_R1117_U309 );
nand NAND2_13475 ( P1_R1117_U311 , P1_R1117_U89 , P1_R1117_U182 );
nand NAND2_13476 ( P1_R1117_U312 , P1_R1117_U132 , P1_R1117_U311 );
nand NAND2_13477 ( P1_R1117_U313 , P1_R1117_U85 , P1_R1117_U182 );
nand NAND2_13478 ( P1_R1117_U314 , P1_R1117_U288 , P1_R1117_U163 );
not NOT1_13479 ( P1_R1117_U315 , P1_R1117_U90 );
nand NAND2_13480 ( P1_R1117_U316 , P1_U3061 , P1_R1117_U48 );
nand NAND2_13481 ( P1_R1117_U317 , P1_R1117_U315 , P1_R1117_U316 );
nand NAND2_13482 ( P1_R1117_U318 , P1_R1117_U136 , P1_R1117_U317 );
nand NAND2_13483 ( P1_R1117_U319 , P1_R1117_U90 , P1_R1117_U181 );
nand NAND2_13484 ( P1_R1117_U320 , P1_U4022 , P1_R1117_U75 );
nand NAND3_13485 ( P1_R1117_U321 , P1_R1117_U320 , P1_R1117_U319 , P1_R1117_U11 );
nand NAND2_13486 ( P1_R1117_U322 , P1_U3061 , P1_R1117_U48 );
nand NAND2_13487 ( P1_R1117_U323 , P1_R1117_U181 , P1_R1117_U322 );
nand NAND2_13488 ( P1_R1117_U324 , P1_R1117_U288 , P1_R1117_U78 );
nand NAND2_13489 ( P1_R1117_U325 , P1_R1117_U262 , P1_R1117_U171 );
not NOT1_13490 ( P1_R1117_U326 , P1_R1117_U91 );
nand NAND2_13491 ( P1_R1117_U327 , P1_U3074 , P1_R1117_U49 );
nand NAND2_13492 ( P1_R1117_U328 , P1_R1117_U326 , P1_R1117_U327 );
nand NAND2_13493 ( P1_R1117_U329 , P1_R1117_U142 , P1_R1117_U328 );
nand NAND2_13494 ( P1_R1117_U330 , P1_R1117_U91 , P1_R1117_U180 );
nand NAND2_13495 ( P1_R1117_U331 , P1_U3506 , P1_R1117_U61 );
nand NAND3_13496 ( P1_R1117_U332 , P1_R1117_U331 , P1_R1117_U330 , P1_R1117_U10 );
nand NAND2_13497 ( P1_R1117_U333 , P1_U3074 , P1_R1117_U49 );
nand NAND2_13498 ( P1_R1117_U334 , P1_R1117_U180 , P1_R1117_U333 );
nand NAND2_13499 ( P1_R1117_U335 , P1_R1117_U262 , P1_R1117_U64 );
nand NAND2_13500 ( P1_R1117_U336 , P1_R1117_U217 , P1_R1117_U148 );
not NOT1_13501 ( P1_R1117_U337 , P1_R1117_U92 );
nand NAND2_13502 ( P1_R1117_U338 , P1_U3062 , P1_R1117_U51 );
nand NAND2_13503 ( P1_R1117_U339 , P1_R1117_U337 , P1_R1117_U338 );
nand NAND2_13504 ( P1_R1117_U340 , P1_R1117_U146 , P1_R1117_U339 );
nand NAND2_13505 ( P1_R1117_U341 , P1_R1117_U92 , P1_R1117_U179 );
nand NAND2_13506 ( P1_R1117_U342 , P1_U3491 , P1_R1117_U52 );
nand NAND2_13507 ( P1_R1117_U343 , P1_R1117_U145 , P1_R1117_U341 );
nand NAND2_13508 ( P1_R1117_U344 , P1_U3062 , P1_R1117_U51 );
nand NAND2_13509 ( P1_R1117_U345 , P1_R1117_U179 , P1_R1117_U344 );
nand NAND2_13510 ( P1_R1117_U346 , P1_U3077 , P1_R1117_U24 );
nand NAND3_13511 ( P1_R1117_U347 , P1_R1117_U89 , P1_R1117_U182 , P1_R1117_U301 );
nand NAND3_13512 ( P1_R1117_U348 , P1_R1117_U12 , P1_R1117_U347 , P1_R1117_U130 );
nand NAND2_13513 ( P1_R1117_U349 , P1_U3485 , P1_R1117_U43 );
nand NAND2_13514 ( P1_R1117_U350 , P1_U3083 , P1_R1117_U42 );
nand NAND2_13515 ( P1_R1117_U351 , P1_R1117_U218 , P1_R1117_U148 );
nand NAND2_13516 ( P1_R1117_U352 , P1_R1117_U216 , P1_R1117_U147 );
nand NAND2_13517 ( P1_R1117_U353 , P1_U3482 , P1_R1117_U41 );
nand NAND2_13518 ( P1_R1117_U354 , P1_U3084 , P1_R1117_U38 );
nand NAND2_13519 ( P1_R1117_U355 , P1_U3482 , P1_R1117_U41 );
nand NAND2_13520 ( P1_R1117_U356 , P1_U3084 , P1_R1117_U38 );
nand NAND2_13521 ( P1_R1117_U357 , P1_R1117_U356 , P1_R1117_U355 );
nand NAND2_13522 ( P1_R1117_U358 , P1_U3479 , P1_R1117_U39 );
nand NAND2_13523 ( P1_R1117_U359 , P1_U3070 , P1_R1117_U22 );
nand NAND2_13524 ( P1_R1117_U360 , P1_R1117_U223 , P1_R1117_U44 );
nand NAND2_13525 ( P1_R1117_U361 , P1_R1117_U149 , P1_R1117_U210 );
nand NAND2_13526 ( P1_R1117_U362 , P1_U3476 , P1_R1117_U34 );
nand NAND2_13527 ( P1_R1117_U363 , P1_U3071 , P1_R1117_U31 );
nand NAND2_13528 ( P1_R1117_U364 , P1_R1117_U363 , P1_R1117_U362 );
nand NAND2_13529 ( P1_R1117_U365 , P1_U3473 , P1_R1117_U35 );
nand NAND2_13530 ( P1_R1117_U366 , P1_U3067 , P1_R1117_U32 );
nand NAND2_13531 ( P1_R1117_U367 , P1_R1117_U233 , P1_R1117_U45 );
nand NAND2_13532 ( P1_R1117_U368 , P1_R1117_U150 , P1_R1117_U225 );
nand NAND2_13533 ( P1_R1117_U369 , P1_U3470 , P1_R1117_U36 );
nand NAND2_13534 ( P1_R1117_U370 , P1_U3060 , P1_R1117_U33 );
nand NAND2_13535 ( P1_R1117_U371 , P1_R1117_U234 , P1_R1117_U152 );
nand NAND2_13536 ( P1_R1117_U372 , P1_R1117_U200 , P1_R1117_U151 );
nand NAND2_13537 ( P1_R1117_U373 , P1_U3467 , P1_R1117_U30 );
nand NAND2_13538 ( P1_R1117_U374 , P1_U3064 , P1_R1117_U27 );
nand NAND2_13539 ( P1_R1117_U375 , P1_U3467 , P1_R1117_U30 );
nand NAND2_13540 ( P1_R1117_U376 , P1_U3064 , P1_R1117_U27 );
nand NAND2_13541 ( P1_R1117_U377 , P1_R1117_U376 , P1_R1117_U375 );
nand NAND2_13542 ( P1_R1117_U378 , P1_U3464 , P1_R1117_U28 );
nand NAND2_13543 ( P1_R1117_U379 , P1_U3068 , P1_R1117_U23 );
nand NAND2_13544 ( P1_R1117_U380 , P1_R1117_U239 , P1_R1117_U46 );
nand NAND2_13545 ( P1_R1117_U381 , P1_R1117_U153 , P1_R1117_U194 );
nand NAND2_13546 ( P1_R1117_U382 , P1_U4028 , P1_R1117_U155 );
nand NAND2_13547 ( P1_R1117_U383 , P1_U3055 , P1_R1117_U154 );
nand NAND2_13548 ( P1_R1117_U384 , P1_U4028 , P1_R1117_U155 );
nand NAND2_13549 ( P1_R1117_U385 , P1_U3055 , P1_R1117_U154 );
nand NAND2_13550 ( P1_R1117_U386 , P1_R1117_U385 , P1_R1117_U384 );
nand NAND3_13551 ( P1_R1117_U387 , P1_U3054 , P1_R1117_U386 , P1_R1117_U87 );
nand NAND3_13552 ( P1_R1117_U388 , P1_R1117_U12 , P1_R1117_U88 , P1_U4017 );
nand NAND2_13553 ( P1_R1117_U389 , P1_U4017 , P1_R1117_U88 );
nand NAND2_13554 ( P1_R1117_U390 , P1_U3054 , P1_R1117_U87 );
not NOT1_13555 ( P1_R1117_U391 , P1_R1117_U131 );
nand NAND2_13556 ( P1_R1117_U392 , P1_R1117_U306 , P1_R1117_U391 );
nand NAND2_13557 ( P1_R1117_U393 , P1_R1117_U131 , P1_R1117_U157 );
nand NAND2_13558 ( P1_R1117_U394 , P1_U4018 , P1_R1117_U86 );
nand NAND2_13559 ( P1_R1117_U395 , P1_U3053 , P1_R1117_U83 );
nand NAND2_13560 ( P1_R1117_U396 , P1_U4018 , P1_R1117_U86 );
nand NAND2_13561 ( P1_R1117_U397 , P1_U3053 , P1_R1117_U83 );
nand NAND2_13562 ( P1_R1117_U398 , P1_R1117_U397 , P1_R1117_U396 );
nand NAND2_13563 ( P1_R1117_U399 , P1_U4019 , P1_R1117_U84 );
nand NAND2_13564 ( P1_R1117_U400 , P1_U3057 , P1_R1117_U47 );
nand NAND2_13565 ( P1_R1117_U401 , P1_R1117_U313 , P1_R1117_U89 );
nand NAND2_13566 ( P1_R1117_U402 , P1_R1117_U158 , P1_R1117_U300 );
nand NAND2_13567 ( P1_R1117_U403 , P1_U4020 , P1_R1117_U82 );
nand NAND2_13568 ( P1_R1117_U404 , P1_U3058 , P1_R1117_U81 );
not NOT1_13569 ( P1_R1117_U405 , P1_R1117_U134 );
nand NAND2_13570 ( P1_R1117_U406 , P1_R1117_U296 , P1_R1117_U405 );
nand NAND2_13571 ( P1_R1117_U407 , P1_R1117_U134 , P1_R1117_U159 );
nand NAND2_13572 ( P1_R1117_U408 , P1_U4021 , P1_R1117_U80 );
nand NAND2_13573 ( P1_R1117_U409 , P1_U3065 , P1_R1117_U79 );
not NOT1_13574 ( P1_R1117_U410 , P1_R1117_U135 );
nand NAND2_13575 ( P1_R1117_U411 , P1_R1117_U292 , P1_R1117_U410 );
nand NAND2_13576 ( P1_R1117_U412 , P1_R1117_U135 , P1_R1117_U160 );
nand NAND2_13577 ( P1_R1117_U413 , P1_U4022 , P1_R1117_U75 );
nand NAND2_13578 ( P1_R1117_U414 , P1_U3066 , P1_R1117_U73 );
nand NAND2_13579 ( P1_R1117_U415 , P1_R1117_U414 , P1_R1117_U413 );
nand NAND2_13580 ( P1_R1117_U416 , P1_U4023 , P1_R1117_U76 );
nand NAND2_13581 ( P1_R1117_U417 , P1_U3061 , P1_R1117_U48 );
nand NAND2_13582 ( P1_R1117_U418 , P1_R1117_U323 , P1_R1117_U90 );
nand NAND2_13583 ( P1_R1117_U419 , P1_R1117_U161 , P1_R1117_U315 );
nand NAND2_13584 ( P1_R1117_U420 , P1_U4024 , P1_R1117_U77 );
nand NAND2_13585 ( P1_R1117_U421 , P1_U3075 , P1_R1117_U74 );
nand NAND2_13586 ( P1_R1117_U422 , P1_R1117_U324 , P1_R1117_U163 );
nand NAND2_13587 ( P1_R1117_U423 , P1_R1117_U282 , P1_R1117_U162 );
nand NAND2_13588 ( P1_R1117_U424 , P1_U4025 , P1_R1117_U72 );
nand NAND2_13589 ( P1_R1117_U425 , P1_U3076 , P1_R1117_U71 );
not NOT1_13590 ( P1_R1117_U426 , P1_R1117_U137 );
nand NAND2_13591 ( P1_R1117_U427 , P1_R1117_U278 , P1_R1117_U426 );
nand NAND2_13592 ( P1_R1117_U428 , P1_R1117_U137 , P1_R1117_U164 );
nand NAND2_13593 ( P1_R1117_U429 , P1_U3461 , P1_R1117_U26 );
nand NAND2_13594 ( P1_R1117_U430 , P1_U3078 , P1_R1117_U165 );
not NOT1_13595 ( P1_R1117_U431 , P1_R1117_U138 );
nand NAND2_13596 ( P1_R1117_U432 , P1_R1117_U431 , P1_R1117_U190 );
nand NAND2_13597 ( P1_R1117_U433 , P1_R1117_U138 , P1_R1117_U25 );
nand NAND2_13598 ( P1_R1117_U434 , P1_U3514 , P1_R1117_U70 );
nand NAND2_13599 ( P1_R1117_U435 , P1_U3081 , P1_R1117_U69 );
not NOT1_13600 ( P1_R1117_U436 , P1_R1117_U139 );
nand NAND2_13601 ( P1_R1117_U437 , P1_R1117_U274 , P1_R1117_U436 );
nand NAND2_13602 ( P1_R1117_U438 , P1_R1117_U139 , P1_R1117_U166 );
nand NAND2_13603 ( P1_R1117_U439 , P1_U3512 , P1_R1117_U68 );
nand NAND2_13604 ( P1_R1117_U440 , P1_U3082 , P1_R1117_U167 );
not NOT1_13605 ( P1_R1117_U441 , P1_R1117_U140 );
nand NAND2_13606 ( P1_R1117_U442 , P1_R1117_U441 , P1_R1117_U270 );
nand NAND2_13607 ( P1_R1117_U443 , P1_R1117_U140 , P1_R1117_U67 );
nand NAND2_13608 ( P1_R1117_U444 , P1_U3509 , P1_R1117_U66 );
nand NAND2_13609 ( P1_R1117_U445 , P1_U3069 , P1_R1117_U65 );
not NOT1_13610 ( P1_R1117_U446 , P1_R1117_U141 );
nand NAND2_13611 ( P1_R1117_U447 , P1_R1117_U266 , P1_R1117_U446 );
nand NAND2_13612 ( P1_R1117_U448 , P1_R1117_U141 , P1_R1117_U168 );
nand NAND2_13613 ( P1_R1117_U449 , P1_U3506 , P1_R1117_U61 );
nand NAND2_13614 ( P1_R1117_U450 , P1_U3073 , P1_R1117_U59 );
nand NAND2_13615 ( P1_R1117_U451 , P1_R1117_U450 , P1_R1117_U449 );
nand NAND2_13616 ( P1_R1117_U452 , P1_U3503 , P1_R1117_U62 );
nand NAND2_13617 ( P1_R1117_U453 , P1_U3074 , P1_R1117_U49 );
nand NAND2_13618 ( P1_R1117_U454 , P1_R1117_U334 , P1_R1117_U91 );
nand NAND2_13619 ( P1_R1117_U455 , P1_R1117_U169 , P1_R1117_U326 );
nand NAND2_13620 ( P1_R1117_U456 , P1_U3500 , P1_R1117_U63 );
nand NAND2_13621 ( P1_R1117_U457 , P1_U3079 , P1_R1117_U60 );
nand NAND2_13622 ( P1_R1117_U458 , P1_R1117_U335 , P1_R1117_U171 );
nand NAND2_13623 ( P1_R1117_U459 , P1_R1117_U256 , P1_R1117_U170 );
nand NAND2_13624 ( P1_R1117_U460 , P1_U3497 , P1_R1117_U58 );
nand NAND2_13625 ( P1_R1117_U461 , P1_U3080 , P1_R1117_U57 );
not NOT1_13626 ( P1_R1117_U462 , P1_R1117_U143 );
nand NAND2_13627 ( P1_R1117_U463 , P1_R1117_U252 , P1_R1117_U462 );
nand NAND2_13628 ( P1_R1117_U464 , P1_R1117_U143 , P1_R1117_U172 );
nand NAND2_13629 ( P1_R1117_U465 , P1_U3494 , P1_R1117_U56 );
nand NAND2_13630 ( P1_R1117_U466 , P1_U3072 , P1_R1117_U55 );
not NOT1_13631 ( P1_R1117_U467 , P1_R1117_U144 );
nand NAND2_13632 ( P1_R1117_U468 , P1_R1117_U248 , P1_R1117_U467 );
nand NAND2_13633 ( P1_R1117_U469 , P1_R1117_U144 , P1_R1117_U173 );
nand NAND2_13634 ( P1_R1117_U470 , P1_U3491 , P1_R1117_U52 );
nand NAND2_13635 ( P1_R1117_U471 , P1_U3063 , P1_R1117_U50 );
nand NAND2_13636 ( P1_R1117_U472 , P1_R1117_U471 , P1_R1117_U470 );
nand NAND2_13637 ( P1_R1117_U473 , P1_U3488 , P1_R1117_U53 );
nand NAND2_13638 ( P1_R1117_U474 , P1_U3062 , P1_R1117_U51 );
nand NAND2_13639 ( P1_R1117_U475 , P1_R1117_U345 , P1_R1117_U92 );
nand NAND2_13640 ( P1_R1117_U476 , P1_R1117_U174 , P1_R1117_U337 );
and AND2_13641 ( P1_R1375_U6 , P1_R1375_U8 , P1_R1375_U191 );
and AND3_13642 ( P1_R1375_U7 , P1_R1375_U190 , P1_R1375_U100 , P1_R1375_U189 );
and AND2_13643 ( P1_R1375_U8 , P1_R1375_U195 , P1_R1375_U194 );
nand NAND2_13644 ( P1_R1375_U9 , P1_R1375_U7 , P1_R1375_U192 );
not NOT1_13645 ( P1_R1375_U10 , P1_U3088 );
not NOT1_13646 ( P1_R1375_U11 , P1_U3087 );
not NOT1_13647 ( P1_R1375_U12 , P1_U3121 );
not NOT1_13648 ( P1_R1375_U13 , P1_U3120 );
not NOT1_13649 ( P1_R1375_U14 , P1_U3152 );
not NOT1_13650 ( P1_R1375_U15 , P1_U3117 );
not NOT1_13651 ( P1_R1375_U16 , P1_U3149 );
not NOT1_13652 ( P1_R1375_U17 , P1_U3148 );
not NOT1_13653 ( P1_R1375_U18 , P1_U3116 );
not NOT1_13654 ( P1_R1375_U19 , P1_U3115 );
not NOT1_13655 ( P1_R1375_U20 , P1_U3147 );
not NOT1_13656 ( P1_R1375_U21 , P1_U3146 );
not NOT1_13657 ( P1_R1375_U22 , P1_U3114 );
not NOT1_13658 ( P1_R1375_U23 , P1_U3113 );
not NOT1_13659 ( P1_R1375_U24 , P1_U3145 );
not NOT1_13660 ( P1_R1375_U25 , P1_U3144 );
not NOT1_13661 ( P1_R1375_U26 , P1_U3112 );
not NOT1_13662 ( P1_R1375_U27 , P1_U3111 );
not NOT1_13663 ( P1_R1375_U28 , P1_U3143 );
not NOT1_13664 ( P1_R1375_U29 , P1_U3142 );
not NOT1_13665 ( P1_R1375_U30 , P1_U3110 );
not NOT1_13666 ( P1_R1375_U31 , P1_U3109 );
not NOT1_13667 ( P1_R1375_U32 , P1_U3141 );
not NOT1_13668 ( P1_R1375_U33 , P1_U3140 );
not NOT1_13669 ( P1_R1375_U34 , P1_U3108 );
not NOT1_13670 ( P1_R1375_U35 , P1_U3107 );
not NOT1_13671 ( P1_R1375_U36 , P1_U3139 );
not NOT1_13672 ( P1_R1375_U37 , P1_U3138 );
not NOT1_13673 ( P1_R1375_U38 , P1_U3106 );
not NOT1_13674 ( P1_R1375_U39 , P1_U3105 );
not NOT1_13675 ( P1_R1375_U40 , P1_U3137 );
not NOT1_13676 ( P1_R1375_U41 , P1_U3136 );
not NOT1_13677 ( P1_R1375_U42 , P1_U3104 );
not NOT1_13678 ( P1_R1375_U43 , P1_U3103 );
not NOT1_13679 ( P1_R1375_U44 , P1_U3135 );
not NOT1_13680 ( P1_R1375_U45 , P1_U3134 );
not NOT1_13681 ( P1_R1375_U46 , P1_U3102 );
not NOT1_13682 ( P1_R1375_U47 , P1_U3101 );
not NOT1_13683 ( P1_R1375_U48 , P1_U3133 );
not NOT1_13684 ( P1_R1375_U49 , P1_U3132 );
not NOT1_13685 ( P1_R1375_U50 , P1_U3100 );
not NOT1_13686 ( P1_R1375_U51 , P1_U3099 );
not NOT1_13687 ( P1_R1375_U52 , P1_U3131 );
not NOT1_13688 ( P1_R1375_U53 , P1_U3130 );
not NOT1_13689 ( P1_R1375_U54 , P1_U3098 );
not NOT1_13690 ( P1_R1375_U55 , P1_U3097 );
not NOT1_13691 ( P1_R1375_U56 , P1_U3129 );
not NOT1_13692 ( P1_R1375_U57 , P1_U3128 );
not NOT1_13693 ( P1_R1375_U58 , P1_U3096 );
not NOT1_13694 ( P1_R1375_U59 , P1_U3095 );
not NOT1_13695 ( P1_R1375_U60 , P1_U3127 );
not NOT1_13696 ( P1_R1375_U61 , P1_U3126 );
not NOT1_13697 ( P1_R1375_U62 , P1_U3094 );
not NOT1_13698 ( P1_R1375_U63 , P1_U3093 );
not NOT1_13699 ( P1_R1375_U64 , P1_U3125 );
not NOT1_13700 ( P1_R1375_U65 , P1_U3124 );
not NOT1_13701 ( P1_R1375_U66 , P1_U3092 );
not NOT1_13702 ( P1_R1375_U67 , P1_U3091 );
not NOT1_13703 ( P1_R1375_U68 , P1_U3123 );
not NOT1_13704 ( P1_R1375_U69 , P1_U3089 );
and AND2_13705 ( P1_R1375_U70 , P1_R1375_U107 , P1_R1375_U108 );
and AND2_13706 ( P1_R1375_U71 , P1_R1375_U110 , P1_R1375_U111 );
and AND2_13707 ( P1_R1375_U72 , P1_R1375_U113 , P1_R1375_U114 );
and AND2_13708 ( P1_R1375_U73 , P1_R1375_U116 , P1_R1375_U117 );
and AND2_13709 ( P1_R1375_U74 , P1_R1375_U119 , P1_R1375_U120 );
and AND2_13710 ( P1_R1375_U75 , P1_R1375_U122 , P1_R1375_U123 );
and AND2_13711 ( P1_R1375_U76 , P1_R1375_U125 , P1_R1375_U126 );
and AND2_13712 ( P1_R1375_U77 , P1_R1375_U128 , P1_R1375_U129 );
and AND2_13713 ( P1_R1375_U78 , P1_R1375_U131 , P1_R1375_U132 );
and AND2_13714 ( P1_R1375_U79 , P1_R1375_U134 , P1_R1375_U135 );
and AND2_13715 ( P1_R1375_U80 , P1_R1375_U137 , P1_R1375_U138 );
and AND2_13716 ( P1_R1375_U81 , P1_R1375_U140 , P1_R1375_U141 );
and AND2_13717 ( P1_R1375_U82 , P1_R1375_U143 , P1_R1375_U144 );
and AND2_13718 ( P1_R1375_U83 , P1_R1375_U146 , P1_R1375_U147 );
and AND2_13719 ( P1_R1375_U84 , P1_R1375_U149 , P1_R1375_U150 );
and AND2_13720 ( P1_R1375_U85 , P1_R1375_U152 , P1_R1375_U153 );
and AND2_13721 ( P1_R1375_U86 , P1_R1375_U155 , P1_R1375_U156 );
and AND2_13722 ( P1_R1375_U87 , P1_R1375_U158 , P1_R1375_U159 );
and AND2_13723 ( P1_R1375_U88 , P1_R1375_U161 , P1_R1375_U162 );
and AND2_13724 ( P1_R1375_U89 , P1_R1375_U164 , P1_R1375_U165 );
and AND2_13725 ( P1_R1375_U90 , P1_R1375_U167 , P1_R1375_U168 );
and AND2_13726 ( P1_R1375_U91 , P1_R1375_U170 , P1_R1375_U171 );
and AND2_13727 ( P1_R1375_U92 , P1_R1375_U173 , P1_R1375_U174 );
and AND2_13728 ( P1_R1375_U93 , P1_R1375_U176 , P1_R1375_U177 );
and AND2_13729 ( P1_R1375_U94 , P1_R1375_U179 , P1_R1375_U180 );
and AND2_13730 ( P1_R1375_U95 , P1_R1375_U182 , P1_R1375_U183 );
and AND2_13731 ( P1_R1375_U96 , P1_R1375_U186 , P1_R1375_U101 );
and AND2_13732 ( P1_R1375_U97 , P1_R1375_U186 , P1_U3090 );
and AND2_13733 ( P1_R1375_U98 , P1_R1375_U187 , P1_R1375_U188 );
not NOT1_13734 ( P1_R1375_U99 , P1_U3119 );
and AND2_13735 ( P1_R1375_U100 , P1_R1375_U197 , P1_R1375_U196 );
not NOT1_13736 ( P1_R1375_U101 , P1_U3122 );
nand NAND2_13737 ( P1_R1375_U102 , P1_U3150 , P1_U3151 );
nand NAND2_13738 ( P1_R1375_U103 , P1_U3118 , P1_R1375_U102 );
or OR2_13739 ( P1_R1375_U104 , P1_U3150 , P1_U3151 );
nand NAND2_13740 ( P1_R1375_U105 , P1_U3117 , P1_R1375_U16 );
nand NAND3_13741 ( P1_R1375_U106 , P1_R1375_U104 , P1_R1375_U105 , P1_R1375_U103 );
nand NAND2_13742 ( P1_R1375_U107 , P1_U3149 , P1_R1375_U15 );
nand NAND2_13743 ( P1_R1375_U108 , P1_U3148 , P1_R1375_U18 );
nand NAND2_13744 ( P1_R1375_U109 , P1_R1375_U70 , P1_R1375_U106 );
nand NAND2_13745 ( P1_R1375_U110 , P1_U3116 , P1_R1375_U17 );
nand NAND2_13746 ( P1_R1375_U111 , P1_U3115 , P1_R1375_U20 );
nand NAND2_13747 ( P1_R1375_U112 , P1_R1375_U71 , P1_R1375_U109 );
nand NAND2_13748 ( P1_R1375_U113 , P1_U3147 , P1_R1375_U19 );
nand NAND2_13749 ( P1_R1375_U114 , P1_U3146 , P1_R1375_U22 );
nand NAND2_13750 ( P1_R1375_U115 , P1_R1375_U72 , P1_R1375_U112 );
nand NAND2_13751 ( P1_R1375_U116 , P1_U3114 , P1_R1375_U21 );
nand NAND2_13752 ( P1_R1375_U117 , P1_U3113 , P1_R1375_U24 );
nand NAND2_13753 ( P1_R1375_U118 , P1_R1375_U73 , P1_R1375_U115 );
nand NAND2_13754 ( P1_R1375_U119 , P1_U3145 , P1_R1375_U23 );
nand NAND2_13755 ( P1_R1375_U120 , P1_U3144 , P1_R1375_U26 );
nand NAND2_13756 ( P1_R1375_U121 , P1_R1375_U74 , P1_R1375_U118 );
nand NAND2_13757 ( P1_R1375_U122 , P1_U3112 , P1_R1375_U25 );
nand NAND2_13758 ( P1_R1375_U123 , P1_U3111 , P1_R1375_U28 );
nand NAND2_13759 ( P1_R1375_U124 , P1_R1375_U75 , P1_R1375_U121 );
nand NAND2_13760 ( P1_R1375_U125 , P1_U3143 , P1_R1375_U27 );
nand NAND2_13761 ( P1_R1375_U126 , P1_U3142 , P1_R1375_U30 );
nand NAND2_13762 ( P1_R1375_U127 , P1_R1375_U76 , P1_R1375_U124 );
nand NAND2_13763 ( P1_R1375_U128 , P1_U3110 , P1_R1375_U29 );
nand NAND2_13764 ( P1_R1375_U129 , P1_U3109 , P1_R1375_U32 );
nand NAND2_13765 ( P1_R1375_U130 , P1_R1375_U77 , P1_R1375_U127 );
nand NAND2_13766 ( P1_R1375_U131 , P1_U3141 , P1_R1375_U31 );
nand NAND2_13767 ( P1_R1375_U132 , P1_U3140 , P1_R1375_U34 );
nand NAND2_13768 ( P1_R1375_U133 , P1_R1375_U78 , P1_R1375_U130 );
nand NAND2_13769 ( P1_R1375_U134 , P1_U3108 , P1_R1375_U33 );
nand NAND2_13770 ( P1_R1375_U135 , P1_U3107 , P1_R1375_U36 );
nand NAND2_13771 ( P1_R1375_U136 , P1_R1375_U79 , P1_R1375_U133 );
nand NAND2_13772 ( P1_R1375_U137 , P1_U3139 , P1_R1375_U35 );
nand NAND2_13773 ( P1_R1375_U138 , P1_U3138 , P1_R1375_U38 );
nand NAND2_13774 ( P1_R1375_U139 , P1_R1375_U80 , P1_R1375_U136 );
nand NAND2_13775 ( P1_R1375_U140 , P1_U3106 , P1_R1375_U37 );
nand NAND2_13776 ( P1_R1375_U141 , P1_U3105 , P1_R1375_U40 );
nand NAND2_13777 ( P1_R1375_U142 , P1_R1375_U81 , P1_R1375_U139 );
nand NAND2_13778 ( P1_R1375_U143 , P1_U3137 , P1_R1375_U39 );
nand NAND2_13779 ( P1_R1375_U144 , P1_U3136 , P1_R1375_U42 );
nand NAND2_13780 ( P1_R1375_U145 , P1_R1375_U82 , P1_R1375_U142 );
nand NAND2_13781 ( P1_R1375_U146 , P1_U3104 , P1_R1375_U41 );
nand NAND2_13782 ( P1_R1375_U147 , P1_U3103 , P1_R1375_U44 );
nand NAND2_13783 ( P1_R1375_U148 , P1_R1375_U83 , P1_R1375_U145 );
nand NAND2_13784 ( P1_R1375_U149 , P1_U3135 , P1_R1375_U43 );
nand NAND2_13785 ( P1_R1375_U150 , P1_U3134 , P1_R1375_U46 );
nand NAND2_13786 ( P1_R1375_U151 , P1_R1375_U84 , P1_R1375_U148 );
nand NAND2_13787 ( P1_R1375_U152 , P1_U3102 , P1_R1375_U45 );
nand NAND2_13788 ( P1_R1375_U153 , P1_U3101 , P1_R1375_U48 );
nand NAND2_13789 ( P1_R1375_U154 , P1_R1375_U85 , P1_R1375_U151 );
nand NAND2_13790 ( P1_R1375_U155 , P1_U3133 , P1_R1375_U47 );
nand NAND2_13791 ( P1_R1375_U156 , P1_U3132 , P1_R1375_U50 );
nand NAND2_13792 ( P1_R1375_U157 , P1_R1375_U86 , P1_R1375_U154 );
nand NAND2_13793 ( P1_R1375_U158 , P1_U3100 , P1_R1375_U49 );
nand NAND2_13794 ( P1_R1375_U159 , P1_U3099 , P1_R1375_U52 );
nand NAND2_13795 ( P1_R1375_U160 , P1_R1375_U87 , P1_R1375_U157 );
nand NAND2_13796 ( P1_R1375_U161 , P1_U3131 , P1_R1375_U51 );
nand NAND2_13797 ( P1_R1375_U162 , P1_U3130 , P1_R1375_U54 );
nand NAND2_13798 ( P1_R1375_U163 , P1_R1375_U88 , P1_R1375_U160 );
nand NAND2_13799 ( P1_R1375_U164 , P1_U3098 , P1_R1375_U53 );
nand NAND2_13800 ( P1_R1375_U165 , P1_U3097 , P1_R1375_U56 );
nand NAND2_13801 ( P1_R1375_U166 , P1_R1375_U89 , P1_R1375_U163 );
nand NAND2_13802 ( P1_R1375_U167 , P1_U3129 , P1_R1375_U55 );
nand NAND2_13803 ( P1_R1375_U168 , P1_U3128 , P1_R1375_U58 );
nand NAND2_13804 ( P1_R1375_U169 , P1_R1375_U90 , P1_R1375_U166 );
nand NAND2_13805 ( P1_R1375_U170 , P1_U3096 , P1_R1375_U57 );
nand NAND2_13806 ( P1_R1375_U171 , P1_U3095 , P1_R1375_U60 );
nand NAND2_13807 ( P1_R1375_U172 , P1_R1375_U91 , P1_R1375_U169 );
nand NAND2_13808 ( P1_R1375_U173 , P1_U3127 , P1_R1375_U59 );
nand NAND2_13809 ( P1_R1375_U174 , P1_U3126 , P1_R1375_U62 );
nand NAND2_13810 ( P1_R1375_U175 , P1_R1375_U92 , P1_R1375_U172 );
nand NAND2_13811 ( P1_R1375_U176 , P1_U3094 , P1_R1375_U61 );
nand NAND2_13812 ( P1_R1375_U177 , P1_U3093 , P1_R1375_U64 );
nand NAND2_13813 ( P1_R1375_U178 , P1_R1375_U93 , P1_R1375_U175 );
nand NAND2_13814 ( P1_R1375_U179 , P1_U3125 , P1_R1375_U63 );
nand NAND2_13815 ( P1_R1375_U180 , P1_U3124 , P1_R1375_U66 );
nand NAND2_13816 ( P1_R1375_U181 , P1_R1375_U94 , P1_R1375_U178 );
nand NAND2_13817 ( P1_R1375_U182 , P1_U3092 , P1_R1375_U65 );
nand NAND2_13818 ( P1_R1375_U183 , P1_U3091 , P1_R1375_U68 );
nand NAND2_13819 ( P1_R1375_U184 , P1_R1375_U95 , P1_R1375_U181 );
nand NAND2_13820 ( P1_R1375_U185 , P1_R1375_U96 , P1_R1375_U184 );
nand NAND2_13821 ( P1_R1375_U186 , P1_U3123 , P1_R1375_U67 );
nand NAND2_13822 ( P1_R1375_U187 , P1_U3090 , P1_R1375_U101 );
nand NAND2_13823 ( P1_R1375_U188 , P1_U3089 , P1_R1375_U12 );
nand NAND4_13824 ( P1_R1375_U189 , P1_R1375_U8 , P1_R1375_U191 , P1_U3121 , P1_R1375_U69 );
nand NAND3_13825 ( P1_R1375_U190 , P1_R1375_U8 , P1_R1375_U10 , P1_U3120 );
nand NAND2_13826 ( P1_R1375_U191 , P1_U3088 , P1_R1375_U13 );
nand NAND4_13827 ( P1_R1375_U192 , P1_R1375_U6 , P1_R1375_U193 , P1_R1375_U98 , P1_R1375_U185 );
nand NAND2_13828 ( P1_R1375_U193 , P1_R1375_U97 , P1_R1375_U184 );
nand NAND2_13829 ( P1_R1375_U194 , P1_U3087 , P1_R1375_U99 );
nand NAND2_13830 ( P1_R1375_U195 , P1_U3119 , P1_R1375_U11 );
nand NAND3_13831 ( P1_R1375_U196 , P1_U3152 , P1_U3087 , P1_R1375_U99 );
nand NAND3_13832 ( P1_R1375_U197 , P1_R1375_U14 , P1_R1375_U11 , P1_U3119 );
and AND2_13833 ( P1_R1352_U6 , P1_U3059 , P1_R1352_U7 );
not NOT1_13834 ( P1_R1352_U7 , P1_U3056 );
and AND2_13835 ( P1_R1207_U6 , P1_R1207_U184 , P1_R1207_U201 );
and AND2_13836 ( P1_R1207_U7 , P1_R1207_U203 , P1_R1207_U202 );
and AND2_13837 ( P1_R1207_U8 , P1_R1207_U179 , P1_R1207_U240 );
and AND2_13838 ( P1_R1207_U9 , P1_R1207_U242 , P1_R1207_U241 );
and AND2_13839 ( P1_R1207_U10 , P1_R1207_U259 , P1_R1207_U258 );
and AND2_13840 ( P1_R1207_U11 , P1_R1207_U285 , P1_R1207_U284 );
and AND2_13841 ( P1_R1207_U12 , P1_R1207_U383 , P1_R1207_U382 );
nand NAND2_13842 ( P1_R1207_U13 , P1_R1207_U340 , P1_R1207_U343 );
nand NAND2_13843 ( P1_R1207_U14 , P1_R1207_U329 , P1_R1207_U332 );
nand NAND2_13844 ( P1_R1207_U15 , P1_R1207_U318 , P1_R1207_U321 );
nand NAND2_13845 ( P1_R1207_U16 , P1_R1207_U310 , P1_R1207_U312 );
nand NAND3_13846 ( P1_R1207_U17 , P1_R1207_U156 , P1_R1207_U175 , P1_R1207_U348 );
nand NAND2_13847 ( P1_R1207_U18 , P1_R1207_U236 , P1_R1207_U238 );
nand NAND2_13848 ( P1_R1207_U19 , P1_R1207_U228 , P1_R1207_U231 );
nand NAND2_13849 ( P1_R1207_U20 , P1_R1207_U220 , P1_R1207_U222 );
nand NAND2_13850 ( P1_R1207_U21 , P1_R1207_U25 , P1_R1207_U346 );
not NOT1_13851 ( P1_R1207_U22 , P1_U3479 );
not NOT1_13852 ( P1_R1207_U23 , P1_U3464 );
not NOT1_13853 ( P1_R1207_U24 , P1_U3456 );
nand NAND2_13854 ( P1_R1207_U25 , P1_U3456 , P1_R1207_U93 );
not NOT1_13855 ( P1_R1207_U26 , P1_U3078 );
not NOT1_13856 ( P1_R1207_U27 , P1_U3467 );
not NOT1_13857 ( P1_R1207_U28 , P1_U3068 );
nand NAND2_13858 ( P1_R1207_U29 , P1_U3068 , P1_R1207_U23 );
not NOT1_13859 ( P1_R1207_U30 , P1_U3064 );
not NOT1_13860 ( P1_R1207_U31 , P1_U3476 );
not NOT1_13861 ( P1_R1207_U32 , P1_U3473 );
not NOT1_13862 ( P1_R1207_U33 , P1_U3470 );
not NOT1_13863 ( P1_R1207_U34 , P1_U3071 );
not NOT1_13864 ( P1_R1207_U35 , P1_U3067 );
not NOT1_13865 ( P1_R1207_U36 , P1_U3060 );
nand NAND2_13866 ( P1_R1207_U37 , P1_U3060 , P1_R1207_U33 );
not NOT1_13867 ( P1_R1207_U38 , P1_U3482 );
not NOT1_13868 ( P1_R1207_U39 , P1_U3070 );
nand NAND2_13869 ( P1_R1207_U40 , P1_U3070 , P1_R1207_U22 );
not NOT1_13870 ( P1_R1207_U41 , P1_U3084 );
not NOT1_13871 ( P1_R1207_U42 , P1_U3485 );
not NOT1_13872 ( P1_R1207_U43 , P1_U3083 );
nand NAND2_13873 ( P1_R1207_U44 , P1_R1207_U209 , P1_R1207_U208 );
nand NAND2_13874 ( P1_R1207_U45 , P1_R1207_U37 , P1_R1207_U224 );
nand NAND2_13875 ( P1_R1207_U46 , P1_R1207_U193 , P1_R1207_U192 );
not NOT1_13876 ( P1_R1207_U47 , P1_U4019 );
not NOT1_13877 ( P1_R1207_U48 , P1_U4023 );
not NOT1_13878 ( P1_R1207_U49 , P1_U3503 );
not NOT1_13879 ( P1_R1207_U50 , P1_U3491 );
not NOT1_13880 ( P1_R1207_U51 , P1_U3488 );
not NOT1_13881 ( P1_R1207_U52 , P1_U3063 );
not NOT1_13882 ( P1_R1207_U53 , P1_U3062 );
nand NAND2_13883 ( P1_R1207_U54 , P1_U3083 , P1_R1207_U42 );
not NOT1_13884 ( P1_R1207_U55 , P1_U3494 );
not NOT1_13885 ( P1_R1207_U56 , P1_U3072 );
not NOT1_13886 ( P1_R1207_U57 , P1_U3497 );
not NOT1_13887 ( P1_R1207_U58 , P1_U3080 );
not NOT1_13888 ( P1_R1207_U59 , P1_U3506 );
not NOT1_13889 ( P1_R1207_U60 , P1_U3500 );
not NOT1_13890 ( P1_R1207_U61 , P1_U3073 );
not NOT1_13891 ( P1_R1207_U62 , P1_U3074 );
not NOT1_13892 ( P1_R1207_U63 , P1_U3079 );
nand NAND2_13893 ( P1_R1207_U64 , P1_U3079 , P1_R1207_U60 );
not NOT1_13894 ( P1_R1207_U65 , P1_U3509 );
not NOT1_13895 ( P1_R1207_U66 , P1_U3069 );
nand NAND2_13896 ( P1_R1207_U67 , P1_R1207_U269 , P1_R1207_U268 );
not NOT1_13897 ( P1_R1207_U68 , P1_U3082 );
not NOT1_13898 ( P1_R1207_U69 , P1_U3514 );
not NOT1_13899 ( P1_R1207_U70 , P1_U3081 );
not NOT1_13900 ( P1_R1207_U71 , P1_U4025 );
not NOT1_13901 ( P1_R1207_U72 , P1_U3076 );
not NOT1_13902 ( P1_R1207_U73 , P1_U4022 );
not NOT1_13903 ( P1_R1207_U74 , P1_U4024 );
not NOT1_13904 ( P1_R1207_U75 , P1_U3066 );
not NOT1_13905 ( P1_R1207_U76 , P1_U3061 );
not NOT1_13906 ( P1_R1207_U77 , P1_U3075 );
nand NAND2_13907 ( P1_R1207_U78 , P1_U3075 , P1_R1207_U74 );
not NOT1_13908 ( P1_R1207_U79 , P1_U4021 );
not NOT1_13909 ( P1_R1207_U80 , P1_U3065 );
not NOT1_13910 ( P1_R1207_U81 , P1_U4020 );
not NOT1_13911 ( P1_R1207_U82 , P1_U3058 );
not NOT1_13912 ( P1_R1207_U83 , P1_U4018 );
not NOT1_13913 ( P1_R1207_U84 , P1_U3057 );
nand NAND2_13914 ( P1_R1207_U85 , P1_U3057 , P1_R1207_U47 );
not NOT1_13915 ( P1_R1207_U86 , P1_U3053 );
not NOT1_13916 ( P1_R1207_U87 , P1_U4017 );
not NOT1_13917 ( P1_R1207_U88 , P1_U3054 );
nand NAND2_13918 ( P1_R1207_U89 , P1_R1207_U299 , P1_R1207_U298 );
nand NAND2_13919 ( P1_R1207_U90 , P1_R1207_U78 , P1_R1207_U314 );
nand NAND2_13920 ( P1_R1207_U91 , P1_R1207_U64 , P1_R1207_U325 );
nand NAND2_13921 ( P1_R1207_U92 , P1_R1207_U54 , P1_R1207_U336 );
not NOT1_13922 ( P1_R1207_U93 , P1_U3077 );
nand NAND2_13923 ( P1_R1207_U94 , P1_R1207_U393 , P1_R1207_U392 );
nand NAND2_13924 ( P1_R1207_U95 , P1_R1207_U407 , P1_R1207_U406 );
nand NAND2_13925 ( P1_R1207_U96 , P1_R1207_U412 , P1_R1207_U411 );
nand NAND2_13926 ( P1_R1207_U97 , P1_R1207_U428 , P1_R1207_U427 );
nand NAND2_13927 ( P1_R1207_U98 , P1_R1207_U433 , P1_R1207_U432 );
nand NAND2_13928 ( P1_R1207_U99 , P1_R1207_U438 , P1_R1207_U437 );
nand NAND2_13929 ( P1_R1207_U100 , P1_R1207_U443 , P1_R1207_U442 );
nand NAND2_13930 ( P1_R1207_U101 , P1_R1207_U448 , P1_R1207_U447 );
nand NAND2_13931 ( P1_R1207_U102 , P1_R1207_U464 , P1_R1207_U463 );
nand NAND2_13932 ( P1_R1207_U103 , P1_R1207_U469 , P1_R1207_U468 );
nand NAND2_13933 ( P1_R1207_U104 , P1_R1207_U352 , P1_R1207_U351 );
nand NAND2_13934 ( P1_R1207_U105 , P1_R1207_U361 , P1_R1207_U360 );
nand NAND2_13935 ( P1_R1207_U106 , P1_R1207_U368 , P1_R1207_U367 );
nand NAND2_13936 ( P1_R1207_U107 , P1_R1207_U372 , P1_R1207_U371 );
nand NAND2_13937 ( P1_R1207_U108 , P1_R1207_U381 , P1_R1207_U380 );
nand NAND2_13938 ( P1_R1207_U109 , P1_R1207_U402 , P1_R1207_U401 );
nand NAND2_13939 ( P1_R1207_U110 , P1_R1207_U419 , P1_R1207_U418 );
nand NAND2_13940 ( P1_R1207_U111 , P1_R1207_U423 , P1_R1207_U422 );
nand NAND2_13941 ( P1_R1207_U112 , P1_R1207_U455 , P1_R1207_U454 );
nand NAND2_13942 ( P1_R1207_U113 , P1_R1207_U459 , P1_R1207_U458 );
nand NAND2_13943 ( P1_R1207_U114 , P1_R1207_U476 , P1_R1207_U475 );
and AND2_13944 ( P1_R1207_U115 , P1_R1207_U195 , P1_R1207_U183 );
and AND2_13945 ( P1_R1207_U116 , P1_R1207_U198 , P1_R1207_U199 );
and AND2_13946 ( P1_R1207_U117 , P1_R1207_U211 , P1_R1207_U185 );
and AND2_13947 ( P1_R1207_U118 , P1_R1207_U214 , P1_R1207_U215 );
and AND3_13948 ( P1_R1207_U119 , P1_R1207_U354 , P1_R1207_U353 , P1_R1207_U40 );
and AND2_13949 ( P1_R1207_U120 , P1_R1207_U357 , P1_R1207_U185 );
and AND2_13950 ( P1_R1207_U121 , P1_R1207_U230 , P1_R1207_U7 );
and AND2_13951 ( P1_R1207_U122 , P1_R1207_U364 , P1_R1207_U184 );
and AND3_13952 ( P1_R1207_U123 , P1_R1207_U374 , P1_R1207_U373 , P1_R1207_U29 );
and AND2_13953 ( P1_R1207_U124 , P1_R1207_U377 , P1_R1207_U183 );
and AND2_13954 ( P1_R1207_U125 , P1_R1207_U217 , P1_R1207_U8 );
and AND2_13955 ( P1_R1207_U126 , P1_R1207_U262 , P1_R1207_U180 );
and AND2_13956 ( P1_R1207_U127 , P1_R1207_U288 , P1_R1207_U181 );
and AND2_13957 ( P1_R1207_U128 , P1_R1207_U304 , P1_R1207_U305 );
and AND2_13958 ( P1_R1207_U129 , P1_R1207_U307 , P1_R1207_U386 );
and AND3_13959 ( P1_R1207_U130 , P1_R1207_U305 , P1_R1207_U304 , P1_R1207_U308 );
nand NAND2_13960 ( P1_R1207_U131 , P1_R1207_U390 , P1_R1207_U389 );
and AND3_13961 ( P1_R1207_U132 , P1_R1207_U395 , P1_R1207_U394 , P1_R1207_U85 );
and AND2_13962 ( P1_R1207_U133 , P1_R1207_U398 , P1_R1207_U182 );
nand NAND2_13963 ( P1_R1207_U134 , P1_R1207_U404 , P1_R1207_U403 );
nand NAND2_13964 ( P1_R1207_U135 , P1_R1207_U409 , P1_R1207_U408 );
and AND2_13965 ( P1_R1207_U136 , P1_R1207_U415 , P1_R1207_U181 );
nand NAND2_13966 ( P1_R1207_U137 , P1_R1207_U425 , P1_R1207_U424 );
nand NAND2_13967 ( P1_R1207_U138 , P1_R1207_U430 , P1_R1207_U429 );
nand NAND2_13968 ( P1_R1207_U139 , P1_R1207_U435 , P1_R1207_U434 );
nand NAND2_13969 ( P1_R1207_U140 , P1_R1207_U440 , P1_R1207_U439 );
nand NAND2_13970 ( P1_R1207_U141 , P1_R1207_U445 , P1_R1207_U444 );
and AND2_13971 ( P1_R1207_U142 , P1_R1207_U451 , P1_R1207_U180 );
nand NAND2_13972 ( P1_R1207_U143 , P1_R1207_U461 , P1_R1207_U460 );
nand NAND2_13973 ( P1_R1207_U144 , P1_R1207_U466 , P1_R1207_U465 );
and AND2_13974 ( P1_R1207_U145 , P1_R1207_U342 , P1_R1207_U9 );
and AND2_13975 ( P1_R1207_U146 , P1_R1207_U472 , P1_R1207_U179 );
and AND2_13976 ( P1_R1207_U147 , P1_R1207_U350 , P1_R1207_U349 );
nand NAND2_13977 ( P1_R1207_U148 , P1_R1207_U118 , P1_R1207_U212 );
and AND2_13978 ( P1_R1207_U149 , P1_R1207_U359 , P1_R1207_U358 );
and AND2_13979 ( P1_R1207_U150 , P1_R1207_U366 , P1_R1207_U365 );
and AND2_13980 ( P1_R1207_U151 , P1_R1207_U370 , P1_R1207_U369 );
nand NAND2_13981 ( P1_R1207_U152 , P1_R1207_U116 , P1_R1207_U196 );
and AND2_13982 ( P1_R1207_U153 , P1_R1207_U379 , P1_R1207_U378 );
not NOT1_13983 ( P1_R1207_U154 , P1_U4028 );
not NOT1_13984 ( P1_R1207_U155 , P1_U3055 );
and AND2_13985 ( P1_R1207_U156 , P1_R1207_U388 , P1_R1207_U387 );
nand NAND2_13986 ( P1_R1207_U157 , P1_R1207_U128 , P1_R1207_U302 );
and AND2_13987 ( P1_R1207_U158 , P1_R1207_U400 , P1_R1207_U399 );
nand NAND2_13988 ( P1_R1207_U159 , P1_R1207_U295 , P1_R1207_U294 );
nand NAND2_13989 ( P1_R1207_U160 , P1_R1207_U291 , P1_R1207_U290 );
and AND2_13990 ( P1_R1207_U161 , P1_R1207_U417 , P1_R1207_U416 );
and AND2_13991 ( P1_R1207_U162 , P1_R1207_U421 , P1_R1207_U420 );
nand NAND2_13992 ( P1_R1207_U163 , P1_R1207_U281 , P1_R1207_U280 );
nand NAND2_13993 ( P1_R1207_U164 , P1_R1207_U277 , P1_R1207_U276 );
not NOT1_13994 ( P1_R1207_U165 , P1_U3461 );
nand NAND2_13995 ( P1_R1207_U166 , P1_R1207_U273 , P1_R1207_U272 );
not NOT1_13996 ( P1_R1207_U167 , P1_U3512 );
nand NAND2_13997 ( P1_R1207_U168 , P1_R1207_U265 , P1_R1207_U264 );
and AND2_13998 ( P1_R1207_U169 , P1_R1207_U453 , P1_R1207_U452 );
and AND2_13999 ( P1_R1207_U170 , P1_R1207_U457 , P1_R1207_U456 );
nand NAND2_14000 ( P1_R1207_U171 , P1_R1207_U255 , P1_R1207_U254 );
nand NAND2_14001 ( P1_R1207_U172 , P1_R1207_U251 , P1_R1207_U250 );
nand NAND2_14002 ( P1_R1207_U173 , P1_R1207_U247 , P1_R1207_U246 );
and AND2_14003 ( P1_R1207_U174 , P1_R1207_U474 , P1_R1207_U473 );
nand NAND2_14004 ( P1_R1207_U175 , P1_R1207_U129 , P1_R1207_U157 );
not NOT1_14005 ( P1_R1207_U176 , P1_R1207_U85 );
not NOT1_14006 ( P1_R1207_U177 , P1_R1207_U29 );
not NOT1_14007 ( P1_R1207_U178 , P1_R1207_U40 );
nand NAND2_14008 ( P1_R1207_U179 , P1_U3488 , P1_R1207_U53 );
nand NAND2_14009 ( P1_R1207_U180 , P1_U3503 , P1_R1207_U62 );
nand NAND2_14010 ( P1_R1207_U181 , P1_U4023 , P1_R1207_U76 );
nand NAND2_14011 ( P1_R1207_U182 , P1_U4019 , P1_R1207_U84 );
nand NAND2_14012 ( P1_R1207_U183 , P1_U3464 , P1_R1207_U28 );
nand NAND2_14013 ( P1_R1207_U184 , P1_U3473 , P1_R1207_U35 );
nand NAND2_14014 ( P1_R1207_U185 , P1_U3479 , P1_R1207_U39 );
not NOT1_14015 ( P1_R1207_U186 , P1_R1207_U64 );
not NOT1_14016 ( P1_R1207_U187 , P1_R1207_U78 );
not NOT1_14017 ( P1_R1207_U188 , P1_R1207_U37 );
not NOT1_14018 ( P1_R1207_U189 , P1_R1207_U54 );
not NOT1_14019 ( P1_R1207_U190 , P1_R1207_U25 );
nand NAND2_14020 ( P1_R1207_U191 , P1_R1207_U190 , P1_R1207_U26 );
nand NAND2_14021 ( P1_R1207_U192 , P1_R1207_U191 , P1_R1207_U165 );
nand NAND2_14022 ( P1_R1207_U193 , P1_U3078 , P1_R1207_U25 );
not NOT1_14023 ( P1_R1207_U194 , P1_R1207_U46 );
nand NAND2_14024 ( P1_R1207_U195 , P1_U3467 , P1_R1207_U30 );
nand NAND2_14025 ( P1_R1207_U196 , P1_R1207_U115 , P1_R1207_U46 );
nand NAND2_14026 ( P1_R1207_U197 , P1_R1207_U30 , P1_R1207_U29 );
nand NAND2_14027 ( P1_R1207_U198 , P1_R1207_U197 , P1_R1207_U27 );
nand NAND2_14028 ( P1_R1207_U199 , P1_U3064 , P1_R1207_U177 );
not NOT1_14029 ( P1_R1207_U200 , P1_R1207_U152 );
nand NAND2_14030 ( P1_R1207_U201 , P1_U3476 , P1_R1207_U34 );
nand NAND2_14031 ( P1_R1207_U202 , P1_U3071 , P1_R1207_U31 );
nand NAND2_14032 ( P1_R1207_U203 , P1_U3067 , P1_R1207_U32 );
nand NAND2_14033 ( P1_R1207_U204 , P1_R1207_U188 , P1_R1207_U6 );
nand NAND2_14034 ( P1_R1207_U205 , P1_R1207_U7 , P1_R1207_U204 );
nand NAND2_14035 ( P1_R1207_U206 , P1_U3470 , P1_R1207_U36 );
nand NAND2_14036 ( P1_R1207_U207 , P1_U3476 , P1_R1207_U34 );
nand NAND3_14037 ( P1_R1207_U208 , P1_R1207_U206 , P1_R1207_U152 , P1_R1207_U6 );
nand NAND2_14038 ( P1_R1207_U209 , P1_R1207_U207 , P1_R1207_U205 );
not NOT1_14039 ( P1_R1207_U210 , P1_R1207_U44 );
nand NAND2_14040 ( P1_R1207_U211 , P1_U3482 , P1_R1207_U41 );
nand NAND2_14041 ( P1_R1207_U212 , P1_R1207_U117 , P1_R1207_U44 );
nand NAND2_14042 ( P1_R1207_U213 , P1_R1207_U41 , P1_R1207_U40 );
nand NAND2_14043 ( P1_R1207_U214 , P1_R1207_U213 , P1_R1207_U38 );
nand NAND2_14044 ( P1_R1207_U215 , P1_U3084 , P1_R1207_U178 );
not NOT1_14045 ( P1_R1207_U216 , P1_R1207_U148 );
nand NAND2_14046 ( P1_R1207_U217 , P1_U3485 , P1_R1207_U43 );
nand NAND2_14047 ( P1_R1207_U218 , P1_R1207_U217 , P1_R1207_U54 );
nand NAND2_14048 ( P1_R1207_U219 , P1_R1207_U210 , P1_R1207_U40 );
nand NAND2_14049 ( P1_R1207_U220 , P1_R1207_U120 , P1_R1207_U219 );
nand NAND2_14050 ( P1_R1207_U221 , P1_R1207_U44 , P1_R1207_U185 );
nand NAND2_14051 ( P1_R1207_U222 , P1_R1207_U119 , P1_R1207_U221 );
nand NAND2_14052 ( P1_R1207_U223 , P1_R1207_U40 , P1_R1207_U185 );
nand NAND2_14053 ( P1_R1207_U224 , P1_R1207_U206 , P1_R1207_U152 );
not NOT1_14054 ( P1_R1207_U225 , P1_R1207_U45 );
nand NAND2_14055 ( P1_R1207_U226 , P1_U3067 , P1_R1207_U32 );
nand NAND2_14056 ( P1_R1207_U227 , P1_R1207_U225 , P1_R1207_U226 );
nand NAND2_14057 ( P1_R1207_U228 , P1_R1207_U122 , P1_R1207_U227 );
nand NAND2_14058 ( P1_R1207_U229 , P1_R1207_U45 , P1_R1207_U184 );
nand NAND2_14059 ( P1_R1207_U230 , P1_U3476 , P1_R1207_U34 );
nand NAND2_14060 ( P1_R1207_U231 , P1_R1207_U121 , P1_R1207_U229 );
nand NAND2_14061 ( P1_R1207_U232 , P1_U3067 , P1_R1207_U32 );
nand NAND2_14062 ( P1_R1207_U233 , P1_R1207_U184 , P1_R1207_U232 );
nand NAND2_14063 ( P1_R1207_U234 , P1_R1207_U206 , P1_R1207_U37 );
nand NAND2_14064 ( P1_R1207_U235 , P1_R1207_U194 , P1_R1207_U29 );
nand NAND2_14065 ( P1_R1207_U236 , P1_R1207_U124 , P1_R1207_U235 );
nand NAND2_14066 ( P1_R1207_U237 , P1_R1207_U46 , P1_R1207_U183 );
nand NAND2_14067 ( P1_R1207_U238 , P1_R1207_U123 , P1_R1207_U237 );
nand NAND2_14068 ( P1_R1207_U239 , P1_R1207_U29 , P1_R1207_U183 );
nand NAND2_14069 ( P1_R1207_U240 , P1_U3491 , P1_R1207_U52 );
nand NAND2_14070 ( P1_R1207_U241 , P1_U3063 , P1_R1207_U50 );
nand NAND2_14071 ( P1_R1207_U242 , P1_U3062 , P1_R1207_U51 );
nand NAND2_14072 ( P1_R1207_U243 , P1_R1207_U189 , P1_R1207_U8 );
nand NAND2_14073 ( P1_R1207_U244 , P1_R1207_U9 , P1_R1207_U243 );
nand NAND2_14074 ( P1_R1207_U245 , P1_U3491 , P1_R1207_U52 );
nand NAND2_14075 ( P1_R1207_U246 , P1_R1207_U125 , P1_R1207_U148 );
nand NAND2_14076 ( P1_R1207_U247 , P1_R1207_U245 , P1_R1207_U244 );
not NOT1_14077 ( P1_R1207_U248 , P1_R1207_U173 );
nand NAND2_14078 ( P1_R1207_U249 , P1_U3494 , P1_R1207_U56 );
nand NAND2_14079 ( P1_R1207_U250 , P1_R1207_U249 , P1_R1207_U173 );
nand NAND2_14080 ( P1_R1207_U251 , P1_U3072 , P1_R1207_U55 );
not NOT1_14081 ( P1_R1207_U252 , P1_R1207_U172 );
nand NAND2_14082 ( P1_R1207_U253 , P1_U3497 , P1_R1207_U58 );
nand NAND2_14083 ( P1_R1207_U254 , P1_R1207_U253 , P1_R1207_U172 );
nand NAND2_14084 ( P1_R1207_U255 , P1_U3080 , P1_R1207_U57 );
not NOT1_14085 ( P1_R1207_U256 , P1_R1207_U171 );
nand NAND2_14086 ( P1_R1207_U257 , P1_U3506 , P1_R1207_U61 );
nand NAND2_14087 ( P1_R1207_U258 , P1_U3073 , P1_R1207_U59 );
nand NAND2_14088 ( P1_R1207_U259 , P1_U3074 , P1_R1207_U49 );
nand NAND2_14089 ( P1_R1207_U260 , P1_R1207_U186 , P1_R1207_U180 );
nand NAND2_14090 ( P1_R1207_U261 , P1_R1207_U10 , P1_R1207_U260 );
nand NAND2_14091 ( P1_R1207_U262 , P1_U3500 , P1_R1207_U63 );
nand NAND2_14092 ( P1_R1207_U263 , P1_U3506 , P1_R1207_U61 );
nand NAND3_14093 ( P1_R1207_U264 , P1_R1207_U171 , P1_R1207_U126 , P1_R1207_U257 );
nand NAND2_14094 ( P1_R1207_U265 , P1_R1207_U263 , P1_R1207_U261 );
not NOT1_14095 ( P1_R1207_U266 , P1_R1207_U168 );
nand NAND2_14096 ( P1_R1207_U267 , P1_U3509 , P1_R1207_U66 );
nand NAND2_14097 ( P1_R1207_U268 , P1_R1207_U267 , P1_R1207_U168 );
nand NAND2_14098 ( P1_R1207_U269 , P1_U3069 , P1_R1207_U65 );
not NOT1_14099 ( P1_R1207_U270 , P1_R1207_U67 );
nand NAND2_14100 ( P1_R1207_U271 , P1_R1207_U270 , P1_R1207_U68 );
nand NAND2_14101 ( P1_R1207_U272 , P1_R1207_U271 , P1_R1207_U167 );
nand NAND2_14102 ( P1_R1207_U273 , P1_U3082 , P1_R1207_U67 );
not NOT1_14103 ( P1_R1207_U274 , P1_R1207_U166 );
nand NAND2_14104 ( P1_R1207_U275 , P1_U3514 , P1_R1207_U70 );
nand NAND2_14105 ( P1_R1207_U276 , P1_R1207_U275 , P1_R1207_U166 );
nand NAND2_14106 ( P1_R1207_U277 , P1_U3081 , P1_R1207_U69 );
not NOT1_14107 ( P1_R1207_U278 , P1_R1207_U164 );
nand NAND2_14108 ( P1_R1207_U279 , P1_U4025 , P1_R1207_U72 );
nand NAND2_14109 ( P1_R1207_U280 , P1_R1207_U279 , P1_R1207_U164 );
nand NAND2_14110 ( P1_R1207_U281 , P1_U3076 , P1_R1207_U71 );
not NOT1_14111 ( P1_R1207_U282 , P1_R1207_U163 );
nand NAND2_14112 ( P1_R1207_U283 , P1_U4022 , P1_R1207_U75 );
nand NAND2_14113 ( P1_R1207_U284 , P1_U3066 , P1_R1207_U73 );
nand NAND2_14114 ( P1_R1207_U285 , P1_U3061 , P1_R1207_U48 );
nand NAND2_14115 ( P1_R1207_U286 , P1_R1207_U187 , P1_R1207_U181 );
nand NAND2_14116 ( P1_R1207_U287 , P1_R1207_U11 , P1_R1207_U286 );
nand NAND2_14117 ( P1_R1207_U288 , P1_U4024 , P1_R1207_U77 );
nand NAND2_14118 ( P1_R1207_U289 , P1_U4022 , P1_R1207_U75 );
nand NAND3_14119 ( P1_R1207_U290 , P1_R1207_U163 , P1_R1207_U127 , P1_R1207_U283 );
nand NAND2_14120 ( P1_R1207_U291 , P1_R1207_U289 , P1_R1207_U287 );
not NOT1_14121 ( P1_R1207_U292 , P1_R1207_U160 );
nand NAND2_14122 ( P1_R1207_U293 , P1_U4021 , P1_R1207_U80 );
nand NAND2_14123 ( P1_R1207_U294 , P1_R1207_U293 , P1_R1207_U160 );
nand NAND2_14124 ( P1_R1207_U295 , P1_U3065 , P1_R1207_U79 );
not NOT1_14125 ( P1_R1207_U296 , P1_R1207_U159 );
nand NAND2_14126 ( P1_R1207_U297 , P1_U4020 , P1_R1207_U82 );
nand NAND2_14127 ( P1_R1207_U298 , P1_R1207_U297 , P1_R1207_U159 );
nand NAND2_14128 ( P1_R1207_U299 , P1_U3058 , P1_R1207_U81 );
not NOT1_14129 ( P1_R1207_U300 , P1_R1207_U89 );
nand NAND2_14130 ( P1_R1207_U301 , P1_U4018 , P1_R1207_U86 );
nand NAND3_14131 ( P1_R1207_U302 , P1_R1207_U89 , P1_R1207_U182 , P1_R1207_U301 );
nand NAND2_14132 ( P1_R1207_U303 , P1_R1207_U86 , P1_R1207_U85 );
nand NAND2_14133 ( P1_R1207_U304 , P1_R1207_U303 , P1_R1207_U83 );
nand NAND2_14134 ( P1_R1207_U305 , P1_U3053 , P1_R1207_U176 );
not NOT1_14135 ( P1_R1207_U306 , P1_R1207_U157 );
nand NAND2_14136 ( P1_R1207_U307 , P1_U4017 , P1_R1207_U88 );
nand NAND2_14137 ( P1_R1207_U308 , P1_U3054 , P1_R1207_U87 );
nand NAND2_14138 ( P1_R1207_U309 , P1_R1207_U300 , P1_R1207_U85 );
nand NAND2_14139 ( P1_R1207_U310 , P1_R1207_U133 , P1_R1207_U309 );
nand NAND2_14140 ( P1_R1207_U311 , P1_R1207_U89 , P1_R1207_U182 );
nand NAND2_14141 ( P1_R1207_U312 , P1_R1207_U132 , P1_R1207_U311 );
nand NAND2_14142 ( P1_R1207_U313 , P1_R1207_U85 , P1_R1207_U182 );
nand NAND2_14143 ( P1_R1207_U314 , P1_R1207_U288 , P1_R1207_U163 );
not NOT1_14144 ( P1_R1207_U315 , P1_R1207_U90 );
nand NAND2_14145 ( P1_R1207_U316 , P1_U3061 , P1_R1207_U48 );
nand NAND2_14146 ( P1_R1207_U317 , P1_R1207_U315 , P1_R1207_U316 );
nand NAND2_14147 ( P1_R1207_U318 , P1_R1207_U136 , P1_R1207_U317 );
nand NAND2_14148 ( P1_R1207_U319 , P1_R1207_U90 , P1_R1207_U181 );
nand NAND2_14149 ( P1_R1207_U320 , P1_U4022 , P1_R1207_U75 );
nand NAND3_14150 ( P1_R1207_U321 , P1_R1207_U320 , P1_R1207_U319 , P1_R1207_U11 );
nand NAND2_14151 ( P1_R1207_U322 , P1_U3061 , P1_R1207_U48 );
nand NAND2_14152 ( P1_R1207_U323 , P1_R1207_U181 , P1_R1207_U322 );
nand NAND2_14153 ( P1_R1207_U324 , P1_R1207_U288 , P1_R1207_U78 );
nand NAND2_14154 ( P1_R1207_U325 , P1_R1207_U262 , P1_R1207_U171 );
not NOT1_14155 ( P1_R1207_U326 , P1_R1207_U91 );
nand NAND2_14156 ( P1_R1207_U327 , P1_U3074 , P1_R1207_U49 );
nand NAND2_14157 ( P1_R1207_U328 , P1_R1207_U326 , P1_R1207_U327 );
nand NAND2_14158 ( P1_R1207_U329 , P1_R1207_U142 , P1_R1207_U328 );
nand NAND2_14159 ( P1_R1207_U330 , P1_R1207_U91 , P1_R1207_U180 );
nand NAND2_14160 ( P1_R1207_U331 , P1_U3506 , P1_R1207_U61 );
nand NAND3_14161 ( P1_R1207_U332 , P1_R1207_U331 , P1_R1207_U330 , P1_R1207_U10 );
nand NAND2_14162 ( P1_R1207_U333 , P1_U3074 , P1_R1207_U49 );
nand NAND2_14163 ( P1_R1207_U334 , P1_R1207_U180 , P1_R1207_U333 );
nand NAND2_14164 ( P1_R1207_U335 , P1_R1207_U262 , P1_R1207_U64 );
nand NAND2_14165 ( P1_R1207_U336 , P1_R1207_U217 , P1_R1207_U148 );
not NOT1_14166 ( P1_R1207_U337 , P1_R1207_U92 );
nand NAND2_14167 ( P1_R1207_U338 , P1_U3062 , P1_R1207_U51 );
nand NAND2_14168 ( P1_R1207_U339 , P1_R1207_U337 , P1_R1207_U338 );
nand NAND2_14169 ( P1_R1207_U340 , P1_R1207_U146 , P1_R1207_U339 );
nand NAND2_14170 ( P1_R1207_U341 , P1_R1207_U92 , P1_R1207_U179 );
nand NAND2_14171 ( P1_R1207_U342 , P1_U3491 , P1_R1207_U52 );
nand NAND2_14172 ( P1_R1207_U343 , P1_R1207_U145 , P1_R1207_U341 );
nand NAND2_14173 ( P1_R1207_U344 , P1_U3062 , P1_R1207_U51 );
nand NAND2_14174 ( P1_R1207_U345 , P1_R1207_U179 , P1_R1207_U344 );
nand NAND2_14175 ( P1_R1207_U346 , P1_U3077 , P1_R1207_U24 );
nand NAND3_14176 ( P1_R1207_U347 , P1_R1207_U89 , P1_R1207_U182 , P1_R1207_U301 );
nand NAND3_14177 ( P1_R1207_U348 , P1_R1207_U12 , P1_R1207_U347 , P1_R1207_U130 );
nand NAND2_14178 ( P1_R1207_U349 , P1_U3485 , P1_R1207_U43 );
nand NAND2_14179 ( P1_R1207_U350 , P1_U3083 , P1_R1207_U42 );
nand NAND2_14180 ( P1_R1207_U351 , P1_R1207_U218 , P1_R1207_U148 );
nand NAND2_14181 ( P1_R1207_U352 , P1_R1207_U216 , P1_R1207_U147 );
nand NAND2_14182 ( P1_R1207_U353 , P1_U3482 , P1_R1207_U41 );
nand NAND2_14183 ( P1_R1207_U354 , P1_U3084 , P1_R1207_U38 );
nand NAND2_14184 ( P1_R1207_U355 , P1_U3482 , P1_R1207_U41 );
nand NAND2_14185 ( P1_R1207_U356 , P1_U3084 , P1_R1207_U38 );
nand NAND2_14186 ( P1_R1207_U357 , P1_R1207_U356 , P1_R1207_U355 );
nand NAND2_14187 ( P1_R1207_U358 , P1_U3479 , P1_R1207_U39 );
nand NAND2_14188 ( P1_R1207_U359 , P1_U3070 , P1_R1207_U22 );
nand NAND2_14189 ( P1_R1207_U360 , P1_R1207_U223 , P1_R1207_U44 );
nand NAND2_14190 ( P1_R1207_U361 , P1_R1207_U149 , P1_R1207_U210 );
nand NAND2_14191 ( P1_R1207_U362 , P1_U3476 , P1_R1207_U34 );
nand NAND2_14192 ( P1_R1207_U363 , P1_U3071 , P1_R1207_U31 );
nand NAND2_14193 ( P1_R1207_U364 , P1_R1207_U363 , P1_R1207_U362 );
nand NAND2_14194 ( P1_R1207_U365 , P1_U3473 , P1_R1207_U35 );
nand NAND2_14195 ( P1_R1207_U366 , P1_U3067 , P1_R1207_U32 );
nand NAND2_14196 ( P1_R1207_U367 , P1_R1207_U233 , P1_R1207_U45 );
nand NAND2_14197 ( P1_R1207_U368 , P1_R1207_U150 , P1_R1207_U225 );
nand NAND2_14198 ( P1_R1207_U369 , P1_U3470 , P1_R1207_U36 );
nand NAND2_14199 ( P1_R1207_U370 , P1_U3060 , P1_R1207_U33 );
nand NAND2_14200 ( P1_R1207_U371 , P1_R1207_U234 , P1_R1207_U152 );
nand NAND2_14201 ( P1_R1207_U372 , P1_R1207_U200 , P1_R1207_U151 );
nand NAND2_14202 ( P1_R1207_U373 , P1_U3467 , P1_R1207_U30 );
nand NAND2_14203 ( P1_R1207_U374 , P1_U3064 , P1_R1207_U27 );
nand NAND2_14204 ( P1_R1207_U375 , P1_U3467 , P1_R1207_U30 );
nand NAND2_14205 ( P1_R1207_U376 , P1_U3064 , P1_R1207_U27 );
nand NAND2_14206 ( P1_R1207_U377 , P1_R1207_U376 , P1_R1207_U375 );
nand NAND2_14207 ( P1_R1207_U378 , P1_U3464 , P1_R1207_U28 );
nand NAND2_14208 ( P1_R1207_U379 , P1_U3068 , P1_R1207_U23 );
nand NAND2_14209 ( P1_R1207_U380 , P1_R1207_U239 , P1_R1207_U46 );
nand NAND2_14210 ( P1_R1207_U381 , P1_R1207_U153 , P1_R1207_U194 );
nand NAND2_14211 ( P1_R1207_U382 , P1_U4028 , P1_R1207_U155 );
nand NAND2_14212 ( P1_R1207_U383 , P1_U3055 , P1_R1207_U154 );
nand NAND2_14213 ( P1_R1207_U384 , P1_U4028 , P1_R1207_U155 );
nand NAND2_14214 ( P1_R1207_U385 , P1_U3055 , P1_R1207_U154 );
nand NAND2_14215 ( P1_R1207_U386 , P1_R1207_U385 , P1_R1207_U384 );
nand NAND3_14216 ( P1_R1207_U387 , P1_U3054 , P1_R1207_U386 , P1_R1207_U87 );
nand NAND3_14217 ( P1_R1207_U388 , P1_R1207_U12 , P1_R1207_U88 , P1_U4017 );
nand NAND2_14218 ( P1_R1207_U389 , P1_U4017 , P1_R1207_U88 );
nand NAND2_14219 ( P1_R1207_U390 , P1_U3054 , P1_R1207_U87 );
not NOT1_14220 ( P1_R1207_U391 , P1_R1207_U131 );
nand NAND2_14221 ( P1_R1207_U392 , P1_R1207_U306 , P1_R1207_U391 );
nand NAND2_14222 ( P1_R1207_U393 , P1_R1207_U131 , P1_R1207_U157 );
nand NAND2_14223 ( P1_R1207_U394 , P1_U4018 , P1_R1207_U86 );
nand NAND2_14224 ( P1_R1207_U395 , P1_U3053 , P1_R1207_U83 );
nand NAND2_14225 ( P1_R1207_U396 , P1_U4018 , P1_R1207_U86 );
nand NAND2_14226 ( P1_R1207_U397 , P1_U3053 , P1_R1207_U83 );
nand NAND2_14227 ( P1_R1207_U398 , P1_R1207_U397 , P1_R1207_U396 );
nand NAND2_14228 ( P1_R1207_U399 , P1_U4019 , P1_R1207_U84 );
nand NAND2_14229 ( P1_R1207_U400 , P1_U3057 , P1_R1207_U47 );
nand NAND2_14230 ( P1_R1207_U401 , P1_R1207_U313 , P1_R1207_U89 );
nand NAND2_14231 ( P1_R1207_U402 , P1_R1207_U158 , P1_R1207_U300 );
nand NAND2_14232 ( P1_R1207_U403 , P1_U4020 , P1_R1207_U82 );
nand NAND2_14233 ( P1_R1207_U404 , P1_U3058 , P1_R1207_U81 );
not NOT1_14234 ( P1_R1207_U405 , P1_R1207_U134 );
nand NAND2_14235 ( P1_R1207_U406 , P1_R1207_U296 , P1_R1207_U405 );
nand NAND2_14236 ( P1_R1207_U407 , P1_R1207_U134 , P1_R1207_U159 );
nand NAND2_14237 ( P1_R1207_U408 , P1_U4021 , P1_R1207_U80 );
nand NAND2_14238 ( P1_R1207_U409 , P1_U3065 , P1_R1207_U79 );
not NOT1_14239 ( P1_R1207_U410 , P1_R1207_U135 );
nand NAND2_14240 ( P1_R1207_U411 , P1_R1207_U292 , P1_R1207_U410 );
nand NAND2_14241 ( P1_R1207_U412 , P1_R1207_U135 , P1_R1207_U160 );
nand NAND2_14242 ( P1_R1207_U413 , P1_U4022 , P1_R1207_U75 );
nand NAND2_14243 ( P1_R1207_U414 , P1_U3066 , P1_R1207_U73 );
nand NAND2_14244 ( P1_R1207_U415 , P1_R1207_U414 , P1_R1207_U413 );
nand NAND2_14245 ( P1_R1207_U416 , P1_U4023 , P1_R1207_U76 );
nand NAND2_14246 ( P1_R1207_U417 , P1_U3061 , P1_R1207_U48 );
nand NAND2_14247 ( P1_R1207_U418 , P1_R1207_U323 , P1_R1207_U90 );
nand NAND2_14248 ( P1_R1207_U419 , P1_R1207_U161 , P1_R1207_U315 );
nand NAND2_14249 ( P1_R1207_U420 , P1_U4024 , P1_R1207_U77 );
nand NAND2_14250 ( P1_R1207_U421 , P1_U3075 , P1_R1207_U74 );
nand NAND2_14251 ( P1_R1207_U422 , P1_R1207_U324 , P1_R1207_U163 );
nand NAND2_14252 ( P1_R1207_U423 , P1_R1207_U282 , P1_R1207_U162 );
nand NAND2_14253 ( P1_R1207_U424 , P1_U4025 , P1_R1207_U72 );
nand NAND2_14254 ( P1_R1207_U425 , P1_U3076 , P1_R1207_U71 );
not NOT1_14255 ( P1_R1207_U426 , P1_R1207_U137 );
nand NAND2_14256 ( P1_R1207_U427 , P1_R1207_U278 , P1_R1207_U426 );
nand NAND2_14257 ( P1_R1207_U428 , P1_R1207_U137 , P1_R1207_U164 );
nand NAND2_14258 ( P1_R1207_U429 , P1_U3461 , P1_R1207_U26 );
nand NAND2_14259 ( P1_R1207_U430 , P1_U3078 , P1_R1207_U165 );
not NOT1_14260 ( P1_R1207_U431 , P1_R1207_U138 );
nand NAND2_14261 ( P1_R1207_U432 , P1_R1207_U431 , P1_R1207_U190 );
nand NAND2_14262 ( P1_R1207_U433 , P1_R1207_U138 , P1_R1207_U25 );
nand NAND2_14263 ( P1_R1207_U434 , P1_U3514 , P1_R1207_U70 );
nand NAND2_14264 ( P1_R1207_U435 , P1_U3081 , P1_R1207_U69 );
not NOT1_14265 ( P1_R1207_U436 , P1_R1207_U139 );
nand NAND2_14266 ( P1_R1207_U437 , P1_R1207_U274 , P1_R1207_U436 );
nand NAND2_14267 ( P1_R1207_U438 , P1_R1207_U139 , P1_R1207_U166 );
nand NAND2_14268 ( P1_R1207_U439 , P1_U3512 , P1_R1207_U68 );
nand NAND2_14269 ( P1_R1207_U440 , P1_U3082 , P1_R1207_U167 );
not NOT1_14270 ( P1_R1207_U441 , P1_R1207_U140 );
nand NAND2_14271 ( P1_R1207_U442 , P1_R1207_U441 , P1_R1207_U270 );
nand NAND2_14272 ( P1_R1207_U443 , P1_R1207_U140 , P1_R1207_U67 );
nand NAND2_14273 ( P1_R1207_U444 , P1_U3509 , P1_R1207_U66 );
nand NAND2_14274 ( P1_R1207_U445 , P1_U3069 , P1_R1207_U65 );
not NOT1_14275 ( P1_R1207_U446 , P1_R1207_U141 );
nand NAND2_14276 ( P1_R1207_U447 , P1_R1207_U266 , P1_R1207_U446 );
nand NAND2_14277 ( P1_R1207_U448 , P1_R1207_U141 , P1_R1207_U168 );
nand NAND2_14278 ( P1_R1207_U449 , P1_U3506 , P1_R1207_U61 );
nand NAND2_14279 ( P1_R1207_U450 , P1_U3073 , P1_R1207_U59 );
nand NAND2_14280 ( P1_R1207_U451 , P1_R1207_U450 , P1_R1207_U449 );
nand NAND2_14281 ( P1_R1207_U452 , P1_U3503 , P1_R1207_U62 );
nand NAND2_14282 ( P1_R1207_U453 , P1_U3074 , P1_R1207_U49 );
nand NAND2_14283 ( P1_R1207_U454 , P1_R1207_U334 , P1_R1207_U91 );
nand NAND2_14284 ( P1_R1207_U455 , P1_R1207_U169 , P1_R1207_U326 );
nand NAND2_14285 ( P1_R1207_U456 , P1_U3500 , P1_R1207_U63 );
nand NAND2_14286 ( P1_R1207_U457 , P1_U3079 , P1_R1207_U60 );
nand NAND2_14287 ( P1_R1207_U458 , P1_R1207_U335 , P1_R1207_U171 );
nand NAND2_14288 ( P1_R1207_U459 , P1_R1207_U256 , P1_R1207_U170 );
nand NAND2_14289 ( P1_R1207_U460 , P1_U3497 , P1_R1207_U58 );
nand NAND2_14290 ( P1_R1207_U461 , P1_U3080 , P1_R1207_U57 );
not NOT1_14291 ( P1_R1207_U462 , P1_R1207_U143 );
nand NAND2_14292 ( P1_R1207_U463 , P1_R1207_U252 , P1_R1207_U462 );
nand NAND2_14293 ( P1_R1207_U464 , P1_R1207_U143 , P1_R1207_U172 );
nand NAND2_14294 ( P1_R1207_U465 , P1_U3494 , P1_R1207_U56 );
nand NAND2_14295 ( P1_R1207_U466 , P1_U3072 , P1_R1207_U55 );
not NOT1_14296 ( P1_R1207_U467 , P1_R1207_U144 );
nand NAND2_14297 ( P1_R1207_U468 , P1_R1207_U248 , P1_R1207_U467 );
nand NAND2_14298 ( P1_R1207_U469 , P1_R1207_U144 , P1_R1207_U173 );
nand NAND2_14299 ( P1_R1207_U470 , P1_U3491 , P1_R1207_U52 );
nand NAND2_14300 ( P1_R1207_U471 , P1_U3063 , P1_R1207_U50 );
nand NAND2_14301 ( P1_R1207_U472 , P1_R1207_U471 , P1_R1207_U470 );
nand NAND2_14302 ( P1_R1207_U473 , P1_U3488 , P1_R1207_U53 );
nand NAND2_14303 ( P1_R1207_U474 , P1_U3062 , P1_R1207_U51 );
nand NAND2_14304 ( P1_R1207_U475 , P1_R1207_U345 , P1_R1207_U92 );
nand NAND2_14305 ( P1_R1207_U476 , P1_R1207_U174 , P1_R1207_U337 );
and AND2_14306 ( P1_R1165_U4 , P1_R1165_U202 , P1_R1165_U201 );
and AND2_14307 ( P1_R1165_U5 , P1_R1165_U217 , P1_R1165_U216 );
and AND2_14308 ( P1_R1165_U6 , P1_R1165_U251 , P1_R1165_U250 );
and AND2_14309 ( P1_R1165_U7 , P1_R1165_U269 , P1_R1165_U268 );
and AND2_14310 ( P1_R1165_U8 , P1_R1165_U281 , P1_R1165_U280 );
and AND2_14311 ( P1_R1165_U9 , P1_R1165_U339 , P1_R1165_U336 );
and AND2_14312 ( P1_R1165_U10 , P1_R1165_U330 , P1_R1165_U327 );
and AND2_14313 ( P1_R1165_U11 , P1_R1165_U323 , P1_R1165_U320 );
and AND2_14314 ( P1_R1165_U12 , P1_R1165_U314 , P1_R1165_U311 );
and AND2_14315 ( P1_R1165_U13 , P1_R1165_U240 , P1_R1165_U237 );
and AND2_14316 ( P1_R1165_U14 , P1_R1165_U233 , P1_R1165_U230 );
not NOT1_14317 ( P1_R1165_U15 , P1_U3211 );
not NOT1_14318 ( P1_R1165_U16 , P1_U3175 );
nand NAND2_14319 ( P1_R1165_U17 , P1_U3175 , P1_R1165_U59 );
not NOT1_14320 ( P1_R1165_U18 , P1_U3174 );
not NOT1_14321 ( P1_R1165_U19 , P1_U3179 );
nand NAND2_14322 ( P1_R1165_U20 , P1_U3179 , P1_R1165_U61 );
not NOT1_14323 ( P1_R1165_U21 , P1_U3178 );
not NOT1_14324 ( P1_R1165_U22 , P1_U3181 );
not NOT1_14325 ( P1_R1165_U23 , P1_U3180 );
nand NAND2_14326 ( P1_R1165_U24 , P1_R1165_U110 , P1_R1165_U206 );
not NOT1_14327 ( P1_R1165_U25 , P1_U3177 );
not NOT1_14328 ( P1_R1165_U26 , P1_U3176 );
not NOT1_14329 ( P1_R1165_U27 , P1_U3173 );
not NOT1_14330 ( P1_R1165_U28 , P1_U3172 );
nand NAND2_14331 ( P1_R1165_U29 , P1_R1165_U226 , P1_R1165_U225 );
nand NAND2_14332 ( P1_R1165_U30 , P1_R1165_U214 , P1_R1165_U213 );
nand NAND2_14333 ( P1_R1165_U31 , P1_R1165_U199 , P1_R1165_U198 );
not NOT1_14334 ( P1_R1165_U32 , P1_U3154 );
not NOT1_14335 ( P1_R1165_U33 , P1_U3155 );
not NOT1_14336 ( P1_R1165_U34 , P1_U3156 );
not NOT1_14337 ( P1_R1165_U35 , P1_U3157 );
not NOT1_14338 ( P1_R1165_U36 , P1_U3160 );
not NOT1_14339 ( P1_R1165_U37 , P1_U3165 );
nand NAND2_14340 ( P1_R1165_U38 , P1_U3165 , P1_R1165_U73 );
not NOT1_14341 ( P1_R1165_U39 , P1_U3164 );
not NOT1_14342 ( P1_R1165_U40 , P1_U3171 );
not NOT1_14343 ( P1_R1165_U41 , P1_U3169 );
not NOT1_14344 ( P1_R1165_U42 , P1_U3170 );
nand NAND2_14345 ( P1_R1165_U43 , P1_U3170 , P1_R1165_U76 );
not NOT1_14346 ( P1_R1165_U44 , P1_U3168 );
not NOT1_14347 ( P1_R1165_U45 , P1_U3167 );
not NOT1_14348 ( P1_R1165_U46 , P1_U3166 );
not NOT1_14349 ( P1_R1165_U47 , P1_U3163 );
not NOT1_14350 ( P1_R1165_U48 , P1_U3162 );
nand NAND2_14351 ( P1_R1165_U49 , P1_U3162 , P1_R1165_U82 );
not NOT1_14352 ( P1_R1165_U50 , P1_U3161 );
not NOT1_14353 ( P1_R1165_U51 , P1_U3159 );
not NOT1_14354 ( P1_R1165_U52 , P1_U3158 );
nand NAND2_14355 ( P1_R1165_U53 , P1_U3155 , P1_R1165_U70 );
nand NAND2_14356 ( P1_R1165_U54 , P1_R1165_U192 , P1_R1165_U307 );
nand NAND2_14357 ( P1_R1165_U55 , P1_R1165_U49 , P1_R1165_U316 );
nand NAND2_14358 ( P1_R1165_U56 , P1_R1165_U266 , P1_R1165_U265 );
nand NAND2_14359 ( P1_R1165_U57 , P1_R1165_U43 , P1_R1165_U332 );
nand NAND2_14360 ( P1_R1165_U58 , P1_R1165_U359 , P1_R1165_U358 );
nand NAND2_14361 ( P1_R1165_U59 , P1_R1165_U388 , P1_R1165_U387 );
nand NAND2_14362 ( P1_R1165_U60 , P1_R1165_U385 , P1_R1165_U384 );
nand NAND2_14363 ( P1_R1165_U61 , P1_R1165_U376 , P1_R1165_U375 );
nand NAND2_14364 ( P1_R1165_U62 , P1_R1165_U373 , P1_R1165_U372 );
nand NAND2_14365 ( P1_R1165_U63 , P1_R1165_U367 , P1_R1165_U366 );
nand NAND2_14366 ( P1_R1165_U64 , P1_R1165_U370 , P1_R1165_U369 );
nand NAND2_14367 ( P1_R1165_U65 , P1_R1165_U379 , P1_R1165_U378 );
nand NAND2_14368 ( P1_R1165_U66 , P1_R1165_U382 , P1_R1165_U381 );
nand NAND2_14369 ( P1_R1165_U67 , P1_R1165_U391 , P1_R1165_U390 );
nand NAND2_14370 ( P1_R1165_U68 , P1_R1165_U431 , P1_R1165_U430 );
nand NAND2_14371 ( P1_R1165_U69 , P1_R1165_U434 , P1_R1165_U433 );
nand NAND2_14372 ( P1_R1165_U70 , P1_R1165_U437 , P1_R1165_U436 );
nand NAND2_14373 ( P1_R1165_U71 , P1_R1165_U440 , P1_R1165_U439 );
nand NAND2_14374 ( P1_R1165_U72 , P1_R1165_U443 , P1_R1165_U442 );
nand NAND2_14375 ( P1_R1165_U73 , P1_R1165_U473 , P1_R1165_U472 );
nand NAND2_14376 ( P1_R1165_U74 , P1_R1165_U470 , P1_R1165_U469 );
nand NAND2_14377 ( P1_R1165_U75 , P1_R1165_U452 , P1_R1165_U451 );
nand NAND2_14378 ( P1_R1165_U76 , P1_R1165_U461 , P1_R1165_U460 );
nand NAND2_14379 ( P1_R1165_U77 , P1_R1165_U455 , P1_R1165_U454 );
nand NAND2_14380 ( P1_R1165_U78 , P1_R1165_U458 , P1_R1165_U457 );
nand NAND2_14381 ( P1_R1165_U79 , P1_R1165_U464 , P1_R1165_U463 );
nand NAND2_14382 ( P1_R1165_U80 , P1_R1165_U467 , P1_R1165_U466 );
nand NAND2_14383 ( P1_R1165_U81 , P1_R1165_U476 , P1_R1165_U475 );
nand NAND2_14384 ( P1_R1165_U82 , P1_R1165_U449 , P1_R1165_U448 );
nand NAND2_14385 ( P1_R1165_U83 , P1_R1165_U446 , P1_R1165_U445 );
nand NAND2_14386 ( P1_R1165_U84 , P1_R1165_U479 , P1_R1165_U478 );
nand NAND2_14387 ( P1_R1165_U85 , P1_R1165_U482 , P1_R1165_U481 );
nand NAND2_14388 ( P1_R1165_U86 , P1_R1165_U488 , P1_R1165_U487 );
nand NAND2_14389 ( P1_R1165_U87 , P1_R1165_U595 , P1_R1165_U594 );
nand NAND2_14390 ( P1_R1165_U88 , P1_R1165_U394 , P1_R1165_U393 );
nand NAND2_14391 ( P1_R1165_U89 , P1_R1165_U401 , P1_R1165_U400 );
nand NAND2_14392 ( P1_R1165_U90 , P1_R1165_U408 , P1_R1165_U407 );
nand NAND2_14393 ( P1_R1165_U91 , P1_R1165_U415 , P1_R1165_U414 );
nand NAND2_14394 ( P1_R1165_U92 , P1_R1165_U422 , P1_R1165_U421 );
nand NAND2_14395 ( P1_R1165_U93 , P1_R1165_U429 , P1_R1165_U428 );
nand NAND2_14396 ( P1_R1165_U94 , P1_R1165_U491 , P1_R1165_U490 );
nand NAND2_14397 ( P1_R1165_U95 , P1_R1165_U498 , P1_R1165_U497 );
nand NAND2_14398 ( P1_R1165_U96 , P1_R1165_U505 , P1_R1165_U504 );
nand NAND2_14399 ( P1_R1165_U97 , P1_R1165_U510 , P1_R1165_U509 );
nand NAND2_14400 ( P1_R1165_U98 , P1_R1165_U517 , P1_R1165_U516 );
nand NAND2_14401 ( P1_R1165_U99 , P1_R1165_U524 , P1_R1165_U523 );
nand NAND2_14402 ( P1_R1165_U100 , P1_R1165_U531 , P1_R1165_U530 );
nand NAND2_14403 ( P1_R1165_U101 , P1_R1165_U538 , P1_R1165_U537 );
nand NAND2_14404 ( P1_R1165_U102 , P1_R1165_U543 , P1_R1165_U542 );
nand NAND2_14405 ( P1_R1165_U103 , P1_R1165_U550 , P1_R1165_U549 );
nand NAND2_14406 ( P1_R1165_U104 , P1_R1165_U557 , P1_R1165_U556 );
nand NAND2_14407 ( P1_R1165_U105 , P1_R1165_U564 , P1_R1165_U563 );
nand NAND2_14408 ( P1_R1165_U106 , P1_R1165_U571 , P1_R1165_U570 );
nand NAND2_14409 ( P1_R1165_U107 , P1_R1165_U578 , P1_R1165_U577 );
nand NAND2_14410 ( P1_R1165_U108 , P1_R1165_U583 , P1_R1165_U582 );
nand NAND2_14411 ( P1_R1165_U109 , P1_R1165_U590 , P1_R1165_U589 );
and AND2_14412 ( P1_R1165_U110 , P1_R1165_U205 , P1_R1165_U204 );
and AND2_14413 ( P1_R1165_U111 , P1_R1165_U221 , P1_R1165_U220 );
and AND3_14414 ( P1_R1165_U112 , P1_R1165_U403 , P1_R1165_U402 , P1_R1165_U17 );
and AND2_14415 ( P1_R1165_U113 , P1_R1165_U232 , P1_R1165_U5 );
and AND3_14416 ( P1_R1165_U114 , P1_R1165_U424 , P1_R1165_U423 , P1_R1165_U20 );
and AND2_14417 ( P1_R1165_U115 , P1_R1165_U239 , P1_R1165_U4 );
and AND2_14418 ( P1_R1165_U116 , P1_R1165_U255 , P1_R1165_U6 );
and AND2_14419 ( P1_R1165_U117 , P1_R1165_U253 , P1_R1165_U187 );
and AND2_14420 ( P1_R1165_U118 , P1_R1165_U273 , P1_R1165_U272 );
and AND2_14421 ( P1_R1165_U119 , P1_R1165_U357 , P1_R1165_U53 );
and AND2_14422 ( P1_R1165_U120 , P1_R1165_U306 , P1_R1165_U301 );
and AND2_14423 ( P1_R1165_U121 , P1_R1165_U354 , P1_R1165_U305 );
nand NAND2_14424 ( P1_R1165_U122 , P1_R1165_U485 , P1_R1165_U484 );
and AND3_14425 ( P1_R1165_U123 , P1_R1165_U500 , P1_R1165_U499 , P1_R1165_U189 );
and AND3_14426 ( P1_R1165_U124 , P1_R1165_U526 , P1_R1165_U525 , P1_R1165_U188 );
and AND3_14427 ( P1_R1165_U125 , P1_R1165_U552 , P1_R1165_U551 , P1_R1165_U38 );
and AND2_14428 ( P1_R1165_U126 , P1_R1165_U329 , P1_R1165_U7 );
and AND3_14429 ( P1_R1165_U127 , P1_R1165_U573 , P1_R1165_U572 , P1_R1165_U187 );
and AND2_14430 ( P1_R1165_U128 , P1_R1165_U338 , P1_R1165_U6 );
nand NAND2_14431 ( P1_R1165_U129 , P1_R1165_U592 , P1_R1165_U591 );
not NOT1_14432 ( P1_R1165_U130 , P1_U3201 );
and AND2_14433 ( P1_R1165_U131 , P1_R1165_U362 , P1_R1165_U361 );
not NOT1_14434 ( P1_R1165_U132 , P1_U3210 );
not NOT1_14435 ( P1_R1165_U133 , P1_U3209 );
not NOT1_14436 ( P1_R1165_U134 , P1_U3207 );
not NOT1_14437 ( P1_R1165_U135 , P1_U3208 );
not NOT1_14438 ( P1_R1165_U136 , P1_U3206 );
not NOT1_14439 ( P1_R1165_U137 , P1_U3205 );
not NOT1_14440 ( P1_R1165_U138 , P1_U3203 );
not NOT1_14441 ( P1_R1165_U139 , P1_U3204 );
not NOT1_14442 ( P1_R1165_U140 , P1_U3202 );
and AND2_14443 ( P1_R1165_U141 , P1_R1165_U396 , P1_R1165_U395 );
nand NAND2_14444 ( P1_R1165_U142 , P1_R1165_U111 , P1_R1165_U222 );
and AND2_14445 ( P1_R1165_U143 , P1_R1165_U410 , P1_R1165_U409 );
nand NAND2_14446 ( P1_R1165_U144 , P1_R1165_U210 , P1_R1165_U209 );
and AND2_14447 ( P1_R1165_U145 , P1_R1165_U417 , P1_R1165_U416 );
not NOT1_14448 ( P1_R1165_U146 , P1_U3183 );
not NOT1_14449 ( P1_R1165_U147 , P1_U3185 );
not NOT1_14450 ( P1_R1165_U148 , P1_U3184 );
not NOT1_14451 ( P1_R1165_U149 , P1_U3186 );
not NOT1_14452 ( P1_R1165_U150 , P1_U3189 );
not NOT1_14453 ( P1_R1165_U151 , P1_U3190 );
not NOT1_14454 ( P1_R1165_U152 , P1_U3191 );
not NOT1_14455 ( P1_R1165_U153 , P1_U3200 );
not NOT1_14456 ( P1_R1165_U154 , P1_U3197 );
not NOT1_14457 ( P1_R1165_U155 , P1_U3198 );
not NOT1_14458 ( P1_R1165_U156 , P1_U3199 );
not NOT1_14459 ( P1_R1165_U157 , P1_U3196 );
not NOT1_14460 ( P1_R1165_U158 , P1_U3195 );
not NOT1_14461 ( P1_R1165_U159 , P1_U3193 );
not NOT1_14462 ( P1_R1165_U160 , P1_U3194 );
not NOT1_14463 ( P1_R1165_U161 , P1_U3192 );
not NOT1_14464 ( P1_R1165_U162 , P1_U3188 );
not NOT1_14465 ( P1_R1165_U163 , P1_U3187 );
not NOT1_14466 ( P1_R1165_U164 , P1_U3153 );
not NOT1_14467 ( P1_R1165_U165 , P1_U3182 );
and AND2_14468 ( P1_R1165_U166 , P1_R1165_U493 , P1_R1165_U492 );
nand NAND3_14469 ( P1_R1165_U167 , P1_R1165_U351 , P1_R1165_U302 , P1_R1165_U53 );
nand NAND2_14470 ( P1_R1165_U168 , P1_R1165_U296 , P1_R1165_U295 );
and AND2_14471 ( P1_R1165_U169 , P1_R1165_U512 , P1_R1165_U511 );
nand NAND2_14472 ( P1_R1165_U170 , P1_R1165_U292 , P1_R1165_U291 );
and AND2_14473 ( P1_R1165_U171 , P1_R1165_U519 , P1_R1165_U518 );
nand NAND3_14474 ( P1_R1165_U172 , P1_R1165_U287 , P1_R1165_U283 , P1_R1165_U288 );
and AND2_14475 ( P1_R1165_U173 , P1_R1165_U533 , P1_R1165_U532 );
nand NAND2_14476 ( P1_R1165_U174 , P1_R1165_U195 , P1_R1165_U194 );
nand NAND2_14477 ( P1_R1165_U175 , P1_R1165_U278 , P1_R1165_U277 );
and AND2_14478 ( P1_R1165_U176 , P1_R1165_U545 , P1_R1165_U544 );
nand NAND2_14479 ( P1_R1165_U177 , P1_R1165_U118 , P1_R1165_U274 );
and AND2_14480 ( P1_R1165_U178 , P1_R1165_U559 , P1_R1165_U558 );
nand NAND2_14481 ( P1_R1165_U179 , P1_R1165_U262 , P1_R1165_U261 );
and AND2_14482 ( P1_R1165_U180 , P1_R1165_U566 , P1_R1165_U565 );
nand NAND2_14483 ( P1_R1165_U181 , P1_R1165_U258 , P1_R1165_U257 );
nand NAND2_14484 ( P1_R1165_U182 , P1_R1165_U248 , P1_R1165_U247 );
and AND2_14485 ( P1_R1165_U183 , P1_R1165_U585 , P1_R1165_U584 );
nand NAND2_14486 ( P1_R1165_U184 , P1_R1165_U244 , P1_R1165_U243 );
nand NAND2_14487 ( P1_R1165_U185 , P1_R1165_U353 , P1_R1165_U352 );
not NOT1_14488 ( P1_R1165_U186 , P1_R1165_U20 );
nand NAND2_14489 ( P1_R1165_U187 , P1_U3169 , P1_R1165_U78 );
nand NAND2_14490 ( P1_R1165_U188 , P1_U3161 , P1_R1165_U83 );
nand NAND2_14491 ( P1_R1165_U189 , P1_U3156 , P1_R1165_U69 );
not NOT1_14492 ( P1_R1165_U190 , P1_R1165_U43 );
not NOT1_14493 ( P1_R1165_U191 , P1_R1165_U49 );
nand NAND2_14494 ( P1_R1165_U192 , P1_U3157 , P1_R1165_U71 );
or OR2_14495 ( P1_R1165_U193 , P1_U3211 , P1_U3181 );
nand NAND2_14496 ( P1_R1165_U194 , P1_R1165_U63 , P1_R1165_U193 );
nand NAND2_14497 ( P1_R1165_U195 , P1_U3181 , P1_U3211 );
not NOT1_14498 ( P1_R1165_U196 , P1_R1165_U174 );
nand NAND2_14499 ( P1_R1165_U197 , P1_R1165_U371 , P1_R1165_U23 );
nand NAND2_14500 ( P1_R1165_U198 , P1_R1165_U197 , P1_R1165_U174 );
nand NAND2_14501 ( P1_R1165_U199 , P1_U3180 , P1_R1165_U64 );
not NOT1_14502 ( P1_R1165_U200 , P1_R1165_U31 );
nand NAND2_14503 ( P1_R1165_U201 , P1_R1165_U374 , P1_R1165_U21 );
nand NAND2_14504 ( P1_R1165_U202 , P1_R1165_U377 , P1_R1165_U19 );
nand NAND2_14505 ( P1_R1165_U203 , P1_R1165_U21 , P1_R1165_U20 );
nand NAND2_14506 ( P1_R1165_U204 , P1_R1165_U62 , P1_R1165_U203 );
nand NAND2_14507 ( P1_R1165_U205 , P1_U3178 , P1_R1165_U186 );
nand NAND2_14508 ( P1_R1165_U206 , P1_R1165_U4 , P1_R1165_U31 );
not NOT1_14509 ( P1_R1165_U207 , P1_R1165_U24 );
nand NAND2_14510 ( P1_R1165_U208 , P1_R1165_U207 , P1_R1165_U25 );
nand NAND2_14511 ( P1_R1165_U209 , P1_R1165_U65 , P1_R1165_U208 );
nand NAND2_14512 ( P1_R1165_U210 , P1_U3177 , P1_R1165_U24 );
not NOT1_14513 ( P1_R1165_U211 , P1_R1165_U144 );
nand NAND2_14514 ( P1_R1165_U212 , P1_R1165_U383 , P1_R1165_U26 );
nand NAND2_14515 ( P1_R1165_U213 , P1_R1165_U212 , P1_R1165_U144 );
nand NAND2_14516 ( P1_R1165_U214 , P1_U3176 , P1_R1165_U66 );
not NOT1_14517 ( P1_R1165_U215 , P1_R1165_U30 );
nand NAND2_14518 ( P1_R1165_U216 , P1_R1165_U386 , P1_R1165_U18 );
nand NAND2_14519 ( P1_R1165_U217 , P1_R1165_U389 , P1_R1165_U16 );
not NOT1_14520 ( P1_R1165_U218 , P1_R1165_U17 );
nand NAND2_14521 ( P1_R1165_U219 , P1_R1165_U18 , P1_R1165_U17 );
nand NAND2_14522 ( P1_R1165_U220 , P1_R1165_U60 , P1_R1165_U219 );
nand NAND2_14523 ( P1_R1165_U221 , P1_U3174 , P1_R1165_U218 );
nand NAND2_14524 ( P1_R1165_U222 , P1_R1165_U5 , P1_R1165_U30 );
not NOT1_14525 ( P1_R1165_U223 , P1_R1165_U142 );
nand NAND2_14526 ( P1_R1165_U224 , P1_R1165_U392 , P1_R1165_U27 );
nand NAND2_14527 ( P1_R1165_U225 , P1_R1165_U224 , P1_R1165_U142 );
nand NAND2_14528 ( P1_R1165_U226 , P1_U3173 , P1_R1165_U67 );
not NOT1_14529 ( P1_R1165_U227 , P1_R1165_U29 );
nand NAND2_14530 ( P1_R1165_U228 , P1_R1165_U389 , P1_R1165_U16 );
nand NAND2_14531 ( P1_R1165_U229 , P1_R1165_U228 , P1_R1165_U30 );
nand NAND2_14532 ( P1_R1165_U230 , P1_R1165_U112 , P1_R1165_U229 );
nand NAND2_14533 ( P1_R1165_U231 , P1_R1165_U215 , P1_R1165_U17 );
nand NAND2_14534 ( P1_R1165_U232 , P1_U3174 , P1_R1165_U60 );
nand NAND2_14535 ( P1_R1165_U233 , P1_R1165_U113 , P1_R1165_U231 );
nand NAND2_14536 ( P1_R1165_U234 , P1_R1165_U389 , P1_R1165_U16 );
nand NAND2_14537 ( P1_R1165_U235 , P1_R1165_U377 , P1_R1165_U19 );
nand NAND2_14538 ( P1_R1165_U236 , P1_R1165_U235 , P1_R1165_U31 );
nand NAND2_14539 ( P1_R1165_U237 , P1_R1165_U114 , P1_R1165_U236 );
nand NAND2_14540 ( P1_R1165_U238 , P1_R1165_U200 , P1_R1165_U20 );
nand NAND2_14541 ( P1_R1165_U239 , P1_U3178 , P1_R1165_U62 );
nand NAND2_14542 ( P1_R1165_U240 , P1_R1165_U115 , P1_R1165_U238 );
nand NAND2_14543 ( P1_R1165_U241 , P1_R1165_U377 , P1_R1165_U19 );
nand NAND2_14544 ( P1_R1165_U242 , P1_R1165_U227 , P1_R1165_U28 );
nand NAND2_14545 ( P1_R1165_U243 , P1_R1165_U58 , P1_R1165_U242 );
nand NAND2_14546 ( P1_R1165_U244 , P1_U3172 , P1_R1165_U29 );
not NOT1_14547 ( P1_R1165_U245 , P1_R1165_U184 );
nand NAND2_14548 ( P1_R1165_U246 , P1_R1165_U453 , P1_R1165_U40 );
nand NAND2_14549 ( P1_R1165_U247 , P1_R1165_U246 , P1_R1165_U184 );
nand NAND2_14550 ( P1_R1165_U248 , P1_U3171 , P1_R1165_U75 );
not NOT1_14551 ( P1_R1165_U249 , P1_R1165_U182 );
nand NAND2_14552 ( P1_R1165_U250 , P1_R1165_U456 , P1_R1165_U44 );
nand NAND2_14553 ( P1_R1165_U251 , P1_R1165_U459 , P1_R1165_U41 );
nand NAND2_14554 ( P1_R1165_U252 , P1_R1165_U190 , P1_R1165_U6 );
nand NAND2_14555 ( P1_R1165_U253 , P1_U3168 , P1_R1165_U77 );
nand NAND2_14556 ( P1_R1165_U254 , P1_R1165_U117 , P1_R1165_U252 );
nand NAND2_14557 ( P1_R1165_U255 , P1_R1165_U462 , P1_R1165_U42 );
nand NAND2_14558 ( P1_R1165_U256 , P1_R1165_U456 , P1_R1165_U44 );
nand NAND2_14559 ( P1_R1165_U257 , P1_R1165_U116 , P1_R1165_U182 );
nand NAND2_14560 ( P1_R1165_U258 , P1_R1165_U256 , P1_R1165_U254 );
not NOT1_14561 ( P1_R1165_U259 , P1_R1165_U181 );
nand NAND2_14562 ( P1_R1165_U260 , P1_R1165_U465 , P1_R1165_U45 );
nand NAND2_14563 ( P1_R1165_U261 , P1_R1165_U260 , P1_R1165_U181 );
nand NAND2_14564 ( P1_R1165_U262 , P1_U3167 , P1_R1165_U79 );
not NOT1_14565 ( P1_R1165_U263 , P1_R1165_U179 );
nand NAND2_14566 ( P1_R1165_U264 , P1_R1165_U468 , P1_R1165_U46 );
nand NAND2_14567 ( P1_R1165_U265 , P1_R1165_U264 , P1_R1165_U179 );
nand NAND2_14568 ( P1_R1165_U266 , P1_U3166 , P1_R1165_U80 );
not NOT1_14569 ( P1_R1165_U267 , P1_R1165_U56 );
nand NAND2_14570 ( P1_R1165_U268 , P1_R1165_U471 , P1_R1165_U39 );
nand NAND2_14571 ( P1_R1165_U269 , P1_R1165_U474 , P1_R1165_U37 );
not NOT1_14572 ( P1_R1165_U270 , P1_R1165_U38 );
nand NAND2_14573 ( P1_R1165_U271 , P1_R1165_U39 , P1_R1165_U38 );
nand NAND2_14574 ( P1_R1165_U272 , P1_R1165_U74 , P1_R1165_U271 );
nand NAND2_14575 ( P1_R1165_U273 , P1_U3164 , P1_R1165_U270 );
nand NAND2_14576 ( P1_R1165_U274 , P1_R1165_U7 , P1_R1165_U56 );
not NOT1_14577 ( P1_R1165_U275 , P1_R1165_U177 );
nand NAND2_14578 ( P1_R1165_U276 , P1_R1165_U477 , P1_R1165_U47 );
nand NAND2_14579 ( P1_R1165_U277 , P1_R1165_U276 , P1_R1165_U177 );
nand NAND2_14580 ( P1_R1165_U278 , P1_U3163 , P1_R1165_U81 );
not NOT1_14581 ( P1_R1165_U279 , P1_R1165_U175 );
nand NAND2_14582 ( P1_R1165_U280 , P1_R1165_U444 , P1_R1165_U36 );
nand NAND2_14583 ( P1_R1165_U281 , P1_R1165_U447 , P1_R1165_U50 );
nand NAND2_14584 ( P1_R1165_U282 , P1_R1165_U191 , P1_R1165_U8 );
nand NAND2_14585 ( P1_R1165_U283 , P1_U3160 , P1_R1165_U72 );
nand NAND2_14586 ( P1_R1165_U284 , P1_R1165_U188 , P1_R1165_U282 );
nand NAND2_14587 ( P1_R1165_U285 , P1_R1165_U450 , P1_R1165_U48 );
nand NAND2_14588 ( P1_R1165_U286 , P1_R1165_U444 , P1_R1165_U36 );
nand NAND3_14589 ( P1_R1165_U287 , P1_R1165_U285 , P1_R1165_U175 , P1_R1165_U8 );
nand NAND2_14590 ( P1_R1165_U288 , P1_R1165_U286 , P1_R1165_U284 );
not NOT1_14591 ( P1_R1165_U289 , P1_R1165_U172 );
nand NAND2_14592 ( P1_R1165_U290 , P1_R1165_U480 , P1_R1165_U51 );
nand NAND2_14593 ( P1_R1165_U291 , P1_R1165_U290 , P1_R1165_U172 );
nand NAND2_14594 ( P1_R1165_U292 , P1_U3159 , P1_R1165_U84 );
not NOT1_14595 ( P1_R1165_U293 , P1_R1165_U170 );
nand NAND2_14596 ( P1_R1165_U294 , P1_R1165_U483 , P1_R1165_U52 );
nand NAND2_14597 ( P1_R1165_U295 , P1_R1165_U294 , P1_R1165_U170 );
nand NAND2_14598 ( P1_R1165_U296 , P1_U3158 , P1_R1165_U85 );
not NOT1_14599 ( P1_R1165_U297 , P1_R1165_U168 );
nand NAND2_14600 ( P1_R1165_U298 , P1_R1165_U435 , P1_R1165_U34 );
nand NAND2_14601 ( P1_R1165_U299 , P1_R1165_U192 , P1_R1165_U189 );
not NOT1_14602 ( P1_R1165_U300 , P1_R1165_U53 );
nand NAND2_14603 ( P1_R1165_U301 , P1_R1165_U441 , P1_R1165_U35 );
nand NAND3_14604 ( P1_R1165_U302 , P1_R1165_U168 , P1_R1165_U301 , P1_R1165_U185 );
not NOT1_14605 ( P1_R1165_U303 , P1_R1165_U167 );
nand NAND2_14606 ( P1_R1165_U304 , P1_R1165_U432 , P1_R1165_U32 );
nand NAND2_14607 ( P1_R1165_U305 , P1_U3154 , P1_R1165_U68 );
nand NAND2_14608 ( P1_R1165_U306 , P1_R1165_U432 , P1_R1165_U32 );
nand NAND2_14609 ( P1_R1165_U307 , P1_R1165_U301 , P1_R1165_U168 );
not NOT1_14610 ( P1_R1165_U308 , P1_R1165_U54 );
nand NAND2_14611 ( P1_R1165_U309 , P1_R1165_U435 , P1_R1165_U34 );
nand NAND2_14612 ( P1_R1165_U310 , P1_R1165_U309 , P1_R1165_U54 );
nand NAND2_14613 ( P1_R1165_U311 , P1_R1165_U123 , P1_R1165_U310 );
nand NAND2_14614 ( P1_R1165_U312 , P1_R1165_U308 , P1_R1165_U189 );
nand NAND2_14615 ( P1_R1165_U313 , P1_U3155 , P1_R1165_U70 );
nand NAND3_14616 ( P1_R1165_U314 , P1_R1165_U312 , P1_R1165_U313 , P1_R1165_U185 );
nand NAND2_14617 ( P1_R1165_U315 , P1_R1165_U435 , P1_R1165_U34 );
nand NAND2_14618 ( P1_R1165_U316 , P1_R1165_U285 , P1_R1165_U175 );
not NOT1_14619 ( P1_R1165_U317 , P1_R1165_U55 );
nand NAND2_14620 ( P1_R1165_U318 , P1_R1165_U447 , P1_R1165_U50 );
nand NAND2_14621 ( P1_R1165_U319 , P1_R1165_U318 , P1_R1165_U55 );
nand NAND2_14622 ( P1_R1165_U320 , P1_R1165_U124 , P1_R1165_U319 );
nand NAND2_14623 ( P1_R1165_U321 , P1_R1165_U317 , P1_R1165_U188 );
nand NAND2_14624 ( P1_R1165_U322 , P1_U3160 , P1_R1165_U72 );
nand NAND3_14625 ( P1_R1165_U323 , P1_R1165_U322 , P1_R1165_U321 , P1_R1165_U8 );
nand NAND2_14626 ( P1_R1165_U324 , P1_R1165_U447 , P1_R1165_U50 );
nand NAND2_14627 ( P1_R1165_U325 , P1_R1165_U474 , P1_R1165_U37 );
nand NAND2_14628 ( P1_R1165_U326 , P1_R1165_U325 , P1_R1165_U56 );
nand NAND2_14629 ( P1_R1165_U327 , P1_R1165_U125 , P1_R1165_U326 );
nand NAND2_14630 ( P1_R1165_U328 , P1_R1165_U267 , P1_R1165_U38 );
nand NAND2_14631 ( P1_R1165_U329 , P1_U3164 , P1_R1165_U74 );
nand NAND2_14632 ( P1_R1165_U330 , P1_R1165_U126 , P1_R1165_U328 );
nand NAND2_14633 ( P1_R1165_U331 , P1_R1165_U474 , P1_R1165_U37 );
nand NAND2_14634 ( P1_R1165_U332 , P1_R1165_U255 , P1_R1165_U182 );
not NOT1_14635 ( P1_R1165_U333 , P1_R1165_U57 );
nand NAND2_14636 ( P1_R1165_U334 , P1_R1165_U459 , P1_R1165_U41 );
nand NAND2_14637 ( P1_R1165_U335 , P1_R1165_U334 , P1_R1165_U57 );
nand NAND2_14638 ( P1_R1165_U336 , P1_R1165_U127 , P1_R1165_U335 );
nand NAND2_14639 ( P1_R1165_U337 , P1_R1165_U333 , P1_R1165_U187 );
nand NAND2_14640 ( P1_R1165_U338 , P1_U3168 , P1_R1165_U77 );
nand NAND2_14641 ( P1_R1165_U339 , P1_R1165_U128 , P1_R1165_U337 );
nand NAND2_14642 ( P1_R1165_U340 , P1_R1165_U459 , P1_R1165_U41 );
nand NAND2_14643 ( P1_R1165_U341 , P1_R1165_U234 , P1_R1165_U17 );
nand NAND2_14644 ( P1_R1165_U342 , P1_R1165_U241 , P1_R1165_U20 );
nand NAND2_14645 ( P1_R1165_U343 , P1_R1165_U315 , P1_R1165_U189 );
nand NAND2_14646 ( P1_R1165_U344 , P1_R1165_U301 , P1_R1165_U192 );
nand NAND2_14647 ( P1_R1165_U345 , P1_R1165_U324 , P1_R1165_U188 );
nand NAND2_14648 ( P1_R1165_U346 , P1_R1165_U285 , P1_R1165_U49 );
nand NAND2_14649 ( P1_R1165_U347 , P1_R1165_U331 , P1_R1165_U38 );
nand NAND2_14650 ( P1_R1165_U348 , P1_R1165_U340 , P1_R1165_U187 );
nand NAND2_14651 ( P1_R1165_U349 , P1_R1165_U255 , P1_R1165_U43 );
nand NAND3_14652 ( P1_R1165_U350 , P1_R1165_U351 , P1_R1165_U302 , P1_R1165_U119 );
nand NAND2_14653 ( P1_R1165_U351 , P1_R1165_U299 , P1_R1165_U185 );
nand NAND2_14654 ( P1_R1165_U352 , P1_R1165_U70 , P1_R1165_U298 );
nand NAND2_14655 ( P1_R1165_U353 , P1_U3155 , P1_R1165_U298 );
nand NAND3_14656 ( P1_R1165_U354 , P1_R1165_U299 , P1_R1165_U185 , P1_R1165_U306 );
nand NAND3_14657 ( P1_R1165_U355 , P1_R1165_U168 , P1_R1165_U185 , P1_R1165_U120 );
nand NAND2_14658 ( P1_R1165_U356 , P1_R1165_U300 , P1_R1165_U306 );
nand NAND2_14659 ( P1_R1165_U357 , P1_U3154 , P1_R1165_U68 );
nand NAND2_14660 ( P1_R1165_U358 , P1_U3211 , P1_R1165_U130 );
nand NAND2_14661 ( P1_R1165_U359 , P1_U3201 , P1_R1165_U15 );
not NOT1_14662 ( P1_R1165_U360 , P1_R1165_U58 );
nand NAND2_14663 ( P1_R1165_U361 , P1_R1165_U360 , P1_U3172 );
nand NAND2_14664 ( P1_R1165_U362 , P1_R1165_U58 , P1_R1165_U28 );
nand NAND2_14665 ( P1_R1165_U363 , P1_R1165_U360 , P1_U3172 );
nand NAND2_14666 ( P1_R1165_U364 , P1_R1165_U58 , P1_R1165_U28 );
nand NAND2_14667 ( P1_R1165_U365 , P1_R1165_U364 , P1_R1165_U363 );
nand NAND2_14668 ( P1_R1165_U366 , P1_U3211 , P1_R1165_U132 );
nand NAND2_14669 ( P1_R1165_U367 , P1_U3210 , P1_R1165_U15 );
not NOT1_14670 ( P1_R1165_U368 , P1_R1165_U63 );
nand NAND2_14671 ( P1_R1165_U369 , P1_U3211 , P1_R1165_U133 );
nand NAND2_14672 ( P1_R1165_U370 , P1_U3209 , P1_R1165_U15 );
not NOT1_14673 ( P1_R1165_U371 , P1_R1165_U64 );
nand NAND2_14674 ( P1_R1165_U372 , P1_U3211 , P1_R1165_U134 );
nand NAND2_14675 ( P1_R1165_U373 , P1_U3207 , P1_R1165_U15 );
not NOT1_14676 ( P1_R1165_U374 , P1_R1165_U62 );
nand NAND2_14677 ( P1_R1165_U375 , P1_U3211 , P1_R1165_U135 );
nand NAND2_14678 ( P1_R1165_U376 , P1_U3208 , P1_R1165_U15 );
not NOT1_14679 ( P1_R1165_U377 , P1_R1165_U61 );
nand NAND2_14680 ( P1_R1165_U378 , P1_U3211 , P1_R1165_U136 );
nand NAND2_14681 ( P1_R1165_U379 , P1_U3206 , P1_R1165_U15 );
not NOT1_14682 ( P1_R1165_U380 , P1_R1165_U65 );
nand NAND2_14683 ( P1_R1165_U381 , P1_U3211 , P1_R1165_U137 );
nand NAND2_14684 ( P1_R1165_U382 , P1_U3205 , P1_R1165_U15 );
not NOT1_14685 ( P1_R1165_U383 , P1_R1165_U66 );
nand NAND2_14686 ( P1_R1165_U384 , P1_U3211 , P1_R1165_U138 );
nand NAND2_14687 ( P1_R1165_U385 , P1_U3203 , P1_R1165_U15 );
not NOT1_14688 ( P1_R1165_U386 , P1_R1165_U60 );
nand NAND2_14689 ( P1_R1165_U387 , P1_U3211 , P1_R1165_U139 );
nand NAND2_14690 ( P1_R1165_U388 , P1_U3204 , P1_R1165_U15 );
not NOT1_14691 ( P1_R1165_U389 , P1_R1165_U59 );
nand NAND2_14692 ( P1_R1165_U390 , P1_U3211 , P1_R1165_U140 );
nand NAND2_14693 ( P1_R1165_U391 , P1_U3202 , P1_R1165_U15 );
not NOT1_14694 ( P1_R1165_U392 , P1_R1165_U67 );
nand NAND2_14695 ( P1_R1165_U393 , P1_R1165_U131 , P1_R1165_U29 );
nand NAND2_14696 ( P1_R1165_U394 , P1_R1165_U365 , P1_R1165_U227 );
nand NAND2_14697 ( P1_R1165_U395 , P1_R1165_U392 , P1_U3173 );
nand NAND2_14698 ( P1_R1165_U396 , P1_R1165_U67 , P1_R1165_U27 );
nand NAND2_14699 ( P1_R1165_U397 , P1_R1165_U392 , P1_U3173 );
nand NAND2_14700 ( P1_R1165_U398 , P1_R1165_U67 , P1_R1165_U27 );
nand NAND2_14701 ( P1_R1165_U399 , P1_R1165_U398 , P1_R1165_U397 );
nand NAND2_14702 ( P1_R1165_U400 , P1_R1165_U141 , P1_R1165_U142 );
nand NAND2_14703 ( P1_R1165_U401 , P1_R1165_U223 , P1_R1165_U399 );
nand NAND2_14704 ( P1_R1165_U402 , P1_R1165_U386 , P1_U3174 );
nand NAND2_14705 ( P1_R1165_U403 , P1_R1165_U60 , P1_R1165_U18 );
nand NAND2_14706 ( P1_R1165_U404 , P1_R1165_U389 , P1_U3175 );
nand NAND2_14707 ( P1_R1165_U405 , P1_R1165_U59 , P1_R1165_U16 );
nand NAND2_14708 ( P1_R1165_U406 , P1_R1165_U405 , P1_R1165_U404 );
nand NAND2_14709 ( P1_R1165_U407 , P1_R1165_U341 , P1_R1165_U30 );
nand NAND2_14710 ( P1_R1165_U408 , P1_R1165_U406 , P1_R1165_U215 );
nand NAND2_14711 ( P1_R1165_U409 , P1_R1165_U383 , P1_U3176 );
nand NAND2_14712 ( P1_R1165_U410 , P1_R1165_U66 , P1_R1165_U26 );
nand NAND2_14713 ( P1_R1165_U411 , P1_R1165_U383 , P1_U3176 );
nand NAND2_14714 ( P1_R1165_U412 , P1_R1165_U66 , P1_R1165_U26 );
nand NAND2_14715 ( P1_R1165_U413 , P1_R1165_U412 , P1_R1165_U411 );
nand NAND2_14716 ( P1_R1165_U414 , P1_R1165_U143 , P1_R1165_U144 );
nand NAND2_14717 ( P1_R1165_U415 , P1_R1165_U211 , P1_R1165_U413 );
nand NAND2_14718 ( P1_R1165_U416 , P1_R1165_U380 , P1_U3177 );
nand NAND2_14719 ( P1_R1165_U417 , P1_R1165_U65 , P1_R1165_U25 );
nand NAND2_14720 ( P1_R1165_U418 , P1_R1165_U380 , P1_U3177 );
nand NAND2_14721 ( P1_R1165_U419 , P1_R1165_U65 , P1_R1165_U25 );
nand NAND2_14722 ( P1_R1165_U420 , P1_R1165_U419 , P1_R1165_U418 );
nand NAND2_14723 ( P1_R1165_U421 , P1_R1165_U145 , P1_R1165_U24 );
nand NAND2_14724 ( P1_R1165_U422 , P1_R1165_U420 , P1_R1165_U207 );
nand NAND2_14725 ( P1_R1165_U423 , P1_R1165_U374 , P1_U3178 );
nand NAND2_14726 ( P1_R1165_U424 , P1_R1165_U62 , P1_R1165_U21 );
nand NAND2_14727 ( P1_R1165_U425 , P1_R1165_U377 , P1_U3179 );
nand NAND2_14728 ( P1_R1165_U426 , P1_R1165_U61 , P1_R1165_U19 );
nand NAND2_14729 ( P1_R1165_U427 , P1_R1165_U426 , P1_R1165_U425 );
nand NAND2_14730 ( P1_R1165_U428 , P1_R1165_U342 , P1_R1165_U31 );
nand NAND2_14731 ( P1_R1165_U429 , P1_R1165_U427 , P1_R1165_U200 );
nand NAND2_14732 ( P1_R1165_U430 , P1_U3211 , P1_R1165_U146 );
nand NAND2_14733 ( P1_R1165_U431 , P1_U3183 , P1_R1165_U15 );
not NOT1_14734 ( P1_R1165_U432 , P1_R1165_U68 );
nand NAND2_14735 ( P1_R1165_U433 , P1_U3211 , P1_R1165_U147 );
nand NAND2_14736 ( P1_R1165_U434 , P1_U3185 , P1_R1165_U15 );
not NOT1_14737 ( P1_R1165_U435 , P1_R1165_U69 );
nand NAND2_14738 ( P1_R1165_U436 , P1_U3211 , P1_R1165_U148 );
nand NAND2_14739 ( P1_R1165_U437 , P1_U3184 , P1_R1165_U15 );
not NOT1_14740 ( P1_R1165_U438 , P1_R1165_U70 );
nand NAND2_14741 ( P1_R1165_U439 , P1_U3211 , P1_R1165_U149 );
nand NAND2_14742 ( P1_R1165_U440 , P1_U3186 , P1_R1165_U15 );
not NOT1_14743 ( P1_R1165_U441 , P1_R1165_U71 );
nand NAND2_14744 ( P1_R1165_U442 , P1_U3211 , P1_R1165_U150 );
nand NAND2_14745 ( P1_R1165_U443 , P1_U3189 , P1_R1165_U15 );
not NOT1_14746 ( P1_R1165_U444 , P1_R1165_U72 );
nand NAND2_14747 ( P1_R1165_U445 , P1_U3211 , P1_R1165_U151 );
nand NAND2_14748 ( P1_R1165_U446 , P1_U3190 , P1_R1165_U15 );
not NOT1_14749 ( P1_R1165_U447 , P1_R1165_U83 );
nand NAND2_14750 ( P1_R1165_U448 , P1_U3211 , P1_R1165_U152 );
nand NAND2_14751 ( P1_R1165_U449 , P1_U3191 , P1_R1165_U15 );
not NOT1_14752 ( P1_R1165_U450 , P1_R1165_U82 );
nand NAND2_14753 ( P1_R1165_U451 , P1_U3211 , P1_R1165_U153 );
nand NAND2_14754 ( P1_R1165_U452 , P1_U3200 , P1_R1165_U15 );
not NOT1_14755 ( P1_R1165_U453 , P1_R1165_U75 );
nand NAND2_14756 ( P1_R1165_U454 , P1_U3211 , P1_R1165_U154 );
nand NAND2_14757 ( P1_R1165_U455 , P1_U3197 , P1_R1165_U15 );
not NOT1_14758 ( P1_R1165_U456 , P1_R1165_U77 );
nand NAND2_14759 ( P1_R1165_U457 , P1_U3211 , P1_R1165_U155 );
nand NAND2_14760 ( P1_R1165_U458 , P1_U3198 , P1_R1165_U15 );
not NOT1_14761 ( P1_R1165_U459 , P1_R1165_U78 );
nand NAND2_14762 ( P1_R1165_U460 , P1_U3211 , P1_R1165_U156 );
nand NAND2_14763 ( P1_R1165_U461 , P1_U3199 , P1_R1165_U15 );
not NOT1_14764 ( P1_R1165_U462 , P1_R1165_U76 );
nand NAND2_14765 ( P1_R1165_U463 , P1_U3211 , P1_R1165_U157 );
nand NAND2_14766 ( P1_R1165_U464 , P1_U3196 , P1_R1165_U15 );
not NOT1_14767 ( P1_R1165_U465 , P1_R1165_U79 );
nand NAND2_14768 ( P1_R1165_U466 , P1_U3211 , P1_R1165_U158 );
nand NAND2_14769 ( P1_R1165_U467 , P1_U3195 , P1_R1165_U15 );
not NOT1_14770 ( P1_R1165_U468 , P1_R1165_U80 );
nand NAND2_14771 ( P1_R1165_U469 , P1_U3211 , P1_R1165_U159 );
nand NAND2_14772 ( P1_R1165_U470 , P1_U3193 , P1_R1165_U15 );
not NOT1_14773 ( P1_R1165_U471 , P1_R1165_U74 );
nand NAND2_14774 ( P1_R1165_U472 , P1_U3211 , P1_R1165_U160 );
nand NAND2_14775 ( P1_R1165_U473 , P1_U3194 , P1_R1165_U15 );
not NOT1_14776 ( P1_R1165_U474 , P1_R1165_U73 );
nand NAND2_14777 ( P1_R1165_U475 , P1_U3211 , P1_R1165_U161 );
nand NAND2_14778 ( P1_R1165_U476 , P1_U3192 , P1_R1165_U15 );
not NOT1_14779 ( P1_R1165_U477 , P1_R1165_U81 );
nand NAND2_14780 ( P1_R1165_U478 , P1_U3211 , P1_R1165_U162 );
nand NAND2_14781 ( P1_R1165_U479 , P1_U3188 , P1_R1165_U15 );
not NOT1_14782 ( P1_R1165_U480 , P1_R1165_U84 );
nand NAND2_14783 ( P1_R1165_U481 , P1_U3211 , P1_R1165_U163 );
nand NAND2_14784 ( P1_R1165_U482 , P1_U3187 , P1_R1165_U15 );
not NOT1_14785 ( P1_R1165_U483 , P1_R1165_U85 );
nand NAND2_14786 ( P1_R1165_U484 , P1_U3211 , P1_R1165_U164 );
nand NAND2_14787 ( P1_R1165_U485 , P1_U3153 , P1_R1165_U15 );
not NOT1_14788 ( P1_R1165_U486 , P1_R1165_U122 );
nand NAND2_14789 ( P1_R1165_U487 , P1_U3182 , P1_R1165_U486 );
nand NAND2_14790 ( P1_R1165_U488 , P1_R1165_U122 , P1_R1165_U165 );
not NOT1_14791 ( P1_R1165_U489 , P1_R1165_U86 );
nand NAND3_14792 ( P1_R1165_U490 , P1_R1165_U350 , P1_R1165_U304 , P1_R1165_U489 );
nand NAND4_14793 ( P1_R1165_U491 , P1_R1165_U356 , P1_R1165_U355 , P1_R1165_U121 , P1_R1165_U86 );
nand NAND2_14794 ( P1_R1165_U492 , P1_R1165_U432 , P1_U3154 );
nand NAND2_14795 ( P1_R1165_U493 , P1_R1165_U68 , P1_R1165_U32 );
nand NAND2_14796 ( P1_R1165_U494 , P1_R1165_U432 , P1_U3154 );
nand NAND2_14797 ( P1_R1165_U495 , P1_R1165_U68 , P1_R1165_U32 );
nand NAND2_14798 ( P1_R1165_U496 , P1_R1165_U495 , P1_R1165_U494 );
nand NAND2_14799 ( P1_R1165_U497 , P1_R1165_U166 , P1_R1165_U167 );
nand NAND2_14800 ( P1_R1165_U498 , P1_R1165_U303 , P1_R1165_U496 );
nand NAND2_14801 ( P1_R1165_U499 , P1_R1165_U438 , P1_U3155 );
nand NAND2_14802 ( P1_R1165_U500 , P1_R1165_U70 , P1_R1165_U33 );
nand NAND2_14803 ( P1_R1165_U501 , P1_R1165_U435 , P1_U3156 );
nand NAND2_14804 ( P1_R1165_U502 , P1_R1165_U69 , P1_R1165_U34 );
nand NAND2_14805 ( P1_R1165_U503 , P1_R1165_U502 , P1_R1165_U501 );
nand NAND2_14806 ( P1_R1165_U504 , P1_R1165_U343 , P1_R1165_U54 );
nand NAND2_14807 ( P1_R1165_U505 , P1_R1165_U503 , P1_R1165_U308 );
nand NAND2_14808 ( P1_R1165_U506 , P1_R1165_U441 , P1_U3157 );
nand NAND2_14809 ( P1_R1165_U507 , P1_R1165_U71 , P1_R1165_U35 );
nand NAND2_14810 ( P1_R1165_U508 , P1_R1165_U507 , P1_R1165_U506 );
nand NAND2_14811 ( P1_R1165_U509 , P1_R1165_U344 , P1_R1165_U168 );
nand NAND2_14812 ( P1_R1165_U510 , P1_R1165_U297 , P1_R1165_U508 );
nand NAND2_14813 ( P1_R1165_U511 , P1_R1165_U483 , P1_U3158 );
nand NAND2_14814 ( P1_R1165_U512 , P1_R1165_U85 , P1_R1165_U52 );
nand NAND2_14815 ( P1_R1165_U513 , P1_R1165_U483 , P1_U3158 );
nand NAND2_14816 ( P1_R1165_U514 , P1_R1165_U85 , P1_R1165_U52 );
nand NAND2_14817 ( P1_R1165_U515 , P1_R1165_U514 , P1_R1165_U513 );
nand NAND2_14818 ( P1_R1165_U516 , P1_R1165_U169 , P1_R1165_U170 );
nand NAND2_14819 ( P1_R1165_U517 , P1_R1165_U293 , P1_R1165_U515 );
nand NAND2_14820 ( P1_R1165_U518 , P1_R1165_U480 , P1_U3159 );
nand NAND2_14821 ( P1_R1165_U519 , P1_R1165_U84 , P1_R1165_U51 );
nand NAND2_14822 ( P1_R1165_U520 , P1_R1165_U480 , P1_U3159 );
nand NAND2_14823 ( P1_R1165_U521 , P1_R1165_U84 , P1_R1165_U51 );
nand NAND2_14824 ( P1_R1165_U522 , P1_R1165_U521 , P1_R1165_U520 );
nand NAND2_14825 ( P1_R1165_U523 , P1_R1165_U171 , P1_R1165_U172 );
nand NAND2_14826 ( P1_R1165_U524 , P1_R1165_U289 , P1_R1165_U522 );
nand NAND2_14827 ( P1_R1165_U525 , P1_R1165_U444 , P1_U3160 );
nand NAND2_14828 ( P1_R1165_U526 , P1_R1165_U72 , P1_R1165_U36 );
nand NAND2_14829 ( P1_R1165_U527 , P1_R1165_U447 , P1_U3161 );
nand NAND2_14830 ( P1_R1165_U528 , P1_R1165_U83 , P1_R1165_U50 );
nand NAND2_14831 ( P1_R1165_U529 , P1_R1165_U528 , P1_R1165_U527 );
nand NAND2_14832 ( P1_R1165_U530 , P1_R1165_U345 , P1_R1165_U55 );
nand NAND2_14833 ( P1_R1165_U531 , P1_R1165_U529 , P1_R1165_U317 );
nand NAND2_14834 ( P1_R1165_U532 , P1_R1165_U371 , P1_U3180 );
nand NAND2_14835 ( P1_R1165_U533 , P1_R1165_U64 , P1_R1165_U23 );
nand NAND2_14836 ( P1_R1165_U534 , P1_R1165_U371 , P1_U3180 );
nand NAND2_14837 ( P1_R1165_U535 , P1_R1165_U64 , P1_R1165_U23 );
nand NAND2_14838 ( P1_R1165_U536 , P1_R1165_U535 , P1_R1165_U534 );
nand NAND2_14839 ( P1_R1165_U537 , P1_R1165_U173 , P1_R1165_U174 );
nand NAND2_14840 ( P1_R1165_U538 , P1_R1165_U196 , P1_R1165_U536 );
nand NAND2_14841 ( P1_R1165_U539 , P1_R1165_U450 , P1_U3162 );
nand NAND2_14842 ( P1_R1165_U540 , P1_R1165_U82 , P1_R1165_U48 );
nand NAND2_14843 ( P1_R1165_U541 , P1_R1165_U540 , P1_R1165_U539 );
nand NAND2_14844 ( P1_R1165_U542 , P1_R1165_U346 , P1_R1165_U175 );
nand NAND2_14845 ( P1_R1165_U543 , P1_R1165_U279 , P1_R1165_U541 );
nand NAND2_14846 ( P1_R1165_U544 , P1_R1165_U477 , P1_U3163 );
nand NAND2_14847 ( P1_R1165_U545 , P1_R1165_U81 , P1_R1165_U47 );
nand NAND2_14848 ( P1_R1165_U546 , P1_R1165_U477 , P1_U3163 );
nand NAND2_14849 ( P1_R1165_U547 , P1_R1165_U81 , P1_R1165_U47 );
nand NAND2_14850 ( P1_R1165_U548 , P1_R1165_U547 , P1_R1165_U546 );
nand NAND2_14851 ( P1_R1165_U549 , P1_R1165_U176 , P1_R1165_U177 );
nand NAND2_14852 ( P1_R1165_U550 , P1_R1165_U275 , P1_R1165_U548 );
nand NAND2_14853 ( P1_R1165_U551 , P1_R1165_U471 , P1_U3164 );
nand NAND2_14854 ( P1_R1165_U552 , P1_R1165_U74 , P1_R1165_U39 );
nand NAND2_14855 ( P1_R1165_U553 , P1_R1165_U474 , P1_U3165 );
nand NAND2_14856 ( P1_R1165_U554 , P1_R1165_U73 , P1_R1165_U37 );
nand NAND2_14857 ( P1_R1165_U555 , P1_R1165_U554 , P1_R1165_U553 );
nand NAND2_14858 ( P1_R1165_U556 , P1_R1165_U347 , P1_R1165_U56 );
nand NAND2_14859 ( P1_R1165_U557 , P1_R1165_U555 , P1_R1165_U267 );
nand NAND2_14860 ( P1_R1165_U558 , P1_R1165_U468 , P1_U3166 );
nand NAND2_14861 ( P1_R1165_U559 , P1_R1165_U80 , P1_R1165_U46 );
nand NAND2_14862 ( P1_R1165_U560 , P1_R1165_U468 , P1_U3166 );
nand NAND2_14863 ( P1_R1165_U561 , P1_R1165_U80 , P1_R1165_U46 );
nand NAND2_14864 ( P1_R1165_U562 , P1_R1165_U561 , P1_R1165_U560 );
nand NAND2_14865 ( P1_R1165_U563 , P1_R1165_U178 , P1_R1165_U179 );
nand NAND2_14866 ( P1_R1165_U564 , P1_R1165_U263 , P1_R1165_U562 );
nand NAND2_14867 ( P1_R1165_U565 , P1_R1165_U465 , P1_U3167 );
nand NAND2_14868 ( P1_R1165_U566 , P1_R1165_U79 , P1_R1165_U45 );
nand NAND2_14869 ( P1_R1165_U567 , P1_R1165_U465 , P1_U3167 );
nand NAND2_14870 ( P1_R1165_U568 , P1_R1165_U79 , P1_R1165_U45 );
nand NAND2_14871 ( P1_R1165_U569 , P1_R1165_U568 , P1_R1165_U567 );
nand NAND2_14872 ( P1_R1165_U570 , P1_R1165_U180 , P1_R1165_U181 );
nand NAND2_14873 ( P1_R1165_U571 , P1_R1165_U259 , P1_R1165_U569 );
nand NAND2_14874 ( P1_R1165_U572 , P1_R1165_U456 , P1_U3168 );
nand NAND2_14875 ( P1_R1165_U573 , P1_R1165_U77 , P1_R1165_U44 );
nand NAND2_14876 ( P1_R1165_U574 , P1_R1165_U459 , P1_U3169 );
nand NAND2_14877 ( P1_R1165_U575 , P1_R1165_U78 , P1_R1165_U41 );
nand NAND2_14878 ( P1_R1165_U576 , P1_R1165_U575 , P1_R1165_U574 );
nand NAND2_14879 ( P1_R1165_U577 , P1_R1165_U348 , P1_R1165_U57 );
nand NAND2_14880 ( P1_R1165_U578 , P1_R1165_U576 , P1_R1165_U333 );
nand NAND2_14881 ( P1_R1165_U579 , P1_R1165_U462 , P1_U3170 );
nand NAND2_14882 ( P1_R1165_U580 , P1_R1165_U76 , P1_R1165_U42 );
nand NAND2_14883 ( P1_R1165_U581 , P1_R1165_U580 , P1_R1165_U579 );
nand NAND2_14884 ( P1_R1165_U582 , P1_R1165_U349 , P1_R1165_U182 );
nand NAND2_14885 ( P1_R1165_U583 , P1_R1165_U249 , P1_R1165_U581 );
nand NAND2_14886 ( P1_R1165_U584 , P1_R1165_U453 , P1_U3171 );
nand NAND2_14887 ( P1_R1165_U585 , P1_R1165_U75 , P1_R1165_U40 );
nand NAND2_14888 ( P1_R1165_U586 , P1_R1165_U453 , P1_U3171 );
nand NAND2_14889 ( P1_R1165_U587 , P1_R1165_U75 , P1_R1165_U40 );
nand NAND2_14890 ( P1_R1165_U588 , P1_R1165_U587 , P1_R1165_U586 );
nand NAND2_14891 ( P1_R1165_U589 , P1_R1165_U183 , P1_R1165_U184 );
nand NAND2_14892 ( P1_R1165_U590 , P1_R1165_U245 , P1_R1165_U588 );
nand NAND2_14893 ( P1_R1165_U591 , P1_U3181 , P1_R1165_U15 );
nand NAND2_14894 ( P1_R1165_U592 , P1_U3211 , P1_R1165_U22 );
not NOT1_14895 ( P1_R1165_U593 , P1_R1165_U129 );
nand NAND2_14896 ( P1_R1165_U594 , P1_R1165_U63 , P1_R1165_U593 );
nand NAND2_14897 ( P1_R1165_U595 , P1_R1165_U129 , P1_R1165_U368 );
and AND2_14898 ( P1_R1150_U6 , P1_R1150_U184 , P1_R1150_U201 );
and AND2_14899 ( P1_R1150_U7 , P1_R1150_U203 , P1_R1150_U202 );
and AND2_14900 ( P1_R1150_U8 , P1_R1150_U179 , P1_R1150_U240 );
and AND2_14901 ( P1_R1150_U9 , P1_R1150_U242 , P1_R1150_U241 );
and AND2_14902 ( P1_R1150_U10 , P1_R1150_U259 , P1_R1150_U258 );
and AND2_14903 ( P1_R1150_U11 , P1_R1150_U285 , P1_R1150_U284 );
and AND2_14904 ( P1_R1150_U12 , P1_R1150_U383 , P1_R1150_U382 );
nand NAND2_14905 ( P1_R1150_U13 , P1_R1150_U340 , P1_R1150_U343 );
nand NAND2_14906 ( P1_R1150_U14 , P1_R1150_U329 , P1_R1150_U332 );
nand NAND2_14907 ( P1_R1150_U15 , P1_R1150_U318 , P1_R1150_U321 );
nand NAND2_14908 ( P1_R1150_U16 , P1_R1150_U310 , P1_R1150_U312 );
nand NAND3_14909 ( P1_R1150_U17 , P1_R1150_U156 , P1_R1150_U175 , P1_R1150_U348 );
nand NAND2_14910 ( P1_R1150_U18 , P1_R1150_U236 , P1_R1150_U238 );
nand NAND2_14911 ( P1_R1150_U19 , P1_R1150_U228 , P1_R1150_U231 );
nand NAND2_14912 ( P1_R1150_U20 , P1_R1150_U220 , P1_R1150_U222 );
nand NAND2_14913 ( P1_R1150_U21 , P1_R1150_U25 , P1_R1150_U346 );
not NOT1_14914 ( P1_R1150_U22 , P1_U3479 );
not NOT1_14915 ( P1_R1150_U23 , P1_U3464 );
not NOT1_14916 ( P1_R1150_U24 , P1_U3456 );
nand NAND2_14917 ( P1_R1150_U25 , P1_U3456 , P1_R1150_U93 );
not NOT1_14918 ( P1_R1150_U26 , P1_U3078 );
not NOT1_14919 ( P1_R1150_U27 , P1_U3467 );
not NOT1_14920 ( P1_R1150_U28 , P1_U3068 );
nand NAND2_14921 ( P1_R1150_U29 , P1_U3068 , P1_R1150_U23 );
not NOT1_14922 ( P1_R1150_U30 , P1_U3064 );
not NOT1_14923 ( P1_R1150_U31 , P1_U3476 );
not NOT1_14924 ( P1_R1150_U32 , P1_U3473 );
not NOT1_14925 ( P1_R1150_U33 , P1_U3470 );
not NOT1_14926 ( P1_R1150_U34 , P1_U3071 );
not NOT1_14927 ( P1_R1150_U35 , P1_U3067 );
not NOT1_14928 ( P1_R1150_U36 , P1_U3060 );
nand NAND2_14929 ( P1_R1150_U37 , P1_U3060 , P1_R1150_U33 );
not NOT1_14930 ( P1_R1150_U38 , P1_U3482 );
not NOT1_14931 ( P1_R1150_U39 , P1_U3070 );
nand NAND2_14932 ( P1_R1150_U40 , P1_U3070 , P1_R1150_U22 );
not NOT1_14933 ( P1_R1150_U41 , P1_U3084 );
not NOT1_14934 ( P1_R1150_U42 , P1_U3485 );
not NOT1_14935 ( P1_R1150_U43 , P1_U3083 );
nand NAND2_14936 ( P1_R1150_U44 , P1_R1150_U209 , P1_R1150_U208 );
nand NAND2_14937 ( P1_R1150_U45 , P1_R1150_U37 , P1_R1150_U224 );
nand NAND2_14938 ( P1_R1150_U46 , P1_R1150_U193 , P1_R1150_U192 );
not NOT1_14939 ( P1_R1150_U47 , P1_U4019 );
not NOT1_14940 ( P1_R1150_U48 , P1_U4023 );
not NOT1_14941 ( P1_R1150_U49 , P1_U3503 );
not NOT1_14942 ( P1_R1150_U50 , P1_U3491 );
not NOT1_14943 ( P1_R1150_U51 , P1_U3488 );
not NOT1_14944 ( P1_R1150_U52 , P1_U3063 );
not NOT1_14945 ( P1_R1150_U53 , P1_U3062 );
nand NAND2_14946 ( P1_R1150_U54 , P1_U3083 , P1_R1150_U42 );
not NOT1_14947 ( P1_R1150_U55 , P1_U3494 );
not NOT1_14948 ( P1_R1150_U56 , P1_U3072 );
not NOT1_14949 ( P1_R1150_U57 , P1_U3497 );
not NOT1_14950 ( P1_R1150_U58 , P1_U3080 );
not NOT1_14951 ( P1_R1150_U59 , P1_U3506 );
not NOT1_14952 ( P1_R1150_U60 , P1_U3500 );
not NOT1_14953 ( P1_R1150_U61 , P1_U3073 );
not NOT1_14954 ( P1_R1150_U62 , P1_U3074 );
not NOT1_14955 ( P1_R1150_U63 , P1_U3079 );
nand NAND2_14956 ( P1_R1150_U64 , P1_U3079 , P1_R1150_U60 );
not NOT1_14957 ( P1_R1150_U65 , P1_U3509 );
not NOT1_14958 ( P1_R1150_U66 , P1_U3069 );
nand NAND2_14959 ( P1_R1150_U67 , P1_R1150_U269 , P1_R1150_U268 );
not NOT1_14960 ( P1_R1150_U68 , P1_U3082 );
not NOT1_14961 ( P1_R1150_U69 , P1_U3514 );
not NOT1_14962 ( P1_R1150_U70 , P1_U3081 );
not NOT1_14963 ( P1_R1150_U71 , P1_U4025 );
not NOT1_14964 ( P1_R1150_U72 , P1_U3076 );
not NOT1_14965 ( P1_R1150_U73 , P1_U4022 );
not NOT1_14966 ( P1_R1150_U74 , P1_U4024 );
not NOT1_14967 ( P1_R1150_U75 , P1_U3066 );
not NOT1_14968 ( P1_R1150_U76 , P1_U3061 );
not NOT1_14969 ( P1_R1150_U77 , P1_U3075 );
nand NAND2_14970 ( P1_R1150_U78 , P1_U3075 , P1_R1150_U74 );
not NOT1_14971 ( P1_R1150_U79 , P1_U4021 );
not NOT1_14972 ( P1_R1150_U80 , P1_U3065 );
not NOT1_14973 ( P1_R1150_U81 , P1_U4020 );
not NOT1_14974 ( P1_R1150_U82 , P1_U3058 );
not NOT1_14975 ( P1_R1150_U83 , P1_U4018 );
not NOT1_14976 ( P1_R1150_U84 , P1_U3057 );
nand NAND2_14977 ( P1_R1150_U85 , P1_U3057 , P1_R1150_U47 );
not NOT1_14978 ( P1_R1150_U86 , P1_U3053 );
not NOT1_14979 ( P1_R1150_U87 , P1_U4017 );
not NOT1_14980 ( P1_R1150_U88 , P1_U3054 );
nand NAND2_14981 ( P1_R1150_U89 , P1_R1150_U299 , P1_R1150_U298 );
nand NAND2_14982 ( P1_R1150_U90 , P1_R1150_U78 , P1_R1150_U314 );
nand NAND2_14983 ( P1_R1150_U91 , P1_R1150_U64 , P1_R1150_U325 );
nand NAND2_14984 ( P1_R1150_U92 , P1_R1150_U54 , P1_R1150_U336 );
not NOT1_14985 ( P1_R1150_U93 , P1_U3077 );
nand NAND2_14986 ( P1_R1150_U94 , P1_R1150_U393 , P1_R1150_U392 );
nand NAND2_14987 ( P1_R1150_U95 , P1_R1150_U407 , P1_R1150_U406 );
nand NAND2_14988 ( P1_R1150_U96 , P1_R1150_U412 , P1_R1150_U411 );
nand NAND2_14989 ( P1_R1150_U97 , P1_R1150_U428 , P1_R1150_U427 );
nand NAND2_14990 ( P1_R1150_U98 , P1_R1150_U433 , P1_R1150_U432 );
nand NAND2_14991 ( P1_R1150_U99 , P1_R1150_U438 , P1_R1150_U437 );
nand NAND2_14992 ( P1_R1150_U100 , P1_R1150_U443 , P1_R1150_U442 );
nand NAND2_14993 ( P1_R1150_U101 , P1_R1150_U448 , P1_R1150_U447 );
nand NAND2_14994 ( P1_R1150_U102 , P1_R1150_U464 , P1_R1150_U463 );
nand NAND2_14995 ( P1_R1150_U103 , P1_R1150_U469 , P1_R1150_U468 );
nand NAND2_14996 ( P1_R1150_U104 , P1_R1150_U352 , P1_R1150_U351 );
nand NAND2_14997 ( P1_R1150_U105 , P1_R1150_U361 , P1_R1150_U360 );
nand NAND2_14998 ( P1_R1150_U106 , P1_R1150_U368 , P1_R1150_U367 );
nand NAND2_14999 ( P1_R1150_U107 , P1_R1150_U372 , P1_R1150_U371 );
nand NAND2_15000 ( P1_R1150_U108 , P1_R1150_U381 , P1_R1150_U380 );
nand NAND2_15001 ( P1_R1150_U109 , P1_R1150_U402 , P1_R1150_U401 );
nand NAND2_15002 ( P1_R1150_U110 , P1_R1150_U419 , P1_R1150_U418 );
nand NAND2_15003 ( P1_R1150_U111 , P1_R1150_U423 , P1_R1150_U422 );
nand NAND2_15004 ( P1_R1150_U112 , P1_R1150_U455 , P1_R1150_U454 );
nand NAND2_15005 ( P1_R1150_U113 , P1_R1150_U459 , P1_R1150_U458 );
nand NAND2_15006 ( P1_R1150_U114 , P1_R1150_U476 , P1_R1150_U475 );
and AND2_15007 ( P1_R1150_U115 , P1_R1150_U195 , P1_R1150_U183 );
and AND2_15008 ( P1_R1150_U116 , P1_R1150_U198 , P1_R1150_U199 );
and AND2_15009 ( P1_R1150_U117 , P1_R1150_U211 , P1_R1150_U185 );
and AND2_15010 ( P1_R1150_U118 , P1_R1150_U214 , P1_R1150_U215 );
and AND3_15011 ( P1_R1150_U119 , P1_R1150_U354 , P1_R1150_U353 , P1_R1150_U40 );
and AND2_15012 ( P1_R1150_U120 , P1_R1150_U357 , P1_R1150_U185 );
and AND2_15013 ( P1_R1150_U121 , P1_R1150_U230 , P1_R1150_U7 );
and AND2_15014 ( P1_R1150_U122 , P1_R1150_U364 , P1_R1150_U184 );
and AND3_15015 ( P1_R1150_U123 , P1_R1150_U374 , P1_R1150_U373 , P1_R1150_U29 );
and AND2_15016 ( P1_R1150_U124 , P1_R1150_U377 , P1_R1150_U183 );
and AND2_15017 ( P1_R1150_U125 , P1_R1150_U217 , P1_R1150_U8 );
and AND2_15018 ( P1_R1150_U126 , P1_R1150_U262 , P1_R1150_U180 );
and AND2_15019 ( P1_R1150_U127 , P1_R1150_U288 , P1_R1150_U181 );
and AND2_15020 ( P1_R1150_U128 , P1_R1150_U304 , P1_R1150_U305 );
and AND2_15021 ( P1_R1150_U129 , P1_R1150_U307 , P1_R1150_U386 );
and AND3_15022 ( P1_R1150_U130 , P1_R1150_U305 , P1_R1150_U304 , P1_R1150_U308 );
nand NAND2_15023 ( P1_R1150_U131 , P1_R1150_U390 , P1_R1150_U389 );
and AND3_15024 ( P1_R1150_U132 , P1_R1150_U395 , P1_R1150_U394 , P1_R1150_U85 );
and AND2_15025 ( P1_R1150_U133 , P1_R1150_U398 , P1_R1150_U182 );
nand NAND2_15026 ( P1_R1150_U134 , P1_R1150_U404 , P1_R1150_U403 );
nand NAND2_15027 ( P1_R1150_U135 , P1_R1150_U409 , P1_R1150_U408 );
and AND2_15028 ( P1_R1150_U136 , P1_R1150_U415 , P1_R1150_U181 );
nand NAND2_15029 ( P1_R1150_U137 , P1_R1150_U425 , P1_R1150_U424 );
nand NAND2_15030 ( P1_R1150_U138 , P1_R1150_U430 , P1_R1150_U429 );
nand NAND2_15031 ( P1_R1150_U139 , P1_R1150_U435 , P1_R1150_U434 );
nand NAND2_15032 ( P1_R1150_U140 , P1_R1150_U440 , P1_R1150_U439 );
nand NAND2_15033 ( P1_R1150_U141 , P1_R1150_U445 , P1_R1150_U444 );
and AND2_15034 ( P1_R1150_U142 , P1_R1150_U451 , P1_R1150_U180 );
nand NAND2_15035 ( P1_R1150_U143 , P1_R1150_U461 , P1_R1150_U460 );
nand NAND2_15036 ( P1_R1150_U144 , P1_R1150_U466 , P1_R1150_U465 );
and AND2_15037 ( P1_R1150_U145 , P1_R1150_U342 , P1_R1150_U9 );
and AND2_15038 ( P1_R1150_U146 , P1_R1150_U472 , P1_R1150_U179 );
and AND2_15039 ( P1_R1150_U147 , P1_R1150_U350 , P1_R1150_U349 );
nand NAND2_15040 ( P1_R1150_U148 , P1_R1150_U118 , P1_R1150_U212 );
and AND2_15041 ( P1_R1150_U149 , P1_R1150_U359 , P1_R1150_U358 );
and AND2_15042 ( P1_R1150_U150 , P1_R1150_U366 , P1_R1150_U365 );
and AND2_15043 ( P1_R1150_U151 , P1_R1150_U370 , P1_R1150_U369 );
nand NAND2_15044 ( P1_R1150_U152 , P1_R1150_U116 , P1_R1150_U196 );
and AND2_15045 ( P1_R1150_U153 , P1_R1150_U379 , P1_R1150_U378 );
not NOT1_15046 ( P1_R1150_U154 , P1_U4028 );
not NOT1_15047 ( P1_R1150_U155 , P1_U3055 );
and AND2_15048 ( P1_R1150_U156 , P1_R1150_U388 , P1_R1150_U387 );
nand NAND2_15049 ( P1_R1150_U157 , P1_R1150_U128 , P1_R1150_U302 );
and AND2_15050 ( P1_R1150_U158 , P1_R1150_U400 , P1_R1150_U399 );
nand NAND2_15051 ( P1_R1150_U159 , P1_R1150_U295 , P1_R1150_U294 );
nand NAND2_15052 ( P1_R1150_U160 , P1_R1150_U291 , P1_R1150_U290 );
and AND2_15053 ( P1_R1150_U161 , P1_R1150_U417 , P1_R1150_U416 );
and AND2_15054 ( P1_R1150_U162 , P1_R1150_U421 , P1_R1150_U420 );
nand NAND2_15055 ( P1_R1150_U163 , P1_R1150_U281 , P1_R1150_U280 );
nand NAND2_15056 ( P1_R1150_U164 , P1_R1150_U277 , P1_R1150_U276 );
not NOT1_15057 ( P1_R1150_U165 , P1_U3461 );
nand NAND2_15058 ( P1_R1150_U166 , P1_R1150_U273 , P1_R1150_U272 );
not NOT1_15059 ( P1_R1150_U167 , P1_U3512 );
nand NAND2_15060 ( P1_R1150_U168 , P1_R1150_U265 , P1_R1150_U264 );
and AND2_15061 ( P1_R1150_U169 , P1_R1150_U453 , P1_R1150_U452 );
and AND2_15062 ( P1_R1150_U170 , P1_R1150_U457 , P1_R1150_U456 );
nand NAND2_15063 ( P1_R1150_U171 , P1_R1150_U255 , P1_R1150_U254 );
nand NAND2_15064 ( P1_R1150_U172 , P1_R1150_U251 , P1_R1150_U250 );
nand NAND2_15065 ( P1_R1150_U173 , P1_R1150_U247 , P1_R1150_U246 );
and AND2_15066 ( P1_R1150_U174 , P1_R1150_U474 , P1_R1150_U473 );
nand NAND2_15067 ( P1_R1150_U175 , P1_R1150_U129 , P1_R1150_U157 );
not NOT1_15068 ( P1_R1150_U176 , P1_R1150_U85 );
not NOT1_15069 ( P1_R1150_U177 , P1_R1150_U29 );
not NOT1_15070 ( P1_R1150_U178 , P1_R1150_U40 );
nand NAND2_15071 ( P1_R1150_U179 , P1_U3488 , P1_R1150_U53 );
nand NAND2_15072 ( P1_R1150_U180 , P1_U3503 , P1_R1150_U62 );
nand NAND2_15073 ( P1_R1150_U181 , P1_U4023 , P1_R1150_U76 );
nand NAND2_15074 ( P1_R1150_U182 , P1_U4019 , P1_R1150_U84 );
nand NAND2_15075 ( P1_R1150_U183 , P1_U3464 , P1_R1150_U28 );
nand NAND2_15076 ( P1_R1150_U184 , P1_U3473 , P1_R1150_U35 );
nand NAND2_15077 ( P1_R1150_U185 , P1_U3479 , P1_R1150_U39 );
not NOT1_15078 ( P1_R1150_U186 , P1_R1150_U64 );
not NOT1_15079 ( P1_R1150_U187 , P1_R1150_U78 );
not NOT1_15080 ( P1_R1150_U188 , P1_R1150_U37 );
not NOT1_15081 ( P1_R1150_U189 , P1_R1150_U54 );
not NOT1_15082 ( P1_R1150_U190 , P1_R1150_U25 );
nand NAND2_15083 ( P1_R1150_U191 , P1_R1150_U190 , P1_R1150_U26 );
nand NAND2_15084 ( P1_R1150_U192 , P1_R1150_U191 , P1_R1150_U165 );
nand NAND2_15085 ( P1_R1150_U193 , P1_U3078 , P1_R1150_U25 );
not NOT1_15086 ( P1_R1150_U194 , P1_R1150_U46 );
nand NAND2_15087 ( P1_R1150_U195 , P1_U3467 , P1_R1150_U30 );
nand NAND2_15088 ( P1_R1150_U196 , P1_R1150_U115 , P1_R1150_U46 );
nand NAND2_15089 ( P1_R1150_U197 , P1_R1150_U30 , P1_R1150_U29 );
nand NAND2_15090 ( P1_R1150_U198 , P1_R1150_U197 , P1_R1150_U27 );
nand NAND2_15091 ( P1_R1150_U199 , P1_U3064 , P1_R1150_U177 );
not NOT1_15092 ( P1_R1150_U200 , P1_R1150_U152 );
nand NAND2_15093 ( P1_R1150_U201 , P1_U3476 , P1_R1150_U34 );
nand NAND2_15094 ( P1_R1150_U202 , P1_U3071 , P1_R1150_U31 );
nand NAND2_15095 ( P1_R1150_U203 , P1_U3067 , P1_R1150_U32 );
nand NAND2_15096 ( P1_R1150_U204 , P1_R1150_U188 , P1_R1150_U6 );
nand NAND2_15097 ( P1_R1150_U205 , P1_R1150_U7 , P1_R1150_U204 );
nand NAND2_15098 ( P1_R1150_U206 , P1_U3470 , P1_R1150_U36 );
nand NAND2_15099 ( P1_R1150_U207 , P1_U3476 , P1_R1150_U34 );
nand NAND3_15100 ( P1_R1150_U208 , P1_R1150_U206 , P1_R1150_U152 , P1_R1150_U6 );
nand NAND2_15101 ( P1_R1150_U209 , P1_R1150_U207 , P1_R1150_U205 );
not NOT1_15102 ( P1_R1150_U210 , P1_R1150_U44 );
nand NAND2_15103 ( P1_R1150_U211 , P1_U3482 , P1_R1150_U41 );
nand NAND2_15104 ( P1_R1150_U212 , P1_R1150_U117 , P1_R1150_U44 );
nand NAND2_15105 ( P1_R1150_U213 , P1_R1150_U41 , P1_R1150_U40 );
nand NAND2_15106 ( P1_R1150_U214 , P1_R1150_U213 , P1_R1150_U38 );
nand NAND2_15107 ( P1_R1150_U215 , P1_U3084 , P1_R1150_U178 );
not NOT1_15108 ( P1_R1150_U216 , P1_R1150_U148 );
nand NAND2_15109 ( P1_R1150_U217 , P1_U3485 , P1_R1150_U43 );
nand NAND2_15110 ( P1_R1150_U218 , P1_R1150_U217 , P1_R1150_U54 );
nand NAND2_15111 ( P1_R1150_U219 , P1_R1150_U210 , P1_R1150_U40 );
nand NAND2_15112 ( P1_R1150_U220 , P1_R1150_U120 , P1_R1150_U219 );
nand NAND2_15113 ( P1_R1150_U221 , P1_R1150_U44 , P1_R1150_U185 );
nand NAND2_15114 ( P1_R1150_U222 , P1_R1150_U119 , P1_R1150_U221 );
nand NAND2_15115 ( P1_R1150_U223 , P1_R1150_U40 , P1_R1150_U185 );
nand NAND2_15116 ( P1_R1150_U224 , P1_R1150_U206 , P1_R1150_U152 );
not NOT1_15117 ( P1_R1150_U225 , P1_R1150_U45 );
nand NAND2_15118 ( P1_R1150_U226 , P1_U3067 , P1_R1150_U32 );
nand NAND2_15119 ( P1_R1150_U227 , P1_R1150_U225 , P1_R1150_U226 );
nand NAND2_15120 ( P1_R1150_U228 , P1_R1150_U122 , P1_R1150_U227 );
nand NAND2_15121 ( P1_R1150_U229 , P1_R1150_U45 , P1_R1150_U184 );
nand NAND2_15122 ( P1_R1150_U230 , P1_U3476 , P1_R1150_U34 );
nand NAND2_15123 ( P1_R1150_U231 , P1_R1150_U121 , P1_R1150_U229 );
nand NAND2_15124 ( P1_R1150_U232 , P1_U3067 , P1_R1150_U32 );
nand NAND2_15125 ( P1_R1150_U233 , P1_R1150_U184 , P1_R1150_U232 );
nand NAND2_15126 ( P1_R1150_U234 , P1_R1150_U206 , P1_R1150_U37 );
nand NAND2_15127 ( P1_R1150_U235 , P1_R1150_U194 , P1_R1150_U29 );
nand NAND2_15128 ( P1_R1150_U236 , P1_R1150_U124 , P1_R1150_U235 );
nand NAND2_15129 ( P1_R1150_U237 , P1_R1150_U46 , P1_R1150_U183 );
nand NAND2_15130 ( P1_R1150_U238 , P1_R1150_U123 , P1_R1150_U237 );
nand NAND2_15131 ( P1_R1150_U239 , P1_R1150_U29 , P1_R1150_U183 );
nand NAND2_15132 ( P1_R1150_U240 , P1_U3491 , P1_R1150_U52 );
nand NAND2_15133 ( P1_R1150_U241 , P1_U3063 , P1_R1150_U50 );
nand NAND2_15134 ( P1_R1150_U242 , P1_U3062 , P1_R1150_U51 );
nand NAND2_15135 ( P1_R1150_U243 , P1_R1150_U189 , P1_R1150_U8 );
nand NAND2_15136 ( P1_R1150_U244 , P1_R1150_U9 , P1_R1150_U243 );
nand NAND2_15137 ( P1_R1150_U245 , P1_U3491 , P1_R1150_U52 );
nand NAND2_15138 ( P1_R1150_U246 , P1_R1150_U125 , P1_R1150_U148 );
nand NAND2_15139 ( P1_R1150_U247 , P1_R1150_U245 , P1_R1150_U244 );
not NOT1_15140 ( P1_R1150_U248 , P1_R1150_U173 );
nand NAND2_15141 ( P1_R1150_U249 , P1_U3494 , P1_R1150_U56 );
nand NAND2_15142 ( P1_R1150_U250 , P1_R1150_U249 , P1_R1150_U173 );
nand NAND2_15143 ( P1_R1150_U251 , P1_U3072 , P1_R1150_U55 );
not NOT1_15144 ( P1_R1150_U252 , P1_R1150_U172 );
nand NAND2_15145 ( P1_R1150_U253 , P1_U3497 , P1_R1150_U58 );
nand NAND2_15146 ( P1_R1150_U254 , P1_R1150_U253 , P1_R1150_U172 );
nand NAND2_15147 ( P1_R1150_U255 , P1_U3080 , P1_R1150_U57 );
not NOT1_15148 ( P1_R1150_U256 , P1_R1150_U171 );
nand NAND2_15149 ( P1_R1150_U257 , P1_U3506 , P1_R1150_U61 );
nand NAND2_15150 ( P1_R1150_U258 , P1_U3073 , P1_R1150_U59 );
nand NAND2_15151 ( P1_R1150_U259 , P1_U3074 , P1_R1150_U49 );
nand NAND2_15152 ( P1_R1150_U260 , P1_R1150_U186 , P1_R1150_U180 );
nand NAND2_15153 ( P1_R1150_U261 , P1_R1150_U10 , P1_R1150_U260 );
nand NAND2_15154 ( P1_R1150_U262 , P1_U3500 , P1_R1150_U63 );
nand NAND2_15155 ( P1_R1150_U263 , P1_U3506 , P1_R1150_U61 );
nand NAND3_15156 ( P1_R1150_U264 , P1_R1150_U171 , P1_R1150_U126 , P1_R1150_U257 );
nand NAND2_15157 ( P1_R1150_U265 , P1_R1150_U263 , P1_R1150_U261 );
not NOT1_15158 ( P1_R1150_U266 , P1_R1150_U168 );
nand NAND2_15159 ( P1_R1150_U267 , P1_U3509 , P1_R1150_U66 );
nand NAND2_15160 ( P1_R1150_U268 , P1_R1150_U267 , P1_R1150_U168 );
nand NAND2_15161 ( P1_R1150_U269 , P1_U3069 , P1_R1150_U65 );
not NOT1_15162 ( P1_R1150_U270 , P1_R1150_U67 );
nand NAND2_15163 ( P1_R1150_U271 , P1_R1150_U270 , P1_R1150_U68 );
nand NAND2_15164 ( P1_R1150_U272 , P1_R1150_U271 , P1_R1150_U167 );
nand NAND2_15165 ( P1_R1150_U273 , P1_U3082 , P1_R1150_U67 );
not NOT1_15166 ( P1_R1150_U274 , P1_R1150_U166 );
nand NAND2_15167 ( P1_R1150_U275 , P1_U3514 , P1_R1150_U70 );
nand NAND2_15168 ( P1_R1150_U276 , P1_R1150_U275 , P1_R1150_U166 );
nand NAND2_15169 ( P1_R1150_U277 , P1_U3081 , P1_R1150_U69 );
not NOT1_15170 ( P1_R1150_U278 , P1_R1150_U164 );
nand NAND2_15171 ( P1_R1150_U279 , P1_U4025 , P1_R1150_U72 );
nand NAND2_15172 ( P1_R1150_U280 , P1_R1150_U279 , P1_R1150_U164 );
nand NAND2_15173 ( P1_R1150_U281 , P1_U3076 , P1_R1150_U71 );
not NOT1_15174 ( P1_R1150_U282 , P1_R1150_U163 );
nand NAND2_15175 ( P1_R1150_U283 , P1_U4022 , P1_R1150_U75 );
nand NAND2_15176 ( P1_R1150_U284 , P1_U3066 , P1_R1150_U73 );
nand NAND2_15177 ( P1_R1150_U285 , P1_U3061 , P1_R1150_U48 );
nand NAND2_15178 ( P1_R1150_U286 , P1_R1150_U187 , P1_R1150_U181 );
nand NAND2_15179 ( P1_R1150_U287 , P1_R1150_U11 , P1_R1150_U286 );
nand NAND2_15180 ( P1_R1150_U288 , P1_U4024 , P1_R1150_U77 );
nand NAND2_15181 ( P1_R1150_U289 , P1_U4022 , P1_R1150_U75 );
nand NAND3_15182 ( P1_R1150_U290 , P1_R1150_U163 , P1_R1150_U127 , P1_R1150_U283 );
nand NAND2_15183 ( P1_R1150_U291 , P1_R1150_U289 , P1_R1150_U287 );
not NOT1_15184 ( P1_R1150_U292 , P1_R1150_U160 );
nand NAND2_15185 ( P1_R1150_U293 , P1_U4021 , P1_R1150_U80 );
nand NAND2_15186 ( P1_R1150_U294 , P1_R1150_U293 , P1_R1150_U160 );
nand NAND2_15187 ( P1_R1150_U295 , P1_U3065 , P1_R1150_U79 );
not NOT1_15188 ( P1_R1150_U296 , P1_R1150_U159 );
nand NAND2_15189 ( P1_R1150_U297 , P1_U4020 , P1_R1150_U82 );
nand NAND2_15190 ( P1_R1150_U298 , P1_R1150_U297 , P1_R1150_U159 );
nand NAND2_15191 ( P1_R1150_U299 , P1_U3058 , P1_R1150_U81 );
not NOT1_15192 ( P1_R1150_U300 , P1_R1150_U89 );
nand NAND2_15193 ( P1_R1150_U301 , P1_U4018 , P1_R1150_U86 );
nand NAND3_15194 ( P1_R1150_U302 , P1_R1150_U89 , P1_R1150_U182 , P1_R1150_U301 );
nand NAND2_15195 ( P1_R1150_U303 , P1_R1150_U86 , P1_R1150_U85 );
nand NAND2_15196 ( P1_R1150_U304 , P1_R1150_U303 , P1_R1150_U83 );
nand NAND2_15197 ( P1_R1150_U305 , P1_U3053 , P1_R1150_U176 );
not NOT1_15198 ( P1_R1150_U306 , P1_R1150_U157 );
nand NAND2_15199 ( P1_R1150_U307 , P1_U4017 , P1_R1150_U88 );
nand NAND2_15200 ( P1_R1150_U308 , P1_U3054 , P1_R1150_U87 );
nand NAND2_15201 ( P1_R1150_U309 , P1_R1150_U300 , P1_R1150_U85 );
nand NAND2_15202 ( P1_R1150_U310 , P1_R1150_U133 , P1_R1150_U309 );
nand NAND2_15203 ( P1_R1150_U311 , P1_R1150_U89 , P1_R1150_U182 );
nand NAND2_15204 ( P1_R1150_U312 , P1_R1150_U132 , P1_R1150_U311 );
nand NAND2_15205 ( P1_R1150_U313 , P1_R1150_U85 , P1_R1150_U182 );
nand NAND2_15206 ( P1_R1150_U314 , P1_R1150_U288 , P1_R1150_U163 );
not NOT1_15207 ( P1_R1150_U315 , P1_R1150_U90 );
nand NAND2_15208 ( P1_R1150_U316 , P1_U3061 , P1_R1150_U48 );
nand NAND2_15209 ( P1_R1150_U317 , P1_R1150_U315 , P1_R1150_U316 );
nand NAND2_15210 ( P1_R1150_U318 , P1_R1150_U136 , P1_R1150_U317 );
nand NAND2_15211 ( P1_R1150_U319 , P1_R1150_U90 , P1_R1150_U181 );
nand NAND2_15212 ( P1_R1150_U320 , P1_U4022 , P1_R1150_U75 );
nand NAND3_15213 ( P1_R1150_U321 , P1_R1150_U320 , P1_R1150_U319 , P1_R1150_U11 );
nand NAND2_15214 ( P1_R1150_U322 , P1_U3061 , P1_R1150_U48 );
nand NAND2_15215 ( P1_R1150_U323 , P1_R1150_U181 , P1_R1150_U322 );
nand NAND2_15216 ( P1_R1150_U324 , P1_R1150_U288 , P1_R1150_U78 );
nand NAND2_15217 ( P1_R1150_U325 , P1_R1150_U262 , P1_R1150_U171 );
not NOT1_15218 ( P1_R1150_U326 , P1_R1150_U91 );
nand NAND2_15219 ( P1_R1150_U327 , P1_U3074 , P1_R1150_U49 );
nand NAND2_15220 ( P1_R1150_U328 , P1_R1150_U326 , P1_R1150_U327 );
nand NAND2_15221 ( P1_R1150_U329 , P1_R1150_U142 , P1_R1150_U328 );
nand NAND2_15222 ( P1_R1150_U330 , P1_R1150_U91 , P1_R1150_U180 );
nand NAND2_15223 ( P1_R1150_U331 , P1_U3506 , P1_R1150_U61 );
nand NAND3_15224 ( P1_R1150_U332 , P1_R1150_U331 , P1_R1150_U330 , P1_R1150_U10 );
nand NAND2_15225 ( P1_R1150_U333 , P1_U3074 , P1_R1150_U49 );
nand NAND2_15226 ( P1_R1150_U334 , P1_R1150_U180 , P1_R1150_U333 );
nand NAND2_15227 ( P1_R1150_U335 , P1_R1150_U262 , P1_R1150_U64 );
nand NAND2_15228 ( P1_R1150_U336 , P1_R1150_U217 , P1_R1150_U148 );
not NOT1_15229 ( P1_R1150_U337 , P1_R1150_U92 );
nand NAND2_15230 ( P1_R1150_U338 , P1_U3062 , P1_R1150_U51 );
nand NAND2_15231 ( P1_R1150_U339 , P1_R1150_U337 , P1_R1150_U338 );
nand NAND2_15232 ( P1_R1150_U340 , P1_R1150_U146 , P1_R1150_U339 );
nand NAND2_15233 ( P1_R1150_U341 , P1_R1150_U92 , P1_R1150_U179 );
nand NAND2_15234 ( P1_R1150_U342 , P1_U3491 , P1_R1150_U52 );
nand NAND2_15235 ( P1_R1150_U343 , P1_R1150_U145 , P1_R1150_U341 );
nand NAND2_15236 ( P1_R1150_U344 , P1_U3062 , P1_R1150_U51 );
nand NAND2_15237 ( P1_R1150_U345 , P1_R1150_U179 , P1_R1150_U344 );
nand NAND2_15238 ( P1_R1150_U346 , P1_U3077 , P1_R1150_U24 );
nand NAND3_15239 ( P1_R1150_U347 , P1_R1150_U89 , P1_R1150_U182 , P1_R1150_U301 );
nand NAND3_15240 ( P1_R1150_U348 , P1_R1150_U12 , P1_R1150_U347 , P1_R1150_U130 );
nand NAND2_15241 ( P1_R1150_U349 , P1_U3485 , P1_R1150_U43 );
nand NAND2_15242 ( P1_R1150_U350 , P1_U3083 , P1_R1150_U42 );
nand NAND2_15243 ( P1_R1150_U351 , P1_R1150_U218 , P1_R1150_U148 );
nand NAND2_15244 ( P1_R1150_U352 , P1_R1150_U216 , P1_R1150_U147 );
nand NAND2_15245 ( P1_R1150_U353 , P1_U3482 , P1_R1150_U41 );
nand NAND2_15246 ( P1_R1150_U354 , P1_U3084 , P1_R1150_U38 );
nand NAND2_15247 ( P1_R1150_U355 , P1_U3482 , P1_R1150_U41 );
nand NAND2_15248 ( P1_R1150_U356 , P1_U3084 , P1_R1150_U38 );
nand NAND2_15249 ( P1_R1150_U357 , P1_R1150_U356 , P1_R1150_U355 );
nand NAND2_15250 ( P1_R1150_U358 , P1_U3479 , P1_R1150_U39 );
nand NAND2_15251 ( P1_R1150_U359 , P1_U3070 , P1_R1150_U22 );
nand NAND2_15252 ( P1_R1150_U360 , P1_R1150_U223 , P1_R1150_U44 );
nand NAND2_15253 ( P1_R1150_U361 , P1_R1150_U149 , P1_R1150_U210 );
nand NAND2_15254 ( P1_R1150_U362 , P1_U3476 , P1_R1150_U34 );
nand NAND2_15255 ( P1_R1150_U363 , P1_U3071 , P1_R1150_U31 );
nand NAND2_15256 ( P1_R1150_U364 , P1_R1150_U363 , P1_R1150_U362 );
nand NAND2_15257 ( P1_R1150_U365 , P1_U3473 , P1_R1150_U35 );
nand NAND2_15258 ( P1_R1150_U366 , P1_U3067 , P1_R1150_U32 );
nand NAND2_15259 ( P1_R1150_U367 , P1_R1150_U233 , P1_R1150_U45 );
nand NAND2_15260 ( P1_R1150_U368 , P1_R1150_U150 , P1_R1150_U225 );
nand NAND2_15261 ( P1_R1150_U369 , P1_U3470 , P1_R1150_U36 );
nand NAND2_15262 ( P1_R1150_U370 , P1_U3060 , P1_R1150_U33 );
nand NAND2_15263 ( P1_R1150_U371 , P1_R1150_U234 , P1_R1150_U152 );
nand NAND2_15264 ( P1_R1150_U372 , P1_R1150_U200 , P1_R1150_U151 );
nand NAND2_15265 ( P1_R1150_U373 , P1_U3467 , P1_R1150_U30 );
nand NAND2_15266 ( P1_R1150_U374 , P1_U3064 , P1_R1150_U27 );
nand NAND2_15267 ( P1_R1150_U375 , P1_U3467 , P1_R1150_U30 );
nand NAND2_15268 ( P1_R1150_U376 , P1_U3064 , P1_R1150_U27 );
nand NAND2_15269 ( P1_R1150_U377 , P1_R1150_U376 , P1_R1150_U375 );
nand NAND2_15270 ( P1_R1150_U378 , P1_U3464 , P1_R1150_U28 );
nand NAND2_15271 ( P1_R1150_U379 , P1_U3068 , P1_R1150_U23 );
nand NAND2_15272 ( P1_R1150_U380 , P1_R1150_U239 , P1_R1150_U46 );
nand NAND2_15273 ( P1_R1150_U381 , P1_R1150_U153 , P1_R1150_U194 );
nand NAND2_15274 ( P1_R1150_U382 , P1_U4028 , P1_R1150_U155 );
nand NAND2_15275 ( P1_R1150_U383 , P1_U3055 , P1_R1150_U154 );
nand NAND2_15276 ( P1_R1150_U384 , P1_U4028 , P1_R1150_U155 );
nand NAND2_15277 ( P1_R1150_U385 , P1_U3055 , P1_R1150_U154 );
nand NAND2_15278 ( P1_R1150_U386 , P1_R1150_U385 , P1_R1150_U384 );
nand NAND3_15279 ( P1_R1150_U387 , P1_U3054 , P1_R1150_U386 , P1_R1150_U87 );
nand NAND3_15280 ( P1_R1150_U388 , P1_R1150_U12 , P1_R1150_U88 , P1_U4017 );
nand NAND2_15281 ( P1_R1150_U389 , P1_U4017 , P1_R1150_U88 );
nand NAND2_15282 ( P1_R1150_U390 , P1_U3054 , P1_R1150_U87 );
not NOT1_15283 ( P1_R1150_U391 , P1_R1150_U131 );
nand NAND2_15284 ( P1_R1150_U392 , P1_R1150_U306 , P1_R1150_U391 );
nand NAND2_15285 ( P1_R1150_U393 , P1_R1150_U131 , P1_R1150_U157 );
nand NAND2_15286 ( P1_R1150_U394 , P1_U4018 , P1_R1150_U86 );
nand NAND2_15287 ( P1_R1150_U395 , P1_U3053 , P1_R1150_U83 );
nand NAND2_15288 ( P1_R1150_U396 , P1_U4018 , P1_R1150_U86 );
nand NAND2_15289 ( P1_R1150_U397 , P1_U3053 , P1_R1150_U83 );
nand NAND2_15290 ( P1_R1150_U398 , P1_R1150_U397 , P1_R1150_U396 );
nand NAND2_15291 ( P1_R1150_U399 , P1_U4019 , P1_R1150_U84 );
nand NAND2_15292 ( P1_R1150_U400 , P1_U3057 , P1_R1150_U47 );
nand NAND2_15293 ( P1_R1150_U401 , P1_R1150_U313 , P1_R1150_U89 );
nand NAND2_15294 ( P1_R1150_U402 , P1_R1150_U158 , P1_R1150_U300 );
nand NAND2_15295 ( P1_R1150_U403 , P1_U4020 , P1_R1150_U82 );
nand NAND2_15296 ( P1_R1150_U404 , P1_U3058 , P1_R1150_U81 );
not NOT1_15297 ( P1_R1150_U405 , P1_R1150_U134 );
nand NAND2_15298 ( P1_R1150_U406 , P1_R1150_U296 , P1_R1150_U405 );
nand NAND2_15299 ( P1_R1150_U407 , P1_R1150_U134 , P1_R1150_U159 );
nand NAND2_15300 ( P1_R1150_U408 , P1_U4021 , P1_R1150_U80 );
nand NAND2_15301 ( P1_R1150_U409 , P1_U3065 , P1_R1150_U79 );
not NOT1_15302 ( P1_R1150_U410 , P1_R1150_U135 );
nand NAND2_15303 ( P1_R1150_U411 , P1_R1150_U292 , P1_R1150_U410 );
nand NAND2_15304 ( P1_R1150_U412 , P1_R1150_U135 , P1_R1150_U160 );
nand NAND2_15305 ( P1_R1150_U413 , P1_U4022 , P1_R1150_U75 );
nand NAND2_15306 ( P1_R1150_U414 , P1_U3066 , P1_R1150_U73 );
nand NAND2_15307 ( P1_R1150_U415 , P1_R1150_U414 , P1_R1150_U413 );
nand NAND2_15308 ( P1_R1150_U416 , P1_U4023 , P1_R1150_U76 );
nand NAND2_15309 ( P1_R1150_U417 , P1_U3061 , P1_R1150_U48 );
nand NAND2_15310 ( P1_R1150_U418 , P1_R1150_U323 , P1_R1150_U90 );
nand NAND2_15311 ( P1_R1150_U419 , P1_R1150_U161 , P1_R1150_U315 );
nand NAND2_15312 ( P1_R1150_U420 , P1_U4024 , P1_R1150_U77 );
nand NAND2_15313 ( P1_R1150_U421 , P1_U3075 , P1_R1150_U74 );
nand NAND2_15314 ( P1_R1150_U422 , P1_R1150_U324 , P1_R1150_U163 );
nand NAND2_15315 ( P1_R1150_U423 , P1_R1150_U282 , P1_R1150_U162 );
nand NAND2_15316 ( P1_R1150_U424 , P1_U4025 , P1_R1150_U72 );
nand NAND2_15317 ( P1_R1150_U425 , P1_U3076 , P1_R1150_U71 );
not NOT1_15318 ( P1_R1150_U426 , P1_R1150_U137 );
nand NAND2_15319 ( P1_R1150_U427 , P1_R1150_U278 , P1_R1150_U426 );
nand NAND2_15320 ( P1_R1150_U428 , P1_R1150_U137 , P1_R1150_U164 );
nand NAND2_15321 ( P1_R1150_U429 , P1_U3461 , P1_R1150_U26 );
nand NAND2_15322 ( P1_R1150_U430 , P1_U3078 , P1_R1150_U165 );
not NOT1_15323 ( P1_R1150_U431 , P1_R1150_U138 );
nand NAND2_15324 ( P1_R1150_U432 , P1_R1150_U431 , P1_R1150_U190 );
nand NAND2_15325 ( P1_R1150_U433 , P1_R1150_U138 , P1_R1150_U25 );
nand NAND2_15326 ( P1_R1150_U434 , P1_U3514 , P1_R1150_U70 );
nand NAND2_15327 ( P1_R1150_U435 , P1_U3081 , P1_R1150_U69 );
not NOT1_15328 ( P1_R1150_U436 , P1_R1150_U139 );
nand NAND2_15329 ( P1_R1150_U437 , P1_R1150_U274 , P1_R1150_U436 );
nand NAND2_15330 ( P1_R1150_U438 , P1_R1150_U139 , P1_R1150_U166 );
nand NAND2_15331 ( P1_R1150_U439 , P1_U3512 , P1_R1150_U68 );
nand NAND2_15332 ( P1_R1150_U440 , P1_U3082 , P1_R1150_U167 );
not NOT1_15333 ( P1_R1150_U441 , P1_R1150_U140 );
nand NAND2_15334 ( P1_R1150_U442 , P1_R1150_U441 , P1_R1150_U270 );
nand NAND2_15335 ( P1_R1150_U443 , P1_R1150_U140 , P1_R1150_U67 );
nand NAND2_15336 ( P1_R1150_U444 , P1_U3509 , P1_R1150_U66 );
nand NAND2_15337 ( P1_R1150_U445 , P1_U3069 , P1_R1150_U65 );
not NOT1_15338 ( P1_R1150_U446 , P1_R1150_U141 );
nand NAND2_15339 ( P1_R1150_U447 , P1_R1150_U266 , P1_R1150_U446 );
nand NAND2_15340 ( P1_R1150_U448 , P1_R1150_U141 , P1_R1150_U168 );
nand NAND2_15341 ( P1_R1150_U449 , P1_U3506 , P1_R1150_U61 );
nand NAND2_15342 ( P1_R1150_U450 , P1_U3073 , P1_R1150_U59 );
nand NAND2_15343 ( P1_R1150_U451 , P1_R1150_U450 , P1_R1150_U449 );
nand NAND2_15344 ( P1_R1150_U452 , P1_U3503 , P1_R1150_U62 );
nand NAND2_15345 ( P1_R1150_U453 , P1_U3074 , P1_R1150_U49 );
nand NAND2_15346 ( P1_R1150_U454 , P1_R1150_U334 , P1_R1150_U91 );
nand NAND2_15347 ( P1_R1150_U455 , P1_R1150_U169 , P1_R1150_U326 );
nand NAND2_15348 ( P1_R1150_U456 , P1_U3500 , P1_R1150_U63 );
nand NAND2_15349 ( P1_R1150_U457 , P1_U3079 , P1_R1150_U60 );
nand NAND2_15350 ( P1_R1150_U458 , P1_R1150_U335 , P1_R1150_U171 );
nand NAND2_15351 ( P1_R1150_U459 , P1_R1150_U256 , P1_R1150_U170 );
nand NAND2_15352 ( P1_R1150_U460 , P1_U3497 , P1_R1150_U58 );
nand NAND2_15353 ( P1_R1150_U461 , P1_U3080 , P1_R1150_U57 );
not NOT1_15354 ( P1_R1150_U462 , P1_R1150_U143 );
nand NAND2_15355 ( P1_R1150_U463 , P1_R1150_U252 , P1_R1150_U462 );
nand NAND2_15356 ( P1_R1150_U464 , P1_R1150_U143 , P1_R1150_U172 );
nand NAND2_15357 ( P1_R1150_U465 , P1_U3494 , P1_R1150_U56 );
nand NAND2_15358 ( P1_R1150_U466 , P1_U3072 , P1_R1150_U55 );
not NOT1_15359 ( P1_R1150_U467 , P1_R1150_U144 );
nand NAND2_15360 ( P1_R1150_U468 , P1_R1150_U248 , P1_R1150_U467 );
nand NAND2_15361 ( P1_R1150_U469 , P1_R1150_U144 , P1_R1150_U173 );
nand NAND2_15362 ( P1_R1150_U470 , P1_U3491 , P1_R1150_U52 );
nand NAND2_15363 ( P1_R1150_U471 , P1_U3063 , P1_R1150_U50 );
nand NAND2_15364 ( P1_R1150_U472 , P1_R1150_U471 , P1_R1150_U470 );
nand NAND2_15365 ( P1_R1150_U473 , P1_U3488 , P1_R1150_U53 );
nand NAND2_15366 ( P1_R1150_U474 , P1_U3062 , P1_R1150_U51 );
nand NAND2_15367 ( P1_R1150_U475 , P1_R1150_U345 , P1_R1150_U92 );
nand NAND2_15368 ( P1_R1150_U476 , P1_R1150_U174 , P1_R1150_U337 );
and AND2_15369 ( P1_R1192_U6 , P1_R1192_U184 , P1_R1192_U201 );
and AND2_15370 ( P1_R1192_U7 , P1_R1192_U203 , P1_R1192_U202 );
and AND2_15371 ( P1_R1192_U8 , P1_R1192_U179 , P1_R1192_U240 );
and AND2_15372 ( P1_R1192_U9 , P1_R1192_U242 , P1_R1192_U241 );
and AND2_15373 ( P1_R1192_U10 , P1_R1192_U259 , P1_R1192_U258 );
and AND2_15374 ( P1_R1192_U11 , P1_R1192_U285 , P1_R1192_U284 );
and AND2_15375 ( P1_R1192_U12 , P1_R1192_U383 , P1_R1192_U382 );
nand NAND2_15376 ( P1_R1192_U13 , P1_R1192_U340 , P1_R1192_U343 );
nand NAND2_15377 ( P1_R1192_U14 , P1_R1192_U329 , P1_R1192_U332 );
nand NAND2_15378 ( P1_R1192_U15 , P1_R1192_U318 , P1_R1192_U321 );
nand NAND2_15379 ( P1_R1192_U16 , P1_R1192_U310 , P1_R1192_U312 );
nand NAND3_15380 ( P1_R1192_U17 , P1_R1192_U156 , P1_R1192_U175 , P1_R1192_U348 );
nand NAND2_15381 ( P1_R1192_U18 , P1_R1192_U236 , P1_R1192_U238 );
nand NAND2_15382 ( P1_R1192_U19 , P1_R1192_U228 , P1_R1192_U231 );
nand NAND2_15383 ( P1_R1192_U20 , P1_R1192_U220 , P1_R1192_U222 );
nand NAND2_15384 ( P1_R1192_U21 , P1_R1192_U25 , P1_R1192_U346 );
not NOT1_15385 ( P1_R1192_U22 , P1_U3479 );
not NOT1_15386 ( P1_R1192_U23 , P1_U3464 );
not NOT1_15387 ( P1_R1192_U24 , P1_U3456 );
nand NAND2_15388 ( P1_R1192_U25 , P1_U3456 , P1_R1192_U93 );
not NOT1_15389 ( P1_R1192_U26 , P1_U3078 );
not NOT1_15390 ( P1_R1192_U27 , P1_U3467 );
not NOT1_15391 ( P1_R1192_U28 , P1_U3068 );
nand NAND2_15392 ( P1_R1192_U29 , P1_U3068 , P1_R1192_U23 );
not NOT1_15393 ( P1_R1192_U30 , P1_U3064 );
not NOT1_15394 ( P1_R1192_U31 , P1_U3476 );
not NOT1_15395 ( P1_R1192_U32 , P1_U3473 );
not NOT1_15396 ( P1_R1192_U33 , P1_U3470 );
not NOT1_15397 ( P1_R1192_U34 , P1_U3071 );
not NOT1_15398 ( P1_R1192_U35 , P1_U3067 );
not NOT1_15399 ( P1_R1192_U36 , P1_U3060 );
nand NAND2_15400 ( P1_R1192_U37 , P1_U3060 , P1_R1192_U33 );
not NOT1_15401 ( P1_R1192_U38 , P1_U3482 );
not NOT1_15402 ( P1_R1192_U39 , P1_U3070 );
nand NAND2_15403 ( P1_R1192_U40 , P1_U3070 , P1_R1192_U22 );
not NOT1_15404 ( P1_R1192_U41 , P1_U3084 );
not NOT1_15405 ( P1_R1192_U42 , P1_U3485 );
not NOT1_15406 ( P1_R1192_U43 , P1_U3083 );
nand NAND2_15407 ( P1_R1192_U44 , P1_R1192_U209 , P1_R1192_U208 );
nand NAND2_15408 ( P1_R1192_U45 , P1_R1192_U37 , P1_R1192_U224 );
nand NAND2_15409 ( P1_R1192_U46 , P1_R1192_U193 , P1_R1192_U192 );
not NOT1_15410 ( P1_R1192_U47 , P1_U4019 );
not NOT1_15411 ( P1_R1192_U48 , P1_U4023 );
not NOT1_15412 ( P1_R1192_U49 , P1_U3503 );
not NOT1_15413 ( P1_R1192_U50 , P1_U3491 );
not NOT1_15414 ( P1_R1192_U51 , P1_U3488 );
not NOT1_15415 ( P1_R1192_U52 , P1_U3063 );
not NOT1_15416 ( P1_R1192_U53 , P1_U3062 );
nand NAND2_15417 ( P1_R1192_U54 , P1_U3083 , P1_R1192_U42 );
not NOT1_15418 ( P1_R1192_U55 , P1_U3494 );
not NOT1_15419 ( P1_R1192_U56 , P1_U3072 );
not NOT1_15420 ( P1_R1192_U57 , P1_U3497 );
not NOT1_15421 ( P1_R1192_U58 , P1_U3080 );
not NOT1_15422 ( P1_R1192_U59 , P1_U3506 );
not NOT1_15423 ( P1_R1192_U60 , P1_U3500 );
not NOT1_15424 ( P1_R1192_U61 , P1_U3073 );
not NOT1_15425 ( P1_R1192_U62 , P1_U3074 );
not NOT1_15426 ( P1_R1192_U63 , P1_U3079 );
nand NAND2_15427 ( P1_R1192_U64 , P1_U3079 , P1_R1192_U60 );
not NOT1_15428 ( P1_R1192_U65 , P1_U3509 );
not NOT1_15429 ( P1_R1192_U66 , P1_U3069 );
nand NAND2_15430 ( P1_R1192_U67 , P1_R1192_U269 , P1_R1192_U268 );
not NOT1_15431 ( P1_R1192_U68 , P1_U3082 );
not NOT1_15432 ( P1_R1192_U69 , P1_U3514 );
not NOT1_15433 ( P1_R1192_U70 , P1_U3081 );
not NOT1_15434 ( P1_R1192_U71 , P1_U4025 );
not NOT1_15435 ( P1_R1192_U72 , P1_U3076 );
not NOT1_15436 ( P1_R1192_U73 , P1_U4022 );
not NOT1_15437 ( P1_R1192_U74 , P1_U4024 );
not NOT1_15438 ( P1_R1192_U75 , P1_U3066 );
not NOT1_15439 ( P1_R1192_U76 , P1_U3061 );
not NOT1_15440 ( P1_R1192_U77 , P1_U3075 );
nand NAND2_15441 ( P1_R1192_U78 , P1_U3075 , P1_R1192_U74 );
not NOT1_15442 ( P1_R1192_U79 , P1_U4021 );
not NOT1_15443 ( P1_R1192_U80 , P1_U3065 );
not NOT1_15444 ( P1_R1192_U81 , P1_U4020 );
not NOT1_15445 ( P1_R1192_U82 , P1_U3058 );
not NOT1_15446 ( P1_R1192_U83 , P1_U4018 );
not NOT1_15447 ( P1_R1192_U84 , P1_U3057 );
nand NAND2_15448 ( P1_R1192_U85 , P1_U3057 , P1_R1192_U47 );
not NOT1_15449 ( P1_R1192_U86 , P1_U3053 );
not NOT1_15450 ( P1_R1192_U87 , P1_U4017 );
not NOT1_15451 ( P1_R1192_U88 , P1_U3054 );
nand NAND2_15452 ( P1_R1192_U89 , P1_R1192_U299 , P1_R1192_U298 );
nand NAND2_15453 ( P1_R1192_U90 , P1_R1192_U78 , P1_R1192_U314 );
nand NAND2_15454 ( P1_R1192_U91 , P1_R1192_U64 , P1_R1192_U325 );
nand NAND2_15455 ( P1_R1192_U92 , P1_R1192_U54 , P1_R1192_U336 );
not NOT1_15456 ( P1_R1192_U93 , P1_U3077 );
nand NAND2_15457 ( P1_R1192_U94 , P1_R1192_U393 , P1_R1192_U392 );
nand NAND2_15458 ( P1_R1192_U95 , P1_R1192_U407 , P1_R1192_U406 );
nand NAND2_15459 ( P1_R1192_U96 , P1_R1192_U412 , P1_R1192_U411 );
nand NAND2_15460 ( P1_R1192_U97 , P1_R1192_U428 , P1_R1192_U427 );
nand NAND2_15461 ( P1_R1192_U98 , P1_R1192_U433 , P1_R1192_U432 );
nand NAND2_15462 ( P1_R1192_U99 , P1_R1192_U438 , P1_R1192_U437 );
nand NAND2_15463 ( P1_R1192_U100 , P1_R1192_U443 , P1_R1192_U442 );
nand NAND2_15464 ( P1_R1192_U101 , P1_R1192_U448 , P1_R1192_U447 );
nand NAND2_15465 ( P1_R1192_U102 , P1_R1192_U464 , P1_R1192_U463 );
nand NAND2_15466 ( P1_R1192_U103 , P1_R1192_U469 , P1_R1192_U468 );
nand NAND2_15467 ( P1_R1192_U104 , P1_R1192_U352 , P1_R1192_U351 );
nand NAND2_15468 ( P1_R1192_U105 , P1_R1192_U361 , P1_R1192_U360 );
nand NAND2_15469 ( P1_R1192_U106 , P1_R1192_U368 , P1_R1192_U367 );
nand NAND2_15470 ( P1_R1192_U107 , P1_R1192_U372 , P1_R1192_U371 );
nand NAND2_15471 ( P1_R1192_U108 , P1_R1192_U381 , P1_R1192_U380 );
nand NAND2_15472 ( P1_R1192_U109 , P1_R1192_U402 , P1_R1192_U401 );
nand NAND2_15473 ( P1_R1192_U110 , P1_R1192_U419 , P1_R1192_U418 );
nand NAND2_15474 ( P1_R1192_U111 , P1_R1192_U423 , P1_R1192_U422 );
nand NAND2_15475 ( P1_R1192_U112 , P1_R1192_U455 , P1_R1192_U454 );
nand NAND2_15476 ( P1_R1192_U113 , P1_R1192_U459 , P1_R1192_U458 );
nand NAND2_15477 ( P1_R1192_U114 , P1_R1192_U476 , P1_R1192_U475 );
and AND2_15478 ( P1_R1192_U115 , P1_R1192_U195 , P1_R1192_U183 );
and AND2_15479 ( P1_R1192_U116 , P1_R1192_U198 , P1_R1192_U199 );
and AND2_15480 ( P1_R1192_U117 , P1_R1192_U211 , P1_R1192_U185 );
and AND2_15481 ( P1_R1192_U118 , P1_R1192_U214 , P1_R1192_U215 );
and AND3_15482 ( P1_R1192_U119 , P1_R1192_U354 , P1_R1192_U353 , P1_R1192_U40 );
and AND2_15483 ( P1_R1192_U120 , P1_R1192_U357 , P1_R1192_U185 );
and AND2_15484 ( P1_R1192_U121 , P1_R1192_U230 , P1_R1192_U7 );
and AND2_15485 ( P1_R1192_U122 , P1_R1192_U364 , P1_R1192_U184 );
and AND3_15486 ( P1_R1192_U123 , P1_R1192_U374 , P1_R1192_U373 , P1_R1192_U29 );
and AND2_15487 ( P1_R1192_U124 , P1_R1192_U377 , P1_R1192_U183 );
and AND2_15488 ( P1_R1192_U125 , P1_R1192_U217 , P1_R1192_U8 );
and AND2_15489 ( P1_R1192_U126 , P1_R1192_U262 , P1_R1192_U180 );
and AND2_15490 ( P1_R1192_U127 , P1_R1192_U288 , P1_R1192_U181 );
and AND2_15491 ( P1_R1192_U128 , P1_R1192_U304 , P1_R1192_U305 );
and AND2_15492 ( P1_R1192_U129 , P1_R1192_U307 , P1_R1192_U386 );
and AND3_15493 ( P1_R1192_U130 , P1_R1192_U305 , P1_R1192_U304 , P1_R1192_U308 );
nand NAND2_15494 ( P1_R1192_U131 , P1_R1192_U390 , P1_R1192_U389 );
and AND3_15495 ( P1_R1192_U132 , P1_R1192_U395 , P1_R1192_U394 , P1_R1192_U85 );
and AND2_15496 ( P1_R1192_U133 , P1_R1192_U398 , P1_R1192_U182 );
nand NAND2_15497 ( P1_R1192_U134 , P1_R1192_U404 , P1_R1192_U403 );
nand NAND2_15498 ( P1_R1192_U135 , P1_R1192_U409 , P1_R1192_U408 );
and AND2_15499 ( P1_R1192_U136 , P1_R1192_U415 , P1_R1192_U181 );
nand NAND2_15500 ( P1_R1192_U137 , P1_R1192_U425 , P1_R1192_U424 );
nand NAND2_15501 ( P1_R1192_U138 , P1_R1192_U430 , P1_R1192_U429 );
nand NAND2_15502 ( P1_R1192_U139 , P1_R1192_U435 , P1_R1192_U434 );
nand NAND2_15503 ( P1_R1192_U140 , P1_R1192_U440 , P1_R1192_U439 );
nand NAND2_15504 ( P1_R1192_U141 , P1_R1192_U445 , P1_R1192_U444 );
and AND2_15505 ( P1_R1192_U142 , P1_R1192_U451 , P1_R1192_U180 );
nand NAND2_15506 ( P1_R1192_U143 , P1_R1192_U461 , P1_R1192_U460 );
nand NAND2_15507 ( P1_R1192_U144 , P1_R1192_U466 , P1_R1192_U465 );
and AND2_15508 ( P1_R1192_U145 , P1_R1192_U342 , P1_R1192_U9 );
and AND2_15509 ( P1_R1192_U146 , P1_R1192_U472 , P1_R1192_U179 );
and AND2_15510 ( P1_R1192_U147 , P1_R1192_U350 , P1_R1192_U349 );
nand NAND2_15511 ( P1_R1192_U148 , P1_R1192_U118 , P1_R1192_U212 );
and AND2_15512 ( P1_R1192_U149 , P1_R1192_U359 , P1_R1192_U358 );
and AND2_15513 ( P1_R1192_U150 , P1_R1192_U366 , P1_R1192_U365 );
and AND2_15514 ( P1_R1192_U151 , P1_R1192_U370 , P1_R1192_U369 );
nand NAND2_15515 ( P1_R1192_U152 , P1_R1192_U116 , P1_R1192_U196 );
and AND2_15516 ( P1_R1192_U153 , P1_R1192_U379 , P1_R1192_U378 );
not NOT1_15517 ( P1_R1192_U154 , P1_U4028 );
not NOT1_15518 ( P1_R1192_U155 , P1_U3055 );
and AND2_15519 ( P1_R1192_U156 , P1_R1192_U388 , P1_R1192_U387 );
nand NAND2_15520 ( P1_R1192_U157 , P1_R1192_U128 , P1_R1192_U302 );
and AND2_15521 ( P1_R1192_U158 , P1_R1192_U400 , P1_R1192_U399 );
nand NAND2_15522 ( P1_R1192_U159 , P1_R1192_U295 , P1_R1192_U294 );
nand NAND2_15523 ( P1_R1192_U160 , P1_R1192_U291 , P1_R1192_U290 );
and AND2_15524 ( P1_R1192_U161 , P1_R1192_U417 , P1_R1192_U416 );
and AND2_15525 ( P1_R1192_U162 , P1_R1192_U421 , P1_R1192_U420 );
nand NAND2_15526 ( P1_R1192_U163 , P1_R1192_U281 , P1_R1192_U280 );
nand NAND2_15527 ( P1_R1192_U164 , P1_R1192_U277 , P1_R1192_U276 );
not NOT1_15528 ( P1_R1192_U165 , P1_U3461 );
nand NAND2_15529 ( P1_R1192_U166 , P1_R1192_U273 , P1_R1192_U272 );
not NOT1_15530 ( P1_R1192_U167 , P1_U3512 );
nand NAND2_15531 ( P1_R1192_U168 , P1_R1192_U265 , P1_R1192_U264 );
and AND2_15532 ( P1_R1192_U169 , P1_R1192_U453 , P1_R1192_U452 );
and AND2_15533 ( P1_R1192_U170 , P1_R1192_U457 , P1_R1192_U456 );
nand NAND2_15534 ( P1_R1192_U171 , P1_R1192_U255 , P1_R1192_U254 );
nand NAND2_15535 ( P1_R1192_U172 , P1_R1192_U251 , P1_R1192_U250 );
nand NAND2_15536 ( P1_R1192_U173 , P1_R1192_U247 , P1_R1192_U246 );
and AND2_15537 ( P1_R1192_U174 , P1_R1192_U474 , P1_R1192_U473 );
nand NAND2_15538 ( P1_R1192_U175 , P1_R1192_U129 , P1_R1192_U157 );
not NOT1_15539 ( P1_R1192_U176 , P1_R1192_U85 );
not NOT1_15540 ( P1_R1192_U177 , P1_R1192_U29 );
not NOT1_15541 ( P1_R1192_U178 , P1_R1192_U40 );
nand NAND2_15542 ( P1_R1192_U179 , P1_U3488 , P1_R1192_U53 );
nand NAND2_15543 ( P1_R1192_U180 , P1_U3503 , P1_R1192_U62 );
nand NAND2_15544 ( P1_R1192_U181 , P1_U4023 , P1_R1192_U76 );
nand NAND2_15545 ( P1_R1192_U182 , P1_U4019 , P1_R1192_U84 );
nand NAND2_15546 ( P1_R1192_U183 , P1_U3464 , P1_R1192_U28 );
nand NAND2_15547 ( P1_R1192_U184 , P1_U3473 , P1_R1192_U35 );
nand NAND2_15548 ( P1_R1192_U185 , P1_U3479 , P1_R1192_U39 );
not NOT1_15549 ( P1_R1192_U186 , P1_R1192_U64 );
not NOT1_15550 ( P1_R1192_U187 , P1_R1192_U78 );
not NOT1_15551 ( P1_R1192_U188 , P1_R1192_U37 );
not NOT1_15552 ( P1_R1192_U189 , P1_R1192_U54 );
not NOT1_15553 ( P1_R1192_U190 , P1_R1192_U25 );
nand NAND2_15554 ( P1_R1192_U191 , P1_R1192_U190 , P1_R1192_U26 );
nand NAND2_15555 ( P1_R1192_U192 , P1_R1192_U191 , P1_R1192_U165 );
nand NAND2_15556 ( P1_R1192_U193 , P1_U3078 , P1_R1192_U25 );
not NOT1_15557 ( P1_R1192_U194 , P1_R1192_U46 );
nand NAND2_15558 ( P1_R1192_U195 , P1_U3467 , P1_R1192_U30 );
nand NAND2_15559 ( P1_R1192_U196 , P1_R1192_U115 , P1_R1192_U46 );
nand NAND2_15560 ( P1_R1192_U197 , P1_R1192_U30 , P1_R1192_U29 );
nand NAND2_15561 ( P1_R1192_U198 , P1_R1192_U197 , P1_R1192_U27 );
nand NAND2_15562 ( P1_R1192_U199 , P1_U3064 , P1_R1192_U177 );
not NOT1_15563 ( P1_R1192_U200 , P1_R1192_U152 );
nand NAND2_15564 ( P1_R1192_U201 , P1_U3476 , P1_R1192_U34 );
nand NAND2_15565 ( P1_R1192_U202 , P1_U3071 , P1_R1192_U31 );
nand NAND2_15566 ( P1_R1192_U203 , P1_U3067 , P1_R1192_U32 );
nand NAND2_15567 ( P1_R1192_U204 , P1_R1192_U188 , P1_R1192_U6 );
nand NAND2_15568 ( P1_R1192_U205 , P1_R1192_U7 , P1_R1192_U204 );
nand NAND2_15569 ( P1_R1192_U206 , P1_U3470 , P1_R1192_U36 );
nand NAND2_15570 ( P1_R1192_U207 , P1_U3476 , P1_R1192_U34 );
nand NAND3_15571 ( P1_R1192_U208 , P1_R1192_U206 , P1_R1192_U152 , P1_R1192_U6 );
nand NAND2_15572 ( P1_R1192_U209 , P1_R1192_U207 , P1_R1192_U205 );
not NOT1_15573 ( P1_R1192_U210 , P1_R1192_U44 );
nand NAND2_15574 ( P1_R1192_U211 , P1_U3482 , P1_R1192_U41 );
nand NAND2_15575 ( P1_R1192_U212 , P1_R1192_U117 , P1_R1192_U44 );
nand NAND2_15576 ( P1_R1192_U213 , P1_R1192_U41 , P1_R1192_U40 );
nand NAND2_15577 ( P1_R1192_U214 , P1_R1192_U213 , P1_R1192_U38 );
nand NAND2_15578 ( P1_R1192_U215 , P1_U3084 , P1_R1192_U178 );
not NOT1_15579 ( P1_R1192_U216 , P1_R1192_U148 );
nand NAND2_15580 ( P1_R1192_U217 , P1_U3485 , P1_R1192_U43 );
nand NAND2_15581 ( P1_R1192_U218 , P1_R1192_U217 , P1_R1192_U54 );
nand NAND2_15582 ( P1_R1192_U219 , P1_R1192_U210 , P1_R1192_U40 );
nand NAND2_15583 ( P1_R1192_U220 , P1_R1192_U120 , P1_R1192_U219 );
nand NAND2_15584 ( P1_R1192_U221 , P1_R1192_U44 , P1_R1192_U185 );
nand NAND2_15585 ( P1_R1192_U222 , P1_R1192_U119 , P1_R1192_U221 );
nand NAND2_15586 ( P1_R1192_U223 , P1_R1192_U40 , P1_R1192_U185 );
nand NAND2_15587 ( P1_R1192_U224 , P1_R1192_U206 , P1_R1192_U152 );
not NOT1_15588 ( P1_R1192_U225 , P1_R1192_U45 );
nand NAND2_15589 ( P1_R1192_U226 , P1_U3067 , P1_R1192_U32 );
nand NAND2_15590 ( P1_R1192_U227 , P1_R1192_U225 , P1_R1192_U226 );
nand NAND2_15591 ( P1_R1192_U228 , P1_R1192_U122 , P1_R1192_U227 );
nand NAND2_15592 ( P1_R1192_U229 , P1_R1192_U45 , P1_R1192_U184 );
nand NAND2_15593 ( P1_R1192_U230 , P1_U3476 , P1_R1192_U34 );
nand NAND2_15594 ( P1_R1192_U231 , P1_R1192_U121 , P1_R1192_U229 );
nand NAND2_15595 ( P1_R1192_U232 , P1_U3067 , P1_R1192_U32 );
nand NAND2_15596 ( P1_R1192_U233 , P1_R1192_U184 , P1_R1192_U232 );
nand NAND2_15597 ( P1_R1192_U234 , P1_R1192_U206 , P1_R1192_U37 );
nand NAND2_15598 ( P1_R1192_U235 , P1_R1192_U194 , P1_R1192_U29 );
nand NAND2_15599 ( P1_R1192_U236 , P1_R1192_U124 , P1_R1192_U235 );
nand NAND2_15600 ( P1_R1192_U237 , P1_R1192_U46 , P1_R1192_U183 );
nand NAND2_15601 ( P1_R1192_U238 , P1_R1192_U123 , P1_R1192_U237 );
nand NAND2_15602 ( P1_R1192_U239 , P1_R1192_U29 , P1_R1192_U183 );
nand NAND2_15603 ( P1_R1192_U240 , P1_U3491 , P1_R1192_U52 );
nand NAND2_15604 ( P1_R1192_U241 , P1_U3063 , P1_R1192_U50 );
nand NAND2_15605 ( P1_R1192_U242 , P1_U3062 , P1_R1192_U51 );
nand NAND2_15606 ( P1_R1192_U243 , P1_R1192_U189 , P1_R1192_U8 );
nand NAND2_15607 ( P1_R1192_U244 , P1_R1192_U9 , P1_R1192_U243 );
nand NAND2_15608 ( P1_R1192_U245 , P1_U3491 , P1_R1192_U52 );
nand NAND2_15609 ( P1_R1192_U246 , P1_R1192_U125 , P1_R1192_U148 );
nand NAND2_15610 ( P1_R1192_U247 , P1_R1192_U245 , P1_R1192_U244 );
not NOT1_15611 ( P1_R1192_U248 , P1_R1192_U173 );
nand NAND2_15612 ( P1_R1192_U249 , P1_U3494 , P1_R1192_U56 );
nand NAND2_15613 ( P1_R1192_U250 , P1_R1192_U249 , P1_R1192_U173 );
nand NAND2_15614 ( P1_R1192_U251 , P1_U3072 , P1_R1192_U55 );
not NOT1_15615 ( P1_R1192_U252 , P1_R1192_U172 );
nand NAND2_15616 ( P1_R1192_U253 , P1_U3497 , P1_R1192_U58 );
nand NAND2_15617 ( P1_R1192_U254 , P1_R1192_U253 , P1_R1192_U172 );
nand NAND2_15618 ( P1_R1192_U255 , P1_U3080 , P1_R1192_U57 );
not NOT1_15619 ( P1_R1192_U256 , P1_R1192_U171 );
nand NAND2_15620 ( P1_R1192_U257 , P1_U3506 , P1_R1192_U61 );
nand NAND2_15621 ( P1_R1192_U258 , P1_U3073 , P1_R1192_U59 );
nand NAND2_15622 ( P1_R1192_U259 , P1_U3074 , P1_R1192_U49 );
nand NAND2_15623 ( P1_R1192_U260 , P1_R1192_U186 , P1_R1192_U180 );
nand NAND2_15624 ( P1_R1192_U261 , P1_R1192_U10 , P1_R1192_U260 );
nand NAND2_15625 ( P1_R1192_U262 , P1_U3500 , P1_R1192_U63 );
nand NAND2_15626 ( P1_R1192_U263 , P1_U3506 , P1_R1192_U61 );
nand NAND3_15627 ( P1_R1192_U264 , P1_R1192_U171 , P1_R1192_U126 , P1_R1192_U257 );
nand NAND2_15628 ( P1_R1192_U265 , P1_R1192_U263 , P1_R1192_U261 );
not NOT1_15629 ( P1_R1192_U266 , P1_R1192_U168 );
nand NAND2_15630 ( P1_R1192_U267 , P1_U3509 , P1_R1192_U66 );
nand NAND2_15631 ( P1_R1192_U268 , P1_R1192_U267 , P1_R1192_U168 );
nand NAND2_15632 ( P1_R1192_U269 , P1_U3069 , P1_R1192_U65 );
not NOT1_15633 ( P1_R1192_U270 , P1_R1192_U67 );
nand NAND2_15634 ( P1_R1192_U271 , P1_R1192_U270 , P1_R1192_U68 );
nand NAND2_15635 ( P1_R1192_U272 , P1_R1192_U271 , P1_R1192_U167 );
nand NAND2_15636 ( P1_R1192_U273 , P1_U3082 , P1_R1192_U67 );
not NOT1_15637 ( P1_R1192_U274 , P1_R1192_U166 );
nand NAND2_15638 ( P1_R1192_U275 , P1_U3514 , P1_R1192_U70 );
nand NAND2_15639 ( P1_R1192_U276 , P1_R1192_U275 , P1_R1192_U166 );
nand NAND2_15640 ( P1_R1192_U277 , P1_U3081 , P1_R1192_U69 );
not NOT1_15641 ( P1_R1192_U278 , P1_R1192_U164 );
nand NAND2_15642 ( P1_R1192_U279 , P1_U4025 , P1_R1192_U72 );
nand NAND2_15643 ( P1_R1192_U280 , P1_R1192_U279 , P1_R1192_U164 );
nand NAND2_15644 ( P1_R1192_U281 , P1_U3076 , P1_R1192_U71 );
not NOT1_15645 ( P1_R1192_U282 , P1_R1192_U163 );
nand NAND2_15646 ( P1_R1192_U283 , P1_U4022 , P1_R1192_U75 );
nand NAND2_15647 ( P1_R1192_U284 , P1_U3066 , P1_R1192_U73 );
nand NAND2_15648 ( P1_R1192_U285 , P1_U3061 , P1_R1192_U48 );
nand NAND2_15649 ( P1_R1192_U286 , P1_R1192_U187 , P1_R1192_U181 );
nand NAND2_15650 ( P1_R1192_U287 , P1_R1192_U11 , P1_R1192_U286 );
nand NAND2_15651 ( P1_R1192_U288 , P1_U4024 , P1_R1192_U77 );
nand NAND2_15652 ( P1_R1192_U289 , P1_U4022 , P1_R1192_U75 );
nand NAND3_15653 ( P1_R1192_U290 , P1_R1192_U163 , P1_R1192_U127 , P1_R1192_U283 );
nand NAND2_15654 ( P1_R1192_U291 , P1_R1192_U289 , P1_R1192_U287 );
not NOT1_15655 ( P1_R1192_U292 , P1_R1192_U160 );
nand NAND2_15656 ( P1_R1192_U293 , P1_U4021 , P1_R1192_U80 );
nand NAND2_15657 ( P1_R1192_U294 , P1_R1192_U293 , P1_R1192_U160 );
nand NAND2_15658 ( P1_R1192_U295 , P1_U3065 , P1_R1192_U79 );
not NOT1_15659 ( P1_R1192_U296 , P1_R1192_U159 );
nand NAND2_15660 ( P1_R1192_U297 , P1_U4020 , P1_R1192_U82 );
nand NAND2_15661 ( P1_R1192_U298 , P1_R1192_U297 , P1_R1192_U159 );
nand NAND2_15662 ( P1_R1192_U299 , P1_U3058 , P1_R1192_U81 );
not NOT1_15663 ( P1_R1192_U300 , P1_R1192_U89 );
nand NAND2_15664 ( P1_R1192_U301 , P1_U4018 , P1_R1192_U86 );
nand NAND3_15665 ( P1_R1192_U302 , P1_R1192_U89 , P1_R1192_U182 , P1_R1192_U301 );
nand NAND2_15666 ( P1_R1192_U303 , P1_R1192_U86 , P1_R1192_U85 );
nand NAND2_15667 ( P1_R1192_U304 , P1_R1192_U303 , P1_R1192_U83 );
nand NAND2_15668 ( P1_R1192_U305 , P1_U3053 , P1_R1192_U176 );
not NOT1_15669 ( P1_R1192_U306 , P1_R1192_U157 );
nand NAND2_15670 ( P1_R1192_U307 , P1_U4017 , P1_R1192_U88 );
nand NAND2_15671 ( P1_R1192_U308 , P1_U3054 , P1_R1192_U87 );
nand NAND2_15672 ( P1_R1192_U309 , P1_R1192_U300 , P1_R1192_U85 );
nand NAND2_15673 ( P1_R1192_U310 , P1_R1192_U133 , P1_R1192_U309 );
nand NAND2_15674 ( P1_R1192_U311 , P1_R1192_U89 , P1_R1192_U182 );
nand NAND2_15675 ( P1_R1192_U312 , P1_R1192_U132 , P1_R1192_U311 );
nand NAND2_15676 ( P1_R1192_U313 , P1_R1192_U85 , P1_R1192_U182 );
nand NAND2_15677 ( P1_R1192_U314 , P1_R1192_U288 , P1_R1192_U163 );
not NOT1_15678 ( P1_R1192_U315 , P1_R1192_U90 );
nand NAND2_15679 ( P1_R1192_U316 , P1_U3061 , P1_R1192_U48 );
nand NAND2_15680 ( P1_R1192_U317 , P1_R1192_U315 , P1_R1192_U316 );
nand NAND2_15681 ( P1_R1192_U318 , P1_R1192_U136 , P1_R1192_U317 );
nand NAND2_15682 ( P1_R1192_U319 , P1_R1192_U90 , P1_R1192_U181 );
nand NAND2_15683 ( P1_R1192_U320 , P1_U4022 , P1_R1192_U75 );
nand NAND3_15684 ( P1_R1192_U321 , P1_R1192_U320 , P1_R1192_U319 , P1_R1192_U11 );
nand NAND2_15685 ( P1_R1192_U322 , P1_U3061 , P1_R1192_U48 );
nand NAND2_15686 ( P1_R1192_U323 , P1_R1192_U181 , P1_R1192_U322 );
nand NAND2_15687 ( P1_R1192_U324 , P1_R1192_U288 , P1_R1192_U78 );
nand NAND2_15688 ( P1_R1192_U325 , P1_R1192_U262 , P1_R1192_U171 );
not NOT1_15689 ( P1_R1192_U326 , P1_R1192_U91 );
nand NAND2_15690 ( P1_R1192_U327 , P1_U3074 , P1_R1192_U49 );
nand NAND2_15691 ( P1_R1192_U328 , P1_R1192_U326 , P1_R1192_U327 );
nand NAND2_15692 ( P1_R1192_U329 , P1_R1192_U142 , P1_R1192_U328 );
nand NAND2_15693 ( P1_R1192_U330 , P1_R1192_U91 , P1_R1192_U180 );
nand NAND2_15694 ( P1_R1192_U331 , P1_U3506 , P1_R1192_U61 );
nand NAND3_15695 ( P1_R1192_U332 , P1_R1192_U331 , P1_R1192_U330 , P1_R1192_U10 );
nand NAND2_15696 ( P1_R1192_U333 , P1_U3074 , P1_R1192_U49 );
nand NAND2_15697 ( P1_R1192_U334 , P1_R1192_U180 , P1_R1192_U333 );
nand NAND2_15698 ( P1_R1192_U335 , P1_R1192_U262 , P1_R1192_U64 );
nand NAND2_15699 ( P1_R1192_U336 , P1_R1192_U217 , P1_R1192_U148 );
not NOT1_15700 ( P1_R1192_U337 , P1_R1192_U92 );
nand NAND2_15701 ( P1_R1192_U338 , P1_U3062 , P1_R1192_U51 );
nand NAND2_15702 ( P1_R1192_U339 , P1_R1192_U337 , P1_R1192_U338 );
nand NAND2_15703 ( P1_R1192_U340 , P1_R1192_U146 , P1_R1192_U339 );
nand NAND2_15704 ( P1_R1192_U341 , P1_R1192_U92 , P1_R1192_U179 );
nand NAND2_15705 ( P1_R1192_U342 , P1_U3491 , P1_R1192_U52 );
nand NAND2_15706 ( P1_R1192_U343 , P1_R1192_U145 , P1_R1192_U341 );
nand NAND2_15707 ( P1_R1192_U344 , P1_U3062 , P1_R1192_U51 );
nand NAND2_15708 ( P1_R1192_U345 , P1_R1192_U179 , P1_R1192_U344 );
nand NAND2_15709 ( P1_R1192_U346 , P1_U3077 , P1_R1192_U24 );
nand NAND3_15710 ( P1_R1192_U347 , P1_R1192_U89 , P1_R1192_U182 , P1_R1192_U301 );
nand NAND3_15711 ( P1_R1192_U348 , P1_R1192_U12 , P1_R1192_U347 , P1_R1192_U130 );
nand NAND2_15712 ( P1_R1192_U349 , P1_U3485 , P1_R1192_U43 );
nand NAND2_15713 ( P1_R1192_U350 , P1_U3083 , P1_R1192_U42 );
nand NAND2_15714 ( P1_R1192_U351 , P1_R1192_U218 , P1_R1192_U148 );
nand NAND2_15715 ( P1_R1192_U352 , P1_R1192_U216 , P1_R1192_U147 );
nand NAND2_15716 ( P1_R1192_U353 , P1_U3482 , P1_R1192_U41 );
nand NAND2_15717 ( P1_R1192_U354 , P1_U3084 , P1_R1192_U38 );
nand NAND2_15718 ( P1_R1192_U355 , P1_U3482 , P1_R1192_U41 );
nand NAND2_15719 ( P1_R1192_U356 , P1_U3084 , P1_R1192_U38 );
nand NAND2_15720 ( P1_R1192_U357 , P1_R1192_U356 , P1_R1192_U355 );
nand NAND2_15721 ( P1_R1192_U358 , P1_U3479 , P1_R1192_U39 );
nand NAND2_15722 ( P1_R1192_U359 , P1_U3070 , P1_R1192_U22 );
nand NAND2_15723 ( P1_R1192_U360 , P1_R1192_U223 , P1_R1192_U44 );
nand NAND2_15724 ( P1_R1192_U361 , P1_R1192_U149 , P1_R1192_U210 );
nand NAND2_15725 ( P1_R1192_U362 , P1_U3476 , P1_R1192_U34 );
nand NAND2_15726 ( P1_R1192_U363 , P1_U3071 , P1_R1192_U31 );
nand NAND2_15727 ( P1_R1192_U364 , P1_R1192_U363 , P1_R1192_U362 );
nand NAND2_15728 ( P1_R1192_U365 , P1_U3473 , P1_R1192_U35 );
nand NAND2_15729 ( P1_R1192_U366 , P1_U3067 , P1_R1192_U32 );
nand NAND2_15730 ( P1_R1192_U367 , P1_R1192_U233 , P1_R1192_U45 );
nand NAND2_15731 ( P1_R1192_U368 , P1_R1192_U150 , P1_R1192_U225 );
nand NAND2_15732 ( P1_R1192_U369 , P1_U3470 , P1_R1192_U36 );
nand NAND2_15733 ( P1_R1192_U370 , P1_U3060 , P1_R1192_U33 );
nand NAND2_15734 ( P1_R1192_U371 , P1_R1192_U234 , P1_R1192_U152 );
nand NAND2_15735 ( P1_R1192_U372 , P1_R1192_U200 , P1_R1192_U151 );
nand NAND2_15736 ( P1_R1192_U373 , P1_U3467 , P1_R1192_U30 );
nand NAND2_15737 ( P1_R1192_U374 , P1_U3064 , P1_R1192_U27 );
nand NAND2_15738 ( P1_R1192_U375 , P1_U3467 , P1_R1192_U30 );
nand NAND2_15739 ( P1_R1192_U376 , P1_U3064 , P1_R1192_U27 );
nand NAND2_15740 ( P1_R1192_U377 , P1_R1192_U376 , P1_R1192_U375 );
nand NAND2_15741 ( P1_R1192_U378 , P1_U3464 , P1_R1192_U28 );
nand NAND2_15742 ( P1_R1192_U379 , P1_U3068 , P1_R1192_U23 );
nand NAND2_15743 ( P1_R1192_U380 , P1_R1192_U239 , P1_R1192_U46 );
nand NAND2_15744 ( P1_R1192_U381 , P1_R1192_U153 , P1_R1192_U194 );
nand NAND2_15745 ( P1_R1192_U382 , P1_U4028 , P1_R1192_U155 );
nand NAND2_15746 ( P1_R1192_U383 , P1_U3055 , P1_R1192_U154 );
nand NAND2_15747 ( P1_R1192_U384 , P1_U4028 , P1_R1192_U155 );
nand NAND2_15748 ( P1_R1192_U385 , P1_U3055 , P1_R1192_U154 );
nand NAND2_15749 ( P1_R1192_U386 , P1_R1192_U385 , P1_R1192_U384 );
nand NAND3_15750 ( P1_R1192_U387 , P1_U3054 , P1_R1192_U386 , P1_R1192_U87 );
nand NAND3_15751 ( P1_R1192_U388 , P1_R1192_U12 , P1_R1192_U88 , P1_U4017 );
nand NAND2_15752 ( P1_R1192_U389 , P1_U4017 , P1_R1192_U88 );
nand NAND2_15753 ( P1_R1192_U390 , P1_U3054 , P1_R1192_U87 );
not NOT1_15754 ( P1_R1192_U391 , P1_R1192_U131 );
nand NAND2_15755 ( P1_R1192_U392 , P1_R1192_U306 , P1_R1192_U391 );
nand NAND2_15756 ( P1_R1192_U393 , P1_R1192_U131 , P1_R1192_U157 );
nand NAND2_15757 ( P1_R1192_U394 , P1_U4018 , P1_R1192_U86 );
nand NAND2_15758 ( P1_R1192_U395 , P1_U3053 , P1_R1192_U83 );
nand NAND2_15759 ( P1_R1192_U396 , P1_U4018 , P1_R1192_U86 );
nand NAND2_15760 ( P1_R1192_U397 , P1_U3053 , P1_R1192_U83 );
nand NAND2_15761 ( P1_R1192_U398 , P1_R1192_U397 , P1_R1192_U396 );
nand NAND2_15762 ( P1_R1192_U399 , P1_U4019 , P1_R1192_U84 );
nand NAND2_15763 ( P1_R1192_U400 , P1_U3057 , P1_R1192_U47 );
nand NAND2_15764 ( P1_R1192_U401 , P1_R1192_U313 , P1_R1192_U89 );
nand NAND2_15765 ( P1_R1192_U402 , P1_R1192_U158 , P1_R1192_U300 );
nand NAND2_15766 ( P1_R1192_U403 , P1_U4020 , P1_R1192_U82 );
nand NAND2_15767 ( P1_R1192_U404 , P1_U3058 , P1_R1192_U81 );
not NOT1_15768 ( P1_R1192_U405 , P1_R1192_U134 );
nand NAND2_15769 ( P1_R1192_U406 , P1_R1192_U296 , P1_R1192_U405 );
nand NAND2_15770 ( P1_R1192_U407 , P1_R1192_U134 , P1_R1192_U159 );
nand NAND2_15771 ( P1_R1192_U408 , P1_U4021 , P1_R1192_U80 );
nand NAND2_15772 ( P1_R1192_U409 , P1_U3065 , P1_R1192_U79 );
not NOT1_15773 ( P1_R1192_U410 , P1_R1192_U135 );
nand NAND2_15774 ( P1_R1192_U411 , P1_R1192_U292 , P1_R1192_U410 );
nand NAND2_15775 ( P1_R1192_U412 , P1_R1192_U135 , P1_R1192_U160 );
nand NAND2_15776 ( P1_R1192_U413 , P1_U4022 , P1_R1192_U75 );
nand NAND2_15777 ( P1_R1192_U414 , P1_U3066 , P1_R1192_U73 );
nand NAND2_15778 ( P1_R1192_U415 , P1_R1192_U414 , P1_R1192_U413 );
nand NAND2_15779 ( P1_R1192_U416 , P1_U4023 , P1_R1192_U76 );
nand NAND2_15780 ( P1_R1192_U417 , P1_U3061 , P1_R1192_U48 );
nand NAND2_15781 ( P1_R1192_U418 , P1_R1192_U323 , P1_R1192_U90 );
nand NAND2_15782 ( P1_R1192_U419 , P1_R1192_U161 , P1_R1192_U315 );
nand NAND2_15783 ( P1_R1192_U420 , P1_U4024 , P1_R1192_U77 );
nand NAND2_15784 ( P1_R1192_U421 , P1_U3075 , P1_R1192_U74 );
nand NAND2_15785 ( P1_R1192_U422 , P1_R1192_U324 , P1_R1192_U163 );
nand NAND2_15786 ( P1_R1192_U423 , P1_R1192_U282 , P1_R1192_U162 );
nand NAND2_15787 ( P1_R1192_U424 , P1_U4025 , P1_R1192_U72 );
nand NAND2_15788 ( P1_R1192_U425 , P1_U3076 , P1_R1192_U71 );
not NOT1_15789 ( P1_R1192_U426 , P1_R1192_U137 );
nand NAND2_15790 ( P1_R1192_U427 , P1_R1192_U278 , P1_R1192_U426 );
nand NAND2_15791 ( P1_R1192_U428 , P1_R1192_U137 , P1_R1192_U164 );
nand NAND2_15792 ( P1_R1192_U429 , P1_U3461 , P1_R1192_U26 );
nand NAND2_15793 ( P1_R1192_U430 , P1_U3078 , P1_R1192_U165 );
not NOT1_15794 ( P1_R1192_U431 , P1_R1192_U138 );
nand NAND2_15795 ( P1_R1192_U432 , P1_R1192_U431 , P1_R1192_U190 );
nand NAND2_15796 ( P1_R1192_U433 , P1_R1192_U138 , P1_R1192_U25 );
nand NAND2_15797 ( P1_R1192_U434 , P1_U3514 , P1_R1192_U70 );
nand NAND2_15798 ( P1_R1192_U435 , P1_U3081 , P1_R1192_U69 );
not NOT1_15799 ( P1_R1192_U436 , P1_R1192_U139 );
nand NAND2_15800 ( P1_R1192_U437 , P1_R1192_U274 , P1_R1192_U436 );
nand NAND2_15801 ( P1_R1192_U438 , P1_R1192_U139 , P1_R1192_U166 );
nand NAND2_15802 ( P1_R1192_U439 , P1_U3512 , P1_R1192_U68 );
nand NAND2_15803 ( P1_R1192_U440 , P1_U3082 , P1_R1192_U167 );
not NOT1_15804 ( P1_R1192_U441 , P1_R1192_U140 );
nand NAND2_15805 ( P1_R1192_U442 , P1_R1192_U441 , P1_R1192_U270 );
nand NAND2_15806 ( P1_R1192_U443 , P1_R1192_U140 , P1_R1192_U67 );
nand NAND2_15807 ( P1_R1192_U444 , P1_U3509 , P1_R1192_U66 );
nand NAND2_15808 ( P1_R1192_U445 , P1_U3069 , P1_R1192_U65 );
not NOT1_15809 ( P1_R1192_U446 , P1_R1192_U141 );
nand NAND2_15810 ( P1_R1192_U447 , P1_R1192_U266 , P1_R1192_U446 );
nand NAND2_15811 ( P1_R1192_U448 , P1_R1192_U141 , P1_R1192_U168 );
nand NAND2_15812 ( P1_R1192_U449 , P1_U3506 , P1_R1192_U61 );
nand NAND2_15813 ( P1_R1192_U450 , P1_U3073 , P1_R1192_U59 );
nand NAND2_15814 ( P1_R1192_U451 , P1_R1192_U450 , P1_R1192_U449 );
nand NAND2_15815 ( P1_R1192_U452 , P1_U3503 , P1_R1192_U62 );
nand NAND2_15816 ( P1_R1192_U453 , P1_U3074 , P1_R1192_U49 );
nand NAND2_15817 ( P1_R1192_U454 , P1_R1192_U334 , P1_R1192_U91 );
nand NAND2_15818 ( P1_R1192_U455 , P1_R1192_U169 , P1_R1192_U326 );
nand NAND2_15819 ( P1_R1192_U456 , P1_U3500 , P1_R1192_U63 );
nand NAND2_15820 ( P1_R1192_U457 , P1_U3079 , P1_R1192_U60 );
nand NAND2_15821 ( P1_R1192_U458 , P1_R1192_U335 , P1_R1192_U171 );
nand NAND2_15822 ( P1_R1192_U459 , P1_R1192_U256 , P1_R1192_U170 );
nand NAND2_15823 ( P1_R1192_U460 , P1_U3497 , P1_R1192_U58 );
nand NAND2_15824 ( P1_R1192_U461 , P1_U3080 , P1_R1192_U57 );
not NOT1_15825 ( P1_R1192_U462 , P1_R1192_U143 );
nand NAND2_15826 ( P1_R1192_U463 , P1_R1192_U252 , P1_R1192_U462 );
nand NAND2_15827 ( P1_R1192_U464 , P1_R1192_U143 , P1_R1192_U172 );
nand NAND2_15828 ( P1_R1192_U465 , P1_U3494 , P1_R1192_U56 );
nand NAND2_15829 ( P1_R1192_U466 , P1_U3072 , P1_R1192_U55 );
not NOT1_15830 ( P1_R1192_U467 , P1_R1192_U144 );
nand NAND2_15831 ( P1_R1192_U468 , P1_R1192_U248 , P1_R1192_U467 );
nand NAND2_15832 ( P1_R1192_U469 , P1_R1192_U144 , P1_R1192_U173 );
nand NAND2_15833 ( P1_R1192_U470 , P1_U3491 , P1_R1192_U52 );
nand NAND2_15834 ( P1_R1192_U471 , P1_U3063 , P1_R1192_U50 );
nand NAND2_15835 ( P1_R1192_U472 , P1_R1192_U471 , P1_R1192_U470 );
nand NAND2_15836 ( P1_R1192_U473 , P1_U3488 , P1_R1192_U53 );
nand NAND2_15837 ( P1_R1192_U474 , P1_U3062 , P1_R1192_U51 );
nand NAND2_15838 ( P1_R1192_U475 , P1_R1192_U345 , P1_R1192_U92 );
nand NAND2_15839 ( P1_R1192_U476 , P1_R1192_U174 , P1_R1192_U337 );
and AND2_15840 ( P1_R1171_U4 , P1_R1171_U176 , P1_R1171_U175 );
and AND2_15841 ( P1_R1171_U5 , P1_R1171_U177 , P1_R1171_U178 );
and AND2_15842 ( P1_R1171_U6 , P1_R1171_U194 , P1_R1171_U193 );
and AND2_15843 ( P1_R1171_U7 , P1_R1171_U234 , P1_R1171_U233 );
and AND2_15844 ( P1_R1171_U8 , P1_R1171_U243 , P1_R1171_U242 );
and AND2_15845 ( P1_R1171_U9 , P1_R1171_U261 , P1_R1171_U260 );
and AND2_15846 ( P1_R1171_U10 , P1_R1171_U269 , P1_R1171_U268 );
and AND2_15847 ( P1_R1171_U11 , P1_R1171_U348 , P1_R1171_U345 );
and AND2_15848 ( P1_R1171_U12 , P1_R1171_U341 , P1_R1171_U338 );
and AND2_15849 ( P1_R1171_U13 , P1_R1171_U332 , P1_R1171_U329 );
and AND2_15850 ( P1_R1171_U14 , P1_R1171_U323 , P1_R1171_U320 );
and AND2_15851 ( P1_R1171_U15 , P1_R1171_U317 , P1_R1171_U315 );
and AND2_15852 ( P1_R1171_U16 , P1_R1171_U310 , P1_R1171_U307 );
and AND2_15853 ( P1_R1171_U17 , P1_R1171_U232 , P1_R1171_U229 );
and AND2_15854 ( P1_R1171_U18 , P1_R1171_U224 , P1_R1171_U221 );
and AND2_15855 ( P1_R1171_U19 , P1_R1171_U210 , P1_R1171_U207 );
not NOT1_15856 ( P1_R1171_U20 , P1_U3476 );
not NOT1_15857 ( P1_R1171_U21 , P1_U3071 );
not NOT1_15858 ( P1_R1171_U22 , P1_U3070 );
nand NAND2_15859 ( P1_R1171_U23 , P1_U3071 , P1_U3476 );
not NOT1_15860 ( P1_R1171_U24 , P1_U3479 );
not NOT1_15861 ( P1_R1171_U25 , P1_U3470 );
not NOT1_15862 ( P1_R1171_U26 , P1_U3060 );
not NOT1_15863 ( P1_R1171_U27 , P1_U3067 );
not NOT1_15864 ( P1_R1171_U28 , P1_U3464 );
not NOT1_15865 ( P1_R1171_U29 , P1_U3068 );
not NOT1_15866 ( P1_R1171_U30 , P1_U3456 );
not NOT1_15867 ( P1_R1171_U31 , P1_U3077 );
nand NAND2_15868 ( P1_R1171_U32 , P1_U3077 , P1_U3456 );
not NOT1_15869 ( P1_R1171_U33 , P1_U3467 );
not NOT1_15870 ( P1_R1171_U34 , P1_U3064 );
nand NAND2_15871 ( P1_R1171_U35 , P1_U3060 , P1_U3470 );
not NOT1_15872 ( P1_R1171_U36 , P1_U3473 );
not NOT1_15873 ( P1_R1171_U37 , P1_U3482 );
not NOT1_15874 ( P1_R1171_U38 , P1_U3084 );
not NOT1_15875 ( P1_R1171_U39 , P1_U3083 );
not NOT1_15876 ( P1_R1171_U40 , P1_U3485 );
nand NAND2_15877 ( P1_R1171_U41 , P1_R1171_U62 , P1_R1171_U202 );
nand NAND2_15878 ( P1_R1171_U42 , P1_R1171_U118 , P1_R1171_U190 );
nand NAND2_15879 ( P1_R1171_U43 , P1_R1171_U179 , P1_R1171_U180 );
nand NAND2_15880 ( P1_R1171_U44 , P1_U3461 , P1_U3078 );
nand NAND2_15881 ( P1_R1171_U45 , P1_R1171_U122 , P1_R1171_U216 );
nand NAND2_15882 ( P1_R1171_U46 , P1_R1171_U213 , P1_R1171_U212 );
not NOT1_15883 ( P1_R1171_U47 , P1_U4018 );
not NOT1_15884 ( P1_R1171_U48 , P1_U3053 );
not NOT1_15885 ( P1_R1171_U49 , P1_U3057 );
not NOT1_15886 ( P1_R1171_U50 , P1_U4019 );
not NOT1_15887 ( P1_R1171_U51 , P1_U4020 );
not NOT1_15888 ( P1_R1171_U52 , P1_U3058 );
not NOT1_15889 ( P1_R1171_U53 , P1_U4021 );
not NOT1_15890 ( P1_R1171_U54 , P1_U3065 );
not NOT1_15891 ( P1_R1171_U55 , P1_U4024 );
not NOT1_15892 ( P1_R1171_U56 , P1_U3075 );
not NOT1_15893 ( P1_R1171_U57 , P1_U3506 );
not NOT1_15894 ( P1_R1171_U58 , P1_U3073 );
not NOT1_15895 ( P1_R1171_U59 , P1_U3069 );
nand NAND2_15896 ( P1_R1171_U60 , P1_U3073 , P1_U3506 );
not NOT1_15897 ( P1_R1171_U61 , P1_U3509 );
nand NAND2_15898 ( P1_R1171_U62 , P1_U3084 , P1_U3482 );
not NOT1_15899 ( P1_R1171_U63 , P1_U3488 );
not NOT1_15900 ( P1_R1171_U64 , P1_U3062 );
not NOT1_15901 ( P1_R1171_U65 , P1_U3494 );
not NOT1_15902 ( P1_R1171_U66 , P1_U3072 );
not NOT1_15903 ( P1_R1171_U67 , P1_U3491 );
not NOT1_15904 ( P1_R1171_U68 , P1_U3063 );
nand NAND2_15905 ( P1_R1171_U69 , P1_U3063 , P1_U3491 );
not NOT1_15906 ( P1_R1171_U70 , P1_U3497 );
not NOT1_15907 ( P1_R1171_U71 , P1_U3080 );
not NOT1_15908 ( P1_R1171_U72 , P1_U3500 );
not NOT1_15909 ( P1_R1171_U73 , P1_U3079 );
not NOT1_15910 ( P1_R1171_U74 , P1_U3503 );
not NOT1_15911 ( P1_R1171_U75 , P1_U3074 );
not NOT1_15912 ( P1_R1171_U76 , P1_U3512 );
not NOT1_15913 ( P1_R1171_U77 , P1_U3082 );
nand NAND2_15914 ( P1_R1171_U78 , P1_U3082 , P1_U3512 );
not NOT1_15915 ( P1_R1171_U79 , P1_U3514 );
not NOT1_15916 ( P1_R1171_U80 , P1_U3081 );
nand NAND2_15917 ( P1_R1171_U81 , P1_U3081 , P1_U3514 );
not NOT1_15918 ( P1_R1171_U82 , P1_U4025 );
not NOT1_15919 ( P1_R1171_U83 , P1_U4023 );
not NOT1_15920 ( P1_R1171_U84 , P1_U3061 );
not NOT1_15921 ( P1_R1171_U85 , P1_U4022 );
not NOT1_15922 ( P1_R1171_U86 , P1_U3066 );
nand NAND2_15923 ( P1_R1171_U87 , P1_U4019 , P1_U3057 );
not NOT1_15924 ( P1_R1171_U88 , P1_U3054 );
not NOT1_15925 ( P1_R1171_U89 , P1_U4017 );
nand NAND2_15926 ( P1_R1171_U90 , P1_R1171_U303 , P1_R1171_U173 );
not NOT1_15927 ( P1_R1171_U91 , P1_U3076 );
nand NAND2_15928 ( P1_R1171_U92 , P1_R1171_U78 , P1_R1171_U312 );
nand NAND2_15929 ( P1_R1171_U93 , P1_R1171_U258 , P1_R1171_U257 );
nand NAND2_15930 ( P1_R1171_U94 , P1_R1171_U69 , P1_R1171_U334 );
nand NAND2_15931 ( P1_R1171_U95 , P1_R1171_U454 , P1_R1171_U453 );
nand NAND2_15932 ( P1_R1171_U96 , P1_R1171_U501 , P1_R1171_U500 );
nand NAND2_15933 ( P1_R1171_U97 , P1_R1171_U372 , P1_R1171_U371 );
nand NAND2_15934 ( P1_R1171_U98 , P1_R1171_U377 , P1_R1171_U376 );
nand NAND2_15935 ( P1_R1171_U99 , P1_R1171_U384 , P1_R1171_U383 );
nand NAND2_15936 ( P1_R1171_U100 , P1_R1171_U391 , P1_R1171_U390 );
nand NAND2_15937 ( P1_R1171_U101 , P1_R1171_U396 , P1_R1171_U395 );
nand NAND2_15938 ( P1_R1171_U102 , P1_R1171_U405 , P1_R1171_U404 );
nand NAND2_15939 ( P1_R1171_U103 , P1_R1171_U412 , P1_R1171_U411 );
nand NAND2_15940 ( P1_R1171_U104 , P1_R1171_U419 , P1_R1171_U418 );
nand NAND2_15941 ( P1_R1171_U105 , P1_R1171_U426 , P1_R1171_U425 );
nand NAND2_15942 ( P1_R1171_U106 , P1_R1171_U431 , P1_R1171_U430 );
nand NAND2_15943 ( P1_R1171_U107 , P1_R1171_U438 , P1_R1171_U437 );
nand NAND2_15944 ( P1_R1171_U108 , P1_R1171_U445 , P1_R1171_U444 );
nand NAND2_15945 ( P1_R1171_U109 , P1_R1171_U459 , P1_R1171_U458 );
nand NAND2_15946 ( P1_R1171_U110 , P1_R1171_U464 , P1_R1171_U463 );
nand NAND2_15947 ( P1_R1171_U111 , P1_R1171_U471 , P1_R1171_U470 );
nand NAND2_15948 ( P1_R1171_U112 , P1_R1171_U478 , P1_R1171_U477 );
nand NAND2_15949 ( P1_R1171_U113 , P1_R1171_U485 , P1_R1171_U484 );
nand NAND2_15950 ( P1_R1171_U114 , P1_R1171_U492 , P1_R1171_U491 );
nand NAND2_15951 ( P1_R1171_U115 , P1_R1171_U497 , P1_R1171_U496 );
and AND2_15952 ( P1_R1171_U116 , P1_U3464 , P1_U3068 );
and AND2_15953 ( P1_R1171_U117 , P1_R1171_U186 , P1_R1171_U184 );
and AND2_15954 ( P1_R1171_U118 , P1_R1171_U191 , P1_R1171_U189 );
and AND2_15955 ( P1_R1171_U119 , P1_R1171_U198 , P1_R1171_U197 );
and AND3_15956 ( P1_R1171_U120 , P1_R1171_U379 , P1_R1171_U378 , P1_R1171_U23 );
and AND2_15957 ( P1_R1171_U121 , P1_R1171_U209 , P1_R1171_U6 );
and AND2_15958 ( P1_R1171_U122 , P1_R1171_U217 , P1_R1171_U215 );
and AND3_15959 ( P1_R1171_U123 , P1_R1171_U386 , P1_R1171_U385 , P1_R1171_U35 );
and AND2_15960 ( P1_R1171_U124 , P1_R1171_U223 , P1_R1171_U4 );
and AND2_15961 ( P1_R1171_U125 , P1_R1171_U231 , P1_R1171_U178 );
and AND2_15962 ( P1_R1171_U126 , P1_R1171_U201 , P1_R1171_U7 );
and AND2_15963 ( P1_R1171_U127 , P1_R1171_U236 , P1_R1171_U168 );
and AND2_15964 ( P1_R1171_U128 , P1_R1171_U245 , P1_R1171_U169 );
and AND2_15965 ( P1_R1171_U129 , P1_R1171_U265 , P1_R1171_U264 );
and AND2_15966 ( P1_R1171_U130 , P1_R1171_U10 , P1_R1171_U279 );
and AND2_15967 ( P1_R1171_U131 , P1_R1171_U282 , P1_R1171_U277 );
and AND2_15968 ( P1_R1171_U132 , P1_R1171_U298 , P1_R1171_U295 );
and AND2_15969 ( P1_R1171_U133 , P1_R1171_U365 , P1_R1171_U299 );
and AND2_15970 ( P1_R1171_U134 , P1_R1171_U156 , P1_R1171_U275 );
and AND3_15971 ( P1_R1171_U135 , P1_R1171_U466 , P1_R1171_U465 , P1_R1171_U60 );
and AND3_15972 ( P1_R1171_U136 , P1_R1171_U487 , P1_R1171_U486 , P1_R1171_U169 );
and AND2_15973 ( P1_R1171_U137 , P1_R1171_U340 , P1_R1171_U8 );
and AND3_15974 ( P1_R1171_U138 , P1_R1171_U499 , P1_R1171_U498 , P1_R1171_U168 );
and AND2_15975 ( P1_R1171_U139 , P1_R1171_U347 , P1_R1171_U7 );
nand NAND2_15976 ( P1_R1171_U140 , P1_R1171_U119 , P1_R1171_U199 );
nand NAND2_15977 ( P1_R1171_U141 , P1_R1171_U214 , P1_R1171_U226 );
not NOT1_15978 ( P1_R1171_U142 , P1_U3055 );
not NOT1_15979 ( P1_R1171_U143 , P1_U4028 );
and AND2_15980 ( P1_R1171_U144 , P1_R1171_U400 , P1_R1171_U399 );
nand NAND3_15981 ( P1_R1171_U145 , P1_R1171_U301 , P1_R1171_U166 , P1_R1171_U361 );
and AND2_15982 ( P1_R1171_U146 , P1_R1171_U407 , P1_R1171_U406 );
nand NAND3_15983 ( P1_R1171_U147 , P1_R1171_U367 , P1_R1171_U366 , P1_R1171_U133 );
and AND2_15984 ( P1_R1171_U148 , P1_R1171_U414 , P1_R1171_U413 );
nand NAND3_15985 ( P1_R1171_U149 , P1_R1171_U362 , P1_R1171_U296 , P1_R1171_U87 );
and AND2_15986 ( P1_R1171_U150 , P1_R1171_U421 , P1_R1171_U420 );
nand NAND2_15987 ( P1_R1171_U151 , P1_R1171_U290 , P1_R1171_U289 );
and AND2_15988 ( P1_R1171_U152 , P1_R1171_U433 , P1_R1171_U432 );
nand NAND2_15989 ( P1_R1171_U153 , P1_R1171_U286 , P1_R1171_U285 );
and AND2_15990 ( P1_R1171_U154 , P1_R1171_U440 , P1_R1171_U439 );
nand NAND2_15991 ( P1_R1171_U155 , P1_R1171_U131 , P1_R1171_U281 );
and AND2_15992 ( P1_R1171_U156 , P1_R1171_U447 , P1_R1171_U446 );
and AND2_15993 ( P1_R1171_U157 , P1_R1171_U452 , P1_R1171_U451 );
nand NAND2_15994 ( P1_R1171_U158 , P1_R1171_U44 , P1_R1171_U324 );
nand NAND2_15995 ( P1_R1171_U159 , P1_R1171_U129 , P1_R1171_U266 );
and AND2_15996 ( P1_R1171_U160 , P1_R1171_U473 , P1_R1171_U472 );
nand NAND2_15997 ( P1_R1171_U161 , P1_R1171_U254 , P1_R1171_U253 );
and AND2_15998 ( P1_R1171_U162 , P1_R1171_U480 , P1_R1171_U479 );
nand NAND2_15999 ( P1_R1171_U163 , P1_R1171_U250 , P1_R1171_U249 );
nand NAND2_16000 ( P1_R1171_U164 , P1_R1171_U240 , P1_R1171_U239 );
nand NAND2_16001 ( P1_R1171_U165 , P1_R1171_U364 , P1_R1171_U363 );
nand NAND2_16002 ( P1_R1171_U166 , P1_U3054 , P1_R1171_U147 );
not NOT1_16003 ( P1_R1171_U167 , P1_R1171_U35 );
nand NAND2_16004 ( P1_R1171_U168 , P1_U3485 , P1_U3083 );
nand NAND2_16005 ( P1_R1171_U169 , P1_U3072 , P1_U3494 );
nand NAND2_16006 ( P1_R1171_U170 , P1_U3058 , P1_U4020 );
not NOT1_16007 ( P1_R1171_U171 , P1_R1171_U69 );
not NOT1_16008 ( P1_R1171_U172 , P1_R1171_U78 );
nand NAND2_16009 ( P1_R1171_U173 , P1_U3065 , P1_U4021 );
not NOT1_16010 ( P1_R1171_U174 , P1_R1171_U62 );
or OR2_16011 ( P1_R1171_U175 , P1_U3067 , P1_U3473 );
or OR2_16012 ( P1_R1171_U176 , P1_U3060 , P1_U3470 );
or OR2_16013 ( P1_R1171_U177 , P1_U3467 , P1_U3064 );
or OR2_16014 ( P1_R1171_U178 , P1_U3464 , P1_U3068 );
not NOT1_16015 ( P1_R1171_U179 , P1_R1171_U32 );
or OR2_16016 ( P1_R1171_U180 , P1_U3461 , P1_U3078 );
not NOT1_16017 ( P1_R1171_U181 , P1_R1171_U43 );
not NOT1_16018 ( P1_R1171_U182 , P1_R1171_U44 );
nand NAND2_16019 ( P1_R1171_U183 , P1_R1171_U43 , P1_R1171_U44 );
nand NAND2_16020 ( P1_R1171_U184 , P1_R1171_U116 , P1_R1171_U177 );
nand NAND2_16021 ( P1_R1171_U185 , P1_R1171_U5 , P1_R1171_U183 );
nand NAND2_16022 ( P1_R1171_U186 , P1_U3064 , P1_U3467 );
nand NAND2_16023 ( P1_R1171_U187 , P1_R1171_U117 , P1_R1171_U185 );
nand NAND2_16024 ( P1_R1171_U188 , P1_R1171_U36 , P1_R1171_U35 );
nand NAND2_16025 ( P1_R1171_U189 , P1_U3067 , P1_R1171_U188 );
nand NAND2_16026 ( P1_R1171_U190 , P1_R1171_U4 , P1_R1171_U187 );
nand NAND2_16027 ( P1_R1171_U191 , P1_U3473 , P1_R1171_U167 );
not NOT1_16028 ( P1_R1171_U192 , P1_R1171_U42 );
or OR2_16029 ( P1_R1171_U193 , P1_U3070 , P1_U3479 );
or OR2_16030 ( P1_R1171_U194 , P1_U3071 , P1_U3476 );
not NOT1_16031 ( P1_R1171_U195 , P1_R1171_U23 );
nand NAND2_16032 ( P1_R1171_U196 , P1_R1171_U24 , P1_R1171_U23 );
nand NAND2_16033 ( P1_R1171_U197 , P1_U3070 , P1_R1171_U196 );
nand NAND2_16034 ( P1_R1171_U198 , P1_U3479 , P1_R1171_U195 );
nand NAND2_16035 ( P1_R1171_U199 , P1_R1171_U6 , P1_R1171_U42 );
not NOT1_16036 ( P1_R1171_U200 , P1_R1171_U140 );
or OR2_16037 ( P1_R1171_U201 , P1_U3482 , P1_U3084 );
nand NAND2_16038 ( P1_R1171_U202 , P1_R1171_U201 , P1_R1171_U140 );
not NOT1_16039 ( P1_R1171_U203 , P1_R1171_U41 );
or OR2_16040 ( P1_R1171_U204 , P1_U3083 , P1_U3485 );
or OR2_16041 ( P1_R1171_U205 , P1_U3476 , P1_U3071 );
nand NAND2_16042 ( P1_R1171_U206 , P1_R1171_U205 , P1_R1171_U42 );
nand NAND2_16043 ( P1_R1171_U207 , P1_R1171_U120 , P1_R1171_U206 );
nand NAND2_16044 ( P1_R1171_U208 , P1_R1171_U192 , P1_R1171_U23 );
nand NAND2_16045 ( P1_R1171_U209 , P1_U3479 , P1_U3070 );
nand NAND2_16046 ( P1_R1171_U210 , P1_R1171_U121 , P1_R1171_U208 );
or OR2_16047 ( P1_R1171_U211 , P1_U3071 , P1_U3476 );
nand NAND2_16048 ( P1_R1171_U212 , P1_R1171_U182 , P1_R1171_U178 );
nand NAND2_16049 ( P1_R1171_U213 , P1_U3068 , P1_U3464 );
not NOT1_16050 ( P1_R1171_U214 , P1_R1171_U46 );
nand NAND2_16051 ( P1_R1171_U215 , P1_R1171_U181 , P1_R1171_U5 );
nand NAND2_16052 ( P1_R1171_U216 , P1_R1171_U46 , P1_R1171_U177 );
nand NAND2_16053 ( P1_R1171_U217 , P1_U3064 , P1_U3467 );
not NOT1_16054 ( P1_R1171_U218 , P1_R1171_U45 );
or OR2_16055 ( P1_R1171_U219 , P1_U3470 , P1_U3060 );
nand NAND2_16056 ( P1_R1171_U220 , P1_R1171_U219 , P1_R1171_U45 );
nand NAND2_16057 ( P1_R1171_U221 , P1_R1171_U123 , P1_R1171_U220 );
nand NAND2_16058 ( P1_R1171_U222 , P1_R1171_U218 , P1_R1171_U35 );
nand NAND2_16059 ( P1_R1171_U223 , P1_U3473 , P1_U3067 );
nand NAND2_16060 ( P1_R1171_U224 , P1_R1171_U124 , P1_R1171_U222 );
or OR2_16061 ( P1_R1171_U225 , P1_U3060 , P1_U3470 );
nand NAND2_16062 ( P1_R1171_U226 , P1_R1171_U181 , P1_R1171_U178 );
not NOT1_16063 ( P1_R1171_U227 , P1_R1171_U141 );
nand NAND2_16064 ( P1_R1171_U228 , P1_U3064 , P1_U3467 );
nand NAND4_16065 ( P1_R1171_U229 , P1_R1171_U398 , P1_R1171_U397 , P1_R1171_U44 , P1_R1171_U43 );
nand NAND2_16066 ( P1_R1171_U230 , P1_R1171_U44 , P1_R1171_U43 );
nand NAND2_16067 ( P1_R1171_U231 , P1_U3068 , P1_U3464 );
nand NAND2_16068 ( P1_R1171_U232 , P1_R1171_U125 , P1_R1171_U230 );
or OR2_16069 ( P1_R1171_U233 , P1_U3083 , P1_U3485 );
or OR2_16070 ( P1_R1171_U234 , P1_U3062 , P1_U3488 );
nand NAND2_16071 ( P1_R1171_U235 , P1_R1171_U174 , P1_R1171_U7 );
nand NAND2_16072 ( P1_R1171_U236 , P1_U3062 , P1_U3488 );
nand NAND2_16073 ( P1_R1171_U237 , P1_R1171_U127 , P1_R1171_U235 );
or OR2_16074 ( P1_R1171_U238 , P1_U3488 , P1_U3062 );
nand NAND2_16075 ( P1_R1171_U239 , P1_R1171_U126 , P1_R1171_U140 );
nand NAND2_16076 ( P1_R1171_U240 , P1_R1171_U238 , P1_R1171_U237 );
not NOT1_16077 ( P1_R1171_U241 , P1_R1171_U164 );
or OR2_16078 ( P1_R1171_U242 , P1_U3080 , P1_U3497 );
or OR2_16079 ( P1_R1171_U243 , P1_U3072 , P1_U3494 );
nand NAND2_16080 ( P1_R1171_U244 , P1_R1171_U171 , P1_R1171_U8 );
nand NAND2_16081 ( P1_R1171_U245 , P1_U3080 , P1_U3497 );
nand NAND2_16082 ( P1_R1171_U246 , P1_R1171_U128 , P1_R1171_U244 );
or OR2_16083 ( P1_R1171_U247 , P1_U3491 , P1_U3063 );
or OR2_16084 ( P1_R1171_U248 , P1_U3497 , P1_U3080 );
nand NAND3_16085 ( P1_R1171_U249 , P1_R1171_U247 , P1_R1171_U164 , P1_R1171_U8 );
nand NAND2_16086 ( P1_R1171_U250 , P1_R1171_U248 , P1_R1171_U246 );
not NOT1_16087 ( P1_R1171_U251 , P1_R1171_U163 );
or OR2_16088 ( P1_R1171_U252 , P1_U3500 , P1_U3079 );
nand NAND2_16089 ( P1_R1171_U253 , P1_R1171_U252 , P1_R1171_U163 );
nand NAND2_16090 ( P1_R1171_U254 , P1_U3079 , P1_U3500 );
not NOT1_16091 ( P1_R1171_U255 , P1_R1171_U161 );
or OR2_16092 ( P1_R1171_U256 , P1_U3503 , P1_U3074 );
nand NAND2_16093 ( P1_R1171_U257 , P1_R1171_U256 , P1_R1171_U161 );
nand NAND2_16094 ( P1_R1171_U258 , P1_U3074 , P1_U3503 );
not NOT1_16095 ( P1_R1171_U259 , P1_R1171_U93 );
or OR2_16096 ( P1_R1171_U260 , P1_U3069 , P1_U3509 );
or OR2_16097 ( P1_R1171_U261 , P1_U3073 , P1_U3506 );
not NOT1_16098 ( P1_R1171_U262 , P1_R1171_U60 );
nand NAND2_16099 ( P1_R1171_U263 , P1_R1171_U61 , P1_R1171_U60 );
nand NAND2_16100 ( P1_R1171_U264 , P1_U3069 , P1_R1171_U263 );
nand NAND2_16101 ( P1_R1171_U265 , P1_U3509 , P1_R1171_U262 );
nand NAND2_16102 ( P1_R1171_U266 , P1_R1171_U9 , P1_R1171_U93 );
not NOT1_16103 ( P1_R1171_U267 , P1_R1171_U159 );
or OR2_16104 ( P1_R1171_U268 , P1_U3076 , P1_U4025 );
or OR2_16105 ( P1_R1171_U269 , P1_U3081 , P1_U3514 );
or OR2_16106 ( P1_R1171_U270 , P1_U3075 , P1_U4024 );
not NOT1_16107 ( P1_R1171_U271 , P1_R1171_U81 );
nand NAND2_16108 ( P1_R1171_U272 , P1_U4025 , P1_R1171_U271 );
nand NAND2_16109 ( P1_R1171_U273 , P1_R1171_U272 , P1_R1171_U91 );
nand NAND2_16110 ( P1_R1171_U274 , P1_R1171_U81 , P1_R1171_U82 );
nand NAND2_16111 ( P1_R1171_U275 , P1_R1171_U274 , P1_R1171_U273 );
nand NAND2_16112 ( P1_R1171_U276 , P1_R1171_U172 , P1_R1171_U10 );
nand NAND2_16113 ( P1_R1171_U277 , P1_U3075 , P1_U4024 );
nand NAND2_16114 ( P1_R1171_U278 , P1_R1171_U275 , P1_R1171_U276 );
or OR2_16115 ( P1_R1171_U279 , P1_U3512 , P1_U3082 );
or OR2_16116 ( P1_R1171_U280 , P1_U4024 , P1_U3075 );
nand NAND3_16117 ( P1_R1171_U281 , P1_R1171_U270 , P1_R1171_U159 , P1_R1171_U130 );
nand NAND2_16118 ( P1_R1171_U282 , P1_R1171_U280 , P1_R1171_U278 );
not NOT1_16119 ( P1_R1171_U283 , P1_R1171_U155 );
or OR2_16120 ( P1_R1171_U284 , P1_U4023 , P1_U3061 );
nand NAND2_16121 ( P1_R1171_U285 , P1_R1171_U284 , P1_R1171_U155 );
nand NAND2_16122 ( P1_R1171_U286 , P1_U3061 , P1_U4023 );
not NOT1_16123 ( P1_R1171_U287 , P1_R1171_U153 );
or OR2_16124 ( P1_R1171_U288 , P1_U4022 , P1_U3066 );
nand NAND2_16125 ( P1_R1171_U289 , P1_R1171_U288 , P1_R1171_U153 );
nand NAND2_16126 ( P1_R1171_U290 , P1_U3066 , P1_U4022 );
not NOT1_16127 ( P1_R1171_U291 , P1_R1171_U151 );
or OR2_16128 ( P1_R1171_U292 , P1_U3058 , P1_U4020 );
nand NAND2_16129 ( P1_R1171_U293 , P1_R1171_U173 , P1_R1171_U170 );
not NOT1_16130 ( P1_R1171_U294 , P1_R1171_U87 );
or OR2_16131 ( P1_R1171_U295 , P1_U4021 , P1_U3065 );
nand NAND3_16132 ( P1_R1171_U296 , P1_R1171_U151 , P1_R1171_U295 , P1_R1171_U165 );
not NOT1_16133 ( P1_R1171_U297 , P1_R1171_U149 );
or OR2_16134 ( P1_R1171_U298 , P1_U4018 , P1_U3053 );
nand NAND2_16135 ( P1_R1171_U299 , P1_U3053 , P1_U4018 );
not NOT1_16136 ( P1_R1171_U300 , P1_R1171_U147 );
nand NAND2_16137 ( P1_R1171_U301 , P1_U4017 , P1_R1171_U147 );
not NOT1_16138 ( P1_R1171_U302 , P1_R1171_U145 );
nand NAND2_16139 ( P1_R1171_U303 , P1_R1171_U295 , P1_R1171_U151 );
not NOT1_16140 ( P1_R1171_U304 , P1_R1171_U90 );
or OR2_16141 ( P1_R1171_U305 , P1_U4020 , P1_U3058 );
nand NAND2_16142 ( P1_R1171_U306 , P1_R1171_U305 , P1_R1171_U90 );
nand NAND3_16143 ( P1_R1171_U307 , P1_R1171_U306 , P1_R1171_U170 , P1_R1171_U150 );
nand NAND2_16144 ( P1_R1171_U308 , P1_R1171_U304 , P1_R1171_U170 );
nand NAND2_16145 ( P1_R1171_U309 , P1_U4019 , P1_U3057 );
nand NAND3_16146 ( P1_R1171_U310 , P1_R1171_U308 , P1_R1171_U309 , P1_R1171_U165 );
or OR2_16147 ( P1_R1171_U311 , P1_U3058 , P1_U4020 );
nand NAND2_16148 ( P1_R1171_U312 , P1_R1171_U279 , P1_R1171_U159 );
not NOT1_16149 ( P1_R1171_U313 , P1_R1171_U92 );
nand NAND2_16150 ( P1_R1171_U314 , P1_R1171_U10 , P1_R1171_U92 );
nand NAND2_16151 ( P1_R1171_U315 , P1_R1171_U134 , P1_R1171_U314 );
nand NAND2_16152 ( P1_R1171_U316 , P1_R1171_U314 , P1_R1171_U275 );
nand NAND2_16153 ( P1_R1171_U317 , P1_R1171_U450 , P1_R1171_U316 );
or OR2_16154 ( P1_R1171_U318 , P1_U3514 , P1_U3081 );
nand NAND2_16155 ( P1_R1171_U319 , P1_R1171_U318 , P1_R1171_U92 );
nand NAND3_16156 ( P1_R1171_U320 , P1_R1171_U319 , P1_R1171_U81 , P1_R1171_U157 );
nand NAND2_16157 ( P1_R1171_U321 , P1_R1171_U313 , P1_R1171_U81 );
nand NAND2_16158 ( P1_R1171_U322 , P1_U3076 , P1_U4025 );
nand NAND3_16159 ( P1_R1171_U323 , P1_R1171_U322 , P1_R1171_U321 , P1_R1171_U10 );
or OR2_16160 ( P1_R1171_U324 , P1_U3461 , P1_U3078 );
not NOT1_16161 ( P1_R1171_U325 , P1_R1171_U158 );
or OR2_16162 ( P1_R1171_U326 , P1_U3081 , P1_U3514 );
or OR2_16163 ( P1_R1171_U327 , P1_U3506 , P1_U3073 );
nand NAND2_16164 ( P1_R1171_U328 , P1_R1171_U327 , P1_R1171_U93 );
nand NAND2_16165 ( P1_R1171_U329 , P1_R1171_U135 , P1_R1171_U328 );
nand NAND2_16166 ( P1_R1171_U330 , P1_R1171_U259 , P1_R1171_U60 );
nand NAND2_16167 ( P1_R1171_U331 , P1_U3509 , P1_U3069 );
nand NAND3_16168 ( P1_R1171_U332 , P1_R1171_U331 , P1_R1171_U330 , P1_R1171_U9 );
or OR2_16169 ( P1_R1171_U333 , P1_U3073 , P1_U3506 );
nand NAND2_16170 ( P1_R1171_U334 , P1_R1171_U247 , P1_R1171_U164 );
not NOT1_16171 ( P1_R1171_U335 , P1_R1171_U94 );
or OR2_16172 ( P1_R1171_U336 , P1_U3494 , P1_U3072 );
nand NAND2_16173 ( P1_R1171_U337 , P1_R1171_U336 , P1_R1171_U94 );
nand NAND2_16174 ( P1_R1171_U338 , P1_R1171_U136 , P1_R1171_U337 );
nand NAND2_16175 ( P1_R1171_U339 , P1_R1171_U335 , P1_R1171_U169 );
nand NAND2_16176 ( P1_R1171_U340 , P1_U3080 , P1_U3497 );
nand NAND2_16177 ( P1_R1171_U341 , P1_R1171_U137 , P1_R1171_U339 );
or OR2_16178 ( P1_R1171_U342 , P1_U3072 , P1_U3494 );
or OR2_16179 ( P1_R1171_U343 , P1_U3485 , P1_U3083 );
nand NAND2_16180 ( P1_R1171_U344 , P1_R1171_U343 , P1_R1171_U41 );
nand NAND2_16181 ( P1_R1171_U345 , P1_R1171_U138 , P1_R1171_U344 );
nand NAND2_16182 ( P1_R1171_U346 , P1_R1171_U203 , P1_R1171_U168 );
nand NAND2_16183 ( P1_R1171_U347 , P1_U3062 , P1_U3488 );
nand NAND2_16184 ( P1_R1171_U348 , P1_R1171_U139 , P1_R1171_U346 );
nand NAND2_16185 ( P1_R1171_U349 , P1_R1171_U204 , P1_R1171_U168 );
nand NAND2_16186 ( P1_R1171_U350 , P1_R1171_U201 , P1_R1171_U62 );
nand NAND2_16187 ( P1_R1171_U351 , P1_R1171_U211 , P1_R1171_U23 );
nand NAND2_16188 ( P1_R1171_U352 , P1_R1171_U225 , P1_R1171_U35 );
nand NAND2_16189 ( P1_R1171_U353 , P1_R1171_U228 , P1_R1171_U177 );
nand NAND2_16190 ( P1_R1171_U354 , P1_R1171_U311 , P1_R1171_U170 );
nand NAND2_16191 ( P1_R1171_U355 , P1_R1171_U295 , P1_R1171_U173 );
nand NAND2_16192 ( P1_R1171_U356 , P1_R1171_U326 , P1_R1171_U81 );
nand NAND2_16193 ( P1_R1171_U357 , P1_R1171_U279 , P1_R1171_U78 );
nand NAND2_16194 ( P1_R1171_U358 , P1_R1171_U333 , P1_R1171_U60 );
nand NAND2_16195 ( P1_R1171_U359 , P1_R1171_U342 , P1_R1171_U169 );
nand NAND2_16196 ( P1_R1171_U360 , P1_R1171_U247 , P1_R1171_U69 );
nand NAND2_16197 ( P1_R1171_U361 , P1_U4017 , P1_U3054 );
nand NAND2_16198 ( P1_R1171_U362 , P1_R1171_U293 , P1_R1171_U165 );
nand NAND2_16199 ( P1_R1171_U363 , P1_U3057 , P1_R1171_U292 );
nand NAND2_16200 ( P1_R1171_U364 , P1_U4019 , P1_R1171_U292 );
nand NAND3_16201 ( P1_R1171_U365 , P1_R1171_U293 , P1_R1171_U165 , P1_R1171_U298 );
nand NAND3_16202 ( P1_R1171_U366 , P1_R1171_U151 , P1_R1171_U165 , P1_R1171_U132 );
nand NAND2_16203 ( P1_R1171_U367 , P1_R1171_U294 , P1_R1171_U298 );
nand NAND2_16204 ( P1_R1171_U368 , P1_U3083 , P1_R1171_U40 );
nand NAND2_16205 ( P1_R1171_U369 , P1_U3485 , P1_R1171_U39 );
nand NAND2_16206 ( P1_R1171_U370 , P1_R1171_U369 , P1_R1171_U368 );
nand NAND2_16207 ( P1_R1171_U371 , P1_R1171_U349 , P1_R1171_U41 );
nand NAND2_16208 ( P1_R1171_U372 , P1_R1171_U370 , P1_R1171_U203 );
nand NAND2_16209 ( P1_R1171_U373 , P1_U3084 , P1_R1171_U37 );
nand NAND2_16210 ( P1_R1171_U374 , P1_U3482 , P1_R1171_U38 );
nand NAND2_16211 ( P1_R1171_U375 , P1_R1171_U374 , P1_R1171_U373 );
nand NAND2_16212 ( P1_R1171_U376 , P1_R1171_U350 , P1_R1171_U140 );
nand NAND2_16213 ( P1_R1171_U377 , P1_R1171_U200 , P1_R1171_U375 );
nand NAND2_16214 ( P1_R1171_U378 , P1_U3070 , P1_R1171_U24 );
nand NAND2_16215 ( P1_R1171_U379 , P1_U3479 , P1_R1171_U22 );
nand NAND2_16216 ( P1_R1171_U380 , P1_U3071 , P1_R1171_U20 );
nand NAND2_16217 ( P1_R1171_U381 , P1_U3476 , P1_R1171_U21 );
nand NAND2_16218 ( P1_R1171_U382 , P1_R1171_U381 , P1_R1171_U380 );
nand NAND2_16219 ( P1_R1171_U383 , P1_R1171_U351 , P1_R1171_U42 );
nand NAND2_16220 ( P1_R1171_U384 , P1_R1171_U382 , P1_R1171_U192 );
nand NAND2_16221 ( P1_R1171_U385 , P1_U3067 , P1_R1171_U36 );
nand NAND2_16222 ( P1_R1171_U386 , P1_U3473 , P1_R1171_U27 );
nand NAND2_16223 ( P1_R1171_U387 , P1_U3060 , P1_R1171_U25 );
nand NAND2_16224 ( P1_R1171_U388 , P1_U3470 , P1_R1171_U26 );
nand NAND2_16225 ( P1_R1171_U389 , P1_R1171_U388 , P1_R1171_U387 );
nand NAND2_16226 ( P1_R1171_U390 , P1_R1171_U352 , P1_R1171_U45 );
nand NAND2_16227 ( P1_R1171_U391 , P1_R1171_U389 , P1_R1171_U218 );
nand NAND2_16228 ( P1_R1171_U392 , P1_U3064 , P1_R1171_U33 );
nand NAND2_16229 ( P1_R1171_U393 , P1_U3467 , P1_R1171_U34 );
nand NAND2_16230 ( P1_R1171_U394 , P1_R1171_U393 , P1_R1171_U392 );
nand NAND2_16231 ( P1_R1171_U395 , P1_R1171_U353 , P1_R1171_U141 );
nand NAND2_16232 ( P1_R1171_U396 , P1_R1171_U227 , P1_R1171_U394 );
nand NAND2_16233 ( P1_R1171_U397 , P1_U3068 , P1_R1171_U28 );
nand NAND2_16234 ( P1_R1171_U398 , P1_U3464 , P1_R1171_U29 );
nand NAND2_16235 ( P1_R1171_U399 , P1_U3055 , P1_R1171_U143 );
nand NAND2_16236 ( P1_R1171_U400 , P1_U4028 , P1_R1171_U142 );
nand NAND2_16237 ( P1_R1171_U401 , P1_U3055 , P1_R1171_U143 );
nand NAND2_16238 ( P1_R1171_U402 , P1_U4028 , P1_R1171_U142 );
nand NAND2_16239 ( P1_R1171_U403 , P1_R1171_U402 , P1_R1171_U401 );
nand NAND2_16240 ( P1_R1171_U404 , P1_R1171_U144 , P1_R1171_U145 );
nand NAND2_16241 ( P1_R1171_U405 , P1_R1171_U302 , P1_R1171_U403 );
nand NAND2_16242 ( P1_R1171_U406 , P1_U3054 , P1_R1171_U89 );
nand NAND2_16243 ( P1_R1171_U407 , P1_U4017 , P1_R1171_U88 );
nand NAND2_16244 ( P1_R1171_U408 , P1_U3054 , P1_R1171_U89 );
nand NAND2_16245 ( P1_R1171_U409 , P1_U4017 , P1_R1171_U88 );
nand NAND2_16246 ( P1_R1171_U410 , P1_R1171_U409 , P1_R1171_U408 );
nand NAND2_16247 ( P1_R1171_U411 , P1_R1171_U146 , P1_R1171_U147 );
nand NAND2_16248 ( P1_R1171_U412 , P1_R1171_U300 , P1_R1171_U410 );
nand NAND2_16249 ( P1_R1171_U413 , P1_U3053 , P1_R1171_U47 );
nand NAND2_16250 ( P1_R1171_U414 , P1_U4018 , P1_R1171_U48 );
nand NAND2_16251 ( P1_R1171_U415 , P1_U3053 , P1_R1171_U47 );
nand NAND2_16252 ( P1_R1171_U416 , P1_U4018 , P1_R1171_U48 );
nand NAND2_16253 ( P1_R1171_U417 , P1_R1171_U416 , P1_R1171_U415 );
nand NAND2_16254 ( P1_R1171_U418 , P1_R1171_U148 , P1_R1171_U149 );
nand NAND2_16255 ( P1_R1171_U419 , P1_R1171_U297 , P1_R1171_U417 );
nand NAND2_16256 ( P1_R1171_U420 , P1_U3057 , P1_R1171_U50 );
nand NAND2_16257 ( P1_R1171_U421 , P1_U4019 , P1_R1171_U49 );
nand NAND2_16258 ( P1_R1171_U422 , P1_U3058 , P1_R1171_U51 );
nand NAND2_16259 ( P1_R1171_U423 , P1_U4020 , P1_R1171_U52 );
nand NAND2_16260 ( P1_R1171_U424 , P1_R1171_U423 , P1_R1171_U422 );
nand NAND2_16261 ( P1_R1171_U425 , P1_R1171_U354 , P1_R1171_U90 );
nand NAND2_16262 ( P1_R1171_U426 , P1_R1171_U424 , P1_R1171_U304 );
nand NAND2_16263 ( P1_R1171_U427 , P1_U3065 , P1_R1171_U53 );
nand NAND2_16264 ( P1_R1171_U428 , P1_U4021 , P1_R1171_U54 );
nand NAND2_16265 ( P1_R1171_U429 , P1_R1171_U428 , P1_R1171_U427 );
nand NAND2_16266 ( P1_R1171_U430 , P1_R1171_U355 , P1_R1171_U151 );
nand NAND2_16267 ( P1_R1171_U431 , P1_R1171_U291 , P1_R1171_U429 );
nand NAND2_16268 ( P1_R1171_U432 , P1_U3066 , P1_R1171_U85 );
nand NAND2_16269 ( P1_R1171_U433 , P1_U4022 , P1_R1171_U86 );
nand NAND2_16270 ( P1_R1171_U434 , P1_U3066 , P1_R1171_U85 );
nand NAND2_16271 ( P1_R1171_U435 , P1_U4022 , P1_R1171_U86 );
nand NAND2_16272 ( P1_R1171_U436 , P1_R1171_U435 , P1_R1171_U434 );
nand NAND2_16273 ( P1_R1171_U437 , P1_R1171_U152 , P1_R1171_U153 );
nand NAND2_16274 ( P1_R1171_U438 , P1_R1171_U287 , P1_R1171_U436 );
nand NAND2_16275 ( P1_R1171_U439 , P1_U3061 , P1_R1171_U83 );
nand NAND2_16276 ( P1_R1171_U440 , P1_U4023 , P1_R1171_U84 );
nand NAND2_16277 ( P1_R1171_U441 , P1_U3061 , P1_R1171_U83 );
nand NAND2_16278 ( P1_R1171_U442 , P1_U4023 , P1_R1171_U84 );
nand NAND2_16279 ( P1_R1171_U443 , P1_R1171_U442 , P1_R1171_U441 );
nand NAND2_16280 ( P1_R1171_U444 , P1_R1171_U154 , P1_R1171_U155 );
nand NAND2_16281 ( P1_R1171_U445 , P1_R1171_U283 , P1_R1171_U443 );
nand NAND2_16282 ( P1_R1171_U446 , P1_U3075 , P1_R1171_U55 );
nand NAND2_16283 ( P1_R1171_U447 , P1_U4024 , P1_R1171_U56 );
nand NAND2_16284 ( P1_R1171_U448 , P1_U3075 , P1_R1171_U55 );
nand NAND2_16285 ( P1_R1171_U449 , P1_U4024 , P1_R1171_U56 );
nand NAND2_16286 ( P1_R1171_U450 , P1_R1171_U449 , P1_R1171_U448 );
nand NAND2_16287 ( P1_R1171_U451 , P1_U3076 , P1_R1171_U82 );
nand NAND2_16288 ( P1_R1171_U452 , P1_U4025 , P1_R1171_U91 );
nand NAND2_16289 ( P1_R1171_U453 , P1_R1171_U179 , P1_R1171_U158 );
nand NAND2_16290 ( P1_R1171_U454 , P1_R1171_U325 , P1_R1171_U32 );
nand NAND2_16291 ( P1_R1171_U455 , P1_U3081 , P1_R1171_U79 );
nand NAND2_16292 ( P1_R1171_U456 , P1_U3514 , P1_R1171_U80 );
nand NAND2_16293 ( P1_R1171_U457 , P1_R1171_U456 , P1_R1171_U455 );
nand NAND2_16294 ( P1_R1171_U458 , P1_R1171_U356 , P1_R1171_U92 );
nand NAND2_16295 ( P1_R1171_U459 , P1_R1171_U457 , P1_R1171_U313 );
nand NAND2_16296 ( P1_R1171_U460 , P1_U3082 , P1_R1171_U76 );
nand NAND2_16297 ( P1_R1171_U461 , P1_U3512 , P1_R1171_U77 );
nand NAND2_16298 ( P1_R1171_U462 , P1_R1171_U461 , P1_R1171_U460 );
nand NAND2_16299 ( P1_R1171_U463 , P1_R1171_U357 , P1_R1171_U159 );
nand NAND2_16300 ( P1_R1171_U464 , P1_R1171_U267 , P1_R1171_U462 );
nand NAND2_16301 ( P1_R1171_U465 , P1_U3069 , P1_R1171_U61 );
nand NAND2_16302 ( P1_R1171_U466 , P1_U3509 , P1_R1171_U59 );
nand NAND2_16303 ( P1_R1171_U467 , P1_U3073 , P1_R1171_U57 );
nand NAND2_16304 ( P1_R1171_U468 , P1_U3506 , P1_R1171_U58 );
nand NAND2_16305 ( P1_R1171_U469 , P1_R1171_U468 , P1_R1171_U467 );
nand NAND2_16306 ( P1_R1171_U470 , P1_R1171_U358 , P1_R1171_U93 );
nand NAND2_16307 ( P1_R1171_U471 , P1_R1171_U469 , P1_R1171_U259 );
nand NAND2_16308 ( P1_R1171_U472 , P1_U3074 , P1_R1171_U74 );
nand NAND2_16309 ( P1_R1171_U473 , P1_U3503 , P1_R1171_U75 );
nand NAND2_16310 ( P1_R1171_U474 , P1_U3074 , P1_R1171_U74 );
nand NAND2_16311 ( P1_R1171_U475 , P1_U3503 , P1_R1171_U75 );
nand NAND2_16312 ( P1_R1171_U476 , P1_R1171_U475 , P1_R1171_U474 );
nand NAND2_16313 ( P1_R1171_U477 , P1_R1171_U160 , P1_R1171_U161 );
nand NAND2_16314 ( P1_R1171_U478 , P1_R1171_U255 , P1_R1171_U476 );
nand NAND2_16315 ( P1_R1171_U479 , P1_U3079 , P1_R1171_U72 );
nand NAND2_16316 ( P1_R1171_U480 , P1_U3500 , P1_R1171_U73 );
nand NAND2_16317 ( P1_R1171_U481 , P1_U3079 , P1_R1171_U72 );
nand NAND2_16318 ( P1_R1171_U482 , P1_U3500 , P1_R1171_U73 );
nand NAND2_16319 ( P1_R1171_U483 , P1_R1171_U482 , P1_R1171_U481 );
nand NAND2_16320 ( P1_R1171_U484 , P1_R1171_U162 , P1_R1171_U163 );
nand NAND2_16321 ( P1_R1171_U485 , P1_R1171_U251 , P1_R1171_U483 );
nand NAND2_16322 ( P1_R1171_U486 , P1_U3080 , P1_R1171_U70 );
nand NAND2_16323 ( P1_R1171_U487 , P1_U3497 , P1_R1171_U71 );
nand NAND2_16324 ( P1_R1171_U488 , P1_U3072 , P1_R1171_U65 );
nand NAND2_16325 ( P1_R1171_U489 , P1_U3494 , P1_R1171_U66 );
nand NAND2_16326 ( P1_R1171_U490 , P1_R1171_U489 , P1_R1171_U488 );
nand NAND2_16327 ( P1_R1171_U491 , P1_R1171_U359 , P1_R1171_U94 );
nand NAND2_16328 ( P1_R1171_U492 , P1_R1171_U490 , P1_R1171_U335 );
nand NAND2_16329 ( P1_R1171_U493 , P1_U3063 , P1_R1171_U67 );
nand NAND2_16330 ( P1_R1171_U494 , P1_U3491 , P1_R1171_U68 );
nand NAND2_16331 ( P1_R1171_U495 , P1_R1171_U494 , P1_R1171_U493 );
nand NAND2_16332 ( P1_R1171_U496 , P1_R1171_U360 , P1_R1171_U164 );
nand NAND2_16333 ( P1_R1171_U497 , P1_R1171_U241 , P1_R1171_U495 );
nand NAND2_16334 ( P1_R1171_U498 , P1_U3062 , P1_R1171_U63 );
nand NAND2_16335 ( P1_R1171_U499 , P1_U3488 , P1_R1171_U64 );
nand NAND2_16336 ( P1_R1171_U500 , P1_U3077 , P1_R1171_U30 );
nand NAND2_16337 ( P1_R1171_U501 , P1_U3456 , P1_R1171_U31 );
and AND2_16338 ( P1_R1138_U4 , P1_R1138_U176 , P1_R1138_U175 );
and AND2_16339 ( P1_R1138_U5 , P1_R1138_U177 , P1_R1138_U178 );
and AND2_16340 ( P1_R1138_U6 , P1_R1138_U194 , P1_R1138_U193 );
and AND2_16341 ( P1_R1138_U7 , P1_R1138_U234 , P1_R1138_U233 );
and AND2_16342 ( P1_R1138_U8 , P1_R1138_U243 , P1_R1138_U242 );
and AND2_16343 ( P1_R1138_U9 , P1_R1138_U261 , P1_R1138_U260 );
and AND2_16344 ( P1_R1138_U10 , P1_R1138_U269 , P1_R1138_U268 );
and AND2_16345 ( P1_R1138_U11 , P1_R1138_U348 , P1_R1138_U345 );
and AND2_16346 ( P1_R1138_U12 , P1_R1138_U341 , P1_R1138_U338 );
and AND2_16347 ( P1_R1138_U13 , P1_R1138_U332 , P1_R1138_U329 );
and AND2_16348 ( P1_R1138_U14 , P1_R1138_U323 , P1_R1138_U320 );
and AND2_16349 ( P1_R1138_U15 , P1_R1138_U317 , P1_R1138_U315 );
and AND2_16350 ( P1_R1138_U16 , P1_R1138_U310 , P1_R1138_U307 );
and AND2_16351 ( P1_R1138_U17 , P1_R1138_U232 , P1_R1138_U229 );
and AND2_16352 ( P1_R1138_U18 , P1_R1138_U224 , P1_R1138_U221 );
and AND2_16353 ( P1_R1138_U19 , P1_R1138_U210 , P1_R1138_U207 );
not NOT1_16354 ( P1_R1138_U20 , P1_U3476 );
not NOT1_16355 ( P1_R1138_U21 , P1_U3071 );
not NOT1_16356 ( P1_R1138_U22 , P1_U3070 );
nand NAND2_16357 ( P1_R1138_U23 , P1_U3071 , P1_U3476 );
not NOT1_16358 ( P1_R1138_U24 , P1_U3479 );
not NOT1_16359 ( P1_R1138_U25 , P1_U3470 );
not NOT1_16360 ( P1_R1138_U26 , P1_U3060 );
not NOT1_16361 ( P1_R1138_U27 , P1_U3067 );
not NOT1_16362 ( P1_R1138_U28 , P1_U3464 );
not NOT1_16363 ( P1_R1138_U29 , P1_U3068 );
not NOT1_16364 ( P1_R1138_U30 , P1_U3456 );
not NOT1_16365 ( P1_R1138_U31 , P1_U3077 );
nand NAND2_16366 ( P1_R1138_U32 , P1_U3077 , P1_U3456 );
not NOT1_16367 ( P1_R1138_U33 , P1_U3467 );
not NOT1_16368 ( P1_R1138_U34 , P1_U3064 );
nand NAND2_16369 ( P1_R1138_U35 , P1_U3060 , P1_U3470 );
not NOT1_16370 ( P1_R1138_U36 , P1_U3473 );
not NOT1_16371 ( P1_R1138_U37 , P1_U3482 );
not NOT1_16372 ( P1_R1138_U38 , P1_U3084 );
not NOT1_16373 ( P1_R1138_U39 , P1_U3083 );
not NOT1_16374 ( P1_R1138_U40 , P1_U3485 );
nand NAND2_16375 ( P1_R1138_U41 , P1_R1138_U62 , P1_R1138_U202 );
nand NAND2_16376 ( P1_R1138_U42 , P1_R1138_U118 , P1_R1138_U190 );
nand NAND2_16377 ( P1_R1138_U43 , P1_R1138_U179 , P1_R1138_U180 );
nand NAND2_16378 ( P1_R1138_U44 , P1_U3461 , P1_U3078 );
nand NAND2_16379 ( P1_R1138_U45 , P1_R1138_U122 , P1_R1138_U216 );
nand NAND2_16380 ( P1_R1138_U46 , P1_R1138_U213 , P1_R1138_U212 );
not NOT1_16381 ( P1_R1138_U47 , P1_U4018 );
not NOT1_16382 ( P1_R1138_U48 , P1_U3053 );
not NOT1_16383 ( P1_R1138_U49 , P1_U3057 );
not NOT1_16384 ( P1_R1138_U50 , P1_U4019 );
not NOT1_16385 ( P1_R1138_U51 , P1_U4020 );
not NOT1_16386 ( P1_R1138_U52 , P1_U3058 );
not NOT1_16387 ( P1_R1138_U53 , P1_U4021 );
not NOT1_16388 ( P1_R1138_U54 , P1_U3065 );
not NOT1_16389 ( P1_R1138_U55 , P1_U4024 );
not NOT1_16390 ( P1_R1138_U56 , P1_U3075 );
not NOT1_16391 ( P1_R1138_U57 , P1_U3506 );
not NOT1_16392 ( P1_R1138_U58 , P1_U3073 );
not NOT1_16393 ( P1_R1138_U59 , P1_U3069 );
nand NAND2_16394 ( P1_R1138_U60 , P1_U3073 , P1_U3506 );
not NOT1_16395 ( P1_R1138_U61 , P1_U3509 );
nand NAND2_16396 ( P1_R1138_U62 , P1_U3084 , P1_U3482 );
not NOT1_16397 ( P1_R1138_U63 , P1_U3488 );
not NOT1_16398 ( P1_R1138_U64 , P1_U3062 );
not NOT1_16399 ( P1_R1138_U65 , P1_U3494 );
not NOT1_16400 ( P1_R1138_U66 , P1_U3072 );
not NOT1_16401 ( P1_R1138_U67 , P1_U3491 );
not NOT1_16402 ( P1_R1138_U68 , P1_U3063 );
nand NAND2_16403 ( P1_R1138_U69 , P1_U3063 , P1_U3491 );
not NOT1_16404 ( P1_R1138_U70 , P1_U3497 );
not NOT1_16405 ( P1_R1138_U71 , P1_U3080 );
not NOT1_16406 ( P1_R1138_U72 , P1_U3500 );
not NOT1_16407 ( P1_R1138_U73 , P1_U3079 );
not NOT1_16408 ( P1_R1138_U74 , P1_U3503 );
not NOT1_16409 ( P1_R1138_U75 , P1_U3074 );
not NOT1_16410 ( P1_R1138_U76 , P1_U3512 );
not NOT1_16411 ( P1_R1138_U77 , P1_U3082 );
nand NAND2_16412 ( P1_R1138_U78 , P1_U3082 , P1_U3512 );
not NOT1_16413 ( P1_R1138_U79 , P1_U3514 );
not NOT1_16414 ( P1_R1138_U80 , P1_U3081 );
nand NAND2_16415 ( P1_R1138_U81 , P1_U3081 , P1_U3514 );
not NOT1_16416 ( P1_R1138_U82 , P1_U4025 );
not NOT1_16417 ( P1_R1138_U83 , P1_U4023 );
not NOT1_16418 ( P1_R1138_U84 , P1_U3061 );
not NOT1_16419 ( P1_R1138_U85 , P1_U4022 );
not NOT1_16420 ( P1_R1138_U86 , P1_U3066 );
nand NAND2_16421 ( P1_R1138_U87 , P1_U4019 , P1_U3057 );
not NOT1_16422 ( P1_R1138_U88 , P1_U3054 );
not NOT1_16423 ( P1_R1138_U89 , P1_U4017 );
nand NAND2_16424 ( P1_R1138_U90 , P1_R1138_U303 , P1_R1138_U173 );
not NOT1_16425 ( P1_R1138_U91 , P1_U3076 );
nand NAND2_16426 ( P1_R1138_U92 , P1_R1138_U78 , P1_R1138_U312 );
nand NAND2_16427 ( P1_R1138_U93 , P1_R1138_U258 , P1_R1138_U257 );
nand NAND2_16428 ( P1_R1138_U94 , P1_R1138_U69 , P1_R1138_U334 );
nand NAND2_16429 ( P1_R1138_U95 , P1_R1138_U454 , P1_R1138_U453 );
nand NAND2_16430 ( P1_R1138_U96 , P1_R1138_U501 , P1_R1138_U500 );
nand NAND2_16431 ( P1_R1138_U97 , P1_R1138_U372 , P1_R1138_U371 );
nand NAND2_16432 ( P1_R1138_U98 , P1_R1138_U377 , P1_R1138_U376 );
nand NAND2_16433 ( P1_R1138_U99 , P1_R1138_U384 , P1_R1138_U383 );
nand NAND2_16434 ( P1_R1138_U100 , P1_R1138_U391 , P1_R1138_U390 );
nand NAND2_16435 ( P1_R1138_U101 , P1_R1138_U396 , P1_R1138_U395 );
nand NAND2_16436 ( P1_R1138_U102 , P1_R1138_U405 , P1_R1138_U404 );
nand NAND2_16437 ( P1_R1138_U103 , P1_R1138_U412 , P1_R1138_U411 );
nand NAND2_16438 ( P1_R1138_U104 , P1_R1138_U419 , P1_R1138_U418 );
nand NAND2_16439 ( P1_R1138_U105 , P1_R1138_U426 , P1_R1138_U425 );
nand NAND2_16440 ( P1_R1138_U106 , P1_R1138_U431 , P1_R1138_U430 );
nand NAND2_16441 ( P1_R1138_U107 , P1_R1138_U438 , P1_R1138_U437 );
nand NAND2_16442 ( P1_R1138_U108 , P1_R1138_U445 , P1_R1138_U444 );
nand NAND2_16443 ( P1_R1138_U109 , P1_R1138_U459 , P1_R1138_U458 );
nand NAND2_16444 ( P1_R1138_U110 , P1_R1138_U464 , P1_R1138_U463 );
nand NAND2_16445 ( P1_R1138_U111 , P1_R1138_U471 , P1_R1138_U470 );
nand NAND2_16446 ( P1_R1138_U112 , P1_R1138_U478 , P1_R1138_U477 );
nand NAND2_16447 ( P1_R1138_U113 , P1_R1138_U485 , P1_R1138_U484 );
nand NAND2_16448 ( P1_R1138_U114 , P1_R1138_U492 , P1_R1138_U491 );
nand NAND2_16449 ( P1_R1138_U115 , P1_R1138_U497 , P1_R1138_U496 );
and AND2_16450 ( P1_R1138_U116 , P1_U3464 , P1_U3068 );
and AND2_16451 ( P1_R1138_U117 , P1_R1138_U186 , P1_R1138_U184 );
and AND2_16452 ( P1_R1138_U118 , P1_R1138_U191 , P1_R1138_U189 );
and AND2_16453 ( P1_R1138_U119 , P1_R1138_U198 , P1_R1138_U197 );
and AND3_16454 ( P1_R1138_U120 , P1_R1138_U379 , P1_R1138_U378 , P1_R1138_U23 );
and AND2_16455 ( P1_R1138_U121 , P1_R1138_U209 , P1_R1138_U6 );
and AND2_16456 ( P1_R1138_U122 , P1_R1138_U217 , P1_R1138_U215 );
and AND3_16457 ( P1_R1138_U123 , P1_R1138_U386 , P1_R1138_U385 , P1_R1138_U35 );
and AND2_16458 ( P1_R1138_U124 , P1_R1138_U223 , P1_R1138_U4 );
and AND2_16459 ( P1_R1138_U125 , P1_R1138_U231 , P1_R1138_U178 );
and AND2_16460 ( P1_R1138_U126 , P1_R1138_U201 , P1_R1138_U7 );
and AND2_16461 ( P1_R1138_U127 , P1_R1138_U236 , P1_R1138_U168 );
and AND2_16462 ( P1_R1138_U128 , P1_R1138_U245 , P1_R1138_U169 );
and AND2_16463 ( P1_R1138_U129 , P1_R1138_U265 , P1_R1138_U264 );
and AND2_16464 ( P1_R1138_U130 , P1_R1138_U10 , P1_R1138_U279 );
and AND2_16465 ( P1_R1138_U131 , P1_R1138_U282 , P1_R1138_U277 );
and AND2_16466 ( P1_R1138_U132 , P1_R1138_U298 , P1_R1138_U295 );
and AND2_16467 ( P1_R1138_U133 , P1_R1138_U365 , P1_R1138_U299 );
and AND2_16468 ( P1_R1138_U134 , P1_R1138_U156 , P1_R1138_U275 );
and AND3_16469 ( P1_R1138_U135 , P1_R1138_U466 , P1_R1138_U465 , P1_R1138_U60 );
and AND3_16470 ( P1_R1138_U136 , P1_R1138_U487 , P1_R1138_U486 , P1_R1138_U169 );
and AND2_16471 ( P1_R1138_U137 , P1_R1138_U340 , P1_R1138_U8 );
and AND3_16472 ( P1_R1138_U138 , P1_R1138_U499 , P1_R1138_U498 , P1_R1138_U168 );
and AND2_16473 ( P1_R1138_U139 , P1_R1138_U347 , P1_R1138_U7 );
nand NAND2_16474 ( P1_R1138_U140 , P1_R1138_U119 , P1_R1138_U199 );
nand NAND2_16475 ( P1_R1138_U141 , P1_R1138_U214 , P1_R1138_U226 );
not NOT1_16476 ( P1_R1138_U142 , P1_U3055 );
not NOT1_16477 ( P1_R1138_U143 , P1_U4028 );
and AND2_16478 ( P1_R1138_U144 , P1_R1138_U400 , P1_R1138_U399 );
nand NAND3_16479 ( P1_R1138_U145 , P1_R1138_U301 , P1_R1138_U166 , P1_R1138_U361 );
and AND2_16480 ( P1_R1138_U146 , P1_R1138_U407 , P1_R1138_U406 );
nand NAND3_16481 ( P1_R1138_U147 , P1_R1138_U367 , P1_R1138_U366 , P1_R1138_U133 );
and AND2_16482 ( P1_R1138_U148 , P1_R1138_U414 , P1_R1138_U413 );
nand NAND3_16483 ( P1_R1138_U149 , P1_R1138_U362 , P1_R1138_U296 , P1_R1138_U87 );
and AND2_16484 ( P1_R1138_U150 , P1_R1138_U421 , P1_R1138_U420 );
nand NAND2_16485 ( P1_R1138_U151 , P1_R1138_U290 , P1_R1138_U289 );
and AND2_16486 ( P1_R1138_U152 , P1_R1138_U433 , P1_R1138_U432 );
nand NAND2_16487 ( P1_R1138_U153 , P1_R1138_U286 , P1_R1138_U285 );
and AND2_16488 ( P1_R1138_U154 , P1_R1138_U440 , P1_R1138_U439 );
nand NAND2_16489 ( P1_R1138_U155 , P1_R1138_U131 , P1_R1138_U281 );
and AND2_16490 ( P1_R1138_U156 , P1_R1138_U447 , P1_R1138_U446 );
and AND2_16491 ( P1_R1138_U157 , P1_R1138_U452 , P1_R1138_U451 );
nand NAND2_16492 ( P1_R1138_U158 , P1_R1138_U44 , P1_R1138_U324 );
nand NAND2_16493 ( P1_R1138_U159 , P1_R1138_U129 , P1_R1138_U266 );
and AND2_16494 ( P1_R1138_U160 , P1_R1138_U473 , P1_R1138_U472 );
nand NAND2_16495 ( P1_R1138_U161 , P1_R1138_U254 , P1_R1138_U253 );
and AND2_16496 ( P1_R1138_U162 , P1_R1138_U480 , P1_R1138_U479 );
nand NAND2_16497 ( P1_R1138_U163 , P1_R1138_U250 , P1_R1138_U249 );
nand NAND2_16498 ( P1_R1138_U164 , P1_R1138_U240 , P1_R1138_U239 );
nand NAND2_16499 ( P1_R1138_U165 , P1_R1138_U364 , P1_R1138_U363 );
nand NAND2_16500 ( P1_R1138_U166 , P1_U3054 , P1_R1138_U147 );
not NOT1_16501 ( P1_R1138_U167 , P1_R1138_U35 );
nand NAND2_16502 ( P1_R1138_U168 , P1_U3485 , P1_U3083 );
nand NAND2_16503 ( P1_R1138_U169 , P1_U3072 , P1_U3494 );
nand NAND2_16504 ( P1_R1138_U170 , P1_U3058 , P1_U4020 );
not NOT1_16505 ( P1_R1138_U171 , P1_R1138_U69 );
not NOT1_16506 ( P1_R1138_U172 , P1_R1138_U78 );
nand NAND2_16507 ( P1_R1138_U173 , P1_U3065 , P1_U4021 );
not NOT1_16508 ( P1_R1138_U174 , P1_R1138_U62 );
or OR2_16509 ( P1_R1138_U175 , P1_U3067 , P1_U3473 );
or OR2_16510 ( P1_R1138_U176 , P1_U3060 , P1_U3470 );
or OR2_16511 ( P1_R1138_U177 , P1_U3467 , P1_U3064 );
or OR2_16512 ( P1_R1138_U178 , P1_U3464 , P1_U3068 );
not NOT1_16513 ( P1_R1138_U179 , P1_R1138_U32 );
or OR2_16514 ( P1_R1138_U180 , P1_U3461 , P1_U3078 );
not NOT1_16515 ( P1_R1138_U181 , P1_R1138_U43 );
not NOT1_16516 ( P1_R1138_U182 , P1_R1138_U44 );
nand NAND2_16517 ( P1_R1138_U183 , P1_R1138_U43 , P1_R1138_U44 );
nand NAND2_16518 ( P1_R1138_U184 , P1_R1138_U116 , P1_R1138_U177 );
nand NAND2_16519 ( P1_R1138_U185 , P1_R1138_U5 , P1_R1138_U183 );
nand NAND2_16520 ( P1_R1138_U186 , P1_U3064 , P1_U3467 );
nand NAND2_16521 ( P1_R1138_U187 , P1_R1138_U117 , P1_R1138_U185 );
nand NAND2_16522 ( P1_R1138_U188 , P1_R1138_U36 , P1_R1138_U35 );
nand NAND2_16523 ( P1_R1138_U189 , P1_U3067 , P1_R1138_U188 );
nand NAND2_16524 ( P1_R1138_U190 , P1_R1138_U4 , P1_R1138_U187 );
nand NAND2_16525 ( P1_R1138_U191 , P1_U3473 , P1_R1138_U167 );
not NOT1_16526 ( P1_R1138_U192 , P1_R1138_U42 );
or OR2_16527 ( P1_R1138_U193 , P1_U3070 , P1_U3479 );
or OR2_16528 ( P1_R1138_U194 , P1_U3071 , P1_U3476 );
not NOT1_16529 ( P1_R1138_U195 , P1_R1138_U23 );
nand NAND2_16530 ( P1_R1138_U196 , P1_R1138_U24 , P1_R1138_U23 );
nand NAND2_16531 ( P1_R1138_U197 , P1_U3070 , P1_R1138_U196 );
nand NAND2_16532 ( P1_R1138_U198 , P1_U3479 , P1_R1138_U195 );
nand NAND2_16533 ( P1_R1138_U199 , P1_R1138_U6 , P1_R1138_U42 );
not NOT1_16534 ( P1_R1138_U200 , P1_R1138_U140 );
or OR2_16535 ( P1_R1138_U201 , P1_U3482 , P1_U3084 );
nand NAND2_16536 ( P1_R1138_U202 , P1_R1138_U201 , P1_R1138_U140 );
not NOT1_16537 ( P1_R1138_U203 , P1_R1138_U41 );
or OR2_16538 ( P1_R1138_U204 , P1_U3083 , P1_U3485 );
or OR2_16539 ( P1_R1138_U205 , P1_U3476 , P1_U3071 );
nand NAND2_16540 ( P1_R1138_U206 , P1_R1138_U205 , P1_R1138_U42 );
nand NAND2_16541 ( P1_R1138_U207 , P1_R1138_U120 , P1_R1138_U206 );
nand NAND2_16542 ( P1_R1138_U208 , P1_R1138_U192 , P1_R1138_U23 );
nand NAND2_16543 ( P1_R1138_U209 , P1_U3479 , P1_U3070 );
nand NAND2_16544 ( P1_R1138_U210 , P1_R1138_U121 , P1_R1138_U208 );
or OR2_16545 ( P1_R1138_U211 , P1_U3071 , P1_U3476 );
nand NAND2_16546 ( P1_R1138_U212 , P1_R1138_U182 , P1_R1138_U178 );
nand NAND2_16547 ( P1_R1138_U213 , P1_U3068 , P1_U3464 );
not NOT1_16548 ( P1_R1138_U214 , P1_R1138_U46 );
nand NAND2_16549 ( P1_R1138_U215 , P1_R1138_U181 , P1_R1138_U5 );
nand NAND2_16550 ( P1_R1138_U216 , P1_R1138_U46 , P1_R1138_U177 );
nand NAND2_16551 ( P1_R1138_U217 , P1_U3064 , P1_U3467 );
not NOT1_16552 ( P1_R1138_U218 , P1_R1138_U45 );
or OR2_16553 ( P1_R1138_U219 , P1_U3470 , P1_U3060 );
nand NAND2_16554 ( P1_R1138_U220 , P1_R1138_U219 , P1_R1138_U45 );
nand NAND2_16555 ( P1_R1138_U221 , P1_R1138_U123 , P1_R1138_U220 );
nand NAND2_16556 ( P1_R1138_U222 , P1_R1138_U218 , P1_R1138_U35 );
nand NAND2_16557 ( P1_R1138_U223 , P1_U3473 , P1_U3067 );
nand NAND2_16558 ( P1_R1138_U224 , P1_R1138_U124 , P1_R1138_U222 );
or OR2_16559 ( P1_R1138_U225 , P1_U3060 , P1_U3470 );
nand NAND2_16560 ( P1_R1138_U226 , P1_R1138_U181 , P1_R1138_U178 );
not NOT1_16561 ( P1_R1138_U227 , P1_R1138_U141 );
nand NAND2_16562 ( P1_R1138_U228 , P1_U3064 , P1_U3467 );
nand NAND4_16563 ( P1_R1138_U229 , P1_R1138_U398 , P1_R1138_U397 , P1_R1138_U44 , P1_R1138_U43 );
nand NAND2_16564 ( P1_R1138_U230 , P1_R1138_U44 , P1_R1138_U43 );
nand NAND2_16565 ( P1_R1138_U231 , P1_U3068 , P1_U3464 );
nand NAND2_16566 ( P1_R1138_U232 , P1_R1138_U125 , P1_R1138_U230 );
or OR2_16567 ( P1_R1138_U233 , P1_U3083 , P1_U3485 );
or OR2_16568 ( P1_R1138_U234 , P1_U3062 , P1_U3488 );
nand NAND2_16569 ( P1_R1138_U235 , P1_R1138_U174 , P1_R1138_U7 );
nand NAND2_16570 ( P1_R1138_U236 , P1_U3062 , P1_U3488 );
nand NAND2_16571 ( P1_R1138_U237 , P1_R1138_U127 , P1_R1138_U235 );
or OR2_16572 ( P1_R1138_U238 , P1_U3488 , P1_U3062 );
nand NAND2_16573 ( P1_R1138_U239 , P1_R1138_U126 , P1_R1138_U140 );
nand NAND2_16574 ( P1_R1138_U240 , P1_R1138_U238 , P1_R1138_U237 );
not NOT1_16575 ( P1_R1138_U241 , P1_R1138_U164 );
or OR2_16576 ( P1_R1138_U242 , P1_U3080 , P1_U3497 );
or OR2_16577 ( P1_R1138_U243 , P1_U3072 , P1_U3494 );
nand NAND2_16578 ( P1_R1138_U244 , P1_R1138_U171 , P1_R1138_U8 );
nand NAND2_16579 ( P1_R1138_U245 , P1_U3080 , P1_U3497 );
nand NAND2_16580 ( P1_R1138_U246 , P1_R1138_U128 , P1_R1138_U244 );
or OR2_16581 ( P1_R1138_U247 , P1_U3491 , P1_U3063 );
or OR2_16582 ( P1_R1138_U248 , P1_U3497 , P1_U3080 );
nand NAND3_16583 ( P1_R1138_U249 , P1_R1138_U247 , P1_R1138_U164 , P1_R1138_U8 );
nand NAND2_16584 ( P1_R1138_U250 , P1_R1138_U248 , P1_R1138_U246 );
not NOT1_16585 ( P1_R1138_U251 , P1_R1138_U163 );
or OR2_16586 ( P1_R1138_U252 , P1_U3500 , P1_U3079 );
nand NAND2_16587 ( P1_R1138_U253 , P1_R1138_U252 , P1_R1138_U163 );
nand NAND2_16588 ( P1_R1138_U254 , P1_U3079 , P1_U3500 );
not NOT1_16589 ( P1_R1138_U255 , P1_R1138_U161 );
or OR2_16590 ( P1_R1138_U256 , P1_U3503 , P1_U3074 );
nand NAND2_16591 ( P1_R1138_U257 , P1_R1138_U256 , P1_R1138_U161 );
nand NAND2_16592 ( P1_R1138_U258 , P1_U3074 , P1_U3503 );
not NOT1_16593 ( P1_R1138_U259 , P1_R1138_U93 );
or OR2_16594 ( P1_R1138_U260 , P1_U3069 , P1_U3509 );
or OR2_16595 ( P1_R1138_U261 , P1_U3073 , P1_U3506 );
not NOT1_16596 ( P1_R1138_U262 , P1_R1138_U60 );
nand NAND2_16597 ( P1_R1138_U263 , P1_R1138_U61 , P1_R1138_U60 );
nand NAND2_16598 ( P1_R1138_U264 , P1_U3069 , P1_R1138_U263 );
nand NAND2_16599 ( P1_R1138_U265 , P1_U3509 , P1_R1138_U262 );
nand NAND2_16600 ( P1_R1138_U266 , P1_R1138_U9 , P1_R1138_U93 );
not NOT1_16601 ( P1_R1138_U267 , P1_R1138_U159 );
or OR2_16602 ( P1_R1138_U268 , P1_U3076 , P1_U4025 );
or OR2_16603 ( P1_R1138_U269 , P1_U3081 , P1_U3514 );
or OR2_16604 ( P1_R1138_U270 , P1_U3075 , P1_U4024 );
not NOT1_16605 ( P1_R1138_U271 , P1_R1138_U81 );
nand NAND2_16606 ( P1_R1138_U272 , P1_U4025 , P1_R1138_U271 );
nand NAND2_16607 ( P1_R1138_U273 , P1_R1138_U272 , P1_R1138_U91 );
nand NAND2_16608 ( P1_R1138_U274 , P1_R1138_U81 , P1_R1138_U82 );
nand NAND2_16609 ( P1_R1138_U275 , P1_R1138_U274 , P1_R1138_U273 );
nand NAND2_16610 ( P1_R1138_U276 , P1_R1138_U172 , P1_R1138_U10 );
nand NAND2_16611 ( P1_R1138_U277 , P1_U3075 , P1_U4024 );
nand NAND2_16612 ( P1_R1138_U278 , P1_R1138_U275 , P1_R1138_U276 );
or OR2_16613 ( P1_R1138_U279 , P1_U3512 , P1_U3082 );
or OR2_16614 ( P1_R1138_U280 , P1_U4024 , P1_U3075 );
nand NAND3_16615 ( P1_R1138_U281 , P1_R1138_U270 , P1_R1138_U159 , P1_R1138_U130 );
nand NAND2_16616 ( P1_R1138_U282 , P1_R1138_U280 , P1_R1138_U278 );
not NOT1_16617 ( P1_R1138_U283 , P1_R1138_U155 );
or OR2_16618 ( P1_R1138_U284 , P1_U4023 , P1_U3061 );
nand NAND2_16619 ( P1_R1138_U285 , P1_R1138_U284 , P1_R1138_U155 );
nand NAND2_16620 ( P1_R1138_U286 , P1_U3061 , P1_U4023 );
not NOT1_16621 ( P1_R1138_U287 , P1_R1138_U153 );
or OR2_16622 ( P1_R1138_U288 , P1_U4022 , P1_U3066 );
nand NAND2_16623 ( P1_R1138_U289 , P1_R1138_U288 , P1_R1138_U153 );
nand NAND2_16624 ( P1_R1138_U290 , P1_U3066 , P1_U4022 );
not NOT1_16625 ( P1_R1138_U291 , P1_R1138_U151 );
or OR2_16626 ( P1_R1138_U292 , P1_U3058 , P1_U4020 );
nand NAND2_16627 ( P1_R1138_U293 , P1_R1138_U173 , P1_R1138_U170 );
not NOT1_16628 ( P1_R1138_U294 , P1_R1138_U87 );
or OR2_16629 ( P1_R1138_U295 , P1_U4021 , P1_U3065 );
nand NAND3_16630 ( P1_R1138_U296 , P1_R1138_U151 , P1_R1138_U295 , P1_R1138_U165 );
not NOT1_16631 ( P1_R1138_U297 , P1_R1138_U149 );
or OR2_16632 ( P1_R1138_U298 , P1_U4018 , P1_U3053 );
nand NAND2_16633 ( P1_R1138_U299 , P1_U3053 , P1_U4018 );
not NOT1_16634 ( P1_R1138_U300 , P1_R1138_U147 );
nand NAND2_16635 ( P1_R1138_U301 , P1_U4017 , P1_R1138_U147 );
not NOT1_16636 ( P1_R1138_U302 , P1_R1138_U145 );
nand NAND2_16637 ( P1_R1138_U303 , P1_R1138_U295 , P1_R1138_U151 );
not NOT1_16638 ( P1_R1138_U304 , P1_R1138_U90 );
or OR2_16639 ( P1_R1138_U305 , P1_U4020 , P1_U3058 );
nand NAND2_16640 ( P1_R1138_U306 , P1_R1138_U305 , P1_R1138_U90 );
nand NAND3_16641 ( P1_R1138_U307 , P1_R1138_U306 , P1_R1138_U170 , P1_R1138_U150 );
nand NAND2_16642 ( P1_R1138_U308 , P1_R1138_U304 , P1_R1138_U170 );
nand NAND2_16643 ( P1_R1138_U309 , P1_U4019 , P1_U3057 );
nand NAND3_16644 ( P1_R1138_U310 , P1_R1138_U308 , P1_R1138_U309 , P1_R1138_U165 );
or OR2_16645 ( P1_R1138_U311 , P1_U3058 , P1_U4020 );
nand NAND2_16646 ( P1_R1138_U312 , P1_R1138_U279 , P1_R1138_U159 );
not NOT1_16647 ( P1_R1138_U313 , P1_R1138_U92 );
nand NAND2_16648 ( P1_R1138_U314 , P1_R1138_U10 , P1_R1138_U92 );
nand NAND2_16649 ( P1_R1138_U315 , P1_R1138_U134 , P1_R1138_U314 );
nand NAND2_16650 ( P1_R1138_U316 , P1_R1138_U314 , P1_R1138_U275 );
nand NAND2_16651 ( P1_R1138_U317 , P1_R1138_U450 , P1_R1138_U316 );
or OR2_16652 ( P1_R1138_U318 , P1_U3514 , P1_U3081 );
nand NAND2_16653 ( P1_R1138_U319 , P1_R1138_U318 , P1_R1138_U92 );
nand NAND3_16654 ( P1_R1138_U320 , P1_R1138_U319 , P1_R1138_U81 , P1_R1138_U157 );
nand NAND2_16655 ( P1_R1138_U321 , P1_R1138_U313 , P1_R1138_U81 );
nand NAND2_16656 ( P1_R1138_U322 , P1_U3076 , P1_U4025 );
nand NAND3_16657 ( P1_R1138_U323 , P1_R1138_U322 , P1_R1138_U321 , P1_R1138_U10 );
or OR2_16658 ( P1_R1138_U324 , P1_U3461 , P1_U3078 );
not NOT1_16659 ( P1_R1138_U325 , P1_R1138_U158 );
or OR2_16660 ( P1_R1138_U326 , P1_U3081 , P1_U3514 );
or OR2_16661 ( P1_R1138_U327 , P1_U3506 , P1_U3073 );
nand NAND2_16662 ( P1_R1138_U328 , P1_R1138_U327 , P1_R1138_U93 );
nand NAND2_16663 ( P1_R1138_U329 , P1_R1138_U135 , P1_R1138_U328 );
nand NAND2_16664 ( P1_R1138_U330 , P1_R1138_U259 , P1_R1138_U60 );
nand NAND2_16665 ( P1_R1138_U331 , P1_U3509 , P1_U3069 );
nand NAND3_16666 ( P1_R1138_U332 , P1_R1138_U331 , P1_R1138_U330 , P1_R1138_U9 );
or OR2_16667 ( P1_R1138_U333 , P1_U3073 , P1_U3506 );
nand NAND2_16668 ( P1_R1138_U334 , P1_R1138_U247 , P1_R1138_U164 );
not NOT1_16669 ( P1_R1138_U335 , P1_R1138_U94 );
or OR2_16670 ( P1_R1138_U336 , P1_U3494 , P1_U3072 );
nand NAND2_16671 ( P1_R1138_U337 , P1_R1138_U336 , P1_R1138_U94 );
nand NAND2_16672 ( P1_R1138_U338 , P1_R1138_U136 , P1_R1138_U337 );
nand NAND2_16673 ( P1_R1138_U339 , P1_R1138_U335 , P1_R1138_U169 );
nand NAND2_16674 ( P1_R1138_U340 , P1_U3080 , P1_U3497 );
nand NAND2_16675 ( P1_R1138_U341 , P1_R1138_U137 , P1_R1138_U339 );
or OR2_16676 ( P1_R1138_U342 , P1_U3072 , P1_U3494 );
or OR2_16677 ( P1_R1138_U343 , P1_U3485 , P1_U3083 );
nand NAND2_16678 ( P1_R1138_U344 , P1_R1138_U343 , P1_R1138_U41 );
nand NAND2_16679 ( P1_R1138_U345 , P1_R1138_U138 , P1_R1138_U344 );
nand NAND2_16680 ( P1_R1138_U346 , P1_R1138_U203 , P1_R1138_U168 );
nand NAND2_16681 ( P1_R1138_U347 , P1_U3062 , P1_U3488 );
nand NAND2_16682 ( P1_R1138_U348 , P1_R1138_U139 , P1_R1138_U346 );
nand NAND2_16683 ( P1_R1138_U349 , P1_R1138_U204 , P1_R1138_U168 );
nand NAND2_16684 ( P1_R1138_U350 , P1_R1138_U201 , P1_R1138_U62 );
nand NAND2_16685 ( P1_R1138_U351 , P1_R1138_U211 , P1_R1138_U23 );
nand NAND2_16686 ( P1_R1138_U352 , P1_R1138_U225 , P1_R1138_U35 );
nand NAND2_16687 ( P1_R1138_U353 , P1_R1138_U228 , P1_R1138_U177 );
nand NAND2_16688 ( P1_R1138_U354 , P1_R1138_U311 , P1_R1138_U170 );
nand NAND2_16689 ( P1_R1138_U355 , P1_R1138_U295 , P1_R1138_U173 );
nand NAND2_16690 ( P1_R1138_U356 , P1_R1138_U326 , P1_R1138_U81 );
nand NAND2_16691 ( P1_R1138_U357 , P1_R1138_U279 , P1_R1138_U78 );
nand NAND2_16692 ( P1_R1138_U358 , P1_R1138_U333 , P1_R1138_U60 );
nand NAND2_16693 ( P1_R1138_U359 , P1_R1138_U342 , P1_R1138_U169 );
nand NAND2_16694 ( P1_R1138_U360 , P1_R1138_U247 , P1_R1138_U69 );
nand NAND2_16695 ( P1_R1138_U361 , P1_U4017 , P1_U3054 );
nand NAND2_16696 ( P1_R1138_U362 , P1_R1138_U293 , P1_R1138_U165 );
nand NAND2_16697 ( P1_R1138_U363 , P1_U3057 , P1_R1138_U292 );
nand NAND2_16698 ( P1_R1138_U364 , P1_U4019 , P1_R1138_U292 );
nand NAND3_16699 ( P1_R1138_U365 , P1_R1138_U293 , P1_R1138_U165 , P1_R1138_U298 );
nand NAND3_16700 ( P1_R1138_U366 , P1_R1138_U151 , P1_R1138_U165 , P1_R1138_U132 );
nand NAND2_16701 ( P1_R1138_U367 , P1_R1138_U294 , P1_R1138_U298 );
nand NAND2_16702 ( P1_R1138_U368 , P1_U3083 , P1_R1138_U40 );
nand NAND2_16703 ( P1_R1138_U369 , P1_U3485 , P1_R1138_U39 );
nand NAND2_16704 ( P1_R1138_U370 , P1_R1138_U369 , P1_R1138_U368 );
nand NAND2_16705 ( P1_R1138_U371 , P1_R1138_U349 , P1_R1138_U41 );
nand NAND2_16706 ( P1_R1138_U372 , P1_R1138_U370 , P1_R1138_U203 );
nand NAND2_16707 ( P1_R1138_U373 , P1_U3084 , P1_R1138_U37 );
nand NAND2_16708 ( P1_R1138_U374 , P1_U3482 , P1_R1138_U38 );
nand NAND2_16709 ( P1_R1138_U375 , P1_R1138_U374 , P1_R1138_U373 );
nand NAND2_16710 ( P1_R1138_U376 , P1_R1138_U350 , P1_R1138_U140 );
nand NAND2_16711 ( P1_R1138_U377 , P1_R1138_U200 , P1_R1138_U375 );
nand NAND2_16712 ( P1_R1138_U378 , P1_U3070 , P1_R1138_U24 );
nand NAND2_16713 ( P1_R1138_U379 , P1_U3479 , P1_R1138_U22 );
nand NAND2_16714 ( P1_R1138_U380 , P1_U3071 , P1_R1138_U20 );
nand NAND2_16715 ( P1_R1138_U381 , P1_U3476 , P1_R1138_U21 );
nand NAND2_16716 ( P1_R1138_U382 , P1_R1138_U381 , P1_R1138_U380 );
nand NAND2_16717 ( P1_R1138_U383 , P1_R1138_U351 , P1_R1138_U42 );
nand NAND2_16718 ( P1_R1138_U384 , P1_R1138_U382 , P1_R1138_U192 );
nand NAND2_16719 ( P1_R1138_U385 , P1_U3067 , P1_R1138_U36 );
nand NAND2_16720 ( P1_R1138_U386 , P1_U3473 , P1_R1138_U27 );
nand NAND2_16721 ( P1_R1138_U387 , P1_U3060 , P1_R1138_U25 );
nand NAND2_16722 ( P1_R1138_U388 , P1_U3470 , P1_R1138_U26 );
nand NAND2_16723 ( P1_R1138_U389 , P1_R1138_U388 , P1_R1138_U387 );
nand NAND2_16724 ( P1_R1138_U390 , P1_R1138_U352 , P1_R1138_U45 );
nand NAND2_16725 ( P1_R1138_U391 , P1_R1138_U389 , P1_R1138_U218 );
nand NAND2_16726 ( P1_R1138_U392 , P1_U3064 , P1_R1138_U33 );
nand NAND2_16727 ( P1_R1138_U393 , P1_U3467 , P1_R1138_U34 );
nand NAND2_16728 ( P1_R1138_U394 , P1_R1138_U393 , P1_R1138_U392 );
nand NAND2_16729 ( P1_R1138_U395 , P1_R1138_U353 , P1_R1138_U141 );
nand NAND2_16730 ( P1_R1138_U396 , P1_R1138_U227 , P1_R1138_U394 );
nand NAND2_16731 ( P1_R1138_U397 , P1_U3068 , P1_R1138_U28 );
nand NAND2_16732 ( P1_R1138_U398 , P1_U3464 , P1_R1138_U29 );
nand NAND2_16733 ( P1_R1138_U399 , P1_U3055 , P1_R1138_U143 );
nand NAND2_16734 ( P1_R1138_U400 , P1_U4028 , P1_R1138_U142 );
nand NAND2_16735 ( P1_R1138_U401 , P1_U3055 , P1_R1138_U143 );
nand NAND2_16736 ( P1_R1138_U402 , P1_U4028 , P1_R1138_U142 );
nand NAND2_16737 ( P1_R1138_U403 , P1_R1138_U402 , P1_R1138_U401 );
nand NAND2_16738 ( P1_R1138_U404 , P1_R1138_U144 , P1_R1138_U145 );
nand NAND2_16739 ( P1_R1138_U405 , P1_R1138_U302 , P1_R1138_U403 );
nand NAND2_16740 ( P1_R1138_U406 , P1_U3054 , P1_R1138_U89 );
nand NAND2_16741 ( P1_R1138_U407 , P1_U4017 , P1_R1138_U88 );
nand NAND2_16742 ( P1_R1138_U408 , P1_U3054 , P1_R1138_U89 );
nand NAND2_16743 ( P1_R1138_U409 , P1_U4017 , P1_R1138_U88 );
nand NAND2_16744 ( P1_R1138_U410 , P1_R1138_U409 , P1_R1138_U408 );
nand NAND2_16745 ( P1_R1138_U411 , P1_R1138_U146 , P1_R1138_U147 );
nand NAND2_16746 ( P1_R1138_U412 , P1_R1138_U300 , P1_R1138_U410 );
nand NAND2_16747 ( P1_R1138_U413 , P1_U3053 , P1_R1138_U47 );
nand NAND2_16748 ( P1_R1138_U414 , P1_U4018 , P1_R1138_U48 );
nand NAND2_16749 ( P1_R1138_U415 , P1_U3053 , P1_R1138_U47 );
nand NAND2_16750 ( P1_R1138_U416 , P1_U4018 , P1_R1138_U48 );
nand NAND2_16751 ( P1_R1138_U417 , P1_R1138_U416 , P1_R1138_U415 );
nand NAND2_16752 ( P1_R1138_U418 , P1_R1138_U148 , P1_R1138_U149 );
nand NAND2_16753 ( P1_R1138_U419 , P1_R1138_U297 , P1_R1138_U417 );
nand NAND2_16754 ( P1_R1138_U420 , P1_U3057 , P1_R1138_U50 );
nand NAND2_16755 ( P1_R1138_U421 , P1_U4019 , P1_R1138_U49 );
nand NAND2_16756 ( P1_R1138_U422 , P1_U3058 , P1_R1138_U51 );
nand NAND2_16757 ( P1_R1138_U423 , P1_U4020 , P1_R1138_U52 );
nand NAND2_16758 ( P1_R1138_U424 , P1_R1138_U423 , P1_R1138_U422 );
nand NAND2_16759 ( P1_R1138_U425 , P1_R1138_U354 , P1_R1138_U90 );
nand NAND2_16760 ( P1_R1138_U426 , P1_R1138_U424 , P1_R1138_U304 );
nand NAND2_16761 ( P1_R1138_U427 , P1_U3065 , P1_R1138_U53 );
nand NAND2_16762 ( P1_R1138_U428 , P1_U4021 , P1_R1138_U54 );
nand NAND2_16763 ( P1_R1138_U429 , P1_R1138_U428 , P1_R1138_U427 );
nand NAND2_16764 ( P1_R1138_U430 , P1_R1138_U355 , P1_R1138_U151 );
nand NAND2_16765 ( P1_R1138_U431 , P1_R1138_U291 , P1_R1138_U429 );
nand NAND2_16766 ( P1_R1138_U432 , P1_U3066 , P1_R1138_U85 );
nand NAND2_16767 ( P1_R1138_U433 , P1_U4022 , P1_R1138_U86 );
nand NAND2_16768 ( P1_R1138_U434 , P1_U3066 , P1_R1138_U85 );
nand NAND2_16769 ( P1_R1138_U435 , P1_U4022 , P1_R1138_U86 );
nand NAND2_16770 ( P1_R1138_U436 , P1_R1138_U435 , P1_R1138_U434 );
nand NAND2_16771 ( P1_R1138_U437 , P1_R1138_U152 , P1_R1138_U153 );
nand NAND2_16772 ( P1_R1138_U438 , P1_R1138_U287 , P1_R1138_U436 );
nand NAND2_16773 ( P1_R1138_U439 , P1_U3061 , P1_R1138_U83 );
nand NAND2_16774 ( P1_R1138_U440 , P1_U4023 , P1_R1138_U84 );
nand NAND2_16775 ( P1_R1138_U441 , P1_U3061 , P1_R1138_U83 );
nand NAND2_16776 ( P1_R1138_U442 , P1_U4023 , P1_R1138_U84 );
nand NAND2_16777 ( P1_R1138_U443 , P1_R1138_U442 , P1_R1138_U441 );
nand NAND2_16778 ( P1_R1138_U444 , P1_R1138_U154 , P1_R1138_U155 );
nand NAND2_16779 ( P1_R1138_U445 , P1_R1138_U283 , P1_R1138_U443 );
nand NAND2_16780 ( P1_R1138_U446 , P1_U3075 , P1_R1138_U55 );
nand NAND2_16781 ( P1_R1138_U447 , P1_U4024 , P1_R1138_U56 );
nand NAND2_16782 ( P1_R1138_U448 , P1_U3075 , P1_R1138_U55 );
nand NAND2_16783 ( P1_R1138_U449 , P1_U4024 , P1_R1138_U56 );
nand NAND2_16784 ( P1_R1138_U450 , P1_R1138_U449 , P1_R1138_U448 );
nand NAND2_16785 ( P1_R1138_U451 , P1_U3076 , P1_R1138_U82 );
nand NAND2_16786 ( P1_R1138_U452 , P1_U4025 , P1_R1138_U91 );
nand NAND2_16787 ( P1_R1138_U453 , P1_R1138_U179 , P1_R1138_U158 );
nand NAND2_16788 ( P1_R1138_U454 , P1_R1138_U325 , P1_R1138_U32 );
nand NAND2_16789 ( P1_R1138_U455 , P1_U3081 , P1_R1138_U79 );
nand NAND2_16790 ( P1_R1138_U456 , P1_U3514 , P1_R1138_U80 );
nand NAND2_16791 ( P1_R1138_U457 , P1_R1138_U456 , P1_R1138_U455 );
nand NAND2_16792 ( P1_R1138_U458 , P1_R1138_U356 , P1_R1138_U92 );
nand NAND2_16793 ( P1_R1138_U459 , P1_R1138_U457 , P1_R1138_U313 );
nand NAND2_16794 ( P1_R1138_U460 , P1_U3082 , P1_R1138_U76 );
nand NAND2_16795 ( P1_R1138_U461 , P1_U3512 , P1_R1138_U77 );
nand NAND2_16796 ( P1_R1138_U462 , P1_R1138_U461 , P1_R1138_U460 );
nand NAND2_16797 ( P1_R1138_U463 , P1_R1138_U357 , P1_R1138_U159 );
nand NAND2_16798 ( P1_R1138_U464 , P1_R1138_U267 , P1_R1138_U462 );
nand NAND2_16799 ( P1_R1138_U465 , P1_U3069 , P1_R1138_U61 );
nand NAND2_16800 ( P1_R1138_U466 , P1_U3509 , P1_R1138_U59 );
nand NAND2_16801 ( P1_R1138_U467 , P1_U3073 , P1_R1138_U57 );
nand NAND2_16802 ( P1_R1138_U468 , P1_U3506 , P1_R1138_U58 );
nand NAND2_16803 ( P1_R1138_U469 , P1_R1138_U468 , P1_R1138_U467 );
nand NAND2_16804 ( P1_R1138_U470 , P1_R1138_U358 , P1_R1138_U93 );
nand NAND2_16805 ( P1_R1138_U471 , P1_R1138_U469 , P1_R1138_U259 );
nand NAND2_16806 ( P1_R1138_U472 , P1_U3074 , P1_R1138_U74 );
nand NAND2_16807 ( P1_R1138_U473 , P1_U3503 , P1_R1138_U75 );
nand NAND2_16808 ( P1_R1138_U474 , P1_U3074 , P1_R1138_U74 );
nand NAND2_16809 ( P1_R1138_U475 , P1_U3503 , P1_R1138_U75 );
nand NAND2_16810 ( P1_R1138_U476 , P1_R1138_U475 , P1_R1138_U474 );
nand NAND2_16811 ( P1_R1138_U477 , P1_R1138_U160 , P1_R1138_U161 );
nand NAND2_16812 ( P1_R1138_U478 , P1_R1138_U255 , P1_R1138_U476 );
nand NAND2_16813 ( P1_R1138_U479 , P1_U3079 , P1_R1138_U72 );
nand NAND2_16814 ( P1_R1138_U480 , P1_U3500 , P1_R1138_U73 );
nand NAND2_16815 ( P1_R1138_U481 , P1_U3079 , P1_R1138_U72 );
nand NAND2_16816 ( P1_R1138_U482 , P1_U3500 , P1_R1138_U73 );
nand NAND2_16817 ( P1_R1138_U483 , P1_R1138_U482 , P1_R1138_U481 );
nand NAND2_16818 ( P1_R1138_U484 , P1_R1138_U162 , P1_R1138_U163 );
nand NAND2_16819 ( P1_R1138_U485 , P1_R1138_U251 , P1_R1138_U483 );
nand NAND2_16820 ( P1_R1138_U486 , P1_U3080 , P1_R1138_U70 );
nand NAND2_16821 ( P1_R1138_U487 , P1_U3497 , P1_R1138_U71 );
nand NAND2_16822 ( P1_R1138_U488 , P1_U3072 , P1_R1138_U65 );
nand NAND2_16823 ( P1_R1138_U489 , P1_U3494 , P1_R1138_U66 );
nand NAND2_16824 ( P1_R1138_U490 , P1_R1138_U489 , P1_R1138_U488 );
nand NAND2_16825 ( P1_R1138_U491 , P1_R1138_U359 , P1_R1138_U94 );
nand NAND2_16826 ( P1_R1138_U492 , P1_R1138_U490 , P1_R1138_U335 );
nand NAND2_16827 ( P1_R1138_U493 , P1_U3063 , P1_R1138_U67 );
nand NAND2_16828 ( P1_R1138_U494 , P1_U3491 , P1_R1138_U68 );
nand NAND2_16829 ( P1_R1138_U495 , P1_R1138_U494 , P1_R1138_U493 );
nand NAND2_16830 ( P1_R1138_U496 , P1_R1138_U360 , P1_R1138_U164 );
nand NAND2_16831 ( P1_R1138_U497 , P1_R1138_U241 , P1_R1138_U495 );
nand NAND2_16832 ( P1_R1138_U498 , P1_U3062 , P1_R1138_U63 );
nand NAND2_16833 ( P1_R1138_U499 , P1_U3488 , P1_R1138_U64 );
nand NAND2_16834 ( P1_R1138_U500 , P1_U3077 , P1_R1138_U30 );
nand NAND2_16835 ( P1_R1138_U501 , P1_U3456 , P1_R1138_U31 );
and AND2_16836 ( P1_R1222_U4 , P1_R1222_U176 , P1_R1222_U175 );
and AND2_16837 ( P1_R1222_U5 , P1_R1222_U177 , P1_R1222_U178 );
and AND2_16838 ( P1_R1222_U6 , P1_R1222_U194 , P1_R1222_U193 );
and AND2_16839 ( P1_R1222_U7 , P1_R1222_U234 , P1_R1222_U233 );
and AND2_16840 ( P1_R1222_U8 , P1_R1222_U243 , P1_R1222_U242 );
and AND2_16841 ( P1_R1222_U9 , P1_R1222_U261 , P1_R1222_U260 );
and AND2_16842 ( P1_R1222_U10 , P1_R1222_U269 , P1_R1222_U268 );
and AND2_16843 ( P1_R1222_U11 , P1_R1222_U348 , P1_R1222_U345 );
and AND2_16844 ( P1_R1222_U12 , P1_R1222_U341 , P1_R1222_U338 );
and AND2_16845 ( P1_R1222_U13 , P1_R1222_U332 , P1_R1222_U329 );
and AND2_16846 ( P1_R1222_U14 , P1_R1222_U323 , P1_R1222_U320 );
and AND2_16847 ( P1_R1222_U15 , P1_R1222_U317 , P1_R1222_U315 );
and AND2_16848 ( P1_R1222_U16 , P1_R1222_U310 , P1_R1222_U307 );
and AND2_16849 ( P1_R1222_U17 , P1_R1222_U232 , P1_R1222_U229 );
and AND2_16850 ( P1_R1222_U18 , P1_R1222_U224 , P1_R1222_U221 );
and AND2_16851 ( P1_R1222_U19 , P1_R1222_U210 , P1_R1222_U207 );
not NOT1_16852 ( P1_R1222_U20 , P1_U3476 );
not NOT1_16853 ( P1_R1222_U21 , P1_U3071 );
not NOT1_16854 ( P1_R1222_U22 , P1_U3070 );
nand NAND2_16855 ( P1_R1222_U23 , P1_U3071 , P1_U3476 );
not NOT1_16856 ( P1_R1222_U24 , P1_U3479 );
not NOT1_16857 ( P1_R1222_U25 , P1_U3470 );
not NOT1_16858 ( P1_R1222_U26 , P1_U3060 );
not NOT1_16859 ( P1_R1222_U27 , P1_U3067 );
not NOT1_16860 ( P1_R1222_U28 , P1_U3464 );
not NOT1_16861 ( P1_R1222_U29 , P1_U3068 );
not NOT1_16862 ( P1_R1222_U30 , P1_U3456 );
not NOT1_16863 ( P1_R1222_U31 , P1_U3077 );
nand NAND2_16864 ( P1_R1222_U32 , P1_U3077 , P1_U3456 );
not NOT1_16865 ( P1_R1222_U33 , P1_U3467 );
not NOT1_16866 ( P1_R1222_U34 , P1_U3064 );
nand NAND2_16867 ( P1_R1222_U35 , P1_U3060 , P1_U3470 );
not NOT1_16868 ( P1_R1222_U36 , P1_U3473 );
not NOT1_16869 ( P1_R1222_U37 , P1_U3482 );
not NOT1_16870 ( P1_R1222_U38 , P1_U3084 );
not NOT1_16871 ( P1_R1222_U39 , P1_U3083 );
not NOT1_16872 ( P1_R1222_U40 , P1_U3485 );
nand NAND2_16873 ( P1_R1222_U41 , P1_R1222_U62 , P1_R1222_U202 );
nand NAND2_16874 ( P1_R1222_U42 , P1_R1222_U118 , P1_R1222_U190 );
nand NAND2_16875 ( P1_R1222_U43 , P1_R1222_U179 , P1_R1222_U180 );
nand NAND2_16876 ( P1_R1222_U44 , P1_U3461 , P1_U3078 );
nand NAND2_16877 ( P1_R1222_U45 , P1_R1222_U122 , P1_R1222_U216 );
nand NAND2_16878 ( P1_R1222_U46 , P1_R1222_U213 , P1_R1222_U212 );
not NOT1_16879 ( P1_R1222_U47 , P1_U4018 );
not NOT1_16880 ( P1_R1222_U48 , P1_U3053 );
not NOT1_16881 ( P1_R1222_U49 , P1_U3057 );
not NOT1_16882 ( P1_R1222_U50 , P1_U4019 );
not NOT1_16883 ( P1_R1222_U51 , P1_U4020 );
not NOT1_16884 ( P1_R1222_U52 , P1_U3058 );
not NOT1_16885 ( P1_R1222_U53 , P1_U4021 );
not NOT1_16886 ( P1_R1222_U54 , P1_U3065 );
not NOT1_16887 ( P1_R1222_U55 , P1_U4024 );
not NOT1_16888 ( P1_R1222_U56 , P1_U3075 );
not NOT1_16889 ( P1_R1222_U57 , P1_U3506 );
not NOT1_16890 ( P1_R1222_U58 , P1_U3073 );
not NOT1_16891 ( P1_R1222_U59 , P1_U3069 );
nand NAND2_16892 ( P1_R1222_U60 , P1_U3073 , P1_U3506 );
not NOT1_16893 ( P1_R1222_U61 , P1_U3509 );
nand NAND2_16894 ( P1_R1222_U62 , P1_U3084 , P1_U3482 );
not NOT1_16895 ( P1_R1222_U63 , P1_U3488 );
not NOT1_16896 ( P1_R1222_U64 , P1_U3062 );
not NOT1_16897 ( P1_R1222_U65 , P1_U3494 );
not NOT1_16898 ( P1_R1222_U66 , P1_U3072 );
not NOT1_16899 ( P1_R1222_U67 , P1_U3491 );
not NOT1_16900 ( P1_R1222_U68 , P1_U3063 );
nand NAND2_16901 ( P1_R1222_U69 , P1_U3063 , P1_U3491 );
not NOT1_16902 ( P1_R1222_U70 , P1_U3497 );
not NOT1_16903 ( P1_R1222_U71 , P1_U3080 );
not NOT1_16904 ( P1_R1222_U72 , P1_U3500 );
not NOT1_16905 ( P1_R1222_U73 , P1_U3079 );
not NOT1_16906 ( P1_R1222_U74 , P1_U3503 );
not NOT1_16907 ( P1_R1222_U75 , P1_U3074 );
not NOT1_16908 ( P1_R1222_U76 , P1_U3512 );
not NOT1_16909 ( P1_R1222_U77 , P1_U3082 );
nand NAND2_16910 ( P1_R1222_U78 , P1_U3082 , P1_U3512 );
not NOT1_16911 ( P1_R1222_U79 , P1_U3514 );
not NOT1_16912 ( P1_R1222_U80 , P1_U3081 );
nand NAND2_16913 ( P1_R1222_U81 , P1_U3081 , P1_U3514 );
not NOT1_16914 ( P1_R1222_U82 , P1_U4025 );
not NOT1_16915 ( P1_R1222_U83 , P1_U4023 );
not NOT1_16916 ( P1_R1222_U84 , P1_U3061 );
not NOT1_16917 ( P1_R1222_U85 , P1_U4022 );
not NOT1_16918 ( P1_R1222_U86 , P1_U3066 );
nand NAND2_16919 ( P1_R1222_U87 , P1_U4019 , P1_U3057 );
not NOT1_16920 ( P1_R1222_U88 , P1_U3054 );
not NOT1_16921 ( P1_R1222_U89 , P1_U4017 );
nand NAND2_16922 ( P1_R1222_U90 , P1_R1222_U303 , P1_R1222_U173 );
not NOT1_16923 ( P1_R1222_U91 , P1_U3076 );
nand NAND2_16924 ( P1_R1222_U92 , P1_R1222_U78 , P1_R1222_U312 );
nand NAND2_16925 ( P1_R1222_U93 , P1_R1222_U258 , P1_R1222_U257 );
nand NAND2_16926 ( P1_R1222_U94 , P1_R1222_U69 , P1_R1222_U334 );
nand NAND2_16927 ( P1_R1222_U95 , P1_R1222_U454 , P1_R1222_U453 );
nand NAND2_16928 ( P1_R1222_U96 , P1_R1222_U501 , P1_R1222_U500 );
nand NAND2_16929 ( P1_R1222_U97 , P1_R1222_U372 , P1_R1222_U371 );
nand NAND2_16930 ( P1_R1222_U98 , P1_R1222_U377 , P1_R1222_U376 );
nand NAND2_16931 ( P1_R1222_U99 , P1_R1222_U384 , P1_R1222_U383 );
nand NAND2_16932 ( P1_R1222_U100 , P1_R1222_U391 , P1_R1222_U390 );
nand NAND2_16933 ( P1_R1222_U101 , P1_R1222_U396 , P1_R1222_U395 );
nand NAND2_16934 ( P1_R1222_U102 , P1_R1222_U405 , P1_R1222_U404 );
nand NAND2_16935 ( P1_R1222_U103 , P1_R1222_U412 , P1_R1222_U411 );
nand NAND2_16936 ( P1_R1222_U104 , P1_R1222_U419 , P1_R1222_U418 );
nand NAND2_16937 ( P1_R1222_U105 , P1_R1222_U426 , P1_R1222_U425 );
nand NAND2_16938 ( P1_R1222_U106 , P1_R1222_U431 , P1_R1222_U430 );
nand NAND2_16939 ( P1_R1222_U107 , P1_R1222_U438 , P1_R1222_U437 );
nand NAND2_16940 ( P1_R1222_U108 , P1_R1222_U445 , P1_R1222_U444 );
nand NAND2_16941 ( P1_R1222_U109 , P1_R1222_U459 , P1_R1222_U458 );
nand NAND2_16942 ( P1_R1222_U110 , P1_R1222_U464 , P1_R1222_U463 );
nand NAND2_16943 ( P1_R1222_U111 , P1_R1222_U471 , P1_R1222_U470 );
nand NAND2_16944 ( P1_R1222_U112 , P1_R1222_U478 , P1_R1222_U477 );
nand NAND2_16945 ( P1_R1222_U113 , P1_R1222_U485 , P1_R1222_U484 );
nand NAND2_16946 ( P1_R1222_U114 , P1_R1222_U492 , P1_R1222_U491 );
nand NAND2_16947 ( P1_R1222_U115 , P1_R1222_U497 , P1_R1222_U496 );
and AND2_16948 ( P1_R1222_U116 , P1_U3464 , P1_U3068 );
and AND2_16949 ( P1_R1222_U117 , P1_R1222_U186 , P1_R1222_U184 );
and AND2_16950 ( P1_R1222_U118 , P1_R1222_U191 , P1_R1222_U189 );
and AND2_16951 ( P1_R1222_U119 , P1_R1222_U198 , P1_R1222_U197 );
and AND3_16952 ( P1_R1222_U120 , P1_R1222_U379 , P1_R1222_U378 , P1_R1222_U23 );
and AND2_16953 ( P1_R1222_U121 , P1_R1222_U209 , P1_R1222_U6 );
and AND2_16954 ( P1_R1222_U122 , P1_R1222_U217 , P1_R1222_U215 );
and AND3_16955 ( P1_R1222_U123 , P1_R1222_U386 , P1_R1222_U385 , P1_R1222_U35 );
and AND2_16956 ( P1_R1222_U124 , P1_R1222_U223 , P1_R1222_U4 );
and AND2_16957 ( P1_R1222_U125 , P1_R1222_U231 , P1_R1222_U178 );
and AND2_16958 ( P1_R1222_U126 , P1_R1222_U201 , P1_R1222_U7 );
and AND2_16959 ( P1_R1222_U127 , P1_R1222_U236 , P1_R1222_U168 );
and AND2_16960 ( P1_R1222_U128 , P1_R1222_U245 , P1_R1222_U169 );
and AND2_16961 ( P1_R1222_U129 , P1_R1222_U265 , P1_R1222_U264 );
and AND2_16962 ( P1_R1222_U130 , P1_R1222_U10 , P1_R1222_U279 );
and AND2_16963 ( P1_R1222_U131 , P1_R1222_U282 , P1_R1222_U277 );
and AND2_16964 ( P1_R1222_U132 , P1_R1222_U298 , P1_R1222_U295 );
and AND2_16965 ( P1_R1222_U133 , P1_R1222_U365 , P1_R1222_U299 );
and AND2_16966 ( P1_R1222_U134 , P1_R1222_U156 , P1_R1222_U275 );
and AND3_16967 ( P1_R1222_U135 , P1_R1222_U466 , P1_R1222_U465 , P1_R1222_U60 );
and AND3_16968 ( P1_R1222_U136 , P1_R1222_U487 , P1_R1222_U486 , P1_R1222_U169 );
and AND2_16969 ( P1_R1222_U137 , P1_R1222_U340 , P1_R1222_U8 );
and AND3_16970 ( P1_R1222_U138 , P1_R1222_U499 , P1_R1222_U498 , P1_R1222_U168 );
and AND2_16971 ( P1_R1222_U139 , P1_R1222_U347 , P1_R1222_U7 );
nand NAND2_16972 ( P1_R1222_U140 , P1_R1222_U119 , P1_R1222_U199 );
nand NAND2_16973 ( P1_R1222_U141 , P1_R1222_U214 , P1_R1222_U226 );
not NOT1_16974 ( P1_R1222_U142 , P1_U3055 );
not NOT1_16975 ( P1_R1222_U143 , P1_U4028 );
and AND2_16976 ( P1_R1222_U144 , P1_R1222_U400 , P1_R1222_U399 );
nand NAND3_16977 ( P1_R1222_U145 , P1_R1222_U301 , P1_R1222_U166 , P1_R1222_U361 );
and AND2_16978 ( P1_R1222_U146 , P1_R1222_U407 , P1_R1222_U406 );
nand NAND3_16979 ( P1_R1222_U147 , P1_R1222_U367 , P1_R1222_U366 , P1_R1222_U133 );
and AND2_16980 ( P1_R1222_U148 , P1_R1222_U414 , P1_R1222_U413 );
nand NAND3_16981 ( P1_R1222_U149 , P1_R1222_U362 , P1_R1222_U296 , P1_R1222_U87 );
and AND2_16982 ( P1_R1222_U150 , P1_R1222_U421 , P1_R1222_U420 );
nand NAND2_16983 ( P1_R1222_U151 , P1_R1222_U290 , P1_R1222_U289 );
and AND2_16984 ( P1_R1222_U152 , P1_R1222_U433 , P1_R1222_U432 );
nand NAND2_16985 ( P1_R1222_U153 , P1_R1222_U286 , P1_R1222_U285 );
and AND2_16986 ( P1_R1222_U154 , P1_R1222_U440 , P1_R1222_U439 );
nand NAND2_16987 ( P1_R1222_U155 , P1_R1222_U131 , P1_R1222_U281 );
and AND2_16988 ( P1_R1222_U156 , P1_R1222_U447 , P1_R1222_U446 );
and AND2_16989 ( P1_R1222_U157 , P1_R1222_U452 , P1_R1222_U451 );
nand NAND2_16990 ( P1_R1222_U158 , P1_R1222_U44 , P1_R1222_U324 );
nand NAND2_16991 ( P1_R1222_U159 , P1_R1222_U129 , P1_R1222_U266 );
and AND2_16992 ( P1_R1222_U160 , P1_R1222_U473 , P1_R1222_U472 );
nand NAND2_16993 ( P1_R1222_U161 , P1_R1222_U254 , P1_R1222_U253 );
and AND2_16994 ( P1_R1222_U162 , P1_R1222_U480 , P1_R1222_U479 );
nand NAND2_16995 ( P1_R1222_U163 , P1_R1222_U250 , P1_R1222_U249 );
nand NAND2_16996 ( P1_R1222_U164 , P1_R1222_U240 , P1_R1222_U239 );
nand NAND2_16997 ( P1_R1222_U165 , P1_R1222_U364 , P1_R1222_U363 );
nand NAND2_16998 ( P1_R1222_U166 , P1_U3054 , P1_R1222_U147 );
not NOT1_16999 ( P1_R1222_U167 , P1_R1222_U35 );
nand NAND2_17000 ( P1_R1222_U168 , P1_U3485 , P1_U3083 );
nand NAND2_17001 ( P1_R1222_U169 , P1_U3072 , P1_U3494 );
nand NAND2_17002 ( P1_R1222_U170 , P1_U3058 , P1_U4020 );
not NOT1_17003 ( P1_R1222_U171 , P1_R1222_U69 );
not NOT1_17004 ( P1_R1222_U172 , P1_R1222_U78 );
nand NAND2_17005 ( P1_R1222_U173 , P1_U3065 , P1_U4021 );
not NOT1_17006 ( P1_R1222_U174 , P1_R1222_U62 );
or OR2_17007 ( P1_R1222_U175 , P1_U3067 , P1_U3473 );
or OR2_17008 ( P1_R1222_U176 , P1_U3060 , P1_U3470 );
or OR2_17009 ( P1_R1222_U177 , P1_U3467 , P1_U3064 );
or OR2_17010 ( P1_R1222_U178 , P1_U3464 , P1_U3068 );
not NOT1_17011 ( P1_R1222_U179 , P1_R1222_U32 );
or OR2_17012 ( P1_R1222_U180 , P1_U3461 , P1_U3078 );
not NOT1_17013 ( P1_R1222_U181 , P1_R1222_U43 );
not NOT1_17014 ( P1_R1222_U182 , P1_R1222_U44 );
nand NAND2_17015 ( P1_R1222_U183 , P1_R1222_U43 , P1_R1222_U44 );
nand NAND2_17016 ( P1_R1222_U184 , P1_R1222_U116 , P1_R1222_U177 );
nand NAND2_17017 ( P1_R1222_U185 , P1_R1222_U5 , P1_R1222_U183 );
nand NAND2_17018 ( P1_R1222_U186 , P1_U3064 , P1_U3467 );
nand NAND2_17019 ( P1_R1222_U187 , P1_R1222_U117 , P1_R1222_U185 );
nand NAND2_17020 ( P1_R1222_U188 , P1_R1222_U36 , P1_R1222_U35 );
nand NAND2_17021 ( P1_R1222_U189 , P1_U3067 , P1_R1222_U188 );
nand NAND2_17022 ( P1_R1222_U190 , P1_R1222_U4 , P1_R1222_U187 );
nand NAND2_17023 ( P1_R1222_U191 , P1_U3473 , P1_R1222_U167 );
not NOT1_17024 ( P1_R1222_U192 , P1_R1222_U42 );
or OR2_17025 ( P1_R1222_U193 , P1_U3070 , P1_U3479 );
or OR2_17026 ( P1_R1222_U194 , P1_U3071 , P1_U3476 );
not NOT1_17027 ( P1_R1222_U195 , P1_R1222_U23 );
nand NAND2_17028 ( P1_R1222_U196 , P1_R1222_U24 , P1_R1222_U23 );
nand NAND2_17029 ( P1_R1222_U197 , P1_U3070 , P1_R1222_U196 );
nand NAND2_17030 ( P1_R1222_U198 , P1_U3479 , P1_R1222_U195 );
nand NAND2_17031 ( P1_R1222_U199 , P1_R1222_U6 , P1_R1222_U42 );
not NOT1_17032 ( P1_R1222_U200 , P1_R1222_U140 );
or OR2_17033 ( P1_R1222_U201 , P1_U3482 , P1_U3084 );
nand NAND2_17034 ( P1_R1222_U202 , P1_R1222_U201 , P1_R1222_U140 );
not NOT1_17035 ( P1_R1222_U203 , P1_R1222_U41 );
or OR2_17036 ( P1_R1222_U204 , P1_U3083 , P1_U3485 );
or OR2_17037 ( P1_R1222_U205 , P1_U3476 , P1_U3071 );
nand NAND2_17038 ( P1_R1222_U206 , P1_R1222_U205 , P1_R1222_U42 );
nand NAND2_17039 ( P1_R1222_U207 , P1_R1222_U120 , P1_R1222_U206 );
nand NAND2_17040 ( P1_R1222_U208 , P1_R1222_U192 , P1_R1222_U23 );
nand NAND2_17041 ( P1_R1222_U209 , P1_U3479 , P1_U3070 );
nand NAND2_17042 ( P1_R1222_U210 , P1_R1222_U121 , P1_R1222_U208 );
or OR2_17043 ( P1_R1222_U211 , P1_U3071 , P1_U3476 );
nand NAND2_17044 ( P1_R1222_U212 , P1_R1222_U182 , P1_R1222_U178 );
nand NAND2_17045 ( P1_R1222_U213 , P1_U3068 , P1_U3464 );
not NOT1_17046 ( P1_R1222_U214 , P1_R1222_U46 );
nand NAND2_17047 ( P1_R1222_U215 , P1_R1222_U181 , P1_R1222_U5 );
nand NAND2_17048 ( P1_R1222_U216 , P1_R1222_U46 , P1_R1222_U177 );
nand NAND2_17049 ( P1_R1222_U217 , P1_U3064 , P1_U3467 );
not NOT1_17050 ( P1_R1222_U218 , P1_R1222_U45 );
or OR2_17051 ( P1_R1222_U219 , P1_U3470 , P1_U3060 );
nand NAND2_17052 ( P1_R1222_U220 , P1_R1222_U219 , P1_R1222_U45 );
nand NAND2_17053 ( P1_R1222_U221 , P1_R1222_U123 , P1_R1222_U220 );
nand NAND2_17054 ( P1_R1222_U222 , P1_R1222_U218 , P1_R1222_U35 );
nand NAND2_17055 ( P1_R1222_U223 , P1_U3473 , P1_U3067 );
nand NAND2_17056 ( P1_R1222_U224 , P1_R1222_U124 , P1_R1222_U222 );
or OR2_17057 ( P1_R1222_U225 , P1_U3060 , P1_U3470 );
nand NAND2_17058 ( P1_R1222_U226 , P1_R1222_U181 , P1_R1222_U178 );
not NOT1_17059 ( P1_R1222_U227 , P1_R1222_U141 );
nand NAND2_17060 ( P1_R1222_U228 , P1_U3064 , P1_U3467 );
nand NAND4_17061 ( P1_R1222_U229 , P1_R1222_U398 , P1_R1222_U397 , P1_R1222_U44 , P1_R1222_U43 );
nand NAND2_17062 ( P1_R1222_U230 , P1_R1222_U44 , P1_R1222_U43 );
nand NAND2_17063 ( P1_R1222_U231 , P1_U3068 , P1_U3464 );
nand NAND2_17064 ( P1_R1222_U232 , P1_R1222_U125 , P1_R1222_U230 );
or OR2_17065 ( P1_R1222_U233 , P1_U3083 , P1_U3485 );
or OR2_17066 ( P1_R1222_U234 , P1_U3062 , P1_U3488 );
nand NAND2_17067 ( P1_R1222_U235 , P1_R1222_U174 , P1_R1222_U7 );
nand NAND2_17068 ( P1_R1222_U236 , P1_U3062 , P1_U3488 );
nand NAND2_17069 ( P1_R1222_U237 , P1_R1222_U127 , P1_R1222_U235 );
or OR2_17070 ( P1_R1222_U238 , P1_U3488 , P1_U3062 );
nand NAND2_17071 ( P1_R1222_U239 , P1_R1222_U126 , P1_R1222_U140 );
nand NAND2_17072 ( P1_R1222_U240 , P1_R1222_U238 , P1_R1222_U237 );
not NOT1_17073 ( P1_R1222_U241 , P1_R1222_U164 );
or OR2_17074 ( P1_R1222_U242 , P1_U3080 , P1_U3497 );
or OR2_17075 ( P1_R1222_U243 , P1_U3072 , P1_U3494 );
nand NAND2_17076 ( P1_R1222_U244 , P1_R1222_U171 , P1_R1222_U8 );
nand NAND2_17077 ( P1_R1222_U245 , P1_U3080 , P1_U3497 );
nand NAND2_17078 ( P1_R1222_U246 , P1_R1222_U128 , P1_R1222_U244 );
or OR2_17079 ( P1_R1222_U247 , P1_U3491 , P1_U3063 );
or OR2_17080 ( P1_R1222_U248 , P1_U3497 , P1_U3080 );
nand NAND3_17081 ( P1_R1222_U249 , P1_R1222_U247 , P1_R1222_U164 , P1_R1222_U8 );
nand NAND2_17082 ( P1_R1222_U250 , P1_R1222_U248 , P1_R1222_U246 );
not NOT1_17083 ( P1_R1222_U251 , P1_R1222_U163 );
or OR2_17084 ( P1_R1222_U252 , P1_U3500 , P1_U3079 );
nand NAND2_17085 ( P1_R1222_U253 , P1_R1222_U252 , P1_R1222_U163 );
nand NAND2_17086 ( P1_R1222_U254 , P1_U3079 , P1_U3500 );
not NOT1_17087 ( P1_R1222_U255 , P1_R1222_U161 );
or OR2_17088 ( P1_R1222_U256 , P1_U3503 , P1_U3074 );
nand NAND2_17089 ( P1_R1222_U257 , P1_R1222_U256 , P1_R1222_U161 );
nand NAND2_17090 ( P1_R1222_U258 , P1_U3074 , P1_U3503 );
not NOT1_17091 ( P1_R1222_U259 , P1_R1222_U93 );
or OR2_17092 ( P1_R1222_U260 , P1_U3069 , P1_U3509 );
or OR2_17093 ( P1_R1222_U261 , P1_U3073 , P1_U3506 );
not NOT1_17094 ( P1_R1222_U262 , P1_R1222_U60 );
nand NAND2_17095 ( P1_R1222_U263 , P1_R1222_U61 , P1_R1222_U60 );
nand NAND2_17096 ( P1_R1222_U264 , P1_U3069 , P1_R1222_U263 );
nand NAND2_17097 ( P1_R1222_U265 , P1_U3509 , P1_R1222_U262 );
nand NAND2_17098 ( P1_R1222_U266 , P1_R1222_U9 , P1_R1222_U93 );
not NOT1_17099 ( P1_R1222_U267 , P1_R1222_U159 );
or OR2_17100 ( P1_R1222_U268 , P1_U3076 , P1_U4025 );
or OR2_17101 ( P1_R1222_U269 , P1_U3081 , P1_U3514 );
or OR2_17102 ( P1_R1222_U270 , P1_U3075 , P1_U4024 );
not NOT1_17103 ( P1_R1222_U271 , P1_R1222_U81 );
nand NAND2_17104 ( P1_R1222_U272 , P1_U4025 , P1_R1222_U271 );
nand NAND2_17105 ( P1_R1222_U273 , P1_R1222_U272 , P1_R1222_U91 );
nand NAND2_17106 ( P1_R1222_U274 , P1_R1222_U81 , P1_R1222_U82 );
nand NAND2_17107 ( P1_R1222_U275 , P1_R1222_U274 , P1_R1222_U273 );
nand NAND2_17108 ( P1_R1222_U276 , P1_R1222_U172 , P1_R1222_U10 );
nand NAND2_17109 ( P1_R1222_U277 , P1_U3075 , P1_U4024 );
nand NAND2_17110 ( P1_R1222_U278 , P1_R1222_U275 , P1_R1222_U276 );
or OR2_17111 ( P1_R1222_U279 , P1_U3512 , P1_U3082 );
or OR2_17112 ( P1_R1222_U280 , P1_U4024 , P1_U3075 );
nand NAND3_17113 ( P1_R1222_U281 , P1_R1222_U270 , P1_R1222_U159 , P1_R1222_U130 );
nand NAND2_17114 ( P1_R1222_U282 , P1_R1222_U280 , P1_R1222_U278 );
not NOT1_17115 ( P1_R1222_U283 , P1_R1222_U155 );
or OR2_17116 ( P1_R1222_U284 , P1_U4023 , P1_U3061 );
nand NAND2_17117 ( P1_R1222_U285 , P1_R1222_U284 , P1_R1222_U155 );
nand NAND2_17118 ( P1_R1222_U286 , P1_U3061 , P1_U4023 );
not NOT1_17119 ( P1_R1222_U287 , P1_R1222_U153 );
or OR2_17120 ( P1_R1222_U288 , P1_U4022 , P1_U3066 );
nand NAND2_17121 ( P1_R1222_U289 , P1_R1222_U288 , P1_R1222_U153 );
nand NAND2_17122 ( P1_R1222_U290 , P1_U3066 , P1_U4022 );
not NOT1_17123 ( P1_R1222_U291 , P1_R1222_U151 );
or OR2_17124 ( P1_R1222_U292 , P1_U3058 , P1_U4020 );
nand NAND2_17125 ( P1_R1222_U293 , P1_R1222_U173 , P1_R1222_U170 );
not NOT1_17126 ( P1_R1222_U294 , P1_R1222_U87 );
or OR2_17127 ( P1_R1222_U295 , P1_U4021 , P1_U3065 );
nand NAND3_17128 ( P1_R1222_U296 , P1_R1222_U151 , P1_R1222_U295 , P1_R1222_U165 );
not NOT1_17129 ( P1_R1222_U297 , P1_R1222_U149 );
or OR2_17130 ( P1_R1222_U298 , P1_U4018 , P1_U3053 );
nand NAND2_17131 ( P1_R1222_U299 , P1_U3053 , P1_U4018 );
not NOT1_17132 ( P1_R1222_U300 , P1_R1222_U147 );
nand NAND2_17133 ( P1_R1222_U301 , P1_U4017 , P1_R1222_U147 );
not NOT1_17134 ( P1_R1222_U302 , P1_R1222_U145 );
nand NAND2_17135 ( P1_R1222_U303 , P1_R1222_U295 , P1_R1222_U151 );
not NOT1_17136 ( P1_R1222_U304 , P1_R1222_U90 );
or OR2_17137 ( P1_R1222_U305 , P1_U4020 , P1_U3058 );
nand NAND2_17138 ( P1_R1222_U306 , P1_R1222_U305 , P1_R1222_U90 );
nand NAND3_17139 ( P1_R1222_U307 , P1_R1222_U306 , P1_R1222_U170 , P1_R1222_U150 );
nand NAND2_17140 ( P1_R1222_U308 , P1_R1222_U304 , P1_R1222_U170 );
nand NAND2_17141 ( P1_R1222_U309 , P1_U4019 , P1_U3057 );
nand NAND3_17142 ( P1_R1222_U310 , P1_R1222_U308 , P1_R1222_U309 , P1_R1222_U165 );
or OR2_17143 ( P1_R1222_U311 , P1_U3058 , P1_U4020 );
nand NAND2_17144 ( P1_R1222_U312 , P1_R1222_U279 , P1_R1222_U159 );
not NOT1_17145 ( P1_R1222_U313 , P1_R1222_U92 );
nand NAND2_17146 ( P1_R1222_U314 , P1_R1222_U10 , P1_R1222_U92 );
nand NAND2_17147 ( P1_R1222_U315 , P1_R1222_U134 , P1_R1222_U314 );
nand NAND2_17148 ( P1_R1222_U316 , P1_R1222_U314 , P1_R1222_U275 );
nand NAND2_17149 ( P1_R1222_U317 , P1_R1222_U450 , P1_R1222_U316 );
or OR2_17150 ( P1_R1222_U318 , P1_U3514 , P1_U3081 );
nand NAND2_17151 ( P1_R1222_U319 , P1_R1222_U318 , P1_R1222_U92 );
nand NAND3_17152 ( P1_R1222_U320 , P1_R1222_U319 , P1_R1222_U81 , P1_R1222_U157 );
nand NAND2_17153 ( P1_R1222_U321 , P1_R1222_U313 , P1_R1222_U81 );
nand NAND2_17154 ( P1_R1222_U322 , P1_U3076 , P1_U4025 );
nand NAND3_17155 ( P1_R1222_U323 , P1_R1222_U322 , P1_R1222_U321 , P1_R1222_U10 );
or OR2_17156 ( P1_R1222_U324 , P1_U3461 , P1_U3078 );
not NOT1_17157 ( P1_R1222_U325 , P1_R1222_U158 );
or OR2_17158 ( P1_R1222_U326 , P1_U3081 , P1_U3514 );
or OR2_17159 ( P1_R1222_U327 , P1_U3506 , P1_U3073 );
nand NAND2_17160 ( P1_R1222_U328 , P1_R1222_U327 , P1_R1222_U93 );
nand NAND2_17161 ( P1_R1222_U329 , P1_R1222_U135 , P1_R1222_U328 );
nand NAND2_17162 ( P1_R1222_U330 , P1_R1222_U259 , P1_R1222_U60 );
nand NAND2_17163 ( P1_R1222_U331 , P1_U3509 , P1_U3069 );
nand NAND3_17164 ( P1_R1222_U332 , P1_R1222_U331 , P1_R1222_U330 , P1_R1222_U9 );
or OR2_17165 ( P1_R1222_U333 , P1_U3073 , P1_U3506 );
nand NAND2_17166 ( P1_R1222_U334 , P1_R1222_U247 , P1_R1222_U164 );
not NOT1_17167 ( P1_R1222_U335 , P1_R1222_U94 );
or OR2_17168 ( P1_R1222_U336 , P1_U3494 , P1_U3072 );
nand NAND2_17169 ( P1_R1222_U337 , P1_R1222_U336 , P1_R1222_U94 );
nand NAND2_17170 ( P1_R1222_U338 , P1_R1222_U136 , P1_R1222_U337 );
nand NAND2_17171 ( P1_R1222_U339 , P1_R1222_U335 , P1_R1222_U169 );
nand NAND2_17172 ( P1_R1222_U340 , P1_U3080 , P1_U3497 );
nand NAND2_17173 ( P1_R1222_U341 , P1_R1222_U137 , P1_R1222_U339 );
or OR2_17174 ( P1_R1222_U342 , P1_U3072 , P1_U3494 );
or OR2_17175 ( P1_R1222_U343 , P1_U3485 , P1_U3083 );
nand NAND2_17176 ( P1_R1222_U344 , P1_R1222_U343 , P1_R1222_U41 );
nand NAND2_17177 ( P1_R1222_U345 , P1_R1222_U138 , P1_R1222_U344 );
nand NAND2_17178 ( P1_R1222_U346 , P1_R1222_U203 , P1_R1222_U168 );
nand NAND2_17179 ( P1_R1222_U347 , P1_U3062 , P1_U3488 );
nand NAND2_17180 ( P1_R1222_U348 , P1_R1222_U139 , P1_R1222_U346 );
nand NAND2_17181 ( P1_R1222_U349 , P1_R1222_U204 , P1_R1222_U168 );
nand NAND2_17182 ( P1_R1222_U350 , P1_R1222_U201 , P1_R1222_U62 );
nand NAND2_17183 ( P1_R1222_U351 , P1_R1222_U211 , P1_R1222_U23 );
nand NAND2_17184 ( P1_R1222_U352 , P1_R1222_U225 , P1_R1222_U35 );
nand NAND2_17185 ( P1_R1222_U353 , P1_R1222_U228 , P1_R1222_U177 );
nand NAND2_17186 ( P1_R1222_U354 , P1_R1222_U311 , P1_R1222_U170 );
nand NAND2_17187 ( P1_R1222_U355 , P1_R1222_U295 , P1_R1222_U173 );
nand NAND2_17188 ( P1_R1222_U356 , P1_R1222_U326 , P1_R1222_U81 );
nand NAND2_17189 ( P1_R1222_U357 , P1_R1222_U279 , P1_R1222_U78 );
nand NAND2_17190 ( P1_R1222_U358 , P1_R1222_U333 , P1_R1222_U60 );
nand NAND2_17191 ( P1_R1222_U359 , P1_R1222_U342 , P1_R1222_U169 );
nand NAND2_17192 ( P1_R1222_U360 , P1_R1222_U247 , P1_R1222_U69 );
nand NAND2_17193 ( P1_R1222_U361 , P1_U4017 , P1_U3054 );
nand NAND2_17194 ( P1_R1222_U362 , P1_R1222_U293 , P1_R1222_U165 );
nand NAND2_17195 ( P1_R1222_U363 , P1_U3057 , P1_R1222_U292 );
nand NAND2_17196 ( P1_R1222_U364 , P1_U4019 , P1_R1222_U292 );
nand NAND3_17197 ( P1_R1222_U365 , P1_R1222_U293 , P1_R1222_U165 , P1_R1222_U298 );
nand NAND3_17198 ( P1_R1222_U366 , P1_R1222_U151 , P1_R1222_U165 , P1_R1222_U132 );
nand NAND2_17199 ( P1_R1222_U367 , P1_R1222_U294 , P1_R1222_U298 );
nand NAND2_17200 ( P1_R1222_U368 , P1_U3083 , P1_R1222_U40 );
nand NAND2_17201 ( P1_R1222_U369 , P1_U3485 , P1_R1222_U39 );
nand NAND2_17202 ( P1_R1222_U370 , P1_R1222_U369 , P1_R1222_U368 );
nand NAND2_17203 ( P1_R1222_U371 , P1_R1222_U349 , P1_R1222_U41 );
nand NAND2_17204 ( P1_R1222_U372 , P1_R1222_U370 , P1_R1222_U203 );
nand NAND2_17205 ( P1_R1222_U373 , P1_U3084 , P1_R1222_U37 );
nand NAND2_17206 ( P1_R1222_U374 , P1_U3482 , P1_R1222_U38 );
nand NAND2_17207 ( P1_R1222_U375 , P1_R1222_U374 , P1_R1222_U373 );
nand NAND2_17208 ( P1_R1222_U376 , P1_R1222_U350 , P1_R1222_U140 );
nand NAND2_17209 ( P1_R1222_U377 , P1_R1222_U200 , P1_R1222_U375 );
nand NAND2_17210 ( P1_R1222_U378 , P1_U3070 , P1_R1222_U24 );
nand NAND2_17211 ( P1_R1222_U379 , P1_U3479 , P1_R1222_U22 );
nand NAND2_17212 ( P1_R1222_U380 , P1_U3071 , P1_R1222_U20 );
nand NAND2_17213 ( P1_R1222_U381 , P1_U3476 , P1_R1222_U21 );
nand NAND2_17214 ( P1_R1222_U382 , P1_R1222_U381 , P1_R1222_U380 );
nand NAND2_17215 ( P1_R1222_U383 , P1_R1222_U351 , P1_R1222_U42 );
nand NAND2_17216 ( P1_R1222_U384 , P1_R1222_U382 , P1_R1222_U192 );
nand NAND2_17217 ( P1_R1222_U385 , P1_U3067 , P1_R1222_U36 );
nand NAND2_17218 ( P1_R1222_U386 , P1_U3473 , P1_R1222_U27 );
nand NAND2_17219 ( P1_R1222_U387 , P1_U3060 , P1_R1222_U25 );
nand NAND2_17220 ( P1_R1222_U388 , P1_U3470 , P1_R1222_U26 );
nand NAND2_17221 ( P1_R1222_U389 , P1_R1222_U388 , P1_R1222_U387 );
nand NAND2_17222 ( P1_R1222_U390 , P1_R1222_U352 , P1_R1222_U45 );
nand NAND2_17223 ( P1_R1222_U391 , P1_R1222_U389 , P1_R1222_U218 );
nand NAND2_17224 ( P1_R1222_U392 , P1_U3064 , P1_R1222_U33 );
nand NAND2_17225 ( P1_R1222_U393 , P1_U3467 , P1_R1222_U34 );
nand NAND2_17226 ( P1_R1222_U394 , P1_R1222_U393 , P1_R1222_U392 );
nand NAND2_17227 ( P1_R1222_U395 , P1_R1222_U353 , P1_R1222_U141 );
nand NAND2_17228 ( P1_R1222_U396 , P1_R1222_U227 , P1_R1222_U394 );
nand NAND2_17229 ( P1_R1222_U397 , P1_U3068 , P1_R1222_U28 );
nand NAND2_17230 ( P1_R1222_U398 , P1_U3464 , P1_R1222_U29 );
nand NAND2_17231 ( P1_R1222_U399 , P1_U3055 , P1_R1222_U143 );
nand NAND2_17232 ( P1_R1222_U400 , P1_U4028 , P1_R1222_U142 );
nand NAND2_17233 ( P1_R1222_U401 , P1_U3055 , P1_R1222_U143 );
nand NAND2_17234 ( P1_R1222_U402 , P1_U4028 , P1_R1222_U142 );
nand NAND2_17235 ( P1_R1222_U403 , P1_R1222_U402 , P1_R1222_U401 );
nand NAND2_17236 ( P1_R1222_U404 , P1_R1222_U144 , P1_R1222_U145 );
nand NAND2_17237 ( P1_R1222_U405 , P1_R1222_U302 , P1_R1222_U403 );
nand NAND2_17238 ( P1_R1222_U406 , P1_U3054 , P1_R1222_U89 );
nand NAND2_17239 ( P1_R1222_U407 , P1_U4017 , P1_R1222_U88 );
nand NAND2_17240 ( P1_R1222_U408 , P1_U3054 , P1_R1222_U89 );
nand NAND2_17241 ( P1_R1222_U409 , P1_U4017 , P1_R1222_U88 );
nand NAND2_17242 ( P1_R1222_U410 , P1_R1222_U409 , P1_R1222_U408 );
nand NAND2_17243 ( P1_R1222_U411 , P1_R1222_U146 , P1_R1222_U147 );
nand NAND2_17244 ( P1_R1222_U412 , P1_R1222_U300 , P1_R1222_U410 );
nand NAND2_17245 ( P1_R1222_U413 , P1_U3053 , P1_R1222_U47 );
nand NAND2_17246 ( P1_R1222_U414 , P1_U4018 , P1_R1222_U48 );
nand NAND2_17247 ( P1_R1222_U415 , P1_U3053 , P1_R1222_U47 );
nand NAND2_17248 ( P1_R1222_U416 , P1_U4018 , P1_R1222_U48 );
nand NAND2_17249 ( P1_R1222_U417 , P1_R1222_U416 , P1_R1222_U415 );
nand NAND2_17250 ( P1_R1222_U418 , P1_R1222_U148 , P1_R1222_U149 );
nand NAND2_17251 ( P1_R1222_U419 , P1_R1222_U297 , P1_R1222_U417 );
nand NAND2_17252 ( P1_R1222_U420 , P1_U3057 , P1_R1222_U50 );
nand NAND2_17253 ( P1_R1222_U421 , P1_U4019 , P1_R1222_U49 );
nand NAND2_17254 ( P1_R1222_U422 , P1_U3058 , P1_R1222_U51 );
nand NAND2_17255 ( P1_R1222_U423 , P1_U4020 , P1_R1222_U52 );
nand NAND2_17256 ( P1_R1222_U424 , P1_R1222_U423 , P1_R1222_U422 );
nand NAND2_17257 ( P1_R1222_U425 , P1_R1222_U354 , P1_R1222_U90 );
nand NAND2_17258 ( P1_R1222_U426 , P1_R1222_U424 , P1_R1222_U304 );
nand NAND2_17259 ( P1_R1222_U427 , P1_U3065 , P1_R1222_U53 );
nand NAND2_17260 ( P1_R1222_U428 , P1_U4021 , P1_R1222_U54 );
nand NAND2_17261 ( P1_R1222_U429 , P1_R1222_U428 , P1_R1222_U427 );
nand NAND2_17262 ( P1_R1222_U430 , P1_R1222_U355 , P1_R1222_U151 );
nand NAND2_17263 ( P1_R1222_U431 , P1_R1222_U291 , P1_R1222_U429 );
nand NAND2_17264 ( P1_R1222_U432 , P1_U3066 , P1_R1222_U85 );
nand NAND2_17265 ( P1_R1222_U433 , P1_U4022 , P1_R1222_U86 );
nand NAND2_17266 ( P1_R1222_U434 , P1_U3066 , P1_R1222_U85 );
nand NAND2_17267 ( P1_R1222_U435 , P1_U4022 , P1_R1222_U86 );
nand NAND2_17268 ( P1_R1222_U436 , P1_R1222_U435 , P1_R1222_U434 );
nand NAND2_17269 ( P1_R1222_U437 , P1_R1222_U152 , P1_R1222_U153 );
nand NAND2_17270 ( P1_R1222_U438 , P1_R1222_U287 , P1_R1222_U436 );
nand NAND2_17271 ( P1_R1222_U439 , P1_U3061 , P1_R1222_U83 );
nand NAND2_17272 ( P1_R1222_U440 , P1_U4023 , P1_R1222_U84 );
nand NAND2_17273 ( P1_R1222_U441 , P1_U3061 , P1_R1222_U83 );
nand NAND2_17274 ( P1_R1222_U442 , P1_U4023 , P1_R1222_U84 );
nand NAND2_17275 ( P1_R1222_U443 , P1_R1222_U442 , P1_R1222_U441 );
nand NAND2_17276 ( P1_R1222_U444 , P1_R1222_U154 , P1_R1222_U155 );
nand NAND2_17277 ( P1_R1222_U445 , P1_R1222_U283 , P1_R1222_U443 );
nand NAND2_17278 ( P1_R1222_U446 , P1_U3075 , P1_R1222_U55 );
nand NAND2_17279 ( P1_R1222_U447 , P1_U4024 , P1_R1222_U56 );
nand NAND2_17280 ( P1_R1222_U448 , P1_U3075 , P1_R1222_U55 );
nand NAND2_17281 ( P1_R1222_U449 , P1_U4024 , P1_R1222_U56 );
nand NAND2_17282 ( P1_R1222_U450 , P1_R1222_U449 , P1_R1222_U448 );
nand NAND2_17283 ( P1_R1222_U451 , P1_U3076 , P1_R1222_U82 );
nand NAND2_17284 ( P1_R1222_U452 , P1_U4025 , P1_R1222_U91 );
nand NAND2_17285 ( P1_R1222_U453 , P1_R1222_U179 , P1_R1222_U158 );
nand NAND2_17286 ( P1_R1222_U454 , P1_R1222_U325 , P1_R1222_U32 );
nand NAND2_17287 ( P1_R1222_U455 , P1_U3081 , P1_R1222_U79 );
nand NAND2_17288 ( P1_R1222_U456 , P1_U3514 , P1_R1222_U80 );
nand NAND2_17289 ( P1_R1222_U457 , P1_R1222_U456 , P1_R1222_U455 );
nand NAND2_17290 ( P1_R1222_U458 , P1_R1222_U356 , P1_R1222_U92 );
nand NAND2_17291 ( P1_R1222_U459 , P1_R1222_U457 , P1_R1222_U313 );
nand NAND2_17292 ( P1_R1222_U460 , P1_U3082 , P1_R1222_U76 );
nand NAND2_17293 ( P1_R1222_U461 , P1_U3512 , P1_R1222_U77 );
nand NAND2_17294 ( P1_R1222_U462 , P1_R1222_U461 , P1_R1222_U460 );
nand NAND2_17295 ( P1_R1222_U463 , P1_R1222_U357 , P1_R1222_U159 );
nand NAND2_17296 ( P1_R1222_U464 , P1_R1222_U267 , P1_R1222_U462 );
nand NAND2_17297 ( P1_R1222_U465 , P1_U3069 , P1_R1222_U61 );
nand NAND2_17298 ( P1_R1222_U466 , P1_U3509 , P1_R1222_U59 );
nand NAND2_17299 ( P1_R1222_U467 , P1_U3073 , P1_R1222_U57 );
nand NAND2_17300 ( P1_R1222_U468 , P1_U3506 , P1_R1222_U58 );
nand NAND2_17301 ( P1_R1222_U469 , P1_R1222_U468 , P1_R1222_U467 );
nand NAND2_17302 ( P1_R1222_U470 , P1_R1222_U358 , P1_R1222_U93 );
nand NAND2_17303 ( P1_R1222_U471 , P1_R1222_U469 , P1_R1222_U259 );
nand NAND2_17304 ( P1_R1222_U472 , P1_U3074 , P1_R1222_U74 );
nand NAND2_17305 ( P1_R1222_U473 , P1_U3503 , P1_R1222_U75 );
nand NAND2_17306 ( P1_R1222_U474 , P1_U3074 , P1_R1222_U74 );
nand NAND2_17307 ( P1_R1222_U475 , P1_U3503 , P1_R1222_U75 );
nand NAND2_17308 ( P1_R1222_U476 , P1_R1222_U475 , P1_R1222_U474 );
nand NAND2_17309 ( P1_R1222_U477 , P1_R1222_U160 , P1_R1222_U161 );
nand NAND2_17310 ( P1_R1222_U478 , P1_R1222_U255 , P1_R1222_U476 );
nand NAND2_17311 ( P1_R1222_U479 , P1_U3079 , P1_R1222_U72 );
nand NAND2_17312 ( P1_R1222_U480 , P1_U3500 , P1_R1222_U73 );
nand NAND2_17313 ( P1_R1222_U481 , P1_U3079 , P1_R1222_U72 );
nand NAND2_17314 ( P1_R1222_U482 , P1_U3500 , P1_R1222_U73 );
nand NAND2_17315 ( P1_R1222_U483 , P1_R1222_U482 , P1_R1222_U481 );
nand NAND2_17316 ( P1_R1222_U484 , P1_R1222_U162 , P1_R1222_U163 );
nand NAND2_17317 ( P1_R1222_U485 , P1_R1222_U251 , P1_R1222_U483 );
nand NAND2_17318 ( P1_R1222_U486 , P1_U3080 , P1_R1222_U70 );
nand NAND2_17319 ( P1_R1222_U487 , P1_U3497 , P1_R1222_U71 );
nand NAND2_17320 ( P1_R1222_U488 , P1_U3072 , P1_R1222_U65 );
nand NAND2_17321 ( P1_R1222_U489 , P1_U3494 , P1_R1222_U66 );
nand NAND2_17322 ( P1_R1222_U490 , P1_R1222_U489 , P1_R1222_U488 );
nand NAND2_17323 ( P1_R1222_U491 , P1_R1222_U359 , P1_R1222_U94 );
nand NAND2_17324 ( P1_R1222_U492 , P1_R1222_U490 , P1_R1222_U335 );
nand NAND2_17325 ( P1_R1222_U493 , P1_U3063 , P1_R1222_U67 );
nand NAND2_17326 ( P1_R1222_U494 , P1_U3491 , P1_R1222_U68 );
nand NAND2_17327 ( P1_R1222_U495 , P1_R1222_U494 , P1_R1222_U493 );
nand NAND2_17328 ( P1_R1222_U496 , P1_R1222_U360 , P1_R1222_U164 );
nand NAND2_17329 ( P1_R1222_U497 , P1_R1222_U241 , P1_R1222_U495 );
nand NAND2_17330 ( P1_R1222_U498 , P1_U3062 , P1_R1222_U63 );
nand NAND2_17331 ( P1_R1222_U499 , P1_U3488 , P1_R1222_U64 );
nand NAND2_17332 ( P1_R1222_U500 , P1_U3077 , P1_R1222_U30 );
nand NAND2_17333 ( P1_R1222_U501 , P1_U3456 , P1_R1222_U31 );
not NOT1_17334 ( P2_ADD_1119_U4 , P2_REG3_REG_3_ );
and AND2_17335 ( P2_ADD_1119_U5 , P2_ADD_1119_U78 , P2_ADD_1119_U106 );
not NOT1_17336 ( P2_ADD_1119_U6 , P2_REG3_REG_5_ );
not NOT1_17337 ( P2_ADD_1119_U7 , P2_REG3_REG_4_ );
nand NAND3_17338 ( P2_ADD_1119_U8 , P2_REG3_REG_5_ , P2_REG3_REG_3_ , P2_REG3_REG_4_ );
not NOT1_17339 ( P2_ADD_1119_U9 , P2_REG3_REG_7_ );
not NOT1_17340 ( P2_ADD_1119_U10 , P2_REG3_REG_6_ );
nand NAND2_17341 ( P2_ADD_1119_U11 , P2_ADD_1119_U75 , P2_ADD_1119_U85 );
not NOT1_17342 ( P2_ADD_1119_U12 , P2_REG3_REG_8_ );
not NOT1_17343 ( P2_ADD_1119_U13 , P2_REG3_REG_9_ );
nand NAND2_17344 ( P2_ADD_1119_U14 , P2_ADD_1119_U76 , P2_ADD_1119_U87 );
not NOT1_17345 ( P2_ADD_1119_U15 , P2_REG3_REG_11_ );
not NOT1_17346 ( P2_ADD_1119_U16 , P2_REG3_REG_10_ );
nand NAND2_17347 ( P2_ADD_1119_U17 , P2_ADD_1119_U77 , P2_ADD_1119_U89 );
not NOT1_17348 ( P2_ADD_1119_U18 , P2_REG3_REG_12_ );
nand NAND2_17349 ( P2_ADD_1119_U19 , P2_REG3_REG_12_ , P2_ADD_1119_U91 );
not NOT1_17350 ( P2_ADD_1119_U20 , P2_REG3_REG_13_ );
nand NAND2_17351 ( P2_ADD_1119_U21 , P2_REG3_REG_13_ , P2_ADD_1119_U92 );
not NOT1_17352 ( P2_ADD_1119_U22 , P2_REG3_REG_14_ );
nand NAND2_17353 ( P2_ADD_1119_U23 , P2_REG3_REG_14_ , P2_ADD_1119_U93 );
not NOT1_17354 ( P2_ADD_1119_U24 , P2_REG3_REG_15_ );
nand NAND2_17355 ( P2_ADD_1119_U25 , P2_REG3_REG_15_ , P2_ADD_1119_U94 );
not NOT1_17356 ( P2_ADD_1119_U26 , P2_REG3_REG_16_ );
nand NAND2_17357 ( P2_ADD_1119_U27 , P2_REG3_REG_16_ , P2_ADD_1119_U95 );
not NOT1_17358 ( P2_ADD_1119_U28 , P2_REG3_REG_17_ );
nand NAND2_17359 ( P2_ADD_1119_U29 , P2_REG3_REG_17_ , P2_ADD_1119_U96 );
not NOT1_17360 ( P2_ADD_1119_U30 , P2_REG3_REG_18_ );
nand NAND2_17361 ( P2_ADD_1119_U31 , P2_REG3_REG_18_ , P2_ADD_1119_U97 );
not NOT1_17362 ( P2_ADD_1119_U32 , P2_REG3_REG_19_ );
nand NAND2_17363 ( P2_ADD_1119_U33 , P2_REG3_REG_19_ , P2_ADD_1119_U98 );
not NOT1_17364 ( P2_ADD_1119_U34 , P2_REG3_REG_20_ );
nand NAND2_17365 ( P2_ADD_1119_U35 , P2_REG3_REG_20_ , P2_ADD_1119_U99 );
not NOT1_17366 ( P2_ADD_1119_U36 , P2_REG3_REG_21_ );
nand NAND2_17367 ( P2_ADD_1119_U37 , P2_REG3_REG_21_ , P2_ADD_1119_U100 );
not NOT1_17368 ( P2_ADD_1119_U38 , P2_REG3_REG_22_ );
nand NAND2_17369 ( P2_ADD_1119_U39 , P2_REG3_REG_22_ , P2_ADD_1119_U101 );
not NOT1_17370 ( P2_ADD_1119_U40 , P2_REG3_REG_23_ );
nand NAND2_17371 ( P2_ADD_1119_U41 , P2_REG3_REG_23_ , P2_ADD_1119_U102 );
not NOT1_17372 ( P2_ADD_1119_U42 , P2_REG3_REG_24_ );
nand NAND2_17373 ( P2_ADD_1119_U43 , P2_REG3_REG_24_ , P2_ADD_1119_U103 );
not NOT1_17374 ( P2_ADD_1119_U44 , P2_REG3_REG_25_ );
nand NAND2_17375 ( P2_ADD_1119_U45 , P2_REG3_REG_25_ , P2_ADD_1119_U104 );
not NOT1_17376 ( P2_ADD_1119_U46 , P2_REG3_REG_26_ );
nand NAND2_17377 ( P2_ADD_1119_U47 , P2_REG3_REG_26_ , P2_ADD_1119_U105 );
not NOT1_17378 ( P2_ADD_1119_U48 , P2_REG3_REG_28_ );
not NOT1_17379 ( P2_ADD_1119_U49 , P2_REG3_REG_27_ );
nand NAND2_17380 ( P2_ADD_1119_U50 , P2_ADD_1119_U109 , P2_ADD_1119_U108 );
nand NAND2_17381 ( P2_ADD_1119_U51 , P2_ADD_1119_U111 , P2_ADD_1119_U110 );
nand NAND2_17382 ( P2_ADD_1119_U52 , P2_ADD_1119_U113 , P2_ADD_1119_U112 );
nand NAND2_17383 ( P2_ADD_1119_U53 , P2_ADD_1119_U115 , P2_ADD_1119_U114 );
nand NAND2_17384 ( P2_ADD_1119_U54 , P2_ADD_1119_U117 , P2_ADD_1119_U116 );
nand NAND2_17385 ( P2_ADD_1119_U55 , P2_ADD_1119_U119 , P2_ADD_1119_U118 );
nand NAND2_17386 ( P2_ADD_1119_U56 , P2_ADD_1119_U121 , P2_ADD_1119_U120 );
nand NAND2_17387 ( P2_ADD_1119_U57 , P2_ADD_1119_U123 , P2_ADD_1119_U122 );
nand NAND2_17388 ( P2_ADD_1119_U58 , P2_ADD_1119_U125 , P2_ADD_1119_U124 );
nand NAND2_17389 ( P2_ADD_1119_U59 , P2_ADD_1119_U127 , P2_ADD_1119_U126 );
nand NAND2_17390 ( P2_ADD_1119_U60 , P2_ADD_1119_U129 , P2_ADD_1119_U128 );
nand NAND2_17391 ( P2_ADD_1119_U61 , P2_ADD_1119_U131 , P2_ADD_1119_U130 );
nand NAND2_17392 ( P2_ADD_1119_U62 , P2_ADD_1119_U133 , P2_ADD_1119_U132 );
nand NAND2_17393 ( P2_ADD_1119_U63 , P2_ADD_1119_U135 , P2_ADD_1119_U134 );
nand NAND2_17394 ( P2_ADD_1119_U64 , P2_ADD_1119_U137 , P2_ADD_1119_U136 );
nand NAND2_17395 ( P2_ADD_1119_U65 , P2_ADD_1119_U139 , P2_ADD_1119_U138 );
nand NAND2_17396 ( P2_ADD_1119_U66 , P2_ADD_1119_U141 , P2_ADD_1119_U140 );
nand NAND2_17397 ( P2_ADD_1119_U67 , P2_ADD_1119_U143 , P2_ADD_1119_U142 );
nand NAND2_17398 ( P2_ADD_1119_U68 , P2_ADD_1119_U145 , P2_ADD_1119_U144 );
nand NAND2_17399 ( P2_ADD_1119_U69 , P2_ADD_1119_U147 , P2_ADD_1119_U146 );
nand NAND2_17400 ( P2_ADD_1119_U70 , P2_ADD_1119_U149 , P2_ADD_1119_U148 );
nand NAND2_17401 ( P2_ADD_1119_U71 , P2_ADD_1119_U151 , P2_ADD_1119_U150 );
nand NAND2_17402 ( P2_ADD_1119_U72 , P2_ADD_1119_U153 , P2_ADD_1119_U152 );
nand NAND2_17403 ( P2_ADD_1119_U73 , P2_ADD_1119_U155 , P2_ADD_1119_U154 );
nand NAND2_17404 ( P2_ADD_1119_U74 , P2_ADD_1119_U157 , P2_ADD_1119_U156 );
and AND2_17405 ( P2_ADD_1119_U75 , P2_REG3_REG_7_ , P2_REG3_REG_6_ );
and AND2_17406 ( P2_ADD_1119_U76 , P2_REG3_REG_8_ , P2_REG3_REG_9_ );
and AND2_17407 ( P2_ADD_1119_U77 , P2_REG3_REG_11_ , P2_REG3_REG_10_ );
and AND2_17408 ( P2_ADD_1119_U78 , P2_REG3_REG_28_ , P2_REG3_REG_27_ );
nand NAND2_17409 ( P2_ADD_1119_U79 , P2_REG3_REG_8_ , P2_ADD_1119_U87 );
nand NAND2_17410 ( P2_ADD_1119_U80 , P2_REG3_REG_6_ , P2_ADD_1119_U85 );
nand NAND2_17411 ( P2_ADD_1119_U81 , P2_REG3_REG_4_ , P2_REG3_REG_3_ );
nand NAND2_17412 ( P2_ADD_1119_U82 , P2_REG3_REG_27_ , P2_ADD_1119_U106 );
nand NAND2_17413 ( P2_ADD_1119_U83 , P2_REG3_REG_10_ , P2_ADD_1119_U89 );
not NOT1_17414 ( P2_ADD_1119_U84 , P2_ADD_1119_U81 );
not NOT1_17415 ( P2_ADD_1119_U85 , P2_ADD_1119_U8 );
not NOT1_17416 ( P2_ADD_1119_U86 , P2_ADD_1119_U80 );
not NOT1_17417 ( P2_ADD_1119_U87 , P2_ADD_1119_U11 );
not NOT1_17418 ( P2_ADD_1119_U88 , P2_ADD_1119_U79 );
not NOT1_17419 ( P2_ADD_1119_U89 , P2_ADD_1119_U14 );
not NOT1_17420 ( P2_ADD_1119_U90 , P2_ADD_1119_U83 );
not NOT1_17421 ( P2_ADD_1119_U91 , P2_ADD_1119_U17 );
not NOT1_17422 ( P2_ADD_1119_U92 , P2_ADD_1119_U19 );
not NOT1_17423 ( P2_ADD_1119_U93 , P2_ADD_1119_U21 );
not NOT1_17424 ( P2_ADD_1119_U94 , P2_ADD_1119_U23 );
not NOT1_17425 ( P2_ADD_1119_U95 , P2_ADD_1119_U25 );
not NOT1_17426 ( P2_ADD_1119_U96 , P2_ADD_1119_U27 );
not NOT1_17427 ( P2_ADD_1119_U97 , P2_ADD_1119_U29 );
not NOT1_17428 ( P2_ADD_1119_U98 , P2_ADD_1119_U31 );
not NOT1_17429 ( P2_ADD_1119_U99 , P2_ADD_1119_U33 );
not NOT1_17430 ( P2_ADD_1119_U100 , P2_ADD_1119_U35 );
not NOT1_17431 ( P2_ADD_1119_U101 , P2_ADD_1119_U37 );
not NOT1_17432 ( P2_ADD_1119_U102 , P2_ADD_1119_U39 );
not NOT1_17433 ( P2_ADD_1119_U103 , P2_ADD_1119_U41 );
not NOT1_17434 ( P2_ADD_1119_U104 , P2_ADD_1119_U43 );
not NOT1_17435 ( P2_ADD_1119_U105 , P2_ADD_1119_U45 );
not NOT1_17436 ( P2_ADD_1119_U106 , P2_ADD_1119_U47 );
not NOT1_17437 ( P2_ADD_1119_U107 , P2_ADD_1119_U82 );
nand NAND2_17438 ( P2_ADD_1119_U108 , P2_REG3_REG_9_ , P2_ADD_1119_U79 );
nand NAND2_17439 ( P2_ADD_1119_U109 , P2_ADD_1119_U88 , P2_ADD_1119_U13 );
nand NAND2_17440 ( P2_ADD_1119_U110 , P2_REG3_REG_8_ , P2_ADD_1119_U11 );
nand NAND2_17441 ( P2_ADD_1119_U111 , P2_ADD_1119_U87 , P2_ADD_1119_U12 );
nand NAND2_17442 ( P2_ADD_1119_U112 , P2_REG3_REG_7_ , P2_ADD_1119_U80 );
nand NAND2_17443 ( P2_ADD_1119_U113 , P2_ADD_1119_U86 , P2_ADD_1119_U9 );
nand NAND2_17444 ( P2_ADD_1119_U114 , P2_REG3_REG_6_ , P2_ADD_1119_U8 );
nand NAND2_17445 ( P2_ADD_1119_U115 , P2_ADD_1119_U85 , P2_ADD_1119_U10 );
nand NAND2_17446 ( P2_ADD_1119_U116 , P2_REG3_REG_5_ , P2_ADD_1119_U81 );
nand NAND2_17447 ( P2_ADD_1119_U117 , P2_ADD_1119_U84 , P2_ADD_1119_U6 );
nand NAND2_17448 ( P2_ADD_1119_U118 , P2_REG3_REG_4_ , P2_ADD_1119_U4 );
nand NAND2_17449 ( P2_ADD_1119_U119 , P2_REG3_REG_3_ , P2_ADD_1119_U7 );
nand NAND2_17450 ( P2_ADD_1119_U120 , P2_REG3_REG_28_ , P2_ADD_1119_U82 );
nand NAND2_17451 ( P2_ADD_1119_U121 , P2_ADD_1119_U107 , P2_ADD_1119_U48 );
nand NAND2_17452 ( P2_ADD_1119_U122 , P2_REG3_REG_27_ , P2_ADD_1119_U47 );
nand NAND2_17453 ( P2_ADD_1119_U123 , P2_ADD_1119_U106 , P2_ADD_1119_U49 );
nand NAND2_17454 ( P2_ADD_1119_U124 , P2_REG3_REG_26_ , P2_ADD_1119_U45 );
nand NAND2_17455 ( P2_ADD_1119_U125 , P2_ADD_1119_U105 , P2_ADD_1119_U46 );
nand NAND2_17456 ( P2_ADD_1119_U126 , P2_REG3_REG_25_ , P2_ADD_1119_U43 );
nand NAND2_17457 ( P2_ADD_1119_U127 , P2_ADD_1119_U104 , P2_ADD_1119_U44 );
nand NAND2_17458 ( P2_ADD_1119_U128 , P2_REG3_REG_24_ , P2_ADD_1119_U41 );
nand NAND2_17459 ( P2_ADD_1119_U129 , P2_ADD_1119_U103 , P2_ADD_1119_U42 );
nand NAND2_17460 ( P2_ADD_1119_U130 , P2_REG3_REG_23_ , P2_ADD_1119_U39 );
nand NAND2_17461 ( P2_ADD_1119_U131 , P2_ADD_1119_U102 , P2_ADD_1119_U40 );
nand NAND2_17462 ( P2_ADD_1119_U132 , P2_REG3_REG_22_ , P2_ADD_1119_U37 );
nand NAND2_17463 ( P2_ADD_1119_U133 , P2_ADD_1119_U101 , P2_ADD_1119_U38 );
nand NAND2_17464 ( P2_ADD_1119_U134 , P2_REG3_REG_21_ , P2_ADD_1119_U35 );
nand NAND2_17465 ( P2_ADD_1119_U135 , P2_ADD_1119_U100 , P2_ADD_1119_U36 );
nand NAND2_17466 ( P2_ADD_1119_U136 , P2_REG3_REG_20_ , P2_ADD_1119_U33 );
nand NAND2_17467 ( P2_ADD_1119_U137 , P2_ADD_1119_U99 , P2_ADD_1119_U34 );
nand NAND2_17468 ( P2_ADD_1119_U138 , P2_REG3_REG_19_ , P2_ADD_1119_U31 );
nand NAND2_17469 ( P2_ADD_1119_U139 , P2_ADD_1119_U98 , P2_ADD_1119_U32 );
nand NAND2_17470 ( P2_ADD_1119_U140 , P2_REG3_REG_18_ , P2_ADD_1119_U29 );
nand NAND2_17471 ( P2_ADD_1119_U141 , P2_ADD_1119_U97 , P2_ADD_1119_U30 );
nand NAND2_17472 ( P2_ADD_1119_U142 , P2_REG3_REG_17_ , P2_ADD_1119_U27 );
nand NAND2_17473 ( P2_ADD_1119_U143 , P2_ADD_1119_U96 , P2_ADD_1119_U28 );
nand NAND2_17474 ( P2_ADD_1119_U144 , P2_REG3_REG_16_ , P2_ADD_1119_U25 );
nand NAND2_17475 ( P2_ADD_1119_U145 , P2_ADD_1119_U95 , P2_ADD_1119_U26 );
nand NAND2_17476 ( P2_ADD_1119_U146 , P2_REG3_REG_15_ , P2_ADD_1119_U23 );
nand NAND2_17477 ( P2_ADD_1119_U147 , P2_ADD_1119_U94 , P2_ADD_1119_U24 );
nand NAND2_17478 ( P2_ADD_1119_U148 , P2_REG3_REG_14_ , P2_ADD_1119_U21 );
nand NAND2_17479 ( P2_ADD_1119_U149 , P2_ADD_1119_U93 , P2_ADD_1119_U22 );
nand NAND2_17480 ( P2_ADD_1119_U150 , P2_REG3_REG_13_ , P2_ADD_1119_U19 );
nand NAND2_17481 ( P2_ADD_1119_U151 , P2_ADD_1119_U92 , P2_ADD_1119_U20 );
nand NAND2_17482 ( P2_ADD_1119_U152 , P2_REG3_REG_12_ , P2_ADD_1119_U17 );
nand NAND2_17483 ( P2_ADD_1119_U153 , P2_ADD_1119_U91 , P2_ADD_1119_U18 );
nand NAND2_17484 ( P2_ADD_1119_U154 , P2_REG3_REG_11_ , P2_ADD_1119_U83 );
nand NAND2_17485 ( P2_ADD_1119_U155 , P2_ADD_1119_U90 , P2_ADD_1119_U15 );
nand NAND2_17486 ( P2_ADD_1119_U156 , P2_REG3_REG_10_ , P2_ADD_1119_U14 );
nand NAND2_17487 ( P2_ADD_1119_U157 , P2_ADD_1119_U89 , P2_ADD_1119_U16 );
and AND2_17488 ( P2_SUB_1108_U6 , P2_SUB_1108_U172 , P2_SUB_1108_U40 );
and AND2_17489 ( P2_SUB_1108_U7 , P2_SUB_1108_U170 , P2_SUB_1108_U140 );
and AND2_17490 ( P2_SUB_1108_U8 , P2_SUB_1108_U169 , P2_SUB_1108_U37 );
and AND2_17491 ( P2_SUB_1108_U9 , P2_SUB_1108_U168 , P2_SUB_1108_U38 );
and AND2_17492 ( P2_SUB_1108_U10 , P2_SUB_1108_U166 , P2_SUB_1108_U143 );
and AND2_17493 ( P2_SUB_1108_U11 , P2_SUB_1108_U165 , P2_SUB_1108_U30 );
and AND2_17494 ( P2_SUB_1108_U12 , P2_SUB_1108_U164 , P2_SUB_1108_U36 );
and AND2_17495 ( P2_SUB_1108_U13 , P2_SUB_1108_U162 , P2_SUB_1108_U32 );
and AND2_17496 ( P2_SUB_1108_U14 , P2_SUB_1108_U160 , P2_SUB_1108_U33 );
and AND2_17497 ( P2_SUB_1108_U15 , P2_SUB_1108_U159 , P2_SUB_1108_U109 );
and AND2_17498 ( P2_SUB_1108_U16 , P2_SUB_1108_U157 , P2_SUB_1108_U29 );
and AND2_17499 ( P2_SUB_1108_U17 , P2_SUB_1108_U155 , P2_SUB_1108_U23 );
and AND2_17500 ( P2_SUB_1108_U18 , P2_SUB_1108_U138 , P2_SUB_1108_U128 );
and AND2_17501 ( P2_SUB_1108_U19 , P2_SUB_1108_U137 , P2_SUB_1108_U25 );
and AND2_17502 ( P2_SUB_1108_U20 , P2_SUB_1108_U136 , P2_SUB_1108_U26 );
and AND2_17503 ( P2_SUB_1108_U21 , P2_SUB_1108_U134 , P2_SUB_1108_U131 );
and AND2_17504 ( P2_SUB_1108_U22 , P2_SUB_1108_U133 , P2_SUB_1108_U24 );
or OR3_17505 ( P2_SUB_1108_U23 , P2_IR_REG_1_ , P2_IR_REG_0_ , P2_IR_REG_2_ );
nand NAND3_17506 ( P2_SUB_1108_U24 , P2_SUB_1108_U45 , P2_SUB_1108_U174 , P2_SUB_1108_U44 );
nand NAND2_17507 ( P2_SUB_1108_U25 , P2_SUB_1108_U46 , P2_SUB_1108_U174 );
nand NAND2_17508 ( P2_SUB_1108_U26 , P2_SUB_1108_U47 , P2_SUB_1108_U129 );
not NOT1_17509 ( P2_SUB_1108_U27 , P2_IR_REG_7_ );
not NOT1_17510 ( P2_SUB_1108_U28 , P2_IR_REG_3_ );
nand NAND2_17511 ( P2_SUB_1108_U29 , P2_SUB_1108_U57 , P2_SUB_1108_U52 );
nand NAND4_17512 ( P2_SUB_1108_U30 , P2_SUB_1108_U91 , P2_SUB_1108_U90 , P2_SUB_1108_U89 , P2_SUB_1108_U88 );
nand NAND2_17513 ( P2_SUB_1108_U31 , P2_SUB_1108_U92 , P2_SUB_1108_U144 );
nand NAND2_17514 ( P2_SUB_1108_U32 , P2_SUB_1108_U93 , P2_SUB_1108_U147 );
nand NAND2_17515 ( P2_SUB_1108_U33 , P2_SUB_1108_U149 , P2_SUB_1108_U34 );
not NOT1_17516 ( P2_SUB_1108_U34 , P2_IR_REG_24_ );
nand NAND2_17517 ( P2_SUB_1108_U35 , P2_SUB_1108_U147 , P2_SUB_1108_U115 );
nand NAND2_17518 ( P2_SUB_1108_U36 , P2_SUB_1108_U94 , P2_SUB_1108_U144 );
nand NAND2_17519 ( P2_SUB_1108_U37 , P2_SUB_1108_U95 , P2_SUB_1108_U132 );
nand NAND2_17520 ( P2_SUB_1108_U38 , P2_SUB_1108_U96 , P2_SUB_1108_U141 );
not NOT1_17521 ( P2_SUB_1108_U39 , P2_IR_REG_15_ );
nand NAND2_17522 ( P2_SUB_1108_U40 , P2_SUB_1108_U97 , P2_SUB_1108_U132 );
not NOT1_17523 ( P2_SUB_1108_U41 , P2_IR_REG_11_ );
nand NAND2_17524 ( P2_SUB_1108_U42 , P2_SUB_1108_U196 , P2_SUB_1108_U195 );
nand NAND2_17525 ( P2_SUB_1108_U43 , P2_SUB_1108_U180 , P2_SUB_1108_U179 );
nor nor_17526 ( P2_SUB_1108_U44 , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ , P2_IR_REG_6_ );
nor nor_17527 ( P2_SUB_1108_U45 , P2_IR_REG_7_ , P2_IR_REG_8_ );
nor nor_17528 ( P2_SUB_1108_U46 , P2_IR_REG_3_ , P2_IR_REG_4_ );
nor nor_17529 ( P2_SUB_1108_U47 , P2_IR_REG_5_ , P2_IR_REG_6_ );
nor nor_17530 ( P2_SUB_1108_U48 , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_ , P2_IR_REG_13_ );
nor nor_17531 ( P2_SUB_1108_U49 , P2_IR_REG_14_ , P2_IR_REG_15_ , P2_IR_REG_16_ , P2_IR_REG_17_ );
nor nor_17532 ( P2_SUB_1108_U50 , P2_IR_REG_18_ , P2_IR_REG_19_ , P2_IR_REG_1_ , P2_IR_REG_0_ );
nor nor_17533 ( P2_SUB_1108_U51 , P2_IR_REG_22_ , P2_IR_REG_20_ , P2_IR_REG_21_ );
and AND4_17534 ( P2_SUB_1108_U52 , P2_SUB_1108_U51 , P2_SUB_1108_U50 , P2_SUB_1108_U49 , P2_SUB_1108_U48 );
nor nor_17535 ( P2_SUB_1108_U53 , P2_IR_REG_23_ , P2_IR_REG_24_ , P2_IR_REG_25_ , P2_IR_REG_26_ );
nor nor_17536 ( P2_SUB_1108_U54 , P2_IR_REG_27_ , P2_IR_REG_28_ , P2_IR_REG_29_ , P2_IR_REG_2_ );
nor nor_17537 ( P2_SUB_1108_U55 , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ , P2_IR_REG_6_ );
nor nor_17538 ( P2_SUB_1108_U56 , P2_IR_REG_9_ , P2_IR_REG_7_ , P2_IR_REG_8_ );
and AND4_17539 ( P2_SUB_1108_U57 , P2_SUB_1108_U56 , P2_SUB_1108_U55 , P2_SUB_1108_U54 , P2_SUB_1108_U53 );
nor nor_17540 ( P2_SUB_1108_U58 , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_ , P2_IR_REG_13_ );
nor nor_17541 ( P2_SUB_1108_U59 , P2_IR_REG_14_ , P2_IR_REG_15_ , P2_IR_REG_16_ , P2_IR_REG_17_ );
nor nor_17542 ( P2_SUB_1108_U60 , P2_IR_REG_18_ , P2_IR_REG_19_ , P2_IR_REG_1_ , P2_IR_REG_0_ );
nor nor_17543 ( P2_SUB_1108_U61 , P2_IR_REG_22_ , P2_IR_REG_20_ , P2_IR_REG_21_ );
and AND4_17544 ( P2_SUB_1108_U62 , P2_SUB_1108_U61 , P2_SUB_1108_U60 , P2_SUB_1108_U59 , P2_SUB_1108_U58 );
nor nor_17545 ( P2_SUB_1108_U63 , P2_IR_REG_23_ , P2_IR_REG_24_ , P2_IR_REG_25_ , P2_IR_REG_26_ );
nor nor_17546 ( P2_SUB_1108_U64 , P2_IR_REG_2_ , P2_IR_REG_27_ , P2_IR_REG_28_ );
nor nor_17547 ( P2_SUB_1108_U65 , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ , P2_IR_REG_6_ );
nor nor_17548 ( P2_SUB_1108_U66 , P2_IR_REG_9_ , P2_IR_REG_7_ , P2_IR_REG_8_ );
and AND4_17549 ( P2_SUB_1108_U67 , P2_SUB_1108_U66 , P2_SUB_1108_U65 , P2_SUB_1108_U64 , P2_SUB_1108_U63 );
nor nor_17550 ( P2_SUB_1108_U68 , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_ , P2_IR_REG_13_ );
nor nor_17551 ( P2_SUB_1108_U69 , P2_IR_REG_16_ , P2_IR_REG_14_ , P2_IR_REG_15_ );
nor nor_17552 ( P2_SUB_1108_U70 , P2_IR_REG_17_ , P2_IR_REG_18_ , P2_IR_REG_19_ , P2_IR_REG_1_ );
nor nor_17553 ( P2_SUB_1108_U71 , P2_IR_REG_21_ , P2_IR_REG_0_ , P2_IR_REG_20_ );
and AND4_17554 ( P2_SUB_1108_U72 , P2_SUB_1108_U71 , P2_SUB_1108_U70 , P2_SUB_1108_U69 , P2_SUB_1108_U68 );
nor nor_17555 ( P2_SUB_1108_U73 , P2_IR_REG_22_ , P2_IR_REG_23_ , P2_IR_REG_24_ , P2_IR_REG_25_ );
nor nor_17556 ( P2_SUB_1108_U74 , P2_IR_REG_2_ , P2_IR_REG_26_ , P2_IR_REG_27_ );
nor nor_17557 ( P2_SUB_1108_U75 , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ , P2_IR_REG_6_ );
nor nor_17558 ( P2_SUB_1108_U76 , P2_IR_REG_9_ , P2_IR_REG_7_ , P2_IR_REG_8_ );
and AND4_17559 ( P2_SUB_1108_U77 , P2_SUB_1108_U76 , P2_SUB_1108_U75 , P2_SUB_1108_U74 , P2_SUB_1108_U73 );
nor nor_17560 ( P2_SUB_1108_U78 , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_ , P2_IR_REG_13_ );
nor nor_17561 ( P2_SUB_1108_U79 , P2_IR_REG_16_ , P2_IR_REG_14_ , P2_IR_REG_15_ );
nor nor_17562 ( P2_SUB_1108_U80 , P2_IR_REG_17_ , P2_IR_REG_18_ , P2_IR_REG_19_ , P2_IR_REG_1_ );
nor nor_17563 ( P2_SUB_1108_U81 , P2_IR_REG_21_ , P2_IR_REG_0_ , P2_IR_REG_20_ );
and AND4_17564 ( P2_SUB_1108_U82 , P2_SUB_1108_U81 , P2_SUB_1108_U80 , P2_SUB_1108_U79 , P2_SUB_1108_U78 );
nor nor_17565 ( P2_SUB_1108_U83 , P2_IR_REG_22_ , P2_IR_REG_23_ , P2_IR_REG_24_ , P2_IR_REG_25_ );
nor nor_17566 ( P2_SUB_1108_U84 , P2_IR_REG_3_ , P2_IR_REG_26_ , P2_IR_REG_2_ );
nor nor_17567 ( P2_SUB_1108_U85 , P2_IR_REG_6_ , P2_IR_REG_4_ , P2_IR_REG_5_ );
nor nor_17568 ( P2_SUB_1108_U86 , P2_IR_REG_9_ , P2_IR_REG_7_ , P2_IR_REG_8_ );
and AND4_17569 ( P2_SUB_1108_U87 , P2_SUB_1108_U86 , P2_SUB_1108_U85 , P2_SUB_1108_U84 , P2_SUB_1108_U83 );
nor nor_17570 ( P2_SUB_1108_U88 , P2_IR_REG_13_ , P2_IR_REG_14_ , P2_IR_REG_12_ , P2_IR_REG_10_ , P2_IR_REG_11_ );
nor nor_17571 ( P2_SUB_1108_U89 , P2_IR_REG_15_ , P2_IR_REG_16_ , P2_IR_REG_1_ , P2_IR_REG_0_ );
nor nor_17572 ( P2_SUB_1108_U90 , P2_IR_REG_2_ , P2_IR_REG_3_ , P2_IR_REG_4_ , P2_IR_REG_5_ );
nor nor_17573 ( P2_SUB_1108_U91 , P2_IR_REG_6_ , P2_IR_REG_7_ , P2_IR_REG_8_ , P2_IR_REG_9_ );
nor nor_17574 ( P2_SUB_1108_U92 , P2_IR_REG_17_ , P2_IR_REG_18_ , P2_IR_REG_19_ , P2_IR_REG_20_ );
nor nor_17575 ( P2_SUB_1108_U93 , P2_IR_REG_23_ , P2_IR_REG_21_ , P2_IR_REG_22_ );
nor nor_17576 ( P2_SUB_1108_U94 , P2_IR_REG_17_ , P2_IR_REG_18_ );
nor nor_17577 ( P2_SUB_1108_U95 , P2_IR_REG_10_ , P2_IR_REG_11_ , P2_IR_REG_12_ , P2_IR_REG_9_ );
nor nor_17578 ( P2_SUB_1108_U96 , P2_IR_REG_13_ , P2_IR_REG_14_ );
nor nor_17579 ( P2_SUB_1108_U97 , P2_IR_REG_10_ , P2_IR_REG_9_ );
not NOT1_17580 ( P2_SUB_1108_U98 , P2_IR_REG_9_ );
and AND2_17581 ( P2_SUB_1108_U99 , P2_SUB_1108_U176 , P2_SUB_1108_U175 );
not NOT1_17582 ( P2_SUB_1108_U100 , P2_IR_REG_5_ );
and AND2_17583 ( P2_SUB_1108_U101 , P2_SUB_1108_U178 , P2_SUB_1108_U177 );
not NOT1_17584 ( P2_SUB_1108_U102 , P2_IR_REG_31_ );
not NOT1_17585 ( P2_SUB_1108_U103 , P2_IR_REG_30_ );
and AND2_17586 ( P2_SUB_1108_U104 , P2_SUB_1108_U182 , P2_SUB_1108_U181 );
not NOT1_17587 ( P2_SUB_1108_U105 , P2_IR_REG_28_ );
nand NAND2_17588 ( P2_SUB_1108_U106 , P2_SUB_1108_U77 , P2_SUB_1108_U72 );
and AND2_17589 ( P2_SUB_1108_U107 , P2_SUB_1108_U184 , P2_SUB_1108_U183 );
not NOT1_17590 ( P2_SUB_1108_U108 , P2_IR_REG_27_ );
nand NAND2_17591 ( P2_SUB_1108_U109 , P2_SUB_1108_U87 , P2_SUB_1108_U82 );
and AND2_17592 ( P2_SUB_1108_U110 , P2_SUB_1108_U186 , P2_SUB_1108_U185 );
not NOT1_17593 ( P2_SUB_1108_U111 , P2_IR_REG_25_ );
and AND2_17594 ( P2_SUB_1108_U112 , P2_SUB_1108_U188 , P2_SUB_1108_U187 );
not NOT1_17595 ( P2_SUB_1108_U113 , P2_IR_REG_22_ );
and AND2_17596 ( P2_SUB_1108_U114 , P2_SUB_1108_U190 , P2_SUB_1108_U189 );
not NOT1_17597 ( P2_SUB_1108_U115 , P2_IR_REG_21_ );
and AND2_17598 ( P2_SUB_1108_U116 , P2_SUB_1108_U192 , P2_SUB_1108_U191 );
not NOT1_17599 ( P2_SUB_1108_U117 , P2_IR_REG_20_ );
nand NAND2_17600 ( P2_SUB_1108_U118 , P2_SUB_1108_U145 , P2_SUB_1108_U122 );
and AND2_17601 ( P2_SUB_1108_U119 , P2_SUB_1108_U194 , P2_SUB_1108_U193 );
not NOT1_17602 ( P2_SUB_1108_U120 , P2_IR_REG_1_ );
not NOT1_17603 ( P2_SUB_1108_U121 , P2_IR_REG_0_ );
not NOT1_17604 ( P2_SUB_1108_U122 , P2_IR_REG_19_ );
and AND2_17605 ( P2_SUB_1108_U123 , P2_SUB_1108_U198 , P2_SUB_1108_U197 );
not NOT1_17606 ( P2_SUB_1108_U124 , P2_IR_REG_17_ );
and AND2_17607 ( P2_SUB_1108_U125 , P2_SUB_1108_U200 , P2_SUB_1108_U199 );
not NOT1_17608 ( P2_SUB_1108_U126 , P2_IR_REG_13_ );
and AND2_17609 ( P2_SUB_1108_U127 , P2_SUB_1108_U202 , P2_SUB_1108_U201 );
nand NAND2_17610 ( P2_SUB_1108_U128 , P2_SUB_1108_U174 , P2_SUB_1108_U28 );
not NOT1_17611 ( P2_SUB_1108_U129 , P2_SUB_1108_U25 );
not NOT1_17612 ( P2_SUB_1108_U130 , P2_SUB_1108_U26 );
nand NAND2_17613 ( P2_SUB_1108_U131 , P2_SUB_1108_U130 , P2_SUB_1108_U27 );
not NOT1_17614 ( P2_SUB_1108_U132 , P2_SUB_1108_U24 );
nand NAND2_17615 ( P2_SUB_1108_U133 , P2_IR_REG_8_ , P2_SUB_1108_U131 );
nand NAND2_17616 ( P2_SUB_1108_U134 , P2_IR_REG_7_ , P2_SUB_1108_U26 );
nand NAND2_17617 ( P2_SUB_1108_U135 , P2_SUB_1108_U129 , P2_SUB_1108_U100 );
nand NAND2_17618 ( P2_SUB_1108_U136 , P2_IR_REG_6_ , P2_SUB_1108_U135 );
nand NAND2_17619 ( P2_SUB_1108_U137 , P2_IR_REG_4_ , P2_SUB_1108_U128 );
nand NAND2_17620 ( P2_SUB_1108_U138 , P2_IR_REG_3_ , P2_SUB_1108_U23 );
not NOT1_17621 ( P2_SUB_1108_U139 , P2_SUB_1108_U40 );
nand NAND2_17622 ( P2_SUB_1108_U140 , P2_SUB_1108_U139 , P2_SUB_1108_U41 );
not NOT1_17623 ( P2_SUB_1108_U141 , P2_SUB_1108_U37 );
not NOT1_17624 ( P2_SUB_1108_U142 , P2_SUB_1108_U38 );
nand NAND2_17625 ( P2_SUB_1108_U143 , P2_SUB_1108_U142 , P2_SUB_1108_U39 );
not NOT1_17626 ( P2_SUB_1108_U144 , P2_SUB_1108_U30 );
not NOT1_17627 ( P2_SUB_1108_U145 , P2_SUB_1108_U36 );
not NOT1_17628 ( P2_SUB_1108_U146 , P2_SUB_1108_U118 );
not NOT1_17629 ( P2_SUB_1108_U147 , P2_SUB_1108_U31 );
not NOT1_17630 ( P2_SUB_1108_U148 , P2_SUB_1108_U35 );
not NOT1_17631 ( P2_SUB_1108_U149 , P2_SUB_1108_U32 );
not NOT1_17632 ( P2_SUB_1108_U150 , P2_SUB_1108_U33 );
not NOT1_17633 ( P2_SUB_1108_U151 , P2_SUB_1108_U109 );
not NOT1_17634 ( P2_SUB_1108_U152 , P2_SUB_1108_U106 );
not NOT1_17635 ( P2_SUB_1108_U153 , P2_SUB_1108_U29 );
or OR2_17636 ( P2_SUB_1108_U154 , P2_IR_REG_1_ , P2_IR_REG_0_ );
nand NAND2_17637 ( P2_SUB_1108_U155 , P2_IR_REG_2_ , P2_SUB_1108_U154 );
nand NAND2_17638 ( P2_SUB_1108_U156 , P2_SUB_1108_U67 , P2_SUB_1108_U62 );
nand NAND2_17639 ( P2_SUB_1108_U157 , P2_IR_REG_29_ , P2_SUB_1108_U156 );
nand NAND2_17640 ( P2_SUB_1108_U158 , P2_SUB_1108_U150 , P2_SUB_1108_U111 );
nand NAND2_17641 ( P2_SUB_1108_U159 , P2_IR_REG_26_ , P2_SUB_1108_U158 );
nand NAND2_17642 ( P2_SUB_1108_U160 , P2_IR_REG_24_ , P2_SUB_1108_U32 );
nand NAND2_17643 ( P2_SUB_1108_U161 , P2_SUB_1108_U148 , P2_SUB_1108_U113 );
nand NAND2_17644 ( P2_SUB_1108_U162 , P2_IR_REG_23_ , P2_SUB_1108_U161 );
nand NAND2_17645 ( P2_SUB_1108_U163 , P2_SUB_1108_U144 , P2_SUB_1108_U124 );
nand NAND2_17646 ( P2_SUB_1108_U164 , P2_IR_REG_18_ , P2_SUB_1108_U163 );
nand NAND2_17647 ( P2_SUB_1108_U165 , P2_IR_REG_16_ , P2_SUB_1108_U143 );
nand NAND2_17648 ( P2_SUB_1108_U166 , P2_IR_REG_15_ , P2_SUB_1108_U38 );
nand NAND2_17649 ( P2_SUB_1108_U167 , P2_SUB_1108_U141 , P2_SUB_1108_U126 );
nand NAND2_17650 ( P2_SUB_1108_U168 , P2_IR_REG_14_ , P2_SUB_1108_U167 );
nand NAND2_17651 ( P2_SUB_1108_U169 , P2_IR_REG_12_ , P2_SUB_1108_U140 );
nand NAND2_17652 ( P2_SUB_1108_U170 , P2_IR_REG_11_ , P2_SUB_1108_U40 );
nand NAND2_17653 ( P2_SUB_1108_U171 , P2_SUB_1108_U132 , P2_SUB_1108_U98 );
nand NAND2_17654 ( P2_SUB_1108_U172 , P2_IR_REG_10_ , P2_SUB_1108_U171 );
nand NAND2_17655 ( P2_SUB_1108_U173 , P2_SUB_1108_U153 , P2_SUB_1108_U103 );
not NOT1_17656 ( P2_SUB_1108_U174 , P2_SUB_1108_U23 );
nand NAND2_17657 ( P2_SUB_1108_U175 , P2_IR_REG_9_ , P2_SUB_1108_U24 );
nand NAND2_17658 ( P2_SUB_1108_U176 , P2_SUB_1108_U132 , P2_SUB_1108_U98 );
nand NAND2_17659 ( P2_SUB_1108_U177 , P2_IR_REG_5_ , P2_SUB_1108_U25 );
nand NAND2_17660 ( P2_SUB_1108_U178 , P2_SUB_1108_U129 , P2_SUB_1108_U100 );
nand NAND2_17661 ( P2_SUB_1108_U179 , P2_SUB_1108_U173 , P2_SUB_1108_U102 );
nand NAND3_17662 ( P2_SUB_1108_U180 , P2_SUB_1108_U153 , P2_SUB_1108_U103 , P2_IR_REG_31_ );
nand NAND2_17663 ( P2_SUB_1108_U181 , P2_IR_REG_30_ , P2_SUB_1108_U29 );
nand NAND2_17664 ( P2_SUB_1108_U182 , P2_SUB_1108_U153 , P2_SUB_1108_U103 );
nand NAND2_17665 ( P2_SUB_1108_U183 , P2_IR_REG_28_ , P2_SUB_1108_U106 );
nand NAND2_17666 ( P2_SUB_1108_U184 , P2_SUB_1108_U152 , P2_SUB_1108_U105 );
nand NAND2_17667 ( P2_SUB_1108_U185 , P2_IR_REG_27_ , P2_SUB_1108_U109 );
nand NAND2_17668 ( P2_SUB_1108_U186 , P2_SUB_1108_U151 , P2_SUB_1108_U108 );
nand NAND2_17669 ( P2_SUB_1108_U187 , P2_IR_REG_25_ , P2_SUB_1108_U33 );
nand NAND2_17670 ( P2_SUB_1108_U188 , P2_SUB_1108_U150 , P2_SUB_1108_U111 );
nand NAND2_17671 ( P2_SUB_1108_U189 , P2_IR_REG_22_ , P2_SUB_1108_U35 );
nand NAND2_17672 ( P2_SUB_1108_U190 , P2_SUB_1108_U148 , P2_SUB_1108_U113 );
nand NAND2_17673 ( P2_SUB_1108_U191 , P2_IR_REG_21_ , P2_SUB_1108_U31 );
nand NAND2_17674 ( P2_SUB_1108_U192 , P2_SUB_1108_U147 , P2_SUB_1108_U115 );
nand NAND2_17675 ( P2_SUB_1108_U193 , P2_IR_REG_20_ , P2_SUB_1108_U118 );
nand NAND2_17676 ( P2_SUB_1108_U194 , P2_SUB_1108_U146 , P2_SUB_1108_U117 );
nand NAND2_17677 ( P2_SUB_1108_U195 , P2_IR_REG_1_ , P2_SUB_1108_U121 );
nand NAND2_17678 ( P2_SUB_1108_U196 , P2_IR_REG_0_ , P2_SUB_1108_U120 );
nand NAND2_17679 ( P2_SUB_1108_U197 , P2_IR_REG_19_ , P2_SUB_1108_U36 );
nand NAND2_17680 ( P2_SUB_1108_U198 , P2_SUB_1108_U145 , P2_SUB_1108_U122 );
nand NAND2_17681 ( P2_SUB_1108_U199 , P2_IR_REG_17_ , P2_SUB_1108_U30 );
nand NAND2_17682 ( P2_SUB_1108_U200 , P2_SUB_1108_U144 , P2_SUB_1108_U124 );
nand NAND2_17683 ( P2_SUB_1108_U201 , P2_IR_REG_13_ , P2_SUB_1108_U37 );
nand NAND2_17684 ( P2_SUB_1108_U202 , P2_SUB_1108_U141 , P2_SUB_1108_U126 );
and AND2_17685 ( P2_R1299_U6 , P2_U3061 , P2_R1299_U7 );
not NOT1_17686 ( P2_R1299_U7 , P2_U3058 );
and AND3_17687 ( P2_R1312_U6 , P2_R1312_U172 , P2_R1312_U170 , P2_R1312_U171 );
and AND2_17688 ( P2_R1312_U7 , P2_R1312_U85 , P2_R1312_U84 );
and AND2_17689 ( P2_R1312_U8 , P2_R1312_U7 , P2_R1312_U173 );
and AND2_17690 ( P2_R1312_U9 , P2_R1312_U183 , P2_R1312_U182 );
and AND2_17691 ( P2_R1312_U10 , P2_R1312_U213 , P2_R1312_U212 );
and AND3_17692 ( P2_R1312_U11 , P2_R1312_U14 , P2_R1312_U82 , P2_R1312_U169 );
and AND4_17693 ( P2_R1312_U12 , P2_R1312_U157 , P2_R1312_U156 , P2_R1312_U155 , P2_R1312_U154 );
and AND4_17694 ( P2_R1312_U13 , P2_R1312_U176 , P2_R1312_U175 , P2_R1312_U174 , P2_R1312_U173 );
and AND3_17695 ( P2_R1312_U14 , P2_R1312_U162 , P2_R1312_U161 , P2_R1312_U164 );
and AND5_17696 ( P2_R1312_U15 , P2_R1312_U6 , P2_R1312_U11 , P2_R1312_U83 , P2_R1312_U165 , P2_R1312_U17 );
and AND2_17697 ( P2_R1312_U16 , P2_R1312_U165 , P2_R1312_U163 );
and AND2_17698 ( P2_R1312_U17 , P2_R1312_U225 , P2_R1312_U224 );
nand NAND5_17699 ( P2_R1312_U18 , P2_R1312_U152 , P2_R1312_U151 , P2_R1312_U150 , P2_R1312_U147 , P2_R1312_U144 );
not NOT1_17700 ( P2_R1312_U19 , P2_U3090 );
not NOT1_17701 ( P2_R1312_U20 , P2_U3093 );
not NOT1_17702 ( P2_R1312_U21 , P2_U3091 );
not NOT1_17703 ( P2_R1312_U22 , P2_U3092 );
not NOT1_17704 ( P2_R1312_U23 , P2_U3126 );
not NOT1_17705 ( P2_R1312_U24 , P2_U3123 );
not NOT1_17706 ( P2_R1312_U25 , P2_U3089 );
not NOT1_17707 ( P2_R1312_U26 , P2_U3121 );
not NOT1_17708 ( P2_R1312_U27 , P2_U3105 );
not NOT1_17709 ( P2_R1312_U28 , P2_U3106 );
not NOT1_17710 ( P2_R1312_U29 , P2_U3108 );
not NOT1_17711 ( P2_R1312_U30 , P2_U3107 );
not NOT1_17712 ( P2_R1312_U31 , P2_U3109 );
not NOT1_17713 ( P2_R1312_U32 , P2_U3110 );
not NOT1_17714 ( P2_R1312_U33 , P2_U3111 );
not NOT1_17715 ( P2_R1312_U34 , P2_U3112 );
not NOT1_17716 ( P2_R1312_U35 , P2_U3115 );
not NOT1_17717 ( P2_R1312_U36 , P2_U3116 );
not NOT1_17718 ( P2_R1312_U37 , P2_U3114 );
not NOT1_17719 ( P2_R1312_U38 , P2_U3113 );
not NOT1_17720 ( P2_R1312_U39 , P2_U3104 );
not NOT1_17721 ( P2_R1312_U40 , P2_U3094 );
not NOT1_17722 ( P2_R1312_U41 , P2_U3102 );
not NOT1_17723 ( P2_R1312_U42 , P2_U3101 );
not NOT1_17724 ( P2_R1312_U43 , P2_U3103 );
not NOT1_17725 ( P2_R1312_U44 , P2_U3100 );
not NOT1_17726 ( P2_R1312_U45 , P2_U3099 );
not NOT1_17727 ( P2_R1312_U46 , P2_U3095 );
not NOT1_17728 ( P2_R1312_U47 , P2_U3097 );
not NOT1_17729 ( P2_R1312_U48 , P2_U3098 );
not NOT1_17730 ( P2_R1312_U49 , P2_U3096 );
not NOT1_17731 ( P2_R1312_U50 , P2_U3149 );
not NOT1_17732 ( P2_R1312_U51 , P2_U3117 );
not NOT1_17733 ( P2_R1312_U52 , P2_U3118 );
not NOT1_17734 ( P2_R1312_U53 , P2_U3119 );
not NOT1_17735 ( P2_R1312_U54 , P2_U3151 );
not NOT1_17736 ( P2_R1312_U55 , P2_U3127 );
not NOT1_17737 ( P2_R1312_U56 , P2_U3125 );
not NOT1_17738 ( P2_R1312_U57 , P2_U3124 );
not NOT1_17739 ( P2_R1312_U58 , P2_U3140 );
not NOT1_17740 ( P2_R1312_U59 , P2_U3141 );
not NOT1_17741 ( P2_R1312_U60 , P2_U3143 );
not NOT1_17742 ( P2_R1312_U61 , P2_U3128 );
not NOT1_17743 ( P2_R1312_U62 , P2_U3129 );
not NOT1_17744 ( P2_R1312_U63 , P2_U3131 );
not NOT1_17745 ( P2_R1312_U64 , P2_U3134 );
not NOT1_17746 ( P2_R1312_U65 , P2_U3135 );
not NOT1_17747 ( P2_R1312_U66 , P2_U3137 );
not NOT1_17748 ( P2_R1312_U67 , P2_U3146 );
not NOT1_17749 ( P2_R1312_U68 , P2_U3147 );
not NOT1_17750 ( P2_R1312_U69 , P2_U3133 );
not NOT1_17751 ( P2_R1312_U70 , P2_U3139 );
not NOT1_17752 ( P2_R1312_U71 , P2_U3145 );
not NOT1_17753 ( P2_R1312_U72 , P2_U3130 );
not NOT1_17754 ( P2_R1312_U73 , P2_U3132 );
not NOT1_17755 ( P2_R1312_U74 , P2_U3136 );
not NOT1_17756 ( P2_R1312_U75 , P2_U3138 );
not NOT1_17757 ( P2_R1312_U76 , P2_U3142 );
not NOT1_17758 ( P2_R1312_U77 , P2_U3144 );
not NOT1_17759 ( P2_R1312_U78 , P2_U3148 );
not NOT1_17760 ( P2_R1312_U79 , P2_U3150 );
not NOT1_17761 ( P2_R1312_U80 , P2_U3122 );
and AND2_17762 ( P2_R1312_U81 , P2_R1312_U17 , P2_R1312_U166 );
and AND2_17763 ( P2_R1312_U82 , P2_R1312_U160 , P2_R1312_U159 );
and AND2_17764 ( P2_R1312_U83 , P2_R1312_U163 , P2_R1312_U158 );
and AND4_17765 ( P2_R1312_U84 , P2_R1312_U177 , P2_R1312_U176 , P2_R1312_U175 , P2_R1312_U174 );
and AND3_17766 ( P2_R1312_U85 , P2_R1312_U179 , P2_R1312_U178 , P2_R1312_U180 );
and AND4_17767 ( P2_R1312_U86 , P2_R1312_U168 , P2_R1312_U51 , P2_R1312_U167 , P2_R1312_U166 );
and AND2_17768 ( P2_R1312_U87 , P2_U3149 , P2_R1312_U12 );
and AND2_17769 ( P2_R1312_U88 , P2_R1312_U186 , P2_R1312_U173 );
and AND5_17770 ( P2_R1312_U89 , P2_R1312_U88 , P2_R1312_U185 , P2_R1312_U168 , P2_R1312_U167 , P2_R1312_U166 );
and AND3_17771 ( P2_R1312_U90 , P2_R1312_U7 , P2_R1312_U187 , P2_R1312_U91 );
and AND2_17772 ( P2_R1312_U91 , P2_R1312_U9 , P2_R1312_U12 );
and AND3_17773 ( P2_R1312_U92 , P2_R1312_U167 , P2_R1312_U53 , P2_R1312_U166 );
and AND3_17774 ( P2_R1312_U93 , P2_U3151 , P2_R1312_U9 , P2_R1312_U12 );
and AND2_17775 ( P2_R1312_U94 , P2_U3127 , P2_R1312_U46 );
and AND2_17776 ( P2_R1312_U95 , P2_R1312_U194 , P2_R1312_U195 );
and AND3_17777 ( P2_R1312_U96 , P2_R1312_U167 , P2_R1312_U168 , P2_R1312_U166 );
and AND4_17778 ( P2_R1312_U97 , P2_R1312_U167 , P2_R1312_U29 , P2_R1312_U173 , P2_R1312_U168 );
and AND3_17779 ( P2_R1312_U98 , P2_R1312_U176 , P2_R1312_U174 , P2_U3140 );
and AND4_17780 ( P2_R1312_U99 , P2_R1312_U168 , P2_R1312_U31 , P2_R1312_U167 , P2_R1312_U166 );
and AND2_17781 ( P2_R1312_U100 , P2_R1312_U13 , P2_U3141 );
and AND4_17782 ( P2_R1312_U101 , P2_R1312_U167 , P2_R1312_U33 , P2_R1312_U177 , P2_R1312_U168 );
and AND2_17783 ( P2_R1312_U102 , P2_R1312_U103 , P2_R1312_U13 );
and AND2_17784 ( P2_R1312_U103 , P2_U3143 , P2_R1312_U178 );
and AND4_17785 ( P2_R1312_U104 , P2_R1312_U168 , P2_R1312_U49 , P2_R1312_U167 , P2_R1312_U166 );
and AND5_17786 ( P2_R1312_U105 , P2_R1312_U164 , P2_R1312_U47 , P2_R1312_U168 , P2_R1312_U167 , P2_R1312_U166 );
and AND4_17787 ( P2_R1312_U106 , P2_R1312_U167 , P2_R1312_U45 , P2_R1312_U169 , P2_R1312_U168 );
and AND2_17788 ( P2_R1312_U107 , P2_U3131 , P2_R1312_U16 );
and AND4_17789 ( P2_R1312_U108 , P2_R1312_U167 , P2_R1312_U41 , P2_R1312_U171 , P2_R1312_U168 );
and AND2_17790 ( P2_R1312_U109 , P2_U3134 , P2_R1312_U16 );
and AND4_17791 ( P2_R1312_U110 , P2_R1312_U167 , P2_R1312_U43 , P2_R1312_U170 , P2_R1312_U168 );
and AND5_17792 ( P2_R1312_U111 , P2_R1312_U11 , P2_R1312_U171 , P2_R1312_U17 , P2_R1312_U112 , P2_R1312_U166 );
and AND2_17793 ( P2_R1312_U112 , P2_U3135 , P2_R1312_U16 );
and AND3_17794 ( P2_R1312_U113 , P2_R1312_U167 , P2_R1312_U27 , P2_R1312_U166 );
and AND2_17795 ( P2_R1312_U114 , P2_U3137 , P2_R1312_U168 );
and AND4_17796 ( P2_R1312_U115 , P2_R1312_U157 , P2_R1312_U37 , P2_R1312_U167 , P2_R1312_U166 );
and AND5_17797 ( P2_R1312_U116 , P2_R1312_U156 , P2_R1312_U35 , P2_R1312_U157 , P2_R1312_U167 , P2_R1312_U166 );
and AND4_17798 ( P2_R1312_U117 , P2_R1312_U168 , P2_R1312_U42 , P2_R1312_U167 , P2_R1312_U166 );
and AND2_17799 ( P2_R1312_U118 , P2_U3133 , P2_R1312_U16 );
and AND4_17800 ( P2_R1312_U119 , P2_R1312_U168 , P2_R1312_U30 , P2_R1312_U167 , P2_R1312_U166 );
and AND3_17801 ( P2_R1312_U120 , P2_R1312_U174 , P2_R1312_U173 , P2_U3139 );
and AND4_17802 ( P2_R1312_U121 , P2_R1312_U168 , P2_R1312_U38 , P2_R1312_U167 , P2_R1312_U166 );
and AND5_17803 ( P2_R1312_U122 , P2_R1312_U161 , P2_R1312_U48 , P2_R1312_U164 , P2_R1312_U167 , P2_R1312_U166 );
and AND2_17804 ( P2_R1312_U123 , P2_R1312_U169 , P2_R1312_U168 );
and AND5_17805 ( P2_R1312_U124 , P2_R1312_U160 , P2_R1312_U44 , P2_R1312_U168 , P2_R1312_U167 , P2_R1312_U166 );
and AND2_17806 ( P2_R1312_U125 , P2_U3132 , P2_R1312_U16 );
and AND2_17807 ( P2_R1312_U126 , P2_R1312_U167 , P2_R1312_U39 );
and AND3_17808 ( P2_R1312_U127 , P2_R1312_U17 , P2_R1312_U168 , P2_R1312_U126 );
and AND2_17809 ( P2_R1312_U128 , P2_R1312_U6 , P2_U3136 );
and AND4_17810 ( P2_R1312_U129 , P2_R1312_U168 , P2_R1312_U28 , P2_R1312_U167 , P2_R1312_U166 );
and AND2_17811 ( P2_R1312_U130 , P2_U3138 , P2_R1312_U173 );
and AND4_17812 ( P2_R1312_U131 , P2_R1312_U168 , P2_R1312_U32 , P2_R1312_U167 , P2_R1312_U166 );
and AND2_17813 ( P2_R1312_U132 , P2_R1312_U133 , P2_R1312_U13 );
and AND2_17814 ( P2_R1312_U133 , P2_U3142 , P2_R1312_U177 );
and AND4_17815 ( P2_R1312_U134 , P2_R1312_U167 , P2_R1312_U34 , P2_R1312_U177 , P2_R1312_U168 );
and AND2_17816 ( P2_R1312_U135 , P2_R1312_U13 , P2_R1312_U136 );
and AND3_17817 ( P2_R1312_U136 , P2_R1312_U179 , P2_R1312_U178 , P2_U3144 );
and AND5_17818 ( P2_R1312_U137 , P2_R1312_U157 , P2_R1312_U156 , P2_R1312_U154 , P2_R1312_U36 , P2_R1312_U166 );
and AND4_17819 ( P2_R1312_U138 , P2_U3148 , P2_R1312_U8 , P2_R1312_U168 , P2_R1312_U167 );
and AND4_17820 ( P2_R1312_U139 , P2_R1312_U167 , P2_R1312_U52 , P2_R1312_U221 , P2_R1312_U168 );
and AND2_17821 ( P2_R1312_U140 , P2_U3150 , P2_R1312_U12 );
and AND2_17822 ( P2_R1312_U141 , P2_R1312_U181 , P2_R1312_U153 );
and AND2_17823 ( P2_R1312_U142 , P2_R1312_U192 , P2_R1312_U188 );
and AND3_17824 ( P2_R1312_U143 , P2_R1312_U199 , P2_R1312_U197 , P2_R1312_U198 );
and AND3_17825 ( P2_R1312_U144 , P2_R1312_U142 , P2_R1312_U141 , P2_R1312_U143 );
and AND2_17826 ( P2_R1312_U145 , P2_R1312_U203 , P2_R1312_U202 );
and AND2_17827 ( P2_R1312_U146 , P2_R1312_U205 , P2_R1312_U204 );
and AND5_17828 ( P2_R1312_U147 , P2_R1312_U201 , P2_R1312_U200 , P2_R1312_U145 , P2_R1312_U146 , P2_R1312_U206 );
and AND2_17829 ( P2_R1312_U148 , P2_R1312_U210 , P2_R1312_U209 );
and AND2_17830 ( P2_R1312_U149 , P2_R1312_U214 , P2_R1312_U215 );
and AND5_17831 ( P2_R1312_U150 , P2_R1312_U208 , P2_R1312_U207 , P2_R1312_U148 , P2_R1312_U149 , P2_R1312_U211 );
and AND4_17832 ( P2_R1312_U151 , P2_R1312_U219 , P2_R1312_U218 , P2_R1312_U217 , P2_R1312_U216 );
and AND3_17833 ( P2_R1312_U152 , P2_R1312_U10 , P2_R1312_U220 , P2_R1312_U222 );
nand NAND2_17834 ( P2_R1312_U153 , P2_R1312_U81 , P2_R1312_U191 );
nand NAND2_17835 ( P2_R1312_U154 , P2_U3115 , P2_R1312_U68 );
nand NAND2_17836 ( P2_R1312_U155 , P2_U3116 , P2_R1312_U78 );
nand NAND2_17837 ( P2_R1312_U156 , P2_U3114 , P2_R1312_U67 );
nand NAND2_17838 ( P2_R1312_U157 , P2_U3113 , P2_R1312_U71 );
nand NAND2_17839 ( P2_R1312_U158 , P2_U3104 , P2_R1312_U74 );
nand NAND2_17840 ( P2_R1312_U159 , P2_U3100 , P2_R1312_U73 );
nand NAND2_17841 ( P2_R1312_U160 , P2_U3099 , P2_R1312_U63 );
nand NAND2_17842 ( P2_R1312_U161 , P2_U3097 , P2_R1312_U62 );
nand NAND2_17843 ( P2_R1312_U162 , P2_U3098 , P2_R1312_U72 );
nand NAND2_17844 ( P2_R1312_U163 , P2_U3094 , P2_R1312_U23 );
nand NAND2_17845 ( P2_R1312_U164 , P2_U3096 , P2_R1312_U61 );
nand NAND2_17846 ( P2_R1312_U165 , P2_U3093 , P2_R1312_U56 );
nand NAND2_17847 ( P2_R1312_U166 , P2_U3090 , P2_R1312_U80 );
nand NAND2_17848 ( P2_R1312_U167 , P2_U3091 , P2_R1312_U24 );
nand NAND2_17849 ( P2_R1312_U168 , P2_U3092 , P2_R1312_U57 );
nand NAND2_17850 ( P2_R1312_U169 , P2_U3095 , P2_R1312_U55 );
nand NAND2_17851 ( P2_R1312_U170 , P2_U3102 , P2_R1312_U64 );
nand NAND2_17852 ( P2_R1312_U171 , P2_U3101 , P2_R1312_U69 );
nand NAND2_17853 ( P2_R1312_U172 , P2_U3103 , P2_R1312_U65 );
nand NAND2_17854 ( P2_R1312_U173 , P2_U3105 , P2_R1312_U66 );
nand NAND2_17855 ( P2_R1312_U174 , P2_U3106 , P2_R1312_U75 );
nand NAND2_17856 ( P2_R1312_U175 , P2_U3108 , P2_R1312_U58 );
nand NAND2_17857 ( P2_R1312_U176 , P2_U3107 , P2_R1312_U70 );
nand NAND2_17858 ( P2_R1312_U177 , P2_U3109 , P2_R1312_U59 );
nand NAND2_17859 ( P2_R1312_U178 , P2_U3110 , P2_R1312_U76 );
nand NAND2_17860 ( P2_R1312_U179 , P2_U3111 , P2_R1312_U60 );
nand NAND2_17861 ( P2_R1312_U180 , P2_U3112 , P2_R1312_U77 );
nand NAND4_17862 ( P2_R1312_U181 , P2_R1312_U8 , P2_R1312_U87 , P2_R1312_U15 , P2_R1312_U86 );
nand NAND2_17863 ( P2_R1312_U182 , P2_U3117 , P2_R1312_U50 );
nand NAND2_17864 ( P2_R1312_U183 , P2_U3118 , P2_R1312_U79 );
nand NAND2_17865 ( P2_R1312_U184 , P2_U3152 , P2_U3153 );
nand NAND2_17866 ( P2_R1312_U185 , P2_U3120 , P2_R1312_U184 );
nand NAND2_17867 ( P2_R1312_U186 , P2_U3119 , P2_R1312_U54 );
or OR2_17868 ( P2_R1312_U187 , P2_U3152 , P2_U3153 );
nand NAND3_17869 ( P2_R1312_U188 , P2_R1312_U15 , P2_R1312_U90 , P2_R1312_U89 );
nand NAND5_17870 ( P2_R1312_U189 , P2_R1312_U165 , P2_R1312_U40 , P2_R1312_U167 , P2_U3126 , P2_R1312_U168 );
nand NAND2_17871 ( P2_R1312_U190 , P2_U3123 , P2_R1312_U21 );
nand NAND2_17872 ( P2_R1312_U191 , P2_R1312_U190 , P2_R1312_U189 );
nand NAND5_17873 ( P2_R1312_U192 , P2_R1312_U8 , P2_R1312_U93 , P2_R1312_U168 , P2_R1312_U15 , P2_R1312_U92 );
nand NAND2_17874 ( P2_R1312_U193 , P2_R1312_U94 , P2_R1312_U16 );
nand NAND2_17875 ( P2_R1312_U194 , P2_U3125 , P2_R1312_U20 );
nand NAND2_17876 ( P2_R1312_U195 , P2_U3124 , P2_R1312_U22 );
nand NAND2_17877 ( P2_R1312_U196 , P2_R1312_U95 , P2_R1312_U193 );
nand NAND3_17878 ( P2_R1312_U197 , P2_R1312_U17 , P2_R1312_U196 , P2_R1312_U96 );
nand NAND4_17879 ( P2_R1312_U198 , P2_R1312_U98 , P2_R1312_U15 , P2_R1312_U166 , P2_R1312_U97 );
nand NAND3_17880 ( P2_R1312_U199 , P2_R1312_U100 , P2_R1312_U15 , P2_R1312_U99 );
nand NAND4_17881 ( P2_R1312_U200 , P2_R1312_U15 , P2_R1312_U102 , P2_R1312_U166 , P2_R1312_U101 );
nand NAND5_17882 ( P2_R1312_U201 , P2_U3128 , P2_R1312_U16 , P2_R1312_U17 , P2_R1312_U169 , P2_R1312_U104 );
nand NAND5_17883 ( P2_R1312_U202 , P2_U3129 , P2_R1312_U16 , P2_R1312_U17 , P2_R1312_U169 , P2_R1312_U105 );
nand NAND5_17884 ( P2_R1312_U203 , P2_R1312_U17 , P2_R1312_U14 , P2_R1312_U107 , P2_R1312_U166 , P2_R1312_U106 );
nand NAND5_17885 ( P2_R1312_U204 , P2_R1312_U17 , P2_R1312_U11 , P2_R1312_U109 , P2_R1312_U166 , P2_R1312_U108 );
nand NAND2_17886 ( P2_R1312_U205 , P2_R1312_U110 , P2_R1312_U111 );
nand NAND3_17887 ( P2_R1312_U206 , P2_R1312_U114 , P2_R1312_U15 , P2_R1312_U113 );
nand NAND5_17888 ( P2_R1312_U207 , P2_U3146 , P2_R1312_U8 , P2_R1312_U168 , P2_R1312_U15 , P2_R1312_U115 );
nand NAND5_17889 ( P2_R1312_U208 , P2_U3147 , P2_R1312_U8 , P2_R1312_U168 , P2_R1312_U15 , P2_R1312_U116 );
nand NAND4_17890 ( P2_R1312_U209 , P2_R1312_U17 , P2_R1312_U11 , P2_R1312_U118 , P2_R1312_U117 );
nand NAND3_17891 ( P2_R1312_U210 , P2_R1312_U120 , P2_R1312_U15 , P2_R1312_U119 );
nand NAND4_17892 ( P2_R1312_U211 , P2_R1312_U8 , P2_U3145 , P2_R1312_U15 , P2_R1312_U121 );
nand NAND3_17893 ( P2_R1312_U212 , P2_R1312_U227 , P2_R1312_U226 , P2_R1312_U223 );
nand NAND3_17894 ( P2_R1312_U213 , P2_R1312_U17 , P2_U3122 , P2_R1312_U19 );
nand NAND5_17895 ( P2_R1312_U214 , P2_U3130 , P2_R1312_U16 , P2_R1312_U17 , P2_R1312_U123 , P2_R1312_U122 );
nand NAND5_17896 ( P2_R1312_U215 , P2_R1312_U14 , P2_R1312_U169 , P2_R1312_U17 , P2_R1312_U125 , P2_R1312_U124 );
nand NAND5_17897 ( P2_R1312_U216 , P2_R1312_U11 , P2_R1312_U128 , P2_R1312_U16 , P2_R1312_U166 , P2_R1312_U127 );
nand NAND3_17898 ( P2_R1312_U217 , P2_R1312_U130 , P2_R1312_U15 , P2_R1312_U129 );
nand NAND3_17899 ( P2_R1312_U218 , P2_R1312_U15 , P2_R1312_U132 , P2_R1312_U131 );
nand NAND4_17900 ( P2_R1312_U219 , P2_R1312_U15 , P2_R1312_U135 , P2_R1312_U166 , P2_R1312_U134 );
nand NAND3_17901 ( P2_R1312_U220 , P2_R1312_U15 , P2_R1312_U138 , P2_R1312_U137 );
nand NAND2_17902 ( P2_R1312_U221 , P2_U3117 , P2_R1312_U50 );
nand NAND5_17903 ( P2_R1312_U222 , P2_R1312_U8 , P2_R1312_U140 , P2_R1312_U15 , P2_R1312_U166 , P2_R1312_U139 );
nand NAND2_17904 ( P2_R1312_U223 , P2_U3121 , P2_U3089 );
nand NAND2_17905 ( P2_R1312_U224 , P2_U3089 , P2_R1312_U26 );
nand NAND2_17906 ( P2_R1312_U225 , P2_U3121 , P2_R1312_U25 );
or OR2_17907 ( P2_R1312_U226 , P2_U3154 , P2_U3121 );
nand NAND2_17908 ( P2_R1312_U227 , P2_U3154 , P2_R1312_U25 );
not NOT1_17909 ( P2_R1335_U6 , P2_U3061 );
not NOT1_17910 ( P2_R1335_U7 , P2_U3058 );
and AND2_17911 ( P2_R1335_U8 , P2_R1335_U10 , P2_R1335_U9 );
nand NAND2_17912 ( P2_R1335_U9 , P2_U3058 , P2_R1335_U6 );
nand NAND2_17913 ( P2_R1335_U10 , P2_U3061 , P2_R1335_U7 );
and AND2_17914 ( P2_R1209_U4 , P2_R1209_U95 , P2_R1209_U94 );
and AND2_17915 ( P2_R1209_U5 , P2_R1209_U96 , P2_R1209_U97 );
and AND2_17916 ( P2_R1209_U6 , P2_R1209_U113 , P2_R1209_U112 );
and AND2_17917 ( P2_R1209_U7 , P2_R1209_U155 , P2_R1209_U154 );
and AND2_17918 ( P2_R1209_U8 , P2_R1209_U164 , P2_R1209_U163 );
and AND2_17919 ( P2_R1209_U9 , P2_R1209_U182 , P2_R1209_U181 );
and AND2_17920 ( P2_R1209_U10 , P2_R1209_U218 , P2_R1209_U215 );
and AND2_17921 ( P2_R1209_U11 , P2_R1209_U211 , P2_R1209_U208 );
and AND2_17922 ( P2_R1209_U12 , P2_R1209_U202 , P2_R1209_U199 );
and AND2_17923 ( P2_R1209_U13 , P2_R1209_U196 , P2_R1209_U192 );
and AND2_17924 ( P2_R1209_U14 , P2_R1209_U151 , P2_R1209_U148 );
and AND2_17925 ( P2_R1209_U15 , P2_R1209_U143 , P2_R1209_U140 );
and AND2_17926 ( P2_R1209_U16 , P2_R1209_U129 , P2_R1209_U126 );
not NOT1_17927 ( P2_R1209_U17 , P2_REG1_REG_6_ );
not NOT1_17928 ( P2_R1209_U18 , P2_U3446 );
not NOT1_17929 ( P2_R1209_U19 , P2_U3449 );
nand NAND2_17930 ( P2_R1209_U20 , P2_U3446 , P2_REG1_REG_6_ );
not NOT1_17931 ( P2_R1209_U21 , P2_REG1_REG_7_ );
not NOT1_17932 ( P2_R1209_U22 , P2_REG1_REG_4_ );
not NOT1_17933 ( P2_R1209_U23 , P2_U3440 );
not NOT1_17934 ( P2_R1209_U24 , P2_U3443 );
not NOT1_17935 ( P2_R1209_U25 , P2_REG1_REG_2_ );
not NOT1_17936 ( P2_R1209_U26 , P2_U3434 );
not NOT1_17937 ( P2_R1209_U27 , P2_REG1_REG_0_ );
not NOT1_17938 ( P2_R1209_U28 , P2_U3425 );
nand NAND2_17939 ( P2_R1209_U29 , P2_U3425 , P2_REG1_REG_0_ );
not NOT1_17940 ( P2_R1209_U30 , P2_REG1_REG_3_ );
not NOT1_17941 ( P2_R1209_U31 , P2_U3437 );
nand NAND2_17942 ( P2_R1209_U32 , P2_U3440 , P2_REG1_REG_4_ );
not NOT1_17943 ( P2_R1209_U33 , P2_REG1_REG_5_ );
not NOT1_17944 ( P2_R1209_U34 , P2_REG1_REG_8_ );
not NOT1_17945 ( P2_R1209_U35 , P2_U3452 );
not NOT1_17946 ( P2_R1209_U36 , P2_U3455 );
not NOT1_17947 ( P2_R1209_U37 , P2_REG1_REG_9_ );
nand NAND2_17948 ( P2_R1209_U38 , P2_R1209_U49 , P2_R1209_U121 );
nand NAND3_17949 ( P2_R1209_U39 , P2_R1209_U110 , P2_R1209_U108 , P2_R1209_U109 );
nand NAND2_17950 ( P2_R1209_U40 , P2_R1209_U98 , P2_R1209_U99 );
nand NAND2_17951 ( P2_R1209_U41 , P2_REG1_REG_1_ , P2_U3431 );
nand NAND3_17952 ( P2_R1209_U42 , P2_R1209_U136 , P2_R1209_U134 , P2_R1209_U135 );
nand NAND2_17953 ( P2_R1209_U43 , P2_R1209_U132 , P2_R1209_U131 );
not NOT1_17954 ( P2_R1209_U44 , P2_REG1_REG_16_ );
not NOT1_17955 ( P2_R1209_U45 , P2_U3476 );
not NOT1_17956 ( P2_R1209_U46 , P2_U3479 );
nand NAND2_17957 ( P2_R1209_U47 , P2_U3476 , P2_REG1_REG_16_ );
not NOT1_17958 ( P2_R1209_U48 , P2_REG1_REG_17_ );
nand NAND2_17959 ( P2_R1209_U49 , P2_U3452 , P2_REG1_REG_8_ );
not NOT1_17960 ( P2_R1209_U50 , P2_REG1_REG_10_ );
not NOT1_17961 ( P2_R1209_U51 , P2_U3458 );
not NOT1_17962 ( P2_R1209_U52 , P2_REG1_REG_12_ );
not NOT1_17963 ( P2_R1209_U53 , P2_U3464 );
not NOT1_17964 ( P2_R1209_U54 , P2_REG1_REG_11_ );
not NOT1_17965 ( P2_R1209_U55 , P2_U3461 );
nand NAND2_17966 ( P2_R1209_U56 , P2_U3461 , P2_REG1_REG_11_ );
not NOT1_17967 ( P2_R1209_U57 , P2_REG1_REG_13_ );
not NOT1_17968 ( P2_R1209_U58 , P2_U3467 );
not NOT1_17969 ( P2_R1209_U59 , P2_REG1_REG_14_ );
not NOT1_17970 ( P2_R1209_U60 , P2_U3470 );
not NOT1_17971 ( P2_R1209_U61 , P2_REG1_REG_15_ );
not NOT1_17972 ( P2_R1209_U62 , P2_U3473 );
not NOT1_17973 ( P2_R1209_U63 , P2_REG1_REG_18_ );
not NOT1_17974 ( P2_R1209_U64 , P2_U3482 );
nand NAND3_17975 ( P2_R1209_U65 , P2_R1209_U186 , P2_R1209_U185 , P2_R1209_U187 );
nand NAND2_17976 ( P2_R1209_U66 , P2_R1209_U179 , P2_R1209_U178 );
nand NAND2_17977 ( P2_R1209_U67 , P2_R1209_U56 , P2_R1209_U204 );
nand NAND2_17978 ( P2_R1209_U68 , P2_R1209_U259 , P2_R1209_U258 );
nand NAND2_17979 ( P2_R1209_U69 , P2_R1209_U308 , P2_R1209_U307 );
nand NAND2_17980 ( P2_R1209_U70 , P2_R1209_U231 , P2_R1209_U230 );
nand NAND2_17981 ( P2_R1209_U71 , P2_R1209_U236 , P2_R1209_U235 );
nand NAND2_17982 ( P2_R1209_U72 , P2_R1209_U243 , P2_R1209_U242 );
nand NAND2_17983 ( P2_R1209_U73 , P2_R1209_U250 , P2_R1209_U249 );
nand NAND2_17984 ( P2_R1209_U74 , P2_R1209_U255 , P2_R1209_U254 );
nand NAND2_17985 ( P2_R1209_U75 , P2_R1209_U271 , P2_R1209_U270 );
nand NAND2_17986 ( P2_R1209_U76 , P2_R1209_U278 , P2_R1209_U277 );
nand NAND2_17987 ( P2_R1209_U77 , P2_R1209_U285 , P2_R1209_U284 );
nand NAND2_17988 ( P2_R1209_U78 , P2_R1209_U292 , P2_R1209_U291 );
nand NAND2_17989 ( P2_R1209_U79 , P2_R1209_U299 , P2_R1209_U298 );
nand NAND2_17990 ( P2_R1209_U80 , P2_R1209_U304 , P2_R1209_U303 );
nand NAND3_17991 ( P2_R1209_U81 , P2_R1209_U117 , P2_R1209_U116 , P2_R1209_U118 );
nand NAND2_17992 ( P2_R1209_U82 , P2_R1209_U133 , P2_R1209_U145 );
nand NAND2_17993 ( P2_R1209_U83 , P2_R1209_U41 , P2_R1209_U152 );
not NOT1_17994 ( P2_R1209_U84 , P2_U3424 );
not NOT1_17995 ( P2_R1209_U85 , P2_REG1_REG_19_ );
nand NAND2_17996 ( P2_R1209_U86 , P2_R1209_U175 , P2_R1209_U174 );
nand NAND2_17997 ( P2_R1209_U87 , P2_R1209_U171 , P2_R1209_U170 );
nand NAND2_17998 ( P2_R1209_U88 , P2_R1209_U161 , P2_R1209_U160 );
not NOT1_17999 ( P2_R1209_U89 , P2_R1209_U32 );
nand NAND2_18000 ( P2_R1209_U90 , P2_REG1_REG_9_ , P2_U3455 );
nand NAND2_18001 ( P2_R1209_U91 , P2_U3464 , P2_REG1_REG_12_ );
not NOT1_18002 ( P2_R1209_U92 , P2_R1209_U56 );
not NOT1_18003 ( P2_R1209_U93 , P2_R1209_U49 );
or OR2_18004 ( P2_R1209_U94 , P2_U3443 , P2_REG1_REG_5_ );
or OR2_18005 ( P2_R1209_U95 , P2_U3440 , P2_REG1_REG_4_ );
or OR2_18006 ( P2_R1209_U96 , P2_REG1_REG_3_ , P2_U3437 );
or OR2_18007 ( P2_R1209_U97 , P2_REG1_REG_2_ , P2_U3434 );
not NOT1_18008 ( P2_R1209_U98 , P2_R1209_U29 );
or OR2_18009 ( P2_R1209_U99 , P2_REG1_REG_1_ , P2_U3431 );
not NOT1_18010 ( P2_R1209_U100 , P2_R1209_U40 );
not NOT1_18011 ( P2_R1209_U101 , P2_R1209_U41 );
nand NAND2_18012 ( P2_R1209_U102 , P2_R1209_U40 , P2_R1209_U41 );
nand NAND3_18013 ( P2_R1209_U103 , P2_REG1_REG_2_ , P2_U3434 , P2_R1209_U96 );
nand NAND2_18014 ( P2_R1209_U104 , P2_R1209_U5 , P2_R1209_U102 );
nand NAND2_18015 ( P2_R1209_U105 , P2_U3437 , P2_REG1_REG_3_ );
nand NAND3_18016 ( P2_R1209_U106 , P2_R1209_U105 , P2_R1209_U103 , P2_R1209_U104 );
nand NAND2_18017 ( P2_R1209_U107 , P2_R1209_U33 , P2_R1209_U32 );
nand NAND2_18018 ( P2_R1209_U108 , P2_U3443 , P2_R1209_U107 );
nand NAND2_18019 ( P2_R1209_U109 , P2_R1209_U4 , P2_R1209_U106 );
nand NAND2_18020 ( P2_R1209_U110 , P2_REG1_REG_5_ , P2_R1209_U89 );
not NOT1_18021 ( P2_R1209_U111 , P2_R1209_U39 );
or OR2_18022 ( P2_R1209_U112 , P2_U3449 , P2_REG1_REG_7_ );
or OR2_18023 ( P2_R1209_U113 , P2_U3446 , P2_REG1_REG_6_ );
not NOT1_18024 ( P2_R1209_U114 , P2_R1209_U20 );
nand NAND2_18025 ( P2_R1209_U115 , P2_R1209_U21 , P2_R1209_U20 );
nand NAND2_18026 ( P2_R1209_U116 , P2_U3449 , P2_R1209_U115 );
nand NAND2_18027 ( P2_R1209_U117 , P2_REG1_REG_7_ , P2_R1209_U114 );
nand NAND2_18028 ( P2_R1209_U118 , P2_R1209_U6 , P2_R1209_U39 );
not NOT1_18029 ( P2_R1209_U119 , P2_R1209_U81 );
or OR2_18030 ( P2_R1209_U120 , P2_REG1_REG_8_ , P2_U3452 );
nand NAND2_18031 ( P2_R1209_U121 , P2_R1209_U120 , P2_R1209_U81 );
not NOT1_18032 ( P2_R1209_U122 , P2_R1209_U38 );
or OR2_18033 ( P2_R1209_U123 , P2_U3455 , P2_REG1_REG_9_ );
or OR2_18034 ( P2_R1209_U124 , P2_REG1_REG_6_ , P2_U3446 );
nand NAND2_18035 ( P2_R1209_U125 , P2_R1209_U124 , P2_R1209_U39 );
nand NAND4_18036 ( P2_R1209_U126 , P2_R1209_U238 , P2_R1209_U237 , P2_R1209_U20 , P2_R1209_U125 );
nand NAND2_18037 ( P2_R1209_U127 , P2_R1209_U111 , P2_R1209_U20 );
nand NAND2_18038 ( P2_R1209_U128 , P2_REG1_REG_7_ , P2_U3449 );
nand NAND3_18039 ( P2_R1209_U129 , P2_R1209_U128 , P2_R1209_U6 , P2_R1209_U127 );
or OR2_18040 ( P2_R1209_U130 , P2_U3446 , P2_REG1_REG_6_ );
nand NAND2_18041 ( P2_R1209_U131 , P2_R1209_U101 , P2_R1209_U97 );
nand NAND2_18042 ( P2_R1209_U132 , P2_U3434 , P2_REG1_REG_2_ );
not NOT1_18043 ( P2_R1209_U133 , P2_R1209_U43 );
nand NAND2_18044 ( P2_R1209_U134 , P2_R1209_U100 , P2_R1209_U5 );
nand NAND2_18045 ( P2_R1209_U135 , P2_R1209_U43 , P2_R1209_U96 );
nand NAND2_18046 ( P2_R1209_U136 , P2_U3437 , P2_REG1_REG_3_ );
not NOT1_18047 ( P2_R1209_U137 , P2_R1209_U42 );
or OR2_18048 ( P2_R1209_U138 , P2_REG1_REG_4_ , P2_U3440 );
nand NAND2_18049 ( P2_R1209_U139 , P2_R1209_U138 , P2_R1209_U42 );
nand NAND4_18050 ( P2_R1209_U140 , P2_R1209_U245 , P2_R1209_U244 , P2_R1209_U32 , P2_R1209_U139 );
nand NAND2_18051 ( P2_R1209_U141 , P2_R1209_U137 , P2_R1209_U32 );
nand NAND2_18052 ( P2_R1209_U142 , P2_REG1_REG_5_ , P2_U3443 );
nand NAND3_18053 ( P2_R1209_U143 , P2_R1209_U142 , P2_R1209_U4 , P2_R1209_U141 );
or OR2_18054 ( P2_R1209_U144 , P2_U3440 , P2_REG1_REG_4_ );
nand NAND2_18055 ( P2_R1209_U145 , P2_R1209_U100 , P2_R1209_U97 );
not NOT1_18056 ( P2_R1209_U146 , P2_R1209_U82 );
nand NAND2_18057 ( P2_R1209_U147 , P2_U3437 , P2_REG1_REG_3_ );
nand NAND4_18058 ( P2_R1209_U148 , P2_R1209_U257 , P2_R1209_U256 , P2_R1209_U41 , P2_R1209_U40 );
nand NAND2_18059 ( P2_R1209_U149 , P2_R1209_U41 , P2_R1209_U40 );
nand NAND2_18060 ( P2_R1209_U150 , P2_U3434 , P2_REG1_REG_2_ );
nand NAND3_18061 ( P2_R1209_U151 , P2_R1209_U150 , P2_R1209_U97 , P2_R1209_U149 );
or OR2_18062 ( P2_R1209_U152 , P2_REG1_REG_1_ , P2_U3431 );
not NOT1_18063 ( P2_R1209_U153 , P2_R1209_U83 );
or OR2_18064 ( P2_R1209_U154 , P2_U3455 , P2_REG1_REG_9_ );
or OR2_18065 ( P2_R1209_U155 , P2_U3458 , P2_REG1_REG_10_ );
nand NAND2_18066 ( P2_R1209_U156 , P2_R1209_U93 , P2_R1209_U7 );
nand NAND2_18067 ( P2_R1209_U157 , P2_U3458 , P2_REG1_REG_10_ );
nand NAND3_18068 ( P2_R1209_U158 , P2_R1209_U157 , P2_R1209_U90 , P2_R1209_U156 );
or OR2_18069 ( P2_R1209_U159 , P2_REG1_REG_10_ , P2_U3458 );
nand NAND3_18070 ( P2_R1209_U160 , P2_R1209_U120 , P2_R1209_U7 , P2_R1209_U81 );
nand NAND2_18071 ( P2_R1209_U161 , P2_R1209_U159 , P2_R1209_U158 );
not NOT1_18072 ( P2_R1209_U162 , P2_R1209_U88 );
or OR2_18073 ( P2_R1209_U163 , P2_U3467 , P2_REG1_REG_13_ );
or OR2_18074 ( P2_R1209_U164 , P2_U3464 , P2_REG1_REG_12_ );
nand NAND2_18075 ( P2_R1209_U165 , P2_R1209_U92 , P2_R1209_U8 );
nand NAND2_18076 ( P2_R1209_U166 , P2_U3467 , P2_REG1_REG_13_ );
nand NAND3_18077 ( P2_R1209_U167 , P2_R1209_U166 , P2_R1209_U91 , P2_R1209_U165 );
or OR2_18078 ( P2_R1209_U168 , P2_REG1_REG_11_ , P2_U3461 );
or OR2_18079 ( P2_R1209_U169 , P2_REG1_REG_13_ , P2_U3467 );
nand NAND3_18080 ( P2_R1209_U170 , P2_R1209_U168 , P2_R1209_U8 , P2_R1209_U88 );
nand NAND2_18081 ( P2_R1209_U171 , P2_R1209_U169 , P2_R1209_U167 );
not NOT1_18082 ( P2_R1209_U172 , P2_R1209_U87 );
or OR2_18083 ( P2_R1209_U173 , P2_REG1_REG_14_ , P2_U3470 );
nand NAND2_18084 ( P2_R1209_U174 , P2_R1209_U173 , P2_R1209_U87 );
nand NAND2_18085 ( P2_R1209_U175 , P2_U3470 , P2_REG1_REG_14_ );
not NOT1_18086 ( P2_R1209_U176 , P2_R1209_U86 );
or OR2_18087 ( P2_R1209_U177 , P2_REG1_REG_15_ , P2_U3473 );
nand NAND2_18088 ( P2_R1209_U178 , P2_R1209_U177 , P2_R1209_U86 );
nand NAND2_18089 ( P2_R1209_U179 , P2_U3473 , P2_REG1_REG_15_ );
not NOT1_18090 ( P2_R1209_U180 , P2_R1209_U66 );
or OR2_18091 ( P2_R1209_U181 , P2_U3479 , P2_REG1_REG_17_ );
or OR2_18092 ( P2_R1209_U182 , P2_U3476 , P2_REG1_REG_16_ );
not NOT1_18093 ( P2_R1209_U183 , P2_R1209_U47 );
nand NAND2_18094 ( P2_R1209_U184 , P2_R1209_U48 , P2_R1209_U47 );
nand NAND2_18095 ( P2_R1209_U185 , P2_U3479 , P2_R1209_U184 );
nand NAND2_18096 ( P2_R1209_U186 , P2_REG1_REG_17_ , P2_R1209_U183 );
nand NAND2_18097 ( P2_R1209_U187 , P2_R1209_U9 , P2_R1209_U66 );
not NOT1_18098 ( P2_R1209_U188 , P2_R1209_U65 );
or OR2_18099 ( P2_R1209_U189 , P2_REG1_REG_18_ , P2_U3482 );
nand NAND2_18100 ( P2_R1209_U190 , P2_R1209_U189 , P2_R1209_U65 );
nand NAND2_18101 ( P2_R1209_U191 , P2_U3482 , P2_REG1_REG_18_ );
nand NAND4_18102 ( P2_R1209_U192 , P2_R1209_U261 , P2_R1209_U260 , P2_R1209_U191 , P2_R1209_U190 );
nand NAND2_18103 ( P2_R1209_U193 , P2_U3482 , P2_REG1_REG_18_ );
nand NAND2_18104 ( P2_R1209_U194 , P2_R1209_U188 , P2_R1209_U193 );
or OR2_18105 ( P2_R1209_U195 , P2_U3482 , P2_REG1_REG_18_ );
nand NAND3_18106 ( P2_R1209_U196 , P2_R1209_U195 , P2_R1209_U264 , P2_R1209_U194 );
or OR2_18107 ( P2_R1209_U197 , P2_REG1_REG_16_ , P2_U3476 );
nand NAND2_18108 ( P2_R1209_U198 , P2_R1209_U197 , P2_R1209_U66 );
nand NAND4_18109 ( P2_R1209_U199 , P2_R1209_U273 , P2_R1209_U272 , P2_R1209_U47 , P2_R1209_U198 );
nand NAND2_18110 ( P2_R1209_U200 , P2_R1209_U180 , P2_R1209_U47 );
nand NAND2_18111 ( P2_R1209_U201 , P2_REG1_REG_17_ , P2_U3479 );
nand NAND3_18112 ( P2_R1209_U202 , P2_R1209_U201 , P2_R1209_U9 , P2_R1209_U200 );
or OR2_18113 ( P2_R1209_U203 , P2_U3476 , P2_REG1_REG_16_ );
nand NAND2_18114 ( P2_R1209_U204 , P2_R1209_U168 , P2_R1209_U88 );
not NOT1_18115 ( P2_R1209_U205 , P2_R1209_U67 );
or OR2_18116 ( P2_R1209_U206 , P2_REG1_REG_12_ , P2_U3464 );
nand NAND2_18117 ( P2_R1209_U207 , P2_R1209_U206 , P2_R1209_U67 );
nand NAND4_18118 ( P2_R1209_U208 , P2_R1209_U294 , P2_R1209_U293 , P2_R1209_U91 , P2_R1209_U207 );
nand NAND2_18119 ( P2_R1209_U209 , P2_R1209_U205 , P2_R1209_U91 );
nand NAND2_18120 ( P2_R1209_U210 , P2_U3467 , P2_REG1_REG_13_ );
nand NAND3_18121 ( P2_R1209_U211 , P2_R1209_U210 , P2_R1209_U8 , P2_R1209_U209 );
or OR2_18122 ( P2_R1209_U212 , P2_U3464 , P2_REG1_REG_12_ );
or OR2_18123 ( P2_R1209_U213 , P2_REG1_REG_9_ , P2_U3455 );
nand NAND2_18124 ( P2_R1209_U214 , P2_R1209_U213 , P2_R1209_U38 );
nand NAND4_18125 ( P2_R1209_U215 , P2_R1209_U306 , P2_R1209_U305 , P2_R1209_U90 , P2_R1209_U214 );
nand NAND2_18126 ( P2_R1209_U216 , P2_R1209_U122 , P2_R1209_U90 );
nand NAND2_18127 ( P2_R1209_U217 , P2_U3458 , P2_REG1_REG_10_ );
nand NAND3_18128 ( P2_R1209_U218 , P2_R1209_U217 , P2_R1209_U7 , P2_R1209_U216 );
nand NAND2_18129 ( P2_R1209_U219 , P2_R1209_U123 , P2_R1209_U90 );
nand NAND2_18130 ( P2_R1209_U220 , P2_R1209_U120 , P2_R1209_U49 );
nand NAND2_18131 ( P2_R1209_U221 , P2_R1209_U130 , P2_R1209_U20 );
nand NAND2_18132 ( P2_R1209_U222 , P2_R1209_U144 , P2_R1209_U32 );
nand NAND2_18133 ( P2_R1209_U223 , P2_R1209_U147 , P2_R1209_U96 );
nand NAND2_18134 ( P2_R1209_U224 , P2_R1209_U203 , P2_R1209_U47 );
nand NAND2_18135 ( P2_R1209_U225 , P2_R1209_U212 , P2_R1209_U91 );
nand NAND2_18136 ( P2_R1209_U226 , P2_R1209_U168 , P2_R1209_U56 );
nand NAND2_18137 ( P2_R1209_U227 , P2_U3455 , P2_R1209_U37 );
nand NAND2_18138 ( P2_R1209_U228 , P2_REG1_REG_9_ , P2_R1209_U36 );
nand NAND2_18139 ( P2_R1209_U229 , P2_R1209_U228 , P2_R1209_U227 );
nand NAND2_18140 ( P2_R1209_U230 , P2_R1209_U219 , P2_R1209_U38 );
nand NAND2_18141 ( P2_R1209_U231 , P2_R1209_U229 , P2_R1209_U122 );
nand NAND2_18142 ( P2_R1209_U232 , P2_U3452 , P2_R1209_U34 );
nand NAND2_18143 ( P2_R1209_U233 , P2_REG1_REG_8_ , P2_R1209_U35 );
nand NAND2_18144 ( P2_R1209_U234 , P2_R1209_U233 , P2_R1209_U232 );
nand NAND2_18145 ( P2_R1209_U235 , P2_R1209_U220 , P2_R1209_U81 );
nand NAND2_18146 ( P2_R1209_U236 , P2_R1209_U119 , P2_R1209_U234 );
nand NAND2_18147 ( P2_R1209_U237 , P2_U3449 , P2_R1209_U21 );
nand NAND2_18148 ( P2_R1209_U238 , P2_REG1_REG_7_ , P2_R1209_U19 );
nand NAND2_18149 ( P2_R1209_U239 , P2_U3446 , P2_R1209_U17 );
nand NAND2_18150 ( P2_R1209_U240 , P2_REG1_REG_6_ , P2_R1209_U18 );
nand NAND2_18151 ( P2_R1209_U241 , P2_R1209_U240 , P2_R1209_U239 );
nand NAND2_18152 ( P2_R1209_U242 , P2_R1209_U221 , P2_R1209_U39 );
nand NAND2_18153 ( P2_R1209_U243 , P2_R1209_U241 , P2_R1209_U111 );
nand NAND2_18154 ( P2_R1209_U244 , P2_U3443 , P2_R1209_U33 );
nand NAND2_18155 ( P2_R1209_U245 , P2_REG1_REG_5_ , P2_R1209_U24 );
nand NAND2_18156 ( P2_R1209_U246 , P2_U3440 , P2_R1209_U22 );
nand NAND2_18157 ( P2_R1209_U247 , P2_REG1_REG_4_ , P2_R1209_U23 );
nand NAND2_18158 ( P2_R1209_U248 , P2_R1209_U247 , P2_R1209_U246 );
nand NAND2_18159 ( P2_R1209_U249 , P2_R1209_U222 , P2_R1209_U42 );
nand NAND2_18160 ( P2_R1209_U250 , P2_R1209_U248 , P2_R1209_U137 );
nand NAND2_18161 ( P2_R1209_U251 , P2_U3437 , P2_R1209_U30 );
nand NAND2_18162 ( P2_R1209_U252 , P2_REG1_REG_3_ , P2_R1209_U31 );
nand NAND2_18163 ( P2_R1209_U253 , P2_R1209_U252 , P2_R1209_U251 );
nand NAND2_18164 ( P2_R1209_U254 , P2_R1209_U223 , P2_R1209_U82 );
nand NAND2_18165 ( P2_R1209_U255 , P2_R1209_U146 , P2_R1209_U253 );
nand NAND2_18166 ( P2_R1209_U256 , P2_U3434 , P2_R1209_U25 );
nand NAND2_18167 ( P2_R1209_U257 , P2_REG1_REG_2_ , P2_R1209_U26 );
nand NAND2_18168 ( P2_R1209_U258 , P2_R1209_U98 , P2_R1209_U83 );
nand NAND2_18169 ( P2_R1209_U259 , P2_R1209_U153 , P2_R1209_U29 );
nand NAND2_18170 ( P2_R1209_U260 , P2_U3424 , P2_R1209_U85 );
nand NAND2_18171 ( P2_R1209_U261 , P2_REG1_REG_19_ , P2_R1209_U84 );
nand NAND2_18172 ( P2_R1209_U262 , P2_U3424 , P2_R1209_U85 );
nand NAND2_18173 ( P2_R1209_U263 , P2_REG1_REG_19_ , P2_R1209_U84 );
nand NAND2_18174 ( P2_R1209_U264 , P2_R1209_U263 , P2_R1209_U262 );
nand NAND2_18175 ( P2_R1209_U265 , P2_U3482 , P2_R1209_U63 );
nand NAND2_18176 ( P2_R1209_U266 , P2_REG1_REG_18_ , P2_R1209_U64 );
nand NAND2_18177 ( P2_R1209_U267 , P2_U3482 , P2_R1209_U63 );
nand NAND2_18178 ( P2_R1209_U268 , P2_REG1_REG_18_ , P2_R1209_U64 );
nand NAND2_18179 ( P2_R1209_U269 , P2_R1209_U268 , P2_R1209_U267 );
nand NAND3_18180 ( P2_R1209_U270 , P2_R1209_U266 , P2_R1209_U265 , P2_R1209_U65 );
nand NAND2_18181 ( P2_R1209_U271 , P2_R1209_U269 , P2_R1209_U188 );
nand NAND2_18182 ( P2_R1209_U272 , P2_U3479 , P2_R1209_U48 );
nand NAND2_18183 ( P2_R1209_U273 , P2_REG1_REG_17_ , P2_R1209_U46 );
nand NAND2_18184 ( P2_R1209_U274 , P2_U3476 , P2_R1209_U44 );
nand NAND2_18185 ( P2_R1209_U275 , P2_REG1_REG_16_ , P2_R1209_U45 );
nand NAND2_18186 ( P2_R1209_U276 , P2_R1209_U275 , P2_R1209_U274 );
nand NAND2_18187 ( P2_R1209_U277 , P2_R1209_U224 , P2_R1209_U66 );
nand NAND2_18188 ( P2_R1209_U278 , P2_R1209_U276 , P2_R1209_U180 );
nand NAND2_18189 ( P2_R1209_U279 , P2_U3473 , P2_R1209_U61 );
nand NAND2_18190 ( P2_R1209_U280 , P2_REG1_REG_15_ , P2_R1209_U62 );
nand NAND2_18191 ( P2_R1209_U281 , P2_U3473 , P2_R1209_U61 );
nand NAND2_18192 ( P2_R1209_U282 , P2_REG1_REG_15_ , P2_R1209_U62 );
nand NAND2_18193 ( P2_R1209_U283 , P2_R1209_U282 , P2_R1209_U281 );
nand NAND3_18194 ( P2_R1209_U284 , P2_R1209_U280 , P2_R1209_U279 , P2_R1209_U86 );
nand NAND2_18195 ( P2_R1209_U285 , P2_R1209_U176 , P2_R1209_U283 );
nand NAND2_18196 ( P2_R1209_U286 , P2_U3470 , P2_R1209_U59 );
nand NAND2_18197 ( P2_R1209_U287 , P2_REG1_REG_14_ , P2_R1209_U60 );
nand NAND2_18198 ( P2_R1209_U288 , P2_U3470 , P2_R1209_U59 );
nand NAND2_18199 ( P2_R1209_U289 , P2_REG1_REG_14_ , P2_R1209_U60 );
nand NAND2_18200 ( P2_R1209_U290 , P2_R1209_U289 , P2_R1209_U288 );
nand NAND3_18201 ( P2_R1209_U291 , P2_R1209_U287 , P2_R1209_U286 , P2_R1209_U87 );
nand NAND2_18202 ( P2_R1209_U292 , P2_R1209_U172 , P2_R1209_U290 );
nand NAND2_18203 ( P2_R1209_U293 , P2_U3467 , P2_R1209_U57 );
nand NAND2_18204 ( P2_R1209_U294 , P2_REG1_REG_13_ , P2_R1209_U58 );
nand NAND2_18205 ( P2_R1209_U295 , P2_U3464 , P2_R1209_U52 );
nand NAND2_18206 ( P2_R1209_U296 , P2_REG1_REG_12_ , P2_R1209_U53 );
nand NAND2_18207 ( P2_R1209_U297 , P2_R1209_U296 , P2_R1209_U295 );
nand NAND2_18208 ( P2_R1209_U298 , P2_R1209_U225 , P2_R1209_U67 );
nand NAND2_18209 ( P2_R1209_U299 , P2_R1209_U297 , P2_R1209_U205 );
nand NAND2_18210 ( P2_R1209_U300 , P2_U3461 , P2_R1209_U54 );
nand NAND2_18211 ( P2_R1209_U301 , P2_REG1_REG_11_ , P2_R1209_U55 );
nand NAND2_18212 ( P2_R1209_U302 , P2_R1209_U301 , P2_R1209_U300 );
nand NAND2_18213 ( P2_R1209_U303 , P2_R1209_U226 , P2_R1209_U88 );
nand NAND2_18214 ( P2_R1209_U304 , P2_R1209_U162 , P2_R1209_U302 );
nand NAND2_18215 ( P2_R1209_U305 , P2_U3458 , P2_R1209_U50 );
nand NAND2_18216 ( P2_R1209_U306 , P2_REG1_REG_10_ , P2_R1209_U51 );
nand NAND2_18217 ( P2_R1209_U307 , P2_U3425 , P2_R1209_U27 );
nand NAND2_18218 ( P2_R1209_U308 , P2_REG1_REG_0_ , P2_R1209_U28 );
and AND2_18219 ( P2_R1170_U4 , P2_R1170_U95 , P2_R1170_U94 );
and AND2_18220 ( P2_R1170_U5 , P2_R1170_U96 , P2_R1170_U97 );
and AND2_18221 ( P2_R1170_U6 , P2_R1170_U113 , P2_R1170_U112 );
and AND2_18222 ( P2_R1170_U7 , P2_R1170_U155 , P2_R1170_U154 );
and AND2_18223 ( P2_R1170_U8 , P2_R1170_U164 , P2_R1170_U163 );
and AND2_18224 ( P2_R1170_U9 , P2_R1170_U182 , P2_R1170_U181 );
and AND2_18225 ( P2_R1170_U10 , P2_R1170_U218 , P2_R1170_U215 );
and AND2_18226 ( P2_R1170_U11 , P2_R1170_U211 , P2_R1170_U208 );
and AND2_18227 ( P2_R1170_U12 , P2_R1170_U202 , P2_R1170_U199 );
and AND2_18228 ( P2_R1170_U13 , P2_R1170_U196 , P2_R1170_U192 );
and AND2_18229 ( P2_R1170_U14 , P2_R1170_U151 , P2_R1170_U148 );
and AND2_18230 ( P2_R1170_U15 , P2_R1170_U143 , P2_R1170_U140 );
and AND2_18231 ( P2_R1170_U16 , P2_R1170_U129 , P2_R1170_U126 );
not NOT1_18232 ( P2_R1170_U17 , P2_REG2_REG_6_ );
not NOT1_18233 ( P2_R1170_U18 , P2_U3446 );
not NOT1_18234 ( P2_R1170_U19 , P2_U3449 );
nand NAND2_18235 ( P2_R1170_U20 , P2_U3446 , P2_REG2_REG_6_ );
not NOT1_18236 ( P2_R1170_U21 , P2_REG2_REG_7_ );
not NOT1_18237 ( P2_R1170_U22 , P2_REG2_REG_4_ );
not NOT1_18238 ( P2_R1170_U23 , P2_U3440 );
not NOT1_18239 ( P2_R1170_U24 , P2_U3443 );
not NOT1_18240 ( P2_R1170_U25 , P2_REG2_REG_2_ );
not NOT1_18241 ( P2_R1170_U26 , P2_U3434 );
not NOT1_18242 ( P2_R1170_U27 , P2_REG2_REG_0_ );
not NOT1_18243 ( P2_R1170_U28 , P2_U3425 );
nand NAND2_18244 ( P2_R1170_U29 , P2_U3425 , P2_REG2_REG_0_ );
not NOT1_18245 ( P2_R1170_U30 , P2_REG2_REG_3_ );
not NOT1_18246 ( P2_R1170_U31 , P2_U3437 );
nand NAND2_18247 ( P2_R1170_U32 , P2_U3440 , P2_REG2_REG_4_ );
not NOT1_18248 ( P2_R1170_U33 , P2_REG2_REG_5_ );
not NOT1_18249 ( P2_R1170_U34 , P2_REG2_REG_8_ );
not NOT1_18250 ( P2_R1170_U35 , P2_U3452 );
not NOT1_18251 ( P2_R1170_U36 , P2_U3455 );
not NOT1_18252 ( P2_R1170_U37 , P2_REG2_REG_9_ );
nand NAND2_18253 ( P2_R1170_U38 , P2_R1170_U49 , P2_R1170_U121 );
nand NAND3_18254 ( P2_R1170_U39 , P2_R1170_U110 , P2_R1170_U108 , P2_R1170_U109 );
nand NAND2_18255 ( P2_R1170_U40 , P2_R1170_U98 , P2_R1170_U99 );
nand NAND2_18256 ( P2_R1170_U41 , P2_REG2_REG_1_ , P2_U3431 );
nand NAND3_18257 ( P2_R1170_U42 , P2_R1170_U136 , P2_R1170_U134 , P2_R1170_U135 );
nand NAND2_18258 ( P2_R1170_U43 , P2_R1170_U132 , P2_R1170_U131 );
not NOT1_18259 ( P2_R1170_U44 , P2_REG2_REG_16_ );
not NOT1_18260 ( P2_R1170_U45 , P2_U3476 );
not NOT1_18261 ( P2_R1170_U46 , P2_U3479 );
nand NAND2_18262 ( P2_R1170_U47 , P2_U3476 , P2_REG2_REG_16_ );
not NOT1_18263 ( P2_R1170_U48 , P2_REG2_REG_17_ );
nand NAND2_18264 ( P2_R1170_U49 , P2_U3452 , P2_REG2_REG_8_ );
not NOT1_18265 ( P2_R1170_U50 , P2_REG2_REG_10_ );
not NOT1_18266 ( P2_R1170_U51 , P2_U3458 );
not NOT1_18267 ( P2_R1170_U52 , P2_REG2_REG_12_ );
not NOT1_18268 ( P2_R1170_U53 , P2_U3464 );
not NOT1_18269 ( P2_R1170_U54 , P2_REG2_REG_11_ );
not NOT1_18270 ( P2_R1170_U55 , P2_U3461 );
nand NAND2_18271 ( P2_R1170_U56 , P2_U3461 , P2_REG2_REG_11_ );
not NOT1_18272 ( P2_R1170_U57 , P2_REG2_REG_13_ );
not NOT1_18273 ( P2_R1170_U58 , P2_U3467 );
not NOT1_18274 ( P2_R1170_U59 , P2_REG2_REG_14_ );
not NOT1_18275 ( P2_R1170_U60 , P2_U3470 );
not NOT1_18276 ( P2_R1170_U61 , P2_REG2_REG_15_ );
not NOT1_18277 ( P2_R1170_U62 , P2_U3473 );
not NOT1_18278 ( P2_R1170_U63 , P2_REG2_REG_18_ );
not NOT1_18279 ( P2_R1170_U64 , P2_U3482 );
nand NAND3_18280 ( P2_R1170_U65 , P2_R1170_U186 , P2_R1170_U185 , P2_R1170_U187 );
nand NAND2_18281 ( P2_R1170_U66 , P2_R1170_U179 , P2_R1170_U178 );
nand NAND2_18282 ( P2_R1170_U67 , P2_R1170_U56 , P2_R1170_U204 );
nand NAND2_18283 ( P2_R1170_U68 , P2_R1170_U259 , P2_R1170_U258 );
nand NAND2_18284 ( P2_R1170_U69 , P2_R1170_U308 , P2_R1170_U307 );
nand NAND2_18285 ( P2_R1170_U70 , P2_R1170_U231 , P2_R1170_U230 );
nand NAND2_18286 ( P2_R1170_U71 , P2_R1170_U236 , P2_R1170_U235 );
nand NAND2_18287 ( P2_R1170_U72 , P2_R1170_U243 , P2_R1170_U242 );
nand NAND2_18288 ( P2_R1170_U73 , P2_R1170_U250 , P2_R1170_U249 );
nand NAND2_18289 ( P2_R1170_U74 , P2_R1170_U255 , P2_R1170_U254 );
nand NAND2_18290 ( P2_R1170_U75 , P2_R1170_U271 , P2_R1170_U270 );
nand NAND2_18291 ( P2_R1170_U76 , P2_R1170_U278 , P2_R1170_U277 );
nand NAND2_18292 ( P2_R1170_U77 , P2_R1170_U285 , P2_R1170_U284 );
nand NAND2_18293 ( P2_R1170_U78 , P2_R1170_U292 , P2_R1170_U291 );
nand NAND2_18294 ( P2_R1170_U79 , P2_R1170_U299 , P2_R1170_U298 );
nand NAND2_18295 ( P2_R1170_U80 , P2_R1170_U304 , P2_R1170_U303 );
nand NAND3_18296 ( P2_R1170_U81 , P2_R1170_U117 , P2_R1170_U116 , P2_R1170_U118 );
nand NAND2_18297 ( P2_R1170_U82 , P2_R1170_U133 , P2_R1170_U145 );
nand NAND2_18298 ( P2_R1170_U83 , P2_R1170_U41 , P2_R1170_U152 );
not NOT1_18299 ( P2_R1170_U84 , P2_U3424 );
not NOT1_18300 ( P2_R1170_U85 , P2_REG2_REG_19_ );
nand NAND2_18301 ( P2_R1170_U86 , P2_R1170_U175 , P2_R1170_U174 );
nand NAND2_18302 ( P2_R1170_U87 , P2_R1170_U171 , P2_R1170_U170 );
nand NAND2_18303 ( P2_R1170_U88 , P2_R1170_U161 , P2_R1170_U160 );
not NOT1_18304 ( P2_R1170_U89 , P2_R1170_U32 );
nand NAND2_18305 ( P2_R1170_U90 , P2_REG2_REG_9_ , P2_U3455 );
nand NAND2_18306 ( P2_R1170_U91 , P2_U3464 , P2_REG2_REG_12_ );
not NOT1_18307 ( P2_R1170_U92 , P2_R1170_U56 );
not NOT1_18308 ( P2_R1170_U93 , P2_R1170_U49 );
or OR2_18309 ( P2_R1170_U94 , P2_U3443 , P2_REG2_REG_5_ );
or OR2_18310 ( P2_R1170_U95 , P2_U3440 , P2_REG2_REG_4_ );
or OR2_18311 ( P2_R1170_U96 , P2_REG2_REG_3_ , P2_U3437 );
or OR2_18312 ( P2_R1170_U97 , P2_REG2_REG_2_ , P2_U3434 );
not NOT1_18313 ( P2_R1170_U98 , P2_R1170_U29 );
or OR2_18314 ( P2_R1170_U99 , P2_REG2_REG_1_ , P2_U3431 );
not NOT1_18315 ( P2_R1170_U100 , P2_R1170_U40 );
not NOT1_18316 ( P2_R1170_U101 , P2_R1170_U41 );
nand NAND2_18317 ( P2_R1170_U102 , P2_R1170_U40 , P2_R1170_U41 );
nand NAND3_18318 ( P2_R1170_U103 , P2_REG2_REG_2_ , P2_U3434 , P2_R1170_U96 );
nand NAND2_18319 ( P2_R1170_U104 , P2_R1170_U5 , P2_R1170_U102 );
nand NAND2_18320 ( P2_R1170_U105 , P2_U3437 , P2_REG2_REG_3_ );
nand NAND3_18321 ( P2_R1170_U106 , P2_R1170_U105 , P2_R1170_U103 , P2_R1170_U104 );
nand NAND2_18322 ( P2_R1170_U107 , P2_R1170_U33 , P2_R1170_U32 );
nand NAND2_18323 ( P2_R1170_U108 , P2_U3443 , P2_R1170_U107 );
nand NAND2_18324 ( P2_R1170_U109 , P2_R1170_U4 , P2_R1170_U106 );
nand NAND2_18325 ( P2_R1170_U110 , P2_REG2_REG_5_ , P2_R1170_U89 );
not NOT1_18326 ( P2_R1170_U111 , P2_R1170_U39 );
or OR2_18327 ( P2_R1170_U112 , P2_U3449 , P2_REG2_REG_7_ );
or OR2_18328 ( P2_R1170_U113 , P2_U3446 , P2_REG2_REG_6_ );
not NOT1_18329 ( P2_R1170_U114 , P2_R1170_U20 );
nand NAND2_18330 ( P2_R1170_U115 , P2_R1170_U21 , P2_R1170_U20 );
nand NAND2_18331 ( P2_R1170_U116 , P2_U3449 , P2_R1170_U115 );
nand NAND2_18332 ( P2_R1170_U117 , P2_REG2_REG_7_ , P2_R1170_U114 );
nand NAND2_18333 ( P2_R1170_U118 , P2_R1170_U6 , P2_R1170_U39 );
not NOT1_18334 ( P2_R1170_U119 , P2_R1170_U81 );
or OR2_18335 ( P2_R1170_U120 , P2_REG2_REG_8_ , P2_U3452 );
nand NAND2_18336 ( P2_R1170_U121 , P2_R1170_U120 , P2_R1170_U81 );
not NOT1_18337 ( P2_R1170_U122 , P2_R1170_U38 );
or OR2_18338 ( P2_R1170_U123 , P2_U3455 , P2_REG2_REG_9_ );
or OR2_18339 ( P2_R1170_U124 , P2_REG2_REG_6_ , P2_U3446 );
nand NAND2_18340 ( P2_R1170_U125 , P2_R1170_U124 , P2_R1170_U39 );
nand NAND4_18341 ( P2_R1170_U126 , P2_R1170_U238 , P2_R1170_U237 , P2_R1170_U20 , P2_R1170_U125 );
nand NAND2_18342 ( P2_R1170_U127 , P2_R1170_U111 , P2_R1170_U20 );
nand NAND2_18343 ( P2_R1170_U128 , P2_REG2_REG_7_ , P2_U3449 );
nand NAND3_18344 ( P2_R1170_U129 , P2_R1170_U128 , P2_R1170_U6 , P2_R1170_U127 );
or OR2_18345 ( P2_R1170_U130 , P2_U3446 , P2_REG2_REG_6_ );
nand NAND2_18346 ( P2_R1170_U131 , P2_R1170_U101 , P2_R1170_U97 );
nand NAND2_18347 ( P2_R1170_U132 , P2_U3434 , P2_REG2_REG_2_ );
not NOT1_18348 ( P2_R1170_U133 , P2_R1170_U43 );
nand NAND2_18349 ( P2_R1170_U134 , P2_R1170_U100 , P2_R1170_U5 );
nand NAND2_18350 ( P2_R1170_U135 , P2_R1170_U43 , P2_R1170_U96 );
nand NAND2_18351 ( P2_R1170_U136 , P2_U3437 , P2_REG2_REG_3_ );
not NOT1_18352 ( P2_R1170_U137 , P2_R1170_U42 );
or OR2_18353 ( P2_R1170_U138 , P2_REG2_REG_4_ , P2_U3440 );
nand NAND2_18354 ( P2_R1170_U139 , P2_R1170_U138 , P2_R1170_U42 );
nand NAND4_18355 ( P2_R1170_U140 , P2_R1170_U245 , P2_R1170_U244 , P2_R1170_U32 , P2_R1170_U139 );
nand NAND2_18356 ( P2_R1170_U141 , P2_R1170_U137 , P2_R1170_U32 );
nand NAND2_18357 ( P2_R1170_U142 , P2_REG2_REG_5_ , P2_U3443 );
nand NAND3_18358 ( P2_R1170_U143 , P2_R1170_U142 , P2_R1170_U4 , P2_R1170_U141 );
or OR2_18359 ( P2_R1170_U144 , P2_U3440 , P2_REG2_REG_4_ );
nand NAND2_18360 ( P2_R1170_U145 , P2_R1170_U100 , P2_R1170_U97 );
not NOT1_18361 ( P2_R1170_U146 , P2_R1170_U82 );
nand NAND2_18362 ( P2_R1170_U147 , P2_U3437 , P2_REG2_REG_3_ );
nand NAND4_18363 ( P2_R1170_U148 , P2_R1170_U257 , P2_R1170_U256 , P2_R1170_U41 , P2_R1170_U40 );
nand NAND2_18364 ( P2_R1170_U149 , P2_R1170_U41 , P2_R1170_U40 );
nand NAND2_18365 ( P2_R1170_U150 , P2_U3434 , P2_REG2_REG_2_ );
nand NAND3_18366 ( P2_R1170_U151 , P2_R1170_U150 , P2_R1170_U97 , P2_R1170_U149 );
or OR2_18367 ( P2_R1170_U152 , P2_REG2_REG_1_ , P2_U3431 );
not NOT1_18368 ( P2_R1170_U153 , P2_R1170_U83 );
or OR2_18369 ( P2_R1170_U154 , P2_U3455 , P2_REG2_REG_9_ );
or OR2_18370 ( P2_R1170_U155 , P2_U3458 , P2_REG2_REG_10_ );
nand NAND2_18371 ( P2_R1170_U156 , P2_R1170_U93 , P2_R1170_U7 );
nand NAND2_18372 ( P2_R1170_U157 , P2_U3458 , P2_REG2_REG_10_ );
nand NAND3_18373 ( P2_R1170_U158 , P2_R1170_U157 , P2_R1170_U90 , P2_R1170_U156 );
or OR2_18374 ( P2_R1170_U159 , P2_REG2_REG_10_ , P2_U3458 );
nand NAND3_18375 ( P2_R1170_U160 , P2_R1170_U120 , P2_R1170_U7 , P2_R1170_U81 );
nand NAND2_18376 ( P2_R1170_U161 , P2_R1170_U159 , P2_R1170_U158 );
not NOT1_18377 ( P2_R1170_U162 , P2_R1170_U88 );
or OR2_18378 ( P2_R1170_U163 , P2_U3467 , P2_REG2_REG_13_ );
or OR2_18379 ( P2_R1170_U164 , P2_U3464 , P2_REG2_REG_12_ );
nand NAND2_18380 ( P2_R1170_U165 , P2_R1170_U92 , P2_R1170_U8 );
nand NAND2_18381 ( P2_R1170_U166 , P2_U3467 , P2_REG2_REG_13_ );
nand NAND3_18382 ( P2_R1170_U167 , P2_R1170_U166 , P2_R1170_U91 , P2_R1170_U165 );
or OR2_18383 ( P2_R1170_U168 , P2_REG2_REG_11_ , P2_U3461 );
or OR2_18384 ( P2_R1170_U169 , P2_REG2_REG_13_ , P2_U3467 );
nand NAND3_18385 ( P2_R1170_U170 , P2_R1170_U168 , P2_R1170_U8 , P2_R1170_U88 );
nand NAND2_18386 ( P2_R1170_U171 , P2_R1170_U169 , P2_R1170_U167 );
not NOT1_18387 ( P2_R1170_U172 , P2_R1170_U87 );
or OR2_18388 ( P2_R1170_U173 , P2_REG2_REG_14_ , P2_U3470 );
nand NAND2_18389 ( P2_R1170_U174 , P2_R1170_U173 , P2_R1170_U87 );
nand NAND2_18390 ( P2_R1170_U175 , P2_U3470 , P2_REG2_REG_14_ );
not NOT1_18391 ( P2_R1170_U176 , P2_R1170_U86 );
or OR2_18392 ( P2_R1170_U177 , P2_REG2_REG_15_ , P2_U3473 );
nand NAND2_18393 ( P2_R1170_U178 , P2_R1170_U177 , P2_R1170_U86 );
nand NAND2_18394 ( P2_R1170_U179 , P2_U3473 , P2_REG2_REG_15_ );
not NOT1_18395 ( P2_R1170_U180 , P2_R1170_U66 );
or OR2_18396 ( P2_R1170_U181 , P2_U3479 , P2_REG2_REG_17_ );
or OR2_18397 ( P2_R1170_U182 , P2_U3476 , P2_REG2_REG_16_ );
not NOT1_18398 ( P2_R1170_U183 , P2_R1170_U47 );
nand NAND2_18399 ( P2_R1170_U184 , P2_R1170_U48 , P2_R1170_U47 );
nand NAND2_18400 ( P2_R1170_U185 , P2_U3479 , P2_R1170_U184 );
nand NAND2_18401 ( P2_R1170_U186 , P2_REG2_REG_17_ , P2_R1170_U183 );
nand NAND2_18402 ( P2_R1170_U187 , P2_R1170_U9 , P2_R1170_U66 );
not NOT1_18403 ( P2_R1170_U188 , P2_R1170_U65 );
or OR2_18404 ( P2_R1170_U189 , P2_REG2_REG_18_ , P2_U3482 );
nand NAND2_18405 ( P2_R1170_U190 , P2_R1170_U189 , P2_R1170_U65 );
nand NAND2_18406 ( P2_R1170_U191 , P2_U3482 , P2_REG2_REG_18_ );
nand NAND4_18407 ( P2_R1170_U192 , P2_R1170_U261 , P2_R1170_U260 , P2_R1170_U191 , P2_R1170_U190 );
nand NAND2_18408 ( P2_R1170_U193 , P2_U3482 , P2_REG2_REG_18_ );
nand NAND2_18409 ( P2_R1170_U194 , P2_R1170_U188 , P2_R1170_U193 );
or OR2_18410 ( P2_R1170_U195 , P2_U3482 , P2_REG2_REG_18_ );
nand NAND3_18411 ( P2_R1170_U196 , P2_R1170_U195 , P2_R1170_U264 , P2_R1170_U194 );
or OR2_18412 ( P2_R1170_U197 , P2_REG2_REG_16_ , P2_U3476 );
nand NAND2_18413 ( P2_R1170_U198 , P2_R1170_U197 , P2_R1170_U66 );
nand NAND4_18414 ( P2_R1170_U199 , P2_R1170_U273 , P2_R1170_U272 , P2_R1170_U47 , P2_R1170_U198 );
nand NAND2_18415 ( P2_R1170_U200 , P2_R1170_U180 , P2_R1170_U47 );
nand NAND2_18416 ( P2_R1170_U201 , P2_REG2_REG_17_ , P2_U3479 );
nand NAND3_18417 ( P2_R1170_U202 , P2_R1170_U201 , P2_R1170_U9 , P2_R1170_U200 );
or OR2_18418 ( P2_R1170_U203 , P2_U3476 , P2_REG2_REG_16_ );
nand NAND2_18419 ( P2_R1170_U204 , P2_R1170_U168 , P2_R1170_U88 );
not NOT1_18420 ( P2_R1170_U205 , P2_R1170_U67 );
or OR2_18421 ( P2_R1170_U206 , P2_REG2_REG_12_ , P2_U3464 );
nand NAND2_18422 ( P2_R1170_U207 , P2_R1170_U206 , P2_R1170_U67 );
nand NAND4_18423 ( P2_R1170_U208 , P2_R1170_U294 , P2_R1170_U293 , P2_R1170_U91 , P2_R1170_U207 );
nand NAND2_18424 ( P2_R1170_U209 , P2_R1170_U205 , P2_R1170_U91 );
nand NAND2_18425 ( P2_R1170_U210 , P2_U3467 , P2_REG2_REG_13_ );
nand NAND3_18426 ( P2_R1170_U211 , P2_R1170_U210 , P2_R1170_U8 , P2_R1170_U209 );
or OR2_18427 ( P2_R1170_U212 , P2_U3464 , P2_REG2_REG_12_ );
or OR2_18428 ( P2_R1170_U213 , P2_REG2_REG_9_ , P2_U3455 );
nand NAND2_18429 ( P2_R1170_U214 , P2_R1170_U213 , P2_R1170_U38 );
nand NAND4_18430 ( P2_R1170_U215 , P2_R1170_U306 , P2_R1170_U305 , P2_R1170_U90 , P2_R1170_U214 );
nand NAND2_18431 ( P2_R1170_U216 , P2_R1170_U122 , P2_R1170_U90 );
nand NAND2_18432 ( P2_R1170_U217 , P2_U3458 , P2_REG2_REG_10_ );
nand NAND3_18433 ( P2_R1170_U218 , P2_R1170_U217 , P2_R1170_U7 , P2_R1170_U216 );
nand NAND2_18434 ( P2_R1170_U219 , P2_R1170_U123 , P2_R1170_U90 );
nand NAND2_18435 ( P2_R1170_U220 , P2_R1170_U120 , P2_R1170_U49 );
nand NAND2_18436 ( P2_R1170_U221 , P2_R1170_U130 , P2_R1170_U20 );
nand NAND2_18437 ( P2_R1170_U222 , P2_R1170_U144 , P2_R1170_U32 );
nand NAND2_18438 ( P2_R1170_U223 , P2_R1170_U147 , P2_R1170_U96 );
nand NAND2_18439 ( P2_R1170_U224 , P2_R1170_U203 , P2_R1170_U47 );
nand NAND2_18440 ( P2_R1170_U225 , P2_R1170_U212 , P2_R1170_U91 );
nand NAND2_18441 ( P2_R1170_U226 , P2_R1170_U168 , P2_R1170_U56 );
nand NAND2_18442 ( P2_R1170_U227 , P2_U3455 , P2_R1170_U37 );
nand NAND2_18443 ( P2_R1170_U228 , P2_REG2_REG_9_ , P2_R1170_U36 );
nand NAND2_18444 ( P2_R1170_U229 , P2_R1170_U228 , P2_R1170_U227 );
nand NAND2_18445 ( P2_R1170_U230 , P2_R1170_U219 , P2_R1170_U38 );
nand NAND2_18446 ( P2_R1170_U231 , P2_R1170_U229 , P2_R1170_U122 );
nand NAND2_18447 ( P2_R1170_U232 , P2_U3452 , P2_R1170_U34 );
nand NAND2_18448 ( P2_R1170_U233 , P2_REG2_REG_8_ , P2_R1170_U35 );
nand NAND2_18449 ( P2_R1170_U234 , P2_R1170_U233 , P2_R1170_U232 );
nand NAND2_18450 ( P2_R1170_U235 , P2_R1170_U220 , P2_R1170_U81 );
nand NAND2_18451 ( P2_R1170_U236 , P2_R1170_U119 , P2_R1170_U234 );
nand NAND2_18452 ( P2_R1170_U237 , P2_U3449 , P2_R1170_U21 );
nand NAND2_18453 ( P2_R1170_U238 , P2_REG2_REG_7_ , P2_R1170_U19 );
nand NAND2_18454 ( P2_R1170_U239 , P2_U3446 , P2_R1170_U17 );
nand NAND2_18455 ( P2_R1170_U240 , P2_REG2_REG_6_ , P2_R1170_U18 );
nand NAND2_18456 ( P2_R1170_U241 , P2_R1170_U240 , P2_R1170_U239 );
nand NAND2_18457 ( P2_R1170_U242 , P2_R1170_U221 , P2_R1170_U39 );
nand NAND2_18458 ( P2_R1170_U243 , P2_R1170_U241 , P2_R1170_U111 );
nand NAND2_18459 ( P2_R1170_U244 , P2_U3443 , P2_R1170_U33 );
nand NAND2_18460 ( P2_R1170_U245 , P2_REG2_REG_5_ , P2_R1170_U24 );
nand NAND2_18461 ( P2_R1170_U246 , P2_U3440 , P2_R1170_U22 );
nand NAND2_18462 ( P2_R1170_U247 , P2_REG2_REG_4_ , P2_R1170_U23 );
nand NAND2_18463 ( P2_R1170_U248 , P2_R1170_U247 , P2_R1170_U246 );
nand NAND2_18464 ( P2_R1170_U249 , P2_R1170_U222 , P2_R1170_U42 );
nand NAND2_18465 ( P2_R1170_U250 , P2_R1170_U248 , P2_R1170_U137 );
nand NAND2_18466 ( P2_R1170_U251 , P2_U3437 , P2_R1170_U30 );
nand NAND2_18467 ( P2_R1170_U252 , P2_REG2_REG_3_ , P2_R1170_U31 );
nand NAND2_18468 ( P2_R1170_U253 , P2_R1170_U252 , P2_R1170_U251 );
nand NAND2_18469 ( P2_R1170_U254 , P2_R1170_U223 , P2_R1170_U82 );
nand NAND2_18470 ( P2_R1170_U255 , P2_R1170_U146 , P2_R1170_U253 );
nand NAND2_18471 ( P2_R1170_U256 , P2_U3434 , P2_R1170_U25 );
nand NAND2_18472 ( P2_R1170_U257 , P2_REG2_REG_2_ , P2_R1170_U26 );
nand NAND2_18473 ( P2_R1170_U258 , P2_R1170_U98 , P2_R1170_U83 );
nand NAND2_18474 ( P2_R1170_U259 , P2_R1170_U153 , P2_R1170_U29 );
nand NAND2_18475 ( P2_R1170_U260 , P2_U3424 , P2_R1170_U85 );
nand NAND2_18476 ( P2_R1170_U261 , P2_REG2_REG_19_ , P2_R1170_U84 );
nand NAND2_18477 ( P2_R1170_U262 , P2_U3424 , P2_R1170_U85 );
nand NAND2_18478 ( P2_R1170_U263 , P2_REG2_REG_19_ , P2_R1170_U84 );
nand NAND2_18479 ( P2_R1170_U264 , P2_R1170_U263 , P2_R1170_U262 );
nand NAND2_18480 ( P2_R1170_U265 , P2_U3482 , P2_R1170_U63 );
nand NAND2_18481 ( P2_R1170_U266 , P2_REG2_REG_18_ , P2_R1170_U64 );
nand NAND2_18482 ( P2_R1170_U267 , P2_U3482 , P2_R1170_U63 );
nand NAND2_18483 ( P2_R1170_U268 , P2_REG2_REG_18_ , P2_R1170_U64 );
nand NAND2_18484 ( P2_R1170_U269 , P2_R1170_U268 , P2_R1170_U267 );
nand NAND3_18485 ( P2_R1170_U270 , P2_R1170_U266 , P2_R1170_U265 , P2_R1170_U65 );
nand NAND2_18486 ( P2_R1170_U271 , P2_R1170_U269 , P2_R1170_U188 );
nand NAND2_18487 ( P2_R1170_U272 , P2_U3479 , P2_R1170_U48 );
nand NAND2_18488 ( P2_R1170_U273 , P2_REG2_REG_17_ , P2_R1170_U46 );
nand NAND2_18489 ( P2_R1170_U274 , P2_U3476 , P2_R1170_U44 );
nand NAND2_18490 ( P2_R1170_U275 , P2_REG2_REG_16_ , P2_R1170_U45 );
nand NAND2_18491 ( P2_R1170_U276 , P2_R1170_U275 , P2_R1170_U274 );
nand NAND2_18492 ( P2_R1170_U277 , P2_R1170_U224 , P2_R1170_U66 );
nand NAND2_18493 ( P2_R1170_U278 , P2_R1170_U276 , P2_R1170_U180 );
nand NAND2_18494 ( P2_R1170_U279 , P2_U3473 , P2_R1170_U61 );
nand NAND2_18495 ( P2_R1170_U280 , P2_REG2_REG_15_ , P2_R1170_U62 );
nand NAND2_18496 ( P2_R1170_U281 , P2_U3473 , P2_R1170_U61 );
nand NAND2_18497 ( P2_R1170_U282 , P2_REG2_REG_15_ , P2_R1170_U62 );
nand NAND2_18498 ( P2_R1170_U283 , P2_R1170_U282 , P2_R1170_U281 );
nand NAND3_18499 ( P2_R1170_U284 , P2_R1170_U280 , P2_R1170_U279 , P2_R1170_U86 );
nand NAND2_18500 ( P2_R1170_U285 , P2_R1170_U176 , P2_R1170_U283 );
nand NAND2_18501 ( P2_R1170_U286 , P2_U3470 , P2_R1170_U59 );
nand NAND2_18502 ( P2_R1170_U287 , P2_REG2_REG_14_ , P2_R1170_U60 );
nand NAND2_18503 ( P2_R1170_U288 , P2_U3470 , P2_R1170_U59 );
nand NAND2_18504 ( P2_R1170_U289 , P2_REG2_REG_14_ , P2_R1170_U60 );
nand NAND2_18505 ( P2_R1170_U290 , P2_R1170_U289 , P2_R1170_U288 );
nand NAND3_18506 ( P2_R1170_U291 , P2_R1170_U287 , P2_R1170_U286 , P2_R1170_U87 );
nand NAND2_18507 ( P2_R1170_U292 , P2_R1170_U172 , P2_R1170_U290 );
nand NAND2_18508 ( P2_R1170_U293 , P2_U3467 , P2_R1170_U57 );
nand NAND2_18509 ( P2_R1170_U294 , P2_REG2_REG_13_ , P2_R1170_U58 );
nand NAND2_18510 ( P2_R1170_U295 , P2_U3464 , P2_R1170_U52 );
nand NAND2_18511 ( P2_R1170_U296 , P2_REG2_REG_12_ , P2_R1170_U53 );
nand NAND2_18512 ( P2_R1170_U297 , P2_R1170_U296 , P2_R1170_U295 );
nand NAND2_18513 ( P2_R1170_U298 , P2_R1170_U225 , P2_R1170_U67 );
nand NAND2_18514 ( P2_R1170_U299 , P2_R1170_U297 , P2_R1170_U205 );
nand NAND2_18515 ( P2_R1170_U300 , P2_U3461 , P2_R1170_U54 );
nand NAND2_18516 ( P2_R1170_U301 , P2_REG2_REG_11_ , P2_R1170_U55 );
nand NAND2_18517 ( P2_R1170_U302 , P2_R1170_U301 , P2_R1170_U300 );
nand NAND2_18518 ( P2_R1170_U303 , P2_R1170_U226 , P2_R1170_U88 );
nand NAND2_18519 ( P2_R1170_U304 , P2_R1170_U162 , P2_R1170_U302 );
nand NAND2_18520 ( P2_R1170_U305 , P2_U3458 , P2_R1170_U50 );
nand NAND2_18521 ( P2_R1170_U306 , P2_REG2_REG_10_ , P2_R1170_U51 );
nand NAND2_18522 ( P2_R1170_U307 , P2_U3425 , P2_R1170_U27 );
nand NAND2_18523 ( P2_R1170_U308 , P2_REG2_REG_0_ , P2_R1170_U28 );
and AND2_18524 ( P2_R1275_U6 , P2_R1275_U135 , P2_R1275_U35 );
and AND2_18525 ( P2_R1275_U7 , P2_R1275_U133 , P2_R1275_U36 );
and AND2_18526 ( P2_R1275_U8 , P2_R1275_U132 , P2_R1275_U37 );
and AND2_18527 ( P2_R1275_U9 , P2_R1275_U131 , P2_R1275_U38 );
and AND2_18528 ( P2_R1275_U10 , P2_R1275_U129 , P2_R1275_U39 );
and AND2_18529 ( P2_R1275_U11 , P2_R1275_U128 , P2_R1275_U40 );
and AND2_18530 ( P2_R1275_U12 , P2_R1275_U127 , P2_R1275_U41 );
and AND2_18531 ( P2_R1275_U13 , P2_R1275_U125 , P2_R1275_U42 );
and AND2_18532 ( P2_R1275_U14 , P2_R1275_U123 , P2_R1275_U43 );
and AND2_18533 ( P2_R1275_U15 , P2_R1275_U121 , P2_R1275_U44 );
and AND2_18534 ( P2_R1275_U16 , P2_R1275_U119 , P2_R1275_U45 );
and AND2_18535 ( P2_R1275_U17 , P2_R1275_U117 , P2_R1275_U46 );
and AND2_18536 ( P2_R1275_U18 , P2_R1275_U115 , P2_R1275_U25 );
and AND2_18537 ( P2_R1275_U19 , P2_R1275_U113 , P2_R1275_U67 );
and AND2_18538 ( P2_R1275_U20 , P2_R1275_U98 , P2_R1275_U26 );
and AND2_18539 ( P2_R1275_U21 , P2_R1275_U97 , P2_R1275_U27 );
and AND2_18540 ( P2_R1275_U22 , P2_R1275_U96 , P2_R1275_U28 );
and AND2_18541 ( P2_R1275_U23 , P2_R1275_U94 , P2_R1275_U29 );
and AND2_18542 ( P2_R1275_U24 , P2_R1275_U93 , P2_R1275_U30 );
or OR3_18543 ( P2_R1275_U25 , P2_U3432 , P2_U3427 , P2_U3435 );
nand NAND2_18544 ( P2_R1275_U26 , P2_R1275_U87 , P2_R1275_U34 );
nand NAND2_18545 ( P2_R1275_U27 , P2_R1275_U88 , P2_R1275_U33 );
nand NAND2_18546 ( P2_R1275_U28 , P2_R1275_U56 , P2_R1275_U89 );
nand NAND2_18547 ( P2_R1275_U29 , P2_R1275_U90 , P2_R1275_U32 );
nand NAND2_18548 ( P2_R1275_U30 , P2_R1275_U91 , P2_R1275_U31 );
not NOT1_18549 ( P2_R1275_U31 , P2_U3453 );
not NOT1_18550 ( P2_R1275_U32 , P2_U3450 );
not NOT1_18551 ( P2_R1275_U33 , P2_U3441 );
not NOT1_18552 ( P2_R1275_U34 , P2_U3438 );
nand NAND2_18553 ( P2_R1275_U35 , P2_R1275_U57 , P2_R1275_U92 );
nand NAND2_18554 ( P2_R1275_U36 , P2_R1275_U99 , P2_R1275_U54 );
nand NAND2_18555 ( P2_R1275_U37 , P2_R1275_U100 , P2_R1275_U53 );
nand NAND2_18556 ( P2_R1275_U38 , P2_R1275_U58 , P2_R1275_U101 );
nand NAND2_18557 ( P2_R1275_U39 , P2_R1275_U102 , P2_R1275_U52 );
nand NAND2_18558 ( P2_R1275_U40 , P2_R1275_U103 , P2_R1275_U51 );
nand NAND2_18559 ( P2_R1275_U41 , P2_R1275_U59 , P2_R1275_U104 );
nand NAND2_18560 ( P2_R1275_U42 , P2_R1275_U60 , P2_R1275_U105 );
nand NAND2_18561 ( P2_R1275_U43 , P2_R1275_U61 , P2_R1275_U106 );
nand NAND3_18562 ( P2_R1275_U44 , P2_R1275_U107 , P2_R1275_U75 , P2_R1275_U50 );
nand NAND3_18563 ( P2_R1275_U45 , P2_R1275_U108 , P2_R1275_U73 , P2_R1275_U49 );
nand NAND3_18564 ( P2_R1275_U46 , P2_R1275_U109 , P2_R1275_U71 , P2_R1275_U48 );
not NOT1_18565 ( P2_R1275_U47 , P2_U3959 );
not NOT1_18566 ( P2_R1275_U48 , P2_U3949 );
not NOT1_18567 ( P2_R1275_U49 , P2_U3951 );
not NOT1_18568 ( P2_R1275_U50 , P2_U3953 );
not NOT1_18569 ( P2_R1275_U51 , P2_U3477 );
not NOT1_18570 ( P2_R1275_U52 , P2_U3474 );
not NOT1_18571 ( P2_R1275_U53 , P2_U3465 );
not NOT1_18572 ( P2_R1275_U54 , P2_U3462 );
nand NAND2_18573 ( P2_R1275_U55 , P2_R1275_U153 , P2_R1275_U152 );
nor nor_18574 ( P2_R1275_U56 , P2_U3444 , P2_U3447 );
nor nor_18575 ( P2_R1275_U57 , P2_U3459 , P2_U3456 );
nor nor_18576 ( P2_R1275_U58 , P2_U3468 , P2_U3471 );
nor nor_18577 ( P2_R1275_U59 , P2_U3480 , P2_U3483 );
nor nor_18578 ( P2_R1275_U60 , P2_U3485 , P2_U3957 );
nor nor_18579 ( P2_R1275_U61 , P2_U3956 , P2_U3955 );
not NOT1_18580 ( P2_R1275_U62 , P2_U3456 );
and AND2_18581 ( P2_R1275_U63 , P2_R1275_U137 , P2_R1275_U136 );
not NOT1_18582 ( P2_R1275_U64 , P2_U3444 );
and AND2_18583 ( P2_R1275_U65 , P2_R1275_U139 , P2_R1275_U138 );
not NOT1_18584 ( P2_R1275_U66 , P2_U3958 );
nand NAND3_18585 ( P2_R1275_U67 , P2_R1275_U110 , P2_R1275_U69 , P2_R1275_U47 );
and AND2_18586 ( P2_R1275_U68 , P2_R1275_U141 , P2_R1275_U140 );
not NOT1_18587 ( P2_R1275_U69 , P2_U3960 );
and AND2_18588 ( P2_R1275_U70 , P2_R1275_U143 , P2_R1275_U142 );
not NOT1_18589 ( P2_R1275_U71 , P2_U3950 );
and AND2_18590 ( P2_R1275_U72 , P2_R1275_U145 , P2_R1275_U144 );
not NOT1_18591 ( P2_R1275_U73 , P2_U3952 );
and AND2_18592 ( P2_R1275_U74 , P2_R1275_U147 , P2_R1275_U146 );
not NOT1_18593 ( P2_R1275_U75 , P2_U3954 );
and AND2_18594 ( P2_R1275_U76 , P2_R1275_U149 , P2_R1275_U148 );
not NOT1_18595 ( P2_R1275_U77 , P2_U3956 );
and AND2_18596 ( P2_R1275_U78 , P2_R1275_U151 , P2_R1275_U150 );
not NOT1_18597 ( P2_R1275_U79 , P2_U3432 );
not NOT1_18598 ( P2_R1275_U80 , P2_U3427 );
not NOT1_18599 ( P2_R1275_U81 , P2_U3485 );
and AND2_18600 ( P2_R1275_U82 , P2_R1275_U155 , P2_R1275_U154 );
not NOT1_18601 ( P2_R1275_U83 , P2_U3480 );
and AND2_18602 ( P2_R1275_U84 , P2_R1275_U157 , P2_R1275_U156 );
not NOT1_18603 ( P2_R1275_U85 , P2_U3468 );
and AND2_18604 ( P2_R1275_U86 , P2_R1275_U159 , P2_R1275_U158 );
not NOT1_18605 ( P2_R1275_U87 , P2_R1275_U25 );
not NOT1_18606 ( P2_R1275_U88 , P2_R1275_U26 );
not NOT1_18607 ( P2_R1275_U89 , P2_R1275_U27 );
not NOT1_18608 ( P2_R1275_U90 , P2_R1275_U28 );
not NOT1_18609 ( P2_R1275_U91 , P2_R1275_U29 );
not NOT1_18610 ( P2_R1275_U92 , P2_R1275_U30 );
nand NAND2_18611 ( P2_R1275_U93 , P2_U3453 , P2_R1275_U29 );
nand NAND2_18612 ( P2_R1275_U94 , P2_U3450 , P2_R1275_U28 );
nand NAND2_18613 ( P2_R1275_U95 , P2_R1275_U89 , P2_R1275_U64 );
nand NAND2_18614 ( P2_R1275_U96 , P2_U3447 , P2_R1275_U95 );
nand NAND2_18615 ( P2_R1275_U97 , P2_U3441 , P2_R1275_U26 );
nand NAND2_18616 ( P2_R1275_U98 , P2_U3438 , P2_R1275_U25 );
not NOT1_18617 ( P2_R1275_U99 , P2_R1275_U35 );
not NOT1_18618 ( P2_R1275_U100 , P2_R1275_U36 );
not NOT1_18619 ( P2_R1275_U101 , P2_R1275_U37 );
not NOT1_18620 ( P2_R1275_U102 , P2_R1275_U38 );
not NOT1_18621 ( P2_R1275_U103 , P2_R1275_U39 );
not NOT1_18622 ( P2_R1275_U104 , P2_R1275_U40 );
not NOT1_18623 ( P2_R1275_U105 , P2_R1275_U41 );
not NOT1_18624 ( P2_R1275_U106 , P2_R1275_U42 );
not NOT1_18625 ( P2_R1275_U107 , P2_R1275_U43 );
not NOT1_18626 ( P2_R1275_U108 , P2_R1275_U44 );
not NOT1_18627 ( P2_R1275_U109 , P2_R1275_U45 );
not NOT1_18628 ( P2_R1275_U110 , P2_R1275_U46 );
not NOT1_18629 ( P2_R1275_U111 , P2_R1275_U67 );
nand NAND2_18630 ( P2_R1275_U112 , P2_R1275_U110 , P2_R1275_U69 );
nand NAND2_18631 ( P2_R1275_U113 , P2_U3959 , P2_R1275_U112 );
or OR2_18632 ( P2_R1275_U114 , P2_U3432 , P2_U3427 );
nand NAND2_18633 ( P2_R1275_U115 , P2_U3435 , P2_R1275_U114 );
nand NAND2_18634 ( P2_R1275_U116 , P2_R1275_U109 , P2_R1275_U71 );
nand NAND2_18635 ( P2_R1275_U117 , P2_U3949 , P2_R1275_U116 );
nand NAND2_18636 ( P2_R1275_U118 , P2_R1275_U108 , P2_R1275_U73 );
nand NAND2_18637 ( P2_R1275_U119 , P2_U3951 , P2_R1275_U118 );
nand NAND2_18638 ( P2_R1275_U120 , P2_R1275_U107 , P2_R1275_U75 );
nand NAND2_18639 ( P2_R1275_U121 , P2_U3953 , P2_R1275_U120 );
nand NAND2_18640 ( P2_R1275_U122 , P2_R1275_U106 , P2_R1275_U77 );
nand NAND2_18641 ( P2_R1275_U123 , P2_U3955 , P2_R1275_U122 );
nand NAND2_18642 ( P2_R1275_U124 , P2_R1275_U105 , P2_R1275_U81 );
nand NAND2_18643 ( P2_R1275_U125 , P2_U3957 , P2_R1275_U124 );
nand NAND2_18644 ( P2_R1275_U126 , P2_R1275_U104 , P2_R1275_U83 );
nand NAND2_18645 ( P2_R1275_U127 , P2_U3483 , P2_R1275_U126 );
nand NAND2_18646 ( P2_R1275_U128 , P2_U3477 , P2_R1275_U39 );
nand NAND2_18647 ( P2_R1275_U129 , P2_U3474 , P2_R1275_U38 );
nand NAND2_18648 ( P2_R1275_U130 , P2_R1275_U101 , P2_R1275_U85 );
nand NAND2_18649 ( P2_R1275_U131 , P2_U3471 , P2_R1275_U130 );
nand NAND2_18650 ( P2_R1275_U132 , P2_U3465 , P2_R1275_U36 );
nand NAND2_18651 ( P2_R1275_U133 , P2_U3462 , P2_R1275_U35 );
nand NAND2_18652 ( P2_R1275_U134 , P2_R1275_U92 , P2_R1275_U62 );
nand NAND2_18653 ( P2_R1275_U135 , P2_U3459 , P2_R1275_U134 );
nand NAND2_18654 ( P2_R1275_U136 , P2_U3456 , P2_R1275_U30 );
nand NAND2_18655 ( P2_R1275_U137 , P2_R1275_U92 , P2_R1275_U62 );
nand NAND2_18656 ( P2_R1275_U138 , P2_U3444 , P2_R1275_U27 );
nand NAND2_18657 ( P2_R1275_U139 , P2_R1275_U89 , P2_R1275_U64 );
nand NAND2_18658 ( P2_R1275_U140 , P2_U3958 , P2_R1275_U67 );
nand NAND2_18659 ( P2_R1275_U141 , P2_R1275_U111 , P2_R1275_U66 );
nand NAND2_18660 ( P2_R1275_U142 , P2_U3960 , P2_R1275_U46 );
nand NAND2_18661 ( P2_R1275_U143 , P2_R1275_U110 , P2_R1275_U69 );
nand NAND2_18662 ( P2_R1275_U144 , P2_U3950 , P2_R1275_U45 );
nand NAND2_18663 ( P2_R1275_U145 , P2_R1275_U109 , P2_R1275_U71 );
nand NAND2_18664 ( P2_R1275_U146 , P2_U3952 , P2_R1275_U44 );
nand NAND2_18665 ( P2_R1275_U147 , P2_R1275_U108 , P2_R1275_U73 );
nand NAND2_18666 ( P2_R1275_U148 , P2_U3954 , P2_R1275_U43 );
nand NAND2_18667 ( P2_R1275_U149 , P2_R1275_U107 , P2_R1275_U75 );
nand NAND2_18668 ( P2_R1275_U150 , P2_U3956 , P2_R1275_U42 );
nand NAND2_18669 ( P2_R1275_U151 , P2_R1275_U106 , P2_R1275_U77 );
nand NAND2_18670 ( P2_R1275_U152 , P2_U3432 , P2_R1275_U80 );
nand NAND2_18671 ( P2_R1275_U153 , P2_U3427 , P2_R1275_U79 );
nand NAND2_18672 ( P2_R1275_U154 , P2_U3485 , P2_R1275_U41 );
nand NAND2_18673 ( P2_R1275_U155 , P2_R1275_U105 , P2_R1275_U81 );
nand NAND2_18674 ( P2_R1275_U156 , P2_U3480 , P2_R1275_U40 );
nand NAND2_18675 ( P2_R1275_U157 , P2_R1275_U104 , P2_R1275_U83 );
nand NAND2_18676 ( P2_R1275_U158 , P2_U3468 , P2_R1275_U37 );
nand NAND2_18677 ( P2_R1275_U159 , P2_R1275_U101 , P2_R1275_U85 );
and AND2_18678 ( P2_R1179_U6 , P2_R1179_U202 , P2_R1179_U201 );
and AND2_18679 ( P2_R1179_U7 , P2_R1179_U241 , P2_R1179_U240 );
and AND2_18680 ( P2_R1179_U8 , P2_R1179_U181 , P2_R1179_U256 );
and AND2_18681 ( P2_R1179_U9 , P2_R1179_U258 , P2_R1179_U257 );
and AND2_18682 ( P2_R1179_U10 , P2_R1179_U182 , P2_R1179_U282 );
and AND2_18683 ( P2_R1179_U11 , P2_R1179_U284 , P2_R1179_U283 );
nand NAND2_18684 ( P2_R1179_U12 , P2_R1179_U344 , P2_R1179_U347 );
nand NAND2_18685 ( P2_R1179_U13 , P2_R1179_U333 , P2_R1179_U336 );
nand NAND2_18686 ( P2_R1179_U14 , P2_R1179_U322 , P2_R1179_U325 );
nand NAND2_18687 ( P2_R1179_U15 , P2_R1179_U314 , P2_R1179_U316 );
nand NAND2_18688 ( P2_R1179_U16 , P2_R1179_U352 , P2_R1179_U312 );
nand NAND2_18689 ( P2_R1179_U17 , P2_R1179_U235 , P2_R1179_U237 );
nand NAND2_18690 ( P2_R1179_U18 , P2_R1179_U227 , P2_R1179_U230 );
nand NAND2_18691 ( P2_R1179_U19 , P2_R1179_U219 , P2_R1179_U221 );
nand NAND2_18692 ( P2_R1179_U20 , P2_R1179_U166 , P2_R1179_U350 );
not NOT1_18693 ( P2_R1179_U21 , P2_U3450 );
not NOT1_18694 ( P2_R1179_U22 , P2_U3444 );
not NOT1_18695 ( P2_R1179_U23 , P2_U3435 );
not NOT1_18696 ( P2_R1179_U24 , P2_U3427 );
not NOT1_18697 ( P2_R1179_U25 , P2_U3080 );
not NOT1_18698 ( P2_R1179_U26 , P2_U3438 );
not NOT1_18699 ( P2_R1179_U27 , P2_U3070 );
nand NAND2_18700 ( P2_R1179_U28 , P2_U3070 , P2_R1179_U23 );
not NOT1_18701 ( P2_R1179_U29 , P2_U3066 );
not NOT1_18702 ( P2_R1179_U30 , P2_U3447 );
not NOT1_18703 ( P2_R1179_U31 , P2_U3441 );
not NOT1_18704 ( P2_R1179_U32 , P2_U3073 );
not NOT1_18705 ( P2_R1179_U33 , P2_U3069 );
not NOT1_18706 ( P2_R1179_U34 , P2_U3062 );
nand NAND2_18707 ( P2_R1179_U35 , P2_U3062 , P2_R1179_U31 );
not NOT1_18708 ( P2_R1179_U36 , P2_U3453 );
not NOT1_18709 ( P2_R1179_U37 , P2_U3072 );
nand NAND2_18710 ( P2_R1179_U38 , P2_U3072 , P2_R1179_U21 );
not NOT1_18711 ( P2_R1179_U39 , P2_U3086 );
not NOT1_18712 ( P2_R1179_U40 , P2_U3456 );
not NOT1_18713 ( P2_R1179_U41 , P2_U3085 );
nand NAND2_18714 ( P2_R1179_U42 , P2_R1179_U208 , P2_R1179_U207 );
nand NAND2_18715 ( P2_R1179_U43 , P2_R1179_U35 , P2_R1179_U223 );
nand NAND3_18716 ( P2_R1179_U44 , P2_R1179_U192 , P2_R1179_U176 , P2_R1179_U351 );
not NOT1_18717 ( P2_R1179_U45 , P2_U3951 );
not NOT1_18718 ( P2_R1179_U46 , P2_U3459 );
not NOT1_18719 ( P2_R1179_U47 , P2_U3462 );
not NOT1_18720 ( P2_R1179_U48 , P2_U3065 );
not NOT1_18721 ( P2_R1179_U49 , P2_U3064 );
nand NAND2_18722 ( P2_R1179_U50 , P2_U3085 , P2_R1179_U40 );
not NOT1_18723 ( P2_R1179_U51 , P2_U3465 );
not NOT1_18724 ( P2_R1179_U52 , P2_U3074 );
not NOT1_18725 ( P2_R1179_U53 , P2_U3468 );
not NOT1_18726 ( P2_R1179_U54 , P2_U3082 );
not NOT1_18727 ( P2_R1179_U55 , P2_U3477 );
not NOT1_18728 ( P2_R1179_U56 , P2_U3474 );
not NOT1_18729 ( P2_R1179_U57 , P2_U3471 );
not NOT1_18730 ( P2_R1179_U58 , P2_U3075 );
not NOT1_18731 ( P2_R1179_U59 , P2_U3076 );
not NOT1_18732 ( P2_R1179_U60 , P2_U3081 );
nand NAND2_18733 ( P2_R1179_U61 , P2_U3081 , P2_R1179_U57 );
not NOT1_18734 ( P2_R1179_U62 , P2_U3480 );
not NOT1_18735 ( P2_R1179_U63 , P2_U3071 );
nand NAND2_18736 ( P2_R1179_U64 , P2_R1179_U268 , P2_R1179_U267 );
not NOT1_18737 ( P2_R1179_U65 , P2_U3084 );
not NOT1_18738 ( P2_R1179_U66 , P2_U3485 );
not NOT1_18739 ( P2_R1179_U67 , P2_U3083 );
not NOT1_18740 ( P2_R1179_U68 , P2_U3957 );
not NOT1_18741 ( P2_R1179_U69 , P2_U3078 );
not NOT1_18742 ( P2_R1179_U70 , P2_U3954 );
not NOT1_18743 ( P2_R1179_U71 , P2_U3955 );
not NOT1_18744 ( P2_R1179_U72 , P2_U3956 );
not NOT1_18745 ( P2_R1179_U73 , P2_U3068 );
not NOT1_18746 ( P2_R1179_U74 , P2_U3063 );
not NOT1_18747 ( P2_R1179_U75 , P2_U3077 );
nand NAND2_18748 ( P2_R1179_U76 , P2_U3077 , P2_R1179_U72 );
not NOT1_18749 ( P2_R1179_U77 , P2_U3953 );
not NOT1_18750 ( P2_R1179_U78 , P2_U3067 );
not NOT1_18751 ( P2_R1179_U79 , P2_U3952 );
not NOT1_18752 ( P2_R1179_U80 , P2_U3060 );
not NOT1_18753 ( P2_R1179_U81 , P2_U3950 );
not NOT1_18754 ( P2_R1179_U82 , P2_U3059 );
nand NAND2_18755 ( P2_R1179_U83 , P2_U3059 , P2_R1179_U45 );
not NOT1_18756 ( P2_R1179_U84 , P2_U3055 );
not NOT1_18757 ( P2_R1179_U85 , P2_U3949 );
not NOT1_18758 ( P2_R1179_U86 , P2_U3056 );
nand NAND2_18759 ( P2_R1179_U87 , P2_R1179_U128 , P2_R1179_U301 );
nand NAND2_18760 ( P2_R1179_U88 , P2_R1179_U298 , P2_R1179_U297 );
nand NAND2_18761 ( P2_R1179_U89 , P2_R1179_U76 , P2_R1179_U318 );
nand NAND2_18762 ( P2_R1179_U90 , P2_R1179_U61 , P2_R1179_U329 );
nand NAND2_18763 ( P2_R1179_U91 , P2_R1179_U50 , P2_R1179_U340 );
not NOT1_18764 ( P2_R1179_U92 , P2_U3079 );
nand NAND2_18765 ( P2_R1179_U93 , P2_R1179_U395 , P2_R1179_U394 );
nand NAND2_18766 ( P2_R1179_U94 , P2_R1179_U409 , P2_R1179_U408 );
nand NAND2_18767 ( P2_R1179_U95 , P2_R1179_U414 , P2_R1179_U413 );
nand NAND2_18768 ( P2_R1179_U96 , P2_R1179_U430 , P2_R1179_U429 );
nand NAND2_18769 ( P2_R1179_U97 , P2_R1179_U435 , P2_R1179_U434 );
nand NAND2_18770 ( P2_R1179_U98 , P2_R1179_U440 , P2_R1179_U439 );
nand NAND2_18771 ( P2_R1179_U99 , P2_R1179_U445 , P2_R1179_U444 );
nand NAND2_18772 ( P2_R1179_U100 , P2_R1179_U450 , P2_R1179_U449 );
nand NAND2_18773 ( P2_R1179_U101 , P2_R1179_U466 , P2_R1179_U465 );
nand NAND2_18774 ( P2_R1179_U102 , P2_R1179_U471 , P2_R1179_U470 );
nand NAND2_18775 ( P2_R1179_U103 , P2_R1179_U356 , P2_R1179_U355 );
nand NAND2_18776 ( P2_R1179_U104 , P2_R1179_U365 , P2_R1179_U364 );
nand NAND2_18777 ( P2_R1179_U105 , P2_R1179_U372 , P2_R1179_U371 );
nand NAND2_18778 ( P2_R1179_U106 , P2_R1179_U376 , P2_R1179_U375 );
nand NAND2_18779 ( P2_R1179_U107 , P2_R1179_U385 , P2_R1179_U384 );
nand NAND2_18780 ( P2_R1179_U108 , P2_R1179_U404 , P2_R1179_U403 );
nand NAND2_18781 ( P2_R1179_U109 , P2_R1179_U421 , P2_R1179_U420 );
nand NAND2_18782 ( P2_R1179_U110 , P2_R1179_U425 , P2_R1179_U424 );
nand NAND2_18783 ( P2_R1179_U111 , P2_R1179_U457 , P2_R1179_U456 );
nand NAND2_18784 ( P2_R1179_U112 , P2_R1179_U461 , P2_R1179_U460 );
nand NAND2_18785 ( P2_R1179_U113 , P2_R1179_U478 , P2_R1179_U477 );
and AND2_18786 ( P2_R1179_U114 , P2_R1179_U194 , P2_R1179_U184 );
and AND2_18787 ( P2_R1179_U115 , P2_R1179_U197 , P2_R1179_U198 );
and AND3_18788 ( P2_R1179_U116 , P2_R1179_U205 , P2_R1179_U200 , P2_R1179_U185 );
and AND2_18789 ( P2_R1179_U117 , P2_R1179_U210 , P2_R1179_U186 );
and AND2_18790 ( P2_R1179_U118 , P2_R1179_U213 , P2_R1179_U214 );
and AND3_18791 ( P2_R1179_U119 , P2_R1179_U358 , P2_R1179_U357 , P2_R1179_U38 );
and AND2_18792 ( P2_R1179_U120 , P2_R1179_U361 , P2_R1179_U186 );
and AND2_18793 ( P2_R1179_U121 , P2_R1179_U229 , P2_R1179_U6 );
and AND2_18794 ( P2_R1179_U122 , P2_R1179_U368 , P2_R1179_U185 );
and AND3_18795 ( P2_R1179_U123 , P2_R1179_U378 , P2_R1179_U377 , P2_R1179_U28 );
and AND2_18796 ( P2_R1179_U124 , P2_R1179_U381 , P2_R1179_U184 );
and AND3_18797 ( P2_R1179_U125 , P2_R1179_U239 , P2_R1179_U216 , P2_R1179_U180 );
and AND2_18798 ( P2_R1179_U126 , P2_R1179_U261 , P2_R1179_U8 );
and AND2_18799 ( P2_R1179_U127 , P2_R1179_U287 , P2_R1179_U10 );
and AND2_18800 ( P2_R1179_U128 , P2_R1179_U303 , P2_R1179_U304 );
and AND3_18801 ( P2_R1179_U129 , P2_R1179_U387 , P2_R1179_U386 , P2_R1179_U311 );
and AND2_18802 ( P2_R1179_U130 , P2_R1179_U308 , P2_R1179_U390 );
nand NAND2_18803 ( P2_R1179_U131 , P2_R1179_U392 , P2_R1179_U391 );
and AND3_18804 ( P2_R1179_U132 , P2_R1179_U397 , P2_R1179_U396 , P2_R1179_U83 );
and AND2_18805 ( P2_R1179_U133 , P2_R1179_U400 , P2_R1179_U183 );
nand NAND2_18806 ( P2_R1179_U134 , P2_R1179_U406 , P2_R1179_U405 );
nand NAND2_18807 ( P2_R1179_U135 , P2_R1179_U411 , P2_R1179_U410 );
and AND2_18808 ( P2_R1179_U136 , P2_R1179_U324 , P2_R1179_U11 );
and AND2_18809 ( P2_R1179_U137 , P2_R1179_U417 , P2_R1179_U182 );
nand NAND2_18810 ( P2_R1179_U138 , P2_R1179_U427 , P2_R1179_U426 );
nand NAND2_18811 ( P2_R1179_U139 , P2_R1179_U432 , P2_R1179_U431 );
nand NAND2_18812 ( P2_R1179_U140 , P2_R1179_U437 , P2_R1179_U436 );
nand NAND2_18813 ( P2_R1179_U141 , P2_R1179_U442 , P2_R1179_U441 );
nand NAND2_18814 ( P2_R1179_U142 , P2_R1179_U447 , P2_R1179_U446 );
and AND2_18815 ( P2_R1179_U143 , P2_R1179_U335 , P2_R1179_U9 );
and AND2_18816 ( P2_R1179_U144 , P2_R1179_U453 , P2_R1179_U181 );
nand NAND2_18817 ( P2_R1179_U145 , P2_R1179_U463 , P2_R1179_U462 );
nand NAND2_18818 ( P2_R1179_U146 , P2_R1179_U468 , P2_R1179_U467 );
and AND2_18819 ( P2_R1179_U147 , P2_R1179_U346 , P2_R1179_U7 );
and AND2_18820 ( P2_R1179_U148 , P2_R1179_U474 , P2_R1179_U180 );
and AND2_18821 ( P2_R1179_U149 , P2_R1179_U354 , P2_R1179_U353 );
nand NAND2_18822 ( P2_R1179_U150 , P2_R1179_U118 , P2_R1179_U211 );
and AND2_18823 ( P2_R1179_U151 , P2_R1179_U363 , P2_R1179_U362 );
and AND2_18824 ( P2_R1179_U152 , P2_R1179_U370 , P2_R1179_U369 );
and AND2_18825 ( P2_R1179_U153 , P2_R1179_U374 , P2_R1179_U373 );
nand NAND2_18826 ( P2_R1179_U154 , P2_R1179_U115 , P2_R1179_U195 );
and AND2_18827 ( P2_R1179_U155 , P2_R1179_U383 , P2_R1179_U382 );
not NOT1_18828 ( P2_R1179_U156 , P2_U3960 );
not NOT1_18829 ( P2_R1179_U157 , P2_U3057 );
and AND2_18830 ( P2_R1179_U158 , P2_R1179_U402 , P2_R1179_U401 );
nand NAND2_18831 ( P2_R1179_U159 , P2_R1179_U294 , P2_R1179_U293 );
nand NAND2_18832 ( P2_R1179_U160 , P2_R1179_U290 , P2_R1179_U289 );
and AND2_18833 ( P2_R1179_U161 , P2_R1179_U419 , P2_R1179_U418 );
and AND2_18834 ( P2_R1179_U162 , P2_R1179_U423 , P2_R1179_U422 );
nand NAND2_18835 ( P2_R1179_U163 , P2_R1179_U280 , P2_R1179_U279 );
nand NAND2_18836 ( P2_R1179_U164 , P2_R1179_U276 , P2_R1179_U275 );
not NOT1_18837 ( P2_R1179_U165 , P2_U3432 );
nand NAND2_18838 ( P2_R1179_U166 , P2_U3427 , P2_R1179_U92 );
nand NAND2_18839 ( P2_R1179_U167 , P2_R1179_U272 , P2_R1179_U271 );
not NOT1_18840 ( P2_R1179_U168 , P2_U3483 );
nand NAND2_18841 ( P2_R1179_U169 , P2_R1179_U264 , P2_R1179_U263 );
and AND2_18842 ( P2_R1179_U170 , P2_R1179_U455 , P2_R1179_U454 );
and AND2_18843 ( P2_R1179_U171 , P2_R1179_U459 , P2_R1179_U458 );
nand NAND2_18844 ( P2_R1179_U172 , P2_R1179_U254 , P2_R1179_U253 );
nand NAND2_18845 ( P2_R1179_U173 , P2_R1179_U250 , P2_R1179_U249 );
nand NAND2_18846 ( P2_R1179_U174 , P2_R1179_U246 , P2_R1179_U245 );
and AND2_18847 ( P2_R1179_U175 , P2_R1179_U476 , P2_R1179_U475 );
nand NAND2_18848 ( P2_R1179_U176 , P2_R1179_U166 , P2_R1179_U165 );
not NOT1_18849 ( P2_R1179_U177 , P2_R1179_U83 );
not NOT1_18850 ( P2_R1179_U178 , P2_R1179_U28 );
not NOT1_18851 ( P2_R1179_U179 , P2_R1179_U38 );
nand NAND2_18852 ( P2_R1179_U180 , P2_U3459 , P2_R1179_U49 );
nand NAND2_18853 ( P2_R1179_U181 , P2_U3474 , P2_R1179_U59 );
nand NAND2_18854 ( P2_R1179_U182 , P2_U3955 , P2_R1179_U74 );
nand NAND2_18855 ( P2_R1179_U183 , P2_U3951 , P2_R1179_U82 );
nand NAND2_18856 ( P2_R1179_U184 , P2_U3435 , P2_R1179_U27 );
nand NAND2_18857 ( P2_R1179_U185 , P2_U3444 , P2_R1179_U33 );
nand NAND2_18858 ( P2_R1179_U186 , P2_U3450 , P2_R1179_U37 );
not NOT1_18859 ( P2_R1179_U187 , P2_R1179_U61 );
not NOT1_18860 ( P2_R1179_U188 , P2_R1179_U76 );
not NOT1_18861 ( P2_R1179_U189 , P2_R1179_U35 );
not NOT1_18862 ( P2_R1179_U190 , P2_R1179_U50 );
not NOT1_18863 ( P2_R1179_U191 , P2_R1179_U166 );
nand NAND2_18864 ( P2_R1179_U192 , P2_U3080 , P2_R1179_U166 );
not NOT1_18865 ( P2_R1179_U193 , P2_R1179_U44 );
nand NAND2_18866 ( P2_R1179_U194 , P2_U3438 , P2_R1179_U29 );
nand NAND2_18867 ( P2_R1179_U195 , P2_R1179_U114 , P2_R1179_U44 );
nand NAND2_18868 ( P2_R1179_U196 , P2_R1179_U29 , P2_R1179_U28 );
nand NAND2_18869 ( P2_R1179_U197 , P2_R1179_U196 , P2_R1179_U26 );
nand NAND2_18870 ( P2_R1179_U198 , P2_U3066 , P2_R1179_U178 );
not NOT1_18871 ( P2_R1179_U199 , P2_R1179_U154 );
nand NAND2_18872 ( P2_R1179_U200 , P2_U3447 , P2_R1179_U32 );
nand NAND2_18873 ( P2_R1179_U201 , P2_U3073 , P2_R1179_U30 );
nand NAND2_18874 ( P2_R1179_U202 , P2_U3069 , P2_R1179_U22 );
nand NAND2_18875 ( P2_R1179_U203 , P2_R1179_U189 , P2_R1179_U185 );
nand NAND2_18876 ( P2_R1179_U204 , P2_R1179_U6 , P2_R1179_U203 );
nand NAND2_18877 ( P2_R1179_U205 , P2_U3441 , P2_R1179_U34 );
nand NAND2_18878 ( P2_R1179_U206 , P2_U3447 , P2_R1179_U32 );
nand NAND2_18879 ( P2_R1179_U207 , P2_R1179_U154 , P2_R1179_U116 );
nand NAND2_18880 ( P2_R1179_U208 , P2_R1179_U206 , P2_R1179_U204 );
not NOT1_18881 ( P2_R1179_U209 , P2_R1179_U42 );
nand NAND2_18882 ( P2_R1179_U210 , P2_U3453 , P2_R1179_U39 );
nand NAND2_18883 ( P2_R1179_U211 , P2_R1179_U117 , P2_R1179_U42 );
nand NAND2_18884 ( P2_R1179_U212 , P2_R1179_U39 , P2_R1179_U38 );
nand NAND2_18885 ( P2_R1179_U213 , P2_R1179_U212 , P2_R1179_U36 );
nand NAND2_18886 ( P2_R1179_U214 , P2_U3086 , P2_R1179_U179 );
not NOT1_18887 ( P2_R1179_U215 , P2_R1179_U150 );
nand NAND2_18888 ( P2_R1179_U216 , P2_U3456 , P2_R1179_U41 );
nand NAND2_18889 ( P2_R1179_U217 , P2_R1179_U216 , P2_R1179_U50 );
nand NAND2_18890 ( P2_R1179_U218 , P2_R1179_U209 , P2_R1179_U38 );
nand NAND2_18891 ( P2_R1179_U219 , P2_R1179_U120 , P2_R1179_U218 );
nand NAND2_18892 ( P2_R1179_U220 , P2_R1179_U42 , P2_R1179_U186 );
nand NAND2_18893 ( P2_R1179_U221 , P2_R1179_U119 , P2_R1179_U220 );
nand NAND2_18894 ( P2_R1179_U222 , P2_R1179_U38 , P2_R1179_U186 );
nand NAND2_18895 ( P2_R1179_U223 , P2_R1179_U205 , P2_R1179_U154 );
not NOT1_18896 ( P2_R1179_U224 , P2_R1179_U43 );
nand NAND2_18897 ( P2_R1179_U225 , P2_U3069 , P2_R1179_U22 );
nand NAND2_18898 ( P2_R1179_U226 , P2_R1179_U224 , P2_R1179_U225 );
nand NAND2_18899 ( P2_R1179_U227 , P2_R1179_U122 , P2_R1179_U226 );
nand NAND2_18900 ( P2_R1179_U228 , P2_R1179_U43 , P2_R1179_U185 );
nand NAND2_18901 ( P2_R1179_U229 , P2_U3447 , P2_R1179_U32 );
nand NAND2_18902 ( P2_R1179_U230 , P2_R1179_U121 , P2_R1179_U228 );
nand NAND2_18903 ( P2_R1179_U231 , P2_U3069 , P2_R1179_U22 );
nand NAND2_18904 ( P2_R1179_U232 , P2_R1179_U185 , P2_R1179_U231 );
nand NAND2_18905 ( P2_R1179_U233 , P2_R1179_U205 , P2_R1179_U35 );
nand NAND2_18906 ( P2_R1179_U234 , P2_R1179_U193 , P2_R1179_U28 );
nand NAND2_18907 ( P2_R1179_U235 , P2_R1179_U124 , P2_R1179_U234 );
nand NAND2_18908 ( P2_R1179_U236 , P2_R1179_U44 , P2_R1179_U184 );
nand NAND2_18909 ( P2_R1179_U237 , P2_R1179_U123 , P2_R1179_U236 );
nand NAND2_18910 ( P2_R1179_U238 , P2_R1179_U28 , P2_R1179_U184 );
nand NAND2_18911 ( P2_R1179_U239 , P2_U3462 , P2_R1179_U48 );
nand NAND2_18912 ( P2_R1179_U240 , P2_U3065 , P2_R1179_U47 );
nand NAND2_18913 ( P2_R1179_U241 , P2_U3064 , P2_R1179_U46 );
nand NAND2_18914 ( P2_R1179_U242 , P2_R1179_U190 , P2_R1179_U180 );
nand NAND2_18915 ( P2_R1179_U243 , P2_R1179_U7 , P2_R1179_U242 );
nand NAND2_18916 ( P2_R1179_U244 , P2_U3462 , P2_R1179_U48 );
nand NAND2_18917 ( P2_R1179_U245 , P2_R1179_U150 , P2_R1179_U125 );
nand NAND2_18918 ( P2_R1179_U246 , P2_R1179_U244 , P2_R1179_U243 );
not NOT1_18919 ( P2_R1179_U247 , P2_R1179_U174 );
nand NAND2_18920 ( P2_R1179_U248 , P2_U3465 , P2_R1179_U52 );
nand NAND2_18921 ( P2_R1179_U249 , P2_R1179_U248 , P2_R1179_U174 );
nand NAND2_18922 ( P2_R1179_U250 , P2_U3074 , P2_R1179_U51 );
not NOT1_18923 ( P2_R1179_U251 , P2_R1179_U173 );
nand NAND2_18924 ( P2_R1179_U252 , P2_U3468 , P2_R1179_U54 );
nand NAND2_18925 ( P2_R1179_U253 , P2_R1179_U252 , P2_R1179_U173 );
nand NAND2_18926 ( P2_R1179_U254 , P2_U3082 , P2_R1179_U53 );
not NOT1_18927 ( P2_R1179_U255 , P2_R1179_U172 );
nand NAND2_18928 ( P2_R1179_U256 , P2_U3477 , P2_R1179_U58 );
nand NAND2_18929 ( P2_R1179_U257 , P2_U3075 , P2_R1179_U55 );
nand NAND2_18930 ( P2_R1179_U258 , P2_U3076 , P2_R1179_U56 );
nand NAND2_18931 ( P2_R1179_U259 , P2_R1179_U187 , P2_R1179_U8 );
nand NAND2_18932 ( P2_R1179_U260 , P2_R1179_U9 , P2_R1179_U259 );
nand NAND2_18933 ( P2_R1179_U261 , P2_U3471 , P2_R1179_U60 );
nand NAND2_18934 ( P2_R1179_U262 , P2_U3477 , P2_R1179_U58 );
nand NAND2_18935 ( P2_R1179_U263 , P2_R1179_U126 , P2_R1179_U172 );
nand NAND2_18936 ( P2_R1179_U264 , P2_R1179_U262 , P2_R1179_U260 );
not NOT1_18937 ( P2_R1179_U265 , P2_R1179_U169 );
nand NAND2_18938 ( P2_R1179_U266 , P2_U3480 , P2_R1179_U63 );
nand NAND2_18939 ( P2_R1179_U267 , P2_R1179_U266 , P2_R1179_U169 );
nand NAND2_18940 ( P2_R1179_U268 , P2_U3071 , P2_R1179_U62 );
not NOT1_18941 ( P2_R1179_U269 , P2_R1179_U64 );
nand NAND2_18942 ( P2_R1179_U270 , P2_R1179_U269 , P2_R1179_U65 );
nand NAND2_18943 ( P2_R1179_U271 , P2_R1179_U270 , P2_R1179_U168 );
nand NAND2_18944 ( P2_R1179_U272 , P2_U3084 , P2_R1179_U64 );
not NOT1_18945 ( P2_R1179_U273 , P2_R1179_U167 );
nand NAND2_18946 ( P2_R1179_U274 , P2_U3485 , P2_R1179_U67 );
nand NAND2_18947 ( P2_R1179_U275 , P2_R1179_U274 , P2_R1179_U167 );
nand NAND2_18948 ( P2_R1179_U276 , P2_U3083 , P2_R1179_U66 );
not NOT1_18949 ( P2_R1179_U277 , P2_R1179_U164 );
nand NAND2_18950 ( P2_R1179_U278 , P2_U3957 , P2_R1179_U69 );
nand NAND2_18951 ( P2_R1179_U279 , P2_R1179_U278 , P2_R1179_U164 );
nand NAND2_18952 ( P2_R1179_U280 , P2_U3078 , P2_R1179_U68 );
not NOT1_18953 ( P2_R1179_U281 , P2_R1179_U163 );
nand NAND2_18954 ( P2_R1179_U282 , P2_U3954 , P2_R1179_U73 );
nand NAND2_18955 ( P2_R1179_U283 , P2_U3068 , P2_R1179_U70 );
nand NAND2_18956 ( P2_R1179_U284 , P2_U3063 , P2_R1179_U71 );
nand NAND2_18957 ( P2_R1179_U285 , P2_R1179_U188 , P2_R1179_U10 );
nand NAND2_18958 ( P2_R1179_U286 , P2_R1179_U11 , P2_R1179_U285 );
nand NAND2_18959 ( P2_R1179_U287 , P2_U3956 , P2_R1179_U75 );
nand NAND2_18960 ( P2_R1179_U288 , P2_U3954 , P2_R1179_U73 );
nand NAND2_18961 ( P2_R1179_U289 , P2_R1179_U127 , P2_R1179_U163 );
nand NAND2_18962 ( P2_R1179_U290 , P2_R1179_U288 , P2_R1179_U286 );
not NOT1_18963 ( P2_R1179_U291 , P2_R1179_U160 );
nand NAND2_18964 ( P2_R1179_U292 , P2_U3953 , P2_R1179_U78 );
nand NAND2_18965 ( P2_R1179_U293 , P2_R1179_U292 , P2_R1179_U160 );
nand NAND2_18966 ( P2_R1179_U294 , P2_U3067 , P2_R1179_U77 );
not NOT1_18967 ( P2_R1179_U295 , P2_R1179_U159 );
nand NAND2_18968 ( P2_R1179_U296 , P2_U3952 , P2_R1179_U80 );
nand NAND2_18969 ( P2_R1179_U297 , P2_R1179_U296 , P2_R1179_U159 );
nand NAND2_18970 ( P2_R1179_U298 , P2_U3060 , P2_R1179_U79 );
not NOT1_18971 ( P2_R1179_U299 , P2_R1179_U88 );
nand NAND2_18972 ( P2_R1179_U300 , P2_U3950 , P2_R1179_U84 );
nand NAND3_18973 ( P2_R1179_U301 , P2_R1179_U88 , P2_R1179_U183 , P2_R1179_U300 );
nand NAND2_18974 ( P2_R1179_U302 , P2_R1179_U84 , P2_R1179_U83 );
nand NAND2_18975 ( P2_R1179_U303 , P2_R1179_U302 , P2_R1179_U81 );
nand NAND2_18976 ( P2_R1179_U304 , P2_U3055 , P2_R1179_U177 );
not NOT1_18977 ( P2_R1179_U305 , P2_R1179_U87 );
nand NAND2_18978 ( P2_R1179_U306 , P2_U3056 , P2_R1179_U85 );
nand NAND2_18979 ( P2_R1179_U307 , P2_R1179_U305 , P2_R1179_U306 );
nand NAND2_18980 ( P2_R1179_U308 , P2_U3949 , P2_R1179_U86 );
nand NAND2_18981 ( P2_R1179_U309 , P2_U3949 , P2_R1179_U86 );
nand NAND2_18982 ( P2_R1179_U310 , P2_R1179_U309 , P2_R1179_U87 );
nand NAND2_18983 ( P2_R1179_U311 , P2_U3056 , P2_R1179_U85 );
nand NAND2_18984 ( P2_R1179_U312 , P2_R1179_U129 , P2_R1179_U310 );
nand NAND2_18985 ( P2_R1179_U313 , P2_R1179_U299 , P2_R1179_U83 );
nand NAND2_18986 ( P2_R1179_U314 , P2_R1179_U133 , P2_R1179_U313 );
nand NAND2_18987 ( P2_R1179_U315 , P2_R1179_U88 , P2_R1179_U183 );
nand NAND2_18988 ( P2_R1179_U316 , P2_R1179_U132 , P2_R1179_U315 );
nand NAND2_18989 ( P2_R1179_U317 , P2_R1179_U83 , P2_R1179_U183 );
nand NAND2_18990 ( P2_R1179_U318 , P2_R1179_U287 , P2_R1179_U163 );
not NOT1_18991 ( P2_R1179_U319 , P2_R1179_U89 );
nand NAND2_18992 ( P2_R1179_U320 , P2_U3063 , P2_R1179_U71 );
nand NAND2_18993 ( P2_R1179_U321 , P2_R1179_U319 , P2_R1179_U320 );
nand NAND2_18994 ( P2_R1179_U322 , P2_R1179_U137 , P2_R1179_U321 );
nand NAND2_18995 ( P2_R1179_U323 , P2_R1179_U89 , P2_R1179_U182 );
nand NAND2_18996 ( P2_R1179_U324 , P2_U3954 , P2_R1179_U73 );
nand NAND2_18997 ( P2_R1179_U325 , P2_R1179_U136 , P2_R1179_U323 );
nand NAND2_18998 ( P2_R1179_U326 , P2_U3063 , P2_R1179_U71 );
nand NAND2_18999 ( P2_R1179_U327 , P2_R1179_U182 , P2_R1179_U326 );
nand NAND2_19000 ( P2_R1179_U328 , P2_R1179_U287 , P2_R1179_U76 );
nand NAND2_19001 ( P2_R1179_U329 , P2_R1179_U261 , P2_R1179_U172 );
not NOT1_19002 ( P2_R1179_U330 , P2_R1179_U90 );
nand NAND2_19003 ( P2_R1179_U331 , P2_U3076 , P2_R1179_U56 );
nand NAND2_19004 ( P2_R1179_U332 , P2_R1179_U330 , P2_R1179_U331 );
nand NAND2_19005 ( P2_R1179_U333 , P2_R1179_U144 , P2_R1179_U332 );
nand NAND2_19006 ( P2_R1179_U334 , P2_R1179_U90 , P2_R1179_U181 );
nand NAND2_19007 ( P2_R1179_U335 , P2_U3477 , P2_R1179_U58 );
nand NAND2_19008 ( P2_R1179_U336 , P2_R1179_U143 , P2_R1179_U334 );
nand NAND2_19009 ( P2_R1179_U337 , P2_U3076 , P2_R1179_U56 );
nand NAND2_19010 ( P2_R1179_U338 , P2_R1179_U181 , P2_R1179_U337 );
nand NAND2_19011 ( P2_R1179_U339 , P2_R1179_U261 , P2_R1179_U61 );
nand NAND2_19012 ( P2_R1179_U340 , P2_R1179_U216 , P2_R1179_U150 );
not NOT1_19013 ( P2_R1179_U341 , P2_R1179_U91 );
nand NAND2_19014 ( P2_R1179_U342 , P2_U3064 , P2_R1179_U46 );
nand NAND2_19015 ( P2_R1179_U343 , P2_R1179_U341 , P2_R1179_U342 );
nand NAND2_19016 ( P2_R1179_U344 , P2_R1179_U148 , P2_R1179_U343 );
nand NAND2_19017 ( P2_R1179_U345 , P2_R1179_U91 , P2_R1179_U180 );
nand NAND2_19018 ( P2_R1179_U346 , P2_U3462 , P2_R1179_U48 );
nand NAND2_19019 ( P2_R1179_U347 , P2_R1179_U147 , P2_R1179_U345 );
nand NAND2_19020 ( P2_R1179_U348 , P2_U3064 , P2_R1179_U46 );
nand NAND2_19021 ( P2_R1179_U349 , P2_R1179_U180 , P2_R1179_U348 );
nand NAND2_19022 ( P2_R1179_U350 , P2_U3079 , P2_R1179_U24 );
nand NAND2_19023 ( P2_R1179_U351 , P2_U3080 , P2_R1179_U165 );
nand NAND2_19024 ( P2_R1179_U352 , P2_R1179_U130 , P2_R1179_U307 );
nand NAND2_19025 ( P2_R1179_U353 , P2_U3456 , P2_R1179_U41 );
nand NAND2_19026 ( P2_R1179_U354 , P2_U3085 , P2_R1179_U40 );
nand NAND2_19027 ( P2_R1179_U355 , P2_R1179_U217 , P2_R1179_U150 );
nand NAND2_19028 ( P2_R1179_U356 , P2_R1179_U215 , P2_R1179_U149 );
nand NAND2_19029 ( P2_R1179_U357 , P2_U3453 , P2_R1179_U39 );
nand NAND2_19030 ( P2_R1179_U358 , P2_U3086 , P2_R1179_U36 );
nand NAND2_19031 ( P2_R1179_U359 , P2_U3453 , P2_R1179_U39 );
nand NAND2_19032 ( P2_R1179_U360 , P2_U3086 , P2_R1179_U36 );
nand NAND2_19033 ( P2_R1179_U361 , P2_R1179_U360 , P2_R1179_U359 );
nand NAND2_19034 ( P2_R1179_U362 , P2_U3450 , P2_R1179_U37 );
nand NAND2_19035 ( P2_R1179_U363 , P2_U3072 , P2_R1179_U21 );
nand NAND2_19036 ( P2_R1179_U364 , P2_R1179_U222 , P2_R1179_U42 );
nand NAND2_19037 ( P2_R1179_U365 , P2_R1179_U151 , P2_R1179_U209 );
nand NAND2_19038 ( P2_R1179_U366 , P2_U3447 , P2_R1179_U32 );
nand NAND2_19039 ( P2_R1179_U367 , P2_U3073 , P2_R1179_U30 );
nand NAND2_19040 ( P2_R1179_U368 , P2_R1179_U367 , P2_R1179_U366 );
nand NAND2_19041 ( P2_R1179_U369 , P2_U3444 , P2_R1179_U33 );
nand NAND2_19042 ( P2_R1179_U370 , P2_U3069 , P2_R1179_U22 );
nand NAND2_19043 ( P2_R1179_U371 , P2_R1179_U232 , P2_R1179_U43 );
nand NAND2_19044 ( P2_R1179_U372 , P2_R1179_U152 , P2_R1179_U224 );
nand NAND2_19045 ( P2_R1179_U373 , P2_U3441 , P2_R1179_U34 );
nand NAND2_19046 ( P2_R1179_U374 , P2_U3062 , P2_R1179_U31 );
nand NAND2_19047 ( P2_R1179_U375 , P2_R1179_U233 , P2_R1179_U154 );
nand NAND2_19048 ( P2_R1179_U376 , P2_R1179_U199 , P2_R1179_U153 );
nand NAND2_19049 ( P2_R1179_U377 , P2_U3438 , P2_R1179_U29 );
nand NAND2_19050 ( P2_R1179_U378 , P2_U3066 , P2_R1179_U26 );
nand NAND2_19051 ( P2_R1179_U379 , P2_U3438 , P2_R1179_U29 );
nand NAND2_19052 ( P2_R1179_U380 , P2_U3066 , P2_R1179_U26 );
nand NAND2_19053 ( P2_R1179_U381 , P2_R1179_U380 , P2_R1179_U379 );
nand NAND2_19054 ( P2_R1179_U382 , P2_U3435 , P2_R1179_U27 );
nand NAND2_19055 ( P2_R1179_U383 , P2_U3070 , P2_R1179_U23 );
nand NAND2_19056 ( P2_R1179_U384 , P2_R1179_U238 , P2_R1179_U44 );
nand NAND2_19057 ( P2_R1179_U385 , P2_R1179_U155 , P2_R1179_U193 );
nand NAND2_19058 ( P2_R1179_U386 , P2_U3960 , P2_R1179_U157 );
nand NAND2_19059 ( P2_R1179_U387 , P2_U3057 , P2_R1179_U156 );
nand NAND2_19060 ( P2_R1179_U388 , P2_U3960 , P2_R1179_U157 );
nand NAND2_19061 ( P2_R1179_U389 , P2_U3057 , P2_R1179_U156 );
nand NAND2_19062 ( P2_R1179_U390 , P2_R1179_U389 , P2_R1179_U388 );
nand NAND2_19063 ( P2_R1179_U391 , P2_U3949 , P2_R1179_U86 );
nand NAND2_19064 ( P2_R1179_U392 , P2_U3056 , P2_R1179_U85 );
not NOT1_19065 ( P2_R1179_U393 , P2_R1179_U131 );
nand NAND2_19066 ( P2_R1179_U394 , P2_R1179_U393 , P2_R1179_U305 );
nand NAND2_19067 ( P2_R1179_U395 , P2_R1179_U131 , P2_R1179_U87 );
nand NAND2_19068 ( P2_R1179_U396 , P2_U3950 , P2_R1179_U84 );
nand NAND2_19069 ( P2_R1179_U397 , P2_U3055 , P2_R1179_U81 );
nand NAND2_19070 ( P2_R1179_U398 , P2_U3950 , P2_R1179_U84 );
nand NAND2_19071 ( P2_R1179_U399 , P2_U3055 , P2_R1179_U81 );
nand NAND2_19072 ( P2_R1179_U400 , P2_R1179_U399 , P2_R1179_U398 );
nand NAND2_19073 ( P2_R1179_U401 , P2_U3951 , P2_R1179_U82 );
nand NAND2_19074 ( P2_R1179_U402 , P2_U3059 , P2_R1179_U45 );
nand NAND2_19075 ( P2_R1179_U403 , P2_R1179_U317 , P2_R1179_U88 );
nand NAND2_19076 ( P2_R1179_U404 , P2_R1179_U158 , P2_R1179_U299 );
nand NAND2_19077 ( P2_R1179_U405 , P2_U3952 , P2_R1179_U80 );
nand NAND2_19078 ( P2_R1179_U406 , P2_U3060 , P2_R1179_U79 );
not NOT1_19079 ( P2_R1179_U407 , P2_R1179_U134 );
nand NAND2_19080 ( P2_R1179_U408 , P2_R1179_U295 , P2_R1179_U407 );
nand NAND2_19081 ( P2_R1179_U409 , P2_R1179_U134 , P2_R1179_U159 );
nand NAND2_19082 ( P2_R1179_U410 , P2_U3953 , P2_R1179_U78 );
nand NAND2_19083 ( P2_R1179_U411 , P2_U3067 , P2_R1179_U77 );
not NOT1_19084 ( P2_R1179_U412 , P2_R1179_U135 );
nand NAND2_19085 ( P2_R1179_U413 , P2_R1179_U291 , P2_R1179_U412 );
nand NAND2_19086 ( P2_R1179_U414 , P2_R1179_U135 , P2_R1179_U160 );
nand NAND2_19087 ( P2_R1179_U415 , P2_U3954 , P2_R1179_U73 );
nand NAND2_19088 ( P2_R1179_U416 , P2_U3068 , P2_R1179_U70 );
nand NAND2_19089 ( P2_R1179_U417 , P2_R1179_U416 , P2_R1179_U415 );
nand NAND2_19090 ( P2_R1179_U418 , P2_U3955 , P2_R1179_U74 );
nand NAND2_19091 ( P2_R1179_U419 , P2_U3063 , P2_R1179_U71 );
nand NAND2_19092 ( P2_R1179_U420 , P2_R1179_U327 , P2_R1179_U89 );
nand NAND2_19093 ( P2_R1179_U421 , P2_R1179_U161 , P2_R1179_U319 );
nand NAND2_19094 ( P2_R1179_U422 , P2_U3956 , P2_R1179_U75 );
nand NAND2_19095 ( P2_R1179_U423 , P2_U3077 , P2_R1179_U72 );
nand NAND2_19096 ( P2_R1179_U424 , P2_R1179_U328 , P2_R1179_U163 );
nand NAND2_19097 ( P2_R1179_U425 , P2_R1179_U281 , P2_R1179_U162 );
nand NAND2_19098 ( P2_R1179_U426 , P2_U3957 , P2_R1179_U69 );
nand NAND2_19099 ( P2_R1179_U427 , P2_U3078 , P2_R1179_U68 );
not NOT1_19100 ( P2_R1179_U428 , P2_R1179_U138 );
nand NAND2_19101 ( P2_R1179_U429 , P2_R1179_U277 , P2_R1179_U428 );
nand NAND2_19102 ( P2_R1179_U430 , P2_R1179_U138 , P2_R1179_U164 );
nand NAND2_19103 ( P2_R1179_U431 , P2_U3432 , P2_R1179_U25 );
nand NAND2_19104 ( P2_R1179_U432 , P2_U3080 , P2_R1179_U165 );
not NOT1_19105 ( P2_R1179_U433 , P2_R1179_U139 );
nand NAND2_19106 ( P2_R1179_U434 , P2_R1179_U191 , P2_R1179_U433 );
nand NAND2_19107 ( P2_R1179_U435 , P2_R1179_U139 , P2_R1179_U166 );
nand NAND2_19108 ( P2_R1179_U436 , P2_U3485 , P2_R1179_U67 );
nand NAND2_19109 ( P2_R1179_U437 , P2_U3083 , P2_R1179_U66 );
not NOT1_19110 ( P2_R1179_U438 , P2_R1179_U140 );
nand NAND2_19111 ( P2_R1179_U439 , P2_R1179_U273 , P2_R1179_U438 );
nand NAND2_19112 ( P2_R1179_U440 , P2_R1179_U140 , P2_R1179_U167 );
nand NAND2_19113 ( P2_R1179_U441 , P2_U3483 , P2_R1179_U65 );
nand NAND2_19114 ( P2_R1179_U442 , P2_U3084 , P2_R1179_U168 );
not NOT1_19115 ( P2_R1179_U443 , P2_R1179_U141 );
nand NAND2_19116 ( P2_R1179_U444 , P2_R1179_U443 , P2_R1179_U269 );
nand NAND2_19117 ( P2_R1179_U445 , P2_R1179_U141 , P2_R1179_U64 );
nand NAND2_19118 ( P2_R1179_U446 , P2_U3480 , P2_R1179_U63 );
nand NAND2_19119 ( P2_R1179_U447 , P2_U3071 , P2_R1179_U62 );
not NOT1_19120 ( P2_R1179_U448 , P2_R1179_U142 );
nand NAND2_19121 ( P2_R1179_U449 , P2_R1179_U265 , P2_R1179_U448 );
nand NAND2_19122 ( P2_R1179_U450 , P2_R1179_U142 , P2_R1179_U169 );
nand NAND2_19123 ( P2_R1179_U451 , P2_U3477 , P2_R1179_U58 );
nand NAND2_19124 ( P2_R1179_U452 , P2_U3075 , P2_R1179_U55 );
nand NAND2_19125 ( P2_R1179_U453 , P2_R1179_U452 , P2_R1179_U451 );
nand NAND2_19126 ( P2_R1179_U454 , P2_U3474 , P2_R1179_U59 );
nand NAND2_19127 ( P2_R1179_U455 , P2_U3076 , P2_R1179_U56 );
nand NAND2_19128 ( P2_R1179_U456 , P2_R1179_U338 , P2_R1179_U90 );
nand NAND2_19129 ( P2_R1179_U457 , P2_R1179_U170 , P2_R1179_U330 );
nand NAND2_19130 ( P2_R1179_U458 , P2_U3471 , P2_R1179_U60 );
nand NAND2_19131 ( P2_R1179_U459 , P2_U3081 , P2_R1179_U57 );
nand NAND2_19132 ( P2_R1179_U460 , P2_R1179_U339 , P2_R1179_U172 );
nand NAND2_19133 ( P2_R1179_U461 , P2_R1179_U255 , P2_R1179_U171 );
nand NAND2_19134 ( P2_R1179_U462 , P2_U3468 , P2_R1179_U54 );
nand NAND2_19135 ( P2_R1179_U463 , P2_U3082 , P2_R1179_U53 );
not NOT1_19136 ( P2_R1179_U464 , P2_R1179_U145 );
nand NAND2_19137 ( P2_R1179_U465 , P2_R1179_U251 , P2_R1179_U464 );
nand NAND2_19138 ( P2_R1179_U466 , P2_R1179_U145 , P2_R1179_U173 );
nand NAND2_19139 ( P2_R1179_U467 , P2_U3465 , P2_R1179_U52 );
nand NAND2_19140 ( P2_R1179_U468 , P2_U3074 , P2_R1179_U51 );
not NOT1_19141 ( P2_R1179_U469 , P2_R1179_U146 );
nand NAND2_19142 ( P2_R1179_U470 , P2_R1179_U247 , P2_R1179_U469 );
nand NAND2_19143 ( P2_R1179_U471 , P2_R1179_U146 , P2_R1179_U174 );
nand NAND2_19144 ( P2_R1179_U472 , P2_U3462 , P2_R1179_U48 );
nand NAND2_19145 ( P2_R1179_U473 , P2_U3065 , P2_R1179_U47 );
nand NAND2_19146 ( P2_R1179_U474 , P2_R1179_U473 , P2_R1179_U472 );
nand NAND2_19147 ( P2_R1179_U475 , P2_U3459 , P2_R1179_U49 );
nand NAND2_19148 ( P2_R1179_U476 , P2_U3064 , P2_R1179_U46 );
nand NAND2_19149 ( P2_R1179_U477 , P2_R1179_U349 , P2_R1179_U91 );
nand NAND2_19150 ( P2_R1179_U478 , P2_R1179_U175 , P2_R1179_U341 );
and AND2_19151 ( P2_R1215_U4 , P2_R1215_U179 , P2_R1215_U178 );
and AND2_19152 ( P2_R1215_U5 , P2_R1215_U180 , P2_R1215_U181 );
and AND2_19153 ( P2_R1215_U6 , P2_R1215_U197 , P2_R1215_U196 );
and AND2_19154 ( P2_R1215_U7 , P2_R1215_U237 , P2_R1215_U236 );
and AND2_19155 ( P2_R1215_U8 , P2_R1215_U246 , P2_R1215_U245 );
and AND2_19156 ( P2_R1215_U9 , P2_R1215_U264 , P2_R1215_U263 );
and AND2_19157 ( P2_R1215_U10 , P2_R1215_U272 , P2_R1215_U271 );
and AND2_19158 ( P2_R1215_U11 , P2_R1215_U351 , P2_R1215_U348 );
and AND2_19159 ( P2_R1215_U12 , P2_R1215_U344 , P2_R1215_U341 );
and AND2_19160 ( P2_R1215_U13 , P2_R1215_U335 , P2_R1215_U332 );
and AND2_19161 ( P2_R1215_U14 , P2_R1215_U326 , P2_R1215_U323 );
and AND2_19162 ( P2_R1215_U15 , P2_R1215_U320 , P2_R1215_U318 );
and AND2_19163 ( P2_R1215_U16 , P2_R1215_U313 , P2_R1215_U310 );
and AND2_19164 ( P2_R1215_U17 , P2_R1215_U235 , P2_R1215_U232 );
and AND2_19165 ( P2_R1215_U18 , P2_R1215_U227 , P2_R1215_U224 );
and AND2_19166 ( P2_R1215_U19 , P2_R1215_U213 , P2_R1215_U210 );
not NOT1_19167 ( P2_R1215_U20 , P2_U3447 );
not NOT1_19168 ( P2_R1215_U21 , P2_U3073 );
not NOT1_19169 ( P2_R1215_U22 , P2_U3072 );
nand NAND2_19170 ( P2_R1215_U23 , P2_U3073 , P2_U3447 );
not NOT1_19171 ( P2_R1215_U24 , P2_U3450 );
not NOT1_19172 ( P2_R1215_U25 , P2_U3441 );
not NOT1_19173 ( P2_R1215_U26 , P2_U3062 );
not NOT1_19174 ( P2_R1215_U27 , P2_U3069 );
not NOT1_19175 ( P2_R1215_U28 , P2_U3435 );
not NOT1_19176 ( P2_R1215_U29 , P2_U3070 );
not NOT1_19177 ( P2_R1215_U30 , P2_U3427 );
not NOT1_19178 ( P2_R1215_U31 , P2_U3079 );
nand NAND2_19179 ( P2_R1215_U32 , P2_U3079 , P2_U3427 );
not NOT1_19180 ( P2_R1215_U33 , P2_U3438 );
not NOT1_19181 ( P2_R1215_U34 , P2_U3066 );
nand NAND2_19182 ( P2_R1215_U35 , P2_U3062 , P2_U3441 );
not NOT1_19183 ( P2_R1215_U36 , P2_U3444 );
not NOT1_19184 ( P2_R1215_U37 , P2_U3453 );
not NOT1_19185 ( P2_R1215_U38 , P2_U3086 );
not NOT1_19186 ( P2_R1215_U39 , P2_U3085 );
not NOT1_19187 ( P2_R1215_U40 , P2_U3456 );
nand NAND2_19188 ( P2_R1215_U41 , P2_R1215_U62 , P2_R1215_U205 );
nand NAND2_19189 ( P2_R1215_U42 , P2_R1215_U118 , P2_R1215_U193 );
nand NAND2_19190 ( P2_R1215_U43 , P2_R1215_U182 , P2_R1215_U183 );
nand NAND2_19191 ( P2_R1215_U44 , P2_U3432 , P2_U3080 );
nand NAND2_19192 ( P2_R1215_U45 , P2_R1215_U122 , P2_R1215_U219 );
nand NAND2_19193 ( P2_R1215_U46 , P2_R1215_U216 , P2_R1215_U215 );
not NOT1_19194 ( P2_R1215_U47 , P2_U3950 );
not NOT1_19195 ( P2_R1215_U48 , P2_U3055 );
not NOT1_19196 ( P2_R1215_U49 , P2_U3059 );
not NOT1_19197 ( P2_R1215_U50 , P2_U3951 );
not NOT1_19198 ( P2_R1215_U51 , P2_U3952 );
not NOT1_19199 ( P2_R1215_U52 , P2_U3060 );
not NOT1_19200 ( P2_R1215_U53 , P2_U3953 );
not NOT1_19201 ( P2_R1215_U54 , P2_U3067 );
not NOT1_19202 ( P2_R1215_U55 , P2_U3956 );
not NOT1_19203 ( P2_R1215_U56 , P2_U3077 );
not NOT1_19204 ( P2_R1215_U57 , P2_U3477 );
not NOT1_19205 ( P2_R1215_U58 , P2_U3075 );
not NOT1_19206 ( P2_R1215_U59 , P2_U3071 );
nand NAND2_19207 ( P2_R1215_U60 , P2_U3075 , P2_U3477 );
not NOT1_19208 ( P2_R1215_U61 , P2_U3480 );
nand NAND2_19209 ( P2_R1215_U62 , P2_U3086 , P2_U3453 );
not NOT1_19210 ( P2_R1215_U63 , P2_U3459 );
not NOT1_19211 ( P2_R1215_U64 , P2_U3064 );
not NOT1_19212 ( P2_R1215_U65 , P2_U3465 );
not NOT1_19213 ( P2_R1215_U66 , P2_U3074 );
not NOT1_19214 ( P2_R1215_U67 , P2_U3462 );
not NOT1_19215 ( P2_R1215_U68 , P2_U3065 );
nand NAND2_19216 ( P2_R1215_U69 , P2_U3065 , P2_U3462 );
not NOT1_19217 ( P2_R1215_U70 , P2_U3468 );
not NOT1_19218 ( P2_R1215_U71 , P2_U3082 );
not NOT1_19219 ( P2_R1215_U72 , P2_U3471 );
not NOT1_19220 ( P2_R1215_U73 , P2_U3081 );
not NOT1_19221 ( P2_R1215_U74 , P2_U3474 );
not NOT1_19222 ( P2_R1215_U75 , P2_U3076 );
not NOT1_19223 ( P2_R1215_U76 , P2_U3483 );
not NOT1_19224 ( P2_R1215_U77 , P2_U3084 );
nand NAND2_19225 ( P2_R1215_U78 , P2_U3084 , P2_U3483 );
not NOT1_19226 ( P2_R1215_U79 , P2_U3485 );
not NOT1_19227 ( P2_R1215_U80 , P2_U3083 );
nand NAND2_19228 ( P2_R1215_U81 , P2_U3083 , P2_U3485 );
not NOT1_19229 ( P2_R1215_U82 , P2_U3957 );
not NOT1_19230 ( P2_R1215_U83 , P2_U3955 );
not NOT1_19231 ( P2_R1215_U84 , P2_U3063 );
not NOT1_19232 ( P2_R1215_U85 , P2_U3954 );
not NOT1_19233 ( P2_R1215_U86 , P2_U3068 );
nand NAND2_19234 ( P2_R1215_U87 , P2_U3951 , P2_U3059 );
not NOT1_19235 ( P2_R1215_U88 , P2_U3056 );
not NOT1_19236 ( P2_R1215_U89 , P2_U3949 );
nand NAND2_19237 ( P2_R1215_U90 , P2_R1215_U306 , P2_R1215_U176 );
not NOT1_19238 ( P2_R1215_U91 , P2_U3078 );
nand NAND2_19239 ( P2_R1215_U92 , P2_R1215_U78 , P2_R1215_U315 );
nand NAND2_19240 ( P2_R1215_U93 , P2_R1215_U261 , P2_R1215_U260 );
nand NAND2_19241 ( P2_R1215_U94 , P2_R1215_U69 , P2_R1215_U337 );
nand NAND2_19242 ( P2_R1215_U95 , P2_R1215_U457 , P2_R1215_U456 );
nand NAND2_19243 ( P2_R1215_U96 , P2_R1215_U504 , P2_R1215_U503 );
nand NAND2_19244 ( P2_R1215_U97 , P2_R1215_U375 , P2_R1215_U374 );
nand NAND2_19245 ( P2_R1215_U98 , P2_R1215_U380 , P2_R1215_U379 );
nand NAND2_19246 ( P2_R1215_U99 , P2_R1215_U387 , P2_R1215_U386 );
nand NAND2_19247 ( P2_R1215_U100 , P2_R1215_U394 , P2_R1215_U393 );
nand NAND2_19248 ( P2_R1215_U101 , P2_R1215_U399 , P2_R1215_U398 );
nand NAND2_19249 ( P2_R1215_U102 , P2_R1215_U408 , P2_R1215_U407 );
nand NAND2_19250 ( P2_R1215_U103 , P2_R1215_U415 , P2_R1215_U414 );
nand NAND2_19251 ( P2_R1215_U104 , P2_R1215_U422 , P2_R1215_U421 );
nand NAND2_19252 ( P2_R1215_U105 , P2_R1215_U429 , P2_R1215_U428 );
nand NAND2_19253 ( P2_R1215_U106 , P2_R1215_U434 , P2_R1215_U433 );
nand NAND2_19254 ( P2_R1215_U107 , P2_R1215_U441 , P2_R1215_U440 );
nand NAND2_19255 ( P2_R1215_U108 , P2_R1215_U448 , P2_R1215_U447 );
nand NAND2_19256 ( P2_R1215_U109 , P2_R1215_U462 , P2_R1215_U461 );
nand NAND2_19257 ( P2_R1215_U110 , P2_R1215_U467 , P2_R1215_U466 );
nand NAND2_19258 ( P2_R1215_U111 , P2_R1215_U474 , P2_R1215_U473 );
nand NAND2_19259 ( P2_R1215_U112 , P2_R1215_U481 , P2_R1215_U480 );
nand NAND2_19260 ( P2_R1215_U113 , P2_R1215_U488 , P2_R1215_U487 );
nand NAND2_19261 ( P2_R1215_U114 , P2_R1215_U495 , P2_R1215_U494 );
nand NAND2_19262 ( P2_R1215_U115 , P2_R1215_U500 , P2_R1215_U499 );
and AND2_19263 ( P2_R1215_U116 , P2_U3435 , P2_U3070 );
and AND2_19264 ( P2_R1215_U117 , P2_R1215_U189 , P2_R1215_U187 );
and AND2_19265 ( P2_R1215_U118 , P2_R1215_U194 , P2_R1215_U192 );
and AND2_19266 ( P2_R1215_U119 , P2_R1215_U201 , P2_R1215_U200 );
and AND3_19267 ( P2_R1215_U120 , P2_R1215_U382 , P2_R1215_U381 , P2_R1215_U23 );
and AND2_19268 ( P2_R1215_U121 , P2_R1215_U212 , P2_R1215_U6 );
and AND2_19269 ( P2_R1215_U122 , P2_R1215_U220 , P2_R1215_U218 );
and AND3_19270 ( P2_R1215_U123 , P2_R1215_U389 , P2_R1215_U388 , P2_R1215_U35 );
and AND2_19271 ( P2_R1215_U124 , P2_R1215_U226 , P2_R1215_U4 );
and AND2_19272 ( P2_R1215_U125 , P2_R1215_U234 , P2_R1215_U181 );
and AND2_19273 ( P2_R1215_U126 , P2_R1215_U204 , P2_R1215_U7 );
and AND2_19274 ( P2_R1215_U127 , P2_R1215_U239 , P2_R1215_U171 );
and AND2_19275 ( P2_R1215_U128 , P2_R1215_U250 , P2_R1215_U8 );
and AND2_19276 ( P2_R1215_U129 , P2_R1215_U248 , P2_R1215_U172 );
and AND2_19277 ( P2_R1215_U130 , P2_R1215_U268 , P2_R1215_U267 );
and AND2_19278 ( P2_R1215_U131 , P2_R1215_U10 , P2_R1215_U282 );
and AND2_19279 ( P2_R1215_U132 , P2_R1215_U285 , P2_R1215_U280 );
and AND2_19280 ( P2_R1215_U133 , P2_R1215_U301 , P2_R1215_U298 );
and AND2_19281 ( P2_R1215_U134 , P2_R1215_U368 , P2_R1215_U302 );
and AND2_19282 ( P2_R1215_U135 , P2_R1215_U160 , P2_R1215_U278 );
and AND3_19283 ( P2_R1215_U136 , P2_R1215_U455 , P2_R1215_U454 , P2_R1215_U81 );
and AND2_19284 ( P2_R1215_U137 , P2_R1215_U325 , P2_R1215_U10 );
and AND3_19285 ( P2_R1215_U138 , P2_R1215_U469 , P2_R1215_U468 , P2_R1215_U60 );
and AND2_19286 ( P2_R1215_U139 , P2_R1215_U334 , P2_R1215_U9 );
and AND3_19287 ( P2_R1215_U140 , P2_R1215_U490 , P2_R1215_U489 , P2_R1215_U172 );
and AND2_19288 ( P2_R1215_U141 , P2_R1215_U343 , P2_R1215_U8 );
and AND3_19289 ( P2_R1215_U142 , P2_R1215_U502 , P2_R1215_U501 , P2_R1215_U171 );
and AND2_19290 ( P2_R1215_U143 , P2_R1215_U350 , P2_R1215_U7 );
nand NAND2_19291 ( P2_R1215_U144 , P2_R1215_U119 , P2_R1215_U202 );
nand NAND2_19292 ( P2_R1215_U145 , P2_R1215_U217 , P2_R1215_U229 );
not NOT1_19293 ( P2_R1215_U146 , P2_U3057 );
not NOT1_19294 ( P2_R1215_U147 , P2_U3960 );
and AND2_19295 ( P2_R1215_U148 , P2_R1215_U403 , P2_R1215_U402 );
nand NAND3_19296 ( P2_R1215_U149 , P2_R1215_U304 , P2_R1215_U169 , P2_R1215_U364 );
and AND2_19297 ( P2_R1215_U150 , P2_R1215_U410 , P2_R1215_U409 );
nand NAND3_19298 ( P2_R1215_U151 , P2_R1215_U370 , P2_R1215_U369 , P2_R1215_U134 );
and AND2_19299 ( P2_R1215_U152 , P2_R1215_U417 , P2_R1215_U416 );
nand NAND3_19300 ( P2_R1215_U153 , P2_R1215_U365 , P2_R1215_U299 , P2_R1215_U87 );
and AND2_19301 ( P2_R1215_U154 , P2_R1215_U424 , P2_R1215_U423 );
nand NAND2_19302 ( P2_R1215_U155 , P2_R1215_U293 , P2_R1215_U292 );
and AND2_19303 ( P2_R1215_U156 , P2_R1215_U436 , P2_R1215_U435 );
nand NAND2_19304 ( P2_R1215_U157 , P2_R1215_U289 , P2_R1215_U288 );
and AND2_19305 ( P2_R1215_U158 , P2_R1215_U443 , P2_R1215_U442 );
nand NAND2_19306 ( P2_R1215_U159 , P2_R1215_U132 , P2_R1215_U284 );
and AND2_19307 ( P2_R1215_U160 , P2_R1215_U450 , P2_R1215_U449 );
nand NAND2_19308 ( P2_R1215_U161 , P2_R1215_U44 , P2_R1215_U327 );
nand NAND2_19309 ( P2_R1215_U162 , P2_R1215_U130 , P2_R1215_U269 );
and AND2_19310 ( P2_R1215_U163 , P2_R1215_U476 , P2_R1215_U475 );
nand NAND2_19311 ( P2_R1215_U164 , P2_R1215_U257 , P2_R1215_U256 );
and AND2_19312 ( P2_R1215_U165 , P2_R1215_U483 , P2_R1215_U482 );
nand NAND2_19313 ( P2_R1215_U166 , P2_R1215_U253 , P2_R1215_U252 );
nand NAND2_19314 ( P2_R1215_U167 , P2_R1215_U243 , P2_R1215_U242 );
nand NAND2_19315 ( P2_R1215_U168 , P2_R1215_U367 , P2_R1215_U366 );
nand NAND2_19316 ( P2_R1215_U169 , P2_U3056 , P2_R1215_U151 );
not NOT1_19317 ( P2_R1215_U170 , P2_R1215_U35 );
nand NAND2_19318 ( P2_R1215_U171 , P2_U3456 , P2_U3085 );
nand NAND2_19319 ( P2_R1215_U172 , P2_U3074 , P2_U3465 );
nand NAND2_19320 ( P2_R1215_U173 , P2_U3060 , P2_U3952 );
not NOT1_19321 ( P2_R1215_U174 , P2_R1215_U69 );
not NOT1_19322 ( P2_R1215_U175 , P2_R1215_U78 );
nand NAND2_19323 ( P2_R1215_U176 , P2_U3067 , P2_U3953 );
not NOT1_19324 ( P2_R1215_U177 , P2_R1215_U62 );
or OR2_19325 ( P2_R1215_U178 , P2_U3069 , P2_U3444 );
or OR2_19326 ( P2_R1215_U179 , P2_U3062 , P2_U3441 );
or OR2_19327 ( P2_R1215_U180 , P2_U3438 , P2_U3066 );
or OR2_19328 ( P2_R1215_U181 , P2_U3435 , P2_U3070 );
not NOT1_19329 ( P2_R1215_U182 , P2_R1215_U32 );
or OR2_19330 ( P2_R1215_U183 , P2_U3432 , P2_U3080 );
not NOT1_19331 ( P2_R1215_U184 , P2_R1215_U43 );
not NOT1_19332 ( P2_R1215_U185 , P2_R1215_U44 );
nand NAND2_19333 ( P2_R1215_U186 , P2_R1215_U43 , P2_R1215_U44 );
nand NAND2_19334 ( P2_R1215_U187 , P2_R1215_U116 , P2_R1215_U180 );
nand NAND2_19335 ( P2_R1215_U188 , P2_R1215_U5 , P2_R1215_U186 );
nand NAND2_19336 ( P2_R1215_U189 , P2_U3066 , P2_U3438 );
nand NAND2_19337 ( P2_R1215_U190 , P2_R1215_U117 , P2_R1215_U188 );
nand NAND2_19338 ( P2_R1215_U191 , P2_R1215_U36 , P2_R1215_U35 );
nand NAND2_19339 ( P2_R1215_U192 , P2_U3069 , P2_R1215_U191 );
nand NAND2_19340 ( P2_R1215_U193 , P2_R1215_U4 , P2_R1215_U190 );
nand NAND2_19341 ( P2_R1215_U194 , P2_U3444 , P2_R1215_U170 );
not NOT1_19342 ( P2_R1215_U195 , P2_R1215_U42 );
or OR2_19343 ( P2_R1215_U196 , P2_U3072 , P2_U3450 );
or OR2_19344 ( P2_R1215_U197 , P2_U3073 , P2_U3447 );
not NOT1_19345 ( P2_R1215_U198 , P2_R1215_U23 );
nand NAND2_19346 ( P2_R1215_U199 , P2_R1215_U24 , P2_R1215_U23 );
nand NAND2_19347 ( P2_R1215_U200 , P2_U3072 , P2_R1215_U199 );
nand NAND2_19348 ( P2_R1215_U201 , P2_U3450 , P2_R1215_U198 );
nand NAND2_19349 ( P2_R1215_U202 , P2_R1215_U6 , P2_R1215_U42 );
not NOT1_19350 ( P2_R1215_U203 , P2_R1215_U144 );
or OR2_19351 ( P2_R1215_U204 , P2_U3453 , P2_U3086 );
nand NAND2_19352 ( P2_R1215_U205 , P2_R1215_U204 , P2_R1215_U144 );
not NOT1_19353 ( P2_R1215_U206 , P2_R1215_U41 );
or OR2_19354 ( P2_R1215_U207 , P2_U3085 , P2_U3456 );
or OR2_19355 ( P2_R1215_U208 , P2_U3447 , P2_U3073 );
nand NAND2_19356 ( P2_R1215_U209 , P2_R1215_U208 , P2_R1215_U42 );
nand NAND2_19357 ( P2_R1215_U210 , P2_R1215_U120 , P2_R1215_U209 );
nand NAND2_19358 ( P2_R1215_U211 , P2_R1215_U195 , P2_R1215_U23 );
nand NAND2_19359 ( P2_R1215_U212 , P2_U3450 , P2_U3072 );
nand NAND2_19360 ( P2_R1215_U213 , P2_R1215_U121 , P2_R1215_U211 );
or OR2_19361 ( P2_R1215_U214 , P2_U3073 , P2_U3447 );
nand NAND2_19362 ( P2_R1215_U215 , P2_R1215_U185 , P2_R1215_U181 );
nand NAND2_19363 ( P2_R1215_U216 , P2_U3070 , P2_U3435 );
not NOT1_19364 ( P2_R1215_U217 , P2_R1215_U46 );
nand NAND2_19365 ( P2_R1215_U218 , P2_R1215_U184 , P2_R1215_U5 );
nand NAND2_19366 ( P2_R1215_U219 , P2_R1215_U46 , P2_R1215_U180 );
nand NAND2_19367 ( P2_R1215_U220 , P2_U3066 , P2_U3438 );
not NOT1_19368 ( P2_R1215_U221 , P2_R1215_U45 );
or OR2_19369 ( P2_R1215_U222 , P2_U3441 , P2_U3062 );
nand NAND2_19370 ( P2_R1215_U223 , P2_R1215_U222 , P2_R1215_U45 );
nand NAND2_19371 ( P2_R1215_U224 , P2_R1215_U123 , P2_R1215_U223 );
nand NAND2_19372 ( P2_R1215_U225 , P2_R1215_U221 , P2_R1215_U35 );
nand NAND2_19373 ( P2_R1215_U226 , P2_U3444 , P2_U3069 );
nand NAND2_19374 ( P2_R1215_U227 , P2_R1215_U124 , P2_R1215_U225 );
or OR2_19375 ( P2_R1215_U228 , P2_U3062 , P2_U3441 );
nand NAND2_19376 ( P2_R1215_U229 , P2_R1215_U184 , P2_R1215_U181 );
not NOT1_19377 ( P2_R1215_U230 , P2_R1215_U145 );
nand NAND2_19378 ( P2_R1215_U231 , P2_U3066 , P2_U3438 );
nand NAND4_19379 ( P2_R1215_U232 , P2_R1215_U401 , P2_R1215_U400 , P2_R1215_U44 , P2_R1215_U43 );
nand NAND2_19380 ( P2_R1215_U233 , P2_R1215_U44 , P2_R1215_U43 );
nand NAND2_19381 ( P2_R1215_U234 , P2_U3070 , P2_U3435 );
nand NAND2_19382 ( P2_R1215_U235 , P2_R1215_U125 , P2_R1215_U233 );
or OR2_19383 ( P2_R1215_U236 , P2_U3085 , P2_U3456 );
or OR2_19384 ( P2_R1215_U237 , P2_U3064 , P2_U3459 );
nand NAND2_19385 ( P2_R1215_U238 , P2_R1215_U177 , P2_R1215_U7 );
nand NAND2_19386 ( P2_R1215_U239 , P2_U3064 , P2_U3459 );
nand NAND2_19387 ( P2_R1215_U240 , P2_R1215_U127 , P2_R1215_U238 );
or OR2_19388 ( P2_R1215_U241 , P2_U3459 , P2_U3064 );
nand NAND2_19389 ( P2_R1215_U242 , P2_R1215_U126 , P2_R1215_U144 );
nand NAND2_19390 ( P2_R1215_U243 , P2_R1215_U241 , P2_R1215_U240 );
not NOT1_19391 ( P2_R1215_U244 , P2_R1215_U167 );
or OR2_19392 ( P2_R1215_U245 , P2_U3082 , P2_U3468 );
or OR2_19393 ( P2_R1215_U246 , P2_U3074 , P2_U3465 );
nand NAND2_19394 ( P2_R1215_U247 , P2_R1215_U174 , P2_R1215_U8 );
nand NAND2_19395 ( P2_R1215_U248 , P2_U3082 , P2_U3468 );
nand NAND2_19396 ( P2_R1215_U249 , P2_R1215_U129 , P2_R1215_U247 );
or OR2_19397 ( P2_R1215_U250 , P2_U3462 , P2_U3065 );
or OR2_19398 ( P2_R1215_U251 , P2_U3468 , P2_U3082 );
nand NAND2_19399 ( P2_R1215_U252 , P2_R1215_U128 , P2_R1215_U167 );
nand NAND2_19400 ( P2_R1215_U253 , P2_R1215_U251 , P2_R1215_U249 );
not NOT1_19401 ( P2_R1215_U254 , P2_R1215_U166 );
or OR2_19402 ( P2_R1215_U255 , P2_U3471 , P2_U3081 );
nand NAND2_19403 ( P2_R1215_U256 , P2_R1215_U255 , P2_R1215_U166 );
nand NAND2_19404 ( P2_R1215_U257 , P2_U3081 , P2_U3471 );
not NOT1_19405 ( P2_R1215_U258 , P2_R1215_U164 );
or OR2_19406 ( P2_R1215_U259 , P2_U3474 , P2_U3076 );
nand NAND2_19407 ( P2_R1215_U260 , P2_R1215_U259 , P2_R1215_U164 );
nand NAND2_19408 ( P2_R1215_U261 , P2_U3076 , P2_U3474 );
not NOT1_19409 ( P2_R1215_U262 , P2_R1215_U93 );
or OR2_19410 ( P2_R1215_U263 , P2_U3071 , P2_U3480 );
or OR2_19411 ( P2_R1215_U264 , P2_U3075 , P2_U3477 );
not NOT1_19412 ( P2_R1215_U265 , P2_R1215_U60 );
nand NAND2_19413 ( P2_R1215_U266 , P2_R1215_U61 , P2_R1215_U60 );
nand NAND2_19414 ( P2_R1215_U267 , P2_U3071 , P2_R1215_U266 );
nand NAND2_19415 ( P2_R1215_U268 , P2_U3480 , P2_R1215_U265 );
nand NAND2_19416 ( P2_R1215_U269 , P2_R1215_U9 , P2_R1215_U93 );
not NOT1_19417 ( P2_R1215_U270 , P2_R1215_U162 );
or OR2_19418 ( P2_R1215_U271 , P2_U3078 , P2_U3957 );
or OR2_19419 ( P2_R1215_U272 , P2_U3083 , P2_U3485 );
or OR2_19420 ( P2_R1215_U273 , P2_U3077 , P2_U3956 );
not NOT1_19421 ( P2_R1215_U274 , P2_R1215_U81 );
nand NAND2_19422 ( P2_R1215_U275 , P2_U3957 , P2_R1215_U274 );
nand NAND2_19423 ( P2_R1215_U276 , P2_R1215_U275 , P2_R1215_U91 );
nand NAND2_19424 ( P2_R1215_U277 , P2_R1215_U81 , P2_R1215_U82 );
nand NAND2_19425 ( P2_R1215_U278 , P2_R1215_U277 , P2_R1215_U276 );
nand NAND2_19426 ( P2_R1215_U279 , P2_R1215_U175 , P2_R1215_U10 );
nand NAND2_19427 ( P2_R1215_U280 , P2_U3077 , P2_U3956 );
nand NAND2_19428 ( P2_R1215_U281 , P2_R1215_U278 , P2_R1215_U279 );
or OR2_19429 ( P2_R1215_U282 , P2_U3483 , P2_U3084 );
or OR2_19430 ( P2_R1215_U283 , P2_U3956 , P2_U3077 );
nand NAND3_19431 ( P2_R1215_U284 , P2_R1215_U273 , P2_R1215_U162 , P2_R1215_U131 );
nand NAND2_19432 ( P2_R1215_U285 , P2_R1215_U283 , P2_R1215_U281 );
not NOT1_19433 ( P2_R1215_U286 , P2_R1215_U159 );
or OR2_19434 ( P2_R1215_U287 , P2_U3955 , P2_U3063 );
nand NAND2_19435 ( P2_R1215_U288 , P2_R1215_U287 , P2_R1215_U159 );
nand NAND2_19436 ( P2_R1215_U289 , P2_U3063 , P2_U3955 );
not NOT1_19437 ( P2_R1215_U290 , P2_R1215_U157 );
or OR2_19438 ( P2_R1215_U291 , P2_U3954 , P2_U3068 );
nand NAND2_19439 ( P2_R1215_U292 , P2_R1215_U291 , P2_R1215_U157 );
nand NAND2_19440 ( P2_R1215_U293 , P2_U3068 , P2_U3954 );
not NOT1_19441 ( P2_R1215_U294 , P2_R1215_U155 );
or OR2_19442 ( P2_R1215_U295 , P2_U3060 , P2_U3952 );
nand NAND2_19443 ( P2_R1215_U296 , P2_R1215_U176 , P2_R1215_U173 );
not NOT1_19444 ( P2_R1215_U297 , P2_R1215_U87 );
or OR2_19445 ( P2_R1215_U298 , P2_U3953 , P2_U3067 );
nand NAND3_19446 ( P2_R1215_U299 , P2_R1215_U155 , P2_R1215_U298 , P2_R1215_U168 );
not NOT1_19447 ( P2_R1215_U300 , P2_R1215_U153 );
or OR2_19448 ( P2_R1215_U301 , P2_U3950 , P2_U3055 );
nand NAND2_19449 ( P2_R1215_U302 , P2_U3055 , P2_U3950 );
not NOT1_19450 ( P2_R1215_U303 , P2_R1215_U151 );
nand NAND2_19451 ( P2_R1215_U304 , P2_U3949 , P2_R1215_U151 );
not NOT1_19452 ( P2_R1215_U305 , P2_R1215_U149 );
nand NAND2_19453 ( P2_R1215_U306 , P2_R1215_U298 , P2_R1215_U155 );
not NOT1_19454 ( P2_R1215_U307 , P2_R1215_U90 );
or OR2_19455 ( P2_R1215_U308 , P2_U3952 , P2_U3060 );
nand NAND2_19456 ( P2_R1215_U309 , P2_R1215_U308 , P2_R1215_U90 );
nand NAND3_19457 ( P2_R1215_U310 , P2_R1215_U309 , P2_R1215_U173 , P2_R1215_U154 );
nand NAND2_19458 ( P2_R1215_U311 , P2_R1215_U307 , P2_R1215_U173 );
nand NAND2_19459 ( P2_R1215_U312 , P2_U3951 , P2_U3059 );
nand NAND3_19460 ( P2_R1215_U313 , P2_R1215_U311 , P2_R1215_U312 , P2_R1215_U168 );
or OR2_19461 ( P2_R1215_U314 , P2_U3060 , P2_U3952 );
nand NAND2_19462 ( P2_R1215_U315 , P2_R1215_U282 , P2_R1215_U162 );
not NOT1_19463 ( P2_R1215_U316 , P2_R1215_U92 );
nand NAND2_19464 ( P2_R1215_U317 , P2_R1215_U10 , P2_R1215_U92 );
nand NAND2_19465 ( P2_R1215_U318 , P2_R1215_U135 , P2_R1215_U317 );
nand NAND2_19466 ( P2_R1215_U319 , P2_R1215_U317 , P2_R1215_U278 );
nand NAND2_19467 ( P2_R1215_U320 , P2_R1215_U453 , P2_R1215_U319 );
or OR2_19468 ( P2_R1215_U321 , P2_U3485 , P2_U3083 );
nand NAND2_19469 ( P2_R1215_U322 , P2_R1215_U321 , P2_R1215_U92 );
nand NAND2_19470 ( P2_R1215_U323 , P2_R1215_U136 , P2_R1215_U322 );
nand NAND2_19471 ( P2_R1215_U324 , P2_R1215_U316 , P2_R1215_U81 );
nand NAND2_19472 ( P2_R1215_U325 , P2_U3078 , P2_U3957 );
nand NAND2_19473 ( P2_R1215_U326 , P2_R1215_U137 , P2_R1215_U324 );
or OR2_19474 ( P2_R1215_U327 , P2_U3432 , P2_U3080 );
not NOT1_19475 ( P2_R1215_U328 , P2_R1215_U161 );
or OR2_19476 ( P2_R1215_U329 , P2_U3083 , P2_U3485 );
or OR2_19477 ( P2_R1215_U330 , P2_U3477 , P2_U3075 );
nand NAND2_19478 ( P2_R1215_U331 , P2_R1215_U330 , P2_R1215_U93 );
nand NAND2_19479 ( P2_R1215_U332 , P2_R1215_U138 , P2_R1215_U331 );
nand NAND2_19480 ( P2_R1215_U333 , P2_R1215_U262 , P2_R1215_U60 );
nand NAND2_19481 ( P2_R1215_U334 , P2_U3480 , P2_U3071 );
nand NAND2_19482 ( P2_R1215_U335 , P2_R1215_U139 , P2_R1215_U333 );
or OR2_19483 ( P2_R1215_U336 , P2_U3075 , P2_U3477 );
nand NAND2_19484 ( P2_R1215_U337 , P2_R1215_U250 , P2_R1215_U167 );
not NOT1_19485 ( P2_R1215_U338 , P2_R1215_U94 );
or OR2_19486 ( P2_R1215_U339 , P2_U3465 , P2_U3074 );
nand NAND2_19487 ( P2_R1215_U340 , P2_R1215_U339 , P2_R1215_U94 );
nand NAND2_19488 ( P2_R1215_U341 , P2_R1215_U140 , P2_R1215_U340 );
nand NAND2_19489 ( P2_R1215_U342 , P2_R1215_U338 , P2_R1215_U172 );
nand NAND2_19490 ( P2_R1215_U343 , P2_U3082 , P2_U3468 );
nand NAND2_19491 ( P2_R1215_U344 , P2_R1215_U141 , P2_R1215_U342 );
or OR2_19492 ( P2_R1215_U345 , P2_U3074 , P2_U3465 );
or OR2_19493 ( P2_R1215_U346 , P2_U3456 , P2_U3085 );
nand NAND2_19494 ( P2_R1215_U347 , P2_R1215_U346 , P2_R1215_U41 );
nand NAND2_19495 ( P2_R1215_U348 , P2_R1215_U142 , P2_R1215_U347 );
nand NAND2_19496 ( P2_R1215_U349 , P2_R1215_U206 , P2_R1215_U171 );
nand NAND2_19497 ( P2_R1215_U350 , P2_U3064 , P2_U3459 );
nand NAND2_19498 ( P2_R1215_U351 , P2_R1215_U143 , P2_R1215_U349 );
nand NAND2_19499 ( P2_R1215_U352 , P2_R1215_U207 , P2_R1215_U171 );
nand NAND2_19500 ( P2_R1215_U353 , P2_R1215_U204 , P2_R1215_U62 );
nand NAND2_19501 ( P2_R1215_U354 , P2_R1215_U214 , P2_R1215_U23 );
nand NAND2_19502 ( P2_R1215_U355 , P2_R1215_U228 , P2_R1215_U35 );
nand NAND2_19503 ( P2_R1215_U356 , P2_R1215_U231 , P2_R1215_U180 );
nand NAND2_19504 ( P2_R1215_U357 , P2_R1215_U314 , P2_R1215_U173 );
nand NAND2_19505 ( P2_R1215_U358 , P2_R1215_U298 , P2_R1215_U176 );
nand NAND2_19506 ( P2_R1215_U359 , P2_R1215_U329 , P2_R1215_U81 );
nand NAND2_19507 ( P2_R1215_U360 , P2_R1215_U282 , P2_R1215_U78 );
nand NAND2_19508 ( P2_R1215_U361 , P2_R1215_U336 , P2_R1215_U60 );
nand NAND2_19509 ( P2_R1215_U362 , P2_R1215_U345 , P2_R1215_U172 );
nand NAND2_19510 ( P2_R1215_U363 , P2_R1215_U250 , P2_R1215_U69 );
nand NAND2_19511 ( P2_R1215_U364 , P2_U3949 , P2_U3056 );
nand NAND2_19512 ( P2_R1215_U365 , P2_R1215_U296 , P2_R1215_U168 );
nand NAND2_19513 ( P2_R1215_U366 , P2_U3059 , P2_R1215_U295 );
nand NAND2_19514 ( P2_R1215_U367 , P2_U3951 , P2_R1215_U295 );
nand NAND3_19515 ( P2_R1215_U368 , P2_R1215_U296 , P2_R1215_U168 , P2_R1215_U301 );
nand NAND3_19516 ( P2_R1215_U369 , P2_R1215_U155 , P2_R1215_U168 , P2_R1215_U133 );
nand NAND2_19517 ( P2_R1215_U370 , P2_R1215_U297 , P2_R1215_U301 );
nand NAND2_19518 ( P2_R1215_U371 , P2_U3085 , P2_R1215_U40 );
nand NAND2_19519 ( P2_R1215_U372 , P2_U3456 , P2_R1215_U39 );
nand NAND2_19520 ( P2_R1215_U373 , P2_R1215_U372 , P2_R1215_U371 );
nand NAND2_19521 ( P2_R1215_U374 , P2_R1215_U352 , P2_R1215_U41 );
nand NAND2_19522 ( P2_R1215_U375 , P2_R1215_U373 , P2_R1215_U206 );
nand NAND2_19523 ( P2_R1215_U376 , P2_U3086 , P2_R1215_U37 );
nand NAND2_19524 ( P2_R1215_U377 , P2_U3453 , P2_R1215_U38 );
nand NAND2_19525 ( P2_R1215_U378 , P2_R1215_U377 , P2_R1215_U376 );
nand NAND2_19526 ( P2_R1215_U379 , P2_R1215_U353 , P2_R1215_U144 );
nand NAND2_19527 ( P2_R1215_U380 , P2_R1215_U203 , P2_R1215_U378 );
nand NAND2_19528 ( P2_R1215_U381 , P2_U3072 , P2_R1215_U24 );
nand NAND2_19529 ( P2_R1215_U382 , P2_U3450 , P2_R1215_U22 );
nand NAND2_19530 ( P2_R1215_U383 , P2_U3073 , P2_R1215_U20 );
nand NAND2_19531 ( P2_R1215_U384 , P2_U3447 , P2_R1215_U21 );
nand NAND2_19532 ( P2_R1215_U385 , P2_R1215_U384 , P2_R1215_U383 );
nand NAND2_19533 ( P2_R1215_U386 , P2_R1215_U354 , P2_R1215_U42 );
nand NAND2_19534 ( P2_R1215_U387 , P2_R1215_U385 , P2_R1215_U195 );
nand NAND2_19535 ( P2_R1215_U388 , P2_U3069 , P2_R1215_U36 );
nand NAND2_19536 ( P2_R1215_U389 , P2_U3444 , P2_R1215_U27 );
nand NAND2_19537 ( P2_R1215_U390 , P2_U3062 , P2_R1215_U25 );
nand NAND2_19538 ( P2_R1215_U391 , P2_U3441 , P2_R1215_U26 );
nand NAND2_19539 ( P2_R1215_U392 , P2_R1215_U391 , P2_R1215_U390 );
nand NAND2_19540 ( P2_R1215_U393 , P2_R1215_U355 , P2_R1215_U45 );
nand NAND2_19541 ( P2_R1215_U394 , P2_R1215_U392 , P2_R1215_U221 );
nand NAND2_19542 ( P2_R1215_U395 , P2_U3066 , P2_R1215_U33 );
nand NAND2_19543 ( P2_R1215_U396 , P2_U3438 , P2_R1215_U34 );
nand NAND2_19544 ( P2_R1215_U397 , P2_R1215_U396 , P2_R1215_U395 );
nand NAND2_19545 ( P2_R1215_U398 , P2_R1215_U356 , P2_R1215_U145 );
nand NAND2_19546 ( P2_R1215_U399 , P2_R1215_U230 , P2_R1215_U397 );
nand NAND2_19547 ( P2_R1215_U400 , P2_U3070 , P2_R1215_U28 );
nand NAND2_19548 ( P2_R1215_U401 , P2_U3435 , P2_R1215_U29 );
nand NAND2_19549 ( P2_R1215_U402 , P2_U3057 , P2_R1215_U147 );
nand NAND2_19550 ( P2_R1215_U403 , P2_U3960 , P2_R1215_U146 );
nand NAND2_19551 ( P2_R1215_U404 , P2_U3057 , P2_R1215_U147 );
nand NAND2_19552 ( P2_R1215_U405 , P2_U3960 , P2_R1215_U146 );
nand NAND2_19553 ( P2_R1215_U406 , P2_R1215_U405 , P2_R1215_U404 );
nand NAND2_19554 ( P2_R1215_U407 , P2_R1215_U148 , P2_R1215_U149 );
nand NAND2_19555 ( P2_R1215_U408 , P2_R1215_U305 , P2_R1215_U406 );
nand NAND2_19556 ( P2_R1215_U409 , P2_U3056 , P2_R1215_U89 );
nand NAND2_19557 ( P2_R1215_U410 , P2_U3949 , P2_R1215_U88 );
nand NAND2_19558 ( P2_R1215_U411 , P2_U3056 , P2_R1215_U89 );
nand NAND2_19559 ( P2_R1215_U412 , P2_U3949 , P2_R1215_U88 );
nand NAND2_19560 ( P2_R1215_U413 , P2_R1215_U412 , P2_R1215_U411 );
nand NAND2_19561 ( P2_R1215_U414 , P2_R1215_U150 , P2_R1215_U151 );
nand NAND2_19562 ( P2_R1215_U415 , P2_R1215_U303 , P2_R1215_U413 );
nand NAND2_19563 ( P2_R1215_U416 , P2_U3055 , P2_R1215_U47 );
nand NAND2_19564 ( P2_R1215_U417 , P2_U3950 , P2_R1215_U48 );
nand NAND2_19565 ( P2_R1215_U418 , P2_U3055 , P2_R1215_U47 );
nand NAND2_19566 ( P2_R1215_U419 , P2_U3950 , P2_R1215_U48 );
nand NAND2_19567 ( P2_R1215_U420 , P2_R1215_U419 , P2_R1215_U418 );
nand NAND2_19568 ( P2_R1215_U421 , P2_R1215_U152 , P2_R1215_U153 );
nand NAND2_19569 ( P2_R1215_U422 , P2_R1215_U300 , P2_R1215_U420 );
nand NAND2_19570 ( P2_R1215_U423 , P2_U3059 , P2_R1215_U50 );
nand NAND2_19571 ( P2_R1215_U424 , P2_U3951 , P2_R1215_U49 );
nand NAND2_19572 ( P2_R1215_U425 , P2_U3060 , P2_R1215_U51 );
nand NAND2_19573 ( P2_R1215_U426 , P2_U3952 , P2_R1215_U52 );
nand NAND2_19574 ( P2_R1215_U427 , P2_R1215_U426 , P2_R1215_U425 );
nand NAND2_19575 ( P2_R1215_U428 , P2_R1215_U357 , P2_R1215_U90 );
nand NAND2_19576 ( P2_R1215_U429 , P2_R1215_U427 , P2_R1215_U307 );
nand NAND2_19577 ( P2_R1215_U430 , P2_U3067 , P2_R1215_U53 );
nand NAND2_19578 ( P2_R1215_U431 , P2_U3953 , P2_R1215_U54 );
nand NAND2_19579 ( P2_R1215_U432 , P2_R1215_U431 , P2_R1215_U430 );
nand NAND2_19580 ( P2_R1215_U433 , P2_R1215_U358 , P2_R1215_U155 );
nand NAND2_19581 ( P2_R1215_U434 , P2_R1215_U294 , P2_R1215_U432 );
nand NAND2_19582 ( P2_R1215_U435 , P2_U3068 , P2_R1215_U85 );
nand NAND2_19583 ( P2_R1215_U436 , P2_U3954 , P2_R1215_U86 );
nand NAND2_19584 ( P2_R1215_U437 , P2_U3068 , P2_R1215_U85 );
nand NAND2_19585 ( P2_R1215_U438 , P2_U3954 , P2_R1215_U86 );
nand NAND2_19586 ( P2_R1215_U439 , P2_R1215_U438 , P2_R1215_U437 );
nand NAND2_19587 ( P2_R1215_U440 , P2_R1215_U156 , P2_R1215_U157 );
nand NAND2_19588 ( P2_R1215_U441 , P2_R1215_U290 , P2_R1215_U439 );
nand NAND2_19589 ( P2_R1215_U442 , P2_U3063 , P2_R1215_U83 );
nand NAND2_19590 ( P2_R1215_U443 , P2_U3955 , P2_R1215_U84 );
nand NAND2_19591 ( P2_R1215_U444 , P2_U3063 , P2_R1215_U83 );
nand NAND2_19592 ( P2_R1215_U445 , P2_U3955 , P2_R1215_U84 );
nand NAND2_19593 ( P2_R1215_U446 , P2_R1215_U445 , P2_R1215_U444 );
nand NAND2_19594 ( P2_R1215_U447 , P2_R1215_U158 , P2_R1215_U159 );
nand NAND2_19595 ( P2_R1215_U448 , P2_R1215_U286 , P2_R1215_U446 );
nand NAND2_19596 ( P2_R1215_U449 , P2_U3077 , P2_R1215_U55 );
nand NAND2_19597 ( P2_R1215_U450 , P2_U3956 , P2_R1215_U56 );
nand NAND2_19598 ( P2_R1215_U451 , P2_U3077 , P2_R1215_U55 );
nand NAND2_19599 ( P2_R1215_U452 , P2_U3956 , P2_R1215_U56 );
nand NAND2_19600 ( P2_R1215_U453 , P2_R1215_U452 , P2_R1215_U451 );
nand NAND2_19601 ( P2_R1215_U454 , P2_U3078 , P2_R1215_U82 );
nand NAND2_19602 ( P2_R1215_U455 , P2_U3957 , P2_R1215_U91 );
nand NAND2_19603 ( P2_R1215_U456 , P2_R1215_U182 , P2_R1215_U161 );
nand NAND2_19604 ( P2_R1215_U457 , P2_R1215_U328 , P2_R1215_U32 );
nand NAND2_19605 ( P2_R1215_U458 , P2_U3083 , P2_R1215_U79 );
nand NAND2_19606 ( P2_R1215_U459 , P2_U3485 , P2_R1215_U80 );
nand NAND2_19607 ( P2_R1215_U460 , P2_R1215_U459 , P2_R1215_U458 );
nand NAND2_19608 ( P2_R1215_U461 , P2_R1215_U359 , P2_R1215_U92 );
nand NAND2_19609 ( P2_R1215_U462 , P2_R1215_U460 , P2_R1215_U316 );
nand NAND2_19610 ( P2_R1215_U463 , P2_U3084 , P2_R1215_U76 );
nand NAND2_19611 ( P2_R1215_U464 , P2_U3483 , P2_R1215_U77 );
nand NAND2_19612 ( P2_R1215_U465 , P2_R1215_U464 , P2_R1215_U463 );
nand NAND2_19613 ( P2_R1215_U466 , P2_R1215_U360 , P2_R1215_U162 );
nand NAND2_19614 ( P2_R1215_U467 , P2_R1215_U270 , P2_R1215_U465 );
nand NAND2_19615 ( P2_R1215_U468 , P2_U3071 , P2_R1215_U61 );
nand NAND2_19616 ( P2_R1215_U469 , P2_U3480 , P2_R1215_U59 );
nand NAND2_19617 ( P2_R1215_U470 , P2_U3075 , P2_R1215_U57 );
nand NAND2_19618 ( P2_R1215_U471 , P2_U3477 , P2_R1215_U58 );
nand NAND2_19619 ( P2_R1215_U472 , P2_R1215_U471 , P2_R1215_U470 );
nand NAND2_19620 ( P2_R1215_U473 , P2_R1215_U361 , P2_R1215_U93 );
nand NAND2_19621 ( P2_R1215_U474 , P2_R1215_U472 , P2_R1215_U262 );
nand NAND2_19622 ( P2_R1215_U475 , P2_U3076 , P2_R1215_U74 );
nand NAND2_19623 ( P2_R1215_U476 , P2_U3474 , P2_R1215_U75 );
nand NAND2_19624 ( P2_R1215_U477 , P2_U3076 , P2_R1215_U74 );
nand NAND2_19625 ( P2_R1215_U478 , P2_U3474 , P2_R1215_U75 );
nand NAND2_19626 ( P2_R1215_U479 , P2_R1215_U478 , P2_R1215_U477 );
nand NAND2_19627 ( P2_R1215_U480 , P2_R1215_U163 , P2_R1215_U164 );
nand NAND2_19628 ( P2_R1215_U481 , P2_R1215_U258 , P2_R1215_U479 );
nand NAND2_19629 ( P2_R1215_U482 , P2_U3081 , P2_R1215_U72 );
nand NAND2_19630 ( P2_R1215_U483 , P2_U3471 , P2_R1215_U73 );
nand NAND2_19631 ( P2_R1215_U484 , P2_U3081 , P2_R1215_U72 );
nand NAND2_19632 ( P2_R1215_U485 , P2_U3471 , P2_R1215_U73 );
nand NAND2_19633 ( P2_R1215_U486 , P2_R1215_U485 , P2_R1215_U484 );
nand NAND2_19634 ( P2_R1215_U487 , P2_R1215_U165 , P2_R1215_U166 );
nand NAND2_19635 ( P2_R1215_U488 , P2_R1215_U254 , P2_R1215_U486 );
nand NAND2_19636 ( P2_R1215_U489 , P2_U3082 , P2_R1215_U70 );
nand NAND2_19637 ( P2_R1215_U490 , P2_U3468 , P2_R1215_U71 );
nand NAND2_19638 ( P2_R1215_U491 , P2_U3074 , P2_R1215_U65 );
nand NAND2_19639 ( P2_R1215_U492 , P2_U3465 , P2_R1215_U66 );
nand NAND2_19640 ( P2_R1215_U493 , P2_R1215_U492 , P2_R1215_U491 );
nand NAND2_19641 ( P2_R1215_U494 , P2_R1215_U362 , P2_R1215_U94 );
nand NAND2_19642 ( P2_R1215_U495 , P2_R1215_U493 , P2_R1215_U338 );
nand NAND2_19643 ( P2_R1215_U496 , P2_U3065 , P2_R1215_U67 );
nand NAND2_19644 ( P2_R1215_U497 , P2_U3462 , P2_R1215_U68 );
nand NAND2_19645 ( P2_R1215_U498 , P2_R1215_U497 , P2_R1215_U496 );
nand NAND2_19646 ( P2_R1215_U499 , P2_R1215_U363 , P2_R1215_U167 );
nand NAND2_19647 ( P2_R1215_U500 , P2_R1215_U244 , P2_R1215_U498 );
nand NAND2_19648 ( P2_R1215_U501 , P2_U3064 , P2_R1215_U63 );
nand NAND2_19649 ( P2_R1215_U502 , P2_U3459 , P2_R1215_U64 );
nand NAND2_19650 ( P2_R1215_U503 , P2_U3079 , P2_R1215_U30 );
nand NAND2_19651 ( P2_R1215_U504 , P2_U3427 , P2_R1215_U31 );
and AND2_19652 ( P2_R1164_U4 , P2_R1164_U179 , P2_R1164_U178 );
and AND2_19653 ( P2_R1164_U5 , P2_R1164_U197 , P2_R1164_U196 );
and AND2_19654 ( P2_R1164_U6 , P2_R1164_U237 , P2_R1164_U236 );
and AND2_19655 ( P2_R1164_U7 , P2_R1164_U246 , P2_R1164_U245 );
and AND2_19656 ( P2_R1164_U8 , P2_R1164_U264 , P2_R1164_U263 );
and AND2_19657 ( P2_R1164_U9 , P2_R1164_U272 , P2_R1164_U271 );
and AND2_19658 ( P2_R1164_U10 , P2_R1164_U351 , P2_R1164_U348 );
and AND2_19659 ( P2_R1164_U11 , P2_R1164_U344 , P2_R1164_U341 );
and AND2_19660 ( P2_R1164_U12 , P2_R1164_U335 , P2_R1164_U332 );
and AND2_19661 ( P2_R1164_U13 , P2_R1164_U326 , P2_R1164_U323 );
and AND2_19662 ( P2_R1164_U14 , P2_R1164_U320 , P2_R1164_U318 );
and AND2_19663 ( P2_R1164_U15 , P2_R1164_U313 , P2_R1164_U310 );
and AND2_19664 ( P2_R1164_U16 , P2_R1164_U235 , P2_R1164_U232 );
and AND2_19665 ( P2_R1164_U17 , P2_R1164_U227 , P2_R1164_U224 );
and AND2_19666 ( P2_R1164_U18 , P2_R1164_U213 , P2_R1164_U210 );
not NOT1_19667 ( P2_R1164_U19 , P2_U3447 );
not NOT1_19668 ( P2_R1164_U20 , P2_U3073 );
not NOT1_19669 ( P2_R1164_U21 , P2_U3072 );
nand NAND2_19670 ( P2_R1164_U22 , P2_U3073 , P2_U3447 );
not NOT1_19671 ( P2_R1164_U23 , P2_U3450 );
not NOT1_19672 ( P2_R1164_U24 , P2_U3441 );
not NOT1_19673 ( P2_R1164_U25 , P2_U3062 );
not NOT1_19674 ( P2_R1164_U26 , P2_U3069 );
not NOT1_19675 ( P2_R1164_U27 , P2_U3435 );
not NOT1_19676 ( P2_R1164_U28 , P2_U3070 );
not NOT1_19677 ( P2_R1164_U29 , P2_U3427 );
not NOT1_19678 ( P2_R1164_U30 , P2_U3079 );
nand NAND2_19679 ( P2_R1164_U31 , P2_U3079 , P2_U3427 );
not NOT1_19680 ( P2_R1164_U32 , P2_U3438 );
not NOT1_19681 ( P2_R1164_U33 , P2_U3066 );
nand NAND2_19682 ( P2_R1164_U34 , P2_U3062 , P2_U3441 );
not NOT1_19683 ( P2_R1164_U35 , P2_U3444 );
not NOT1_19684 ( P2_R1164_U36 , P2_U3453 );
not NOT1_19685 ( P2_R1164_U37 , P2_U3086 );
not NOT1_19686 ( P2_R1164_U38 , P2_U3085 );
not NOT1_19687 ( P2_R1164_U39 , P2_U3456 );
nand NAND2_19688 ( P2_R1164_U40 , P2_R1164_U61 , P2_R1164_U205 );
nand NAND2_19689 ( P2_R1164_U41 , P2_R1164_U117 , P2_R1164_U193 );
nand NAND2_19690 ( P2_R1164_U42 , P2_R1164_U182 , P2_R1164_U183 );
nand NAND2_19691 ( P2_R1164_U43 , P2_U3432 , P2_U3080 );
nand NAND2_19692 ( P2_R1164_U44 , P2_R1164_U122 , P2_R1164_U219 );
nand NAND2_19693 ( P2_R1164_U45 , P2_R1164_U216 , P2_R1164_U215 );
not NOT1_19694 ( P2_R1164_U46 , P2_U3950 );
not NOT1_19695 ( P2_R1164_U47 , P2_U3055 );
not NOT1_19696 ( P2_R1164_U48 , P2_U3059 );
not NOT1_19697 ( P2_R1164_U49 , P2_U3951 );
not NOT1_19698 ( P2_R1164_U50 , P2_U3952 );
not NOT1_19699 ( P2_R1164_U51 , P2_U3060 );
not NOT1_19700 ( P2_R1164_U52 , P2_U3953 );
not NOT1_19701 ( P2_R1164_U53 , P2_U3067 );
not NOT1_19702 ( P2_R1164_U54 , P2_U3956 );
not NOT1_19703 ( P2_R1164_U55 , P2_U3077 );
not NOT1_19704 ( P2_R1164_U56 , P2_U3477 );
not NOT1_19705 ( P2_R1164_U57 , P2_U3075 );
not NOT1_19706 ( P2_R1164_U58 , P2_U3071 );
nand NAND2_19707 ( P2_R1164_U59 , P2_U3075 , P2_U3477 );
not NOT1_19708 ( P2_R1164_U60 , P2_U3480 );
nand NAND2_19709 ( P2_R1164_U61 , P2_U3086 , P2_U3453 );
not NOT1_19710 ( P2_R1164_U62 , P2_U3459 );
not NOT1_19711 ( P2_R1164_U63 , P2_U3064 );
not NOT1_19712 ( P2_R1164_U64 , P2_U3465 );
not NOT1_19713 ( P2_R1164_U65 , P2_U3074 );
not NOT1_19714 ( P2_R1164_U66 , P2_U3462 );
not NOT1_19715 ( P2_R1164_U67 , P2_U3065 );
nand NAND2_19716 ( P2_R1164_U68 , P2_U3065 , P2_U3462 );
not NOT1_19717 ( P2_R1164_U69 , P2_U3468 );
not NOT1_19718 ( P2_R1164_U70 , P2_U3082 );
not NOT1_19719 ( P2_R1164_U71 , P2_U3471 );
not NOT1_19720 ( P2_R1164_U72 , P2_U3081 );
not NOT1_19721 ( P2_R1164_U73 , P2_U3474 );
not NOT1_19722 ( P2_R1164_U74 , P2_U3076 );
not NOT1_19723 ( P2_R1164_U75 , P2_U3483 );
not NOT1_19724 ( P2_R1164_U76 , P2_U3084 );
nand NAND2_19725 ( P2_R1164_U77 , P2_U3084 , P2_U3483 );
not NOT1_19726 ( P2_R1164_U78 , P2_U3485 );
not NOT1_19727 ( P2_R1164_U79 , P2_U3083 );
nand NAND2_19728 ( P2_R1164_U80 , P2_U3083 , P2_U3485 );
not NOT1_19729 ( P2_R1164_U81 , P2_U3957 );
not NOT1_19730 ( P2_R1164_U82 , P2_U3955 );
not NOT1_19731 ( P2_R1164_U83 , P2_U3063 );
not NOT1_19732 ( P2_R1164_U84 , P2_U3954 );
not NOT1_19733 ( P2_R1164_U85 , P2_U3068 );
nand NAND2_19734 ( P2_R1164_U86 , P2_U3951 , P2_U3059 );
not NOT1_19735 ( P2_R1164_U87 , P2_U3056 );
not NOT1_19736 ( P2_R1164_U88 , P2_U3949 );
nand NAND2_19737 ( P2_R1164_U89 , P2_R1164_U306 , P2_R1164_U176 );
not NOT1_19738 ( P2_R1164_U90 , P2_U3078 );
nand NAND2_19739 ( P2_R1164_U91 , P2_R1164_U77 , P2_R1164_U315 );
nand NAND2_19740 ( P2_R1164_U92 , P2_R1164_U261 , P2_R1164_U260 );
nand NAND2_19741 ( P2_R1164_U93 , P2_R1164_U68 , P2_R1164_U337 );
nand NAND2_19742 ( P2_R1164_U94 , P2_R1164_U457 , P2_R1164_U456 );
nand NAND2_19743 ( P2_R1164_U95 , P2_R1164_U504 , P2_R1164_U503 );
nand NAND2_19744 ( P2_R1164_U96 , P2_R1164_U375 , P2_R1164_U374 );
nand NAND2_19745 ( P2_R1164_U97 , P2_R1164_U380 , P2_R1164_U379 );
nand NAND2_19746 ( P2_R1164_U98 , P2_R1164_U387 , P2_R1164_U386 );
nand NAND2_19747 ( P2_R1164_U99 , P2_R1164_U394 , P2_R1164_U393 );
nand NAND2_19748 ( P2_R1164_U100 , P2_R1164_U399 , P2_R1164_U398 );
nand NAND2_19749 ( P2_R1164_U101 , P2_R1164_U408 , P2_R1164_U407 );
nand NAND2_19750 ( P2_R1164_U102 , P2_R1164_U415 , P2_R1164_U414 );
nand NAND2_19751 ( P2_R1164_U103 , P2_R1164_U422 , P2_R1164_U421 );
nand NAND2_19752 ( P2_R1164_U104 , P2_R1164_U429 , P2_R1164_U428 );
nand NAND2_19753 ( P2_R1164_U105 , P2_R1164_U434 , P2_R1164_U433 );
nand NAND2_19754 ( P2_R1164_U106 , P2_R1164_U441 , P2_R1164_U440 );
nand NAND2_19755 ( P2_R1164_U107 , P2_R1164_U448 , P2_R1164_U447 );
nand NAND2_19756 ( P2_R1164_U108 , P2_R1164_U462 , P2_R1164_U461 );
nand NAND2_19757 ( P2_R1164_U109 , P2_R1164_U467 , P2_R1164_U466 );
nand NAND2_19758 ( P2_R1164_U110 , P2_R1164_U474 , P2_R1164_U473 );
nand NAND2_19759 ( P2_R1164_U111 , P2_R1164_U481 , P2_R1164_U480 );
nand NAND2_19760 ( P2_R1164_U112 , P2_R1164_U488 , P2_R1164_U487 );
nand NAND2_19761 ( P2_R1164_U113 , P2_R1164_U495 , P2_R1164_U494 );
nand NAND2_19762 ( P2_R1164_U114 , P2_R1164_U500 , P2_R1164_U499 );
and AND2_19763 ( P2_R1164_U115 , P2_R1164_U189 , P2_R1164_U187 );
and AND2_19764 ( P2_R1164_U116 , P2_R1164_U4 , P2_R1164_U180 );
and AND2_19765 ( P2_R1164_U117 , P2_R1164_U194 , P2_R1164_U192 );
and AND2_19766 ( P2_R1164_U118 , P2_R1164_U201 , P2_R1164_U200 );
and AND3_19767 ( P2_R1164_U119 , P2_R1164_U382 , P2_R1164_U381 , P2_R1164_U22 );
and AND2_19768 ( P2_R1164_U120 , P2_R1164_U212 , P2_R1164_U5 );
and AND2_19769 ( P2_R1164_U121 , P2_R1164_U181 , P2_R1164_U180 );
and AND2_19770 ( P2_R1164_U122 , P2_R1164_U220 , P2_R1164_U218 );
and AND3_19771 ( P2_R1164_U123 , P2_R1164_U389 , P2_R1164_U388 , P2_R1164_U34 );
and AND2_19772 ( P2_R1164_U124 , P2_R1164_U226 , P2_R1164_U4 );
and AND2_19773 ( P2_R1164_U125 , P2_R1164_U234 , P2_R1164_U181 );
and AND2_19774 ( P2_R1164_U126 , P2_R1164_U204 , P2_R1164_U6 );
and AND2_19775 ( P2_R1164_U127 , P2_R1164_U239 , P2_R1164_U171 );
and AND2_19776 ( P2_R1164_U128 , P2_R1164_U250 , P2_R1164_U7 );
and AND2_19777 ( P2_R1164_U129 , P2_R1164_U248 , P2_R1164_U172 );
and AND2_19778 ( P2_R1164_U130 , P2_R1164_U268 , P2_R1164_U267 );
and AND2_19779 ( P2_R1164_U131 , P2_R1164_U9 , P2_R1164_U282 );
and AND2_19780 ( P2_R1164_U132 , P2_R1164_U285 , P2_R1164_U280 );
and AND2_19781 ( P2_R1164_U133 , P2_R1164_U301 , P2_R1164_U298 );
and AND2_19782 ( P2_R1164_U134 , P2_R1164_U368 , P2_R1164_U302 );
and AND2_19783 ( P2_R1164_U135 , P2_R1164_U160 , P2_R1164_U278 );
and AND3_19784 ( P2_R1164_U136 , P2_R1164_U455 , P2_R1164_U454 , P2_R1164_U80 );
and AND2_19785 ( P2_R1164_U137 , P2_R1164_U325 , P2_R1164_U9 );
and AND3_19786 ( P2_R1164_U138 , P2_R1164_U469 , P2_R1164_U468 , P2_R1164_U59 );
and AND2_19787 ( P2_R1164_U139 , P2_R1164_U334 , P2_R1164_U8 );
and AND3_19788 ( P2_R1164_U140 , P2_R1164_U490 , P2_R1164_U489 , P2_R1164_U172 );
and AND2_19789 ( P2_R1164_U141 , P2_R1164_U343 , P2_R1164_U7 );
and AND3_19790 ( P2_R1164_U142 , P2_R1164_U502 , P2_R1164_U501 , P2_R1164_U171 );
and AND2_19791 ( P2_R1164_U143 , P2_R1164_U350 , P2_R1164_U6 );
nand NAND2_19792 ( P2_R1164_U144 , P2_R1164_U118 , P2_R1164_U202 );
nand NAND2_19793 ( P2_R1164_U145 , P2_R1164_U217 , P2_R1164_U229 );
not NOT1_19794 ( P2_R1164_U146 , P2_U3057 );
not NOT1_19795 ( P2_R1164_U147 , P2_U3960 );
and AND2_19796 ( P2_R1164_U148 , P2_R1164_U403 , P2_R1164_U402 );
nand NAND3_19797 ( P2_R1164_U149 , P2_R1164_U304 , P2_R1164_U169 , P2_R1164_U364 );
and AND2_19798 ( P2_R1164_U150 , P2_R1164_U410 , P2_R1164_U409 );
nand NAND3_19799 ( P2_R1164_U151 , P2_R1164_U370 , P2_R1164_U369 , P2_R1164_U134 );
and AND2_19800 ( P2_R1164_U152 , P2_R1164_U417 , P2_R1164_U416 );
nand NAND3_19801 ( P2_R1164_U153 , P2_R1164_U365 , P2_R1164_U299 , P2_R1164_U86 );
and AND2_19802 ( P2_R1164_U154 , P2_R1164_U424 , P2_R1164_U423 );
nand NAND2_19803 ( P2_R1164_U155 , P2_R1164_U293 , P2_R1164_U292 );
and AND2_19804 ( P2_R1164_U156 , P2_R1164_U436 , P2_R1164_U435 );
nand NAND2_19805 ( P2_R1164_U157 , P2_R1164_U289 , P2_R1164_U288 );
and AND2_19806 ( P2_R1164_U158 , P2_R1164_U443 , P2_R1164_U442 );
nand NAND2_19807 ( P2_R1164_U159 , P2_R1164_U132 , P2_R1164_U284 );
and AND2_19808 ( P2_R1164_U160 , P2_R1164_U450 , P2_R1164_U449 );
nand NAND2_19809 ( P2_R1164_U161 , P2_R1164_U43 , P2_R1164_U327 );
nand NAND2_19810 ( P2_R1164_U162 , P2_R1164_U130 , P2_R1164_U269 );
and AND2_19811 ( P2_R1164_U163 , P2_R1164_U476 , P2_R1164_U475 );
nand NAND2_19812 ( P2_R1164_U164 , P2_R1164_U257 , P2_R1164_U256 );
and AND2_19813 ( P2_R1164_U165 , P2_R1164_U483 , P2_R1164_U482 );
nand NAND2_19814 ( P2_R1164_U166 , P2_R1164_U253 , P2_R1164_U252 );
nand NAND2_19815 ( P2_R1164_U167 , P2_R1164_U243 , P2_R1164_U242 );
nand NAND2_19816 ( P2_R1164_U168 , P2_R1164_U367 , P2_R1164_U366 );
nand NAND2_19817 ( P2_R1164_U169 , P2_U3056 , P2_R1164_U151 );
not NOT1_19818 ( P2_R1164_U170 , P2_R1164_U34 );
nand NAND2_19819 ( P2_R1164_U171 , P2_U3456 , P2_U3085 );
nand NAND2_19820 ( P2_R1164_U172 , P2_U3074 , P2_U3465 );
nand NAND2_19821 ( P2_R1164_U173 , P2_U3060 , P2_U3952 );
not NOT1_19822 ( P2_R1164_U174 , P2_R1164_U68 );
not NOT1_19823 ( P2_R1164_U175 , P2_R1164_U77 );
nand NAND2_19824 ( P2_R1164_U176 , P2_U3067 , P2_U3953 );
not NOT1_19825 ( P2_R1164_U177 , P2_R1164_U61 );
or OR2_19826 ( P2_R1164_U178 , P2_U3069 , P2_U3444 );
or OR2_19827 ( P2_R1164_U179 , P2_U3062 , P2_U3441 );
or OR2_19828 ( P2_R1164_U180 , P2_U3438 , P2_U3066 );
or OR2_19829 ( P2_R1164_U181 , P2_U3435 , P2_U3070 );
not NOT1_19830 ( P2_R1164_U182 , P2_R1164_U31 );
or OR2_19831 ( P2_R1164_U183 , P2_U3432 , P2_U3080 );
not NOT1_19832 ( P2_R1164_U184 , P2_R1164_U42 );
not NOT1_19833 ( P2_R1164_U185 , P2_R1164_U43 );
nand NAND2_19834 ( P2_R1164_U186 , P2_R1164_U42 , P2_R1164_U43 );
nand NAND2_19835 ( P2_R1164_U187 , P2_U3070 , P2_U3435 );
nand NAND2_19836 ( P2_R1164_U188 , P2_R1164_U186 , P2_R1164_U181 );
nand NAND2_19837 ( P2_R1164_U189 , P2_U3066 , P2_U3438 );
nand NAND2_19838 ( P2_R1164_U190 , P2_R1164_U115 , P2_R1164_U188 );
nand NAND2_19839 ( P2_R1164_U191 , P2_R1164_U35 , P2_R1164_U34 );
nand NAND2_19840 ( P2_R1164_U192 , P2_U3069 , P2_R1164_U191 );
nand NAND2_19841 ( P2_R1164_U193 , P2_R1164_U116 , P2_R1164_U190 );
nand NAND2_19842 ( P2_R1164_U194 , P2_U3444 , P2_R1164_U170 );
not NOT1_19843 ( P2_R1164_U195 , P2_R1164_U41 );
or OR2_19844 ( P2_R1164_U196 , P2_U3072 , P2_U3450 );
or OR2_19845 ( P2_R1164_U197 , P2_U3073 , P2_U3447 );
not NOT1_19846 ( P2_R1164_U198 , P2_R1164_U22 );
nand NAND2_19847 ( P2_R1164_U199 , P2_R1164_U23 , P2_R1164_U22 );
nand NAND2_19848 ( P2_R1164_U200 , P2_U3072 , P2_R1164_U199 );
nand NAND2_19849 ( P2_R1164_U201 , P2_U3450 , P2_R1164_U198 );
nand NAND2_19850 ( P2_R1164_U202 , P2_R1164_U5 , P2_R1164_U41 );
not NOT1_19851 ( P2_R1164_U203 , P2_R1164_U144 );
or OR2_19852 ( P2_R1164_U204 , P2_U3453 , P2_U3086 );
nand NAND2_19853 ( P2_R1164_U205 , P2_R1164_U204 , P2_R1164_U144 );
not NOT1_19854 ( P2_R1164_U206 , P2_R1164_U40 );
or OR2_19855 ( P2_R1164_U207 , P2_U3085 , P2_U3456 );
or OR2_19856 ( P2_R1164_U208 , P2_U3447 , P2_U3073 );
nand NAND2_19857 ( P2_R1164_U209 , P2_R1164_U208 , P2_R1164_U41 );
nand NAND2_19858 ( P2_R1164_U210 , P2_R1164_U119 , P2_R1164_U209 );
nand NAND2_19859 ( P2_R1164_U211 , P2_R1164_U195 , P2_R1164_U22 );
nand NAND2_19860 ( P2_R1164_U212 , P2_U3450 , P2_U3072 );
nand NAND2_19861 ( P2_R1164_U213 , P2_R1164_U120 , P2_R1164_U211 );
or OR2_19862 ( P2_R1164_U214 , P2_U3073 , P2_U3447 );
nand NAND2_19863 ( P2_R1164_U215 , P2_R1164_U185 , P2_R1164_U181 );
nand NAND2_19864 ( P2_R1164_U216 , P2_U3070 , P2_U3435 );
not NOT1_19865 ( P2_R1164_U217 , P2_R1164_U45 );
nand NAND2_19866 ( P2_R1164_U218 , P2_R1164_U121 , P2_R1164_U184 );
nand NAND2_19867 ( P2_R1164_U219 , P2_R1164_U45 , P2_R1164_U180 );
nand NAND2_19868 ( P2_R1164_U220 , P2_U3066 , P2_U3438 );
not NOT1_19869 ( P2_R1164_U221 , P2_R1164_U44 );
or OR2_19870 ( P2_R1164_U222 , P2_U3441 , P2_U3062 );
nand NAND2_19871 ( P2_R1164_U223 , P2_R1164_U222 , P2_R1164_U44 );
nand NAND2_19872 ( P2_R1164_U224 , P2_R1164_U123 , P2_R1164_U223 );
nand NAND2_19873 ( P2_R1164_U225 , P2_R1164_U221 , P2_R1164_U34 );
nand NAND2_19874 ( P2_R1164_U226 , P2_U3444 , P2_U3069 );
nand NAND2_19875 ( P2_R1164_U227 , P2_R1164_U124 , P2_R1164_U225 );
or OR2_19876 ( P2_R1164_U228 , P2_U3062 , P2_U3441 );
nand NAND2_19877 ( P2_R1164_U229 , P2_R1164_U184 , P2_R1164_U181 );
not NOT1_19878 ( P2_R1164_U230 , P2_R1164_U145 );
nand NAND2_19879 ( P2_R1164_U231 , P2_U3066 , P2_U3438 );
nand NAND4_19880 ( P2_R1164_U232 , P2_R1164_U401 , P2_R1164_U400 , P2_R1164_U43 , P2_R1164_U42 );
nand NAND2_19881 ( P2_R1164_U233 , P2_R1164_U43 , P2_R1164_U42 );
nand NAND2_19882 ( P2_R1164_U234 , P2_U3070 , P2_U3435 );
nand NAND2_19883 ( P2_R1164_U235 , P2_R1164_U125 , P2_R1164_U233 );
or OR2_19884 ( P2_R1164_U236 , P2_U3085 , P2_U3456 );
or OR2_19885 ( P2_R1164_U237 , P2_U3064 , P2_U3459 );
nand NAND2_19886 ( P2_R1164_U238 , P2_R1164_U177 , P2_R1164_U6 );
nand NAND2_19887 ( P2_R1164_U239 , P2_U3064 , P2_U3459 );
nand NAND2_19888 ( P2_R1164_U240 , P2_R1164_U127 , P2_R1164_U238 );
or OR2_19889 ( P2_R1164_U241 , P2_U3459 , P2_U3064 );
nand NAND2_19890 ( P2_R1164_U242 , P2_R1164_U126 , P2_R1164_U144 );
nand NAND2_19891 ( P2_R1164_U243 , P2_R1164_U241 , P2_R1164_U240 );
not NOT1_19892 ( P2_R1164_U244 , P2_R1164_U167 );
or OR2_19893 ( P2_R1164_U245 , P2_U3082 , P2_U3468 );
or OR2_19894 ( P2_R1164_U246 , P2_U3074 , P2_U3465 );
nand NAND2_19895 ( P2_R1164_U247 , P2_R1164_U174 , P2_R1164_U7 );
nand NAND2_19896 ( P2_R1164_U248 , P2_U3082 , P2_U3468 );
nand NAND2_19897 ( P2_R1164_U249 , P2_R1164_U129 , P2_R1164_U247 );
or OR2_19898 ( P2_R1164_U250 , P2_U3462 , P2_U3065 );
or OR2_19899 ( P2_R1164_U251 , P2_U3468 , P2_U3082 );
nand NAND2_19900 ( P2_R1164_U252 , P2_R1164_U128 , P2_R1164_U167 );
nand NAND2_19901 ( P2_R1164_U253 , P2_R1164_U251 , P2_R1164_U249 );
not NOT1_19902 ( P2_R1164_U254 , P2_R1164_U166 );
or OR2_19903 ( P2_R1164_U255 , P2_U3471 , P2_U3081 );
nand NAND2_19904 ( P2_R1164_U256 , P2_R1164_U255 , P2_R1164_U166 );
nand NAND2_19905 ( P2_R1164_U257 , P2_U3081 , P2_U3471 );
not NOT1_19906 ( P2_R1164_U258 , P2_R1164_U164 );
or OR2_19907 ( P2_R1164_U259 , P2_U3474 , P2_U3076 );
nand NAND2_19908 ( P2_R1164_U260 , P2_R1164_U259 , P2_R1164_U164 );
nand NAND2_19909 ( P2_R1164_U261 , P2_U3076 , P2_U3474 );
not NOT1_19910 ( P2_R1164_U262 , P2_R1164_U92 );
or OR2_19911 ( P2_R1164_U263 , P2_U3071 , P2_U3480 );
or OR2_19912 ( P2_R1164_U264 , P2_U3075 , P2_U3477 );
not NOT1_19913 ( P2_R1164_U265 , P2_R1164_U59 );
nand NAND2_19914 ( P2_R1164_U266 , P2_R1164_U60 , P2_R1164_U59 );
nand NAND2_19915 ( P2_R1164_U267 , P2_U3071 , P2_R1164_U266 );
nand NAND2_19916 ( P2_R1164_U268 , P2_U3480 , P2_R1164_U265 );
nand NAND2_19917 ( P2_R1164_U269 , P2_R1164_U8 , P2_R1164_U92 );
not NOT1_19918 ( P2_R1164_U270 , P2_R1164_U162 );
or OR2_19919 ( P2_R1164_U271 , P2_U3078 , P2_U3957 );
or OR2_19920 ( P2_R1164_U272 , P2_U3083 , P2_U3485 );
or OR2_19921 ( P2_R1164_U273 , P2_U3077 , P2_U3956 );
not NOT1_19922 ( P2_R1164_U274 , P2_R1164_U80 );
nand NAND2_19923 ( P2_R1164_U275 , P2_U3957 , P2_R1164_U274 );
nand NAND2_19924 ( P2_R1164_U276 , P2_R1164_U275 , P2_R1164_U90 );
nand NAND2_19925 ( P2_R1164_U277 , P2_R1164_U80 , P2_R1164_U81 );
nand NAND2_19926 ( P2_R1164_U278 , P2_R1164_U277 , P2_R1164_U276 );
nand NAND2_19927 ( P2_R1164_U279 , P2_R1164_U175 , P2_R1164_U9 );
nand NAND2_19928 ( P2_R1164_U280 , P2_U3077 , P2_U3956 );
nand NAND2_19929 ( P2_R1164_U281 , P2_R1164_U278 , P2_R1164_U279 );
or OR2_19930 ( P2_R1164_U282 , P2_U3483 , P2_U3084 );
or OR2_19931 ( P2_R1164_U283 , P2_U3956 , P2_U3077 );
nand NAND3_19932 ( P2_R1164_U284 , P2_R1164_U273 , P2_R1164_U162 , P2_R1164_U131 );
nand NAND2_19933 ( P2_R1164_U285 , P2_R1164_U283 , P2_R1164_U281 );
not NOT1_19934 ( P2_R1164_U286 , P2_R1164_U159 );
or OR2_19935 ( P2_R1164_U287 , P2_U3955 , P2_U3063 );
nand NAND2_19936 ( P2_R1164_U288 , P2_R1164_U287 , P2_R1164_U159 );
nand NAND2_19937 ( P2_R1164_U289 , P2_U3063 , P2_U3955 );
not NOT1_19938 ( P2_R1164_U290 , P2_R1164_U157 );
or OR2_19939 ( P2_R1164_U291 , P2_U3954 , P2_U3068 );
nand NAND2_19940 ( P2_R1164_U292 , P2_R1164_U291 , P2_R1164_U157 );
nand NAND2_19941 ( P2_R1164_U293 , P2_U3068 , P2_U3954 );
not NOT1_19942 ( P2_R1164_U294 , P2_R1164_U155 );
or OR2_19943 ( P2_R1164_U295 , P2_U3060 , P2_U3952 );
nand NAND2_19944 ( P2_R1164_U296 , P2_R1164_U176 , P2_R1164_U173 );
not NOT1_19945 ( P2_R1164_U297 , P2_R1164_U86 );
or OR2_19946 ( P2_R1164_U298 , P2_U3953 , P2_U3067 );
nand NAND3_19947 ( P2_R1164_U299 , P2_R1164_U155 , P2_R1164_U298 , P2_R1164_U168 );
not NOT1_19948 ( P2_R1164_U300 , P2_R1164_U153 );
or OR2_19949 ( P2_R1164_U301 , P2_U3950 , P2_U3055 );
nand NAND2_19950 ( P2_R1164_U302 , P2_U3055 , P2_U3950 );
not NOT1_19951 ( P2_R1164_U303 , P2_R1164_U151 );
nand NAND2_19952 ( P2_R1164_U304 , P2_U3949 , P2_R1164_U151 );
not NOT1_19953 ( P2_R1164_U305 , P2_R1164_U149 );
nand NAND2_19954 ( P2_R1164_U306 , P2_R1164_U298 , P2_R1164_U155 );
not NOT1_19955 ( P2_R1164_U307 , P2_R1164_U89 );
or OR2_19956 ( P2_R1164_U308 , P2_U3952 , P2_U3060 );
nand NAND2_19957 ( P2_R1164_U309 , P2_R1164_U308 , P2_R1164_U89 );
nand NAND3_19958 ( P2_R1164_U310 , P2_R1164_U309 , P2_R1164_U173 , P2_R1164_U154 );
nand NAND2_19959 ( P2_R1164_U311 , P2_R1164_U307 , P2_R1164_U173 );
nand NAND2_19960 ( P2_R1164_U312 , P2_U3951 , P2_U3059 );
nand NAND3_19961 ( P2_R1164_U313 , P2_R1164_U311 , P2_R1164_U312 , P2_R1164_U168 );
or OR2_19962 ( P2_R1164_U314 , P2_U3060 , P2_U3952 );
nand NAND2_19963 ( P2_R1164_U315 , P2_R1164_U282 , P2_R1164_U162 );
not NOT1_19964 ( P2_R1164_U316 , P2_R1164_U91 );
nand NAND2_19965 ( P2_R1164_U317 , P2_R1164_U9 , P2_R1164_U91 );
nand NAND2_19966 ( P2_R1164_U318 , P2_R1164_U135 , P2_R1164_U317 );
nand NAND2_19967 ( P2_R1164_U319 , P2_R1164_U317 , P2_R1164_U278 );
nand NAND2_19968 ( P2_R1164_U320 , P2_R1164_U453 , P2_R1164_U319 );
or OR2_19969 ( P2_R1164_U321 , P2_U3485 , P2_U3083 );
nand NAND2_19970 ( P2_R1164_U322 , P2_R1164_U321 , P2_R1164_U91 );
nand NAND2_19971 ( P2_R1164_U323 , P2_R1164_U136 , P2_R1164_U322 );
nand NAND2_19972 ( P2_R1164_U324 , P2_R1164_U316 , P2_R1164_U80 );
nand NAND2_19973 ( P2_R1164_U325 , P2_U3078 , P2_U3957 );
nand NAND2_19974 ( P2_R1164_U326 , P2_R1164_U137 , P2_R1164_U324 );
or OR2_19975 ( P2_R1164_U327 , P2_U3432 , P2_U3080 );
not NOT1_19976 ( P2_R1164_U328 , P2_R1164_U161 );
or OR2_19977 ( P2_R1164_U329 , P2_U3083 , P2_U3485 );
or OR2_19978 ( P2_R1164_U330 , P2_U3477 , P2_U3075 );
nand NAND2_19979 ( P2_R1164_U331 , P2_R1164_U330 , P2_R1164_U92 );
nand NAND2_19980 ( P2_R1164_U332 , P2_R1164_U138 , P2_R1164_U331 );
nand NAND2_19981 ( P2_R1164_U333 , P2_R1164_U262 , P2_R1164_U59 );
nand NAND2_19982 ( P2_R1164_U334 , P2_U3480 , P2_U3071 );
nand NAND2_19983 ( P2_R1164_U335 , P2_R1164_U139 , P2_R1164_U333 );
or OR2_19984 ( P2_R1164_U336 , P2_U3075 , P2_U3477 );
nand NAND2_19985 ( P2_R1164_U337 , P2_R1164_U250 , P2_R1164_U167 );
not NOT1_19986 ( P2_R1164_U338 , P2_R1164_U93 );
or OR2_19987 ( P2_R1164_U339 , P2_U3465 , P2_U3074 );
nand NAND2_19988 ( P2_R1164_U340 , P2_R1164_U339 , P2_R1164_U93 );
nand NAND2_19989 ( P2_R1164_U341 , P2_R1164_U140 , P2_R1164_U340 );
nand NAND2_19990 ( P2_R1164_U342 , P2_R1164_U338 , P2_R1164_U172 );
nand NAND2_19991 ( P2_R1164_U343 , P2_U3082 , P2_U3468 );
nand NAND2_19992 ( P2_R1164_U344 , P2_R1164_U141 , P2_R1164_U342 );
or OR2_19993 ( P2_R1164_U345 , P2_U3074 , P2_U3465 );
or OR2_19994 ( P2_R1164_U346 , P2_U3456 , P2_U3085 );
nand NAND2_19995 ( P2_R1164_U347 , P2_R1164_U346 , P2_R1164_U40 );
nand NAND2_19996 ( P2_R1164_U348 , P2_R1164_U142 , P2_R1164_U347 );
nand NAND2_19997 ( P2_R1164_U349 , P2_R1164_U206 , P2_R1164_U171 );
nand NAND2_19998 ( P2_R1164_U350 , P2_U3064 , P2_U3459 );
nand NAND2_19999 ( P2_R1164_U351 , P2_R1164_U143 , P2_R1164_U349 );
nand NAND2_20000 ( P2_R1164_U352 , P2_R1164_U207 , P2_R1164_U171 );
nand NAND2_20001 ( P2_R1164_U353 , P2_R1164_U204 , P2_R1164_U61 );
nand NAND2_20002 ( P2_R1164_U354 , P2_R1164_U214 , P2_R1164_U22 );
nand NAND2_20003 ( P2_R1164_U355 , P2_R1164_U228 , P2_R1164_U34 );
nand NAND2_20004 ( P2_R1164_U356 , P2_R1164_U231 , P2_R1164_U180 );
nand NAND2_20005 ( P2_R1164_U357 , P2_R1164_U314 , P2_R1164_U173 );
nand NAND2_20006 ( P2_R1164_U358 , P2_R1164_U298 , P2_R1164_U176 );
nand NAND2_20007 ( P2_R1164_U359 , P2_R1164_U329 , P2_R1164_U80 );
nand NAND2_20008 ( P2_R1164_U360 , P2_R1164_U282 , P2_R1164_U77 );
nand NAND2_20009 ( P2_R1164_U361 , P2_R1164_U336 , P2_R1164_U59 );
nand NAND2_20010 ( P2_R1164_U362 , P2_R1164_U345 , P2_R1164_U172 );
nand NAND2_20011 ( P2_R1164_U363 , P2_R1164_U250 , P2_R1164_U68 );
nand NAND2_20012 ( P2_R1164_U364 , P2_U3949 , P2_U3056 );
nand NAND2_20013 ( P2_R1164_U365 , P2_R1164_U296 , P2_R1164_U168 );
nand NAND2_20014 ( P2_R1164_U366 , P2_U3059 , P2_R1164_U295 );
nand NAND2_20015 ( P2_R1164_U367 , P2_U3951 , P2_R1164_U295 );
nand NAND3_20016 ( P2_R1164_U368 , P2_R1164_U296 , P2_R1164_U168 , P2_R1164_U301 );
nand NAND3_20017 ( P2_R1164_U369 , P2_R1164_U155 , P2_R1164_U168 , P2_R1164_U133 );
nand NAND2_20018 ( P2_R1164_U370 , P2_R1164_U297 , P2_R1164_U301 );
nand NAND2_20019 ( P2_R1164_U371 , P2_U3085 , P2_R1164_U39 );
nand NAND2_20020 ( P2_R1164_U372 , P2_U3456 , P2_R1164_U38 );
nand NAND2_20021 ( P2_R1164_U373 , P2_R1164_U372 , P2_R1164_U371 );
nand NAND2_20022 ( P2_R1164_U374 , P2_R1164_U352 , P2_R1164_U40 );
nand NAND2_20023 ( P2_R1164_U375 , P2_R1164_U373 , P2_R1164_U206 );
nand NAND2_20024 ( P2_R1164_U376 , P2_U3086 , P2_R1164_U36 );
nand NAND2_20025 ( P2_R1164_U377 , P2_U3453 , P2_R1164_U37 );
nand NAND2_20026 ( P2_R1164_U378 , P2_R1164_U377 , P2_R1164_U376 );
nand NAND2_20027 ( P2_R1164_U379 , P2_R1164_U353 , P2_R1164_U144 );
nand NAND2_20028 ( P2_R1164_U380 , P2_R1164_U203 , P2_R1164_U378 );
nand NAND2_20029 ( P2_R1164_U381 , P2_U3072 , P2_R1164_U23 );
nand NAND2_20030 ( P2_R1164_U382 , P2_U3450 , P2_R1164_U21 );
nand NAND2_20031 ( P2_R1164_U383 , P2_U3073 , P2_R1164_U19 );
nand NAND2_20032 ( P2_R1164_U384 , P2_U3447 , P2_R1164_U20 );
nand NAND2_20033 ( P2_R1164_U385 , P2_R1164_U384 , P2_R1164_U383 );
nand NAND2_20034 ( P2_R1164_U386 , P2_R1164_U354 , P2_R1164_U41 );
nand NAND2_20035 ( P2_R1164_U387 , P2_R1164_U385 , P2_R1164_U195 );
nand NAND2_20036 ( P2_R1164_U388 , P2_U3069 , P2_R1164_U35 );
nand NAND2_20037 ( P2_R1164_U389 , P2_U3444 , P2_R1164_U26 );
nand NAND2_20038 ( P2_R1164_U390 , P2_U3062 , P2_R1164_U24 );
nand NAND2_20039 ( P2_R1164_U391 , P2_U3441 , P2_R1164_U25 );
nand NAND2_20040 ( P2_R1164_U392 , P2_R1164_U391 , P2_R1164_U390 );
nand NAND2_20041 ( P2_R1164_U393 , P2_R1164_U355 , P2_R1164_U44 );
nand NAND2_20042 ( P2_R1164_U394 , P2_R1164_U392 , P2_R1164_U221 );
nand NAND2_20043 ( P2_R1164_U395 , P2_U3066 , P2_R1164_U32 );
nand NAND2_20044 ( P2_R1164_U396 , P2_U3438 , P2_R1164_U33 );
nand NAND2_20045 ( P2_R1164_U397 , P2_R1164_U396 , P2_R1164_U395 );
nand NAND2_20046 ( P2_R1164_U398 , P2_R1164_U356 , P2_R1164_U145 );
nand NAND2_20047 ( P2_R1164_U399 , P2_R1164_U230 , P2_R1164_U397 );
nand NAND2_20048 ( P2_R1164_U400 , P2_U3070 , P2_R1164_U27 );
nand NAND2_20049 ( P2_R1164_U401 , P2_U3435 , P2_R1164_U28 );
nand NAND2_20050 ( P2_R1164_U402 , P2_U3057 , P2_R1164_U147 );
nand NAND2_20051 ( P2_R1164_U403 , P2_U3960 , P2_R1164_U146 );
nand NAND2_20052 ( P2_R1164_U404 , P2_U3057 , P2_R1164_U147 );
nand NAND2_20053 ( P2_R1164_U405 , P2_U3960 , P2_R1164_U146 );
nand NAND2_20054 ( P2_R1164_U406 , P2_R1164_U405 , P2_R1164_U404 );
nand NAND2_20055 ( P2_R1164_U407 , P2_R1164_U148 , P2_R1164_U149 );
nand NAND2_20056 ( P2_R1164_U408 , P2_R1164_U305 , P2_R1164_U406 );
nand NAND2_20057 ( P2_R1164_U409 , P2_U3056 , P2_R1164_U88 );
nand NAND2_20058 ( P2_R1164_U410 , P2_U3949 , P2_R1164_U87 );
nand NAND2_20059 ( P2_R1164_U411 , P2_U3056 , P2_R1164_U88 );
nand NAND2_20060 ( P2_R1164_U412 , P2_U3949 , P2_R1164_U87 );
nand NAND2_20061 ( P2_R1164_U413 , P2_R1164_U412 , P2_R1164_U411 );
nand NAND2_20062 ( P2_R1164_U414 , P2_R1164_U150 , P2_R1164_U151 );
nand NAND2_20063 ( P2_R1164_U415 , P2_R1164_U303 , P2_R1164_U413 );
nand NAND2_20064 ( P2_R1164_U416 , P2_U3055 , P2_R1164_U46 );
nand NAND2_20065 ( P2_R1164_U417 , P2_U3950 , P2_R1164_U47 );
nand NAND2_20066 ( P2_R1164_U418 , P2_U3055 , P2_R1164_U46 );
nand NAND2_20067 ( P2_R1164_U419 , P2_U3950 , P2_R1164_U47 );
nand NAND2_20068 ( P2_R1164_U420 , P2_R1164_U419 , P2_R1164_U418 );
nand NAND2_20069 ( P2_R1164_U421 , P2_R1164_U152 , P2_R1164_U153 );
nand NAND2_20070 ( P2_R1164_U422 , P2_R1164_U300 , P2_R1164_U420 );
nand NAND2_20071 ( P2_R1164_U423 , P2_U3059 , P2_R1164_U49 );
nand NAND2_20072 ( P2_R1164_U424 , P2_U3951 , P2_R1164_U48 );
nand NAND2_20073 ( P2_R1164_U425 , P2_U3060 , P2_R1164_U50 );
nand NAND2_20074 ( P2_R1164_U426 , P2_U3952 , P2_R1164_U51 );
nand NAND2_20075 ( P2_R1164_U427 , P2_R1164_U426 , P2_R1164_U425 );
nand NAND2_20076 ( P2_R1164_U428 , P2_R1164_U357 , P2_R1164_U89 );
nand NAND2_20077 ( P2_R1164_U429 , P2_R1164_U427 , P2_R1164_U307 );
nand NAND2_20078 ( P2_R1164_U430 , P2_U3067 , P2_R1164_U52 );
nand NAND2_20079 ( P2_R1164_U431 , P2_U3953 , P2_R1164_U53 );
nand NAND2_20080 ( P2_R1164_U432 , P2_R1164_U431 , P2_R1164_U430 );
nand NAND2_20081 ( P2_R1164_U433 , P2_R1164_U358 , P2_R1164_U155 );
nand NAND2_20082 ( P2_R1164_U434 , P2_R1164_U294 , P2_R1164_U432 );
nand NAND2_20083 ( P2_R1164_U435 , P2_U3068 , P2_R1164_U84 );
nand NAND2_20084 ( P2_R1164_U436 , P2_U3954 , P2_R1164_U85 );
nand NAND2_20085 ( P2_R1164_U437 , P2_U3068 , P2_R1164_U84 );
nand NAND2_20086 ( P2_R1164_U438 , P2_U3954 , P2_R1164_U85 );
nand NAND2_20087 ( P2_R1164_U439 , P2_R1164_U438 , P2_R1164_U437 );
nand NAND2_20088 ( P2_R1164_U440 , P2_R1164_U156 , P2_R1164_U157 );
nand NAND2_20089 ( P2_R1164_U441 , P2_R1164_U290 , P2_R1164_U439 );
nand NAND2_20090 ( P2_R1164_U442 , P2_U3063 , P2_R1164_U82 );
nand NAND2_20091 ( P2_R1164_U443 , P2_U3955 , P2_R1164_U83 );
nand NAND2_20092 ( P2_R1164_U444 , P2_U3063 , P2_R1164_U82 );
nand NAND2_20093 ( P2_R1164_U445 , P2_U3955 , P2_R1164_U83 );
nand NAND2_20094 ( P2_R1164_U446 , P2_R1164_U445 , P2_R1164_U444 );
nand NAND2_20095 ( P2_R1164_U447 , P2_R1164_U158 , P2_R1164_U159 );
nand NAND2_20096 ( P2_R1164_U448 , P2_R1164_U286 , P2_R1164_U446 );
nand NAND2_20097 ( P2_R1164_U449 , P2_U3077 , P2_R1164_U54 );
nand NAND2_20098 ( P2_R1164_U450 , P2_U3956 , P2_R1164_U55 );
nand NAND2_20099 ( P2_R1164_U451 , P2_U3077 , P2_R1164_U54 );
nand NAND2_20100 ( P2_R1164_U452 , P2_U3956 , P2_R1164_U55 );
nand NAND2_20101 ( P2_R1164_U453 , P2_R1164_U452 , P2_R1164_U451 );
nand NAND2_20102 ( P2_R1164_U454 , P2_U3078 , P2_R1164_U81 );
nand NAND2_20103 ( P2_R1164_U455 , P2_U3957 , P2_R1164_U90 );
nand NAND2_20104 ( P2_R1164_U456 , P2_R1164_U182 , P2_R1164_U161 );
nand NAND2_20105 ( P2_R1164_U457 , P2_R1164_U328 , P2_R1164_U31 );
nand NAND2_20106 ( P2_R1164_U458 , P2_U3083 , P2_R1164_U78 );
nand NAND2_20107 ( P2_R1164_U459 , P2_U3485 , P2_R1164_U79 );
nand NAND2_20108 ( P2_R1164_U460 , P2_R1164_U459 , P2_R1164_U458 );
nand NAND2_20109 ( P2_R1164_U461 , P2_R1164_U359 , P2_R1164_U91 );
nand NAND2_20110 ( P2_R1164_U462 , P2_R1164_U460 , P2_R1164_U316 );
nand NAND2_20111 ( P2_R1164_U463 , P2_U3084 , P2_R1164_U75 );
nand NAND2_20112 ( P2_R1164_U464 , P2_U3483 , P2_R1164_U76 );
nand NAND2_20113 ( P2_R1164_U465 , P2_R1164_U464 , P2_R1164_U463 );
nand NAND2_20114 ( P2_R1164_U466 , P2_R1164_U360 , P2_R1164_U162 );
nand NAND2_20115 ( P2_R1164_U467 , P2_R1164_U270 , P2_R1164_U465 );
nand NAND2_20116 ( P2_R1164_U468 , P2_U3071 , P2_R1164_U60 );
nand NAND2_20117 ( P2_R1164_U469 , P2_U3480 , P2_R1164_U58 );
nand NAND2_20118 ( P2_R1164_U470 , P2_U3075 , P2_R1164_U56 );
nand NAND2_20119 ( P2_R1164_U471 , P2_U3477 , P2_R1164_U57 );
nand NAND2_20120 ( P2_R1164_U472 , P2_R1164_U471 , P2_R1164_U470 );
nand NAND2_20121 ( P2_R1164_U473 , P2_R1164_U361 , P2_R1164_U92 );
nand NAND2_20122 ( P2_R1164_U474 , P2_R1164_U472 , P2_R1164_U262 );
nand NAND2_20123 ( P2_R1164_U475 , P2_U3076 , P2_R1164_U73 );
nand NAND2_20124 ( P2_R1164_U476 , P2_U3474 , P2_R1164_U74 );
nand NAND2_20125 ( P2_R1164_U477 , P2_U3076 , P2_R1164_U73 );
nand NAND2_20126 ( P2_R1164_U478 , P2_U3474 , P2_R1164_U74 );
nand NAND2_20127 ( P2_R1164_U479 , P2_R1164_U478 , P2_R1164_U477 );
nand NAND2_20128 ( P2_R1164_U480 , P2_R1164_U163 , P2_R1164_U164 );
nand NAND2_20129 ( P2_R1164_U481 , P2_R1164_U258 , P2_R1164_U479 );
nand NAND2_20130 ( P2_R1164_U482 , P2_U3081 , P2_R1164_U71 );
nand NAND2_20131 ( P2_R1164_U483 , P2_U3471 , P2_R1164_U72 );
nand NAND2_20132 ( P2_R1164_U484 , P2_U3081 , P2_R1164_U71 );
nand NAND2_20133 ( P2_R1164_U485 , P2_U3471 , P2_R1164_U72 );
nand NAND2_20134 ( P2_R1164_U486 , P2_R1164_U485 , P2_R1164_U484 );
nand NAND2_20135 ( P2_R1164_U487 , P2_R1164_U165 , P2_R1164_U166 );
nand NAND2_20136 ( P2_R1164_U488 , P2_R1164_U254 , P2_R1164_U486 );
nand NAND2_20137 ( P2_R1164_U489 , P2_U3082 , P2_R1164_U69 );
nand NAND2_20138 ( P2_R1164_U490 , P2_U3468 , P2_R1164_U70 );
nand NAND2_20139 ( P2_R1164_U491 , P2_U3074 , P2_R1164_U64 );
nand NAND2_20140 ( P2_R1164_U492 , P2_U3465 , P2_R1164_U65 );
nand NAND2_20141 ( P2_R1164_U493 , P2_R1164_U492 , P2_R1164_U491 );
nand NAND2_20142 ( P2_R1164_U494 , P2_R1164_U362 , P2_R1164_U93 );
nand NAND2_20143 ( P2_R1164_U495 , P2_R1164_U493 , P2_R1164_U338 );
nand NAND2_20144 ( P2_R1164_U496 , P2_U3065 , P2_R1164_U66 );
nand NAND2_20145 ( P2_R1164_U497 , P2_U3462 , P2_R1164_U67 );
nand NAND2_20146 ( P2_R1164_U498 , P2_R1164_U497 , P2_R1164_U496 );
nand NAND2_20147 ( P2_R1164_U499 , P2_R1164_U363 , P2_R1164_U167 );
nand NAND2_20148 ( P2_R1164_U500 , P2_R1164_U244 , P2_R1164_U498 );
nand NAND2_20149 ( P2_R1164_U501 , P2_U3064 , P2_R1164_U62 );
nand NAND2_20150 ( P2_R1164_U502 , P2_U3459 , P2_R1164_U63 );
nand NAND2_20151 ( P2_R1164_U503 , P2_U3079 , P2_R1164_U29 );
nand NAND2_20152 ( P2_R1164_U504 , P2_U3427 , P2_R1164_U30 );
and AND2_20153 ( P2_R1233_U4 , P2_R1233_U179 , P2_R1233_U178 );
and AND2_20154 ( P2_R1233_U5 , P2_R1233_U197 , P2_R1233_U196 );
and AND2_20155 ( P2_R1233_U6 , P2_R1233_U237 , P2_R1233_U236 );
and AND2_20156 ( P2_R1233_U7 , P2_R1233_U246 , P2_R1233_U245 );
and AND2_20157 ( P2_R1233_U8 , P2_R1233_U264 , P2_R1233_U263 );
and AND2_20158 ( P2_R1233_U9 , P2_R1233_U272 , P2_R1233_U271 );
and AND2_20159 ( P2_R1233_U10 , P2_R1233_U351 , P2_R1233_U348 );
and AND2_20160 ( P2_R1233_U11 , P2_R1233_U344 , P2_R1233_U341 );
and AND2_20161 ( P2_R1233_U12 , P2_R1233_U335 , P2_R1233_U332 );
and AND2_20162 ( P2_R1233_U13 , P2_R1233_U326 , P2_R1233_U323 );
and AND2_20163 ( P2_R1233_U14 , P2_R1233_U320 , P2_R1233_U318 );
and AND2_20164 ( P2_R1233_U15 , P2_R1233_U313 , P2_R1233_U310 );
and AND2_20165 ( P2_R1233_U16 , P2_R1233_U235 , P2_R1233_U232 );
and AND2_20166 ( P2_R1233_U17 , P2_R1233_U227 , P2_R1233_U224 );
and AND2_20167 ( P2_R1233_U18 , P2_R1233_U213 , P2_R1233_U210 );
not NOT1_20168 ( P2_R1233_U19 , P2_U3447 );
not NOT1_20169 ( P2_R1233_U20 , P2_U3073 );
not NOT1_20170 ( P2_R1233_U21 , P2_U3072 );
nand NAND2_20171 ( P2_R1233_U22 , P2_U3073 , P2_U3447 );
not NOT1_20172 ( P2_R1233_U23 , P2_U3450 );
not NOT1_20173 ( P2_R1233_U24 , P2_U3441 );
not NOT1_20174 ( P2_R1233_U25 , P2_U3062 );
not NOT1_20175 ( P2_R1233_U26 , P2_U3069 );
not NOT1_20176 ( P2_R1233_U27 , P2_U3435 );
not NOT1_20177 ( P2_R1233_U28 , P2_U3070 );
not NOT1_20178 ( P2_R1233_U29 , P2_U3427 );
not NOT1_20179 ( P2_R1233_U30 , P2_U3079 );
nand NAND2_20180 ( P2_R1233_U31 , P2_U3079 , P2_U3427 );
not NOT1_20181 ( P2_R1233_U32 , P2_U3438 );
not NOT1_20182 ( P2_R1233_U33 , P2_U3066 );
nand NAND2_20183 ( P2_R1233_U34 , P2_U3062 , P2_U3441 );
not NOT1_20184 ( P2_R1233_U35 , P2_U3444 );
not NOT1_20185 ( P2_R1233_U36 , P2_U3453 );
not NOT1_20186 ( P2_R1233_U37 , P2_U3086 );
not NOT1_20187 ( P2_R1233_U38 , P2_U3085 );
not NOT1_20188 ( P2_R1233_U39 , P2_U3456 );
nand NAND2_20189 ( P2_R1233_U40 , P2_R1233_U61 , P2_R1233_U205 );
nand NAND2_20190 ( P2_R1233_U41 , P2_R1233_U117 , P2_R1233_U193 );
nand NAND2_20191 ( P2_R1233_U42 , P2_R1233_U182 , P2_R1233_U183 );
nand NAND2_20192 ( P2_R1233_U43 , P2_U3432 , P2_U3080 );
nand NAND2_20193 ( P2_R1233_U44 , P2_R1233_U122 , P2_R1233_U219 );
nand NAND2_20194 ( P2_R1233_U45 , P2_R1233_U216 , P2_R1233_U215 );
not NOT1_20195 ( P2_R1233_U46 , P2_U3950 );
not NOT1_20196 ( P2_R1233_U47 , P2_U3055 );
not NOT1_20197 ( P2_R1233_U48 , P2_U3059 );
not NOT1_20198 ( P2_R1233_U49 , P2_U3951 );
not NOT1_20199 ( P2_R1233_U50 , P2_U3952 );
not NOT1_20200 ( P2_R1233_U51 , P2_U3060 );
not NOT1_20201 ( P2_R1233_U52 , P2_U3953 );
not NOT1_20202 ( P2_R1233_U53 , P2_U3067 );
not NOT1_20203 ( P2_R1233_U54 , P2_U3956 );
not NOT1_20204 ( P2_R1233_U55 , P2_U3077 );
not NOT1_20205 ( P2_R1233_U56 , P2_U3477 );
not NOT1_20206 ( P2_R1233_U57 , P2_U3075 );
not NOT1_20207 ( P2_R1233_U58 , P2_U3071 );
nand NAND2_20208 ( P2_R1233_U59 , P2_U3075 , P2_U3477 );
not NOT1_20209 ( P2_R1233_U60 , P2_U3480 );
nand NAND2_20210 ( P2_R1233_U61 , P2_U3086 , P2_U3453 );
not NOT1_20211 ( P2_R1233_U62 , P2_U3459 );
not NOT1_20212 ( P2_R1233_U63 , P2_U3064 );
not NOT1_20213 ( P2_R1233_U64 , P2_U3465 );
not NOT1_20214 ( P2_R1233_U65 , P2_U3074 );
not NOT1_20215 ( P2_R1233_U66 , P2_U3462 );
not NOT1_20216 ( P2_R1233_U67 , P2_U3065 );
nand NAND2_20217 ( P2_R1233_U68 , P2_U3065 , P2_U3462 );
not NOT1_20218 ( P2_R1233_U69 , P2_U3468 );
not NOT1_20219 ( P2_R1233_U70 , P2_U3082 );
not NOT1_20220 ( P2_R1233_U71 , P2_U3471 );
not NOT1_20221 ( P2_R1233_U72 , P2_U3081 );
not NOT1_20222 ( P2_R1233_U73 , P2_U3474 );
not NOT1_20223 ( P2_R1233_U74 , P2_U3076 );
not NOT1_20224 ( P2_R1233_U75 , P2_U3483 );
not NOT1_20225 ( P2_R1233_U76 , P2_U3084 );
nand NAND2_20226 ( P2_R1233_U77 , P2_U3084 , P2_U3483 );
not NOT1_20227 ( P2_R1233_U78 , P2_U3485 );
not NOT1_20228 ( P2_R1233_U79 , P2_U3083 );
nand NAND2_20229 ( P2_R1233_U80 , P2_U3083 , P2_U3485 );
not NOT1_20230 ( P2_R1233_U81 , P2_U3957 );
not NOT1_20231 ( P2_R1233_U82 , P2_U3955 );
not NOT1_20232 ( P2_R1233_U83 , P2_U3063 );
not NOT1_20233 ( P2_R1233_U84 , P2_U3954 );
not NOT1_20234 ( P2_R1233_U85 , P2_U3068 );
nand NAND2_20235 ( P2_R1233_U86 , P2_U3951 , P2_U3059 );
not NOT1_20236 ( P2_R1233_U87 , P2_U3056 );
not NOT1_20237 ( P2_R1233_U88 , P2_U3949 );
nand NAND2_20238 ( P2_R1233_U89 , P2_R1233_U306 , P2_R1233_U176 );
not NOT1_20239 ( P2_R1233_U90 , P2_U3078 );
nand NAND2_20240 ( P2_R1233_U91 , P2_R1233_U77 , P2_R1233_U315 );
nand NAND2_20241 ( P2_R1233_U92 , P2_R1233_U261 , P2_R1233_U260 );
nand NAND2_20242 ( P2_R1233_U93 , P2_R1233_U68 , P2_R1233_U337 );
nand NAND2_20243 ( P2_R1233_U94 , P2_R1233_U457 , P2_R1233_U456 );
nand NAND2_20244 ( P2_R1233_U95 , P2_R1233_U504 , P2_R1233_U503 );
nand NAND2_20245 ( P2_R1233_U96 , P2_R1233_U375 , P2_R1233_U374 );
nand NAND2_20246 ( P2_R1233_U97 , P2_R1233_U380 , P2_R1233_U379 );
nand NAND2_20247 ( P2_R1233_U98 , P2_R1233_U387 , P2_R1233_U386 );
nand NAND2_20248 ( P2_R1233_U99 , P2_R1233_U394 , P2_R1233_U393 );
nand NAND2_20249 ( P2_R1233_U100 , P2_R1233_U399 , P2_R1233_U398 );
nand NAND2_20250 ( P2_R1233_U101 , P2_R1233_U408 , P2_R1233_U407 );
nand NAND2_20251 ( P2_R1233_U102 , P2_R1233_U415 , P2_R1233_U414 );
nand NAND2_20252 ( P2_R1233_U103 , P2_R1233_U422 , P2_R1233_U421 );
nand NAND2_20253 ( P2_R1233_U104 , P2_R1233_U429 , P2_R1233_U428 );
nand NAND2_20254 ( P2_R1233_U105 , P2_R1233_U434 , P2_R1233_U433 );
nand NAND2_20255 ( P2_R1233_U106 , P2_R1233_U441 , P2_R1233_U440 );
nand NAND2_20256 ( P2_R1233_U107 , P2_R1233_U448 , P2_R1233_U447 );
nand NAND2_20257 ( P2_R1233_U108 , P2_R1233_U462 , P2_R1233_U461 );
nand NAND2_20258 ( P2_R1233_U109 , P2_R1233_U467 , P2_R1233_U466 );
nand NAND2_20259 ( P2_R1233_U110 , P2_R1233_U474 , P2_R1233_U473 );
nand NAND2_20260 ( P2_R1233_U111 , P2_R1233_U481 , P2_R1233_U480 );
nand NAND2_20261 ( P2_R1233_U112 , P2_R1233_U488 , P2_R1233_U487 );
nand NAND2_20262 ( P2_R1233_U113 , P2_R1233_U495 , P2_R1233_U494 );
nand NAND2_20263 ( P2_R1233_U114 , P2_R1233_U500 , P2_R1233_U499 );
and AND2_20264 ( P2_R1233_U115 , P2_R1233_U189 , P2_R1233_U187 );
and AND2_20265 ( P2_R1233_U116 , P2_R1233_U4 , P2_R1233_U180 );
and AND2_20266 ( P2_R1233_U117 , P2_R1233_U194 , P2_R1233_U192 );
and AND2_20267 ( P2_R1233_U118 , P2_R1233_U201 , P2_R1233_U200 );
and AND3_20268 ( P2_R1233_U119 , P2_R1233_U382 , P2_R1233_U381 , P2_R1233_U22 );
and AND2_20269 ( P2_R1233_U120 , P2_R1233_U212 , P2_R1233_U5 );
and AND2_20270 ( P2_R1233_U121 , P2_R1233_U181 , P2_R1233_U180 );
and AND2_20271 ( P2_R1233_U122 , P2_R1233_U220 , P2_R1233_U218 );
and AND3_20272 ( P2_R1233_U123 , P2_R1233_U389 , P2_R1233_U388 , P2_R1233_U34 );
and AND2_20273 ( P2_R1233_U124 , P2_R1233_U226 , P2_R1233_U4 );
and AND2_20274 ( P2_R1233_U125 , P2_R1233_U234 , P2_R1233_U181 );
and AND2_20275 ( P2_R1233_U126 , P2_R1233_U204 , P2_R1233_U6 );
and AND2_20276 ( P2_R1233_U127 , P2_R1233_U239 , P2_R1233_U171 );
and AND2_20277 ( P2_R1233_U128 , P2_R1233_U250 , P2_R1233_U7 );
and AND2_20278 ( P2_R1233_U129 , P2_R1233_U248 , P2_R1233_U172 );
and AND2_20279 ( P2_R1233_U130 , P2_R1233_U268 , P2_R1233_U267 );
and AND2_20280 ( P2_R1233_U131 , P2_R1233_U9 , P2_R1233_U282 );
and AND2_20281 ( P2_R1233_U132 , P2_R1233_U285 , P2_R1233_U280 );
and AND2_20282 ( P2_R1233_U133 , P2_R1233_U301 , P2_R1233_U298 );
and AND2_20283 ( P2_R1233_U134 , P2_R1233_U368 , P2_R1233_U302 );
and AND2_20284 ( P2_R1233_U135 , P2_R1233_U160 , P2_R1233_U278 );
and AND3_20285 ( P2_R1233_U136 , P2_R1233_U455 , P2_R1233_U454 , P2_R1233_U80 );
and AND2_20286 ( P2_R1233_U137 , P2_R1233_U325 , P2_R1233_U9 );
and AND3_20287 ( P2_R1233_U138 , P2_R1233_U469 , P2_R1233_U468 , P2_R1233_U59 );
and AND2_20288 ( P2_R1233_U139 , P2_R1233_U334 , P2_R1233_U8 );
and AND3_20289 ( P2_R1233_U140 , P2_R1233_U490 , P2_R1233_U489 , P2_R1233_U172 );
and AND2_20290 ( P2_R1233_U141 , P2_R1233_U343 , P2_R1233_U7 );
and AND3_20291 ( P2_R1233_U142 , P2_R1233_U502 , P2_R1233_U501 , P2_R1233_U171 );
and AND2_20292 ( P2_R1233_U143 , P2_R1233_U350 , P2_R1233_U6 );
nand NAND2_20293 ( P2_R1233_U144 , P2_R1233_U118 , P2_R1233_U202 );
nand NAND2_20294 ( P2_R1233_U145 , P2_R1233_U217 , P2_R1233_U229 );
not NOT1_20295 ( P2_R1233_U146 , P2_U3057 );
not NOT1_20296 ( P2_R1233_U147 , P2_U3960 );
and AND2_20297 ( P2_R1233_U148 , P2_R1233_U403 , P2_R1233_U402 );
nand NAND3_20298 ( P2_R1233_U149 , P2_R1233_U304 , P2_R1233_U169 , P2_R1233_U364 );
and AND2_20299 ( P2_R1233_U150 , P2_R1233_U410 , P2_R1233_U409 );
nand NAND3_20300 ( P2_R1233_U151 , P2_R1233_U370 , P2_R1233_U369 , P2_R1233_U134 );
and AND2_20301 ( P2_R1233_U152 , P2_R1233_U417 , P2_R1233_U416 );
nand NAND3_20302 ( P2_R1233_U153 , P2_R1233_U365 , P2_R1233_U299 , P2_R1233_U86 );
and AND2_20303 ( P2_R1233_U154 , P2_R1233_U424 , P2_R1233_U423 );
nand NAND2_20304 ( P2_R1233_U155 , P2_R1233_U293 , P2_R1233_U292 );
and AND2_20305 ( P2_R1233_U156 , P2_R1233_U436 , P2_R1233_U435 );
nand NAND2_20306 ( P2_R1233_U157 , P2_R1233_U289 , P2_R1233_U288 );
and AND2_20307 ( P2_R1233_U158 , P2_R1233_U443 , P2_R1233_U442 );
nand NAND2_20308 ( P2_R1233_U159 , P2_R1233_U132 , P2_R1233_U284 );
and AND2_20309 ( P2_R1233_U160 , P2_R1233_U450 , P2_R1233_U449 );
nand NAND2_20310 ( P2_R1233_U161 , P2_R1233_U43 , P2_R1233_U327 );
nand NAND2_20311 ( P2_R1233_U162 , P2_R1233_U130 , P2_R1233_U269 );
and AND2_20312 ( P2_R1233_U163 , P2_R1233_U476 , P2_R1233_U475 );
nand NAND2_20313 ( P2_R1233_U164 , P2_R1233_U257 , P2_R1233_U256 );
and AND2_20314 ( P2_R1233_U165 , P2_R1233_U483 , P2_R1233_U482 );
nand NAND2_20315 ( P2_R1233_U166 , P2_R1233_U253 , P2_R1233_U252 );
nand NAND2_20316 ( P2_R1233_U167 , P2_R1233_U243 , P2_R1233_U242 );
nand NAND2_20317 ( P2_R1233_U168 , P2_R1233_U367 , P2_R1233_U366 );
nand NAND2_20318 ( P2_R1233_U169 , P2_U3056 , P2_R1233_U151 );
not NOT1_20319 ( P2_R1233_U170 , P2_R1233_U34 );
nand NAND2_20320 ( P2_R1233_U171 , P2_U3456 , P2_U3085 );
nand NAND2_20321 ( P2_R1233_U172 , P2_U3074 , P2_U3465 );
nand NAND2_20322 ( P2_R1233_U173 , P2_U3060 , P2_U3952 );
not NOT1_20323 ( P2_R1233_U174 , P2_R1233_U68 );
not NOT1_20324 ( P2_R1233_U175 , P2_R1233_U77 );
nand NAND2_20325 ( P2_R1233_U176 , P2_U3067 , P2_U3953 );
not NOT1_20326 ( P2_R1233_U177 , P2_R1233_U61 );
or OR2_20327 ( P2_R1233_U178 , P2_U3069 , P2_U3444 );
or OR2_20328 ( P2_R1233_U179 , P2_U3062 , P2_U3441 );
or OR2_20329 ( P2_R1233_U180 , P2_U3438 , P2_U3066 );
or OR2_20330 ( P2_R1233_U181 , P2_U3435 , P2_U3070 );
not NOT1_20331 ( P2_R1233_U182 , P2_R1233_U31 );
or OR2_20332 ( P2_R1233_U183 , P2_U3432 , P2_U3080 );
not NOT1_20333 ( P2_R1233_U184 , P2_R1233_U42 );
not NOT1_20334 ( P2_R1233_U185 , P2_R1233_U43 );
nand NAND2_20335 ( P2_R1233_U186 , P2_R1233_U42 , P2_R1233_U43 );
nand NAND2_20336 ( P2_R1233_U187 , P2_U3070 , P2_U3435 );
nand NAND2_20337 ( P2_R1233_U188 , P2_R1233_U186 , P2_R1233_U181 );
nand NAND2_20338 ( P2_R1233_U189 , P2_U3066 , P2_U3438 );
nand NAND2_20339 ( P2_R1233_U190 , P2_R1233_U115 , P2_R1233_U188 );
nand NAND2_20340 ( P2_R1233_U191 , P2_R1233_U35 , P2_R1233_U34 );
nand NAND2_20341 ( P2_R1233_U192 , P2_U3069 , P2_R1233_U191 );
nand NAND2_20342 ( P2_R1233_U193 , P2_R1233_U116 , P2_R1233_U190 );
nand NAND2_20343 ( P2_R1233_U194 , P2_U3444 , P2_R1233_U170 );
not NOT1_20344 ( P2_R1233_U195 , P2_R1233_U41 );
or OR2_20345 ( P2_R1233_U196 , P2_U3072 , P2_U3450 );
or OR2_20346 ( P2_R1233_U197 , P2_U3073 , P2_U3447 );
not NOT1_20347 ( P2_R1233_U198 , P2_R1233_U22 );
nand NAND2_20348 ( P2_R1233_U199 , P2_R1233_U23 , P2_R1233_U22 );
nand NAND2_20349 ( P2_R1233_U200 , P2_U3072 , P2_R1233_U199 );
nand NAND2_20350 ( P2_R1233_U201 , P2_U3450 , P2_R1233_U198 );
nand NAND2_20351 ( P2_R1233_U202 , P2_R1233_U5 , P2_R1233_U41 );
not NOT1_20352 ( P2_R1233_U203 , P2_R1233_U144 );
or OR2_20353 ( P2_R1233_U204 , P2_U3453 , P2_U3086 );
nand NAND2_20354 ( P2_R1233_U205 , P2_R1233_U204 , P2_R1233_U144 );
not NOT1_20355 ( P2_R1233_U206 , P2_R1233_U40 );
or OR2_20356 ( P2_R1233_U207 , P2_U3085 , P2_U3456 );
or OR2_20357 ( P2_R1233_U208 , P2_U3447 , P2_U3073 );
nand NAND2_20358 ( P2_R1233_U209 , P2_R1233_U208 , P2_R1233_U41 );
nand NAND2_20359 ( P2_R1233_U210 , P2_R1233_U119 , P2_R1233_U209 );
nand NAND2_20360 ( P2_R1233_U211 , P2_R1233_U195 , P2_R1233_U22 );
nand NAND2_20361 ( P2_R1233_U212 , P2_U3450 , P2_U3072 );
nand NAND2_20362 ( P2_R1233_U213 , P2_R1233_U120 , P2_R1233_U211 );
or OR2_20363 ( P2_R1233_U214 , P2_U3073 , P2_U3447 );
nand NAND2_20364 ( P2_R1233_U215 , P2_R1233_U185 , P2_R1233_U181 );
nand NAND2_20365 ( P2_R1233_U216 , P2_U3070 , P2_U3435 );
not NOT1_20366 ( P2_R1233_U217 , P2_R1233_U45 );
nand NAND2_20367 ( P2_R1233_U218 , P2_R1233_U121 , P2_R1233_U184 );
nand NAND2_20368 ( P2_R1233_U219 , P2_R1233_U45 , P2_R1233_U180 );
nand NAND2_20369 ( P2_R1233_U220 , P2_U3066 , P2_U3438 );
not NOT1_20370 ( P2_R1233_U221 , P2_R1233_U44 );
or OR2_20371 ( P2_R1233_U222 , P2_U3441 , P2_U3062 );
nand NAND2_20372 ( P2_R1233_U223 , P2_R1233_U222 , P2_R1233_U44 );
nand NAND2_20373 ( P2_R1233_U224 , P2_R1233_U123 , P2_R1233_U223 );
nand NAND2_20374 ( P2_R1233_U225 , P2_R1233_U221 , P2_R1233_U34 );
nand NAND2_20375 ( P2_R1233_U226 , P2_U3444 , P2_U3069 );
nand NAND2_20376 ( P2_R1233_U227 , P2_R1233_U124 , P2_R1233_U225 );
or OR2_20377 ( P2_R1233_U228 , P2_U3062 , P2_U3441 );
nand NAND2_20378 ( P2_R1233_U229 , P2_R1233_U184 , P2_R1233_U181 );
not NOT1_20379 ( P2_R1233_U230 , P2_R1233_U145 );
nand NAND2_20380 ( P2_R1233_U231 , P2_U3066 , P2_U3438 );
nand NAND4_20381 ( P2_R1233_U232 , P2_R1233_U401 , P2_R1233_U400 , P2_R1233_U43 , P2_R1233_U42 );
nand NAND2_20382 ( P2_R1233_U233 , P2_R1233_U43 , P2_R1233_U42 );
nand NAND2_20383 ( P2_R1233_U234 , P2_U3070 , P2_U3435 );
nand NAND2_20384 ( P2_R1233_U235 , P2_R1233_U125 , P2_R1233_U233 );
or OR2_20385 ( P2_R1233_U236 , P2_U3085 , P2_U3456 );
or OR2_20386 ( P2_R1233_U237 , P2_U3064 , P2_U3459 );
nand NAND2_20387 ( P2_R1233_U238 , P2_R1233_U177 , P2_R1233_U6 );
nand NAND2_20388 ( P2_R1233_U239 , P2_U3064 , P2_U3459 );
nand NAND2_20389 ( P2_R1233_U240 , P2_R1233_U127 , P2_R1233_U238 );
or OR2_20390 ( P2_R1233_U241 , P2_U3459 , P2_U3064 );
nand NAND2_20391 ( P2_R1233_U242 , P2_R1233_U126 , P2_R1233_U144 );
nand NAND2_20392 ( P2_R1233_U243 , P2_R1233_U241 , P2_R1233_U240 );
not NOT1_20393 ( P2_R1233_U244 , P2_R1233_U167 );
or OR2_20394 ( P2_R1233_U245 , P2_U3082 , P2_U3468 );
or OR2_20395 ( P2_R1233_U246 , P2_U3074 , P2_U3465 );
nand NAND2_20396 ( P2_R1233_U247 , P2_R1233_U174 , P2_R1233_U7 );
nand NAND2_20397 ( P2_R1233_U248 , P2_U3082 , P2_U3468 );
nand NAND2_20398 ( P2_R1233_U249 , P2_R1233_U129 , P2_R1233_U247 );
or OR2_20399 ( P2_R1233_U250 , P2_U3462 , P2_U3065 );
or OR2_20400 ( P2_R1233_U251 , P2_U3468 , P2_U3082 );
nand NAND2_20401 ( P2_R1233_U252 , P2_R1233_U128 , P2_R1233_U167 );
nand NAND2_20402 ( P2_R1233_U253 , P2_R1233_U251 , P2_R1233_U249 );
not NOT1_20403 ( P2_R1233_U254 , P2_R1233_U166 );
or OR2_20404 ( P2_R1233_U255 , P2_U3471 , P2_U3081 );
nand NAND2_20405 ( P2_R1233_U256 , P2_R1233_U255 , P2_R1233_U166 );
nand NAND2_20406 ( P2_R1233_U257 , P2_U3081 , P2_U3471 );
not NOT1_20407 ( P2_R1233_U258 , P2_R1233_U164 );
or OR2_20408 ( P2_R1233_U259 , P2_U3474 , P2_U3076 );
nand NAND2_20409 ( P2_R1233_U260 , P2_R1233_U259 , P2_R1233_U164 );
nand NAND2_20410 ( P2_R1233_U261 , P2_U3076 , P2_U3474 );
not NOT1_20411 ( P2_R1233_U262 , P2_R1233_U92 );
or OR2_20412 ( P2_R1233_U263 , P2_U3071 , P2_U3480 );
or OR2_20413 ( P2_R1233_U264 , P2_U3075 , P2_U3477 );
not NOT1_20414 ( P2_R1233_U265 , P2_R1233_U59 );
nand NAND2_20415 ( P2_R1233_U266 , P2_R1233_U60 , P2_R1233_U59 );
nand NAND2_20416 ( P2_R1233_U267 , P2_U3071 , P2_R1233_U266 );
nand NAND2_20417 ( P2_R1233_U268 , P2_U3480 , P2_R1233_U265 );
nand NAND2_20418 ( P2_R1233_U269 , P2_R1233_U8 , P2_R1233_U92 );
not NOT1_20419 ( P2_R1233_U270 , P2_R1233_U162 );
or OR2_20420 ( P2_R1233_U271 , P2_U3078 , P2_U3957 );
or OR2_20421 ( P2_R1233_U272 , P2_U3083 , P2_U3485 );
or OR2_20422 ( P2_R1233_U273 , P2_U3077 , P2_U3956 );
not NOT1_20423 ( P2_R1233_U274 , P2_R1233_U80 );
nand NAND2_20424 ( P2_R1233_U275 , P2_U3957 , P2_R1233_U274 );
nand NAND2_20425 ( P2_R1233_U276 , P2_R1233_U275 , P2_R1233_U90 );
nand NAND2_20426 ( P2_R1233_U277 , P2_R1233_U80 , P2_R1233_U81 );
nand NAND2_20427 ( P2_R1233_U278 , P2_R1233_U277 , P2_R1233_U276 );
nand NAND2_20428 ( P2_R1233_U279 , P2_R1233_U175 , P2_R1233_U9 );
nand NAND2_20429 ( P2_R1233_U280 , P2_U3077 , P2_U3956 );
nand NAND2_20430 ( P2_R1233_U281 , P2_R1233_U278 , P2_R1233_U279 );
or OR2_20431 ( P2_R1233_U282 , P2_U3483 , P2_U3084 );
or OR2_20432 ( P2_R1233_U283 , P2_U3956 , P2_U3077 );
nand NAND3_20433 ( P2_R1233_U284 , P2_R1233_U273 , P2_R1233_U162 , P2_R1233_U131 );
nand NAND2_20434 ( P2_R1233_U285 , P2_R1233_U283 , P2_R1233_U281 );
not NOT1_20435 ( P2_R1233_U286 , P2_R1233_U159 );
or OR2_20436 ( P2_R1233_U287 , P2_U3955 , P2_U3063 );
nand NAND2_20437 ( P2_R1233_U288 , P2_R1233_U287 , P2_R1233_U159 );
nand NAND2_20438 ( P2_R1233_U289 , P2_U3063 , P2_U3955 );
not NOT1_20439 ( P2_R1233_U290 , P2_R1233_U157 );
or OR2_20440 ( P2_R1233_U291 , P2_U3954 , P2_U3068 );
nand NAND2_20441 ( P2_R1233_U292 , P2_R1233_U291 , P2_R1233_U157 );
nand NAND2_20442 ( P2_R1233_U293 , P2_U3068 , P2_U3954 );
not NOT1_20443 ( P2_R1233_U294 , P2_R1233_U155 );
or OR2_20444 ( P2_R1233_U295 , P2_U3060 , P2_U3952 );
nand NAND2_20445 ( P2_R1233_U296 , P2_R1233_U176 , P2_R1233_U173 );
not NOT1_20446 ( P2_R1233_U297 , P2_R1233_U86 );
or OR2_20447 ( P2_R1233_U298 , P2_U3953 , P2_U3067 );
nand NAND3_20448 ( P2_R1233_U299 , P2_R1233_U155 , P2_R1233_U298 , P2_R1233_U168 );
not NOT1_20449 ( P2_R1233_U300 , P2_R1233_U153 );
or OR2_20450 ( P2_R1233_U301 , P2_U3950 , P2_U3055 );
nand NAND2_20451 ( P2_R1233_U302 , P2_U3055 , P2_U3950 );
not NOT1_20452 ( P2_R1233_U303 , P2_R1233_U151 );
nand NAND2_20453 ( P2_R1233_U304 , P2_U3949 , P2_R1233_U151 );
not NOT1_20454 ( P2_R1233_U305 , P2_R1233_U149 );
nand NAND2_20455 ( P2_R1233_U306 , P2_R1233_U298 , P2_R1233_U155 );
not NOT1_20456 ( P2_R1233_U307 , P2_R1233_U89 );
or OR2_20457 ( P2_R1233_U308 , P2_U3952 , P2_U3060 );
nand NAND2_20458 ( P2_R1233_U309 , P2_R1233_U308 , P2_R1233_U89 );
nand NAND3_20459 ( P2_R1233_U310 , P2_R1233_U309 , P2_R1233_U173 , P2_R1233_U154 );
nand NAND2_20460 ( P2_R1233_U311 , P2_R1233_U307 , P2_R1233_U173 );
nand NAND2_20461 ( P2_R1233_U312 , P2_U3951 , P2_U3059 );
nand NAND3_20462 ( P2_R1233_U313 , P2_R1233_U311 , P2_R1233_U312 , P2_R1233_U168 );
or OR2_20463 ( P2_R1233_U314 , P2_U3060 , P2_U3952 );
nand NAND2_20464 ( P2_R1233_U315 , P2_R1233_U282 , P2_R1233_U162 );
not NOT1_20465 ( P2_R1233_U316 , P2_R1233_U91 );
nand NAND2_20466 ( P2_R1233_U317 , P2_R1233_U9 , P2_R1233_U91 );
nand NAND2_20467 ( P2_R1233_U318 , P2_R1233_U135 , P2_R1233_U317 );
nand NAND2_20468 ( P2_R1233_U319 , P2_R1233_U317 , P2_R1233_U278 );
nand NAND2_20469 ( P2_R1233_U320 , P2_R1233_U453 , P2_R1233_U319 );
or OR2_20470 ( P2_R1233_U321 , P2_U3485 , P2_U3083 );
nand NAND2_20471 ( P2_R1233_U322 , P2_R1233_U321 , P2_R1233_U91 );
nand NAND2_20472 ( P2_R1233_U323 , P2_R1233_U136 , P2_R1233_U322 );
nand NAND2_20473 ( P2_R1233_U324 , P2_R1233_U316 , P2_R1233_U80 );
nand NAND2_20474 ( P2_R1233_U325 , P2_U3078 , P2_U3957 );
nand NAND2_20475 ( P2_R1233_U326 , P2_R1233_U137 , P2_R1233_U324 );
or OR2_20476 ( P2_R1233_U327 , P2_U3432 , P2_U3080 );
not NOT1_20477 ( P2_R1233_U328 , P2_R1233_U161 );
or OR2_20478 ( P2_R1233_U329 , P2_U3083 , P2_U3485 );
or OR2_20479 ( P2_R1233_U330 , P2_U3477 , P2_U3075 );
nand NAND2_20480 ( P2_R1233_U331 , P2_R1233_U330 , P2_R1233_U92 );
nand NAND2_20481 ( P2_R1233_U332 , P2_R1233_U138 , P2_R1233_U331 );
nand NAND2_20482 ( P2_R1233_U333 , P2_R1233_U262 , P2_R1233_U59 );
nand NAND2_20483 ( P2_R1233_U334 , P2_U3480 , P2_U3071 );
nand NAND2_20484 ( P2_R1233_U335 , P2_R1233_U139 , P2_R1233_U333 );
or OR2_20485 ( P2_R1233_U336 , P2_U3075 , P2_U3477 );
nand NAND2_20486 ( P2_R1233_U337 , P2_R1233_U250 , P2_R1233_U167 );
not NOT1_20487 ( P2_R1233_U338 , P2_R1233_U93 );
or OR2_20488 ( P2_R1233_U339 , P2_U3465 , P2_U3074 );
nand NAND2_20489 ( P2_R1233_U340 , P2_R1233_U339 , P2_R1233_U93 );
nand NAND2_20490 ( P2_R1233_U341 , P2_R1233_U140 , P2_R1233_U340 );
nand NAND2_20491 ( P2_R1233_U342 , P2_R1233_U338 , P2_R1233_U172 );
nand NAND2_20492 ( P2_R1233_U343 , P2_U3082 , P2_U3468 );
nand NAND2_20493 ( P2_R1233_U344 , P2_R1233_U141 , P2_R1233_U342 );
or OR2_20494 ( P2_R1233_U345 , P2_U3074 , P2_U3465 );
or OR2_20495 ( P2_R1233_U346 , P2_U3456 , P2_U3085 );
nand NAND2_20496 ( P2_R1233_U347 , P2_R1233_U346 , P2_R1233_U40 );
nand NAND2_20497 ( P2_R1233_U348 , P2_R1233_U142 , P2_R1233_U347 );
nand NAND2_20498 ( P2_R1233_U349 , P2_R1233_U206 , P2_R1233_U171 );
nand NAND2_20499 ( P2_R1233_U350 , P2_U3064 , P2_U3459 );
nand NAND2_20500 ( P2_R1233_U351 , P2_R1233_U143 , P2_R1233_U349 );
nand NAND2_20501 ( P2_R1233_U352 , P2_R1233_U207 , P2_R1233_U171 );
nand NAND2_20502 ( P2_R1233_U353 , P2_R1233_U204 , P2_R1233_U61 );
nand NAND2_20503 ( P2_R1233_U354 , P2_R1233_U214 , P2_R1233_U22 );
nand NAND2_20504 ( P2_R1233_U355 , P2_R1233_U228 , P2_R1233_U34 );
nand NAND2_20505 ( P2_R1233_U356 , P2_R1233_U231 , P2_R1233_U180 );
nand NAND2_20506 ( P2_R1233_U357 , P2_R1233_U314 , P2_R1233_U173 );
nand NAND2_20507 ( P2_R1233_U358 , P2_R1233_U298 , P2_R1233_U176 );
nand NAND2_20508 ( P2_R1233_U359 , P2_R1233_U329 , P2_R1233_U80 );
nand NAND2_20509 ( P2_R1233_U360 , P2_R1233_U282 , P2_R1233_U77 );
nand NAND2_20510 ( P2_R1233_U361 , P2_R1233_U336 , P2_R1233_U59 );
nand NAND2_20511 ( P2_R1233_U362 , P2_R1233_U345 , P2_R1233_U172 );
nand NAND2_20512 ( P2_R1233_U363 , P2_R1233_U250 , P2_R1233_U68 );
nand NAND2_20513 ( P2_R1233_U364 , P2_U3949 , P2_U3056 );
nand NAND2_20514 ( P2_R1233_U365 , P2_R1233_U296 , P2_R1233_U168 );
nand NAND2_20515 ( P2_R1233_U366 , P2_U3059 , P2_R1233_U295 );
nand NAND2_20516 ( P2_R1233_U367 , P2_U3951 , P2_R1233_U295 );
nand NAND3_20517 ( P2_R1233_U368 , P2_R1233_U296 , P2_R1233_U168 , P2_R1233_U301 );
nand NAND3_20518 ( P2_R1233_U369 , P2_R1233_U155 , P2_R1233_U168 , P2_R1233_U133 );
nand NAND2_20519 ( P2_R1233_U370 , P2_R1233_U297 , P2_R1233_U301 );
nand NAND2_20520 ( P2_R1233_U371 , P2_U3085 , P2_R1233_U39 );
nand NAND2_20521 ( P2_R1233_U372 , P2_U3456 , P2_R1233_U38 );
nand NAND2_20522 ( P2_R1233_U373 , P2_R1233_U372 , P2_R1233_U371 );
nand NAND2_20523 ( P2_R1233_U374 , P2_R1233_U352 , P2_R1233_U40 );
nand NAND2_20524 ( P2_R1233_U375 , P2_R1233_U373 , P2_R1233_U206 );
nand NAND2_20525 ( P2_R1233_U376 , P2_U3086 , P2_R1233_U36 );
nand NAND2_20526 ( P2_R1233_U377 , P2_U3453 , P2_R1233_U37 );
nand NAND2_20527 ( P2_R1233_U378 , P2_R1233_U377 , P2_R1233_U376 );
nand NAND2_20528 ( P2_R1233_U379 , P2_R1233_U353 , P2_R1233_U144 );
nand NAND2_20529 ( P2_R1233_U380 , P2_R1233_U203 , P2_R1233_U378 );
nand NAND2_20530 ( P2_R1233_U381 , P2_U3072 , P2_R1233_U23 );
nand NAND2_20531 ( P2_R1233_U382 , P2_U3450 , P2_R1233_U21 );
nand NAND2_20532 ( P2_R1233_U383 , P2_U3073 , P2_R1233_U19 );
nand NAND2_20533 ( P2_R1233_U384 , P2_U3447 , P2_R1233_U20 );
nand NAND2_20534 ( P2_R1233_U385 , P2_R1233_U384 , P2_R1233_U383 );
nand NAND2_20535 ( P2_R1233_U386 , P2_R1233_U354 , P2_R1233_U41 );
nand NAND2_20536 ( P2_R1233_U387 , P2_R1233_U385 , P2_R1233_U195 );
nand NAND2_20537 ( P2_R1233_U388 , P2_U3069 , P2_R1233_U35 );
nand NAND2_20538 ( P2_R1233_U389 , P2_U3444 , P2_R1233_U26 );
nand NAND2_20539 ( P2_R1233_U390 , P2_U3062 , P2_R1233_U24 );
nand NAND2_20540 ( P2_R1233_U391 , P2_U3441 , P2_R1233_U25 );
nand NAND2_20541 ( P2_R1233_U392 , P2_R1233_U391 , P2_R1233_U390 );
nand NAND2_20542 ( P2_R1233_U393 , P2_R1233_U355 , P2_R1233_U44 );
nand NAND2_20543 ( P2_R1233_U394 , P2_R1233_U392 , P2_R1233_U221 );
nand NAND2_20544 ( P2_R1233_U395 , P2_U3066 , P2_R1233_U32 );
nand NAND2_20545 ( P2_R1233_U396 , P2_U3438 , P2_R1233_U33 );
nand NAND2_20546 ( P2_R1233_U397 , P2_R1233_U396 , P2_R1233_U395 );
nand NAND2_20547 ( P2_R1233_U398 , P2_R1233_U356 , P2_R1233_U145 );
nand NAND2_20548 ( P2_R1233_U399 , P2_R1233_U230 , P2_R1233_U397 );
nand NAND2_20549 ( P2_R1233_U400 , P2_U3070 , P2_R1233_U27 );
nand NAND2_20550 ( P2_R1233_U401 , P2_U3435 , P2_R1233_U28 );
nand NAND2_20551 ( P2_R1233_U402 , P2_U3057 , P2_R1233_U147 );
nand NAND2_20552 ( P2_R1233_U403 , P2_U3960 , P2_R1233_U146 );
nand NAND2_20553 ( P2_R1233_U404 , P2_U3057 , P2_R1233_U147 );
nand NAND2_20554 ( P2_R1233_U405 , P2_U3960 , P2_R1233_U146 );
nand NAND2_20555 ( P2_R1233_U406 , P2_R1233_U405 , P2_R1233_U404 );
nand NAND2_20556 ( P2_R1233_U407 , P2_R1233_U148 , P2_R1233_U149 );
nand NAND2_20557 ( P2_R1233_U408 , P2_R1233_U305 , P2_R1233_U406 );
nand NAND2_20558 ( P2_R1233_U409 , P2_U3056 , P2_R1233_U88 );
nand NAND2_20559 ( P2_R1233_U410 , P2_U3949 , P2_R1233_U87 );
nand NAND2_20560 ( P2_R1233_U411 , P2_U3056 , P2_R1233_U88 );
nand NAND2_20561 ( P2_R1233_U412 , P2_U3949 , P2_R1233_U87 );
nand NAND2_20562 ( P2_R1233_U413 , P2_R1233_U412 , P2_R1233_U411 );
nand NAND2_20563 ( P2_R1233_U414 , P2_R1233_U150 , P2_R1233_U151 );
nand NAND2_20564 ( P2_R1233_U415 , P2_R1233_U303 , P2_R1233_U413 );
nand NAND2_20565 ( P2_R1233_U416 , P2_U3055 , P2_R1233_U46 );
nand NAND2_20566 ( P2_R1233_U417 , P2_U3950 , P2_R1233_U47 );
nand NAND2_20567 ( P2_R1233_U418 , P2_U3055 , P2_R1233_U46 );
nand NAND2_20568 ( P2_R1233_U419 , P2_U3950 , P2_R1233_U47 );
nand NAND2_20569 ( P2_R1233_U420 , P2_R1233_U419 , P2_R1233_U418 );
nand NAND2_20570 ( P2_R1233_U421 , P2_R1233_U152 , P2_R1233_U153 );
nand NAND2_20571 ( P2_R1233_U422 , P2_R1233_U300 , P2_R1233_U420 );
nand NAND2_20572 ( P2_R1233_U423 , P2_U3059 , P2_R1233_U49 );
nand NAND2_20573 ( P2_R1233_U424 , P2_U3951 , P2_R1233_U48 );
nand NAND2_20574 ( P2_R1233_U425 , P2_U3060 , P2_R1233_U50 );
nand NAND2_20575 ( P2_R1233_U426 , P2_U3952 , P2_R1233_U51 );
nand NAND2_20576 ( P2_R1233_U427 , P2_R1233_U426 , P2_R1233_U425 );
nand NAND2_20577 ( P2_R1233_U428 , P2_R1233_U357 , P2_R1233_U89 );
nand NAND2_20578 ( P2_R1233_U429 , P2_R1233_U427 , P2_R1233_U307 );
nand NAND2_20579 ( P2_R1233_U430 , P2_U3067 , P2_R1233_U52 );
nand NAND2_20580 ( P2_R1233_U431 , P2_U3953 , P2_R1233_U53 );
nand NAND2_20581 ( P2_R1233_U432 , P2_R1233_U431 , P2_R1233_U430 );
nand NAND2_20582 ( P2_R1233_U433 , P2_R1233_U358 , P2_R1233_U155 );
nand NAND2_20583 ( P2_R1233_U434 , P2_R1233_U294 , P2_R1233_U432 );
nand NAND2_20584 ( P2_R1233_U435 , P2_U3068 , P2_R1233_U84 );
nand NAND2_20585 ( P2_R1233_U436 , P2_U3954 , P2_R1233_U85 );
nand NAND2_20586 ( P2_R1233_U437 , P2_U3068 , P2_R1233_U84 );
nand NAND2_20587 ( P2_R1233_U438 , P2_U3954 , P2_R1233_U85 );
nand NAND2_20588 ( P2_R1233_U439 , P2_R1233_U438 , P2_R1233_U437 );
nand NAND2_20589 ( P2_R1233_U440 , P2_R1233_U156 , P2_R1233_U157 );
nand NAND2_20590 ( P2_R1233_U441 , P2_R1233_U290 , P2_R1233_U439 );
nand NAND2_20591 ( P2_R1233_U442 , P2_U3063 , P2_R1233_U82 );
nand NAND2_20592 ( P2_R1233_U443 , P2_U3955 , P2_R1233_U83 );
nand NAND2_20593 ( P2_R1233_U444 , P2_U3063 , P2_R1233_U82 );
nand NAND2_20594 ( P2_R1233_U445 , P2_U3955 , P2_R1233_U83 );
nand NAND2_20595 ( P2_R1233_U446 , P2_R1233_U445 , P2_R1233_U444 );
nand NAND2_20596 ( P2_R1233_U447 , P2_R1233_U158 , P2_R1233_U159 );
nand NAND2_20597 ( P2_R1233_U448 , P2_R1233_U286 , P2_R1233_U446 );
nand NAND2_20598 ( P2_R1233_U449 , P2_U3077 , P2_R1233_U54 );
nand NAND2_20599 ( P2_R1233_U450 , P2_U3956 , P2_R1233_U55 );
nand NAND2_20600 ( P2_R1233_U451 , P2_U3077 , P2_R1233_U54 );
nand NAND2_20601 ( P2_R1233_U452 , P2_U3956 , P2_R1233_U55 );
nand NAND2_20602 ( P2_R1233_U453 , P2_R1233_U452 , P2_R1233_U451 );
nand NAND2_20603 ( P2_R1233_U454 , P2_U3078 , P2_R1233_U81 );
nand NAND2_20604 ( P2_R1233_U455 , P2_U3957 , P2_R1233_U90 );
nand NAND2_20605 ( P2_R1233_U456 , P2_R1233_U182 , P2_R1233_U161 );
nand NAND2_20606 ( P2_R1233_U457 , P2_R1233_U328 , P2_R1233_U31 );
nand NAND2_20607 ( P2_R1233_U458 , P2_U3083 , P2_R1233_U78 );
nand NAND2_20608 ( P2_R1233_U459 , P2_U3485 , P2_R1233_U79 );
nand NAND2_20609 ( P2_R1233_U460 , P2_R1233_U459 , P2_R1233_U458 );
nand NAND2_20610 ( P2_R1233_U461 , P2_R1233_U359 , P2_R1233_U91 );
nand NAND2_20611 ( P2_R1233_U462 , P2_R1233_U460 , P2_R1233_U316 );
nand NAND2_20612 ( P2_R1233_U463 , P2_U3084 , P2_R1233_U75 );
nand NAND2_20613 ( P2_R1233_U464 , P2_U3483 , P2_R1233_U76 );
nand NAND2_20614 ( P2_R1233_U465 , P2_R1233_U464 , P2_R1233_U463 );
nand NAND2_20615 ( P2_R1233_U466 , P2_R1233_U360 , P2_R1233_U162 );
nand NAND2_20616 ( P2_R1233_U467 , P2_R1233_U270 , P2_R1233_U465 );
nand NAND2_20617 ( P2_R1233_U468 , P2_U3071 , P2_R1233_U60 );
nand NAND2_20618 ( P2_R1233_U469 , P2_U3480 , P2_R1233_U58 );
nand NAND2_20619 ( P2_R1233_U470 , P2_U3075 , P2_R1233_U56 );
nand NAND2_20620 ( P2_R1233_U471 , P2_U3477 , P2_R1233_U57 );
nand NAND2_20621 ( P2_R1233_U472 , P2_R1233_U471 , P2_R1233_U470 );
nand NAND2_20622 ( P2_R1233_U473 , P2_R1233_U361 , P2_R1233_U92 );
nand NAND2_20623 ( P2_R1233_U474 , P2_R1233_U472 , P2_R1233_U262 );
nand NAND2_20624 ( P2_R1233_U475 , P2_U3076 , P2_R1233_U73 );
nand NAND2_20625 ( P2_R1233_U476 , P2_U3474 , P2_R1233_U74 );
nand NAND2_20626 ( P2_R1233_U477 , P2_U3076 , P2_R1233_U73 );
nand NAND2_20627 ( P2_R1233_U478 , P2_U3474 , P2_R1233_U74 );
nand NAND2_20628 ( P2_R1233_U479 , P2_R1233_U478 , P2_R1233_U477 );
nand NAND2_20629 ( P2_R1233_U480 , P2_R1233_U163 , P2_R1233_U164 );
nand NAND2_20630 ( P2_R1233_U481 , P2_R1233_U258 , P2_R1233_U479 );
nand NAND2_20631 ( P2_R1233_U482 , P2_U3081 , P2_R1233_U71 );
nand NAND2_20632 ( P2_R1233_U483 , P2_U3471 , P2_R1233_U72 );
nand NAND2_20633 ( P2_R1233_U484 , P2_U3081 , P2_R1233_U71 );
nand NAND2_20634 ( P2_R1233_U485 , P2_U3471 , P2_R1233_U72 );
nand NAND2_20635 ( P2_R1233_U486 , P2_R1233_U485 , P2_R1233_U484 );
nand NAND2_20636 ( P2_R1233_U487 , P2_R1233_U165 , P2_R1233_U166 );
nand NAND2_20637 ( P2_R1233_U488 , P2_R1233_U254 , P2_R1233_U486 );
nand NAND2_20638 ( P2_R1233_U489 , P2_U3082 , P2_R1233_U69 );
nand NAND2_20639 ( P2_R1233_U490 , P2_U3468 , P2_R1233_U70 );
nand NAND2_20640 ( P2_R1233_U491 , P2_U3074 , P2_R1233_U64 );
nand NAND2_20641 ( P2_R1233_U492 , P2_U3465 , P2_R1233_U65 );
nand NAND2_20642 ( P2_R1233_U493 , P2_R1233_U492 , P2_R1233_U491 );
nand NAND2_20643 ( P2_R1233_U494 , P2_R1233_U362 , P2_R1233_U93 );
nand NAND2_20644 ( P2_R1233_U495 , P2_R1233_U493 , P2_R1233_U338 );
nand NAND2_20645 ( P2_R1233_U496 , P2_U3065 , P2_R1233_U66 );
nand NAND2_20646 ( P2_R1233_U497 , P2_U3462 , P2_R1233_U67 );
nand NAND2_20647 ( P2_R1233_U498 , P2_R1233_U497 , P2_R1233_U496 );
nand NAND2_20648 ( P2_R1233_U499 , P2_R1233_U363 , P2_R1233_U167 );
nand NAND2_20649 ( P2_R1233_U500 , P2_R1233_U244 , P2_R1233_U498 );
nand NAND2_20650 ( P2_R1233_U501 , P2_U3064 , P2_R1233_U62 );
nand NAND2_20651 ( P2_R1233_U502 , P2_U3459 , P2_R1233_U63 );
nand NAND2_20652 ( P2_R1233_U503 , P2_U3079 , P2_R1233_U29 );
nand NAND2_20653 ( P2_R1233_U504 , P2_U3427 , P2_R1233_U30 );
and AND2_20654 ( P2_R1176_U4 , P2_R1176_U221 , P2_R1176_U220 );
and AND2_20655 ( P2_R1176_U5 , P2_R1176_U234 , P2_R1176_U233 );
and AND2_20656 ( P2_R1176_U6 , P2_R1176_U264 , P2_R1176_U263 );
and AND2_20657 ( P2_R1176_U7 , P2_R1176_U280 , P2_R1176_U279 );
and AND2_20658 ( P2_R1176_U8 , P2_R1176_U292 , P2_R1176_U291 );
and AND2_20659 ( P2_R1176_U9 , P2_R1176_U6 , P2_R1176_U268 );
and AND2_20660 ( P2_R1176_U10 , P2_R1176_U5 , P2_R1176_U229 );
and AND2_20661 ( P2_R1176_U11 , P2_R1176_U9 , P2_R1176_U259 );
and AND2_20662 ( P2_R1176_U12 , P2_R1176_U528 , P2_R1176_U527 );
and AND2_20663 ( P2_R1176_U13 , P2_R1176_U351 , P2_R1176_U348 );
and AND2_20664 ( P2_R1176_U14 , P2_R1176_U342 , P2_R1176_U339 );
and AND2_20665 ( P2_R1176_U15 , P2_R1176_U335 , P2_R1176_U332 );
and AND3_20666 ( P2_R1176_U16 , P2_R1176_U326 , P2_R1176_U323 , P2_R1176_U385 );
and AND2_20667 ( P2_R1176_U17 , P2_R1176_U255 , P2_R1176_U252 );
and AND2_20668 ( P2_R1176_U18 , P2_R1176_U248 , P2_R1176_U245 );
not NOT1_20669 ( P2_R1176_U19 , P2_U3184 );
not NOT1_20670 ( P2_R1176_U20 , P2_U3175 );
not NOT1_20671 ( P2_R1176_U21 , P2_U3181 );
nand NAND2_20672 ( P2_R1176_U22 , P2_U3181 , P2_R1176_U66 );
not NOT1_20673 ( P2_R1176_U23 , P2_U3180 );
not NOT1_20674 ( P2_R1176_U24 , P2_U3182 );
not NOT1_20675 ( P2_R1176_U25 , P2_U3183 );
nand NAND2_20676 ( P2_R1176_U26 , P2_U3184 , P2_R1176_U69 );
not NOT1_20677 ( P2_R1176_U27 , P2_U3179 );
not NOT1_20678 ( P2_R1176_U28 , P2_U3177 );
nand NAND2_20679 ( P2_R1176_U29 , P2_U3177 , P2_R1176_U73 );
not NOT1_20680 ( P2_R1176_U30 , P2_U3176 );
not NOT1_20681 ( P2_R1176_U31 , P2_U3178 );
nand NAND2_20682 ( P2_R1176_U32 , P2_U3178 , P2_R1176_U71 );
not NOT1_20683 ( P2_R1176_U33 , P2_U3174 );
nand NAND3_20684 ( P2_R1176_U34 , P2_R1176_U238 , P2_R1176_U237 , P2_R1176_U369 );
nand NAND2_20685 ( P2_R1176_U35 , P2_R1176_U32 , P2_R1176_U230 );
nand NAND3_20686 ( P2_R1176_U36 , P2_R1176_U366 , P2_R1176_U218 , P2_R1176_U365 );
not NOT1_20687 ( P2_R1176_U37 , P2_U3156 );
not NOT1_20688 ( P2_R1176_U38 , P2_U3158 );
not NOT1_20689 ( P2_R1176_U39 , P2_U3159 );
not NOT1_20690 ( P2_R1176_U40 , P2_U3157 );
not NOT1_20691 ( P2_R1176_U41 , P2_U3167 );
nand NAND2_20692 ( P2_R1176_U42 , P2_U3167 , P2_R1176_U78 );
not NOT1_20693 ( P2_R1176_U43 , P2_U3166 );
not NOT1_20694 ( P2_R1176_U44 , P2_U3169 );
not NOT1_20695 ( P2_R1176_U45 , P2_U3171 );
not NOT1_20696 ( P2_R1176_U46 , P2_U3172 );
nand NAND2_20697 ( P2_R1176_U47 , P2_U3172 , P2_R1176_U82 );
not NOT1_20698 ( P2_R1176_U48 , P2_U3170 );
not NOT1_20699 ( P2_R1176_U49 , P2_U3173 );
nand NAND2_20700 ( P2_R1176_U50 , P2_U3173 , P2_R1176_U81 );
not NOT1_20701 ( P2_R1176_U51 , P2_U3168 );
not NOT1_20702 ( P2_R1176_U52 , P2_U3165 );
not NOT1_20703 ( P2_R1176_U53 , P2_U3163 );
not NOT1_20704 ( P2_R1176_U54 , P2_U3164 );
nand NAND2_20705 ( P2_R1176_U55 , P2_U3164 , P2_R1176_U87 );
not NOT1_20706 ( P2_R1176_U56 , P2_U3162 );
not NOT1_20707 ( P2_R1176_U57 , P2_U3161 );
not NOT1_20708 ( P2_R1176_U58 , P2_U3160 );
nand NAND2_20709 ( P2_R1176_U59 , P2_R1176_U212 , P2_R1176_U321 );
nand NAND2_20710 ( P2_R1176_U60 , P2_R1176_U55 , P2_R1176_U328 );
nand NAND2_20711 ( P2_R1176_U61 , P2_R1176_U277 , P2_R1176_U276 );
nand NAND2_20712 ( P2_R1176_U62 , P2_R1176_U374 , P2_R1176_U270 );
nand NAND2_20713 ( P2_R1176_U63 , P2_R1176_U47 , P2_R1176_U344 );
nand NAND2_20714 ( P2_R1176_U64 , P2_R1176_U387 , P2_R1176_U386 );
nand NAND2_20715 ( P2_R1176_U65 , P2_R1176_U419 , P2_R1176_U418 );
nand NAND2_20716 ( P2_R1176_U66 , P2_R1176_U407 , P2_R1176_U406 );
nand NAND2_20717 ( P2_R1176_U67 , P2_R1176_U404 , P2_R1176_U403 );
nand NAND2_20718 ( P2_R1176_U68 , P2_R1176_U398 , P2_R1176_U397 );
nand NAND2_20719 ( P2_R1176_U69 , P2_R1176_U401 , P2_R1176_U400 );
nand NAND2_20720 ( P2_R1176_U70 , P2_R1176_U395 , P2_R1176_U394 );
nand NAND2_20721 ( P2_R1176_U71 , P2_R1176_U410 , P2_R1176_U409 );
nand NAND2_20722 ( P2_R1176_U72 , P2_R1176_U413 , P2_R1176_U412 );
nand NAND2_20723 ( P2_R1176_U73 , P2_R1176_U416 , P2_R1176_U415 );
nand NAND2_20724 ( P2_R1176_U74 , P2_R1176_U459 , P2_R1176_U458 );
nand NAND2_20725 ( P2_R1176_U75 , P2_R1176_U507 , P2_R1176_U506 );
nand NAND2_20726 ( P2_R1176_U76 , P2_R1176_U510 , P2_R1176_U509 );
nand NAND2_20727 ( P2_R1176_U77 , P2_R1176_U462 , P2_R1176_U461 );
nand NAND2_20728 ( P2_R1176_U78 , P2_R1176_U486 , P2_R1176_U485 );
nand NAND2_20729 ( P2_R1176_U79 , P2_R1176_U483 , P2_R1176_U482 );
nand NAND2_20730 ( P2_R1176_U80 , P2_R1176_U477 , P2_R1176_U476 );
nand NAND2_20731 ( P2_R1176_U81 , P2_R1176_U465 , P2_R1176_U464 );
nand NAND2_20732 ( P2_R1176_U82 , P2_R1176_U468 , P2_R1176_U467 );
nand NAND2_20733 ( P2_R1176_U83 , P2_R1176_U471 , P2_R1176_U470 );
nand NAND2_20734 ( P2_R1176_U84 , P2_R1176_U474 , P2_R1176_U473 );
nand NAND2_20735 ( P2_R1176_U85 , P2_R1176_U480 , P2_R1176_U479 );
nand NAND2_20736 ( P2_R1176_U86 , P2_R1176_U489 , P2_R1176_U488 );
nand NAND2_20737 ( P2_R1176_U87 , P2_R1176_U498 , P2_R1176_U497 );
nand NAND2_20738 ( P2_R1176_U88 , P2_R1176_U492 , P2_R1176_U491 );
nand NAND2_20739 ( P2_R1176_U89 , P2_R1176_U495 , P2_R1176_U494 );
nand NAND2_20740 ( P2_R1176_U90 , P2_R1176_U501 , P2_R1176_U500 );
nand NAND2_20741 ( P2_R1176_U91 , P2_R1176_U504 , P2_R1176_U503 );
nand NAND2_20742 ( P2_R1176_U92 , P2_R1176_U516 , P2_R1176_U515 );
nand NAND2_20743 ( P2_R1176_U93 , P2_R1176_U623 , P2_R1176_U622 );
nand NAND2_20744 ( P2_R1176_U94 , P2_R1176_U422 , P2_R1176_U421 );
nand NAND2_20745 ( P2_R1176_U95 , P2_R1176_U429 , P2_R1176_U428 );
nand NAND2_20746 ( P2_R1176_U96 , P2_R1176_U436 , P2_R1176_U435 );
nand NAND2_20747 ( P2_R1176_U97 , P2_R1176_U443 , P2_R1176_U442 );
nand NAND2_20748 ( P2_R1176_U98 , P2_R1176_U450 , P2_R1176_U449 );
nand NAND2_20749 ( P2_R1176_U99 , P2_R1176_U457 , P2_R1176_U456 );
nand NAND2_20750 ( P2_R1176_U100 , P2_R1176_U519 , P2_R1176_U518 );
nand NAND2_20751 ( P2_R1176_U101 , P2_R1176_U526 , P2_R1176_U525 );
nand NAND2_20752 ( P2_R1176_U102 , P2_R1176_U533 , P2_R1176_U532 );
nand NAND2_20753 ( P2_R1176_U103 , P2_R1176_U538 , P2_R1176_U537 );
nand NAND2_20754 ( P2_R1176_U104 , P2_R1176_U545 , P2_R1176_U544 );
nand NAND2_20755 ( P2_R1176_U105 , P2_R1176_U552 , P2_R1176_U551 );
nand NAND2_20756 ( P2_R1176_U106 , P2_R1176_U559 , P2_R1176_U558 );
nand NAND2_20757 ( P2_R1176_U107 , P2_R1176_U566 , P2_R1176_U565 );
nand NAND2_20758 ( P2_R1176_U108 , P2_R1176_U571 , P2_R1176_U570 );
nand NAND2_20759 ( P2_R1176_U109 , P2_R1176_U578 , P2_R1176_U577 );
nand NAND2_20760 ( P2_R1176_U110 , P2_R1176_U585 , P2_R1176_U584 );
nand NAND2_20761 ( P2_R1176_U111 , P2_R1176_U592 , P2_R1176_U591 );
nand NAND2_20762 ( P2_R1176_U112 , P2_R1176_U599 , P2_R1176_U598 );
nand NAND2_20763 ( P2_R1176_U113 , P2_R1176_U606 , P2_R1176_U605 );
nand NAND2_20764 ( P2_R1176_U114 , P2_R1176_U611 , P2_R1176_U610 );
nand NAND2_20765 ( P2_R1176_U115 , P2_R1176_U618 , P2_R1176_U617 );
and AND2_20766 ( P2_R1176_U116 , P2_R1176_U224 , P2_R1176_U223 );
and AND2_20767 ( P2_R1176_U117 , P2_R1176_U240 , P2_R1176_U10 );
and AND2_20768 ( P2_R1176_U118 , P2_R1176_U372 , P2_R1176_U241 );
and AND3_20769 ( P2_R1176_U119 , P2_R1176_U431 , P2_R1176_U430 , P2_R1176_U29 );
and AND2_20770 ( P2_R1176_U120 , P2_R1176_U247 , P2_R1176_U5 );
and AND3_20771 ( P2_R1176_U121 , P2_R1176_U452 , P2_R1176_U451 , P2_R1176_U22 );
and AND2_20772 ( P2_R1176_U122 , P2_R1176_U254 , P2_R1176_U4 );
and AND2_20773 ( P2_R1176_U123 , P2_R1176_U272 , P2_R1176_U11 );
and AND2_20774 ( P2_R1176_U124 , P2_R1176_U266 , P2_R1176_U207 );
and AND2_20775 ( P2_R1176_U125 , P2_R1176_U380 , P2_R1176_U273 );
and AND2_20776 ( P2_R1176_U126 , P2_R1176_U284 , P2_R1176_U283 );
and AND2_20777 ( P2_R1176_U127 , P2_R1176_U296 , P2_R1176_U8 );
and AND2_20778 ( P2_R1176_U128 , P2_R1176_U294 , P2_R1176_U208 );
and AND2_20779 ( P2_R1176_U129 , P2_R1176_U312 , P2_R1176_U203 );
and AND2_20780 ( P2_R1176_U130 , P2_R1176_U383 , P2_R1176_U318 );
and AND2_20781 ( P2_R1176_U131 , P2_R1176_U320 , P2_R1176_U310 );
and AND2_20782 ( P2_R1176_U132 , P2_R1176_U320 , P2_R1176_U312 );
and AND2_20783 ( P2_R1176_U133 , P2_R1176_U381 , P2_R1176_U319 );
nand NAND2_20784 ( P2_R1176_U134 , P2_R1176_U513 , P2_R1176_U512 );
and AND2_20785 ( P2_R1176_U135 , P2_R1176_U508 , P2_R1176_U38 );
and AND2_20786 ( P2_R1176_U136 , P2_R1176_U212 , P2_R1176_U209 );
and AND2_20787 ( P2_R1176_U137 , P2_R1176_U325 , P2_R1176_U203 );
and AND2_20788 ( P2_R1176_U138 , P2_R1176_U12 , P2_R1176_U209 );
and AND3_20789 ( P2_R1176_U139 , P2_R1176_U554 , P2_R1176_U553 , P2_R1176_U208 );
and AND2_20790 ( P2_R1176_U140 , P2_R1176_U334 , P2_R1176_U8 );
and AND3_20791 ( P2_R1176_U141 , P2_R1176_U580 , P2_R1176_U579 , P2_R1176_U42 );
and AND2_20792 ( P2_R1176_U142 , P2_R1176_U341 , P2_R1176_U7 );
and AND3_20793 ( P2_R1176_U143 , P2_R1176_U601 , P2_R1176_U600 , P2_R1176_U207 );
and AND2_20794 ( P2_R1176_U144 , P2_R1176_U350 , P2_R1176_U6 );
nand NAND2_20795 ( P2_R1176_U145 , P2_R1176_U620 , P2_R1176_U619 );
not NOT1_20796 ( P2_R1176_U146 , P2_U3456 );
and AND2_20797 ( P2_R1176_U147 , P2_R1176_U390 , P2_R1176_U389 );
not NOT1_20798 ( P2_R1176_U148 , P2_U3441 );
not NOT1_20799 ( P2_R1176_U149 , P2_U3432 );
not NOT1_20800 ( P2_R1176_U150 , P2_U3427 );
not NOT1_20801 ( P2_R1176_U151 , P2_U3438 );
not NOT1_20802 ( P2_R1176_U152 , P2_U3435 );
not NOT1_20803 ( P2_R1176_U153 , P2_U3444 );
not NOT1_20804 ( P2_R1176_U154 , P2_U3450 );
not NOT1_20805 ( P2_R1176_U155 , P2_U3447 );
not NOT1_20806 ( P2_R1176_U156 , P2_U3453 );
nand NAND2_20807 ( P2_R1176_U157 , P2_R1176_U118 , P2_R1176_U371 );
and AND2_20808 ( P2_R1176_U158 , P2_R1176_U424 , P2_R1176_U423 );
nand NAND2_20809 ( P2_R1176_U159 , P2_R1176_U370 , P2_R1176_U368 );
and AND2_20810 ( P2_R1176_U160 , P2_R1176_U438 , P2_R1176_U437 );
nand NAND3_20811 ( P2_R1176_U161 , P2_R1176_U227 , P2_R1176_U205 , P2_R1176_U362 );
and AND2_20812 ( P2_R1176_U162 , P2_R1176_U445 , P2_R1176_U444 );
nand NAND2_20813 ( P2_R1176_U163 , P2_R1176_U116 , P2_R1176_U225 );
not NOT1_20814 ( P2_R1176_U164 , P2_U3950 );
not NOT1_20815 ( P2_R1176_U165 , P2_U3951 );
not NOT1_20816 ( P2_R1176_U166 , P2_U3459 );
not NOT1_20817 ( P2_R1176_U167 , P2_U3462 );
not NOT1_20818 ( P2_R1176_U168 , P2_U3468 );
not NOT1_20819 ( P2_R1176_U169 , P2_U3465 );
not NOT1_20820 ( P2_R1176_U170 , P2_U3471 );
not NOT1_20821 ( P2_R1176_U171 , P2_U3474 );
not NOT1_20822 ( P2_R1176_U172 , P2_U3480 );
not NOT1_20823 ( P2_R1176_U173 , P2_U3477 );
not NOT1_20824 ( P2_R1176_U174 , P2_U3483 );
not NOT1_20825 ( P2_R1176_U175 , P2_U3956 );
not NOT1_20826 ( P2_R1176_U176 , P2_U3957 );
not NOT1_20827 ( P2_R1176_U177 , P2_U3485 );
not NOT1_20828 ( P2_R1176_U178 , P2_U3955 );
not NOT1_20829 ( P2_R1176_U179 , P2_U3954 );
not NOT1_20830 ( P2_R1176_U180 , P2_U3952 );
not NOT1_20831 ( P2_R1176_U181 , P2_U3953 );
not NOT1_20832 ( P2_R1176_U182 , P2_U3949 );
not NOT1_20833 ( P2_R1176_U183 , P2_U3155 );
and AND2_20834 ( P2_R1176_U184 , P2_R1176_U521 , P2_R1176_U520 );
nand NAND2_20835 ( P2_R1176_U185 , P2_R1176_U315 , P2_R1176_U314 );
nand NAND2_20836 ( P2_R1176_U186 , P2_R1176_U307 , P2_R1176_U306 );
and AND2_20837 ( P2_R1176_U187 , P2_R1176_U540 , P2_R1176_U539 );
nand NAND2_20838 ( P2_R1176_U188 , P2_R1176_U303 , P2_R1176_U302 );
and AND2_20839 ( P2_R1176_U189 , P2_R1176_U547 , P2_R1176_U546 );
nand NAND2_20840 ( P2_R1176_U190 , P2_R1176_U299 , P2_R1176_U298 );
and AND2_20841 ( P2_R1176_U191 , P2_R1176_U561 , P2_R1176_U560 );
nand NAND2_20842 ( P2_R1176_U192 , P2_R1176_U26 , P2_R1176_U214 );
nand NAND2_20843 ( P2_R1176_U193 , P2_R1176_U289 , P2_R1176_U288 );
and AND2_20844 ( P2_R1176_U194 , P2_R1176_U573 , P2_R1176_U572 );
nand NAND2_20845 ( P2_R1176_U195 , P2_R1176_U126 , P2_R1176_U285 );
and AND2_20846 ( P2_R1176_U196 , P2_R1176_U587 , P2_R1176_U586 );
nand NAND2_20847 ( P2_R1176_U197 , P2_R1176_U125 , P2_R1176_U379 );
and AND2_20848 ( P2_R1176_U198 , P2_R1176_U594 , P2_R1176_U593 );
nand NAND2_20849 ( P2_R1176_U199 , P2_R1176_U378 , P2_R1176_U373 );
nand NAND2_20850 ( P2_R1176_U200 , P2_R1176_U50 , P2_R1176_U260 );
and AND2_20851 ( P2_R1176_U201 , P2_R1176_U613 , P2_R1176_U612 );
nand NAND3_20852 ( P2_R1176_U202 , P2_R1176_U257 , P2_R1176_U204 , P2_R1176_U363 );
nand NAND2_20853 ( P2_R1176_U203 , P2_R1176_U377 , P2_R1176_U376 );
nand NAND2_20854 ( P2_R1176_U204 , P2_R1176_U64 , P2_R1176_U157 );
nand NAND2_20855 ( P2_R1176_U205 , P2_R1176_U70 , P2_R1176_U163 );
not NOT1_20856 ( P2_R1176_U206 , P2_R1176_U22 );
nand NAND2_20857 ( P2_R1176_U207 , P2_U3171 , P2_R1176_U84 );
nand NAND2_20858 ( P2_R1176_U208 , P2_U3163 , P2_R1176_U89 );
nand NAND2_20859 ( P2_R1176_U209 , P2_U3158 , P2_R1176_U75 );
not NOT1_20860 ( P2_R1176_U210 , P2_R1176_U47 );
not NOT1_20861 ( P2_R1176_U211 , P2_R1176_U55 );
nand NAND2_20862 ( P2_R1176_U212 , P2_U3159 , P2_R1176_U76 );
nand NAND2_20863 ( P2_R1176_U213 , P2_R1176_U402 , P2_R1176_U19 );
nand NAND2_20864 ( P2_R1176_U214 , P2_U3183 , P2_R1176_U213 );
not NOT1_20865 ( P2_R1176_U215 , P2_R1176_U26 );
not NOT1_20866 ( P2_R1176_U216 , P2_R1176_U192 );
nand NAND2_20867 ( P2_R1176_U217 , P2_R1176_U399 , P2_R1176_U24 );
nand NAND2_20868 ( P2_R1176_U218 , P2_U3182 , P2_R1176_U68 );
not NOT1_20869 ( P2_R1176_U219 , P2_R1176_U36 );
nand NAND2_20870 ( P2_R1176_U220 , P2_R1176_U405 , P2_R1176_U23 );
nand NAND2_20871 ( P2_R1176_U221 , P2_R1176_U408 , P2_R1176_U21 );
nand NAND2_20872 ( P2_R1176_U222 , P2_R1176_U23 , P2_R1176_U22 );
nand NAND2_20873 ( P2_R1176_U223 , P2_R1176_U67 , P2_R1176_U222 );
nand NAND2_20874 ( P2_R1176_U224 , P2_U3180 , P2_R1176_U206 );
nand NAND2_20875 ( P2_R1176_U225 , P2_R1176_U4 , P2_R1176_U36 );
not NOT1_20876 ( P2_R1176_U226 , P2_R1176_U163 );
nand NAND2_20877 ( P2_R1176_U227 , P2_U3179 , P2_R1176_U163 );
not NOT1_20878 ( P2_R1176_U228 , P2_R1176_U161 );
nand NAND2_20879 ( P2_R1176_U229 , P2_R1176_U411 , P2_R1176_U31 );
nand NAND2_20880 ( P2_R1176_U230 , P2_R1176_U229 , P2_R1176_U161 );
not NOT1_20881 ( P2_R1176_U231 , P2_R1176_U32 );
not NOT1_20882 ( P2_R1176_U232 , P2_R1176_U35 );
nand NAND2_20883 ( P2_R1176_U233 , P2_R1176_U414 , P2_R1176_U30 );
nand NAND2_20884 ( P2_R1176_U234 , P2_R1176_U417 , P2_R1176_U28 );
not NOT1_20885 ( P2_R1176_U235 , P2_R1176_U29 );
nand NAND2_20886 ( P2_R1176_U236 , P2_R1176_U30 , P2_R1176_U29 );
nand NAND2_20887 ( P2_R1176_U237 , P2_R1176_U72 , P2_R1176_U236 );
nand NAND2_20888 ( P2_R1176_U238 , P2_U3176 , P2_R1176_U235 );
not NOT1_20889 ( P2_R1176_U239 , P2_R1176_U159 );
nand NAND2_20890 ( P2_R1176_U240 , P2_R1176_U420 , P2_R1176_U20 );
nand NAND2_20891 ( P2_R1176_U241 , P2_U3175 , P2_R1176_U65 );
not NOT1_20892 ( P2_R1176_U242 , P2_R1176_U157 );
nand NAND2_20893 ( P2_R1176_U243 , P2_R1176_U417 , P2_R1176_U28 );
nand NAND2_20894 ( P2_R1176_U244 , P2_R1176_U243 , P2_R1176_U35 );
nand NAND2_20895 ( P2_R1176_U245 , P2_R1176_U119 , P2_R1176_U244 );
nand NAND2_20896 ( P2_R1176_U246 , P2_R1176_U232 , P2_R1176_U29 );
nand NAND2_20897 ( P2_R1176_U247 , P2_U3176 , P2_R1176_U72 );
nand NAND2_20898 ( P2_R1176_U248 , P2_R1176_U120 , P2_R1176_U246 );
nand NAND2_20899 ( P2_R1176_U249 , P2_R1176_U417 , P2_R1176_U28 );
nand NAND2_20900 ( P2_R1176_U250 , P2_R1176_U408 , P2_R1176_U21 );
nand NAND2_20901 ( P2_R1176_U251 , P2_R1176_U250 , P2_R1176_U36 );
nand NAND2_20902 ( P2_R1176_U252 , P2_R1176_U121 , P2_R1176_U251 );
nand NAND2_20903 ( P2_R1176_U253 , P2_R1176_U219 , P2_R1176_U22 );
nand NAND2_20904 ( P2_R1176_U254 , P2_U3180 , P2_R1176_U67 );
nand NAND2_20905 ( P2_R1176_U255 , P2_R1176_U122 , P2_R1176_U253 );
nand NAND2_20906 ( P2_R1176_U256 , P2_R1176_U408 , P2_R1176_U21 );
nand NAND2_20907 ( P2_R1176_U257 , P2_U3174 , P2_R1176_U157 );
not NOT1_20908 ( P2_R1176_U258 , P2_R1176_U202 );
nand NAND2_20909 ( P2_R1176_U259 , P2_R1176_U466 , P2_R1176_U49 );
nand NAND2_20910 ( P2_R1176_U260 , P2_R1176_U259 , P2_R1176_U202 );
not NOT1_20911 ( P2_R1176_U261 , P2_R1176_U50 );
not NOT1_20912 ( P2_R1176_U262 , P2_R1176_U200 );
nand NAND2_20913 ( P2_R1176_U263 , P2_R1176_U472 , P2_R1176_U48 );
nand NAND2_20914 ( P2_R1176_U264 , P2_R1176_U475 , P2_R1176_U45 );
nand NAND2_20915 ( P2_R1176_U265 , P2_R1176_U210 , P2_R1176_U6 );
nand NAND2_20916 ( P2_R1176_U266 , P2_U3170 , P2_R1176_U83 );
nand NAND2_20917 ( P2_R1176_U267 , P2_R1176_U124 , P2_R1176_U265 );
nand NAND2_20918 ( P2_R1176_U268 , P2_R1176_U469 , P2_R1176_U46 );
nand NAND2_20919 ( P2_R1176_U269 , P2_R1176_U472 , P2_R1176_U48 );
nand NAND2_20920 ( P2_R1176_U270 , P2_R1176_U269 , P2_R1176_U267 );
not NOT1_20921 ( P2_R1176_U271 , P2_R1176_U199 );
nand NAND2_20922 ( P2_R1176_U272 , P2_R1176_U478 , P2_R1176_U44 );
nand NAND2_20923 ( P2_R1176_U273 , P2_U3169 , P2_R1176_U80 );
not NOT1_20924 ( P2_R1176_U274 , P2_R1176_U197 );
nand NAND2_20925 ( P2_R1176_U275 , P2_R1176_U481 , P2_R1176_U51 );
nand NAND2_20926 ( P2_R1176_U276 , P2_R1176_U275 , P2_R1176_U197 );
nand NAND2_20927 ( P2_R1176_U277 , P2_U3168 , P2_R1176_U85 );
not NOT1_20928 ( P2_R1176_U278 , P2_R1176_U61 );
nand NAND2_20929 ( P2_R1176_U279 , P2_R1176_U484 , P2_R1176_U43 );
nand NAND2_20930 ( P2_R1176_U280 , P2_R1176_U487 , P2_R1176_U41 );
not NOT1_20931 ( P2_R1176_U281 , P2_R1176_U42 );
nand NAND2_20932 ( P2_R1176_U282 , P2_R1176_U43 , P2_R1176_U42 );
nand NAND2_20933 ( P2_R1176_U283 , P2_R1176_U79 , P2_R1176_U282 );
nand NAND2_20934 ( P2_R1176_U284 , P2_U3166 , P2_R1176_U281 );
nand NAND2_20935 ( P2_R1176_U285 , P2_R1176_U7 , P2_R1176_U61 );
not NOT1_20936 ( P2_R1176_U286 , P2_R1176_U195 );
nand NAND2_20937 ( P2_R1176_U287 , P2_R1176_U490 , P2_R1176_U52 );
nand NAND2_20938 ( P2_R1176_U288 , P2_R1176_U287 , P2_R1176_U195 );
nand NAND2_20939 ( P2_R1176_U289 , P2_U3165 , P2_R1176_U86 );
not NOT1_20940 ( P2_R1176_U290 , P2_R1176_U193 );
nand NAND2_20941 ( P2_R1176_U291 , P2_R1176_U493 , P2_R1176_U56 );
nand NAND2_20942 ( P2_R1176_U292 , P2_R1176_U496 , P2_R1176_U53 );
nand NAND2_20943 ( P2_R1176_U293 , P2_R1176_U211 , P2_R1176_U8 );
nand NAND2_20944 ( P2_R1176_U294 , P2_U3162 , P2_R1176_U88 );
nand NAND2_20945 ( P2_R1176_U295 , P2_R1176_U128 , P2_R1176_U293 );
nand NAND2_20946 ( P2_R1176_U296 , P2_R1176_U499 , P2_R1176_U54 );
nand NAND2_20947 ( P2_R1176_U297 , P2_R1176_U493 , P2_R1176_U56 );
nand NAND2_20948 ( P2_R1176_U298 , P2_R1176_U127 , P2_R1176_U193 );
nand NAND2_20949 ( P2_R1176_U299 , P2_R1176_U297 , P2_R1176_U295 );
not NOT1_20950 ( P2_R1176_U300 , P2_R1176_U190 );
nand NAND2_20951 ( P2_R1176_U301 , P2_R1176_U502 , P2_R1176_U57 );
nand NAND2_20952 ( P2_R1176_U302 , P2_R1176_U301 , P2_R1176_U190 );
nand NAND2_20953 ( P2_R1176_U303 , P2_U3161 , P2_R1176_U90 );
not NOT1_20954 ( P2_R1176_U304 , P2_R1176_U188 );
nand NAND2_20955 ( P2_R1176_U305 , P2_R1176_U505 , P2_R1176_U58 );
nand NAND2_20956 ( P2_R1176_U306 , P2_R1176_U305 , P2_R1176_U188 );
nand NAND2_20957 ( P2_R1176_U307 , P2_U3160 , P2_R1176_U91 );
not NOT1_20958 ( P2_R1176_U308 , P2_R1176_U186 );
nand NAND2_20959 ( P2_R1176_U309 , P2_R1176_U508 , P2_R1176_U38 );
nand NAND3_20960 ( P2_R1176_U310 , P2_R1176_U212 , P2_R1176_U209 , P2_R1176_U311 );
nand NAND2_20961 ( P2_R1176_U311 , P2_U3157 , P2_R1176_U77 );
nand NAND2_20962 ( P2_R1176_U312 , P2_R1176_U511 , P2_R1176_U39 );
nand NAND2_20963 ( P2_R1176_U313 , P2_R1176_U463 , P2_R1176_U40 );
nand NAND2_20964 ( P2_R1176_U314 , P2_R1176_U129 , P2_R1176_U186 );
nand NAND2_20965 ( P2_R1176_U315 , P2_R1176_U375 , P2_R1176_U310 );
not NOT1_20966 ( P2_R1176_U316 , P2_R1176_U185 );
nand NAND2_20967 ( P2_R1176_U317 , P2_R1176_U460 , P2_R1176_U37 );
nand NAND2_20968 ( P2_R1176_U318 , P2_U3156 , P2_R1176_U74 );
nand NAND2_20969 ( P2_R1176_U319 , P2_U3156 , P2_R1176_U74 );
nand NAND2_20970 ( P2_R1176_U320 , P2_R1176_U460 , P2_R1176_U37 );
nand NAND2_20971 ( P2_R1176_U321 , P2_R1176_U312 , P2_R1176_U186 );
not NOT1_20972 ( P2_R1176_U322 , P2_R1176_U59 );
nand NAND2_20973 ( P2_R1176_U323 , P2_R1176_U135 , P2_R1176_U12 );
nand NAND2_20974 ( P2_R1176_U324 , P2_R1176_U136 , P2_R1176_U321 );
nand NAND2_20975 ( P2_R1176_U325 , P2_U3157 , P2_R1176_U77 );
nand NAND2_20976 ( P2_R1176_U326 , P2_R1176_U137 , P2_R1176_U324 );
nand NAND2_20977 ( P2_R1176_U327 , P2_R1176_U508 , P2_R1176_U38 );
nand NAND2_20978 ( P2_R1176_U328 , P2_R1176_U296 , P2_R1176_U193 );
not NOT1_20979 ( P2_R1176_U329 , P2_R1176_U60 );
nand NAND2_20980 ( P2_R1176_U330 , P2_R1176_U496 , P2_R1176_U53 );
nand NAND2_20981 ( P2_R1176_U331 , P2_R1176_U330 , P2_R1176_U60 );
nand NAND2_20982 ( P2_R1176_U332 , P2_R1176_U139 , P2_R1176_U331 );
nand NAND2_20983 ( P2_R1176_U333 , P2_R1176_U329 , P2_R1176_U208 );
nand NAND2_20984 ( P2_R1176_U334 , P2_U3162 , P2_R1176_U88 );
nand NAND2_20985 ( P2_R1176_U335 , P2_R1176_U140 , P2_R1176_U333 );
nand NAND2_20986 ( P2_R1176_U336 , P2_R1176_U496 , P2_R1176_U53 );
nand NAND2_20987 ( P2_R1176_U337 , P2_R1176_U487 , P2_R1176_U41 );
nand NAND2_20988 ( P2_R1176_U338 , P2_R1176_U337 , P2_R1176_U61 );
nand NAND2_20989 ( P2_R1176_U339 , P2_R1176_U141 , P2_R1176_U338 );
nand NAND2_20990 ( P2_R1176_U340 , P2_R1176_U278 , P2_R1176_U42 );
nand NAND2_20991 ( P2_R1176_U341 , P2_U3166 , P2_R1176_U79 );
nand NAND2_20992 ( P2_R1176_U342 , P2_R1176_U142 , P2_R1176_U340 );
nand NAND2_20993 ( P2_R1176_U343 , P2_R1176_U487 , P2_R1176_U41 );
nand NAND2_20994 ( P2_R1176_U344 , P2_R1176_U268 , P2_R1176_U200 );
not NOT1_20995 ( P2_R1176_U345 , P2_R1176_U63 );
nand NAND2_20996 ( P2_R1176_U346 , P2_R1176_U475 , P2_R1176_U45 );
nand NAND2_20997 ( P2_R1176_U347 , P2_R1176_U346 , P2_R1176_U63 );
nand NAND2_20998 ( P2_R1176_U348 , P2_R1176_U143 , P2_R1176_U347 );
nand NAND2_20999 ( P2_R1176_U349 , P2_R1176_U345 , P2_R1176_U207 );
nand NAND2_21000 ( P2_R1176_U350 , P2_U3170 , P2_R1176_U83 );
nand NAND2_21001 ( P2_R1176_U351 , P2_R1176_U144 , P2_R1176_U349 );
nand NAND2_21002 ( P2_R1176_U352 , P2_R1176_U475 , P2_R1176_U45 );
nand NAND2_21003 ( P2_R1176_U353 , P2_R1176_U249 , P2_R1176_U29 );
nand NAND2_21004 ( P2_R1176_U354 , P2_R1176_U256 , P2_R1176_U22 );
nand NAND2_21005 ( P2_R1176_U355 , P2_R1176_U327 , P2_R1176_U209 );
nand NAND2_21006 ( P2_R1176_U356 , P2_R1176_U312 , P2_R1176_U212 );
nand NAND2_21007 ( P2_R1176_U357 , P2_R1176_U336 , P2_R1176_U208 );
nand NAND2_21008 ( P2_R1176_U358 , P2_R1176_U296 , P2_R1176_U55 );
nand NAND2_21009 ( P2_R1176_U359 , P2_R1176_U343 , P2_R1176_U42 );
nand NAND2_21010 ( P2_R1176_U360 , P2_R1176_U352 , P2_R1176_U207 );
nand NAND2_21011 ( P2_R1176_U361 , P2_R1176_U268 , P2_R1176_U47 );
nand NAND2_21012 ( P2_R1176_U362 , P2_U3179 , P2_R1176_U70 );
nand NAND2_21013 ( P2_R1176_U363 , P2_U3174 , P2_R1176_U64 );
nand NAND3_21014 ( P2_R1176_U364 , P2_R1176_U314 , P2_R1176_U311 , P2_R1176_U130 );
nand NAND3_21015 ( P2_R1176_U365 , P2_U3183 , P2_R1176_U213 , P2_R1176_U367 );
nand NAND2_21016 ( P2_R1176_U366 , P2_R1176_U215 , P2_R1176_U217 );
nand NAND2_21017 ( P2_R1176_U367 , P2_R1176_U399 , P2_R1176_U24 );
nand NAND2_21018 ( P2_R1176_U368 , P2_R1176_U10 , P2_R1176_U161 );
nand NAND2_21019 ( P2_R1176_U369 , P2_R1176_U231 , P2_R1176_U5 );
not NOT1_21020 ( P2_R1176_U370 , P2_R1176_U34 );
nand NAND2_21021 ( P2_R1176_U371 , P2_R1176_U117 , P2_R1176_U161 );
nand NAND2_21022 ( P2_R1176_U372 , P2_R1176_U34 , P2_R1176_U240 );
nand NAND2_21023 ( P2_R1176_U373 , P2_R1176_U11 , P2_R1176_U202 );
nand NAND2_21024 ( P2_R1176_U374 , P2_R1176_U261 , P2_R1176_U9 );
nand NAND3_21025 ( P2_R1176_U375 , P2_R1176_U376 , P2_R1176_U311 , P2_R1176_U377 );
nand NAND2_21026 ( P2_R1176_U376 , P2_R1176_U77 , P2_R1176_U309 );
nand NAND2_21027 ( P2_R1176_U377 , P2_U3157 , P2_R1176_U309 );
not NOT1_21028 ( P2_R1176_U378 , P2_R1176_U62 );
nand NAND2_21029 ( P2_R1176_U379 , P2_R1176_U123 , P2_R1176_U202 );
nand NAND2_21030 ( P2_R1176_U380 , P2_R1176_U62 , P2_R1176_U272 );
nand NAND2_21031 ( P2_R1176_U381 , P2_R1176_U131 , P2_R1176_U375 );
nand NAND3_21032 ( P2_R1176_U382 , P2_R1176_U186 , P2_R1176_U203 , P2_R1176_U132 );
nand NAND3_21033 ( P2_R1176_U383 , P2_R1176_U384 , P2_R1176_U309 , P2_R1176_U313 );
nand NAND2_21034 ( P2_R1176_U384 , P2_R1176_U212 , P2_R1176_U209 );
nand NAND2_21035 ( P2_R1176_U385 , P2_R1176_U138 , P2_R1176_U322 );
nand NAND2_21036 ( P2_R1176_U386 , P2_U3184 , P2_R1176_U146 );
nand NAND2_21037 ( P2_R1176_U387 , P2_U3456 , P2_R1176_U19 );
not NOT1_21038 ( P2_R1176_U388 , P2_R1176_U64 );
nand NAND2_21039 ( P2_R1176_U389 , P2_R1176_U388 , P2_U3174 );
nand NAND2_21040 ( P2_R1176_U390 , P2_R1176_U64 , P2_R1176_U33 );
nand NAND2_21041 ( P2_R1176_U391 , P2_R1176_U388 , P2_U3174 );
nand NAND2_21042 ( P2_R1176_U392 , P2_R1176_U64 , P2_R1176_U33 );
nand NAND2_21043 ( P2_R1176_U393 , P2_R1176_U392 , P2_R1176_U391 );
nand NAND2_21044 ( P2_R1176_U394 , P2_U3184 , P2_R1176_U148 );
nand NAND2_21045 ( P2_R1176_U395 , P2_U3441 , P2_R1176_U19 );
not NOT1_21046 ( P2_R1176_U396 , P2_R1176_U70 );
nand NAND2_21047 ( P2_R1176_U397 , P2_U3184 , P2_R1176_U149 );
nand NAND2_21048 ( P2_R1176_U398 , P2_U3432 , P2_R1176_U19 );
not NOT1_21049 ( P2_R1176_U399 , P2_R1176_U68 );
nand NAND2_21050 ( P2_R1176_U400 , P2_U3184 , P2_R1176_U150 );
nand NAND2_21051 ( P2_R1176_U401 , P2_U3427 , P2_R1176_U19 );
not NOT1_21052 ( P2_R1176_U402 , P2_R1176_U69 );
nand NAND2_21053 ( P2_R1176_U403 , P2_U3184 , P2_R1176_U151 );
nand NAND2_21054 ( P2_R1176_U404 , P2_U3438 , P2_R1176_U19 );
not NOT1_21055 ( P2_R1176_U405 , P2_R1176_U67 );
nand NAND2_21056 ( P2_R1176_U406 , P2_U3184 , P2_R1176_U152 );
nand NAND2_21057 ( P2_R1176_U407 , P2_U3435 , P2_R1176_U19 );
not NOT1_21058 ( P2_R1176_U408 , P2_R1176_U66 );
nand NAND2_21059 ( P2_R1176_U409 , P2_U3184 , P2_R1176_U153 );
nand NAND2_21060 ( P2_R1176_U410 , P2_U3444 , P2_R1176_U19 );
not NOT1_21061 ( P2_R1176_U411 , P2_R1176_U71 );
nand NAND2_21062 ( P2_R1176_U412 , P2_U3184 , P2_R1176_U154 );
nand NAND2_21063 ( P2_R1176_U413 , P2_U3450 , P2_R1176_U19 );
not NOT1_21064 ( P2_R1176_U414 , P2_R1176_U72 );
nand NAND2_21065 ( P2_R1176_U415 , P2_U3184 , P2_R1176_U155 );
nand NAND2_21066 ( P2_R1176_U416 , P2_U3447 , P2_R1176_U19 );
not NOT1_21067 ( P2_R1176_U417 , P2_R1176_U73 );
nand NAND2_21068 ( P2_R1176_U418 , P2_U3184 , P2_R1176_U156 );
nand NAND2_21069 ( P2_R1176_U419 , P2_U3453 , P2_R1176_U19 );
not NOT1_21070 ( P2_R1176_U420 , P2_R1176_U65 );
nand NAND2_21071 ( P2_R1176_U421 , P2_R1176_U147 , P2_R1176_U157 );
nand NAND2_21072 ( P2_R1176_U422 , P2_R1176_U242 , P2_R1176_U393 );
nand NAND2_21073 ( P2_R1176_U423 , P2_R1176_U420 , P2_U3175 );
nand NAND2_21074 ( P2_R1176_U424 , P2_R1176_U65 , P2_R1176_U20 );
nand NAND2_21075 ( P2_R1176_U425 , P2_R1176_U420 , P2_U3175 );
nand NAND2_21076 ( P2_R1176_U426 , P2_R1176_U65 , P2_R1176_U20 );
nand NAND2_21077 ( P2_R1176_U427 , P2_R1176_U426 , P2_R1176_U425 );
nand NAND2_21078 ( P2_R1176_U428 , P2_R1176_U158 , P2_R1176_U159 );
nand NAND2_21079 ( P2_R1176_U429 , P2_R1176_U239 , P2_R1176_U427 );
nand NAND2_21080 ( P2_R1176_U430 , P2_R1176_U414 , P2_U3176 );
nand NAND2_21081 ( P2_R1176_U431 , P2_R1176_U72 , P2_R1176_U30 );
nand NAND2_21082 ( P2_R1176_U432 , P2_R1176_U417 , P2_U3177 );
nand NAND2_21083 ( P2_R1176_U433 , P2_R1176_U73 , P2_R1176_U28 );
nand NAND2_21084 ( P2_R1176_U434 , P2_R1176_U433 , P2_R1176_U432 );
nand NAND2_21085 ( P2_R1176_U435 , P2_R1176_U353 , P2_R1176_U35 );
nand NAND2_21086 ( P2_R1176_U436 , P2_R1176_U434 , P2_R1176_U232 );
nand NAND2_21087 ( P2_R1176_U437 , P2_R1176_U411 , P2_U3178 );
nand NAND2_21088 ( P2_R1176_U438 , P2_R1176_U71 , P2_R1176_U31 );
nand NAND2_21089 ( P2_R1176_U439 , P2_R1176_U411 , P2_U3178 );
nand NAND2_21090 ( P2_R1176_U440 , P2_R1176_U71 , P2_R1176_U31 );
nand NAND2_21091 ( P2_R1176_U441 , P2_R1176_U440 , P2_R1176_U439 );
nand NAND2_21092 ( P2_R1176_U442 , P2_R1176_U160 , P2_R1176_U161 );
nand NAND2_21093 ( P2_R1176_U443 , P2_R1176_U228 , P2_R1176_U441 );
nand NAND2_21094 ( P2_R1176_U444 , P2_R1176_U396 , P2_U3179 );
nand NAND2_21095 ( P2_R1176_U445 , P2_R1176_U70 , P2_R1176_U27 );
nand NAND2_21096 ( P2_R1176_U446 , P2_R1176_U396 , P2_U3179 );
nand NAND2_21097 ( P2_R1176_U447 , P2_R1176_U70 , P2_R1176_U27 );
nand NAND2_21098 ( P2_R1176_U448 , P2_R1176_U447 , P2_R1176_U446 );
nand NAND2_21099 ( P2_R1176_U449 , P2_R1176_U162 , P2_R1176_U163 );
nand NAND2_21100 ( P2_R1176_U450 , P2_R1176_U226 , P2_R1176_U448 );
nand NAND2_21101 ( P2_R1176_U451 , P2_R1176_U405 , P2_U3180 );
nand NAND2_21102 ( P2_R1176_U452 , P2_R1176_U67 , P2_R1176_U23 );
nand NAND2_21103 ( P2_R1176_U453 , P2_R1176_U408 , P2_U3181 );
nand NAND2_21104 ( P2_R1176_U454 , P2_R1176_U66 , P2_R1176_U21 );
nand NAND2_21105 ( P2_R1176_U455 , P2_R1176_U454 , P2_R1176_U453 );
nand NAND2_21106 ( P2_R1176_U456 , P2_R1176_U354 , P2_R1176_U36 );
nand NAND2_21107 ( P2_R1176_U457 , P2_R1176_U455 , P2_R1176_U219 );
nand NAND2_21108 ( P2_R1176_U458 , P2_U3184 , P2_R1176_U164 );
nand NAND2_21109 ( P2_R1176_U459 , P2_U3950 , P2_R1176_U19 );
not NOT1_21110 ( P2_R1176_U460 , P2_R1176_U74 );
nand NAND2_21111 ( P2_R1176_U461 , P2_U3184 , P2_R1176_U165 );
nand NAND2_21112 ( P2_R1176_U462 , P2_U3951 , P2_R1176_U19 );
not NOT1_21113 ( P2_R1176_U463 , P2_R1176_U77 );
nand NAND2_21114 ( P2_R1176_U464 , P2_U3184 , P2_R1176_U166 );
nand NAND2_21115 ( P2_R1176_U465 , P2_U3459 , P2_R1176_U19 );
not NOT1_21116 ( P2_R1176_U466 , P2_R1176_U81 );
nand NAND2_21117 ( P2_R1176_U467 , P2_U3184 , P2_R1176_U167 );
nand NAND2_21118 ( P2_R1176_U468 , P2_U3462 , P2_R1176_U19 );
not NOT1_21119 ( P2_R1176_U469 , P2_R1176_U82 );
nand NAND2_21120 ( P2_R1176_U470 , P2_U3184 , P2_R1176_U168 );
nand NAND2_21121 ( P2_R1176_U471 , P2_U3468 , P2_R1176_U19 );
not NOT1_21122 ( P2_R1176_U472 , P2_R1176_U83 );
nand NAND2_21123 ( P2_R1176_U473 , P2_U3184 , P2_R1176_U169 );
nand NAND2_21124 ( P2_R1176_U474 , P2_U3465 , P2_R1176_U19 );
not NOT1_21125 ( P2_R1176_U475 , P2_R1176_U84 );
nand NAND2_21126 ( P2_R1176_U476 , P2_U3184 , P2_R1176_U170 );
nand NAND2_21127 ( P2_R1176_U477 , P2_U3471 , P2_R1176_U19 );
not NOT1_21128 ( P2_R1176_U478 , P2_R1176_U80 );
nand NAND2_21129 ( P2_R1176_U479 , P2_U3184 , P2_R1176_U171 );
nand NAND2_21130 ( P2_R1176_U480 , P2_U3474 , P2_R1176_U19 );
not NOT1_21131 ( P2_R1176_U481 , P2_R1176_U85 );
nand NAND2_21132 ( P2_R1176_U482 , P2_U3184 , P2_R1176_U172 );
nand NAND2_21133 ( P2_R1176_U483 , P2_U3480 , P2_R1176_U19 );
not NOT1_21134 ( P2_R1176_U484 , P2_R1176_U79 );
nand NAND2_21135 ( P2_R1176_U485 , P2_U3184 , P2_R1176_U173 );
nand NAND2_21136 ( P2_R1176_U486 , P2_U3477 , P2_R1176_U19 );
not NOT1_21137 ( P2_R1176_U487 , P2_R1176_U78 );
nand NAND2_21138 ( P2_R1176_U488 , P2_U3184 , P2_R1176_U174 );
nand NAND2_21139 ( P2_R1176_U489 , P2_U3483 , P2_R1176_U19 );
not NOT1_21140 ( P2_R1176_U490 , P2_R1176_U86 );
nand NAND2_21141 ( P2_R1176_U491 , P2_U3184 , P2_R1176_U175 );
nand NAND2_21142 ( P2_R1176_U492 , P2_U3956 , P2_R1176_U19 );
not NOT1_21143 ( P2_R1176_U493 , P2_R1176_U88 );
nand NAND2_21144 ( P2_R1176_U494 , P2_U3184 , P2_R1176_U176 );
nand NAND2_21145 ( P2_R1176_U495 , P2_U3957 , P2_R1176_U19 );
not NOT1_21146 ( P2_R1176_U496 , P2_R1176_U89 );
nand NAND2_21147 ( P2_R1176_U497 , P2_U3184 , P2_R1176_U177 );
nand NAND2_21148 ( P2_R1176_U498 , P2_U3485 , P2_R1176_U19 );
not NOT1_21149 ( P2_R1176_U499 , P2_R1176_U87 );
nand NAND2_21150 ( P2_R1176_U500 , P2_U3184 , P2_R1176_U178 );
nand NAND2_21151 ( P2_R1176_U501 , P2_U3955 , P2_R1176_U19 );
not NOT1_21152 ( P2_R1176_U502 , P2_R1176_U90 );
nand NAND2_21153 ( P2_R1176_U503 , P2_U3184 , P2_R1176_U179 );
nand NAND2_21154 ( P2_R1176_U504 , P2_U3954 , P2_R1176_U19 );
not NOT1_21155 ( P2_R1176_U505 , P2_R1176_U91 );
nand NAND2_21156 ( P2_R1176_U506 , P2_U3184 , P2_R1176_U180 );
nand NAND2_21157 ( P2_R1176_U507 , P2_U3952 , P2_R1176_U19 );
not NOT1_21158 ( P2_R1176_U508 , P2_R1176_U75 );
nand NAND2_21159 ( P2_R1176_U509 , P2_U3184 , P2_R1176_U181 );
nand NAND2_21160 ( P2_R1176_U510 , P2_U3953 , P2_R1176_U19 );
not NOT1_21161 ( P2_R1176_U511 , P2_R1176_U76 );
nand NAND2_21162 ( P2_R1176_U512 , P2_U3184 , P2_R1176_U182 );
nand NAND2_21163 ( P2_R1176_U513 , P2_U3949 , P2_R1176_U19 );
not NOT1_21164 ( P2_R1176_U514 , P2_R1176_U134 );
nand NAND2_21165 ( P2_R1176_U515 , P2_U3155 , P2_R1176_U514 );
nand NAND2_21166 ( P2_R1176_U516 , P2_R1176_U134 , P2_R1176_U183 );
not NOT1_21167 ( P2_R1176_U517 , P2_R1176_U92 );
nand NAND3_21168 ( P2_R1176_U518 , P2_R1176_U364 , P2_R1176_U317 , P2_R1176_U517 );
nand NAND3_21169 ( P2_R1176_U519 , P2_R1176_U133 , P2_R1176_U382 , P2_R1176_U92 );
nand NAND2_21170 ( P2_R1176_U520 , P2_R1176_U460 , P2_U3156 );
nand NAND2_21171 ( P2_R1176_U521 , P2_R1176_U74 , P2_R1176_U37 );
nand NAND2_21172 ( P2_R1176_U522 , P2_R1176_U460 , P2_U3156 );
nand NAND2_21173 ( P2_R1176_U523 , P2_R1176_U74 , P2_R1176_U37 );
nand NAND2_21174 ( P2_R1176_U524 , P2_R1176_U523 , P2_R1176_U522 );
nand NAND2_21175 ( P2_R1176_U525 , P2_R1176_U184 , P2_R1176_U185 );
nand NAND2_21176 ( P2_R1176_U526 , P2_R1176_U316 , P2_R1176_U524 );
nand NAND2_21177 ( P2_R1176_U527 , P2_R1176_U463 , P2_U3157 );
nand NAND2_21178 ( P2_R1176_U528 , P2_R1176_U77 , P2_R1176_U40 );
nand NAND2_21179 ( P2_R1176_U529 , P2_R1176_U508 , P2_U3158 );
nand NAND2_21180 ( P2_R1176_U530 , P2_R1176_U75 , P2_R1176_U38 );
nand NAND2_21181 ( P2_R1176_U531 , P2_R1176_U530 , P2_R1176_U529 );
nand NAND2_21182 ( P2_R1176_U532 , P2_R1176_U355 , P2_R1176_U59 );
nand NAND2_21183 ( P2_R1176_U533 , P2_R1176_U531 , P2_R1176_U322 );
nand NAND2_21184 ( P2_R1176_U534 , P2_R1176_U511 , P2_U3159 );
nand NAND2_21185 ( P2_R1176_U535 , P2_R1176_U76 , P2_R1176_U39 );
nand NAND2_21186 ( P2_R1176_U536 , P2_R1176_U535 , P2_R1176_U534 );
nand NAND2_21187 ( P2_R1176_U537 , P2_R1176_U356 , P2_R1176_U186 );
nand NAND2_21188 ( P2_R1176_U538 , P2_R1176_U308 , P2_R1176_U536 );
nand NAND2_21189 ( P2_R1176_U539 , P2_R1176_U505 , P2_U3160 );
nand NAND2_21190 ( P2_R1176_U540 , P2_R1176_U91 , P2_R1176_U58 );
nand NAND2_21191 ( P2_R1176_U541 , P2_R1176_U505 , P2_U3160 );
nand NAND2_21192 ( P2_R1176_U542 , P2_R1176_U91 , P2_R1176_U58 );
nand NAND2_21193 ( P2_R1176_U543 , P2_R1176_U542 , P2_R1176_U541 );
nand NAND2_21194 ( P2_R1176_U544 , P2_R1176_U187 , P2_R1176_U188 );
nand NAND2_21195 ( P2_R1176_U545 , P2_R1176_U304 , P2_R1176_U543 );
nand NAND2_21196 ( P2_R1176_U546 , P2_R1176_U502 , P2_U3161 );
nand NAND2_21197 ( P2_R1176_U547 , P2_R1176_U90 , P2_R1176_U57 );
nand NAND2_21198 ( P2_R1176_U548 , P2_R1176_U502 , P2_U3161 );
nand NAND2_21199 ( P2_R1176_U549 , P2_R1176_U90 , P2_R1176_U57 );
nand NAND2_21200 ( P2_R1176_U550 , P2_R1176_U549 , P2_R1176_U548 );
nand NAND2_21201 ( P2_R1176_U551 , P2_R1176_U189 , P2_R1176_U190 );
nand NAND2_21202 ( P2_R1176_U552 , P2_R1176_U300 , P2_R1176_U550 );
nand NAND2_21203 ( P2_R1176_U553 , P2_R1176_U493 , P2_U3162 );
nand NAND2_21204 ( P2_R1176_U554 , P2_R1176_U88 , P2_R1176_U56 );
nand NAND2_21205 ( P2_R1176_U555 , P2_R1176_U496 , P2_U3163 );
nand NAND2_21206 ( P2_R1176_U556 , P2_R1176_U89 , P2_R1176_U53 );
nand NAND2_21207 ( P2_R1176_U557 , P2_R1176_U556 , P2_R1176_U555 );
nand NAND2_21208 ( P2_R1176_U558 , P2_R1176_U357 , P2_R1176_U60 );
nand NAND2_21209 ( P2_R1176_U559 , P2_R1176_U557 , P2_R1176_U329 );
nand NAND2_21210 ( P2_R1176_U560 , P2_R1176_U399 , P2_U3182 );
nand NAND2_21211 ( P2_R1176_U561 , P2_R1176_U68 , P2_R1176_U24 );
nand NAND2_21212 ( P2_R1176_U562 , P2_R1176_U399 , P2_U3182 );
nand NAND2_21213 ( P2_R1176_U563 , P2_R1176_U68 , P2_R1176_U24 );
nand NAND2_21214 ( P2_R1176_U564 , P2_R1176_U563 , P2_R1176_U562 );
nand NAND2_21215 ( P2_R1176_U565 , P2_R1176_U191 , P2_R1176_U192 );
nand NAND2_21216 ( P2_R1176_U566 , P2_R1176_U216 , P2_R1176_U564 );
nand NAND2_21217 ( P2_R1176_U567 , P2_R1176_U499 , P2_U3164 );
nand NAND2_21218 ( P2_R1176_U568 , P2_R1176_U87 , P2_R1176_U54 );
nand NAND2_21219 ( P2_R1176_U569 , P2_R1176_U568 , P2_R1176_U567 );
nand NAND2_21220 ( P2_R1176_U570 , P2_R1176_U358 , P2_R1176_U193 );
nand NAND2_21221 ( P2_R1176_U571 , P2_R1176_U290 , P2_R1176_U569 );
nand NAND2_21222 ( P2_R1176_U572 , P2_R1176_U490 , P2_U3165 );
nand NAND2_21223 ( P2_R1176_U573 , P2_R1176_U86 , P2_R1176_U52 );
nand NAND2_21224 ( P2_R1176_U574 , P2_R1176_U490 , P2_U3165 );
nand NAND2_21225 ( P2_R1176_U575 , P2_R1176_U86 , P2_R1176_U52 );
nand NAND2_21226 ( P2_R1176_U576 , P2_R1176_U575 , P2_R1176_U574 );
nand NAND2_21227 ( P2_R1176_U577 , P2_R1176_U194 , P2_R1176_U195 );
nand NAND2_21228 ( P2_R1176_U578 , P2_R1176_U286 , P2_R1176_U576 );
nand NAND2_21229 ( P2_R1176_U579 , P2_R1176_U484 , P2_U3166 );
nand NAND2_21230 ( P2_R1176_U580 , P2_R1176_U79 , P2_R1176_U43 );
nand NAND2_21231 ( P2_R1176_U581 , P2_R1176_U487 , P2_U3167 );
nand NAND2_21232 ( P2_R1176_U582 , P2_R1176_U78 , P2_R1176_U41 );
nand NAND2_21233 ( P2_R1176_U583 , P2_R1176_U582 , P2_R1176_U581 );
nand NAND2_21234 ( P2_R1176_U584 , P2_R1176_U359 , P2_R1176_U61 );
nand NAND2_21235 ( P2_R1176_U585 , P2_R1176_U583 , P2_R1176_U278 );
nand NAND2_21236 ( P2_R1176_U586 , P2_R1176_U481 , P2_U3168 );
nand NAND2_21237 ( P2_R1176_U587 , P2_R1176_U85 , P2_R1176_U51 );
nand NAND2_21238 ( P2_R1176_U588 , P2_R1176_U481 , P2_U3168 );
nand NAND2_21239 ( P2_R1176_U589 , P2_R1176_U85 , P2_R1176_U51 );
nand NAND2_21240 ( P2_R1176_U590 , P2_R1176_U589 , P2_R1176_U588 );
nand NAND2_21241 ( P2_R1176_U591 , P2_R1176_U196 , P2_R1176_U197 );
nand NAND2_21242 ( P2_R1176_U592 , P2_R1176_U274 , P2_R1176_U590 );
nand NAND2_21243 ( P2_R1176_U593 , P2_R1176_U478 , P2_U3169 );
nand NAND2_21244 ( P2_R1176_U594 , P2_R1176_U80 , P2_R1176_U44 );
nand NAND2_21245 ( P2_R1176_U595 , P2_R1176_U478 , P2_U3169 );
nand NAND2_21246 ( P2_R1176_U596 , P2_R1176_U80 , P2_R1176_U44 );
nand NAND2_21247 ( P2_R1176_U597 , P2_R1176_U596 , P2_R1176_U595 );
nand NAND2_21248 ( P2_R1176_U598 , P2_R1176_U198 , P2_R1176_U199 );
nand NAND2_21249 ( P2_R1176_U599 , P2_R1176_U271 , P2_R1176_U597 );
nand NAND2_21250 ( P2_R1176_U600 , P2_R1176_U472 , P2_U3170 );
nand NAND2_21251 ( P2_R1176_U601 , P2_R1176_U83 , P2_R1176_U48 );
nand NAND2_21252 ( P2_R1176_U602 , P2_R1176_U475 , P2_U3171 );
nand NAND2_21253 ( P2_R1176_U603 , P2_R1176_U84 , P2_R1176_U45 );
nand NAND2_21254 ( P2_R1176_U604 , P2_R1176_U603 , P2_R1176_U602 );
nand NAND2_21255 ( P2_R1176_U605 , P2_R1176_U360 , P2_R1176_U63 );
nand NAND2_21256 ( P2_R1176_U606 , P2_R1176_U604 , P2_R1176_U345 );
nand NAND2_21257 ( P2_R1176_U607 , P2_R1176_U469 , P2_U3172 );
nand NAND2_21258 ( P2_R1176_U608 , P2_R1176_U82 , P2_R1176_U46 );
nand NAND2_21259 ( P2_R1176_U609 , P2_R1176_U608 , P2_R1176_U607 );
nand NAND2_21260 ( P2_R1176_U610 , P2_R1176_U361 , P2_R1176_U200 );
nand NAND2_21261 ( P2_R1176_U611 , P2_R1176_U262 , P2_R1176_U609 );
nand NAND2_21262 ( P2_R1176_U612 , P2_R1176_U466 , P2_U3173 );
nand NAND2_21263 ( P2_R1176_U613 , P2_R1176_U81 , P2_R1176_U49 );
nand NAND2_21264 ( P2_R1176_U614 , P2_R1176_U466 , P2_U3173 );
nand NAND2_21265 ( P2_R1176_U615 , P2_R1176_U81 , P2_R1176_U49 );
nand NAND2_21266 ( P2_R1176_U616 , P2_R1176_U615 , P2_R1176_U614 );
nand NAND2_21267 ( P2_R1176_U617 , P2_R1176_U201 , P2_R1176_U202 );
nand NAND2_21268 ( P2_R1176_U618 , P2_R1176_U258 , P2_R1176_U616 );
nand NAND2_21269 ( P2_R1176_U619 , P2_R1176_U69 , P2_R1176_U19 );
nand NAND2_21270 ( P2_R1176_U620 , P2_R1176_U402 , P2_U3184 );
not NOT1_21271 ( P2_R1176_U621 , P2_R1176_U145 );
nand NAND2_21272 ( P2_R1176_U622 , P2_R1176_U621 , P2_U3183 );
nand NAND2_21273 ( P2_R1176_U623 , P2_R1176_U145 , P2_R1176_U25 );
and AND2_21274 ( P2_R1131_U4 , P2_R1131_U179 , P2_R1131_U178 );
and AND2_21275 ( P2_R1131_U5 , P2_R1131_U197 , P2_R1131_U196 );
and AND2_21276 ( P2_R1131_U6 , P2_R1131_U237 , P2_R1131_U236 );
and AND2_21277 ( P2_R1131_U7 , P2_R1131_U246 , P2_R1131_U245 );
and AND2_21278 ( P2_R1131_U8 , P2_R1131_U264 , P2_R1131_U263 );
and AND2_21279 ( P2_R1131_U9 , P2_R1131_U272 , P2_R1131_U271 );
and AND2_21280 ( P2_R1131_U10 , P2_R1131_U351 , P2_R1131_U348 );
and AND2_21281 ( P2_R1131_U11 , P2_R1131_U344 , P2_R1131_U341 );
and AND2_21282 ( P2_R1131_U12 , P2_R1131_U335 , P2_R1131_U332 );
and AND2_21283 ( P2_R1131_U13 , P2_R1131_U326 , P2_R1131_U323 );
and AND2_21284 ( P2_R1131_U14 , P2_R1131_U320 , P2_R1131_U318 );
and AND2_21285 ( P2_R1131_U15 , P2_R1131_U313 , P2_R1131_U310 );
and AND2_21286 ( P2_R1131_U16 , P2_R1131_U235 , P2_R1131_U232 );
and AND2_21287 ( P2_R1131_U17 , P2_R1131_U227 , P2_R1131_U224 );
and AND2_21288 ( P2_R1131_U18 , P2_R1131_U213 , P2_R1131_U210 );
not NOT1_21289 ( P2_R1131_U19 , P2_U3447 );
not NOT1_21290 ( P2_R1131_U20 , P2_U3073 );
not NOT1_21291 ( P2_R1131_U21 , P2_U3072 );
nand NAND2_21292 ( P2_R1131_U22 , P2_U3073 , P2_U3447 );
not NOT1_21293 ( P2_R1131_U23 , P2_U3450 );
not NOT1_21294 ( P2_R1131_U24 , P2_U3441 );
not NOT1_21295 ( P2_R1131_U25 , P2_U3062 );
not NOT1_21296 ( P2_R1131_U26 , P2_U3069 );
not NOT1_21297 ( P2_R1131_U27 , P2_U3435 );
not NOT1_21298 ( P2_R1131_U28 , P2_U3070 );
not NOT1_21299 ( P2_R1131_U29 , P2_U3427 );
not NOT1_21300 ( P2_R1131_U30 , P2_U3079 );
nand NAND2_21301 ( P2_R1131_U31 , P2_U3079 , P2_U3427 );
not NOT1_21302 ( P2_R1131_U32 , P2_U3438 );
not NOT1_21303 ( P2_R1131_U33 , P2_U3066 );
nand NAND2_21304 ( P2_R1131_U34 , P2_U3062 , P2_U3441 );
not NOT1_21305 ( P2_R1131_U35 , P2_U3444 );
not NOT1_21306 ( P2_R1131_U36 , P2_U3453 );
not NOT1_21307 ( P2_R1131_U37 , P2_U3086 );
not NOT1_21308 ( P2_R1131_U38 , P2_U3085 );
not NOT1_21309 ( P2_R1131_U39 , P2_U3456 );
nand NAND2_21310 ( P2_R1131_U40 , P2_R1131_U61 , P2_R1131_U205 );
nand NAND2_21311 ( P2_R1131_U41 , P2_R1131_U117 , P2_R1131_U193 );
nand NAND2_21312 ( P2_R1131_U42 , P2_R1131_U182 , P2_R1131_U183 );
nand NAND2_21313 ( P2_R1131_U43 , P2_U3432 , P2_U3080 );
nand NAND2_21314 ( P2_R1131_U44 , P2_R1131_U122 , P2_R1131_U219 );
nand NAND2_21315 ( P2_R1131_U45 , P2_R1131_U216 , P2_R1131_U215 );
not NOT1_21316 ( P2_R1131_U46 , P2_U3950 );
not NOT1_21317 ( P2_R1131_U47 , P2_U3055 );
not NOT1_21318 ( P2_R1131_U48 , P2_U3059 );
not NOT1_21319 ( P2_R1131_U49 , P2_U3951 );
not NOT1_21320 ( P2_R1131_U50 , P2_U3952 );
not NOT1_21321 ( P2_R1131_U51 , P2_U3060 );
not NOT1_21322 ( P2_R1131_U52 , P2_U3953 );
not NOT1_21323 ( P2_R1131_U53 , P2_U3067 );
not NOT1_21324 ( P2_R1131_U54 , P2_U3956 );
not NOT1_21325 ( P2_R1131_U55 , P2_U3077 );
not NOT1_21326 ( P2_R1131_U56 , P2_U3477 );
not NOT1_21327 ( P2_R1131_U57 , P2_U3075 );
not NOT1_21328 ( P2_R1131_U58 , P2_U3071 );
nand NAND2_21329 ( P2_R1131_U59 , P2_U3075 , P2_U3477 );
not NOT1_21330 ( P2_R1131_U60 , P2_U3480 );
nand NAND2_21331 ( P2_R1131_U61 , P2_U3086 , P2_U3453 );
not NOT1_21332 ( P2_R1131_U62 , P2_U3459 );
not NOT1_21333 ( P2_R1131_U63 , P2_U3064 );
not NOT1_21334 ( P2_R1131_U64 , P2_U3465 );
not NOT1_21335 ( P2_R1131_U65 , P2_U3074 );
not NOT1_21336 ( P2_R1131_U66 , P2_U3462 );
not NOT1_21337 ( P2_R1131_U67 , P2_U3065 );
nand NAND2_21338 ( P2_R1131_U68 , P2_U3065 , P2_U3462 );
not NOT1_21339 ( P2_R1131_U69 , P2_U3468 );
not NOT1_21340 ( P2_R1131_U70 , P2_U3082 );
not NOT1_21341 ( P2_R1131_U71 , P2_U3471 );
not NOT1_21342 ( P2_R1131_U72 , P2_U3081 );
not NOT1_21343 ( P2_R1131_U73 , P2_U3474 );
not NOT1_21344 ( P2_R1131_U74 , P2_U3076 );
not NOT1_21345 ( P2_R1131_U75 , P2_U3483 );
not NOT1_21346 ( P2_R1131_U76 , P2_U3084 );
nand NAND2_21347 ( P2_R1131_U77 , P2_U3084 , P2_U3483 );
not NOT1_21348 ( P2_R1131_U78 , P2_U3485 );
not NOT1_21349 ( P2_R1131_U79 , P2_U3083 );
nand NAND2_21350 ( P2_R1131_U80 , P2_U3083 , P2_U3485 );
not NOT1_21351 ( P2_R1131_U81 , P2_U3957 );
not NOT1_21352 ( P2_R1131_U82 , P2_U3955 );
not NOT1_21353 ( P2_R1131_U83 , P2_U3063 );
not NOT1_21354 ( P2_R1131_U84 , P2_U3954 );
not NOT1_21355 ( P2_R1131_U85 , P2_U3068 );
nand NAND2_21356 ( P2_R1131_U86 , P2_U3951 , P2_U3059 );
not NOT1_21357 ( P2_R1131_U87 , P2_U3056 );
not NOT1_21358 ( P2_R1131_U88 , P2_U3949 );
nand NAND2_21359 ( P2_R1131_U89 , P2_R1131_U306 , P2_R1131_U176 );
not NOT1_21360 ( P2_R1131_U90 , P2_U3078 );
nand NAND2_21361 ( P2_R1131_U91 , P2_R1131_U77 , P2_R1131_U315 );
nand NAND2_21362 ( P2_R1131_U92 , P2_R1131_U261 , P2_R1131_U260 );
nand NAND2_21363 ( P2_R1131_U93 , P2_R1131_U68 , P2_R1131_U337 );
nand NAND2_21364 ( P2_R1131_U94 , P2_R1131_U457 , P2_R1131_U456 );
nand NAND2_21365 ( P2_R1131_U95 , P2_R1131_U504 , P2_R1131_U503 );
nand NAND2_21366 ( P2_R1131_U96 , P2_R1131_U375 , P2_R1131_U374 );
nand NAND2_21367 ( P2_R1131_U97 , P2_R1131_U380 , P2_R1131_U379 );
nand NAND2_21368 ( P2_R1131_U98 , P2_R1131_U387 , P2_R1131_U386 );
nand NAND2_21369 ( P2_R1131_U99 , P2_R1131_U394 , P2_R1131_U393 );
nand NAND2_21370 ( P2_R1131_U100 , P2_R1131_U399 , P2_R1131_U398 );
nand NAND2_21371 ( P2_R1131_U101 , P2_R1131_U408 , P2_R1131_U407 );
nand NAND2_21372 ( P2_R1131_U102 , P2_R1131_U415 , P2_R1131_U414 );
nand NAND2_21373 ( P2_R1131_U103 , P2_R1131_U422 , P2_R1131_U421 );
nand NAND2_21374 ( P2_R1131_U104 , P2_R1131_U429 , P2_R1131_U428 );
nand NAND2_21375 ( P2_R1131_U105 , P2_R1131_U434 , P2_R1131_U433 );
nand NAND2_21376 ( P2_R1131_U106 , P2_R1131_U441 , P2_R1131_U440 );
nand NAND2_21377 ( P2_R1131_U107 , P2_R1131_U448 , P2_R1131_U447 );
nand NAND2_21378 ( P2_R1131_U108 , P2_R1131_U462 , P2_R1131_U461 );
nand NAND2_21379 ( P2_R1131_U109 , P2_R1131_U467 , P2_R1131_U466 );
nand NAND2_21380 ( P2_R1131_U110 , P2_R1131_U474 , P2_R1131_U473 );
nand NAND2_21381 ( P2_R1131_U111 , P2_R1131_U481 , P2_R1131_U480 );
nand NAND2_21382 ( P2_R1131_U112 , P2_R1131_U488 , P2_R1131_U487 );
nand NAND2_21383 ( P2_R1131_U113 , P2_R1131_U495 , P2_R1131_U494 );
nand NAND2_21384 ( P2_R1131_U114 , P2_R1131_U500 , P2_R1131_U499 );
and AND2_21385 ( P2_R1131_U115 , P2_R1131_U189 , P2_R1131_U187 );
and AND2_21386 ( P2_R1131_U116 , P2_R1131_U4 , P2_R1131_U180 );
and AND2_21387 ( P2_R1131_U117 , P2_R1131_U194 , P2_R1131_U192 );
and AND2_21388 ( P2_R1131_U118 , P2_R1131_U201 , P2_R1131_U200 );
and AND3_21389 ( P2_R1131_U119 , P2_R1131_U382 , P2_R1131_U381 , P2_R1131_U22 );
and AND2_21390 ( P2_R1131_U120 , P2_R1131_U212 , P2_R1131_U5 );
and AND2_21391 ( P2_R1131_U121 , P2_R1131_U181 , P2_R1131_U180 );
and AND2_21392 ( P2_R1131_U122 , P2_R1131_U220 , P2_R1131_U218 );
and AND3_21393 ( P2_R1131_U123 , P2_R1131_U389 , P2_R1131_U388 , P2_R1131_U34 );
and AND2_21394 ( P2_R1131_U124 , P2_R1131_U226 , P2_R1131_U4 );
and AND2_21395 ( P2_R1131_U125 , P2_R1131_U234 , P2_R1131_U181 );
and AND2_21396 ( P2_R1131_U126 , P2_R1131_U204 , P2_R1131_U6 );
and AND2_21397 ( P2_R1131_U127 , P2_R1131_U239 , P2_R1131_U171 );
and AND2_21398 ( P2_R1131_U128 , P2_R1131_U250 , P2_R1131_U7 );
and AND2_21399 ( P2_R1131_U129 , P2_R1131_U248 , P2_R1131_U172 );
and AND2_21400 ( P2_R1131_U130 , P2_R1131_U268 , P2_R1131_U267 );
and AND2_21401 ( P2_R1131_U131 , P2_R1131_U9 , P2_R1131_U282 );
and AND2_21402 ( P2_R1131_U132 , P2_R1131_U285 , P2_R1131_U280 );
and AND2_21403 ( P2_R1131_U133 , P2_R1131_U301 , P2_R1131_U298 );
and AND2_21404 ( P2_R1131_U134 , P2_R1131_U368 , P2_R1131_U302 );
and AND2_21405 ( P2_R1131_U135 , P2_R1131_U160 , P2_R1131_U278 );
and AND3_21406 ( P2_R1131_U136 , P2_R1131_U455 , P2_R1131_U454 , P2_R1131_U80 );
and AND2_21407 ( P2_R1131_U137 , P2_R1131_U325 , P2_R1131_U9 );
and AND3_21408 ( P2_R1131_U138 , P2_R1131_U469 , P2_R1131_U468 , P2_R1131_U59 );
and AND2_21409 ( P2_R1131_U139 , P2_R1131_U334 , P2_R1131_U8 );
and AND3_21410 ( P2_R1131_U140 , P2_R1131_U490 , P2_R1131_U489 , P2_R1131_U172 );
and AND2_21411 ( P2_R1131_U141 , P2_R1131_U343 , P2_R1131_U7 );
and AND3_21412 ( P2_R1131_U142 , P2_R1131_U502 , P2_R1131_U501 , P2_R1131_U171 );
and AND2_21413 ( P2_R1131_U143 , P2_R1131_U350 , P2_R1131_U6 );
nand NAND2_21414 ( P2_R1131_U144 , P2_R1131_U118 , P2_R1131_U202 );
nand NAND2_21415 ( P2_R1131_U145 , P2_R1131_U217 , P2_R1131_U229 );
not NOT1_21416 ( P2_R1131_U146 , P2_U3057 );
not NOT1_21417 ( P2_R1131_U147 , P2_U3960 );
and AND2_21418 ( P2_R1131_U148 , P2_R1131_U403 , P2_R1131_U402 );
nand NAND3_21419 ( P2_R1131_U149 , P2_R1131_U304 , P2_R1131_U169 , P2_R1131_U364 );
and AND2_21420 ( P2_R1131_U150 , P2_R1131_U410 , P2_R1131_U409 );
nand NAND3_21421 ( P2_R1131_U151 , P2_R1131_U370 , P2_R1131_U369 , P2_R1131_U134 );
and AND2_21422 ( P2_R1131_U152 , P2_R1131_U417 , P2_R1131_U416 );
nand NAND3_21423 ( P2_R1131_U153 , P2_R1131_U365 , P2_R1131_U299 , P2_R1131_U86 );
and AND2_21424 ( P2_R1131_U154 , P2_R1131_U424 , P2_R1131_U423 );
nand NAND2_21425 ( P2_R1131_U155 , P2_R1131_U293 , P2_R1131_U292 );
and AND2_21426 ( P2_R1131_U156 , P2_R1131_U436 , P2_R1131_U435 );
nand NAND2_21427 ( P2_R1131_U157 , P2_R1131_U289 , P2_R1131_U288 );
and AND2_21428 ( P2_R1131_U158 , P2_R1131_U443 , P2_R1131_U442 );
nand NAND2_21429 ( P2_R1131_U159 , P2_R1131_U132 , P2_R1131_U284 );
and AND2_21430 ( P2_R1131_U160 , P2_R1131_U450 , P2_R1131_U449 );
nand NAND2_21431 ( P2_R1131_U161 , P2_R1131_U43 , P2_R1131_U327 );
nand NAND2_21432 ( P2_R1131_U162 , P2_R1131_U130 , P2_R1131_U269 );
and AND2_21433 ( P2_R1131_U163 , P2_R1131_U476 , P2_R1131_U475 );
nand NAND2_21434 ( P2_R1131_U164 , P2_R1131_U257 , P2_R1131_U256 );
and AND2_21435 ( P2_R1131_U165 , P2_R1131_U483 , P2_R1131_U482 );
nand NAND2_21436 ( P2_R1131_U166 , P2_R1131_U253 , P2_R1131_U252 );
nand NAND2_21437 ( P2_R1131_U167 , P2_R1131_U243 , P2_R1131_U242 );
nand NAND2_21438 ( P2_R1131_U168 , P2_R1131_U367 , P2_R1131_U366 );
nand NAND2_21439 ( P2_R1131_U169 , P2_U3056 , P2_R1131_U151 );
not NOT1_21440 ( P2_R1131_U170 , P2_R1131_U34 );
nand NAND2_21441 ( P2_R1131_U171 , P2_U3456 , P2_U3085 );
nand NAND2_21442 ( P2_R1131_U172 , P2_U3074 , P2_U3465 );
nand NAND2_21443 ( P2_R1131_U173 , P2_U3060 , P2_U3952 );
not NOT1_21444 ( P2_R1131_U174 , P2_R1131_U68 );
not NOT1_21445 ( P2_R1131_U175 , P2_R1131_U77 );
nand NAND2_21446 ( P2_R1131_U176 , P2_U3067 , P2_U3953 );
not NOT1_21447 ( P2_R1131_U177 , P2_R1131_U61 );
or OR2_21448 ( P2_R1131_U178 , P2_U3069 , P2_U3444 );
or OR2_21449 ( P2_R1131_U179 , P2_U3062 , P2_U3441 );
or OR2_21450 ( P2_R1131_U180 , P2_U3438 , P2_U3066 );
or OR2_21451 ( P2_R1131_U181 , P2_U3435 , P2_U3070 );
not NOT1_21452 ( P2_R1131_U182 , P2_R1131_U31 );
or OR2_21453 ( P2_R1131_U183 , P2_U3432 , P2_U3080 );
not NOT1_21454 ( P2_R1131_U184 , P2_R1131_U42 );
not NOT1_21455 ( P2_R1131_U185 , P2_R1131_U43 );
nand NAND2_21456 ( P2_R1131_U186 , P2_R1131_U42 , P2_R1131_U43 );
nand NAND2_21457 ( P2_R1131_U187 , P2_U3070 , P2_U3435 );
nand NAND2_21458 ( P2_R1131_U188 , P2_R1131_U186 , P2_R1131_U181 );
nand NAND2_21459 ( P2_R1131_U189 , P2_U3066 , P2_U3438 );
nand NAND2_21460 ( P2_R1131_U190 , P2_R1131_U115 , P2_R1131_U188 );
nand NAND2_21461 ( P2_R1131_U191 , P2_R1131_U35 , P2_R1131_U34 );
nand NAND2_21462 ( P2_R1131_U192 , P2_U3069 , P2_R1131_U191 );
nand NAND2_21463 ( P2_R1131_U193 , P2_R1131_U116 , P2_R1131_U190 );
nand NAND2_21464 ( P2_R1131_U194 , P2_U3444 , P2_R1131_U170 );
not NOT1_21465 ( P2_R1131_U195 , P2_R1131_U41 );
or OR2_21466 ( P2_R1131_U196 , P2_U3072 , P2_U3450 );
or OR2_21467 ( P2_R1131_U197 , P2_U3073 , P2_U3447 );
not NOT1_21468 ( P2_R1131_U198 , P2_R1131_U22 );
nand NAND2_21469 ( P2_R1131_U199 , P2_R1131_U23 , P2_R1131_U22 );
nand NAND2_21470 ( P2_R1131_U200 , P2_U3072 , P2_R1131_U199 );
nand NAND2_21471 ( P2_R1131_U201 , P2_U3450 , P2_R1131_U198 );
nand NAND2_21472 ( P2_R1131_U202 , P2_R1131_U5 , P2_R1131_U41 );
not NOT1_21473 ( P2_R1131_U203 , P2_R1131_U144 );
or OR2_21474 ( P2_R1131_U204 , P2_U3453 , P2_U3086 );
nand NAND2_21475 ( P2_R1131_U205 , P2_R1131_U204 , P2_R1131_U144 );
not NOT1_21476 ( P2_R1131_U206 , P2_R1131_U40 );
or OR2_21477 ( P2_R1131_U207 , P2_U3085 , P2_U3456 );
or OR2_21478 ( P2_R1131_U208 , P2_U3447 , P2_U3073 );
nand NAND2_21479 ( P2_R1131_U209 , P2_R1131_U208 , P2_R1131_U41 );
nand NAND2_21480 ( P2_R1131_U210 , P2_R1131_U119 , P2_R1131_U209 );
nand NAND2_21481 ( P2_R1131_U211 , P2_R1131_U195 , P2_R1131_U22 );
nand NAND2_21482 ( P2_R1131_U212 , P2_U3450 , P2_U3072 );
nand NAND2_21483 ( P2_R1131_U213 , P2_R1131_U120 , P2_R1131_U211 );
or OR2_21484 ( P2_R1131_U214 , P2_U3073 , P2_U3447 );
nand NAND2_21485 ( P2_R1131_U215 , P2_R1131_U185 , P2_R1131_U181 );
nand NAND2_21486 ( P2_R1131_U216 , P2_U3070 , P2_U3435 );
not NOT1_21487 ( P2_R1131_U217 , P2_R1131_U45 );
nand NAND2_21488 ( P2_R1131_U218 , P2_R1131_U121 , P2_R1131_U184 );
nand NAND2_21489 ( P2_R1131_U219 , P2_R1131_U45 , P2_R1131_U180 );
nand NAND2_21490 ( P2_R1131_U220 , P2_U3066 , P2_U3438 );
not NOT1_21491 ( P2_R1131_U221 , P2_R1131_U44 );
or OR2_21492 ( P2_R1131_U222 , P2_U3441 , P2_U3062 );
nand NAND2_21493 ( P2_R1131_U223 , P2_R1131_U222 , P2_R1131_U44 );
nand NAND2_21494 ( P2_R1131_U224 , P2_R1131_U123 , P2_R1131_U223 );
nand NAND2_21495 ( P2_R1131_U225 , P2_R1131_U221 , P2_R1131_U34 );
nand NAND2_21496 ( P2_R1131_U226 , P2_U3444 , P2_U3069 );
nand NAND2_21497 ( P2_R1131_U227 , P2_R1131_U124 , P2_R1131_U225 );
or OR2_21498 ( P2_R1131_U228 , P2_U3062 , P2_U3441 );
nand NAND2_21499 ( P2_R1131_U229 , P2_R1131_U184 , P2_R1131_U181 );
not NOT1_21500 ( P2_R1131_U230 , P2_R1131_U145 );
nand NAND2_21501 ( P2_R1131_U231 , P2_U3066 , P2_U3438 );
nand NAND4_21502 ( P2_R1131_U232 , P2_R1131_U401 , P2_R1131_U400 , P2_R1131_U43 , P2_R1131_U42 );
nand NAND2_21503 ( P2_R1131_U233 , P2_R1131_U43 , P2_R1131_U42 );
nand NAND2_21504 ( P2_R1131_U234 , P2_U3070 , P2_U3435 );
nand NAND2_21505 ( P2_R1131_U235 , P2_R1131_U125 , P2_R1131_U233 );
or OR2_21506 ( P2_R1131_U236 , P2_U3085 , P2_U3456 );
or OR2_21507 ( P2_R1131_U237 , P2_U3064 , P2_U3459 );
nand NAND2_21508 ( P2_R1131_U238 , P2_R1131_U177 , P2_R1131_U6 );
nand NAND2_21509 ( P2_R1131_U239 , P2_U3064 , P2_U3459 );
nand NAND2_21510 ( P2_R1131_U240 , P2_R1131_U127 , P2_R1131_U238 );
or OR2_21511 ( P2_R1131_U241 , P2_U3459 , P2_U3064 );
nand NAND2_21512 ( P2_R1131_U242 , P2_R1131_U126 , P2_R1131_U144 );
nand NAND2_21513 ( P2_R1131_U243 , P2_R1131_U241 , P2_R1131_U240 );
not NOT1_21514 ( P2_R1131_U244 , P2_R1131_U167 );
or OR2_21515 ( P2_R1131_U245 , P2_U3082 , P2_U3468 );
or OR2_21516 ( P2_R1131_U246 , P2_U3074 , P2_U3465 );
nand NAND2_21517 ( P2_R1131_U247 , P2_R1131_U174 , P2_R1131_U7 );
nand NAND2_21518 ( P2_R1131_U248 , P2_U3082 , P2_U3468 );
nand NAND2_21519 ( P2_R1131_U249 , P2_R1131_U129 , P2_R1131_U247 );
or OR2_21520 ( P2_R1131_U250 , P2_U3462 , P2_U3065 );
or OR2_21521 ( P2_R1131_U251 , P2_U3468 , P2_U3082 );
nand NAND2_21522 ( P2_R1131_U252 , P2_R1131_U128 , P2_R1131_U167 );
nand NAND2_21523 ( P2_R1131_U253 , P2_R1131_U251 , P2_R1131_U249 );
not NOT1_21524 ( P2_R1131_U254 , P2_R1131_U166 );
or OR2_21525 ( P2_R1131_U255 , P2_U3471 , P2_U3081 );
nand NAND2_21526 ( P2_R1131_U256 , P2_R1131_U255 , P2_R1131_U166 );
nand NAND2_21527 ( P2_R1131_U257 , P2_U3081 , P2_U3471 );
not NOT1_21528 ( P2_R1131_U258 , P2_R1131_U164 );
or OR2_21529 ( P2_R1131_U259 , P2_U3474 , P2_U3076 );
nand NAND2_21530 ( P2_R1131_U260 , P2_R1131_U259 , P2_R1131_U164 );
nand NAND2_21531 ( P2_R1131_U261 , P2_U3076 , P2_U3474 );
not NOT1_21532 ( P2_R1131_U262 , P2_R1131_U92 );
or OR2_21533 ( P2_R1131_U263 , P2_U3071 , P2_U3480 );
or OR2_21534 ( P2_R1131_U264 , P2_U3075 , P2_U3477 );
not NOT1_21535 ( P2_R1131_U265 , P2_R1131_U59 );
nand NAND2_21536 ( P2_R1131_U266 , P2_R1131_U60 , P2_R1131_U59 );
nand NAND2_21537 ( P2_R1131_U267 , P2_U3071 , P2_R1131_U266 );
nand NAND2_21538 ( P2_R1131_U268 , P2_U3480 , P2_R1131_U265 );
nand NAND2_21539 ( P2_R1131_U269 , P2_R1131_U8 , P2_R1131_U92 );
not NOT1_21540 ( P2_R1131_U270 , P2_R1131_U162 );
or OR2_21541 ( P2_R1131_U271 , P2_U3078 , P2_U3957 );
or OR2_21542 ( P2_R1131_U272 , P2_U3083 , P2_U3485 );
or OR2_21543 ( P2_R1131_U273 , P2_U3077 , P2_U3956 );
not NOT1_21544 ( P2_R1131_U274 , P2_R1131_U80 );
nand NAND2_21545 ( P2_R1131_U275 , P2_U3957 , P2_R1131_U274 );
nand NAND2_21546 ( P2_R1131_U276 , P2_R1131_U275 , P2_R1131_U90 );
nand NAND2_21547 ( P2_R1131_U277 , P2_R1131_U80 , P2_R1131_U81 );
nand NAND2_21548 ( P2_R1131_U278 , P2_R1131_U277 , P2_R1131_U276 );
nand NAND2_21549 ( P2_R1131_U279 , P2_R1131_U175 , P2_R1131_U9 );
nand NAND2_21550 ( P2_R1131_U280 , P2_U3077 , P2_U3956 );
nand NAND2_21551 ( P2_R1131_U281 , P2_R1131_U278 , P2_R1131_U279 );
or OR2_21552 ( P2_R1131_U282 , P2_U3483 , P2_U3084 );
or OR2_21553 ( P2_R1131_U283 , P2_U3956 , P2_U3077 );
nand NAND3_21554 ( P2_R1131_U284 , P2_R1131_U273 , P2_R1131_U162 , P2_R1131_U131 );
nand NAND2_21555 ( P2_R1131_U285 , P2_R1131_U283 , P2_R1131_U281 );
not NOT1_21556 ( P2_R1131_U286 , P2_R1131_U159 );
or OR2_21557 ( P2_R1131_U287 , P2_U3955 , P2_U3063 );
nand NAND2_21558 ( P2_R1131_U288 , P2_R1131_U287 , P2_R1131_U159 );
nand NAND2_21559 ( P2_R1131_U289 , P2_U3063 , P2_U3955 );
not NOT1_21560 ( P2_R1131_U290 , P2_R1131_U157 );
or OR2_21561 ( P2_R1131_U291 , P2_U3954 , P2_U3068 );
nand NAND2_21562 ( P2_R1131_U292 , P2_R1131_U291 , P2_R1131_U157 );
nand NAND2_21563 ( P2_R1131_U293 , P2_U3068 , P2_U3954 );
not NOT1_21564 ( P2_R1131_U294 , P2_R1131_U155 );
or OR2_21565 ( P2_R1131_U295 , P2_U3060 , P2_U3952 );
nand NAND2_21566 ( P2_R1131_U296 , P2_R1131_U176 , P2_R1131_U173 );
not NOT1_21567 ( P2_R1131_U297 , P2_R1131_U86 );
or OR2_21568 ( P2_R1131_U298 , P2_U3953 , P2_U3067 );
nand NAND3_21569 ( P2_R1131_U299 , P2_R1131_U155 , P2_R1131_U298 , P2_R1131_U168 );
not NOT1_21570 ( P2_R1131_U300 , P2_R1131_U153 );
or OR2_21571 ( P2_R1131_U301 , P2_U3950 , P2_U3055 );
nand NAND2_21572 ( P2_R1131_U302 , P2_U3055 , P2_U3950 );
not NOT1_21573 ( P2_R1131_U303 , P2_R1131_U151 );
nand NAND2_21574 ( P2_R1131_U304 , P2_U3949 , P2_R1131_U151 );
not NOT1_21575 ( P2_R1131_U305 , P2_R1131_U149 );
nand NAND2_21576 ( P2_R1131_U306 , P2_R1131_U298 , P2_R1131_U155 );
not NOT1_21577 ( P2_R1131_U307 , P2_R1131_U89 );
or OR2_21578 ( P2_R1131_U308 , P2_U3952 , P2_U3060 );
nand NAND2_21579 ( P2_R1131_U309 , P2_R1131_U308 , P2_R1131_U89 );
nand NAND3_21580 ( P2_R1131_U310 , P2_R1131_U309 , P2_R1131_U173 , P2_R1131_U154 );
nand NAND2_21581 ( P2_R1131_U311 , P2_R1131_U307 , P2_R1131_U173 );
nand NAND2_21582 ( P2_R1131_U312 , P2_U3951 , P2_U3059 );
nand NAND3_21583 ( P2_R1131_U313 , P2_R1131_U311 , P2_R1131_U312 , P2_R1131_U168 );
or OR2_21584 ( P2_R1131_U314 , P2_U3060 , P2_U3952 );
nand NAND2_21585 ( P2_R1131_U315 , P2_R1131_U282 , P2_R1131_U162 );
not NOT1_21586 ( P2_R1131_U316 , P2_R1131_U91 );
nand NAND2_21587 ( P2_R1131_U317 , P2_R1131_U9 , P2_R1131_U91 );
nand NAND2_21588 ( P2_R1131_U318 , P2_R1131_U135 , P2_R1131_U317 );
nand NAND2_21589 ( P2_R1131_U319 , P2_R1131_U317 , P2_R1131_U278 );
nand NAND2_21590 ( P2_R1131_U320 , P2_R1131_U453 , P2_R1131_U319 );
or OR2_21591 ( P2_R1131_U321 , P2_U3485 , P2_U3083 );
nand NAND2_21592 ( P2_R1131_U322 , P2_R1131_U321 , P2_R1131_U91 );
nand NAND2_21593 ( P2_R1131_U323 , P2_R1131_U136 , P2_R1131_U322 );
nand NAND2_21594 ( P2_R1131_U324 , P2_R1131_U316 , P2_R1131_U80 );
nand NAND2_21595 ( P2_R1131_U325 , P2_U3078 , P2_U3957 );
nand NAND2_21596 ( P2_R1131_U326 , P2_R1131_U137 , P2_R1131_U324 );
or OR2_21597 ( P2_R1131_U327 , P2_U3432 , P2_U3080 );
not NOT1_21598 ( P2_R1131_U328 , P2_R1131_U161 );
or OR2_21599 ( P2_R1131_U329 , P2_U3083 , P2_U3485 );
or OR2_21600 ( P2_R1131_U330 , P2_U3477 , P2_U3075 );
nand NAND2_21601 ( P2_R1131_U331 , P2_R1131_U330 , P2_R1131_U92 );
nand NAND2_21602 ( P2_R1131_U332 , P2_R1131_U138 , P2_R1131_U331 );
nand NAND2_21603 ( P2_R1131_U333 , P2_R1131_U262 , P2_R1131_U59 );
nand NAND2_21604 ( P2_R1131_U334 , P2_U3480 , P2_U3071 );
nand NAND2_21605 ( P2_R1131_U335 , P2_R1131_U139 , P2_R1131_U333 );
or OR2_21606 ( P2_R1131_U336 , P2_U3075 , P2_U3477 );
nand NAND2_21607 ( P2_R1131_U337 , P2_R1131_U250 , P2_R1131_U167 );
not NOT1_21608 ( P2_R1131_U338 , P2_R1131_U93 );
or OR2_21609 ( P2_R1131_U339 , P2_U3465 , P2_U3074 );
nand NAND2_21610 ( P2_R1131_U340 , P2_R1131_U339 , P2_R1131_U93 );
nand NAND2_21611 ( P2_R1131_U341 , P2_R1131_U140 , P2_R1131_U340 );
nand NAND2_21612 ( P2_R1131_U342 , P2_R1131_U338 , P2_R1131_U172 );
nand NAND2_21613 ( P2_R1131_U343 , P2_U3082 , P2_U3468 );
nand NAND2_21614 ( P2_R1131_U344 , P2_R1131_U141 , P2_R1131_U342 );
or OR2_21615 ( P2_R1131_U345 , P2_U3074 , P2_U3465 );
or OR2_21616 ( P2_R1131_U346 , P2_U3456 , P2_U3085 );
nand NAND2_21617 ( P2_R1131_U347 , P2_R1131_U346 , P2_R1131_U40 );
nand NAND2_21618 ( P2_R1131_U348 , P2_R1131_U142 , P2_R1131_U347 );
nand NAND2_21619 ( P2_R1131_U349 , P2_R1131_U206 , P2_R1131_U171 );
nand NAND2_21620 ( P2_R1131_U350 , P2_U3064 , P2_U3459 );
nand NAND2_21621 ( P2_R1131_U351 , P2_R1131_U143 , P2_R1131_U349 );
nand NAND2_21622 ( P2_R1131_U352 , P2_R1131_U207 , P2_R1131_U171 );
nand NAND2_21623 ( P2_R1131_U353 , P2_R1131_U204 , P2_R1131_U61 );
nand NAND2_21624 ( P2_R1131_U354 , P2_R1131_U214 , P2_R1131_U22 );
nand NAND2_21625 ( P2_R1131_U355 , P2_R1131_U228 , P2_R1131_U34 );
nand NAND2_21626 ( P2_R1131_U356 , P2_R1131_U231 , P2_R1131_U180 );
nand NAND2_21627 ( P2_R1131_U357 , P2_R1131_U314 , P2_R1131_U173 );
nand NAND2_21628 ( P2_R1131_U358 , P2_R1131_U298 , P2_R1131_U176 );
nand NAND2_21629 ( P2_R1131_U359 , P2_R1131_U329 , P2_R1131_U80 );
nand NAND2_21630 ( P2_R1131_U360 , P2_R1131_U282 , P2_R1131_U77 );
nand NAND2_21631 ( P2_R1131_U361 , P2_R1131_U336 , P2_R1131_U59 );
nand NAND2_21632 ( P2_R1131_U362 , P2_R1131_U345 , P2_R1131_U172 );
nand NAND2_21633 ( P2_R1131_U363 , P2_R1131_U250 , P2_R1131_U68 );
nand NAND2_21634 ( P2_R1131_U364 , P2_U3949 , P2_U3056 );
nand NAND2_21635 ( P2_R1131_U365 , P2_R1131_U296 , P2_R1131_U168 );
nand NAND2_21636 ( P2_R1131_U366 , P2_U3059 , P2_R1131_U295 );
nand NAND2_21637 ( P2_R1131_U367 , P2_U3951 , P2_R1131_U295 );
nand NAND3_21638 ( P2_R1131_U368 , P2_R1131_U296 , P2_R1131_U168 , P2_R1131_U301 );
nand NAND3_21639 ( P2_R1131_U369 , P2_R1131_U155 , P2_R1131_U168 , P2_R1131_U133 );
nand NAND2_21640 ( P2_R1131_U370 , P2_R1131_U297 , P2_R1131_U301 );
nand NAND2_21641 ( P2_R1131_U371 , P2_U3085 , P2_R1131_U39 );
nand NAND2_21642 ( P2_R1131_U372 , P2_U3456 , P2_R1131_U38 );
nand NAND2_21643 ( P2_R1131_U373 , P2_R1131_U372 , P2_R1131_U371 );
nand NAND2_21644 ( P2_R1131_U374 , P2_R1131_U352 , P2_R1131_U40 );
nand NAND2_21645 ( P2_R1131_U375 , P2_R1131_U373 , P2_R1131_U206 );
nand NAND2_21646 ( P2_R1131_U376 , P2_U3086 , P2_R1131_U36 );
nand NAND2_21647 ( P2_R1131_U377 , P2_U3453 , P2_R1131_U37 );
nand NAND2_21648 ( P2_R1131_U378 , P2_R1131_U377 , P2_R1131_U376 );
nand NAND2_21649 ( P2_R1131_U379 , P2_R1131_U353 , P2_R1131_U144 );
nand NAND2_21650 ( P2_R1131_U380 , P2_R1131_U203 , P2_R1131_U378 );
nand NAND2_21651 ( P2_R1131_U381 , P2_U3072 , P2_R1131_U23 );
nand NAND2_21652 ( P2_R1131_U382 , P2_U3450 , P2_R1131_U21 );
nand NAND2_21653 ( P2_R1131_U383 , P2_U3073 , P2_R1131_U19 );
nand NAND2_21654 ( P2_R1131_U384 , P2_U3447 , P2_R1131_U20 );
nand NAND2_21655 ( P2_R1131_U385 , P2_R1131_U384 , P2_R1131_U383 );
nand NAND2_21656 ( P2_R1131_U386 , P2_R1131_U354 , P2_R1131_U41 );
nand NAND2_21657 ( P2_R1131_U387 , P2_R1131_U385 , P2_R1131_U195 );
nand NAND2_21658 ( P2_R1131_U388 , P2_U3069 , P2_R1131_U35 );
nand NAND2_21659 ( P2_R1131_U389 , P2_U3444 , P2_R1131_U26 );
nand NAND2_21660 ( P2_R1131_U390 , P2_U3062 , P2_R1131_U24 );
nand NAND2_21661 ( P2_R1131_U391 , P2_U3441 , P2_R1131_U25 );
nand NAND2_21662 ( P2_R1131_U392 , P2_R1131_U391 , P2_R1131_U390 );
nand NAND2_21663 ( P2_R1131_U393 , P2_R1131_U355 , P2_R1131_U44 );
nand NAND2_21664 ( P2_R1131_U394 , P2_R1131_U392 , P2_R1131_U221 );
nand NAND2_21665 ( P2_R1131_U395 , P2_U3066 , P2_R1131_U32 );
nand NAND2_21666 ( P2_R1131_U396 , P2_U3438 , P2_R1131_U33 );
nand NAND2_21667 ( P2_R1131_U397 , P2_R1131_U396 , P2_R1131_U395 );
nand NAND2_21668 ( P2_R1131_U398 , P2_R1131_U356 , P2_R1131_U145 );
nand NAND2_21669 ( P2_R1131_U399 , P2_R1131_U230 , P2_R1131_U397 );
nand NAND2_21670 ( P2_R1131_U400 , P2_U3070 , P2_R1131_U27 );
nand NAND2_21671 ( P2_R1131_U401 , P2_U3435 , P2_R1131_U28 );
nand NAND2_21672 ( P2_R1131_U402 , P2_U3057 , P2_R1131_U147 );
nand NAND2_21673 ( P2_R1131_U403 , P2_U3960 , P2_R1131_U146 );
nand NAND2_21674 ( P2_R1131_U404 , P2_U3057 , P2_R1131_U147 );
nand NAND2_21675 ( P2_R1131_U405 , P2_U3960 , P2_R1131_U146 );
nand NAND2_21676 ( P2_R1131_U406 , P2_R1131_U405 , P2_R1131_U404 );
nand NAND2_21677 ( P2_R1131_U407 , P2_R1131_U148 , P2_R1131_U149 );
nand NAND2_21678 ( P2_R1131_U408 , P2_R1131_U305 , P2_R1131_U406 );
nand NAND2_21679 ( P2_R1131_U409 , P2_U3056 , P2_R1131_U88 );
nand NAND2_21680 ( P2_R1131_U410 , P2_U3949 , P2_R1131_U87 );
nand NAND2_21681 ( P2_R1131_U411 , P2_U3056 , P2_R1131_U88 );
nand NAND2_21682 ( P2_R1131_U412 , P2_U3949 , P2_R1131_U87 );
nand NAND2_21683 ( P2_R1131_U413 , P2_R1131_U412 , P2_R1131_U411 );
nand NAND2_21684 ( P2_R1131_U414 , P2_R1131_U150 , P2_R1131_U151 );
nand NAND2_21685 ( P2_R1131_U415 , P2_R1131_U303 , P2_R1131_U413 );
nand NAND2_21686 ( P2_R1131_U416 , P2_U3055 , P2_R1131_U46 );
nand NAND2_21687 ( P2_R1131_U417 , P2_U3950 , P2_R1131_U47 );
nand NAND2_21688 ( P2_R1131_U418 , P2_U3055 , P2_R1131_U46 );
nand NAND2_21689 ( P2_R1131_U419 , P2_U3950 , P2_R1131_U47 );
nand NAND2_21690 ( P2_R1131_U420 , P2_R1131_U419 , P2_R1131_U418 );
nand NAND2_21691 ( P2_R1131_U421 , P2_R1131_U152 , P2_R1131_U153 );
nand NAND2_21692 ( P2_R1131_U422 , P2_R1131_U300 , P2_R1131_U420 );
nand NAND2_21693 ( P2_R1131_U423 , P2_U3059 , P2_R1131_U49 );
nand NAND2_21694 ( P2_R1131_U424 , P2_U3951 , P2_R1131_U48 );
nand NAND2_21695 ( P2_R1131_U425 , P2_U3060 , P2_R1131_U50 );
nand NAND2_21696 ( P2_R1131_U426 , P2_U3952 , P2_R1131_U51 );
nand NAND2_21697 ( P2_R1131_U427 , P2_R1131_U426 , P2_R1131_U425 );
nand NAND2_21698 ( P2_R1131_U428 , P2_R1131_U357 , P2_R1131_U89 );
nand NAND2_21699 ( P2_R1131_U429 , P2_R1131_U427 , P2_R1131_U307 );
nand NAND2_21700 ( P2_R1131_U430 , P2_U3067 , P2_R1131_U52 );
nand NAND2_21701 ( P2_R1131_U431 , P2_U3953 , P2_R1131_U53 );
nand NAND2_21702 ( P2_R1131_U432 , P2_R1131_U431 , P2_R1131_U430 );
nand NAND2_21703 ( P2_R1131_U433 , P2_R1131_U358 , P2_R1131_U155 );
nand NAND2_21704 ( P2_R1131_U434 , P2_R1131_U294 , P2_R1131_U432 );
nand NAND2_21705 ( P2_R1131_U435 , P2_U3068 , P2_R1131_U84 );
nand NAND2_21706 ( P2_R1131_U436 , P2_U3954 , P2_R1131_U85 );
nand NAND2_21707 ( P2_R1131_U437 , P2_U3068 , P2_R1131_U84 );
nand NAND2_21708 ( P2_R1131_U438 , P2_U3954 , P2_R1131_U85 );
nand NAND2_21709 ( P2_R1131_U439 , P2_R1131_U438 , P2_R1131_U437 );
nand NAND2_21710 ( P2_R1131_U440 , P2_R1131_U156 , P2_R1131_U157 );
nand NAND2_21711 ( P2_R1131_U441 , P2_R1131_U290 , P2_R1131_U439 );
nand NAND2_21712 ( P2_R1131_U442 , P2_U3063 , P2_R1131_U82 );
nand NAND2_21713 ( P2_R1131_U443 , P2_U3955 , P2_R1131_U83 );
nand NAND2_21714 ( P2_R1131_U444 , P2_U3063 , P2_R1131_U82 );
nand NAND2_21715 ( P2_R1131_U445 , P2_U3955 , P2_R1131_U83 );
nand NAND2_21716 ( P2_R1131_U446 , P2_R1131_U445 , P2_R1131_U444 );
nand NAND2_21717 ( P2_R1131_U447 , P2_R1131_U158 , P2_R1131_U159 );
nand NAND2_21718 ( P2_R1131_U448 , P2_R1131_U286 , P2_R1131_U446 );
nand NAND2_21719 ( P2_R1131_U449 , P2_U3077 , P2_R1131_U54 );
nand NAND2_21720 ( P2_R1131_U450 , P2_U3956 , P2_R1131_U55 );
nand NAND2_21721 ( P2_R1131_U451 , P2_U3077 , P2_R1131_U54 );
nand NAND2_21722 ( P2_R1131_U452 , P2_U3956 , P2_R1131_U55 );
nand NAND2_21723 ( P2_R1131_U453 , P2_R1131_U452 , P2_R1131_U451 );
nand NAND2_21724 ( P2_R1131_U454 , P2_U3078 , P2_R1131_U81 );
nand NAND2_21725 ( P2_R1131_U455 , P2_U3957 , P2_R1131_U90 );
nand NAND2_21726 ( P2_R1131_U456 , P2_R1131_U182 , P2_R1131_U161 );
nand NAND2_21727 ( P2_R1131_U457 , P2_R1131_U328 , P2_R1131_U31 );
nand NAND2_21728 ( P2_R1131_U458 , P2_U3083 , P2_R1131_U78 );
nand NAND2_21729 ( P2_R1131_U459 , P2_U3485 , P2_R1131_U79 );
nand NAND2_21730 ( P2_R1131_U460 , P2_R1131_U459 , P2_R1131_U458 );
nand NAND2_21731 ( P2_R1131_U461 , P2_R1131_U359 , P2_R1131_U91 );
nand NAND2_21732 ( P2_R1131_U462 , P2_R1131_U460 , P2_R1131_U316 );
nand NAND2_21733 ( P2_R1131_U463 , P2_U3084 , P2_R1131_U75 );
nand NAND2_21734 ( P2_R1131_U464 , P2_U3483 , P2_R1131_U76 );
nand NAND2_21735 ( P2_R1131_U465 , P2_R1131_U464 , P2_R1131_U463 );
nand NAND2_21736 ( P2_R1131_U466 , P2_R1131_U360 , P2_R1131_U162 );
nand NAND2_21737 ( P2_R1131_U467 , P2_R1131_U270 , P2_R1131_U465 );
nand NAND2_21738 ( P2_R1131_U468 , P2_U3071 , P2_R1131_U60 );
nand NAND2_21739 ( P2_R1131_U469 , P2_U3480 , P2_R1131_U58 );
nand NAND2_21740 ( P2_R1131_U470 , P2_U3075 , P2_R1131_U56 );
nand NAND2_21741 ( P2_R1131_U471 , P2_U3477 , P2_R1131_U57 );
nand NAND2_21742 ( P2_R1131_U472 , P2_R1131_U471 , P2_R1131_U470 );
nand NAND2_21743 ( P2_R1131_U473 , P2_R1131_U361 , P2_R1131_U92 );
nand NAND2_21744 ( P2_R1131_U474 , P2_R1131_U472 , P2_R1131_U262 );
nand NAND2_21745 ( P2_R1131_U475 , P2_U3076 , P2_R1131_U73 );
nand NAND2_21746 ( P2_R1131_U476 , P2_U3474 , P2_R1131_U74 );
nand NAND2_21747 ( P2_R1131_U477 , P2_U3076 , P2_R1131_U73 );
nand NAND2_21748 ( P2_R1131_U478 , P2_U3474 , P2_R1131_U74 );
nand NAND2_21749 ( P2_R1131_U479 , P2_R1131_U478 , P2_R1131_U477 );
nand NAND2_21750 ( P2_R1131_U480 , P2_R1131_U163 , P2_R1131_U164 );
nand NAND2_21751 ( P2_R1131_U481 , P2_R1131_U258 , P2_R1131_U479 );
nand NAND2_21752 ( P2_R1131_U482 , P2_U3081 , P2_R1131_U71 );
nand NAND2_21753 ( P2_R1131_U483 , P2_U3471 , P2_R1131_U72 );
nand NAND2_21754 ( P2_R1131_U484 , P2_U3081 , P2_R1131_U71 );
nand NAND2_21755 ( P2_R1131_U485 , P2_U3471 , P2_R1131_U72 );
nand NAND2_21756 ( P2_R1131_U486 , P2_R1131_U485 , P2_R1131_U484 );
nand NAND2_21757 ( P2_R1131_U487 , P2_R1131_U165 , P2_R1131_U166 );
nand NAND2_21758 ( P2_R1131_U488 , P2_R1131_U254 , P2_R1131_U486 );
nand NAND2_21759 ( P2_R1131_U489 , P2_U3082 , P2_R1131_U69 );
nand NAND2_21760 ( P2_R1131_U490 , P2_U3468 , P2_R1131_U70 );
nand NAND2_21761 ( P2_R1131_U491 , P2_U3074 , P2_R1131_U64 );
nand NAND2_21762 ( P2_R1131_U492 , P2_U3465 , P2_R1131_U65 );
nand NAND2_21763 ( P2_R1131_U493 , P2_R1131_U492 , P2_R1131_U491 );
nand NAND2_21764 ( P2_R1131_U494 , P2_R1131_U362 , P2_R1131_U93 );
nand NAND2_21765 ( P2_R1131_U495 , P2_R1131_U493 , P2_R1131_U338 );
nand NAND2_21766 ( P2_R1131_U496 , P2_U3065 , P2_R1131_U66 );
nand NAND2_21767 ( P2_R1131_U497 , P2_U3462 , P2_R1131_U67 );
nand NAND2_21768 ( P2_R1131_U498 , P2_R1131_U497 , P2_R1131_U496 );
nand NAND2_21769 ( P2_R1131_U499 , P2_R1131_U363 , P2_R1131_U167 );
nand NAND2_21770 ( P2_R1131_U500 , P2_R1131_U244 , P2_R1131_U498 );
nand NAND2_21771 ( P2_R1131_U501 , P2_U3064 , P2_R1131_U62 );
nand NAND2_21772 ( P2_R1131_U502 , P2_U3459 , P2_R1131_U63 );
nand NAND2_21773 ( P2_R1131_U503 , P2_U3079 , P2_R1131_U29 );
nand NAND2_21774 ( P2_R1131_U504 , P2_U3427 , P2_R1131_U30 );
and AND2_21775 ( P2_R1146_U6 , P2_R1146_U202 , P2_R1146_U201 );
and AND2_21776 ( P2_R1146_U7 , P2_R1146_U241 , P2_R1146_U240 );
and AND2_21777 ( P2_R1146_U8 , P2_R1146_U181 , P2_R1146_U256 );
and AND2_21778 ( P2_R1146_U9 , P2_R1146_U258 , P2_R1146_U257 );
and AND2_21779 ( P2_R1146_U10 , P2_R1146_U182 , P2_R1146_U282 );
and AND2_21780 ( P2_R1146_U11 , P2_R1146_U284 , P2_R1146_U283 );
nand NAND2_21781 ( P2_R1146_U12 , P2_R1146_U344 , P2_R1146_U347 );
nand NAND2_21782 ( P2_R1146_U13 , P2_R1146_U333 , P2_R1146_U336 );
nand NAND2_21783 ( P2_R1146_U14 , P2_R1146_U322 , P2_R1146_U325 );
nand NAND2_21784 ( P2_R1146_U15 , P2_R1146_U314 , P2_R1146_U316 );
nand NAND2_21785 ( P2_R1146_U16 , P2_R1146_U352 , P2_R1146_U312 );
nand NAND2_21786 ( P2_R1146_U17 , P2_R1146_U235 , P2_R1146_U237 );
nand NAND2_21787 ( P2_R1146_U18 , P2_R1146_U227 , P2_R1146_U230 );
nand NAND2_21788 ( P2_R1146_U19 , P2_R1146_U219 , P2_R1146_U221 );
nand NAND2_21789 ( P2_R1146_U20 , P2_R1146_U166 , P2_R1146_U350 );
not NOT1_21790 ( P2_R1146_U21 , P2_U3450 );
not NOT1_21791 ( P2_R1146_U22 , P2_U3444 );
not NOT1_21792 ( P2_R1146_U23 , P2_U3435 );
not NOT1_21793 ( P2_R1146_U24 , P2_U3427 );
not NOT1_21794 ( P2_R1146_U25 , P2_U3080 );
not NOT1_21795 ( P2_R1146_U26 , P2_U3438 );
not NOT1_21796 ( P2_R1146_U27 , P2_U3070 );
nand NAND2_21797 ( P2_R1146_U28 , P2_U3070 , P2_R1146_U23 );
not NOT1_21798 ( P2_R1146_U29 , P2_U3066 );
not NOT1_21799 ( P2_R1146_U30 , P2_U3447 );
not NOT1_21800 ( P2_R1146_U31 , P2_U3441 );
not NOT1_21801 ( P2_R1146_U32 , P2_U3073 );
not NOT1_21802 ( P2_R1146_U33 , P2_U3069 );
not NOT1_21803 ( P2_R1146_U34 , P2_U3062 );
nand NAND2_21804 ( P2_R1146_U35 , P2_U3062 , P2_R1146_U31 );
not NOT1_21805 ( P2_R1146_U36 , P2_U3453 );
not NOT1_21806 ( P2_R1146_U37 , P2_U3072 );
nand NAND2_21807 ( P2_R1146_U38 , P2_U3072 , P2_R1146_U21 );
not NOT1_21808 ( P2_R1146_U39 , P2_U3086 );
not NOT1_21809 ( P2_R1146_U40 , P2_U3456 );
not NOT1_21810 ( P2_R1146_U41 , P2_U3085 );
nand NAND2_21811 ( P2_R1146_U42 , P2_R1146_U208 , P2_R1146_U207 );
nand NAND2_21812 ( P2_R1146_U43 , P2_R1146_U35 , P2_R1146_U223 );
nand NAND3_21813 ( P2_R1146_U44 , P2_R1146_U192 , P2_R1146_U176 , P2_R1146_U351 );
not NOT1_21814 ( P2_R1146_U45 , P2_U3951 );
not NOT1_21815 ( P2_R1146_U46 , P2_U3459 );
not NOT1_21816 ( P2_R1146_U47 , P2_U3462 );
not NOT1_21817 ( P2_R1146_U48 , P2_U3065 );
not NOT1_21818 ( P2_R1146_U49 , P2_U3064 );
nand NAND2_21819 ( P2_R1146_U50 , P2_U3085 , P2_R1146_U40 );
not NOT1_21820 ( P2_R1146_U51 , P2_U3465 );
not NOT1_21821 ( P2_R1146_U52 , P2_U3074 );
not NOT1_21822 ( P2_R1146_U53 , P2_U3468 );
not NOT1_21823 ( P2_R1146_U54 , P2_U3082 );
not NOT1_21824 ( P2_R1146_U55 , P2_U3477 );
not NOT1_21825 ( P2_R1146_U56 , P2_U3474 );
not NOT1_21826 ( P2_R1146_U57 , P2_U3471 );
not NOT1_21827 ( P2_R1146_U58 , P2_U3075 );
not NOT1_21828 ( P2_R1146_U59 , P2_U3076 );
not NOT1_21829 ( P2_R1146_U60 , P2_U3081 );
nand NAND2_21830 ( P2_R1146_U61 , P2_U3081 , P2_R1146_U57 );
not NOT1_21831 ( P2_R1146_U62 , P2_U3480 );
not NOT1_21832 ( P2_R1146_U63 , P2_U3071 );
nand NAND2_21833 ( P2_R1146_U64 , P2_R1146_U268 , P2_R1146_U267 );
not NOT1_21834 ( P2_R1146_U65 , P2_U3084 );
not NOT1_21835 ( P2_R1146_U66 , P2_U3485 );
not NOT1_21836 ( P2_R1146_U67 , P2_U3083 );
not NOT1_21837 ( P2_R1146_U68 , P2_U3957 );
not NOT1_21838 ( P2_R1146_U69 , P2_U3078 );
not NOT1_21839 ( P2_R1146_U70 , P2_U3954 );
not NOT1_21840 ( P2_R1146_U71 , P2_U3955 );
not NOT1_21841 ( P2_R1146_U72 , P2_U3956 );
not NOT1_21842 ( P2_R1146_U73 , P2_U3068 );
not NOT1_21843 ( P2_R1146_U74 , P2_U3063 );
not NOT1_21844 ( P2_R1146_U75 , P2_U3077 );
nand NAND2_21845 ( P2_R1146_U76 , P2_U3077 , P2_R1146_U72 );
not NOT1_21846 ( P2_R1146_U77 , P2_U3953 );
not NOT1_21847 ( P2_R1146_U78 , P2_U3067 );
not NOT1_21848 ( P2_R1146_U79 , P2_U3952 );
not NOT1_21849 ( P2_R1146_U80 , P2_U3060 );
not NOT1_21850 ( P2_R1146_U81 , P2_U3950 );
not NOT1_21851 ( P2_R1146_U82 , P2_U3059 );
nand NAND2_21852 ( P2_R1146_U83 , P2_U3059 , P2_R1146_U45 );
not NOT1_21853 ( P2_R1146_U84 , P2_U3055 );
not NOT1_21854 ( P2_R1146_U85 , P2_U3949 );
not NOT1_21855 ( P2_R1146_U86 , P2_U3056 );
nand NAND2_21856 ( P2_R1146_U87 , P2_R1146_U128 , P2_R1146_U301 );
nand NAND2_21857 ( P2_R1146_U88 , P2_R1146_U298 , P2_R1146_U297 );
nand NAND2_21858 ( P2_R1146_U89 , P2_R1146_U76 , P2_R1146_U318 );
nand NAND2_21859 ( P2_R1146_U90 , P2_R1146_U61 , P2_R1146_U329 );
nand NAND2_21860 ( P2_R1146_U91 , P2_R1146_U50 , P2_R1146_U340 );
not NOT1_21861 ( P2_R1146_U92 , P2_U3079 );
nand NAND2_21862 ( P2_R1146_U93 , P2_R1146_U395 , P2_R1146_U394 );
nand NAND2_21863 ( P2_R1146_U94 , P2_R1146_U409 , P2_R1146_U408 );
nand NAND2_21864 ( P2_R1146_U95 , P2_R1146_U414 , P2_R1146_U413 );
nand NAND2_21865 ( P2_R1146_U96 , P2_R1146_U430 , P2_R1146_U429 );
nand NAND2_21866 ( P2_R1146_U97 , P2_R1146_U435 , P2_R1146_U434 );
nand NAND2_21867 ( P2_R1146_U98 , P2_R1146_U440 , P2_R1146_U439 );
nand NAND2_21868 ( P2_R1146_U99 , P2_R1146_U445 , P2_R1146_U444 );
nand NAND2_21869 ( P2_R1146_U100 , P2_R1146_U450 , P2_R1146_U449 );
nand NAND2_21870 ( P2_R1146_U101 , P2_R1146_U466 , P2_R1146_U465 );
nand NAND2_21871 ( P2_R1146_U102 , P2_R1146_U471 , P2_R1146_U470 );
nand NAND2_21872 ( P2_R1146_U103 , P2_R1146_U356 , P2_R1146_U355 );
nand NAND2_21873 ( P2_R1146_U104 , P2_R1146_U365 , P2_R1146_U364 );
nand NAND2_21874 ( P2_R1146_U105 , P2_R1146_U372 , P2_R1146_U371 );
nand NAND2_21875 ( P2_R1146_U106 , P2_R1146_U376 , P2_R1146_U375 );
nand NAND2_21876 ( P2_R1146_U107 , P2_R1146_U385 , P2_R1146_U384 );
nand NAND2_21877 ( P2_R1146_U108 , P2_R1146_U404 , P2_R1146_U403 );
nand NAND2_21878 ( P2_R1146_U109 , P2_R1146_U421 , P2_R1146_U420 );
nand NAND2_21879 ( P2_R1146_U110 , P2_R1146_U425 , P2_R1146_U424 );
nand NAND2_21880 ( P2_R1146_U111 , P2_R1146_U457 , P2_R1146_U456 );
nand NAND2_21881 ( P2_R1146_U112 , P2_R1146_U461 , P2_R1146_U460 );
nand NAND2_21882 ( P2_R1146_U113 , P2_R1146_U478 , P2_R1146_U477 );
and AND2_21883 ( P2_R1146_U114 , P2_R1146_U194 , P2_R1146_U184 );
and AND2_21884 ( P2_R1146_U115 , P2_R1146_U197 , P2_R1146_U198 );
and AND3_21885 ( P2_R1146_U116 , P2_R1146_U205 , P2_R1146_U200 , P2_R1146_U185 );
and AND2_21886 ( P2_R1146_U117 , P2_R1146_U210 , P2_R1146_U186 );
and AND2_21887 ( P2_R1146_U118 , P2_R1146_U213 , P2_R1146_U214 );
and AND3_21888 ( P2_R1146_U119 , P2_R1146_U358 , P2_R1146_U357 , P2_R1146_U38 );
and AND2_21889 ( P2_R1146_U120 , P2_R1146_U361 , P2_R1146_U186 );
and AND2_21890 ( P2_R1146_U121 , P2_R1146_U229 , P2_R1146_U6 );
and AND2_21891 ( P2_R1146_U122 , P2_R1146_U368 , P2_R1146_U185 );
and AND3_21892 ( P2_R1146_U123 , P2_R1146_U378 , P2_R1146_U377 , P2_R1146_U28 );
and AND2_21893 ( P2_R1146_U124 , P2_R1146_U381 , P2_R1146_U184 );
and AND3_21894 ( P2_R1146_U125 , P2_R1146_U239 , P2_R1146_U216 , P2_R1146_U180 );
and AND2_21895 ( P2_R1146_U126 , P2_R1146_U261 , P2_R1146_U8 );
and AND2_21896 ( P2_R1146_U127 , P2_R1146_U287 , P2_R1146_U10 );
and AND2_21897 ( P2_R1146_U128 , P2_R1146_U303 , P2_R1146_U304 );
and AND3_21898 ( P2_R1146_U129 , P2_R1146_U387 , P2_R1146_U386 , P2_R1146_U311 );
and AND2_21899 ( P2_R1146_U130 , P2_R1146_U308 , P2_R1146_U390 );
nand NAND2_21900 ( P2_R1146_U131 , P2_R1146_U392 , P2_R1146_U391 );
and AND3_21901 ( P2_R1146_U132 , P2_R1146_U397 , P2_R1146_U396 , P2_R1146_U83 );
and AND2_21902 ( P2_R1146_U133 , P2_R1146_U400 , P2_R1146_U183 );
nand NAND2_21903 ( P2_R1146_U134 , P2_R1146_U406 , P2_R1146_U405 );
nand NAND2_21904 ( P2_R1146_U135 , P2_R1146_U411 , P2_R1146_U410 );
and AND2_21905 ( P2_R1146_U136 , P2_R1146_U324 , P2_R1146_U11 );
and AND2_21906 ( P2_R1146_U137 , P2_R1146_U417 , P2_R1146_U182 );
nand NAND2_21907 ( P2_R1146_U138 , P2_R1146_U427 , P2_R1146_U426 );
nand NAND2_21908 ( P2_R1146_U139 , P2_R1146_U432 , P2_R1146_U431 );
nand NAND2_21909 ( P2_R1146_U140 , P2_R1146_U437 , P2_R1146_U436 );
nand NAND2_21910 ( P2_R1146_U141 , P2_R1146_U442 , P2_R1146_U441 );
nand NAND2_21911 ( P2_R1146_U142 , P2_R1146_U447 , P2_R1146_U446 );
and AND2_21912 ( P2_R1146_U143 , P2_R1146_U335 , P2_R1146_U9 );
and AND2_21913 ( P2_R1146_U144 , P2_R1146_U453 , P2_R1146_U181 );
nand NAND2_21914 ( P2_R1146_U145 , P2_R1146_U463 , P2_R1146_U462 );
nand NAND2_21915 ( P2_R1146_U146 , P2_R1146_U468 , P2_R1146_U467 );
and AND2_21916 ( P2_R1146_U147 , P2_R1146_U346 , P2_R1146_U7 );
and AND2_21917 ( P2_R1146_U148 , P2_R1146_U474 , P2_R1146_U180 );
and AND2_21918 ( P2_R1146_U149 , P2_R1146_U354 , P2_R1146_U353 );
nand NAND2_21919 ( P2_R1146_U150 , P2_R1146_U118 , P2_R1146_U211 );
and AND2_21920 ( P2_R1146_U151 , P2_R1146_U363 , P2_R1146_U362 );
and AND2_21921 ( P2_R1146_U152 , P2_R1146_U370 , P2_R1146_U369 );
and AND2_21922 ( P2_R1146_U153 , P2_R1146_U374 , P2_R1146_U373 );
nand NAND2_21923 ( P2_R1146_U154 , P2_R1146_U115 , P2_R1146_U195 );
and AND2_21924 ( P2_R1146_U155 , P2_R1146_U383 , P2_R1146_U382 );
not NOT1_21925 ( P2_R1146_U156 , P2_U3960 );
not NOT1_21926 ( P2_R1146_U157 , P2_U3057 );
and AND2_21927 ( P2_R1146_U158 , P2_R1146_U402 , P2_R1146_U401 );
nand NAND2_21928 ( P2_R1146_U159 , P2_R1146_U294 , P2_R1146_U293 );
nand NAND2_21929 ( P2_R1146_U160 , P2_R1146_U290 , P2_R1146_U289 );
and AND2_21930 ( P2_R1146_U161 , P2_R1146_U419 , P2_R1146_U418 );
and AND2_21931 ( P2_R1146_U162 , P2_R1146_U423 , P2_R1146_U422 );
nand NAND2_21932 ( P2_R1146_U163 , P2_R1146_U280 , P2_R1146_U279 );
nand NAND2_21933 ( P2_R1146_U164 , P2_R1146_U276 , P2_R1146_U275 );
not NOT1_21934 ( P2_R1146_U165 , P2_U3432 );
nand NAND2_21935 ( P2_R1146_U166 , P2_U3427 , P2_R1146_U92 );
nand NAND2_21936 ( P2_R1146_U167 , P2_R1146_U272 , P2_R1146_U271 );
not NOT1_21937 ( P2_R1146_U168 , P2_U3483 );
nand NAND2_21938 ( P2_R1146_U169 , P2_R1146_U264 , P2_R1146_U263 );
and AND2_21939 ( P2_R1146_U170 , P2_R1146_U455 , P2_R1146_U454 );
and AND2_21940 ( P2_R1146_U171 , P2_R1146_U459 , P2_R1146_U458 );
nand NAND2_21941 ( P2_R1146_U172 , P2_R1146_U254 , P2_R1146_U253 );
nand NAND2_21942 ( P2_R1146_U173 , P2_R1146_U250 , P2_R1146_U249 );
nand NAND2_21943 ( P2_R1146_U174 , P2_R1146_U246 , P2_R1146_U245 );
and AND2_21944 ( P2_R1146_U175 , P2_R1146_U476 , P2_R1146_U475 );
nand NAND2_21945 ( P2_R1146_U176 , P2_R1146_U166 , P2_R1146_U165 );
not NOT1_21946 ( P2_R1146_U177 , P2_R1146_U83 );
not NOT1_21947 ( P2_R1146_U178 , P2_R1146_U28 );
not NOT1_21948 ( P2_R1146_U179 , P2_R1146_U38 );
nand NAND2_21949 ( P2_R1146_U180 , P2_U3459 , P2_R1146_U49 );
nand NAND2_21950 ( P2_R1146_U181 , P2_U3474 , P2_R1146_U59 );
nand NAND2_21951 ( P2_R1146_U182 , P2_U3955 , P2_R1146_U74 );
nand NAND2_21952 ( P2_R1146_U183 , P2_U3951 , P2_R1146_U82 );
nand NAND2_21953 ( P2_R1146_U184 , P2_U3435 , P2_R1146_U27 );
nand NAND2_21954 ( P2_R1146_U185 , P2_U3444 , P2_R1146_U33 );
nand NAND2_21955 ( P2_R1146_U186 , P2_U3450 , P2_R1146_U37 );
not NOT1_21956 ( P2_R1146_U187 , P2_R1146_U61 );
not NOT1_21957 ( P2_R1146_U188 , P2_R1146_U76 );
not NOT1_21958 ( P2_R1146_U189 , P2_R1146_U35 );
not NOT1_21959 ( P2_R1146_U190 , P2_R1146_U50 );
not NOT1_21960 ( P2_R1146_U191 , P2_R1146_U166 );
nand NAND2_21961 ( P2_R1146_U192 , P2_U3080 , P2_R1146_U166 );
not NOT1_21962 ( P2_R1146_U193 , P2_R1146_U44 );
nand NAND2_21963 ( P2_R1146_U194 , P2_U3438 , P2_R1146_U29 );
nand NAND2_21964 ( P2_R1146_U195 , P2_R1146_U114 , P2_R1146_U44 );
nand NAND2_21965 ( P2_R1146_U196 , P2_R1146_U29 , P2_R1146_U28 );
nand NAND2_21966 ( P2_R1146_U197 , P2_R1146_U196 , P2_R1146_U26 );
nand NAND2_21967 ( P2_R1146_U198 , P2_U3066 , P2_R1146_U178 );
not NOT1_21968 ( P2_R1146_U199 , P2_R1146_U154 );
nand NAND2_21969 ( P2_R1146_U200 , P2_U3447 , P2_R1146_U32 );
nand NAND2_21970 ( P2_R1146_U201 , P2_U3073 , P2_R1146_U30 );
nand NAND2_21971 ( P2_R1146_U202 , P2_U3069 , P2_R1146_U22 );
nand NAND2_21972 ( P2_R1146_U203 , P2_R1146_U189 , P2_R1146_U185 );
nand NAND2_21973 ( P2_R1146_U204 , P2_R1146_U6 , P2_R1146_U203 );
nand NAND2_21974 ( P2_R1146_U205 , P2_U3441 , P2_R1146_U34 );
nand NAND2_21975 ( P2_R1146_U206 , P2_U3447 , P2_R1146_U32 );
nand NAND2_21976 ( P2_R1146_U207 , P2_R1146_U154 , P2_R1146_U116 );
nand NAND2_21977 ( P2_R1146_U208 , P2_R1146_U206 , P2_R1146_U204 );
not NOT1_21978 ( P2_R1146_U209 , P2_R1146_U42 );
nand NAND2_21979 ( P2_R1146_U210 , P2_U3453 , P2_R1146_U39 );
nand NAND2_21980 ( P2_R1146_U211 , P2_R1146_U117 , P2_R1146_U42 );
nand NAND2_21981 ( P2_R1146_U212 , P2_R1146_U39 , P2_R1146_U38 );
nand NAND2_21982 ( P2_R1146_U213 , P2_R1146_U212 , P2_R1146_U36 );
nand NAND2_21983 ( P2_R1146_U214 , P2_U3086 , P2_R1146_U179 );
not NOT1_21984 ( P2_R1146_U215 , P2_R1146_U150 );
nand NAND2_21985 ( P2_R1146_U216 , P2_U3456 , P2_R1146_U41 );
nand NAND2_21986 ( P2_R1146_U217 , P2_R1146_U216 , P2_R1146_U50 );
nand NAND2_21987 ( P2_R1146_U218 , P2_R1146_U209 , P2_R1146_U38 );
nand NAND2_21988 ( P2_R1146_U219 , P2_R1146_U120 , P2_R1146_U218 );
nand NAND2_21989 ( P2_R1146_U220 , P2_R1146_U42 , P2_R1146_U186 );
nand NAND2_21990 ( P2_R1146_U221 , P2_R1146_U119 , P2_R1146_U220 );
nand NAND2_21991 ( P2_R1146_U222 , P2_R1146_U38 , P2_R1146_U186 );
nand NAND2_21992 ( P2_R1146_U223 , P2_R1146_U205 , P2_R1146_U154 );
not NOT1_21993 ( P2_R1146_U224 , P2_R1146_U43 );
nand NAND2_21994 ( P2_R1146_U225 , P2_U3069 , P2_R1146_U22 );
nand NAND2_21995 ( P2_R1146_U226 , P2_R1146_U224 , P2_R1146_U225 );
nand NAND2_21996 ( P2_R1146_U227 , P2_R1146_U122 , P2_R1146_U226 );
nand NAND2_21997 ( P2_R1146_U228 , P2_R1146_U43 , P2_R1146_U185 );
nand NAND2_21998 ( P2_R1146_U229 , P2_U3447 , P2_R1146_U32 );
nand NAND2_21999 ( P2_R1146_U230 , P2_R1146_U121 , P2_R1146_U228 );
nand NAND2_22000 ( P2_R1146_U231 , P2_U3069 , P2_R1146_U22 );
nand NAND2_22001 ( P2_R1146_U232 , P2_R1146_U185 , P2_R1146_U231 );
nand NAND2_22002 ( P2_R1146_U233 , P2_R1146_U205 , P2_R1146_U35 );
nand NAND2_22003 ( P2_R1146_U234 , P2_R1146_U193 , P2_R1146_U28 );
nand NAND2_22004 ( P2_R1146_U235 , P2_R1146_U124 , P2_R1146_U234 );
nand NAND2_22005 ( P2_R1146_U236 , P2_R1146_U44 , P2_R1146_U184 );
nand NAND2_22006 ( P2_R1146_U237 , P2_R1146_U123 , P2_R1146_U236 );
nand NAND2_22007 ( P2_R1146_U238 , P2_R1146_U28 , P2_R1146_U184 );
nand NAND2_22008 ( P2_R1146_U239 , P2_U3462 , P2_R1146_U48 );
nand NAND2_22009 ( P2_R1146_U240 , P2_U3065 , P2_R1146_U47 );
nand NAND2_22010 ( P2_R1146_U241 , P2_U3064 , P2_R1146_U46 );
nand NAND2_22011 ( P2_R1146_U242 , P2_R1146_U190 , P2_R1146_U180 );
nand NAND2_22012 ( P2_R1146_U243 , P2_R1146_U7 , P2_R1146_U242 );
nand NAND2_22013 ( P2_R1146_U244 , P2_U3462 , P2_R1146_U48 );
nand NAND2_22014 ( P2_R1146_U245 , P2_R1146_U150 , P2_R1146_U125 );
nand NAND2_22015 ( P2_R1146_U246 , P2_R1146_U244 , P2_R1146_U243 );
not NOT1_22016 ( P2_R1146_U247 , P2_R1146_U174 );
nand NAND2_22017 ( P2_R1146_U248 , P2_U3465 , P2_R1146_U52 );
nand NAND2_22018 ( P2_R1146_U249 , P2_R1146_U248 , P2_R1146_U174 );
nand NAND2_22019 ( P2_R1146_U250 , P2_U3074 , P2_R1146_U51 );
not NOT1_22020 ( P2_R1146_U251 , P2_R1146_U173 );
nand NAND2_22021 ( P2_R1146_U252 , P2_U3468 , P2_R1146_U54 );
nand NAND2_22022 ( P2_R1146_U253 , P2_R1146_U252 , P2_R1146_U173 );
nand NAND2_22023 ( P2_R1146_U254 , P2_U3082 , P2_R1146_U53 );
not NOT1_22024 ( P2_R1146_U255 , P2_R1146_U172 );
nand NAND2_22025 ( P2_R1146_U256 , P2_U3477 , P2_R1146_U58 );
nand NAND2_22026 ( P2_R1146_U257 , P2_U3075 , P2_R1146_U55 );
nand NAND2_22027 ( P2_R1146_U258 , P2_U3076 , P2_R1146_U56 );
nand NAND2_22028 ( P2_R1146_U259 , P2_R1146_U187 , P2_R1146_U8 );
nand NAND2_22029 ( P2_R1146_U260 , P2_R1146_U9 , P2_R1146_U259 );
nand NAND2_22030 ( P2_R1146_U261 , P2_U3471 , P2_R1146_U60 );
nand NAND2_22031 ( P2_R1146_U262 , P2_U3477 , P2_R1146_U58 );
nand NAND2_22032 ( P2_R1146_U263 , P2_R1146_U126 , P2_R1146_U172 );
nand NAND2_22033 ( P2_R1146_U264 , P2_R1146_U262 , P2_R1146_U260 );
not NOT1_22034 ( P2_R1146_U265 , P2_R1146_U169 );
nand NAND2_22035 ( P2_R1146_U266 , P2_U3480 , P2_R1146_U63 );
nand NAND2_22036 ( P2_R1146_U267 , P2_R1146_U266 , P2_R1146_U169 );
nand NAND2_22037 ( P2_R1146_U268 , P2_U3071 , P2_R1146_U62 );
not NOT1_22038 ( P2_R1146_U269 , P2_R1146_U64 );
nand NAND2_22039 ( P2_R1146_U270 , P2_R1146_U269 , P2_R1146_U65 );
nand NAND2_22040 ( P2_R1146_U271 , P2_R1146_U270 , P2_R1146_U168 );
nand NAND2_22041 ( P2_R1146_U272 , P2_U3084 , P2_R1146_U64 );
not NOT1_22042 ( P2_R1146_U273 , P2_R1146_U167 );
nand NAND2_22043 ( P2_R1146_U274 , P2_U3485 , P2_R1146_U67 );
nand NAND2_22044 ( P2_R1146_U275 , P2_R1146_U274 , P2_R1146_U167 );
nand NAND2_22045 ( P2_R1146_U276 , P2_U3083 , P2_R1146_U66 );
not NOT1_22046 ( P2_R1146_U277 , P2_R1146_U164 );
nand NAND2_22047 ( P2_R1146_U278 , P2_U3957 , P2_R1146_U69 );
nand NAND2_22048 ( P2_R1146_U279 , P2_R1146_U278 , P2_R1146_U164 );
nand NAND2_22049 ( P2_R1146_U280 , P2_U3078 , P2_R1146_U68 );
not NOT1_22050 ( P2_R1146_U281 , P2_R1146_U163 );
nand NAND2_22051 ( P2_R1146_U282 , P2_U3954 , P2_R1146_U73 );
nand NAND2_22052 ( P2_R1146_U283 , P2_U3068 , P2_R1146_U70 );
nand NAND2_22053 ( P2_R1146_U284 , P2_U3063 , P2_R1146_U71 );
nand NAND2_22054 ( P2_R1146_U285 , P2_R1146_U188 , P2_R1146_U10 );
nand NAND2_22055 ( P2_R1146_U286 , P2_R1146_U11 , P2_R1146_U285 );
nand NAND2_22056 ( P2_R1146_U287 , P2_U3956 , P2_R1146_U75 );
nand NAND2_22057 ( P2_R1146_U288 , P2_U3954 , P2_R1146_U73 );
nand NAND2_22058 ( P2_R1146_U289 , P2_R1146_U127 , P2_R1146_U163 );
nand NAND2_22059 ( P2_R1146_U290 , P2_R1146_U288 , P2_R1146_U286 );
not NOT1_22060 ( P2_R1146_U291 , P2_R1146_U160 );
nand NAND2_22061 ( P2_R1146_U292 , P2_U3953 , P2_R1146_U78 );
nand NAND2_22062 ( P2_R1146_U293 , P2_R1146_U292 , P2_R1146_U160 );
nand NAND2_22063 ( P2_R1146_U294 , P2_U3067 , P2_R1146_U77 );
not NOT1_22064 ( P2_R1146_U295 , P2_R1146_U159 );
nand NAND2_22065 ( P2_R1146_U296 , P2_U3952 , P2_R1146_U80 );
nand NAND2_22066 ( P2_R1146_U297 , P2_R1146_U296 , P2_R1146_U159 );
nand NAND2_22067 ( P2_R1146_U298 , P2_U3060 , P2_R1146_U79 );
not NOT1_22068 ( P2_R1146_U299 , P2_R1146_U88 );
nand NAND2_22069 ( P2_R1146_U300 , P2_U3950 , P2_R1146_U84 );
nand NAND3_22070 ( P2_R1146_U301 , P2_R1146_U88 , P2_R1146_U183 , P2_R1146_U300 );
nand NAND2_22071 ( P2_R1146_U302 , P2_R1146_U84 , P2_R1146_U83 );
nand NAND2_22072 ( P2_R1146_U303 , P2_R1146_U302 , P2_R1146_U81 );
nand NAND2_22073 ( P2_R1146_U304 , P2_U3055 , P2_R1146_U177 );
not NOT1_22074 ( P2_R1146_U305 , P2_R1146_U87 );
nand NAND2_22075 ( P2_R1146_U306 , P2_U3056 , P2_R1146_U85 );
nand NAND2_22076 ( P2_R1146_U307 , P2_R1146_U305 , P2_R1146_U306 );
nand NAND2_22077 ( P2_R1146_U308 , P2_U3949 , P2_R1146_U86 );
nand NAND2_22078 ( P2_R1146_U309 , P2_U3949 , P2_R1146_U86 );
nand NAND2_22079 ( P2_R1146_U310 , P2_R1146_U309 , P2_R1146_U87 );
nand NAND2_22080 ( P2_R1146_U311 , P2_U3056 , P2_R1146_U85 );
nand NAND2_22081 ( P2_R1146_U312 , P2_R1146_U129 , P2_R1146_U310 );
nand NAND2_22082 ( P2_R1146_U313 , P2_R1146_U299 , P2_R1146_U83 );
nand NAND2_22083 ( P2_R1146_U314 , P2_R1146_U133 , P2_R1146_U313 );
nand NAND2_22084 ( P2_R1146_U315 , P2_R1146_U88 , P2_R1146_U183 );
nand NAND2_22085 ( P2_R1146_U316 , P2_R1146_U132 , P2_R1146_U315 );
nand NAND2_22086 ( P2_R1146_U317 , P2_R1146_U83 , P2_R1146_U183 );
nand NAND2_22087 ( P2_R1146_U318 , P2_R1146_U287 , P2_R1146_U163 );
not NOT1_22088 ( P2_R1146_U319 , P2_R1146_U89 );
nand NAND2_22089 ( P2_R1146_U320 , P2_U3063 , P2_R1146_U71 );
nand NAND2_22090 ( P2_R1146_U321 , P2_R1146_U319 , P2_R1146_U320 );
nand NAND2_22091 ( P2_R1146_U322 , P2_R1146_U137 , P2_R1146_U321 );
nand NAND2_22092 ( P2_R1146_U323 , P2_R1146_U89 , P2_R1146_U182 );
nand NAND2_22093 ( P2_R1146_U324 , P2_U3954 , P2_R1146_U73 );
nand NAND2_22094 ( P2_R1146_U325 , P2_R1146_U136 , P2_R1146_U323 );
nand NAND2_22095 ( P2_R1146_U326 , P2_U3063 , P2_R1146_U71 );
nand NAND2_22096 ( P2_R1146_U327 , P2_R1146_U182 , P2_R1146_U326 );
nand NAND2_22097 ( P2_R1146_U328 , P2_R1146_U287 , P2_R1146_U76 );
nand NAND2_22098 ( P2_R1146_U329 , P2_R1146_U261 , P2_R1146_U172 );
not NOT1_22099 ( P2_R1146_U330 , P2_R1146_U90 );
nand NAND2_22100 ( P2_R1146_U331 , P2_U3076 , P2_R1146_U56 );
nand NAND2_22101 ( P2_R1146_U332 , P2_R1146_U330 , P2_R1146_U331 );
nand NAND2_22102 ( P2_R1146_U333 , P2_R1146_U144 , P2_R1146_U332 );
nand NAND2_22103 ( P2_R1146_U334 , P2_R1146_U90 , P2_R1146_U181 );
nand NAND2_22104 ( P2_R1146_U335 , P2_U3477 , P2_R1146_U58 );
nand NAND2_22105 ( P2_R1146_U336 , P2_R1146_U143 , P2_R1146_U334 );
nand NAND2_22106 ( P2_R1146_U337 , P2_U3076 , P2_R1146_U56 );
nand NAND2_22107 ( P2_R1146_U338 , P2_R1146_U181 , P2_R1146_U337 );
nand NAND2_22108 ( P2_R1146_U339 , P2_R1146_U261 , P2_R1146_U61 );
nand NAND2_22109 ( P2_R1146_U340 , P2_R1146_U216 , P2_R1146_U150 );
not NOT1_22110 ( P2_R1146_U341 , P2_R1146_U91 );
nand NAND2_22111 ( P2_R1146_U342 , P2_U3064 , P2_R1146_U46 );
nand NAND2_22112 ( P2_R1146_U343 , P2_R1146_U341 , P2_R1146_U342 );
nand NAND2_22113 ( P2_R1146_U344 , P2_R1146_U148 , P2_R1146_U343 );
nand NAND2_22114 ( P2_R1146_U345 , P2_R1146_U91 , P2_R1146_U180 );
nand NAND2_22115 ( P2_R1146_U346 , P2_U3462 , P2_R1146_U48 );
nand NAND2_22116 ( P2_R1146_U347 , P2_R1146_U147 , P2_R1146_U345 );
nand NAND2_22117 ( P2_R1146_U348 , P2_U3064 , P2_R1146_U46 );
nand NAND2_22118 ( P2_R1146_U349 , P2_R1146_U180 , P2_R1146_U348 );
nand NAND2_22119 ( P2_R1146_U350 , P2_U3079 , P2_R1146_U24 );
nand NAND2_22120 ( P2_R1146_U351 , P2_U3080 , P2_R1146_U165 );
nand NAND2_22121 ( P2_R1146_U352 , P2_R1146_U130 , P2_R1146_U307 );
nand NAND2_22122 ( P2_R1146_U353 , P2_U3456 , P2_R1146_U41 );
nand NAND2_22123 ( P2_R1146_U354 , P2_U3085 , P2_R1146_U40 );
nand NAND2_22124 ( P2_R1146_U355 , P2_R1146_U217 , P2_R1146_U150 );
nand NAND2_22125 ( P2_R1146_U356 , P2_R1146_U215 , P2_R1146_U149 );
nand NAND2_22126 ( P2_R1146_U357 , P2_U3453 , P2_R1146_U39 );
nand NAND2_22127 ( P2_R1146_U358 , P2_U3086 , P2_R1146_U36 );
nand NAND2_22128 ( P2_R1146_U359 , P2_U3453 , P2_R1146_U39 );
nand NAND2_22129 ( P2_R1146_U360 , P2_U3086 , P2_R1146_U36 );
nand NAND2_22130 ( P2_R1146_U361 , P2_R1146_U360 , P2_R1146_U359 );
nand NAND2_22131 ( P2_R1146_U362 , P2_U3450 , P2_R1146_U37 );
nand NAND2_22132 ( P2_R1146_U363 , P2_U3072 , P2_R1146_U21 );
nand NAND2_22133 ( P2_R1146_U364 , P2_R1146_U222 , P2_R1146_U42 );
nand NAND2_22134 ( P2_R1146_U365 , P2_R1146_U151 , P2_R1146_U209 );
nand NAND2_22135 ( P2_R1146_U366 , P2_U3447 , P2_R1146_U32 );
nand NAND2_22136 ( P2_R1146_U367 , P2_U3073 , P2_R1146_U30 );
nand NAND2_22137 ( P2_R1146_U368 , P2_R1146_U367 , P2_R1146_U366 );
nand NAND2_22138 ( P2_R1146_U369 , P2_U3444 , P2_R1146_U33 );
nand NAND2_22139 ( P2_R1146_U370 , P2_U3069 , P2_R1146_U22 );
nand NAND2_22140 ( P2_R1146_U371 , P2_R1146_U232 , P2_R1146_U43 );
nand NAND2_22141 ( P2_R1146_U372 , P2_R1146_U152 , P2_R1146_U224 );
nand NAND2_22142 ( P2_R1146_U373 , P2_U3441 , P2_R1146_U34 );
nand NAND2_22143 ( P2_R1146_U374 , P2_U3062 , P2_R1146_U31 );
nand NAND2_22144 ( P2_R1146_U375 , P2_R1146_U233 , P2_R1146_U154 );
nand NAND2_22145 ( P2_R1146_U376 , P2_R1146_U199 , P2_R1146_U153 );
nand NAND2_22146 ( P2_R1146_U377 , P2_U3438 , P2_R1146_U29 );
nand NAND2_22147 ( P2_R1146_U378 , P2_U3066 , P2_R1146_U26 );
nand NAND2_22148 ( P2_R1146_U379 , P2_U3438 , P2_R1146_U29 );
nand NAND2_22149 ( P2_R1146_U380 , P2_U3066 , P2_R1146_U26 );
nand NAND2_22150 ( P2_R1146_U381 , P2_R1146_U380 , P2_R1146_U379 );
nand NAND2_22151 ( P2_R1146_U382 , P2_U3435 , P2_R1146_U27 );
nand NAND2_22152 ( P2_R1146_U383 , P2_U3070 , P2_R1146_U23 );
nand NAND2_22153 ( P2_R1146_U384 , P2_R1146_U238 , P2_R1146_U44 );
nand NAND2_22154 ( P2_R1146_U385 , P2_R1146_U155 , P2_R1146_U193 );
nand NAND2_22155 ( P2_R1146_U386 , P2_U3960 , P2_R1146_U157 );
nand NAND2_22156 ( P2_R1146_U387 , P2_U3057 , P2_R1146_U156 );
nand NAND2_22157 ( P2_R1146_U388 , P2_U3960 , P2_R1146_U157 );
nand NAND2_22158 ( P2_R1146_U389 , P2_U3057 , P2_R1146_U156 );
nand NAND2_22159 ( P2_R1146_U390 , P2_R1146_U389 , P2_R1146_U388 );
nand NAND2_22160 ( P2_R1146_U391 , P2_U3949 , P2_R1146_U86 );
nand NAND2_22161 ( P2_R1146_U392 , P2_U3056 , P2_R1146_U85 );
not NOT1_22162 ( P2_R1146_U393 , P2_R1146_U131 );
nand NAND2_22163 ( P2_R1146_U394 , P2_R1146_U393 , P2_R1146_U305 );
nand NAND2_22164 ( P2_R1146_U395 , P2_R1146_U131 , P2_R1146_U87 );
nand NAND2_22165 ( P2_R1146_U396 , P2_U3950 , P2_R1146_U84 );
nand NAND2_22166 ( P2_R1146_U397 , P2_U3055 , P2_R1146_U81 );
nand NAND2_22167 ( P2_R1146_U398 , P2_U3950 , P2_R1146_U84 );
nand NAND2_22168 ( P2_R1146_U399 , P2_U3055 , P2_R1146_U81 );
nand NAND2_22169 ( P2_R1146_U400 , P2_R1146_U399 , P2_R1146_U398 );
nand NAND2_22170 ( P2_R1146_U401 , P2_U3951 , P2_R1146_U82 );
nand NAND2_22171 ( P2_R1146_U402 , P2_U3059 , P2_R1146_U45 );
nand NAND2_22172 ( P2_R1146_U403 , P2_R1146_U317 , P2_R1146_U88 );
nand NAND2_22173 ( P2_R1146_U404 , P2_R1146_U158 , P2_R1146_U299 );
nand NAND2_22174 ( P2_R1146_U405 , P2_U3952 , P2_R1146_U80 );
nand NAND2_22175 ( P2_R1146_U406 , P2_U3060 , P2_R1146_U79 );
not NOT1_22176 ( P2_R1146_U407 , P2_R1146_U134 );
nand NAND2_22177 ( P2_R1146_U408 , P2_R1146_U295 , P2_R1146_U407 );
nand NAND2_22178 ( P2_R1146_U409 , P2_R1146_U134 , P2_R1146_U159 );
nand NAND2_22179 ( P2_R1146_U410 , P2_U3953 , P2_R1146_U78 );
nand NAND2_22180 ( P2_R1146_U411 , P2_U3067 , P2_R1146_U77 );
not NOT1_22181 ( P2_R1146_U412 , P2_R1146_U135 );
nand NAND2_22182 ( P2_R1146_U413 , P2_R1146_U291 , P2_R1146_U412 );
nand NAND2_22183 ( P2_R1146_U414 , P2_R1146_U135 , P2_R1146_U160 );
nand NAND2_22184 ( P2_R1146_U415 , P2_U3954 , P2_R1146_U73 );
nand NAND2_22185 ( P2_R1146_U416 , P2_U3068 , P2_R1146_U70 );
nand NAND2_22186 ( P2_R1146_U417 , P2_R1146_U416 , P2_R1146_U415 );
nand NAND2_22187 ( P2_R1146_U418 , P2_U3955 , P2_R1146_U74 );
nand NAND2_22188 ( P2_R1146_U419 , P2_U3063 , P2_R1146_U71 );
nand NAND2_22189 ( P2_R1146_U420 , P2_R1146_U327 , P2_R1146_U89 );
nand NAND2_22190 ( P2_R1146_U421 , P2_R1146_U161 , P2_R1146_U319 );
nand NAND2_22191 ( P2_R1146_U422 , P2_U3956 , P2_R1146_U75 );
nand NAND2_22192 ( P2_R1146_U423 , P2_U3077 , P2_R1146_U72 );
nand NAND2_22193 ( P2_R1146_U424 , P2_R1146_U328 , P2_R1146_U163 );
nand NAND2_22194 ( P2_R1146_U425 , P2_R1146_U281 , P2_R1146_U162 );
nand NAND2_22195 ( P2_R1146_U426 , P2_U3957 , P2_R1146_U69 );
nand NAND2_22196 ( P2_R1146_U427 , P2_U3078 , P2_R1146_U68 );
not NOT1_22197 ( P2_R1146_U428 , P2_R1146_U138 );
nand NAND2_22198 ( P2_R1146_U429 , P2_R1146_U277 , P2_R1146_U428 );
nand NAND2_22199 ( P2_R1146_U430 , P2_R1146_U138 , P2_R1146_U164 );
nand NAND2_22200 ( P2_R1146_U431 , P2_U3432 , P2_R1146_U25 );
nand NAND2_22201 ( P2_R1146_U432 , P2_U3080 , P2_R1146_U165 );
not NOT1_22202 ( P2_R1146_U433 , P2_R1146_U139 );
nand NAND2_22203 ( P2_R1146_U434 , P2_R1146_U191 , P2_R1146_U433 );
nand NAND2_22204 ( P2_R1146_U435 , P2_R1146_U139 , P2_R1146_U166 );
nand NAND2_22205 ( P2_R1146_U436 , P2_U3485 , P2_R1146_U67 );
nand NAND2_22206 ( P2_R1146_U437 , P2_U3083 , P2_R1146_U66 );
not NOT1_22207 ( P2_R1146_U438 , P2_R1146_U140 );
nand NAND2_22208 ( P2_R1146_U439 , P2_R1146_U273 , P2_R1146_U438 );
nand NAND2_22209 ( P2_R1146_U440 , P2_R1146_U140 , P2_R1146_U167 );
nand NAND2_22210 ( P2_R1146_U441 , P2_U3483 , P2_R1146_U65 );
nand NAND2_22211 ( P2_R1146_U442 , P2_U3084 , P2_R1146_U168 );
not NOT1_22212 ( P2_R1146_U443 , P2_R1146_U141 );
nand NAND2_22213 ( P2_R1146_U444 , P2_R1146_U443 , P2_R1146_U269 );
nand NAND2_22214 ( P2_R1146_U445 , P2_R1146_U141 , P2_R1146_U64 );
nand NAND2_22215 ( P2_R1146_U446 , P2_U3480 , P2_R1146_U63 );
nand NAND2_22216 ( P2_R1146_U447 , P2_U3071 , P2_R1146_U62 );
not NOT1_22217 ( P2_R1146_U448 , P2_R1146_U142 );
nand NAND2_22218 ( P2_R1146_U449 , P2_R1146_U265 , P2_R1146_U448 );
nand NAND2_22219 ( P2_R1146_U450 , P2_R1146_U142 , P2_R1146_U169 );
nand NAND2_22220 ( P2_R1146_U451 , P2_U3477 , P2_R1146_U58 );
nand NAND2_22221 ( P2_R1146_U452 , P2_U3075 , P2_R1146_U55 );
nand NAND2_22222 ( P2_R1146_U453 , P2_R1146_U452 , P2_R1146_U451 );
nand NAND2_22223 ( P2_R1146_U454 , P2_U3474 , P2_R1146_U59 );
nand NAND2_22224 ( P2_R1146_U455 , P2_U3076 , P2_R1146_U56 );
nand NAND2_22225 ( P2_R1146_U456 , P2_R1146_U338 , P2_R1146_U90 );
nand NAND2_22226 ( P2_R1146_U457 , P2_R1146_U170 , P2_R1146_U330 );
nand NAND2_22227 ( P2_R1146_U458 , P2_U3471 , P2_R1146_U60 );
nand NAND2_22228 ( P2_R1146_U459 , P2_U3081 , P2_R1146_U57 );
nand NAND2_22229 ( P2_R1146_U460 , P2_R1146_U339 , P2_R1146_U172 );
nand NAND2_22230 ( P2_R1146_U461 , P2_R1146_U255 , P2_R1146_U171 );
nand NAND2_22231 ( P2_R1146_U462 , P2_U3468 , P2_R1146_U54 );
nand NAND2_22232 ( P2_R1146_U463 , P2_U3082 , P2_R1146_U53 );
not NOT1_22233 ( P2_R1146_U464 , P2_R1146_U145 );
nand NAND2_22234 ( P2_R1146_U465 , P2_R1146_U251 , P2_R1146_U464 );
nand NAND2_22235 ( P2_R1146_U466 , P2_R1146_U145 , P2_R1146_U173 );
nand NAND2_22236 ( P2_R1146_U467 , P2_U3465 , P2_R1146_U52 );
nand NAND2_22237 ( P2_R1146_U468 , P2_U3074 , P2_R1146_U51 );
not NOT1_22238 ( P2_R1146_U469 , P2_R1146_U146 );
nand NAND2_22239 ( P2_R1146_U470 , P2_R1146_U247 , P2_R1146_U469 );
nand NAND2_22240 ( P2_R1146_U471 , P2_R1146_U146 , P2_R1146_U174 );
nand NAND2_22241 ( P2_R1146_U472 , P2_U3462 , P2_R1146_U48 );
nand NAND2_22242 ( P2_R1146_U473 , P2_U3065 , P2_R1146_U47 );
nand NAND2_22243 ( P2_R1146_U474 , P2_R1146_U473 , P2_R1146_U472 );
nand NAND2_22244 ( P2_R1146_U475 , P2_U3459 , P2_R1146_U49 );
nand NAND2_22245 ( P2_R1146_U476 , P2_U3064 , P2_R1146_U46 );
nand NAND2_22246 ( P2_R1146_U477 , P2_R1146_U349 , P2_R1146_U91 );
nand NAND2_22247 ( P2_R1146_U478 , P2_R1146_U175 , P2_R1146_U341 );
and AND2_22248 ( P2_R1203_U6 , P2_R1203_U202 , P2_R1203_U201 );
and AND2_22249 ( P2_R1203_U7 , P2_R1203_U241 , P2_R1203_U240 );
and AND2_22250 ( P2_R1203_U8 , P2_R1203_U181 , P2_R1203_U256 );
and AND2_22251 ( P2_R1203_U9 , P2_R1203_U258 , P2_R1203_U257 );
and AND2_22252 ( P2_R1203_U10 , P2_R1203_U182 , P2_R1203_U282 );
and AND2_22253 ( P2_R1203_U11 , P2_R1203_U284 , P2_R1203_U283 );
nand NAND2_22254 ( P2_R1203_U12 , P2_R1203_U344 , P2_R1203_U347 );
nand NAND2_22255 ( P2_R1203_U13 , P2_R1203_U333 , P2_R1203_U336 );
nand NAND2_22256 ( P2_R1203_U14 , P2_R1203_U322 , P2_R1203_U325 );
nand NAND2_22257 ( P2_R1203_U15 , P2_R1203_U314 , P2_R1203_U316 );
nand NAND2_22258 ( P2_R1203_U16 , P2_R1203_U352 , P2_R1203_U312 );
nand NAND2_22259 ( P2_R1203_U17 , P2_R1203_U235 , P2_R1203_U237 );
nand NAND2_22260 ( P2_R1203_U18 , P2_R1203_U227 , P2_R1203_U230 );
nand NAND2_22261 ( P2_R1203_U19 , P2_R1203_U219 , P2_R1203_U221 );
nand NAND2_22262 ( P2_R1203_U20 , P2_R1203_U166 , P2_R1203_U350 );
not NOT1_22263 ( P2_R1203_U21 , P2_U3450 );
not NOT1_22264 ( P2_R1203_U22 , P2_U3444 );
not NOT1_22265 ( P2_R1203_U23 , P2_U3435 );
not NOT1_22266 ( P2_R1203_U24 , P2_U3427 );
not NOT1_22267 ( P2_R1203_U25 , P2_U3080 );
not NOT1_22268 ( P2_R1203_U26 , P2_U3438 );
not NOT1_22269 ( P2_R1203_U27 , P2_U3070 );
nand NAND2_22270 ( P2_R1203_U28 , P2_U3070 , P2_R1203_U23 );
not NOT1_22271 ( P2_R1203_U29 , P2_U3066 );
not NOT1_22272 ( P2_R1203_U30 , P2_U3447 );
not NOT1_22273 ( P2_R1203_U31 , P2_U3441 );
not NOT1_22274 ( P2_R1203_U32 , P2_U3073 );
not NOT1_22275 ( P2_R1203_U33 , P2_U3069 );
not NOT1_22276 ( P2_R1203_U34 , P2_U3062 );
nand NAND2_22277 ( P2_R1203_U35 , P2_U3062 , P2_R1203_U31 );
not NOT1_22278 ( P2_R1203_U36 , P2_U3453 );
not NOT1_22279 ( P2_R1203_U37 , P2_U3072 );
nand NAND2_22280 ( P2_R1203_U38 , P2_U3072 , P2_R1203_U21 );
not NOT1_22281 ( P2_R1203_U39 , P2_U3086 );
not NOT1_22282 ( P2_R1203_U40 , P2_U3456 );
not NOT1_22283 ( P2_R1203_U41 , P2_U3085 );
nand NAND2_22284 ( P2_R1203_U42 , P2_R1203_U208 , P2_R1203_U207 );
nand NAND2_22285 ( P2_R1203_U43 , P2_R1203_U35 , P2_R1203_U223 );
nand NAND3_22286 ( P2_R1203_U44 , P2_R1203_U192 , P2_R1203_U176 , P2_R1203_U351 );
not NOT1_22287 ( P2_R1203_U45 , P2_U3951 );
not NOT1_22288 ( P2_R1203_U46 , P2_U3459 );
not NOT1_22289 ( P2_R1203_U47 , P2_U3462 );
not NOT1_22290 ( P2_R1203_U48 , P2_U3065 );
not NOT1_22291 ( P2_R1203_U49 , P2_U3064 );
nand NAND2_22292 ( P2_R1203_U50 , P2_U3085 , P2_R1203_U40 );
not NOT1_22293 ( P2_R1203_U51 , P2_U3465 );
not NOT1_22294 ( P2_R1203_U52 , P2_U3074 );
not NOT1_22295 ( P2_R1203_U53 , P2_U3468 );
not NOT1_22296 ( P2_R1203_U54 , P2_U3082 );
not NOT1_22297 ( P2_R1203_U55 , P2_U3477 );
not NOT1_22298 ( P2_R1203_U56 , P2_U3474 );
not NOT1_22299 ( P2_R1203_U57 , P2_U3471 );
not NOT1_22300 ( P2_R1203_U58 , P2_U3075 );
not NOT1_22301 ( P2_R1203_U59 , P2_U3076 );
not NOT1_22302 ( P2_R1203_U60 , P2_U3081 );
nand NAND2_22303 ( P2_R1203_U61 , P2_U3081 , P2_R1203_U57 );
not NOT1_22304 ( P2_R1203_U62 , P2_U3480 );
not NOT1_22305 ( P2_R1203_U63 , P2_U3071 );
nand NAND2_22306 ( P2_R1203_U64 , P2_R1203_U268 , P2_R1203_U267 );
not NOT1_22307 ( P2_R1203_U65 , P2_U3084 );
not NOT1_22308 ( P2_R1203_U66 , P2_U3485 );
not NOT1_22309 ( P2_R1203_U67 , P2_U3083 );
not NOT1_22310 ( P2_R1203_U68 , P2_U3957 );
not NOT1_22311 ( P2_R1203_U69 , P2_U3078 );
not NOT1_22312 ( P2_R1203_U70 , P2_U3954 );
not NOT1_22313 ( P2_R1203_U71 , P2_U3955 );
not NOT1_22314 ( P2_R1203_U72 , P2_U3956 );
not NOT1_22315 ( P2_R1203_U73 , P2_U3068 );
not NOT1_22316 ( P2_R1203_U74 , P2_U3063 );
not NOT1_22317 ( P2_R1203_U75 , P2_U3077 );
nand NAND2_22318 ( P2_R1203_U76 , P2_U3077 , P2_R1203_U72 );
not NOT1_22319 ( P2_R1203_U77 , P2_U3953 );
not NOT1_22320 ( P2_R1203_U78 , P2_U3067 );
not NOT1_22321 ( P2_R1203_U79 , P2_U3952 );
not NOT1_22322 ( P2_R1203_U80 , P2_U3060 );
not NOT1_22323 ( P2_R1203_U81 , P2_U3950 );
not NOT1_22324 ( P2_R1203_U82 , P2_U3059 );
nand NAND2_22325 ( P2_R1203_U83 , P2_U3059 , P2_R1203_U45 );
not NOT1_22326 ( P2_R1203_U84 , P2_U3055 );
not NOT1_22327 ( P2_R1203_U85 , P2_U3949 );
not NOT1_22328 ( P2_R1203_U86 , P2_U3056 );
nand NAND2_22329 ( P2_R1203_U87 , P2_R1203_U128 , P2_R1203_U301 );
nand NAND2_22330 ( P2_R1203_U88 , P2_R1203_U298 , P2_R1203_U297 );
nand NAND2_22331 ( P2_R1203_U89 , P2_R1203_U76 , P2_R1203_U318 );
nand NAND2_22332 ( P2_R1203_U90 , P2_R1203_U61 , P2_R1203_U329 );
nand NAND2_22333 ( P2_R1203_U91 , P2_R1203_U50 , P2_R1203_U340 );
not NOT1_22334 ( P2_R1203_U92 , P2_U3079 );
nand NAND2_22335 ( P2_R1203_U93 , P2_R1203_U395 , P2_R1203_U394 );
nand NAND2_22336 ( P2_R1203_U94 , P2_R1203_U409 , P2_R1203_U408 );
nand NAND2_22337 ( P2_R1203_U95 , P2_R1203_U414 , P2_R1203_U413 );
nand NAND2_22338 ( P2_R1203_U96 , P2_R1203_U430 , P2_R1203_U429 );
nand NAND2_22339 ( P2_R1203_U97 , P2_R1203_U435 , P2_R1203_U434 );
nand NAND2_22340 ( P2_R1203_U98 , P2_R1203_U440 , P2_R1203_U439 );
nand NAND2_22341 ( P2_R1203_U99 , P2_R1203_U445 , P2_R1203_U444 );
nand NAND2_22342 ( P2_R1203_U100 , P2_R1203_U450 , P2_R1203_U449 );
nand NAND2_22343 ( P2_R1203_U101 , P2_R1203_U466 , P2_R1203_U465 );
nand NAND2_22344 ( P2_R1203_U102 , P2_R1203_U471 , P2_R1203_U470 );
nand NAND2_22345 ( P2_R1203_U103 , P2_R1203_U356 , P2_R1203_U355 );
nand NAND2_22346 ( P2_R1203_U104 , P2_R1203_U365 , P2_R1203_U364 );
nand NAND2_22347 ( P2_R1203_U105 , P2_R1203_U372 , P2_R1203_U371 );
nand NAND2_22348 ( P2_R1203_U106 , P2_R1203_U376 , P2_R1203_U375 );
nand NAND2_22349 ( P2_R1203_U107 , P2_R1203_U385 , P2_R1203_U384 );
nand NAND2_22350 ( P2_R1203_U108 , P2_R1203_U404 , P2_R1203_U403 );
nand NAND2_22351 ( P2_R1203_U109 , P2_R1203_U421 , P2_R1203_U420 );
nand NAND2_22352 ( P2_R1203_U110 , P2_R1203_U425 , P2_R1203_U424 );
nand NAND2_22353 ( P2_R1203_U111 , P2_R1203_U457 , P2_R1203_U456 );
nand NAND2_22354 ( P2_R1203_U112 , P2_R1203_U461 , P2_R1203_U460 );
nand NAND2_22355 ( P2_R1203_U113 , P2_R1203_U478 , P2_R1203_U477 );
and AND2_22356 ( P2_R1203_U114 , P2_R1203_U194 , P2_R1203_U184 );
and AND2_22357 ( P2_R1203_U115 , P2_R1203_U197 , P2_R1203_U198 );
and AND3_22358 ( P2_R1203_U116 , P2_R1203_U205 , P2_R1203_U200 , P2_R1203_U185 );
and AND2_22359 ( P2_R1203_U117 , P2_R1203_U210 , P2_R1203_U186 );
and AND2_22360 ( P2_R1203_U118 , P2_R1203_U213 , P2_R1203_U214 );
and AND3_22361 ( P2_R1203_U119 , P2_R1203_U358 , P2_R1203_U357 , P2_R1203_U38 );
and AND2_22362 ( P2_R1203_U120 , P2_R1203_U361 , P2_R1203_U186 );
and AND2_22363 ( P2_R1203_U121 , P2_R1203_U229 , P2_R1203_U6 );
and AND2_22364 ( P2_R1203_U122 , P2_R1203_U368 , P2_R1203_U185 );
and AND3_22365 ( P2_R1203_U123 , P2_R1203_U378 , P2_R1203_U377 , P2_R1203_U28 );
and AND2_22366 ( P2_R1203_U124 , P2_R1203_U381 , P2_R1203_U184 );
and AND3_22367 ( P2_R1203_U125 , P2_R1203_U239 , P2_R1203_U216 , P2_R1203_U180 );
and AND2_22368 ( P2_R1203_U126 , P2_R1203_U261 , P2_R1203_U8 );
and AND2_22369 ( P2_R1203_U127 , P2_R1203_U287 , P2_R1203_U10 );
and AND2_22370 ( P2_R1203_U128 , P2_R1203_U303 , P2_R1203_U304 );
and AND3_22371 ( P2_R1203_U129 , P2_R1203_U387 , P2_R1203_U386 , P2_R1203_U311 );
and AND2_22372 ( P2_R1203_U130 , P2_R1203_U308 , P2_R1203_U390 );
nand NAND2_22373 ( P2_R1203_U131 , P2_R1203_U392 , P2_R1203_U391 );
and AND3_22374 ( P2_R1203_U132 , P2_R1203_U397 , P2_R1203_U396 , P2_R1203_U83 );
and AND2_22375 ( P2_R1203_U133 , P2_R1203_U400 , P2_R1203_U183 );
nand NAND2_22376 ( P2_R1203_U134 , P2_R1203_U406 , P2_R1203_U405 );
nand NAND2_22377 ( P2_R1203_U135 , P2_R1203_U411 , P2_R1203_U410 );
and AND2_22378 ( P2_R1203_U136 , P2_R1203_U324 , P2_R1203_U11 );
and AND2_22379 ( P2_R1203_U137 , P2_R1203_U417 , P2_R1203_U182 );
nand NAND2_22380 ( P2_R1203_U138 , P2_R1203_U427 , P2_R1203_U426 );
nand NAND2_22381 ( P2_R1203_U139 , P2_R1203_U432 , P2_R1203_U431 );
nand NAND2_22382 ( P2_R1203_U140 , P2_R1203_U437 , P2_R1203_U436 );
nand NAND2_22383 ( P2_R1203_U141 , P2_R1203_U442 , P2_R1203_U441 );
nand NAND2_22384 ( P2_R1203_U142 , P2_R1203_U447 , P2_R1203_U446 );
and AND2_22385 ( P2_R1203_U143 , P2_R1203_U335 , P2_R1203_U9 );
and AND2_22386 ( P2_R1203_U144 , P2_R1203_U453 , P2_R1203_U181 );
nand NAND2_22387 ( P2_R1203_U145 , P2_R1203_U463 , P2_R1203_U462 );
nand NAND2_22388 ( P2_R1203_U146 , P2_R1203_U468 , P2_R1203_U467 );
and AND2_22389 ( P2_R1203_U147 , P2_R1203_U346 , P2_R1203_U7 );
and AND2_22390 ( P2_R1203_U148 , P2_R1203_U474 , P2_R1203_U180 );
and AND2_22391 ( P2_R1203_U149 , P2_R1203_U354 , P2_R1203_U353 );
nand NAND2_22392 ( P2_R1203_U150 , P2_R1203_U118 , P2_R1203_U211 );
and AND2_22393 ( P2_R1203_U151 , P2_R1203_U363 , P2_R1203_U362 );
and AND2_22394 ( P2_R1203_U152 , P2_R1203_U370 , P2_R1203_U369 );
and AND2_22395 ( P2_R1203_U153 , P2_R1203_U374 , P2_R1203_U373 );
nand NAND2_22396 ( P2_R1203_U154 , P2_R1203_U115 , P2_R1203_U195 );
and AND2_22397 ( P2_R1203_U155 , P2_R1203_U383 , P2_R1203_U382 );
not NOT1_22398 ( P2_R1203_U156 , P2_U3960 );
not NOT1_22399 ( P2_R1203_U157 , P2_U3057 );
and AND2_22400 ( P2_R1203_U158 , P2_R1203_U402 , P2_R1203_U401 );
nand NAND2_22401 ( P2_R1203_U159 , P2_R1203_U294 , P2_R1203_U293 );
nand NAND2_22402 ( P2_R1203_U160 , P2_R1203_U290 , P2_R1203_U289 );
and AND2_22403 ( P2_R1203_U161 , P2_R1203_U419 , P2_R1203_U418 );
and AND2_22404 ( P2_R1203_U162 , P2_R1203_U423 , P2_R1203_U422 );
nand NAND2_22405 ( P2_R1203_U163 , P2_R1203_U280 , P2_R1203_U279 );
nand NAND2_22406 ( P2_R1203_U164 , P2_R1203_U276 , P2_R1203_U275 );
not NOT1_22407 ( P2_R1203_U165 , P2_U3432 );
nand NAND2_22408 ( P2_R1203_U166 , P2_U3427 , P2_R1203_U92 );
nand NAND2_22409 ( P2_R1203_U167 , P2_R1203_U272 , P2_R1203_U271 );
not NOT1_22410 ( P2_R1203_U168 , P2_U3483 );
nand NAND2_22411 ( P2_R1203_U169 , P2_R1203_U264 , P2_R1203_U263 );
and AND2_22412 ( P2_R1203_U170 , P2_R1203_U455 , P2_R1203_U454 );
and AND2_22413 ( P2_R1203_U171 , P2_R1203_U459 , P2_R1203_U458 );
nand NAND2_22414 ( P2_R1203_U172 , P2_R1203_U254 , P2_R1203_U253 );
nand NAND2_22415 ( P2_R1203_U173 , P2_R1203_U250 , P2_R1203_U249 );
nand NAND2_22416 ( P2_R1203_U174 , P2_R1203_U246 , P2_R1203_U245 );
and AND2_22417 ( P2_R1203_U175 , P2_R1203_U476 , P2_R1203_U475 );
nand NAND2_22418 ( P2_R1203_U176 , P2_R1203_U166 , P2_R1203_U165 );
not NOT1_22419 ( P2_R1203_U177 , P2_R1203_U83 );
not NOT1_22420 ( P2_R1203_U178 , P2_R1203_U28 );
not NOT1_22421 ( P2_R1203_U179 , P2_R1203_U38 );
nand NAND2_22422 ( P2_R1203_U180 , P2_U3459 , P2_R1203_U49 );
nand NAND2_22423 ( P2_R1203_U181 , P2_U3474 , P2_R1203_U59 );
nand NAND2_22424 ( P2_R1203_U182 , P2_U3955 , P2_R1203_U74 );
nand NAND2_22425 ( P2_R1203_U183 , P2_U3951 , P2_R1203_U82 );
nand NAND2_22426 ( P2_R1203_U184 , P2_U3435 , P2_R1203_U27 );
nand NAND2_22427 ( P2_R1203_U185 , P2_U3444 , P2_R1203_U33 );
nand NAND2_22428 ( P2_R1203_U186 , P2_U3450 , P2_R1203_U37 );
not NOT1_22429 ( P2_R1203_U187 , P2_R1203_U61 );
not NOT1_22430 ( P2_R1203_U188 , P2_R1203_U76 );
not NOT1_22431 ( P2_R1203_U189 , P2_R1203_U35 );
not NOT1_22432 ( P2_R1203_U190 , P2_R1203_U50 );
not NOT1_22433 ( P2_R1203_U191 , P2_R1203_U166 );
nand NAND2_22434 ( P2_R1203_U192 , P2_U3080 , P2_R1203_U166 );
not NOT1_22435 ( P2_R1203_U193 , P2_R1203_U44 );
nand NAND2_22436 ( P2_R1203_U194 , P2_U3438 , P2_R1203_U29 );
nand NAND2_22437 ( P2_R1203_U195 , P2_R1203_U114 , P2_R1203_U44 );
nand NAND2_22438 ( P2_R1203_U196 , P2_R1203_U29 , P2_R1203_U28 );
nand NAND2_22439 ( P2_R1203_U197 , P2_R1203_U196 , P2_R1203_U26 );
nand NAND2_22440 ( P2_R1203_U198 , P2_U3066 , P2_R1203_U178 );
not NOT1_22441 ( P2_R1203_U199 , P2_R1203_U154 );
nand NAND2_22442 ( P2_R1203_U200 , P2_U3447 , P2_R1203_U32 );
nand NAND2_22443 ( P2_R1203_U201 , P2_U3073 , P2_R1203_U30 );
nand NAND2_22444 ( P2_R1203_U202 , P2_U3069 , P2_R1203_U22 );
nand NAND2_22445 ( P2_R1203_U203 , P2_R1203_U189 , P2_R1203_U185 );
nand NAND2_22446 ( P2_R1203_U204 , P2_R1203_U6 , P2_R1203_U203 );
nand NAND2_22447 ( P2_R1203_U205 , P2_U3441 , P2_R1203_U34 );
nand NAND2_22448 ( P2_R1203_U206 , P2_U3447 , P2_R1203_U32 );
nand NAND2_22449 ( P2_R1203_U207 , P2_R1203_U154 , P2_R1203_U116 );
nand NAND2_22450 ( P2_R1203_U208 , P2_R1203_U206 , P2_R1203_U204 );
not NOT1_22451 ( P2_R1203_U209 , P2_R1203_U42 );
nand NAND2_22452 ( P2_R1203_U210 , P2_U3453 , P2_R1203_U39 );
nand NAND2_22453 ( P2_R1203_U211 , P2_R1203_U117 , P2_R1203_U42 );
nand NAND2_22454 ( P2_R1203_U212 , P2_R1203_U39 , P2_R1203_U38 );
nand NAND2_22455 ( P2_R1203_U213 , P2_R1203_U212 , P2_R1203_U36 );
nand NAND2_22456 ( P2_R1203_U214 , P2_U3086 , P2_R1203_U179 );
not NOT1_22457 ( P2_R1203_U215 , P2_R1203_U150 );
nand NAND2_22458 ( P2_R1203_U216 , P2_U3456 , P2_R1203_U41 );
nand NAND2_22459 ( P2_R1203_U217 , P2_R1203_U216 , P2_R1203_U50 );
nand NAND2_22460 ( P2_R1203_U218 , P2_R1203_U209 , P2_R1203_U38 );
nand NAND2_22461 ( P2_R1203_U219 , P2_R1203_U120 , P2_R1203_U218 );
nand NAND2_22462 ( P2_R1203_U220 , P2_R1203_U42 , P2_R1203_U186 );
nand NAND2_22463 ( P2_R1203_U221 , P2_R1203_U119 , P2_R1203_U220 );
nand NAND2_22464 ( P2_R1203_U222 , P2_R1203_U38 , P2_R1203_U186 );
nand NAND2_22465 ( P2_R1203_U223 , P2_R1203_U205 , P2_R1203_U154 );
not NOT1_22466 ( P2_R1203_U224 , P2_R1203_U43 );
nand NAND2_22467 ( P2_R1203_U225 , P2_U3069 , P2_R1203_U22 );
nand NAND2_22468 ( P2_R1203_U226 , P2_R1203_U224 , P2_R1203_U225 );
nand NAND2_22469 ( P2_R1203_U227 , P2_R1203_U122 , P2_R1203_U226 );
nand NAND2_22470 ( P2_R1203_U228 , P2_R1203_U43 , P2_R1203_U185 );
nand NAND2_22471 ( P2_R1203_U229 , P2_U3447 , P2_R1203_U32 );
nand NAND2_22472 ( P2_R1203_U230 , P2_R1203_U121 , P2_R1203_U228 );
nand NAND2_22473 ( P2_R1203_U231 , P2_U3069 , P2_R1203_U22 );
nand NAND2_22474 ( P2_R1203_U232 , P2_R1203_U185 , P2_R1203_U231 );
nand NAND2_22475 ( P2_R1203_U233 , P2_R1203_U205 , P2_R1203_U35 );
nand NAND2_22476 ( P2_R1203_U234 , P2_R1203_U193 , P2_R1203_U28 );
nand NAND2_22477 ( P2_R1203_U235 , P2_R1203_U124 , P2_R1203_U234 );
nand NAND2_22478 ( P2_R1203_U236 , P2_R1203_U44 , P2_R1203_U184 );
nand NAND2_22479 ( P2_R1203_U237 , P2_R1203_U123 , P2_R1203_U236 );
nand NAND2_22480 ( P2_R1203_U238 , P2_R1203_U28 , P2_R1203_U184 );
nand NAND2_22481 ( P2_R1203_U239 , P2_U3462 , P2_R1203_U48 );
nand NAND2_22482 ( P2_R1203_U240 , P2_U3065 , P2_R1203_U47 );
nand NAND2_22483 ( P2_R1203_U241 , P2_U3064 , P2_R1203_U46 );
nand NAND2_22484 ( P2_R1203_U242 , P2_R1203_U190 , P2_R1203_U180 );
nand NAND2_22485 ( P2_R1203_U243 , P2_R1203_U7 , P2_R1203_U242 );
nand NAND2_22486 ( P2_R1203_U244 , P2_U3462 , P2_R1203_U48 );
nand NAND2_22487 ( P2_R1203_U245 , P2_R1203_U150 , P2_R1203_U125 );
nand NAND2_22488 ( P2_R1203_U246 , P2_R1203_U244 , P2_R1203_U243 );
not NOT1_22489 ( P2_R1203_U247 , P2_R1203_U174 );
nand NAND2_22490 ( P2_R1203_U248 , P2_U3465 , P2_R1203_U52 );
nand NAND2_22491 ( P2_R1203_U249 , P2_R1203_U248 , P2_R1203_U174 );
nand NAND2_22492 ( P2_R1203_U250 , P2_U3074 , P2_R1203_U51 );
not NOT1_22493 ( P2_R1203_U251 , P2_R1203_U173 );
nand NAND2_22494 ( P2_R1203_U252 , P2_U3468 , P2_R1203_U54 );
nand NAND2_22495 ( P2_R1203_U253 , P2_R1203_U252 , P2_R1203_U173 );
nand NAND2_22496 ( P2_R1203_U254 , P2_U3082 , P2_R1203_U53 );
not NOT1_22497 ( P2_R1203_U255 , P2_R1203_U172 );
nand NAND2_22498 ( P2_R1203_U256 , P2_U3477 , P2_R1203_U58 );
nand NAND2_22499 ( P2_R1203_U257 , P2_U3075 , P2_R1203_U55 );
nand NAND2_22500 ( P2_R1203_U258 , P2_U3076 , P2_R1203_U56 );
nand NAND2_22501 ( P2_R1203_U259 , P2_R1203_U187 , P2_R1203_U8 );
nand NAND2_22502 ( P2_R1203_U260 , P2_R1203_U9 , P2_R1203_U259 );
nand NAND2_22503 ( P2_R1203_U261 , P2_U3471 , P2_R1203_U60 );
nand NAND2_22504 ( P2_R1203_U262 , P2_U3477 , P2_R1203_U58 );
nand NAND2_22505 ( P2_R1203_U263 , P2_R1203_U126 , P2_R1203_U172 );
nand NAND2_22506 ( P2_R1203_U264 , P2_R1203_U262 , P2_R1203_U260 );
not NOT1_22507 ( P2_R1203_U265 , P2_R1203_U169 );
nand NAND2_22508 ( P2_R1203_U266 , P2_U3480 , P2_R1203_U63 );
nand NAND2_22509 ( P2_R1203_U267 , P2_R1203_U266 , P2_R1203_U169 );
nand NAND2_22510 ( P2_R1203_U268 , P2_U3071 , P2_R1203_U62 );
not NOT1_22511 ( P2_R1203_U269 , P2_R1203_U64 );
nand NAND2_22512 ( P2_R1203_U270 , P2_R1203_U269 , P2_R1203_U65 );
nand NAND2_22513 ( P2_R1203_U271 , P2_R1203_U270 , P2_R1203_U168 );
nand NAND2_22514 ( P2_R1203_U272 , P2_U3084 , P2_R1203_U64 );
not NOT1_22515 ( P2_R1203_U273 , P2_R1203_U167 );
nand NAND2_22516 ( P2_R1203_U274 , P2_U3485 , P2_R1203_U67 );
nand NAND2_22517 ( P2_R1203_U275 , P2_R1203_U274 , P2_R1203_U167 );
nand NAND2_22518 ( P2_R1203_U276 , P2_U3083 , P2_R1203_U66 );
not NOT1_22519 ( P2_R1203_U277 , P2_R1203_U164 );
nand NAND2_22520 ( P2_R1203_U278 , P2_U3957 , P2_R1203_U69 );
nand NAND2_22521 ( P2_R1203_U279 , P2_R1203_U278 , P2_R1203_U164 );
nand NAND2_22522 ( P2_R1203_U280 , P2_U3078 , P2_R1203_U68 );
not NOT1_22523 ( P2_R1203_U281 , P2_R1203_U163 );
nand NAND2_22524 ( P2_R1203_U282 , P2_U3954 , P2_R1203_U73 );
nand NAND2_22525 ( P2_R1203_U283 , P2_U3068 , P2_R1203_U70 );
nand NAND2_22526 ( P2_R1203_U284 , P2_U3063 , P2_R1203_U71 );
nand NAND2_22527 ( P2_R1203_U285 , P2_R1203_U188 , P2_R1203_U10 );
nand NAND2_22528 ( P2_R1203_U286 , P2_R1203_U11 , P2_R1203_U285 );
nand NAND2_22529 ( P2_R1203_U287 , P2_U3956 , P2_R1203_U75 );
nand NAND2_22530 ( P2_R1203_U288 , P2_U3954 , P2_R1203_U73 );
nand NAND2_22531 ( P2_R1203_U289 , P2_R1203_U127 , P2_R1203_U163 );
nand NAND2_22532 ( P2_R1203_U290 , P2_R1203_U288 , P2_R1203_U286 );
not NOT1_22533 ( P2_R1203_U291 , P2_R1203_U160 );
nand NAND2_22534 ( P2_R1203_U292 , P2_U3953 , P2_R1203_U78 );
nand NAND2_22535 ( P2_R1203_U293 , P2_R1203_U292 , P2_R1203_U160 );
nand NAND2_22536 ( P2_R1203_U294 , P2_U3067 , P2_R1203_U77 );
not NOT1_22537 ( P2_R1203_U295 , P2_R1203_U159 );
nand NAND2_22538 ( P2_R1203_U296 , P2_U3952 , P2_R1203_U80 );
nand NAND2_22539 ( P2_R1203_U297 , P2_R1203_U296 , P2_R1203_U159 );
nand NAND2_22540 ( P2_R1203_U298 , P2_U3060 , P2_R1203_U79 );
not NOT1_22541 ( P2_R1203_U299 , P2_R1203_U88 );
nand NAND2_22542 ( P2_R1203_U300 , P2_U3950 , P2_R1203_U84 );
nand NAND3_22543 ( P2_R1203_U301 , P2_R1203_U88 , P2_R1203_U183 , P2_R1203_U300 );
nand NAND2_22544 ( P2_R1203_U302 , P2_R1203_U84 , P2_R1203_U83 );
nand NAND2_22545 ( P2_R1203_U303 , P2_R1203_U302 , P2_R1203_U81 );
nand NAND2_22546 ( P2_R1203_U304 , P2_U3055 , P2_R1203_U177 );
not NOT1_22547 ( P2_R1203_U305 , P2_R1203_U87 );
nand NAND2_22548 ( P2_R1203_U306 , P2_U3056 , P2_R1203_U85 );
nand NAND2_22549 ( P2_R1203_U307 , P2_R1203_U305 , P2_R1203_U306 );
nand NAND2_22550 ( P2_R1203_U308 , P2_U3949 , P2_R1203_U86 );
nand NAND2_22551 ( P2_R1203_U309 , P2_U3949 , P2_R1203_U86 );
nand NAND2_22552 ( P2_R1203_U310 , P2_R1203_U309 , P2_R1203_U87 );
nand NAND2_22553 ( P2_R1203_U311 , P2_U3056 , P2_R1203_U85 );
nand NAND2_22554 ( P2_R1203_U312 , P2_R1203_U129 , P2_R1203_U310 );
nand NAND2_22555 ( P2_R1203_U313 , P2_R1203_U299 , P2_R1203_U83 );
nand NAND2_22556 ( P2_R1203_U314 , P2_R1203_U133 , P2_R1203_U313 );
nand NAND2_22557 ( P2_R1203_U315 , P2_R1203_U88 , P2_R1203_U183 );
nand NAND2_22558 ( P2_R1203_U316 , P2_R1203_U132 , P2_R1203_U315 );
nand NAND2_22559 ( P2_R1203_U317 , P2_R1203_U83 , P2_R1203_U183 );
nand NAND2_22560 ( P2_R1203_U318 , P2_R1203_U287 , P2_R1203_U163 );
not NOT1_22561 ( P2_R1203_U319 , P2_R1203_U89 );
nand NAND2_22562 ( P2_R1203_U320 , P2_U3063 , P2_R1203_U71 );
nand NAND2_22563 ( P2_R1203_U321 , P2_R1203_U319 , P2_R1203_U320 );
nand NAND2_22564 ( P2_R1203_U322 , P2_R1203_U137 , P2_R1203_U321 );
nand NAND2_22565 ( P2_R1203_U323 , P2_R1203_U89 , P2_R1203_U182 );
nand NAND2_22566 ( P2_R1203_U324 , P2_U3954 , P2_R1203_U73 );
nand NAND2_22567 ( P2_R1203_U325 , P2_R1203_U136 , P2_R1203_U323 );
nand NAND2_22568 ( P2_R1203_U326 , P2_U3063 , P2_R1203_U71 );
nand NAND2_22569 ( P2_R1203_U327 , P2_R1203_U182 , P2_R1203_U326 );
nand NAND2_22570 ( P2_R1203_U328 , P2_R1203_U287 , P2_R1203_U76 );
nand NAND2_22571 ( P2_R1203_U329 , P2_R1203_U261 , P2_R1203_U172 );
not NOT1_22572 ( P2_R1203_U330 , P2_R1203_U90 );
nand NAND2_22573 ( P2_R1203_U331 , P2_U3076 , P2_R1203_U56 );
nand NAND2_22574 ( P2_R1203_U332 , P2_R1203_U330 , P2_R1203_U331 );
nand NAND2_22575 ( P2_R1203_U333 , P2_R1203_U144 , P2_R1203_U332 );
nand NAND2_22576 ( P2_R1203_U334 , P2_R1203_U90 , P2_R1203_U181 );
nand NAND2_22577 ( P2_R1203_U335 , P2_U3477 , P2_R1203_U58 );
nand NAND2_22578 ( P2_R1203_U336 , P2_R1203_U143 , P2_R1203_U334 );
nand NAND2_22579 ( P2_R1203_U337 , P2_U3076 , P2_R1203_U56 );
nand NAND2_22580 ( P2_R1203_U338 , P2_R1203_U181 , P2_R1203_U337 );
nand NAND2_22581 ( P2_R1203_U339 , P2_R1203_U261 , P2_R1203_U61 );
nand NAND2_22582 ( P2_R1203_U340 , P2_R1203_U216 , P2_R1203_U150 );
not NOT1_22583 ( P2_R1203_U341 , P2_R1203_U91 );
nand NAND2_22584 ( P2_R1203_U342 , P2_U3064 , P2_R1203_U46 );
nand NAND2_22585 ( P2_R1203_U343 , P2_R1203_U341 , P2_R1203_U342 );
nand NAND2_22586 ( P2_R1203_U344 , P2_R1203_U148 , P2_R1203_U343 );
nand NAND2_22587 ( P2_R1203_U345 , P2_R1203_U91 , P2_R1203_U180 );
nand NAND2_22588 ( P2_R1203_U346 , P2_U3462 , P2_R1203_U48 );
nand NAND2_22589 ( P2_R1203_U347 , P2_R1203_U147 , P2_R1203_U345 );
nand NAND2_22590 ( P2_R1203_U348 , P2_U3064 , P2_R1203_U46 );
nand NAND2_22591 ( P2_R1203_U349 , P2_R1203_U180 , P2_R1203_U348 );
nand NAND2_22592 ( P2_R1203_U350 , P2_U3079 , P2_R1203_U24 );
nand NAND2_22593 ( P2_R1203_U351 , P2_U3080 , P2_R1203_U165 );
nand NAND2_22594 ( P2_R1203_U352 , P2_R1203_U130 , P2_R1203_U307 );
nand NAND2_22595 ( P2_R1203_U353 , P2_U3456 , P2_R1203_U41 );
nand NAND2_22596 ( P2_R1203_U354 , P2_U3085 , P2_R1203_U40 );
nand NAND2_22597 ( P2_R1203_U355 , P2_R1203_U217 , P2_R1203_U150 );
nand NAND2_22598 ( P2_R1203_U356 , P2_R1203_U215 , P2_R1203_U149 );
nand NAND2_22599 ( P2_R1203_U357 , P2_U3453 , P2_R1203_U39 );
nand NAND2_22600 ( P2_R1203_U358 , P2_U3086 , P2_R1203_U36 );
nand NAND2_22601 ( P2_R1203_U359 , P2_U3453 , P2_R1203_U39 );
nand NAND2_22602 ( P2_R1203_U360 , P2_U3086 , P2_R1203_U36 );
nand NAND2_22603 ( P2_R1203_U361 , P2_R1203_U360 , P2_R1203_U359 );
nand NAND2_22604 ( P2_R1203_U362 , P2_U3450 , P2_R1203_U37 );
nand NAND2_22605 ( P2_R1203_U363 , P2_U3072 , P2_R1203_U21 );
nand NAND2_22606 ( P2_R1203_U364 , P2_R1203_U222 , P2_R1203_U42 );
nand NAND2_22607 ( P2_R1203_U365 , P2_R1203_U151 , P2_R1203_U209 );
nand NAND2_22608 ( P2_R1203_U366 , P2_U3447 , P2_R1203_U32 );
nand NAND2_22609 ( P2_R1203_U367 , P2_U3073 , P2_R1203_U30 );
nand NAND2_22610 ( P2_R1203_U368 , P2_R1203_U367 , P2_R1203_U366 );
nand NAND2_22611 ( P2_R1203_U369 , P2_U3444 , P2_R1203_U33 );
nand NAND2_22612 ( P2_R1203_U370 , P2_U3069 , P2_R1203_U22 );
nand NAND2_22613 ( P2_R1203_U371 , P2_R1203_U232 , P2_R1203_U43 );
nand NAND2_22614 ( P2_R1203_U372 , P2_R1203_U152 , P2_R1203_U224 );
nand NAND2_22615 ( P2_R1203_U373 , P2_U3441 , P2_R1203_U34 );
nand NAND2_22616 ( P2_R1203_U374 , P2_U3062 , P2_R1203_U31 );
nand NAND2_22617 ( P2_R1203_U375 , P2_R1203_U233 , P2_R1203_U154 );
nand NAND2_22618 ( P2_R1203_U376 , P2_R1203_U199 , P2_R1203_U153 );
nand NAND2_22619 ( P2_R1203_U377 , P2_U3438 , P2_R1203_U29 );
nand NAND2_22620 ( P2_R1203_U378 , P2_U3066 , P2_R1203_U26 );
nand NAND2_22621 ( P2_R1203_U379 , P2_U3438 , P2_R1203_U29 );
nand NAND2_22622 ( P2_R1203_U380 , P2_U3066 , P2_R1203_U26 );
nand NAND2_22623 ( P2_R1203_U381 , P2_R1203_U380 , P2_R1203_U379 );
nand NAND2_22624 ( P2_R1203_U382 , P2_U3435 , P2_R1203_U27 );
nand NAND2_22625 ( P2_R1203_U383 , P2_U3070 , P2_R1203_U23 );
nand NAND2_22626 ( P2_R1203_U384 , P2_R1203_U238 , P2_R1203_U44 );
nand NAND2_22627 ( P2_R1203_U385 , P2_R1203_U155 , P2_R1203_U193 );
nand NAND2_22628 ( P2_R1203_U386 , P2_U3960 , P2_R1203_U157 );
nand NAND2_22629 ( P2_R1203_U387 , P2_U3057 , P2_R1203_U156 );
nand NAND2_22630 ( P2_R1203_U388 , P2_U3960 , P2_R1203_U157 );
nand NAND2_22631 ( P2_R1203_U389 , P2_U3057 , P2_R1203_U156 );
nand NAND2_22632 ( P2_R1203_U390 , P2_R1203_U389 , P2_R1203_U388 );
nand NAND2_22633 ( P2_R1203_U391 , P2_U3949 , P2_R1203_U86 );
nand NAND2_22634 ( P2_R1203_U392 , P2_U3056 , P2_R1203_U85 );
not NOT1_22635 ( P2_R1203_U393 , P2_R1203_U131 );
nand NAND2_22636 ( P2_R1203_U394 , P2_R1203_U393 , P2_R1203_U305 );
nand NAND2_22637 ( P2_R1203_U395 , P2_R1203_U131 , P2_R1203_U87 );
nand NAND2_22638 ( P2_R1203_U396 , P2_U3950 , P2_R1203_U84 );
nand NAND2_22639 ( P2_R1203_U397 , P2_U3055 , P2_R1203_U81 );
nand NAND2_22640 ( P2_R1203_U398 , P2_U3950 , P2_R1203_U84 );
nand NAND2_22641 ( P2_R1203_U399 , P2_U3055 , P2_R1203_U81 );
nand NAND2_22642 ( P2_R1203_U400 , P2_R1203_U399 , P2_R1203_U398 );
nand NAND2_22643 ( P2_R1203_U401 , P2_U3951 , P2_R1203_U82 );
nand NAND2_22644 ( P2_R1203_U402 , P2_U3059 , P2_R1203_U45 );
nand NAND2_22645 ( P2_R1203_U403 , P2_R1203_U317 , P2_R1203_U88 );
nand NAND2_22646 ( P2_R1203_U404 , P2_R1203_U158 , P2_R1203_U299 );
nand NAND2_22647 ( P2_R1203_U405 , P2_U3952 , P2_R1203_U80 );
nand NAND2_22648 ( P2_R1203_U406 , P2_U3060 , P2_R1203_U79 );
not NOT1_22649 ( P2_R1203_U407 , P2_R1203_U134 );
nand NAND2_22650 ( P2_R1203_U408 , P2_R1203_U295 , P2_R1203_U407 );
nand NAND2_22651 ( P2_R1203_U409 , P2_R1203_U134 , P2_R1203_U159 );
nand NAND2_22652 ( P2_R1203_U410 , P2_U3953 , P2_R1203_U78 );
nand NAND2_22653 ( P2_R1203_U411 , P2_U3067 , P2_R1203_U77 );
not NOT1_22654 ( P2_R1203_U412 , P2_R1203_U135 );
nand NAND2_22655 ( P2_R1203_U413 , P2_R1203_U291 , P2_R1203_U412 );
nand NAND2_22656 ( P2_R1203_U414 , P2_R1203_U135 , P2_R1203_U160 );
nand NAND2_22657 ( P2_R1203_U415 , P2_U3954 , P2_R1203_U73 );
nand NAND2_22658 ( P2_R1203_U416 , P2_U3068 , P2_R1203_U70 );
nand NAND2_22659 ( P2_R1203_U417 , P2_R1203_U416 , P2_R1203_U415 );
nand NAND2_22660 ( P2_R1203_U418 , P2_U3955 , P2_R1203_U74 );
nand NAND2_22661 ( P2_R1203_U419 , P2_U3063 , P2_R1203_U71 );
nand NAND2_22662 ( P2_R1203_U420 , P2_R1203_U327 , P2_R1203_U89 );
nand NAND2_22663 ( P2_R1203_U421 , P2_R1203_U161 , P2_R1203_U319 );
nand NAND2_22664 ( P2_R1203_U422 , P2_U3956 , P2_R1203_U75 );
nand NAND2_22665 ( P2_R1203_U423 , P2_U3077 , P2_R1203_U72 );
nand NAND2_22666 ( P2_R1203_U424 , P2_R1203_U328 , P2_R1203_U163 );
nand NAND2_22667 ( P2_R1203_U425 , P2_R1203_U281 , P2_R1203_U162 );
nand NAND2_22668 ( P2_R1203_U426 , P2_U3957 , P2_R1203_U69 );
nand NAND2_22669 ( P2_R1203_U427 , P2_U3078 , P2_R1203_U68 );
not NOT1_22670 ( P2_R1203_U428 , P2_R1203_U138 );
nand NAND2_22671 ( P2_R1203_U429 , P2_R1203_U277 , P2_R1203_U428 );
nand NAND2_22672 ( P2_R1203_U430 , P2_R1203_U138 , P2_R1203_U164 );
nand NAND2_22673 ( P2_R1203_U431 , P2_U3432 , P2_R1203_U25 );
nand NAND2_22674 ( P2_R1203_U432 , P2_U3080 , P2_R1203_U165 );
not NOT1_22675 ( P2_R1203_U433 , P2_R1203_U139 );
nand NAND2_22676 ( P2_R1203_U434 , P2_R1203_U191 , P2_R1203_U433 );
nand NAND2_22677 ( P2_R1203_U435 , P2_R1203_U139 , P2_R1203_U166 );
nand NAND2_22678 ( P2_R1203_U436 , P2_U3485 , P2_R1203_U67 );
nand NAND2_22679 ( P2_R1203_U437 , P2_U3083 , P2_R1203_U66 );
not NOT1_22680 ( P2_R1203_U438 , P2_R1203_U140 );
nand NAND2_22681 ( P2_R1203_U439 , P2_R1203_U273 , P2_R1203_U438 );
nand NAND2_22682 ( P2_R1203_U440 , P2_R1203_U140 , P2_R1203_U167 );
nand NAND2_22683 ( P2_R1203_U441 , P2_U3483 , P2_R1203_U65 );
nand NAND2_22684 ( P2_R1203_U442 , P2_U3084 , P2_R1203_U168 );
not NOT1_22685 ( P2_R1203_U443 , P2_R1203_U141 );
nand NAND2_22686 ( P2_R1203_U444 , P2_R1203_U443 , P2_R1203_U269 );
nand NAND2_22687 ( P2_R1203_U445 , P2_R1203_U141 , P2_R1203_U64 );
nand NAND2_22688 ( P2_R1203_U446 , P2_U3480 , P2_R1203_U63 );
nand NAND2_22689 ( P2_R1203_U447 , P2_U3071 , P2_R1203_U62 );
not NOT1_22690 ( P2_R1203_U448 , P2_R1203_U142 );
nand NAND2_22691 ( P2_R1203_U449 , P2_R1203_U265 , P2_R1203_U448 );
nand NAND2_22692 ( P2_R1203_U450 , P2_R1203_U142 , P2_R1203_U169 );
nand NAND2_22693 ( P2_R1203_U451 , P2_U3477 , P2_R1203_U58 );
nand NAND2_22694 ( P2_R1203_U452 , P2_U3075 , P2_R1203_U55 );
nand NAND2_22695 ( P2_R1203_U453 , P2_R1203_U452 , P2_R1203_U451 );
nand NAND2_22696 ( P2_R1203_U454 , P2_U3474 , P2_R1203_U59 );
nand NAND2_22697 ( P2_R1203_U455 , P2_U3076 , P2_R1203_U56 );
nand NAND2_22698 ( P2_R1203_U456 , P2_R1203_U338 , P2_R1203_U90 );
nand NAND2_22699 ( P2_R1203_U457 , P2_R1203_U170 , P2_R1203_U330 );
nand NAND2_22700 ( P2_R1203_U458 , P2_U3471 , P2_R1203_U60 );
nand NAND2_22701 ( P2_R1203_U459 , P2_U3081 , P2_R1203_U57 );
nand NAND2_22702 ( P2_R1203_U460 , P2_R1203_U339 , P2_R1203_U172 );
nand NAND2_22703 ( P2_R1203_U461 , P2_R1203_U255 , P2_R1203_U171 );
nand NAND2_22704 ( P2_R1203_U462 , P2_U3468 , P2_R1203_U54 );
nand NAND2_22705 ( P2_R1203_U463 , P2_U3082 , P2_R1203_U53 );
not NOT1_22706 ( P2_R1203_U464 , P2_R1203_U145 );
nand NAND2_22707 ( P2_R1203_U465 , P2_R1203_U251 , P2_R1203_U464 );
nand NAND2_22708 ( P2_R1203_U466 , P2_R1203_U145 , P2_R1203_U173 );
nand NAND2_22709 ( P2_R1203_U467 , P2_U3465 , P2_R1203_U52 );
nand NAND2_22710 ( P2_R1203_U468 , P2_U3074 , P2_R1203_U51 );
not NOT1_22711 ( P2_R1203_U469 , P2_R1203_U146 );
nand NAND2_22712 ( P2_R1203_U470 , P2_R1203_U247 , P2_R1203_U469 );
nand NAND2_22713 ( P2_R1203_U471 , P2_R1203_U146 , P2_R1203_U174 );
nand NAND2_22714 ( P2_R1203_U472 , P2_U3462 , P2_R1203_U48 );
nand NAND2_22715 ( P2_R1203_U473 , P2_U3065 , P2_R1203_U47 );
nand NAND2_22716 ( P2_R1203_U474 , P2_R1203_U473 , P2_R1203_U472 );
nand NAND2_22717 ( P2_R1203_U475 , P2_U3459 , P2_R1203_U49 );
nand NAND2_22718 ( P2_R1203_U476 , P2_U3064 , P2_R1203_U46 );
nand NAND2_22719 ( P2_R1203_U477 , P2_R1203_U349 , P2_R1203_U91 );
nand NAND2_22720 ( P2_R1203_U478 , P2_R1203_U175 , P2_R1203_U341 );
and AND2_22721 ( P2_R1113_U6 , P2_R1113_U202 , P2_R1113_U201 );
and AND2_22722 ( P2_R1113_U7 , P2_R1113_U241 , P2_R1113_U240 );
and AND2_22723 ( P2_R1113_U8 , P2_R1113_U181 , P2_R1113_U256 );
and AND2_22724 ( P2_R1113_U9 , P2_R1113_U258 , P2_R1113_U257 );
and AND2_22725 ( P2_R1113_U10 , P2_R1113_U182 , P2_R1113_U282 );
and AND2_22726 ( P2_R1113_U11 , P2_R1113_U284 , P2_R1113_U283 );
nand NAND2_22727 ( P2_R1113_U12 , P2_R1113_U344 , P2_R1113_U347 );
nand NAND2_22728 ( P2_R1113_U13 , P2_R1113_U333 , P2_R1113_U336 );
nand NAND2_22729 ( P2_R1113_U14 , P2_R1113_U322 , P2_R1113_U325 );
nand NAND2_22730 ( P2_R1113_U15 , P2_R1113_U314 , P2_R1113_U316 );
nand NAND2_22731 ( P2_R1113_U16 , P2_R1113_U352 , P2_R1113_U312 );
nand NAND2_22732 ( P2_R1113_U17 , P2_R1113_U235 , P2_R1113_U237 );
nand NAND2_22733 ( P2_R1113_U18 , P2_R1113_U227 , P2_R1113_U230 );
nand NAND2_22734 ( P2_R1113_U19 , P2_R1113_U219 , P2_R1113_U221 );
nand NAND2_22735 ( P2_R1113_U20 , P2_R1113_U166 , P2_R1113_U350 );
not NOT1_22736 ( P2_R1113_U21 , P2_U3450 );
not NOT1_22737 ( P2_R1113_U22 , P2_U3444 );
not NOT1_22738 ( P2_R1113_U23 , P2_U3435 );
not NOT1_22739 ( P2_R1113_U24 , P2_U3427 );
not NOT1_22740 ( P2_R1113_U25 , P2_U3080 );
not NOT1_22741 ( P2_R1113_U26 , P2_U3438 );
not NOT1_22742 ( P2_R1113_U27 , P2_U3070 );
nand NAND2_22743 ( P2_R1113_U28 , P2_U3070 , P2_R1113_U23 );
not NOT1_22744 ( P2_R1113_U29 , P2_U3066 );
not NOT1_22745 ( P2_R1113_U30 , P2_U3447 );
not NOT1_22746 ( P2_R1113_U31 , P2_U3441 );
not NOT1_22747 ( P2_R1113_U32 , P2_U3073 );
not NOT1_22748 ( P2_R1113_U33 , P2_U3069 );
not NOT1_22749 ( P2_R1113_U34 , P2_U3062 );
nand NAND2_22750 ( P2_R1113_U35 , P2_U3062 , P2_R1113_U31 );
not NOT1_22751 ( P2_R1113_U36 , P2_U3453 );
not NOT1_22752 ( P2_R1113_U37 , P2_U3072 );
nand NAND2_22753 ( P2_R1113_U38 , P2_U3072 , P2_R1113_U21 );
not NOT1_22754 ( P2_R1113_U39 , P2_U3086 );
not NOT1_22755 ( P2_R1113_U40 , P2_U3456 );
not NOT1_22756 ( P2_R1113_U41 , P2_U3085 );
nand NAND2_22757 ( P2_R1113_U42 , P2_R1113_U208 , P2_R1113_U207 );
nand NAND2_22758 ( P2_R1113_U43 , P2_R1113_U35 , P2_R1113_U223 );
nand NAND3_22759 ( P2_R1113_U44 , P2_R1113_U192 , P2_R1113_U176 , P2_R1113_U351 );
not NOT1_22760 ( P2_R1113_U45 , P2_U3951 );
not NOT1_22761 ( P2_R1113_U46 , P2_U3459 );
not NOT1_22762 ( P2_R1113_U47 , P2_U3462 );
not NOT1_22763 ( P2_R1113_U48 , P2_U3065 );
not NOT1_22764 ( P2_R1113_U49 , P2_U3064 );
nand NAND2_22765 ( P2_R1113_U50 , P2_U3085 , P2_R1113_U40 );
not NOT1_22766 ( P2_R1113_U51 , P2_U3465 );
not NOT1_22767 ( P2_R1113_U52 , P2_U3074 );
not NOT1_22768 ( P2_R1113_U53 , P2_U3468 );
not NOT1_22769 ( P2_R1113_U54 , P2_U3082 );
not NOT1_22770 ( P2_R1113_U55 , P2_U3477 );
not NOT1_22771 ( P2_R1113_U56 , P2_U3474 );
not NOT1_22772 ( P2_R1113_U57 , P2_U3471 );
not NOT1_22773 ( P2_R1113_U58 , P2_U3075 );
not NOT1_22774 ( P2_R1113_U59 , P2_U3076 );
not NOT1_22775 ( P2_R1113_U60 , P2_U3081 );
nand NAND2_22776 ( P2_R1113_U61 , P2_U3081 , P2_R1113_U57 );
not NOT1_22777 ( P2_R1113_U62 , P2_U3480 );
not NOT1_22778 ( P2_R1113_U63 , P2_U3071 );
nand NAND2_22779 ( P2_R1113_U64 , P2_R1113_U268 , P2_R1113_U267 );
not NOT1_22780 ( P2_R1113_U65 , P2_U3084 );
not NOT1_22781 ( P2_R1113_U66 , P2_U3485 );
not NOT1_22782 ( P2_R1113_U67 , P2_U3083 );
not NOT1_22783 ( P2_R1113_U68 , P2_U3957 );
not NOT1_22784 ( P2_R1113_U69 , P2_U3078 );
not NOT1_22785 ( P2_R1113_U70 , P2_U3954 );
not NOT1_22786 ( P2_R1113_U71 , P2_U3955 );
not NOT1_22787 ( P2_R1113_U72 , P2_U3956 );
not NOT1_22788 ( P2_R1113_U73 , P2_U3068 );
not NOT1_22789 ( P2_R1113_U74 , P2_U3063 );
not NOT1_22790 ( P2_R1113_U75 , P2_U3077 );
nand NAND2_22791 ( P2_R1113_U76 , P2_U3077 , P2_R1113_U72 );
not NOT1_22792 ( P2_R1113_U77 , P2_U3953 );
not NOT1_22793 ( P2_R1113_U78 , P2_U3067 );
not NOT1_22794 ( P2_R1113_U79 , P2_U3952 );
not NOT1_22795 ( P2_R1113_U80 , P2_U3060 );
not NOT1_22796 ( P2_R1113_U81 , P2_U3950 );
not NOT1_22797 ( P2_R1113_U82 , P2_U3059 );
nand NAND2_22798 ( P2_R1113_U83 , P2_U3059 , P2_R1113_U45 );
not NOT1_22799 ( P2_R1113_U84 , P2_U3055 );
not NOT1_22800 ( P2_R1113_U85 , P2_U3949 );
not NOT1_22801 ( P2_R1113_U86 , P2_U3056 );
nand NAND2_22802 ( P2_R1113_U87 , P2_R1113_U128 , P2_R1113_U301 );
nand NAND2_22803 ( P2_R1113_U88 , P2_R1113_U298 , P2_R1113_U297 );
nand NAND2_22804 ( P2_R1113_U89 , P2_R1113_U76 , P2_R1113_U318 );
nand NAND2_22805 ( P2_R1113_U90 , P2_R1113_U61 , P2_R1113_U329 );
nand NAND2_22806 ( P2_R1113_U91 , P2_R1113_U50 , P2_R1113_U340 );
not NOT1_22807 ( P2_R1113_U92 , P2_U3079 );
nand NAND2_22808 ( P2_R1113_U93 , P2_R1113_U395 , P2_R1113_U394 );
nand NAND2_22809 ( P2_R1113_U94 , P2_R1113_U409 , P2_R1113_U408 );
nand NAND2_22810 ( P2_R1113_U95 , P2_R1113_U414 , P2_R1113_U413 );
nand NAND2_22811 ( P2_R1113_U96 , P2_R1113_U430 , P2_R1113_U429 );
nand NAND2_22812 ( P2_R1113_U97 , P2_R1113_U435 , P2_R1113_U434 );
nand NAND2_22813 ( P2_R1113_U98 , P2_R1113_U440 , P2_R1113_U439 );
nand NAND2_22814 ( P2_R1113_U99 , P2_R1113_U445 , P2_R1113_U444 );
nand NAND2_22815 ( P2_R1113_U100 , P2_R1113_U450 , P2_R1113_U449 );
nand NAND2_22816 ( P2_R1113_U101 , P2_R1113_U466 , P2_R1113_U465 );
nand NAND2_22817 ( P2_R1113_U102 , P2_R1113_U471 , P2_R1113_U470 );
nand NAND2_22818 ( P2_R1113_U103 , P2_R1113_U356 , P2_R1113_U355 );
nand NAND2_22819 ( P2_R1113_U104 , P2_R1113_U365 , P2_R1113_U364 );
nand NAND2_22820 ( P2_R1113_U105 , P2_R1113_U372 , P2_R1113_U371 );
nand NAND2_22821 ( P2_R1113_U106 , P2_R1113_U376 , P2_R1113_U375 );
nand NAND2_22822 ( P2_R1113_U107 , P2_R1113_U385 , P2_R1113_U384 );
nand NAND2_22823 ( P2_R1113_U108 , P2_R1113_U404 , P2_R1113_U403 );
nand NAND2_22824 ( P2_R1113_U109 , P2_R1113_U421 , P2_R1113_U420 );
nand NAND2_22825 ( P2_R1113_U110 , P2_R1113_U425 , P2_R1113_U424 );
nand NAND2_22826 ( P2_R1113_U111 , P2_R1113_U457 , P2_R1113_U456 );
nand NAND2_22827 ( P2_R1113_U112 , P2_R1113_U461 , P2_R1113_U460 );
nand NAND2_22828 ( P2_R1113_U113 , P2_R1113_U478 , P2_R1113_U477 );
and AND2_22829 ( P2_R1113_U114 , P2_R1113_U194 , P2_R1113_U184 );
and AND2_22830 ( P2_R1113_U115 , P2_R1113_U197 , P2_R1113_U198 );
and AND3_22831 ( P2_R1113_U116 , P2_R1113_U205 , P2_R1113_U200 , P2_R1113_U185 );
and AND2_22832 ( P2_R1113_U117 , P2_R1113_U210 , P2_R1113_U186 );
and AND2_22833 ( P2_R1113_U118 , P2_R1113_U213 , P2_R1113_U214 );
and AND3_22834 ( P2_R1113_U119 , P2_R1113_U358 , P2_R1113_U357 , P2_R1113_U38 );
and AND2_22835 ( P2_R1113_U120 , P2_R1113_U361 , P2_R1113_U186 );
and AND2_22836 ( P2_R1113_U121 , P2_R1113_U229 , P2_R1113_U6 );
and AND2_22837 ( P2_R1113_U122 , P2_R1113_U368 , P2_R1113_U185 );
and AND3_22838 ( P2_R1113_U123 , P2_R1113_U378 , P2_R1113_U377 , P2_R1113_U28 );
and AND2_22839 ( P2_R1113_U124 , P2_R1113_U381 , P2_R1113_U184 );
and AND3_22840 ( P2_R1113_U125 , P2_R1113_U239 , P2_R1113_U216 , P2_R1113_U180 );
and AND2_22841 ( P2_R1113_U126 , P2_R1113_U261 , P2_R1113_U8 );
and AND2_22842 ( P2_R1113_U127 , P2_R1113_U287 , P2_R1113_U10 );
and AND2_22843 ( P2_R1113_U128 , P2_R1113_U303 , P2_R1113_U304 );
and AND3_22844 ( P2_R1113_U129 , P2_R1113_U387 , P2_R1113_U386 , P2_R1113_U311 );
and AND2_22845 ( P2_R1113_U130 , P2_R1113_U308 , P2_R1113_U390 );
nand NAND2_22846 ( P2_R1113_U131 , P2_R1113_U392 , P2_R1113_U391 );
and AND3_22847 ( P2_R1113_U132 , P2_R1113_U397 , P2_R1113_U396 , P2_R1113_U83 );
and AND2_22848 ( P2_R1113_U133 , P2_R1113_U400 , P2_R1113_U183 );
nand NAND2_22849 ( P2_R1113_U134 , P2_R1113_U406 , P2_R1113_U405 );
nand NAND2_22850 ( P2_R1113_U135 , P2_R1113_U411 , P2_R1113_U410 );
and AND2_22851 ( P2_R1113_U136 , P2_R1113_U324 , P2_R1113_U11 );
and AND2_22852 ( P2_R1113_U137 , P2_R1113_U417 , P2_R1113_U182 );
nand NAND2_22853 ( P2_R1113_U138 , P2_R1113_U427 , P2_R1113_U426 );
nand NAND2_22854 ( P2_R1113_U139 , P2_R1113_U432 , P2_R1113_U431 );
nand NAND2_22855 ( P2_R1113_U140 , P2_R1113_U437 , P2_R1113_U436 );
nand NAND2_22856 ( P2_R1113_U141 , P2_R1113_U442 , P2_R1113_U441 );
nand NAND2_22857 ( P2_R1113_U142 , P2_R1113_U447 , P2_R1113_U446 );
and AND2_22858 ( P2_R1113_U143 , P2_R1113_U335 , P2_R1113_U9 );
and AND2_22859 ( P2_R1113_U144 , P2_R1113_U453 , P2_R1113_U181 );
nand NAND2_22860 ( P2_R1113_U145 , P2_R1113_U463 , P2_R1113_U462 );
nand NAND2_22861 ( P2_R1113_U146 , P2_R1113_U468 , P2_R1113_U467 );
and AND2_22862 ( P2_R1113_U147 , P2_R1113_U346 , P2_R1113_U7 );
and AND2_22863 ( P2_R1113_U148 , P2_R1113_U474 , P2_R1113_U180 );
and AND2_22864 ( P2_R1113_U149 , P2_R1113_U354 , P2_R1113_U353 );
nand NAND2_22865 ( P2_R1113_U150 , P2_R1113_U118 , P2_R1113_U211 );
and AND2_22866 ( P2_R1113_U151 , P2_R1113_U363 , P2_R1113_U362 );
and AND2_22867 ( P2_R1113_U152 , P2_R1113_U370 , P2_R1113_U369 );
and AND2_22868 ( P2_R1113_U153 , P2_R1113_U374 , P2_R1113_U373 );
nand NAND2_22869 ( P2_R1113_U154 , P2_R1113_U115 , P2_R1113_U195 );
and AND2_22870 ( P2_R1113_U155 , P2_R1113_U383 , P2_R1113_U382 );
not NOT1_22871 ( P2_R1113_U156 , P2_U3960 );
not NOT1_22872 ( P2_R1113_U157 , P2_U3057 );
and AND2_22873 ( P2_R1113_U158 , P2_R1113_U402 , P2_R1113_U401 );
nand NAND2_22874 ( P2_R1113_U159 , P2_R1113_U294 , P2_R1113_U293 );
nand NAND2_22875 ( P2_R1113_U160 , P2_R1113_U290 , P2_R1113_U289 );
and AND2_22876 ( P2_R1113_U161 , P2_R1113_U419 , P2_R1113_U418 );
and AND2_22877 ( P2_R1113_U162 , P2_R1113_U423 , P2_R1113_U422 );
nand NAND2_22878 ( P2_R1113_U163 , P2_R1113_U280 , P2_R1113_U279 );
nand NAND2_22879 ( P2_R1113_U164 , P2_R1113_U276 , P2_R1113_U275 );
not NOT1_22880 ( P2_R1113_U165 , P2_U3432 );
nand NAND2_22881 ( P2_R1113_U166 , P2_U3427 , P2_R1113_U92 );
nand NAND2_22882 ( P2_R1113_U167 , P2_R1113_U272 , P2_R1113_U271 );
not NOT1_22883 ( P2_R1113_U168 , P2_U3483 );
nand NAND2_22884 ( P2_R1113_U169 , P2_R1113_U264 , P2_R1113_U263 );
and AND2_22885 ( P2_R1113_U170 , P2_R1113_U455 , P2_R1113_U454 );
and AND2_22886 ( P2_R1113_U171 , P2_R1113_U459 , P2_R1113_U458 );
nand NAND2_22887 ( P2_R1113_U172 , P2_R1113_U254 , P2_R1113_U253 );
nand NAND2_22888 ( P2_R1113_U173 , P2_R1113_U250 , P2_R1113_U249 );
nand NAND2_22889 ( P2_R1113_U174 , P2_R1113_U246 , P2_R1113_U245 );
and AND2_22890 ( P2_R1113_U175 , P2_R1113_U476 , P2_R1113_U475 );
nand NAND2_22891 ( P2_R1113_U176 , P2_R1113_U166 , P2_R1113_U165 );
not NOT1_22892 ( P2_R1113_U177 , P2_R1113_U83 );
not NOT1_22893 ( P2_R1113_U178 , P2_R1113_U28 );
not NOT1_22894 ( P2_R1113_U179 , P2_R1113_U38 );
nand NAND2_22895 ( P2_R1113_U180 , P2_U3459 , P2_R1113_U49 );
nand NAND2_22896 ( P2_R1113_U181 , P2_U3474 , P2_R1113_U59 );
nand NAND2_22897 ( P2_R1113_U182 , P2_U3955 , P2_R1113_U74 );
nand NAND2_22898 ( P2_R1113_U183 , P2_U3951 , P2_R1113_U82 );
nand NAND2_22899 ( P2_R1113_U184 , P2_U3435 , P2_R1113_U27 );
nand NAND2_22900 ( P2_R1113_U185 , P2_U3444 , P2_R1113_U33 );
nand NAND2_22901 ( P2_R1113_U186 , P2_U3450 , P2_R1113_U37 );
not NOT1_22902 ( P2_R1113_U187 , P2_R1113_U61 );
not NOT1_22903 ( P2_R1113_U188 , P2_R1113_U76 );
not NOT1_22904 ( P2_R1113_U189 , P2_R1113_U35 );
not NOT1_22905 ( P2_R1113_U190 , P2_R1113_U50 );
not NOT1_22906 ( P2_R1113_U191 , P2_R1113_U166 );
nand NAND2_22907 ( P2_R1113_U192 , P2_U3080 , P2_R1113_U166 );
not NOT1_22908 ( P2_R1113_U193 , P2_R1113_U44 );
nand NAND2_22909 ( P2_R1113_U194 , P2_U3438 , P2_R1113_U29 );
nand NAND2_22910 ( P2_R1113_U195 , P2_R1113_U114 , P2_R1113_U44 );
nand NAND2_22911 ( P2_R1113_U196 , P2_R1113_U29 , P2_R1113_U28 );
nand NAND2_22912 ( P2_R1113_U197 , P2_R1113_U196 , P2_R1113_U26 );
nand NAND2_22913 ( P2_R1113_U198 , P2_U3066 , P2_R1113_U178 );
not NOT1_22914 ( P2_R1113_U199 , P2_R1113_U154 );
nand NAND2_22915 ( P2_R1113_U200 , P2_U3447 , P2_R1113_U32 );
nand NAND2_22916 ( P2_R1113_U201 , P2_U3073 , P2_R1113_U30 );
nand NAND2_22917 ( P2_R1113_U202 , P2_U3069 , P2_R1113_U22 );
nand NAND2_22918 ( P2_R1113_U203 , P2_R1113_U189 , P2_R1113_U185 );
nand NAND2_22919 ( P2_R1113_U204 , P2_R1113_U6 , P2_R1113_U203 );
nand NAND2_22920 ( P2_R1113_U205 , P2_U3441 , P2_R1113_U34 );
nand NAND2_22921 ( P2_R1113_U206 , P2_U3447 , P2_R1113_U32 );
nand NAND2_22922 ( P2_R1113_U207 , P2_R1113_U154 , P2_R1113_U116 );
nand NAND2_22923 ( P2_R1113_U208 , P2_R1113_U206 , P2_R1113_U204 );
not NOT1_22924 ( P2_R1113_U209 , P2_R1113_U42 );
nand NAND2_22925 ( P2_R1113_U210 , P2_U3453 , P2_R1113_U39 );
nand NAND2_22926 ( P2_R1113_U211 , P2_R1113_U117 , P2_R1113_U42 );
nand NAND2_22927 ( P2_R1113_U212 , P2_R1113_U39 , P2_R1113_U38 );
nand NAND2_22928 ( P2_R1113_U213 , P2_R1113_U212 , P2_R1113_U36 );
nand NAND2_22929 ( P2_R1113_U214 , P2_U3086 , P2_R1113_U179 );
not NOT1_22930 ( P2_R1113_U215 , P2_R1113_U150 );
nand NAND2_22931 ( P2_R1113_U216 , P2_U3456 , P2_R1113_U41 );
nand NAND2_22932 ( P2_R1113_U217 , P2_R1113_U216 , P2_R1113_U50 );
nand NAND2_22933 ( P2_R1113_U218 , P2_R1113_U209 , P2_R1113_U38 );
nand NAND2_22934 ( P2_R1113_U219 , P2_R1113_U120 , P2_R1113_U218 );
nand NAND2_22935 ( P2_R1113_U220 , P2_R1113_U42 , P2_R1113_U186 );
nand NAND2_22936 ( P2_R1113_U221 , P2_R1113_U119 , P2_R1113_U220 );
nand NAND2_22937 ( P2_R1113_U222 , P2_R1113_U38 , P2_R1113_U186 );
nand NAND2_22938 ( P2_R1113_U223 , P2_R1113_U205 , P2_R1113_U154 );
not NOT1_22939 ( P2_R1113_U224 , P2_R1113_U43 );
nand NAND2_22940 ( P2_R1113_U225 , P2_U3069 , P2_R1113_U22 );
nand NAND2_22941 ( P2_R1113_U226 , P2_R1113_U224 , P2_R1113_U225 );
nand NAND2_22942 ( P2_R1113_U227 , P2_R1113_U122 , P2_R1113_U226 );
nand NAND2_22943 ( P2_R1113_U228 , P2_R1113_U43 , P2_R1113_U185 );
nand NAND2_22944 ( P2_R1113_U229 , P2_U3447 , P2_R1113_U32 );
nand NAND2_22945 ( P2_R1113_U230 , P2_R1113_U121 , P2_R1113_U228 );
nand NAND2_22946 ( P2_R1113_U231 , P2_U3069 , P2_R1113_U22 );
nand NAND2_22947 ( P2_R1113_U232 , P2_R1113_U185 , P2_R1113_U231 );
nand NAND2_22948 ( P2_R1113_U233 , P2_R1113_U205 , P2_R1113_U35 );
nand NAND2_22949 ( P2_R1113_U234 , P2_R1113_U193 , P2_R1113_U28 );
nand NAND2_22950 ( P2_R1113_U235 , P2_R1113_U124 , P2_R1113_U234 );
nand NAND2_22951 ( P2_R1113_U236 , P2_R1113_U44 , P2_R1113_U184 );
nand NAND2_22952 ( P2_R1113_U237 , P2_R1113_U123 , P2_R1113_U236 );
nand NAND2_22953 ( P2_R1113_U238 , P2_R1113_U28 , P2_R1113_U184 );
nand NAND2_22954 ( P2_R1113_U239 , P2_U3462 , P2_R1113_U48 );
nand NAND2_22955 ( P2_R1113_U240 , P2_U3065 , P2_R1113_U47 );
nand NAND2_22956 ( P2_R1113_U241 , P2_U3064 , P2_R1113_U46 );
nand NAND2_22957 ( P2_R1113_U242 , P2_R1113_U190 , P2_R1113_U180 );
nand NAND2_22958 ( P2_R1113_U243 , P2_R1113_U7 , P2_R1113_U242 );
nand NAND2_22959 ( P2_R1113_U244 , P2_U3462 , P2_R1113_U48 );
nand NAND2_22960 ( P2_R1113_U245 , P2_R1113_U150 , P2_R1113_U125 );
nand NAND2_22961 ( P2_R1113_U246 , P2_R1113_U244 , P2_R1113_U243 );
not NOT1_22962 ( P2_R1113_U247 , P2_R1113_U174 );
nand NAND2_22963 ( P2_R1113_U248 , P2_U3465 , P2_R1113_U52 );
nand NAND2_22964 ( P2_R1113_U249 , P2_R1113_U248 , P2_R1113_U174 );
nand NAND2_22965 ( P2_R1113_U250 , P2_U3074 , P2_R1113_U51 );
not NOT1_22966 ( P2_R1113_U251 , P2_R1113_U173 );
nand NAND2_22967 ( P2_R1113_U252 , P2_U3468 , P2_R1113_U54 );
nand NAND2_22968 ( P2_R1113_U253 , P2_R1113_U252 , P2_R1113_U173 );
nand NAND2_22969 ( P2_R1113_U254 , P2_U3082 , P2_R1113_U53 );
not NOT1_22970 ( P2_R1113_U255 , P2_R1113_U172 );
nand NAND2_22971 ( P2_R1113_U256 , P2_U3477 , P2_R1113_U58 );
nand NAND2_22972 ( P2_R1113_U257 , P2_U3075 , P2_R1113_U55 );
nand NAND2_22973 ( P2_R1113_U258 , P2_U3076 , P2_R1113_U56 );
nand NAND2_22974 ( P2_R1113_U259 , P2_R1113_U187 , P2_R1113_U8 );
nand NAND2_22975 ( P2_R1113_U260 , P2_R1113_U9 , P2_R1113_U259 );
nand NAND2_22976 ( P2_R1113_U261 , P2_U3471 , P2_R1113_U60 );
nand NAND2_22977 ( P2_R1113_U262 , P2_U3477 , P2_R1113_U58 );
nand NAND2_22978 ( P2_R1113_U263 , P2_R1113_U126 , P2_R1113_U172 );
nand NAND2_22979 ( P2_R1113_U264 , P2_R1113_U262 , P2_R1113_U260 );
not NOT1_22980 ( P2_R1113_U265 , P2_R1113_U169 );
nand NAND2_22981 ( P2_R1113_U266 , P2_U3480 , P2_R1113_U63 );
nand NAND2_22982 ( P2_R1113_U267 , P2_R1113_U266 , P2_R1113_U169 );
nand NAND2_22983 ( P2_R1113_U268 , P2_U3071 , P2_R1113_U62 );
not NOT1_22984 ( P2_R1113_U269 , P2_R1113_U64 );
nand NAND2_22985 ( P2_R1113_U270 , P2_R1113_U269 , P2_R1113_U65 );
nand NAND2_22986 ( P2_R1113_U271 , P2_R1113_U270 , P2_R1113_U168 );
nand NAND2_22987 ( P2_R1113_U272 , P2_U3084 , P2_R1113_U64 );
not NOT1_22988 ( P2_R1113_U273 , P2_R1113_U167 );
nand NAND2_22989 ( P2_R1113_U274 , P2_U3485 , P2_R1113_U67 );
nand NAND2_22990 ( P2_R1113_U275 , P2_R1113_U274 , P2_R1113_U167 );
nand NAND2_22991 ( P2_R1113_U276 , P2_U3083 , P2_R1113_U66 );
not NOT1_22992 ( P2_R1113_U277 , P2_R1113_U164 );
nand NAND2_22993 ( P2_R1113_U278 , P2_U3957 , P2_R1113_U69 );
nand NAND2_22994 ( P2_R1113_U279 , P2_R1113_U278 , P2_R1113_U164 );
nand NAND2_22995 ( P2_R1113_U280 , P2_U3078 , P2_R1113_U68 );
not NOT1_22996 ( P2_R1113_U281 , P2_R1113_U163 );
nand NAND2_22997 ( P2_R1113_U282 , P2_U3954 , P2_R1113_U73 );
nand NAND2_22998 ( P2_R1113_U283 , P2_U3068 , P2_R1113_U70 );
nand NAND2_22999 ( P2_R1113_U284 , P2_U3063 , P2_R1113_U71 );
nand NAND2_23000 ( P2_R1113_U285 , P2_R1113_U188 , P2_R1113_U10 );
nand NAND2_23001 ( P2_R1113_U286 , P2_R1113_U11 , P2_R1113_U285 );
nand NAND2_23002 ( P2_R1113_U287 , P2_U3956 , P2_R1113_U75 );
nand NAND2_23003 ( P2_R1113_U288 , P2_U3954 , P2_R1113_U73 );
nand NAND2_23004 ( P2_R1113_U289 , P2_R1113_U127 , P2_R1113_U163 );
nand NAND2_23005 ( P2_R1113_U290 , P2_R1113_U288 , P2_R1113_U286 );
not NOT1_23006 ( P2_R1113_U291 , P2_R1113_U160 );
nand NAND2_23007 ( P2_R1113_U292 , P2_U3953 , P2_R1113_U78 );
nand NAND2_23008 ( P2_R1113_U293 , P2_R1113_U292 , P2_R1113_U160 );
nand NAND2_23009 ( P2_R1113_U294 , P2_U3067 , P2_R1113_U77 );
not NOT1_23010 ( P2_R1113_U295 , P2_R1113_U159 );
nand NAND2_23011 ( P2_R1113_U296 , P2_U3952 , P2_R1113_U80 );
nand NAND2_23012 ( P2_R1113_U297 , P2_R1113_U296 , P2_R1113_U159 );
nand NAND2_23013 ( P2_R1113_U298 , P2_U3060 , P2_R1113_U79 );
not NOT1_23014 ( P2_R1113_U299 , P2_R1113_U88 );
nand NAND2_23015 ( P2_R1113_U300 , P2_U3950 , P2_R1113_U84 );
nand NAND3_23016 ( P2_R1113_U301 , P2_R1113_U88 , P2_R1113_U183 , P2_R1113_U300 );
nand NAND2_23017 ( P2_R1113_U302 , P2_R1113_U84 , P2_R1113_U83 );
nand NAND2_23018 ( P2_R1113_U303 , P2_R1113_U302 , P2_R1113_U81 );
nand NAND2_23019 ( P2_R1113_U304 , P2_U3055 , P2_R1113_U177 );
not NOT1_23020 ( P2_R1113_U305 , P2_R1113_U87 );
nand NAND2_23021 ( P2_R1113_U306 , P2_U3056 , P2_R1113_U85 );
nand NAND2_23022 ( P2_R1113_U307 , P2_R1113_U305 , P2_R1113_U306 );
nand NAND2_23023 ( P2_R1113_U308 , P2_U3949 , P2_R1113_U86 );
nand NAND2_23024 ( P2_R1113_U309 , P2_U3949 , P2_R1113_U86 );
nand NAND2_23025 ( P2_R1113_U310 , P2_R1113_U309 , P2_R1113_U87 );
nand NAND2_23026 ( P2_R1113_U311 , P2_U3056 , P2_R1113_U85 );
nand NAND2_23027 ( P2_R1113_U312 , P2_R1113_U129 , P2_R1113_U310 );
nand NAND2_23028 ( P2_R1113_U313 , P2_R1113_U299 , P2_R1113_U83 );
nand NAND2_23029 ( P2_R1113_U314 , P2_R1113_U133 , P2_R1113_U313 );
nand NAND2_23030 ( P2_R1113_U315 , P2_R1113_U88 , P2_R1113_U183 );
nand NAND2_23031 ( P2_R1113_U316 , P2_R1113_U132 , P2_R1113_U315 );
nand NAND2_23032 ( P2_R1113_U317 , P2_R1113_U83 , P2_R1113_U183 );
nand NAND2_23033 ( P2_R1113_U318 , P2_R1113_U287 , P2_R1113_U163 );
not NOT1_23034 ( P2_R1113_U319 , P2_R1113_U89 );
nand NAND2_23035 ( P2_R1113_U320 , P2_U3063 , P2_R1113_U71 );
nand NAND2_23036 ( P2_R1113_U321 , P2_R1113_U319 , P2_R1113_U320 );
nand NAND2_23037 ( P2_R1113_U322 , P2_R1113_U137 , P2_R1113_U321 );
nand NAND2_23038 ( P2_R1113_U323 , P2_R1113_U89 , P2_R1113_U182 );
nand NAND2_23039 ( P2_R1113_U324 , P2_U3954 , P2_R1113_U73 );
nand NAND2_23040 ( P2_R1113_U325 , P2_R1113_U136 , P2_R1113_U323 );
nand NAND2_23041 ( P2_R1113_U326 , P2_U3063 , P2_R1113_U71 );
nand NAND2_23042 ( P2_R1113_U327 , P2_R1113_U182 , P2_R1113_U326 );
nand NAND2_23043 ( P2_R1113_U328 , P2_R1113_U287 , P2_R1113_U76 );
nand NAND2_23044 ( P2_R1113_U329 , P2_R1113_U261 , P2_R1113_U172 );
not NOT1_23045 ( P2_R1113_U330 , P2_R1113_U90 );
nand NAND2_23046 ( P2_R1113_U331 , P2_U3076 , P2_R1113_U56 );
nand NAND2_23047 ( P2_R1113_U332 , P2_R1113_U330 , P2_R1113_U331 );
nand NAND2_23048 ( P2_R1113_U333 , P2_R1113_U144 , P2_R1113_U332 );
nand NAND2_23049 ( P2_R1113_U334 , P2_R1113_U90 , P2_R1113_U181 );
nand NAND2_23050 ( P2_R1113_U335 , P2_U3477 , P2_R1113_U58 );
nand NAND2_23051 ( P2_R1113_U336 , P2_R1113_U143 , P2_R1113_U334 );
nand NAND2_23052 ( P2_R1113_U337 , P2_U3076 , P2_R1113_U56 );
nand NAND2_23053 ( P2_R1113_U338 , P2_R1113_U181 , P2_R1113_U337 );
nand NAND2_23054 ( P2_R1113_U339 , P2_R1113_U261 , P2_R1113_U61 );
nand NAND2_23055 ( P2_R1113_U340 , P2_R1113_U216 , P2_R1113_U150 );
not NOT1_23056 ( P2_R1113_U341 , P2_R1113_U91 );
nand NAND2_23057 ( P2_R1113_U342 , P2_U3064 , P2_R1113_U46 );
nand NAND2_23058 ( P2_R1113_U343 , P2_R1113_U341 , P2_R1113_U342 );
nand NAND2_23059 ( P2_R1113_U344 , P2_R1113_U148 , P2_R1113_U343 );
nand NAND2_23060 ( P2_R1113_U345 , P2_R1113_U91 , P2_R1113_U180 );
nand NAND2_23061 ( P2_R1113_U346 , P2_U3462 , P2_R1113_U48 );
nand NAND2_23062 ( P2_R1113_U347 , P2_R1113_U147 , P2_R1113_U345 );
nand NAND2_23063 ( P2_R1113_U348 , P2_U3064 , P2_R1113_U46 );
nand NAND2_23064 ( P2_R1113_U349 , P2_R1113_U180 , P2_R1113_U348 );
nand NAND2_23065 ( P2_R1113_U350 , P2_U3079 , P2_R1113_U24 );
nand NAND2_23066 ( P2_R1113_U351 , P2_U3080 , P2_R1113_U165 );
nand NAND2_23067 ( P2_R1113_U352 , P2_R1113_U130 , P2_R1113_U307 );
nand NAND2_23068 ( P2_R1113_U353 , P2_U3456 , P2_R1113_U41 );
nand NAND2_23069 ( P2_R1113_U354 , P2_U3085 , P2_R1113_U40 );
nand NAND2_23070 ( P2_R1113_U355 , P2_R1113_U217 , P2_R1113_U150 );
nand NAND2_23071 ( P2_R1113_U356 , P2_R1113_U215 , P2_R1113_U149 );
nand NAND2_23072 ( P2_R1113_U357 , P2_U3453 , P2_R1113_U39 );
nand NAND2_23073 ( P2_R1113_U358 , P2_U3086 , P2_R1113_U36 );
nand NAND2_23074 ( P2_R1113_U359 , P2_U3453 , P2_R1113_U39 );
nand NAND2_23075 ( P2_R1113_U360 , P2_U3086 , P2_R1113_U36 );
nand NAND2_23076 ( P2_R1113_U361 , P2_R1113_U360 , P2_R1113_U359 );
nand NAND2_23077 ( P2_R1113_U362 , P2_U3450 , P2_R1113_U37 );
nand NAND2_23078 ( P2_R1113_U363 , P2_U3072 , P2_R1113_U21 );
nand NAND2_23079 ( P2_R1113_U364 , P2_R1113_U222 , P2_R1113_U42 );
nand NAND2_23080 ( P2_R1113_U365 , P2_R1113_U151 , P2_R1113_U209 );
nand NAND2_23081 ( P2_R1113_U366 , P2_U3447 , P2_R1113_U32 );
nand NAND2_23082 ( P2_R1113_U367 , P2_U3073 , P2_R1113_U30 );
nand NAND2_23083 ( P2_R1113_U368 , P2_R1113_U367 , P2_R1113_U366 );
nand NAND2_23084 ( P2_R1113_U369 , P2_U3444 , P2_R1113_U33 );
nand NAND2_23085 ( P2_R1113_U370 , P2_U3069 , P2_R1113_U22 );
nand NAND2_23086 ( P2_R1113_U371 , P2_R1113_U232 , P2_R1113_U43 );
nand NAND2_23087 ( P2_R1113_U372 , P2_R1113_U152 , P2_R1113_U224 );
nand NAND2_23088 ( P2_R1113_U373 , P2_U3441 , P2_R1113_U34 );
nand NAND2_23089 ( P2_R1113_U374 , P2_U3062 , P2_R1113_U31 );
nand NAND2_23090 ( P2_R1113_U375 , P2_R1113_U233 , P2_R1113_U154 );
nand NAND2_23091 ( P2_R1113_U376 , P2_R1113_U199 , P2_R1113_U153 );
nand NAND2_23092 ( P2_R1113_U377 , P2_U3438 , P2_R1113_U29 );
nand NAND2_23093 ( P2_R1113_U378 , P2_U3066 , P2_R1113_U26 );
nand NAND2_23094 ( P2_R1113_U379 , P2_U3438 , P2_R1113_U29 );
nand NAND2_23095 ( P2_R1113_U380 , P2_U3066 , P2_R1113_U26 );
nand NAND2_23096 ( P2_R1113_U381 , P2_R1113_U380 , P2_R1113_U379 );
nand NAND2_23097 ( P2_R1113_U382 , P2_U3435 , P2_R1113_U27 );
nand NAND2_23098 ( P2_R1113_U383 , P2_U3070 , P2_R1113_U23 );
nand NAND2_23099 ( P2_R1113_U384 , P2_R1113_U238 , P2_R1113_U44 );
nand NAND2_23100 ( P2_R1113_U385 , P2_R1113_U155 , P2_R1113_U193 );
nand NAND2_23101 ( P2_R1113_U386 , P2_U3960 , P2_R1113_U157 );
nand NAND2_23102 ( P2_R1113_U387 , P2_U3057 , P2_R1113_U156 );
nand NAND2_23103 ( P2_R1113_U388 , P2_U3960 , P2_R1113_U157 );
nand NAND2_23104 ( P2_R1113_U389 , P2_U3057 , P2_R1113_U156 );
nand NAND2_23105 ( P2_R1113_U390 , P2_R1113_U389 , P2_R1113_U388 );
nand NAND2_23106 ( P2_R1113_U391 , P2_U3949 , P2_R1113_U86 );
nand NAND2_23107 ( P2_R1113_U392 , P2_U3056 , P2_R1113_U85 );
not NOT1_23108 ( P2_R1113_U393 , P2_R1113_U131 );
nand NAND2_23109 ( P2_R1113_U394 , P2_R1113_U393 , P2_R1113_U305 );
nand NAND2_23110 ( P2_R1113_U395 , P2_R1113_U131 , P2_R1113_U87 );
nand NAND2_23111 ( P2_R1113_U396 , P2_U3950 , P2_R1113_U84 );
nand NAND2_23112 ( P2_R1113_U397 , P2_U3055 , P2_R1113_U81 );
nand NAND2_23113 ( P2_R1113_U398 , P2_U3950 , P2_R1113_U84 );
nand NAND2_23114 ( P2_R1113_U399 , P2_U3055 , P2_R1113_U81 );
nand NAND2_23115 ( P2_R1113_U400 , P2_R1113_U399 , P2_R1113_U398 );
nand NAND2_23116 ( P2_R1113_U401 , P2_U3951 , P2_R1113_U82 );
nand NAND2_23117 ( P2_R1113_U402 , P2_U3059 , P2_R1113_U45 );
nand NAND2_23118 ( P2_R1113_U403 , P2_R1113_U317 , P2_R1113_U88 );
nand NAND2_23119 ( P2_R1113_U404 , P2_R1113_U158 , P2_R1113_U299 );
nand NAND2_23120 ( P2_R1113_U405 , P2_U3952 , P2_R1113_U80 );
nand NAND2_23121 ( P2_R1113_U406 , P2_U3060 , P2_R1113_U79 );
not NOT1_23122 ( P2_R1113_U407 , P2_R1113_U134 );
nand NAND2_23123 ( P2_R1113_U408 , P2_R1113_U295 , P2_R1113_U407 );
nand NAND2_23124 ( P2_R1113_U409 , P2_R1113_U134 , P2_R1113_U159 );
nand NAND2_23125 ( P2_R1113_U410 , P2_U3953 , P2_R1113_U78 );
nand NAND2_23126 ( P2_R1113_U411 , P2_U3067 , P2_R1113_U77 );
not NOT1_23127 ( P2_R1113_U412 , P2_R1113_U135 );
nand NAND2_23128 ( P2_R1113_U413 , P2_R1113_U291 , P2_R1113_U412 );
nand NAND2_23129 ( P2_R1113_U414 , P2_R1113_U135 , P2_R1113_U160 );
nand NAND2_23130 ( P2_R1113_U415 , P2_U3954 , P2_R1113_U73 );
nand NAND2_23131 ( P2_R1113_U416 , P2_U3068 , P2_R1113_U70 );
nand NAND2_23132 ( P2_R1113_U417 , P2_R1113_U416 , P2_R1113_U415 );
nand NAND2_23133 ( P2_R1113_U418 , P2_U3955 , P2_R1113_U74 );
nand NAND2_23134 ( P2_R1113_U419 , P2_U3063 , P2_R1113_U71 );
nand NAND2_23135 ( P2_R1113_U420 , P2_R1113_U327 , P2_R1113_U89 );
nand NAND2_23136 ( P2_R1113_U421 , P2_R1113_U161 , P2_R1113_U319 );
nand NAND2_23137 ( P2_R1113_U422 , P2_U3956 , P2_R1113_U75 );
nand NAND2_23138 ( P2_R1113_U423 , P2_U3077 , P2_R1113_U72 );
nand NAND2_23139 ( P2_R1113_U424 , P2_R1113_U328 , P2_R1113_U163 );
nand NAND2_23140 ( P2_R1113_U425 , P2_R1113_U281 , P2_R1113_U162 );
nand NAND2_23141 ( P2_R1113_U426 , P2_U3957 , P2_R1113_U69 );
nand NAND2_23142 ( P2_R1113_U427 , P2_U3078 , P2_R1113_U68 );
not NOT1_23143 ( P2_R1113_U428 , P2_R1113_U138 );
nand NAND2_23144 ( P2_R1113_U429 , P2_R1113_U277 , P2_R1113_U428 );
nand NAND2_23145 ( P2_R1113_U430 , P2_R1113_U138 , P2_R1113_U164 );
nand NAND2_23146 ( P2_R1113_U431 , P2_U3432 , P2_R1113_U25 );
nand NAND2_23147 ( P2_R1113_U432 , P2_U3080 , P2_R1113_U165 );
not NOT1_23148 ( P2_R1113_U433 , P2_R1113_U139 );
nand NAND2_23149 ( P2_R1113_U434 , P2_R1113_U191 , P2_R1113_U433 );
nand NAND2_23150 ( P2_R1113_U435 , P2_R1113_U139 , P2_R1113_U166 );
nand NAND2_23151 ( P2_R1113_U436 , P2_U3485 , P2_R1113_U67 );
nand NAND2_23152 ( P2_R1113_U437 , P2_U3083 , P2_R1113_U66 );
not NOT1_23153 ( P2_R1113_U438 , P2_R1113_U140 );
nand NAND2_23154 ( P2_R1113_U439 , P2_R1113_U273 , P2_R1113_U438 );
nand NAND2_23155 ( P2_R1113_U440 , P2_R1113_U140 , P2_R1113_U167 );
nand NAND2_23156 ( P2_R1113_U441 , P2_U3483 , P2_R1113_U65 );
nand NAND2_23157 ( P2_R1113_U442 , P2_U3084 , P2_R1113_U168 );
not NOT1_23158 ( P2_R1113_U443 , P2_R1113_U141 );
nand NAND2_23159 ( P2_R1113_U444 , P2_R1113_U443 , P2_R1113_U269 );
nand NAND2_23160 ( P2_R1113_U445 , P2_R1113_U141 , P2_R1113_U64 );
nand NAND2_23161 ( P2_R1113_U446 , P2_U3480 , P2_R1113_U63 );
nand NAND2_23162 ( P2_R1113_U447 , P2_U3071 , P2_R1113_U62 );
not NOT1_23163 ( P2_R1113_U448 , P2_R1113_U142 );
nand NAND2_23164 ( P2_R1113_U449 , P2_R1113_U265 , P2_R1113_U448 );
nand NAND2_23165 ( P2_R1113_U450 , P2_R1113_U142 , P2_R1113_U169 );
nand NAND2_23166 ( P2_R1113_U451 , P2_U3477 , P2_R1113_U58 );
nand NAND2_23167 ( P2_R1113_U452 , P2_U3075 , P2_R1113_U55 );
nand NAND2_23168 ( P2_R1113_U453 , P2_R1113_U452 , P2_R1113_U451 );
nand NAND2_23169 ( P2_R1113_U454 , P2_U3474 , P2_R1113_U59 );
nand NAND2_23170 ( P2_R1113_U455 , P2_U3076 , P2_R1113_U56 );
nand NAND2_23171 ( P2_R1113_U456 , P2_R1113_U338 , P2_R1113_U90 );
nand NAND2_23172 ( P2_R1113_U457 , P2_R1113_U170 , P2_R1113_U330 );
nand NAND2_23173 ( P2_R1113_U458 , P2_U3471 , P2_R1113_U60 );
nand NAND2_23174 ( P2_R1113_U459 , P2_U3081 , P2_R1113_U57 );
nand NAND2_23175 ( P2_R1113_U460 , P2_R1113_U339 , P2_R1113_U172 );
nand NAND2_23176 ( P2_R1113_U461 , P2_R1113_U255 , P2_R1113_U171 );
nand NAND2_23177 ( P2_R1113_U462 , P2_U3468 , P2_R1113_U54 );
nand NAND2_23178 ( P2_R1113_U463 , P2_U3082 , P2_R1113_U53 );
not NOT1_23179 ( P2_R1113_U464 , P2_R1113_U145 );
nand NAND2_23180 ( P2_R1113_U465 , P2_R1113_U251 , P2_R1113_U464 );
nand NAND2_23181 ( P2_R1113_U466 , P2_R1113_U145 , P2_R1113_U173 );
nand NAND2_23182 ( P2_R1113_U467 , P2_U3465 , P2_R1113_U52 );
nand NAND2_23183 ( P2_R1113_U468 , P2_U3074 , P2_R1113_U51 );
not NOT1_23184 ( P2_R1113_U469 , P2_R1113_U146 );
nand NAND2_23185 ( P2_R1113_U470 , P2_R1113_U247 , P2_R1113_U469 );
nand NAND2_23186 ( P2_R1113_U471 , P2_R1113_U146 , P2_R1113_U174 );
nand NAND2_23187 ( P2_R1113_U472 , P2_U3462 , P2_R1113_U48 );
nand NAND2_23188 ( P2_R1113_U473 , P2_U3065 , P2_R1113_U47 );
nand NAND2_23189 ( P2_R1113_U474 , P2_R1113_U473 , P2_R1113_U472 );
nand NAND2_23190 ( P2_R1113_U475 , P2_U3459 , P2_R1113_U49 );
nand NAND2_23191 ( P2_R1113_U476 , P2_U3064 , P2_R1113_U46 );
nand NAND2_23192 ( P2_R1113_U477 , P2_R1113_U349 , P2_R1113_U91 );
nand NAND2_23193 ( P2_R1113_U478 , P2_R1113_U175 , P2_R1113_U341 );
nor nor_23194 ( P3_SUB_598_U6 , P3_IR_REG_19_ , P3_IR_REG_20_ , P3_IR_REG_17_ , P3_IR_REG_18_ );
and AND2_23195 ( P3_SUB_598_U7 , P3_SUB_598_U136 , P3_SUB_598_U49 );
and AND2_23196 ( P3_SUB_598_U8 , P3_SUB_598_U134 , P3_SUB_598_U102 );
and AND2_23197 ( P3_SUB_598_U9 , P3_SUB_598_U133 , P3_SUB_598_U46 );
and AND2_23198 ( P3_SUB_598_U10 , P3_SUB_598_U132 , P3_SUB_598_U47 );
and AND2_23199 ( P3_SUB_598_U11 , P3_SUB_598_U130 , P3_SUB_598_U105 );
and AND2_23200 ( P3_SUB_598_U12 , P3_SUB_598_U129 , P3_SUB_598_U34 );
and AND2_23201 ( P3_SUB_598_U13 , P3_SUB_598_U128 , P3_SUB_598_U44 );
and AND2_23202 ( P3_SUB_598_U14 , P3_SUB_598_U126 , P3_SUB_598_U108 );
and AND2_23203 ( P3_SUB_598_U15 , P3_SUB_598_U125 , P3_SUB_598_U40 );
and AND2_23204 ( P3_SUB_598_U16 , P3_SUB_598_U124 , P3_SUB_598_U41 );
and AND2_23205 ( P3_SUB_598_U17 , P3_SUB_598_U122 , P3_SUB_598_U111 );
and AND2_23206 ( P3_SUB_598_U18 , P3_SUB_598_U121 , P3_SUB_598_U35 );
and AND2_23207 ( P3_SUB_598_U19 , P3_SUB_598_U120 , P3_SUB_598_U78 );
and AND2_23208 ( P3_SUB_598_U20 , P3_SUB_598_U65 , P3_SUB_598_U139 );
and AND2_23209 ( P3_SUB_598_U21 , P3_SUB_598_U118 , P3_SUB_598_U37 );
and AND2_23210 ( P3_SUB_598_U22 , P3_SUB_598_U117 , P3_SUB_598_U28 );
and AND2_23211 ( P3_SUB_598_U23 , P3_SUB_598_U100 , P3_SUB_598_U90 );
and AND2_23212 ( P3_SUB_598_U24 , P3_SUB_598_U99 , P3_SUB_598_U30 );
and AND2_23213 ( P3_SUB_598_U25 , P3_SUB_598_U98 , P3_SUB_598_U31 );
and AND2_23214 ( P3_SUB_598_U26 , P3_SUB_598_U96 , P3_SUB_598_U93 );
and AND2_23215 ( P3_SUB_598_U27 , P3_SUB_598_U95 , P3_SUB_598_U29 );
or OR3_23216 ( P3_SUB_598_U28 , P3_IR_REG_1_ , P3_IR_REG_0_ , P3_IR_REG_2_ );
nand NAND3_23217 ( P3_SUB_598_U29 , P3_SUB_598_U54 , P3_SUB_598_U140 , P3_SUB_598_U53 );
nand NAND2_23218 ( P3_SUB_598_U30 , P3_SUB_598_U55 , P3_SUB_598_U140 );
nand NAND2_23219 ( P3_SUB_598_U31 , P3_SUB_598_U56 , P3_SUB_598_U91 );
not NOT1_23220 ( P3_SUB_598_U32 , P3_IR_REG_7_ );
not NOT1_23221 ( P3_SUB_598_U33 , P3_IR_REG_3_ );
nand NAND4_23222 ( P3_SUB_598_U34 , P3_SUB_598_U60 , P3_SUB_598_U59 , P3_SUB_598_U58 , P3_SUB_598_U57 );
nand NAND2_23223 ( P3_SUB_598_U35 , P3_SUB_598_U62 , P3_SUB_598_U106 );
nand NAND2_23224 ( P3_SUB_598_U36 , P3_SUB_598_U63 , P3_SUB_598_U112 );
nand NAND2_23225 ( P3_SUB_598_U37 , P3_SUB_598_U114 , P3_SUB_598_U38 );
not NOT1_23226 ( P3_SUB_598_U38 , P3_IR_REG_29_ );
not NOT1_23227 ( P3_SUB_598_U39 , P3_IR_REG_27_ );
nand NAND2_23228 ( P3_SUB_598_U40 , P3_SUB_598_U106 , P3_SUB_598_U6 );
nand NAND2_23229 ( P3_SUB_598_U41 , P3_SUB_598_U66 , P3_SUB_598_U109 );
not NOT1_23230 ( P3_SUB_598_U42 , P3_IR_REG_24_ );
not NOT1_23231 ( P3_SUB_598_U43 , P3_IR_REG_23_ );
nand NAND2_23232 ( P3_SUB_598_U44 , P3_SUB_598_U67 , P3_SUB_598_U106 );
not NOT1_23233 ( P3_SUB_598_U45 , P3_IR_REG_19_ );
nand NAND2_23234 ( P3_SUB_598_U46 , P3_SUB_598_U68 , P3_SUB_598_U94 );
nand NAND2_23235 ( P3_SUB_598_U47 , P3_SUB_598_U69 , P3_SUB_598_U103 );
not NOT1_23236 ( P3_SUB_598_U48 , P3_IR_REG_15_ );
nand NAND2_23237 ( P3_SUB_598_U49 , P3_SUB_598_U70 , P3_SUB_598_U94 );
not NOT1_23238 ( P3_SUB_598_U50 , P3_IR_REG_11_ );
nand NAND2_23239 ( P3_SUB_598_U51 , P3_SUB_598_U156 , P3_SUB_598_U155 );
nand NAND2_23240 ( P3_SUB_598_U52 , P3_SUB_598_U146 , P3_SUB_598_U145 );
nor nor_23241 ( P3_SUB_598_U53 , P3_IR_REG_3_ , P3_IR_REG_4_ , P3_IR_REG_5_ , P3_IR_REG_6_ );
nor nor_23242 ( P3_SUB_598_U54 , P3_IR_REG_7_ , P3_IR_REG_8_ );
nor nor_23243 ( P3_SUB_598_U55 , P3_IR_REG_3_ , P3_IR_REG_4_ );
nor nor_23244 ( P3_SUB_598_U56 , P3_IR_REG_5_ , P3_IR_REG_6_ );
nor nor_23245 ( P3_SUB_598_U57 , P3_IR_REG_13_ , P3_IR_REG_14_ , P3_IR_REG_12_ , P3_IR_REG_10_ , P3_IR_REG_11_ );
nor nor_23246 ( P3_SUB_598_U58 , P3_IR_REG_15_ , P3_IR_REG_16_ , P3_IR_REG_1_ , P3_IR_REG_0_ );
nor nor_23247 ( P3_SUB_598_U59 , P3_IR_REG_2_ , P3_IR_REG_3_ , P3_IR_REG_4_ , P3_IR_REG_5_ );
nor nor_23248 ( P3_SUB_598_U60 , P3_IR_REG_6_ , P3_IR_REG_7_ , P3_IR_REG_8_ , P3_IR_REG_9_ );
nor nor_23249 ( P3_SUB_598_U61 , P3_IR_REG_23_ , P3_IR_REG_21_ , P3_IR_REG_22_ );
and AND3_23250 ( P3_SUB_598_U62 , P3_SUB_598_U6 , P3_SUB_598_U42 , P3_SUB_598_U61 );
nor nor_23251 ( P3_SUB_598_U63 , P3_IR_REG_25_ , P3_IR_REG_26_ , P3_IR_REG_27_ , P3_IR_REG_28_ );
nor nor_23252 ( P3_SUB_598_U64 , P3_IR_REG_25_ , P3_IR_REG_26_ );
and AND2_23253 ( P3_SUB_598_U65 , P3_SUB_598_U138 , P3_SUB_598_U36 );
nor nor_23254 ( P3_SUB_598_U66 , P3_IR_REG_21_ , P3_IR_REG_22_ );
nor nor_23255 ( P3_SUB_598_U67 , P3_IR_REG_17_ , P3_IR_REG_18_ );
nor nor_23256 ( P3_SUB_598_U68 , P3_IR_REG_10_ , P3_IR_REG_11_ , P3_IR_REG_12_ , P3_IR_REG_9_ );
nor nor_23257 ( P3_SUB_598_U69 , P3_IR_REG_13_ , P3_IR_REG_14_ );
nor nor_23258 ( P3_SUB_598_U70 , P3_IR_REG_10_ , P3_IR_REG_9_ );
not NOT1_23259 ( P3_SUB_598_U71 , P3_IR_REG_9_ );
and AND2_23260 ( P3_SUB_598_U72 , P3_SUB_598_U142 , P3_SUB_598_U141 );
not NOT1_23261 ( P3_SUB_598_U73 , P3_IR_REG_5_ );
and AND2_23262 ( P3_SUB_598_U74 , P3_SUB_598_U144 , P3_SUB_598_U143 );
not NOT1_23263 ( P3_SUB_598_U75 , P3_IR_REG_31_ );
not NOT1_23264 ( P3_SUB_598_U76 , P3_IR_REG_30_ );
and AND2_23265 ( P3_SUB_598_U77 , P3_SUB_598_U148 , P3_SUB_598_U147 );
nand NAND2_23266 ( P3_SUB_598_U78 , P3_SUB_598_U64 , P3_SUB_598_U112 );
and AND2_23267 ( P3_SUB_598_U79 , P3_SUB_598_U150 , P3_SUB_598_U149 );
not NOT1_23268 ( P3_SUB_598_U80 , P3_IR_REG_25_ );
and AND2_23269 ( P3_SUB_598_U81 , P3_SUB_598_U152 , P3_SUB_598_U151 );
not NOT1_23270 ( P3_SUB_598_U82 , P3_IR_REG_21_ );
and AND2_23271 ( P3_SUB_598_U83 , P3_SUB_598_U154 , P3_SUB_598_U153 );
not NOT1_23272 ( P3_SUB_598_U84 , P3_IR_REG_1_ );
not NOT1_23273 ( P3_SUB_598_U85 , P3_IR_REG_0_ );
not NOT1_23274 ( P3_SUB_598_U86 , P3_IR_REG_17_ );
and AND2_23275 ( P3_SUB_598_U87 , P3_SUB_598_U158 , P3_SUB_598_U157 );
not NOT1_23276 ( P3_SUB_598_U88 , P3_IR_REG_13_ );
and AND2_23277 ( P3_SUB_598_U89 , P3_SUB_598_U160 , P3_SUB_598_U159 );
nand NAND2_23278 ( P3_SUB_598_U90 , P3_SUB_598_U140 , P3_SUB_598_U33 );
not NOT1_23279 ( P3_SUB_598_U91 , P3_SUB_598_U30 );
not NOT1_23280 ( P3_SUB_598_U92 , P3_SUB_598_U31 );
nand NAND2_23281 ( P3_SUB_598_U93 , P3_SUB_598_U92 , P3_SUB_598_U32 );
not NOT1_23282 ( P3_SUB_598_U94 , P3_SUB_598_U29 );
nand NAND2_23283 ( P3_SUB_598_U95 , P3_IR_REG_8_ , P3_SUB_598_U93 );
nand NAND2_23284 ( P3_SUB_598_U96 , P3_IR_REG_7_ , P3_SUB_598_U31 );
nand NAND2_23285 ( P3_SUB_598_U97 , P3_SUB_598_U91 , P3_SUB_598_U73 );
nand NAND2_23286 ( P3_SUB_598_U98 , P3_IR_REG_6_ , P3_SUB_598_U97 );
nand NAND2_23287 ( P3_SUB_598_U99 , P3_IR_REG_4_ , P3_SUB_598_U90 );
nand NAND2_23288 ( P3_SUB_598_U100 , P3_IR_REG_3_ , P3_SUB_598_U28 );
not NOT1_23289 ( P3_SUB_598_U101 , P3_SUB_598_U49 );
nand NAND2_23290 ( P3_SUB_598_U102 , P3_SUB_598_U101 , P3_SUB_598_U50 );
not NOT1_23291 ( P3_SUB_598_U103 , P3_SUB_598_U46 );
not NOT1_23292 ( P3_SUB_598_U104 , P3_SUB_598_U47 );
nand NAND2_23293 ( P3_SUB_598_U105 , P3_SUB_598_U104 , P3_SUB_598_U48 );
not NOT1_23294 ( P3_SUB_598_U106 , P3_SUB_598_U34 );
not NOT1_23295 ( P3_SUB_598_U107 , P3_SUB_598_U44 );
nand NAND2_23296 ( P3_SUB_598_U108 , P3_SUB_598_U107 , P3_SUB_598_U45 );
not NOT1_23297 ( P3_SUB_598_U109 , P3_SUB_598_U40 );
not NOT1_23298 ( P3_SUB_598_U110 , P3_SUB_598_U41 );
nand NAND2_23299 ( P3_SUB_598_U111 , P3_SUB_598_U110 , P3_SUB_598_U43 );
not NOT1_23300 ( P3_SUB_598_U112 , P3_SUB_598_U35 );
not NOT1_23301 ( P3_SUB_598_U113 , P3_SUB_598_U78 );
not NOT1_23302 ( P3_SUB_598_U114 , P3_SUB_598_U36 );
not NOT1_23303 ( P3_SUB_598_U115 , P3_SUB_598_U37 );
or OR2_23304 ( P3_SUB_598_U116 , P3_IR_REG_1_ , P3_IR_REG_0_ );
nand NAND2_23305 ( P3_SUB_598_U117 , P3_IR_REG_2_ , P3_SUB_598_U116 );
nand NAND2_23306 ( P3_SUB_598_U118 , P3_IR_REG_29_ , P3_SUB_598_U36 );
nand NAND2_23307 ( P3_SUB_598_U119 , P3_SUB_598_U112 , P3_SUB_598_U80 );
nand NAND2_23308 ( P3_SUB_598_U120 , P3_IR_REG_26_ , P3_SUB_598_U119 );
nand NAND2_23309 ( P3_SUB_598_U121 , P3_IR_REG_24_ , P3_SUB_598_U111 );
nand NAND2_23310 ( P3_SUB_598_U122 , P3_IR_REG_23_ , P3_SUB_598_U41 );
nand NAND2_23311 ( P3_SUB_598_U123 , P3_SUB_598_U109 , P3_SUB_598_U82 );
nand NAND2_23312 ( P3_SUB_598_U124 , P3_IR_REG_22_ , P3_SUB_598_U123 );
nand NAND2_23313 ( P3_SUB_598_U125 , P3_IR_REG_20_ , P3_SUB_598_U108 );
nand NAND2_23314 ( P3_SUB_598_U126 , P3_IR_REG_19_ , P3_SUB_598_U44 );
nand NAND2_23315 ( P3_SUB_598_U127 , P3_SUB_598_U106 , P3_SUB_598_U86 );
nand NAND2_23316 ( P3_SUB_598_U128 , P3_IR_REG_18_ , P3_SUB_598_U127 );
nand NAND2_23317 ( P3_SUB_598_U129 , P3_IR_REG_16_ , P3_SUB_598_U105 );
nand NAND2_23318 ( P3_SUB_598_U130 , P3_IR_REG_15_ , P3_SUB_598_U47 );
nand NAND2_23319 ( P3_SUB_598_U131 , P3_SUB_598_U103 , P3_SUB_598_U88 );
nand NAND2_23320 ( P3_SUB_598_U132 , P3_IR_REG_14_ , P3_SUB_598_U131 );
nand NAND2_23321 ( P3_SUB_598_U133 , P3_IR_REG_12_ , P3_SUB_598_U102 );
nand NAND2_23322 ( P3_SUB_598_U134 , P3_IR_REG_11_ , P3_SUB_598_U49 );
nand NAND2_23323 ( P3_SUB_598_U135 , P3_SUB_598_U94 , P3_SUB_598_U71 );
nand NAND2_23324 ( P3_SUB_598_U136 , P3_IR_REG_10_ , P3_SUB_598_U135 );
nand NAND2_23325 ( P3_SUB_598_U137 , P3_SUB_598_U115 , P3_SUB_598_U76 );
nand NAND2_23326 ( P3_SUB_598_U138 , P3_IR_REG_27_ , P3_IR_REG_28_ );
nand NAND2_23327 ( P3_SUB_598_U139 , P3_IR_REG_28_ , P3_SUB_598_U78 );
not NOT1_23328 ( P3_SUB_598_U140 , P3_SUB_598_U28 );
nand NAND2_23329 ( P3_SUB_598_U141 , P3_IR_REG_9_ , P3_SUB_598_U29 );
nand NAND2_23330 ( P3_SUB_598_U142 , P3_SUB_598_U94 , P3_SUB_598_U71 );
nand NAND2_23331 ( P3_SUB_598_U143 , P3_IR_REG_5_ , P3_SUB_598_U30 );
nand NAND2_23332 ( P3_SUB_598_U144 , P3_SUB_598_U91 , P3_SUB_598_U73 );
nand NAND2_23333 ( P3_SUB_598_U145 , P3_SUB_598_U137 , P3_SUB_598_U75 );
nand NAND3_23334 ( P3_SUB_598_U146 , P3_SUB_598_U115 , P3_SUB_598_U76 , P3_IR_REG_31_ );
nand NAND2_23335 ( P3_SUB_598_U147 , P3_IR_REG_30_ , P3_SUB_598_U37 );
nand NAND2_23336 ( P3_SUB_598_U148 , P3_SUB_598_U115 , P3_SUB_598_U76 );
nand NAND2_23337 ( P3_SUB_598_U149 , P3_IR_REG_27_ , P3_SUB_598_U78 );
nand NAND2_23338 ( P3_SUB_598_U150 , P3_SUB_598_U113 , P3_SUB_598_U39 );
nand NAND2_23339 ( P3_SUB_598_U151 , P3_IR_REG_25_ , P3_SUB_598_U35 );
nand NAND2_23340 ( P3_SUB_598_U152 , P3_SUB_598_U112 , P3_SUB_598_U80 );
nand NAND2_23341 ( P3_SUB_598_U153 , P3_IR_REG_21_ , P3_SUB_598_U40 );
nand NAND2_23342 ( P3_SUB_598_U154 , P3_SUB_598_U109 , P3_SUB_598_U82 );
nand NAND2_23343 ( P3_SUB_598_U155 , P3_IR_REG_1_ , P3_SUB_598_U85 );
nand NAND2_23344 ( P3_SUB_598_U156 , P3_IR_REG_0_ , P3_SUB_598_U84 );
nand NAND2_23345 ( P3_SUB_598_U157 , P3_IR_REG_17_ , P3_SUB_598_U34 );
nand NAND2_23346 ( P3_SUB_598_U158 , P3_SUB_598_U106 , P3_SUB_598_U86 );
nand NAND2_23347 ( P3_SUB_598_U159 , P3_IR_REG_13_ , P3_SUB_598_U46 );
nand NAND2_23348 ( P3_SUB_598_U160 , P3_SUB_598_U103 , P3_SUB_598_U88 );
and AND2_23349 ( P3_R693_U6 , P3_R693_U113 , P3_R693_U114 );
and AND2_23350 ( P3_R693_U7 , P3_R693_U115 , P3_R693_U116 );
and AND4_23351 ( P3_R693_U8 , P3_R693_U80 , P3_R693_U118 , P3_R693_U120 , P3_R693_U7 );
and AND2_23352 ( P3_R693_U9 , P3_R693_U126 , P3_R693_U125 );
and AND2_23353 ( P3_R693_U10 , P3_R693_U130 , P3_R693_U131 );
and AND2_23354 ( P3_R693_U11 , P3_R693_U84 , P3_R693_U10 );
and AND2_23355 ( P3_R693_U12 , P3_R693_U142 , P3_R693_U141 );
and AND3_23356 ( P3_R693_U13 , P3_R693_U178 , P3_R693_U179 , P3_R693_U177 );
and AND4_23357 ( P3_R693_U14 , P3_R693_U189 , P3_R693_U188 , P3_R693_U108 , P3_R693_U109 );
not NOT1_23358 ( P3_R693_U15 , P3_U3529 );
not NOT1_23359 ( P3_R693_U16 , P3_U3537 );
not NOT1_23360 ( P3_R693_U17 , P3_U3536 );
not NOT1_23361 ( P3_R693_U18 , P3_U3905 );
not NOT1_23362 ( P3_R693_U19 , P3_U3540 );
not NOT1_23363 ( P3_R693_U20 , P3_U3906 );
not NOT1_23364 ( P3_R693_U21 , P3_U3541 );
not NOT1_23365 ( P3_R693_U22 , P3_U3543 );
not NOT1_23366 ( P3_R693_U23 , P3_U3443 );
not NOT1_23367 ( P3_R693_U24 , P3_U3544 );
not NOT1_23368 ( P3_R693_U25 , P3_U3440 );
not NOT1_23369 ( P3_R693_U26 , P3_U3445 );
not NOT1_23370 ( P3_R693_U27 , P3_U3907 );
not NOT1_23371 ( P3_R693_U28 , P3_U3545 );
not NOT1_23372 ( P3_R693_U29 , P3_U3546 );
not NOT1_23373 ( P3_R693_U30 , P3_U3437 );
not NOT1_23374 ( P3_R693_U31 , P3_U3434 );
not NOT1_23375 ( P3_R693_U32 , P3_U3526 );
not NOT1_23376 ( P3_R693_U33 , P3_U3525 );
not NOT1_23377 ( P3_R693_U34 , P3_U3404 );
not NOT1_23378 ( P3_R693_U35 , P3_U3407 );
not NOT1_23379 ( P3_R693_U36 , P3_U3416 );
not NOT1_23380 ( P3_R693_U37 , P3_U3419 );
not NOT1_23381 ( P3_R693_U38 , P3_U3410 );
not NOT1_23382 ( P3_R693_U39 , P3_U3413 );
not NOT1_23383 ( P3_R693_U40 , P3_U3398 );
not NOT1_23384 ( P3_R693_U41 , P3_U3401 );
not NOT1_23385 ( P3_R693_U42 , P3_U3553 );
not NOT1_23386 ( P3_R693_U43 , P3_U3395 );
not NOT1_23387 ( P3_R693_U44 , P3_U3392 );
not NOT1_23388 ( P3_R693_U45 , P3_U3550 );
not NOT1_23389 ( P3_R693_U46 , P3_U3549 );
not NOT1_23390 ( P3_R693_U47 , P3_U3542 );
not NOT1_23391 ( P3_R693_U48 , P3_U3531 );
not NOT1_23392 ( P3_R693_U49 , P3_U3528 );
not NOT1_23393 ( P3_R693_U50 , P3_U3527 );
not NOT1_23394 ( P3_R693_U51 , P3_U3523 );
not NOT1_23395 ( P3_R693_U52 , P3_U3524 );
not NOT1_23396 ( P3_R693_U53 , P3_U3552 );
not NOT1_23397 ( P3_R693_U54 , P3_U3551 );
not NOT1_23398 ( P3_R693_U55 , P3_U3425 );
not NOT1_23399 ( P3_R693_U56 , P3_U3422 );
not NOT1_23400 ( P3_R693_U57 , P3_U3431 );
not NOT1_23401 ( P3_R693_U58 , P3_U3428 );
not NOT1_23402 ( P3_R693_U59 , P3_U3548 );
not NOT1_23403 ( P3_R693_U60 , P3_U3547 );
not NOT1_23404 ( P3_R693_U61 , P3_U3539 );
not NOT1_23405 ( P3_R693_U62 , P3_U3538 );
not NOT1_23406 ( P3_R693_U63 , P3_U3908 );
not NOT1_23407 ( P3_R693_U64 , P3_U3900 );
not NOT1_23408 ( P3_R693_U65 , P3_U3899 );
not NOT1_23409 ( P3_R693_U66 , P3_U3904 );
not NOT1_23410 ( P3_R693_U67 , P3_U3903 );
not NOT1_23411 ( P3_R693_U68 , P3_U3902 );
not NOT1_23412 ( P3_R693_U69 , P3_U3901 );
not NOT1_23413 ( P3_R693_U70 , P3_U3533 );
not NOT1_23414 ( P3_R693_U71 , P3_U3534 );
not NOT1_23415 ( P3_R693_U72 , P3_U3872 );
not NOT1_23416 ( P3_R693_U73 , P3_U3532 );
not NOT1_23417 ( P3_R693_U74 , P3_U3535 );
and AND2_23418 ( P3_R693_U75 , P3_U3540 , P3_R693_U20 );
and AND2_23419 ( P3_R693_U76 , P3_U3541 , P3_R693_U27 );
and AND2_23420 ( P3_R693_U77 , P3_R693_U168 , P3_R693_U167 );
and AND2_23421 ( P3_R693_U78 , P3_U3443 , P3_R693_U24 );
and AND2_23422 ( P3_R693_U79 , P3_U3440 , P3_R693_U28 );
and AND2_23423 ( P3_R693_U80 , P3_R693_U119 , P3_R693_U117 );
and AND2_23424 ( P3_R693_U81 , P3_U3404 , P3_R693_U50 );
and AND2_23425 ( P3_R693_U82 , P3_U3407 , P3_R693_U32 );
and AND2_23426 ( P3_R693_U83 , P3_U3387 , P3_R693_U111 );
and AND2_23427 ( P3_R693_U84 , P3_R693_U133 , P3_R693_U132 );
and AND2_23428 ( P3_R693_U85 , P3_R693_U129 , P3_R693_U86 );
and AND2_23429 ( P3_R693_U86 , P3_R693_U135 , P3_R693_U134 );
and AND2_23430 ( P3_R693_U87 , P3_R693_U138 , P3_R693_U137 );
and AND2_23431 ( P3_R693_U88 , P3_R693_U135 , P3_R693_U134 );
and AND2_23432 ( P3_R693_U89 , P3_R693_U9 , P3_R693_U148 );
and AND3_23433 ( P3_R693_U90 , P3_R693_U129 , P3_R693_U127 , P3_R693_U11 );
and AND2_23434 ( P3_R693_U91 , P3_U3523 , P3_R693_U36 );
and AND2_23435 ( P3_R693_U92 , P3_U3524 , P3_R693_U39 );
and AND3_23436 ( P3_R693_U93 , P3_R693_U152 , P3_R693_U151 , P3_R693_U95 );
and AND2_23437 ( P3_R693_U94 , P3_R693_U154 , P3_R693_U153 );
and AND2_23438 ( P3_R693_U95 , P3_R693_U94 , P3_R693_U12 );
and AND2_23439 ( P3_R693_U96 , P3_U3425 , P3_R693_U45 );
and AND2_23440 ( P3_R693_U97 , P3_U3422 , P3_R693_U54 );
and AND2_23441 ( P3_R693_U98 , P3_R693_U157 , P3_R693_U100 );
and AND2_23442 ( P3_R693_U99 , P3_R693_U98 , P3_R693_U158 );
and AND2_23443 ( P3_R693_U100 , P3_R693_U160 , P3_R693_U159 );
and AND4_23444 ( P3_R693_U101 , P3_R693_U171 , P3_R693_U170 , P3_R693_U122 , P3_R693_U123 );
and AND2_23445 ( P3_R693_U102 , P3_R693_U175 , P3_R693_U174 );
and AND2_23446 ( P3_R693_U103 , P3_R693_U187 , P3_R693_U186 );
and AND2_23447 ( P3_R693_U104 , P3_R693_U103 , P3_R693_U13 );
and AND2_23448 ( P3_R693_U105 , P3_R693_U106 , P3_R693_U190 );
and AND2_23449 ( P3_R693_U106 , P3_U3533 , P3_R693_U65 );
and AND2_23450 ( P3_R693_U107 , P3_U3532 , P3_R693_U63 );
and AND2_23451 ( P3_R693_U108 , P3_R693_U192 , P3_R693_U191 );
and AND3_23452 ( P3_R693_U109 , P3_R693_U194 , P3_R693_U193 , P3_R693_U195 );
not NOT1_23453 ( P3_R693_U110 , P3_U3873 );
not NOT1_23454 ( P3_R693_U111 , P3_U3554 );
nand NAND2_23455 ( P3_R693_U112 , P3_R693_U181 , P3_R693_U196 );
nand NAND2_23456 ( P3_R693_U113 , P3_U3543 , P3_R693_U26 );
nand NAND2_23457 ( P3_R693_U114 , P3_U3544 , P3_R693_U23 );
nand NAND2_23458 ( P3_R693_U115 , P3_U3905 , P3_R693_U61 );
nand NAND2_23459 ( P3_R693_U116 , P3_U3906 , P3_R693_U19 );
nand NAND2_23460 ( P3_R693_U117 , P3_R693_U78 , P3_R693_U113 );
nand NAND2_23461 ( P3_R693_U118 , P3_R693_U79 , P3_R693_U6 );
nand NAND2_23462 ( P3_R693_U119 , P3_U3445 , P3_R693_U22 );
nand NAND2_23463 ( P3_R693_U120 , P3_U3907 , P3_R693_U21 );
nand NAND2_23464 ( P3_R693_U121 , P3_U3437 , P3_R693_U29 );
nand NAND2_23465 ( P3_R693_U122 , P3_U3537 , P3_R693_U67 );
nand NAND2_23466 ( P3_R693_U123 , P3_U3536 , P3_R693_U68 );
nand NAND2_23467 ( P3_R693_U124 , P3_U3434 , P3_R693_U60 );
nand NAND2_23468 ( P3_R693_U125 , P3_U3526 , P3_R693_U35 );
nand NAND2_23469 ( P3_R693_U126 , P3_U3525 , P3_R693_U38 );
nand NAND2_23470 ( P3_R693_U127 , P3_R693_U81 , P3_R693_U9 );
nand NAND2_23471 ( P3_R693_U128 , P3_U3525 , P3_R693_U38 );
nand NAND2_23472 ( P3_R693_U129 , P3_R693_U82 , P3_R693_U128 );
nand NAND2_23473 ( P3_R693_U130 , P3_U3419 , P3_R693_U53 );
nand NAND2_23474 ( P3_R693_U131 , P3_U3416 , P3_R693_U51 );
nand NAND2_23475 ( P3_R693_U132 , P3_U3410 , P3_R693_U33 );
nand NAND2_23476 ( P3_R693_U133 , P3_U3413 , P3_R693_U52 );
nand NAND2_23477 ( P3_R693_U134 , P3_U3398 , P3_R693_U48 );
nand NAND2_23478 ( P3_R693_U135 , P3_U3401 , P3_R693_U49 );
nand NAND2_23479 ( P3_R693_U136 , P3_U3553 , P3_R693_U44 );
nand NAND2_23480 ( P3_R693_U137 , P3_R693_U83 , P3_R693_U136 );
nand NAND2_23481 ( P3_R693_U138 , P3_U3395 , P3_R693_U47 );
nand NAND2_23482 ( P3_R693_U139 , P3_U3392 , P3_R693_U42 );
nand NAND5_23483 ( P3_R693_U140 , P3_R693_U11 , P3_R693_U139 , P3_R693_U87 , P3_R693_U127 , P3_R693_U85 );
nand NAND2_23484 ( P3_R693_U141 , P3_U3550 , P3_R693_U55 );
nand NAND2_23485 ( P3_R693_U142 , P3_U3549 , P3_R693_U58 );
nand NAND2_23486 ( P3_R693_U143 , P3_U3542 , P3_R693_U43 );
nand NAND2_23487 ( P3_R693_U144 , P3_U3531 , P3_R693_U40 );
nand NAND2_23488 ( P3_R693_U145 , P3_R693_U144 , P3_R693_U143 );
nand NAND2_23489 ( P3_R693_U146 , P3_R693_U88 , P3_R693_U145 );
nand NAND2_23490 ( P3_R693_U147 , P3_U3528 , P3_R693_U41 );
nand NAND2_23491 ( P3_R693_U148 , P3_U3527 , P3_R693_U34 );
nand NAND3_23492 ( P3_R693_U149 , P3_R693_U147 , P3_R693_U146 , P3_R693_U89 );
nand NAND2_23493 ( P3_R693_U150 , P3_R693_U90 , P3_R693_U149 );
nand NAND2_23494 ( P3_R693_U151 , P3_R693_U91 , P3_R693_U130 );
nand NAND2_23495 ( P3_R693_U152 , P3_R693_U92 , P3_R693_U10 );
nand NAND2_23496 ( P3_R693_U153 , P3_U3552 , P3_R693_U37 );
nand NAND2_23497 ( P3_R693_U154 , P3_U3551 , P3_R693_U56 );
nand NAND3_23498 ( P3_R693_U155 , P3_R693_U150 , P3_R693_U140 , P3_R693_U93 );
nand NAND2_23499 ( P3_R693_U156 , P3_U3549 , P3_R693_U58 );
nand NAND2_23500 ( P3_R693_U157 , P3_R693_U96 , P3_R693_U156 );
nand NAND2_23501 ( P3_R693_U158 , P3_R693_U97 , P3_R693_U12 );
nand NAND2_23502 ( P3_R693_U159 , P3_U3431 , P3_R693_U59 );
nand NAND2_23503 ( P3_R693_U160 , P3_U3428 , P3_R693_U46 );
nand NAND2_23504 ( P3_R693_U161 , P3_R693_U155 , P3_R693_U99 );
nand NAND2_23505 ( P3_R693_U162 , P3_U3548 , P3_R693_U57 );
nand NAND2_23506 ( P3_R693_U163 , P3_R693_U162 , P3_R693_U161 );
nand NAND2_23507 ( P3_R693_U164 , P3_R693_U163 , P3_R693_U124 );
nand NAND2_23508 ( P3_R693_U165 , P3_U3547 , P3_R693_U31 );
nand NAND2_23509 ( P3_R693_U166 , P3_R693_U165 , P3_R693_U164 );
nand NAND2_23510 ( P3_R693_U167 , P3_U3545 , P3_R693_U25 );
nand NAND2_23511 ( P3_R693_U168 , P3_U3546 , P3_R693_U30 );
nand NAND2_23512 ( P3_R693_U169 , P3_R693_U77 , P3_R693_U6 );
nand NAND2_23513 ( P3_R693_U170 , P3_R693_U75 , P3_R693_U115 );
nand NAND2_23514 ( P3_R693_U171 , P3_R693_U76 , P3_R693_U7 );
nand NAND2_23515 ( P3_R693_U172 , P3_R693_U8 , P3_R693_U169 );
nand NAND3_23516 ( P3_R693_U173 , P3_R693_U166 , P3_R693_U121 , P3_R693_U8 );
nand NAND2_23517 ( P3_R693_U174 , P3_U3539 , P3_R693_U18 );
nand NAND2_23518 ( P3_R693_U175 , P3_U3538 , P3_R693_U66 );
nand NAND4_23519 ( P3_R693_U176 , P3_R693_U173 , P3_R693_U172 , P3_R693_U102 , P3_R693_U101 );
nand NAND2_23520 ( P3_R693_U177 , P3_U3908 , P3_R693_U73 );
nand NAND2_23521 ( P3_R693_U178 , P3_U3900 , P3_R693_U71 );
nand NAND2_23522 ( P3_R693_U179 , P3_U3899 , P3_R693_U70 );
nand NAND2_23523 ( P3_R693_U180 , P3_U3529 , P3_R693_U72 );
nand NAND2_23524 ( P3_R693_U181 , P3_R693_U180 , P3_R693_U110 );
nand NAND2_23525 ( P3_R693_U182 , P3_U3904 , P3_R693_U62 );
nand NAND2_23526 ( P3_R693_U183 , P3_U3903 , P3_R693_U16 );
nand NAND2_23527 ( P3_R693_U184 , P3_R693_U183 , P3_R693_U182 );
nand NAND3_23528 ( P3_R693_U185 , P3_R693_U184 , P3_R693_U122 , P3_R693_U123 );
nand NAND2_23529 ( P3_R693_U186 , P3_U3902 , P3_R693_U17 );
nand NAND2_23530 ( P3_R693_U187 , P3_U3901 , P3_R693_U74 );
nand NAND4_23531 ( P3_R693_U188 , P3_R693_U176 , P3_R693_U185 , P3_R693_U112 , P3_R693_U104 );
nand NAND3_23532 ( P3_R693_U189 , P3_R693_U180 , P3_U3530 , P3_R693_U110 );
nand NAND2_23533 ( P3_R693_U190 , P3_U3908 , P3_R693_U73 );
nand NAND2_23534 ( P3_R693_U191 , P3_R693_U112 , P3_R693_U105 );
nand NAND4_23535 ( P3_R693_U192 , P3_U3534 , P3_R693_U13 , P3_R693_U112 , P3_R693_U64 );
nand NAND2_23536 ( P3_R693_U193 , P3_U3872 , P3_R693_U15 );
nand NAND2_23537 ( P3_R693_U194 , P3_R693_U107 , P3_R693_U112 );
nand NAND4_23538 ( P3_R693_U195 , P3_U3535 , P3_R693_U13 , P3_R693_U112 , P3_R693_U69 );
nand NAND2_23539 ( P3_R693_U196 , P3_U3530 , P3_R693_U180 );
nand NAND2_23540 ( P3_SUB_609_U6 , P3_SUB_609_U40 , P3_SUB_609_U98 );
nand NAND2_23541 ( P3_SUB_609_U7 , P3_SUB_609_U79 , P3_SUB_609_U105 );
nand NAND2_23542 ( P3_SUB_609_U8 , P3_SUB_609_U65 , P3_SUB_609_U113 );
nand NAND2_23543 ( P3_SUB_609_U9 , P3_SUB_609_U34 , P3_SUB_609_U110 );
nand NAND2_23544 ( P3_SUB_609_U10 , P3_SUB_609_U87 , P3_SUB_609_U97 );
nand NAND2_23545 ( P3_SUB_609_U11 , P3_SUB_609_U81 , P3_SUB_609_U103 );
nand NAND2_23546 ( P3_SUB_609_U12 , P3_SUB_609_U67 , P3_SUB_609_U70 );
nand NAND2_23547 ( P3_SUB_609_U13 , P3_SUB_609_U73 , P3_SUB_609_U111 );
nand NAND2_23548 ( P3_SUB_609_U14 , P3_SUB_609_U33 , P3_SUB_609_U69 );
nand NAND2_23549 ( P3_SUB_609_U15 , P3_SUB_609_U38 , P3_SUB_609_U102 );
nand NAND2_23550 ( P3_SUB_609_U16 , P3_SUB_609_U41 , P3_SUB_609_U96 );
nand NAND2_23551 ( P3_SUB_609_U17 , P3_SUB_609_U85 , P3_SUB_609_U99 );
nand NAND2_23552 ( P3_SUB_609_U18 , P3_SUB_609_U31 , P3_SUB_609_U71 );
nand NAND2_23553 ( P3_SUB_609_U19 , P3_SUB_609_U37 , P3_SUB_609_U104 );
nand NAND2_23554 ( P3_SUB_609_U20 , P3_SUB_609_U83 , P3_SUB_609_U101 );
nand NAND2_23555 ( P3_SUB_609_U21 , P3_SUB_609_U36 , P3_SUB_609_U106 );
nand NAND2_23556 ( P3_SUB_609_U22 , P3_SUB_609_U42 , P3_SUB_609_U94 );
nand NAND2_23557 ( P3_SUB_609_U23 , P3_SUB_609_U75 , P3_SUB_609_U109 );
nand NAND2_23558 ( P3_SUB_609_U24 , P3_SUB_609_U35 , P3_SUB_609_U108 );
not NOT1_23559 ( P3_SUB_609_U25 , P3_REG3_REG_3_ );
nand NAND2_23560 ( P3_SUB_609_U26 , P3_SUB_609_U89 , P3_SUB_609_U95 );
nand NAND2_23561 ( P3_SUB_609_U27 , P3_SUB_609_U39 , P3_SUB_609_U100 );
nand NAND2_23562 ( P3_SUB_609_U28 , P3_SUB_609_U91 , P3_SUB_609_U93 );
nand NAND2_23563 ( P3_SUB_609_U29 , P3_SUB_609_U64 , P3_SUB_609_U72 );
nand NAND2_23564 ( P3_SUB_609_U30 , P3_SUB_609_U77 , P3_SUB_609_U107 );
or OR5_23565 ( P3_SUB_609_U31 , P3_REG3_REG_4_ , P3_REG3_REG_3_ , P3_REG3_REG_5_ , P3_REG3_REG_6_ , P3_REG3_REG_7_ );
not NOT1_23566 ( P3_SUB_609_U32 , P3_REG3_REG_8_ );
nand NAND2_23567 ( P3_SUB_609_U33 , P3_SUB_609_U54 , P3_SUB_609_U66 );
nand NAND2_23568 ( P3_SUB_609_U34 , P3_SUB_609_U55 , P3_SUB_609_U68 );
nand NAND2_23569 ( P3_SUB_609_U35 , P3_SUB_609_U56 , P3_SUB_609_U74 );
nand NAND2_23570 ( P3_SUB_609_U36 , P3_SUB_609_U57 , P3_SUB_609_U76 );
nand NAND2_23571 ( P3_SUB_609_U37 , P3_SUB_609_U58 , P3_SUB_609_U78 );
nand NAND2_23572 ( P3_SUB_609_U38 , P3_SUB_609_U59 , P3_SUB_609_U80 );
nand NAND2_23573 ( P3_SUB_609_U39 , P3_SUB_609_U60 , P3_SUB_609_U82 );
nand NAND2_23574 ( P3_SUB_609_U40 , P3_SUB_609_U61 , P3_SUB_609_U84 );
nand NAND2_23575 ( P3_SUB_609_U41 , P3_SUB_609_U62 , P3_SUB_609_U86 );
nand NAND2_23576 ( P3_SUB_609_U42 , P3_SUB_609_U63 , P3_SUB_609_U88 );
not NOT1_23577 ( P3_SUB_609_U43 , P3_REG3_REG_28_ );
not NOT1_23578 ( P3_SUB_609_U44 , P3_REG3_REG_26_ );
not NOT1_23579 ( P3_SUB_609_U45 , P3_REG3_REG_24_ );
not NOT1_23580 ( P3_SUB_609_U46 , P3_REG3_REG_22_ );
not NOT1_23581 ( P3_SUB_609_U47 , P3_REG3_REG_20_ );
not NOT1_23582 ( P3_SUB_609_U48 , P3_REG3_REG_18_ );
not NOT1_23583 ( P3_SUB_609_U49 , P3_REG3_REG_16_ );
not NOT1_23584 ( P3_SUB_609_U50 , P3_REG3_REG_14_ );
not NOT1_23585 ( P3_SUB_609_U51 , P3_REG3_REG_12_ );
not NOT1_23586 ( P3_SUB_609_U52 , P3_REG3_REG_10_ );
nand NAND2_23587 ( P3_SUB_609_U53 , P3_SUB_609_U115 , P3_SUB_609_U114 );
nor nor_23588 ( P3_SUB_609_U54 , P3_REG3_REG_8_ , P3_REG3_REG_9_ );
nor nor_23589 ( P3_SUB_609_U55 , P3_REG3_REG_10_ , P3_REG3_REG_11_ );
nor nor_23590 ( P3_SUB_609_U56 , P3_REG3_REG_12_ , P3_REG3_REG_13_ );
nor nor_23591 ( P3_SUB_609_U57 , P3_REG3_REG_14_ , P3_REG3_REG_15_ );
nor nor_23592 ( P3_SUB_609_U58 , P3_REG3_REG_16_ , P3_REG3_REG_17_ );
nor nor_23593 ( P3_SUB_609_U59 , P3_REG3_REG_18_ , P3_REG3_REG_19_ );
nor nor_23594 ( P3_SUB_609_U60 , P3_REG3_REG_20_ , P3_REG3_REG_21_ );
nor nor_23595 ( P3_SUB_609_U61 , P3_REG3_REG_22_ , P3_REG3_REG_23_ );
nor nor_23596 ( P3_SUB_609_U62 , P3_REG3_REG_24_ , P3_REG3_REG_25_ );
nor nor_23597 ( P3_SUB_609_U63 , P3_REG3_REG_26_ , P3_REG3_REG_27_ );
or OR2_23598 ( P3_SUB_609_U64 , P3_REG3_REG_3_ , P3_REG3_REG_4_ );
or OR4_23599 ( P3_SUB_609_U65 , P3_REG3_REG_5_ , P3_REG3_REG_6_ , P3_REG3_REG_4_ , P3_REG3_REG_3_ );
not NOT1_23600 ( P3_SUB_609_U66 , P3_SUB_609_U31 );
nand NAND2_23601 ( P3_SUB_609_U67 , P3_SUB_609_U66 , P3_SUB_609_U32 );
not NOT1_23602 ( P3_SUB_609_U68 , P3_SUB_609_U33 );
nand NAND2_23603 ( P3_SUB_609_U69 , P3_REG3_REG_9_ , P3_SUB_609_U67 );
nand NAND2_23604 ( P3_SUB_609_U70 , P3_REG3_REG_8_ , P3_SUB_609_U31 );
nand NAND2_23605 ( P3_SUB_609_U71 , P3_REG3_REG_7_ , P3_SUB_609_U65 );
nand NAND2_23606 ( P3_SUB_609_U72 , P3_REG3_REG_4_ , P3_REG3_REG_3_ );
nand NAND2_23607 ( P3_SUB_609_U73 , P3_SUB_609_U68 , P3_SUB_609_U52 );
not NOT1_23608 ( P3_SUB_609_U74 , P3_SUB_609_U34 );
nand NAND2_23609 ( P3_SUB_609_U75 , P3_SUB_609_U74 , P3_SUB_609_U51 );
not NOT1_23610 ( P3_SUB_609_U76 , P3_SUB_609_U35 );
nand NAND2_23611 ( P3_SUB_609_U77 , P3_SUB_609_U76 , P3_SUB_609_U50 );
not NOT1_23612 ( P3_SUB_609_U78 , P3_SUB_609_U36 );
nand NAND2_23613 ( P3_SUB_609_U79 , P3_SUB_609_U78 , P3_SUB_609_U49 );
not NOT1_23614 ( P3_SUB_609_U80 , P3_SUB_609_U37 );
nand NAND2_23615 ( P3_SUB_609_U81 , P3_SUB_609_U80 , P3_SUB_609_U48 );
not NOT1_23616 ( P3_SUB_609_U82 , P3_SUB_609_U38 );
nand NAND2_23617 ( P3_SUB_609_U83 , P3_SUB_609_U82 , P3_SUB_609_U47 );
not NOT1_23618 ( P3_SUB_609_U84 , P3_SUB_609_U39 );
nand NAND2_23619 ( P3_SUB_609_U85 , P3_SUB_609_U84 , P3_SUB_609_U46 );
not NOT1_23620 ( P3_SUB_609_U86 , P3_SUB_609_U40 );
nand NAND2_23621 ( P3_SUB_609_U87 , P3_SUB_609_U86 , P3_SUB_609_U45 );
not NOT1_23622 ( P3_SUB_609_U88 , P3_SUB_609_U41 );
nand NAND2_23623 ( P3_SUB_609_U89 , P3_SUB_609_U88 , P3_SUB_609_U44 );
not NOT1_23624 ( P3_SUB_609_U90 , P3_SUB_609_U42 );
nand NAND2_23625 ( P3_SUB_609_U91 , P3_SUB_609_U90 , P3_SUB_609_U43 );
not NOT1_23626 ( P3_SUB_609_U92 , P3_SUB_609_U91 );
nand NAND2_23627 ( P3_SUB_609_U93 , P3_REG3_REG_28_ , P3_SUB_609_U42 );
nand NAND2_23628 ( P3_SUB_609_U94 , P3_REG3_REG_27_ , P3_SUB_609_U89 );
nand NAND2_23629 ( P3_SUB_609_U95 , P3_REG3_REG_26_ , P3_SUB_609_U41 );
nand NAND2_23630 ( P3_SUB_609_U96 , P3_REG3_REG_25_ , P3_SUB_609_U87 );
nand NAND2_23631 ( P3_SUB_609_U97 , P3_REG3_REG_24_ , P3_SUB_609_U40 );
nand NAND2_23632 ( P3_SUB_609_U98 , P3_REG3_REG_23_ , P3_SUB_609_U85 );
nand NAND2_23633 ( P3_SUB_609_U99 , P3_REG3_REG_22_ , P3_SUB_609_U39 );
nand NAND2_23634 ( P3_SUB_609_U100 , P3_REG3_REG_21_ , P3_SUB_609_U83 );
nand NAND2_23635 ( P3_SUB_609_U101 , P3_REG3_REG_20_ , P3_SUB_609_U38 );
nand NAND2_23636 ( P3_SUB_609_U102 , P3_REG3_REG_19_ , P3_SUB_609_U81 );
nand NAND2_23637 ( P3_SUB_609_U103 , P3_REG3_REG_18_ , P3_SUB_609_U37 );
nand NAND2_23638 ( P3_SUB_609_U104 , P3_REG3_REG_17_ , P3_SUB_609_U79 );
nand NAND2_23639 ( P3_SUB_609_U105 , P3_REG3_REG_16_ , P3_SUB_609_U36 );
nand NAND2_23640 ( P3_SUB_609_U106 , P3_REG3_REG_15_ , P3_SUB_609_U77 );
nand NAND2_23641 ( P3_SUB_609_U107 , P3_REG3_REG_14_ , P3_SUB_609_U35 );
nand NAND2_23642 ( P3_SUB_609_U108 , P3_REG3_REG_13_ , P3_SUB_609_U75 );
nand NAND2_23643 ( P3_SUB_609_U109 , P3_REG3_REG_12_ , P3_SUB_609_U34 );
nand NAND2_23644 ( P3_SUB_609_U110 , P3_REG3_REG_11_ , P3_SUB_609_U73 );
nand NAND2_23645 ( P3_SUB_609_U111 , P3_REG3_REG_10_ , P3_SUB_609_U33 );
or OR3_23646 ( P3_SUB_609_U112 , P3_REG3_REG_4_ , P3_REG3_REG_3_ , P3_REG3_REG_5_ );
nand NAND2_23647 ( P3_SUB_609_U113 , P3_REG3_REG_6_ , P3_SUB_609_U112 );
nand NAND2_23648 ( P3_SUB_609_U114 , P3_REG3_REG_5_ , P3_SUB_609_U64 );
or OR3_23649 ( P3_SUB_609_U115 , P3_REG3_REG_4_ , P3_REG3_REG_3_ , P3_REG3_REG_5_ );
and AND2_23650 ( P3_R1095_U6 , P3_R1095_U210 , P3_R1095_U209 );
and AND2_23651 ( P3_R1095_U7 , P3_R1095_U189 , P3_R1095_U245 );
and AND2_23652 ( P3_R1095_U8 , P3_R1095_U247 , P3_R1095_U246 );
and AND2_23653 ( P3_R1095_U9 , P3_R1095_U190 , P3_R1095_U262 );
and AND2_23654 ( P3_R1095_U10 , P3_R1095_U264 , P3_R1095_U263 );
and AND2_23655 ( P3_R1095_U11 , P3_R1095_U191 , P3_R1095_U286 );
and AND2_23656 ( P3_R1095_U12 , P3_R1095_U288 , P3_R1095_U287 );
and AND3_23657 ( P3_R1095_U13 , P3_R1095_U208 , P3_R1095_U194 , P3_R1095_U213 );
and AND2_23658 ( P3_R1095_U14 , P3_R1095_U218 , P3_R1095_U195 );
and AND2_23659 ( P3_R1095_U15 , P3_R1095_U392 , P3_R1095_U391 );
nand NAND2_23660 ( P3_R1095_U16 , P3_R1095_U342 , P3_R1095_U345 );
nand NAND2_23661 ( P3_R1095_U17 , P3_R1095_U331 , P3_R1095_U334 );
nand NAND2_23662 ( P3_R1095_U18 , P3_R1095_U320 , P3_R1095_U323 );
nand NAND2_23663 ( P3_R1095_U19 , P3_R1095_U312 , P3_R1095_U314 );
nand NAND3_23664 ( P3_R1095_U20 , P3_R1095_U162 , P3_R1095_U183 , P3_R1095_U351 );
nand NAND2_23665 ( P3_R1095_U21 , P3_R1095_U241 , P3_R1095_U243 );
nand NAND2_23666 ( P3_R1095_U22 , P3_R1095_U233 , P3_R1095_U236 );
nand NAND2_23667 ( P3_R1095_U23 , P3_R1095_U225 , P3_R1095_U227 );
nand NAND2_23668 ( P3_R1095_U24 , P3_R1095_U172 , P3_R1095_U348 );
not NOT1_23669 ( P3_R1095_U25 , P3_U3069 );
nand NAND2_23670 ( P3_R1095_U26 , P3_U3069 , P3_R1095_U39 );
not NOT1_23671 ( P3_R1095_U27 , P3_U3083 );
not NOT1_23672 ( P3_R1095_U28 , P3_U3413 );
not NOT1_23673 ( P3_R1095_U29 , P3_U3395 );
not NOT1_23674 ( P3_R1095_U30 , P3_U3387 );
not NOT1_23675 ( P3_R1095_U31 , P3_U3077 );
not NOT1_23676 ( P3_R1095_U32 , P3_U3398 );
not NOT1_23677 ( P3_R1095_U33 , P3_U3067 );
nand NAND2_23678 ( P3_R1095_U34 , P3_U3067 , P3_R1095_U29 );
not NOT1_23679 ( P3_R1095_U35 , P3_U3063 );
not NOT1_23680 ( P3_R1095_U36 , P3_U3404 );
not NOT1_23681 ( P3_R1095_U37 , P3_U3407 );
not NOT1_23682 ( P3_R1095_U38 , P3_U3401 );
not NOT1_23683 ( P3_R1095_U39 , P3_U3410 );
not NOT1_23684 ( P3_R1095_U40 , P3_U3070 );
not NOT1_23685 ( P3_R1095_U41 , P3_U3066 );
not NOT1_23686 ( P3_R1095_U42 , P3_U3059 );
nand NAND2_23687 ( P3_R1095_U43 , P3_U3059 , P3_R1095_U38 );
nand NAND2_23688 ( P3_R1095_U44 , P3_R1095_U214 , P3_R1095_U212 );
not NOT1_23689 ( P3_R1095_U45 , P3_U3416 );
not NOT1_23690 ( P3_R1095_U46 , P3_U3082 );
nand NAND2_23691 ( P3_R1095_U47 , P3_R1095_U44 , P3_R1095_U215 );
nand NAND2_23692 ( P3_R1095_U48 , P3_R1095_U43 , P3_R1095_U229 );
nand NAND3_23693 ( P3_R1095_U49 , P3_R1095_U201 , P3_R1095_U185 , P3_R1095_U349 );
not NOT1_23694 ( P3_R1095_U50 , P3_U3901 );
not NOT1_23695 ( P3_R1095_U51 , P3_U3422 );
not NOT1_23696 ( P3_R1095_U52 , P3_U3419 );
not NOT1_23697 ( P3_R1095_U53 , P3_U3062 );
not NOT1_23698 ( P3_R1095_U54 , P3_U3061 );
nand NAND2_23699 ( P3_R1095_U55 , P3_U3082 , P3_R1095_U45 );
not NOT1_23700 ( P3_R1095_U56 , P3_U3425 );
not NOT1_23701 ( P3_R1095_U57 , P3_U3071 );
not NOT1_23702 ( P3_R1095_U58 , P3_U3428 );
not NOT1_23703 ( P3_R1095_U59 , P3_U3079 );
not NOT1_23704 ( P3_R1095_U60 , P3_U3437 );
not NOT1_23705 ( P3_R1095_U61 , P3_U3434 );
not NOT1_23706 ( P3_R1095_U62 , P3_U3431 );
not NOT1_23707 ( P3_R1095_U63 , P3_U3072 );
not NOT1_23708 ( P3_R1095_U64 , P3_U3073 );
not NOT1_23709 ( P3_R1095_U65 , P3_U3078 );
nand NAND2_23710 ( P3_R1095_U66 , P3_U3078 , P3_R1095_U62 );
not NOT1_23711 ( P3_R1095_U67 , P3_U3440 );
not NOT1_23712 ( P3_R1095_U68 , P3_U3068 );
not NOT1_23713 ( P3_R1095_U69 , P3_U3081 );
not NOT1_23714 ( P3_R1095_U70 , P3_U3445 );
not NOT1_23715 ( P3_R1095_U71 , P3_U3080 );
not NOT1_23716 ( P3_R1095_U72 , P3_U3907 );
not NOT1_23717 ( P3_R1095_U73 , P3_U3075 );
not NOT1_23718 ( P3_R1095_U74 , P3_U3904 );
not NOT1_23719 ( P3_R1095_U75 , P3_U3905 );
not NOT1_23720 ( P3_R1095_U76 , P3_U3906 );
not NOT1_23721 ( P3_R1095_U77 , P3_U3065 );
not NOT1_23722 ( P3_R1095_U78 , P3_U3060 );
not NOT1_23723 ( P3_R1095_U79 , P3_U3074 );
nand NAND2_23724 ( P3_R1095_U80 , P3_U3074 , P3_R1095_U76 );
not NOT1_23725 ( P3_R1095_U81 , P3_U3903 );
not NOT1_23726 ( P3_R1095_U82 , P3_U3064 );
not NOT1_23727 ( P3_R1095_U83 , P3_U3902 );
not NOT1_23728 ( P3_R1095_U84 , P3_U3057 );
not NOT1_23729 ( P3_R1095_U85 , P3_U3900 );
not NOT1_23730 ( P3_R1095_U86 , P3_U3056 );
nand NAND2_23731 ( P3_R1095_U87 , P3_U3056 , P3_R1095_U50 );
not NOT1_23732 ( P3_R1095_U88 , P3_U3052 );
not NOT1_23733 ( P3_R1095_U89 , P3_U3899 );
not NOT1_23734 ( P3_R1095_U90 , P3_U3053 );
nand NAND2_23735 ( P3_R1095_U91 , P3_R1095_U302 , P3_R1095_U301 );
nand NAND2_23736 ( P3_R1095_U92 , P3_R1095_U80 , P3_R1095_U316 );
nand NAND2_23737 ( P3_R1095_U93 , P3_R1095_U66 , P3_R1095_U327 );
nand NAND2_23738 ( P3_R1095_U94 , P3_R1095_U55 , P3_R1095_U338 );
not NOT1_23739 ( P3_R1095_U95 , P3_U3076 );
nand NAND2_23740 ( P3_R1095_U96 , P3_R1095_U402 , P3_R1095_U401 );
nand NAND2_23741 ( P3_R1095_U97 , P3_R1095_U416 , P3_R1095_U415 );
nand NAND2_23742 ( P3_R1095_U98 , P3_R1095_U421 , P3_R1095_U420 );
nand NAND2_23743 ( P3_R1095_U99 , P3_R1095_U437 , P3_R1095_U436 );
nand NAND2_23744 ( P3_R1095_U100 , P3_R1095_U442 , P3_R1095_U441 );
nand NAND2_23745 ( P3_R1095_U101 , P3_R1095_U447 , P3_R1095_U446 );
nand NAND2_23746 ( P3_R1095_U102 , P3_R1095_U452 , P3_R1095_U451 );
nand NAND2_23747 ( P3_R1095_U103 , P3_R1095_U457 , P3_R1095_U456 );
nand NAND2_23748 ( P3_R1095_U104 , P3_R1095_U473 , P3_R1095_U472 );
nand NAND2_23749 ( P3_R1095_U105 , P3_R1095_U478 , P3_R1095_U477 );
nand NAND2_23750 ( P3_R1095_U106 , P3_R1095_U361 , P3_R1095_U360 );
nand NAND2_23751 ( P3_R1095_U107 , P3_R1095_U370 , P3_R1095_U369 );
nand NAND2_23752 ( P3_R1095_U108 , P3_R1095_U377 , P3_R1095_U376 );
nand NAND2_23753 ( P3_R1095_U109 , P3_R1095_U381 , P3_R1095_U380 );
nand NAND2_23754 ( P3_R1095_U110 , P3_R1095_U390 , P3_R1095_U389 );
nand NAND2_23755 ( P3_R1095_U111 , P3_R1095_U411 , P3_R1095_U410 );
nand NAND2_23756 ( P3_R1095_U112 , P3_R1095_U428 , P3_R1095_U427 );
nand NAND2_23757 ( P3_R1095_U113 , P3_R1095_U432 , P3_R1095_U431 );
nand NAND2_23758 ( P3_R1095_U114 , P3_R1095_U464 , P3_R1095_U463 );
nand NAND2_23759 ( P3_R1095_U115 , P3_R1095_U468 , P3_R1095_U467 );
nand NAND2_23760 ( P3_R1095_U116 , P3_R1095_U485 , P3_R1095_U484 );
and AND2_23761 ( P3_R1095_U117 , P3_R1095_U352 , P3_R1095_U193 );
and AND2_23762 ( P3_R1095_U118 , P3_R1095_U205 , P3_R1095_U206 );
and AND2_23763 ( P3_R1095_U119 , P3_R1095_U14 , P3_R1095_U13 );
and AND2_23764 ( P3_R1095_U120 , P3_R1095_U357 , P3_R1095_U354 );
and AND3_23765 ( P3_R1095_U121 , P3_R1095_U363 , P3_R1095_U362 , P3_R1095_U26 );
and AND2_23766 ( P3_R1095_U122 , P3_R1095_U366 , P3_R1095_U195 );
and AND2_23767 ( P3_R1095_U123 , P3_R1095_U235 , P3_R1095_U6 );
and AND2_23768 ( P3_R1095_U124 , P3_R1095_U373 , P3_R1095_U194 );
and AND3_23769 ( P3_R1095_U125 , P3_R1095_U383 , P3_R1095_U382 , P3_R1095_U34 );
and AND2_23770 ( P3_R1095_U126 , P3_R1095_U386 , P3_R1095_U193 );
and AND2_23771 ( P3_R1095_U127 , P3_R1095_U222 , P3_R1095_U7 );
and AND2_23772 ( P3_R1095_U128 , P3_R1095_U267 , P3_R1095_U9 );
and AND2_23773 ( P3_R1095_U129 , P3_R1095_U291 , P3_R1095_U11 );
and AND2_23774 ( P3_R1095_U130 , P3_R1095_U355 , P3_R1095_U192 );
and AND2_23775 ( P3_R1095_U131 , P3_R1095_U306 , P3_R1095_U307 );
and AND2_23776 ( P3_R1095_U132 , P3_R1095_U309 , P3_R1095_U395 );
and AND2_23777 ( P3_R1095_U133 , P3_R1095_U306 , P3_R1095_U307 );
and AND2_23778 ( P3_R1095_U134 , P3_R1095_U15 , P3_R1095_U310 );
nand NAND2_23779 ( P3_R1095_U135 , P3_R1095_U399 , P3_R1095_U398 );
and AND3_23780 ( P3_R1095_U136 , P3_R1095_U404 , P3_R1095_U403 , P3_R1095_U87 );
and AND2_23781 ( P3_R1095_U137 , P3_R1095_U407 , P3_R1095_U192 );
nand NAND2_23782 ( P3_R1095_U138 , P3_R1095_U413 , P3_R1095_U412 );
nand NAND2_23783 ( P3_R1095_U139 , P3_R1095_U418 , P3_R1095_U417 );
and AND2_23784 ( P3_R1095_U140 , P3_R1095_U322 , P3_R1095_U12 );
and AND2_23785 ( P3_R1095_U141 , P3_R1095_U424 , P3_R1095_U191 );
nand NAND2_23786 ( P3_R1095_U142 , P3_R1095_U434 , P3_R1095_U433 );
nand NAND2_23787 ( P3_R1095_U143 , P3_R1095_U439 , P3_R1095_U438 );
nand NAND2_23788 ( P3_R1095_U144 , P3_R1095_U444 , P3_R1095_U443 );
nand NAND2_23789 ( P3_R1095_U145 , P3_R1095_U449 , P3_R1095_U448 );
nand NAND2_23790 ( P3_R1095_U146 , P3_R1095_U454 , P3_R1095_U453 );
and AND2_23791 ( P3_R1095_U147 , P3_R1095_U333 , P3_R1095_U10 );
and AND2_23792 ( P3_R1095_U148 , P3_R1095_U460 , P3_R1095_U190 );
nand NAND2_23793 ( P3_R1095_U149 , P3_R1095_U470 , P3_R1095_U469 );
nand NAND2_23794 ( P3_R1095_U150 , P3_R1095_U475 , P3_R1095_U474 );
and AND2_23795 ( P3_R1095_U151 , P3_R1095_U344 , P3_R1095_U8 );
and AND2_23796 ( P3_R1095_U152 , P3_R1095_U481 , P3_R1095_U189 );
and AND2_23797 ( P3_R1095_U153 , P3_R1095_U359 , P3_R1095_U358 );
nand NAND2_23798 ( P3_R1095_U154 , P3_R1095_U120 , P3_R1095_U356 );
and AND2_23799 ( P3_R1095_U155 , P3_R1095_U368 , P3_R1095_U367 );
and AND2_23800 ( P3_R1095_U156 , P3_R1095_U375 , P3_R1095_U374 );
and AND2_23801 ( P3_R1095_U157 , P3_R1095_U379 , P3_R1095_U378 );
nand NAND2_23802 ( P3_R1095_U158 , P3_R1095_U118 , P3_R1095_U203 );
and AND2_23803 ( P3_R1095_U159 , P3_R1095_U388 , P3_R1095_U387 );
not NOT1_23804 ( P3_R1095_U160 , P3_U3908 );
not NOT1_23805 ( P3_R1095_U161 , P3_U3054 );
and AND2_23806 ( P3_R1095_U162 , P3_R1095_U397 , P3_R1095_U396 );
nand NAND2_23807 ( P3_R1095_U163 , P3_R1095_U131 , P3_R1095_U304 );
and AND2_23808 ( P3_R1095_U164 , P3_R1095_U409 , P3_R1095_U408 );
nand NAND2_23809 ( P3_R1095_U165 , P3_R1095_U298 , P3_R1095_U297 );
nand NAND2_23810 ( P3_R1095_U166 , P3_R1095_U294 , P3_R1095_U293 );
and AND2_23811 ( P3_R1095_U167 , P3_R1095_U426 , P3_R1095_U425 );
and AND2_23812 ( P3_R1095_U168 , P3_R1095_U430 , P3_R1095_U429 );
nand NAND2_23813 ( P3_R1095_U169 , P3_R1095_U284 , P3_R1095_U283 );
nand NAND2_23814 ( P3_R1095_U170 , P3_R1095_U280 , P3_R1095_U279 );
not NOT1_23815 ( P3_R1095_U171 , P3_U3392 );
nand NAND2_23816 ( P3_R1095_U172 , P3_U3387 , P3_R1095_U95 );
nand NAND3_23817 ( P3_R1095_U173 , P3_R1095_U276 , P3_R1095_U184 , P3_R1095_U350 );
not NOT1_23818 ( P3_R1095_U174 , P3_U3443 );
nand NAND2_23819 ( P3_R1095_U175 , P3_R1095_U274 , P3_R1095_U273 );
nand NAND2_23820 ( P3_R1095_U176 , P3_R1095_U270 , P3_R1095_U269 );
and AND2_23821 ( P3_R1095_U177 , P3_R1095_U462 , P3_R1095_U461 );
and AND2_23822 ( P3_R1095_U178 , P3_R1095_U466 , P3_R1095_U465 );
nand NAND2_23823 ( P3_R1095_U179 , P3_R1095_U260 , P3_R1095_U259 );
nand NAND2_23824 ( P3_R1095_U180 , P3_R1095_U256 , P3_R1095_U255 );
nand NAND2_23825 ( P3_R1095_U181 , P3_R1095_U252 , P3_R1095_U251 );
and AND2_23826 ( P3_R1095_U182 , P3_R1095_U483 , P3_R1095_U482 );
nand NAND2_23827 ( P3_R1095_U183 , P3_R1095_U132 , P3_R1095_U163 );
nand NAND2_23828 ( P3_R1095_U184 , P3_R1095_U175 , P3_R1095_U174 );
nand NAND2_23829 ( P3_R1095_U185 , P3_R1095_U172 , P3_R1095_U171 );
not NOT1_23830 ( P3_R1095_U186 , P3_R1095_U87 );
not NOT1_23831 ( P3_R1095_U187 , P3_R1095_U34 );
not NOT1_23832 ( P3_R1095_U188 , P3_R1095_U26 );
nand NAND2_23833 ( P3_R1095_U189 , P3_U3419 , P3_R1095_U54 );
nand NAND2_23834 ( P3_R1095_U190 , P3_U3434 , P3_R1095_U64 );
nand NAND2_23835 ( P3_R1095_U191 , P3_U3905 , P3_R1095_U78 );
nand NAND2_23836 ( P3_R1095_U192 , P3_U3901 , P3_R1095_U86 );
nand NAND2_23837 ( P3_R1095_U193 , P3_U3395 , P3_R1095_U33 );
nand NAND2_23838 ( P3_R1095_U194 , P3_U3404 , P3_R1095_U41 );
nand NAND2_23839 ( P3_R1095_U195 , P3_U3410 , P3_R1095_U25 );
not NOT1_23840 ( P3_R1095_U196 , P3_R1095_U66 );
not NOT1_23841 ( P3_R1095_U197 , P3_R1095_U80 );
not NOT1_23842 ( P3_R1095_U198 , P3_R1095_U43 );
not NOT1_23843 ( P3_R1095_U199 , P3_R1095_U55 );
not NOT1_23844 ( P3_R1095_U200 , P3_R1095_U172 );
nand NAND2_23845 ( P3_R1095_U201 , P3_U3077 , P3_R1095_U172 );
not NOT1_23846 ( P3_R1095_U202 , P3_R1095_U49 );
nand NAND2_23847 ( P3_R1095_U203 , P3_R1095_U117 , P3_R1095_U49 );
nand NAND2_23848 ( P3_R1095_U204 , P3_R1095_U35 , P3_R1095_U34 );
nand NAND2_23849 ( P3_R1095_U205 , P3_R1095_U204 , P3_R1095_U32 );
nand NAND2_23850 ( P3_R1095_U206 , P3_U3063 , P3_R1095_U187 );
not NOT1_23851 ( P3_R1095_U207 , P3_R1095_U158 );
nand NAND2_23852 ( P3_R1095_U208 , P3_U3407 , P3_R1095_U40 );
nand NAND2_23853 ( P3_R1095_U209 , P3_U3070 , P3_R1095_U37 );
nand NAND2_23854 ( P3_R1095_U210 , P3_U3066 , P3_R1095_U36 );
nand NAND2_23855 ( P3_R1095_U211 , P3_R1095_U198 , P3_R1095_U194 );
nand NAND2_23856 ( P3_R1095_U212 , P3_R1095_U6 , P3_R1095_U211 );
nand NAND2_23857 ( P3_R1095_U213 , P3_U3401 , P3_R1095_U42 );
nand NAND2_23858 ( P3_R1095_U214 , P3_U3407 , P3_R1095_U40 );
nand NAND2_23859 ( P3_R1095_U215 , P3_R1095_U13 , P3_R1095_U158 );
not NOT1_23860 ( P3_R1095_U216 , P3_R1095_U44 );
not NOT1_23861 ( P3_R1095_U217 , P3_R1095_U47 );
nand NAND2_23862 ( P3_R1095_U218 , P3_U3413 , P3_R1095_U27 );
nand NAND2_23863 ( P3_R1095_U219 , P3_R1095_U27 , P3_R1095_U26 );
nand NAND2_23864 ( P3_R1095_U220 , P3_U3083 , P3_R1095_U188 );
not NOT1_23865 ( P3_R1095_U221 , P3_R1095_U154 );
nand NAND2_23866 ( P3_R1095_U222 , P3_U3416 , P3_R1095_U46 );
nand NAND2_23867 ( P3_R1095_U223 , P3_R1095_U222 , P3_R1095_U55 );
nand NAND2_23868 ( P3_R1095_U224 , P3_R1095_U217 , P3_R1095_U26 );
nand NAND2_23869 ( P3_R1095_U225 , P3_R1095_U122 , P3_R1095_U224 );
nand NAND2_23870 ( P3_R1095_U226 , P3_R1095_U47 , P3_R1095_U195 );
nand NAND2_23871 ( P3_R1095_U227 , P3_R1095_U121 , P3_R1095_U226 );
nand NAND2_23872 ( P3_R1095_U228 , P3_R1095_U26 , P3_R1095_U195 );
nand NAND2_23873 ( P3_R1095_U229 , P3_R1095_U213 , P3_R1095_U158 );
not NOT1_23874 ( P3_R1095_U230 , P3_R1095_U48 );
nand NAND2_23875 ( P3_R1095_U231 , P3_U3066 , P3_R1095_U36 );
nand NAND2_23876 ( P3_R1095_U232 , P3_R1095_U230 , P3_R1095_U231 );
nand NAND2_23877 ( P3_R1095_U233 , P3_R1095_U124 , P3_R1095_U232 );
nand NAND2_23878 ( P3_R1095_U234 , P3_R1095_U48 , P3_R1095_U194 );
nand NAND2_23879 ( P3_R1095_U235 , P3_U3407 , P3_R1095_U40 );
nand NAND2_23880 ( P3_R1095_U236 , P3_R1095_U123 , P3_R1095_U234 );
nand NAND2_23881 ( P3_R1095_U237 , P3_U3066 , P3_R1095_U36 );
nand NAND2_23882 ( P3_R1095_U238 , P3_R1095_U194 , P3_R1095_U237 );
nand NAND2_23883 ( P3_R1095_U239 , P3_R1095_U213 , P3_R1095_U43 );
nand NAND2_23884 ( P3_R1095_U240 , P3_R1095_U202 , P3_R1095_U34 );
nand NAND2_23885 ( P3_R1095_U241 , P3_R1095_U126 , P3_R1095_U240 );
nand NAND2_23886 ( P3_R1095_U242 , P3_R1095_U49 , P3_R1095_U193 );
nand NAND2_23887 ( P3_R1095_U243 , P3_R1095_U125 , P3_R1095_U242 );
nand NAND2_23888 ( P3_R1095_U244 , P3_R1095_U193 , P3_R1095_U34 );
nand NAND2_23889 ( P3_R1095_U245 , P3_U3422 , P3_R1095_U53 );
nand NAND2_23890 ( P3_R1095_U246 , P3_U3062 , P3_R1095_U51 );
nand NAND2_23891 ( P3_R1095_U247 , P3_U3061 , P3_R1095_U52 );
nand NAND2_23892 ( P3_R1095_U248 , P3_R1095_U199 , P3_R1095_U7 );
nand NAND2_23893 ( P3_R1095_U249 , P3_R1095_U8 , P3_R1095_U248 );
nand NAND2_23894 ( P3_R1095_U250 , P3_U3422 , P3_R1095_U53 );
nand NAND2_23895 ( P3_R1095_U251 , P3_R1095_U127 , P3_R1095_U154 );
nand NAND2_23896 ( P3_R1095_U252 , P3_R1095_U250 , P3_R1095_U249 );
not NOT1_23897 ( P3_R1095_U253 , P3_R1095_U181 );
nand NAND2_23898 ( P3_R1095_U254 , P3_U3425 , P3_R1095_U57 );
nand NAND2_23899 ( P3_R1095_U255 , P3_R1095_U254 , P3_R1095_U181 );
nand NAND2_23900 ( P3_R1095_U256 , P3_U3071 , P3_R1095_U56 );
not NOT1_23901 ( P3_R1095_U257 , P3_R1095_U180 );
nand NAND2_23902 ( P3_R1095_U258 , P3_U3428 , P3_R1095_U59 );
nand NAND2_23903 ( P3_R1095_U259 , P3_R1095_U258 , P3_R1095_U180 );
nand NAND2_23904 ( P3_R1095_U260 , P3_U3079 , P3_R1095_U58 );
not NOT1_23905 ( P3_R1095_U261 , P3_R1095_U179 );
nand NAND2_23906 ( P3_R1095_U262 , P3_U3437 , P3_R1095_U63 );
nand NAND2_23907 ( P3_R1095_U263 , P3_U3072 , P3_R1095_U60 );
nand NAND2_23908 ( P3_R1095_U264 , P3_U3073 , P3_R1095_U61 );
nand NAND2_23909 ( P3_R1095_U265 , P3_R1095_U196 , P3_R1095_U9 );
nand NAND2_23910 ( P3_R1095_U266 , P3_R1095_U10 , P3_R1095_U265 );
nand NAND2_23911 ( P3_R1095_U267 , P3_U3431 , P3_R1095_U65 );
nand NAND2_23912 ( P3_R1095_U268 , P3_U3437 , P3_R1095_U63 );
nand NAND2_23913 ( P3_R1095_U269 , P3_R1095_U128 , P3_R1095_U179 );
nand NAND2_23914 ( P3_R1095_U270 , P3_R1095_U268 , P3_R1095_U266 );
not NOT1_23915 ( P3_R1095_U271 , P3_R1095_U176 );
nand NAND2_23916 ( P3_R1095_U272 , P3_U3440 , P3_R1095_U68 );
nand NAND2_23917 ( P3_R1095_U273 , P3_R1095_U272 , P3_R1095_U176 );
nand NAND2_23918 ( P3_R1095_U274 , P3_U3068 , P3_R1095_U67 );
not NOT1_23919 ( P3_R1095_U275 , P3_R1095_U175 );
nand NAND2_23920 ( P3_R1095_U276 , P3_U3081 , P3_R1095_U175 );
not NOT1_23921 ( P3_R1095_U277 , P3_R1095_U173 );
nand NAND2_23922 ( P3_R1095_U278 , P3_U3445 , P3_R1095_U71 );
nand NAND2_23923 ( P3_R1095_U279 , P3_R1095_U278 , P3_R1095_U173 );
nand NAND2_23924 ( P3_R1095_U280 , P3_U3080 , P3_R1095_U70 );
not NOT1_23925 ( P3_R1095_U281 , P3_R1095_U170 );
nand NAND2_23926 ( P3_R1095_U282 , P3_U3907 , P3_R1095_U73 );
nand NAND2_23927 ( P3_R1095_U283 , P3_R1095_U282 , P3_R1095_U170 );
nand NAND2_23928 ( P3_R1095_U284 , P3_U3075 , P3_R1095_U72 );
not NOT1_23929 ( P3_R1095_U285 , P3_R1095_U169 );
nand NAND2_23930 ( P3_R1095_U286 , P3_U3904 , P3_R1095_U77 );
nand NAND2_23931 ( P3_R1095_U287 , P3_U3065 , P3_R1095_U74 );
nand NAND2_23932 ( P3_R1095_U288 , P3_U3060 , P3_R1095_U75 );
nand NAND2_23933 ( P3_R1095_U289 , P3_R1095_U197 , P3_R1095_U11 );
nand NAND2_23934 ( P3_R1095_U290 , P3_R1095_U12 , P3_R1095_U289 );
nand NAND2_23935 ( P3_R1095_U291 , P3_U3906 , P3_R1095_U79 );
nand NAND2_23936 ( P3_R1095_U292 , P3_U3904 , P3_R1095_U77 );
nand NAND2_23937 ( P3_R1095_U293 , P3_R1095_U129 , P3_R1095_U169 );
nand NAND2_23938 ( P3_R1095_U294 , P3_R1095_U292 , P3_R1095_U290 );
not NOT1_23939 ( P3_R1095_U295 , P3_R1095_U166 );
nand NAND2_23940 ( P3_R1095_U296 , P3_U3903 , P3_R1095_U82 );
nand NAND2_23941 ( P3_R1095_U297 , P3_R1095_U296 , P3_R1095_U166 );
nand NAND2_23942 ( P3_R1095_U298 , P3_U3064 , P3_R1095_U81 );
not NOT1_23943 ( P3_R1095_U299 , P3_R1095_U165 );
nand NAND2_23944 ( P3_R1095_U300 , P3_U3902 , P3_R1095_U84 );
nand NAND2_23945 ( P3_R1095_U301 , P3_R1095_U300 , P3_R1095_U165 );
nand NAND2_23946 ( P3_R1095_U302 , P3_U3057 , P3_R1095_U83 );
not NOT1_23947 ( P3_R1095_U303 , P3_R1095_U91 );
nand NAND2_23948 ( P3_R1095_U304 , P3_R1095_U130 , P3_R1095_U91 );
nand NAND2_23949 ( P3_R1095_U305 , P3_R1095_U88 , P3_R1095_U87 );
nand NAND2_23950 ( P3_R1095_U306 , P3_R1095_U305 , P3_R1095_U85 );
nand NAND2_23951 ( P3_R1095_U307 , P3_U3052 , P3_R1095_U186 );
not NOT1_23952 ( P3_R1095_U308 , P3_R1095_U163 );
nand NAND2_23953 ( P3_R1095_U309 , P3_U3899 , P3_R1095_U90 );
nand NAND2_23954 ( P3_R1095_U310 , P3_U3053 , P3_R1095_U89 );
nand NAND2_23955 ( P3_R1095_U311 , P3_R1095_U303 , P3_R1095_U87 );
nand NAND2_23956 ( P3_R1095_U312 , P3_R1095_U137 , P3_R1095_U311 );
nand NAND2_23957 ( P3_R1095_U313 , P3_R1095_U91 , P3_R1095_U192 );
nand NAND2_23958 ( P3_R1095_U314 , P3_R1095_U136 , P3_R1095_U313 );
nand NAND2_23959 ( P3_R1095_U315 , P3_R1095_U192 , P3_R1095_U87 );
nand NAND2_23960 ( P3_R1095_U316 , P3_R1095_U291 , P3_R1095_U169 );
not NOT1_23961 ( P3_R1095_U317 , P3_R1095_U92 );
nand NAND2_23962 ( P3_R1095_U318 , P3_U3060 , P3_R1095_U75 );
nand NAND2_23963 ( P3_R1095_U319 , P3_R1095_U317 , P3_R1095_U318 );
nand NAND2_23964 ( P3_R1095_U320 , P3_R1095_U141 , P3_R1095_U319 );
nand NAND2_23965 ( P3_R1095_U321 , P3_R1095_U92 , P3_R1095_U191 );
nand NAND2_23966 ( P3_R1095_U322 , P3_U3904 , P3_R1095_U77 );
nand NAND2_23967 ( P3_R1095_U323 , P3_R1095_U140 , P3_R1095_U321 );
nand NAND2_23968 ( P3_R1095_U324 , P3_U3060 , P3_R1095_U75 );
nand NAND2_23969 ( P3_R1095_U325 , P3_R1095_U191 , P3_R1095_U324 );
nand NAND2_23970 ( P3_R1095_U326 , P3_R1095_U291 , P3_R1095_U80 );
nand NAND2_23971 ( P3_R1095_U327 , P3_R1095_U267 , P3_R1095_U179 );
not NOT1_23972 ( P3_R1095_U328 , P3_R1095_U93 );
nand NAND2_23973 ( P3_R1095_U329 , P3_U3073 , P3_R1095_U61 );
nand NAND2_23974 ( P3_R1095_U330 , P3_R1095_U328 , P3_R1095_U329 );
nand NAND2_23975 ( P3_R1095_U331 , P3_R1095_U148 , P3_R1095_U330 );
nand NAND2_23976 ( P3_R1095_U332 , P3_R1095_U93 , P3_R1095_U190 );
nand NAND2_23977 ( P3_R1095_U333 , P3_U3437 , P3_R1095_U63 );
nand NAND2_23978 ( P3_R1095_U334 , P3_R1095_U147 , P3_R1095_U332 );
nand NAND2_23979 ( P3_R1095_U335 , P3_U3073 , P3_R1095_U61 );
nand NAND2_23980 ( P3_R1095_U336 , P3_R1095_U190 , P3_R1095_U335 );
nand NAND2_23981 ( P3_R1095_U337 , P3_R1095_U267 , P3_R1095_U66 );
nand NAND2_23982 ( P3_R1095_U338 , P3_R1095_U222 , P3_R1095_U154 );
not NOT1_23983 ( P3_R1095_U339 , P3_R1095_U94 );
nand NAND2_23984 ( P3_R1095_U340 , P3_U3061 , P3_R1095_U52 );
nand NAND2_23985 ( P3_R1095_U341 , P3_R1095_U339 , P3_R1095_U340 );
nand NAND2_23986 ( P3_R1095_U342 , P3_R1095_U152 , P3_R1095_U341 );
nand NAND2_23987 ( P3_R1095_U343 , P3_R1095_U94 , P3_R1095_U189 );
nand NAND2_23988 ( P3_R1095_U344 , P3_U3422 , P3_R1095_U53 );
nand NAND2_23989 ( P3_R1095_U345 , P3_R1095_U151 , P3_R1095_U343 );
nand NAND2_23990 ( P3_R1095_U346 , P3_U3061 , P3_R1095_U52 );
nand NAND2_23991 ( P3_R1095_U347 , P3_R1095_U189 , P3_R1095_U346 );
nand NAND2_23992 ( P3_R1095_U348 , P3_U3076 , P3_R1095_U30 );
nand NAND2_23993 ( P3_R1095_U349 , P3_U3077 , P3_R1095_U171 );
nand NAND2_23994 ( P3_R1095_U350 , P3_U3081 , P3_R1095_U174 );
nand NAND3_23995 ( P3_R1095_U351 , P3_R1095_U133 , P3_R1095_U304 , P3_R1095_U134 );
nand NAND2_23996 ( P3_R1095_U352 , P3_U3398 , P3_R1095_U35 );
nand NAND2_23997 ( P3_R1095_U353 , P3_U3413 , P3_R1095_U220 );
nand NAND2_23998 ( P3_R1095_U354 , P3_R1095_U353 , P3_R1095_U219 );
nand NAND2_23999 ( P3_R1095_U355 , P3_U3900 , P3_R1095_U88 );
nand NAND2_24000 ( P3_R1095_U356 , P3_R1095_U119 , P3_R1095_U158 );
nand NAND2_24001 ( P3_R1095_U357 , P3_R1095_U216 , P3_R1095_U14 );
nand NAND2_24002 ( P3_R1095_U358 , P3_U3416 , P3_R1095_U46 );
nand NAND2_24003 ( P3_R1095_U359 , P3_U3082 , P3_R1095_U45 );
nand NAND2_24004 ( P3_R1095_U360 , P3_R1095_U223 , P3_R1095_U154 );
nand NAND2_24005 ( P3_R1095_U361 , P3_R1095_U221 , P3_R1095_U153 );
nand NAND2_24006 ( P3_R1095_U362 , P3_U3413 , P3_R1095_U27 );
nand NAND2_24007 ( P3_R1095_U363 , P3_U3083 , P3_R1095_U28 );
nand NAND2_24008 ( P3_R1095_U364 , P3_U3413 , P3_R1095_U27 );
nand NAND2_24009 ( P3_R1095_U365 , P3_U3083 , P3_R1095_U28 );
nand NAND2_24010 ( P3_R1095_U366 , P3_R1095_U365 , P3_R1095_U364 );
nand NAND2_24011 ( P3_R1095_U367 , P3_U3410 , P3_R1095_U25 );
nand NAND2_24012 ( P3_R1095_U368 , P3_U3069 , P3_R1095_U39 );
nand NAND2_24013 ( P3_R1095_U369 , P3_R1095_U228 , P3_R1095_U47 );
nand NAND2_24014 ( P3_R1095_U370 , P3_R1095_U155 , P3_R1095_U217 );
nand NAND2_24015 ( P3_R1095_U371 , P3_U3407 , P3_R1095_U40 );
nand NAND2_24016 ( P3_R1095_U372 , P3_U3070 , P3_R1095_U37 );
nand NAND2_24017 ( P3_R1095_U373 , P3_R1095_U372 , P3_R1095_U371 );
nand NAND2_24018 ( P3_R1095_U374 , P3_U3404 , P3_R1095_U41 );
nand NAND2_24019 ( P3_R1095_U375 , P3_U3066 , P3_R1095_U36 );
nand NAND2_24020 ( P3_R1095_U376 , P3_R1095_U238 , P3_R1095_U48 );
nand NAND2_24021 ( P3_R1095_U377 , P3_R1095_U156 , P3_R1095_U230 );
nand NAND2_24022 ( P3_R1095_U378 , P3_U3401 , P3_R1095_U42 );
nand NAND2_24023 ( P3_R1095_U379 , P3_U3059 , P3_R1095_U38 );
nand NAND2_24024 ( P3_R1095_U380 , P3_R1095_U239 , P3_R1095_U158 );
nand NAND2_24025 ( P3_R1095_U381 , P3_R1095_U207 , P3_R1095_U157 );
nand NAND2_24026 ( P3_R1095_U382 , P3_U3398 , P3_R1095_U35 );
nand NAND2_24027 ( P3_R1095_U383 , P3_U3063 , P3_R1095_U32 );
nand NAND2_24028 ( P3_R1095_U384 , P3_U3398 , P3_R1095_U35 );
nand NAND2_24029 ( P3_R1095_U385 , P3_U3063 , P3_R1095_U32 );
nand NAND2_24030 ( P3_R1095_U386 , P3_R1095_U385 , P3_R1095_U384 );
nand NAND2_24031 ( P3_R1095_U387 , P3_U3395 , P3_R1095_U33 );
nand NAND2_24032 ( P3_R1095_U388 , P3_U3067 , P3_R1095_U29 );
nand NAND2_24033 ( P3_R1095_U389 , P3_R1095_U244 , P3_R1095_U49 );
nand NAND2_24034 ( P3_R1095_U390 , P3_R1095_U159 , P3_R1095_U202 );
nand NAND2_24035 ( P3_R1095_U391 , P3_U3908 , P3_R1095_U161 );
nand NAND2_24036 ( P3_R1095_U392 , P3_U3054 , P3_R1095_U160 );
nand NAND2_24037 ( P3_R1095_U393 , P3_U3908 , P3_R1095_U161 );
nand NAND2_24038 ( P3_R1095_U394 , P3_U3054 , P3_R1095_U160 );
nand NAND2_24039 ( P3_R1095_U395 , P3_R1095_U394 , P3_R1095_U393 );
nand NAND3_24040 ( P3_R1095_U396 , P3_U3053 , P3_R1095_U395 , P3_R1095_U89 );
nand NAND3_24041 ( P3_R1095_U397 , P3_R1095_U15 , P3_R1095_U90 , P3_U3899 );
nand NAND2_24042 ( P3_R1095_U398 , P3_U3899 , P3_R1095_U90 );
nand NAND2_24043 ( P3_R1095_U399 , P3_U3053 , P3_R1095_U89 );
not NOT1_24044 ( P3_R1095_U400 , P3_R1095_U135 );
nand NAND2_24045 ( P3_R1095_U401 , P3_R1095_U308 , P3_R1095_U400 );
nand NAND2_24046 ( P3_R1095_U402 , P3_R1095_U135 , P3_R1095_U163 );
nand NAND2_24047 ( P3_R1095_U403 , P3_U3900 , P3_R1095_U88 );
nand NAND2_24048 ( P3_R1095_U404 , P3_U3052 , P3_R1095_U85 );
nand NAND2_24049 ( P3_R1095_U405 , P3_U3900 , P3_R1095_U88 );
nand NAND2_24050 ( P3_R1095_U406 , P3_U3052 , P3_R1095_U85 );
nand NAND2_24051 ( P3_R1095_U407 , P3_R1095_U406 , P3_R1095_U405 );
nand NAND2_24052 ( P3_R1095_U408 , P3_U3901 , P3_R1095_U86 );
nand NAND2_24053 ( P3_R1095_U409 , P3_U3056 , P3_R1095_U50 );
nand NAND2_24054 ( P3_R1095_U410 , P3_R1095_U315 , P3_R1095_U91 );
nand NAND2_24055 ( P3_R1095_U411 , P3_R1095_U164 , P3_R1095_U303 );
nand NAND2_24056 ( P3_R1095_U412 , P3_U3902 , P3_R1095_U84 );
nand NAND2_24057 ( P3_R1095_U413 , P3_U3057 , P3_R1095_U83 );
not NOT1_24058 ( P3_R1095_U414 , P3_R1095_U138 );
nand NAND2_24059 ( P3_R1095_U415 , P3_R1095_U299 , P3_R1095_U414 );
nand NAND2_24060 ( P3_R1095_U416 , P3_R1095_U138 , P3_R1095_U165 );
nand NAND2_24061 ( P3_R1095_U417 , P3_U3903 , P3_R1095_U82 );
nand NAND2_24062 ( P3_R1095_U418 , P3_U3064 , P3_R1095_U81 );
not NOT1_24063 ( P3_R1095_U419 , P3_R1095_U139 );
nand NAND2_24064 ( P3_R1095_U420 , P3_R1095_U295 , P3_R1095_U419 );
nand NAND2_24065 ( P3_R1095_U421 , P3_R1095_U139 , P3_R1095_U166 );
nand NAND2_24066 ( P3_R1095_U422 , P3_U3904 , P3_R1095_U77 );
nand NAND2_24067 ( P3_R1095_U423 , P3_U3065 , P3_R1095_U74 );
nand NAND2_24068 ( P3_R1095_U424 , P3_R1095_U423 , P3_R1095_U422 );
nand NAND2_24069 ( P3_R1095_U425 , P3_U3905 , P3_R1095_U78 );
nand NAND2_24070 ( P3_R1095_U426 , P3_U3060 , P3_R1095_U75 );
nand NAND2_24071 ( P3_R1095_U427 , P3_R1095_U325 , P3_R1095_U92 );
nand NAND2_24072 ( P3_R1095_U428 , P3_R1095_U167 , P3_R1095_U317 );
nand NAND2_24073 ( P3_R1095_U429 , P3_U3906 , P3_R1095_U79 );
nand NAND2_24074 ( P3_R1095_U430 , P3_U3074 , P3_R1095_U76 );
nand NAND2_24075 ( P3_R1095_U431 , P3_R1095_U326 , P3_R1095_U169 );
nand NAND2_24076 ( P3_R1095_U432 , P3_R1095_U285 , P3_R1095_U168 );
nand NAND2_24077 ( P3_R1095_U433 , P3_U3907 , P3_R1095_U73 );
nand NAND2_24078 ( P3_R1095_U434 , P3_U3075 , P3_R1095_U72 );
not NOT1_24079 ( P3_R1095_U435 , P3_R1095_U142 );
nand NAND2_24080 ( P3_R1095_U436 , P3_R1095_U281 , P3_R1095_U435 );
nand NAND2_24081 ( P3_R1095_U437 , P3_R1095_U142 , P3_R1095_U170 );
nand NAND2_24082 ( P3_R1095_U438 , P3_U3392 , P3_R1095_U31 );
nand NAND2_24083 ( P3_R1095_U439 , P3_U3077 , P3_R1095_U171 );
not NOT1_24084 ( P3_R1095_U440 , P3_R1095_U143 );
nand NAND2_24085 ( P3_R1095_U441 , P3_R1095_U200 , P3_R1095_U440 );
nand NAND2_24086 ( P3_R1095_U442 , P3_R1095_U143 , P3_R1095_U172 );
nand NAND2_24087 ( P3_R1095_U443 , P3_U3445 , P3_R1095_U71 );
nand NAND2_24088 ( P3_R1095_U444 , P3_U3080 , P3_R1095_U70 );
not NOT1_24089 ( P3_R1095_U445 , P3_R1095_U144 );
nand NAND2_24090 ( P3_R1095_U446 , P3_R1095_U277 , P3_R1095_U445 );
nand NAND2_24091 ( P3_R1095_U447 , P3_R1095_U144 , P3_R1095_U173 );
nand NAND2_24092 ( P3_R1095_U448 , P3_U3443 , P3_R1095_U69 );
nand NAND2_24093 ( P3_R1095_U449 , P3_U3081 , P3_R1095_U174 );
not NOT1_24094 ( P3_R1095_U450 , P3_R1095_U145 );
nand NAND2_24095 ( P3_R1095_U451 , P3_R1095_U275 , P3_R1095_U450 );
nand NAND2_24096 ( P3_R1095_U452 , P3_R1095_U145 , P3_R1095_U175 );
nand NAND2_24097 ( P3_R1095_U453 , P3_U3440 , P3_R1095_U68 );
nand NAND2_24098 ( P3_R1095_U454 , P3_U3068 , P3_R1095_U67 );
not NOT1_24099 ( P3_R1095_U455 , P3_R1095_U146 );
nand NAND2_24100 ( P3_R1095_U456 , P3_R1095_U271 , P3_R1095_U455 );
nand NAND2_24101 ( P3_R1095_U457 , P3_R1095_U146 , P3_R1095_U176 );
nand NAND2_24102 ( P3_R1095_U458 , P3_U3437 , P3_R1095_U63 );
nand NAND2_24103 ( P3_R1095_U459 , P3_U3072 , P3_R1095_U60 );
nand NAND2_24104 ( P3_R1095_U460 , P3_R1095_U459 , P3_R1095_U458 );
nand NAND2_24105 ( P3_R1095_U461 , P3_U3434 , P3_R1095_U64 );
nand NAND2_24106 ( P3_R1095_U462 , P3_U3073 , P3_R1095_U61 );
nand NAND2_24107 ( P3_R1095_U463 , P3_R1095_U336 , P3_R1095_U93 );
nand NAND2_24108 ( P3_R1095_U464 , P3_R1095_U177 , P3_R1095_U328 );
nand NAND2_24109 ( P3_R1095_U465 , P3_U3431 , P3_R1095_U65 );
nand NAND2_24110 ( P3_R1095_U466 , P3_U3078 , P3_R1095_U62 );
nand NAND2_24111 ( P3_R1095_U467 , P3_R1095_U337 , P3_R1095_U179 );
nand NAND2_24112 ( P3_R1095_U468 , P3_R1095_U261 , P3_R1095_U178 );
nand NAND2_24113 ( P3_R1095_U469 , P3_U3428 , P3_R1095_U59 );
nand NAND2_24114 ( P3_R1095_U470 , P3_U3079 , P3_R1095_U58 );
not NOT1_24115 ( P3_R1095_U471 , P3_R1095_U149 );
nand NAND2_24116 ( P3_R1095_U472 , P3_R1095_U257 , P3_R1095_U471 );
nand NAND2_24117 ( P3_R1095_U473 , P3_R1095_U149 , P3_R1095_U180 );
nand NAND2_24118 ( P3_R1095_U474 , P3_U3425 , P3_R1095_U57 );
nand NAND2_24119 ( P3_R1095_U475 , P3_U3071 , P3_R1095_U56 );
not NOT1_24120 ( P3_R1095_U476 , P3_R1095_U150 );
nand NAND2_24121 ( P3_R1095_U477 , P3_R1095_U253 , P3_R1095_U476 );
nand NAND2_24122 ( P3_R1095_U478 , P3_R1095_U150 , P3_R1095_U181 );
nand NAND2_24123 ( P3_R1095_U479 , P3_U3422 , P3_R1095_U53 );
nand NAND2_24124 ( P3_R1095_U480 , P3_U3062 , P3_R1095_U51 );
nand NAND2_24125 ( P3_R1095_U481 , P3_R1095_U480 , P3_R1095_U479 );
nand NAND2_24126 ( P3_R1095_U482 , P3_U3419 , P3_R1095_U54 );
nand NAND2_24127 ( P3_R1095_U483 , P3_U3061 , P3_R1095_U52 );
nand NAND2_24128 ( P3_R1095_U484 , P3_R1095_U347 , P3_R1095_U94 );
nand NAND2_24129 ( P3_R1095_U485 , P3_R1095_U182 , P3_R1095_U339 );
nand NAND2_24130 ( P3_R1212_U6 , P3_R1212_U176 , P3_R1212_U180 );
nand NAND2_24131 ( P3_R1212_U7 , P3_R1212_U9 , P3_R1212_U181 );
not NOT1_24132 ( P3_R1212_U8 , P3_REG2_REG_0_ );
nand NAND2_24133 ( P3_R1212_U9 , P3_REG2_REG_0_ , P3_R1212_U48 );
not NOT1_24134 ( P3_R1212_U10 , P3_REG2_REG_1_ );
not NOT1_24135 ( P3_R1212_U11 , P3_U3391 );
not NOT1_24136 ( P3_R1212_U12 , P3_REG2_REG_2_ );
not NOT1_24137 ( P3_R1212_U13 , P3_U3394 );
not NOT1_24138 ( P3_R1212_U14 , P3_REG2_REG_3_ );
not NOT1_24139 ( P3_R1212_U15 , P3_U3397 );
not NOT1_24140 ( P3_R1212_U16 , P3_REG2_REG_4_ );
not NOT1_24141 ( P3_R1212_U17 , P3_U3400 );
not NOT1_24142 ( P3_R1212_U18 , P3_REG2_REG_5_ );
not NOT1_24143 ( P3_R1212_U19 , P3_U3403 );
not NOT1_24144 ( P3_R1212_U20 , P3_REG2_REG_6_ );
not NOT1_24145 ( P3_R1212_U21 , P3_U3406 );
not NOT1_24146 ( P3_R1212_U22 , P3_REG2_REG_7_ );
not NOT1_24147 ( P3_R1212_U23 , P3_U3409 );
not NOT1_24148 ( P3_R1212_U24 , P3_REG2_REG_8_ );
not NOT1_24149 ( P3_R1212_U25 , P3_U3412 );
not NOT1_24150 ( P3_R1212_U26 , P3_REG2_REG_9_ );
not NOT1_24151 ( P3_R1212_U27 , P3_U3415 );
not NOT1_24152 ( P3_R1212_U28 , P3_REG2_REG_10_ );
not NOT1_24153 ( P3_R1212_U29 , P3_U3418 );
not NOT1_24154 ( P3_R1212_U30 , P3_REG2_REG_11_ );
not NOT1_24155 ( P3_R1212_U31 , P3_U3421 );
not NOT1_24156 ( P3_R1212_U32 , P3_REG2_REG_12_ );
not NOT1_24157 ( P3_R1212_U33 , P3_U3424 );
not NOT1_24158 ( P3_R1212_U34 , P3_REG2_REG_13_ );
not NOT1_24159 ( P3_R1212_U35 , P3_U3427 );
not NOT1_24160 ( P3_R1212_U36 , P3_REG2_REG_14_ );
not NOT1_24161 ( P3_R1212_U37 , P3_U3430 );
nand NAND2_24162 ( P3_R1212_U38 , P3_R1212_U159 , P3_R1212_U158 );
not NOT1_24163 ( P3_R1212_U39 , P3_REG2_REG_15_ );
not NOT1_24164 ( P3_R1212_U40 , P3_U3433 );
not NOT1_24165 ( P3_R1212_U41 , P3_REG2_REG_16_ );
not NOT1_24166 ( P3_R1212_U42 , P3_U3436 );
not NOT1_24167 ( P3_R1212_U43 , P3_REG2_REG_17_ );
not NOT1_24168 ( P3_R1212_U44 , P3_U3439 );
not NOT1_24169 ( P3_R1212_U45 , P3_REG2_REG_18_ );
not NOT1_24170 ( P3_R1212_U46 , P3_U3442 );
nand NAND2_24171 ( P3_R1212_U47 , P3_R1212_U171 , P3_R1212_U170 );
not NOT1_24172 ( P3_R1212_U48 , P3_U3386 );
nand NAND2_24173 ( P3_R1212_U49 , P3_R1212_U186 , P3_R1212_U185 );
nand NAND2_24174 ( P3_R1212_U50 , P3_R1212_U191 , P3_R1212_U190 );
nand NAND2_24175 ( P3_R1212_U51 , P3_R1212_U196 , P3_R1212_U195 );
nand NAND2_24176 ( P3_R1212_U52 , P3_R1212_U201 , P3_R1212_U200 );
nand NAND2_24177 ( P3_R1212_U53 , P3_R1212_U206 , P3_R1212_U205 );
nand NAND2_24178 ( P3_R1212_U54 , P3_R1212_U211 , P3_R1212_U210 );
nand NAND2_24179 ( P3_R1212_U55 , P3_R1212_U216 , P3_R1212_U215 );
nand NAND2_24180 ( P3_R1212_U56 , P3_R1212_U221 , P3_R1212_U220 );
nand NAND2_24181 ( P3_R1212_U57 , P3_R1212_U226 , P3_R1212_U225 );
nand NAND2_24182 ( P3_R1212_U58 , P3_R1212_U236 , P3_R1212_U235 );
nand NAND2_24183 ( P3_R1212_U59 , P3_R1212_U241 , P3_R1212_U240 );
nand NAND2_24184 ( P3_R1212_U60 , P3_R1212_U246 , P3_R1212_U245 );
nand NAND2_24185 ( P3_R1212_U61 , P3_R1212_U251 , P3_R1212_U250 );
nand NAND2_24186 ( P3_R1212_U62 , P3_R1212_U256 , P3_R1212_U255 );
nand NAND2_24187 ( P3_R1212_U63 , P3_R1212_U261 , P3_R1212_U260 );
nand NAND2_24188 ( P3_R1212_U64 , P3_R1212_U266 , P3_R1212_U265 );
nand NAND2_24189 ( P3_R1212_U65 , P3_R1212_U271 , P3_R1212_U270 );
nand NAND2_24190 ( P3_R1212_U66 , P3_R1212_U276 , P3_R1212_U275 );
nand NAND2_24191 ( P3_R1212_U67 , P3_R1212_U183 , P3_R1212_U182 );
nand NAND2_24192 ( P3_R1212_U68 , P3_R1212_U188 , P3_R1212_U187 );
nand NAND2_24193 ( P3_R1212_U69 , P3_R1212_U193 , P3_R1212_U192 );
nand NAND2_24194 ( P3_R1212_U70 , P3_R1212_U198 , P3_R1212_U197 );
nand NAND2_24195 ( P3_R1212_U71 , P3_R1212_U203 , P3_R1212_U202 );
nand NAND2_24196 ( P3_R1212_U72 , P3_R1212_U208 , P3_R1212_U207 );
nand NAND2_24197 ( P3_R1212_U73 , P3_R1212_U213 , P3_R1212_U212 );
nand NAND2_24198 ( P3_R1212_U74 , P3_R1212_U218 , P3_R1212_U217 );
nand NAND2_24199 ( P3_R1212_U75 , P3_R1212_U223 , P3_R1212_U222 );
and AND3_24200 ( P3_R1212_U76 , P3_R1212_U228 , P3_R1212_U227 , P3_R1212_U179 );
and AND2_24201 ( P3_R1212_U77 , P3_R1212_U175 , P3_R1212_U231 );
nand NAND2_24202 ( P3_R1212_U78 , P3_R1212_U233 , P3_R1212_U232 );
nand NAND2_24203 ( P3_R1212_U79 , P3_R1212_U238 , P3_R1212_U237 );
nand NAND2_24204 ( P3_R1212_U80 , P3_R1212_U243 , P3_R1212_U242 );
nand NAND2_24205 ( P3_R1212_U81 , P3_R1212_U248 , P3_R1212_U247 );
nand NAND2_24206 ( P3_R1212_U82 , P3_R1212_U253 , P3_R1212_U252 );
nand NAND2_24207 ( P3_R1212_U83 , P3_R1212_U258 , P3_R1212_U257 );
nand NAND2_24208 ( P3_R1212_U84 , P3_R1212_U263 , P3_R1212_U262 );
nand NAND2_24209 ( P3_R1212_U85 , P3_R1212_U268 , P3_R1212_U267 );
nand NAND2_24210 ( P3_R1212_U86 , P3_R1212_U273 , P3_R1212_U272 );
nand NAND2_24211 ( P3_R1212_U87 , P3_R1212_U135 , P3_R1212_U134 );
nand NAND2_24212 ( P3_R1212_U88 , P3_R1212_U131 , P3_R1212_U130 );
nand NAND2_24213 ( P3_R1212_U89 , P3_R1212_U127 , P3_R1212_U126 );
nand NAND2_24214 ( P3_R1212_U90 , P3_R1212_U123 , P3_R1212_U122 );
nand NAND2_24215 ( P3_R1212_U91 , P3_R1212_U119 , P3_R1212_U118 );
nand NAND2_24216 ( P3_R1212_U92 , P3_R1212_U115 , P3_R1212_U114 );
nand NAND2_24217 ( P3_R1212_U93 , P3_R1212_U111 , P3_R1212_U110 );
nand NAND2_24218 ( P3_R1212_U94 , P3_R1212_U107 , P3_R1212_U106 );
not NOT1_24219 ( P3_R1212_U95 , P3_REG2_REG_19_ );
not NOT1_24220 ( P3_R1212_U96 , P3_U3379 );
nand NAND2_24221 ( P3_R1212_U97 , P3_R1212_U167 , P3_R1212_U166 );
nand NAND2_24222 ( P3_R1212_U98 , P3_R1212_U163 , P3_R1212_U162 );
nand NAND2_24223 ( P3_R1212_U99 , P3_R1212_U155 , P3_R1212_U154 );
nand NAND2_24224 ( P3_R1212_U100 , P3_R1212_U151 , P3_R1212_U150 );
nand NAND2_24225 ( P3_R1212_U101 , P3_R1212_U147 , P3_R1212_U146 );
nand NAND2_24226 ( P3_R1212_U102 , P3_R1212_U143 , P3_R1212_U142 );
nand NAND2_24227 ( P3_R1212_U103 , P3_R1212_U139 , P3_R1212_U138 );
not NOT1_24228 ( P3_R1212_U104 , P3_R1212_U9 );
nand NAND2_24229 ( P3_R1212_U105 , P3_REG2_REG_1_ , P3_R1212_U104 );
nand NAND2_24230 ( P3_R1212_U106 , P3_U3391 , P3_R1212_U105 );
nand NAND2_24231 ( P3_R1212_U107 , P3_R1212_U9 , P3_R1212_U10 );
not NOT1_24232 ( P3_R1212_U108 , P3_R1212_U94 );
nand NAND2_24233 ( P3_R1212_U109 , P3_REG2_REG_2_ , P3_R1212_U13 );
nand NAND2_24234 ( P3_R1212_U110 , P3_R1212_U109 , P3_R1212_U94 );
nand NAND2_24235 ( P3_R1212_U111 , P3_U3394 , P3_R1212_U12 );
not NOT1_24236 ( P3_R1212_U112 , P3_R1212_U93 );
nand NAND2_24237 ( P3_R1212_U113 , P3_REG2_REG_3_ , P3_R1212_U15 );
nand NAND2_24238 ( P3_R1212_U114 , P3_R1212_U113 , P3_R1212_U93 );
nand NAND2_24239 ( P3_R1212_U115 , P3_U3397 , P3_R1212_U14 );
not NOT1_24240 ( P3_R1212_U116 , P3_R1212_U92 );
nand NAND2_24241 ( P3_R1212_U117 , P3_REG2_REG_4_ , P3_R1212_U17 );
nand NAND2_24242 ( P3_R1212_U118 , P3_R1212_U117 , P3_R1212_U92 );
nand NAND2_24243 ( P3_R1212_U119 , P3_U3400 , P3_R1212_U16 );
not NOT1_24244 ( P3_R1212_U120 , P3_R1212_U91 );
nand NAND2_24245 ( P3_R1212_U121 , P3_REG2_REG_5_ , P3_R1212_U19 );
nand NAND2_24246 ( P3_R1212_U122 , P3_R1212_U121 , P3_R1212_U91 );
nand NAND2_24247 ( P3_R1212_U123 , P3_U3403 , P3_R1212_U18 );
not NOT1_24248 ( P3_R1212_U124 , P3_R1212_U90 );
nand NAND2_24249 ( P3_R1212_U125 , P3_REG2_REG_6_ , P3_R1212_U21 );
nand NAND2_24250 ( P3_R1212_U126 , P3_R1212_U125 , P3_R1212_U90 );
nand NAND2_24251 ( P3_R1212_U127 , P3_U3406 , P3_R1212_U20 );
not NOT1_24252 ( P3_R1212_U128 , P3_R1212_U89 );
nand NAND2_24253 ( P3_R1212_U129 , P3_REG2_REG_7_ , P3_R1212_U23 );
nand NAND2_24254 ( P3_R1212_U130 , P3_R1212_U129 , P3_R1212_U89 );
nand NAND2_24255 ( P3_R1212_U131 , P3_U3409 , P3_R1212_U22 );
not NOT1_24256 ( P3_R1212_U132 , P3_R1212_U88 );
nand NAND2_24257 ( P3_R1212_U133 , P3_REG2_REG_8_ , P3_R1212_U25 );
nand NAND2_24258 ( P3_R1212_U134 , P3_R1212_U133 , P3_R1212_U88 );
nand NAND2_24259 ( P3_R1212_U135 , P3_U3412 , P3_R1212_U24 );
not NOT1_24260 ( P3_R1212_U136 , P3_R1212_U87 );
nand NAND2_24261 ( P3_R1212_U137 , P3_REG2_REG_9_ , P3_R1212_U27 );
nand NAND2_24262 ( P3_R1212_U138 , P3_R1212_U137 , P3_R1212_U87 );
nand NAND2_24263 ( P3_R1212_U139 , P3_U3415 , P3_R1212_U26 );
not NOT1_24264 ( P3_R1212_U140 , P3_R1212_U103 );
nand NAND2_24265 ( P3_R1212_U141 , P3_REG2_REG_10_ , P3_R1212_U29 );
nand NAND2_24266 ( P3_R1212_U142 , P3_R1212_U141 , P3_R1212_U103 );
nand NAND2_24267 ( P3_R1212_U143 , P3_U3418 , P3_R1212_U28 );
not NOT1_24268 ( P3_R1212_U144 , P3_R1212_U102 );
nand NAND2_24269 ( P3_R1212_U145 , P3_REG2_REG_11_ , P3_R1212_U31 );
nand NAND2_24270 ( P3_R1212_U146 , P3_R1212_U145 , P3_R1212_U102 );
nand NAND2_24271 ( P3_R1212_U147 , P3_U3421 , P3_R1212_U30 );
not NOT1_24272 ( P3_R1212_U148 , P3_R1212_U101 );
nand NAND2_24273 ( P3_R1212_U149 , P3_REG2_REG_12_ , P3_R1212_U33 );
nand NAND2_24274 ( P3_R1212_U150 , P3_R1212_U149 , P3_R1212_U101 );
nand NAND2_24275 ( P3_R1212_U151 , P3_U3424 , P3_R1212_U32 );
not NOT1_24276 ( P3_R1212_U152 , P3_R1212_U100 );
nand NAND2_24277 ( P3_R1212_U153 , P3_REG2_REG_13_ , P3_R1212_U35 );
nand NAND2_24278 ( P3_R1212_U154 , P3_R1212_U153 , P3_R1212_U100 );
nand NAND2_24279 ( P3_R1212_U155 , P3_U3427 , P3_R1212_U34 );
not NOT1_24280 ( P3_R1212_U156 , P3_R1212_U99 );
nand NAND2_24281 ( P3_R1212_U157 , P3_REG2_REG_14_ , P3_R1212_U37 );
nand NAND2_24282 ( P3_R1212_U158 , P3_R1212_U157 , P3_R1212_U99 );
nand NAND2_24283 ( P3_R1212_U159 , P3_U3430 , P3_R1212_U36 );
not NOT1_24284 ( P3_R1212_U160 , P3_R1212_U38 );
nand NAND2_24285 ( P3_R1212_U161 , P3_REG2_REG_15_ , P3_R1212_U160 );
nand NAND2_24286 ( P3_R1212_U162 , P3_U3433 , P3_R1212_U161 );
nand NAND2_24287 ( P3_R1212_U163 , P3_R1212_U38 , P3_R1212_U39 );
not NOT1_24288 ( P3_R1212_U164 , P3_R1212_U98 );
nand NAND2_24289 ( P3_R1212_U165 , P3_REG2_REG_16_ , P3_R1212_U42 );
nand NAND2_24290 ( P3_R1212_U166 , P3_R1212_U165 , P3_R1212_U98 );
nand NAND2_24291 ( P3_R1212_U167 , P3_U3436 , P3_R1212_U41 );
not NOT1_24292 ( P3_R1212_U168 , P3_R1212_U97 );
nand NAND2_24293 ( P3_R1212_U169 , P3_REG2_REG_17_ , P3_R1212_U44 );
nand NAND2_24294 ( P3_R1212_U170 , P3_R1212_U169 , P3_R1212_U97 );
nand NAND2_24295 ( P3_R1212_U171 , P3_U3439 , P3_R1212_U43 );
not NOT1_24296 ( P3_R1212_U172 , P3_R1212_U47 );
nand NAND2_24297 ( P3_R1212_U173 , P3_U3442 , P3_R1212_U45 );
nand NAND2_24298 ( P3_R1212_U174 , P3_R1212_U172 , P3_R1212_U173 );
nand NAND2_24299 ( P3_R1212_U175 , P3_REG2_REG_18_ , P3_R1212_U46 );
nand NAND2_24300 ( P3_R1212_U176 , P3_R1212_U77 , P3_R1212_U174 );
nand NAND2_24301 ( P3_R1212_U177 , P3_REG2_REG_18_ , P3_R1212_U46 );
nand NAND2_24302 ( P3_R1212_U178 , P3_R1212_U177 , P3_R1212_U47 );
nand NAND2_24303 ( P3_R1212_U179 , P3_U3442 , P3_R1212_U45 );
nand NAND2_24304 ( P3_R1212_U180 , P3_R1212_U76 , P3_R1212_U178 );
nand NAND2_24305 ( P3_R1212_U181 , P3_U3386 , P3_R1212_U8 );
nand NAND2_24306 ( P3_R1212_U182 , P3_REG2_REG_9_ , P3_R1212_U27 );
nand NAND2_24307 ( P3_R1212_U183 , P3_U3415 , P3_R1212_U26 );
not NOT1_24308 ( P3_R1212_U184 , P3_R1212_U67 );
nand NAND2_24309 ( P3_R1212_U185 , P3_R1212_U136 , P3_R1212_U184 );
nand NAND2_24310 ( P3_R1212_U186 , P3_R1212_U67 , P3_R1212_U87 );
nand NAND2_24311 ( P3_R1212_U187 , P3_REG2_REG_8_ , P3_R1212_U25 );
nand NAND2_24312 ( P3_R1212_U188 , P3_U3412 , P3_R1212_U24 );
not NOT1_24313 ( P3_R1212_U189 , P3_R1212_U68 );
nand NAND2_24314 ( P3_R1212_U190 , P3_R1212_U132 , P3_R1212_U189 );
nand NAND2_24315 ( P3_R1212_U191 , P3_R1212_U68 , P3_R1212_U88 );
nand NAND2_24316 ( P3_R1212_U192 , P3_REG2_REG_7_ , P3_R1212_U23 );
nand NAND2_24317 ( P3_R1212_U193 , P3_U3409 , P3_R1212_U22 );
not NOT1_24318 ( P3_R1212_U194 , P3_R1212_U69 );
nand NAND2_24319 ( P3_R1212_U195 , P3_R1212_U128 , P3_R1212_U194 );
nand NAND2_24320 ( P3_R1212_U196 , P3_R1212_U69 , P3_R1212_U89 );
nand NAND2_24321 ( P3_R1212_U197 , P3_REG2_REG_6_ , P3_R1212_U21 );
nand NAND2_24322 ( P3_R1212_U198 , P3_U3406 , P3_R1212_U20 );
not NOT1_24323 ( P3_R1212_U199 , P3_R1212_U70 );
nand NAND2_24324 ( P3_R1212_U200 , P3_R1212_U124 , P3_R1212_U199 );
nand NAND2_24325 ( P3_R1212_U201 , P3_R1212_U70 , P3_R1212_U90 );
nand NAND2_24326 ( P3_R1212_U202 , P3_REG2_REG_5_ , P3_R1212_U19 );
nand NAND2_24327 ( P3_R1212_U203 , P3_U3403 , P3_R1212_U18 );
not NOT1_24328 ( P3_R1212_U204 , P3_R1212_U71 );
nand NAND2_24329 ( P3_R1212_U205 , P3_R1212_U120 , P3_R1212_U204 );
nand NAND2_24330 ( P3_R1212_U206 , P3_R1212_U71 , P3_R1212_U91 );
nand NAND2_24331 ( P3_R1212_U207 , P3_REG2_REG_4_ , P3_R1212_U17 );
nand NAND2_24332 ( P3_R1212_U208 , P3_U3400 , P3_R1212_U16 );
not NOT1_24333 ( P3_R1212_U209 , P3_R1212_U72 );
nand NAND2_24334 ( P3_R1212_U210 , P3_R1212_U116 , P3_R1212_U209 );
nand NAND2_24335 ( P3_R1212_U211 , P3_R1212_U72 , P3_R1212_U92 );
nand NAND2_24336 ( P3_R1212_U212 , P3_REG2_REG_3_ , P3_R1212_U15 );
nand NAND2_24337 ( P3_R1212_U213 , P3_U3397 , P3_R1212_U14 );
not NOT1_24338 ( P3_R1212_U214 , P3_R1212_U73 );
nand NAND2_24339 ( P3_R1212_U215 , P3_R1212_U112 , P3_R1212_U214 );
nand NAND2_24340 ( P3_R1212_U216 , P3_R1212_U73 , P3_R1212_U93 );
nand NAND2_24341 ( P3_R1212_U217 , P3_REG2_REG_2_ , P3_R1212_U13 );
nand NAND2_24342 ( P3_R1212_U218 , P3_U3394 , P3_R1212_U12 );
not NOT1_24343 ( P3_R1212_U219 , P3_R1212_U74 );
nand NAND2_24344 ( P3_R1212_U220 , P3_R1212_U108 , P3_R1212_U219 );
nand NAND2_24345 ( P3_R1212_U221 , P3_R1212_U74 , P3_R1212_U94 );
nand NAND2_24346 ( P3_R1212_U222 , P3_R1212_U104 , P3_R1212_U10 );
nand NAND2_24347 ( P3_R1212_U223 , P3_REG2_REG_1_ , P3_R1212_U9 );
not NOT1_24348 ( P3_R1212_U224 , P3_R1212_U75 );
nand NAND2_24349 ( P3_R1212_U225 , P3_R1212_U224 , P3_U3391 );
nand NAND2_24350 ( P3_R1212_U226 , P3_R1212_U75 , P3_R1212_U11 );
nand NAND2_24351 ( P3_R1212_U227 , P3_REG2_REG_19_ , P3_R1212_U96 );
nand NAND2_24352 ( P3_R1212_U228 , P3_U3379 , P3_R1212_U95 );
nand NAND2_24353 ( P3_R1212_U229 , P3_REG2_REG_19_ , P3_R1212_U96 );
nand NAND2_24354 ( P3_R1212_U230 , P3_U3379 , P3_R1212_U95 );
nand NAND2_24355 ( P3_R1212_U231 , P3_R1212_U230 , P3_R1212_U229 );
nand NAND2_24356 ( P3_R1212_U232 , P3_REG2_REG_18_ , P3_R1212_U46 );
nand NAND2_24357 ( P3_R1212_U233 , P3_U3442 , P3_R1212_U45 );
not NOT1_24358 ( P3_R1212_U234 , P3_R1212_U78 );
nand NAND2_24359 ( P3_R1212_U235 , P3_R1212_U234 , P3_R1212_U172 );
nand NAND2_24360 ( P3_R1212_U236 , P3_R1212_U78 , P3_R1212_U47 );
nand NAND2_24361 ( P3_R1212_U237 , P3_REG2_REG_17_ , P3_R1212_U44 );
nand NAND2_24362 ( P3_R1212_U238 , P3_U3439 , P3_R1212_U43 );
not NOT1_24363 ( P3_R1212_U239 , P3_R1212_U79 );
nand NAND2_24364 ( P3_R1212_U240 , P3_R1212_U168 , P3_R1212_U239 );
nand NAND2_24365 ( P3_R1212_U241 , P3_R1212_U79 , P3_R1212_U97 );
nand NAND2_24366 ( P3_R1212_U242 , P3_REG2_REG_16_ , P3_R1212_U42 );
nand NAND2_24367 ( P3_R1212_U243 , P3_U3436 , P3_R1212_U41 );
not NOT1_24368 ( P3_R1212_U244 , P3_R1212_U80 );
nand NAND2_24369 ( P3_R1212_U245 , P3_R1212_U164 , P3_R1212_U244 );
nand NAND2_24370 ( P3_R1212_U246 , P3_R1212_U80 , P3_R1212_U98 );
nand NAND2_24371 ( P3_R1212_U247 , P3_U3433 , P3_R1212_U39 );
nand NAND2_24372 ( P3_R1212_U248 , P3_REG2_REG_15_ , P3_R1212_U40 );
not NOT1_24373 ( P3_R1212_U249 , P3_R1212_U81 );
nand NAND2_24374 ( P3_R1212_U250 , P3_R1212_U249 , P3_R1212_U160 );
nand NAND2_24375 ( P3_R1212_U251 , P3_R1212_U81 , P3_R1212_U38 );
nand NAND2_24376 ( P3_R1212_U252 , P3_REG2_REG_14_ , P3_R1212_U37 );
nand NAND2_24377 ( P3_R1212_U253 , P3_U3430 , P3_R1212_U36 );
not NOT1_24378 ( P3_R1212_U254 , P3_R1212_U82 );
nand NAND2_24379 ( P3_R1212_U255 , P3_R1212_U156 , P3_R1212_U254 );
nand NAND2_24380 ( P3_R1212_U256 , P3_R1212_U82 , P3_R1212_U99 );
nand NAND2_24381 ( P3_R1212_U257 , P3_REG2_REG_13_ , P3_R1212_U35 );
nand NAND2_24382 ( P3_R1212_U258 , P3_U3427 , P3_R1212_U34 );
not NOT1_24383 ( P3_R1212_U259 , P3_R1212_U83 );
nand NAND2_24384 ( P3_R1212_U260 , P3_R1212_U152 , P3_R1212_U259 );
nand NAND2_24385 ( P3_R1212_U261 , P3_R1212_U83 , P3_R1212_U100 );
nand NAND2_24386 ( P3_R1212_U262 , P3_REG2_REG_12_ , P3_R1212_U33 );
nand NAND2_24387 ( P3_R1212_U263 , P3_U3424 , P3_R1212_U32 );
not NOT1_24388 ( P3_R1212_U264 , P3_R1212_U84 );
nand NAND2_24389 ( P3_R1212_U265 , P3_R1212_U148 , P3_R1212_U264 );
nand NAND2_24390 ( P3_R1212_U266 , P3_R1212_U84 , P3_R1212_U101 );
nand NAND2_24391 ( P3_R1212_U267 , P3_REG2_REG_11_ , P3_R1212_U31 );
nand NAND2_24392 ( P3_R1212_U268 , P3_U3421 , P3_R1212_U30 );
not NOT1_24393 ( P3_R1212_U269 , P3_R1212_U85 );
nand NAND2_24394 ( P3_R1212_U270 , P3_R1212_U144 , P3_R1212_U269 );
nand NAND2_24395 ( P3_R1212_U271 , P3_R1212_U85 , P3_R1212_U102 );
nand NAND2_24396 ( P3_R1212_U272 , P3_REG2_REG_10_ , P3_R1212_U29 );
nand NAND2_24397 ( P3_R1212_U273 , P3_U3418 , P3_R1212_U28 );
not NOT1_24398 ( P3_R1212_U274 , P3_R1212_U86 );
nand NAND2_24399 ( P3_R1212_U275 , P3_R1212_U140 , P3_R1212_U274 );
nand NAND2_24400 ( P3_R1212_U276 , P3_R1212_U86 , P3_R1212_U103 );
nand NAND2_24401 ( P3_R1209_U6 , P3_R1209_U176 , P3_R1209_U180 );
nand NAND2_24402 ( P3_R1209_U7 , P3_R1209_U9 , P3_R1209_U181 );
not NOT1_24403 ( P3_R1209_U8 , P3_REG1_REG_0_ );
nand NAND2_24404 ( P3_R1209_U9 , P3_REG1_REG_0_ , P3_R1209_U48 );
not NOT1_24405 ( P3_R1209_U10 , P3_REG1_REG_1_ );
not NOT1_24406 ( P3_R1209_U11 , P3_U3391 );
not NOT1_24407 ( P3_R1209_U12 , P3_REG1_REG_2_ );
not NOT1_24408 ( P3_R1209_U13 , P3_U3394 );
not NOT1_24409 ( P3_R1209_U14 , P3_REG1_REG_3_ );
not NOT1_24410 ( P3_R1209_U15 , P3_U3397 );
not NOT1_24411 ( P3_R1209_U16 , P3_REG1_REG_4_ );
not NOT1_24412 ( P3_R1209_U17 , P3_U3400 );
not NOT1_24413 ( P3_R1209_U18 , P3_REG1_REG_5_ );
not NOT1_24414 ( P3_R1209_U19 , P3_U3403 );
not NOT1_24415 ( P3_R1209_U20 , P3_REG1_REG_6_ );
not NOT1_24416 ( P3_R1209_U21 , P3_U3406 );
not NOT1_24417 ( P3_R1209_U22 , P3_REG1_REG_7_ );
not NOT1_24418 ( P3_R1209_U23 , P3_U3409 );
not NOT1_24419 ( P3_R1209_U24 , P3_REG1_REG_8_ );
not NOT1_24420 ( P3_R1209_U25 , P3_U3412 );
not NOT1_24421 ( P3_R1209_U26 , P3_REG1_REG_9_ );
not NOT1_24422 ( P3_R1209_U27 , P3_U3415 );
not NOT1_24423 ( P3_R1209_U28 , P3_REG1_REG_10_ );
not NOT1_24424 ( P3_R1209_U29 , P3_U3418 );
not NOT1_24425 ( P3_R1209_U30 , P3_REG1_REG_11_ );
not NOT1_24426 ( P3_R1209_U31 , P3_U3421 );
not NOT1_24427 ( P3_R1209_U32 , P3_REG1_REG_12_ );
not NOT1_24428 ( P3_R1209_U33 , P3_U3424 );
not NOT1_24429 ( P3_R1209_U34 , P3_REG1_REG_13_ );
not NOT1_24430 ( P3_R1209_U35 , P3_U3427 );
not NOT1_24431 ( P3_R1209_U36 , P3_REG1_REG_14_ );
not NOT1_24432 ( P3_R1209_U37 , P3_U3430 );
nand NAND2_24433 ( P3_R1209_U38 , P3_R1209_U159 , P3_R1209_U158 );
not NOT1_24434 ( P3_R1209_U39 , P3_REG1_REG_15_ );
not NOT1_24435 ( P3_R1209_U40 , P3_U3433 );
not NOT1_24436 ( P3_R1209_U41 , P3_REG1_REG_16_ );
not NOT1_24437 ( P3_R1209_U42 , P3_U3436 );
not NOT1_24438 ( P3_R1209_U43 , P3_REG1_REG_17_ );
not NOT1_24439 ( P3_R1209_U44 , P3_U3439 );
not NOT1_24440 ( P3_R1209_U45 , P3_REG1_REG_18_ );
not NOT1_24441 ( P3_R1209_U46 , P3_U3442 );
nand NAND2_24442 ( P3_R1209_U47 , P3_R1209_U171 , P3_R1209_U170 );
not NOT1_24443 ( P3_R1209_U48 , P3_U3386 );
nand NAND2_24444 ( P3_R1209_U49 , P3_R1209_U186 , P3_R1209_U185 );
nand NAND2_24445 ( P3_R1209_U50 , P3_R1209_U191 , P3_R1209_U190 );
nand NAND2_24446 ( P3_R1209_U51 , P3_R1209_U196 , P3_R1209_U195 );
nand NAND2_24447 ( P3_R1209_U52 , P3_R1209_U201 , P3_R1209_U200 );
nand NAND2_24448 ( P3_R1209_U53 , P3_R1209_U206 , P3_R1209_U205 );
nand NAND2_24449 ( P3_R1209_U54 , P3_R1209_U211 , P3_R1209_U210 );
nand NAND2_24450 ( P3_R1209_U55 , P3_R1209_U216 , P3_R1209_U215 );
nand NAND2_24451 ( P3_R1209_U56 , P3_R1209_U221 , P3_R1209_U220 );
nand NAND2_24452 ( P3_R1209_U57 , P3_R1209_U226 , P3_R1209_U225 );
nand NAND2_24453 ( P3_R1209_U58 , P3_R1209_U236 , P3_R1209_U235 );
nand NAND2_24454 ( P3_R1209_U59 , P3_R1209_U241 , P3_R1209_U240 );
nand NAND2_24455 ( P3_R1209_U60 , P3_R1209_U246 , P3_R1209_U245 );
nand NAND2_24456 ( P3_R1209_U61 , P3_R1209_U251 , P3_R1209_U250 );
nand NAND2_24457 ( P3_R1209_U62 , P3_R1209_U256 , P3_R1209_U255 );
nand NAND2_24458 ( P3_R1209_U63 , P3_R1209_U261 , P3_R1209_U260 );
nand NAND2_24459 ( P3_R1209_U64 , P3_R1209_U266 , P3_R1209_U265 );
nand NAND2_24460 ( P3_R1209_U65 , P3_R1209_U271 , P3_R1209_U270 );
nand NAND2_24461 ( P3_R1209_U66 , P3_R1209_U276 , P3_R1209_U275 );
nand NAND2_24462 ( P3_R1209_U67 , P3_R1209_U183 , P3_R1209_U182 );
nand NAND2_24463 ( P3_R1209_U68 , P3_R1209_U188 , P3_R1209_U187 );
nand NAND2_24464 ( P3_R1209_U69 , P3_R1209_U193 , P3_R1209_U192 );
nand NAND2_24465 ( P3_R1209_U70 , P3_R1209_U198 , P3_R1209_U197 );
nand NAND2_24466 ( P3_R1209_U71 , P3_R1209_U203 , P3_R1209_U202 );
nand NAND2_24467 ( P3_R1209_U72 , P3_R1209_U208 , P3_R1209_U207 );
nand NAND2_24468 ( P3_R1209_U73 , P3_R1209_U213 , P3_R1209_U212 );
nand NAND2_24469 ( P3_R1209_U74 , P3_R1209_U218 , P3_R1209_U217 );
nand NAND2_24470 ( P3_R1209_U75 , P3_R1209_U223 , P3_R1209_U222 );
and AND3_24471 ( P3_R1209_U76 , P3_R1209_U228 , P3_R1209_U227 , P3_R1209_U179 );
and AND2_24472 ( P3_R1209_U77 , P3_R1209_U175 , P3_R1209_U231 );
nand NAND2_24473 ( P3_R1209_U78 , P3_R1209_U233 , P3_R1209_U232 );
nand NAND2_24474 ( P3_R1209_U79 , P3_R1209_U238 , P3_R1209_U237 );
nand NAND2_24475 ( P3_R1209_U80 , P3_R1209_U243 , P3_R1209_U242 );
nand NAND2_24476 ( P3_R1209_U81 , P3_R1209_U248 , P3_R1209_U247 );
nand NAND2_24477 ( P3_R1209_U82 , P3_R1209_U253 , P3_R1209_U252 );
nand NAND2_24478 ( P3_R1209_U83 , P3_R1209_U258 , P3_R1209_U257 );
nand NAND2_24479 ( P3_R1209_U84 , P3_R1209_U263 , P3_R1209_U262 );
nand NAND2_24480 ( P3_R1209_U85 , P3_R1209_U268 , P3_R1209_U267 );
nand NAND2_24481 ( P3_R1209_U86 , P3_R1209_U273 , P3_R1209_U272 );
nand NAND2_24482 ( P3_R1209_U87 , P3_R1209_U135 , P3_R1209_U134 );
nand NAND2_24483 ( P3_R1209_U88 , P3_R1209_U131 , P3_R1209_U130 );
nand NAND2_24484 ( P3_R1209_U89 , P3_R1209_U127 , P3_R1209_U126 );
nand NAND2_24485 ( P3_R1209_U90 , P3_R1209_U123 , P3_R1209_U122 );
nand NAND2_24486 ( P3_R1209_U91 , P3_R1209_U119 , P3_R1209_U118 );
nand NAND2_24487 ( P3_R1209_U92 , P3_R1209_U115 , P3_R1209_U114 );
nand NAND2_24488 ( P3_R1209_U93 , P3_R1209_U111 , P3_R1209_U110 );
nand NAND2_24489 ( P3_R1209_U94 , P3_R1209_U107 , P3_R1209_U106 );
not NOT1_24490 ( P3_R1209_U95 , P3_REG1_REG_19_ );
not NOT1_24491 ( P3_R1209_U96 , P3_U3379 );
nand NAND2_24492 ( P3_R1209_U97 , P3_R1209_U167 , P3_R1209_U166 );
nand NAND2_24493 ( P3_R1209_U98 , P3_R1209_U163 , P3_R1209_U162 );
nand NAND2_24494 ( P3_R1209_U99 , P3_R1209_U155 , P3_R1209_U154 );
nand NAND2_24495 ( P3_R1209_U100 , P3_R1209_U151 , P3_R1209_U150 );
nand NAND2_24496 ( P3_R1209_U101 , P3_R1209_U147 , P3_R1209_U146 );
nand NAND2_24497 ( P3_R1209_U102 , P3_R1209_U143 , P3_R1209_U142 );
nand NAND2_24498 ( P3_R1209_U103 , P3_R1209_U139 , P3_R1209_U138 );
not NOT1_24499 ( P3_R1209_U104 , P3_R1209_U9 );
nand NAND2_24500 ( P3_R1209_U105 , P3_REG1_REG_1_ , P3_R1209_U104 );
nand NAND2_24501 ( P3_R1209_U106 , P3_U3391 , P3_R1209_U105 );
nand NAND2_24502 ( P3_R1209_U107 , P3_R1209_U9 , P3_R1209_U10 );
not NOT1_24503 ( P3_R1209_U108 , P3_R1209_U94 );
nand NAND2_24504 ( P3_R1209_U109 , P3_REG1_REG_2_ , P3_R1209_U13 );
nand NAND2_24505 ( P3_R1209_U110 , P3_R1209_U109 , P3_R1209_U94 );
nand NAND2_24506 ( P3_R1209_U111 , P3_U3394 , P3_R1209_U12 );
not NOT1_24507 ( P3_R1209_U112 , P3_R1209_U93 );
nand NAND2_24508 ( P3_R1209_U113 , P3_REG1_REG_3_ , P3_R1209_U15 );
nand NAND2_24509 ( P3_R1209_U114 , P3_R1209_U113 , P3_R1209_U93 );
nand NAND2_24510 ( P3_R1209_U115 , P3_U3397 , P3_R1209_U14 );
not NOT1_24511 ( P3_R1209_U116 , P3_R1209_U92 );
nand NAND2_24512 ( P3_R1209_U117 , P3_REG1_REG_4_ , P3_R1209_U17 );
nand NAND2_24513 ( P3_R1209_U118 , P3_R1209_U117 , P3_R1209_U92 );
nand NAND2_24514 ( P3_R1209_U119 , P3_U3400 , P3_R1209_U16 );
not NOT1_24515 ( P3_R1209_U120 , P3_R1209_U91 );
nand NAND2_24516 ( P3_R1209_U121 , P3_REG1_REG_5_ , P3_R1209_U19 );
nand NAND2_24517 ( P3_R1209_U122 , P3_R1209_U121 , P3_R1209_U91 );
nand NAND2_24518 ( P3_R1209_U123 , P3_U3403 , P3_R1209_U18 );
not NOT1_24519 ( P3_R1209_U124 , P3_R1209_U90 );
nand NAND2_24520 ( P3_R1209_U125 , P3_REG1_REG_6_ , P3_R1209_U21 );
nand NAND2_24521 ( P3_R1209_U126 , P3_R1209_U125 , P3_R1209_U90 );
nand NAND2_24522 ( P3_R1209_U127 , P3_U3406 , P3_R1209_U20 );
not NOT1_24523 ( P3_R1209_U128 , P3_R1209_U89 );
nand NAND2_24524 ( P3_R1209_U129 , P3_REG1_REG_7_ , P3_R1209_U23 );
nand NAND2_24525 ( P3_R1209_U130 , P3_R1209_U129 , P3_R1209_U89 );
nand NAND2_24526 ( P3_R1209_U131 , P3_U3409 , P3_R1209_U22 );
not NOT1_24527 ( P3_R1209_U132 , P3_R1209_U88 );
nand NAND2_24528 ( P3_R1209_U133 , P3_REG1_REG_8_ , P3_R1209_U25 );
nand NAND2_24529 ( P3_R1209_U134 , P3_R1209_U133 , P3_R1209_U88 );
nand NAND2_24530 ( P3_R1209_U135 , P3_U3412 , P3_R1209_U24 );
not NOT1_24531 ( P3_R1209_U136 , P3_R1209_U87 );
nand NAND2_24532 ( P3_R1209_U137 , P3_REG1_REG_9_ , P3_R1209_U27 );
nand NAND2_24533 ( P3_R1209_U138 , P3_R1209_U137 , P3_R1209_U87 );
nand NAND2_24534 ( P3_R1209_U139 , P3_U3415 , P3_R1209_U26 );
not NOT1_24535 ( P3_R1209_U140 , P3_R1209_U103 );
nand NAND2_24536 ( P3_R1209_U141 , P3_REG1_REG_10_ , P3_R1209_U29 );
nand NAND2_24537 ( P3_R1209_U142 , P3_R1209_U141 , P3_R1209_U103 );
nand NAND2_24538 ( P3_R1209_U143 , P3_U3418 , P3_R1209_U28 );
not NOT1_24539 ( P3_R1209_U144 , P3_R1209_U102 );
nand NAND2_24540 ( P3_R1209_U145 , P3_REG1_REG_11_ , P3_R1209_U31 );
nand NAND2_24541 ( P3_R1209_U146 , P3_R1209_U145 , P3_R1209_U102 );
nand NAND2_24542 ( P3_R1209_U147 , P3_U3421 , P3_R1209_U30 );
not NOT1_24543 ( P3_R1209_U148 , P3_R1209_U101 );
nand NAND2_24544 ( P3_R1209_U149 , P3_REG1_REG_12_ , P3_R1209_U33 );
nand NAND2_24545 ( P3_R1209_U150 , P3_R1209_U149 , P3_R1209_U101 );
nand NAND2_24546 ( P3_R1209_U151 , P3_U3424 , P3_R1209_U32 );
not NOT1_24547 ( P3_R1209_U152 , P3_R1209_U100 );
nand NAND2_24548 ( P3_R1209_U153 , P3_REG1_REG_13_ , P3_R1209_U35 );
nand NAND2_24549 ( P3_R1209_U154 , P3_R1209_U153 , P3_R1209_U100 );
nand NAND2_24550 ( P3_R1209_U155 , P3_U3427 , P3_R1209_U34 );
not NOT1_24551 ( P3_R1209_U156 , P3_R1209_U99 );
nand NAND2_24552 ( P3_R1209_U157 , P3_REG1_REG_14_ , P3_R1209_U37 );
nand NAND2_24553 ( P3_R1209_U158 , P3_R1209_U157 , P3_R1209_U99 );
nand NAND2_24554 ( P3_R1209_U159 , P3_U3430 , P3_R1209_U36 );
not NOT1_24555 ( P3_R1209_U160 , P3_R1209_U38 );
nand NAND2_24556 ( P3_R1209_U161 , P3_REG1_REG_15_ , P3_R1209_U160 );
nand NAND2_24557 ( P3_R1209_U162 , P3_U3433 , P3_R1209_U161 );
nand NAND2_24558 ( P3_R1209_U163 , P3_R1209_U38 , P3_R1209_U39 );
not NOT1_24559 ( P3_R1209_U164 , P3_R1209_U98 );
nand NAND2_24560 ( P3_R1209_U165 , P3_REG1_REG_16_ , P3_R1209_U42 );
nand NAND2_24561 ( P3_R1209_U166 , P3_R1209_U165 , P3_R1209_U98 );
nand NAND2_24562 ( P3_R1209_U167 , P3_U3436 , P3_R1209_U41 );
not NOT1_24563 ( P3_R1209_U168 , P3_R1209_U97 );
nand NAND2_24564 ( P3_R1209_U169 , P3_REG1_REG_17_ , P3_R1209_U44 );
nand NAND2_24565 ( P3_R1209_U170 , P3_R1209_U169 , P3_R1209_U97 );
nand NAND2_24566 ( P3_R1209_U171 , P3_U3439 , P3_R1209_U43 );
not NOT1_24567 ( P3_R1209_U172 , P3_R1209_U47 );
nand NAND2_24568 ( P3_R1209_U173 , P3_U3442 , P3_R1209_U45 );
nand NAND2_24569 ( P3_R1209_U174 , P3_R1209_U172 , P3_R1209_U173 );
nand NAND2_24570 ( P3_R1209_U175 , P3_REG1_REG_18_ , P3_R1209_U46 );
nand NAND2_24571 ( P3_R1209_U176 , P3_R1209_U77 , P3_R1209_U174 );
nand NAND2_24572 ( P3_R1209_U177 , P3_REG1_REG_18_ , P3_R1209_U46 );
nand NAND2_24573 ( P3_R1209_U178 , P3_R1209_U177 , P3_R1209_U47 );
nand NAND2_24574 ( P3_R1209_U179 , P3_U3442 , P3_R1209_U45 );
nand NAND2_24575 ( P3_R1209_U180 , P3_R1209_U76 , P3_R1209_U178 );
nand NAND2_24576 ( P3_R1209_U181 , P3_U3386 , P3_R1209_U8 );
nand NAND2_24577 ( P3_R1209_U182 , P3_REG1_REG_9_ , P3_R1209_U27 );
nand NAND2_24578 ( P3_R1209_U183 , P3_U3415 , P3_R1209_U26 );
not NOT1_24579 ( P3_R1209_U184 , P3_R1209_U67 );
nand NAND2_24580 ( P3_R1209_U185 , P3_R1209_U136 , P3_R1209_U184 );
nand NAND2_24581 ( P3_R1209_U186 , P3_R1209_U67 , P3_R1209_U87 );
nand NAND2_24582 ( P3_R1209_U187 , P3_REG1_REG_8_ , P3_R1209_U25 );
nand NAND2_24583 ( P3_R1209_U188 , P3_U3412 , P3_R1209_U24 );
not NOT1_24584 ( P3_R1209_U189 , P3_R1209_U68 );
nand NAND2_24585 ( P3_R1209_U190 , P3_R1209_U132 , P3_R1209_U189 );
nand NAND2_24586 ( P3_R1209_U191 , P3_R1209_U68 , P3_R1209_U88 );
nand NAND2_24587 ( P3_R1209_U192 , P3_REG1_REG_7_ , P3_R1209_U23 );
nand NAND2_24588 ( P3_R1209_U193 , P3_U3409 , P3_R1209_U22 );
not NOT1_24589 ( P3_R1209_U194 , P3_R1209_U69 );
nand NAND2_24590 ( P3_R1209_U195 , P3_R1209_U128 , P3_R1209_U194 );
nand NAND2_24591 ( P3_R1209_U196 , P3_R1209_U69 , P3_R1209_U89 );
nand NAND2_24592 ( P3_R1209_U197 , P3_REG1_REG_6_ , P3_R1209_U21 );
nand NAND2_24593 ( P3_R1209_U198 , P3_U3406 , P3_R1209_U20 );
not NOT1_24594 ( P3_R1209_U199 , P3_R1209_U70 );
nand NAND2_24595 ( P3_R1209_U200 , P3_R1209_U124 , P3_R1209_U199 );
nand NAND2_24596 ( P3_R1209_U201 , P3_R1209_U70 , P3_R1209_U90 );
nand NAND2_24597 ( P3_R1209_U202 , P3_REG1_REG_5_ , P3_R1209_U19 );
nand NAND2_24598 ( P3_R1209_U203 , P3_U3403 , P3_R1209_U18 );
not NOT1_24599 ( P3_R1209_U204 , P3_R1209_U71 );
nand NAND2_24600 ( P3_R1209_U205 , P3_R1209_U120 , P3_R1209_U204 );
nand NAND2_24601 ( P3_R1209_U206 , P3_R1209_U71 , P3_R1209_U91 );
nand NAND2_24602 ( P3_R1209_U207 , P3_REG1_REG_4_ , P3_R1209_U17 );
nand NAND2_24603 ( P3_R1209_U208 , P3_U3400 , P3_R1209_U16 );
not NOT1_24604 ( P3_R1209_U209 , P3_R1209_U72 );
nand NAND2_24605 ( P3_R1209_U210 , P3_R1209_U116 , P3_R1209_U209 );
nand NAND2_24606 ( P3_R1209_U211 , P3_R1209_U72 , P3_R1209_U92 );
nand NAND2_24607 ( P3_R1209_U212 , P3_REG1_REG_3_ , P3_R1209_U15 );
nand NAND2_24608 ( P3_R1209_U213 , P3_U3397 , P3_R1209_U14 );
not NOT1_24609 ( P3_R1209_U214 , P3_R1209_U73 );
nand NAND2_24610 ( P3_R1209_U215 , P3_R1209_U112 , P3_R1209_U214 );
nand NAND2_24611 ( P3_R1209_U216 , P3_R1209_U73 , P3_R1209_U93 );
nand NAND2_24612 ( P3_R1209_U217 , P3_REG1_REG_2_ , P3_R1209_U13 );
nand NAND2_24613 ( P3_R1209_U218 , P3_U3394 , P3_R1209_U12 );
not NOT1_24614 ( P3_R1209_U219 , P3_R1209_U74 );
nand NAND2_24615 ( P3_R1209_U220 , P3_R1209_U108 , P3_R1209_U219 );
nand NAND2_24616 ( P3_R1209_U221 , P3_R1209_U74 , P3_R1209_U94 );
nand NAND2_24617 ( P3_R1209_U222 , P3_R1209_U104 , P3_R1209_U10 );
nand NAND2_24618 ( P3_R1209_U223 , P3_REG1_REG_1_ , P3_R1209_U9 );
not NOT1_24619 ( P3_R1209_U224 , P3_R1209_U75 );
nand NAND2_24620 ( P3_R1209_U225 , P3_R1209_U224 , P3_U3391 );
nand NAND2_24621 ( P3_R1209_U226 , P3_R1209_U75 , P3_R1209_U11 );
nand NAND2_24622 ( P3_R1209_U227 , P3_REG1_REG_19_ , P3_R1209_U96 );
nand NAND2_24623 ( P3_R1209_U228 , P3_U3379 , P3_R1209_U95 );
nand NAND2_24624 ( P3_R1209_U229 , P3_REG1_REG_19_ , P3_R1209_U96 );
nand NAND2_24625 ( P3_R1209_U230 , P3_U3379 , P3_R1209_U95 );
nand NAND2_24626 ( P3_R1209_U231 , P3_R1209_U230 , P3_R1209_U229 );
nand NAND2_24627 ( P3_R1209_U232 , P3_REG1_REG_18_ , P3_R1209_U46 );
nand NAND2_24628 ( P3_R1209_U233 , P3_U3442 , P3_R1209_U45 );
not NOT1_24629 ( P3_R1209_U234 , P3_R1209_U78 );
nand NAND2_24630 ( P3_R1209_U235 , P3_R1209_U234 , P3_R1209_U172 );
nand NAND2_24631 ( P3_R1209_U236 , P3_R1209_U78 , P3_R1209_U47 );
nand NAND2_24632 ( P3_R1209_U237 , P3_REG1_REG_17_ , P3_R1209_U44 );
nand NAND2_24633 ( P3_R1209_U238 , P3_U3439 , P3_R1209_U43 );
not NOT1_24634 ( P3_R1209_U239 , P3_R1209_U79 );
nand NAND2_24635 ( P3_R1209_U240 , P3_R1209_U168 , P3_R1209_U239 );
nand NAND2_24636 ( P3_R1209_U241 , P3_R1209_U79 , P3_R1209_U97 );
nand NAND2_24637 ( P3_R1209_U242 , P3_REG1_REG_16_ , P3_R1209_U42 );
nand NAND2_24638 ( P3_R1209_U243 , P3_U3436 , P3_R1209_U41 );
not NOT1_24639 ( P3_R1209_U244 , P3_R1209_U80 );
nand NAND2_24640 ( P3_R1209_U245 , P3_R1209_U164 , P3_R1209_U244 );
nand NAND2_24641 ( P3_R1209_U246 , P3_R1209_U80 , P3_R1209_U98 );
nand NAND2_24642 ( P3_R1209_U247 , P3_U3433 , P3_R1209_U39 );
nand NAND2_24643 ( P3_R1209_U248 , P3_REG1_REG_15_ , P3_R1209_U40 );
not NOT1_24644 ( P3_R1209_U249 , P3_R1209_U81 );
nand NAND2_24645 ( P3_R1209_U250 , P3_R1209_U249 , P3_R1209_U160 );
nand NAND2_24646 ( P3_R1209_U251 , P3_R1209_U81 , P3_R1209_U38 );
nand NAND2_24647 ( P3_R1209_U252 , P3_REG1_REG_14_ , P3_R1209_U37 );
nand NAND2_24648 ( P3_R1209_U253 , P3_U3430 , P3_R1209_U36 );
not NOT1_24649 ( P3_R1209_U254 , P3_R1209_U82 );
nand NAND2_24650 ( P3_R1209_U255 , P3_R1209_U156 , P3_R1209_U254 );
nand NAND2_24651 ( P3_R1209_U256 , P3_R1209_U82 , P3_R1209_U99 );
nand NAND2_24652 ( P3_R1209_U257 , P3_REG1_REG_13_ , P3_R1209_U35 );
nand NAND2_24653 ( P3_R1209_U258 , P3_U3427 , P3_R1209_U34 );
not NOT1_24654 ( P3_R1209_U259 , P3_R1209_U83 );
nand NAND2_24655 ( P3_R1209_U260 , P3_R1209_U152 , P3_R1209_U259 );
nand NAND2_24656 ( P3_R1209_U261 , P3_R1209_U83 , P3_R1209_U100 );
nand NAND2_24657 ( P3_R1209_U262 , P3_REG1_REG_12_ , P3_R1209_U33 );
nand NAND2_24658 ( P3_R1209_U263 , P3_U3424 , P3_R1209_U32 );
not NOT1_24659 ( P3_R1209_U264 , P3_R1209_U84 );
nand NAND2_24660 ( P3_R1209_U265 , P3_R1209_U148 , P3_R1209_U264 );
nand NAND2_24661 ( P3_R1209_U266 , P3_R1209_U84 , P3_R1209_U101 );
nand NAND2_24662 ( P3_R1209_U267 , P3_REG1_REG_11_ , P3_R1209_U31 );
nand NAND2_24663 ( P3_R1209_U268 , P3_U3421 , P3_R1209_U30 );
not NOT1_24664 ( P3_R1209_U269 , P3_R1209_U85 );
nand NAND2_24665 ( P3_R1209_U270 , P3_R1209_U144 , P3_R1209_U269 );
nand NAND2_24666 ( P3_R1209_U271 , P3_R1209_U85 , P3_R1209_U102 );
nand NAND2_24667 ( P3_R1209_U272 , P3_REG1_REG_10_ , P3_R1209_U29 );
nand NAND2_24668 ( P3_R1209_U273 , P3_U3418 , P3_R1209_U28 );
not NOT1_24669 ( P3_R1209_U274 , P3_R1209_U86 );
nand NAND2_24670 ( P3_R1209_U275 , P3_R1209_U140 , P3_R1209_U274 );
nand NAND2_24671 ( P3_R1209_U276 , P3_R1209_U86 , P3_R1209_U103 );
not NOT1_24672 ( P3_R1300_U6 , P3_U3058 );
not NOT1_24673 ( P3_R1300_U7 , P3_U3055 );
and AND2_24674 ( P3_R1300_U8 , P3_R1300_U10 , P3_R1300_U9 );
nand NAND2_24675 ( P3_R1300_U9 , P3_U3055 , P3_R1300_U6 );
nand NAND2_24676 ( P3_R1300_U10 , P3_U3058 , P3_R1300_U7 );
and AND2_24677 ( P3_R1200_U6 , P3_R1200_U210 , P3_R1200_U209 );
and AND2_24678 ( P3_R1200_U7 , P3_R1200_U189 , P3_R1200_U245 );
and AND2_24679 ( P3_R1200_U8 , P3_R1200_U247 , P3_R1200_U246 );
and AND2_24680 ( P3_R1200_U9 , P3_R1200_U190 , P3_R1200_U262 );
and AND2_24681 ( P3_R1200_U10 , P3_R1200_U264 , P3_R1200_U263 );
and AND2_24682 ( P3_R1200_U11 , P3_R1200_U191 , P3_R1200_U286 );
and AND2_24683 ( P3_R1200_U12 , P3_R1200_U288 , P3_R1200_U287 );
and AND3_24684 ( P3_R1200_U13 , P3_R1200_U208 , P3_R1200_U194 , P3_R1200_U213 );
and AND2_24685 ( P3_R1200_U14 , P3_R1200_U218 , P3_R1200_U195 );
and AND2_24686 ( P3_R1200_U15 , P3_R1200_U392 , P3_R1200_U391 );
nand NAND2_24687 ( P3_R1200_U16 , P3_R1200_U342 , P3_R1200_U345 );
nand NAND2_24688 ( P3_R1200_U17 , P3_R1200_U331 , P3_R1200_U334 );
nand NAND2_24689 ( P3_R1200_U18 , P3_R1200_U320 , P3_R1200_U323 );
nand NAND2_24690 ( P3_R1200_U19 , P3_R1200_U312 , P3_R1200_U314 );
nand NAND3_24691 ( P3_R1200_U20 , P3_R1200_U162 , P3_R1200_U183 , P3_R1200_U351 );
nand NAND2_24692 ( P3_R1200_U21 , P3_R1200_U241 , P3_R1200_U243 );
nand NAND2_24693 ( P3_R1200_U22 , P3_R1200_U233 , P3_R1200_U236 );
nand NAND2_24694 ( P3_R1200_U23 , P3_R1200_U225 , P3_R1200_U227 );
nand NAND2_24695 ( P3_R1200_U24 , P3_R1200_U172 , P3_R1200_U348 );
not NOT1_24696 ( P3_R1200_U25 , P3_U3069 );
nand NAND2_24697 ( P3_R1200_U26 , P3_U3069 , P3_R1200_U39 );
not NOT1_24698 ( P3_R1200_U27 , P3_U3083 );
not NOT1_24699 ( P3_R1200_U28 , P3_U3413 );
not NOT1_24700 ( P3_R1200_U29 , P3_U3395 );
not NOT1_24701 ( P3_R1200_U30 , P3_U3387 );
not NOT1_24702 ( P3_R1200_U31 , P3_U3077 );
not NOT1_24703 ( P3_R1200_U32 , P3_U3398 );
not NOT1_24704 ( P3_R1200_U33 , P3_U3067 );
nand NAND2_24705 ( P3_R1200_U34 , P3_U3067 , P3_R1200_U29 );
not NOT1_24706 ( P3_R1200_U35 , P3_U3063 );
not NOT1_24707 ( P3_R1200_U36 , P3_U3404 );
not NOT1_24708 ( P3_R1200_U37 , P3_U3407 );
not NOT1_24709 ( P3_R1200_U38 , P3_U3401 );
not NOT1_24710 ( P3_R1200_U39 , P3_U3410 );
not NOT1_24711 ( P3_R1200_U40 , P3_U3070 );
not NOT1_24712 ( P3_R1200_U41 , P3_U3066 );
not NOT1_24713 ( P3_R1200_U42 , P3_U3059 );
nand NAND2_24714 ( P3_R1200_U43 , P3_U3059 , P3_R1200_U38 );
nand NAND2_24715 ( P3_R1200_U44 , P3_R1200_U214 , P3_R1200_U212 );
not NOT1_24716 ( P3_R1200_U45 , P3_U3416 );
not NOT1_24717 ( P3_R1200_U46 , P3_U3082 );
nand NAND2_24718 ( P3_R1200_U47 , P3_R1200_U44 , P3_R1200_U215 );
nand NAND2_24719 ( P3_R1200_U48 , P3_R1200_U43 , P3_R1200_U229 );
nand NAND3_24720 ( P3_R1200_U49 , P3_R1200_U201 , P3_R1200_U185 , P3_R1200_U349 );
not NOT1_24721 ( P3_R1200_U50 , P3_U3901 );
not NOT1_24722 ( P3_R1200_U51 , P3_U3422 );
not NOT1_24723 ( P3_R1200_U52 , P3_U3419 );
not NOT1_24724 ( P3_R1200_U53 , P3_U3062 );
not NOT1_24725 ( P3_R1200_U54 , P3_U3061 );
nand NAND2_24726 ( P3_R1200_U55 , P3_U3082 , P3_R1200_U45 );
not NOT1_24727 ( P3_R1200_U56 , P3_U3425 );
not NOT1_24728 ( P3_R1200_U57 , P3_U3071 );
not NOT1_24729 ( P3_R1200_U58 , P3_U3428 );
not NOT1_24730 ( P3_R1200_U59 , P3_U3079 );
not NOT1_24731 ( P3_R1200_U60 , P3_U3437 );
not NOT1_24732 ( P3_R1200_U61 , P3_U3434 );
not NOT1_24733 ( P3_R1200_U62 , P3_U3431 );
not NOT1_24734 ( P3_R1200_U63 , P3_U3072 );
not NOT1_24735 ( P3_R1200_U64 , P3_U3073 );
not NOT1_24736 ( P3_R1200_U65 , P3_U3078 );
nand NAND2_24737 ( P3_R1200_U66 , P3_U3078 , P3_R1200_U62 );
not NOT1_24738 ( P3_R1200_U67 , P3_U3440 );
not NOT1_24739 ( P3_R1200_U68 , P3_U3068 );
not NOT1_24740 ( P3_R1200_U69 , P3_U3081 );
not NOT1_24741 ( P3_R1200_U70 , P3_U3445 );
not NOT1_24742 ( P3_R1200_U71 , P3_U3080 );
not NOT1_24743 ( P3_R1200_U72 , P3_U3907 );
not NOT1_24744 ( P3_R1200_U73 , P3_U3075 );
not NOT1_24745 ( P3_R1200_U74 , P3_U3904 );
not NOT1_24746 ( P3_R1200_U75 , P3_U3905 );
not NOT1_24747 ( P3_R1200_U76 , P3_U3906 );
not NOT1_24748 ( P3_R1200_U77 , P3_U3065 );
not NOT1_24749 ( P3_R1200_U78 , P3_U3060 );
not NOT1_24750 ( P3_R1200_U79 , P3_U3074 );
nand NAND2_24751 ( P3_R1200_U80 , P3_U3074 , P3_R1200_U76 );
not NOT1_24752 ( P3_R1200_U81 , P3_U3903 );
not NOT1_24753 ( P3_R1200_U82 , P3_U3064 );
not NOT1_24754 ( P3_R1200_U83 , P3_U3902 );
not NOT1_24755 ( P3_R1200_U84 , P3_U3057 );
not NOT1_24756 ( P3_R1200_U85 , P3_U3900 );
not NOT1_24757 ( P3_R1200_U86 , P3_U3056 );
nand NAND2_24758 ( P3_R1200_U87 , P3_U3056 , P3_R1200_U50 );
not NOT1_24759 ( P3_R1200_U88 , P3_U3052 );
not NOT1_24760 ( P3_R1200_U89 , P3_U3899 );
not NOT1_24761 ( P3_R1200_U90 , P3_U3053 );
nand NAND2_24762 ( P3_R1200_U91 , P3_R1200_U302 , P3_R1200_U301 );
nand NAND2_24763 ( P3_R1200_U92 , P3_R1200_U80 , P3_R1200_U316 );
nand NAND2_24764 ( P3_R1200_U93 , P3_R1200_U66 , P3_R1200_U327 );
nand NAND2_24765 ( P3_R1200_U94 , P3_R1200_U55 , P3_R1200_U338 );
not NOT1_24766 ( P3_R1200_U95 , P3_U3076 );
nand NAND2_24767 ( P3_R1200_U96 , P3_R1200_U402 , P3_R1200_U401 );
nand NAND2_24768 ( P3_R1200_U97 , P3_R1200_U416 , P3_R1200_U415 );
nand NAND2_24769 ( P3_R1200_U98 , P3_R1200_U421 , P3_R1200_U420 );
nand NAND2_24770 ( P3_R1200_U99 , P3_R1200_U437 , P3_R1200_U436 );
nand NAND2_24771 ( P3_R1200_U100 , P3_R1200_U442 , P3_R1200_U441 );
nand NAND2_24772 ( P3_R1200_U101 , P3_R1200_U447 , P3_R1200_U446 );
nand NAND2_24773 ( P3_R1200_U102 , P3_R1200_U452 , P3_R1200_U451 );
nand NAND2_24774 ( P3_R1200_U103 , P3_R1200_U457 , P3_R1200_U456 );
nand NAND2_24775 ( P3_R1200_U104 , P3_R1200_U473 , P3_R1200_U472 );
nand NAND2_24776 ( P3_R1200_U105 , P3_R1200_U478 , P3_R1200_U477 );
nand NAND2_24777 ( P3_R1200_U106 , P3_R1200_U361 , P3_R1200_U360 );
nand NAND2_24778 ( P3_R1200_U107 , P3_R1200_U370 , P3_R1200_U369 );
nand NAND2_24779 ( P3_R1200_U108 , P3_R1200_U377 , P3_R1200_U376 );
nand NAND2_24780 ( P3_R1200_U109 , P3_R1200_U381 , P3_R1200_U380 );
nand NAND2_24781 ( P3_R1200_U110 , P3_R1200_U390 , P3_R1200_U389 );
nand NAND2_24782 ( P3_R1200_U111 , P3_R1200_U411 , P3_R1200_U410 );
nand NAND2_24783 ( P3_R1200_U112 , P3_R1200_U428 , P3_R1200_U427 );
nand NAND2_24784 ( P3_R1200_U113 , P3_R1200_U432 , P3_R1200_U431 );
nand NAND2_24785 ( P3_R1200_U114 , P3_R1200_U464 , P3_R1200_U463 );
nand NAND2_24786 ( P3_R1200_U115 , P3_R1200_U468 , P3_R1200_U467 );
nand NAND2_24787 ( P3_R1200_U116 , P3_R1200_U485 , P3_R1200_U484 );
and AND2_24788 ( P3_R1200_U117 , P3_R1200_U352 , P3_R1200_U193 );
and AND2_24789 ( P3_R1200_U118 , P3_R1200_U205 , P3_R1200_U206 );
and AND2_24790 ( P3_R1200_U119 , P3_R1200_U14 , P3_R1200_U13 );
and AND2_24791 ( P3_R1200_U120 , P3_R1200_U357 , P3_R1200_U354 );
and AND3_24792 ( P3_R1200_U121 , P3_R1200_U363 , P3_R1200_U362 , P3_R1200_U26 );
and AND2_24793 ( P3_R1200_U122 , P3_R1200_U366 , P3_R1200_U195 );
and AND2_24794 ( P3_R1200_U123 , P3_R1200_U235 , P3_R1200_U6 );
and AND2_24795 ( P3_R1200_U124 , P3_R1200_U373 , P3_R1200_U194 );
and AND3_24796 ( P3_R1200_U125 , P3_R1200_U383 , P3_R1200_U382 , P3_R1200_U34 );
and AND2_24797 ( P3_R1200_U126 , P3_R1200_U386 , P3_R1200_U193 );
and AND2_24798 ( P3_R1200_U127 , P3_R1200_U222 , P3_R1200_U7 );
and AND2_24799 ( P3_R1200_U128 , P3_R1200_U267 , P3_R1200_U9 );
and AND2_24800 ( P3_R1200_U129 , P3_R1200_U291 , P3_R1200_U11 );
and AND2_24801 ( P3_R1200_U130 , P3_R1200_U355 , P3_R1200_U192 );
and AND2_24802 ( P3_R1200_U131 , P3_R1200_U306 , P3_R1200_U307 );
and AND2_24803 ( P3_R1200_U132 , P3_R1200_U309 , P3_R1200_U395 );
and AND2_24804 ( P3_R1200_U133 , P3_R1200_U306 , P3_R1200_U307 );
and AND2_24805 ( P3_R1200_U134 , P3_R1200_U15 , P3_R1200_U310 );
nand NAND2_24806 ( P3_R1200_U135 , P3_R1200_U399 , P3_R1200_U398 );
and AND3_24807 ( P3_R1200_U136 , P3_R1200_U404 , P3_R1200_U403 , P3_R1200_U87 );
and AND2_24808 ( P3_R1200_U137 , P3_R1200_U407 , P3_R1200_U192 );
nand NAND2_24809 ( P3_R1200_U138 , P3_R1200_U413 , P3_R1200_U412 );
nand NAND2_24810 ( P3_R1200_U139 , P3_R1200_U418 , P3_R1200_U417 );
and AND2_24811 ( P3_R1200_U140 , P3_R1200_U322 , P3_R1200_U12 );
and AND2_24812 ( P3_R1200_U141 , P3_R1200_U424 , P3_R1200_U191 );
nand NAND2_24813 ( P3_R1200_U142 , P3_R1200_U434 , P3_R1200_U433 );
nand NAND2_24814 ( P3_R1200_U143 , P3_R1200_U439 , P3_R1200_U438 );
nand NAND2_24815 ( P3_R1200_U144 , P3_R1200_U444 , P3_R1200_U443 );
nand NAND2_24816 ( P3_R1200_U145 , P3_R1200_U449 , P3_R1200_U448 );
nand NAND2_24817 ( P3_R1200_U146 , P3_R1200_U454 , P3_R1200_U453 );
and AND2_24818 ( P3_R1200_U147 , P3_R1200_U333 , P3_R1200_U10 );
and AND2_24819 ( P3_R1200_U148 , P3_R1200_U460 , P3_R1200_U190 );
nand NAND2_24820 ( P3_R1200_U149 , P3_R1200_U470 , P3_R1200_U469 );
nand NAND2_24821 ( P3_R1200_U150 , P3_R1200_U475 , P3_R1200_U474 );
and AND2_24822 ( P3_R1200_U151 , P3_R1200_U344 , P3_R1200_U8 );
and AND2_24823 ( P3_R1200_U152 , P3_R1200_U481 , P3_R1200_U189 );
and AND2_24824 ( P3_R1200_U153 , P3_R1200_U359 , P3_R1200_U358 );
nand NAND2_24825 ( P3_R1200_U154 , P3_R1200_U120 , P3_R1200_U356 );
and AND2_24826 ( P3_R1200_U155 , P3_R1200_U368 , P3_R1200_U367 );
and AND2_24827 ( P3_R1200_U156 , P3_R1200_U375 , P3_R1200_U374 );
and AND2_24828 ( P3_R1200_U157 , P3_R1200_U379 , P3_R1200_U378 );
nand NAND2_24829 ( P3_R1200_U158 , P3_R1200_U118 , P3_R1200_U203 );
and AND2_24830 ( P3_R1200_U159 , P3_R1200_U388 , P3_R1200_U387 );
not NOT1_24831 ( P3_R1200_U160 , P3_U3908 );
not NOT1_24832 ( P3_R1200_U161 , P3_U3054 );
and AND2_24833 ( P3_R1200_U162 , P3_R1200_U397 , P3_R1200_U396 );
nand NAND2_24834 ( P3_R1200_U163 , P3_R1200_U131 , P3_R1200_U304 );
and AND2_24835 ( P3_R1200_U164 , P3_R1200_U409 , P3_R1200_U408 );
nand NAND2_24836 ( P3_R1200_U165 , P3_R1200_U298 , P3_R1200_U297 );
nand NAND2_24837 ( P3_R1200_U166 , P3_R1200_U294 , P3_R1200_U293 );
and AND2_24838 ( P3_R1200_U167 , P3_R1200_U426 , P3_R1200_U425 );
and AND2_24839 ( P3_R1200_U168 , P3_R1200_U430 , P3_R1200_U429 );
nand NAND2_24840 ( P3_R1200_U169 , P3_R1200_U284 , P3_R1200_U283 );
nand NAND2_24841 ( P3_R1200_U170 , P3_R1200_U280 , P3_R1200_U279 );
not NOT1_24842 ( P3_R1200_U171 , P3_U3392 );
nand NAND2_24843 ( P3_R1200_U172 , P3_U3387 , P3_R1200_U95 );
nand NAND3_24844 ( P3_R1200_U173 , P3_R1200_U276 , P3_R1200_U184 , P3_R1200_U350 );
not NOT1_24845 ( P3_R1200_U174 , P3_U3443 );
nand NAND2_24846 ( P3_R1200_U175 , P3_R1200_U274 , P3_R1200_U273 );
nand NAND2_24847 ( P3_R1200_U176 , P3_R1200_U270 , P3_R1200_U269 );
and AND2_24848 ( P3_R1200_U177 , P3_R1200_U462 , P3_R1200_U461 );
and AND2_24849 ( P3_R1200_U178 , P3_R1200_U466 , P3_R1200_U465 );
nand NAND2_24850 ( P3_R1200_U179 , P3_R1200_U260 , P3_R1200_U259 );
nand NAND2_24851 ( P3_R1200_U180 , P3_R1200_U256 , P3_R1200_U255 );
nand NAND2_24852 ( P3_R1200_U181 , P3_R1200_U252 , P3_R1200_U251 );
and AND2_24853 ( P3_R1200_U182 , P3_R1200_U483 , P3_R1200_U482 );
nand NAND2_24854 ( P3_R1200_U183 , P3_R1200_U132 , P3_R1200_U163 );
nand NAND2_24855 ( P3_R1200_U184 , P3_R1200_U175 , P3_R1200_U174 );
nand NAND2_24856 ( P3_R1200_U185 , P3_R1200_U172 , P3_R1200_U171 );
not NOT1_24857 ( P3_R1200_U186 , P3_R1200_U87 );
not NOT1_24858 ( P3_R1200_U187 , P3_R1200_U34 );
not NOT1_24859 ( P3_R1200_U188 , P3_R1200_U26 );
nand NAND2_24860 ( P3_R1200_U189 , P3_U3419 , P3_R1200_U54 );
nand NAND2_24861 ( P3_R1200_U190 , P3_U3434 , P3_R1200_U64 );
nand NAND2_24862 ( P3_R1200_U191 , P3_U3905 , P3_R1200_U78 );
nand NAND2_24863 ( P3_R1200_U192 , P3_U3901 , P3_R1200_U86 );
nand NAND2_24864 ( P3_R1200_U193 , P3_U3395 , P3_R1200_U33 );
nand NAND2_24865 ( P3_R1200_U194 , P3_U3404 , P3_R1200_U41 );
nand NAND2_24866 ( P3_R1200_U195 , P3_U3410 , P3_R1200_U25 );
not NOT1_24867 ( P3_R1200_U196 , P3_R1200_U66 );
not NOT1_24868 ( P3_R1200_U197 , P3_R1200_U80 );
not NOT1_24869 ( P3_R1200_U198 , P3_R1200_U43 );
not NOT1_24870 ( P3_R1200_U199 , P3_R1200_U55 );
not NOT1_24871 ( P3_R1200_U200 , P3_R1200_U172 );
nand NAND2_24872 ( P3_R1200_U201 , P3_U3077 , P3_R1200_U172 );
not NOT1_24873 ( P3_R1200_U202 , P3_R1200_U49 );
nand NAND2_24874 ( P3_R1200_U203 , P3_R1200_U117 , P3_R1200_U49 );
nand NAND2_24875 ( P3_R1200_U204 , P3_R1200_U35 , P3_R1200_U34 );
nand NAND2_24876 ( P3_R1200_U205 , P3_R1200_U204 , P3_R1200_U32 );
nand NAND2_24877 ( P3_R1200_U206 , P3_U3063 , P3_R1200_U187 );
not NOT1_24878 ( P3_R1200_U207 , P3_R1200_U158 );
nand NAND2_24879 ( P3_R1200_U208 , P3_U3407 , P3_R1200_U40 );
nand NAND2_24880 ( P3_R1200_U209 , P3_U3070 , P3_R1200_U37 );
nand NAND2_24881 ( P3_R1200_U210 , P3_U3066 , P3_R1200_U36 );
nand NAND2_24882 ( P3_R1200_U211 , P3_R1200_U198 , P3_R1200_U194 );
nand NAND2_24883 ( P3_R1200_U212 , P3_R1200_U6 , P3_R1200_U211 );
nand NAND2_24884 ( P3_R1200_U213 , P3_U3401 , P3_R1200_U42 );
nand NAND2_24885 ( P3_R1200_U214 , P3_U3407 , P3_R1200_U40 );
nand NAND2_24886 ( P3_R1200_U215 , P3_R1200_U13 , P3_R1200_U158 );
not NOT1_24887 ( P3_R1200_U216 , P3_R1200_U44 );
not NOT1_24888 ( P3_R1200_U217 , P3_R1200_U47 );
nand NAND2_24889 ( P3_R1200_U218 , P3_U3413 , P3_R1200_U27 );
nand NAND2_24890 ( P3_R1200_U219 , P3_R1200_U27 , P3_R1200_U26 );
nand NAND2_24891 ( P3_R1200_U220 , P3_U3083 , P3_R1200_U188 );
not NOT1_24892 ( P3_R1200_U221 , P3_R1200_U154 );
nand NAND2_24893 ( P3_R1200_U222 , P3_U3416 , P3_R1200_U46 );
nand NAND2_24894 ( P3_R1200_U223 , P3_R1200_U222 , P3_R1200_U55 );
nand NAND2_24895 ( P3_R1200_U224 , P3_R1200_U217 , P3_R1200_U26 );
nand NAND2_24896 ( P3_R1200_U225 , P3_R1200_U122 , P3_R1200_U224 );
nand NAND2_24897 ( P3_R1200_U226 , P3_R1200_U47 , P3_R1200_U195 );
nand NAND2_24898 ( P3_R1200_U227 , P3_R1200_U121 , P3_R1200_U226 );
nand NAND2_24899 ( P3_R1200_U228 , P3_R1200_U26 , P3_R1200_U195 );
nand NAND2_24900 ( P3_R1200_U229 , P3_R1200_U213 , P3_R1200_U158 );
not NOT1_24901 ( P3_R1200_U230 , P3_R1200_U48 );
nand NAND2_24902 ( P3_R1200_U231 , P3_U3066 , P3_R1200_U36 );
nand NAND2_24903 ( P3_R1200_U232 , P3_R1200_U230 , P3_R1200_U231 );
nand NAND2_24904 ( P3_R1200_U233 , P3_R1200_U124 , P3_R1200_U232 );
nand NAND2_24905 ( P3_R1200_U234 , P3_R1200_U48 , P3_R1200_U194 );
nand NAND2_24906 ( P3_R1200_U235 , P3_U3407 , P3_R1200_U40 );
nand NAND2_24907 ( P3_R1200_U236 , P3_R1200_U123 , P3_R1200_U234 );
nand NAND2_24908 ( P3_R1200_U237 , P3_U3066 , P3_R1200_U36 );
nand NAND2_24909 ( P3_R1200_U238 , P3_R1200_U194 , P3_R1200_U237 );
nand NAND2_24910 ( P3_R1200_U239 , P3_R1200_U213 , P3_R1200_U43 );
nand NAND2_24911 ( P3_R1200_U240 , P3_R1200_U202 , P3_R1200_U34 );
nand NAND2_24912 ( P3_R1200_U241 , P3_R1200_U126 , P3_R1200_U240 );
nand NAND2_24913 ( P3_R1200_U242 , P3_R1200_U49 , P3_R1200_U193 );
nand NAND2_24914 ( P3_R1200_U243 , P3_R1200_U125 , P3_R1200_U242 );
nand NAND2_24915 ( P3_R1200_U244 , P3_R1200_U193 , P3_R1200_U34 );
nand NAND2_24916 ( P3_R1200_U245 , P3_U3422 , P3_R1200_U53 );
nand NAND2_24917 ( P3_R1200_U246 , P3_U3062 , P3_R1200_U51 );
nand NAND2_24918 ( P3_R1200_U247 , P3_U3061 , P3_R1200_U52 );
nand NAND2_24919 ( P3_R1200_U248 , P3_R1200_U199 , P3_R1200_U7 );
nand NAND2_24920 ( P3_R1200_U249 , P3_R1200_U8 , P3_R1200_U248 );
nand NAND2_24921 ( P3_R1200_U250 , P3_U3422 , P3_R1200_U53 );
nand NAND2_24922 ( P3_R1200_U251 , P3_R1200_U127 , P3_R1200_U154 );
nand NAND2_24923 ( P3_R1200_U252 , P3_R1200_U250 , P3_R1200_U249 );
not NOT1_24924 ( P3_R1200_U253 , P3_R1200_U181 );
nand NAND2_24925 ( P3_R1200_U254 , P3_U3425 , P3_R1200_U57 );
nand NAND2_24926 ( P3_R1200_U255 , P3_R1200_U254 , P3_R1200_U181 );
nand NAND2_24927 ( P3_R1200_U256 , P3_U3071 , P3_R1200_U56 );
not NOT1_24928 ( P3_R1200_U257 , P3_R1200_U180 );
nand NAND2_24929 ( P3_R1200_U258 , P3_U3428 , P3_R1200_U59 );
nand NAND2_24930 ( P3_R1200_U259 , P3_R1200_U258 , P3_R1200_U180 );
nand NAND2_24931 ( P3_R1200_U260 , P3_U3079 , P3_R1200_U58 );
not NOT1_24932 ( P3_R1200_U261 , P3_R1200_U179 );
nand NAND2_24933 ( P3_R1200_U262 , P3_U3437 , P3_R1200_U63 );
nand NAND2_24934 ( P3_R1200_U263 , P3_U3072 , P3_R1200_U60 );
nand NAND2_24935 ( P3_R1200_U264 , P3_U3073 , P3_R1200_U61 );
nand NAND2_24936 ( P3_R1200_U265 , P3_R1200_U196 , P3_R1200_U9 );
nand NAND2_24937 ( P3_R1200_U266 , P3_R1200_U10 , P3_R1200_U265 );
nand NAND2_24938 ( P3_R1200_U267 , P3_U3431 , P3_R1200_U65 );
nand NAND2_24939 ( P3_R1200_U268 , P3_U3437 , P3_R1200_U63 );
nand NAND2_24940 ( P3_R1200_U269 , P3_R1200_U128 , P3_R1200_U179 );
nand NAND2_24941 ( P3_R1200_U270 , P3_R1200_U268 , P3_R1200_U266 );
not NOT1_24942 ( P3_R1200_U271 , P3_R1200_U176 );
nand NAND2_24943 ( P3_R1200_U272 , P3_U3440 , P3_R1200_U68 );
nand NAND2_24944 ( P3_R1200_U273 , P3_R1200_U272 , P3_R1200_U176 );
nand NAND2_24945 ( P3_R1200_U274 , P3_U3068 , P3_R1200_U67 );
not NOT1_24946 ( P3_R1200_U275 , P3_R1200_U175 );
nand NAND2_24947 ( P3_R1200_U276 , P3_U3081 , P3_R1200_U175 );
not NOT1_24948 ( P3_R1200_U277 , P3_R1200_U173 );
nand NAND2_24949 ( P3_R1200_U278 , P3_U3445 , P3_R1200_U71 );
nand NAND2_24950 ( P3_R1200_U279 , P3_R1200_U278 , P3_R1200_U173 );
nand NAND2_24951 ( P3_R1200_U280 , P3_U3080 , P3_R1200_U70 );
not NOT1_24952 ( P3_R1200_U281 , P3_R1200_U170 );
nand NAND2_24953 ( P3_R1200_U282 , P3_U3907 , P3_R1200_U73 );
nand NAND2_24954 ( P3_R1200_U283 , P3_R1200_U282 , P3_R1200_U170 );
nand NAND2_24955 ( P3_R1200_U284 , P3_U3075 , P3_R1200_U72 );
not NOT1_24956 ( P3_R1200_U285 , P3_R1200_U169 );
nand NAND2_24957 ( P3_R1200_U286 , P3_U3904 , P3_R1200_U77 );
nand NAND2_24958 ( P3_R1200_U287 , P3_U3065 , P3_R1200_U74 );
nand NAND2_24959 ( P3_R1200_U288 , P3_U3060 , P3_R1200_U75 );
nand NAND2_24960 ( P3_R1200_U289 , P3_R1200_U197 , P3_R1200_U11 );
nand NAND2_24961 ( P3_R1200_U290 , P3_R1200_U12 , P3_R1200_U289 );
nand NAND2_24962 ( P3_R1200_U291 , P3_U3906 , P3_R1200_U79 );
nand NAND2_24963 ( P3_R1200_U292 , P3_U3904 , P3_R1200_U77 );
nand NAND2_24964 ( P3_R1200_U293 , P3_R1200_U129 , P3_R1200_U169 );
nand NAND2_24965 ( P3_R1200_U294 , P3_R1200_U292 , P3_R1200_U290 );
not NOT1_24966 ( P3_R1200_U295 , P3_R1200_U166 );
nand NAND2_24967 ( P3_R1200_U296 , P3_U3903 , P3_R1200_U82 );
nand NAND2_24968 ( P3_R1200_U297 , P3_R1200_U296 , P3_R1200_U166 );
nand NAND2_24969 ( P3_R1200_U298 , P3_U3064 , P3_R1200_U81 );
not NOT1_24970 ( P3_R1200_U299 , P3_R1200_U165 );
nand NAND2_24971 ( P3_R1200_U300 , P3_U3902 , P3_R1200_U84 );
nand NAND2_24972 ( P3_R1200_U301 , P3_R1200_U300 , P3_R1200_U165 );
nand NAND2_24973 ( P3_R1200_U302 , P3_U3057 , P3_R1200_U83 );
not NOT1_24974 ( P3_R1200_U303 , P3_R1200_U91 );
nand NAND2_24975 ( P3_R1200_U304 , P3_R1200_U130 , P3_R1200_U91 );
nand NAND2_24976 ( P3_R1200_U305 , P3_R1200_U88 , P3_R1200_U87 );
nand NAND2_24977 ( P3_R1200_U306 , P3_R1200_U305 , P3_R1200_U85 );
nand NAND2_24978 ( P3_R1200_U307 , P3_U3052 , P3_R1200_U186 );
not NOT1_24979 ( P3_R1200_U308 , P3_R1200_U163 );
nand NAND2_24980 ( P3_R1200_U309 , P3_U3899 , P3_R1200_U90 );
nand NAND2_24981 ( P3_R1200_U310 , P3_U3053 , P3_R1200_U89 );
nand NAND2_24982 ( P3_R1200_U311 , P3_R1200_U303 , P3_R1200_U87 );
nand NAND2_24983 ( P3_R1200_U312 , P3_R1200_U137 , P3_R1200_U311 );
nand NAND2_24984 ( P3_R1200_U313 , P3_R1200_U91 , P3_R1200_U192 );
nand NAND2_24985 ( P3_R1200_U314 , P3_R1200_U136 , P3_R1200_U313 );
nand NAND2_24986 ( P3_R1200_U315 , P3_R1200_U192 , P3_R1200_U87 );
nand NAND2_24987 ( P3_R1200_U316 , P3_R1200_U291 , P3_R1200_U169 );
not NOT1_24988 ( P3_R1200_U317 , P3_R1200_U92 );
nand NAND2_24989 ( P3_R1200_U318 , P3_U3060 , P3_R1200_U75 );
nand NAND2_24990 ( P3_R1200_U319 , P3_R1200_U317 , P3_R1200_U318 );
nand NAND2_24991 ( P3_R1200_U320 , P3_R1200_U141 , P3_R1200_U319 );
nand NAND2_24992 ( P3_R1200_U321 , P3_R1200_U92 , P3_R1200_U191 );
nand NAND2_24993 ( P3_R1200_U322 , P3_U3904 , P3_R1200_U77 );
nand NAND2_24994 ( P3_R1200_U323 , P3_R1200_U140 , P3_R1200_U321 );
nand NAND2_24995 ( P3_R1200_U324 , P3_U3060 , P3_R1200_U75 );
nand NAND2_24996 ( P3_R1200_U325 , P3_R1200_U191 , P3_R1200_U324 );
nand NAND2_24997 ( P3_R1200_U326 , P3_R1200_U291 , P3_R1200_U80 );
nand NAND2_24998 ( P3_R1200_U327 , P3_R1200_U267 , P3_R1200_U179 );
not NOT1_24999 ( P3_R1200_U328 , P3_R1200_U93 );
nand NAND2_25000 ( P3_R1200_U329 , P3_U3073 , P3_R1200_U61 );
nand NAND2_25001 ( P3_R1200_U330 , P3_R1200_U328 , P3_R1200_U329 );
nand NAND2_25002 ( P3_R1200_U331 , P3_R1200_U148 , P3_R1200_U330 );
nand NAND2_25003 ( P3_R1200_U332 , P3_R1200_U93 , P3_R1200_U190 );
nand NAND2_25004 ( P3_R1200_U333 , P3_U3437 , P3_R1200_U63 );
nand NAND2_25005 ( P3_R1200_U334 , P3_R1200_U147 , P3_R1200_U332 );
nand NAND2_25006 ( P3_R1200_U335 , P3_U3073 , P3_R1200_U61 );
nand NAND2_25007 ( P3_R1200_U336 , P3_R1200_U190 , P3_R1200_U335 );
nand NAND2_25008 ( P3_R1200_U337 , P3_R1200_U267 , P3_R1200_U66 );
nand NAND2_25009 ( P3_R1200_U338 , P3_R1200_U222 , P3_R1200_U154 );
not NOT1_25010 ( P3_R1200_U339 , P3_R1200_U94 );
nand NAND2_25011 ( P3_R1200_U340 , P3_U3061 , P3_R1200_U52 );
nand NAND2_25012 ( P3_R1200_U341 , P3_R1200_U339 , P3_R1200_U340 );
nand NAND2_25013 ( P3_R1200_U342 , P3_R1200_U152 , P3_R1200_U341 );
nand NAND2_25014 ( P3_R1200_U343 , P3_R1200_U94 , P3_R1200_U189 );
nand NAND2_25015 ( P3_R1200_U344 , P3_U3422 , P3_R1200_U53 );
nand NAND2_25016 ( P3_R1200_U345 , P3_R1200_U151 , P3_R1200_U343 );
nand NAND2_25017 ( P3_R1200_U346 , P3_U3061 , P3_R1200_U52 );
nand NAND2_25018 ( P3_R1200_U347 , P3_R1200_U189 , P3_R1200_U346 );
nand NAND2_25019 ( P3_R1200_U348 , P3_U3076 , P3_R1200_U30 );
nand NAND2_25020 ( P3_R1200_U349 , P3_U3077 , P3_R1200_U171 );
nand NAND2_25021 ( P3_R1200_U350 , P3_U3081 , P3_R1200_U174 );
nand NAND3_25022 ( P3_R1200_U351 , P3_R1200_U133 , P3_R1200_U304 , P3_R1200_U134 );
nand NAND2_25023 ( P3_R1200_U352 , P3_U3398 , P3_R1200_U35 );
nand NAND2_25024 ( P3_R1200_U353 , P3_U3413 , P3_R1200_U220 );
nand NAND2_25025 ( P3_R1200_U354 , P3_R1200_U353 , P3_R1200_U219 );
nand NAND2_25026 ( P3_R1200_U355 , P3_U3900 , P3_R1200_U88 );
nand NAND2_25027 ( P3_R1200_U356 , P3_R1200_U119 , P3_R1200_U158 );
nand NAND2_25028 ( P3_R1200_U357 , P3_R1200_U216 , P3_R1200_U14 );
nand NAND2_25029 ( P3_R1200_U358 , P3_U3416 , P3_R1200_U46 );
nand NAND2_25030 ( P3_R1200_U359 , P3_U3082 , P3_R1200_U45 );
nand NAND2_25031 ( P3_R1200_U360 , P3_R1200_U223 , P3_R1200_U154 );
nand NAND2_25032 ( P3_R1200_U361 , P3_R1200_U221 , P3_R1200_U153 );
nand NAND2_25033 ( P3_R1200_U362 , P3_U3413 , P3_R1200_U27 );
nand NAND2_25034 ( P3_R1200_U363 , P3_U3083 , P3_R1200_U28 );
nand NAND2_25035 ( P3_R1200_U364 , P3_U3413 , P3_R1200_U27 );
nand NAND2_25036 ( P3_R1200_U365 , P3_U3083 , P3_R1200_U28 );
nand NAND2_25037 ( P3_R1200_U366 , P3_R1200_U365 , P3_R1200_U364 );
nand NAND2_25038 ( P3_R1200_U367 , P3_U3410 , P3_R1200_U25 );
nand NAND2_25039 ( P3_R1200_U368 , P3_U3069 , P3_R1200_U39 );
nand NAND2_25040 ( P3_R1200_U369 , P3_R1200_U228 , P3_R1200_U47 );
nand NAND2_25041 ( P3_R1200_U370 , P3_R1200_U155 , P3_R1200_U217 );
nand NAND2_25042 ( P3_R1200_U371 , P3_U3407 , P3_R1200_U40 );
nand NAND2_25043 ( P3_R1200_U372 , P3_U3070 , P3_R1200_U37 );
nand NAND2_25044 ( P3_R1200_U373 , P3_R1200_U372 , P3_R1200_U371 );
nand NAND2_25045 ( P3_R1200_U374 , P3_U3404 , P3_R1200_U41 );
nand NAND2_25046 ( P3_R1200_U375 , P3_U3066 , P3_R1200_U36 );
nand NAND2_25047 ( P3_R1200_U376 , P3_R1200_U238 , P3_R1200_U48 );
nand NAND2_25048 ( P3_R1200_U377 , P3_R1200_U156 , P3_R1200_U230 );
nand NAND2_25049 ( P3_R1200_U378 , P3_U3401 , P3_R1200_U42 );
nand NAND2_25050 ( P3_R1200_U379 , P3_U3059 , P3_R1200_U38 );
nand NAND2_25051 ( P3_R1200_U380 , P3_R1200_U239 , P3_R1200_U158 );
nand NAND2_25052 ( P3_R1200_U381 , P3_R1200_U207 , P3_R1200_U157 );
nand NAND2_25053 ( P3_R1200_U382 , P3_U3398 , P3_R1200_U35 );
nand NAND2_25054 ( P3_R1200_U383 , P3_U3063 , P3_R1200_U32 );
nand NAND2_25055 ( P3_R1200_U384 , P3_U3398 , P3_R1200_U35 );
nand NAND2_25056 ( P3_R1200_U385 , P3_U3063 , P3_R1200_U32 );
nand NAND2_25057 ( P3_R1200_U386 , P3_R1200_U385 , P3_R1200_U384 );
nand NAND2_25058 ( P3_R1200_U387 , P3_U3395 , P3_R1200_U33 );
nand NAND2_25059 ( P3_R1200_U388 , P3_U3067 , P3_R1200_U29 );
nand NAND2_25060 ( P3_R1200_U389 , P3_R1200_U244 , P3_R1200_U49 );
nand NAND2_25061 ( P3_R1200_U390 , P3_R1200_U159 , P3_R1200_U202 );
nand NAND2_25062 ( P3_R1200_U391 , P3_U3908 , P3_R1200_U161 );
nand NAND2_25063 ( P3_R1200_U392 , P3_U3054 , P3_R1200_U160 );
nand NAND2_25064 ( P3_R1200_U393 , P3_U3908 , P3_R1200_U161 );
nand NAND2_25065 ( P3_R1200_U394 , P3_U3054 , P3_R1200_U160 );
nand NAND2_25066 ( P3_R1200_U395 , P3_R1200_U394 , P3_R1200_U393 );
nand NAND3_25067 ( P3_R1200_U396 , P3_U3053 , P3_R1200_U395 , P3_R1200_U89 );
nand NAND3_25068 ( P3_R1200_U397 , P3_R1200_U15 , P3_R1200_U90 , P3_U3899 );
nand NAND2_25069 ( P3_R1200_U398 , P3_U3899 , P3_R1200_U90 );
nand NAND2_25070 ( P3_R1200_U399 , P3_U3053 , P3_R1200_U89 );
not NOT1_25071 ( P3_R1200_U400 , P3_R1200_U135 );
nand NAND2_25072 ( P3_R1200_U401 , P3_R1200_U308 , P3_R1200_U400 );
nand NAND2_25073 ( P3_R1200_U402 , P3_R1200_U135 , P3_R1200_U163 );
nand NAND2_25074 ( P3_R1200_U403 , P3_U3900 , P3_R1200_U88 );
nand NAND2_25075 ( P3_R1200_U404 , P3_U3052 , P3_R1200_U85 );
nand NAND2_25076 ( P3_R1200_U405 , P3_U3900 , P3_R1200_U88 );
nand NAND2_25077 ( P3_R1200_U406 , P3_U3052 , P3_R1200_U85 );
nand NAND2_25078 ( P3_R1200_U407 , P3_R1200_U406 , P3_R1200_U405 );
nand NAND2_25079 ( P3_R1200_U408 , P3_U3901 , P3_R1200_U86 );
nand NAND2_25080 ( P3_R1200_U409 , P3_U3056 , P3_R1200_U50 );
nand NAND2_25081 ( P3_R1200_U410 , P3_R1200_U315 , P3_R1200_U91 );
nand NAND2_25082 ( P3_R1200_U411 , P3_R1200_U164 , P3_R1200_U303 );
nand NAND2_25083 ( P3_R1200_U412 , P3_U3902 , P3_R1200_U84 );
nand NAND2_25084 ( P3_R1200_U413 , P3_U3057 , P3_R1200_U83 );
not NOT1_25085 ( P3_R1200_U414 , P3_R1200_U138 );
nand NAND2_25086 ( P3_R1200_U415 , P3_R1200_U299 , P3_R1200_U414 );
nand NAND2_25087 ( P3_R1200_U416 , P3_R1200_U138 , P3_R1200_U165 );
nand NAND2_25088 ( P3_R1200_U417 , P3_U3903 , P3_R1200_U82 );
nand NAND2_25089 ( P3_R1200_U418 , P3_U3064 , P3_R1200_U81 );
not NOT1_25090 ( P3_R1200_U419 , P3_R1200_U139 );
nand NAND2_25091 ( P3_R1200_U420 , P3_R1200_U295 , P3_R1200_U419 );
nand NAND2_25092 ( P3_R1200_U421 , P3_R1200_U139 , P3_R1200_U166 );
nand NAND2_25093 ( P3_R1200_U422 , P3_U3904 , P3_R1200_U77 );
nand NAND2_25094 ( P3_R1200_U423 , P3_U3065 , P3_R1200_U74 );
nand NAND2_25095 ( P3_R1200_U424 , P3_R1200_U423 , P3_R1200_U422 );
nand NAND2_25096 ( P3_R1200_U425 , P3_U3905 , P3_R1200_U78 );
nand NAND2_25097 ( P3_R1200_U426 , P3_U3060 , P3_R1200_U75 );
nand NAND2_25098 ( P3_R1200_U427 , P3_R1200_U325 , P3_R1200_U92 );
nand NAND2_25099 ( P3_R1200_U428 , P3_R1200_U167 , P3_R1200_U317 );
nand NAND2_25100 ( P3_R1200_U429 , P3_U3906 , P3_R1200_U79 );
nand NAND2_25101 ( P3_R1200_U430 , P3_U3074 , P3_R1200_U76 );
nand NAND2_25102 ( P3_R1200_U431 , P3_R1200_U326 , P3_R1200_U169 );
nand NAND2_25103 ( P3_R1200_U432 , P3_R1200_U285 , P3_R1200_U168 );
nand NAND2_25104 ( P3_R1200_U433 , P3_U3907 , P3_R1200_U73 );
nand NAND2_25105 ( P3_R1200_U434 , P3_U3075 , P3_R1200_U72 );
not NOT1_25106 ( P3_R1200_U435 , P3_R1200_U142 );
nand NAND2_25107 ( P3_R1200_U436 , P3_R1200_U281 , P3_R1200_U435 );
nand NAND2_25108 ( P3_R1200_U437 , P3_R1200_U142 , P3_R1200_U170 );
nand NAND2_25109 ( P3_R1200_U438 , P3_U3392 , P3_R1200_U31 );
nand NAND2_25110 ( P3_R1200_U439 , P3_U3077 , P3_R1200_U171 );
not NOT1_25111 ( P3_R1200_U440 , P3_R1200_U143 );
nand NAND2_25112 ( P3_R1200_U441 , P3_R1200_U200 , P3_R1200_U440 );
nand NAND2_25113 ( P3_R1200_U442 , P3_R1200_U143 , P3_R1200_U172 );
nand NAND2_25114 ( P3_R1200_U443 , P3_U3445 , P3_R1200_U71 );
nand NAND2_25115 ( P3_R1200_U444 , P3_U3080 , P3_R1200_U70 );
not NOT1_25116 ( P3_R1200_U445 , P3_R1200_U144 );
nand NAND2_25117 ( P3_R1200_U446 , P3_R1200_U277 , P3_R1200_U445 );
nand NAND2_25118 ( P3_R1200_U447 , P3_R1200_U144 , P3_R1200_U173 );
nand NAND2_25119 ( P3_R1200_U448 , P3_U3443 , P3_R1200_U69 );
nand NAND2_25120 ( P3_R1200_U449 , P3_U3081 , P3_R1200_U174 );
not NOT1_25121 ( P3_R1200_U450 , P3_R1200_U145 );
nand NAND2_25122 ( P3_R1200_U451 , P3_R1200_U275 , P3_R1200_U450 );
nand NAND2_25123 ( P3_R1200_U452 , P3_R1200_U145 , P3_R1200_U175 );
nand NAND2_25124 ( P3_R1200_U453 , P3_U3440 , P3_R1200_U68 );
nand NAND2_25125 ( P3_R1200_U454 , P3_U3068 , P3_R1200_U67 );
not NOT1_25126 ( P3_R1200_U455 , P3_R1200_U146 );
nand NAND2_25127 ( P3_R1200_U456 , P3_R1200_U271 , P3_R1200_U455 );
nand NAND2_25128 ( P3_R1200_U457 , P3_R1200_U146 , P3_R1200_U176 );
nand NAND2_25129 ( P3_R1200_U458 , P3_U3437 , P3_R1200_U63 );
nand NAND2_25130 ( P3_R1200_U459 , P3_U3072 , P3_R1200_U60 );
nand NAND2_25131 ( P3_R1200_U460 , P3_R1200_U459 , P3_R1200_U458 );
nand NAND2_25132 ( P3_R1200_U461 , P3_U3434 , P3_R1200_U64 );
nand NAND2_25133 ( P3_R1200_U462 , P3_U3073 , P3_R1200_U61 );
nand NAND2_25134 ( P3_R1200_U463 , P3_R1200_U336 , P3_R1200_U93 );
nand NAND2_25135 ( P3_R1200_U464 , P3_R1200_U177 , P3_R1200_U328 );
nand NAND2_25136 ( P3_R1200_U465 , P3_U3431 , P3_R1200_U65 );
nand NAND2_25137 ( P3_R1200_U466 , P3_U3078 , P3_R1200_U62 );
nand NAND2_25138 ( P3_R1200_U467 , P3_R1200_U337 , P3_R1200_U179 );
nand NAND2_25139 ( P3_R1200_U468 , P3_R1200_U261 , P3_R1200_U178 );
nand NAND2_25140 ( P3_R1200_U469 , P3_U3428 , P3_R1200_U59 );
nand NAND2_25141 ( P3_R1200_U470 , P3_U3079 , P3_R1200_U58 );
not NOT1_25142 ( P3_R1200_U471 , P3_R1200_U149 );
nand NAND2_25143 ( P3_R1200_U472 , P3_R1200_U257 , P3_R1200_U471 );
nand NAND2_25144 ( P3_R1200_U473 , P3_R1200_U149 , P3_R1200_U180 );
nand NAND2_25145 ( P3_R1200_U474 , P3_U3425 , P3_R1200_U57 );
nand NAND2_25146 ( P3_R1200_U475 , P3_U3071 , P3_R1200_U56 );
not NOT1_25147 ( P3_R1200_U476 , P3_R1200_U150 );
nand NAND2_25148 ( P3_R1200_U477 , P3_R1200_U253 , P3_R1200_U476 );
nand NAND2_25149 ( P3_R1200_U478 , P3_R1200_U150 , P3_R1200_U181 );
nand NAND2_25150 ( P3_R1200_U479 , P3_U3422 , P3_R1200_U53 );
nand NAND2_25151 ( P3_R1200_U480 , P3_U3062 , P3_R1200_U51 );
nand NAND2_25152 ( P3_R1200_U481 , P3_R1200_U480 , P3_R1200_U479 );
nand NAND2_25153 ( P3_R1200_U482 , P3_U3419 , P3_R1200_U54 );
nand NAND2_25154 ( P3_R1200_U483 , P3_U3061 , P3_R1200_U52 );
nand NAND2_25155 ( P3_R1200_U484 , P3_R1200_U347 , P3_R1200_U94 );
nand NAND2_25156 ( P3_R1200_U485 , P3_R1200_U182 , P3_R1200_U339 );
and AND2_25157 ( P3_R1179_U6 , P3_R1179_U210 , P3_R1179_U209 );
and AND2_25158 ( P3_R1179_U7 , P3_R1179_U189 , P3_R1179_U245 );
and AND2_25159 ( P3_R1179_U8 , P3_R1179_U247 , P3_R1179_U246 );
and AND2_25160 ( P3_R1179_U9 , P3_R1179_U190 , P3_R1179_U262 );
and AND2_25161 ( P3_R1179_U10 , P3_R1179_U264 , P3_R1179_U263 );
and AND2_25162 ( P3_R1179_U11 , P3_R1179_U191 , P3_R1179_U286 );
and AND2_25163 ( P3_R1179_U12 , P3_R1179_U288 , P3_R1179_U287 );
and AND3_25164 ( P3_R1179_U13 , P3_R1179_U208 , P3_R1179_U194 , P3_R1179_U213 );
and AND2_25165 ( P3_R1179_U14 , P3_R1179_U218 , P3_R1179_U195 );
and AND2_25166 ( P3_R1179_U15 , P3_R1179_U392 , P3_R1179_U391 );
nand NAND2_25167 ( P3_R1179_U16 , P3_R1179_U342 , P3_R1179_U345 );
nand NAND2_25168 ( P3_R1179_U17 , P3_R1179_U331 , P3_R1179_U334 );
nand NAND2_25169 ( P3_R1179_U18 , P3_R1179_U320 , P3_R1179_U323 );
nand NAND2_25170 ( P3_R1179_U19 , P3_R1179_U312 , P3_R1179_U314 );
nand NAND3_25171 ( P3_R1179_U20 , P3_R1179_U162 , P3_R1179_U183 , P3_R1179_U351 );
nand NAND2_25172 ( P3_R1179_U21 , P3_R1179_U241 , P3_R1179_U243 );
nand NAND2_25173 ( P3_R1179_U22 , P3_R1179_U233 , P3_R1179_U236 );
nand NAND2_25174 ( P3_R1179_U23 , P3_R1179_U225 , P3_R1179_U227 );
nand NAND2_25175 ( P3_R1179_U24 , P3_R1179_U172 , P3_R1179_U348 );
not NOT1_25176 ( P3_R1179_U25 , P3_U3069 );
nand NAND2_25177 ( P3_R1179_U26 , P3_U3069 , P3_R1179_U39 );
not NOT1_25178 ( P3_R1179_U27 , P3_U3083 );
not NOT1_25179 ( P3_R1179_U28 , P3_U3413 );
not NOT1_25180 ( P3_R1179_U29 , P3_U3395 );
not NOT1_25181 ( P3_R1179_U30 , P3_U3387 );
not NOT1_25182 ( P3_R1179_U31 , P3_U3077 );
not NOT1_25183 ( P3_R1179_U32 , P3_U3398 );
not NOT1_25184 ( P3_R1179_U33 , P3_U3067 );
nand NAND2_25185 ( P3_R1179_U34 , P3_U3067 , P3_R1179_U29 );
not NOT1_25186 ( P3_R1179_U35 , P3_U3063 );
not NOT1_25187 ( P3_R1179_U36 , P3_U3404 );
not NOT1_25188 ( P3_R1179_U37 , P3_U3407 );
not NOT1_25189 ( P3_R1179_U38 , P3_U3401 );
not NOT1_25190 ( P3_R1179_U39 , P3_U3410 );
not NOT1_25191 ( P3_R1179_U40 , P3_U3070 );
not NOT1_25192 ( P3_R1179_U41 , P3_U3066 );
not NOT1_25193 ( P3_R1179_U42 , P3_U3059 );
nand NAND2_25194 ( P3_R1179_U43 , P3_U3059 , P3_R1179_U38 );
nand NAND2_25195 ( P3_R1179_U44 , P3_R1179_U214 , P3_R1179_U212 );
not NOT1_25196 ( P3_R1179_U45 , P3_U3416 );
not NOT1_25197 ( P3_R1179_U46 , P3_U3082 );
nand NAND2_25198 ( P3_R1179_U47 , P3_R1179_U44 , P3_R1179_U215 );
nand NAND2_25199 ( P3_R1179_U48 , P3_R1179_U43 , P3_R1179_U229 );
nand NAND3_25200 ( P3_R1179_U49 , P3_R1179_U201 , P3_R1179_U185 , P3_R1179_U349 );
not NOT1_25201 ( P3_R1179_U50 , P3_U3901 );
not NOT1_25202 ( P3_R1179_U51 , P3_U3422 );
not NOT1_25203 ( P3_R1179_U52 , P3_U3419 );
not NOT1_25204 ( P3_R1179_U53 , P3_U3062 );
not NOT1_25205 ( P3_R1179_U54 , P3_U3061 );
nand NAND2_25206 ( P3_R1179_U55 , P3_U3082 , P3_R1179_U45 );
not NOT1_25207 ( P3_R1179_U56 , P3_U3425 );
not NOT1_25208 ( P3_R1179_U57 , P3_U3071 );
not NOT1_25209 ( P3_R1179_U58 , P3_U3428 );
not NOT1_25210 ( P3_R1179_U59 , P3_U3079 );
not NOT1_25211 ( P3_R1179_U60 , P3_U3437 );
not NOT1_25212 ( P3_R1179_U61 , P3_U3434 );
not NOT1_25213 ( P3_R1179_U62 , P3_U3431 );
not NOT1_25214 ( P3_R1179_U63 , P3_U3072 );
not NOT1_25215 ( P3_R1179_U64 , P3_U3073 );
not NOT1_25216 ( P3_R1179_U65 , P3_U3078 );
nand NAND2_25217 ( P3_R1179_U66 , P3_U3078 , P3_R1179_U62 );
not NOT1_25218 ( P3_R1179_U67 , P3_U3440 );
not NOT1_25219 ( P3_R1179_U68 , P3_U3068 );
not NOT1_25220 ( P3_R1179_U69 , P3_U3081 );
not NOT1_25221 ( P3_R1179_U70 , P3_U3445 );
not NOT1_25222 ( P3_R1179_U71 , P3_U3080 );
not NOT1_25223 ( P3_R1179_U72 , P3_U3907 );
not NOT1_25224 ( P3_R1179_U73 , P3_U3075 );
not NOT1_25225 ( P3_R1179_U74 , P3_U3904 );
not NOT1_25226 ( P3_R1179_U75 , P3_U3905 );
not NOT1_25227 ( P3_R1179_U76 , P3_U3906 );
not NOT1_25228 ( P3_R1179_U77 , P3_U3065 );
not NOT1_25229 ( P3_R1179_U78 , P3_U3060 );
not NOT1_25230 ( P3_R1179_U79 , P3_U3074 );
nand NAND2_25231 ( P3_R1179_U80 , P3_U3074 , P3_R1179_U76 );
not NOT1_25232 ( P3_R1179_U81 , P3_U3903 );
not NOT1_25233 ( P3_R1179_U82 , P3_U3064 );
not NOT1_25234 ( P3_R1179_U83 , P3_U3902 );
not NOT1_25235 ( P3_R1179_U84 , P3_U3057 );
not NOT1_25236 ( P3_R1179_U85 , P3_U3900 );
not NOT1_25237 ( P3_R1179_U86 , P3_U3056 );
nand NAND2_25238 ( P3_R1179_U87 , P3_U3056 , P3_R1179_U50 );
not NOT1_25239 ( P3_R1179_U88 , P3_U3052 );
not NOT1_25240 ( P3_R1179_U89 , P3_U3899 );
not NOT1_25241 ( P3_R1179_U90 , P3_U3053 );
nand NAND2_25242 ( P3_R1179_U91 , P3_R1179_U302 , P3_R1179_U301 );
nand NAND2_25243 ( P3_R1179_U92 , P3_R1179_U80 , P3_R1179_U316 );
nand NAND2_25244 ( P3_R1179_U93 , P3_R1179_U66 , P3_R1179_U327 );
nand NAND2_25245 ( P3_R1179_U94 , P3_R1179_U55 , P3_R1179_U338 );
not NOT1_25246 ( P3_R1179_U95 , P3_U3076 );
nand NAND2_25247 ( P3_R1179_U96 , P3_R1179_U402 , P3_R1179_U401 );
nand NAND2_25248 ( P3_R1179_U97 , P3_R1179_U416 , P3_R1179_U415 );
nand NAND2_25249 ( P3_R1179_U98 , P3_R1179_U421 , P3_R1179_U420 );
nand NAND2_25250 ( P3_R1179_U99 , P3_R1179_U437 , P3_R1179_U436 );
nand NAND2_25251 ( P3_R1179_U100 , P3_R1179_U442 , P3_R1179_U441 );
nand NAND2_25252 ( P3_R1179_U101 , P3_R1179_U447 , P3_R1179_U446 );
nand NAND2_25253 ( P3_R1179_U102 , P3_R1179_U452 , P3_R1179_U451 );
nand NAND2_25254 ( P3_R1179_U103 , P3_R1179_U457 , P3_R1179_U456 );
nand NAND2_25255 ( P3_R1179_U104 , P3_R1179_U473 , P3_R1179_U472 );
nand NAND2_25256 ( P3_R1179_U105 , P3_R1179_U478 , P3_R1179_U477 );
nand NAND2_25257 ( P3_R1179_U106 , P3_R1179_U361 , P3_R1179_U360 );
nand NAND2_25258 ( P3_R1179_U107 , P3_R1179_U370 , P3_R1179_U369 );
nand NAND2_25259 ( P3_R1179_U108 , P3_R1179_U377 , P3_R1179_U376 );
nand NAND2_25260 ( P3_R1179_U109 , P3_R1179_U381 , P3_R1179_U380 );
nand NAND2_25261 ( P3_R1179_U110 , P3_R1179_U390 , P3_R1179_U389 );
nand NAND2_25262 ( P3_R1179_U111 , P3_R1179_U411 , P3_R1179_U410 );
nand NAND2_25263 ( P3_R1179_U112 , P3_R1179_U428 , P3_R1179_U427 );
nand NAND2_25264 ( P3_R1179_U113 , P3_R1179_U432 , P3_R1179_U431 );
nand NAND2_25265 ( P3_R1179_U114 , P3_R1179_U464 , P3_R1179_U463 );
nand NAND2_25266 ( P3_R1179_U115 , P3_R1179_U468 , P3_R1179_U467 );
nand NAND2_25267 ( P3_R1179_U116 , P3_R1179_U485 , P3_R1179_U484 );
and AND2_25268 ( P3_R1179_U117 , P3_R1179_U352 , P3_R1179_U193 );
and AND2_25269 ( P3_R1179_U118 , P3_R1179_U205 , P3_R1179_U206 );
and AND2_25270 ( P3_R1179_U119 , P3_R1179_U14 , P3_R1179_U13 );
and AND2_25271 ( P3_R1179_U120 , P3_R1179_U357 , P3_R1179_U354 );
and AND3_25272 ( P3_R1179_U121 , P3_R1179_U363 , P3_R1179_U362 , P3_R1179_U26 );
and AND2_25273 ( P3_R1179_U122 , P3_R1179_U366 , P3_R1179_U195 );
and AND2_25274 ( P3_R1179_U123 , P3_R1179_U235 , P3_R1179_U6 );
and AND2_25275 ( P3_R1179_U124 , P3_R1179_U373 , P3_R1179_U194 );
and AND3_25276 ( P3_R1179_U125 , P3_R1179_U383 , P3_R1179_U382 , P3_R1179_U34 );
and AND2_25277 ( P3_R1179_U126 , P3_R1179_U386 , P3_R1179_U193 );
and AND2_25278 ( P3_R1179_U127 , P3_R1179_U222 , P3_R1179_U7 );
and AND2_25279 ( P3_R1179_U128 , P3_R1179_U267 , P3_R1179_U9 );
and AND2_25280 ( P3_R1179_U129 , P3_R1179_U291 , P3_R1179_U11 );
and AND2_25281 ( P3_R1179_U130 , P3_R1179_U355 , P3_R1179_U192 );
and AND2_25282 ( P3_R1179_U131 , P3_R1179_U306 , P3_R1179_U307 );
and AND2_25283 ( P3_R1179_U132 , P3_R1179_U309 , P3_R1179_U395 );
and AND2_25284 ( P3_R1179_U133 , P3_R1179_U306 , P3_R1179_U307 );
and AND2_25285 ( P3_R1179_U134 , P3_R1179_U15 , P3_R1179_U310 );
nand NAND2_25286 ( P3_R1179_U135 , P3_R1179_U399 , P3_R1179_U398 );
and AND3_25287 ( P3_R1179_U136 , P3_R1179_U404 , P3_R1179_U403 , P3_R1179_U87 );
and AND2_25288 ( P3_R1179_U137 , P3_R1179_U407 , P3_R1179_U192 );
nand NAND2_25289 ( P3_R1179_U138 , P3_R1179_U413 , P3_R1179_U412 );
nand NAND2_25290 ( P3_R1179_U139 , P3_R1179_U418 , P3_R1179_U417 );
and AND2_25291 ( P3_R1179_U140 , P3_R1179_U322 , P3_R1179_U12 );
and AND2_25292 ( P3_R1179_U141 , P3_R1179_U424 , P3_R1179_U191 );
nand NAND2_25293 ( P3_R1179_U142 , P3_R1179_U434 , P3_R1179_U433 );
nand NAND2_25294 ( P3_R1179_U143 , P3_R1179_U439 , P3_R1179_U438 );
nand NAND2_25295 ( P3_R1179_U144 , P3_R1179_U444 , P3_R1179_U443 );
nand NAND2_25296 ( P3_R1179_U145 , P3_R1179_U449 , P3_R1179_U448 );
nand NAND2_25297 ( P3_R1179_U146 , P3_R1179_U454 , P3_R1179_U453 );
and AND2_25298 ( P3_R1179_U147 , P3_R1179_U333 , P3_R1179_U10 );
and AND2_25299 ( P3_R1179_U148 , P3_R1179_U460 , P3_R1179_U190 );
nand NAND2_25300 ( P3_R1179_U149 , P3_R1179_U470 , P3_R1179_U469 );
nand NAND2_25301 ( P3_R1179_U150 , P3_R1179_U475 , P3_R1179_U474 );
and AND2_25302 ( P3_R1179_U151 , P3_R1179_U344 , P3_R1179_U8 );
and AND2_25303 ( P3_R1179_U152 , P3_R1179_U481 , P3_R1179_U189 );
and AND2_25304 ( P3_R1179_U153 , P3_R1179_U359 , P3_R1179_U358 );
nand NAND2_25305 ( P3_R1179_U154 , P3_R1179_U120 , P3_R1179_U356 );
and AND2_25306 ( P3_R1179_U155 , P3_R1179_U368 , P3_R1179_U367 );
and AND2_25307 ( P3_R1179_U156 , P3_R1179_U375 , P3_R1179_U374 );
and AND2_25308 ( P3_R1179_U157 , P3_R1179_U379 , P3_R1179_U378 );
nand NAND2_25309 ( P3_R1179_U158 , P3_R1179_U118 , P3_R1179_U203 );
and AND2_25310 ( P3_R1179_U159 , P3_R1179_U388 , P3_R1179_U387 );
not NOT1_25311 ( P3_R1179_U160 , P3_U3908 );
not NOT1_25312 ( P3_R1179_U161 , P3_U3054 );
and AND2_25313 ( P3_R1179_U162 , P3_R1179_U397 , P3_R1179_U396 );
nand NAND2_25314 ( P3_R1179_U163 , P3_R1179_U131 , P3_R1179_U304 );
and AND2_25315 ( P3_R1179_U164 , P3_R1179_U409 , P3_R1179_U408 );
nand NAND2_25316 ( P3_R1179_U165 , P3_R1179_U298 , P3_R1179_U297 );
nand NAND2_25317 ( P3_R1179_U166 , P3_R1179_U294 , P3_R1179_U293 );
and AND2_25318 ( P3_R1179_U167 , P3_R1179_U426 , P3_R1179_U425 );
and AND2_25319 ( P3_R1179_U168 , P3_R1179_U430 , P3_R1179_U429 );
nand NAND2_25320 ( P3_R1179_U169 , P3_R1179_U284 , P3_R1179_U283 );
nand NAND2_25321 ( P3_R1179_U170 , P3_R1179_U280 , P3_R1179_U279 );
not NOT1_25322 ( P3_R1179_U171 , P3_U3392 );
nand NAND2_25323 ( P3_R1179_U172 , P3_U3387 , P3_R1179_U95 );
nand NAND3_25324 ( P3_R1179_U173 , P3_R1179_U276 , P3_R1179_U184 , P3_R1179_U350 );
not NOT1_25325 ( P3_R1179_U174 , P3_U3443 );
nand NAND2_25326 ( P3_R1179_U175 , P3_R1179_U274 , P3_R1179_U273 );
nand NAND2_25327 ( P3_R1179_U176 , P3_R1179_U270 , P3_R1179_U269 );
and AND2_25328 ( P3_R1179_U177 , P3_R1179_U462 , P3_R1179_U461 );
and AND2_25329 ( P3_R1179_U178 , P3_R1179_U466 , P3_R1179_U465 );
nand NAND2_25330 ( P3_R1179_U179 , P3_R1179_U260 , P3_R1179_U259 );
nand NAND2_25331 ( P3_R1179_U180 , P3_R1179_U256 , P3_R1179_U255 );
nand NAND2_25332 ( P3_R1179_U181 , P3_R1179_U252 , P3_R1179_U251 );
and AND2_25333 ( P3_R1179_U182 , P3_R1179_U483 , P3_R1179_U482 );
nand NAND2_25334 ( P3_R1179_U183 , P3_R1179_U132 , P3_R1179_U163 );
nand NAND2_25335 ( P3_R1179_U184 , P3_R1179_U175 , P3_R1179_U174 );
nand NAND2_25336 ( P3_R1179_U185 , P3_R1179_U172 , P3_R1179_U171 );
not NOT1_25337 ( P3_R1179_U186 , P3_R1179_U87 );
not NOT1_25338 ( P3_R1179_U187 , P3_R1179_U34 );
not NOT1_25339 ( P3_R1179_U188 , P3_R1179_U26 );
nand NAND2_25340 ( P3_R1179_U189 , P3_U3419 , P3_R1179_U54 );
nand NAND2_25341 ( P3_R1179_U190 , P3_U3434 , P3_R1179_U64 );
nand NAND2_25342 ( P3_R1179_U191 , P3_U3905 , P3_R1179_U78 );
nand NAND2_25343 ( P3_R1179_U192 , P3_U3901 , P3_R1179_U86 );
nand NAND2_25344 ( P3_R1179_U193 , P3_U3395 , P3_R1179_U33 );
nand NAND2_25345 ( P3_R1179_U194 , P3_U3404 , P3_R1179_U41 );
nand NAND2_25346 ( P3_R1179_U195 , P3_U3410 , P3_R1179_U25 );
not NOT1_25347 ( P3_R1179_U196 , P3_R1179_U66 );
not NOT1_25348 ( P3_R1179_U197 , P3_R1179_U80 );
not NOT1_25349 ( P3_R1179_U198 , P3_R1179_U43 );
not NOT1_25350 ( P3_R1179_U199 , P3_R1179_U55 );
not NOT1_25351 ( P3_R1179_U200 , P3_R1179_U172 );
nand NAND2_25352 ( P3_R1179_U201 , P3_U3077 , P3_R1179_U172 );
not NOT1_25353 ( P3_R1179_U202 , P3_R1179_U49 );
nand NAND2_25354 ( P3_R1179_U203 , P3_R1179_U117 , P3_R1179_U49 );
nand NAND2_25355 ( P3_R1179_U204 , P3_R1179_U35 , P3_R1179_U34 );
nand NAND2_25356 ( P3_R1179_U205 , P3_R1179_U204 , P3_R1179_U32 );
nand NAND2_25357 ( P3_R1179_U206 , P3_U3063 , P3_R1179_U187 );
not NOT1_25358 ( P3_R1179_U207 , P3_R1179_U158 );
nand NAND2_25359 ( P3_R1179_U208 , P3_U3407 , P3_R1179_U40 );
nand NAND2_25360 ( P3_R1179_U209 , P3_U3070 , P3_R1179_U37 );
nand NAND2_25361 ( P3_R1179_U210 , P3_U3066 , P3_R1179_U36 );
nand NAND2_25362 ( P3_R1179_U211 , P3_R1179_U198 , P3_R1179_U194 );
nand NAND2_25363 ( P3_R1179_U212 , P3_R1179_U6 , P3_R1179_U211 );
nand NAND2_25364 ( P3_R1179_U213 , P3_U3401 , P3_R1179_U42 );
nand NAND2_25365 ( P3_R1179_U214 , P3_U3407 , P3_R1179_U40 );
nand NAND2_25366 ( P3_R1179_U215 , P3_R1179_U13 , P3_R1179_U158 );
not NOT1_25367 ( P3_R1179_U216 , P3_R1179_U44 );
not NOT1_25368 ( P3_R1179_U217 , P3_R1179_U47 );
nand NAND2_25369 ( P3_R1179_U218 , P3_U3413 , P3_R1179_U27 );
nand NAND2_25370 ( P3_R1179_U219 , P3_R1179_U27 , P3_R1179_U26 );
nand NAND2_25371 ( P3_R1179_U220 , P3_U3083 , P3_R1179_U188 );
not NOT1_25372 ( P3_R1179_U221 , P3_R1179_U154 );
nand NAND2_25373 ( P3_R1179_U222 , P3_U3416 , P3_R1179_U46 );
nand NAND2_25374 ( P3_R1179_U223 , P3_R1179_U222 , P3_R1179_U55 );
nand NAND2_25375 ( P3_R1179_U224 , P3_R1179_U217 , P3_R1179_U26 );
nand NAND2_25376 ( P3_R1179_U225 , P3_R1179_U122 , P3_R1179_U224 );
nand NAND2_25377 ( P3_R1179_U226 , P3_R1179_U47 , P3_R1179_U195 );
nand NAND2_25378 ( P3_R1179_U227 , P3_R1179_U121 , P3_R1179_U226 );
nand NAND2_25379 ( P3_R1179_U228 , P3_R1179_U26 , P3_R1179_U195 );
nand NAND2_25380 ( P3_R1179_U229 , P3_R1179_U213 , P3_R1179_U158 );
not NOT1_25381 ( P3_R1179_U230 , P3_R1179_U48 );
nand NAND2_25382 ( P3_R1179_U231 , P3_U3066 , P3_R1179_U36 );
nand NAND2_25383 ( P3_R1179_U232 , P3_R1179_U230 , P3_R1179_U231 );
nand NAND2_25384 ( P3_R1179_U233 , P3_R1179_U124 , P3_R1179_U232 );
nand NAND2_25385 ( P3_R1179_U234 , P3_R1179_U48 , P3_R1179_U194 );
nand NAND2_25386 ( P3_R1179_U235 , P3_U3407 , P3_R1179_U40 );
nand NAND2_25387 ( P3_R1179_U236 , P3_R1179_U123 , P3_R1179_U234 );
nand NAND2_25388 ( P3_R1179_U237 , P3_U3066 , P3_R1179_U36 );
nand NAND2_25389 ( P3_R1179_U238 , P3_R1179_U194 , P3_R1179_U237 );
nand NAND2_25390 ( P3_R1179_U239 , P3_R1179_U213 , P3_R1179_U43 );
nand NAND2_25391 ( P3_R1179_U240 , P3_R1179_U202 , P3_R1179_U34 );
nand NAND2_25392 ( P3_R1179_U241 , P3_R1179_U126 , P3_R1179_U240 );
nand NAND2_25393 ( P3_R1179_U242 , P3_R1179_U49 , P3_R1179_U193 );
nand NAND2_25394 ( P3_R1179_U243 , P3_R1179_U125 , P3_R1179_U242 );
nand NAND2_25395 ( P3_R1179_U244 , P3_R1179_U193 , P3_R1179_U34 );
nand NAND2_25396 ( P3_R1179_U245 , P3_U3422 , P3_R1179_U53 );
nand NAND2_25397 ( P3_R1179_U246 , P3_U3062 , P3_R1179_U51 );
nand NAND2_25398 ( P3_R1179_U247 , P3_U3061 , P3_R1179_U52 );
nand NAND2_25399 ( P3_R1179_U248 , P3_R1179_U199 , P3_R1179_U7 );
nand NAND2_25400 ( P3_R1179_U249 , P3_R1179_U8 , P3_R1179_U248 );
nand NAND2_25401 ( P3_R1179_U250 , P3_U3422 , P3_R1179_U53 );
nand NAND2_25402 ( P3_R1179_U251 , P3_R1179_U127 , P3_R1179_U154 );
nand NAND2_25403 ( P3_R1179_U252 , P3_R1179_U250 , P3_R1179_U249 );
not NOT1_25404 ( P3_R1179_U253 , P3_R1179_U181 );
nand NAND2_25405 ( P3_R1179_U254 , P3_U3425 , P3_R1179_U57 );
nand NAND2_25406 ( P3_R1179_U255 , P3_R1179_U254 , P3_R1179_U181 );
nand NAND2_25407 ( P3_R1179_U256 , P3_U3071 , P3_R1179_U56 );
not NOT1_25408 ( P3_R1179_U257 , P3_R1179_U180 );
nand NAND2_25409 ( P3_R1179_U258 , P3_U3428 , P3_R1179_U59 );
nand NAND2_25410 ( P3_R1179_U259 , P3_R1179_U258 , P3_R1179_U180 );
nand NAND2_25411 ( P3_R1179_U260 , P3_U3079 , P3_R1179_U58 );
not NOT1_25412 ( P3_R1179_U261 , P3_R1179_U179 );
nand NAND2_25413 ( P3_R1179_U262 , P3_U3437 , P3_R1179_U63 );
nand NAND2_25414 ( P3_R1179_U263 , P3_U3072 , P3_R1179_U60 );
nand NAND2_25415 ( P3_R1179_U264 , P3_U3073 , P3_R1179_U61 );
nand NAND2_25416 ( P3_R1179_U265 , P3_R1179_U196 , P3_R1179_U9 );
nand NAND2_25417 ( P3_R1179_U266 , P3_R1179_U10 , P3_R1179_U265 );
nand NAND2_25418 ( P3_R1179_U267 , P3_U3431 , P3_R1179_U65 );
nand NAND2_25419 ( P3_R1179_U268 , P3_U3437 , P3_R1179_U63 );
nand NAND2_25420 ( P3_R1179_U269 , P3_R1179_U128 , P3_R1179_U179 );
nand NAND2_25421 ( P3_R1179_U270 , P3_R1179_U268 , P3_R1179_U266 );
not NOT1_25422 ( P3_R1179_U271 , P3_R1179_U176 );
nand NAND2_25423 ( P3_R1179_U272 , P3_U3440 , P3_R1179_U68 );
nand NAND2_25424 ( P3_R1179_U273 , P3_R1179_U272 , P3_R1179_U176 );
nand NAND2_25425 ( P3_R1179_U274 , P3_U3068 , P3_R1179_U67 );
not NOT1_25426 ( P3_R1179_U275 , P3_R1179_U175 );
nand NAND2_25427 ( P3_R1179_U276 , P3_U3081 , P3_R1179_U175 );
not NOT1_25428 ( P3_R1179_U277 , P3_R1179_U173 );
nand NAND2_25429 ( P3_R1179_U278 , P3_U3445 , P3_R1179_U71 );
nand NAND2_25430 ( P3_R1179_U279 , P3_R1179_U278 , P3_R1179_U173 );
nand NAND2_25431 ( P3_R1179_U280 , P3_U3080 , P3_R1179_U70 );
not NOT1_25432 ( P3_R1179_U281 , P3_R1179_U170 );
nand NAND2_25433 ( P3_R1179_U282 , P3_U3907 , P3_R1179_U73 );
nand NAND2_25434 ( P3_R1179_U283 , P3_R1179_U282 , P3_R1179_U170 );
nand NAND2_25435 ( P3_R1179_U284 , P3_U3075 , P3_R1179_U72 );
not NOT1_25436 ( P3_R1179_U285 , P3_R1179_U169 );
nand NAND2_25437 ( P3_R1179_U286 , P3_U3904 , P3_R1179_U77 );
nand NAND2_25438 ( P3_R1179_U287 , P3_U3065 , P3_R1179_U74 );
nand NAND2_25439 ( P3_R1179_U288 , P3_U3060 , P3_R1179_U75 );
nand NAND2_25440 ( P3_R1179_U289 , P3_R1179_U197 , P3_R1179_U11 );
nand NAND2_25441 ( P3_R1179_U290 , P3_R1179_U12 , P3_R1179_U289 );
nand NAND2_25442 ( P3_R1179_U291 , P3_U3906 , P3_R1179_U79 );
nand NAND2_25443 ( P3_R1179_U292 , P3_U3904 , P3_R1179_U77 );
nand NAND2_25444 ( P3_R1179_U293 , P3_R1179_U129 , P3_R1179_U169 );
nand NAND2_25445 ( P3_R1179_U294 , P3_R1179_U292 , P3_R1179_U290 );
not NOT1_25446 ( P3_R1179_U295 , P3_R1179_U166 );
nand NAND2_25447 ( P3_R1179_U296 , P3_U3903 , P3_R1179_U82 );
nand NAND2_25448 ( P3_R1179_U297 , P3_R1179_U296 , P3_R1179_U166 );
nand NAND2_25449 ( P3_R1179_U298 , P3_U3064 , P3_R1179_U81 );
not NOT1_25450 ( P3_R1179_U299 , P3_R1179_U165 );
nand NAND2_25451 ( P3_R1179_U300 , P3_U3902 , P3_R1179_U84 );
nand NAND2_25452 ( P3_R1179_U301 , P3_R1179_U300 , P3_R1179_U165 );
nand NAND2_25453 ( P3_R1179_U302 , P3_U3057 , P3_R1179_U83 );
not NOT1_25454 ( P3_R1179_U303 , P3_R1179_U91 );
nand NAND2_25455 ( P3_R1179_U304 , P3_R1179_U130 , P3_R1179_U91 );
nand NAND2_25456 ( P3_R1179_U305 , P3_R1179_U88 , P3_R1179_U87 );
nand NAND2_25457 ( P3_R1179_U306 , P3_R1179_U305 , P3_R1179_U85 );
nand NAND2_25458 ( P3_R1179_U307 , P3_U3052 , P3_R1179_U186 );
not NOT1_25459 ( P3_R1179_U308 , P3_R1179_U163 );
nand NAND2_25460 ( P3_R1179_U309 , P3_U3899 , P3_R1179_U90 );
nand NAND2_25461 ( P3_R1179_U310 , P3_U3053 , P3_R1179_U89 );
nand NAND2_25462 ( P3_R1179_U311 , P3_R1179_U303 , P3_R1179_U87 );
nand NAND2_25463 ( P3_R1179_U312 , P3_R1179_U137 , P3_R1179_U311 );
nand NAND2_25464 ( P3_R1179_U313 , P3_R1179_U91 , P3_R1179_U192 );
nand NAND2_25465 ( P3_R1179_U314 , P3_R1179_U136 , P3_R1179_U313 );
nand NAND2_25466 ( P3_R1179_U315 , P3_R1179_U192 , P3_R1179_U87 );
nand NAND2_25467 ( P3_R1179_U316 , P3_R1179_U291 , P3_R1179_U169 );
not NOT1_25468 ( P3_R1179_U317 , P3_R1179_U92 );
nand NAND2_25469 ( P3_R1179_U318 , P3_U3060 , P3_R1179_U75 );
nand NAND2_25470 ( P3_R1179_U319 , P3_R1179_U317 , P3_R1179_U318 );
nand NAND2_25471 ( P3_R1179_U320 , P3_R1179_U141 , P3_R1179_U319 );
nand NAND2_25472 ( P3_R1179_U321 , P3_R1179_U92 , P3_R1179_U191 );
nand NAND2_25473 ( P3_R1179_U322 , P3_U3904 , P3_R1179_U77 );
nand NAND2_25474 ( P3_R1179_U323 , P3_R1179_U140 , P3_R1179_U321 );
nand NAND2_25475 ( P3_R1179_U324 , P3_U3060 , P3_R1179_U75 );
nand NAND2_25476 ( P3_R1179_U325 , P3_R1179_U191 , P3_R1179_U324 );
nand NAND2_25477 ( P3_R1179_U326 , P3_R1179_U291 , P3_R1179_U80 );
nand NAND2_25478 ( P3_R1179_U327 , P3_R1179_U267 , P3_R1179_U179 );
not NOT1_25479 ( P3_R1179_U328 , P3_R1179_U93 );
nand NAND2_25480 ( P3_R1179_U329 , P3_U3073 , P3_R1179_U61 );
nand NAND2_25481 ( P3_R1179_U330 , P3_R1179_U328 , P3_R1179_U329 );
nand NAND2_25482 ( P3_R1179_U331 , P3_R1179_U148 , P3_R1179_U330 );
nand NAND2_25483 ( P3_R1179_U332 , P3_R1179_U93 , P3_R1179_U190 );
nand NAND2_25484 ( P3_R1179_U333 , P3_U3437 , P3_R1179_U63 );
nand NAND2_25485 ( P3_R1179_U334 , P3_R1179_U147 , P3_R1179_U332 );
nand NAND2_25486 ( P3_R1179_U335 , P3_U3073 , P3_R1179_U61 );
nand NAND2_25487 ( P3_R1179_U336 , P3_R1179_U190 , P3_R1179_U335 );
nand NAND2_25488 ( P3_R1179_U337 , P3_R1179_U267 , P3_R1179_U66 );
nand NAND2_25489 ( P3_R1179_U338 , P3_R1179_U222 , P3_R1179_U154 );
not NOT1_25490 ( P3_R1179_U339 , P3_R1179_U94 );
nand NAND2_25491 ( P3_R1179_U340 , P3_U3061 , P3_R1179_U52 );
nand NAND2_25492 ( P3_R1179_U341 , P3_R1179_U339 , P3_R1179_U340 );
nand NAND2_25493 ( P3_R1179_U342 , P3_R1179_U152 , P3_R1179_U341 );
nand NAND2_25494 ( P3_R1179_U343 , P3_R1179_U94 , P3_R1179_U189 );
nand NAND2_25495 ( P3_R1179_U344 , P3_U3422 , P3_R1179_U53 );
nand NAND2_25496 ( P3_R1179_U345 , P3_R1179_U151 , P3_R1179_U343 );
nand NAND2_25497 ( P3_R1179_U346 , P3_U3061 , P3_R1179_U52 );
nand NAND2_25498 ( P3_R1179_U347 , P3_R1179_U189 , P3_R1179_U346 );
nand NAND2_25499 ( P3_R1179_U348 , P3_U3076 , P3_R1179_U30 );
nand NAND2_25500 ( P3_R1179_U349 , P3_U3077 , P3_R1179_U171 );
nand NAND2_25501 ( P3_R1179_U350 , P3_U3081 , P3_R1179_U174 );
nand NAND3_25502 ( P3_R1179_U351 , P3_R1179_U133 , P3_R1179_U304 , P3_R1179_U134 );
nand NAND2_25503 ( P3_R1179_U352 , P3_U3398 , P3_R1179_U35 );
nand NAND2_25504 ( P3_R1179_U353 , P3_U3413 , P3_R1179_U220 );
nand NAND2_25505 ( P3_R1179_U354 , P3_R1179_U353 , P3_R1179_U219 );
nand NAND2_25506 ( P3_R1179_U355 , P3_U3900 , P3_R1179_U88 );
nand NAND2_25507 ( P3_R1179_U356 , P3_R1179_U119 , P3_R1179_U158 );
nand NAND2_25508 ( P3_R1179_U357 , P3_R1179_U216 , P3_R1179_U14 );
nand NAND2_25509 ( P3_R1179_U358 , P3_U3416 , P3_R1179_U46 );
nand NAND2_25510 ( P3_R1179_U359 , P3_U3082 , P3_R1179_U45 );
nand NAND2_25511 ( P3_R1179_U360 , P3_R1179_U223 , P3_R1179_U154 );
nand NAND2_25512 ( P3_R1179_U361 , P3_R1179_U221 , P3_R1179_U153 );
nand NAND2_25513 ( P3_R1179_U362 , P3_U3413 , P3_R1179_U27 );
nand NAND2_25514 ( P3_R1179_U363 , P3_U3083 , P3_R1179_U28 );
nand NAND2_25515 ( P3_R1179_U364 , P3_U3413 , P3_R1179_U27 );
nand NAND2_25516 ( P3_R1179_U365 , P3_U3083 , P3_R1179_U28 );
nand NAND2_25517 ( P3_R1179_U366 , P3_R1179_U365 , P3_R1179_U364 );
nand NAND2_25518 ( P3_R1179_U367 , P3_U3410 , P3_R1179_U25 );
nand NAND2_25519 ( P3_R1179_U368 , P3_U3069 , P3_R1179_U39 );
nand NAND2_25520 ( P3_R1179_U369 , P3_R1179_U228 , P3_R1179_U47 );
nand NAND2_25521 ( P3_R1179_U370 , P3_R1179_U155 , P3_R1179_U217 );
nand NAND2_25522 ( P3_R1179_U371 , P3_U3407 , P3_R1179_U40 );
nand NAND2_25523 ( P3_R1179_U372 , P3_U3070 , P3_R1179_U37 );
nand NAND2_25524 ( P3_R1179_U373 , P3_R1179_U372 , P3_R1179_U371 );
nand NAND2_25525 ( P3_R1179_U374 , P3_U3404 , P3_R1179_U41 );
nand NAND2_25526 ( P3_R1179_U375 , P3_U3066 , P3_R1179_U36 );
nand NAND2_25527 ( P3_R1179_U376 , P3_R1179_U238 , P3_R1179_U48 );
nand NAND2_25528 ( P3_R1179_U377 , P3_R1179_U156 , P3_R1179_U230 );
nand NAND2_25529 ( P3_R1179_U378 , P3_U3401 , P3_R1179_U42 );
nand NAND2_25530 ( P3_R1179_U379 , P3_U3059 , P3_R1179_U38 );
nand NAND2_25531 ( P3_R1179_U380 , P3_R1179_U239 , P3_R1179_U158 );
nand NAND2_25532 ( P3_R1179_U381 , P3_R1179_U207 , P3_R1179_U157 );
nand NAND2_25533 ( P3_R1179_U382 , P3_U3398 , P3_R1179_U35 );
nand NAND2_25534 ( P3_R1179_U383 , P3_U3063 , P3_R1179_U32 );
nand NAND2_25535 ( P3_R1179_U384 , P3_U3398 , P3_R1179_U35 );
nand NAND2_25536 ( P3_R1179_U385 , P3_U3063 , P3_R1179_U32 );
nand NAND2_25537 ( P3_R1179_U386 , P3_R1179_U385 , P3_R1179_U384 );
nand NAND2_25538 ( P3_R1179_U387 , P3_U3395 , P3_R1179_U33 );
nand NAND2_25539 ( P3_R1179_U388 , P3_U3067 , P3_R1179_U29 );
nand NAND2_25540 ( P3_R1179_U389 , P3_R1179_U244 , P3_R1179_U49 );
nand NAND2_25541 ( P3_R1179_U390 , P3_R1179_U159 , P3_R1179_U202 );
nand NAND2_25542 ( P3_R1179_U391 , P3_U3908 , P3_R1179_U161 );
nand NAND2_25543 ( P3_R1179_U392 , P3_U3054 , P3_R1179_U160 );
nand NAND2_25544 ( P3_R1179_U393 , P3_U3908 , P3_R1179_U161 );
nand NAND2_25545 ( P3_R1179_U394 , P3_U3054 , P3_R1179_U160 );
nand NAND2_25546 ( P3_R1179_U395 , P3_R1179_U394 , P3_R1179_U393 );
nand NAND3_25547 ( P3_R1179_U396 , P3_U3053 , P3_R1179_U395 , P3_R1179_U89 );
nand NAND3_25548 ( P3_R1179_U397 , P3_R1179_U15 , P3_R1179_U90 , P3_U3899 );
nand NAND2_25549 ( P3_R1179_U398 , P3_U3899 , P3_R1179_U90 );
nand NAND2_25550 ( P3_R1179_U399 , P3_U3053 , P3_R1179_U89 );
not NOT1_25551 ( P3_R1179_U400 , P3_R1179_U135 );
nand NAND2_25552 ( P3_R1179_U401 , P3_R1179_U308 , P3_R1179_U400 );
nand NAND2_25553 ( P3_R1179_U402 , P3_R1179_U135 , P3_R1179_U163 );
nand NAND2_25554 ( P3_R1179_U403 , P3_U3900 , P3_R1179_U88 );
nand NAND2_25555 ( P3_R1179_U404 , P3_U3052 , P3_R1179_U85 );
nand NAND2_25556 ( P3_R1179_U405 , P3_U3900 , P3_R1179_U88 );
nand NAND2_25557 ( P3_R1179_U406 , P3_U3052 , P3_R1179_U85 );
nand NAND2_25558 ( P3_R1179_U407 , P3_R1179_U406 , P3_R1179_U405 );
nand NAND2_25559 ( P3_R1179_U408 , P3_U3901 , P3_R1179_U86 );
nand NAND2_25560 ( P3_R1179_U409 , P3_U3056 , P3_R1179_U50 );
nand NAND2_25561 ( P3_R1179_U410 , P3_R1179_U315 , P3_R1179_U91 );
nand NAND2_25562 ( P3_R1179_U411 , P3_R1179_U164 , P3_R1179_U303 );
nand NAND2_25563 ( P3_R1179_U412 , P3_U3902 , P3_R1179_U84 );
nand NAND2_25564 ( P3_R1179_U413 , P3_U3057 , P3_R1179_U83 );
not NOT1_25565 ( P3_R1179_U414 , P3_R1179_U138 );
nand NAND2_25566 ( P3_R1179_U415 , P3_R1179_U299 , P3_R1179_U414 );
nand NAND2_25567 ( P3_R1179_U416 , P3_R1179_U138 , P3_R1179_U165 );
nand NAND2_25568 ( P3_R1179_U417 , P3_U3903 , P3_R1179_U82 );
nand NAND2_25569 ( P3_R1179_U418 , P3_U3064 , P3_R1179_U81 );
not NOT1_25570 ( P3_R1179_U419 , P3_R1179_U139 );
nand NAND2_25571 ( P3_R1179_U420 , P3_R1179_U295 , P3_R1179_U419 );
nand NAND2_25572 ( P3_R1179_U421 , P3_R1179_U139 , P3_R1179_U166 );
nand NAND2_25573 ( P3_R1179_U422 , P3_U3904 , P3_R1179_U77 );
nand NAND2_25574 ( P3_R1179_U423 , P3_U3065 , P3_R1179_U74 );
nand NAND2_25575 ( P3_R1179_U424 , P3_R1179_U423 , P3_R1179_U422 );
nand NAND2_25576 ( P3_R1179_U425 , P3_U3905 , P3_R1179_U78 );
nand NAND2_25577 ( P3_R1179_U426 , P3_U3060 , P3_R1179_U75 );
nand NAND2_25578 ( P3_R1179_U427 , P3_R1179_U325 , P3_R1179_U92 );
nand NAND2_25579 ( P3_R1179_U428 , P3_R1179_U167 , P3_R1179_U317 );
nand NAND2_25580 ( P3_R1179_U429 , P3_U3906 , P3_R1179_U79 );
nand NAND2_25581 ( P3_R1179_U430 , P3_U3074 , P3_R1179_U76 );
nand NAND2_25582 ( P3_R1179_U431 , P3_R1179_U326 , P3_R1179_U169 );
nand NAND2_25583 ( P3_R1179_U432 , P3_R1179_U285 , P3_R1179_U168 );
nand NAND2_25584 ( P3_R1179_U433 , P3_U3907 , P3_R1179_U73 );
nand NAND2_25585 ( P3_R1179_U434 , P3_U3075 , P3_R1179_U72 );
not NOT1_25586 ( P3_R1179_U435 , P3_R1179_U142 );
nand NAND2_25587 ( P3_R1179_U436 , P3_R1179_U281 , P3_R1179_U435 );
nand NAND2_25588 ( P3_R1179_U437 , P3_R1179_U142 , P3_R1179_U170 );
nand NAND2_25589 ( P3_R1179_U438 , P3_U3392 , P3_R1179_U31 );
nand NAND2_25590 ( P3_R1179_U439 , P3_U3077 , P3_R1179_U171 );
not NOT1_25591 ( P3_R1179_U440 , P3_R1179_U143 );
nand NAND2_25592 ( P3_R1179_U441 , P3_R1179_U200 , P3_R1179_U440 );
nand NAND2_25593 ( P3_R1179_U442 , P3_R1179_U143 , P3_R1179_U172 );
nand NAND2_25594 ( P3_R1179_U443 , P3_U3445 , P3_R1179_U71 );
nand NAND2_25595 ( P3_R1179_U444 , P3_U3080 , P3_R1179_U70 );
not NOT1_25596 ( P3_R1179_U445 , P3_R1179_U144 );
nand NAND2_25597 ( P3_R1179_U446 , P3_R1179_U277 , P3_R1179_U445 );
nand NAND2_25598 ( P3_R1179_U447 , P3_R1179_U144 , P3_R1179_U173 );
nand NAND2_25599 ( P3_R1179_U448 , P3_U3443 , P3_R1179_U69 );
nand NAND2_25600 ( P3_R1179_U449 , P3_U3081 , P3_R1179_U174 );
not NOT1_25601 ( P3_R1179_U450 , P3_R1179_U145 );
nand NAND2_25602 ( P3_R1179_U451 , P3_R1179_U275 , P3_R1179_U450 );
nand NAND2_25603 ( P3_R1179_U452 , P3_R1179_U145 , P3_R1179_U175 );
nand NAND2_25604 ( P3_R1179_U453 , P3_U3440 , P3_R1179_U68 );
nand NAND2_25605 ( P3_R1179_U454 , P3_U3068 , P3_R1179_U67 );
not NOT1_25606 ( P3_R1179_U455 , P3_R1179_U146 );
nand NAND2_25607 ( P3_R1179_U456 , P3_R1179_U271 , P3_R1179_U455 );
nand NAND2_25608 ( P3_R1179_U457 , P3_R1179_U146 , P3_R1179_U176 );
nand NAND2_25609 ( P3_R1179_U458 , P3_U3437 , P3_R1179_U63 );
nand NAND2_25610 ( P3_R1179_U459 , P3_U3072 , P3_R1179_U60 );
nand NAND2_25611 ( P3_R1179_U460 , P3_R1179_U459 , P3_R1179_U458 );
nand NAND2_25612 ( P3_R1179_U461 , P3_U3434 , P3_R1179_U64 );
nand NAND2_25613 ( P3_R1179_U462 , P3_U3073 , P3_R1179_U61 );
nand NAND2_25614 ( P3_R1179_U463 , P3_R1179_U336 , P3_R1179_U93 );
nand NAND2_25615 ( P3_R1179_U464 , P3_R1179_U177 , P3_R1179_U328 );
nand NAND2_25616 ( P3_R1179_U465 , P3_U3431 , P3_R1179_U65 );
nand NAND2_25617 ( P3_R1179_U466 , P3_U3078 , P3_R1179_U62 );
nand NAND2_25618 ( P3_R1179_U467 , P3_R1179_U337 , P3_R1179_U179 );
nand NAND2_25619 ( P3_R1179_U468 , P3_R1179_U261 , P3_R1179_U178 );
nand NAND2_25620 ( P3_R1179_U469 , P3_U3428 , P3_R1179_U59 );
nand NAND2_25621 ( P3_R1179_U470 , P3_U3079 , P3_R1179_U58 );
not NOT1_25622 ( P3_R1179_U471 , P3_R1179_U149 );
nand NAND2_25623 ( P3_R1179_U472 , P3_R1179_U257 , P3_R1179_U471 );
nand NAND2_25624 ( P3_R1179_U473 , P3_R1179_U149 , P3_R1179_U180 );
nand NAND2_25625 ( P3_R1179_U474 , P3_U3425 , P3_R1179_U57 );
nand NAND2_25626 ( P3_R1179_U475 , P3_U3071 , P3_R1179_U56 );
not NOT1_25627 ( P3_R1179_U476 , P3_R1179_U150 );
nand NAND2_25628 ( P3_R1179_U477 , P3_R1179_U253 , P3_R1179_U476 );
nand NAND2_25629 ( P3_R1179_U478 , P3_R1179_U150 , P3_R1179_U181 );
nand NAND2_25630 ( P3_R1179_U479 , P3_U3422 , P3_R1179_U53 );
nand NAND2_25631 ( P3_R1179_U480 , P3_U3062 , P3_R1179_U51 );
nand NAND2_25632 ( P3_R1179_U481 , P3_R1179_U480 , P3_R1179_U479 );
nand NAND2_25633 ( P3_R1179_U482 , P3_U3419 , P3_R1179_U54 );
nand NAND2_25634 ( P3_R1179_U483 , P3_U3061 , P3_R1179_U52 );
nand NAND2_25635 ( P3_R1179_U484 , P3_R1179_U347 , P3_R1179_U94 );
nand NAND2_25636 ( P3_R1179_U485 , P3_R1179_U182 , P3_R1179_U339 );
and AND2_25637 ( P3_R1269_U6 , P3_R1269_U107 , P3_R1269_U108 );
and AND2_25638 ( P3_R1269_U7 , P3_R1269_U118 , P3_R1269_U117 );
and AND2_25639 ( P3_R1269_U8 , P3_R1269_U142 , P3_R1269_U141 );
and AND2_25640 ( P3_R1269_U9 , P3_R1269_U200 , P3_R1269_U199 );
and AND2_25641 ( P3_R1269_U10 , P3_R1269_U202 , P3_R1269_U201 );
nand NAND3_25642 ( P3_R1269_U11 , P3_R1269_U10 , P3_R1269_U194 , P3_R1269_U196 );
not NOT1_25643 ( P3_R1269_U12 , P3_U3116 );
not NOT1_25644 ( P3_R1269_U13 , P3_U3094 );
not NOT1_25645 ( P3_R1269_U14 , P3_U3095 );
not NOT1_25646 ( P3_R1269_U15 , P3_U3130 );
not NOT1_25647 ( P3_R1269_U16 , P3_U3136 );
not NOT1_25648 ( P3_R1269_U17 , P3_U3135 );
not NOT1_25649 ( P3_R1269_U18 , P3_U3106 );
not NOT1_25650 ( P3_R1269_U19 , P3_U3107 );
not NOT1_25651 ( P3_R1269_U20 , P3_U3112 );
not NOT1_25652 ( P3_R1269_U21 , P3_U3113 );
not NOT1_25653 ( P3_R1269_U22 , P3_U3114 );
not NOT1_25654 ( P3_R1269_U23 , P3_U3142 );
not NOT1_25655 ( P3_R1269_U24 , P3_U3141 );
not NOT1_25656 ( P3_R1269_U25 , P3_U3146 );
not NOT1_25657 ( P3_R1269_U26 , P3_U3145 );
not NOT1_25658 ( P3_R1269_U27 , P3_U3144 );
not NOT1_25659 ( P3_R1269_U28 , P3_U3143 );
not NOT1_25660 ( P3_R1269_U29 , P3_U3111 );
not NOT1_25661 ( P3_R1269_U30 , P3_U3109 );
not NOT1_25662 ( P3_R1269_U31 , P3_U3110 );
not NOT1_25663 ( P3_R1269_U32 , P3_U3108 );
not NOT1_25664 ( P3_R1269_U33 , P3_U3140 );
not NOT1_25665 ( P3_R1269_U34 , P3_U3139 );
not NOT1_25666 ( P3_R1269_U35 , P3_U3138 );
not NOT1_25667 ( P3_R1269_U36 , P3_U3137 );
not NOT1_25668 ( P3_R1269_U37 , P3_U3101 );
not NOT1_25669 ( P3_R1269_U38 , P3_U3100 );
not NOT1_25670 ( P3_R1269_U39 , P3_U3104 );
not NOT1_25671 ( P3_R1269_U40 , P3_U3105 );
not NOT1_25672 ( P3_R1269_U41 , P3_U3103 );
not NOT1_25673 ( P3_R1269_U42 , P3_U3102 );
not NOT1_25674 ( P3_R1269_U43 , P3_U3134 );
not NOT1_25675 ( P3_R1269_U44 , P3_U3133 );
not NOT1_25676 ( P3_R1269_U45 , P3_U3132 );
not NOT1_25677 ( P3_R1269_U46 , P3_U3131 );
not NOT1_25678 ( P3_R1269_U47 , P3_U3099 );
not NOT1_25679 ( P3_R1269_U48 , P3_U3098 );
nand NAND2_25680 ( P3_R1269_U49 , P3_R1269_U157 , P3_R1269_U156 );
not NOT1_25681 ( P3_R1269_U50 , P3_U3129 );
not NOT1_25682 ( P3_R1269_U51 , P3_U3096 );
not NOT1_25683 ( P3_R1269_U52 , P3_U3123 );
not NOT1_25684 ( P3_R1269_U53 , P3_U3124 );
not NOT1_25685 ( P3_R1269_U54 , P3_U3128 );
not NOT1_25686 ( P3_R1269_U55 , P3_U3127 );
not NOT1_25687 ( P3_R1269_U56 , P3_U3126 );
not NOT1_25688 ( P3_R1269_U57 , P3_U3125 );
not NOT1_25689 ( P3_R1269_U58 , P3_U3087 );
not NOT1_25690 ( P3_R1269_U59 , P3_U3089 );
not NOT1_25691 ( P3_R1269_U60 , P3_U3088 );
not NOT1_25692 ( P3_R1269_U61 , P3_U3086 );
not NOT1_25693 ( P3_R1269_U62 , P3_U3093 );
not NOT1_25694 ( P3_R1269_U63 , P3_U3092 );
not NOT1_25695 ( P3_R1269_U64 , P3_U3090 );
not NOT1_25696 ( P3_R1269_U65 , P3_U3091 );
not NOT1_25697 ( P3_R1269_U66 , P3_U3120 );
not NOT1_25698 ( P3_R1269_U67 , P3_U3119 );
nand NAND2_25699 ( P3_R1269_U68 , P3_R1269_U178 , P3_R1269_U177 );
not NOT1_25700 ( P3_R1269_U69 , P3_U3121 );
not NOT1_25701 ( P3_R1269_U70 , P3_U3122 );
not NOT1_25702 ( P3_R1269_U71 , P3_U3118 );
not NOT1_25703 ( P3_R1269_U72 , P3_U3149 );
and AND2_25704 ( P3_R1269_U73 , P3_R1269_U111 , P3_R1269_U110 );
and AND2_25705 ( P3_R1269_U74 , P3_R1269_U7 , P3_R1269_U124 );
and AND2_25706 ( P3_R1269_U75 , P3_U3111 , P3_R1269_U28 );
and AND2_25707 ( P3_R1269_U76 , P3_U3110 , P3_R1269_U23 );
and AND3_25708 ( P3_R1269_U77 , P3_R1269_U126 , P3_R1269_U127 , P3_R1269_U78 );
and AND2_25709 ( P3_R1269_U78 , P3_R1269_U130 , P3_R1269_U129 );
and AND2_25710 ( P3_R1269_U79 , P3_R1269_U6 , P3_R1269_U80 );
and AND2_25711 ( P3_R1269_U80 , P3_R1269_U138 , P3_R1269_U139 );
and AND2_25712 ( P3_R1269_U81 , P3_U3104 , P3_R1269_U16 );
and AND2_25713 ( P3_R1269_U82 , P3_U3105 , P3_R1269_U36 );
and AND3_25714 ( P3_R1269_U83 , P3_R1269_U143 , P3_R1269_U144 , P3_R1269_U85 );
and AND2_25715 ( P3_R1269_U84 , P3_R1269_U146 , P3_R1269_U145 );
and AND2_25716 ( P3_R1269_U85 , P3_R1269_U84 , P3_R1269_U8 );
and AND2_25717 ( P3_R1269_U86 , P3_U3134 , P3_R1269_U42 );
and AND2_25718 ( P3_R1269_U87 , P3_U3133 , P3_R1269_U37 );
and AND3_25719 ( P3_R1269_U88 , P3_R1269_U148 , P3_R1269_U150 , P3_R1269_U89 );
and AND2_25720 ( P3_R1269_U89 , P3_R1269_U152 , P3_R1269_U151 );
and AND2_25721 ( P3_R1269_U90 , P3_R1269_U104 , P3_R1269_U103 );
and AND2_25722 ( P3_R1269_U91 , P3_R1269_U162 , P3_R1269_U161 );
and AND2_25723 ( P3_R1269_U92 , P3_U3128 , P3_R1269_U51 );
and AND4_25724 ( P3_R1269_U93 , P3_R1269_U170 , P3_R1269_U169 , P3_R1269_U171 , P3_R1269_U165 );
and AND2_25725 ( P3_R1269_U94 , P3_R1269_U175 , P3_R1269_U174 );
and AND5_25726 ( P3_R1269_U95 , P3_R1269_U172 , P3_R1269_U94 , P3_R1269_U173 , P3_R1269_U96 , P3_R1269_U176 );
and AND3_25727 ( P3_R1269_U96 , P3_R1269_U193 , P3_R1269_U191 , P3_R1269_U192 );
and AND2_25728 ( P3_R1269_U97 , P3_U3120 , P3_R1269_U60 );
and AND2_25729 ( P3_R1269_U98 , P3_R1269_U174 , P3_R1269_U175 );
and AND2_25730 ( P3_R1269_U99 , P3_R1269_U198 , P3_R1269_U186 );
not NOT1_25731 ( P3_R1269_U100 , P3_U3084 );
not NOT1_25732 ( P3_R1269_U101 , P3_U3085 );
nand NAND2_25733 ( P3_R1269_U102 , P3_R1269_U187 , P3_R1269_U195 );
nand NAND2_25734 ( P3_R1269_U103 , P3_U3094 , P3_R1269_U56 );
nand NAND2_25735 ( P3_R1269_U104 , P3_U3095 , P3_R1269_U55 );
nand NAND2_25736 ( P3_R1269_U105 , P3_U3130 , P3_R1269_U48 );
nand NAND2_25737 ( P3_R1269_U106 , P3_U3106 , P3_R1269_U35 );
nand NAND2_25738 ( P3_R1269_U107 , P3_U3135 , P3_R1269_U41 );
nand NAND2_25739 ( P3_R1269_U108 , P3_U3136 , P3_R1269_U39 );
nand NAND2_25740 ( P3_R1269_U109 , P3_U3107 , P3_R1269_U34 );
nand NAND2_25741 ( P3_R1269_U110 , P3_U3112 , P3_R1269_U27 );
nand NAND2_25742 ( P3_R1269_U111 , P3_U3113 , P3_R1269_U26 );
nand NAND2_25743 ( P3_R1269_U112 , P3_U3147 , P3_U3148 );
nand NAND2_25744 ( P3_R1269_U113 , P3_U3115 , P3_R1269_U112 );
or OR2_25745 ( P3_R1269_U114 , P3_U3147 , P3_U3148 );
nand NAND2_25746 ( P3_R1269_U115 , P3_U3114 , P3_R1269_U25 );
nand NAND5_25747 ( P3_R1269_U116 , P3_R1269_U111 , P3_R1269_U110 , P3_R1269_U113 , P3_R1269_U115 , P3_R1269_U114 );
nand NAND2_25748 ( P3_R1269_U117 , P3_U3142 , P3_R1269_U31 );
nand NAND2_25749 ( P3_R1269_U118 , P3_U3141 , P3_R1269_U30 );
nand NAND2_25750 ( P3_R1269_U119 , P3_U3146 , P3_R1269_U22 );
nand NAND2_25751 ( P3_R1269_U120 , P3_U3145 , P3_R1269_U21 );
nand NAND2_25752 ( P3_R1269_U121 , P3_R1269_U120 , P3_R1269_U119 );
nand NAND2_25753 ( P3_R1269_U122 , P3_R1269_U73 , P3_R1269_U121 );
nand NAND2_25754 ( P3_R1269_U123 , P3_U3144 , P3_R1269_U20 );
nand NAND2_25755 ( P3_R1269_U124 , P3_U3143 , P3_R1269_U29 );
nand NAND4_25756 ( P3_R1269_U125 , P3_R1269_U122 , P3_R1269_U123 , P3_R1269_U116 , P3_R1269_U74 );
nand NAND2_25757 ( P3_R1269_U126 , P3_R1269_U75 , P3_R1269_U7 );
nand NAND2_25758 ( P3_R1269_U127 , P3_U3109 , P3_R1269_U24 );
nand NAND2_25759 ( P3_R1269_U128 , P3_U3141 , P3_R1269_U30 );
nand NAND2_25760 ( P3_R1269_U129 , P3_R1269_U76 , P3_R1269_U128 );
nand NAND2_25761 ( P3_R1269_U130 , P3_U3108 , P3_R1269_U33 );
nand NAND2_25762 ( P3_R1269_U131 , P3_R1269_U125 , P3_R1269_U77 );
nand NAND2_25763 ( P3_R1269_U132 , P3_U3140 , P3_R1269_U32 );
nand NAND2_25764 ( P3_R1269_U133 , P3_R1269_U132 , P3_R1269_U131 );
nand NAND2_25765 ( P3_R1269_U134 , P3_R1269_U133 , P3_R1269_U109 );
nand NAND2_25766 ( P3_R1269_U135 , P3_U3139 , P3_R1269_U19 );
nand NAND2_25767 ( P3_R1269_U136 , P3_R1269_U135 , P3_R1269_U134 );
nand NAND2_25768 ( P3_R1269_U137 , P3_R1269_U136 , P3_R1269_U106 );
nand NAND2_25769 ( P3_R1269_U138 , P3_U3138 , P3_R1269_U18 );
nand NAND2_25770 ( P3_R1269_U139 , P3_U3137 , P3_R1269_U40 );
nand NAND2_25771 ( P3_R1269_U140 , P3_R1269_U137 , P3_R1269_U79 );
nand NAND2_25772 ( P3_R1269_U141 , P3_U3101 , P3_R1269_U44 );
nand NAND2_25773 ( P3_R1269_U142 , P3_U3100 , P3_R1269_U45 );
nand NAND2_25774 ( P3_R1269_U143 , P3_R1269_U81 , P3_R1269_U107 );
nand NAND2_25775 ( P3_R1269_U144 , P3_R1269_U82 , P3_R1269_U6 );
nand NAND2_25776 ( P3_R1269_U145 , P3_U3103 , P3_R1269_U17 );
nand NAND2_25777 ( P3_R1269_U146 , P3_U3102 , P3_R1269_U43 );
nand NAND2_25778 ( P3_R1269_U147 , P3_R1269_U140 , P3_R1269_U83 );
nand NAND2_25779 ( P3_R1269_U148 , P3_R1269_U86 , P3_R1269_U8 );
nand NAND2_25780 ( P3_R1269_U149 , P3_U3100 , P3_R1269_U45 );
nand NAND2_25781 ( P3_R1269_U150 , P3_R1269_U87 , P3_R1269_U149 );
nand NAND2_25782 ( P3_R1269_U151 , P3_U3132 , P3_R1269_U38 );
nand NAND2_25783 ( P3_R1269_U152 , P3_U3131 , P3_R1269_U47 );
nand NAND2_25784 ( P3_R1269_U153 , P3_R1269_U147 , P3_R1269_U88 );
nand NAND2_25785 ( P3_R1269_U154 , P3_U3099 , P3_R1269_U46 );
nand NAND2_25786 ( P3_R1269_U155 , P3_R1269_U154 , P3_R1269_U153 );
nand NAND2_25787 ( P3_R1269_U156 , P3_R1269_U155 , P3_R1269_U105 );
nand NAND2_25788 ( P3_R1269_U157 , P3_U3098 , P3_R1269_U15 );
not NOT1_25789 ( P3_R1269_U158 , P3_R1269_U49 );
nand NAND2_25790 ( P3_R1269_U159 , P3_U3129 , P3_R1269_U158 );
nand NAND2_25791 ( P3_R1269_U160 , P3_U3097 , P3_R1269_U159 );
nand NAND2_25792 ( P3_R1269_U161 , P3_R1269_U49 , P3_R1269_U50 );
nand NAND2_25793 ( P3_R1269_U162 , P3_U3096 , P3_R1269_U54 );
nand NAND3_25794 ( P3_R1269_U163 , P3_R1269_U90 , P3_R1269_U160 , P3_R1269_U91 );
nand NAND2_25795 ( P3_R1269_U164 , P3_U3123 , P3_R1269_U65 );
nand NAND2_25796 ( P3_R1269_U165 , P3_U3124 , P3_R1269_U63 );
nand NAND2_25797 ( P3_R1269_U166 , P3_R1269_U92 , P3_R1269_U104 );
nand NAND2_25798 ( P3_R1269_U167 , P3_U3127 , P3_R1269_U14 );
nand NAND2_25799 ( P3_R1269_U168 , P3_R1269_U167 , P3_R1269_U166 );
nand NAND2_25800 ( P3_R1269_U169 , P3_R1269_U168 , P3_R1269_U103 );
nand NAND2_25801 ( P3_R1269_U170 , P3_U3126 , P3_R1269_U13 );
nand NAND2_25802 ( P3_R1269_U171 , P3_U3125 , P3_R1269_U62 );
nand NAND3_25803 ( P3_R1269_U172 , P3_R1269_U93 , P3_R1269_U163 , P3_R1269_U164 );
nand NAND2_25804 ( P3_R1269_U173 , P3_U3087 , P3_R1269_U67 );
nand NAND2_25805 ( P3_R1269_U174 , P3_U3089 , P3_R1269_U69 );
nand NAND2_25806 ( P3_R1269_U175 , P3_U3088 , P3_R1269_U66 );
nand NAND2_25807 ( P3_R1269_U176 , P3_U3086 , P3_R1269_U71 );
nand NAND2_25808 ( P3_R1269_U177 , P3_R1269_U97 , P3_R1269_U173 );
nand NAND2_25809 ( P3_R1269_U178 , P3_U3119 , P3_R1269_U58 );
not NOT1_25810 ( P3_R1269_U179 , P3_R1269_U68 );
nand NAND2_25811 ( P3_R1269_U180 , P3_U3121 , P3_R1269_U59 );
nand NAND2_25812 ( P3_R1269_U181 , P3_U3122 , P3_R1269_U64 );
nand NAND2_25813 ( P3_R1269_U182 , P3_R1269_U181 , P3_R1269_U180 );
nand NAND2_25814 ( P3_R1269_U183 , P3_R1269_U179 , P3_R1269_U71 );
nand NAND2_25815 ( P3_R1269_U184 , P3_R1269_U183 , P3_R1269_U61 );
nand NAND4_25816 ( P3_R1269_U185 , P3_R1269_U98 , P3_R1269_U182 , P3_R1269_U173 , P3_R1269_U176 );
nand NAND2_25817 ( P3_R1269_U186 , P3_U3118 , P3_R1269_U68 );
nand NAND2_25818 ( P3_R1269_U187 , P3_R1269_U9 , P3_R1269_U101 );
nand NAND2_25819 ( P3_R1269_U188 , P3_U3093 , P3_R1269_U57 );
nand NAND2_25820 ( P3_R1269_U189 , P3_U3092 , P3_R1269_U53 );
nand NAND2_25821 ( P3_R1269_U190 , P3_R1269_U189 , P3_R1269_U188 );
nand NAND3_25822 ( P3_R1269_U191 , P3_R1269_U165 , P3_R1269_U190 , P3_R1269_U164 );
nand NAND2_25823 ( P3_R1269_U192 , P3_U3090 , P3_R1269_U70 );
nand NAND2_25824 ( P3_R1269_U193 , P3_U3091 , P3_R1269_U52 );
nand NAND2_25825 ( P3_R1269_U194 , P3_R1269_U102 , P3_R1269_U95 );
nand NAND2_25826 ( P3_R1269_U195 , P3_U3117 , P3_R1269_U9 );
nand NAND2_25827 ( P3_R1269_U196 , P3_R1269_U197 , P3_R1269_U102 );
nand NAND3_25828 ( P3_R1269_U197 , P3_R1269_U185 , P3_R1269_U184 , P3_R1269_U99 );
nand NAND2_25829 ( P3_R1269_U198 , P3_U3117 , P3_R1269_U101 );
nand NAND2_25830 ( P3_R1269_U199 , P3_U3084 , P3_R1269_U12 );
nand NAND2_25831 ( P3_R1269_U200 , P3_U3116 , P3_R1269_U100 );
nand NAND3_25832 ( P3_R1269_U201 , P3_U3116 , P3_R1269_U72 , P3_R1269_U100 );
nand NAND3_25833 ( P3_R1269_U202 , P3_U3149 , P3_R1269_U12 , P3_U3084 );
and AND2_25834 ( P3_R1110_U4 , P3_R1110_U179 , P3_R1110_U178 );
and AND2_25835 ( P3_R1110_U5 , P3_R1110_U197 , P3_R1110_U196 );
and AND2_25836 ( P3_R1110_U6 , P3_R1110_U237 , P3_R1110_U236 );
and AND2_25837 ( P3_R1110_U7 , P3_R1110_U246 , P3_R1110_U245 );
and AND2_25838 ( P3_R1110_U8 , P3_R1110_U264 , P3_R1110_U263 );
and AND2_25839 ( P3_R1110_U9 , P3_R1110_U272 , P3_R1110_U271 );
and AND2_25840 ( P3_R1110_U10 , P3_R1110_U351 , P3_R1110_U348 );
and AND2_25841 ( P3_R1110_U11 , P3_R1110_U344 , P3_R1110_U341 );
and AND2_25842 ( P3_R1110_U12 , P3_R1110_U335 , P3_R1110_U332 );
and AND2_25843 ( P3_R1110_U13 , P3_R1110_U326 , P3_R1110_U323 );
and AND2_25844 ( P3_R1110_U14 , P3_R1110_U320 , P3_R1110_U318 );
and AND2_25845 ( P3_R1110_U15 , P3_R1110_U313 , P3_R1110_U310 );
and AND2_25846 ( P3_R1110_U16 , P3_R1110_U235 , P3_R1110_U232 );
and AND2_25847 ( P3_R1110_U17 , P3_R1110_U227 , P3_R1110_U224 );
and AND2_25848 ( P3_R1110_U18 , P3_R1110_U213 , P3_R1110_U210 );
not NOT1_25849 ( P3_R1110_U19 , P3_U3407 );
not NOT1_25850 ( P3_R1110_U20 , P3_U3070 );
not NOT1_25851 ( P3_R1110_U21 , P3_U3069 );
nand NAND2_25852 ( P3_R1110_U22 , P3_U3070 , P3_U3407 );
not NOT1_25853 ( P3_R1110_U23 , P3_U3410 );
not NOT1_25854 ( P3_R1110_U24 , P3_U3401 );
not NOT1_25855 ( P3_R1110_U25 , P3_U3059 );
not NOT1_25856 ( P3_R1110_U26 , P3_U3066 );
not NOT1_25857 ( P3_R1110_U27 , P3_U3395 );
not NOT1_25858 ( P3_R1110_U28 , P3_U3067 );
not NOT1_25859 ( P3_R1110_U29 , P3_U3387 );
not NOT1_25860 ( P3_R1110_U30 , P3_U3076 );
nand NAND2_25861 ( P3_R1110_U31 , P3_U3076 , P3_U3387 );
not NOT1_25862 ( P3_R1110_U32 , P3_U3398 );
not NOT1_25863 ( P3_R1110_U33 , P3_U3063 );
nand NAND2_25864 ( P3_R1110_U34 , P3_U3059 , P3_U3401 );
not NOT1_25865 ( P3_R1110_U35 , P3_U3404 );
not NOT1_25866 ( P3_R1110_U36 , P3_U3413 );
not NOT1_25867 ( P3_R1110_U37 , P3_U3083 );
not NOT1_25868 ( P3_R1110_U38 , P3_U3082 );
not NOT1_25869 ( P3_R1110_U39 , P3_U3416 );
nand NAND2_25870 ( P3_R1110_U40 , P3_R1110_U61 , P3_R1110_U205 );
nand NAND2_25871 ( P3_R1110_U41 , P3_R1110_U117 , P3_R1110_U193 );
nand NAND2_25872 ( P3_R1110_U42 , P3_R1110_U182 , P3_R1110_U183 );
nand NAND2_25873 ( P3_R1110_U43 , P3_U3392 , P3_U3077 );
nand NAND2_25874 ( P3_R1110_U44 , P3_R1110_U122 , P3_R1110_U219 );
nand NAND2_25875 ( P3_R1110_U45 , P3_R1110_U216 , P3_R1110_U215 );
not NOT1_25876 ( P3_R1110_U46 , P3_U3900 );
not NOT1_25877 ( P3_R1110_U47 , P3_U3052 );
not NOT1_25878 ( P3_R1110_U48 , P3_U3056 );
not NOT1_25879 ( P3_R1110_U49 , P3_U3901 );
not NOT1_25880 ( P3_R1110_U50 , P3_U3902 );
not NOT1_25881 ( P3_R1110_U51 , P3_U3057 );
not NOT1_25882 ( P3_R1110_U52 , P3_U3903 );
not NOT1_25883 ( P3_R1110_U53 , P3_U3064 );
not NOT1_25884 ( P3_R1110_U54 , P3_U3906 );
not NOT1_25885 ( P3_R1110_U55 , P3_U3074 );
not NOT1_25886 ( P3_R1110_U56 , P3_U3437 );
not NOT1_25887 ( P3_R1110_U57 , P3_U3072 );
not NOT1_25888 ( P3_R1110_U58 , P3_U3068 );
nand NAND2_25889 ( P3_R1110_U59 , P3_U3072 , P3_U3437 );
not NOT1_25890 ( P3_R1110_U60 , P3_U3440 );
nand NAND2_25891 ( P3_R1110_U61 , P3_U3083 , P3_U3413 );
not NOT1_25892 ( P3_R1110_U62 , P3_U3419 );
not NOT1_25893 ( P3_R1110_U63 , P3_U3061 );
not NOT1_25894 ( P3_R1110_U64 , P3_U3425 );
not NOT1_25895 ( P3_R1110_U65 , P3_U3071 );
not NOT1_25896 ( P3_R1110_U66 , P3_U3422 );
not NOT1_25897 ( P3_R1110_U67 , P3_U3062 );
nand NAND2_25898 ( P3_R1110_U68 , P3_U3062 , P3_U3422 );
not NOT1_25899 ( P3_R1110_U69 , P3_U3428 );
not NOT1_25900 ( P3_R1110_U70 , P3_U3079 );
not NOT1_25901 ( P3_R1110_U71 , P3_U3431 );
not NOT1_25902 ( P3_R1110_U72 , P3_U3078 );
not NOT1_25903 ( P3_R1110_U73 , P3_U3434 );
not NOT1_25904 ( P3_R1110_U74 , P3_U3073 );
not NOT1_25905 ( P3_R1110_U75 , P3_U3443 );
not NOT1_25906 ( P3_R1110_U76 , P3_U3081 );
nand NAND2_25907 ( P3_R1110_U77 , P3_U3081 , P3_U3443 );
not NOT1_25908 ( P3_R1110_U78 , P3_U3445 );
not NOT1_25909 ( P3_R1110_U79 , P3_U3080 );
nand NAND2_25910 ( P3_R1110_U80 , P3_U3080 , P3_U3445 );
not NOT1_25911 ( P3_R1110_U81 , P3_U3907 );
not NOT1_25912 ( P3_R1110_U82 , P3_U3905 );
not NOT1_25913 ( P3_R1110_U83 , P3_U3060 );
not NOT1_25914 ( P3_R1110_U84 , P3_U3904 );
not NOT1_25915 ( P3_R1110_U85 , P3_U3065 );
nand NAND2_25916 ( P3_R1110_U86 , P3_U3901 , P3_U3056 );
not NOT1_25917 ( P3_R1110_U87 , P3_U3053 );
not NOT1_25918 ( P3_R1110_U88 , P3_U3899 );
nand NAND2_25919 ( P3_R1110_U89 , P3_R1110_U306 , P3_R1110_U176 );
not NOT1_25920 ( P3_R1110_U90 , P3_U3075 );
nand NAND2_25921 ( P3_R1110_U91 , P3_R1110_U77 , P3_R1110_U315 );
nand NAND2_25922 ( P3_R1110_U92 , P3_R1110_U261 , P3_R1110_U260 );
nand NAND2_25923 ( P3_R1110_U93 , P3_R1110_U68 , P3_R1110_U337 );
nand NAND2_25924 ( P3_R1110_U94 , P3_R1110_U457 , P3_R1110_U456 );
nand NAND2_25925 ( P3_R1110_U95 , P3_R1110_U504 , P3_R1110_U503 );
nand NAND2_25926 ( P3_R1110_U96 , P3_R1110_U375 , P3_R1110_U374 );
nand NAND2_25927 ( P3_R1110_U97 , P3_R1110_U380 , P3_R1110_U379 );
nand NAND2_25928 ( P3_R1110_U98 , P3_R1110_U387 , P3_R1110_U386 );
nand NAND2_25929 ( P3_R1110_U99 , P3_R1110_U394 , P3_R1110_U393 );
nand NAND2_25930 ( P3_R1110_U100 , P3_R1110_U399 , P3_R1110_U398 );
nand NAND2_25931 ( P3_R1110_U101 , P3_R1110_U408 , P3_R1110_U407 );
nand NAND2_25932 ( P3_R1110_U102 , P3_R1110_U415 , P3_R1110_U414 );
nand NAND2_25933 ( P3_R1110_U103 , P3_R1110_U422 , P3_R1110_U421 );
nand NAND2_25934 ( P3_R1110_U104 , P3_R1110_U429 , P3_R1110_U428 );
nand NAND2_25935 ( P3_R1110_U105 , P3_R1110_U434 , P3_R1110_U433 );
nand NAND2_25936 ( P3_R1110_U106 , P3_R1110_U441 , P3_R1110_U440 );
nand NAND2_25937 ( P3_R1110_U107 , P3_R1110_U448 , P3_R1110_U447 );
nand NAND2_25938 ( P3_R1110_U108 , P3_R1110_U462 , P3_R1110_U461 );
nand NAND2_25939 ( P3_R1110_U109 , P3_R1110_U467 , P3_R1110_U466 );
nand NAND2_25940 ( P3_R1110_U110 , P3_R1110_U474 , P3_R1110_U473 );
nand NAND2_25941 ( P3_R1110_U111 , P3_R1110_U481 , P3_R1110_U480 );
nand NAND2_25942 ( P3_R1110_U112 , P3_R1110_U488 , P3_R1110_U487 );
nand NAND2_25943 ( P3_R1110_U113 , P3_R1110_U495 , P3_R1110_U494 );
nand NAND2_25944 ( P3_R1110_U114 , P3_R1110_U500 , P3_R1110_U499 );
and AND2_25945 ( P3_R1110_U115 , P3_R1110_U189 , P3_R1110_U187 );
and AND2_25946 ( P3_R1110_U116 , P3_R1110_U4 , P3_R1110_U180 );
and AND2_25947 ( P3_R1110_U117 , P3_R1110_U194 , P3_R1110_U192 );
and AND2_25948 ( P3_R1110_U118 , P3_R1110_U201 , P3_R1110_U200 );
and AND3_25949 ( P3_R1110_U119 , P3_R1110_U382 , P3_R1110_U381 , P3_R1110_U22 );
and AND2_25950 ( P3_R1110_U120 , P3_R1110_U212 , P3_R1110_U5 );
and AND2_25951 ( P3_R1110_U121 , P3_R1110_U181 , P3_R1110_U180 );
and AND2_25952 ( P3_R1110_U122 , P3_R1110_U220 , P3_R1110_U218 );
and AND3_25953 ( P3_R1110_U123 , P3_R1110_U389 , P3_R1110_U388 , P3_R1110_U34 );
and AND2_25954 ( P3_R1110_U124 , P3_R1110_U226 , P3_R1110_U4 );
and AND2_25955 ( P3_R1110_U125 , P3_R1110_U234 , P3_R1110_U181 );
and AND2_25956 ( P3_R1110_U126 , P3_R1110_U204 , P3_R1110_U6 );
and AND2_25957 ( P3_R1110_U127 , P3_R1110_U239 , P3_R1110_U171 );
and AND2_25958 ( P3_R1110_U128 , P3_R1110_U250 , P3_R1110_U7 );
and AND2_25959 ( P3_R1110_U129 , P3_R1110_U248 , P3_R1110_U172 );
and AND2_25960 ( P3_R1110_U130 , P3_R1110_U268 , P3_R1110_U267 );
and AND3_25961 ( P3_R1110_U131 , P3_R1110_U9 , P3_R1110_U282 , P3_R1110_U273 );
and AND2_25962 ( P3_R1110_U132 , P3_R1110_U285 , P3_R1110_U280 );
and AND2_25963 ( P3_R1110_U133 , P3_R1110_U301 , P3_R1110_U298 );
and AND2_25964 ( P3_R1110_U134 , P3_R1110_U368 , P3_R1110_U302 );
and AND2_25965 ( P3_R1110_U135 , P3_R1110_U160 , P3_R1110_U278 );
and AND3_25966 ( P3_R1110_U136 , P3_R1110_U455 , P3_R1110_U454 , P3_R1110_U80 );
and AND2_25967 ( P3_R1110_U137 , P3_R1110_U325 , P3_R1110_U9 );
and AND3_25968 ( P3_R1110_U138 , P3_R1110_U469 , P3_R1110_U468 , P3_R1110_U59 );
and AND2_25969 ( P3_R1110_U139 , P3_R1110_U334 , P3_R1110_U8 );
and AND3_25970 ( P3_R1110_U140 , P3_R1110_U490 , P3_R1110_U489 , P3_R1110_U172 );
and AND2_25971 ( P3_R1110_U141 , P3_R1110_U343 , P3_R1110_U7 );
and AND3_25972 ( P3_R1110_U142 , P3_R1110_U502 , P3_R1110_U501 , P3_R1110_U171 );
and AND2_25973 ( P3_R1110_U143 , P3_R1110_U350 , P3_R1110_U6 );
nand NAND2_25974 ( P3_R1110_U144 , P3_R1110_U118 , P3_R1110_U202 );
nand NAND2_25975 ( P3_R1110_U145 , P3_R1110_U217 , P3_R1110_U229 );
not NOT1_25976 ( P3_R1110_U146 , P3_U3054 );
not NOT1_25977 ( P3_R1110_U147 , P3_U3908 );
and AND2_25978 ( P3_R1110_U148 , P3_R1110_U403 , P3_R1110_U402 );
nand NAND3_25979 ( P3_R1110_U149 , P3_R1110_U304 , P3_R1110_U169 , P3_R1110_U364 );
and AND2_25980 ( P3_R1110_U150 , P3_R1110_U410 , P3_R1110_U409 );
nand NAND3_25981 ( P3_R1110_U151 , P3_R1110_U370 , P3_R1110_U369 , P3_R1110_U134 );
and AND2_25982 ( P3_R1110_U152 , P3_R1110_U417 , P3_R1110_U416 );
nand NAND3_25983 ( P3_R1110_U153 , P3_R1110_U365 , P3_R1110_U299 , P3_R1110_U86 );
and AND2_25984 ( P3_R1110_U154 , P3_R1110_U424 , P3_R1110_U423 );
nand NAND2_25985 ( P3_R1110_U155 , P3_R1110_U293 , P3_R1110_U292 );
and AND2_25986 ( P3_R1110_U156 , P3_R1110_U436 , P3_R1110_U435 );
nand NAND2_25987 ( P3_R1110_U157 , P3_R1110_U289 , P3_R1110_U288 );
and AND2_25988 ( P3_R1110_U158 , P3_R1110_U443 , P3_R1110_U442 );
nand NAND2_25989 ( P3_R1110_U159 , P3_R1110_U132 , P3_R1110_U284 );
and AND2_25990 ( P3_R1110_U160 , P3_R1110_U450 , P3_R1110_U449 );
nand NAND2_25991 ( P3_R1110_U161 , P3_R1110_U43 , P3_R1110_U327 );
nand NAND2_25992 ( P3_R1110_U162 , P3_R1110_U130 , P3_R1110_U269 );
and AND2_25993 ( P3_R1110_U163 , P3_R1110_U476 , P3_R1110_U475 );
nand NAND2_25994 ( P3_R1110_U164 , P3_R1110_U257 , P3_R1110_U256 );
and AND2_25995 ( P3_R1110_U165 , P3_R1110_U483 , P3_R1110_U482 );
nand NAND2_25996 ( P3_R1110_U166 , P3_R1110_U253 , P3_R1110_U252 );
nand NAND2_25997 ( P3_R1110_U167 , P3_R1110_U243 , P3_R1110_U242 );
nand NAND2_25998 ( P3_R1110_U168 , P3_R1110_U367 , P3_R1110_U366 );
nand NAND2_25999 ( P3_R1110_U169 , P3_U3053 , P3_R1110_U151 );
not NOT1_26000 ( P3_R1110_U170 , P3_R1110_U34 );
nand NAND2_26001 ( P3_R1110_U171 , P3_U3416 , P3_U3082 );
nand NAND2_26002 ( P3_R1110_U172 , P3_U3071 , P3_U3425 );
nand NAND2_26003 ( P3_R1110_U173 , P3_U3057 , P3_U3902 );
not NOT1_26004 ( P3_R1110_U174 , P3_R1110_U68 );
not NOT1_26005 ( P3_R1110_U175 , P3_R1110_U77 );
nand NAND2_26006 ( P3_R1110_U176 , P3_U3064 , P3_U3903 );
not NOT1_26007 ( P3_R1110_U177 , P3_R1110_U61 );
or OR2_26008 ( P3_R1110_U178 , P3_U3066 , P3_U3404 );
or OR2_26009 ( P3_R1110_U179 , P3_U3059 , P3_U3401 );
or OR2_26010 ( P3_R1110_U180 , P3_U3398 , P3_U3063 );
or OR2_26011 ( P3_R1110_U181 , P3_U3395 , P3_U3067 );
not NOT1_26012 ( P3_R1110_U182 , P3_R1110_U31 );
or OR2_26013 ( P3_R1110_U183 , P3_U3392 , P3_U3077 );
not NOT1_26014 ( P3_R1110_U184 , P3_R1110_U42 );
not NOT1_26015 ( P3_R1110_U185 , P3_R1110_U43 );
nand NAND2_26016 ( P3_R1110_U186 , P3_R1110_U42 , P3_R1110_U43 );
nand NAND2_26017 ( P3_R1110_U187 , P3_U3067 , P3_U3395 );
nand NAND2_26018 ( P3_R1110_U188 , P3_R1110_U186 , P3_R1110_U181 );
nand NAND2_26019 ( P3_R1110_U189 , P3_U3063 , P3_U3398 );
nand NAND2_26020 ( P3_R1110_U190 , P3_R1110_U115 , P3_R1110_U188 );
nand NAND2_26021 ( P3_R1110_U191 , P3_R1110_U35 , P3_R1110_U34 );
nand NAND2_26022 ( P3_R1110_U192 , P3_U3066 , P3_R1110_U191 );
nand NAND2_26023 ( P3_R1110_U193 , P3_R1110_U116 , P3_R1110_U190 );
nand NAND2_26024 ( P3_R1110_U194 , P3_U3404 , P3_R1110_U170 );
not NOT1_26025 ( P3_R1110_U195 , P3_R1110_U41 );
or OR2_26026 ( P3_R1110_U196 , P3_U3069 , P3_U3410 );
or OR2_26027 ( P3_R1110_U197 , P3_U3070 , P3_U3407 );
not NOT1_26028 ( P3_R1110_U198 , P3_R1110_U22 );
nand NAND2_26029 ( P3_R1110_U199 , P3_R1110_U23 , P3_R1110_U22 );
nand NAND2_26030 ( P3_R1110_U200 , P3_U3069 , P3_R1110_U199 );
nand NAND2_26031 ( P3_R1110_U201 , P3_U3410 , P3_R1110_U198 );
nand NAND2_26032 ( P3_R1110_U202 , P3_R1110_U5 , P3_R1110_U41 );
not NOT1_26033 ( P3_R1110_U203 , P3_R1110_U144 );
or OR2_26034 ( P3_R1110_U204 , P3_U3413 , P3_U3083 );
nand NAND2_26035 ( P3_R1110_U205 , P3_R1110_U204 , P3_R1110_U144 );
not NOT1_26036 ( P3_R1110_U206 , P3_R1110_U40 );
or OR2_26037 ( P3_R1110_U207 , P3_U3082 , P3_U3416 );
or OR2_26038 ( P3_R1110_U208 , P3_U3407 , P3_U3070 );
nand NAND2_26039 ( P3_R1110_U209 , P3_R1110_U208 , P3_R1110_U41 );
nand NAND2_26040 ( P3_R1110_U210 , P3_R1110_U119 , P3_R1110_U209 );
nand NAND2_26041 ( P3_R1110_U211 , P3_R1110_U195 , P3_R1110_U22 );
nand NAND2_26042 ( P3_R1110_U212 , P3_U3410 , P3_U3069 );
nand NAND2_26043 ( P3_R1110_U213 , P3_R1110_U120 , P3_R1110_U211 );
or OR2_26044 ( P3_R1110_U214 , P3_U3070 , P3_U3407 );
nand NAND2_26045 ( P3_R1110_U215 , P3_R1110_U185 , P3_R1110_U181 );
nand NAND2_26046 ( P3_R1110_U216 , P3_U3067 , P3_U3395 );
not NOT1_26047 ( P3_R1110_U217 , P3_R1110_U45 );
nand NAND2_26048 ( P3_R1110_U218 , P3_R1110_U121 , P3_R1110_U184 );
nand NAND2_26049 ( P3_R1110_U219 , P3_R1110_U45 , P3_R1110_U180 );
nand NAND2_26050 ( P3_R1110_U220 , P3_U3063 , P3_U3398 );
not NOT1_26051 ( P3_R1110_U221 , P3_R1110_U44 );
or OR2_26052 ( P3_R1110_U222 , P3_U3401 , P3_U3059 );
nand NAND2_26053 ( P3_R1110_U223 , P3_R1110_U222 , P3_R1110_U44 );
nand NAND2_26054 ( P3_R1110_U224 , P3_R1110_U123 , P3_R1110_U223 );
nand NAND2_26055 ( P3_R1110_U225 , P3_R1110_U221 , P3_R1110_U34 );
nand NAND2_26056 ( P3_R1110_U226 , P3_U3404 , P3_U3066 );
nand NAND2_26057 ( P3_R1110_U227 , P3_R1110_U124 , P3_R1110_U225 );
or OR2_26058 ( P3_R1110_U228 , P3_U3059 , P3_U3401 );
nand NAND2_26059 ( P3_R1110_U229 , P3_R1110_U184 , P3_R1110_U181 );
not NOT1_26060 ( P3_R1110_U230 , P3_R1110_U145 );
nand NAND2_26061 ( P3_R1110_U231 , P3_U3063 , P3_U3398 );
nand NAND4_26062 ( P3_R1110_U232 , P3_R1110_U401 , P3_R1110_U400 , P3_R1110_U43 , P3_R1110_U42 );
nand NAND2_26063 ( P3_R1110_U233 , P3_R1110_U43 , P3_R1110_U42 );
nand NAND2_26064 ( P3_R1110_U234 , P3_U3067 , P3_U3395 );
nand NAND2_26065 ( P3_R1110_U235 , P3_R1110_U125 , P3_R1110_U233 );
or OR2_26066 ( P3_R1110_U236 , P3_U3082 , P3_U3416 );
or OR2_26067 ( P3_R1110_U237 , P3_U3061 , P3_U3419 );
nand NAND2_26068 ( P3_R1110_U238 , P3_R1110_U177 , P3_R1110_U6 );
nand NAND2_26069 ( P3_R1110_U239 , P3_U3061 , P3_U3419 );
nand NAND2_26070 ( P3_R1110_U240 , P3_R1110_U127 , P3_R1110_U238 );
or OR2_26071 ( P3_R1110_U241 , P3_U3419 , P3_U3061 );
nand NAND2_26072 ( P3_R1110_U242 , P3_R1110_U126 , P3_R1110_U144 );
nand NAND2_26073 ( P3_R1110_U243 , P3_R1110_U241 , P3_R1110_U240 );
not NOT1_26074 ( P3_R1110_U244 , P3_R1110_U167 );
or OR2_26075 ( P3_R1110_U245 , P3_U3079 , P3_U3428 );
or OR2_26076 ( P3_R1110_U246 , P3_U3071 , P3_U3425 );
nand NAND2_26077 ( P3_R1110_U247 , P3_R1110_U174 , P3_R1110_U7 );
nand NAND2_26078 ( P3_R1110_U248 , P3_U3079 , P3_U3428 );
nand NAND2_26079 ( P3_R1110_U249 , P3_R1110_U129 , P3_R1110_U247 );
or OR2_26080 ( P3_R1110_U250 , P3_U3422 , P3_U3062 );
or OR2_26081 ( P3_R1110_U251 , P3_U3428 , P3_U3079 );
nand NAND2_26082 ( P3_R1110_U252 , P3_R1110_U128 , P3_R1110_U167 );
nand NAND2_26083 ( P3_R1110_U253 , P3_R1110_U251 , P3_R1110_U249 );
not NOT1_26084 ( P3_R1110_U254 , P3_R1110_U166 );
or OR2_26085 ( P3_R1110_U255 , P3_U3431 , P3_U3078 );
nand NAND2_26086 ( P3_R1110_U256 , P3_R1110_U255 , P3_R1110_U166 );
nand NAND2_26087 ( P3_R1110_U257 , P3_U3078 , P3_U3431 );
not NOT1_26088 ( P3_R1110_U258 , P3_R1110_U164 );
or OR2_26089 ( P3_R1110_U259 , P3_U3434 , P3_U3073 );
nand NAND2_26090 ( P3_R1110_U260 , P3_R1110_U259 , P3_R1110_U164 );
nand NAND2_26091 ( P3_R1110_U261 , P3_U3073 , P3_U3434 );
not NOT1_26092 ( P3_R1110_U262 , P3_R1110_U92 );
or OR2_26093 ( P3_R1110_U263 , P3_U3068 , P3_U3440 );
or OR2_26094 ( P3_R1110_U264 , P3_U3072 , P3_U3437 );
not NOT1_26095 ( P3_R1110_U265 , P3_R1110_U59 );
nand NAND2_26096 ( P3_R1110_U266 , P3_R1110_U60 , P3_R1110_U59 );
nand NAND2_26097 ( P3_R1110_U267 , P3_U3068 , P3_R1110_U266 );
nand NAND2_26098 ( P3_R1110_U268 , P3_U3440 , P3_R1110_U265 );
nand NAND2_26099 ( P3_R1110_U269 , P3_R1110_U8 , P3_R1110_U92 );
not NOT1_26100 ( P3_R1110_U270 , P3_R1110_U162 );
or OR2_26101 ( P3_R1110_U271 , P3_U3075 , P3_U3907 );
or OR2_26102 ( P3_R1110_U272 , P3_U3080 , P3_U3445 );
or OR2_26103 ( P3_R1110_U273 , P3_U3074 , P3_U3906 );
not NOT1_26104 ( P3_R1110_U274 , P3_R1110_U80 );
nand NAND2_26105 ( P3_R1110_U275 , P3_U3907 , P3_R1110_U274 );
nand NAND2_26106 ( P3_R1110_U276 , P3_R1110_U275 , P3_R1110_U90 );
nand NAND2_26107 ( P3_R1110_U277 , P3_R1110_U80 , P3_R1110_U81 );
nand NAND2_26108 ( P3_R1110_U278 , P3_R1110_U277 , P3_R1110_U276 );
nand NAND2_26109 ( P3_R1110_U279 , P3_R1110_U175 , P3_R1110_U9 );
nand NAND2_26110 ( P3_R1110_U280 , P3_U3074 , P3_U3906 );
nand NAND2_26111 ( P3_R1110_U281 , P3_R1110_U278 , P3_R1110_U279 );
or OR2_26112 ( P3_R1110_U282 , P3_U3443 , P3_U3081 );
or OR2_26113 ( P3_R1110_U283 , P3_U3906 , P3_U3074 );
nand NAND2_26114 ( P3_R1110_U284 , P3_R1110_U162 , P3_R1110_U131 );
nand NAND2_26115 ( P3_R1110_U285 , P3_R1110_U283 , P3_R1110_U281 );
not NOT1_26116 ( P3_R1110_U286 , P3_R1110_U159 );
or OR2_26117 ( P3_R1110_U287 , P3_U3905 , P3_U3060 );
nand NAND2_26118 ( P3_R1110_U288 , P3_R1110_U287 , P3_R1110_U159 );
nand NAND2_26119 ( P3_R1110_U289 , P3_U3060 , P3_U3905 );
not NOT1_26120 ( P3_R1110_U290 , P3_R1110_U157 );
or OR2_26121 ( P3_R1110_U291 , P3_U3904 , P3_U3065 );
nand NAND2_26122 ( P3_R1110_U292 , P3_R1110_U291 , P3_R1110_U157 );
nand NAND2_26123 ( P3_R1110_U293 , P3_U3065 , P3_U3904 );
not NOT1_26124 ( P3_R1110_U294 , P3_R1110_U155 );
or OR2_26125 ( P3_R1110_U295 , P3_U3057 , P3_U3902 );
nand NAND2_26126 ( P3_R1110_U296 , P3_R1110_U176 , P3_R1110_U173 );
not NOT1_26127 ( P3_R1110_U297 , P3_R1110_U86 );
or OR2_26128 ( P3_R1110_U298 , P3_U3903 , P3_U3064 );
nand NAND3_26129 ( P3_R1110_U299 , P3_R1110_U155 , P3_R1110_U298 , P3_R1110_U168 );
not NOT1_26130 ( P3_R1110_U300 , P3_R1110_U153 );
or OR2_26131 ( P3_R1110_U301 , P3_U3900 , P3_U3052 );
nand NAND2_26132 ( P3_R1110_U302 , P3_U3052 , P3_U3900 );
not NOT1_26133 ( P3_R1110_U303 , P3_R1110_U151 );
nand NAND2_26134 ( P3_R1110_U304 , P3_U3899 , P3_R1110_U151 );
not NOT1_26135 ( P3_R1110_U305 , P3_R1110_U149 );
nand NAND2_26136 ( P3_R1110_U306 , P3_R1110_U298 , P3_R1110_U155 );
not NOT1_26137 ( P3_R1110_U307 , P3_R1110_U89 );
or OR2_26138 ( P3_R1110_U308 , P3_U3902 , P3_U3057 );
nand NAND2_26139 ( P3_R1110_U309 , P3_R1110_U308 , P3_R1110_U89 );
nand NAND3_26140 ( P3_R1110_U310 , P3_R1110_U309 , P3_R1110_U173 , P3_R1110_U154 );
nand NAND2_26141 ( P3_R1110_U311 , P3_R1110_U307 , P3_R1110_U173 );
nand NAND2_26142 ( P3_R1110_U312 , P3_U3901 , P3_U3056 );
nand NAND3_26143 ( P3_R1110_U313 , P3_R1110_U311 , P3_R1110_U312 , P3_R1110_U168 );
or OR2_26144 ( P3_R1110_U314 , P3_U3057 , P3_U3902 );
nand NAND2_26145 ( P3_R1110_U315 , P3_R1110_U282 , P3_R1110_U162 );
not NOT1_26146 ( P3_R1110_U316 , P3_R1110_U91 );
nand NAND2_26147 ( P3_R1110_U317 , P3_R1110_U9 , P3_R1110_U91 );
nand NAND2_26148 ( P3_R1110_U318 , P3_R1110_U135 , P3_R1110_U317 );
nand NAND2_26149 ( P3_R1110_U319 , P3_R1110_U317 , P3_R1110_U278 );
nand NAND2_26150 ( P3_R1110_U320 , P3_R1110_U453 , P3_R1110_U319 );
or OR2_26151 ( P3_R1110_U321 , P3_U3445 , P3_U3080 );
nand NAND2_26152 ( P3_R1110_U322 , P3_R1110_U321 , P3_R1110_U91 );
nand NAND2_26153 ( P3_R1110_U323 , P3_R1110_U136 , P3_R1110_U322 );
nand NAND2_26154 ( P3_R1110_U324 , P3_R1110_U316 , P3_R1110_U80 );
nand NAND2_26155 ( P3_R1110_U325 , P3_U3075 , P3_U3907 );
nand NAND2_26156 ( P3_R1110_U326 , P3_R1110_U137 , P3_R1110_U324 );
or OR2_26157 ( P3_R1110_U327 , P3_U3392 , P3_U3077 );
not NOT1_26158 ( P3_R1110_U328 , P3_R1110_U161 );
or OR2_26159 ( P3_R1110_U329 , P3_U3080 , P3_U3445 );
or OR2_26160 ( P3_R1110_U330 , P3_U3437 , P3_U3072 );
nand NAND2_26161 ( P3_R1110_U331 , P3_R1110_U330 , P3_R1110_U92 );
nand NAND2_26162 ( P3_R1110_U332 , P3_R1110_U138 , P3_R1110_U331 );
nand NAND2_26163 ( P3_R1110_U333 , P3_R1110_U262 , P3_R1110_U59 );
nand NAND2_26164 ( P3_R1110_U334 , P3_U3440 , P3_U3068 );
nand NAND2_26165 ( P3_R1110_U335 , P3_R1110_U139 , P3_R1110_U333 );
or OR2_26166 ( P3_R1110_U336 , P3_U3072 , P3_U3437 );
nand NAND2_26167 ( P3_R1110_U337 , P3_R1110_U250 , P3_R1110_U167 );
not NOT1_26168 ( P3_R1110_U338 , P3_R1110_U93 );
or OR2_26169 ( P3_R1110_U339 , P3_U3425 , P3_U3071 );
nand NAND2_26170 ( P3_R1110_U340 , P3_R1110_U339 , P3_R1110_U93 );
nand NAND2_26171 ( P3_R1110_U341 , P3_R1110_U140 , P3_R1110_U340 );
nand NAND2_26172 ( P3_R1110_U342 , P3_R1110_U338 , P3_R1110_U172 );
nand NAND2_26173 ( P3_R1110_U343 , P3_U3079 , P3_U3428 );
nand NAND2_26174 ( P3_R1110_U344 , P3_R1110_U141 , P3_R1110_U342 );
or OR2_26175 ( P3_R1110_U345 , P3_U3071 , P3_U3425 );
or OR2_26176 ( P3_R1110_U346 , P3_U3416 , P3_U3082 );
nand NAND2_26177 ( P3_R1110_U347 , P3_R1110_U346 , P3_R1110_U40 );
nand NAND2_26178 ( P3_R1110_U348 , P3_R1110_U142 , P3_R1110_U347 );
nand NAND2_26179 ( P3_R1110_U349 , P3_R1110_U206 , P3_R1110_U171 );
nand NAND2_26180 ( P3_R1110_U350 , P3_U3061 , P3_U3419 );
nand NAND2_26181 ( P3_R1110_U351 , P3_R1110_U143 , P3_R1110_U349 );
nand NAND2_26182 ( P3_R1110_U352 , P3_R1110_U207 , P3_R1110_U171 );
nand NAND2_26183 ( P3_R1110_U353 , P3_R1110_U204 , P3_R1110_U61 );
nand NAND2_26184 ( P3_R1110_U354 , P3_R1110_U214 , P3_R1110_U22 );
nand NAND2_26185 ( P3_R1110_U355 , P3_R1110_U228 , P3_R1110_U34 );
nand NAND2_26186 ( P3_R1110_U356 , P3_R1110_U231 , P3_R1110_U180 );
nand NAND2_26187 ( P3_R1110_U357 , P3_R1110_U314 , P3_R1110_U173 );
nand NAND2_26188 ( P3_R1110_U358 , P3_R1110_U298 , P3_R1110_U176 );
nand NAND2_26189 ( P3_R1110_U359 , P3_R1110_U329 , P3_R1110_U80 );
nand NAND2_26190 ( P3_R1110_U360 , P3_R1110_U282 , P3_R1110_U77 );
nand NAND2_26191 ( P3_R1110_U361 , P3_R1110_U336 , P3_R1110_U59 );
nand NAND2_26192 ( P3_R1110_U362 , P3_R1110_U345 , P3_R1110_U172 );
nand NAND2_26193 ( P3_R1110_U363 , P3_R1110_U250 , P3_R1110_U68 );
nand NAND2_26194 ( P3_R1110_U364 , P3_U3899 , P3_U3053 );
nand NAND2_26195 ( P3_R1110_U365 , P3_R1110_U296 , P3_R1110_U168 );
nand NAND2_26196 ( P3_R1110_U366 , P3_U3056 , P3_R1110_U295 );
nand NAND2_26197 ( P3_R1110_U367 , P3_U3901 , P3_R1110_U295 );
nand NAND3_26198 ( P3_R1110_U368 , P3_R1110_U296 , P3_R1110_U168 , P3_R1110_U301 );
nand NAND3_26199 ( P3_R1110_U369 , P3_R1110_U155 , P3_R1110_U168 , P3_R1110_U133 );
nand NAND2_26200 ( P3_R1110_U370 , P3_R1110_U297 , P3_R1110_U301 );
nand NAND2_26201 ( P3_R1110_U371 , P3_U3082 , P3_R1110_U39 );
nand NAND2_26202 ( P3_R1110_U372 , P3_U3416 , P3_R1110_U38 );
nand NAND2_26203 ( P3_R1110_U373 , P3_R1110_U372 , P3_R1110_U371 );
nand NAND2_26204 ( P3_R1110_U374 , P3_R1110_U352 , P3_R1110_U40 );
nand NAND2_26205 ( P3_R1110_U375 , P3_R1110_U373 , P3_R1110_U206 );
nand NAND2_26206 ( P3_R1110_U376 , P3_U3083 , P3_R1110_U36 );
nand NAND2_26207 ( P3_R1110_U377 , P3_U3413 , P3_R1110_U37 );
nand NAND2_26208 ( P3_R1110_U378 , P3_R1110_U377 , P3_R1110_U376 );
nand NAND2_26209 ( P3_R1110_U379 , P3_R1110_U353 , P3_R1110_U144 );
nand NAND2_26210 ( P3_R1110_U380 , P3_R1110_U203 , P3_R1110_U378 );
nand NAND2_26211 ( P3_R1110_U381 , P3_U3069 , P3_R1110_U23 );
nand NAND2_26212 ( P3_R1110_U382 , P3_U3410 , P3_R1110_U21 );
nand NAND2_26213 ( P3_R1110_U383 , P3_U3070 , P3_R1110_U19 );
nand NAND2_26214 ( P3_R1110_U384 , P3_U3407 , P3_R1110_U20 );
nand NAND2_26215 ( P3_R1110_U385 , P3_R1110_U384 , P3_R1110_U383 );
nand NAND2_26216 ( P3_R1110_U386 , P3_R1110_U354 , P3_R1110_U41 );
nand NAND2_26217 ( P3_R1110_U387 , P3_R1110_U385 , P3_R1110_U195 );
nand NAND2_26218 ( P3_R1110_U388 , P3_U3066 , P3_R1110_U35 );
nand NAND2_26219 ( P3_R1110_U389 , P3_U3404 , P3_R1110_U26 );
nand NAND2_26220 ( P3_R1110_U390 , P3_U3059 , P3_R1110_U24 );
nand NAND2_26221 ( P3_R1110_U391 , P3_U3401 , P3_R1110_U25 );
nand NAND2_26222 ( P3_R1110_U392 , P3_R1110_U391 , P3_R1110_U390 );
nand NAND2_26223 ( P3_R1110_U393 , P3_R1110_U355 , P3_R1110_U44 );
nand NAND2_26224 ( P3_R1110_U394 , P3_R1110_U392 , P3_R1110_U221 );
nand NAND2_26225 ( P3_R1110_U395 , P3_U3063 , P3_R1110_U32 );
nand NAND2_26226 ( P3_R1110_U396 , P3_U3398 , P3_R1110_U33 );
nand NAND2_26227 ( P3_R1110_U397 , P3_R1110_U396 , P3_R1110_U395 );
nand NAND2_26228 ( P3_R1110_U398 , P3_R1110_U356 , P3_R1110_U145 );
nand NAND2_26229 ( P3_R1110_U399 , P3_R1110_U230 , P3_R1110_U397 );
nand NAND2_26230 ( P3_R1110_U400 , P3_U3067 , P3_R1110_U27 );
nand NAND2_26231 ( P3_R1110_U401 , P3_U3395 , P3_R1110_U28 );
nand NAND2_26232 ( P3_R1110_U402 , P3_U3054 , P3_R1110_U147 );
nand NAND2_26233 ( P3_R1110_U403 , P3_U3908 , P3_R1110_U146 );
nand NAND2_26234 ( P3_R1110_U404 , P3_U3054 , P3_R1110_U147 );
nand NAND2_26235 ( P3_R1110_U405 , P3_U3908 , P3_R1110_U146 );
nand NAND2_26236 ( P3_R1110_U406 , P3_R1110_U405 , P3_R1110_U404 );
nand NAND2_26237 ( P3_R1110_U407 , P3_R1110_U148 , P3_R1110_U149 );
nand NAND2_26238 ( P3_R1110_U408 , P3_R1110_U305 , P3_R1110_U406 );
nand NAND2_26239 ( P3_R1110_U409 , P3_U3053 , P3_R1110_U88 );
nand NAND2_26240 ( P3_R1110_U410 , P3_U3899 , P3_R1110_U87 );
nand NAND2_26241 ( P3_R1110_U411 , P3_U3053 , P3_R1110_U88 );
nand NAND2_26242 ( P3_R1110_U412 , P3_U3899 , P3_R1110_U87 );
nand NAND2_26243 ( P3_R1110_U413 , P3_R1110_U412 , P3_R1110_U411 );
nand NAND2_26244 ( P3_R1110_U414 , P3_R1110_U150 , P3_R1110_U151 );
nand NAND2_26245 ( P3_R1110_U415 , P3_R1110_U303 , P3_R1110_U413 );
nand NAND2_26246 ( P3_R1110_U416 , P3_U3052 , P3_R1110_U46 );
nand NAND2_26247 ( P3_R1110_U417 , P3_U3900 , P3_R1110_U47 );
nand NAND2_26248 ( P3_R1110_U418 , P3_U3052 , P3_R1110_U46 );
nand NAND2_26249 ( P3_R1110_U419 , P3_U3900 , P3_R1110_U47 );
nand NAND2_26250 ( P3_R1110_U420 , P3_R1110_U419 , P3_R1110_U418 );
nand NAND2_26251 ( P3_R1110_U421 , P3_R1110_U152 , P3_R1110_U153 );
nand NAND2_26252 ( P3_R1110_U422 , P3_R1110_U300 , P3_R1110_U420 );
nand NAND2_26253 ( P3_R1110_U423 , P3_U3056 , P3_R1110_U49 );
nand NAND2_26254 ( P3_R1110_U424 , P3_U3901 , P3_R1110_U48 );
nand NAND2_26255 ( P3_R1110_U425 , P3_U3057 , P3_R1110_U50 );
nand NAND2_26256 ( P3_R1110_U426 , P3_U3902 , P3_R1110_U51 );
nand NAND2_26257 ( P3_R1110_U427 , P3_R1110_U426 , P3_R1110_U425 );
nand NAND2_26258 ( P3_R1110_U428 , P3_R1110_U357 , P3_R1110_U89 );
nand NAND2_26259 ( P3_R1110_U429 , P3_R1110_U427 , P3_R1110_U307 );
nand NAND2_26260 ( P3_R1110_U430 , P3_U3064 , P3_R1110_U52 );
nand NAND2_26261 ( P3_R1110_U431 , P3_U3903 , P3_R1110_U53 );
nand NAND2_26262 ( P3_R1110_U432 , P3_R1110_U431 , P3_R1110_U430 );
nand NAND2_26263 ( P3_R1110_U433 , P3_R1110_U358 , P3_R1110_U155 );
nand NAND2_26264 ( P3_R1110_U434 , P3_R1110_U294 , P3_R1110_U432 );
nand NAND2_26265 ( P3_R1110_U435 , P3_U3065 , P3_R1110_U84 );
nand NAND2_26266 ( P3_R1110_U436 , P3_U3904 , P3_R1110_U85 );
nand NAND2_26267 ( P3_R1110_U437 , P3_U3065 , P3_R1110_U84 );
nand NAND2_26268 ( P3_R1110_U438 , P3_U3904 , P3_R1110_U85 );
nand NAND2_26269 ( P3_R1110_U439 , P3_R1110_U438 , P3_R1110_U437 );
nand NAND2_26270 ( P3_R1110_U440 , P3_R1110_U156 , P3_R1110_U157 );
nand NAND2_26271 ( P3_R1110_U441 , P3_R1110_U290 , P3_R1110_U439 );
nand NAND2_26272 ( P3_R1110_U442 , P3_U3060 , P3_R1110_U82 );
nand NAND2_26273 ( P3_R1110_U443 , P3_U3905 , P3_R1110_U83 );
nand NAND2_26274 ( P3_R1110_U444 , P3_U3060 , P3_R1110_U82 );
nand NAND2_26275 ( P3_R1110_U445 , P3_U3905 , P3_R1110_U83 );
nand NAND2_26276 ( P3_R1110_U446 , P3_R1110_U445 , P3_R1110_U444 );
nand NAND2_26277 ( P3_R1110_U447 , P3_R1110_U158 , P3_R1110_U159 );
nand NAND2_26278 ( P3_R1110_U448 , P3_R1110_U286 , P3_R1110_U446 );
nand NAND2_26279 ( P3_R1110_U449 , P3_U3074 , P3_R1110_U54 );
nand NAND2_26280 ( P3_R1110_U450 , P3_U3906 , P3_R1110_U55 );
nand NAND2_26281 ( P3_R1110_U451 , P3_U3074 , P3_R1110_U54 );
nand NAND2_26282 ( P3_R1110_U452 , P3_U3906 , P3_R1110_U55 );
nand NAND2_26283 ( P3_R1110_U453 , P3_R1110_U452 , P3_R1110_U451 );
nand NAND2_26284 ( P3_R1110_U454 , P3_U3075 , P3_R1110_U81 );
nand NAND2_26285 ( P3_R1110_U455 , P3_U3907 , P3_R1110_U90 );
nand NAND2_26286 ( P3_R1110_U456 , P3_R1110_U182 , P3_R1110_U161 );
nand NAND2_26287 ( P3_R1110_U457 , P3_R1110_U328 , P3_R1110_U31 );
nand NAND2_26288 ( P3_R1110_U458 , P3_U3080 , P3_R1110_U78 );
nand NAND2_26289 ( P3_R1110_U459 , P3_U3445 , P3_R1110_U79 );
nand NAND2_26290 ( P3_R1110_U460 , P3_R1110_U459 , P3_R1110_U458 );
nand NAND2_26291 ( P3_R1110_U461 , P3_R1110_U359 , P3_R1110_U91 );
nand NAND2_26292 ( P3_R1110_U462 , P3_R1110_U460 , P3_R1110_U316 );
nand NAND2_26293 ( P3_R1110_U463 , P3_U3081 , P3_R1110_U75 );
nand NAND2_26294 ( P3_R1110_U464 , P3_U3443 , P3_R1110_U76 );
nand NAND2_26295 ( P3_R1110_U465 , P3_R1110_U464 , P3_R1110_U463 );
nand NAND2_26296 ( P3_R1110_U466 , P3_R1110_U360 , P3_R1110_U162 );
nand NAND2_26297 ( P3_R1110_U467 , P3_R1110_U270 , P3_R1110_U465 );
nand NAND2_26298 ( P3_R1110_U468 , P3_U3068 , P3_R1110_U60 );
nand NAND2_26299 ( P3_R1110_U469 , P3_U3440 , P3_R1110_U58 );
nand NAND2_26300 ( P3_R1110_U470 , P3_U3072 , P3_R1110_U56 );
nand NAND2_26301 ( P3_R1110_U471 , P3_U3437 , P3_R1110_U57 );
nand NAND2_26302 ( P3_R1110_U472 , P3_R1110_U471 , P3_R1110_U470 );
nand NAND2_26303 ( P3_R1110_U473 , P3_R1110_U361 , P3_R1110_U92 );
nand NAND2_26304 ( P3_R1110_U474 , P3_R1110_U472 , P3_R1110_U262 );
nand NAND2_26305 ( P3_R1110_U475 , P3_U3073 , P3_R1110_U73 );
nand NAND2_26306 ( P3_R1110_U476 , P3_U3434 , P3_R1110_U74 );
nand NAND2_26307 ( P3_R1110_U477 , P3_U3073 , P3_R1110_U73 );
nand NAND2_26308 ( P3_R1110_U478 , P3_U3434 , P3_R1110_U74 );
nand NAND2_26309 ( P3_R1110_U479 , P3_R1110_U478 , P3_R1110_U477 );
nand NAND2_26310 ( P3_R1110_U480 , P3_R1110_U163 , P3_R1110_U164 );
nand NAND2_26311 ( P3_R1110_U481 , P3_R1110_U258 , P3_R1110_U479 );
nand NAND2_26312 ( P3_R1110_U482 , P3_U3078 , P3_R1110_U71 );
nand NAND2_26313 ( P3_R1110_U483 , P3_U3431 , P3_R1110_U72 );
nand NAND2_26314 ( P3_R1110_U484 , P3_U3078 , P3_R1110_U71 );
nand NAND2_26315 ( P3_R1110_U485 , P3_U3431 , P3_R1110_U72 );
nand NAND2_26316 ( P3_R1110_U486 , P3_R1110_U485 , P3_R1110_U484 );
nand NAND2_26317 ( P3_R1110_U487 , P3_R1110_U165 , P3_R1110_U166 );
nand NAND2_26318 ( P3_R1110_U488 , P3_R1110_U254 , P3_R1110_U486 );
nand NAND2_26319 ( P3_R1110_U489 , P3_U3079 , P3_R1110_U69 );
nand NAND2_26320 ( P3_R1110_U490 , P3_U3428 , P3_R1110_U70 );
nand NAND2_26321 ( P3_R1110_U491 , P3_U3071 , P3_R1110_U64 );
nand NAND2_26322 ( P3_R1110_U492 , P3_U3425 , P3_R1110_U65 );
nand NAND2_26323 ( P3_R1110_U493 , P3_R1110_U492 , P3_R1110_U491 );
nand NAND2_26324 ( P3_R1110_U494 , P3_R1110_U362 , P3_R1110_U93 );
nand NAND2_26325 ( P3_R1110_U495 , P3_R1110_U493 , P3_R1110_U338 );
nand NAND2_26326 ( P3_R1110_U496 , P3_U3062 , P3_R1110_U66 );
nand NAND2_26327 ( P3_R1110_U497 , P3_U3422 , P3_R1110_U67 );
nand NAND2_26328 ( P3_R1110_U498 , P3_R1110_U497 , P3_R1110_U496 );
nand NAND2_26329 ( P3_R1110_U499 , P3_R1110_U363 , P3_R1110_U167 );
nand NAND2_26330 ( P3_R1110_U500 , P3_R1110_U244 , P3_R1110_U498 );
nand NAND2_26331 ( P3_R1110_U501 , P3_U3061 , P3_R1110_U62 );
nand NAND2_26332 ( P3_R1110_U502 , P3_U3419 , P3_R1110_U63 );
nand NAND2_26333 ( P3_R1110_U503 , P3_U3076 , P3_R1110_U29 );
nand NAND2_26334 ( P3_R1110_U504 , P3_U3387 , P3_R1110_U30 );
and AND2_26335 ( P3_R1297_U6 , P3_U3058 , P3_R1297_U7 );
not NOT1_26336 ( P3_R1297_U7 , P3_U3055 );
and AND2_26337 ( P3_R1077_U4 , P3_R1077_U179 , P3_R1077_U178 );
and AND2_26338 ( P3_R1077_U5 , P3_R1077_U197 , P3_R1077_U196 );
and AND2_26339 ( P3_R1077_U6 , P3_R1077_U237 , P3_R1077_U236 );
and AND2_26340 ( P3_R1077_U7 , P3_R1077_U246 , P3_R1077_U245 );
and AND2_26341 ( P3_R1077_U8 , P3_R1077_U264 , P3_R1077_U263 );
and AND2_26342 ( P3_R1077_U9 , P3_R1077_U272 , P3_R1077_U271 );
and AND2_26343 ( P3_R1077_U10 , P3_R1077_U351 , P3_R1077_U348 );
and AND2_26344 ( P3_R1077_U11 , P3_R1077_U344 , P3_R1077_U341 );
and AND2_26345 ( P3_R1077_U12 , P3_R1077_U335 , P3_R1077_U332 );
and AND2_26346 ( P3_R1077_U13 , P3_R1077_U326 , P3_R1077_U323 );
and AND2_26347 ( P3_R1077_U14 , P3_R1077_U320 , P3_R1077_U318 );
and AND2_26348 ( P3_R1077_U15 , P3_R1077_U313 , P3_R1077_U310 );
and AND2_26349 ( P3_R1077_U16 , P3_R1077_U235 , P3_R1077_U232 );
and AND2_26350 ( P3_R1077_U17 , P3_R1077_U227 , P3_R1077_U224 );
and AND2_26351 ( P3_R1077_U18 , P3_R1077_U213 , P3_R1077_U210 );
not NOT1_26352 ( P3_R1077_U19 , P3_U3407 );
not NOT1_26353 ( P3_R1077_U20 , P3_U3070 );
not NOT1_26354 ( P3_R1077_U21 , P3_U3069 );
nand NAND2_26355 ( P3_R1077_U22 , P3_U3070 , P3_U3407 );
not NOT1_26356 ( P3_R1077_U23 , P3_U3410 );
not NOT1_26357 ( P3_R1077_U24 , P3_U3401 );
not NOT1_26358 ( P3_R1077_U25 , P3_U3059 );
not NOT1_26359 ( P3_R1077_U26 , P3_U3066 );
not NOT1_26360 ( P3_R1077_U27 , P3_U3395 );
not NOT1_26361 ( P3_R1077_U28 , P3_U3067 );
not NOT1_26362 ( P3_R1077_U29 , P3_U3387 );
not NOT1_26363 ( P3_R1077_U30 , P3_U3076 );
nand NAND2_26364 ( P3_R1077_U31 , P3_U3076 , P3_U3387 );
not NOT1_26365 ( P3_R1077_U32 , P3_U3398 );
not NOT1_26366 ( P3_R1077_U33 , P3_U3063 );
nand NAND2_26367 ( P3_R1077_U34 , P3_U3059 , P3_U3401 );
not NOT1_26368 ( P3_R1077_U35 , P3_U3404 );
not NOT1_26369 ( P3_R1077_U36 , P3_U3413 );
not NOT1_26370 ( P3_R1077_U37 , P3_U3083 );
not NOT1_26371 ( P3_R1077_U38 , P3_U3082 );
not NOT1_26372 ( P3_R1077_U39 , P3_U3416 );
nand NAND2_26373 ( P3_R1077_U40 , P3_R1077_U61 , P3_R1077_U205 );
nand NAND2_26374 ( P3_R1077_U41 , P3_R1077_U117 , P3_R1077_U193 );
nand NAND2_26375 ( P3_R1077_U42 , P3_R1077_U182 , P3_R1077_U183 );
nand NAND2_26376 ( P3_R1077_U43 , P3_U3392 , P3_U3077 );
nand NAND2_26377 ( P3_R1077_U44 , P3_R1077_U122 , P3_R1077_U219 );
nand NAND2_26378 ( P3_R1077_U45 , P3_R1077_U216 , P3_R1077_U215 );
not NOT1_26379 ( P3_R1077_U46 , P3_U3900 );
not NOT1_26380 ( P3_R1077_U47 , P3_U3052 );
not NOT1_26381 ( P3_R1077_U48 , P3_U3056 );
not NOT1_26382 ( P3_R1077_U49 , P3_U3901 );
not NOT1_26383 ( P3_R1077_U50 , P3_U3902 );
not NOT1_26384 ( P3_R1077_U51 , P3_U3057 );
not NOT1_26385 ( P3_R1077_U52 , P3_U3903 );
not NOT1_26386 ( P3_R1077_U53 , P3_U3064 );
not NOT1_26387 ( P3_R1077_U54 , P3_U3906 );
not NOT1_26388 ( P3_R1077_U55 , P3_U3074 );
not NOT1_26389 ( P3_R1077_U56 , P3_U3437 );
not NOT1_26390 ( P3_R1077_U57 , P3_U3072 );
not NOT1_26391 ( P3_R1077_U58 , P3_U3068 );
nand NAND2_26392 ( P3_R1077_U59 , P3_U3072 , P3_U3437 );
not NOT1_26393 ( P3_R1077_U60 , P3_U3440 );
nand NAND2_26394 ( P3_R1077_U61 , P3_U3083 , P3_U3413 );
not NOT1_26395 ( P3_R1077_U62 , P3_U3419 );
not NOT1_26396 ( P3_R1077_U63 , P3_U3061 );
not NOT1_26397 ( P3_R1077_U64 , P3_U3425 );
not NOT1_26398 ( P3_R1077_U65 , P3_U3071 );
not NOT1_26399 ( P3_R1077_U66 , P3_U3422 );
not NOT1_26400 ( P3_R1077_U67 , P3_U3062 );
nand NAND2_26401 ( P3_R1077_U68 , P3_U3062 , P3_U3422 );
not NOT1_26402 ( P3_R1077_U69 , P3_U3428 );
not NOT1_26403 ( P3_R1077_U70 , P3_U3079 );
not NOT1_26404 ( P3_R1077_U71 , P3_U3431 );
not NOT1_26405 ( P3_R1077_U72 , P3_U3078 );
not NOT1_26406 ( P3_R1077_U73 , P3_U3434 );
not NOT1_26407 ( P3_R1077_U74 , P3_U3073 );
not NOT1_26408 ( P3_R1077_U75 , P3_U3443 );
not NOT1_26409 ( P3_R1077_U76 , P3_U3081 );
nand NAND2_26410 ( P3_R1077_U77 , P3_U3081 , P3_U3443 );
not NOT1_26411 ( P3_R1077_U78 , P3_U3445 );
not NOT1_26412 ( P3_R1077_U79 , P3_U3080 );
nand NAND2_26413 ( P3_R1077_U80 , P3_U3080 , P3_U3445 );
not NOT1_26414 ( P3_R1077_U81 , P3_U3907 );
not NOT1_26415 ( P3_R1077_U82 , P3_U3905 );
not NOT1_26416 ( P3_R1077_U83 , P3_U3060 );
not NOT1_26417 ( P3_R1077_U84 , P3_U3904 );
not NOT1_26418 ( P3_R1077_U85 , P3_U3065 );
nand NAND2_26419 ( P3_R1077_U86 , P3_U3901 , P3_U3056 );
not NOT1_26420 ( P3_R1077_U87 , P3_U3053 );
not NOT1_26421 ( P3_R1077_U88 , P3_U3899 );
nand NAND2_26422 ( P3_R1077_U89 , P3_R1077_U306 , P3_R1077_U176 );
not NOT1_26423 ( P3_R1077_U90 , P3_U3075 );
nand NAND2_26424 ( P3_R1077_U91 , P3_R1077_U77 , P3_R1077_U315 );
nand NAND2_26425 ( P3_R1077_U92 , P3_R1077_U261 , P3_R1077_U260 );
nand NAND2_26426 ( P3_R1077_U93 , P3_R1077_U68 , P3_R1077_U337 );
nand NAND2_26427 ( P3_R1077_U94 , P3_R1077_U457 , P3_R1077_U456 );
nand NAND2_26428 ( P3_R1077_U95 , P3_R1077_U504 , P3_R1077_U503 );
nand NAND2_26429 ( P3_R1077_U96 , P3_R1077_U375 , P3_R1077_U374 );
nand NAND2_26430 ( P3_R1077_U97 , P3_R1077_U380 , P3_R1077_U379 );
nand NAND2_26431 ( P3_R1077_U98 , P3_R1077_U387 , P3_R1077_U386 );
nand NAND2_26432 ( P3_R1077_U99 , P3_R1077_U394 , P3_R1077_U393 );
nand NAND2_26433 ( P3_R1077_U100 , P3_R1077_U399 , P3_R1077_U398 );
nand NAND2_26434 ( P3_R1077_U101 , P3_R1077_U408 , P3_R1077_U407 );
nand NAND2_26435 ( P3_R1077_U102 , P3_R1077_U415 , P3_R1077_U414 );
nand NAND2_26436 ( P3_R1077_U103 , P3_R1077_U422 , P3_R1077_U421 );
nand NAND2_26437 ( P3_R1077_U104 , P3_R1077_U429 , P3_R1077_U428 );
nand NAND2_26438 ( P3_R1077_U105 , P3_R1077_U434 , P3_R1077_U433 );
nand NAND2_26439 ( P3_R1077_U106 , P3_R1077_U441 , P3_R1077_U440 );
nand NAND2_26440 ( P3_R1077_U107 , P3_R1077_U448 , P3_R1077_U447 );
nand NAND2_26441 ( P3_R1077_U108 , P3_R1077_U462 , P3_R1077_U461 );
nand NAND2_26442 ( P3_R1077_U109 , P3_R1077_U467 , P3_R1077_U466 );
nand NAND2_26443 ( P3_R1077_U110 , P3_R1077_U474 , P3_R1077_U473 );
nand NAND2_26444 ( P3_R1077_U111 , P3_R1077_U481 , P3_R1077_U480 );
nand NAND2_26445 ( P3_R1077_U112 , P3_R1077_U488 , P3_R1077_U487 );
nand NAND2_26446 ( P3_R1077_U113 , P3_R1077_U495 , P3_R1077_U494 );
nand NAND2_26447 ( P3_R1077_U114 , P3_R1077_U500 , P3_R1077_U499 );
and AND2_26448 ( P3_R1077_U115 , P3_R1077_U189 , P3_R1077_U187 );
and AND2_26449 ( P3_R1077_U116 , P3_R1077_U4 , P3_R1077_U180 );
and AND2_26450 ( P3_R1077_U117 , P3_R1077_U194 , P3_R1077_U192 );
and AND2_26451 ( P3_R1077_U118 , P3_R1077_U201 , P3_R1077_U200 );
and AND3_26452 ( P3_R1077_U119 , P3_R1077_U382 , P3_R1077_U381 , P3_R1077_U22 );
and AND2_26453 ( P3_R1077_U120 , P3_R1077_U212 , P3_R1077_U5 );
and AND2_26454 ( P3_R1077_U121 , P3_R1077_U181 , P3_R1077_U180 );
and AND2_26455 ( P3_R1077_U122 , P3_R1077_U220 , P3_R1077_U218 );
and AND3_26456 ( P3_R1077_U123 , P3_R1077_U389 , P3_R1077_U388 , P3_R1077_U34 );
and AND2_26457 ( P3_R1077_U124 , P3_R1077_U226 , P3_R1077_U4 );
and AND2_26458 ( P3_R1077_U125 , P3_R1077_U234 , P3_R1077_U181 );
and AND2_26459 ( P3_R1077_U126 , P3_R1077_U204 , P3_R1077_U6 );
and AND2_26460 ( P3_R1077_U127 , P3_R1077_U239 , P3_R1077_U171 );
and AND2_26461 ( P3_R1077_U128 , P3_R1077_U250 , P3_R1077_U7 );
and AND2_26462 ( P3_R1077_U129 , P3_R1077_U248 , P3_R1077_U172 );
and AND2_26463 ( P3_R1077_U130 , P3_R1077_U268 , P3_R1077_U267 );
and AND3_26464 ( P3_R1077_U131 , P3_R1077_U9 , P3_R1077_U282 , P3_R1077_U273 );
and AND2_26465 ( P3_R1077_U132 , P3_R1077_U285 , P3_R1077_U280 );
and AND2_26466 ( P3_R1077_U133 , P3_R1077_U301 , P3_R1077_U298 );
and AND2_26467 ( P3_R1077_U134 , P3_R1077_U368 , P3_R1077_U302 );
and AND2_26468 ( P3_R1077_U135 , P3_R1077_U160 , P3_R1077_U278 );
and AND3_26469 ( P3_R1077_U136 , P3_R1077_U455 , P3_R1077_U454 , P3_R1077_U80 );
and AND2_26470 ( P3_R1077_U137 , P3_R1077_U325 , P3_R1077_U9 );
and AND3_26471 ( P3_R1077_U138 , P3_R1077_U469 , P3_R1077_U468 , P3_R1077_U59 );
and AND2_26472 ( P3_R1077_U139 , P3_R1077_U334 , P3_R1077_U8 );
and AND3_26473 ( P3_R1077_U140 , P3_R1077_U490 , P3_R1077_U489 , P3_R1077_U172 );
and AND2_26474 ( P3_R1077_U141 , P3_R1077_U343 , P3_R1077_U7 );
and AND3_26475 ( P3_R1077_U142 , P3_R1077_U502 , P3_R1077_U501 , P3_R1077_U171 );
and AND2_26476 ( P3_R1077_U143 , P3_R1077_U350 , P3_R1077_U6 );
nand NAND2_26477 ( P3_R1077_U144 , P3_R1077_U118 , P3_R1077_U202 );
nand NAND2_26478 ( P3_R1077_U145 , P3_R1077_U217 , P3_R1077_U229 );
not NOT1_26479 ( P3_R1077_U146 , P3_U3054 );
not NOT1_26480 ( P3_R1077_U147 , P3_U3908 );
and AND2_26481 ( P3_R1077_U148 , P3_R1077_U403 , P3_R1077_U402 );
nand NAND3_26482 ( P3_R1077_U149 , P3_R1077_U304 , P3_R1077_U169 , P3_R1077_U364 );
and AND2_26483 ( P3_R1077_U150 , P3_R1077_U410 , P3_R1077_U409 );
nand NAND3_26484 ( P3_R1077_U151 , P3_R1077_U370 , P3_R1077_U369 , P3_R1077_U134 );
and AND2_26485 ( P3_R1077_U152 , P3_R1077_U417 , P3_R1077_U416 );
nand NAND3_26486 ( P3_R1077_U153 , P3_R1077_U365 , P3_R1077_U299 , P3_R1077_U86 );
and AND2_26487 ( P3_R1077_U154 , P3_R1077_U424 , P3_R1077_U423 );
nand NAND2_26488 ( P3_R1077_U155 , P3_R1077_U293 , P3_R1077_U292 );
and AND2_26489 ( P3_R1077_U156 , P3_R1077_U436 , P3_R1077_U435 );
nand NAND2_26490 ( P3_R1077_U157 , P3_R1077_U289 , P3_R1077_U288 );
and AND2_26491 ( P3_R1077_U158 , P3_R1077_U443 , P3_R1077_U442 );
nand NAND2_26492 ( P3_R1077_U159 , P3_R1077_U132 , P3_R1077_U284 );
and AND2_26493 ( P3_R1077_U160 , P3_R1077_U450 , P3_R1077_U449 );
nand NAND2_26494 ( P3_R1077_U161 , P3_R1077_U43 , P3_R1077_U327 );
nand NAND2_26495 ( P3_R1077_U162 , P3_R1077_U130 , P3_R1077_U269 );
and AND2_26496 ( P3_R1077_U163 , P3_R1077_U476 , P3_R1077_U475 );
nand NAND2_26497 ( P3_R1077_U164 , P3_R1077_U257 , P3_R1077_U256 );
and AND2_26498 ( P3_R1077_U165 , P3_R1077_U483 , P3_R1077_U482 );
nand NAND2_26499 ( P3_R1077_U166 , P3_R1077_U253 , P3_R1077_U252 );
nand NAND2_26500 ( P3_R1077_U167 , P3_R1077_U243 , P3_R1077_U242 );
nand NAND2_26501 ( P3_R1077_U168 , P3_R1077_U367 , P3_R1077_U366 );
nand NAND2_26502 ( P3_R1077_U169 , P3_U3053 , P3_R1077_U151 );
not NOT1_26503 ( P3_R1077_U170 , P3_R1077_U34 );
nand NAND2_26504 ( P3_R1077_U171 , P3_U3416 , P3_U3082 );
nand NAND2_26505 ( P3_R1077_U172 , P3_U3071 , P3_U3425 );
nand NAND2_26506 ( P3_R1077_U173 , P3_U3057 , P3_U3902 );
not NOT1_26507 ( P3_R1077_U174 , P3_R1077_U68 );
not NOT1_26508 ( P3_R1077_U175 , P3_R1077_U77 );
nand NAND2_26509 ( P3_R1077_U176 , P3_U3064 , P3_U3903 );
not NOT1_26510 ( P3_R1077_U177 , P3_R1077_U61 );
or OR2_26511 ( P3_R1077_U178 , P3_U3066 , P3_U3404 );
or OR2_26512 ( P3_R1077_U179 , P3_U3059 , P3_U3401 );
or OR2_26513 ( P3_R1077_U180 , P3_U3398 , P3_U3063 );
or OR2_26514 ( P3_R1077_U181 , P3_U3395 , P3_U3067 );
not NOT1_26515 ( P3_R1077_U182 , P3_R1077_U31 );
or OR2_26516 ( P3_R1077_U183 , P3_U3392 , P3_U3077 );
not NOT1_26517 ( P3_R1077_U184 , P3_R1077_U42 );
not NOT1_26518 ( P3_R1077_U185 , P3_R1077_U43 );
nand NAND2_26519 ( P3_R1077_U186 , P3_R1077_U42 , P3_R1077_U43 );
nand NAND2_26520 ( P3_R1077_U187 , P3_U3067 , P3_U3395 );
nand NAND2_26521 ( P3_R1077_U188 , P3_R1077_U186 , P3_R1077_U181 );
nand NAND2_26522 ( P3_R1077_U189 , P3_U3063 , P3_U3398 );
nand NAND2_26523 ( P3_R1077_U190 , P3_R1077_U115 , P3_R1077_U188 );
nand NAND2_26524 ( P3_R1077_U191 , P3_R1077_U35 , P3_R1077_U34 );
nand NAND2_26525 ( P3_R1077_U192 , P3_U3066 , P3_R1077_U191 );
nand NAND2_26526 ( P3_R1077_U193 , P3_R1077_U116 , P3_R1077_U190 );
nand NAND2_26527 ( P3_R1077_U194 , P3_U3404 , P3_R1077_U170 );
not NOT1_26528 ( P3_R1077_U195 , P3_R1077_U41 );
or OR2_26529 ( P3_R1077_U196 , P3_U3069 , P3_U3410 );
or OR2_26530 ( P3_R1077_U197 , P3_U3070 , P3_U3407 );
not NOT1_26531 ( P3_R1077_U198 , P3_R1077_U22 );
nand NAND2_26532 ( P3_R1077_U199 , P3_R1077_U23 , P3_R1077_U22 );
nand NAND2_26533 ( P3_R1077_U200 , P3_U3069 , P3_R1077_U199 );
nand NAND2_26534 ( P3_R1077_U201 , P3_U3410 , P3_R1077_U198 );
nand NAND2_26535 ( P3_R1077_U202 , P3_R1077_U5 , P3_R1077_U41 );
not NOT1_26536 ( P3_R1077_U203 , P3_R1077_U144 );
or OR2_26537 ( P3_R1077_U204 , P3_U3413 , P3_U3083 );
nand NAND2_26538 ( P3_R1077_U205 , P3_R1077_U204 , P3_R1077_U144 );
not NOT1_26539 ( P3_R1077_U206 , P3_R1077_U40 );
or OR2_26540 ( P3_R1077_U207 , P3_U3082 , P3_U3416 );
or OR2_26541 ( P3_R1077_U208 , P3_U3407 , P3_U3070 );
nand NAND2_26542 ( P3_R1077_U209 , P3_R1077_U208 , P3_R1077_U41 );
nand NAND2_26543 ( P3_R1077_U210 , P3_R1077_U119 , P3_R1077_U209 );
nand NAND2_26544 ( P3_R1077_U211 , P3_R1077_U195 , P3_R1077_U22 );
nand NAND2_26545 ( P3_R1077_U212 , P3_U3410 , P3_U3069 );
nand NAND2_26546 ( P3_R1077_U213 , P3_R1077_U120 , P3_R1077_U211 );
or OR2_26547 ( P3_R1077_U214 , P3_U3070 , P3_U3407 );
nand NAND2_26548 ( P3_R1077_U215 , P3_R1077_U185 , P3_R1077_U181 );
nand NAND2_26549 ( P3_R1077_U216 , P3_U3067 , P3_U3395 );
not NOT1_26550 ( P3_R1077_U217 , P3_R1077_U45 );
nand NAND2_26551 ( P3_R1077_U218 , P3_R1077_U121 , P3_R1077_U184 );
nand NAND2_26552 ( P3_R1077_U219 , P3_R1077_U45 , P3_R1077_U180 );
nand NAND2_26553 ( P3_R1077_U220 , P3_U3063 , P3_U3398 );
not NOT1_26554 ( P3_R1077_U221 , P3_R1077_U44 );
or OR2_26555 ( P3_R1077_U222 , P3_U3401 , P3_U3059 );
nand NAND2_26556 ( P3_R1077_U223 , P3_R1077_U222 , P3_R1077_U44 );
nand NAND2_26557 ( P3_R1077_U224 , P3_R1077_U123 , P3_R1077_U223 );
nand NAND2_26558 ( P3_R1077_U225 , P3_R1077_U221 , P3_R1077_U34 );
nand NAND2_26559 ( P3_R1077_U226 , P3_U3404 , P3_U3066 );
nand NAND2_26560 ( P3_R1077_U227 , P3_R1077_U124 , P3_R1077_U225 );
or OR2_26561 ( P3_R1077_U228 , P3_U3059 , P3_U3401 );
nand NAND2_26562 ( P3_R1077_U229 , P3_R1077_U184 , P3_R1077_U181 );
not NOT1_26563 ( P3_R1077_U230 , P3_R1077_U145 );
nand NAND2_26564 ( P3_R1077_U231 , P3_U3063 , P3_U3398 );
nand NAND4_26565 ( P3_R1077_U232 , P3_R1077_U401 , P3_R1077_U400 , P3_R1077_U43 , P3_R1077_U42 );
nand NAND2_26566 ( P3_R1077_U233 , P3_R1077_U43 , P3_R1077_U42 );
nand NAND2_26567 ( P3_R1077_U234 , P3_U3067 , P3_U3395 );
nand NAND2_26568 ( P3_R1077_U235 , P3_R1077_U125 , P3_R1077_U233 );
or OR2_26569 ( P3_R1077_U236 , P3_U3082 , P3_U3416 );
or OR2_26570 ( P3_R1077_U237 , P3_U3061 , P3_U3419 );
nand NAND2_26571 ( P3_R1077_U238 , P3_R1077_U177 , P3_R1077_U6 );
nand NAND2_26572 ( P3_R1077_U239 , P3_U3061 , P3_U3419 );
nand NAND2_26573 ( P3_R1077_U240 , P3_R1077_U127 , P3_R1077_U238 );
or OR2_26574 ( P3_R1077_U241 , P3_U3419 , P3_U3061 );
nand NAND2_26575 ( P3_R1077_U242 , P3_R1077_U126 , P3_R1077_U144 );
nand NAND2_26576 ( P3_R1077_U243 , P3_R1077_U241 , P3_R1077_U240 );
not NOT1_26577 ( P3_R1077_U244 , P3_R1077_U167 );
or OR2_26578 ( P3_R1077_U245 , P3_U3079 , P3_U3428 );
or OR2_26579 ( P3_R1077_U246 , P3_U3071 , P3_U3425 );
nand NAND2_26580 ( P3_R1077_U247 , P3_R1077_U174 , P3_R1077_U7 );
nand NAND2_26581 ( P3_R1077_U248 , P3_U3079 , P3_U3428 );
nand NAND2_26582 ( P3_R1077_U249 , P3_R1077_U129 , P3_R1077_U247 );
or OR2_26583 ( P3_R1077_U250 , P3_U3422 , P3_U3062 );
or OR2_26584 ( P3_R1077_U251 , P3_U3428 , P3_U3079 );
nand NAND2_26585 ( P3_R1077_U252 , P3_R1077_U128 , P3_R1077_U167 );
nand NAND2_26586 ( P3_R1077_U253 , P3_R1077_U251 , P3_R1077_U249 );
not NOT1_26587 ( P3_R1077_U254 , P3_R1077_U166 );
or OR2_26588 ( P3_R1077_U255 , P3_U3431 , P3_U3078 );
nand NAND2_26589 ( P3_R1077_U256 , P3_R1077_U255 , P3_R1077_U166 );
nand NAND2_26590 ( P3_R1077_U257 , P3_U3078 , P3_U3431 );
not NOT1_26591 ( P3_R1077_U258 , P3_R1077_U164 );
or OR2_26592 ( P3_R1077_U259 , P3_U3434 , P3_U3073 );
nand NAND2_26593 ( P3_R1077_U260 , P3_R1077_U259 , P3_R1077_U164 );
nand NAND2_26594 ( P3_R1077_U261 , P3_U3073 , P3_U3434 );
not NOT1_26595 ( P3_R1077_U262 , P3_R1077_U92 );
or OR2_26596 ( P3_R1077_U263 , P3_U3068 , P3_U3440 );
or OR2_26597 ( P3_R1077_U264 , P3_U3072 , P3_U3437 );
not NOT1_26598 ( P3_R1077_U265 , P3_R1077_U59 );
nand NAND2_26599 ( P3_R1077_U266 , P3_R1077_U60 , P3_R1077_U59 );
nand NAND2_26600 ( P3_R1077_U267 , P3_U3068 , P3_R1077_U266 );
nand NAND2_26601 ( P3_R1077_U268 , P3_U3440 , P3_R1077_U265 );
nand NAND2_26602 ( P3_R1077_U269 , P3_R1077_U8 , P3_R1077_U92 );
not NOT1_26603 ( P3_R1077_U270 , P3_R1077_U162 );
or OR2_26604 ( P3_R1077_U271 , P3_U3075 , P3_U3907 );
or OR2_26605 ( P3_R1077_U272 , P3_U3080 , P3_U3445 );
or OR2_26606 ( P3_R1077_U273 , P3_U3074 , P3_U3906 );
not NOT1_26607 ( P3_R1077_U274 , P3_R1077_U80 );
nand NAND2_26608 ( P3_R1077_U275 , P3_U3907 , P3_R1077_U274 );
nand NAND2_26609 ( P3_R1077_U276 , P3_R1077_U275 , P3_R1077_U90 );
nand NAND2_26610 ( P3_R1077_U277 , P3_R1077_U80 , P3_R1077_U81 );
nand NAND2_26611 ( P3_R1077_U278 , P3_R1077_U277 , P3_R1077_U276 );
nand NAND2_26612 ( P3_R1077_U279 , P3_R1077_U175 , P3_R1077_U9 );
nand NAND2_26613 ( P3_R1077_U280 , P3_U3074 , P3_U3906 );
nand NAND2_26614 ( P3_R1077_U281 , P3_R1077_U278 , P3_R1077_U279 );
or OR2_26615 ( P3_R1077_U282 , P3_U3443 , P3_U3081 );
or OR2_26616 ( P3_R1077_U283 , P3_U3906 , P3_U3074 );
nand NAND2_26617 ( P3_R1077_U284 , P3_R1077_U162 , P3_R1077_U131 );
nand NAND2_26618 ( P3_R1077_U285 , P3_R1077_U283 , P3_R1077_U281 );
not NOT1_26619 ( P3_R1077_U286 , P3_R1077_U159 );
or OR2_26620 ( P3_R1077_U287 , P3_U3905 , P3_U3060 );
nand NAND2_26621 ( P3_R1077_U288 , P3_R1077_U287 , P3_R1077_U159 );
nand NAND2_26622 ( P3_R1077_U289 , P3_U3060 , P3_U3905 );
not NOT1_26623 ( P3_R1077_U290 , P3_R1077_U157 );
or OR2_26624 ( P3_R1077_U291 , P3_U3904 , P3_U3065 );
nand NAND2_26625 ( P3_R1077_U292 , P3_R1077_U291 , P3_R1077_U157 );
nand NAND2_26626 ( P3_R1077_U293 , P3_U3065 , P3_U3904 );
not NOT1_26627 ( P3_R1077_U294 , P3_R1077_U155 );
or OR2_26628 ( P3_R1077_U295 , P3_U3057 , P3_U3902 );
nand NAND2_26629 ( P3_R1077_U296 , P3_R1077_U176 , P3_R1077_U173 );
not NOT1_26630 ( P3_R1077_U297 , P3_R1077_U86 );
or OR2_26631 ( P3_R1077_U298 , P3_U3903 , P3_U3064 );
nand NAND3_26632 ( P3_R1077_U299 , P3_R1077_U155 , P3_R1077_U298 , P3_R1077_U168 );
not NOT1_26633 ( P3_R1077_U300 , P3_R1077_U153 );
or OR2_26634 ( P3_R1077_U301 , P3_U3900 , P3_U3052 );
nand NAND2_26635 ( P3_R1077_U302 , P3_U3052 , P3_U3900 );
not NOT1_26636 ( P3_R1077_U303 , P3_R1077_U151 );
nand NAND2_26637 ( P3_R1077_U304 , P3_U3899 , P3_R1077_U151 );
not NOT1_26638 ( P3_R1077_U305 , P3_R1077_U149 );
nand NAND2_26639 ( P3_R1077_U306 , P3_R1077_U298 , P3_R1077_U155 );
not NOT1_26640 ( P3_R1077_U307 , P3_R1077_U89 );
or OR2_26641 ( P3_R1077_U308 , P3_U3902 , P3_U3057 );
nand NAND2_26642 ( P3_R1077_U309 , P3_R1077_U308 , P3_R1077_U89 );
nand NAND3_26643 ( P3_R1077_U310 , P3_R1077_U309 , P3_R1077_U173 , P3_R1077_U154 );
nand NAND2_26644 ( P3_R1077_U311 , P3_R1077_U307 , P3_R1077_U173 );
nand NAND2_26645 ( P3_R1077_U312 , P3_U3901 , P3_U3056 );
nand NAND3_26646 ( P3_R1077_U313 , P3_R1077_U311 , P3_R1077_U312 , P3_R1077_U168 );
or OR2_26647 ( P3_R1077_U314 , P3_U3057 , P3_U3902 );
nand NAND2_26648 ( P3_R1077_U315 , P3_R1077_U282 , P3_R1077_U162 );
not NOT1_26649 ( P3_R1077_U316 , P3_R1077_U91 );
nand NAND2_26650 ( P3_R1077_U317 , P3_R1077_U9 , P3_R1077_U91 );
nand NAND2_26651 ( P3_R1077_U318 , P3_R1077_U135 , P3_R1077_U317 );
nand NAND2_26652 ( P3_R1077_U319 , P3_R1077_U317 , P3_R1077_U278 );
nand NAND2_26653 ( P3_R1077_U320 , P3_R1077_U453 , P3_R1077_U319 );
or OR2_26654 ( P3_R1077_U321 , P3_U3445 , P3_U3080 );
nand NAND2_26655 ( P3_R1077_U322 , P3_R1077_U321 , P3_R1077_U91 );
nand NAND2_26656 ( P3_R1077_U323 , P3_R1077_U136 , P3_R1077_U322 );
nand NAND2_26657 ( P3_R1077_U324 , P3_R1077_U316 , P3_R1077_U80 );
nand NAND2_26658 ( P3_R1077_U325 , P3_U3075 , P3_U3907 );
nand NAND2_26659 ( P3_R1077_U326 , P3_R1077_U137 , P3_R1077_U324 );
or OR2_26660 ( P3_R1077_U327 , P3_U3392 , P3_U3077 );
not NOT1_26661 ( P3_R1077_U328 , P3_R1077_U161 );
or OR2_26662 ( P3_R1077_U329 , P3_U3080 , P3_U3445 );
or OR2_26663 ( P3_R1077_U330 , P3_U3437 , P3_U3072 );
nand NAND2_26664 ( P3_R1077_U331 , P3_R1077_U330 , P3_R1077_U92 );
nand NAND2_26665 ( P3_R1077_U332 , P3_R1077_U138 , P3_R1077_U331 );
nand NAND2_26666 ( P3_R1077_U333 , P3_R1077_U262 , P3_R1077_U59 );
nand NAND2_26667 ( P3_R1077_U334 , P3_U3440 , P3_U3068 );
nand NAND2_26668 ( P3_R1077_U335 , P3_R1077_U139 , P3_R1077_U333 );
or OR2_26669 ( P3_R1077_U336 , P3_U3072 , P3_U3437 );
nand NAND2_26670 ( P3_R1077_U337 , P3_R1077_U250 , P3_R1077_U167 );
not NOT1_26671 ( P3_R1077_U338 , P3_R1077_U93 );
or OR2_26672 ( P3_R1077_U339 , P3_U3425 , P3_U3071 );
nand NAND2_26673 ( P3_R1077_U340 , P3_R1077_U339 , P3_R1077_U93 );
nand NAND2_26674 ( P3_R1077_U341 , P3_R1077_U140 , P3_R1077_U340 );
nand NAND2_26675 ( P3_R1077_U342 , P3_R1077_U338 , P3_R1077_U172 );
nand NAND2_26676 ( P3_R1077_U343 , P3_U3079 , P3_U3428 );
nand NAND2_26677 ( P3_R1077_U344 , P3_R1077_U141 , P3_R1077_U342 );
or OR2_26678 ( P3_R1077_U345 , P3_U3071 , P3_U3425 );
or OR2_26679 ( P3_R1077_U346 , P3_U3416 , P3_U3082 );
nand NAND2_26680 ( P3_R1077_U347 , P3_R1077_U346 , P3_R1077_U40 );
nand NAND2_26681 ( P3_R1077_U348 , P3_R1077_U142 , P3_R1077_U347 );
nand NAND2_26682 ( P3_R1077_U349 , P3_R1077_U206 , P3_R1077_U171 );
nand NAND2_26683 ( P3_R1077_U350 , P3_U3061 , P3_U3419 );
nand NAND2_26684 ( P3_R1077_U351 , P3_R1077_U143 , P3_R1077_U349 );
nand NAND2_26685 ( P3_R1077_U352 , P3_R1077_U207 , P3_R1077_U171 );
nand NAND2_26686 ( P3_R1077_U353 , P3_R1077_U204 , P3_R1077_U61 );
nand NAND2_26687 ( P3_R1077_U354 , P3_R1077_U214 , P3_R1077_U22 );
nand NAND2_26688 ( P3_R1077_U355 , P3_R1077_U228 , P3_R1077_U34 );
nand NAND2_26689 ( P3_R1077_U356 , P3_R1077_U231 , P3_R1077_U180 );
nand NAND2_26690 ( P3_R1077_U357 , P3_R1077_U314 , P3_R1077_U173 );
nand NAND2_26691 ( P3_R1077_U358 , P3_R1077_U298 , P3_R1077_U176 );
nand NAND2_26692 ( P3_R1077_U359 , P3_R1077_U329 , P3_R1077_U80 );
nand NAND2_26693 ( P3_R1077_U360 , P3_R1077_U282 , P3_R1077_U77 );
nand NAND2_26694 ( P3_R1077_U361 , P3_R1077_U336 , P3_R1077_U59 );
nand NAND2_26695 ( P3_R1077_U362 , P3_R1077_U345 , P3_R1077_U172 );
nand NAND2_26696 ( P3_R1077_U363 , P3_R1077_U250 , P3_R1077_U68 );
nand NAND2_26697 ( P3_R1077_U364 , P3_U3899 , P3_U3053 );
nand NAND2_26698 ( P3_R1077_U365 , P3_R1077_U296 , P3_R1077_U168 );
nand NAND2_26699 ( P3_R1077_U366 , P3_U3056 , P3_R1077_U295 );
nand NAND2_26700 ( P3_R1077_U367 , P3_U3901 , P3_R1077_U295 );
nand NAND3_26701 ( P3_R1077_U368 , P3_R1077_U296 , P3_R1077_U168 , P3_R1077_U301 );
nand NAND3_26702 ( P3_R1077_U369 , P3_R1077_U155 , P3_R1077_U168 , P3_R1077_U133 );
nand NAND2_26703 ( P3_R1077_U370 , P3_R1077_U297 , P3_R1077_U301 );
nand NAND2_26704 ( P3_R1077_U371 , P3_U3082 , P3_R1077_U39 );
nand NAND2_26705 ( P3_R1077_U372 , P3_U3416 , P3_R1077_U38 );
nand NAND2_26706 ( P3_R1077_U373 , P3_R1077_U372 , P3_R1077_U371 );
nand NAND2_26707 ( P3_R1077_U374 , P3_R1077_U352 , P3_R1077_U40 );
nand NAND2_26708 ( P3_R1077_U375 , P3_R1077_U373 , P3_R1077_U206 );
nand NAND2_26709 ( P3_R1077_U376 , P3_U3083 , P3_R1077_U36 );
nand NAND2_26710 ( P3_R1077_U377 , P3_U3413 , P3_R1077_U37 );
nand NAND2_26711 ( P3_R1077_U378 , P3_R1077_U377 , P3_R1077_U376 );
nand NAND2_26712 ( P3_R1077_U379 , P3_R1077_U353 , P3_R1077_U144 );
nand NAND2_26713 ( P3_R1077_U380 , P3_R1077_U203 , P3_R1077_U378 );
nand NAND2_26714 ( P3_R1077_U381 , P3_U3069 , P3_R1077_U23 );
nand NAND2_26715 ( P3_R1077_U382 , P3_U3410 , P3_R1077_U21 );
nand NAND2_26716 ( P3_R1077_U383 , P3_U3070 , P3_R1077_U19 );
nand NAND2_26717 ( P3_R1077_U384 , P3_U3407 , P3_R1077_U20 );
nand NAND2_26718 ( P3_R1077_U385 , P3_R1077_U384 , P3_R1077_U383 );
nand NAND2_26719 ( P3_R1077_U386 , P3_R1077_U354 , P3_R1077_U41 );
nand NAND2_26720 ( P3_R1077_U387 , P3_R1077_U385 , P3_R1077_U195 );
nand NAND2_26721 ( P3_R1077_U388 , P3_U3066 , P3_R1077_U35 );
nand NAND2_26722 ( P3_R1077_U389 , P3_U3404 , P3_R1077_U26 );
nand NAND2_26723 ( P3_R1077_U390 , P3_U3059 , P3_R1077_U24 );
nand NAND2_26724 ( P3_R1077_U391 , P3_U3401 , P3_R1077_U25 );
nand NAND2_26725 ( P3_R1077_U392 , P3_R1077_U391 , P3_R1077_U390 );
nand NAND2_26726 ( P3_R1077_U393 , P3_R1077_U355 , P3_R1077_U44 );
nand NAND2_26727 ( P3_R1077_U394 , P3_R1077_U392 , P3_R1077_U221 );
nand NAND2_26728 ( P3_R1077_U395 , P3_U3063 , P3_R1077_U32 );
nand NAND2_26729 ( P3_R1077_U396 , P3_U3398 , P3_R1077_U33 );
nand NAND2_26730 ( P3_R1077_U397 , P3_R1077_U396 , P3_R1077_U395 );
nand NAND2_26731 ( P3_R1077_U398 , P3_R1077_U356 , P3_R1077_U145 );
nand NAND2_26732 ( P3_R1077_U399 , P3_R1077_U230 , P3_R1077_U397 );
nand NAND2_26733 ( P3_R1077_U400 , P3_U3067 , P3_R1077_U27 );
nand NAND2_26734 ( P3_R1077_U401 , P3_U3395 , P3_R1077_U28 );
nand NAND2_26735 ( P3_R1077_U402 , P3_U3054 , P3_R1077_U147 );
nand NAND2_26736 ( P3_R1077_U403 , P3_U3908 , P3_R1077_U146 );
nand NAND2_26737 ( P3_R1077_U404 , P3_U3054 , P3_R1077_U147 );
nand NAND2_26738 ( P3_R1077_U405 , P3_U3908 , P3_R1077_U146 );
nand NAND2_26739 ( P3_R1077_U406 , P3_R1077_U405 , P3_R1077_U404 );
nand NAND2_26740 ( P3_R1077_U407 , P3_R1077_U148 , P3_R1077_U149 );
nand NAND2_26741 ( P3_R1077_U408 , P3_R1077_U305 , P3_R1077_U406 );
nand NAND2_26742 ( P3_R1077_U409 , P3_U3053 , P3_R1077_U88 );
nand NAND2_26743 ( P3_R1077_U410 , P3_U3899 , P3_R1077_U87 );
nand NAND2_26744 ( P3_R1077_U411 , P3_U3053 , P3_R1077_U88 );
nand NAND2_26745 ( P3_R1077_U412 , P3_U3899 , P3_R1077_U87 );
nand NAND2_26746 ( P3_R1077_U413 , P3_R1077_U412 , P3_R1077_U411 );
nand NAND2_26747 ( P3_R1077_U414 , P3_R1077_U150 , P3_R1077_U151 );
nand NAND2_26748 ( P3_R1077_U415 , P3_R1077_U303 , P3_R1077_U413 );
nand NAND2_26749 ( P3_R1077_U416 , P3_U3052 , P3_R1077_U46 );
nand NAND2_26750 ( P3_R1077_U417 , P3_U3900 , P3_R1077_U47 );
nand NAND2_26751 ( P3_R1077_U418 , P3_U3052 , P3_R1077_U46 );
nand NAND2_26752 ( P3_R1077_U419 , P3_U3900 , P3_R1077_U47 );
nand NAND2_26753 ( P3_R1077_U420 , P3_R1077_U419 , P3_R1077_U418 );
nand NAND2_26754 ( P3_R1077_U421 , P3_R1077_U152 , P3_R1077_U153 );
nand NAND2_26755 ( P3_R1077_U422 , P3_R1077_U300 , P3_R1077_U420 );
nand NAND2_26756 ( P3_R1077_U423 , P3_U3056 , P3_R1077_U49 );
nand NAND2_26757 ( P3_R1077_U424 , P3_U3901 , P3_R1077_U48 );
nand NAND2_26758 ( P3_R1077_U425 , P3_U3057 , P3_R1077_U50 );
nand NAND2_26759 ( P3_R1077_U426 , P3_U3902 , P3_R1077_U51 );
nand NAND2_26760 ( P3_R1077_U427 , P3_R1077_U426 , P3_R1077_U425 );
nand NAND2_26761 ( P3_R1077_U428 , P3_R1077_U357 , P3_R1077_U89 );
nand NAND2_26762 ( P3_R1077_U429 , P3_R1077_U427 , P3_R1077_U307 );
nand NAND2_26763 ( P3_R1077_U430 , P3_U3064 , P3_R1077_U52 );
nand NAND2_26764 ( P3_R1077_U431 , P3_U3903 , P3_R1077_U53 );
nand NAND2_26765 ( P3_R1077_U432 , P3_R1077_U431 , P3_R1077_U430 );
nand NAND2_26766 ( P3_R1077_U433 , P3_R1077_U358 , P3_R1077_U155 );
nand NAND2_26767 ( P3_R1077_U434 , P3_R1077_U294 , P3_R1077_U432 );
nand NAND2_26768 ( P3_R1077_U435 , P3_U3065 , P3_R1077_U84 );
nand NAND2_26769 ( P3_R1077_U436 , P3_U3904 , P3_R1077_U85 );
nand NAND2_26770 ( P3_R1077_U437 , P3_U3065 , P3_R1077_U84 );
nand NAND2_26771 ( P3_R1077_U438 , P3_U3904 , P3_R1077_U85 );
nand NAND2_26772 ( P3_R1077_U439 , P3_R1077_U438 , P3_R1077_U437 );
nand NAND2_26773 ( P3_R1077_U440 , P3_R1077_U156 , P3_R1077_U157 );
nand NAND2_26774 ( P3_R1077_U441 , P3_R1077_U290 , P3_R1077_U439 );
nand NAND2_26775 ( P3_R1077_U442 , P3_U3060 , P3_R1077_U82 );
nand NAND2_26776 ( P3_R1077_U443 , P3_U3905 , P3_R1077_U83 );
nand NAND2_26777 ( P3_R1077_U444 , P3_U3060 , P3_R1077_U82 );
nand NAND2_26778 ( P3_R1077_U445 , P3_U3905 , P3_R1077_U83 );
nand NAND2_26779 ( P3_R1077_U446 , P3_R1077_U445 , P3_R1077_U444 );
nand NAND2_26780 ( P3_R1077_U447 , P3_R1077_U158 , P3_R1077_U159 );
nand NAND2_26781 ( P3_R1077_U448 , P3_R1077_U286 , P3_R1077_U446 );
nand NAND2_26782 ( P3_R1077_U449 , P3_U3074 , P3_R1077_U54 );
nand NAND2_26783 ( P3_R1077_U450 , P3_U3906 , P3_R1077_U55 );
nand NAND2_26784 ( P3_R1077_U451 , P3_U3074 , P3_R1077_U54 );
nand NAND2_26785 ( P3_R1077_U452 , P3_U3906 , P3_R1077_U55 );
nand NAND2_26786 ( P3_R1077_U453 , P3_R1077_U452 , P3_R1077_U451 );
nand NAND2_26787 ( P3_R1077_U454 , P3_U3075 , P3_R1077_U81 );
nand NAND2_26788 ( P3_R1077_U455 , P3_U3907 , P3_R1077_U90 );
nand NAND2_26789 ( P3_R1077_U456 , P3_R1077_U182 , P3_R1077_U161 );
nand NAND2_26790 ( P3_R1077_U457 , P3_R1077_U328 , P3_R1077_U31 );
nand NAND2_26791 ( P3_R1077_U458 , P3_U3080 , P3_R1077_U78 );
nand NAND2_26792 ( P3_R1077_U459 , P3_U3445 , P3_R1077_U79 );
nand NAND2_26793 ( P3_R1077_U460 , P3_R1077_U459 , P3_R1077_U458 );
nand NAND2_26794 ( P3_R1077_U461 , P3_R1077_U359 , P3_R1077_U91 );
nand NAND2_26795 ( P3_R1077_U462 , P3_R1077_U460 , P3_R1077_U316 );
nand NAND2_26796 ( P3_R1077_U463 , P3_U3081 , P3_R1077_U75 );
nand NAND2_26797 ( P3_R1077_U464 , P3_U3443 , P3_R1077_U76 );
nand NAND2_26798 ( P3_R1077_U465 , P3_R1077_U464 , P3_R1077_U463 );
nand NAND2_26799 ( P3_R1077_U466 , P3_R1077_U360 , P3_R1077_U162 );
nand NAND2_26800 ( P3_R1077_U467 , P3_R1077_U270 , P3_R1077_U465 );
nand NAND2_26801 ( P3_R1077_U468 , P3_U3068 , P3_R1077_U60 );
nand NAND2_26802 ( P3_R1077_U469 , P3_U3440 , P3_R1077_U58 );
nand NAND2_26803 ( P3_R1077_U470 , P3_U3072 , P3_R1077_U56 );
nand NAND2_26804 ( P3_R1077_U471 , P3_U3437 , P3_R1077_U57 );
nand NAND2_26805 ( P3_R1077_U472 , P3_R1077_U471 , P3_R1077_U470 );
nand NAND2_26806 ( P3_R1077_U473 , P3_R1077_U361 , P3_R1077_U92 );
nand NAND2_26807 ( P3_R1077_U474 , P3_R1077_U472 , P3_R1077_U262 );
nand NAND2_26808 ( P3_R1077_U475 , P3_U3073 , P3_R1077_U73 );
nand NAND2_26809 ( P3_R1077_U476 , P3_U3434 , P3_R1077_U74 );
nand NAND2_26810 ( P3_R1077_U477 , P3_U3073 , P3_R1077_U73 );
nand NAND2_26811 ( P3_R1077_U478 , P3_U3434 , P3_R1077_U74 );
nand NAND2_26812 ( P3_R1077_U479 , P3_R1077_U478 , P3_R1077_U477 );
nand NAND2_26813 ( P3_R1077_U480 , P3_R1077_U163 , P3_R1077_U164 );
nand NAND2_26814 ( P3_R1077_U481 , P3_R1077_U258 , P3_R1077_U479 );
nand NAND2_26815 ( P3_R1077_U482 , P3_U3078 , P3_R1077_U71 );
nand NAND2_26816 ( P3_R1077_U483 , P3_U3431 , P3_R1077_U72 );
nand NAND2_26817 ( P3_R1077_U484 , P3_U3078 , P3_R1077_U71 );
nand NAND2_26818 ( P3_R1077_U485 , P3_U3431 , P3_R1077_U72 );
nand NAND2_26819 ( P3_R1077_U486 , P3_R1077_U485 , P3_R1077_U484 );
nand NAND2_26820 ( P3_R1077_U487 , P3_R1077_U165 , P3_R1077_U166 );
nand NAND2_26821 ( P3_R1077_U488 , P3_R1077_U254 , P3_R1077_U486 );
nand NAND2_26822 ( P3_R1077_U489 , P3_U3079 , P3_R1077_U69 );
nand NAND2_26823 ( P3_R1077_U490 , P3_U3428 , P3_R1077_U70 );
nand NAND2_26824 ( P3_R1077_U491 , P3_U3071 , P3_R1077_U64 );
nand NAND2_26825 ( P3_R1077_U492 , P3_U3425 , P3_R1077_U65 );
nand NAND2_26826 ( P3_R1077_U493 , P3_R1077_U492 , P3_R1077_U491 );
nand NAND2_26827 ( P3_R1077_U494 , P3_R1077_U362 , P3_R1077_U93 );
nand NAND2_26828 ( P3_R1077_U495 , P3_R1077_U493 , P3_R1077_U338 );
nand NAND2_26829 ( P3_R1077_U496 , P3_U3062 , P3_R1077_U66 );
nand NAND2_26830 ( P3_R1077_U497 , P3_U3422 , P3_R1077_U67 );
nand NAND2_26831 ( P3_R1077_U498 , P3_R1077_U497 , P3_R1077_U496 );
nand NAND2_26832 ( P3_R1077_U499 , P3_R1077_U363 , P3_R1077_U167 );
nand NAND2_26833 ( P3_R1077_U500 , P3_R1077_U244 , P3_R1077_U498 );
nand NAND2_26834 ( P3_R1077_U501 , P3_U3061 , P3_R1077_U62 );
nand NAND2_26835 ( P3_R1077_U502 , P3_U3419 , P3_R1077_U63 );
nand NAND2_26836 ( P3_R1077_U503 , P3_U3076 , P3_R1077_U29 );
nand NAND2_26837 ( P3_R1077_U504 , P3_U3387 , P3_R1077_U30 );
and AND2_26838 ( P3_R1143_U4 , P3_R1143_U179 , P3_R1143_U178 );
and AND2_26839 ( P3_R1143_U5 , P3_R1143_U197 , P3_R1143_U196 );
and AND2_26840 ( P3_R1143_U6 , P3_R1143_U237 , P3_R1143_U236 );
and AND2_26841 ( P3_R1143_U7 , P3_R1143_U246 , P3_R1143_U245 );
and AND2_26842 ( P3_R1143_U8 , P3_R1143_U264 , P3_R1143_U263 );
and AND2_26843 ( P3_R1143_U9 , P3_R1143_U272 , P3_R1143_U271 );
and AND2_26844 ( P3_R1143_U10 , P3_R1143_U351 , P3_R1143_U348 );
and AND2_26845 ( P3_R1143_U11 , P3_R1143_U344 , P3_R1143_U341 );
and AND2_26846 ( P3_R1143_U12 , P3_R1143_U335 , P3_R1143_U332 );
and AND2_26847 ( P3_R1143_U13 , P3_R1143_U326 , P3_R1143_U323 );
and AND2_26848 ( P3_R1143_U14 , P3_R1143_U320 , P3_R1143_U318 );
and AND2_26849 ( P3_R1143_U15 , P3_R1143_U313 , P3_R1143_U310 );
and AND2_26850 ( P3_R1143_U16 , P3_R1143_U235 , P3_R1143_U232 );
and AND2_26851 ( P3_R1143_U17 , P3_R1143_U227 , P3_R1143_U224 );
and AND2_26852 ( P3_R1143_U18 , P3_R1143_U213 , P3_R1143_U210 );
not NOT1_26853 ( P3_R1143_U19 , P3_U3407 );
not NOT1_26854 ( P3_R1143_U20 , P3_U3070 );
not NOT1_26855 ( P3_R1143_U21 , P3_U3069 );
nand NAND2_26856 ( P3_R1143_U22 , P3_U3070 , P3_U3407 );
not NOT1_26857 ( P3_R1143_U23 , P3_U3410 );
not NOT1_26858 ( P3_R1143_U24 , P3_U3401 );
not NOT1_26859 ( P3_R1143_U25 , P3_U3059 );
not NOT1_26860 ( P3_R1143_U26 , P3_U3066 );
not NOT1_26861 ( P3_R1143_U27 , P3_U3395 );
not NOT1_26862 ( P3_R1143_U28 , P3_U3067 );
not NOT1_26863 ( P3_R1143_U29 , P3_U3387 );
not NOT1_26864 ( P3_R1143_U30 , P3_U3076 );
nand NAND2_26865 ( P3_R1143_U31 , P3_U3076 , P3_U3387 );
not NOT1_26866 ( P3_R1143_U32 , P3_U3398 );
not NOT1_26867 ( P3_R1143_U33 , P3_U3063 );
nand NAND2_26868 ( P3_R1143_U34 , P3_U3059 , P3_U3401 );
not NOT1_26869 ( P3_R1143_U35 , P3_U3404 );
not NOT1_26870 ( P3_R1143_U36 , P3_U3413 );
not NOT1_26871 ( P3_R1143_U37 , P3_U3083 );
not NOT1_26872 ( P3_R1143_U38 , P3_U3082 );
not NOT1_26873 ( P3_R1143_U39 , P3_U3416 );
nand NAND2_26874 ( P3_R1143_U40 , P3_R1143_U63 , P3_R1143_U205 );
nand NAND2_26875 ( P3_R1143_U41 , P3_R1143_U117 , P3_R1143_U193 );
nand NAND2_26876 ( P3_R1143_U42 , P3_R1143_U182 , P3_R1143_U183 );
nand NAND2_26877 ( P3_R1143_U43 , P3_U3392 , P3_U3077 );
nand NAND2_26878 ( P3_R1143_U44 , P3_R1143_U122 , P3_R1143_U219 );
nand NAND2_26879 ( P3_R1143_U45 , P3_R1143_U216 , P3_R1143_U215 );
not NOT1_26880 ( P3_R1143_U46 , P3_U3900 );
not NOT1_26881 ( P3_R1143_U47 , P3_U3052 );
not NOT1_26882 ( P3_R1143_U48 , P3_U3056 );
not NOT1_26883 ( P3_R1143_U49 , P3_U3901 );
not NOT1_26884 ( P3_R1143_U50 , P3_U3902 );
not NOT1_26885 ( P3_R1143_U51 , P3_U3057 );
not NOT1_26886 ( P3_R1143_U52 , P3_U3903 );
not NOT1_26887 ( P3_R1143_U53 , P3_U3064 );
not NOT1_26888 ( P3_R1143_U54 , P3_U3906 );
not NOT1_26889 ( P3_R1143_U55 , P3_U3074 );
not NOT1_26890 ( P3_R1143_U56 , P3_U3437 );
not NOT1_26891 ( P3_R1143_U57 , P3_U3072 );
not NOT1_26892 ( P3_R1143_U58 , P3_U3068 );
nand NAND2_26893 ( P3_R1143_U59 , P3_U3072 , P3_U3437 );
not NOT1_26894 ( P3_R1143_U60 , P3_U3440 );
not NOT1_26895 ( P3_R1143_U61 , P3_U3419 );
not NOT1_26896 ( P3_R1143_U62 , P3_U3061 );
nand NAND2_26897 ( P3_R1143_U63 , P3_U3083 , P3_U3413 );
not NOT1_26898 ( P3_R1143_U64 , P3_U3425 );
not NOT1_26899 ( P3_R1143_U65 , P3_U3071 );
not NOT1_26900 ( P3_R1143_U66 , P3_U3422 );
not NOT1_26901 ( P3_R1143_U67 , P3_U3062 );
nand NAND2_26902 ( P3_R1143_U68 , P3_U3062 , P3_U3422 );
not NOT1_26903 ( P3_R1143_U69 , P3_U3428 );
not NOT1_26904 ( P3_R1143_U70 , P3_U3079 );
not NOT1_26905 ( P3_R1143_U71 , P3_U3431 );
not NOT1_26906 ( P3_R1143_U72 , P3_U3078 );
not NOT1_26907 ( P3_R1143_U73 , P3_U3434 );
not NOT1_26908 ( P3_R1143_U74 , P3_U3073 );
not NOT1_26909 ( P3_R1143_U75 , P3_U3443 );
not NOT1_26910 ( P3_R1143_U76 , P3_U3081 );
nand NAND2_26911 ( P3_R1143_U77 , P3_U3081 , P3_U3443 );
not NOT1_26912 ( P3_R1143_U78 , P3_U3445 );
not NOT1_26913 ( P3_R1143_U79 , P3_U3080 );
nand NAND2_26914 ( P3_R1143_U80 , P3_U3080 , P3_U3445 );
not NOT1_26915 ( P3_R1143_U81 , P3_U3907 );
not NOT1_26916 ( P3_R1143_U82 , P3_U3905 );
not NOT1_26917 ( P3_R1143_U83 , P3_U3060 );
not NOT1_26918 ( P3_R1143_U84 , P3_U3904 );
not NOT1_26919 ( P3_R1143_U85 , P3_U3065 );
nand NAND2_26920 ( P3_R1143_U86 , P3_U3901 , P3_U3056 );
not NOT1_26921 ( P3_R1143_U87 , P3_U3053 );
not NOT1_26922 ( P3_R1143_U88 , P3_U3899 );
nand NAND2_26923 ( P3_R1143_U89 , P3_R1143_U306 , P3_R1143_U176 );
not NOT1_26924 ( P3_R1143_U90 , P3_U3075 );
nand NAND2_26925 ( P3_R1143_U91 , P3_R1143_U77 , P3_R1143_U315 );
nand NAND2_26926 ( P3_R1143_U92 , P3_R1143_U261 , P3_R1143_U260 );
nand NAND2_26927 ( P3_R1143_U93 , P3_R1143_U68 , P3_R1143_U337 );
nand NAND2_26928 ( P3_R1143_U94 , P3_R1143_U457 , P3_R1143_U456 );
nand NAND2_26929 ( P3_R1143_U95 , P3_R1143_U504 , P3_R1143_U503 );
nand NAND2_26930 ( P3_R1143_U96 , P3_R1143_U375 , P3_R1143_U374 );
nand NAND2_26931 ( P3_R1143_U97 , P3_R1143_U380 , P3_R1143_U379 );
nand NAND2_26932 ( P3_R1143_U98 , P3_R1143_U387 , P3_R1143_U386 );
nand NAND2_26933 ( P3_R1143_U99 , P3_R1143_U394 , P3_R1143_U393 );
nand NAND2_26934 ( P3_R1143_U100 , P3_R1143_U399 , P3_R1143_U398 );
nand NAND2_26935 ( P3_R1143_U101 , P3_R1143_U408 , P3_R1143_U407 );
nand NAND2_26936 ( P3_R1143_U102 , P3_R1143_U415 , P3_R1143_U414 );
nand NAND2_26937 ( P3_R1143_U103 , P3_R1143_U422 , P3_R1143_U421 );
nand NAND2_26938 ( P3_R1143_U104 , P3_R1143_U429 , P3_R1143_U428 );
nand NAND2_26939 ( P3_R1143_U105 , P3_R1143_U434 , P3_R1143_U433 );
nand NAND2_26940 ( P3_R1143_U106 , P3_R1143_U441 , P3_R1143_U440 );
nand NAND2_26941 ( P3_R1143_U107 , P3_R1143_U448 , P3_R1143_U447 );
nand NAND2_26942 ( P3_R1143_U108 , P3_R1143_U462 , P3_R1143_U461 );
nand NAND2_26943 ( P3_R1143_U109 , P3_R1143_U467 , P3_R1143_U466 );
nand NAND2_26944 ( P3_R1143_U110 , P3_R1143_U474 , P3_R1143_U473 );
nand NAND2_26945 ( P3_R1143_U111 , P3_R1143_U481 , P3_R1143_U480 );
nand NAND2_26946 ( P3_R1143_U112 , P3_R1143_U488 , P3_R1143_U487 );
nand NAND2_26947 ( P3_R1143_U113 , P3_R1143_U495 , P3_R1143_U494 );
nand NAND2_26948 ( P3_R1143_U114 , P3_R1143_U500 , P3_R1143_U499 );
and AND2_26949 ( P3_R1143_U115 , P3_R1143_U189 , P3_R1143_U187 );
and AND2_26950 ( P3_R1143_U116 , P3_R1143_U4 , P3_R1143_U180 );
and AND2_26951 ( P3_R1143_U117 , P3_R1143_U194 , P3_R1143_U192 );
and AND2_26952 ( P3_R1143_U118 , P3_R1143_U201 , P3_R1143_U200 );
and AND3_26953 ( P3_R1143_U119 , P3_R1143_U382 , P3_R1143_U381 , P3_R1143_U22 );
and AND2_26954 ( P3_R1143_U120 , P3_R1143_U212 , P3_R1143_U5 );
and AND2_26955 ( P3_R1143_U121 , P3_R1143_U181 , P3_R1143_U180 );
and AND2_26956 ( P3_R1143_U122 , P3_R1143_U220 , P3_R1143_U218 );
and AND3_26957 ( P3_R1143_U123 , P3_R1143_U389 , P3_R1143_U388 , P3_R1143_U34 );
and AND2_26958 ( P3_R1143_U124 , P3_R1143_U226 , P3_R1143_U4 );
and AND2_26959 ( P3_R1143_U125 , P3_R1143_U234 , P3_R1143_U181 );
and AND2_26960 ( P3_R1143_U126 , P3_R1143_U204 , P3_R1143_U6 );
and AND2_26961 ( P3_R1143_U127 , P3_R1143_U243 , P3_R1143_U239 );
and AND2_26962 ( P3_R1143_U128 , P3_R1143_U250 , P3_R1143_U7 );
and AND2_26963 ( P3_R1143_U129 , P3_R1143_U248 , P3_R1143_U172 );
and AND2_26964 ( P3_R1143_U130 , P3_R1143_U268 , P3_R1143_U267 );
and AND3_26965 ( P3_R1143_U131 , P3_R1143_U9 , P3_R1143_U282 , P3_R1143_U273 );
and AND2_26966 ( P3_R1143_U132 , P3_R1143_U285 , P3_R1143_U280 );
and AND2_26967 ( P3_R1143_U133 , P3_R1143_U301 , P3_R1143_U298 );
and AND2_26968 ( P3_R1143_U134 , P3_R1143_U368 , P3_R1143_U302 );
and AND2_26969 ( P3_R1143_U135 , P3_R1143_U160 , P3_R1143_U278 );
and AND3_26970 ( P3_R1143_U136 , P3_R1143_U455 , P3_R1143_U454 , P3_R1143_U80 );
and AND2_26971 ( P3_R1143_U137 , P3_R1143_U325 , P3_R1143_U9 );
and AND3_26972 ( P3_R1143_U138 , P3_R1143_U469 , P3_R1143_U468 , P3_R1143_U59 );
and AND2_26973 ( P3_R1143_U139 , P3_R1143_U334 , P3_R1143_U8 );
and AND3_26974 ( P3_R1143_U140 , P3_R1143_U490 , P3_R1143_U489 , P3_R1143_U172 );
and AND2_26975 ( P3_R1143_U141 , P3_R1143_U343 , P3_R1143_U7 );
and AND3_26976 ( P3_R1143_U142 , P3_R1143_U502 , P3_R1143_U501 , P3_R1143_U171 );
and AND2_26977 ( P3_R1143_U143 , P3_R1143_U350 , P3_R1143_U6 );
nand NAND2_26978 ( P3_R1143_U144 , P3_R1143_U118 , P3_R1143_U202 );
nand NAND2_26979 ( P3_R1143_U145 , P3_R1143_U217 , P3_R1143_U229 );
not NOT1_26980 ( P3_R1143_U146 , P3_U3054 );
not NOT1_26981 ( P3_R1143_U147 , P3_U3908 );
and AND2_26982 ( P3_R1143_U148 , P3_R1143_U403 , P3_R1143_U402 );
nand NAND3_26983 ( P3_R1143_U149 , P3_R1143_U304 , P3_R1143_U169 , P3_R1143_U364 );
and AND2_26984 ( P3_R1143_U150 , P3_R1143_U410 , P3_R1143_U409 );
nand NAND3_26985 ( P3_R1143_U151 , P3_R1143_U370 , P3_R1143_U369 , P3_R1143_U134 );
and AND2_26986 ( P3_R1143_U152 , P3_R1143_U417 , P3_R1143_U416 );
nand NAND3_26987 ( P3_R1143_U153 , P3_R1143_U365 , P3_R1143_U299 , P3_R1143_U86 );
and AND2_26988 ( P3_R1143_U154 , P3_R1143_U424 , P3_R1143_U423 );
nand NAND2_26989 ( P3_R1143_U155 , P3_R1143_U293 , P3_R1143_U292 );
and AND2_26990 ( P3_R1143_U156 , P3_R1143_U436 , P3_R1143_U435 );
nand NAND2_26991 ( P3_R1143_U157 , P3_R1143_U289 , P3_R1143_U288 );
and AND2_26992 ( P3_R1143_U158 , P3_R1143_U443 , P3_R1143_U442 );
nand NAND2_26993 ( P3_R1143_U159 , P3_R1143_U132 , P3_R1143_U284 );
and AND2_26994 ( P3_R1143_U160 , P3_R1143_U450 , P3_R1143_U449 );
nand NAND2_26995 ( P3_R1143_U161 , P3_R1143_U43 , P3_R1143_U327 );
nand NAND2_26996 ( P3_R1143_U162 , P3_R1143_U130 , P3_R1143_U269 );
and AND2_26997 ( P3_R1143_U163 , P3_R1143_U476 , P3_R1143_U475 );
nand NAND2_26998 ( P3_R1143_U164 , P3_R1143_U257 , P3_R1143_U256 );
and AND2_26999 ( P3_R1143_U165 , P3_R1143_U483 , P3_R1143_U482 );
nand NAND2_27000 ( P3_R1143_U166 , P3_R1143_U253 , P3_R1143_U252 );
nand NAND2_27001 ( P3_R1143_U167 , P3_R1143_U127 , P3_R1143_U242 );
nand NAND2_27002 ( P3_R1143_U168 , P3_R1143_U367 , P3_R1143_U366 );
nand NAND2_27003 ( P3_R1143_U169 , P3_U3053 , P3_R1143_U151 );
not NOT1_27004 ( P3_R1143_U170 , P3_R1143_U34 );
nand NAND2_27005 ( P3_R1143_U171 , P3_U3416 , P3_U3082 );
nand NAND2_27006 ( P3_R1143_U172 , P3_U3071 , P3_U3425 );
nand NAND2_27007 ( P3_R1143_U173 , P3_U3057 , P3_U3902 );
not NOT1_27008 ( P3_R1143_U174 , P3_R1143_U68 );
not NOT1_27009 ( P3_R1143_U175 , P3_R1143_U77 );
nand NAND2_27010 ( P3_R1143_U176 , P3_U3064 , P3_U3903 );
not NOT1_27011 ( P3_R1143_U177 , P3_R1143_U63 );
or OR2_27012 ( P3_R1143_U178 , P3_U3066 , P3_U3404 );
or OR2_27013 ( P3_R1143_U179 , P3_U3059 , P3_U3401 );
or OR2_27014 ( P3_R1143_U180 , P3_U3398 , P3_U3063 );
or OR2_27015 ( P3_R1143_U181 , P3_U3395 , P3_U3067 );
not NOT1_27016 ( P3_R1143_U182 , P3_R1143_U31 );
or OR2_27017 ( P3_R1143_U183 , P3_U3392 , P3_U3077 );
not NOT1_27018 ( P3_R1143_U184 , P3_R1143_U42 );
not NOT1_27019 ( P3_R1143_U185 , P3_R1143_U43 );
nand NAND2_27020 ( P3_R1143_U186 , P3_R1143_U42 , P3_R1143_U43 );
nand NAND2_27021 ( P3_R1143_U187 , P3_U3067 , P3_U3395 );
nand NAND2_27022 ( P3_R1143_U188 , P3_R1143_U186 , P3_R1143_U181 );
nand NAND2_27023 ( P3_R1143_U189 , P3_U3063 , P3_U3398 );
nand NAND2_27024 ( P3_R1143_U190 , P3_R1143_U115 , P3_R1143_U188 );
nand NAND2_27025 ( P3_R1143_U191 , P3_R1143_U35 , P3_R1143_U34 );
nand NAND2_27026 ( P3_R1143_U192 , P3_U3066 , P3_R1143_U191 );
nand NAND2_27027 ( P3_R1143_U193 , P3_R1143_U116 , P3_R1143_U190 );
nand NAND2_27028 ( P3_R1143_U194 , P3_U3404 , P3_R1143_U170 );
not NOT1_27029 ( P3_R1143_U195 , P3_R1143_U41 );
or OR2_27030 ( P3_R1143_U196 , P3_U3069 , P3_U3410 );
or OR2_27031 ( P3_R1143_U197 , P3_U3070 , P3_U3407 );
not NOT1_27032 ( P3_R1143_U198 , P3_R1143_U22 );
nand NAND2_27033 ( P3_R1143_U199 , P3_R1143_U23 , P3_R1143_U22 );
nand NAND2_27034 ( P3_R1143_U200 , P3_U3069 , P3_R1143_U199 );
nand NAND2_27035 ( P3_R1143_U201 , P3_U3410 , P3_R1143_U198 );
nand NAND2_27036 ( P3_R1143_U202 , P3_R1143_U5 , P3_R1143_U41 );
not NOT1_27037 ( P3_R1143_U203 , P3_R1143_U144 );
or OR2_27038 ( P3_R1143_U204 , P3_U3413 , P3_U3083 );
nand NAND2_27039 ( P3_R1143_U205 , P3_R1143_U204 , P3_R1143_U144 );
not NOT1_27040 ( P3_R1143_U206 , P3_R1143_U40 );
or OR2_27041 ( P3_R1143_U207 , P3_U3082 , P3_U3416 );
or OR2_27042 ( P3_R1143_U208 , P3_U3407 , P3_U3070 );
nand NAND2_27043 ( P3_R1143_U209 , P3_R1143_U208 , P3_R1143_U41 );
nand NAND2_27044 ( P3_R1143_U210 , P3_R1143_U119 , P3_R1143_U209 );
nand NAND2_27045 ( P3_R1143_U211 , P3_R1143_U195 , P3_R1143_U22 );
nand NAND2_27046 ( P3_R1143_U212 , P3_U3410 , P3_U3069 );
nand NAND2_27047 ( P3_R1143_U213 , P3_R1143_U120 , P3_R1143_U211 );
or OR2_27048 ( P3_R1143_U214 , P3_U3070 , P3_U3407 );
nand NAND2_27049 ( P3_R1143_U215 , P3_R1143_U185 , P3_R1143_U181 );
nand NAND2_27050 ( P3_R1143_U216 , P3_U3067 , P3_U3395 );
not NOT1_27051 ( P3_R1143_U217 , P3_R1143_U45 );
nand NAND2_27052 ( P3_R1143_U218 , P3_R1143_U121 , P3_R1143_U184 );
nand NAND2_27053 ( P3_R1143_U219 , P3_R1143_U45 , P3_R1143_U180 );
nand NAND2_27054 ( P3_R1143_U220 , P3_U3063 , P3_U3398 );
not NOT1_27055 ( P3_R1143_U221 , P3_R1143_U44 );
or OR2_27056 ( P3_R1143_U222 , P3_U3401 , P3_U3059 );
nand NAND2_27057 ( P3_R1143_U223 , P3_R1143_U222 , P3_R1143_U44 );
nand NAND2_27058 ( P3_R1143_U224 , P3_R1143_U123 , P3_R1143_U223 );
nand NAND2_27059 ( P3_R1143_U225 , P3_R1143_U221 , P3_R1143_U34 );
nand NAND2_27060 ( P3_R1143_U226 , P3_U3404 , P3_U3066 );
nand NAND2_27061 ( P3_R1143_U227 , P3_R1143_U124 , P3_R1143_U225 );
or OR2_27062 ( P3_R1143_U228 , P3_U3059 , P3_U3401 );
nand NAND2_27063 ( P3_R1143_U229 , P3_R1143_U184 , P3_R1143_U181 );
not NOT1_27064 ( P3_R1143_U230 , P3_R1143_U145 );
nand NAND2_27065 ( P3_R1143_U231 , P3_U3063 , P3_U3398 );
nand NAND4_27066 ( P3_R1143_U232 , P3_R1143_U401 , P3_R1143_U400 , P3_R1143_U43 , P3_R1143_U42 );
nand NAND2_27067 ( P3_R1143_U233 , P3_R1143_U43 , P3_R1143_U42 );
nand NAND2_27068 ( P3_R1143_U234 , P3_U3067 , P3_U3395 );
nand NAND2_27069 ( P3_R1143_U235 , P3_R1143_U125 , P3_R1143_U233 );
or OR2_27070 ( P3_R1143_U236 , P3_U3082 , P3_U3416 );
or OR2_27071 ( P3_R1143_U237 , P3_U3061 , P3_U3419 );
nand NAND2_27072 ( P3_R1143_U238 , P3_R1143_U177 , P3_R1143_U6 );
nand NAND2_27073 ( P3_R1143_U239 , P3_U3061 , P3_U3419 );
nand NAND2_27074 ( P3_R1143_U240 , P3_R1143_U171 , P3_R1143_U238 );
or OR2_27075 ( P3_R1143_U241 , P3_U3419 , P3_U3061 );
nand NAND2_27076 ( P3_R1143_U242 , P3_R1143_U126 , P3_R1143_U144 );
nand NAND2_27077 ( P3_R1143_U243 , P3_R1143_U241 , P3_R1143_U240 );
not NOT1_27078 ( P3_R1143_U244 , P3_R1143_U167 );
or OR2_27079 ( P3_R1143_U245 , P3_U3079 , P3_U3428 );
or OR2_27080 ( P3_R1143_U246 , P3_U3071 , P3_U3425 );
nand NAND2_27081 ( P3_R1143_U247 , P3_R1143_U174 , P3_R1143_U7 );
nand NAND2_27082 ( P3_R1143_U248 , P3_U3079 , P3_U3428 );
nand NAND2_27083 ( P3_R1143_U249 , P3_R1143_U129 , P3_R1143_U247 );
or OR2_27084 ( P3_R1143_U250 , P3_U3422 , P3_U3062 );
or OR2_27085 ( P3_R1143_U251 , P3_U3428 , P3_U3079 );
nand NAND2_27086 ( P3_R1143_U252 , P3_R1143_U128 , P3_R1143_U167 );
nand NAND2_27087 ( P3_R1143_U253 , P3_R1143_U251 , P3_R1143_U249 );
not NOT1_27088 ( P3_R1143_U254 , P3_R1143_U166 );
or OR2_27089 ( P3_R1143_U255 , P3_U3431 , P3_U3078 );
nand NAND2_27090 ( P3_R1143_U256 , P3_R1143_U255 , P3_R1143_U166 );
nand NAND2_27091 ( P3_R1143_U257 , P3_U3078 , P3_U3431 );
not NOT1_27092 ( P3_R1143_U258 , P3_R1143_U164 );
or OR2_27093 ( P3_R1143_U259 , P3_U3434 , P3_U3073 );
nand NAND2_27094 ( P3_R1143_U260 , P3_R1143_U259 , P3_R1143_U164 );
nand NAND2_27095 ( P3_R1143_U261 , P3_U3073 , P3_U3434 );
not NOT1_27096 ( P3_R1143_U262 , P3_R1143_U92 );
or OR2_27097 ( P3_R1143_U263 , P3_U3068 , P3_U3440 );
or OR2_27098 ( P3_R1143_U264 , P3_U3072 , P3_U3437 );
not NOT1_27099 ( P3_R1143_U265 , P3_R1143_U59 );
nand NAND2_27100 ( P3_R1143_U266 , P3_R1143_U60 , P3_R1143_U59 );
nand NAND2_27101 ( P3_R1143_U267 , P3_U3068 , P3_R1143_U266 );
nand NAND2_27102 ( P3_R1143_U268 , P3_U3440 , P3_R1143_U265 );
nand NAND2_27103 ( P3_R1143_U269 , P3_R1143_U8 , P3_R1143_U92 );
not NOT1_27104 ( P3_R1143_U270 , P3_R1143_U162 );
or OR2_27105 ( P3_R1143_U271 , P3_U3075 , P3_U3907 );
or OR2_27106 ( P3_R1143_U272 , P3_U3080 , P3_U3445 );
or OR2_27107 ( P3_R1143_U273 , P3_U3074 , P3_U3906 );
not NOT1_27108 ( P3_R1143_U274 , P3_R1143_U80 );
nand NAND2_27109 ( P3_R1143_U275 , P3_U3907 , P3_R1143_U274 );
nand NAND2_27110 ( P3_R1143_U276 , P3_R1143_U275 , P3_R1143_U90 );
nand NAND2_27111 ( P3_R1143_U277 , P3_R1143_U80 , P3_R1143_U81 );
nand NAND2_27112 ( P3_R1143_U278 , P3_R1143_U277 , P3_R1143_U276 );
nand NAND2_27113 ( P3_R1143_U279 , P3_R1143_U175 , P3_R1143_U9 );
nand NAND2_27114 ( P3_R1143_U280 , P3_U3074 , P3_U3906 );
nand NAND2_27115 ( P3_R1143_U281 , P3_R1143_U278 , P3_R1143_U279 );
or OR2_27116 ( P3_R1143_U282 , P3_U3443 , P3_U3081 );
or OR2_27117 ( P3_R1143_U283 , P3_U3906 , P3_U3074 );
nand NAND2_27118 ( P3_R1143_U284 , P3_R1143_U162 , P3_R1143_U131 );
nand NAND2_27119 ( P3_R1143_U285 , P3_R1143_U283 , P3_R1143_U281 );
not NOT1_27120 ( P3_R1143_U286 , P3_R1143_U159 );
or OR2_27121 ( P3_R1143_U287 , P3_U3905 , P3_U3060 );
nand NAND2_27122 ( P3_R1143_U288 , P3_R1143_U287 , P3_R1143_U159 );
nand NAND2_27123 ( P3_R1143_U289 , P3_U3060 , P3_U3905 );
not NOT1_27124 ( P3_R1143_U290 , P3_R1143_U157 );
or OR2_27125 ( P3_R1143_U291 , P3_U3904 , P3_U3065 );
nand NAND2_27126 ( P3_R1143_U292 , P3_R1143_U291 , P3_R1143_U157 );
nand NAND2_27127 ( P3_R1143_U293 , P3_U3065 , P3_U3904 );
not NOT1_27128 ( P3_R1143_U294 , P3_R1143_U155 );
or OR2_27129 ( P3_R1143_U295 , P3_U3057 , P3_U3902 );
nand NAND2_27130 ( P3_R1143_U296 , P3_R1143_U176 , P3_R1143_U173 );
not NOT1_27131 ( P3_R1143_U297 , P3_R1143_U86 );
or OR2_27132 ( P3_R1143_U298 , P3_U3903 , P3_U3064 );
nand NAND3_27133 ( P3_R1143_U299 , P3_R1143_U155 , P3_R1143_U298 , P3_R1143_U168 );
not NOT1_27134 ( P3_R1143_U300 , P3_R1143_U153 );
or OR2_27135 ( P3_R1143_U301 , P3_U3900 , P3_U3052 );
nand NAND2_27136 ( P3_R1143_U302 , P3_U3052 , P3_U3900 );
not NOT1_27137 ( P3_R1143_U303 , P3_R1143_U151 );
nand NAND2_27138 ( P3_R1143_U304 , P3_U3899 , P3_R1143_U151 );
not NOT1_27139 ( P3_R1143_U305 , P3_R1143_U149 );
nand NAND2_27140 ( P3_R1143_U306 , P3_R1143_U298 , P3_R1143_U155 );
not NOT1_27141 ( P3_R1143_U307 , P3_R1143_U89 );
or OR2_27142 ( P3_R1143_U308 , P3_U3902 , P3_U3057 );
nand NAND2_27143 ( P3_R1143_U309 , P3_R1143_U308 , P3_R1143_U89 );
nand NAND3_27144 ( P3_R1143_U310 , P3_R1143_U309 , P3_R1143_U173 , P3_R1143_U154 );
nand NAND2_27145 ( P3_R1143_U311 , P3_R1143_U307 , P3_R1143_U173 );
nand NAND2_27146 ( P3_R1143_U312 , P3_U3901 , P3_U3056 );
nand NAND3_27147 ( P3_R1143_U313 , P3_R1143_U311 , P3_R1143_U312 , P3_R1143_U168 );
or OR2_27148 ( P3_R1143_U314 , P3_U3057 , P3_U3902 );
nand NAND2_27149 ( P3_R1143_U315 , P3_R1143_U282 , P3_R1143_U162 );
not NOT1_27150 ( P3_R1143_U316 , P3_R1143_U91 );
nand NAND2_27151 ( P3_R1143_U317 , P3_R1143_U9 , P3_R1143_U91 );
nand NAND2_27152 ( P3_R1143_U318 , P3_R1143_U135 , P3_R1143_U317 );
nand NAND2_27153 ( P3_R1143_U319 , P3_R1143_U317 , P3_R1143_U278 );
nand NAND2_27154 ( P3_R1143_U320 , P3_R1143_U453 , P3_R1143_U319 );
or OR2_27155 ( P3_R1143_U321 , P3_U3445 , P3_U3080 );
nand NAND2_27156 ( P3_R1143_U322 , P3_R1143_U321 , P3_R1143_U91 );
nand NAND2_27157 ( P3_R1143_U323 , P3_R1143_U136 , P3_R1143_U322 );
nand NAND2_27158 ( P3_R1143_U324 , P3_R1143_U316 , P3_R1143_U80 );
nand NAND2_27159 ( P3_R1143_U325 , P3_U3075 , P3_U3907 );
nand NAND2_27160 ( P3_R1143_U326 , P3_R1143_U137 , P3_R1143_U324 );
or OR2_27161 ( P3_R1143_U327 , P3_U3392 , P3_U3077 );
not NOT1_27162 ( P3_R1143_U328 , P3_R1143_U161 );
or OR2_27163 ( P3_R1143_U329 , P3_U3080 , P3_U3445 );
or OR2_27164 ( P3_R1143_U330 , P3_U3437 , P3_U3072 );
nand NAND2_27165 ( P3_R1143_U331 , P3_R1143_U330 , P3_R1143_U92 );
nand NAND2_27166 ( P3_R1143_U332 , P3_R1143_U138 , P3_R1143_U331 );
nand NAND2_27167 ( P3_R1143_U333 , P3_R1143_U262 , P3_R1143_U59 );
nand NAND2_27168 ( P3_R1143_U334 , P3_U3440 , P3_U3068 );
nand NAND2_27169 ( P3_R1143_U335 , P3_R1143_U139 , P3_R1143_U333 );
or OR2_27170 ( P3_R1143_U336 , P3_U3072 , P3_U3437 );
nand NAND2_27171 ( P3_R1143_U337 , P3_R1143_U250 , P3_R1143_U167 );
not NOT1_27172 ( P3_R1143_U338 , P3_R1143_U93 );
or OR2_27173 ( P3_R1143_U339 , P3_U3425 , P3_U3071 );
nand NAND2_27174 ( P3_R1143_U340 , P3_R1143_U339 , P3_R1143_U93 );
nand NAND2_27175 ( P3_R1143_U341 , P3_R1143_U140 , P3_R1143_U340 );
nand NAND2_27176 ( P3_R1143_U342 , P3_R1143_U338 , P3_R1143_U172 );
nand NAND2_27177 ( P3_R1143_U343 , P3_U3079 , P3_U3428 );
nand NAND2_27178 ( P3_R1143_U344 , P3_R1143_U141 , P3_R1143_U342 );
or OR2_27179 ( P3_R1143_U345 , P3_U3071 , P3_U3425 );
or OR2_27180 ( P3_R1143_U346 , P3_U3416 , P3_U3082 );
nand NAND2_27181 ( P3_R1143_U347 , P3_R1143_U346 , P3_R1143_U40 );
nand NAND2_27182 ( P3_R1143_U348 , P3_R1143_U142 , P3_R1143_U347 );
nand NAND2_27183 ( P3_R1143_U349 , P3_R1143_U206 , P3_R1143_U171 );
nand NAND2_27184 ( P3_R1143_U350 , P3_U3061 , P3_U3419 );
nand NAND2_27185 ( P3_R1143_U351 , P3_R1143_U143 , P3_R1143_U349 );
nand NAND2_27186 ( P3_R1143_U352 , P3_R1143_U207 , P3_R1143_U171 );
nand NAND2_27187 ( P3_R1143_U353 , P3_R1143_U204 , P3_R1143_U63 );
nand NAND2_27188 ( P3_R1143_U354 , P3_R1143_U214 , P3_R1143_U22 );
nand NAND2_27189 ( P3_R1143_U355 , P3_R1143_U228 , P3_R1143_U34 );
nand NAND2_27190 ( P3_R1143_U356 , P3_R1143_U231 , P3_R1143_U180 );
nand NAND2_27191 ( P3_R1143_U357 , P3_R1143_U314 , P3_R1143_U173 );
nand NAND2_27192 ( P3_R1143_U358 , P3_R1143_U298 , P3_R1143_U176 );
nand NAND2_27193 ( P3_R1143_U359 , P3_R1143_U329 , P3_R1143_U80 );
nand NAND2_27194 ( P3_R1143_U360 , P3_R1143_U282 , P3_R1143_U77 );
nand NAND2_27195 ( P3_R1143_U361 , P3_R1143_U336 , P3_R1143_U59 );
nand NAND2_27196 ( P3_R1143_U362 , P3_R1143_U345 , P3_R1143_U172 );
nand NAND2_27197 ( P3_R1143_U363 , P3_R1143_U250 , P3_R1143_U68 );
nand NAND2_27198 ( P3_R1143_U364 , P3_U3899 , P3_U3053 );
nand NAND2_27199 ( P3_R1143_U365 , P3_R1143_U296 , P3_R1143_U168 );
nand NAND2_27200 ( P3_R1143_U366 , P3_U3056 , P3_R1143_U295 );
nand NAND2_27201 ( P3_R1143_U367 , P3_U3901 , P3_R1143_U295 );
nand NAND3_27202 ( P3_R1143_U368 , P3_R1143_U296 , P3_R1143_U168 , P3_R1143_U301 );
nand NAND3_27203 ( P3_R1143_U369 , P3_R1143_U155 , P3_R1143_U168 , P3_R1143_U133 );
nand NAND2_27204 ( P3_R1143_U370 , P3_R1143_U297 , P3_R1143_U301 );
nand NAND2_27205 ( P3_R1143_U371 , P3_U3082 , P3_R1143_U39 );
nand NAND2_27206 ( P3_R1143_U372 , P3_U3416 , P3_R1143_U38 );
nand NAND2_27207 ( P3_R1143_U373 , P3_R1143_U372 , P3_R1143_U371 );
nand NAND2_27208 ( P3_R1143_U374 , P3_R1143_U352 , P3_R1143_U40 );
nand NAND2_27209 ( P3_R1143_U375 , P3_R1143_U373 , P3_R1143_U206 );
nand NAND2_27210 ( P3_R1143_U376 , P3_U3083 , P3_R1143_U36 );
nand NAND2_27211 ( P3_R1143_U377 , P3_U3413 , P3_R1143_U37 );
nand NAND2_27212 ( P3_R1143_U378 , P3_R1143_U377 , P3_R1143_U376 );
nand NAND2_27213 ( P3_R1143_U379 , P3_R1143_U353 , P3_R1143_U144 );
nand NAND2_27214 ( P3_R1143_U380 , P3_R1143_U203 , P3_R1143_U378 );
nand NAND2_27215 ( P3_R1143_U381 , P3_U3069 , P3_R1143_U23 );
nand NAND2_27216 ( P3_R1143_U382 , P3_U3410 , P3_R1143_U21 );
nand NAND2_27217 ( P3_R1143_U383 , P3_U3070 , P3_R1143_U19 );
nand NAND2_27218 ( P3_R1143_U384 , P3_U3407 , P3_R1143_U20 );
nand NAND2_27219 ( P3_R1143_U385 , P3_R1143_U384 , P3_R1143_U383 );
nand NAND2_27220 ( P3_R1143_U386 , P3_R1143_U354 , P3_R1143_U41 );
nand NAND2_27221 ( P3_R1143_U387 , P3_R1143_U385 , P3_R1143_U195 );
nand NAND2_27222 ( P3_R1143_U388 , P3_U3066 , P3_R1143_U35 );
nand NAND2_27223 ( P3_R1143_U389 , P3_U3404 , P3_R1143_U26 );
nand NAND2_27224 ( P3_R1143_U390 , P3_U3059 , P3_R1143_U24 );
nand NAND2_27225 ( P3_R1143_U391 , P3_U3401 , P3_R1143_U25 );
nand NAND2_27226 ( P3_R1143_U392 , P3_R1143_U391 , P3_R1143_U390 );
nand NAND2_27227 ( P3_R1143_U393 , P3_R1143_U355 , P3_R1143_U44 );
nand NAND2_27228 ( P3_R1143_U394 , P3_R1143_U392 , P3_R1143_U221 );
nand NAND2_27229 ( P3_R1143_U395 , P3_U3063 , P3_R1143_U32 );
nand NAND2_27230 ( P3_R1143_U396 , P3_U3398 , P3_R1143_U33 );
nand NAND2_27231 ( P3_R1143_U397 , P3_R1143_U396 , P3_R1143_U395 );
nand NAND2_27232 ( P3_R1143_U398 , P3_R1143_U356 , P3_R1143_U145 );
nand NAND2_27233 ( P3_R1143_U399 , P3_R1143_U230 , P3_R1143_U397 );
nand NAND2_27234 ( P3_R1143_U400 , P3_U3067 , P3_R1143_U27 );
nand NAND2_27235 ( P3_R1143_U401 , P3_U3395 , P3_R1143_U28 );
nand NAND2_27236 ( P3_R1143_U402 , P3_U3054 , P3_R1143_U147 );
nand NAND2_27237 ( P3_R1143_U403 , P3_U3908 , P3_R1143_U146 );
nand NAND2_27238 ( P3_R1143_U404 , P3_U3054 , P3_R1143_U147 );
nand NAND2_27239 ( P3_R1143_U405 , P3_U3908 , P3_R1143_U146 );
nand NAND2_27240 ( P3_R1143_U406 , P3_R1143_U405 , P3_R1143_U404 );
nand NAND2_27241 ( P3_R1143_U407 , P3_R1143_U148 , P3_R1143_U149 );
nand NAND2_27242 ( P3_R1143_U408 , P3_R1143_U305 , P3_R1143_U406 );
nand NAND2_27243 ( P3_R1143_U409 , P3_U3053 , P3_R1143_U88 );
nand NAND2_27244 ( P3_R1143_U410 , P3_U3899 , P3_R1143_U87 );
nand NAND2_27245 ( P3_R1143_U411 , P3_U3053 , P3_R1143_U88 );
nand NAND2_27246 ( P3_R1143_U412 , P3_U3899 , P3_R1143_U87 );
nand NAND2_27247 ( P3_R1143_U413 , P3_R1143_U412 , P3_R1143_U411 );
nand NAND2_27248 ( P3_R1143_U414 , P3_R1143_U150 , P3_R1143_U151 );
nand NAND2_27249 ( P3_R1143_U415 , P3_R1143_U303 , P3_R1143_U413 );
nand NAND2_27250 ( P3_R1143_U416 , P3_U3052 , P3_R1143_U46 );
nand NAND2_27251 ( P3_R1143_U417 , P3_U3900 , P3_R1143_U47 );
nand NAND2_27252 ( P3_R1143_U418 , P3_U3052 , P3_R1143_U46 );
nand NAND2_27253 ( P3_R1143_U419 , P3_U3900 , P3_R1143_U47 );
nand NAND2_27254 ( P3_R1143_U420 , P3_R1143_U419 , P3_R1143_U418 );
nand NAND2_27255 ( P3_R1143_U421 , P3_R1143_U152 , P3_R1143_U153 );
nand NAND2_27256 ( P3_R1143_U422 , P3_R1143_U300 , P3_R1143_U420 );
nand NAND2_27257 ( P3_R1143_U423 , P3_U3056 , P3_R1143_U49 );
nand NAND2_27258 ( P3_R1143_U424 , P3_U3901 , P3_R1143_U48 );
nand NAND2_27259 ( P3_R1143_U425 , P3_U3057 , P3_R1143_U50 );
nand NAND2_27260 ( P3_R1143_U426 , P3_U3902 , P3_R1143_U51 );
nand NAND2_27261 ( P3_R1143_U427 , P3_R1143_U426 , P3_R1143_U425 );
nand NAND2_27262 ( P3_R1143_U428 , P3_R1143_U357 , P3_R1143_U89 );
nand NAND2_27263 ( P3_R1143_U429 , P3_R1143_U427 , P3_R1143_U307 );
nand NAND2_27264 ( P3_R1143_U430 , P3_U3064 , P3_R1143_U52 );
nand NAND2_27265 ( P3_R1143_U431 , P3_U3903 , P3_R1143_U53 );
nand NAND2_27266 ( P3_R1143_U432 , P3_R1143_U431 , P3_R1143_U430 );
nand NAND2_27267 ( P3_R1143_U433 , P3_R1143_U358 , P3_R1143_U155 );
nand NAND2_27268 ( P3_R1143_U434 , P3_R1143_U294 , P3_R1143_U432 );
nand NAND2_27269 ( P3_R1143_U435 , P3_U3065 , P3_R1143_U84 );
nand NAND2_27270 ( P3_R1143_U436 , P3_U3904 , P3_R1143_U85 );
nand NAND2_27271 ( P3_R1143_U437 , P3_U3065 , P3_R1143_U84 );
nand NAND2_27272 ( P3_R1143_U438 , P3_U3904 , P3_R1143_U85 );
nand NAND2_27273 ( P3_R1143_U439 , P3_R1143_U438 , P3_R1143_U437 );
nand NAND2_27274 ( P3_R1143_U440 , P3_R1143_U156 , P3_R1143_U157 );
nand NAND2_27275 ( P3_R1143_U441 , P3_R1143_U290 , P3_R1143_U439 );
nand NAND2_27276 ( P3_R1143_U442 , P3_U3060 , P3_R1143_U82 );
nand NAND2_27277 ( P3_R1143_U443 , P3_U3905 , P3_R1143_U83 );
nand NAND2_27278 ( P3_R1143_U444 , P3_U3060 , P3_R1143_U82 );
nand NAND2_27279 ( P3_R1143_U445 , P3_U3905 , P3_R1143_U83 );
nand NAND2_27280 ( P3_R1143_U446 , P3_R1143_U445 , P3_R1143_U444 );
nand NAND2_27281 ( P3_R1143_U447 , P3_R1143_U158 , P3_R1143_U159 );
nand NAND2_27282 ( P3_R1143_U448 , P3_R1143_U286 , P3_R1143_U446 );
nand NAND2_27283 ( P3_R1143_U449 , P3_U3074 , P3_R1143_U54 );
nand NAND2_27284 ( P3_R1143_U450 , P3_U3906 , P3_R1143_U55 );
nand NAND2_27285 ( P3_R1143_U451 , P3_U3074 , P3_R1143_U54 );
nand NAND2_27286 ( P3_R1143_U452 , P3_U3906 , P3_R1143_U55 );
nand NAND2_27287 ( P3_R1143_U453 , P3_R1143_U452 , P3_R1143_U451 );
nand NAND2_27288 ( P3_R1143_U454 , P3_U3075 , P3_R1143_U81 );
nand NAND2_27289 ( P3_R1143_U455 , P3_U3907 , P3_R1143_U90 );
nand NAND2_27290 ( P3_R1143_U456 , P3_R1143_U182 , P3_R1143_U161 );
nand NAND2_27291 ( P3_R1143_U457 , P3_R1143_U328 , P3_R1143_U31 );
nand NAND2_27292 ( P3_R1143_U458 , P3_U3080 , P3_R1143_U78 );
nand NAND2_27293 ( P3_R1143_U459 , P3_U3445 , P3_R1143_U79 );
nand NAND2_27294 ( P3_R1143_U460 , P3_R1143_U459 , P3_R1143_U458 );
nand NAND2_27295 ( P3_R1143_U461 , P3_R1143_U359 , P3_R1143_U91 );
nand NAND2_27296 ( P3_R1143_U462 , P3_R1143_U460 , P3_R1143_U316 );
nand NAND2_27297 ( P3_R1143_U463 , P3_U3081 , P3_R1143_U75 );
nand NAND2_27298 ( P3_R1143_U464 , P3_U3443 , P3_R1143_U76 );
nand NAND2_27299 ( P3_R1143_U465 , P3_R1143_U464 , P3_R1143_U463 );
nand NAND2_27300 ( P3_R1143_U466 , P3_R1143_U360 , P3_R1143_U162 );
nand NAND2_27301 ( P3_R1143_U467 , P3_R1143_U270 , P3_R1143_U465 );
nand NAND2_27302 ( P3_R1143_U468 , P3_U3068 , P3_R1143_U60 );
nand NAND2_27303 ( P3_R1143_U469 , P3_U3440 , P3_R1143_U58 );
nand NAND2_27304 ( P3_R1143_U470 , P3_U3072 , P3_R1143_U56 );
nand NAND2_27305 ( P3_R1143_U471 , P3_U3437 , P3_R1143_U57 );
nand NAND2_27306 ( P3_R1143_U472 , P3_R1143_U471 , P3_R1143_U470 );
nand NAND2_27307 ( P3_R1143_U473 , P3_R1143_U361 , P3_R1143_U92 );
nand NAND2_27308 ( P3_R1143_U474 , P3_R1143_U472 , P3_R1143_U262 );
nand NAND2_27309 ( P3_R1143_U475 , P3_U3073 , P3_R1143_U73 );
nand NAND2_27310 ( P3_R1143_U476 , P3_U3434 , P3_R1143_U74 );
nand NAND2_27311 ( P3_R1143_U477 , P3_U3073 , P3_R1143_U73 );
nand NAND2_27312 ( P3_R1143_U478 , P3_U3434 , P3_R1143_U74 );
nand NAND2_27313 ( P3_R1143_U479 , P3_R1143_U478 , P3_R1143_U477 );
nand NAND2_27314 ( P3_R1143_U480 , P3_R1143_U163 , P3_R1143_U164 );
nand NAND2_27315 ( P3_R1143_U481 , P3_R1143_U258 , P3_R1143_U479 );
nand NAND2_27316 ( P3_R1143_U482 , P3_U3078 , P3_R1143_U71 );
nand NAND2_27317 ( P3_R1143_U483 , P3_U3431 , P3_R1143_U72 );
nand NAND2_27318 ( P3_R1143_U484 , P3_U3078 , P3_R1143_U71 );
nand NAND2_27319 ( P3_R1143_U485 , P3_U3431 , P3_R1143_U72 );
nand NAND2_27320 ( P3_R1143_U486 , P3_R1143_U485 , P3_R1143_U484 );
nand NAND2_27321 ( P3_R1143_U487 , P3_R1143_U165 , P3_R1143_U166 );
nand NAND2_27322 ( P3_R1143_U488 , P3_R1143_U254 , P3_R1143_U486 );
nand NAND2_27323 ( P3_R1143_U489 , P3_U3079 , P3_R1143_U69 );
nand NAND2_27324 ( P3_R1143_U490 , P3_U3428 , P3_R1143_U70 );
nand NAND2_27325 ( P3_R1143_U491 , P3_U3071 , P3_R1143_U64 );
nand NAND2_27326 ( P3_R1143_U492 , P3_U3425 , P3_R1143_U65 );
nand NAND2_27327 ( P3_R1143_U493 , P3_R1143_U492 , P3_R1143_U491 );
nand NAND2_27328 ( P3_R1143_U494 , P3_R1143_U362 , P3_R1143_U93 );
nand NAND2_27329 ( P3_R1143_U495 , P3_R1143_U493 , P3_R1143_U338 );
nand NAND2_27330 ( P3_R1143_U496 , P3_U3062 , P3_R1143_U66 );
nand NAND2_27331 ( P3_R1143_U497 , P3_U3422 , P3_R1143_U67 );
nand NAND2_27332 ( P3_R1143_U498 , P3_R1143_U497 , P3_R1143_U496 );
nand NAND2_27333 ( P3_R1143_U499 , P3_R1143_U363 , P3_R1143_U167 );
nand NAND2_27334 ( P3_R1143_U500 , P3_R1143_U244 , P3_R1143_U498 );
nand NAND2_27335 ( P3_R1143_U501 , P3_U3061 , P3_R1143_U61 );
nand NAND2_27336 ( P3_R1143_U502 , P3_U3419 , P3_R1143_U62 );
nand NAND2_27337 ( P3_R1143_U503 , P3_U3076 , P3_R1143_U29 );
nand NAND2_27338 ( P3_R1143_U504 , P3_U3387 , P3_R1143_U30 );
and AND2_27339 ( P3_R1158_U4 , P3_R1158_U227 , P3_R1158_U226 );
and AND2_27340 ( P3_R1158_U5 , P3_R1158_U238 , P3_R1158_U237 );
and AND2_27341 ( P3_R1158_U6 , P3_R1158_U263 , P3_R1158_U262 );
and AND2_27342 ( P3_R1158_U7 , P3_R1158_U277 , P3_R1158_U276 );
and AND2_27343 ( P3_R1158_U8 , P3_R1158_U289 , P3_R1158_U288 );
and AND2_27344 ( P3_R1158_U9 , P3_R1158_U6 , P3_R1158_U267 );
and AND2_27345 ( P3_R1158_U10 , P3_R1158_U5 , P3_R1158_U235 );
and AND2_27346 ( P3_R1158_U11 , P3_R1158_U9 , P3_R1158_U260 );
and AND2_27347 ( P3_R1158_U12 , P3_R1158_U535 , P3_R1158_U534 );
and AND2_27348 ( P3_R1158_U13 , P3_R1158_U345 , P3_R1158_U342 );
and AND2_27349 ( P3_R1158_U14 , P3_R1158_U336 , P3_R1158_U333 );
and AND2_27350 ( P3_R1158_U15 , P3_R1158_U329 , P3_R1158_U326 );
and AND3_27351 ( P3_R1158_U16 , P3_R1158_U537 , P3_R1158_U536 , P3_R1158_U142 );
and AND2_27352 ( P3_R1158_U17 , P3_R1158_U256 , P3_R1158_U253 );
and AND2_27353 ( P3_R1158_U18 , P3_R1158_U249 , P3_R1158_U246 );
nand NAND2_27354 ( P3_R1158_U19 , P3_U3056 , P3_R1158_U306 );
not NOT1_27355 ( P3_R1158_U20 , P3_U3152 );
not NOT1_27356 ( P3_R1158_U21 , P3_U3083 );
not NOT1_27357 ( P3_R1158_U22 , P3_U3070 );
nand NAND2_27358 ( P3_R1158_U23 , P3_U3070 , P3_R1158_U67 );
not NOT1_27359 ( P3_R1158_U24 , P3_U3069 );
not NOT1_27360 ( P3_R1158_U25 , P3_U3066 );
nand NAND2_27361 ( P3_R1158_U26 , P3_U3066 , P3_R1158_U69 );
not NOT1_27362 ( P3_R1158_U27 , P3_U3067 );
nand NAND2_27363 ( P3_R1158_U28 , P3_U3067 , P3_R1158_U70 );
not NOT1_27364 ( P3_R1158_U29 , P3_U3063 );
not NOT1_27365 ( P3_R1158_U30 , P3_U3077 );
not NOT1_27366 ( P3_R1158_U31 , P3_U3076 );
not NOT1_27367 ( P3_R1158_U32 , P3_U3059 );
not NOT1_27368 ( P3_R1158_U33 , P3_U3082 );
nand NAND3_27369 ( P3_R1158_U34 , P3_R1158_U359 , P3_R1158_U241 , P3_R1158_U362 );
nand NAND2_27370 ( P3_R1158_U35 , P3_R1158_U379 , P3_R1158_U26 );
nand NAND3_27371 ( P3_R1158_U36 , P3_R1158_U361 , P3_R1158_U224 , P3_R1158_U360 );
not NOT1_27372 ( P3_R1158_U37 , P3_U3052 );
not NOT1_27373 ( P3_R1158_U38 , P3_U3057 );
not NOT1_27374 ( P3_R1158_U39 , P3_U3064 );
not NOT1_27375 ( P3_R1158_U40 , P3_U3056 );
not NOT1_27376 ( P3_R1158_U41 , P3_U3072 );
nand NAND2_27377 ( P3_R1158_U42 , P3_U3072 , P3_R1158_U79 );
not NOT1_27378 ( P3_R1158_U43 , P3_U3068 );
not NOT1_27379 ( P3_R1158_U44 , P3_U3078 );
not NOT1_27380 ( P3_R1158_U45 , P3_U3071 );
not NOT1_27381 ( P3_R1158_U46 , P3_U3062 );
nand NAND2_27382 ( P3_R1158_U47 , P3_U3062 , P3_R1158_U84 );
not NOT1_27383 ( P3_R1158_U48 , P3_U3079 );
not NOT1_27384 ( P3_R1158_U49 , P3_U3061 );
nand NAND2_27385 ( P3_R1158_U50 , P3_U3061 , P3_R1158_U85 );
not NOT1_27386 ( P3_R1158_U51 , P3_U3073 );
not NOT1_27387 ( P3_R1158_U52 , P3_U3081 );
not NOT1_27388 ( P3_R1158_U53 , P3_U3075 );
not NOT1_27389 ( P3_R1158_U54 , P3_U3080 );
nand NAND2_27390 ( P3_R1158_U55 , P3_U3080 , P3_R1158_U88 );
not NOT1_27391 ( P3_R1158_U56 , P3_U3074 );
not NOT1_27392 ( P3_R1158_U57 , P3_U3060 );
not NOT1_27393 ( P3_R1158_U58 , P3_U3065 );
nand NAND2_27394 ( P3_R1158_U59 , P3_U3057 , P3_R1158_U76 );
nand NAND2_27395 ( P3_R1158_U60 , P3_U3064 , P3_R1158_U77 );
nand NAND2_27396 ( P3_R1158_U61 , P3_R1158_U55 , P3_R1158_U322 );
nand NAND2_27397 ( P3_R1158_U62 , P3_R1158_U274 , P3_R1158_U273 );
nand NAND2_27398 ( P3_R1158_U63 , P3_R1158_U365 , P3_R1158_U269 );
nand NAND2_27399 ( P3_R1158_U64 , P3_R1158_U47 , P3_R1158_U338 );
nand NAND2_27400 ( P3_R1158_U65 , P3_R1158_U394 , P3_R1158_U393 );
nand NAND2_27401 ( P3_R1158_U66 , P3_R1158_U426 , P3_R1158_U425 );
nand NAND2_27402 ( P3_R1158_U67 , P3_R1158_U423 , P3_R1158_U422 );
nand NAND2_27403 ( P3_R1158_U68 , P3_R1158_U420 , P3_R1158_U419 );
nand NAND2_27404 ( P3_R1158_U69 , P3_R1158_U417 , P3_R1158_U416 );
nand NAND2_27405 ( P3_R1158_U70 , P3_R1158_U414 , P3_R1158_U413 );
nand NAND2_27406 ( P3_R1158_U71 , P3_R1158_U411 , P3_R1158_U410 );
nand NAND2_27407 ( P3_R1158_U72 , P3_R1158_U405 , P3_R1158_U404 );
nand NAND2_27408 ( P3_R1158_U73 , P3_R1158_U408 , P3_R1158_U407 );
nand NAND2_27409 ( P3_R1158_U74 , P3_R1158_U402 , P3_R1158_U401 );
nand NAND2_27410 ( P3_R1158_U75 , P3_R1158_U466 , P3_R1158_U465 );
nand NAND2_27411 ( P3_R1158_U76 , P3_R1158_U514 , P3_R1158_U513 );
nand NAND2_27412 ( P3_R1158_U77 , P3_R1158_U517 , P3_R1158_U516 );
nand NAND2_27413 ( P3_R1158_U78 , P3_R1158_U511 , P3_R1158_U510 );
nand NAND2_27414 ( P3_R1158_U79 , P3_R1158_U490 , P3_R1158_U489 );
nand NAND2_27415 ( P3_R1158_U80 , P3_R1158_U487 , P3_R1158_U486 );
nand NAND2_27416 ( P3_R1158_U81 , P3_R1158_U481 , P3_R1158_U480 );
nand NAND2_27417 ( P3_R1158_U82 , P3_R1158_U478 , P3_R1158_U477 );
nand NAND2_27418 ( P3_R1158_U83 , P3_R1158_U475 , P3_R1158_U474 );
nand NAND2_27419 ( P3_R1158_U84 , P3_R1158_U472 , P3_R1158_U471 );
nand NAND2_27420 ( P3_R1158_U85 , P3_R1158_U469 , P3_R1158_U468 );
nand NAND2_27421 ( P3_R1158_U86 , P3_R1158_U484 , P3_R1158_U483 );
nand NAND2_27422 ( P3_R1158_U87 , P3_R1158_U493 , P3_R1158_U492 );
nand NAND2_27423 ( P3_R1158_U88 , P3_R1158_U502 , P3_R1158_U501 );
nand NAND2_27424 ( P3_R1158_U89 , P3_R1158_U496 , P3_R1158_U495 );
nand NAND2_27425 ( P3_R1158_U90 , P3_R1158_U499 , P3_R1158_U498 );
nand NAND2_27426 ( P3_R1158_U91 , P3_R1158_U505 , P3_R1158_U504 );
nand NAND2_27427 ( P3_R1158_U92 , P3_R1158_U508 , P3_R1158_U507 );
nand NAND2_27428 ( P3_R1158_U93 , P3_R1158_U523 , P3_R1158_U522 );
nand NAND2_27429 ( P3_R1158_U94 , P3_R1158_U632 , P3_R1158_U631 );
nand NAND2_27430 ( P3_R1158_U95 , P3_R1158_U429 , P3_R1158_U428 );
nand NAND2_27431 ( P3_R1158_U96 , P3_R1158_U436 , P3_R1158_U435 );
nand NAND2_27432 ( P3_R1158_U97 , P3_R1158_U443 , P3_R1158_U442 );
nand NAND2_27433 ( P3_R1158_U98 , P3_R1158_U450 , P3_R1158_U449 );
nand NAND2_27434 ( P3_R1158_U99 , P3_R1158_U457 , P3_R1158_U456 );
nand NAND2_27435 ( P3_R1158_U100 , P3_R1158_U464 , P3_R1158_U463 );
nand NAND2_27436 ( P3_R1158_U101 , P3_R1158_U526 , P3_R1158_U525 );
nand NAND2_27437 ( P3_R1158_U102 , P3_R1158_U533 , P3_R1158_U532 );
and AND2_27438 ( P3_R1158_U103 , P3_R1158_U320 , P3_R1158_U209 );
and AND2_27439 ( P3_R1158_U104 , P3_R1158_U141 , P3_R1158_U12 );
nand NAND2_27440 ( P3_R1158_U105 , P3_R1158_U542 , P3_R1158_U541 );
nand NAND2_27441 ( P3_R1158_U106 , P3_R1158_U547 , P3_R1158_U546 );
nand NAND2_27442 ( P3_R1158_U107 , P3_R1158_U554 , P3_R1158_U553 );
nand NAND2_27443 ( P3_R1158_U108 , P3_R1158_U561 , P3_R1158_U560 );
nand NAND2_27444 ( P3_R1158_U109 , P3_R1158_U568 , P3_R1158_U567 );
nand NAND2_27445 ( P3_R1158_U110 , P3_R1158_U575 , P3_R1158_U574 );
nand NAND2_27446 ( P3_R1158_U111 , P3_R1158_U580 , P3_R1158_U579 );
nand NAND2_27447 ( P3_R1158_U112 , P3_R1158_U587 , P3_R1158_U586 );
nand NAND2_27448 ( P3_R1158_U113 , P3_R1158_U594 , P3_R1158_U593 );
nand NAND2_27449 ( P3_R1158_U114 , P3_R1158_U601 , P3_R1158_U600 );
nand NAND2_27450 ( P3_R1158_U115 , P3_R1158_U608 , P3_R1158_U607 );
nand NAND2_27451 ( P3_R1158_U116 , P3_R1158_U615 , P3_R1158_U614 );
nand NAND2_27452 ( P3_R1158_U117 , P3_R1158_U620 , P3_R1158_U619 );
nand NAND2_27453 ( P3_R1158_U118 , P3_R1158_U627 , P3_R1158_U626 );
and AND2_27454 ( P3_R1158_U119 , P3_R1158_U73 , P3_U3152 );
and AND2_27455 ( P3_R1158_U120 , P3_R1158_U230 , P3_R1158_U229 );
and AND2_27456 ( P3_R1158_U121 , P3_R1158_U242 , P3_R1158_U10 );
and AND2_27457 ( P3_R1158_U122 , P3_R1158_U364 , P3_R1158_U243 );
and AND3_27458 ( P3_R1158_U123 , P3_R1158_U438 , P3_R1158_U437 , P3_R1158_U23 );
and AND2_27459 ( P3_R1158_U124 , P3_R1158_U248 , P3_R1158_U5 );
and AND3_27460 ( P3_R1158_U125 , P3_R1158_U459 , P3_R1158_U458 , P3_R1158_U28 );
and AND2_27461 ( P3_R1158_U126 , P3_R1158_U255 , P3_R1158_U4 );
and AND2_27462 ( P3_R1158_U127 , P3_R1158_U265 , P3_R1158_U213 );
and AND2_27463 ( P3_R1158_U128 , P3_R1158_U270 , P3_R1158_U11 );
and AND2_27464 ( P3_R1158_U129 , P3_R1158_U373 , P3_R1158_U271 );
and AND2_27465 ( P3_R1158_U130 , P3_R1158_U281 , P3_R1158_U280 );
and AND2_27466 ( P3_R1158_U131 , P3_R1158_U293 , P3_R1158_U8 );
and AND2_27467 ( P3_R1158_U132 , P3_R1158_U291 , P3_R1158_U214 );
and AND2_27468 ( P3_R1158_U133 , P3_R1158_U314 , P3_R1158_U376 );
and AND2_27469 ( P3_R1158_U134 , P3_R1158_U316 , P3_R1158_U307 );
and AND2_27470 ( P3_R1158_U135 , P3_R1158_U316 , P3_R1158_U369 );
and AND2_27471 ( P3_R1158_U136 , P3_R1158_U374 , P3_R1158_U315 );
nand NAND2_27472 ( P3_R1158_U137 , P3_R1158_U520 , P3_R1158_U519 );
and AND2_27473 ( P3_R1158_U138 , P3_R1158_U515 , P3_R1158_U38 );
and AND2_27474 ( P3_R1158_U139 , P3_R1158_U320 , P3_R1158_U215 );
and AND2_27475 ( P3_R1158_U140 , P3_R1158_U320 , P3_R1158_U218 );
and AND2_27476 ( P3_R1158_U141 , P3_R1158_U60 , P3_R1158_U59 );
and AND3_27477 ( P3_R1158_U142 , P3_R1158_U391 , P3_R1158_U319 , P3_R1158_U392 );
and AND3_27478 ( P3_R1158_U143 , P3_R1158_U563 , P3_R1158_U562 , P3_R1158_U214 );
and AND2_27479 ( P3_R1158_U144 , P3_R1158_U328 , P3_R1158_U8 );
and AND3_27480 ( P3_R1158_U145 , P3_R1158_U589 , P3_R1158_U588 , P3_R1158_U42 );
and AND2_27481 ( P3_R1158_U146 , P3_R1158_U335 , P3_R1158_U7 );
and AND3_27482 ( P3_R1158_U147 , P3_R1158_U610 , P3_R1158_U609 , P3_R1158_U213 );
and AND2_27483 ( P3_R1158_U148 , P3_R1158_U344 , P3_R1158_U6 );
nand NAND2_27484 ( P3_R1158_U149 , P3_R1158_U629 , P3_R1158_U628 );
not NOT1_27485 ( P3_R1158_U150 , P3_U3416 );
and AND2_27486 ( P3_R1158_U151 , P3_R1158_U397 , P3_R1158_U396 );
not NOT1_27487 ( P3_R1158_U152 , P3_U3401 );
not NOT1_27488 ( P3_R1158_U153 , P3_U3392 );
not NOT1_27489 ( P3_R1158_U154 , P3_U3387 );
not NOT1_27490 ( P3_R1158_U155 , P3_U3398 );
not NOT1_27491 ( P3_R1158_U156 , P3_U3395 );
not NOT1_27492 ( P3_R1158_U157 , P3_U3404 );
not NOT1_27493 ( P3_R1158_U158 , P3_U3410 );
not NOT1_27494 ( P3_R1158_U159 , P3_U3407 );
not NOT1_27495 ( P3_R1158_U160 , P3_U3413 );
nand NAND2_27496 ( P3_R1158_U161 , P3_R1158_U122 , P3_R1158_U383 );
and AND2_27497 ( P3_R1158_U162 , P3_R1158_U431 , P3_R1158_U430 );
nand NAND2_27498 ( P3_R1158_U163 , P3_R1158_U363 , P3_R1158_U381 );
and AND2_27499 ( P3_R1158_U164 , P3_R1158_U445 , P3_R1158_U444 );
nand NAND3_27500 ( P3_R1158_U165 , P3_R1158_U233 , P3_R1158_U211 , P3_R1158_U356 );
and AND2_27501 ( P3_R1158_U166 , P3_R1158_U452 , P3_R1158_U451 );
nand NAND2_27502 ( P3_R1158_U167 , P3_R1158_U120 , P3_R1158_U231 );
not NOT1_27503 ( P3_R1158_U168 , P3_U3900 );
not NOT1_27504 ( P3_R1158_U169 , P3_U3419 );
not NOT1_27505 ( P3_R1158_U170 , P3_U3422 );
not NOT1_27506 ( P3_R1158_U171 , P3_U3428 );
not NOT1_27507 ( P3_R1158_U172 , P3_U3425 );
not NOT1_27508 ( P3_R1158_U173 , P3_U3431 );
not NOT1_27509 ( P3_R1158_U174 , P3_U3434 );
not NOT1_27510 ( P3_R1158_U175 , P3_U3440 );
not NOT1_27511 ( P3_R1158_U176 , P3_U3437 );
not NOT1_27512 ( P3_R1158_U177 , P3_U3443 );
not NOT1_27513 ( P3_R1158_U178 , P3_U3906 );
not NOT1_27514 ( P3_R1158_U179 , P3_U3907 );
not NOT1_27515 ( P3_R1158_U180 , P3_U3445 );
not NOT1_27516 ( P3_R1158_U181 , P3_U3905 );
not NOT1_27517 ( P3_R1158_U182 , P3_U3904 );
not NOT1_27518 ( P3_R1158_U183 , P3_U3901 );
not NOT1_27519 ( P3_R1158_U184 , P3_U3902 );
not NOT1_27520 ( P3_R1158_U185 , P3_U3903 );
not NOT1_27521 ( P3_R1158_U186 , P3_U3053 );
not NOT1_27522 ( P3_R1158_U187 , P3_U3899 );
and AND2_27523 ( P3_R1158_U188 , P3_R1158_U528 , P3_R1158_U527 );
nand NAND2_27524 ( P3_R1158_U189 , P3_R1158_U311 , P3_R1158_U310 );
nand NAND2_27525 ( P3_R1158_U190 , P3_R1158_U309 , P3_R1158_U192 );
nand NAND2_27526 ( P3_R1158_U191 , P3_R1158_U60 , P3_R1158_U190 );
nand NAND2_27527 ( P3_R1158_U192 , P3_R1158_U304 , P3_R1158_U303 );
and AND2_27528 ( P3_R1158_U193 , P3_R1158_U549 , P3_R1158_U548 );
nand NAND2_27529 ( P3_R1158_U194 , P3_R1158_U300 , P3_R1158_U299 );
and AND2_27530 ( P3_R1158_U195 , P3_R1158_U556 , P3_R1158_U555 );
nand NAND2_27531 ( P3_R1158_U196 , P3_R1158_U296 , P3_R1158_U295 );
and AND2_27532 ( P3_R1158_U197 , P3_R1158_U570 , P3_R1158_U569 );
nand NAND2_27533 ( P3_R1158_U198 , P3_R1158_U221 , P3_R1158_U220 );
nand NAND2_27534 ( P3_R1158_U199 , P3_R1158_U286 , P3_R1158_U285 );
and AND2_27535 ( P3_R1158_U200 , P3_R1158_U582 , P3_R1158_U581 );
nand NAND2_27536 ( P3_R1158_U201 , P3_R1158_U130 , P3_R1158_U282 );
and AND2_27537 ( P3_R1158_U202 , P3_R1158_U596 , P3_R1158_U595 );
nand NAND2_27538 ( P3_R1158_U203 , P3_R1158_U129 , P3_R1158_U389 );
and AND2_27539 ( P3_R1158_U204 , P3_R1158_U603 , P3_R1158_U602 );
nand NAND2_27540 ( P3_R1158_U205 , P3_R1158_U372 , P3_R1158_U387 );
nand NAND2_27541 ( P3_R1158_U206 , P3_R1158_U385 , P3_R1158_U50 );
and AND2_27542 ( P3_R1158_U207 , P3_R1158_U622 , P3_R1158_U621 );
nand NAND3_27543 ( P3_R1158_U208 , P3_R1158_U258 , P3_R1158_U210 , P3_R1158_U357 );
nand NAND2_27544 ( P3_R1158_U209 , P3_R1158_U19 , P3_R1158_U367 );
nand NAND2_27545 ( P3_R1158_U210 , P3_R1158_U65 , P3_R1158_U161 );
nand NAND2_27546 ( P3_R1158_U211 , P3_R1158_U74 , P3_R1158_U167 );
not NOT1_27547 ( P3_R1158_U212 , P3_R1158_U28 );
nand NAND2_27548 ( P3_R1158_U213 , P3_U3071 , P3_R1158_U82 );
nand NAND2_27549 ( P3_R1158_U214 , P3_U3075 , P3_R1158_U90 );
not NOT1_27550 ( P3_R1158_U215 , P3_R1158_U59 );
not NOT1_27551 ( P3_R1158_U216 , P3_R1158_U47 );
not NOT1_27552 ( P3_R1158_U217 , P3_R1158_U55 );
not NOT1_27553 ( P3_R1158_U218 , P3_R1158_U60 );
nand NAND2_27554 ( P3_R1158_U219 , P3_R1158_U409 , P3_R1158_U20 );
nand NAND2_27555 ( P3_R1158_U220 , P3_U3076 , P3_R1158_U219 );
nand NAND2_27556 ( P3_R1158_U221 , P3_U3152 , P3_R1158_U73 );
not NOT1_27557 ( P3_R1158_U222 , P3_R1158_U198 );
nand NAND2_27558 ( P3_R1158_U223 , P3_R1158_U406 , P3_R1158_U30 );
nand NAND2_27559 ( P3_R1158_U224 , P3_U3077 , P3_R1158_U72 );
not NOT1_27560 ( P3_R1158_U225 , P3_R1158_U36 );
nand NAND2_27561 ( P3_R1158_U226 , P3_R1158_U412 , P3_R1158_U29 );
nand NAND2_27562 ( P3_R1158_U227 , P3_R1158_U415 , P3_R1158_U27 );
nand NAND2_27563 ( P3_R1158_U228 , P3_R1158_U29 , P3_R1158_U28 );
nand NAND2_27564 ( P3_R1158_U229 , P3_R1158_U71 , P3_R1158_U228 );
nand NAND2_27565 ( P3_R1158_U230 , P3_U3063 , P3_R1158_U212 );
nand NAND2_27566 ( P3_R1158_U231 , P3_R1158_U4 , P3_R1158_U36 );
not NOT1_27567 ( P3_R1158_U232 , P3_R1158_U167 );
nand NAND2_27568 ( P3_R1158_U233 , P3_U3059 , P3_R1158_U167 );
not NOT1_27569 ( P3_R1158_U234 , P3_R1158_U165 );
nand NAND2_27570 ( P3_R1158_U235 , P3_R1158_U418 , P3_R1158_U25 );
not NOT1_27571 ( P3_R1158_U236 , P3_R1158_U26 );
nand NAND2_27572 ( P3_R1158_U237 , P3_R1158_U421 , P3_R1158_U24 );
nand NAND2_27573 ( P3_R1158_U238 , P3_R1158_U424 , P3_R1158_U22 );
not NOT1_27574 ( P3_R1158_U239 , P3_R1158_U23 );
nand NAND2_27575 ( P3_R1158_U240 , P3_R1158_U24 , P3_R1158_U23 );
nand NAND2_27576 ( P3_R1158_U241 , P3_U3069 , P3_R1158_U239 );
nand NAND2_27577 ( P3_R1158_U242 , P3_R1158_U427 , P3_R1158_U21 );
nand NAND2_27578 ( P3_R1158_U243 , P3_U3083 , P3_R1158_U66 );
nand NAND2_27579 ( P3_R1158_U244 , P3_R1158_U424 , P3_R1158_U22 );
nand NAND2_27580 ( P3_R1158_U245 , P3_R1158_U244 , P3_R1158_U35 );
nand NAND2_27581 ( P3_R1158_U246 , P3_R1158_U123 , P3_R1158_U245 );
nand NAND2_27582 ( P3_R1158_U247 , P3_R1158_U380 , P3_R1158_U23 );
nand NAND2_27583 ( P3_R1158_U248 , P3_U3069 , P3_R1158_U68 );
nand NAND2_27584 ( P3_R1158_U249 , P3_R1158_U124 , P3_R1158_U247 );
nand NAND2_27585 ( P3_R1158_U250 , P3_R1158_U424 , P3_R1158_U22 );
nand NAND2_27586 ( P3_R1158_U251 , P3_R1158_U415 , P3_R1158_U27 );
nand NAND2_27587 ( P3_R1158_U252 , P3_R1158_U251 , P3_R1158_U36 );
nand NAND2_27588 ( P3_R1158_U253 , P3_R1158_U125 , P3_R1158_U252 );
nand NAND2_27589 ( P3_R1158_U254 , P3_R1158_U225 , P3_R1158_U28 );
nand NAND2_27590 ( P3_R1158_U255 , P3_U3063 , P3_R1158_U71 );
nand NAND2_27591 ( P3_R1158_U256 , P3_R1158_U126 , P3_R1158_U254 );
nand NAND2_27592 ( P3_R1158_U257 , P3_R1158_U415 , P3_R1158_U27 );
nand NAND2_27593 ( P3_R1158_U258 , P3_U3082 , P3_R1158_U161 );
not NOT1_27594 ( P3_R1158_U259 , P3_R1158_U208 );
nand NAND2_27595 ( P3_R1158_U260 , P3_R1158_U470 , P3_R1158_U49 );
not NOT1_27596 ( P3_R1158_U261 , P3_R1158_U50 );
nand NAND2_27597 ( P3_R1158_U262 , P3_R1158_U476 , P3_R1158_U48 );
nand NAND2_27598 ( P3_R1158_U263 , P3_R1158_U479 , P3_R1158_U45 );
nand NAND2_27599 ( P3_R1158_U264 , P3_R1158_U216 , P3_R1158_U6 );
nand NAND2_27600 ( P3_R1158_U265 , P3_U3079 , P3_R1158_U83 );
nand NAND2_27601 ( P3_R1158_U266 , P3_R1158_U127 , P3_R1158_U264 );
nand NAND2_27602 ( P3_R1158_U267 , P3_R1158_U473 , P3_R1158_U46 );
nand NAND2_27603 ( P3_R1158_U268 , P3_R1158_U476 , P3_R1158_U48 );
nand NAND2_27604 ( P3_R1158_U269 , P3_R1158_U268 , P3_R1158_U266 );
nand NAND2_27605 ( P3_R1158_U270 , P3_R1158_U482 , P3_R1158_U44 );
nand NAND2_27606 ( P3_R1158_U271 , P3_U3078 , P3_R1158_U81 );
nand NAND2_27607 ( P3_R1158_U272 , P3_R1158_U485 , P3_R1158_U51 );
nand NAND2_27608 ( P3_R1158_U273 , P3_R1158_U272 , P3_R1158_U203 );
nand NAND2_27609 ( P3_R1158_U274 , P3_U3073 , P3_R1158_U86 );
not NOT1_27610 ( P3_R1158_U275 , P3_R1158_U62 );
nand NAND2_27611 ( P3_R1158_U276 , P3_R1158_U488 , P3_R1158_U43 );
nand NAND2_27612 ( P3_R1158_U277 , P3_R1158_U491 , P3_R1158_U41 );
not NOT1_27613 ( P3_R1158_U278 , P3_R1158_U42 );
nand NAND2_27614 ( P3_R1158_U279 , P3_R1158_U43 , P3_R1158_U42 );
nand NAND2_27615 ( P3_R1158_U280 , P3_R1158_U80 , P3_R1158_U279 );
nand NAND2_27616 ( P3_R1158_U281 , P3_U3068 , P3_R1158_U278 );
nand NAND2_27617 ( P3_R1158_U282 , P3_R1158_U7 , P3_R1158_U62 );
not NOT1_27618 ( P3_R1158_U283 , P3_R1158_U201 );
nand NAND2_27619 ( P3_R1158_U284 , P3_R1158_U494 , P3_R1158_U52 );
nand NAND2_27620 ( P3_R1158_U285 , P3_R1158_U284 , P3_R1158_U201 );
nand NAND2_27621 ( P3_R1158_U286 , P3_U3081 , P3_R1158_U87 );
not NOT1_27622 ( P3_R1158_U287 , P3_R1158_U199 );
nand NAND2_27623 ( P3_R1158_U288 , P3_R1158_U497 , P3_R1158_U56 );
nand NAND2_27624 ( P3_R1158_U289 , P3_R1158_U500 , P3_R1158_U53 );
nand NAND2_27625 ( P3_R1158_U290 , P3_R1158_U217 , P3_R1158_U8 );
nand NAND2_27626 ( P3_R1158_U291 , P3_U3074 , P3_R1158_U89 );
nand NAND2_27627 ( P3_R1158_U292 , P3_R1158_U132 , P3_R1158_U290 );
nand NAND2_27628 ( P3_R1158_U293 , P3_R1158_U503 , P3_R1158_U54 );
nand NAND2_27629 ( P3_R1158_U294 , P3_R1158_U497 , P3_R1158_U56 );
nand NAND2_27630 ( P3_R1158_U295 , P3_R1158_U131 , P3_R1158_U199 );
nand NAND2_27631 ( P3_R1158_U296 , P3_R1158_U294 , P3_R1158_U292 );
not NOT1_27632 ( P3_R1158_U297 , P3_R1158_U196 );
nand NAND2_27633 ( P3_R1158_U298 , P3_R1158_U506 , P3_R1158_U57 );
nand NAND2_27634 ( P3_R1158_U299 , P3_R1158_U298 , P3_R1158_U196 );
nand NAND2_27635 ( P3_R1158_U300 , P3_U3060 , P3_R1158_U91 );
not NOT1_27636 ( P3_R1158_U301 , P3_R1158_U194 );
nand NAND2_27637 ( P3_R1158_U302 , P3_R1158_U509 , P3_R1158_U58 );
nand NAND2_27638 ( P3_R1158_U303 , P3_R1158_U302 , P3_R1158_U194 );
nand NAND2_27639 ( P3_R1158_U304 , P3_U3065 , P3_R1158_U92 );
not NOT1_27640 ( P3_R1158_U305 , P3_R1158_U192 );
nand NAND2_27641 ( P3_R1158_U306 , P3_R1158_U515 , P3_R1158_U38 );
nand NAND3_27642 ( P3_R1158_U307 , P3_R1158_U60 , P3_R1158_U59 , P3_R1158_U308 );
nand NAND2_27643 ( P3_R1158_U308 , P3_U3056 , P3_R1158_U78 );
nand NAND2_27644 ( P3_R1158_U309 , P3_R1158_U518 , P3_R1158_U39 );
nand NAND2_27645 ( P3_R1158_U310 , P3_R1158_U369 , P3_R1158_U192 );
nand NAND2_27646 ( P3_R1158_U311 , P3_R1158_U366 , P3_R1158_U307 );
not NOT1_27647 ( P3_R1158_U312 , P3_R1158_U189 );
nand NAND2_27648 ( P3_R1158_U313 , P3_R1158_U467 , P3_R1158_U37 );
nand NAND2_27649 ( P3_R1158_U314 , P3_U3052 , P3_R1158_U75 );
nand NAND2_27650 ( P3_R1158_U315 , P3_U3052 , P3_R1158_U75 );
nand NAND2_27651 ( P3_R1158_U316 , P3_R1158_U467 , P3_R1158_U37 );
not NOT1_27652 ( P3_R1158_U317 , P3_R1158_U190 );
not NOT1_27653 ( P3_R1158_U318 , P3_R1158_U191 );
nand NAND2_27654 ( P3_R1158_U319 , P3_R1158_U138 , P3_R1158_U12 );
nand NAND2_27655 ( P3_R1158_U320 , P3_U3056 , P3_R1158_U78 );
nand NAND2_27656 ( P3_R1158_U321 , P3_R1158_U515 , P3_R1158_U38 );
nand NAND2_27657 ( P3_R1158_U322 , P3_R1158_U293 , P3_R1158_U199 );
not NOT1_27658 ( P3_R1158_U323 , P3_R1158_U61 );
nand NAND2_27659 ( P3_R1158_U324 , P3_R1158_U500 , P3_R1158_U53 );
nand NAND2_27660 ( P3_R1158_U325 , P3_R1158_U324 , P3_R1158_U61 );
nand NAND2_27661 ( P3_R1158_U326 , P3_R1158_U143 , P3_R1158_U325 );
nand NAND2_27662 ( P3_R1158_U327 , P3_R1158_U323 , P3_R1158_U214 );
nand NAND2_27663 ( P3_R1158_U328 , P3_U3074 , P3_R1158_U89 );
nand NAND2_27664 ( P3_R1158_U329 , P3_R1158_U144 , P3_R1158_U327 );
nand NAND2_27665 ( P3_R1158_U330 , P3_R1158_U500 , P3_R1158_U53 );
nand NAND2_27666 ( P3_R1158_U331 , P3_R1158_U491 , P3_R1158_U41 );
nand NAND2_27667 ( P3_R1158_U332 , P3_R1158_U331 , P3_R1158_U62 );
nand NAND2_27668 ( P3_R1158_U333 , P3_R1158_U145 , P3_R1158_U332 );
nand NAND2_27669 ( P3_R1158_U334 , P3_R1158_U275 , P3_R1158_U42 );
nand NAND2_27670 ( P3_R1158_U335 , P3_U3068 , P3_R1158_U80 );
nand NAND2_27671 ( P3_R1158_U336 , P3_R1158_U146 , P3_R1158_U334 );
nand NAND2_27672 ( P3_R1158_U337 , P3_R1158_U491 , P3_R1158_U41 );
nand NAND2_27673 ( P3_R1158_U338 , P3_R1158_U267 , P3_R1158_U206 );
not NOT1_27674 ( P3_R1158_U339 , P3_R1158_U64 );
nand NAND2_27675 ( P3_R1158_U340 , P3_R1158_U479 , P3_R1158_U45 );
nand NAND2_27676 ( P3_R1158_U341 , P3_R1158_U340 , P3_R1158_U64 );
nand NAND2_27677 ( P3_R1158_U342 , P3_R1158_U147 , P3_R1158_U341 );
nand NAND2_27678 ( P3_R1158_U343 , P3_R1158_U339 , P3_R1158_U213 );
nand NAND2_27679 ( P3_R1158_U344 , P3_U3079 , P3_R1158_U83 );
nand NAND2_27680 ( P3_R1158_U345 , P3_R1158_U148 , P3_R1158_U343 );
nand NAND2_27681 ( P3_R1158_U346 , P3_R1158_U479 , P3_R1158_U45 );
nand NAND2_27682 ( P3_R1158_U347 , P3_R1158_U250 , P3_R1158_U23 );
nand NAND2_27683 ( P3_R1158_U348 , P3_R1158_U257 , P3_R1158_U28 );
nand NAND2_27684 ( P3_R1158_U349 , P3_R1158_U321 , P3_R1158_U59 );
nand NAND2_27685 ( P3_R1158_U350 , P3_R1158_U309 , P3_R1158_U60 );
nand NAND2_27686 ( P3_R1158_U351 , P3_R1158_U330 , P3_R1158_U214 );
nand NAND2_27687 ( P3_R1158_U352 , P3_R1158_U293 , P3_R1158_U55 );
nand NAND2_27688 ( P3_R1158_U353 , P3_R1158_U337 , P3_R1158_U42 );
nand NAND2_27689 ( P3_R1158_U354 , P3_R1158_U346 , P3_R1158_U213 );
nand NAND2_27690 ( P3_R1158_U355 , P3_R1158_U267 , P3_R1158_U47 );
nand NAND2_27691 ( P3_R1158_U356 , P3_U3059 , P3_R1158_U74 );
nand NAND2_27692 ( P3_R1158_U357 , P3_U3082 , P3_R1158_U65 );
nand NAND2_27693 ( P3_R1158_U358 , P3_R1158_U133 , P3_R1158_U310 );
nand NAND2_27694 ( P3_R1158_U359 , P3_R1158_U68 , P3_R1158_U240 );
nand NAND3_27695 ( P3_R1158_U360 , P3_U3076 , P3_R1158_U219 , P3_R1158_U223 );
nand NAND2_27696 ( P3_R1158_U361 , P3_R1158_U119 , P3_R1158_U223 );
nand NAND2_27697 ( P3_R1158_U362 , P3_R1158_U236 , P3_R1158_U5 );
not NOT1_27698 ( P3_R1158_U363 , P3_R1158_U34 );
nand NAND2_27699 ( P3_R1158_U364 , P3_R1158_U34 , P3_R1158_U242 );
nand NAND2_27700 ( P3_R1158_U365 , P3_R1158_U261 , P3_R1158_U9 );
nand NAND3_27701 ( P3_R1158_U366 , P3_R1158_U367 , P3_R1158_U308 , P3_R1158_U19 );
nand NAND2_27702 ( P3_R1158_U367 , P3_R1158_U78 , P3_R1158_U306 );
not NOT1_27703 ( P3_R1158_U368 , P3_R1158_U19 );
nand NAND2_27704 ( P3_R1158_U369 , P3_R1158_U371 , P3_R1158_U370 );
nand NAND3_27705 ( P3_R1158_U370 , P3_R1158_U309 , P3_R1158_U306 , P3_R1158_U78 );
nand NAND2_27706 ( P3_R1158_U371 , P3_R1158_U368 , P3_R1158_U309 );
not NOT1_27707 ( P3_R1158_U372 , P3_R1158_U63 );
nand NAND2_27708 ( P3_R1158_U373 , P3_R1158_U63 , P3_R1158_U270 );
nand NAND2_27709 ( P3_R1158_U374 , P3_R1158_U134 , P3_R1158_U366 );
nand NAND2_27710 ( P3_R1158_U375 , P3_R1158_U135 , P3_R1158_U192 );
nand NAND2_27711 ( P3_R1158_U376 , P3_R1158_U378 , P3_R1158_U377 );
nand NAND3_27712 ( P3_R1158_U377 , P3_R1158_U60 , P3_R1158_U59 , P3_R1158_U308 );
nand NAND3_27713 ( P3_R1158_U378 , P3_R1158_U367 , P3_R1158_U308 , P3_R1158_U19 );
nand NAND2_27714 ( P3_R1158_U379 , P3_R1158_U235 , P3_R1158_U165 );
not NOT1_27715 ( P3_R1158_U380 , P3_R1158_U35 );
nand NAND2_27716 ( P3_R1158_U381 , P3_R1158_U10 , P3_R1158_U165 );
not NOT1_27717 ( P3_R1158_U382 , P3_R1158_U163 );
nand NAND2_27718 ( P3_R1158_U383 , P3_R1158_U121 , P3_R1158_U165 );
not NOT1_27719 ( P3_R1158_U384 , P3_R1158_U161 );
nand NAND2_27720 ( P3_R1158_U385 , P3_R1158_U260 , P3_R1158_U208 );
not NOT1_27721 ( P3_R1158_U386 , P3_R1158_U206 );
nand NAND2_27722 ( P3_R1158_U387 , P3_R1158_U11 , P3_R1158_U208 );
not NOT1_27723 ( P3_R1158_U388 , P3_R1158_U205 );
nand NAND2_27724 ( P3_R1158_U389 , P3_R1158_U128 , P3_R1158_U208 );
not NOT1_27725 ( P3_R1158_U390 , P3_R1158_U203 );
nand NAND2_27726 ( P3_R1158_U391 , P3_R1158_U139 , P3_R1158_U209 );
nand NAND2_27727 ( P3_R1158_U392 , P3_R1158_U140 , P3_R1158_U209 );
nand NAND2_27728 ( P3_R1158_U393 , P3_U3152 , P3_R1158_U150 );
nand NAND2_27729 ( P3_R1158_U394 , P3_U3416 , P3_R1158_U20 );
not NOT1_27730 ( P3_R1158_U395 , P3_R1158_U65 );
nand NAND2_27731 ( P3_R1158_U396 , P3_R1158_U395 , P3_U3082 );
nand NAND2_27732 ( P3_R1158_U397 , P3_R1158_U65 , P3_R1158_U33 );
nand NAND2_27733 ( P3_R1158_U398 , P3_R1158_U395 , P3_U3082 );
nand NAND2_27734 ( P3_R1158_U399 , P3_R1158_U65 , P3_R1158_U33 );
nand NAND2_27735 ( P3_R1158_U400 , P3_R1158_U399 , P3_R1158_U398 );
nand NAND2_27736 ( P3_R1158_U401 , P3_U3152 , P3_R1158_U152 );
nand NAND2_27737 ( P3_R1158_U402 , P3_U3401 , P3_R1158_U20 );
not NOT1_27738 ( P3_R1158_U403 , P3_R1158_U74 );
nand NAND2_27739 ( P3_R1158_U404 , P3_U3152 , P3_R1158_U153 );
nand NAND2_27740 ( P3_R1158_U405 , P3_U3392 , P3_R1158_U20 );
not NOT1_27741 ( P3_R1158_U406 , P3_R1158_U72 );
nand NAND2_27742 ( P3_R1158_U407 , P3_U3152 , P3_R1158_U154 );
nand NAND2_27743 ( P3_R1158_U408 , P3_U3387 , P3_R1158_U20 );
not NOT1_27744 ( P3_R1158_U409 , P3_R1158_U73 );
nand NAND2_27745 ( P3_R1158_U410 , P3_U3152 , P3_R1158_U155 );
nand NAND2_27746 ( P3_R1158_U411 , P3_U3398 , P3_R1158_U20 );
not NOT1_27747 ( P3_R1158_U412 , P3_R1158_U71 );
nand NAND2_27748 ( P3_R1158_U413 , P3_U3152 , P3_R1158_U156 );
nand NAND2_27749 ( P3_R1158_U414 , P3_U3395 , P3_R1158_U20 );
not NOT1_27750 ( P3_R1158_U415 , P3_R1158_U70 );
nand NAND2_27751 ( P3_R1158_U416 , P3_U3152 , P3_R1158_U157 );
nand NAND2_27752 ( P3_R1158_U417 , P3_U3404 , P3_R1158_U20 );
not NOT1_27753 ( P3_R1158_U418 , P3_R1158_U69 );
nand NAND2_27754 ( P3_R1158_U419 , P3_U3152 , P3_R1158_U158 );
nand NAND2_27755 ( P3_R1158_U420 , P3_U3410 , P3_R1158_U20 );
not NOT1_27756 ( P3_R1158_U421 , P3_R1158_U68 );
nand NAND2_27757 ( P3_R1158_U422 , P3_U3152 , P3_R1158_U159 );
nand NAND2_27758 ( P3_R1158_U423 , P3_U3407 , P3_R1158_U20 );
not NOT1_27759 ( P3_R1158_U424 , P3_R1158_U67 );
nand NAND2_27760 ( P3_R1158_U425 , P3_U3152 , P3_R1158_U160 );
nand NAND2_27761 ( P3_R1158_U426 , P3_U3413 , P3_R1158_U20 );
not NOT1_27762 ( P3_R1158_U427 , P3_R1158_U66 );
nand NAND2_27763 ( P3_R1158_U428 , P3_R1158_U151 , P3_R1158_U161 );
nand NAND2_27764 ( P3_R1158_U429 , P3_R1158_U384 , P3_R1158_U400 );
nand NAND2_27765 ( P3_R1158_U430 , P3_R1158_U427 , P3_U3083 );
nand NAND2_27766 ( P3_R1158_U431 , P3_R1158_U66 , P3_R1158_U21 );
nand NAND2_27767 ( P3_R1158_U432 , P3_R1158_U427 , P3_U3083 );
nand NAND2_27768 ( P3_R1158_U433 , P3_R1158_U66 , P3_R1158_U21 );
nand NAND2_27769 ( P3_R1158_U434 , P3_R1158_U433 , P3_R1158_U432 );
nand NAND2_27770 ( P3_R1158_U435 , P3_R1158_U162 , P3_R1158_U163 );
nand NAND2_27771 ( P3_R1158_U436 , P3_R1158_U382 , P3_R1158_U434 );
nand NAND2_27772 ( P3_R1158_U437 , P3_R1158_U421 , P3_U3069 );
nand NAND2_27773 ( P3_R1158_U438 , P3_R1158_U68 , P3_R1158_U24 );
nand NAND2_27774 ( P3_R1158_U439 , P3_R1158_U424 , P3_U3070 );
nand NAND2_27775 ( P3_R1158_U440 , P3_R1158_U67 , P3_R1158_U22 );
nand NAND2_27776 ( P3_R1158_U441 , P3_R1158_U440 , P3_R1158_U439 );
nand NAND2_27777 ( P3_R1158_U442 , P3_R1158_U35 , P3_R1158_U347 );
nand NAND2_27778 ( P3_R1158_U443 , P3_R1158_U441 , P3_R1158_U380 );
nand NAND2_27779 ( P3_R1158_U444 , P3_R1158_U418 , P3_U3066 );
nand NAND2_27780 ( P3_R1158_U445 , P3_R1158_U69 , P3_R1158_U25 );
nand NAND2_27781 ( P3_R1158_U446 , P3_R1158_U418 , P3_U3066 );
nand NAND2_27782 ( P3_R1158_U447 , P3_R1158_U69 , P3_R1158_U25 );
nand NAND2_27783 ( P3_R1158_U448 , P3_R1158_U447 , P3_R1158_U446 );
nand NAND2_27784 ( P3_R1158_U449 , P3_R1158_U164 , P3_R1158_U165 );
nand NAND2_27785 ( P3_R1158_U450 , P3_R1158_U234 , P3_R1158_U448 );
nand NAND2_27786 ( P3_R1158_U451 , P3_R1158_U403 , P3_U3059 );
nand NAND2_27787 ( P3_R1158_U452 , P3_R1158_U74 , P3_R1158_U32 );
nand NAND2_27788 ( P3_R1158_U453 , P3_R1158_U403 , P3_U3059 );
nand NAND2_27789 ( P3_R1158_U454 , P3_R1158_U74 , P3_R1158_U32 );
nand NAND2_27790 ( P3_R1158_U455 , P3_R1158_U454 , P3_R1158_U453 );
nand NAND2_27791 ( P3_R1158_U456 , P3_R1158_U166 , P3_R1158_U167 );
nand NAND2_27792 ( P3_R1158_U457 , P3_R1158_U232 , P3_R1158_U455 );
nand NAND2_27793 ( P3_R1158_U458 , P3_R1158_U412 , P3_U3063 );
nand NAND2_27794 ( P3_R1158_U459 , P3_R1158_U71 , P3_R1158_U29 );
nand NAND2_27795 ( P3_R1158_U460 , P3_R1158_U415 , P3_U3067 );
nand NAND2_27796 ( P3_R1158_U461 , P3_R1158_U70 , P3_R1158_U27 );
nand NAND2_27797 ( P3_R1158_U462 , P3_R1158_U461 , P3_R1158_U460 );
nand NAND2_27798 ( P3_R1158_U463 , P3_R1158_U348 , P3_R1158_U36 );
nand NAND2_27799 ( P3_R1158_U464 , P3_R1158_U462 , P3_R1158_U225 );
nand NAND2_27800 ( P3_R1158_U465 , P3_U3152 , P3_R1158_U168 );
nand NAND2_27801 ( P3_R1158_U466 , P3_U3900 , P3_R1158_U20 );
not NOT1_27802 ( P3_R1158_U467 , P3_R1158_U75 );
nand NAND2_27803 ( P3_R1158_U468 , P3_U3152 , P3_R1158_U169 );
nand NAND2_27804 ( P3_R1158_U469 , P3_U3419 , P3_R1158_U20 );
not NOT1_27805 ( P3_R1158_U470 , P3_R1158_U85 );
nand NAND2_27806 ( P3_R1158_U471 , P3_U3152 , P3_R1158_U170 );
nand NAND2_27807 ( P3_R1158_U472 , P3_U3422 , P3_R1158_U20 );
not NOT1_27808 ( P3_R1158_U473 , P3_R1158_U84 );
nand NAND2_27809 ( P3_R1158_U474 , P3_U3152 , P3_R1158_U171 );
nand NAND2_27810 ( P3_R1158_U475 , P3_U3428 , P3_R1158_U20 );
not NOT1_27811 ( P3_R1158_U476 , P3_R1158_U83 );
nand NAND2_27812 ( P3_R1158_U477 , P3_U3152 , P3_R1158_U172 );
nand NAND2_27813 ( P3_R1158_U478 , P3_U3425 , P3_R1158_U20 );
not NOT1_27814 ( P3_R1158_U479 , P3_R1158_U82 );
nand NAND2_27815 ( P3_R1158_U480 , P3_U3152 , P3_R1158_U173 );
nand NAND2_27816 ( P3_R1158_U481 , P3_U3431 , P3_R1158_U20 );
not NOT1_27817 ( P3_R1158_U482 , P3_R1158_U81 );
nand NAND2_27818 ( P3_R1158_U483 , P3_U3152 , P3_R1158_U174 );
nand NAND2_27819 ( P3_R1158_U484 , P3_U3434 , P3_R1158_U20 );
not NOT1_27820 ( P3_R1158_U485 , P3_R1158_U86 );
nand NAND2_27821 ( P3_R1158_U486 , P3_U3152 , P3_R1158_U175 );
nand NAND2_27822 ( P3_R1158_U487 , P3_U3440 , P3_R1158_U20 );
not NOT1_27823 ( P3_R1158_U488 , P3_R1158_U80 );
nand NAND2_27824 ( P3_R1158_U489 , P3_U3152 , P3_R1158_U176 );
nand NAND2_27825 ( P3_R1158_U490 , P3_U3437 , P3_R1158_U20 );
not NOT1_27826 ( P3_R1158_U491 , P3_R1158_U79 );
nand NAND2_27827 ( P3_R1158_U492 , P3_U3152 , P3_R1158_U177 );
nand NAND2_27828 ( P3_R1158_U493 , P3_U3443 , P3_R1158_U20 );
not NOT1_27829 ( P3_R1158_U494 , P3_R1158_U87 );
nand NAND2_27830 ( P3_R1158_U495 , P3_U3152 , P3_R1158_U178 );
nand NAND2_27831 ( P3_R1158_U496 , P3_U3906 , P3_R1158_U20 );
not NOT1_27832 ( P3_R1158_U497 , P3_R1158_U89 );
nand NAND2_27833 ( P3_R1158_U498 , P3_U3152 , P3_R1158_U179 );
nand NAND2_27834 ( P3_R1158_U499 , P3_U3907 , P3_R1158_U20 );
not NOT1_27835 ( P3_R1158_U500 , P3_R1158_U90 );
nand NAND2_27836 ( P3_R1158_U501 , P3_U3152 , P3_R1158_U180 );
nand NAND2_27837 ( P3_R1158_U502 , P3_U3445 , P3_R1158_U20 );
not NOT1_27838 ( P3_R1158_U503 , P3_R1158_U88 );
nand NAND2_27839 ( P3_R1158_U504 , P3_U3152 , P3_R1158_U181 );
nand NAND2_27840 ( P3_R1158_U505 , P3_U3905 , P3_R1158_U20 );
not NOT1_27841 ( P3_R1158_U506 , P3_R1158_U91 );
nand NAND2_27842 ( P3_R1158_U507 , P3_U3152 , P3_R1158_U182 );
nand NAND2_27843 ( P3_R1158_U508 , P3_U3904 , P3_R1158_U20 );
not NOT1_27844 ( P3_R1158_U509 , P3_R1158_U92 );
nand NAND2_27845 ( P3_R1158_U510 , P3_U3152 , P3_R1158_U183 );
nand NAND2_27846 ( P3_R1158_U511 , P3_U3901 , P3_R1158_U20 );
not NOT1_27847 ( P3_R1158_U512 , P3_R1158_U78 );
nand NAND2_27848 ( P3_R1158_U513 , P3_U3152 , P3_R1158_U184 );
nand NAND2_27849 ( P3_R1158_U514 , P3_U3902 , P3_R1158_U20 );
not NOT1_27850 ( P3_R1158_U515 , P3_R1158_U76 );
nand NAND2_27851 ( P3_R1158_U516 , P3_U3152 , P3_R1158_U185 );
nand NAND2_27852 ( P3_R1158_U517 , P3_U3903 , P3_R1158_U20 );
not NOT1_27853 ( P3_R1158_U518 , P3_R1158_U77 );
nand NAND2_27854 ( P3_R1158_U519 , P3_U3152 , P3_R1158_U186 );
nand NAND2_27855 ( P3_R1158_U520 , P3_U3053 , P3_R1158_U20 );
not NOT1_27856 ( P3_R1158_U521 , P3_R1158_U137 );
nand NAND2_27857 ( P3_R1158_U522 , P3_U3899 , P3_R1158_U521 );
nand NAND2_27858 ( P3_R1158_U523 , P3_R1158_U137 , P3_R1158_U187 );
not NOT1_27859 ( P3_R1158_U524 , P3_R1158_U93 );
nand NAND3_27860 ( P3_R1158_U525 , P3_R1158_U358 , P3_R1158_U313 , P3_R1158_U524 );
nand NAND3_27861 ( P3_R1158_U526 , P3_R1158_U136 , P3_R1158_U375 , P3_R1158_U93 );
nand NAND2_27862 ( P3_R1158_U527 , P3_R1158_U467 , P3_U3052 );
nand NAND2_27863 ( P3_R1158_U528 , P3_R1158_U75 , P3_R1158_U37 );
nand NAND2_27864 ( P3_R1158_U529 , P3_R1158_U467 , P3_U3052 );
nand NAND2_27865 ( P3_R1158_U530 , P3_R1158_U75 , P3_R1158_U37 );
nand NAND2_27866 ( P3_R1158_U531 , P3_R1158_U530 , P3_R1158_U529 );
nand NAND2_27867 ( P3_R1158_U532 , P3_R1158_U188 , P3_R1158_U189 );
nand NAND2_27868 ( P3_R1158_U533 , P3_R1158_U312 , P3_R1158_U531 );
nand NAND2_27869 ( P3_R1158_U534 , P3_R1158_U512 , P3_U3056 );
nand NAND2_27870 ( P3_R1158_U535 , P3_R1158_U78 , P3_R1158_U40 );
nand NAND2_27871 ( P3_R1158_U536 , P3_R1158_U104 , P3_R1158_U190 );
nand NAND2_27872 ( P3_R1158_U537 , P3_R1158_U103 , P3_R1158_U317 );
nand NAND2_27873 ( P3_R1158_U538 , P3_R1158_U515 , P3_U3057 );
nand NAND2_27874 ( P3_R1158_U539 , P3_R1158_U76 , P3_R1158_U38 );
nand NAND2_27875 ( P3_R1158_U540 , P3_R1158_U539 , P3_R1158_U538 );
nand NAND2_27876 ( P3_R1158_U541 , P3_R1158_U349 , P3_R1158_U191 );
nand NAND2_27877 ( P3_R1158_U542 , P3_R1158_U318 , P3_R1158_U540 );
nand NAND2_27878 ( P3_R1158_U543 , P3_R1158_U518 , P3_U3064 );
nand NAND2_27879 ( P3_R1158_U544 , P3_R1158_U77 , P3_R1158_U39 );
nand NAND2_27880 ( P3_R1158_U545 , P3_R1158_U544 , P3_R1158_U543 );
nand NAND2_27881 ( P3_R1158_U546 , P3_R1158_U350 , P3_R1158_U192 );
nand NAND2_27882 ( P3_R1158_U547 , P3_R1158_U305 , P3_R1158_U545 );
nand NAND2_27883 ( P3_R1158_U548 , P3_R1158_U509 , P3_U3065 );
nand NAND2_27884 ( P3_R1158_U549 , P3_R1158_U92 , P3_R1158_U58 );
nand NAND2_27885 ( P3_R1158_U550 , P3_R1158_U509 , P3_U3065 );
nand NAND2_27886 ( P3_R1158_U551 , P3_R1158_U92 , P3_R1158_U58 );
nand NAND2_27887 ( P3_R1158_U552 , P3_R1158_U551 , P3_R1158_U550 );
nand NAND2_27888 ( P3_R1158_U553 , P3_R1158_U193 , P3_R1158_U194 );
nand NAND2_27889 ( P3_R1158_U554 , P3_R1158_U301 , P3_R1158_U552 );
nand NAND2_27890 ( P3_R1158_U555 , P3_R1158_U506 , P3_U3060 );
nand NAND2_27891 ( P3_R1158_U556 , P3_R1158_U91 , P3_R1158_U57 );
nand NAND2_27892 ( P3_R1158_U557 , P3_R1158_U506 , P3_U3060 );
nand NAND2_27893 ( P3_R1158_U558 , P3_R1158_U91 , P3_R1158_U57 );
nand NAND2_27894 ( P3_R1158_U559 , P3_R1158_U558 , P3_R1158_U557 );
nand NAND2_27895 ( P3_R1158_U560 , P3_R1158_U195 , P3_R1158_U196 );
nand NAND2_27896 ( P3_R1158_U561 , P3_R1158_U297 , P3_R1158_U559 );
nand NAND2_27897 ( P3_R1158_U562 , P3_R1158_U497 , P3_U3074 );
nand NAND2_27898 ( P3_R1158_U563 , P3_R1158_U89 , P3_R1158_U56 );
nand NAND2_27899 ( P3_R1158_U564 , P3_R1158_U500 , P3_U3075 );
nand NAND2_27900 ( P3_R1158_U565 , P3_R1158_U90 , P3_R1158_U53 );
nand NAND2_27901 ( P3_R1158_U566 , P3_R1158_U565 , P3_R1158_U564 );
nand NAND2_27902 ( P3_R1158_U567 , P3_R1158_U351 , P3_R1158_U61 );
nand NAND2_27903 ( P3_R1158_U568 , P3_R1158_U566 , P3_R1158_U323 );
nand NAND2_27904 ( P3_R1158_U569 , P3_R1158_U406 , P3_U3077 );
nand NAND2_27905 ( P3_R1158_U570 , P3_R1158_U72 , P3_R1158_U30 );
nand NAND2_27906 ( P3_R1158_U571 , P3_R1158_U406 , P3_U3077 );
nand NAND2_27907 ( P3_R1158_U572 , P3_R1158_U72 , P3_R1158_U30 );
nand NAND2_27908 ( P3_R1158_U573 , P3_R1158_U572 , P3_R1158_U571 );
nand NAND2_27909 ( P3_R1158_U574 , P3_R1158_U197 , P3_R1158_U198 );
nand NAND2_27910 ( P3_R1158_U575 , P3_R1158_U222 , P3_R1158_U573 );
nand NAND2_27911 ( P3_R1158_U576 , P3_R1158_U503 , P3_U3080 );
nand NAND2_27912 ( P3_R1158_U577 , P3_R1158_U88 , P3_R1158_U54 );
nand NAND2_27913 ( P3_R1158_U578 , P3_R1158_U577 , P3_R1158_U576 );
nand NAND2_27914 ( P3_R1158_U579 , P3_R1158_U352 , P3_R1158_U199 );
nand NAND2_27915 ( P3_R1158_U580 , P3_R1158_U287 , P3_R1158_U578 );
nand NAND2_27916 ( P3_R1158_U581 , P3_R1158_U494 , P3_U3081 );
nand NAND2_27917 ( P3_R1158_U582 , P3_R1158_U87 , P3_R1158_U52 );
nand NAND2_27918 ( P3_R1158_U583 , P3_R1158_U494 , P3_U3081 );
nand NAND2_27919 ( P3_R1158_U584 , P3_R1158_U87 , P3_R1158_U52 );
nand NAND2_27920 ( P3_R1158_U585 , P3_R1158_U584 , P3_R1158_U583 );
nand NAND2_27921 ( P3_R1158_U586 , P3_R1158_U200 , P3_R1158_U201 );
nand NAND2_27922 ( P3_R1158_U587 , P3_R1158_U283 , P3_R1158_U585 );
nand NAND2_27923 ( P3_R1158_U588 , P3_R1158_U488 , P3_U3068 );
nand NAND2_27924 ( P3_R1158_U589 , P3_R1158_U80 , P3_R1158_U43 );
nand NAND2_27925 ( P3_R1158_U590 , P3_R1158_U491 , P3_U3072 );
nand NAND2_27926 ( P3_R1158_U591 , P3_R1158_U79 , P3_R1158_U41 );
nand NAND2_27927 ( P3_R1158_U592 , P3_R1158_U591 , P3_R1158_U590 );
nand NAND2_27928 ( P3_R1158_U593 , P3_R1158_U353 , P3_R1158_U62 );
nand NAND2_27929 ( P3_R1158_U594 , P3_R1158_U592 , P3_R1158_U275 );
nand NAND2_27930 ( P3_R1158_U595 , P3_R1158_U485 , P3_U3073 );
nand NAND2_27931 ( P3_R1158_U596 , P3_R1158_U86 , P3_R1158_U51 );
nand NAND2_27932 ( P3_R1158_U597 , P3_R1158_U485 , P3_U3073 );
nand NAND2_27933 ( P3_R1158_U598 , P3_R1158_U86 , P3_R1158_U51 );
nand NAND2_27934 ( P3_R1158_U599 , P3_R1158_U598 , P3_R1158_U597 );
nand NAND2_27935 ( P3_R1158_U600 , P3_R1158_U202 , P3_R1158_U203 );
nand NAND2_27936 ( P3_R1158_U601 , P3_R1158_U390 , P3_R1158_U599 );
nand NAND2_27937 ( P3_R1158_U602 , P3_R1158_U482 , P3_U3078 );
nand NAND2_27938 ( P3_R1158_U603 , P3_R1158_U81 , P3_R1158_U44 );
nand NAND2_27939 ( P3_R1158_U604 , P3_R1158_U482 , P3_U3078 );
nand NAND2_27940 ( P3_R1158_U605 , P3_R1158_U81 , P3_R1158_U44 );
nand NAND2_27941 ( P3_R1158_U606 , P3_R1158_U605 , P3_R1158_U604 );
nand NAND2_27942 ( P3_R1158_U607 , P3_R1158_U204 , P3_R1158_U205 );
nand NAND2_27943 ( P3_R1158_U608 , P3_R1158_U388 , P3_R1158_U606 );
nand NAND2_27944 ( P3_R1158_U609 , P3_R1158_U476 , P3_U3079 );
nand NAND2_27945 ( P3_R1158_U610 , P3_R1158_U83 , P3_R1158_U48 );
nand NAND2_27946 ( P3_R1158_U611 , P3_R1158_U479 , P3_U3071 );
nand NAND2_27947 ( P3_R1158_U612 , P3_R1158_U82 , P3_R1158_U45 );
nand NAND2_27948 ( P3_R1158_U613 , P3_R1158_U612 , P3_R1158_U611 );
nand NAND2_27949 ( P3_R1158_U614 , P3_R1158_U354 , P3_R1158_U64 );
nand NAND2_27950 ( P3_R1158_U615 , P3_R1158_U613 , P3_R1158_U339 );
nand NAND2_27951 ( P3_R1158_U616 , P3_R1158_U473 , P3_U3062 );
nand NAND2_27952 ( P3_R1158_U617 , P3_R1158_U84 , P3_R1158_U46 );
nand NAND2_27953 ( P3_R1158_U618 , P3_R1158_U617 , P3_R1158_U616 );
nand NAND2_27954 ( P3_R1158_U619 , P3_R1158_U206 , P3_R1158_U355 );
nand NAND2_27955 ( P3_R1158_U620 , P3_R1158_U386 , P3_R1158_U618 );
nand NAND2_27956 ( P3_R1158_U621 , P3_R1158_U470 , P3_U3061 );
nand NAND2_27957 ( P3_R1158_U622 , P3_R1158_U85 , P3_R1158_U49 );
nand NAND2_27958 ( P3_R1158_U623 , P3_R1158_U470 , P3_U3061 );
nand NAND2_27959 ( P3_R1158_U624 , P3_R1158_U85 , P3_R1158_U49 );
nand NAND2_27960 ( P3_R1158_U625 , P3_R1158_U624 , P3_R1158_U623 );
nand NAND2_27961 ( P3_R1158_U626 , P3_R1158_U207 , P3_R1158_U208 );
nand NAND2_27962 ( P3_R1158_U627 , P3_R1158_U259 , P3_R1158_U625 );
nand NAND2_27963 ( P3_R1158_U628 , P3_R1158_U73 , P3_R1158_U20 );
nand NAND2_27964 ( P3_R1158_U629 , P3_R1158_U409 , P3_U3152 );
not NOT1_27965 ( P3_R1158_U630 , P3_R1158_U149 );
nand NAND2_27966 ( P3_R1158_U631 , P3_R1158_U630 , P3_U3076 );
nand NAND2_27967 ( P3_R1158_U632 , P3_R1158_U149 , P3_R1158_U31 );
and AND2_27968 ( P3_R1131_U6 , P3_R1131_U210 , P3_R1131_U209 );
and AND2_27969 ( P3_R1131_U7 , P3_R1131_U189 , P3_R1131_U245 );
and AND2_27970 ( P3_R1131_U8 , P3_R1131_U247 , P3_R1131_U246 );
and AND2_27971 ( P3_R1131_U9 , P3_R1131_U190 , P3_R1131_U262 );
and AND2_27972 ( P3_R1131_U10 , P3_R1131_U264 , P3_R1131_U263 );
and AND2_27973 ( P3_R1131_U11 , P3_R1131_U191 , P3_R1131_U286 );
and AND2_27974 ( P3_R1131_U12 , P3_R1131_U288 , P3_R1131_U287 );
and AND3_27975 ( P3_R1131_U13 , P3_R1131_U208 , P3_R1131_U194 , P3_R1131_U213 );
and AND2_27976 ( P3_R1131_U14 , P3_R1131_U218 , P3_R1131_U195 );
and AND2_27977 ( P3_R1131_U15 , P3_R1131_U392 , P3_R1131_U391 );
nand NAND2_27978 ( P3_R1131_U16 , P3_R1131_U342 , P3_R1131_U345 );
nand NAND2_27979 ( P3_R1131_U17 , P3_R1131_U331 , P3_R1131_U334 );
nand NAND2_27980 ( P3_R1131_U18 , P3_R1131_U320 , P3_R1131_U323 );
nand NAND2_27981 ( P3_R1131_U19 , P3_R1131_U312 , P3_R1131_U314 );
nand NAND3_27982 ( P3_R1131_U20 , P3_R1131_U162 , P3_R1131_U183 , P3_R1131_U351 );
nand NAND2_27983 ( P3_R1131_U21 , P3_R1131_U241 , P3_R1131_U243 );
nand NAND2_27984 ( P3_R1131_U22 , P3_R1131_U233 , P3_R1131_U236 );
nand NAND2_27985 ( P3_R1131_U23 , P3_R1131_U225 , P3_R1131_U227 );
nand NAND2_27986 ( P3_R1131_U24 , P3_R1131_U172 , P3_R1131_U348 );
not NOT1_27987 ( P3_R1131_U25 , P3_U3069 );
nand NAND2_27988 ( P3_R1131_U26 , P3_U3069 , P3_R1131_U39 );
not NOT1_27989 ( P3_R1131_U27 , P3_U3083 );
not NOT1_27990 ( P3_R1131_U28 , P3_U3413 );
not NOT1_27991 ( P3_R1131_U29 , P3_U3395 );
not NOT1_27992 ( P3_R1131_U30 , P3_U3387 );
not NOT1_27993 ( P3_R1131_U31 , P3_U3077 );
not NOT1_27994 ( P3_R1131_U32 , P3_U3398 );
not NOT1_27995 ( P3_R1131_U33 , P3_U3067 );
nand NAND2_27996 ( P3_R1131_U34 , P3_U3067 , P3_R1131_U29 );
not NOT1_27997 ( P3_R1131_U35 , P3_U3063 );
not NOT1_27998 ( P3_R1131_U36 , P3_U3404 );
not NOT1_27999 ( P3_R1131_U37 , P3_U3407 );
not NOT1_28000 ( P3_R1131_U38 , P3_U3401 );
not NOT1_28001 ( P3_R1131_U39 , P3_U3410 );
not NOT1_28002 ( P3_R1131_U40 , P3_U3070 );
not NOT1_28003 ( P3_R1131_U41 , P3_U3066 );
not NOT1_28004 ( P3_R1131_U42 , P3_U3059 );
nand NAND2_28005 ( P3_R1131_U43 , P3_U3059 , P3_R1131_U38 );
nand NAND2_28006 ( P3_R1131_U44 , P3_R1131_U214 , P3_R1131_U212 );
not NOT1_28007 ( P3_R1131_U45 , P3_U3416 );
not NOT1_28008 ( P3_R1131_U46 , P3_U3082 );
nand NAND2_28009 ( P3_R1131_U47 , P3_R1131_U44 , P3_R1131_U215 );
nand NAND2_28010 ( P3_R1131_U48 , P3_R1131_U43 , P3_R1131_U229 );
nand NAND3_28011 ( P3_R1131_U49 , P3_R1131_U201 , P3_R1131_U185 , P3_R1131_U349 );
not NOT1_28012 ( P3_R1131_U50 , P3_U3901 );
not NOT1_28013 ( P3_R1131_U51 , P3_U3422 );
not NOT1_28014 ( P3_R1131_U52 , P3_U3419 );
not NOT1_28015 ( P3_R1131_U53 , P3_U3062 );
not NOT1_28016 ( P3_R1131_U54 , P3_U3061 );
nand NAND2_28017 ( P3_R1131_U55 , P3_U3082 , P3_R1131_U45 );
not NOT1_28018 ( P3_R1131_U56 , P3_U3425 );
not NOT1_28019 ( P3_R1131_U57 , P3_U3071 );
not NOT1_28020 ( P3_R1131_U58 , P3_U3428 );
not NOT1_28021 ( P3_R1131_U59 , P3_U3079 );
not NOT1_28022 ( P3_R1131_U60 , P3_U3437 );
not NOT1_28023 ( P3_R1131_U61 , P3_U3434 );
not NOT1_28024 ( P3_R1131_U62 , P3_U3431 );
not NOT1_28025 ( P3_R1131_U63 , P3_U3072 );
not NOT1_28026 ( P3_R1131_U64 , P3_U3073 );
not NOT1_28027 ( P3_R1131_U65 , P3_U3078 );
nand NAND2_28028 ( P3_R1131_U66 , P3_U3078 , P3_R1131_U62 );
not NOT1_28029 ( P3_R1131_U67 , P3_U3440 );
not NOT1_28030 ( P3_R1131_U68 , P3_U3068 );
not NOT1_28031 ( P3_R1131_U69 , P3_U3081 );
not NOT1_28032 ( P3_R1131_U70 , P3_U3445 );
not NOT1_28033 ( P3_R1131_U71 , P3_U3080 );
not NOT1_28034 ( P3_R1131_U72 , P3_U3907 );
not NOT1_28035 ( P3_R1131_U73 , P3_U3075 );
not NOT1_28036 ( P3_R1131_U74 , P3_U3904 );
not NOT1_28037 ( P3_R1131_U75 , P3_U3905 );
not NOT1_28038 ( P3_R1131_U76 , P3_U3906 );
not NOT1_28039 ( P3_R1131_U77 , P3_U3065 );
not NOT1_28040 ( P3_R1131_U78 , P3_U3060 );
not NOT1_28041 ( P3_R1131_U79 , P3_U3074 );
nand NAND2_28042 ( P3_R1131_U80 , P3_U3074 , P3_R1131_U76 );
not NOT1_28043 ( P3_R1131_U81 , P3_U3903 );
not NOT1_28044 ( P3_R1131_U82 , P3_U3064 );
not NOT1_28045 ( P3_R1131_U83 , P3_U3902 );
not NOT1_28046 ( P3_R1131_U84 , P3_U3057 );
not NOT1_28047 ( P3_R1131_U85 , P3_U3900 );
not NOT1_28048 ( P3_R1131_U86 , P3_U3056 );
nand NAND2_28049 ( P3_R1131_U87 , P3_U3056 , P3_R1131_U50 );
not NOT1_28050 ( P3_R1131_U88 , P3_U3052 );
not NOT1_28051 ( P3_R1131_U89 , P3_U3899 );
not NOT1_28052 ( P3_R1131_U90 , P3_U3053 );
nand NAND2_28053 ( P3_R1131_U91 , P3_R1131_U302 , P3_R1131_U301 );
nand NAND2_28054 ( P3_R1131_U92 , P3_R1131_U80 , P3_R1131_U316 );
nand NAND2_28055 ( P3_R1131_U93 , P3_R1131_U66 , P3_R1131_U327 );
nand NAND2_28056 ( P3_R1131_U94 , P3_R1131_U55 , P3_R1131_U338 );
not NOT1_28057 ( P3_R1131_U95 , P3_U3076 );
nand NAND2_28058 ( P3_R1131_U96 , P3_R1131_U402 , P3_R1131_U401 );
nand NAND2_28059 ( P3_R1131_U97 , P3_R1131_U416 , P3_R1131_U415 );
nand NAND2_28060 ( P3_R1131_U98 , P3_R1131_U421 , P3_R1131_U420 );
nand NAND2_28061 ( P3_R1131_U99 , P3_R1131_U437 , P3_R1131_U436 );
nand NAND2_28062 ( P3_R1131_U100 , P3_R1131_U442 , P3_R1131_U441 );
nand NAND2_28063 ( P3_R1131_U101 , P3_R1131_U447 , P3_R1131_U446 );
nand NAND2_28064 ( P3_R1131_U102 , P3_R1131_U452 , P3_R1131_U451 );
nand NAND2_28065 ( P3_R1131_U103 , P3_R1131_U457 , P3_R1131_U456 );
nand NAND2_28066 ( P3_R1131_U104 , P3_R1131_U473 , P3_R1131_U472 );
nand NAND2_28067 ( P3_R1131_U105 , P3_R1131_U478 , P3_R1131_U477 );
nand NAND2_28068 ( P3_R1131_U106 , P3_R1131_U361 , P3_R1131_U360 );
nand NAND2_28069 ( P3_R1131_U107 , P3_R1131_U370 , P3_R1131_U369 );
nand NAND2_28070 ( P3_R1131_U108 , P3_R1131_U377 , P3_R1131_U376 );
nand NAND2_28071 ( P3_R1131_U109 , P3_R1131_U381 , P3_R1131_U380 );
nand NAND2_28072 ( P3_R1131_U110 , P3_R1131_U390 , P3_R1131_U389 );
nand NAND2_28073 ( P3_R1131_U111 , P3_R1131_U411 , P3_R1131_U410 );
nand NAND2_28074 ( P3_R1131_U112 , P3_R1131_U428 , P3_R1131_U427 );
nand NAND2_28075 ( P3_R1131_U113 , P3_R1131_U432 , P3_R1131_U431 );
nand NAND2_28076 ( P3_R1131_U114 , P3_R1131_U464 , P3_R1131_U463 );
nand NAND2_28077 ( P3_R1131_U115 , P3_R1131_U468 , P3_R1131_U467 );
nand NAND2_28078 ( P3_R1131_U116 , P3_R1131_U485 , P3_R1131_U484 );
and AND2_28079 ( P3_R1131_U117 , P3_R1131_U352 , P3_R1131_U193 );
and AND2_28080 ( P3_R1131_U118 , P3_R1131_U205 , P3_R1131_U206 );
and AND2_28081 ( P3_R1131_U119 , P3_R1131_U14 , P3_R1131_U13 );
and AND2_28082 ( P3_R1131_U120 , P3_R1131_U357 , P3_R1131_U354 );
and AND3_28083 ( P3_R1131_U121 , P3_R1131_U363 , P3_R1131_U362 , P3_R1131_U26 );
and AND2_28084 ( P3_R1131_U122 , P3_R1131_U366 , P3_R1131_U195 );
and AND2_28085 ( P3_R1131_U123 , P3_R1131_U235 , P3_R1131_U6 );
and AND2_28086 ( P3_R1131_U124 , P3_R1131_U373 , P3_R1131_U194 );
and AND3_28087 ( P3_R1131_U125 , P3_R1131_U383 , P3_R1131_U382 , P3_R1131_U34 );
and AND2_28088 ( P3_R1131_U126 , P3_R1131_U386 , P3_R1131_U193 );
and AND2_28089 ( P3_R1131_U127 , P3_R1131_U222 , P3_R1131_U7 );
and AND2_28090 ( P3_R1131_U128 , P3_R1131_U267 , P3_R1131_U9 );
and AND2_28091 ( P3_R1131_U129 , P3_R1131_U291 , P3_R1131_U11 );
and AND2_28092 ( P3_R1131_U130 , P3_R1131_U355 , P3_R1131_U192 );
and AND2_28093 ( P3_R1131_U131 , P3_R1131_U306 , P3_R1131_U307 );
and AND2_28094 ( P3_R1131_U132 , P3_R1131_U309 , P3_R1131_U395 );
and AND2_28095 ( P3_R1131_U133 , P3_R1131_U306 , P3_R1131_U307 );
and AND2_28096 ( P3_R1131_U134 , P3_R1131_U15 , P3_R1131_U310 );
nand NAND2_28097 ( P3_R1131_U135 , P3_R1131_U399 , P3_R1131_U398 );
and AND3_28098 ( P3_R1131_U136 , P3_R1131_U404 , P3_R1131_U403 , P3_R1131_U87 );
and AND2_28099 ( P3_R1131_U137 , P3_R1131_U407 , P3_R1131_U192 );
nand NAND2_28100 ( P3_R1131_U138 , P3_R1131_U413 , P3_R1131_U412 );
nand NAND2_28101 ( P3_R1131_U139 , P3_R1131_U418 , P3_R1131_U417 );
and AND2_28102 ( P3_R1131_U140 , P3_R1131_U322 , P3_R1131_U12 );
and AND2_28103 ( P3_R1131_U141 , P3_R1131_U424 , P3_R1131_U191 );
nand NAND2_28104 ( P3_R1131_U142 , P3_R1131_U434 , P3_R1131_U433 );
nand NAND2_28105 ( P3_R1131_U143 , P3_R1131_U439 , P3_R1131_U438 );
nand NAND2_28106 ( P3_R1131_U144 , P3_R1131_U444 , P3_R1131_U443 );
nand NAND2_28107 ( P3_R1131_U145 , P3_R1131_U449 , P3_R1131_U448 );
nand NAND2_28108 ( P3_R1131_U146 , P3_R1131_U454 , P3_R1131_U453 );
and AND2_28109 ( P3_R1131_U147 , P3_R1131_U333 , P3_R1131_U10 );
and AND2_28110 ( P3_R1131_U148 , P3_R1131_U460 , P3_R1131_U190 );
nand NAND2_28111 ( P3_R1131_U149 , P3_R1131_U470 , P3_R1131_U469 );
nand NAND2_28112 ( P3_R1131_U150 , P3_R1131_U475 , P3_R1131_U474 );
and AND2_28113 ( P3_R1131_U151 , P3_R1131_U344 , P3_R1131_U8 );
and AND2_28114 ( P3_R1131_U152 , P3_R1131_U481 , P3_R1131_U189 );
and AND2_28115 ( P3_R1131_U153 , P3_R1131_U359 , P3_R1131_U358 );
nand NAND2_28116 ( P3_R1131_U154 , P3_R1131_U120 , P3_R1131_U356 );
and AND2_28117 ( P3_R1131_U155 , P3_R1131_U368 , P3_R1131_U367 );
and AND2_28118 ( P3_R1131_U156 , P3_R1131_U375 , P3_R1131_U374 );
and AND2_28119 ( P3_R1131_U157 , P3_R1131_U379 , P3_R1131_U378 );
nand NAND2_28120 ( P3_R1131_U158 , P3_R1131_U118 , P3_R1131_U203 );
and AND2_28121 ( P3_R1131_U159 , P3_R1131_U388 , P3_R1131_U387 );
not NOT1_28122 ( P3_R1131_U160 , P3_U3908 );
not NOT1_28123 ( P3_R1131_U161 , P3_U3054 );
and AND2_28124 ( P3_R1131_U162 , P3_R1131_U397 , P3_R1131_U396 );
nand NAND2_28125 ( P3_R1131_U163 , P3_R1131_U131 , P3_R1131_U304 );
and AND2_28126 ( P3_R1131_U164 , P3_R1131_U409 , P3_R1131_U408 );
nand NAND2_28127 ( P3_R1131_U165 , P3_R1131_U298 , P3_R1131_U297 );
nand NAND2_28128 ( P3_R1131_U166 , P3_R1131_U294 , P3_R1131_U293 );
and AND2_28129 ( P3_R1131_U167 , P3_R1131_U426 , P3_R1131_U425 );
and AND2_28130 ( P3_R1131_U168 , P3_R1131_U430 , P3_R1131_U429 );
nand NAND2_28131 ( P3_R1131_U169 , P3_R1131_U284 , P3_R1131_U283 );
nand NAND2_28132 ( P3_R1131_U170 , P3_R1131_U280 , P3_R1131_U279 );
not NOT1_28133 ( P3_R1131_U171 , P3_U3392 );
nand NAND2_28134 ( P3_R1131_U172 , P3_U3387 , P3_R1131_U95 );
nand NAND3_28135 ( P3_R1131_U173 , P3_R1131_U276 , P3_R1131_U184 , P3_R1131_U350 );
not NOT1_28136 ( P3_R1131_U174 , P3_U3443 );
nand NAND2_28137 ( P3_R1131_U175 , P3_R1131_U274 , P3_R1131_U273 );
nand NAND2_28138 ( P3_R1131_U176 , P3_R1131_U270 , P3_R1131_U269 );
and AND2_28139 ( P3_R1131_U177 , P3_R1131_U462 , P3_R1131_U461 );
and AND2_28140 ( P3_R1131_U178 , P3_R1131_U466 , P3_R1131_U465 );
nand NAND2_28141 ( P3_R1131_U179 , P3_R1131_U260 , P3_R1131_U259 );
nand NAND2_28142 ( P3_R1131_U180 , P3_R1131_U256 , P3_R1131_U255 );
nand NAND2_28143 ( P3_R1131_U181 , P3_R1131_U252 , P3_R1131_U251 );
and AND2_28144 ( P3_R1131_U182 , P3_R1131_U483 , P3_R1131_U482 );
nand NAND2_28145 ( P3_R1131_U183 , P3_R1131_U132 , P3_R1131_U163 );
nand NAND2_28146 ( P3_R1131_U184 , P3_R1131_U175 , P3_R1131_U174 );
nand NAND2_28147 ( P3_R1131_U185 , P3_R1131_U172 , P3_R1131_U171 );
not NOT1_28148 ( P3_R1131_U186 , P3_R1131_U87 );
not NOT1_28149 ( P3_R1131_U187 , P3_R1131_U34 );
not NOT1_28150 ( P3_R1131_U188 , P3_R1131_U26 );
nand NAND2_28151 ( P3_R1131_U189 , P3_U3419 , P3_R1131_U54 );
nand NAND2_28152 ( P3_R1131_U190 , P3_U3434 , P3_R1131_U64 );
nand NAND2_28153 ( P3_R1131_U191 , P3_U3905 , P3_R1131_U78 );
nand NAND2_28154 ( P3_R1131_U192 , P3_U3901 , P3_R1131_U86 );
nand NAND2_28155 ( P3_R1131_U193 , P3_U3395 , P3_R1131_U33 );
nand NAND2_28156 ( P3_R1131_U194 , P3_U3404 , P3_R1131_U41 );
nand NAND2_28157 ( P3_R1131_U195 , P3_U3410 , P3_R1131_U25 );
not NOT1_28158 ( P3_R1131_U196 , P3_R1131_U66 );
not NOT1_28159 ( P3_R1131_U197 , P3_R1131_U80 );
not NOT1_28160 ( P3_R1131_U198 , P3_R1131_U43 );
not NOT1_28161 ( P3_R1131_U199 , P3_R1131_U55 );
not NOT1_28162 ( P3_R1131_U200 , P3_R1131_U172 );
nand NAND2_28163 ( P3_R1131_U201 , P3_U3077 , P3_R1131_U172 );
not NOT1_28164 ( P3_R1131_U202 , P3_R1131_U49 );
nand NAND2_28165 ( P3_R1131_U203 , P3_R1131_U117 , P3_R1131_U49 );
nand NAND2_28166 ( P3_R1131_U204 , P3_R1131_U35 , P3_R1131_U34 );
nand NAND2_28167 ( P3_R1131_U205 , P3_R1131_U204 , P3_R1131_U32 );
nand NAND2_28168 ( P3_R1131_U206 , P3_U3063 , P3_R1131_U187 );
not NOT1_28169 ( P3_R1131_U207 , P3_R1131_U158 );
nand NAND2_28170 ( P3_R1131_U208 , P3_U3407 , P3_R1131_U40 );
nand NAND2_28171 ( P3_R1131_U209 , P3_U3070 , P3_R1131_U37 );
nand NAND2_28172 ( P3_R1131_U210 , P3_U3066 , P3_R1131_U36 );
nand NAND2_28173 ( P3_R1131_U211 , P3_R1131_U198 , P3_R1131_U194 );
nand NAND2_28174 ( P3_R1131_U212 , P3_R1131_U6 , P3_R1131_U211 );
nand NAND2_28175 ( P3_R1131_U213 , P3_U3401 , P3_R1131_U42 );
nand NAND2_28176 ( P3_R1131_U214 , P3_U3407 , P3_R1131_U40 );
nand NAND2_28177 ( P3_R1131_U215 , P3_R1131_U13 , P3_R1131_U158 );
not NOT1_28178 ( P3_R1131_U216 , P3_R1131_U44 );
not NOT1_28179 ( P3_R1131_U217 , P3_R1131_U47 );
nand NAND2_28180 ( P3_R1131_U218 , P3_U3413 , P3_R1131_U27 );
nand NAND2_28181 ( P3_R1131_U219 , P3_R1131_U27 , P3_R1131_U26 );
nand NAND2_28182 ( P3_R1131_U220 , P3_U3083 , P3_R1131_U188 );
not NOT1_28183 ( P3_R1131_U221 , P3_R1131_U154 );
nand NAND2_28184 ( P3_R1131_U222 , P3_U3416 , P3_R1131_U46 );
nand NAND2_28185 ( P3_R1131_U223 , P3_R1131_U222 , P3_R1131_U55 );
nand NAND2_28186 ( P3_R1131_U224 , P3_R1131_U217 , P3_R1131_U26 );
nand NAND2_28187 ( P3_R1131_U225 , P3_R1131_U122 , P3_R1131_U224 );
nand NAND2_28188 ( P3_R1131_U226 , P3_R1131_U47 , P3_R1131_U195 );
nand NAND2_28189 ( P3_R1131_U227 , P3_R1131_U121 , P3_R1131_U226 );
nand NAND2_28190 ( P3_R1131_U228 , P3_R1131_U26 , P3_R1131_U195 );
nand NAND2_28191 ( P3_R1131_U229 , P3_R1131_U213 , P3_R1131_U158 );
not NOT1_28192 ( P3_R1131_U230 , P3_R1131_U48 );
nand NAND2_28193 ( P3_R1131_U231 , P3_U3066 , P3_R1131_U36 );
nand NAND2_28194 ( P3_R1131_U232 , P3_R1131_U230 , P3_R1131_U231 );
nand NAND2_28195 ( P3_R1131_U233 , P3_R1131_U124 , P3_R1131_U232 );
nand NAND2_28196 ( P3_R1131_U234 , P3_R1131_U48 , P3_R1131_U194 );
nand NAND2_28197 ( P3_R1131_U235 , P3_U3407 , P3_R1131_U40 );
nand NAND2_28198 ( P3_R1131_U236 , P3_R1131_U123 , P3_R1131_U234 );
nand NAND2_28199 ( P3_R1131_U237 , P3_U3066 , P3_R1131_U36 );
nand NAND2_28200 ( P3_R1131_U238 , P3_R1131_U194 , P3_R1131_U237 );
nand NAND2_28201 ( P3_R1131_U239 , P3_R1131_U213 , P3_R1131_U43 );
nand NAND2_28202 ( P3_R1131_U240 , P3_R1131_U202 , P3_R1131_U34 );
nand NAND2_28203 ( P3_R1131_U241 , P3_R1131_U126 , P3_R1131_U240 );
nand NAND2_28204 ( P3_R1131_U242 , P3_R1131_U49 , P3_R1131_U193 );
nand NAND2_28205 ( P3_R1131_U243 , P3_R1131_U125 , P3_R1131_U242 );
nand NAND2_28206 ( P3_R1131_U244 , P3_R1131_U193 , P3_R1131_U34 );
nand NAND2_28207 ( P3_R1131_U245 , P3_U3422 , P3_R1131_U53 );
nand NAND2_28208 ( P3_R1131_U246 , P3_U3062 , P3_R1131_U51 );
nand NAND2_28209 ( P3_R1131_U247 , P3_U3061 , P3_R1131_U52 );
nand NAND2_28210 ( P3_R1131_U248 , P3_R1131_U199 , P3_R1131_U7 );
nand NAND2_28211 ( P3_R1131_U249 , P3_R1131_U8 , P3_R1131_U248 );
nand NAND2_28212 ( P3_R1131_U250 , P3_U3422 , P3_R1131_U53 );
nand NAND2_28213 ( P3_R1131_U251 , P3_R1131_U127 , P3_R1131_U154 );
nand NAND2_28214 ( P3_R1131_U252 , P3_R1131_U250 , P3_R1131_U249 );
not NOT1_28215 ( P3_R1131_U253 , P3_R1131_U181 );
nand NAND2_28216 ( P3_R1131_U254 , P3_U3425 , P3_R1131_U57 );
nand NAND2_28217 ( P3_R1131_U255 , P3_R1131_U254 , P3_R1131_U181 );
nand NAND2_28218 ( P3_R1131_U256 , P3_U3071 , P3_R1131_U56 );
not NOT1_28219 ( P3_R1131_U257 , P3_R1131_U180 );
nand NAND2_28220 ( P3_R1131_U258 , P3_U3428 , P3_R1131_U59 );
nand NAND2_28221 ( P3_R1131_U259 , P3_R1131_U258 , P3_R1131_U180 );
nand NAND2_28222 ( P3_R1131_U260 , P3_U3079 , P3_R1131_U58 );
not NOT1_28223 ( P3_R1131_U261 , P3_R1131_U179 );
nand NAND2_28224 ( P3_R1131_U262 , P3_U3437 , P3_R1131_U63 );
nand NAND2_28225 ( P3_R1131_U263 , P3_U3072 , P3_R1131_U60 );
nand NAND2_28226 ( P3_R1131_U264 , P3_U3073 , P3_R1131_U61 );
nand NAND2_28227 ( P3_R1131_U265 , P3_R1131_U196 , P3_R1131_U9 );
nand NAND2_28228 ( P3_R1131_U266 , P3_R1131_U10 , P3_R1131_U265 );
nand NAND2_28229 ( P3_R1131_U267 , P3_U3431 , P3_R1131_U65 );
nand NAND2_28230 ( P3_R1131_U268 , P3_U3437 , P3_R1131_U63 );
nand NAND2_28231 ( P3_R1131_U269 , P3_R1131_U128 , P3_R1131_U179 );
nand NAND2_28232 ( P3_R1131_U270 , P3_R1131_U268 , P3_R1131_U266 );
not NOT1_28233 ( P3_R1131_U271 , P3_R1131_U176 );
nand NAND2_28234 ( P3_R1131_U272 , P3_U3440 , P3_R1131_U68 );
nand NAND2_28235 ( P3_R1131_U273 , P3_R1131_U272 , P3_R1131_U176 );
nand NAND2_28236 ( P3_R1131_U274 , P3_U3068 , P3_R1131_U67 );
not NOT1_28237 ( P3_R1131_U275 , P3_R1131_U175 );
nand NAND2_28238 ( P3_R1131_U276 , P3_U3081 , P3_R1131_U175 );
not NOT1_28239 ( P3_R1131_U277 , P3_R1131_U173 );
nand NAND2_28240 ( P3_R1131_U278 , P3_U3445 , P3_R1131_U71 );
nand NAND2_28241 ( P3_R1131_U279 , P3_R1131_U278 , P3_R1131_U173 );
nand NAND2_28242 ( P3_R1131_U280 , P3_U3080 , P3_R1131_U70 );
not NOT1_28243 ( P3_R1131_U281 , P3_R1131_U170 );
nand NAND2_28244 ( P3_R1131_U282 , P3_U3907 , P3_R1131_U73 );
nand NAND2_28245 ( P3_R1131_U283 , P3_R1131_U282 , P3_R1131_U170 );
nand NAND2_28246 ( P3_R1131_U284 , P3_U3075 , P3_R1131_U72 );
not NOT1_28247 ( P3_R1131_U285 , P3_R1131_U169 );
nand NAND2_28248 ( P3_R1131_U286 , P3_U3904 , P3_R1131_U77 );
nand NAND2_28249 ( P3_R1131_U287 , P3_U3065 , P3_R1131_U74 );
nand NAND2_28250 ( P3_R1131_U288 , P3_U3060 , P3_R1131_U75 );
nand NAND2_28251 ( P3_R1131_U289 , P3_R1131_U197 , P3_R1131_U11 );
nand NAND2_28252 ( P3_R1131_U290 , P3_R1131_U12 , P3_R1131_U289 );
nand NAND2_28253 ( P3_R1131_U291 , P3_U3906 , P3_R1131_U79 );
nand NAND2_28254 ( P3_R1131_U292 , P3_U3904 , P3_R1131_U77 );
nand NAND2_28255 ( P3_R1131_U293 , P3_R1131_U129 , P3_R1131_U169 );
nand NAND2_28256 ( P3_R1131_U294 , P3_R1131_U292 , P3_R1131_U290 );
not NOT1_28257 ( P3_R1131_U295 , P3_R1131_U166 );
nand NAND2_28258 ( P3_R1131_U296 , P3_U3903 , P3_R1131_U82 );
nand NAND2_28259 ( P3_R1131_U297 , P3_R1131_U296 , P3_R1131_U166 );
nand NAND2_28260 ( P3_R1131_U298 , P3_U3064 , P3_R1131_U81 );
not NOT1_28261 ( P3_R1131_U299 , P3_R1131_U165 );
nand NAND2_28262 ( P3_R1131_U300 , P3_U3902 , P3_R1131_U84 );
nand NAND2_28263 ( P3_R1131_U301 , P3_R1131_U300 , P3_R1131_U165 );
nand NAND2_28264 ( P3_R1131_U302 , P3_U3057 , P3_R1131_U83 );
not NOT1_28265 ( P3_R1131_U303 , P3_R1131_U91 );
nand NAND2_28266 ( P3_R1131_U304 , P3_R1131_U130 , P3_R1131_U91 );
nand NAND2_28267 ( P3_R1131_U305 , P3_R1131_U88 , P3_R1131_U87 );
nand NAND2_28268 ( P3_R1131_U306 , P3_R1131_U305 , P3_R1131_U85 );
nand NAND2_28269 ( P3_R1131_U307 , P3_U3052 , P3_R1131_U186 );
not NOT1_28270 ( P3_R1131_U308 , P3_R1131_U163 );
nand NAND2_28271 ( P3_R1131_U309 , P3_U3899 , P3_R1131_U90 );
nand NAND2_28272 ( P3_R1131_U310 , P3_U3053 , P3_R1131_U89 );
nand NAND2_28273 ( P3_R1131_U311 , P3_R1131_U303 , P3_R1131_U87 );
nand NAND2_28274 ( P3_R1131_U312 , P3_R1131_U137 , P3_R1131_U311 );
nand NAND2_28275 ( P3_R1131_U313 , P3_R1131_U91 , P3_R1131_U192 );
nand NAND2_28276 ( P3_R1131_U314 , P3_R1131_U136 , P3_R1131_U313 );
nand NAND2_28277 ( P3_R1131_U315 , P3_R1131_U192 , P3_R1131_U87 );
nand NAND2_28278 ( P3_R1131_U316 , P3_R1131_U291 , P3_R1131_U169 );
not NOT1_28279 ( P3_R1131_U317 , P3_R1131_U92 );
nand NAND2_28280 ( P3_R1131_U318 , P3_U3060 , P3_R1131_U75 );
nand NAND2_28281 ( P3_R1131_U319 , P3_R1131_U317 , P3_R1131_U318 );
nand NAND2_28282 ( P3_R1131_U320 , P3_R1131_U141 , P3_R1131_U319 );
nand NAND2_28283 ( P3_R1131_U321 , P3_R1131_U92 , P3_R1131_U191 );
nand NAND2_28284 ( P3_R1131_U322 , P3_U3904 , P3_R1131_U77 );
nand NAND2_28285 ( P3_R1131_U323 , P3_R1131_U140 , P3_R1131_U321 );
nand NAND2_28286 ( P3_R1131_U324 , P3_U3060 , P3_R1131_U75 );
nand NAND2_28287 ( P3_R1131_U325 , P3_R1131_U191 , P3_R1131_U324 );
nand NAND2_28288 ( P3_R1131_U326 , P3_R1131_U291 , P3_R1131_U80 );
nand NAND2_28289 ( P3_R1131_U327 , P3_R1131_U267 , P3_R1131_U179 );
not NOT1_28290 ( P3_R1131_U328 , P3_R1131_U93 );
nand NAND2_28291 ( P3_R1131_U329 , P3_U3073 , P3_R1131_U61 );
nand NAND2_28292 ( P3_R1131_U330 , P3_R1131_U328 , P3_R1131_U329 );
nand NAND2_28293 ( P3_R1131_U331 , P3_R1131_U148 , P3_R1131_U330 );
nand NAND2_28294 ( P3_R1131_U332 , P3_R1131_U93 , P3_R1131_U190 );
nand NAND2_28295 ( P3_R1131_U333 , P3_U3437 , P3_R1131_U63 );
nand NAND2_28296 ( P3_R1131_U334 , P3_R1131_U147 , P3_R1131_U332 );
nand NAND2_28297 ( P3_R1131_U335 , P3_U3073 , P3_R1131_U61 );
nand NAND2_28298 ( P3_R1131_U336 , P3_R1131_U190 , P3_R1131_U335 );
nand NAND2_28299 ( P3_R1131_U337 , P3_R1131_U267 , P3_R1131_U66 );
nand NAND2_28300 ( P3_R1131_U338 , P3_R1131_U222 , P3_R1131_U154 );
not NOT1_28301 ( P3_R1131_U339 , P3_R1131_U94 );
nand NAND2_28302 ( P3_R1131_U340 , P3_U3061 , P3_R1131_U52 );
nand NAND2_28303 ( P3_R1131_U341 , P3_R1131_U339 , P3_R1131_U340 );
nand NAND2_28304 ( P3_R1131_U342 , P3_R1131_U152 , P3_R1131_U341 );
nand NAND2_28305 ( P3_R1131_U343 , P3_R1131_U94 , P3_R1131_U189 );
nand NAND2_28306 ( P3_R1131_U344 , P3_U3422 , P3_R1131_U53 );
nand NAND2_28307 ( P3_R1131_U345 , P3_R1131_U151 , P3_R1131_U343 );
nand NAND2_28308 ( P3_R1131_U346 , P3_U3061 , P3_R1131_U52 );
nand NAND2_28309 ( P3_R1131_U347 , P3_R1131_U189 , P3_R1131_U346 );
nand NAND2_28310 ( P3_R1131_U348 , P3_U3076 , P3_R1131_U30 );
nand NAND2_28311 ( P3_R1131_U349 , P3_U3077 , P3_R1131_U171 );
nand NAND2_28312 ( P3_R1131_U350 , P3_U3081 , P3_R1131_U174 );
nand NAND3_28313 ( P3_R1131_U351 , P3_R1131_U133 , P3_R1131_U304 , P3_R1131_U134 );
nand NAND2_28314 ( P3_R1131_U352 , P3_U3398 , P3_R1131_U35 );
nand NAND2_28315 ( P3_R1131_U353 , P3_U3413 , P3_R1131_U220 );
nand NAND2_28316 ( P3_R1131_U354 , P3_R1131_U353 , P3_R1131_U219 );
nand NAND2_28317 ( P3_R1131_U355 , P3_U3900 , P3_R1131_U88 );
nand NAND2_28318 ( P3_R1131_U356 , P3_R1131_U119 , P3_R1131_U158 );
nand NAND2_28319 ( P3_R1131_U357 , P3_R1131_U216 , P3_R1131_U14 );
nand NAND2_28320 ( P3_R1131_U358 , P3_U3416 , P3_R1131_U46 );
nand NAND2_28321 ( P3_R1131_U359 , P3_U3082 , P3_R1131_U45 );
nand NAND2_28322 ( P3_R1131_U360 , P3_R1131_U223 , P3_R1131_U154 );
nand NAND2_28323 ( P3_R1131_U361 , P3_R1131_U221 , P3_R1131_U153 );
nand NAND2_28324 ( P3_R1131_U362 , P3_U3413 , P3_R1131_U27 );
nand NAND2_28325 ( P3_R1131_U363 , P3_U3083 , P3_R1131_U28 );
nand NAND2_28326 ( P3_R1131_U364 , P3_U3413 , P3_R1131_U27 );
nand NAND2_28327 ( P3_R1131_U365 , P3_U3083 , P3_R1131_U28 );
nand NAND2_28328 ( P3_R1131_U366 , P3_R1131_U365 , P3_R1131_U364 );
nand NAND2_28329 ( P3_R1131_U367 , P3_U3410 , P3_R1131_U25 );
nand NAND2_28330 ( P3_R1131_U368 , P3_U3069 , P3_R1131_U39 );
nand NAND2_28331 ( P3_R1131_U369 , P3_R1131_U228 , P3_R1131_U47 );
nand NAND2_28332 ( P3_R1131_U370 , P3_R1131_U155 , P3_R1131_U217 );
nand NAND2_28333 ( P3_R1131_U371 , P3_U3407 , P3_R1131_U40 );
nand NAND2_28334 ( P3_R1131_U372 , P3_U3070 , P3_R1131_U37 );
nand NAND2_28335 ( P3_R1131_U373 , P3_R1131_U372 , P3_R1131_U371 );
nand NAND2_28336 ( P3_R1131_U374 , P3_U3404 , P3_R1131_U41 );
nand NAND2_28337 ( P3_R1131_U375 , P3_U3066 , P3_R1131_U36 );
nand NAND2_28338 ( P3_R1131_U376 , P3_R1131_U238 , P3_R1131_U48 );
nand NAND2_28339 ( P3_R1131_U377 , P3_R1131_U156 , P3_R1131_U230 );
nand NAND2_28340 ( P3_R1131_U378 , P3_U3401 , P3_R1131_U42 );
nand NAND2_28341 ( P3_R1131_U379 , P3_U3059 , P3_R1131_U38 );
nand NAND2_28342 ( P3_R1131_U380 , P3_R1131_U239 , P3_R1131_U158 );
nand NAND2_28343 ( P3_R1131_U381 , P3_R1131_U207 , P3_R1131_U157 );
nand NAND2_28344 ( P3_R1131_U382 , P3_U3398 , P3_R1131_U35 );
nand NAND2_28345 ( P3_R1131_U383 , P3_U3063 , P3_R1131_U32 );
nand NAND2_28346 ( P3_R1131_U384 , P3_U3398 , P3_R1131_U35 );
nand NAND2_28347 ( P3_R1131_U385 , P3_U3063 , P3_R1131_U32 );
nand NAND2_28348 ( P3_R1131_U386 , P3_R1131_U385 , P3_R1131_U384 );
nand NAND2_28349 ( P3_R1131_U387 , P3_U3395 , P3_R1131_U33 );
nand NAND2_28350 ( P3_R1131_U388 , P3_U3067 , P3_R1131_U29 );
nand NAND2_28351 ( P3_R1131_U389 , P3_R1131_U244 , P3_R1131_U49 );
nand NAND2_28352 ( P3_R1131_U390 , P3_R1131_U159 , P3_R1131_U202 );
nand NAND2_28353 ( P3_R1131_U391 , P3_U3908 , P3_R1131_U161 );
nand NAND2_28354 ( P3_R1131_U392 , P3_U3054 , P3_R1131_U160 );
nand NAND2_28355 ( P3_R1131_U393 , P3_U3908 , P3_R1131_U161 );
nand NAND2_28356 ( P3_R1131_U394 , P3_U3054 , P3_R1131_U160 );
nand NAND2_28357 ( P3_R1131_U395 , P3_R1131_U394 , P3_R1131_U393 );
nand NAND3_28358 ( P3_R1131_U396 , P3_U3053 , P3_R1131_U395 , P3_R1131_U89 );
nand NAND3_28359 ( P3_R1131_U397 , P3_R1131_U15 , P3_R1131_U90 , P3_U3899 );
nand NAND2_28360 ( P3_R1131_U398 , P3_U3899 , P3_R1131_U90 );
nand NAND2_28361 ( P3_R1131_U399 , P3_U3053 , P3_R1131_U89 );
not NOT1_28362 ( P3_R1131_U400 , P3_R1131_U135 );
nand NAND2_28363 ( P3_R1131_U401 , P3_R1131_U308 , P3_R1131_U400 );
nand NAND2_28364 ( P3_R1131_U402 , P3_R1131_U135 , P3_R1131_U163 );
nand NAND2_28365 ( P3_R1131_U403 , P3_U3900 , P3_R1131_U88 );
nand NAND2_28366 ( P3_R1131_U404 , P3_U3052 , P3_R1131_U85 );
nand NAND2_28367 ( P3_R1131_U405 , P3_U3900 , P3_R1131_U88 );
nand NAND2_28368 ( P3_R1131_U406 , P3_U3052 , P3_R1131_U85 );
nand NAND2_28369 ( P3_R1131_U407 , P3_R1131_U406 , P3_R1131_U405 );
nand NAND2_28370 ( P3_R1131_U408 , P3_U3901 , P3_R1131_U86 );
nand NAND2_28371 ( P3_R1131_U409 , P3_U3056 , P3_R1131_U50 );
nand NAND2_28372 ( P3_R1131_U410 , P3_R1131_U315 , P3_R1131_U91 );
nand NAND2_28373 ( P3_R1131_U411 , P3_R1131_U164 , P3_R1131_U303 );
nand NAND2_28374 ( P3_R1131_U412 , P3_U3902 , P3_R1131_U84 );
nand NAND2_28375 ( P3_R1131_U413 , P3_U3057 , P3_R1131_U83 );
not NOT1_28376 ( P3_R1131_U414 , P3_R1131_U138 );
nand NAND2_28377 ( P3_R1131_U415 , P3_R1131_U299 , P3_R1131_U414 );
nand NAND2_28378 ( P3_R1131_U416 , P3_R1131_U138 , P3_R1131_U165 );
nand NAND2_28379 ( P3_R1131_U417 , P3_U3903 , P3_R1131_U82 );
nand NAND2_28380 ( P3_R1131_U418 , P3_U3064 , P3_R1131_U81 );
not NOT1_28381 ( P3_R1131_U419 , P3_R1131_U139 );
nand NAND2_28382 ( P3_R1131_U420 , P3_R1131_U295 , P3_R1131_U419 );
nand NAND2_28383 ( P3_R1131_U421 , P3_R1131_U139 , P3_R1131_U166 );
nand NAND2_28384 ( P3_R1131_U422 , P3_U3904 , P3_R1131_U77 );
nand NAND2_28385 ( P3_R1131_U423 , P3_U3065 , P3_R1131_U74 );
nand NAND2_28386 ( P3_R1131_U424 , P3_R1131_U423 , P3_R1131_U422 );
nand NAND2_28387 ( P3_R1131_U425 , P3_U3905 , P3_R1131_U78 );
nand NAND2_28388 ( P3_R1131_U426 , P3_U3060 , P3_R1131_U75 );
nand NAND2_28389 ( P3_R1131_U427 , P3_R1131_U325 , P3_R1131_U92 );
nand NAND2_28390 ( P3_R1131_U428 , P3_R1131_U167 , P3_R1131_U317 );
nand NAND2_28391 ( P3_R1131_U429 , P3_U3906 , P3_R1131_U79 );
nand NAND2_28392 ( P3_R1131_U430 , P3_U3074 , P3_R1131_U76 );
nand NAND2_28393 ( P3_R1131_U431 , P3_R1131_U326 , P3_R1131_U169 );
nand NAND2_28394 ( P3_R1131_U432 , P3_R1131_U285 , P3_R1131_U168 );
nand NAND2_28395 ( P3_R1131_U433 , P3_U3907 , P3_R1131_U73 );
nand NAND2_28396 ( P3_R1131_U434 , P3_U3075 , P3_R1131_U72 );
not NOT1_28397 ( P3_R1131_U435 , P3_R1131_U142 );
nand NAND2_28398 ( P3_R1131_U436 , P3_R1131_U281 , P3_R1131_U435 );
nand NAND2_28399 ( P3_R1131_U437 , P3_R1131_U142 , P3_R1131_U170 );
nand NAND2_28400 ( P3_R1131_U438 , P3_U3392 , P3_R1131_U31 );
nand NAND2_28401 ( P3_R1131_U439 , P3_U3077 , P3_R1131_U171 );
not NOT1_28402 ( P3_R1131_U440 , P3_R1131_U143 );
nand NAND2_28403 ( P3_R1131_U441 , P3_R1131_U200 , P3_R1131_U440 );
nand NAND2_28404 ( P3_R1131_U442 , P3_R1131_U143 , P3_R1131_U172 );
nand NAND2_28405 ( P3_R1131_U443 , P3_U3445 , P3_R1131_U71 );
nand NAND2_28406 ( P3_R1131_U444 , P3_U3080 , P3_R1131_U70 );
not NOT1_28407 ( P3_R1131_U445 , P3_R1131_U144 );
nand NAND2_28408 ( P3_R1131_U446 , P3_R1131_U277 , P3_R1131_U445 );
nand NAND2_28409 ( P3_R1131_U447 , P3_R1131_U144 , P3_R1131_U173 );
nand NAND2_28410 ( P3_R1131_U448 , P3_U3443 , P3_R1131_U69 );
nand NAND2_28411 ( P3_R1131_U449 , P3_U3081 , P3_R1131_U174 );
not NOT1_28412 ( P3_R1131_U450 , P3_R1131_U145 );
nand NAND2_28413 ( P3_R1131_U451 , P3_R1131_U275 , P3_R1131_U450 );
nand NAND2_28414 ( P3_R1131_U452 , P3_R1131_U145 , P3_R1131_U175 );
nand NAND2_28415 ( P3_R1131_U453 , P3_U3440 , P3_R1131_U68 );
nand NAND2_28416 ( P3_R1131_U454 , P3_U3068 , P3_R1131_U67 );
not NOT1_28417 ( P3_R1131_U455 , P3_R1131_U146 );
nand NAND2_28418 ( P3_R1131_U456 , P3_R1131_U271 , P3_R1131_U455 );
nand NAND2_28419 ( P3_R1131_U457 , P3_R1131_U146 , P3_R1131_U176 );
nand NAND2_28420 ( P3_R1131_U458 , P3_U3437 , P3_R1131_U63 );
nand NAND2_28421 ( P3_R1131_U459 , P3_U3072 , P3_R1131_U60 );
nand NAND2_28422 ( P3_R1131_U460 , P3_R1131_U459 , P3_R1131_U458 );
nand NAND2_28423 ( P3_R1131_U461 , P3_U3434 , P3_R1131_U64 );
nand NAND2_28424 ( P3_R1131_U462 , P3_U3073 , P3_R1131_U61 );
nand NAND2_28425 ( P3_R1131_U463 , P3_R1131_U336 , P3_R1131_U93 );
nand NAND2_28426 ( P3_R1131_U464 , P3_R1131_U177 , P3_R1131_U328 );
nand NAND2_28427 ( P3_R1131_U465 , P3_U3431 , P3_R1131_U65 );
nand NAND2_28428 ( P3_R1131_U466 , P3_U3078 , P3_R1131_U62 );
nand NAND2_28429 ( P3_R1131_U467 , P3_R1131_U337 , P3_R1131_U179 );
nand NAND2_28430 ( P3_R1131_U468 , P3_R1131_U261 , P3_R1131_U178 );
nand NAND2_28431 ( P3_R1131_U469 , P3_U3428 , P3_R1131_U59 );
nand NAND2_28432 ( P3_R1131_U470 , P3_U3079 , P3_R1131_U58 );
not NOT1_28433 ( P3_R1131_U471 , P3_R1131_U149 );
nand NAND2_28434 ( P3_R1131_U472 , P3_R1131_U257 , P3_R1131_U471 );
nand NAND2_28435 ( P3_R1131_U473 , P3_R1131_U149 , P3_R1131_U180 );
nand NAND2_28436 ( P3_R1131_U474 , P3_U3425 , P3_R1131_U57 );
nand NAND2_28437 ( P3_R1131_U475 , P3_U3071 , P3_R1131_U56 );
not NOT1_28438 ( P3_R1131_U476 , P3_R1131_U150 );
nand NAND2_28439 ( P3_R1131_U477 , P3_R1131_U253 , P3_R1131_U476 );
nand NAND2_28440 ( P3_R1131_U478 , P3_R1131_U150 , P3_R1131_U181 );
nand NAND2_28441 ( P3_R1131_U479 , P3_U3422 , P3_R1131_U53 );
nand NAND2_28442 ( P3_R1131_U480 , P3_U3062 , P3_R1131_U51 );
nand NAND2_28443 ( P3_R1131_U481 , P3_R1131_U480 , P3_R1131_U479 );
nand NAND2_28444 ( P3_R1131_U482 , P3_U3419 , P3_R1131_U54 );
nand NAND2_28445 ( P3_R1131_U483 , P3_U3061 , P3_R1131_U52 );
nand NAND2_28446 ( P3_R1131_U484 , P3_R1131_U347 , P3_R1131_U94 );
nand NAND2_28447 ( P3_R1131_U485 , P3_R1131_U182 , P3_R1131_U339 );
and AND2_28448 ( P3_R1054_U6 , P3_R1054_U102 , P3_R1054_U118 );
and AND2_28449 ( P3_R1054_U7 , P3_R1054_U120 , P3_R1054_U119 );
and AND2_28450 ( P3_R1054_U8 , P3_R1054_U99 , P3_R1054_U157 );
and AND2_28451 ( P3_R1054_U9 , P3_R1054_U159 , P3_R1054_U158 );
and AND2_28452 ( P3_R1054_U10 , P3_R1054_U100 , P3_R1054_U174 );
and AND2_28453 ( P3_R1054_U11 , P3_R1054_U176 , P3_R1054_U175 );
nand NAND2_28454 ( P3_R1054_U12 , P3_R1054_U207 , P3_R1054_U210 );
nand NAND2_28455 ( P3_R1054_U13 , P3_R1054_U196 , P3_R1054_U199 );
nand NAND2_28456 ( P3_R1054_U14 , P3_R1054_U153 , P3_R1054_U155 );
nand NAND2_28457 ( P3_R1054_U15 , P3_R1054_U145 , P3_R1054_U148 );
nand NAND2_28458 ( P3_R1054_U16 , P3_R1054_U137 , P3_R1054_U139 );
nand NAND2_28459 ( P3_R1054_U17 , P3_R1054_U21 , P3_R1054_U213 );
not NOT1_28460 ( P3_R1054_U18 , P3_U3409 );
not NOT1_28461 ( P3_R1054_U19 , P3_U3394 );
not NOT1_28462 ( P3_R1054_U20 , P3_U3386 );
nand NAND2_28463 ( P3_R1054_U21 , P3_U3386 , P3_R1054_U65 );
not NOT1_28464 ( P3_R1054_U22 , P3_U3573 );
not NOT1_28465 ( P3_R1054_U23 , P3_U3397 );
not NOT1_28466 ( P3_R1054_U24 , P3_U3562 );
nand NAND2_28467 ( P3_R1054_U25 , P3_U3562 , P3_R1054_U19 );
not NOT1_28468 ( P3_R1054_U26 , P3_U3561 );
not NOT1_28469 ( P3_R1054_U27 , P3_U3406 );
not NOT1_28470 ( P3_R1054_U28 , P3_U3403 );
not NOT1_28471 ( P3_R1054_U29 , P3_U3400 );
not NOT1_28472 ( P3_R1054_U30 , P3_U3558 );
not NOT1_28473 ( P3_R1054_U31 , P3_U3559 );
not NOT1_28474 ( P3_R1054_U32 , P3_U3560 );
nand NAND2_28475 ( P3_R1054_U33 , P3_U3560 , P3_R1054_U29 );
not NOT1_28476 ( P3_R1054_U34 , P3_U3412 );
not NOT1_28477 ( P3_R1054_U35 , P3_U3557 );
nand NAND2_28478 ( P3_R1054_U36 , P3_U3557 , P3_R1054_U18 );
not NOT1_28479 ( P3_R1054_U37 , P3_U3556 );
not NOT1_28480 ( P3_R1054_U38 , P3_U3415 );
not NOT1_28481 ( P3_R1054_U39 , P3_U3555 );
nand NAND2_28482 ( P3_R1054_U40 , P3_R1054_U126 , P3_R1054_U125 );
nand NAND2_28483 ( P3_R1054_U41 , P3_R1054_U33 , P3_R1054_U141 );
nand NAND2_28484 ( P3_R1054_U42 , P3_R1054_U110 , P3_R1054_U109 );
not NOT1_28485 ( P3_R1054_U43 , P3_U3421 );
not NOT1_28486 ( P3_R1054_U44 , P3_U3418 );
not NOT1_28487 ( P3_R1054_U45 , P3_U3571 );
not NOT1_28488 ( P3_R1054_U46 , P3_U3572 );
nand NAND2_28489 ( P3_R1054_U47 , P3_U3555 , P3_R1054_U38 );
not NOT1_28490 ( P3_R1054_U48 , P3_U3424 );
not NOT1_28491 ( P3_R1054_U49 , P3_U3570 );
not NOT1_28492 ( P3_R1054_U50 , P3_U3427 );
not NOT1_28493 ( P3_R1054_U51 , P3_U3569 );
not NOT1_28494 ( P3_R1054_U52 , P3_U3436 );
not NOT1_28495 ( P3_R1054_U53 , P3_U3433 );
not NOT1_28496 ( P3_R1054_U54 , P3_U3430 );
not NOT1_28497 ( P3_R1054_U55 , P3_U3566 );
not NOT1_28498 ( P3_R1054_U56 , P3_U3567 );
not NOT1_28499 ( P3_R1054_U57 , P3_U3568 );
nand NAND2_28500 ( P3_R1054_U58 , P3_U3568 , P3_R1054_U54 );
not NOT1_28501 ( P3_R1054_U59 , P3_U3439 );
not NOT1_28502 ( P3_R1054_U60 , P3_U3565 );
nand NAND2_28503 ( P3_R1054_U61 , P3_R1054_U186 , P3_R1054_U185 );
not NOT1_28504 ( P3_R1054_U62 , P3_U3564 );
nand NAND2_28505 ( P3_R1054_U63 , P3_R1054_U58 , P3_R1054_U192 );
nand NAND2_28506 ( P3_R1054_U64 , P3_R1054_U47 , P3_R1054_U203 );
not NOT1_28507 ( P3_R1054_U65 , P3_U3574 );
nand NAND2_28508 ( P3_R1054_U66 , P3_R1054_U251 , P3_R1054_U250 );
nand NAND2_28509 ( P3_R1054_U67 , P3_R1054_U256 , P3_R1054_U255 );
nand NAND2_28510 ( P3_R1054_U68 , P3_R1054_U261 , P3_R1054_U260 );
nand NAND2_28511 ( P3_R1054_U69 , P3_R1054_U266 , P3_R1054_U265 );
nand NAND2_28512 ( P3_R1054_U70 , P3_R1054_U282 , P3_R1054_U281 );
nand NAND2_28513 ( P3_R1054_U71 , P3_R1054_U287 , P3_R1054_U286 );
nand NAND2_28514 ( P3_R1054_U72 , P3_R1054_U217 , P3_R1054_U216 );
nand NAND2_28515 ( P3_R1054_U73 , P3_R1054_U226 , P3_R1054_U225 );
nand NAND2_28516 ( P3_R1054_U74 , P3_R1054_U233 , P3_R1054_U232 );
nand NAND2_28517 ( P3_R1054_U75 , P3_R1054_U237 , P3_R1054_U236 );
nand NAND2_28518 ( P3_R1054_U76 , P3_R1054_U246 , P3_R1054_U245 );
nand NAND2_28519 ( P3_R1054_U77 , P3_R1054_U273 , P3_R1054_U272 );
nand NAND2_28520 ( P3_R1054_U78 , P3_R1054_U277 , P3_R1054_U276 );
nand NAND2_28521 ( P3_R1054_U79 , P3_R1054_U294 , P3_R1054_U293 );
nand NAND2_28522 ( P3_R1054_U80 , P3_R1054_U248 , P3_R1054_U247 );
nand NAND2_28523 ( P3_R1054_U81 , P3_R1054_U253 , P3_R1054_U252 );
nand NAND2_28524 ( P3_R1054_U82 , P3_R1054_U258 , P3_R1054_U257 );
nand NAND2_28525 ( P3_R1054_U83 , P3_R1054_U263 , P3_R1054_U262 );
nand NAND2_28526 ( P3_R1054_U84 , P3_R1054_U279 , P3_R1054_U278 );
nand NAND2_28527 ( P3_R1054_U85 , P3_R1054_U284 , P3_R1054_U283 );
nand NAND3_28528 ( P3_R1054_U86 , P3_R1054_U131 , P3_R1054_U132 , P3_R1054_U129 );
nand NAND3_28529 ( P3_R1054_U87 , P3_R1054_U115 , P3_R1054_U116 , P3_R1054_U113 );
not NOT1_28530 ( P3_R1054_U88 , P3_U3391 );
not NOT1_28531 ( P3_R1054_U89 , P3_U3379 );
not NOT1_28532 ( P3_R1054_U90 , P3_U3563 );
nand NAND2_28533 ( P3_R1054_U91 , P3_R1054_U190 , P3_R1054_U189 );
not NOT1_28534 ( P3_R1054_U92 , P3_U3442 );
nand NAND2_28535 ( P3_R1054_U93 , P3_R1054_U182 , P3_R1054_U181 );
nand NAND2_28536 ( P3_R1054_U94 , P3_R1054_U172 , P3_R1054_U171 );
nand NAND2_28537 ( P3_R1054_U95 , P3_R1054_U168 , P3_R1054_U167 );
nand NAND2_28538 ( P3_R1054_U96 , P3_R1054_U164 , P3_R1054_U163 );
not NOT1_28539 ( P3_R1054_U97 , P3_R1054_U25 );
not NOT1_28540 ( P3_R1054_U98 , P3_R1054_U36 );
nand NAND2_28541 ( P3_R1054_U99 , P3_U3418 , P3_R1054_U46 );
nand NAND2_28542 ( P3_R1054_U100 , P3_U3433 , P3_R1054_U56 );
nand NAND2_28543 ( P3_R1054_U101 , P3_U3394 , P3_R1054_U24 );
nand NAND2_28544 ( P3_R1054_U102 , P3_U3403 , P3_R1054_U31 );
nand NAND2_28545 ( P3_R1054_U103 , P3_U3409 , P3_R1054_U35 );
not NOT1_28546 ( P3_R1054_U104 , P3_R1054_U58 );
not NOT1_28547 ( P3_R1054_U105 , P3_R1054_U33 );
not NOT1_28548 ( P3_R1054_U106 , P3_R1054_U47 );
not NOT1_28549 ( P3_R1054_U107 , P3_R1054_U21 );
nand NAND2_28550 ( P3_R1054_U108 , P3_R1054_U107 , P3_R1054_U22 );
nand NAND2_28551 ( P3_R1054_U109 , P3_R1054_U108 , P3_R1054_U88 );
nand NAND2_28552 ( P3_R1054_U110 , P3_U3573 , P3_R1054_U21 );
not NOT1_28553 ( P3_R1054_U111 , P3_R1054_U42 );
nand NAND2_28554 ( P3_R1054_U112 , P3_U3397 , P3_R1054_U26 );
nand NAND3_28555 ( P3_R1054_U113 , P3_R1054_U112 , P3_R1054_U101 , P3_R1054_U42 );
nand NAND2_28556 ( P3_R1054_U114 , P3_R1054_U26 , P3_R1054_U25 );
nand NAND2_28557 ( P3_R1054_U115 , P3_R1054_U114 , P3_R1054_U23 );
nand NAND2_28558 ( P3_R1054_U116 , P3_U3561 , P3_R1054_U97 );
not NOT1_28559 ( P3_R1054_U117 , P3_R1054_U87 );
nand NAND2_28560 ( P3_R1054_U118 , P3_U3406 , P3_R1054_U30 );
nand NAND2_28561 ( P3_R1054_U119 , P3_U3558 , P3_R1054_U27 );
nand NAND2_28562 ( P3_R1054_U120 , P3_U3559 , P3_R1054_U28 );
nand NAND2_28563 ( P3_R1054_U121 , P3_R1054_U105 , P3_R1054_U6 );
nand NAND2_28564 ( P3_R1054_U122 , P3_R1054_U7 , P3_R1054_U121 );
nand NAND2_28565 ( P3_R1054_U123 , P3_U3400 , P3_R1054_U32 );
nand NAND2_28566 ( P3_R1054_U124 , P3_U3406 , P3_R1054_U30 );
nand NAND3_28567 ( P3_R1054_U125 , P3_R1054_U123 , P3_R1054_U6 , P3_R1054_U87 );
nand NAND2_28568 ( P3_R1054_U126 , P3_R1054_U124 , P3_R1054_U122 );
not NOT1_28569 ( P3_R1054_U127 , P3_R1054_U40 );
nand NAND2_28570 ( P3_R1054_U128 , P3_U3412 , P3_R1054_U37 );
nand NAND3_28571 ( P3_R1054_U129 , P3_R1054_U128 , P3_R1054_U103 , P3_R1054_U40 );
nand NAND2_28572 ( P3_R1054_U130 , P3_R1054_U37 , P3_R1054_U36 );
nand NAND2_28573 ( P3_R1054_U131 , P3_R1054_U130 , P3_R1054_U34 );
nand NAND2_28574 ( P3_R1054_U132 , P3_U3556 , P3_R1054_U98 );
not NOT1_28575 ( P3_R1054_U133 , P3_R1054_U86 );
nand NAND2_28576 ( P3_R1054_U134 , P3_U3415 , P3_R1054_U39 );
nand NAND2_28577 ( P3_R1054_U135 , P3_R1054_U134 , P3_R1054_U47 );
nand NAND2_28578 ( P3_R1054_U136 , P3_R1054_U127 , P3_R1054_U36 );
nand NAND3_28579 ( P3_R1054_U137 , P3_R1054_U222 , P3_R1054_U103 , P3_R1054_U136 );
nand NAND2_28580 ( P3_R1054_U138 , P3_R1054_U40 , P3_R1054_U103 );
nand NAND4_28581 ( P3_R1054_U139 , P3_R1054_U219 , P3_R1054_U218 , P3_R1054_U36 , P3_R1054_U138 );
nand NAND2_28582 ( P3_R1054_U140 , P3_R1054_U36 , P3_R1054_U103 );
nand NAND2_28583 ( P3_R1054_U141 , P3_R1054_U123 , P3_R1054_U87 );
not NOT1_28584 ( P3_R1054_U142 , P3_R1054_U41 );
nand NAND2_28585 ( P3_R1054_U143 , P3_U3559 , P3_R1054_U28 );
nand NAND2_28586 ( P3_R1054_U144 , P3_R1054_U142 , P3_R1054_U143 );
nand NAND3_28587 ( P3_R1054_U145 , P3_R1054_U229 , P3_R1054_U102 , P3_R1054_U144 );
nand NAND2_28588 ( P3_R1054_U146 , P3_R1054_U41 , P3_R1054_U102 );
nand NAND2_28589 ( P3_R1054_U147 , P3_U3406 , P3_R1054_U30 );
nand NAND3_28590 ( P3_R1054_U148 , P3_R1054_U147 , P3_R1054_U7 , P3_R1054_U146 );
nand NAND2_28591 ( P3_R1054_U149 , P3_U3559 , P3_R1054_U28 );
nand NAND2_28592 ( P3_R1054_U150 , P3_R1054_U102 , P3_R1054_U149 );
nand NAND2_28593 ( P3_R1054_U151 , P3_R1054_U123 , P3_R1054_U33 );
nand NAND2_28594 ( P3_R1054_U152 , P3_R1054_U111 , P3_R1054_U25 );
nand NAND3_28595 ( P3_R1054_U153 , P3_R1054_U242 , P3_R1054_U101 , P3_R1054_U152 );
nand NAND2_28596 ( P3_R1054_U154 , P3_R1054_U42 , P3_R1054_U101 );
nand NAND4_28597 ( P3_R1054_U155 , P3_R1054_U239 , P3_R1054_U238 , P3_R1054_U25 , P3_R1054_U154 );
nand NAND2_28598 ( P3_R1054_U156 , P3_R1054_U25 , P3_R1054_U101 );
nand NAND2_28599 ( P3_R1054_U157 , P3_U3421 , P3_R1054_U45 );
nand NAND2_28600 ( P3_R1054_U158 , P3_U3571 , P3_R1054_U43 );
nand NAND2_28601 ( P3_R1054_U159 , P3_U3572 , P3_R1054_U44 );
nand NAND2_28602 ( P3_R1054_U160 , P3_R1054_U106 , P3_R1054_U8 );
nand NAND2_28603 ( P3_R1054_U161 , P3_R1054_U9 , P3_R1054_U160 );
nand NAND2_28604 ( P3_R1054_U162 , P3_U3421 , P3_R1054_U45 );
nand NAND3_28605 ( P3_R1054_U163 , P3_R1054_U134 , P3_R1054_U8 , P3_R1054_U86 );
nand NAND2_28606 ( P3_R1054_U164 , P3_R1054_U162 , P3_R1054_U161 );
not NOT1_28607 ( P3_R1054_U165 , P3_R1054_U96 );
nand NAND2_28608 ( P3_R1054_U166 , P3_U3424 , P3_R1054_U49 );
nand NAND2_28609 ( P3_R1054_U167 , P3_R1054_U166 , P3_R1054_U96 );
nand NAND2_28610 ( P3_R1054_U168 , P3_U3570 , P3_R1054_U48 );
not NOT1_28611 ( P3_R1054_U169 , P3_R1054_U95 );
nand NAND2_28612 ( P3_R1054_U170 , P3_U3427 , P3_R1054_U51 );
nand NAND2_28613 ( P3_R1054_U171 , P3_R1054_U170 , P3_R1054_U95 );
nand NAND2_28614 ( P3_R1054_U172 , P3_U3569 , P3_R1054_U50 );
not NOT1_28615 ( P3_R1054_U173 , P3_R1054_U94 );
nand NAND2_28616 ( P3_R1054_U174 , P3_U3436 , P3_R1054_U55 );
nand NAND2_28617 ( P3_R1054_U175 , P3_U3566 , P3_R1054_U52 );
nand NAND2_28618 ( P3_R1054_U176 , P3_U3567 , P3_R1054_U53 );
nand NAND2_28619 ( P3_R1054_U177 , P3_R1054_U104 , P3_R1054_U10 );
nand NAND2_28620 ( P3_R1054_U178 , P3_R1054_U11 , P3_R1054_U177 );
nand NAND2_28621 ( P3_R1054_U179 , P3_U3430 , P3_R1054_U57 );
nand NAND2_28622 ( P3_R1054_U180 , P3_U3436 , P3_R1054_U55 );
nand NAND3_28623 ( P3_R1054_U181 , P3_R1054_U179 , P3_R1054_U10 , P3_R1054_U94 );
nand NAND2_28624 ( P3_R1054_U182 , P3_R1054_U180 , P3_R1054_U178 );
not NOT1_28625 ( P3_R1054_U183 , P3_R1054_U93 );
nand NAND2_28626 ( P3_R1054_U184 , P3_U3439 , P3_R1054_U60 );
nand NAND2_28627 ( P3_R1054_U185 , P3_R1054_U184 , P3_R1054_U93 );
nand NAND2_28628 ( P3_R1054_U186 , P3_U3565 , P3_R1054_U59 );
not NOT1_28629 ( P3_R1054_U187 , P3_R1054_U61 );
nand NAND2_28630 ( P3_R1054_U188 , P3_R1054_U187 , P3_R1054_U62 );
nand NAND2_28631 ( P3_R1054_U189 , P3_R1054_U188 , P3_R1054_U92 );
nand NAND2_28632 ( P3_R1054_U190 , P3_U3564 , P3_R1054_U61 );
not NOT1_28633 ( P3_R1054_U191 , P3_R1054_U91 );
nand NAND2_28634 ( P3_R1054_U192 , P3_R1054_U179 , P3_R1054_U94 );
not NOT1_28635 ( P3_R1054_U193 , P3_R1054_U63 );
nand NAND2_28636 ( P3_R1054_U194 , P3_U3567 , P3_R1054_U53 );
nand NAND2_28637 ( P3_R1054_U195 , P3_R1054_U193 , P3_R1054_U194 );
nand NAND3_28638 ( P3_R1054_U196 , P3_R1054_U269 , P3_R1054_U100 , P3_R1054_U195 );
nand NAND2_28639 ( P3_R1054_U197 , P3_R1054_U63 , P3_R1054_U100 );
nand NAND2_28640 ( P3_R1054_U198 , P3_U3436 , P3_R1054_U55 );
nand NAND3_28641 ( P3_R1054_U199 , P3_R1054_U198 , P3_R1054_U11 , P3_R1054_U197 );
nand NAND2_28642 ( P3_R1054_U200 , P3_U3567 , P3_R1054_U53 );
nand NAND2_28643 ( P3_R1054_U201 , P3_R1054_U100 , P3_R1054_U200 );
nand NAND2_28644 ( P3_R1054_U202 , P3_R1054_U179 , P3_R1054_U58 );
nand NAND2_28645 ( P3_R1054_U203 , P3_R1054_U134 , P3_R1054_U86 );
not NOT1_28646 ( P3_R1054_U204 , P3_R1054_U64 );
nand NAND2_28647 ( P3_R1054_U205 , P3_U3572 , P3_R1054_U44 );
nand NAND2_28648 ( P3_R1054_U206 , P3_R1054_U204 , P3_R1054_U205 );
nand NAND3_28649 ( P3_R1054_U207 , P3_R1054_U290 , P3_R1054_U99 , P3_R1054_U206 );
nand NAND2_28650 ( P3_R1054_U208 , P3_R1054_U64 , P3_R1054_U99 );
nand NAND2_28651 ( P3_R1054_U209 , P3_U3421 , P3_R1054_U45 );
nand NAND3_28652 ( P3_R1054_U210 , P3_R1054_U209 , P3_R1054_U9 , P3_R1054_U208 );
nand NAND2_28653 ( P3_R1054_U211 , P3_U3572 , P3_R1054_U44 );
nand NAND2_28654 ( P3_R1054_U212 , P3_R1054_U99 , P3_R1054_U211 );
nand NAND2_28655 ( P3_R1054_U213 , P3_U3574 , P3_R1054_U20 );
nand NAND2_28656 ( P3_R1054_U214 , P3_U3415 , P3_R1054_U39 );
nand NAND2_28657 ( P3_R1054_U215 , P3_U3555 , P3_R1054_U38 );
nand NAND2_28658 ( P3_R1054_U216 , P3_R1054_U135 , P3_R1054_U86 );
nand NAND3_28659 ( P3_R1054_U217 , P3_R1054_U215 , P3_R1054_U214 , P3_R1054_U133 );
nand NAND2_28660 ( P3_R1054_U218 , P3_U3412 , P3_R1054_U37 );
nand NAND2_28661 ( P3_R1054_U219 , P3_U3556 , P3_R1054_U34 );
nand NAND2_28662 ( P3_R1054_U220 , P3_U3412 , P3_R1054_U37 );
nand NAND2_28663 ( P3_R1054_U221 , P3_U3556 , P3_R1054_U34 );
nand NAND2_28664 ( P3_R1054_U222 , P3_R1054_U221 , P3_R1054_U220 );
nand NAND2_28665 ( P3_R1054_U223 , P3_U3409 , P3_R1054_U35 );
nand NAND2_28666 ( P3_R1054_U224 , P3_U3557 , P3_R1054_U18 );
nand NAND2_28667 ( P3_R1054_U225 , P3_R1054_U140 , P3_R1054_U40 );
nand NAND3_28668 ( P3_R1054_U226 , P3_R1054_U224 , P3_R1054_U223 , P3_R1054_U127 );
nand NAND2_28669 ( P3_R1054_U227 , P3_U3406 , P3_R1054_U30 );
nand NAND2_28670 ( P3_R1054_U228 , P3_U3558 , P3_R1054_U27 );
nand NAND2_28671 ( P3_R1054_U229 , P3_R1054_U228 , P3_R1054_U227 );
nand NAND2_28672 ( P3_R1054_U230 , P3_U3403 , P3_R1054_U31 );
nand NAND2_28673 ( P3_R1054_U231 , P3_U3559 , P3_R1054_U28 );
nand NAND2_28674 ( P3_R1054_U232 , P3_R1054_U150 , P3_R1054_U41 );
nand NAND3_28675 ( P3_R1054_U233 , P3_R1054_U231 , P3_R1054_U230 , P3_R1054_U142 );
nand NAND2_28676 ( P3_R1054_U234 , P3_U3400 , P3_R1054_U32 );
nand NAND2_28677 ( P3_R1054_U235 , P3_U3560 , P3_R1054_U29 );
nand NAND2_28678 ( P3_R1054_U236 , P3_R1054_U151 , P3_R1054_U87 );
nand NAND3_28679 ( P3_R1054_U237 , P3_R1054_U235 , P3_R1054_U234 , P3_R1054_U117 );
nand NAND2_28680 ( P3_R1054_U238 , P3_U3397 , P3_R1054_U26 );
nand NAND2_28681 ( P3_R1054_U239 , P3_U3561 , P3_R1054_U23 );
nand NAND2_28682 ( P3_R1054_U240 , P3_U3397 , P3_R1054_U26 );
nand NAND2_28683 ( P3_R1054_U241 , P3_U3561 , P3_R1054_U23 );
nand NAND2_28684 ( P3_R1054_U242 , P3_R1054_U241 , P3_R1054_U240 );
nand NAND2_28685 ( P3_R1054_U243 , P3_U3394 , P3_R1054_U24 );
nand NAND2_28686 ( P3_R1054_U244 , P3_U3562 , P3_R1054_U19 );
nand NAND2_28687 ( P3_R1054_U245 , P3_R1054_U156 , P3_R1054_U42 );
nand NAND3_28688 ( P3_R1054_U246 , P3_R1054_U244 , P3_R1054_U243 , P3_R1054_U111 );
nand NAND2_28689 ( P3_R1054_U247 , P3_U3391 , P3_R1054_U22 );
nand NAND2_28690 ( P3_R1054_U248 , P3_U3573 , P3_R1054_U88 );
not NOT1_28691 ( P3_R1054_U249 , P3_R1054_U80 );
nand NAND2_28692 ( P3_R1054_U250 , P3_R1054_U249 , P3_R1054_U107 );
nand NAND2_28693 ( P3_R1054_U251 , P3_R1054_U80 , P3_R1054_U21 );
nand NAND2_28694 ( P3_R1054_U252 , P3_U3379 , P3_R1054_U90 );
nand NAND2_28695 ( P3_R1054_U253 , P3_U3563 , P3_R1054_U89 );
not NOT1_28696 ( P3_R1054_U254 , P3_R1054_U81 );
nand NAND2_28697 ( P3_R1054_U255 , P3_R1054_U191 , P3_R1054_U254 );
nand NAND2_28698 ( P3_R1054_U256 , P3_R1054_U81 , P3_R1054_U91 );
nand NAND2_28699 ( P3_R1054_U257 , P3_U3442 , P3_R1054_U62 );
nand NAND2_28700 ( P3_R1054_U258 , P3_U3564 , P3_R1054_U92 );
not NOT1_28701 ( P3_R1054_U259 , P3_R1054_U82 );
nand NAND2_28702 ( P3_R1054_U260 , P3_R1054_U259 , P3_R1054_U187 );
nand NAND2_28703 ( P3_R1054_U261 , P3_R1054_U82 , P3_R1054_U61 );
nand NAND2_28704 ( P3_R1054_U262 , P3_U3439 , P3_R1054_U60 );
nand NAND2_28705 ( P3_R1054_U263 , P3_U3565 , P3_R1054_U59 );
not NOT1_28706 ( P3_R1054_U264 , P3_R1054_U83 );
nand NAND2_28707 ( P3_R1054_U265 , P3_R1054_U183 , P3_R1054_U264 );
nand NAND2_28708 ( P3_R1054_U266 , P3_R1054_U83 , P3_R1054_U93 );
nand NAND2_28709 ( P3_R1054_U267 , P3_U3436 , P3_R1054_U55 );
nand NAND2_28710 ( P3_R1054_U268 , P3_U3566 , P3_R1054_U52 );
nand NAND2_28711 ( P3_R1054_U269 , P3_R1054_U268 , P3_R1054_U267 );
nand NAND2_28712 ( P3_R1054_U270 , P3_U3433 , P3_R1054_U56 );
nand NAND2_28713 ( P3_R1054_U271 , P3_U3567 , P3_R1054_U53 );
nand NAND2_28714 ( P3_R1054_U272 , P3_R1054_U201 , P3_R1054_U63 );
nand NAND3_28715 ( P3_R1054_U273 , P3_R1054_U271 , P3_R1054_U270 , P3_R1054_U193 );
nand NAND2_28716 ( P3_R1054_U274 , P3_U3430 , P3_R1054_U57 );
nand NAND2_28717 ( P3_R1054_U275 , P3_U3568 , P3_R1054_U54 );
nand NAND2_28718 ( P3_R1054_U276 , P3_R1054_U202 , P3_R1054_U94 );
nand NAND3_28719 ( P3_R1054_U277 , P3_R1054_U275 , P3_R1054_U274 , P3_R1054_U173 );
nand NAND2_28720 ( P3_R1054_U278 , P3_U3427 , P3_R1054_U51 );
nand NAND2_28721 ( P3_R1054_U279 , P3_U3569 , P3_R1054_U50 );
not NOT1_28722 ( P3_R1054_U280 , P3_R1054_U84 );
nand NAND2_28723 ( P3_R1054_U281 , P3_R1054_U169 , P3_R1054_U280 );
nand NAND2_28724 ( P3_R1054_U282 , P3_R1054_U84 , P3_R1054_U95 );
nand NAND2_28725 ( P3_R1054_U283 , P3_U3424 , P3_R1054_U49 );
nand NAND2_28726 ( P3_R1054_U284 , P3_U3570 , P3_R1054_U48 );
not NOT1_28727 ( P3_R1054_U285 , P3_R1054_U85 );
nand NAND2_28728 ( P3_R1054_U286 , P3_R1054_U165 , P3_R1054_U285 );
nand NAND2_28729 ( P3_R1054_U287 , P3_R1054_U85 , P3_R1054_U96 );
nand NAND2_28730 ( P3_R1054_U288 , P3_U3421 , P3_R1054_U45 );
nand NAND2_28731 ( P3_R1054_U289 , P3_U3571 , P3_R1054_U43 );
nand NAND2_28732 ( P3_R1054_U290 , P3_R1054_U289 , P3_R1054_U288 );
nand NAND2_28733 ( P3_R1054_U291 , P3_U3418 , P3_R1054_U46 );
nand NAND2_28734 ( P3_R1054_U292 , P3_U3572 , P3_R1054_U44 );
nand NAND2_28735 ( P3_R1054_U293 , P3_R1054_U212 , P3_R1054_U64 );
nand NAND3_28736 ( P3_R1054_U294 , P3_R1054_U292 , P3_R1054_U291 , P3_R1054_U204 );
and AND2_28737 ( P3_R1161_U4 , P3_R1161_U179 , P3_R1161_U178 );
and AND2_28738 ( P3_R1161_U5 , P3_R1161_U197 , P3_R1161_U196 );
and AND2_28739 ( P3_R1161_U6 , P3_R1161_U237 , P3_R1161_U236 );
and AND2_28740 ( P3_R1161_U7 , P3_R1161_U246 , P3_R1161_U245 );
and AND2_28741 ( P3_R1161_U8 , P3_R1161_U264 , P3_R1161_U263 );
and AND2_28742 ( P3_R1161_U9 , P3_R1161_U272 , P3_R1161_U271 );
and AND2_28743 ( P3_R1161_U10 , P3_R1161_U351 , P3_R1161_U348 );
and AND2_28744 ( P3_R1161_U11 , P3_R1161_U344 , P3_R1161_U341 );
and AND2_28745 ( P3_R1161_U12 , P3_R1161_U335 , P3_R1161_U332 );
and AND2_28746 ( P3_R1161_U13 , P3_R1161_U326 , P3_R1161_U323 );
and AND2_28747 ( P3_R1161_U14 , P3_R1161_U320 , P3_R1161_U318 );
and AND2_28748 ( P3_R1161_U15 , P3_R1161_U313 , P3_R1161_U310 );
and AND2_28749 ( P3_R1161_U16 , P3_R1161_U235 , P3_R1161_U232 );
and AND2_28750 ( P3_R1161_U17 , P3_R1161_U227 , P3_R1161_U224 );
and AND2_28751 ( P3_R1161_U18 , P3_R1161_U213 , P3_R1161_U210 );
not NOT1_28752 ( P3_R1161_U19 , P3_U3407 );
not NOT1_28753 ( P3_R1161_U20 , P3_U3070 );
not NOT1_28754 ( P3_R1161_U21 , P3_U3069 );
nand NAND2_28755 ( P3_R1161_U22 , P3_U3070 , P3_U3407 );
not NOT1_28756 ( P3_R1161_U23 , P3_U3410 );
not NOT1_28757 ( P3_R1161_U24 , P3_U3401 );
not NOT1_28758 ( P3_R1161_U25 , P3_U3059 );
not NOT1_28759 ( P3_R1161_U26 , P3_U3066 );
not NOT1_28760 ( P3_R1161_U27 , P3_U3395 );
not NOT1_28761 ( P3_R1161_U28 , P3_U3067 );
not NOT1_28762 ( P3_R1161_U29 , P3_U3387 );
not NOT1_28763 ( P3_R1161_U30 , P3_U3076 );
nand NAND2_28764 ( P3_R1161_U31 , P3_U3076 , P3_U3387 );
not NOT1_28765 ( P3_R1161_U32 , P3_U3398 );
not NOT1_28766 ( P3_R1161_U33 , P3_U3063 );
nand NAND2_28767 ( P3_R1161_U34 , P3_U3059 , P3_U3401 );
not NOT1_28768 ( P3_R1161_U35 , P3_U3404 );
not NOT1_28769 ( P3_R1161_U36 , P3_U3413 );
not NOT1_28770 ( P3_R1161_U37 , P3_U3083 );
not NOT1_28771 ( P3_R1161_U38 , P3_U3082 );
not NOT1_28772 ( P3_R1161_U39 , P3_U3416 );
nand NAND2_28773 ( P3_R1161_U40 , P3_R1161_U63 , P3_R1161_U205 );
nand NAND2_28774 ( P3_R1161_U41 , P3_R1161_U117 , P3_R1161_U193 );
nand NAND2_28775 ( P3_R1161_U42 , P3_R1161_U182 , P3_R1161_U183 );
nand NAND2_28776 ( P3_R1161_U43 , P3_U3392 , P3_U3077 );
nand NAND2_28777 ( P3_R1161_U44 , P3_R1161_U122 , P3_R1161_U219 );
nand NAND2_28778 ( P3_R1161_U45 , P3_R1161_U216 , P3_R1161_U215 );
not NOT1_28779 ( P3_R1161_U46 , P3_U3900 );
not NOT1_28780 ( P3_R1161_U47 , P3_U3052 );
not NOT1_28781 ( P3_R1161_U48 , P3_U3056 );
not NOT1_28782 ( P3_R1161_U49 , P3_U3901 );
not NOT1_28783 ( P3_R1161_U50 , P3_U3902 );
not NOT1_28784 ( P3_R1161_U51 , P3_U3057 );
not NOT1_28785 ( P3_R1161_U52 , P3_U3903 );
not NOT1_28786 ( P3_R1161_U53 , P3_U3064 );
not NOT1_28787 ( P3_R1161_U54 , P3_U3906 );
not NOT1_28788 ( P3_R1161_U55 , P3_U3074 );
not NOT1_28789 ( P3_R1161_U56 , P3_U3437 );
not NOT1_28790 ( P3_R1161_U57 , P3_U3072 );
not NOT1_28791 ( P3_R1161_U58 , P3_U3068 );
nand NAND2_28792 ( P3_R1161_U59 , P3_U3072 , P3_U3437 );
not NOT1_28793 ( P3_R1161_U60 , P3_U3440 );
not NOT1_28794 ( P3_R1161_U61 , P3_U3419 );
not NOT1_28795 ( P3_R1161_U62 , P3_U3061 );
nand NAND2_28796 ( P3_R1161_U63 , P3_U3083 , P3_U3413 );
not NOT1_28797 ( P3_R1161_U64 , P3_U3425 );
not NOT1_28798 ( P3_R1161_U65 , P3_U3071 );
not NOT1_28799 ( P3_R1161_U66 , P3_U3422 );
not NOT1_28800 ( P3_R1161_U67 , P3_U3062 );
nand NAND2_28801 ( P3_R1161_U68 , P3_U3062 , P3_U3422 );
not NOT1_28802 ( P3_R1161_U69 , P3_U3428 );
not NOT1_28803 ( P3_R1161_U70 , P3_U3079 );
not NOT1_28804 ( P3_R1161_U71 , P3_U3431 );
not NOT1_28805 ( P3_R1161_U72 , P3_U3078 );
not NOT1_28806 ( P3_R1161_U73 , P3_U3434 );
not NOT1_28807 ( P3_R1161_U74 , P3_U3073 );
not NOT1_28808 ( P3_R1161_U75 , P3_U3443 );
not NOT1_28809 ( P3_R1161_U76 , P3_U3081 );
nand NAND2_28810 ( P3_R1161_U77 , P3_U3081 , P3_U3443 );
not NOT1_28811 ( P3_R1161_U78 , P3_U3445 );
not NOT1_28812 ( P3_R1161_U79 , P3_U3080 );
nand NAND2_28813 ( P3_R1161_U80 , P3_U3080 , P3_U3445 );
not NOT1_28814 ( P3_R1161_U81 , P3_U3907 );
not NOT1_28815 ( P3_R1161_U82 , P3_U3905 );
not NOT1_28816 ( P3_R1161_U83 , P3_U3060 );
not NOT1_28817 ( P3_R1161_U84 , P3_U3904 );
not NOT1_28818 ( P3_R1161_U85 , P3_U3065 );
nand NAND2_28819 ( P3_R1161_U86 , P3_U3901 , P3_U3056 );
not NOT1_28820 ( P3_R1161_U87 , P3_U3053 );
not NOT1_28821 ( P3_R1161_U88 , P3_U3899 );
nand NAND2_28822 ( P3_R1161_U89 , P3_R1161_U306 , P3_R1161_U176 );
not NOT1_28823 ( P3_R1161_U90 , P3_U3075 );
nand NAND2_28824 ( P3_R1161_U91 , P3_R1161_U77 , P3_R1161_U315 );
nand NAND2_28825 ( P3_R1161_U92 , P3_R1161_U261 , P3_R1161_U260 );
nand NAND2_28826 ( P3_R1161_U93 , P3_R1161_U68 , P3_R1161_U337 );
nand NAND2_28827 ( P3_R1161_U94 , P3_R1161_U457 , P3_R1161_U456 );
nand NAND2_28828 ( P3_R1161_U95 , P3_R1161_U504 , P3_R1161_U503 );
nand NAND2_28829 ( P3_R1161_U96 , P3_R1161_U375 , P3_R1161_U374 );
nand NAND2_28830 ( P3_R1161_U97 , P3_R1161_U380 , P3_R1161_U379 );
nand NAND2_28831 ( P3_R1161_U98 , P3_R1161_U387 , P3_R1161_U386 );
nand NAND2_28832 ( P3_R1161_U99 , P3_R1161_U394 , P3_R1161_U393 );
nand NAND2_28833 ( P3_R1161_U100 , P3_R1161_U399 , P3_R1161_U398 );
nand NAND2_28834 ( P3_R1161_U101 , P3_R1161_U408 , P3_R1161_U407 );
nand NAND2_28835 ( P3_R1161_U102 , P3_R1161_U415 , P3_R1161_U414 );
nand NAND2_28836 ( P3_R1161_U103 , P3_R1161_U422 , P3_R1161_U421 );
nand NAND2_28837 ( P3_R1161_U104 , P3_R1161_U429 , P3_R1161_U428 );
nand NAND2_28838 ( P3_R1161_U105 , P3_R1161_U434 , P3_R1161_U433 );
nand NAND2_28839 ( P3_R1161_U106 , P3_R1161_U441 , P3_R1161_U440 );
nand NAND2_28840 ( P3_R1161_U107 , P3_R1161_U448 , P3_R1161_U447 );
nand NAND2_28841 ( P3_R1161_U108 , P3_R1161_U462 , P3_R1161_U461 );
nand NAND2_28842 ( P3_R1161_U109 , P3_R1161_U467 , P3_R1161_U466 );
nand NAND2_28843 ( P3_R1161_U110 , P3_R1161_U474 , P3_R1161_U473 );
nand NAND2_28844 ( P3_R1161_U111 , P3_R1161_U481 , P3_R1161_U480 );
nand NAND2_28845 ( P3_R1161_U112 , P3_R1161_U488 , P3_R1161_U487 );
nand NAND2_28846 ( P3_R1161_U113 , P3_R1161_U495 , P3_R1161_U494 );
nand NAND2_28847 ( P3_R1161_U114 , P3_R1161_U500 , P3_R1161_U499 );
and AND2_28848 ( P3_R1161_U115 , P3_R1161_U189 , P3_R1161_U187 );
and AND2_28849 ( P3_R1161_U116 , P3_R1161_U4 , P3_R1161_U180 );
and AND2_28850 ( P3_R1161_U117 , P3_R1161_U194 , P3_R1161_U192 );
and AND2_28851 ( P3_R1161_U118 , P3_R1161_U201 , P3_R1161_U200 );
and AND3_28852 ( P3_R1161_U119 , P3_R1161_U382 , P3_R1161_U381 , P3_R1161_U22 );
and AND2_28853 ( P3_R1161_U120 , P3_R1161_U212 , P3_R1161_U5 );
and AND2_28854 ( P3_R1161_U121 , P3_R1161_U181 , P3_R1161_U180 );
and AND2_28855 ( P3_R1161_U122 , P3_R1161_U220 , P3_R1161_U218 );
and AND3_28856 ( P3_R1161_U123 , P3_R1161_U389 , P3_R1161_U388 , P3_R1161_U34 );
and AND2_28857 ( P3_R1161_U124 , P3_R1161_U226 , P3_R1161_U4 );
and AND2_28858 ( P3_R1161_U125 , P3_R1161_U234 , P3_R1161_U181 );
and AND2_28859 ( P3_R1161_U126 , P3_R1161_U204 , P3_R1161_U6 );
and AND2_28860 ( P3_R1161_U127 , P3_R1161_U243 , P3_R1161_U239 );
and AND2_28861 ( P3_R1161_U128 , P3_R1161_U250 , P3_R1161_U7 );
and AND2_28862 ( P3_R1161_U129 , P3_R1161_U248 , P3_R1161_U172 );
and AND2_28863 ( P3_R1161_U130 , P3_R1161_U268 , P3_R1161_U267 );
and AND3_28864 ( P3_R1161_U131 , P3_R1161_U9 , P3_R1161_U282 , P3_R1161_U273 );
and AND2_28865 ( P3_R1161_U132 , P3_R1161_U285 , P3_R1161_U280 );
and AND2_28866 ( P3_R1161_U133 , P3_R1161_U301 , P3_R1161_U298 );
and AND2_28867 ( P3_R1161_U134 , P3_R1161_U368 , P3_R1161_U302 );
and AND2_28868 ( P3_R1161_U135 , P3_R1161_U160 , P3_R1161_U278 );
and AND3_28869 ( P3_R1161_U136 , P3_R1161_U455 , P3_R1161_U454 , P3_R1161_U80 );
and AND2_28870 ( P3_R1161_U137 , P3_R1161_U325 , P3_R1161_U9 );
and AND3_28871 ( P3_R1161_U138 , P3_R1161_U469 , P3_R1161_U468 , P3_R1161_U59 );
and AND2_28872 ( P3_R1161_U139 , P3_R1161_U334 , P3_R1161_U8 );
and AND3_28873 ( P3_R1161_U140 , P3_R1161_U490 , P3_R1161_U489 , P3_R1161_U172 );
and AND2_28874 ( P3_R1161_U141 , P3_R1161_U343 , P3_R1161_U7 );
and AND3_28875 ( P3_R1161_U142 , P3_R1161_U502 , P3_R1161_U501 , P3_R1161_U171 );
and AND2_28876 ( P3_R1161_U143 , P3_R1161_U350 , P3_R1161_U6 );
nand NAND2_28877 ( P3_R1161_U144 , P3_R1161_U118 , P3_R1161_U202 );
nand NAND2_28878 ( P3_R1161_U145 , P3_R1161_U217 , P3_R1161_U229 );
not NOT1_28879 ( P3_R1161_U146 , P3_U3054 );
not NOT1_28880 ( P3_R1161_U147 , P3_U3908 );
and AND2_28881 ( P3_R1161_U148 , P3_R1161_U403 , P3_R1161_U402 );
nand NAND3_28882 ( P3_R1161_U149 , P3_R1161_U304 , P3_R1161_U169 , P3_R1161_U364 );
and AND2_28883 ( P3_R1161_U150 , P3_R1161_U410 , P3_R1161_U409 );
nand NAND3_28884 ( P3_R1161_U151 , P3_R1161_U370 , P3_R1161_U369 , P3_R1161_U134 );
and AND2_28885 ( P3_R1161_U152 , P3_R1161_U417 , P3_R1161_U416 );
nand NAND3_28886 ( P3_R1161_U153 , P3_R1161_U365 , P3_R1161_U299 , P3_R1161_U86 );
and AND2_28887 ( P3_R1161_U154 , P3_R1161_U424 , P3_R1161_U423 );
nand NAND2_28888 ( P3_R1161_U155 , P3_R1161_U293 , P3_R1161_U292 );
and AND2_28889 ( P3_R1161_U156 , P3_R1161_U436 , P3_R1161_U435 );
nand NAND2_28890 ( P3_R1161_U157 , P3_R1161_U289 , P3_R1161_U288 );
and AND2_28891 ( P3_R1161_U158 , P3_R1161_U443 , P3_R1161_U442 );
nand NAND2_28892 ( P3_R1161_U159 , P3_R1161_U132 , P3_R1161_U284 );
and AND2_28893 ( P3_R1161_U160 , P3_R1161_U450 , P3_R1161_U449 );
nand NAND2_28894 ( P3_R1161_U161 , P3_R1161_U43 , P3_R1161_U327 );
nand NAND2_28895 ( P3_R1161_U162 , P3_R1161_U130 , P3_R1161_U269 );
and AND2_28896 ( P3_R1161_U163 , P3_R1161_U476 , P3_R1161_U475 );
nand NAND2_28897 ( P3_R1161_U164 , P3_R1161_U257 , P3_R1161_U256 );
and AND2_28898 ( P3_R1161_U165 , P3_R1161_U483 , P3_R1161_U482 );
nand NAND2_28899 ( P3_R1161_U166 , P3_R1161_U253 , P3_R1161_U252 );
nand NAND2_28900 ( P3_R1161_U167 , P3_R1161_U127 , P3_R1161_U242 );
nand NAND2_28901 ( P3_R1161_U168 , P3_R1161_U367 , P3_R1161_U366 );
nand NAND2_28902 ( P3_R1161_U169 , P3_U3053 , P3_R1161_U151 );
not NOT1_28903 ( P3_R1161_U170 , P3_R1161_U34 );
nand NAND2_28904 ( P3_R1161_U171 , P3_U3416 , P3_U3082 );
nand NAND2_28905 ( P3_R1161_U172 , P3_U3071 , P3_U3425 );
nand NAND2_28906 ( P3_R1161_U173 , P3_U3057 , P3_U3902 );
not NOT1_28907 ( P3_R1161_U174 , P3_R1161_U68 );
not NOT1_28908 ( P3_R1161_U175 , P3_R1161_U77 );
nand NAND2_28909 ( P3_R1161_U176 , P3_U3064 , P3_U3903 );
not NOT1_28910 ( P3_R1161_U177 , P3_R1161_U63 );
or OR2_28911 ( P3_R1161_U178 , P3_U3066 , P3_U3404 );
or OR2_28912 ( P3_R1161_U179 , P3_U3059 , P3_U3401 );
or OR2_28913 ( P3_R1161_U180 , P3_U3398 , P3_U3063 );
or OR2_28914 ( P3_R1161_U181 , P3_U3395 , P3_U3067 );
not NOT1_28915 ( P3_R1161_U182 , P3_R1161_U31 );
or OR2_28916 ( P3_R1161_U183 , P3_U3392 , P3_U3077 );
not NOT1_28917 ( P3_R1161_U184 , P3_R1161_U42 );
not NOT1_28918 ( P3_R1161_U185 , P3_R1161_U43 );
nand NAND2_28919 ( P3_R1161_U186 , P3_R1161_U42 , P3_R1161_U43 );
nand NAND2_28920 ( P3_R1161_U187 , P3_U3067 , P3_U3395 );
nand NAND2_28921 ( P3_R1161_U188 , P3_R1161_U186 , P3_R1161_U181 );
nand NAND2_28922 ( P3_R1161_U189 , P3_U3063 , P3_U3398 );
nand NAND2_28923 ( P3_R1161_U190 , P3_R1161_U115 , P3_R1161_U188 );
nand NAND2_28924 ( P3_R1161_U191 , P3_R1161_U35 , P3_R1161_U34 );
nand NAND2_28925 ( P3_R1161_U192 , P3_U3066 , P3_R1161_U191 );
nand NAND2_28926 ( P3_R1161_U193 , P3_R1161_U116 , P3_R1161_U190 );
nand NAND2_28927 ( P3_R1161_U194 , P3_U3404 , P3_R1161_U170 );
not NOT1_28928 ( P3_R1161_U195 , P3_R1161_U41 );
or OR2_28929 ( P3_R1161_U196 , P3_U3069 , P3_U3410 );
or OR2_28930 ( P3_R1161_U197 , P3_U3070 , P3_U3407 );
not NOT1_28931 ( P3_R1161_U198 , P3_R1161_U22 );
nand NAND2_28932 ( P3_R1161_U199 , P3_R1161_U23 , P3_R1161_U22 );
nand NAND2_28933 ( P3_R1161_U200 , P3_U3069 , P3_R1161_U199 );
nand NAND2_28934 ( P3_R1161_U201 , P3_U3410 , P3_R1161_U198 );
nand NAND2_28935 ( P3_R1161_U202 , P3_R1161_U5 , P3_R1161_U41 );
not NOT1_28936 ( P3_R1161_U203 , P3_R1161_U144 );
or OR2_28937 ( P3_R1161_U204 , P3_U3413 , P3_U3083 );
nand NAND2_28938 ( P3_R1161_U205 , P3_R1161_U204 , P3_R1161_U144 );
not NOT1_28939 ( P3_R1161_U206 , P3_R1161_U40 );
or OR2_28940 ( P3_R1161_U207 , P3_U3082 , P3_U3416 );
or OR2_28941 ( P3_R1161_U208 , P3_U3407 , P3_U3070 );
nand NAND2_28942 ( P3_R1161_U209 , P3_R1161_U208 , P3_R1161_U41 );
nand NAND2_28943 ( P3_R1161_U210 , P3_R1161_U119 , P3_R1161_U209 );
nand NAND2_28944 ( P3_R1161_U211 , P3_R1161_U195 , P3_R1161_U22 );
nand NAND2_28945 ( P3_R1161_U212 , P3_U3410 , P3_U3069 );
nand NAND2_28946 ( P3_R1161_U213 , P3_R1161_U120 , P3_R1161_U211 );
or OR2_28947 ( P3_R1161_U214 , P3_U3070 , P3_U3407 );
nand NAND2_28948 ( P3_R1161_U215 , P3_R1161_U185 , P3_R1161_U181 );
nand NAND2_28949 ( P3_R1161_U216 , P3_U3067 , P3_U3395 );
not NOT1_28950 ( P3_R1161_U217 , P3_R1161_U45 );
nand NAND2_28951 ( P3_R1161_U218 , P3_R1161_U121 , P3_R1161_U184 );
nand NAND2_28952 ( P3_R1161_U219 , P3_R1161_U45 , P3_R1161_U180 );
nand NAND2_28953 ( P3_R1161_U220 , P3_U3063 , P3_U3398 );
not NOT1_28954 ( P3_R1161_U221 , P3_R1161_U44 );
or OR2_28955 ( P3_R1161_U222 , P3_U3401 , P3_U3059 );
nand NAND2_28956 ( P3_R1161_U223 , P3_R1161_U222 , P3_R1161_U44 );
nand NAND2_28957 ( P3_R1161_U224 , P3_R1161_U123 , P3_R1161_U223 );
nand NAND2_28958 ( P3_R1161_U225 , P3_R1161_U221 , P3_R1161_U34 );
nand NAND2_28959 ( P3_R1161_U226 , P3_U3404 , P3_U3066 );
nand NAND2_28960 ( P3_R1161_U227 , P3_R1161_U124 , P3_R1161_U225 );
or OR2_28961 ( P3_R1161_U228 , P3_U3059 , P3_U3401 );
nand NAND2_28962 ( P3_R1161_U229 , P3_R1161_U184 , P3_R1161_U181 );
not NOT1_28963 ( P3_R1161_U230 , P3_R1161_U145 );
nand NAND2_28964 ( P3_R1161_U231 , P3_U3063 , P3_U3398 );
nand NAND4_28965 ( P3_R1161_U232 , P3_R1161_U401 , P3_R1161_U400 , P3_R1161_U43 , P3_R1161_U42 );
nand NAND2_28966 ( P3_R1161_U233 , P3_R1161_U43 , P3_R1161_U42 );
nand NAND2_28967 ( P3_R1161_U234 , P3_U3067 , P3_U3395 );
nand NAND2_28968 ( P3_R1161_U235 , P3_R1161_U125 , P3_R1161_U233 );
or OR2_28969 ( P3_R1161_U236 , P3_U3082 , P3_U3416 );
or OR2_28970 ( P3_R1161_U237 , P3_U3061 , P3_U3419 );
nand NAND2_28971 ( P3_R1161_U238 , P3_R1161_U177 , P3_R1161_U6 );
nand NAND2_28972 ( P3_R1161_U239 , P3_U3061 , P3_U3419 );
nand NAND2_28973 ( P3_R1161_U240 , P3_R1161_U171 , P3_R1161_U238 );
or OR2_28974 ( P3_R1161_U241 , P3_U3419 , P3_U3061 );
nand NAND2_28975 ( P3_R1161_U242 , P3_R1161_U126 , P3_R1161_U144 );
nand NAND2_28976 ( P3_R1161_U243 , P3_R1161_U241 , P3_R1161_U240 );
not NOT1_28977 ( P3_R1161_U244 , P3_R1161_U167 );
or OR2_28978 ( P3_R1161_U245 , P3_U3079 , P3_U3428 );
or OR2_28979 ( P3_R1161_U246 , P3_U3071 , P3_U3425 );
nand NAND2_28980 ( P3_R1161_U247 , P3_R1161_U174 , P3_R1161_U7 );
nand NAND2_28981 ( P3_R1161_U248 , P3_U3079 , P3_U3428 );
nand NAND2_28982 ( P3_R1161_U249 , P3_R1161_U129 , P3_R1161_U247 );
or OR2_28983 ( P3_R1161_U250 , P3_U3422 , P3_U3062 );
or OR2_28984 ( P3_R1161_U251 , P3_U3428 , P3_U3079 );
nand NAND2_28985 ( P3_R1161_U252 , P3_R1161_U128 , P3_R1161_U167 );
nand NAND2_28986 ( P3_R1161_U253 , P3_R1161_U251 , P3_R1161_U249 );
not NOT1_28987 ( P3_R1161_U254 , P3_R1161_U166 );
or OR2_28988 ( P3_R1161_U255 , P3_U3431 , P3_U3078 );
nand NAND2_28989 ( P3_R1161_U256 , P3_R1161_U255 , P3_R1161_U166 );
nand NAND2_28990 ( P3_R1161_U257 , P3_U3078 , P3_U3431 );
not NOT1_28991 ( P3_R1161_U258 , P3_R1161_U164 );
or OR2_28992 ( P3_R1161_U259 , P3_U3434 , P3_U3073 );
nand NAND2_28993 ( P3_R1161_U260 , P3_R1161_U259 , P3_R1161_U164 );
nand NAND2_28994 ( P3_R1161_U261 , P3_U3073 , P3_U3434 );
not NOT1_28995 ( P3_R1161_U262 , P3_R1161_U92 );
or OR2_28996 ( P3_R1161_U263 , P3_U3068 , P3_U3440 );
or OR2_28997 ( P3_R1161_U264 , P3_U3072 , P3_U3437 );
not NOT1_28998 ( P3_R1161_U265 , P3_R1161_U59 );
nand NAND2_28999 ( P3_R1161_U266 , P3_R1161_U60 , P3_R1161_U59 );
nand NAND2_29000 ( P3_R1161_U267 , P3_U3068 , P3_R1161_U266 );
nand NAND2_29001 ( P3_R1161_U268 , P3_U3440 , P3_R1161_U265 );
nand NAND2_29002 ( P3_R1161_U269 , P3_R1161_U8 , P3_R1161_U92 );
not NOT1_29003 ( P3_R1161_U270 , P3_R1161_U162 );
or OR2_29004 ( P3_R1161_U271 , P3_U3075 , P3_U3907 );
or OR2_29005 ( P3_R1161_U272 , P3_U3080 , P3_U3445 );
or OR2_29006 ( P3_R1161_U273 , P3_U3074 , P3_U3906 );
not NOT1_29007 ( P3_R1161_U274 , P3_R1161_U80 );
nand NAND2_29008 ( P3_R1161_U275 , P3_U3907 , P3_R1161_U274 );
nand NAND2_29009 ( P3_R1161_U276 , P3_R1161_U275 , P3_R1161_U90 );
nand NAND2_29010 ( P3_R1161_U277 , P3_R1161_U80 , P3_R1161_U81 );
nand NAND2_29011 ( P3_R1161_U278 , P3_R1161_U277 , P3_R1161_U276 );
nand NAND2_29012 ( P3_R1161_U279 , P3_R1161_U175 , P3_R1161_U9 );
nand NAND2_29013 ( P3_R1161_U280 , P3_U3074 , P3_U3906 );
nand NAND2_29014 ( P3_R1161_U281 , P3_R1161_U278 , P3_R1161_U279 );
or OR2_29015 ( P3_R1161_U282 , P3_U3443 , P3_U3081 );
or OR2_29016 ( P3_R1161_U283 , P3_U3906 , P3_U3074 );
nand NAND2_29017 ( P3_R1161_U284 , P3_R1161_U162 , P3_R1161_U131 );
nand NAND2_29018 ( P3_R1161_U285 , P3_R1161_U283 , P3_R1161_U281 );
not NOT1_29019 ( P3_R1161_U286 , P3_R1161_U159 );
or OR2_29020 ( P3_R1161_U287 , P3_U3905 , P3_U3060 );
nand NAND2_29021 ( P3_R1161_U288 , P3_R1161_U287 , P3_R1161_U159 );
nand NAND2_29022 ( P3_R1161_U289 , P3_U3060 , P3_U3905 );
not NOT1_29023 ( P3_R1161_U290 , P3_R1161_U157 );
or OR2_29024 ( P3_R1161_U291 , P3_U3904 , P3_U3065 );
nand NAND2_29025 ( P3_R1161_U292 , P3_R1161_U291 , P3_R1161_U157 );
nand NAND2_29026 ( P3_R1161_U293 , P3_U3065 , P3_U3904 );
not NOT1_29027 ( P3_R1161_U294 , P3_R1161_U155 );
or OR2_29028 ( P3_R1161_U295 , P3_U3057 , P3_U3902 );
nand NAND2_29029 ( P3_R1161_U296 , P3_R1161_U176 , P3_R1161_U173 );
not NOT1_29030 ( P3_R1161_U297 , P3_R1161_U86 );
or OR2_29031 ( P3_R1161_U298 , P3_U3903 , P3_U3064 );
nand NAND3_29032 ( P3_R1161_U299 , P3_R1161_U155 , P3_R1161_U298 , P3_R1161_U168 );
not NOT1_29033 ( P3_R1161_U300 , P3_R1161_U153 );
or OR2_29034 ( P3_R1161_U301 , P3_U3900 , P3_U3052 );
nand NAND2_29035 ( P3_R1161_U302 , P3_U3052 , P3_U3900 );
not NOT1_29036 ( P3_R1161_U303 , P3_R1161_U151 );
nand NAND2_29037 ( P3_R1161_U304 , P3_U3899 , P3_R1161_U151 );
not NOT1_29038 ( P3_R1161_U305 , P3_R1161_U149 );
nand NAND2_29039 ( P3_R1161_U306 , P3_R1161_U298 , P3_R1161_U155 );
not NOT1_29040 ( P3_R1161_U307 , P3_R1161_U89 );
or OR2_29041 ( P3_R1161_U308 , P3_U3902 , P3_U3057 );
nand NAND2_29042 ( P3_R1161_U309 , P3_R1161_U308 , P3_R1161_U89 );
nand NAND3_29043 ( P3_R1161_U310 , P3_R1161_U309 , P3_R1161_U173 , P3_R1161_U154 );
nand NAND2_29044 ( P3_R1161_U311 , P3_R1161_U307 , P3_R1161_U173 );
nand NAND2_29045 ( P3_R1161_U312 , P3_U3901 , P3_U3056 );
nand NAND3_29046 ( P3_R1161_U313 , P3_R1161_U311 , P3_R1161_U312 , P3_R1161_U168 );
or OR2_29047 ( P3_R1161_U314 , P3_U3057 , P3_U3902 );
nand NAND2_29048 ( P3_R1161_U315 , P3_R1161_U282 , P3_R1161_U162 );
not NOT1_29049 ( P3_R1161_U316 , P3_R1161_U91 );
nand NAND2_29050 ( P3_R1161_U317 , P3_R1161_U9 , P3_R1161_U91 );
nand NAND2_29051 ( P3_R1161_U318 , P3_R1161_U135 , P3_R1161_U317 );
nand NAND2_29052 ( P3_R1161_U319 , P3_R1161_U317 , P3_R1161_U278 );
nand NAND2_29053 ( P3_R1161_U320 , P3_R1161_U453 , P3_R1161_U319 );
or OR2_29054 ( P3_R1161_U321 , P3_U3445 , P3_U3080 );
nand NAND2_29055 ( P3_R1161_U322 , P3_R1161_U321 , P3_R1161_U91 );
nand NAND2_29056 ( P3_R1161_U323 , P3_R1161_U136 , P3_R1161_U322 );
nand NAND2_29057 ( P3_R1161_U324 , P3_R1161_U316 , P3_R1161_U80 );
nand NAND2_29058 ( P3_R1161_U325 , P3_U3075 , P3_U3907 );
nand NAND2_29059 ( P3_R1161_U326 , P3_R1161_U137 , P3_R1161_U324 );
or OR2_29060 ( P3_R1161_U327 , P3_U3392 , P3_U3077 );
not NOT1_29061 ( P3_R1161_U328 , P3_R1161_U161 );
or OR2_29062 ( P3_R1161_U329 , P3_U3080 , P3_U3445 );
or OR2_29063 ( P3_R1161_U330 , P3_U3437 , P3_U3072 );
nand NAND2_29064 ( P3_R1161_U331 , P3_R1161_U330 , P3_R1161_U92 );
nand NAND2_29065 ( P3_R1161_U332 , P3_R1161_U138 , P3_R1161_U331 );
nand NAND2_29066 ( P3_R1161_U333 , P3_R1161_U262 , P3_R1161_U59 );
nand NAND2_29067 ( P3_R1161_U334 , P3_U3440 , P3_U3068 );
nand NAND2_29068 ( P3_R1161_U335 , P3_R1161_U139 , P3_R1161_U333 );
or OR2_29069 ( P3_R1161_U336 , P3_U3072 , P3_U3437 );
nand NAND2_29070 ( P3_R1161_U337 , P3_R1161_U250 , P3_R1161_U167 );
not NOT1_29071 ( P3_R1161_U338 , P3_R1161_U93 );
or OR2_29072 ( P3_R1161_U339 , P3_U3425 , P3_U3071 );
nand NAND2_29073 ( P3_R1161_U340 , P3_R1161_U339 , P3_R1161_U93 );
nand NAND2_29074 ( P3_R1161_U341 , P3_R1161_U140 , P3_R1161_U340 );
nand NAND2_29075 ( P3_R1161_U342 , P3_R1161_U338 , P3_R1161_U172 );
nand NAND2_29076 ( P3_R1161_U343 , P3_U3079 , P3_U3428 );
nand NAND2_29077 ( P3_R1161_U344 , P3_R1161_U141 , P3_R1161_U342 );
or OR2_29078 ( P3_R1161_U345 , P3_U3071 , P3_U3425 );
or OR2_29079 ( P3_R1161_U346 , P3_U3416 , P3_U3082 );
nand NAND2_29080 ( P3_R1161_U347 , P3_R1161_U346 , P3_R1161_U40 );
nand NAND2_29081 ( P3_R1161_U348 , P3_R1161_U142 , P3_R1161_U347 );
nand NAND2_29082 ( P3_R1161_U349 , P3_R1161_U206 , P3_R1161_U171 );
nand NAND2_29083 ( P3_R1161_U350 , P3_U3061 , P3_U3419 );
nand NAND2_29084 ( P3_R1161_U351 , P3_R1161_U143 , P3_R1161_U349 );
nand NAND2_29085 ( P3_R1161_U352 , P3_R1161_U207 , P3_R1161_U171 );
nand NAND2_29086 ( P3_R1161_U353 , P3_R1161_U204 , P3_R1161_U63 );
nand NAND2_29087 ( P3_R1161_U354 , P3_R1161_U214 , P3_R1161_U22 );
nand NAND2_29088 ( P3_R1161_U355 , P3_R1161_U228 , P3_R1161_U34 );
nand NAND2_29089 ( P3_R1161_U356 , P3_R1161_U231 , P3_R1161_U180 );
nand NAND2_29090 ( P3_R1161_U357 , P3_R1161_U314 , P3_R1161_U173 );
nand NAND2_29091 ( P3_R1161_U358 , P3_R1161_U298 , P3_R1161_U176 );
nand NAND2_29092 ( P3_R1161_U359 , P3_R1161_U329 , P3_R1161_U80 );
nand NAND2_29093 ( P3_R1161_U360 , P3_R1161_U282 , P3_R1161_U77 );
nand NAND2_29094 ( P3_R1161_U361 , P3_R1161_U336 , P3_R1161_U59 );
nand NAND2_29095 ( P3_R1161_U362 , P3_R1161_U345 , P3_R1161_U172 );
nand NAND2_29096 ( P3_R1161_U363 , P3_R1161_U250 , P3_R1161_U68 );
nand NAND2_29097 ( P3_R1161_U364 , P3_U3899 , P3_U3053 );
nand NAND2_29098 ( P3_R1161_U365 , P3_R1161_U296 , P3_R1161_U168 );
nand NAND2_29099 ( P3_R1161_U366 , P3_U3056 , P3_R1161_U295 );
nand NAND2_29100 ( P3_R1161_U367 , P3_U3901 , P3_R1161_U295 );
nand NAND3_29101 ( P3_R1161_U368 , P3_R1161_U296 , P3_R1161_U168 , P3_R1161_U301 );
nand NAND3_29102 ( P3_R1161_U369 , P3_R1161_U155 , P3_R1161_U168 , P3_R1161_U133 );
nand NAND2_29103 ( P3_R1161_U370 , P3_R1161_U297 , P3_R1161_U301 );
nand NAND2_29104 ( P3_R1161_U371 , P3_U3082 , P3_R1161_U39 );
nand NAND2_29105 ( P3_R1161_U372 , P3_U3416 , P3_R1161_U38 );
nand NAND2_29106 ( P3_R1161_U373 , P3_R1161_U372 , P3_R1161_U371 );
nand NAND2_29107 ( P3_R1161_U374 , P3_R1161_U352 , P3_R1161_U40 );
nand NAND2_29108 ( P3_R1161_U375 , P3_R1161_U373 , P3_R1161_U206 );
nand NAND2_29109 ( P3_R1161_U376 , P3_U3083 , P3_R1161_U36 );
nand NAND2_29110 ( P3_R1161_U377 , P3_U3413 , P3_R1161_U37 );
nand NAND2_29111 ( P3_R1161_U378 , P3_R1161_U377 , P3_R1161_U376 );
nand NAND2_29112 ( P3_R1161_U379 , P3_R1161_U353 , P3_R1161_U144 );
nand NAND2_29113 ( P3_R1161_U380 , P3_R1161_U203 , P3_R1161_U378 );
nand NAND2_29114 ( P3_R1161_U381 , P3_U3069 , P3_R1161_U23 );
nand NAND2_29115 ( P3_R1161_U382 , P3_U3410 , P3_R1161_U21 );
nand NAND2_29116 ( P3_R1161_U383 , P3_U3070 , P3_R1161_U19 );
nand NAND2_29117 ( P3_R1161_U384 , P3_U3407 , P3_R1161_U20 );
nand NAND2_29118 ( P3_R1161_U385 , P3_R1161_U384 , P3_R1161_U383 );
nand NAND2_29119 ( P3_R1161_U386 , P3_R1161_U354 , P3_R1161_U41 );
nand NAND2_29120 ( P3_R1161_U387 , P3_R1161_U385 , P3_R1161_U195 );
nand NAND2_29121 ( P3_R1161_U388 , P3_U3066 , P3_R1161_U35 );
nand NAND2_29122 ( P3_R1161_U389 , P3_U3404 , P3_R1161_U26 );
nand NAND2_29123 ( P3_R1161_U390 , P3_U3059 , P3_R1161_U24 );
nand NAND2_29124 ( P3_R1161_U391 , P3_U3401 , P3_R1161_U25 );
nand NAND2_29125 ( P3_R1161_U392 , P3_R1161_U391 , P3_R1161_U390 );
nand NAND2_29126 ( P3_R1161_U393 , P3_R1161_U355 , P3_R1161_U44 );
nand NAND2_29127 ( P3_R1161_U394 , P3_R1161_U392 , P3_R1161_U221 );
nand NAND2_29128 ( P3_R1161_U395 , P3_U3063 , P3_R1161_U32 );
nand NAND2_29129 ( P3_R1161_U396 , P3_U3398 , P3_R1161_U33 );
nand NAND2_29130 ( P3_R1161_U397 , P3_R1161_U396 , P3_R1161_U395 );
nand NAND2_29131 ( P3_R1161_U398 , P3_R1161_U356 , P3_R1161_U145 );
nand NAND2_29132 ( P3_R1161_U399 , P3_R1161_U230 , P3_R1161_U397 );
nand NAND2_29133 ( P3_R1161_U400 , P3_U3067 , P3_R1161_U27 );
nand NAND2_29134 ( P3_R1161_U401 , P3_U3395 , P3_R1161_U28 );
nand NAND2_29135 ( P3_R1161_U402 , P3_U3054 , P3_R1161_U147 );
nand NAND2_29136 ( P3_R1161_U403 , P3_U3908 , P3_R1161_U146 );
nand NAND2_29137 ( P3_R1161_U404 , P3_U3054 , P3_R1161_U147 );
nand NAND2_29138 ( P3_R1161_U405 , P3_U3908 , P3_R1161_U146 );
nand NAND2_29139 ( P3_R1161_U406 , P3_R1161_U405 , P3_R1161_U404 );
nand NAND2_29140 ( P3_R1161_U407 , P3_R1161_U148 , P3_R1161_U149 );
nand NAND2_29141 ( P3_R1161_U408 , P3_R1161_U305 , P3_R1161_U406 );
nand NAND2_29142 ( P3_R1161_U409 , P3_U3053 , P3_R1161_U88 );
nand NAND2_29143 ( P3_R1161_U410 , P3_U3899 , P3_R1161_U87 );
nand NAND2_29144 ( P3_R1161_U411 , P3_U3053 , P3_R1161_U88 );
nand NAND2_29145 ( P3_R1161_U412 , P3_U3899 , P3_R1161_U87 );
nand NAND2_29146 ( P3_R1161_U413 , P3_R1161_U412 , P3_R1161_U411 );
nand NAND2_29147 ( P3_R1161_U414 , P3_R1161_U150 , P3_R1161_U151 );
nand NAND2_29148 ( P3_R1161_U415 , P3_R1161_U303 , P3_R1161_U413 );
nand NAND2_29149 ( P3_R1161_U416 , P3_U3052 , P3_R1161_U46 );
nand NAND2_29150 ( P3_R1161_U417 , P3_U3900 , P3_R1161_U47 );
nand NAND2_29151 ( P3_R1161_U418 , P3_U3052 , P3_R1161_U46 );
nand NAND2_29152 ( P3_R1161_U419 , P3_U3900 , P3_R1161_U47 );
nand NAND2_29153 ( P3_R1161_U420 , P3_R1161_U419 , P3_R1161_U418 );
nand NAND2_29154 ( P3_R1161_U421 , P3_R1161_U152 , P3_R1161_U153 );
nand NAND2_29155 ( P3_R1161_U422 , P3_R1161_U300 , P3_R1161_U420 );
nand NAND2_29156 ( P3_R1161_U423 , P3_U3056 , P3_R1161_U49 );
nand NAND2_29157 ( P3_R1161_U424 , P3_U3901 , P3_R1161_U48 );
nand NAND2_29158 ( P3_R1161_U425 , P3_U3057 , P3_R1161_U50 );
nand NAND2_29159 ( P3_R1161_U426 , P3_U3902 , P3_R1161_U51 );
nand NAND2_29160 ( P3_R1161_U427 , P3_R1161_U426 , P3_R1161_U425 );
nand NAND2_29161 ( P3_R1161_U428 , P3_R1161_U357 , P3_R1161_U89 );
nand NAND2_29162 ( P3_R1161_U429 , P3_R1161_U427 , P3_R1161_U307 );

endmodule
