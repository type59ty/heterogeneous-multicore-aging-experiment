`timescale 1ns/10ps

`define cycle 10.0
`define terminate_cycle 400000//200000 // Modify your terminate ycle here

module c5315d_testfixture;

`define in_file "c5315d/rand_input_vector_c5315d_0.out"
`define out_file "c5315d/rand_output_vector_c5315d_0.out"

parameter vec_width = 356;
parameter vec_length = 4;

reg clk = 0;


reg [vec_width-1:0] input_vec_mem [0:vec_length-1];
reg [vec_width-1:0] vec;

wire n1709, n1816, n11066, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11147, n11152, n11153, n11154, n11155, n11972, n12054, n12060, n12061, n12139, n12142, n12309, n12387, n12527, n12584, n12590, n12623, n13357, n13358, n13359, n13360, n13604, n13613, n14272, n14275, n14278, n14279, n14737, n14738, n14739, n14740, n15240, n15388, n16641, n16643, n16646, n16648, n16716, n16877, n16924, n16925, n16926, n16927, n17015, n17363, n17365, n17432, n17449, n17465, n17466, n17467, n17469, n17470, n17471, n17472, n17473, n17474, n17476, n17503, n17504, n17506, n17511, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17626, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n18075, n18076, n18123, n18124, n18127, n18128, n2709, n2816, n21066, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21147, n21152, n21153, n21154, n21155, n21972, n22054, n22060, n22061, n22139, n22142, n22309, n22387, n22527, n22584, n22590, n22623, n23357, n23358, n23359, n23360, n23604, n23613, n24272, n24275, n24278, n24279, n24737, n24738, n24739, n24740, n25240, n25388, n26641, n26643, n26646, n26648, n26716, n26877, n26924, n26925, n26926, n26927, n27015, n27363, n27365, n27432, n27449, n27465, n27466, n27467, n27469, n27470, n27471, n27472, n27473, n27474, n27476, n27503, n27504, n27506, n27511, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27626, n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761, n28075, n28076, n28123, n28124, n28127, n28128;
initial begin
	$readmemb(`in_file, input_vec_mem );
end

always #(`cycle/2) clk = ~clk;

c5315d cc (.N11(vec[355]), .N14(vec[354]), .N111(vec[353]), .N114(vec[352]), .N117(vec[351]), .N120(vec[350]), .N123(vec[349]), .N124(vec[348]), .N125(vec[347]), .N126(vec[346]), .N127(vec[345]), .N131(vec[344]), .N134(vec[343]), .N137(vec[342]), .N140(vec[341]), .N143(vec[340]), .N146(vec[339]), .N149(vec[338]), .N152(vec[337]), .N153(vec[336]), .N154(vec[335]), .N161(vec[334]), .N164(vec[333]), .N167(vec[332]), .N170(vec[331]), .N173(vec[330]), .N176(vec[329]), .N179(vec[328]), .N180(vec[327]), .N181(vec[326]), .N182(vec[325]), .N183(vec[324]), .N186(vec[323]), .N187(vec[322]), .N188(vec[321]), .N191(vec[320]), .N194(vec[319]), .N197(vec[318]), .N1100(vec[317]), .N1103(vec[316]), .N1106(vec[315]), .N1109(vec[314]), .N1112(vec[313]), .N1113(vec[312]), .N1114(vec[311]), .N1115(vec[310]), .N1116(vec[309]), .N1117(vec[308]), .N1118(vec[307]), .N1119(vec[306]), .N1120(vec[305]), .N1121(vec[304]), .N1122(vec[303]), .N1123(vec[302]), .N1126(vec[301]), .N1127(vec[300]), .N1128(vec[299]), .N1129(vec[298]), .N1130(vec[297]), .N1131(vec[296]), .N1132(vec[295]), .N1135(vec[294]), .N1136(vec[293]), .N1137(vec[292]), .N1140(vec[291]), .N1141(vec[290]), .N1145(vec[289]), .N1146(vec[288]), .N1149(vec[287]), .N1152(vec[286]), .N1155(vec[285]), .N1158(vec[284]), .N1161(vec[283]), .N1164(vec[282]), .N1167(vec[281]), .N1170(vec[280]), .N1173(vec[279]), .N1176(vec[278]), .N1179(vec[277]), .N1182(vec[276]), .N1185(vec[275]), .N1188(vec[274]), .N1191(vec[273]), .N1194(vec[272]), .N1197(vec[271]), .N1200(vec[270]), .N1203(vec[269]), .N1206(vec[268]), .N1209(vec[267]), .N1210(vec[266]), .N1217(vec[265]), .N1218(vec[264]), .N1225(vec[263]), .N1226(vec[262]), .N1233(vec[261]), .N1234(vec[260]), .N1241(vec[259]), .N1242(vec[258]), .N1245(vec[257]), .N1248(vec[256]), .N1251(vec[255]), .N1254(vec[254]), .N1257(vec[253]), .N1264(vec[252]), .N1265(vec[251]), .N1272(vec[250]), .N1273(vec[249]), .N1280(vec[248]), .N1281(vec[247]), .N1288(vec[246]), .N1289(vec[245]), .N1292(vec[244]), .N1293(vec[243]), .N1299(vec[242]), .N1302(vec[241]), .N1307(vec[240]), .N1308(vec[239]), .N1315(vec[238]), .N1316(vec[237]), .N1323(vec[236]), .N1324(vec[235]), .N1331(vec[234]), .N1332(vec[233]), .N1335(vec[232]), .N1338(vec[231]), .N1341(vec[230]), .N1348(vec[229]), .N1351(vec[228]), .N1358(vec[227]), .N1361(vec[226]), .N1366(vec[225]), .N1369(vec[224]), .N1372(vec[223]), .N1373(vec[222]), .N1374(vec[221]), .N1386(vec[220]), .N1389(vec[219]), .N1400(vec[218]), .N1411(vec[217]), .N1422(vec[216]), .N1435(vec[215]), .N1446(vec[214]), .N1457(vec[213]), .N1468(vec[212]), .N1479(vec[211]), .N1490(vec[210]), .N1503(vec[209]), .N1514(vec[208]), .N1523(vec[207]), .N1534(vec[206]), .N1545(vec[205]), .N1549(vec[204]), .N1552(vec[203]), .N1556(vec[202]), .N1559(vec[201]), .N1562(vec[200]), .N1566(vec[199]), .N1571(vec[198]), .N1574(vec[197]), .N1577(vec[196]), .N1580(vec[195]), .N1583(vec[194]), .N1588(vec[193]), .N1591(vec[192]), .N1592(vec[191]), .N1595(vec[190]), .N1596(vec[189]), .N1597(vec[188]), .N1598(vec[187]), .N1599(vec[186]), .N1603(vec[185]), .N1607(vec[184]), .N1610(vec[183]), .N1613(vec[182]), .N1616(vec[181]), .N1619(vec[180]), .N1625(vec[179]), .N1631(vec[178]), .N21(vec[177]), .N24(vec[176]), .N211(vec[175]), .N214(vec[174]), .N217(vec[173]), .N220(vec[172]), .N223(vec[171]), .N224(vec[170]), .N225(vec[169]), .N226(vec[168]), .N227(vec[167]), .N231(vec[166]), .N234(vec[165]), .N237(vec[164]), .N240(vec[163]), .N243(vec[162]), .N246(vec[161]), .N249(vec[160]), .N252(vec[159]), .N253(vec[158]), .N254(vec[157]), .N261(vec[156]), .N264(vec[155]), .N267(vec[154]), .N270(vec[153]), .N273(vec[152]), .N276(vec[151]), .N279(vec[150]), .N280(vec[149]), .N281(vec[148]), .N282(vec[147]), .N283(vec[146]), .N286(vec[145]), .N287(vec[144]), .N288(vec[143]), .N291(vec[142]), .N294(vec[141]), .N297(vec[140]), .N2100(vec[139]), .N2103(vec[138]), .N2106(vec[137]), .N2109(vec[136]), .N2112(vec[135]), .N2113(vec[134]), .N2114(vec[133]), .N2115(vec[132]), .N2116(vec[131]), .N2117(vec[130]), .N2118(vec[129]), .N2119(vec[128]), .N2120(vec[127]), .N2121(vec[126]), .N2122(vec[125]), .N2123(vec[124]), .N2126(vec[123]), .N2127(vec[122]), .N2128(vec[121]), .N2129(vec[120]), .N2130(vec[119]), .N2131(vec[118]), .N2132(vec[117]), .N2135(vec[116]), .N2136(vec[115]), .N2137(vec[114]), .N2140(vec[113]), .N2141(vec[112]), .N2145(vec[111]), .N2146(vec[110]), .N2149(vec[109]), .N2152(vec[108]), .N2155(vec[107]), .N2158(vec[106]), .N2161(vec[105]), .N2164(vec[104]), .N2167(vec[103]), .N2170(vec[102]), .N2173(vec[101]), .N2176(vec[100]), .N2179(vec[99]), .N2182(vec[98]), .N2185(vec[97]), .N2188(vec[96]), .N2191(vec[95]), .N2194(vec[94]), .N2197(vec[93]), .N2200(vec[92]), .N2203(vec[91]), .N2206(vec[90]), .N2209(vec[89]), .N2210(vec[88]), .N2217(vec[87]), .N2218(vec[86]), .N2225(vec[85]), .N2226(vec[84]), .N2233(vec[83]), .N2234(vec[82]), .N2241(vec[81]), .N2242(vec[80]), .N2245(vec[79]), .N2248(vec[78]), .N2251(vec[77]), .N2254(vec[76]), .N2257(vec[75]), .N2264(vec[74]), .N2265(vec[73]), .N2272(vec[72]), .N2273(vec[71]), .N2280(vec[70]), .N2281(vec[69]), .N2288(vec[68]), .N2289(vec[67]), .N2292(vec[66]), .N2293(vec[65]), .N2299(vec[64]), .N2302(vec[63]), .N2307(vec[62]), .N2308(vec[61]), .N2315(vec[60]), .N2316(vec[59]), .N2323(vec[58]), .N2324(vec[57]), .N2331(vec[56]), .N2332(vec[55]), .N2335(vec[54]), .N2338(vec[53]), .N2341(vec[52]), .N2348(vec[51]), .N2351(vec[50]), .N2358(vec[49]), .N2361(vec[48]), .N2366(vec[47]), .N2369(vec[46]), .N2372(vec[45]), .N2373(vec[44]), .N2374(vec[43]), .N2386(vec[42]), .N2389(vec[41]), .N2400(vec[40]), .N2411(vec[39]), .N2422(vec[38]), .N2435(vec[37]), .N2446(vec[36]), .N2457(vec[35]), .N2468(vec[34]), .N2479(vec[33]), .N2490(vec[32]), .N2503(vec[31]), .N2514(vec[30]), .N2523(vec[29]), .N2534(vec[28]), .N2545(vec[27]), .N2549(vec[26]), .N2552(vec[25]), .N2556(vec[24]), .N2559(vec[23]), .N2562(vec[22]), .N2566(vec[21]), .N2571(vec[20]), .N2574(vec[19]), .N2577(vec[18]), .N2580(vec[17]), .N2583(vec[16]), .N2588(vec[15]), .N2591(vec[14]), .N2592(vec[13]), .N2595(vec[12]), .N2596(vec[11]), .N2597(vec[10]), .N2598(vec[9]), .N2599(vec[8]), .N2603(vec[7]), .N2607(vec[6]), .N2610(vec[5]), .N2613(vec[4]), .N2616(vec[3]), .N2619(vec[2]), .N2625(vec[1]), .N2631(vec[0]), .N1709(n1709), .N1816(n1816), .N11066(n11066), .N11137(n11137), .N11138(n11138), .N11139(n11139), .N11140(n11140), .N11141(n11141), .N11142(n11142), .N11143(n11143), .N11144(n11144), .N11145(n11145), .N11147(n11147), .N11152(n11152), .N11153(n11153), .N11154(n11154), .N11155(n11155), .N11972(n11972), .N12054(n12054), .N12060(n12060), .N12061(n12061), .N12139(n12139), .N12142(n12142), .N12309(n12309), .N12387(n12387), .N12527(n12527), .N12584(n12584), .N12590(n12590), .N12623(n12623), .N13357(n13357), .N13358(n13358), .N13359(n13359), .N13360(n13360), .N13604(n13604), .N13613(n13613), .N14272(n14272), .N14275(n14275), .N14278(n14278), .N14279(n14279), .N14737(n14737), .N14738(n14738), .N14739(n14739), .N14740(n14740), .N15240(n15240), .N15388(n15388), .N16641(n16641), .N16643(n16643), .N16646(n16646), .N16648(n16648), .N16716(n16716), .N16877(n16877), .N16924(n16924), .N16925(n16925), .N16926(n16926), .N16927(n16927), .N17015(n17015), .N17363(n17363), .N17365(n17365), .N17432(n17432), .N17449(n17449), .N17465(n17465), .N17466(n17466), .N17467(n17467), .N17469(n17469), .N17470(n17470), .N17471(n17471), .N17472(n17472), .N17473(n17473), .N17474(n17474), .N17476(n17476), .N17503(n17503), .N17504(n17504), .N17506(n17506), .N17511(n17511), .N17515(n17515), .N17516(n17516), .N17517(n17517), .N17518(n17518), .N17519(n17519), .N17520(n17520), .N17521(n17521), .N17522(n17522), .N17600(n17600), .N17601(n17601), .N17602(n17602), .N17603(n17603), .N17604(n17604), .N17605(n17605), .N17606(n17606), .N17607(n17607), .N17626(n17626), .N17698(n17698), .N17699(n17699), .N17700(n17700), .N17701(n17701), .N17702(n17702), .N17703(n17703), .N17704(n17704), .N17705(n17705), .N17706(n17706), .N17707(n17707), .N17735(n17735), .N17736(n17736), .N17737(n17737), .N17738(n17738), .N17739(n17739), .N17740(n17740), .N17741(n17741), .N17742(n17742), .N17754(n17754), .N17755(n17755), .N17756(n17756), .N17757(n17757), .N17758(n17758), .N17759(n17759), .N17760(n17760), .N17761(n17761), .N18075(n18075), .N18076(n18076), .N18123(n18123), .N18124(n18124), .N18127(n18127), .N18128(n18128), .N2709(n2709), .N2816(n2816), .N21066(n21066), .N21137(n21137), .N21138(n21138), .N21139(n21139), .N21140(n21140), .N21141(n21141), .N21142(n21142), .N21143(n21143), .N21144(n21144), .N21145(n21145), .N21147(n21147), .N21152(n21152), .N21153(n21153), .N21154(n21154), .N21155(n21155), .N21972(n21972), .N22054(n22054), .N22060(n22060), .N22061(n22061), .N22139(n22139), .N22142(n22142), .N22309(n22309), .N22387(n22387), .N22527(n22527), .N22584(n22584), .N22590(n22590), .N22623(n22623), .N23357(n23357), .N23358(n23358), .N23359(n23359), .N23360(n23360), .N23604(n23604), .N23613(n23613), .N24272(n24272), .N24275(n24275), .N24278(n24278), .N24279(n24279), .N24737(n24737), .N24738(n24738), .N24739(n24739), .N24740(n24740), .N25240(n25240), .N25388(n25388), .N26641(n26641), .N26643(n26643), .N26646(n26646), .N26648(n26648), .N26716(n26716), .N26877(n26877), .N26924(n26924), .N26925(n26925), .N26926(n26926), .N26927(n26927), .N27015(n27015), .N27363(n27363), .N27365(n27365), .N27432(n27432), .N27449(n27449), .N27465(n27465), .N27466(n27466), .N27467(n27467), .N27469(n27469), .N27470(n27470), .N27471(n27471), .N27472(n27472), .N27473(n27473), .N27474(n27474), .N27476(n27476), .N27503(n27503), .N27504(n27504), .N27506(n27506), .N27511(n27511), .N27515(n27515), .N27516(n27516), .N27517(n27517), .N27518(n27518), .N27519(n27519), .N27520(n27520), .N27521(n27521), .N27522(n27522), .N27600(n27600), .N27601(n27601), .N27602(n27602), .N27603(n27603), .N27604(n27604), .N27605(n27605), .N27606(n27606), .N27607(n27607), .N27626(n27626), .N27698(n27698), .N27699(n27699), .N27700(n27700), .N27701(n27701), .N27702(n27702), .N27703(n27703), .N27704(n27704), .N27705(n27705), .N27706(n27706), .N27707(n27707), .N27735(n27735), .N27736(n27736), .N27737(n27737), .N27738(n27738), .N27739(n27739), .N27740(n27740), .N27741(n27741), .N27742(n27742), .N27754(n27754), .N27755(n27755), .N27756(n27756), .N27757(n27757), .N27758(n27758), .N27759(n27759), .N27760(n27760), .N27761(n27761), .N28075(n28075), .N28076(n28076), .N28123(n28123), .N28124(n28124), .N28127(n28127), .N28128(n28128));

integer i=0;
always @ (posedge clk) begin
	vec = input_vec_mem[i];
	$monitor(vec);
	i = i + 1;

end

always @ (negedge clk)begin
	$fdisplay ( fh_w, n1709, n1816, n11066, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11147, n11152, n11153, n11154, n11155, n11972, n12054, n12060, n12061, n12139, n12142, n12309, n12387, n12527, n12584, n12590, n12623, n13357, n13358, n13359, n13360, n13604, n13613, n14272, n14275, n14278, n14279, n14737, n14738, n14739, n14740, n15240, n15388, n16641, n16643, n16646, n16648, n16716, n16877, n16924, n16925, n16926, n16927, n17015, n17363, n17365, n17432, n17449, n17465, n17466, n17467, n17469, n17470, n17471, n17472, n17473, n17474, n17476, n17503, n17504, n17506, n17511, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17626, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n18075, n18076, n18123, n18124, n18127, n18128, n2709, n2816, n21066, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21147, n21152, n21153, n21154, n21155, n21972, n22054, n22060, n22061, n22139, n22142, n22309, n22387, n22527, n22584, n22590, n22623, n23357, n23358, n23359, n23360, n23604, n23613, n24272, n24275, n24278, n24279, n24737, n24738, n24739, n24740, n25240, n25388, n26641, n26643, n26646, n26648, n26716, n26877, n26924, n26925, n26926, n26927, n27015, n27363, n27365, n27432, n27449, n27465, n27466, n27467, n27469, n27470, n27471, n27472, n27473, n27474, n27476, n27503, n27504, n27506, n27511, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27626, n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761, n28075, n28076, n28123, n28124, n28127, n28128);
	if(i == vec_length)begin
		$finish;
	end
end

integer fh_w;
initial begin
	fh_w = $fopen(`out_file, "w");
end
 
initial begin
	//$fsdbDumpfile("SET.fsdb");
	//$fsdbDumpvars;
	//$fsdbDumpMDA;
	$dumpfile("test_result.vcd");
    $dumpvars;

end
endmodule
