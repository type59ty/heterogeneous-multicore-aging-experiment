// b15
// 485 inputs  (36 PIs + 449 PPIs)
// 519 outputs (70 POs + 449 PPOs)
// 8437 gates (7367 gates + 1000 inverters + 70 buffers )
// ( 1232 AND + 54 OR + 6041 NAND + 40 NOR + 70 BUFF )
// Time: Wed Mar 25 17:47:21 2009
// All copyrigh from NCKU EE TestLAB, Taiwan. [2008.12. WCL]

module b15_ras ( U3445 , U3446 , U3447 , U3448 , U3213 , U3212 ,
             U3211 , U3210 , U3209 , U3208 , U3207 , U3206 ,
             U3205 , U3204 , U3203 , U3202 , U3201 , U3200 ,
             U3199 , U3198 , U3197 , U3196 , U3195 , U3194 ,
             U3193 , U3192 , U3191 , U3190 , U3189 , U3188 ,
             U3187 , U3186 , U3185 , U3184 , U3183 , U3182 ,
             U3181 , U3451 , U3452 , U3180 , U3179 , U3178 ,
             U3177 , U3176 , U3175 , U3174 , U3173 , U3172 ,
             U3171 , U3170 , U3169 , U3168 , U3167 , U3166 ,
             U3165 , U3164 , U3163 , U3162 , U3161 , U3160 ,
             U3159 , U3158 , U3157 , U3156 , U3155 , U3154 ,
             U3153 , U3152 , U3151 , U3453 , U3150 , U3149 ,
             U3148 , U3147 , U3146 , U3145 , U3144 , U3143 ,
             U3142 , U3141 , U3140 , U3139 , U3138 , U3137 ,
             U3136 , U3135 , U3134 , U3133 , U3132 , U3131 ,
             U3130 , U3129 , U3128 , U3127 , U3126 , U3125 ,
             U3124 , U3123 , U3122 , U3121 , U3120 , U3119 ,
             U3118 , U3117 , U3116 , U3115 , U3114 , U3113 ,
             U3112 , U3111 , U3110 , U3109 , U3108 , U3107 ,
             U3106 , U3105 , U3104 , U3103 , U3102 , U3101 ,
             U3100 , U3099 , U3098 , U3097 , U3096 , U3095 ,
             U3094 , U3093 , U3092 , U3091 , U3090 , U3089 ,
             U3088 , U3087 , U3086 , U3085 , U3084 , U3083 ,
             U3082 , U3081 , U3080 , U3079 , U3078 , U3077 ,
             U3076 , U3075 , U3074 , U3073 , U3072 , U3071 ,
             U3070 , U3069 , U3068 , U3067 , U3066 , U3065 ,
             U3064 , U3063 , U3062 , U3061 , U3060 , U3059 ,
             U3058 , U3057 , U3056 , U3055 , U3054 , U3053 ,
             U3052 , U3051 , U3050 , U3049 , U3048 , U3047 ,
             U3046 , U3045 , U3044 , U3043 , U3042 , U3041 ,
             U3040 , U3039 , U3038 , U3037 , U3036 , U3035 ,
             U3034 , U3033 , U3032 , U3031 , U3030 , U3029 ,
             U3028 , U3027 , U3026 , U3025 , U3024 , U3023 ,
             U3022 , U3021 , U3020 , U3455 , U3456 , U3459 ,
             U3460 , U3461 , U3019 , U3462 , U3463 , U3464 ,
             U3465 , U3018 , U3017 , U3016 , U3015 , U3014 ,
             U3013 , U3012 , U3011 , U3010 , U3009 , U3008 ,
             U3007 , U3006 , U3005 , U3004 , U3003 , U3002 ,
             U3001 , U3000 , U2999 , U2998 , U2997 , U2996 ,
             U2995 , U2994 , U2993 , U2992 , U2991 , U2990 ,
             U2989 , U2988 , U2987 , U2986 , U2985 , U2984 ,
             U2983 , U2982 , U2981 , U2980 , U2979 , U2978 ,
             U2977 , U2976 , U2975 , U2974 , U2973 , U2972 ,
             U2971 , U2970 , U2969 , U2968 , U2967 , U2966 ,
             U2965 , U2964 , U2963 , U2962 , U2961 , U2960 ,
             U2959 , U2958 , U2957 , U2956 , U2955 , U2954 ,
             U2953 , U2952 , U2951 , U2950 , U2949 , U2948 ,
             U2947 , U2946 , U2945 , U2944 , U2943 , U2942 ,
             U2941 , U2940 , U2939 , U2938 , U2937 , U2936 ,
             U2935 , U2934 , U2933 , U2932 , U2931 , U2930 ,
             U2929 , U2928 , U2927 , U2926 , U2925 , U2924 ,
             U2923 , U2922 , U2921 , U2920 , U2919 , U2918 ,
             U2917 , U2916 , U2915 , U2914 , U2913 , U2912 ,
             U2911 , U2910 , U2909 , U2908 , U2907 , U2906 ,
             U2905 , U2904 , U2903 , U2902 , U2901 , U2900 ,
             U2899 , U2898 , U2897 , U2896 , U2895 , U2894 ,
             U2893 , U2892 , U2891 , U2890 , U2889 , U2888 ,
             U2887 , U2886 , U2885 , U2884 , U2883 , U2882 ,
             U2881 , U2880 , U2879 , U2878 , U2877 , U2876 ,
             U2875 , U2874 , U2873 , U2872 , U2871 , U2870 ,
             U2869 , U2868 , U2867 , U2866 , U2865 , U2864 ,
             U2863 , U2862 , U2861 , U2860 , U2859 , U2858 ,
             U2857 , U2856 , U2855 , U2854 , U2853 , U2852 ,
             U2851 , U2850 , U2849 , U2848 , U2847 , U2846 ,
             U2845 , U2844 , U2843 , U2842 , U2841 , U2840 ,
             U2839 , U2838 , U2837 , U2836 , U2835 , U2834 ,
             U2833 , U2832 , U2831 , U2830 , U2829 , U2828 ,
             U2827 , U2826 , U2825 , U2824 , U2823 , U2822 ,
             U2821 , U2820 , U2819 , U2818 , U2817 , U2816 ,
             U2815 , U2814 , U2813 , U2812 , U2811 , U2810 ,
             U2809 , U2808 , U2807 , U2806 , U2805 , U2804 ,
             U2803 , U2802 , U2801 , U2800 , U2799 , U2798 ,
             U2797 , U2796 , U2795 , U3468 , U2794 , U3469 ,
             U3470 , U2793 , U3471 , U2792 , U3472 , U2791 ,
             U3473 , U2790 , U2789 , U3474 , U2788 , BE_N_REG_3_ ,
             BE_N_REG_2_ , BE_N_REG_1_ , BE_N_REG_0_ , ADDRESS_REG_29_ , ADDRESS_REG_28_ , ADDRESS_REG_27_ ,
             ADDRESS_REG_26_ , ADDRESS_REG_25_ , ADDRESS_REG_24_ , ADDRESS_REG_23_ , ADDRESS_REG_22_ , ADDRESS_REG_21_ ,
             ADDRESS_REG_20_ , ADDRESS_REG_19_ , ADDRESS_REG_18_ , ADDRESS_REG_17_ , ADDRESS_REG_16_ , ADDRESS_REG_15_ ,
             ADDRESS_REG_14_ , ADDRESS_REG_13_ , ADDRESS_REG_12_ , ADDRESS_REG_11_ , ADDRESS_REG_10_ , ADDRESS_REG_9_ ,
             ADDRESS_REG_8_ , ADDRESS_REG_7_ , ADDRESS_REG_6_ , ADDRESS_REG_5_ , ADDRESS_REG_4_ , ADDRESS_REG_3_ ,
             ADDRESS_REG_2_ , ADDRESS_REG_1_ , ADDRESS_REG_0_ , W_R_N_REG , D_C_N_REG , M_IO_N_REG ,
             ADS_N_REG , DATAO_REG_31_ , DATAO_REG_30_ , DATAO_REG_29_ , DATAO_REG_28_ , DATAO_REG_27_ ,
             DATAO_REG_26_ , DATAO_REG_25_ , DATAO_REG_24_ , DATAO_REG_23_ , DATAO_REG_22_ , DATAO_REG_21_ ,
             DATAO_REG_20_ , DATAO_REG_19_ , DATAO_REG_18_ , DATAO_REG_17_ , DATAO_REG_16_ , DATAO_REG_15_ ,
             DATAO_REG_14_ , DATAO_REG_13_ , DATAO_REG_12_ , DATAO_REG_11_ , DATAO_REG_10_ , DATAO_REG_9_ ,
             DATAO_REG_8_ , DATAO_REG_7_ , DATAO_REG_6_ , DATAO_REG_5_ , DATAO_REG_4_ , DATAO_REG_3_ ,
             DATAO_REG_2_ , DATAO_REG_1_ , DATAO_REG_0_ ,
						 
             BE_N_REG_3__EXTRA , BE_N_REG_2__EXTRA , BE_N_REG_1__EXTRA , BE_N_REG_0__EXTRA , ADDRESS_REG_29__EXTRA , ADDRESS_REG_28__EXTRA ,
             ADDRESS_REG_27__EXTRA , ADDRESS_REG_26__EXTRA , ADDRESS_REG_25__EXTRA , ADDRESS_REG_24__EXTRA , ADDRESS_REG_23__EXTRA , ADDRESS_REG_22__EXTRA ,
             ADDRESS_REG_21__EXTRA , ADDRESS_REG_20__EXTRA , ADDRESS_REG_19__EXTRA , ADDRESS_REG_18__EXTRA , ADDRESS_REG_17__EXTRA , ADDRESS_REG_16__EXTRA ,
             ADDRESS_REG_15__EXTRA , ADDRESS_REG_14__EXTRA , ADDRESS_REG_13__EXTRA , ADDRESS_REG_12__EXTRA , ADDRESS_REG_11__EXTRA , ADDRESS_REG_10__EXTRA ,
             ADDRESS_REG_9__EXTRA , ADDRESS_REG_8__EXTRA , ADDRESS_REG_7__EXTRA , ADDRESS_REG_6__EXTRA , ADDRESS_REG_5__EXTRA , ADDRESS_REG_4__EXTRA ,
             ADDRESS_REG_3__EXTRA , ADDRESS_REG_2__EXTRA , ADDRESS_REG_1__EXTRA , ADDRESS_REG_0__EXTRA , STATE_REG_2_ , STATE_REG_1_ ,
             STATE_REG_0_ , DATAWIDTH_REG_0_ , DATAWIDTH_REG_1_ , DATAWIDTH_REG_2_ , DATAWIDTH_REG_3_ , DATAWIDTH_REG_4_ ,
             DATAWIDTH_REG_5_ , DATAWIDTH_REG_6_ , DATAWIDTH_REG_7_ , DATAWIDTH_REG_8_ , DATAWIDTH_REG_9_ , DATAWIDTH_REG_10_ ,
             DATAWIDTH_REG_11_ , DATAWIDTH_REG_12_ , DATAWIDTH_REG_13_ , DATAWIDTH_REG_14_ , DATAWIDTH_REG_15_ , DATAWIDTH_REG_16_ ,
             DATAWIDTH_REG_17_ , DATAWIDTH_REG_18_ , DATAWIDTH_REG_19_ , DATAWIDTH_REG_20_ , DATAWIDTH_REG_21_ , DATAWIDTH_REG_22_ ,
             DATAWIDTH_REG_23_ , DATAWIDTH_REG_24_ , DATAWIDTH_REG_25_ , DATAWIDTH_REG_26_ , DATAWIDTH_REG_27_ , DATAWIDTH_REG_28_ ,
             DATAWIDTH_REG_29_ , DATAWIDTH_REG_30_ , DATAWIDTH_REG_31_ , STATE2_REG_3_ , STATE2_REG_2_ , STATE2_REG_1_ ,
             STATE2_REG_0_ , INSTQUEUE_REG_15__7_ , INSTQUEUE_REG_15__6_ , INSTQUEUE_REG_15__5_ , INSTQUEUE_REG_15__4_ , INSTQUEUE_REG_15__3_ ,
             INSTQUEUE_REG_15__2_ , INSTQUEUE_REG_15__1_ , INSTQUEUE_REG_15__0_ , INSTQUEUE_REG_14__7_ , INSTQUEUE_REG_14__6_ , INSTQUEUE_REG_14__5_ ,
             INSTQUEUE_REG_14__4_ , INSTQUEUE_REG_14__3_ , INSTQUEUE_REG_14__2_ , INSTQUEUE_REG_14__1_ , INSTQUEUE_REG_14__0_ , INSTQUEUE_REG_13__7_ ,
             INSTQUEUE_REG_13__6_ , INSTQUEUE_REG_13__5_ , INSTQUEUE_REG_13__4_ , INSTQUEUE_REG_13__3_ , INSTQUEUE_REG_13__2_ , INSTQUEUE_REG_13__1_ ,
             INSTQUEUE_REG_13__0_ , INSTQUEUE_REG_12__7_ , INSTQUEUE_REG_12__6_ , INSTQUEUE_REG_12__5_ , INSTQUEUE_REG_12__4_ , INSTQUEUE_REG_12__3_ ,
             INSTQUEUE_REG_12__2_ , INSTQUEUE_REG_12__1_ , INSTQUEUE_REG_12__0_ , INSTQUEUE_REG_11__7_ , INSTQUEUE_REG_11__6_ , INSTQUEUE_REG_11__5_ ,
             INSTQUEUE_REG_11__4_ , INSTQUEUE_REG_11__3_ , INSTQUEUE_REG_11__2_ , INSTQUEUE_REG_11__1_ , INSTQUEUE_REG_11__0_ , INSTQUEUE_REG_10__7_ ,
             INSTQUEUE_REG_10__6_ , INSTQUEUE_REG_10__5_ , INSTQUEUE_REG_10__4_ , INSTQUEUE_REG_10__3_ , INSTQUEUE_REG_10__2_ , INSTQUEUE_REG_10__1_ ,
             INSTQUEUE_REG_10__0_ , INSTQUEUE_REG_9__7_ , INSTQUEUE_REG_9__6_ , INSTQUEUE_REG_9__5_ , INSTQUEUE_REG_9__4_ , INSTQUEUE_REG_9__3_ ,
             INSTQUEUE_REG_9__2_ , INSTQUEUE_REG_9__1_ , INSTQUEUE_REG_9__0_ , INSTQUEUE_REG_8__7_ , INSTQUEUE_REG_8__6_ , INSTQUEUE_REG_8__5_ ,
             INSTQUEUE_REG_8__4_ , INSTQUEUE_REG_8__3_ , INSTQUEUE_REG_8__2_ , INSTQUEUE_REG_8__1_ , INSTQUEUE_REG_8__0_ , INSTQUEUE_REG_7__7_ ,
             INSTQUEUE_REG_7__6_ , INSTQUEUE_REG_7__5_ , INSTQUEUE_REG_7__4_ , INSTQUEUE_REG_7__3_ , INSTQUEUE_REG_7__2_ , INSTQUEUE_REG_7__1_ ,
             INSTQUEUE_REG_7__0_ , INSTQUEUE_REG_6__7_ , INSTQUEUE_REG_6__6_ , INSTQUEUE_REG_6__5_ , INSTQUEUE_REG_6__4_ , INSTQUEUE_REG_6__3_ ,
             INSTQUEUE_REG_6__2_ , INSTQUEUE_REG_6__1_ , INSTQUEUE_REG_6__0_ , INSTQUEUE_REG_5__7_ , INSTQUEUE_REG_5__6_ , INSTQUEUE_REG_5__5_ ,
             INSTQUEUE_REG_5__4_ , INSTQUEUE_REG_5__3_ , INSTQUEUE_REG_5__2_ , INSTQUEUE_REG_5__1_ , INSTQUEUE_REG_5__0_ , INSTQUEUE_REG_4__7_ ,
             INSTQUEUE_REG_4__6_ , INSTQUEUE_REG_4__5_ , INSTQUEUE_REG_4__4_ , INSTQUEUE_REG_4__3_ , INSTQUEUE_REG_4__2_ , INSTQUEUE_REG_4__1_ ,
             INSTQUEUE_REG_4__0_ , INSTQUEUE_REG_3__7_ , INSTQUEUE_REG_3__6_ , INSTQUEUE_REG_3__5_ , INSTQUEUE_REG_3__4_ , INSTQUEUE_REG_3__3_ ,
             INSTQUEUE_REG_3__2_ , INSTQUEUE_REG_3__1_ , INSTQUEUE_REG_3__0_ , INSTQUEUE_REG_2__7_ , INSTQUEUE_REG_2__6_ , INSTQUEUE_REG_2__5_ ,
             INSTQUEUE_REG_2__4_ , INSTQUEUE_REG_2__3_ , INSTQUEUE_REG_2__2_ , INSTQUEUE_REG_2__1_ , INSTQUEUE_REG_2__0_ , INSTQUEUE_REG_1__7_ ,
             INSTQUEUE_REG_1__6_ , INSTQUEUE_REG_1__5_ , INSTQUEUE_REG_1__4_ , INSTQUEUE_REG_1__3_ , INSTQUEUE_REG_1__2_ , INSTQUEUE_REG_1__1_ ,
             INSTQUEUE_REG_1__0_ , INSTQUEUE_REG_0__7_ , INSTQUEUE_REG_0__6_ , INSTQUEUE_REG_0__5_ , INSTQUEUE_REG_0__4_ , INSTQUEUE_REG_0__3_ ,
             INSTQUEUE_REG_0__2_ , INSTQUEUE_REG_0__1_ , INSTQUEUE_REG_0__0_ , INSTQUEUERD_ADDR_REG_4_ , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_2_ ,
             INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUEWR_ADDR_REG_4_ , INSTQUEUEWR_ADDR_REG_3_ , INSTQUEUEWR_ADDR_REG_2_ , INSTQUEUEWR_ADDR_REG_1_ ,
             INSTQUEUEWR_ADDR_REG_0_ , INSTADDRPOINTER_REG_0_ , INSTADDRPOINTER_REG_1_ , INSTADDRPOINTER_REG_2_ , INSTADDRPOINTER_REG_3_ , INSTADDRPOINTER_REG_4_ ,
             INSTADDRPOINTER_REG_5_ , INSTADDRPOINTER_REG_6_ , INSTADDRPOINTER_REG_7_ , INSTADDRPOINTER_REG_8_ , INSTADDRPOINTER_REG_9_ , INSTADDRPOINTER_REG_10_ ,
             INSTADDRPOINTER_REG_11_ , INSTADDRPOINTER_REG_12_ , INSTADDRPOINTER_REG_13_ , INSTADDRPOINTER_REG_14_ , INSTADDRPOINTER_REG_15_ , INSTADDRPOINTER_REG_16_ ,
             INSTADDRPOINTER_REG_17_ , INSTADDRPOINTER_REG_18_ , INSTADDRPOINTER_REG_19_ , INSTADDRPOINTER_REG_20_ , INSTADDRPOINTER_REG_21_ , INSTADDRPOINTER_REG_22_ ,
             INSTADDRPOINTER_REG_23_ , INSTADDRPOINTER_REG_24_ , INSTADDRPOINTER_REG_25_ , INSTADDRPOINTER_REG_26_ , INSTADDRPOINTER_REG_27_ , INSTADDRPOINTER_REG_28_ ,
             INSTADDRPOINTER_REG_29_ , INSTADDRPOINTER_REG_30_ , INSTADDRPOINTER_REG_31_ , PHYADDRPOINTER_REG_0_ , PHYADDRPOINTER_REG_1_ , PHYADDRPOINTER_REG_2_ ,
             PHYADDRPOINTER_REG_3_ , PHYADDRPOINTER_REG_4_ , PHYADDRPOINTER_REG_5_ , PHYADDRPOINTER_REG_6_ , PHYADDRPOINTER_REG_7_ , PHYADDRPOINTER_REG_8_ ,
             PHYADDRPOINTER_REG_9_ , PHYADDRPOINTER_REG_10_ , PHYADDRPOINTER_REG_11_ , PHYADDRPOINTER_REG_12_ , PHYADDRPOINTER_REG_13_ , PHYADDRPOINTER_REG_14_ ,
             PHYADDRPOINTER_REG_15_ , PHYADDRPOINTER_REG_16_ , PHYADDRPOINTER_REG_17_ , PHYADDRPOINTER_REG_18_ , PHYADDRPOINTER_REG_19_ , PHYADDRPOINTER_REG_20_ ,
             PHYADDRPOINTER_REG_21_ , PHYADDRPOINTER_REG_22_ , PHYADDRPOINTER_REG_23_ , PHYADDRPOINTER_REG_24_ , PHYADDRPOINTER_REG_25_ , PHYADDRPOINTER_REG_26_ ,
             PHYADDRPOINTER_REG_27_ , PHYADDRPOINTER_REG_28_ , PHYADDRPOINTER_REG_29_ , PHYADDRPOINTER_REG_30_ , PHYADDRPOINTER_REG_31_ , LWORD_REG_15_ ,
             LWORD_REG_14_ , LWORD_REG_13_ , LWORD_REG_12_ , LWORD_REG_11_ , LWORD_REG_10_ , LWORD_REG_9_ ,
             LWORD_REG_8_ , LWORD_REG_7_ , LWORD_REG_6_ , LWORD_REG_5_ , LWORD_REG_4_ , LWORD_REG_3_ ,
             LWORD_REG_2_ , LWORD_REG_1_ , LWORD_REG_0_ , UWORD_REG_14_ , UWORD_REG_13_ , UWORD_REG_12_ ,
             UWORD_REG_11_ , UWORD_REG_10_ , UWORD_REG_9_ , UWORD_REG_8_ , UWORD_REG_7_ , UWORD_REG_6_ ,
             UWORD_REG_5_ , UWORD_REG_4_ , UWORD_REG_3_ , UWORD_REG_2_ , UWORD_REG_1_ , UWORD_REG_0_ ,
             DATAO_REG_0__EXTRA , DATAO_REG_1__EXTRA , DATAO_REG_2__EXTRA , DATAO_REG_3__EXTRA , DATAO_REG_4__EXTRA , DATAO_REG_5__EXTRA ,
             DATAO_REG_6__EXTRA , DATAO_REG_7__EXTRA , DATAO_REG_8__EXTRA , DATAO_REG_9__EXTRA , DATAO_REG_10__EXTRA , DATAO_REG_11__EXTRA ,
             DATAO_REG_12__EXTRA , DATAO_REG_13__EXTRA , DATAO_REG_14__EXTRA , DATAO_REG_15__EXTRA , DATAO_REG_16__EXTRA , DATAO_REG_17__EXTRA ,
             DATAO_REG_18__EXTRA , DATAO_REG_19__EXTRA , DATAO_REG_20__EXTRA , DATAO_REG_21__EXTRA , DATAO_REG_22__EXTRA , DATAO_REG_23__EXTRA ,
             DATAO_REG_24__EXTRA , DATAO_REG_25__EXTRA , DATAO_REG_26__EXTRA , DATAO_REG_27__EXTRA , DATAO_REG_28__EXTRA , DATAO_REG_29__EXTRA ,
             DATAO_REG_30__EXTRA , DATAO_REG_31__EXTRA , EAX_REG_0_ , EAX_REG_1_ , EAX_REG_2_ , EAX_REG_3_ ,
             EAX_REG_4_ , EAX_REG_5_ , EAX_REG_6_ , EAX_REG_7_ , EAX_REG_8_ , EAX_REG_9_ ,
             EAX_REG_10_ , EAX_REG_11_ , EAX_REG_12_ , EAX_REG_13_ , EAX_REG_14_ , EAX_REG_15_ ,
             EAX_REG_16_ , EAX_REG_17_ , EAX_REG_18_ , EAX_REG_19_ , EAX_REG_20_ , EAX_REG_21_ ,
             EAX_REG_22_ , EAX_REG_23_ , EAX_REG_24_ , EAX_REG_25_ , EAX_REG_26_ , EAX_REG_27_ ,
             EAX_REG_28_ , EAX_REG_29_ , EAX_REG_30_ , EAX_REG_31_ , EBX_REG_0_ , EBX_REG_1_ ,
             EBX_REG_2_ , EBX_REG_3_ , EBX_REG_4_ , EBX_REG_5_ , EBX_REG_6_ , EBX_REG_7_ ,
             EBX_REG_8_ , EBX_REG_9_ , EBX_REG_10_ , EBX_REG_11_ , EBX_REG_12_ , EBX_REG_13_ ,
             EBX_REG_14_ , EBX_REG_15_ , EBX_REG_16_ , EBX_REG_17_ , EBX_REG_18_ , EBX_REG_19_ ,
             EBX_REG_20_ , EBX_REG_21_ , EBX_REG_22_ , EBX_REG_23_ , EBX_REG_24_ , EBX_REG_25_ ,
             EBX_REG_26_ , EBX_REG_27_ , EBX_REG_28_ , EBX_REG_29_ , EBX_REG_30_ , EBX_REG_31_ ,
             REIP_REG_0_ , REIP_REG_1_ , REIP_REG_2_ , REIP_REG_3_ , REIP_REG_4_ , REIP_REG_5_ ,
             REIP_REG_6_ , REIP_REG_7_ , REIP_REG_8_ , REIP_REG_9_ , REIP_REG_10_ , REIP_REG_11_ ,
             REIP_REG_12_ , REIP_REG_13_ , REIP_REG_14_ , REIP_REG_15_ , REIP_REG_16_ , REIP_REG_17_ ,
             REIP_REG_18_ , REIP_REG_19_ , REIP_REG_20_ , REIP_REG_21_ , REIP_REG_22_ , REIP_REG_23_ ,
             REIP_REG_24_ , REIP_REG_25_ , REIP_REG_26_ , REIP_REG_27_ , REIP_REG_28_ , REIP_REG_29_ ,
             REIP_REG_30_ , REIP_REG_31_ , BYTEENABLE_REG_3_ , BYTEENABLE_REG_2_ , BYTEENABLE_REG_1_ , BYTEENABLE_REG_0_ ,
             W_R_N_REG_EXTRA , FLUSH_REG , MORE_REG , STATEBS16_REG , REQUESTPENDING_REG , D_C_N_REG_EXTRA ,
             M_IO_N_REG_EXTRA , CODEFETCH_REG , ADS_N_REG_EXTRA , READREQUEST_REG , MEMORYFETCH_REG , DATAI_31_ ,
             DATAI_30_ , DATAI_29_ , DATAI_28_ , DATAI_27_ , DATAI_26_ , DATAI_25_ ,
             DATAI_24_ , DATAI_23_ , DATAI_22_ , DATAI_21_ , DATAI_20_ , DATAI_19_ ,
             DATAI_18_ , DATAI_17_ , DATAI_16_ , DATAI_15_ , DATAI_14_ , DATAI_13_ ,
             DATAI_12_ , DATAI_11_ , DATAI_10_ , DATAI_9_ , DATAI_8_ , DATAI_7_ ,
             DATAI_6_ , DATAI_5_ , DATAI_4_ , DATAI_3_ , DATAI_2_ , DATAI_1_ ,
             DATAI_0_ , NA_N , BS16_N , READY_N , HOLD );

output U3445 , U3446 , U3447 , U3448 , U3213 , U3212 , U3211;
output U3210 , U3209 , U3208 , U3207 , U3206 , U3205 , U3204;
output U3203 , U3202 , U3201 , U3200 , U3199 , U3198 , U3197;
output U3196 , U3195 , U3194 , U3193 , U3192 , U3191 , U3190;
output U3189 , U3188 , U3187 , U3186 , U3185 , U3184 , U3183;
output U3182 , U3181 , U3451 , U3452 , U3180 , U3179 , U3178;
output U3177 , U3176 , U3175 , U3174 , U3173 , U3172 , U3171;
output U3170 , U3169 , U3168 , U3167 , U3166 , U3165 , U3164;
output U3163 , U3162 , U3161 , U3160 , U3159 , U3158 , U3157;
output U3156 , U3155 , U3154 , U3153 , U3152 , U3151 , U3453;
output U3150 , U3149 , U3148 , U3147 , U3146 , U3145 , U3144;
output U3143 , U3142 , U3141 , U3140 , U3139 , U3138 , U3137;
output U3136 , U3135 , U3134 , U3133 , U3132 , U3131 , U3130;
output U3129 , U3128 , U3127 , U3126 , U3125 , U3124 , U3123;
output U3122 , U3121 , U3120 , U3119 , U3118 , U3117 , U3116;
output U3115 , U3114 , U3113 , U3112 , U3111 , U3110 , U3109;
output U3108 , U3107 , U3106 , U3105 , U3104 , U3103 , U3102;
output U3101 , U3100 , U3099 , U3098 , U3097 , U3096 , U3095;
output U3094 , U3093 , U3092 , U3091 , U3090 , U3089 , U3088;
output U3087 , U3086 , U3085 , U3084 , U3083 , U3082 , U3081;
output U3080 , U3079 , U3078 , U3077 , U3076 , U3075 , U3074;
output U3073 , U3072 , U3071 , U3070 , U3069 , U3068 , U3067;
output U3066 , U3065 , U3064 , U3063 , U3062 , U3061 , U3060;
output U3059 , U3058 , U3057 , U3056 , U3055 , U3054 , U3053;
output U3052 , U3051 , U3050 , U3049 , U3048 , U3047 , U3046;
output U3045 , U3044 , U3043 , U3042 , U3041 , U3040 , U3039;
output U3038 , U3037 , U3036 , U3035 , U3034 , U3033 , U3032;
output U3031 , U3030 , U3029 , U3028 , U3027 , U3026 , U3025;
output U3024 , U3023 , U3022 , U3021 , U3020 , U3455 , U3456;
output U3459 , U3460 , U3461 , U3019 , U3462 , U3463 , U3464;
output U3465 , U3018 , U3017 , U3016 , U3015 , U3014 , U3013;
output U3012 , U3011 , U3010 , U3009 , U3008 , U3007 , U3006;
output U3005 , U3004 , U3003 , U3002 , U3001 , U3000 , U2999;
output U2998 , U2997 , U2996 , U2995 , U2994 , U2993 , U2992;
output U2991 , U2990 , U2989 , U2988 , U2987 , U2986 , U2985;
output U2984 , U2983 , U2982 , U2981 , U2980 , U2979 , U2978;
output U2977 , U2976 , U2975 , U2974 , U2973 , U2972 , U2971;
output U2970 , U2969 , U2968 , U2967 , U2966 , U2965 , U2964;
output U2963 , U2962 , U2961 , U2960 , U2959 , U2958 , U2957;
output U2956 , U2955 , U2954 , U2953 , U2952 , U2951 , U2950;
output U2949 , U2948 , U2947 , U2946 , U2945 , U2944 , U2943;
output U2942 , U2941 , U2940 , U2939 , U2938 , U2937 , U2936;
output U2935 , U2934 , U2933 , U2932 , U2931 , U2930 , U2929;
output U2928 , U2927 , U2926 , U2925 , U2924 , U2923 , U2922;
output U2921 , U2920 , U2919 , U2918 , U2917 , U2916 , U2915;
output U2914 , U2913 , U2912 , U2911 , U2910 , U2909 , U2908;
output U2907 , U2906 , U2905 , U2904 , U2903 , U2902 , U2901;
output U2900 , U2899 , U2898 , U2897 , U2896 , U2895 , U2894;
output U2893 , U2892 , U2891 , U2890 , U2889 , U2888 , U2887;
output U2886 , U2885 , U2884 , U2883 , U2882 , U2881 , U2880;
output U2879 , U2878 , U2877 , U2876 , U2875 , U2874 , U2873;
output U2872 , U2871 , U2870 , U2869 , U2868 , U2867 , U2866;
output U2865 , U2864 , U2863 , U2862 , U2861 , U2860 , U2859;
output U2858 , U2857 , U2856 , U2855 , U2854 , U2853 , U2852;
output U2851 , U2850 , U2849 , U2848 , U2847 , U2846 , U2845;
output U2844 , U2843 , U2842 , U2841 , U2840 , U2839 , U2838;
output U2837 , U2836 , U2835 , U2834 , U2833 , U2832 , U2831;
output U2830 , U2829 , U2828 , U2827 , U2826 , U2825 , U2824;
output U2823 , U2822 , U2821 , U2820 , U2819 , U2818 , U2817;
output U2816 , U2815 , U2814 , U2813 , U2812 , U2811 , U2810;
output U2809 , U2808 , U2807 , U2806 , U2805 , U2804 , U2803;
output U2802 , U2801 , U2800 , U2799 , U2798 , U2797 , U2796;
output U2795 , U3468 , U2794 , U3469 , U3470 , U2793 , U3471;
output U2792 , U3472 , U2791 , U3473 , U2790 , U2789 , U3474;
output U2788;
output BE_N_REG_3_ , BE_N_REG_2_ , BE_N_REG_1_ , BE_N_REG_0_ , ADDRESS_REG_29_ , ADDRESS_REG_28_;
output ADDRESS_REG_27_ , ADDRESS_REG_26_ , ADDRESS_REG_25_ , ADDRESS_REG_24_ , ADDRESS_REG_23_ , ADDRESS_REG_22_;
output ADDRESS_REG_21_ , ADDRESS_REG_20_ , ADDRESS_REG_19_ , ADDRESS_REG_18_ , ADDRESS_REG_17_ , ADDRESS_REG_16_;
output ADDRESS_REG_15_ , ADDRESS_REG_14_ , ADDRESS_REG_13_ , ADDRESS_REG_12_ , ADDRESS_REG_11_ , ADDRESS_REG_10_;
output ADDRESS_REG_9_ , ADDRESS_REG_8_ , ADDRESS_REG_7_ , ADDRESS_REG_6_ , ADDRESS_REG_5_ , ADDRESS_REG_4_;
output ADDRESS_REG_3_ , ADDRESS_REG_2_ , ADDRESS_REG_1_ , ADDRESS_REG_0_ , W_R_N_REG , D_C_N_REG;
output M_IO_N_REG , ADS_N_REG , DATAO_REG_31_ , DATAO_REG_30_ , DATAO_REG_29_ , DATAO_REG_28_;
output DATAO_REG_27_ , DATAO_REG_26_ , DATAO_REG_25_ , DATAO_REG_24_ , DATAO_REG_23_ , DATAO_REG_22_;
output DATAO_REG_21_ , DATAO_REG_20_ , DATAO_REG_19_ , DATAO_REG_18_ , DATAO_REG_17_ , DATAO_REG_16_;
output DATAO_REG_15_ , DATAO_REG_14_ , DATAO_REG_13_ , DATAO_REG_12_ , DATAO_REG_11_ , DATAO_REG_10_;
output DATAO_REG_9_ , DATAO_REG_8_ , DATAO_REG_7_ , DATAO_REG_6_ , DATAO_REG_5_ , DATAO_REG_4_;
output DATAO_REG_3_ , DATAO_REG_2_ , DATAO_REG_1_ , DATAO_REG_0_;

input BE_N_REG_3__EXTRA , BE_N_REG_2__EXTRA , BE_N_REG_1__EXTRA , BE_N_REG_0__EXTRA , ADDRESS_REG_29__EXTRA , ADDRESS_REG_28__EXTRA;
input ADDRESS_REG_27__EXTRA , ADDRESS_REG_26__EXTRA , ADDRESS_REG_25__EXTRA , ADDRESS_REG_24__EXTRA , ADDRESS_REG_23__EXTRA , ADDRESS_REG_22__EXTRA;
input ADDRESS_REG_21__EXTRA , ADDRESS_REG_20__EXTRA , ADDRESS_REG_19__EXTRA , ADDRESS_REG_18__EXTRA , ADDRESS_REG_17__EXTRA , ADDRESS_REG_16__EXTRA;
input ADDRESS_REG_15__EXTRA , ADDRESS_REG_14__EXTRA , ADDRESS_REG_13__EXTRA , ADDRESS_REG_12__EXTRA , ADDRESS_REG_11__EXTRA , ADDRESS_REG_10__EXTRA;
input ADDRESS_REG_9__EXTRA , ADDRESS_REG_8__EXTRA , ADDRESS_REG_7__EXTRA , ADDRESS_REG_6__EXTRA , ADDRESS_REG_5__EXTRA , ADDRESS_REG_4__EXTRA;
input ADDRESS_REG_3__EXTRA , ADDRESS_REG_2__EXTRA , ADDRESS_REG_1__EXTRA , ADDRESS_REG_0__EXTRA , STATE_REG_2_ , STATE_REG_1_;
input STATE_REG_0_ , DATAWIDTH_REG_0_ , DATAWIDTH_REG_1_ , DATAWIDTH_REG_2_ , DATAWIDTH_REG_3_ , DATAWIDTH_REG_4_;
input DATAWIDTH_REG_5_ , DATAWIDTH_REG_6_ , DATAWIDTH_REG_7_ , DATAWIDTH_REG_8_ , DATAWIDTH_REG_9_ , DATAWIDTH_REG_10_;
input DATAWIDTH_REG_11_ , DATAWIDTH_REG_12_ , DATAWIDTH_REG_13_ , DATAWIDTH_REG_14_ , DATAWIDTH_REG_15_ , DATAWIDTH_REG_16_;
input DATAWIDTH_REG_17_ , DATAWIDTH_REG_18_ , DATAWIDTH_REG_19_ , DATAWIDTH_REG_20_ , DATAWIDTH_REG_21_ , DATAWIDTH_REG_22_;
input DATAWIDTH_REG_23_ , DATAWIDTH_REG_24_ , DATAWIDTH_REG_25_ , DATAWIDTH_REG_26_ , DATAWIDTH_REG_27_ , DATAWIDTH_REG_28_;
input DATAWIDTH_REG_29_ , DATAWIDTH_REG_30_ , DATAWIDTH_REG_31_ , STATE2_REG_3_ , STATE2_REG_2_ , STATE2_REG_1_;
input STATE2_REG_0_ , INSTQUEUE_REG_15__7_ , INSTQUEUE_REG_15__6_ , INSTQUEUE_REG_15__5_ , INSTQUEUE_REG_15__4_ , INSTQUEUE_REG_15__3_;
input INSTQUEUE_REG_15__2_ , INSTQUEUE_REG_15__1_ , INSTQUEUE_REG_15__0_ , INSTQUEUE_REG_14__7_ , INSTQUEUE_REG_14__6_ , INSTQUEUE_REG_14__5_;
input INSTQUEUE_REG_14__4_ , INSTQUEUE_REG_14__3_ , INSTQUEUE_REG_14__2_ , INSTQUEUE_REG_14__1_ , INSTQUEUE_REG_14__0_ , INSTQUEUE_REG_13__7_;
input INSTQUEUE_REG_13__6_ , INSTQUEUE_REG_13__5_ , INSTQUEUE_REG_13__4_ , INSTQUEUE_REG_13__3_ , INSTQUEUE_REG_13__2_ , INSTQUEUE_REG_13__1_;
input INSTQUEUE_REG_13__0_ , INSTQUEUE_REG_12__7_ , INSTQUEUE_REG_12__6_ , INSTQUEUE_REG_12__5_ , INSTQUEUE_REG_12__4_ , INSTQUEUE_REG_12__3_;
input INSTQUEUE_REG_12__2_ , INSTQUEUE_REG_12__1_ , INSTQUEUE_REG_12__0_ , INSTQUEUE_REG_11__7_ , INSTQUEUE_REG_11__6_ , INSTQUEUE_REG_11__5_;
input INSTQUEUE_REG_11__4_ , INSTQUEUE_REG_11__3_ , INSTQUEUE_REG_11__2_ , INSTQUEUE_REG_11__1_ , INSTQUEUE_REG_11__0_ , INSTQUEUE_REG_10__7_;
input INSTQUEUE_REG_10__6_ , INSTQUEUE_REG_10__5_ , INSTQUEUE_REG_10__4_ , INSTQUEUE_REG_10__3_ , INSTQUEUE_REG_10__2_ , INSTQUEUE_REG_10__1_;
input INSTQUEUE_REG_10__0_ , INSTQUEUE_REG_9__7_ , INSTQUEUE_REG_9__6_ , INSTQUEUE_REG_9__5_ , INSTQUEUE_REG_9__4_ , INSTQUEUE_REG_9__3_;
input INSTQUEUE_REG_9__2_ , INSTQUEUE_REG_9__1_ , INSTQUEUE_REG_9__0_ , INSTQUEUE_REG_8__7_ , INSTQUEUE_REG_8__6_ , INSTQUEUE_REG_8__5_;
input INSTQUEUE_REG_8__4_ , INSTQUEUE_REG_8__3_ , INSTQUEUE_REG_8__2_ , INSTQUEUE_REG_8__1_ , INSTQUEUE_REG_8__0_ , INSTQUEUE_REG_7__7_;
input INSTQUEUE_REG_7__6_ , INSTQUEUE_REG_7__5_ , INSTQUEUE_REG_7__4_ , INSTQUEUE_REG_7__3_ , INSTQUEUE_REG_7__2_ , INSTQUEUE_REG_7__1_;
input INSTQUEUE_REG_7__0_ , INSTQUEUE_REG_6__7_ , INSTQUEUE_REG_6__6_ , INSTQUEUE_REG_6__5_ , INSTQUEUE_REG_6__4_ , INSTQUEUE_REG_6__3_;
input INSTQUEUE_REG_6__2_ , INSTQUEUE_REG_6__1_ , INSTQUEUE_REG_6__0_ , INSTQUEUE_REG_5__7_ , INSTQUEUE_REG_5__6_ , INSTQUEUE_REG_5__5_;
input INSTQUEUE_REG_5__4_ , INSTQUEUE_REG_5__3_ , INSTQUEUE_REG_5__2_ , INSTQUEUE_REG_5__1_ , INSTQUEUE_REG_5__0_ , INSTQUEUE_REG_4__7_;
input INSTQUEUE_REG_4__6_ , INSTQUEUE_REG_4__5_ , INSTQUEUE_REG_4__4_ , INSTQUEUE_REG_4__3_ , INSTQUEUE_REG_4__2_ , INSTQUEUE_REG_4__1_;
input INSTQUEUE_REG_4__0_ , INSTQUEUE_REG_3__7_ , INSTQUEUE_REG_3__6_ , INSTQUEUE_REG_3__5_ , INSTQUEUE_REG_3__4_ , INSTQUEUE_REG_3__3_;
input INSTQUEUE_REG_3__2_ , INSTQUEUE_REG_3__1_ , INSTQUEUE_REG_3__0_ , INSTQUEUE_REG_2__7_ , INSTQUEUE_REG_2__6_ , INSTQUEUE_REG_2__5_;
input INSTQUEUE_REG_2__4_ , INSTQUEUE_REG_2__3_ , INSTQUEUE_REG_2__2_ , INSTQUEUE_REG_2__1_ , INSTQUEUE_REG_2__0_ , INSTQUEUE_REG_1__7_;
input INSTQUEUE_REG_1__6_ , INSTQUEUE_REG_1__5_ , INSTQUEUE_REG_1__4_ , INSTQUEUE_REG_1__3_ , INSTQUEUE_REG_1__2_ , INSTQUEUE_REG_1__1_;
input INSTQUEUE_REG_1__0_ , INSTQUEUE_REG_0__7_ , INSTQUEUE_REG_0__6_ , INSTQUEUE_REG_0__5_ , INSTQUEUE_REG_0__4_ , INSTQUEUE_REG_0__3_;
input INSTQUEUE_REG_0__2_ , INSTQUEUE_REG_0__1_ , INSTQUEUE_REG_0__0_ , INSTQUEUERD_ADDR_REG_4_ , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_2_;
input INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUEWR_ADDR_REG_4_ , INSTQUEUEWR_ADDR_REG_3_ , INSTQUEUEWR_ADDR_REG_2_ , INSTQUEUEWR_ADDR_REG_1_;
input INSTQUEUEWR_ADDR_REG_0_ , INSTADDRPOINTER_REG_0_ , INSTADDRPOINTER_REG_1_ , INSTADDRPOINTER_REG_2_ , INSTADDRPOINTER_REG_3_ , INSTADDRPOINTER_REG_4_;
input INSTADDRPOINTER_REG_5_ , INSTADDRPOINTER_REG_6_ , INSTADDRPOINTER_REG_7_ , INSTADDRPOINTER_REG_8_ , INSTADDRPOINTER_REG_9_ , INSTADDRPOINTER_REG_10_;
input INSTADDRPOINTER_REG_11_ , INSTADDRPOINTER_REG_12_ , INSTADDRPOINTER_REG_13_ , INSTADDRPOINTER_REG_14_ , INSTADDRPOINTER_REG_15_ , INSTADDRPOINTER_REG_16_;
input INSTADDRPOINTER_REG_17_ , INSTADDRPOINTER_REG_18_ , INSTADDRPOINTER_REG_19_ , INSTADDRPOINTER_REG_20_ , INSTADDRPOINTER_REG_21_ , INSTADDRPOINTER_REG_22_;
input INSTADDRPOINTER_REG_23_ , INSTADDRPOINTER_REG_24_ , INSTADDRPOINTER_REG_25_ , INSTADDRPOINTER_REG_26_ , INSTADDRPOINTER_REG_27_ , INSTADDRPOINTER_REG_28_;
input INSTADDRPOINTER_REG_29_ , INSTADDRPOINTER_REG_30_ , INSTADDRPOINTER_REG_31_ , PHYADDRPOINTER_REG_0_ , PHYADDRPOINTER_REG_1_ , PHYADDRPOINTER_REG_2_;
input PHYADDRPOINTER_REG_3_ , PHYADDRPOINTER_REG_4_ , PHYADDRPOINTER_REG_5_ , PHYADDRPOINTER_REG_6_ , PHYADDRPOINTER_REG_7_ , PHYADDRPOINTER_REG_8_;
input PHYADDRPOINTER_REG_9_ , PHYADDRPOINTER_REG_10_ , PHYADDRPOINTER_REG_11_ , PHYADDRPOINTER_REG_12_ , PHYADDRPOINTER_REG_13_ , PHYADDRPOINTER_REG_14_;
input PHYADDRPOINTER_REG_15_ , PHYADDRPOINTER_REG_16_ , PHYADDRPOINTER_REG_17_ , PHYADDRPOINTER_REG_18_ , PHYADDRPOINTER_REG_19_ , PHYADDRPOINTER_REG_20_;
input PHYADDRPOINTER_REG_21_ , PHYADDRPOINTER_REG_22_ , PHYADDRPOINTER_REG_23_ , PHYADDRPOINTER_REG_24_ , PHYADDRPOINTER_REG_25_ , PHYADDRPOINTER_REG_26_;
input PHYADDRPOINTER_REG_27_ , PHYADDRPOINTER_REG_28_ , PHYADDRPOINTER_REG_29_ , PHYADDRPOINTER_REG_30_ , PHYADDRPOINTER_REG_31_ , LWORD_REG_15_;
input LWORD_REG_14_ , LWORD_REG_13_ , LWORD_REG_12_ , LWORD_REG_11_ , LWORD_REG_10_ , LWORD_REG_9_;
input LWORD_REG_8_ , LWORD_REG_7_ , LWORD_REG_6_ , LWORD_REG_5_ , LWORD_REG_4_ , LWORD_REG_3_;
input LWORD_REG_2_ , LWORD_REG_1_ , LWORD_REG_0_ , UWORD_REG_14_ , UWORD_REG_13_ , UWORD_REG_12_;
input UWORD_REG_11_ , UWORD_REG_10_ , UWORD_REG_9_ , UWORD_REG_8_ , UWORD_REG_7_ , UWORD_REG_6_;
input UWORD_REG_5_ , UWORD_REG_4_ , UWORD_REG_3_ , UWORD_REG_2_ , UWORD_REG_1_ , UWORD_REG_0_;
input DATAO_REG_0__EXTRA , DATAO_REG_1__EXTRA , DATAO_REG_2__EXTRA , DATAO_REG_3__EXTRA , DATAO_REG_4__EXTRA , DATAO_REG_5__EXTRA;
input DATAO_REG_6__EXTRA , DATAO_REG_7__EXTRA , DATAO_REG_8__EXTRA , DATAO_REG_9__EXTRA , DATAO_REG_10__EXTRA , DATAO_REG_11__EXTRA;
input DATAO_REG_12__EXTRA , DATAO_REG_13__EXTRA , DATAO_REG_14__EXTRA , DATAO_REG_15__EXTRA , DATAO_REG_16__EXTRA , DATAO_REG_17__EXTRA;
input DATAO_REG_18__EXTRA , DATAO_REG_19__EXTRA , DATAO_REG_20__EXTRA , DATAO_REG_21__EXTRA , DATAO_REG_22__EXTRA , DATAO_REG_23__EXTRA;
input DATAO_REG_24__EXTRA , DATAO_REG_25__EXTRA , DATAO_REG_26__EXTRA , DATAO_REG_27__EXTRA , DATAO_REG_28__EXTRA , DATAO_REG_29__EXTRA;
input DATAO_REG_30__EXTRA , DATAO_REG_31__EXTRA , EAX_REG_0_ , EAX_REG_1_ , EAX_REG_2_ , EAX_REG_3_;
input EAX_REG_4_ , EAX_REG_5_ , EAX_REG_6_ , EAX_REG_7_ , EAX_REG_8_ , EAX_REG_9_;
input EAX_REG_10_ , EAX_REG_11_ , EAX_REG_12_ , EAX_REG_13_ , EAX_REG_14_ , EAX_REG_15_;
input EAX_REG_16_ , EAX_REG_17_ , EAX_REG_18_ , EAX_REG_19_ , EAX_REG_20_ , EAX_REG_21_;
input EAX_REG_22_ , EAX_REG_23_ , EAX_REG_24_ , EAX_REG_25_ , EAX_REG_26_ , EAX_REG_27_;
input EAX_REG_28_ , EAX_REG_29_ , EAX_REG_30_ , EAX_REG_31_ , EBX_REG_0_ , EBX_REG_1_;
input EBX_REG_2_ , EBX_REG_3_ , EBX_REG_4_ , EBX_REG_5_ , EBX_REG_6_ , EBX_REG_7_;
input EBX_REG_8_ , EBX_REG_9_ , EBX_REG_10_ , EBX_REG_11_ , EBX_REG_12_ , EBX_REG_13_;
input EBX_REG_14_ , EBX_REG_15_ , EBX_REG_16_ , EBX_REG_17_ , EBX_REG_18_ , EBX_REG_19_;
input EBX_REG_20_ , EBX_REG_21_ , EBX_REG_22_ , EBX_REG_23_ , EBX_REG_24_ , EBX_REG_25_;
input EBX_REG_26_ , EBX_REG_27_ , EBX_REG_28_ , EBX_REG_29_ , EBX_REG_30_ , EBX_REG_31_;
input REIP_REG_0_ , REIP_REG_1_ , REIP_REG_2_ , REIP_REG_3_ , REIP_REG_4_ , REIP_REG_5_;
input REIP_REG_6_ , REIP_REG_7_ , REIP_REG_8_ , REIP_REG_9_ , REIP_REG_10_ , REIP_REG_11_;
input REIP_REG_12_ , REIP_REG_13_ , REIP_REG_14_ , REIP_REG_15_ , REIP_REG_16_ , REIP_REG_17_;
input REIP_REG_18_ , REIP_REG_19_ , REIP_REG_20_ , REIP_REG_21_ , REIP_REG_22_ , REIP_REG_23_;
input REIP_REG_24_ , REIP_REG_25_ , REIP_REG_26_ , REIP_REG_27_ , REIP_REG_28_ , REIP_REG_29_;
input REIP_REG_30_ , REIP_REG_31_ , BYTEENABLE_REG_3_ , BYTEENABLE_REG_2_ , BYTEENABLE_REG_1_ , BYTEENABLE_REG_0_;
input W_R_N_REG_EXTRA , FLUSH_REG , MORE_REG , STATEBS16_REG , REQUESTPENDING_REG , D_C_N_REG_EXTRA;
input M_IO_N_REG_EXTRA , CODEFETCH_REG , ADS_N_REG_EXTRA , READREQUEST_REG , MEMORYFETCH_REG;
input DATAI_31_ , DATAI_30_ , DATAI_29_ , DATAI_28_ , DATAI_27_ , DATAI_26_;
input DATAI_25_ , DATAI_24_ , DATAI_23_ , DATAI_22_ , DATAI_21_ , DATAI_20_;
input DATAI_19_ , DATAI_18_ , DATAI_17_ , DATAI_16_ , DATAI_15_ , DATAI_14_;
input DATAI_13_ , DATAI_12_ , DATAI_11_ , DATAI_10_ , DATAI_9_ , DATAI_8_;
input DATAI_7_ , DATAI_6_ , DATAI_5_ , DATAI_4_ , DATAI_3_ , DATAI_2_;
input DATAI_1_ , DATAI_0_ , NA_N , BS16_N , READY_N , HOLD;



wire ADD_515_U182 , ADD_515_U181 , ADD_515_U180 , U2352 , U2353 , U2354 , U2355 , U2356 , U2357 , U2358;
wire U2359 , U2360 , U2361 , U2362 , U2363 , U2364 , U2365 , U2366 , U2367 , U2368;
wire U2369 , U2370 , U2371 , U2372 , U2373 , U2374 , U2375 , U2376 , U2377 , U2378;
wire U2379 , U2380 , U2381 , U2382 , U2383 , U2384 , U2385 , U2386 , U2387 , U2388;
wire U2389 , U2390 , U2391 , U2392 , U2393 , U2394 , U2395 , U2396 , U2397 , U2398;
wire U2399 , U2400 , U2401 , U2402 , U2403 , U2404 , U2405 , U2406 , U2407 , U2408;
wire U2409 , U2410 , U2411 , U2412 , U2413 , U2414 , U2415 , U2416 , U2417 , U2418;
wire U2419 , U2420 , U2421 , U2422 , U2423 , U2424 , U2425 , U2426 , U2427 , U2428;
wire U2429 , U2430 , U2431 , U2432 , U2433 , U2434 , U2435 , U2436 , U2437 , U2438;
wire U2439 , U2440 , U2441 , U2442 , U2443 , U2444 , U2445 , U2446 , U2447 , U2448;
wire U2449 , U2450 , U2451 , U2452 , U2453 , U2454 , U2455 , U2456 , U2457 , U2458;
wire U2459 , U2460 , U2461 , U2462 , U2463 , U2464 , U2465 , U2466 , U2467 , U2468;
wire U2469 , U2470 , U2471 , U2472 , U2473 , U2474 , U2475 , U2476 , U2477 , U2478;
wire U2479 , U2480 , U2481 , U2482 , U2483 , U2484 , U2485 , U2486 , U2487 , U2488;
wire U2489 , U2490 , U2491 , U2492 , U2493 , U2494 , U2495 , U2496 , U2497 , U2498;
wire U2499 , U2500 , U2501 , U2502 , U2503 , U2504 , U2505 , U2506 , U2507 , U2508;
wire U2509 , U2510 , U2511 , U2512 , U2513 , U2514 , U2515 , U2516 , U2517 , U2518;
wire U2519 , U2520 , U2521 , U2522 , U2523 , U2524 , U2525 , U2526 , U2527 , U2528;
wire U2529 , U2530 , U2531 , U2532 , U2533 , U2534 , U2535 , U2536 , U2537 , U2538;
wire U2539 , U2540 , U2541 , U2542 , U2543 , U2544 , U2545 , U2546 , U2547 , U2548;
wire U2549 , U2550 , U2551 , U2552 , U2553 , U2554 , U2555 , U2556 , U2557 , U2558;
wire U2559 , U2560 , U2561 , U2562 , U2563 , U2564 , U2565 , U2566 , U2567 , U2568;
wire U2569 , U2570 , U2571 , U2572 , U2573 , U2574 , U2575 , U2576 , U2577 , U2578;
wire U2579 , U2580 , U2581 , U2582 , U2583 , U2584 , U2585 , U2586 , U2587 , U2588;
wire U2589 , U2590 , U2591 , U2592 , U2593 , U2594 , U2595 , U2596 , U2597 , U2598;
wire U2599 , U2600 , U2601 , U2602 , U2603 , U2604 , U2605 , U2606 , U2607 , U2608;
wire U2609 , U2610 , U2611 , U2612 , U2613 , U2614 , U2615 , U2616 , U2617 , U2618;
wire ADD_515_U179 , U2620 , U2621 , U2622 , U2623 , U2624 , U2625 , U2626 , U2627 , U2628;
wire U2629 , U2630 , U2631 , U2632 , U2633 , U2634 , U2635 , U2636 , U2637 , U2638;
wire U2639 , U2640 , U2641 , U2642 , U2643 , U2644 , U2645 , U2646 , U2647 , U2648;
wire U2649 , U2650 , U2651 , U2652 , U2653 , U2654 , U2655 , U2656 , U2657 , U2658;
wire U2659 , U2660 , U2661 , U2662 , U2663 , U2664 , U2665 , U2666 , U2667 , U2668;
wire U2669 , U2670 , U2671 , U2672 , U2673 , U2674 , U2675 , U2676 , U2677 , U2678;
wire U2679 , U2680 , U2681 , U2682 , U2683 , U2684 , U2685 , U2686 , U2687 , U2688;
wire U2689 , U2690 , U2691 , U2692 , U2693 , U2694 , U2695 , U2696 , U2697 , U2698;
wire U2699 , U2700 , U2701 , U2702 , U2703 , U2704 , U2705 , U2706 , U2707 , U2708;
wire U2709 , U2710 , U2711 , U2712 , U2713 , U2714 , U2715 , U2716 , U2717 , U2718;
wire U2719 , U2720 , U2721 , U2722 , U2723 , U2724 , U2725 , U2726 , U2727 , U2728;
wire U2729 , U2730 , U2731 , U2732 , U2733 , U2734 , U2735 , U2736 , U2737 , U2738;
wire U2739 , U2740 , U2741 , U2742 , U2743 , U2744 , U2745 , U2746 , U2747 , U2748;
wire U2749 , U2750 , U2751 , U2752 , U2753 , U2754 , U2755 , U2756 , U2757 , U2758;
wire U2759 , U2760 , U2761 , U2762 , U2763 , U2764 , U2765 , U2766 , U2767 , U2768;
wire U2769 , U2770 , U2771 , U2772 , U2773 , U2774 , U2775 , U2776 , U2777 , U2778;
wire U2779 , U2780 , U2781 , U2782 , U2783 , U2784 , U2785 , U2786 , U2787 , U3214;
wire U3215 , U3216 , U3217 , U3218 , U3219 , U3220 , U3221 , U3222 , U3223 , U3224;
wire U3225 , U3226 , U3227 , U3228 , U3229 , U3230 , U3231 , U3232 , U3233 , U3234;
wire U3235 , U3236 , U3237 , U3238 , U3239 , U3240 , U3241 , U3242 , U3243 , U3244;
wire U3245 , U3246 , U3247 , U3248 , U3249 , U3250 , U3251 , U3252 , U3253 , U3254;
wire U3255 , U3256 , U3257 , U3258 , U3259 , U3260 , U3261 , U3262 , U3263 , U3264;
wire U3265 , U3266 , U3267 , U3268 , U3269 , U3270 , U3271 , U3272 , U3273 , U3274;
wire U3275 , U3276 , U3277 , U3278 , U3279 , U3280 , U3281 , U3282 , U3283 , U3284;
wire U3285 , U3286 , U3287 , U3288 , U3289 , U3290 , U3291 , U3292 , U3293 , U3294;
wire U3295 , U3296 , U3297 , U3298 , U3299 , U3300 , U3301 , U3302 , U3303 , U3304;
wire U3305 , U3306 , U3307 , U3308 , U3309 , U3310 , U3311 , U3312 , U3313 , U3314;
wire U3315 , U3316 , U3317 , U3318 , U3319 , U3320 , U3321 , U3322 , U3323 , U3324;
wire U3325 , U3326 , U3327 , U3328 , U3329 , U3330 , U3331 , U3332 , U3333 , U3334;
wire U3335 , U3336 , U3337 , U3338 , U3339 , U3340 , U3341 , U3342 , U3343 , U3344;
wire U3345 , U3346 , U3347 , U3348 , U3349 , U3350 , U3351 , U3352 , U3353 , U3354;
wire U3355 , U3356 , U3357 , U3358 , U3359 , U3360 , U3361 , U3362 , U3363 , U3364;
wire U3365 , U3366 , U3367 , U3368 , U3369 , U3370 , U3371 , U3372 , U3373 , U3374;
wire U3375 , U3376 , U3377 , U3378 , U3379 , U3380 , U3381 , U3382 , U3383 , U3384;
wire U3385 , U3386 , U3387 , U3388 , U3389 , U3390 , U3391 , U3392 , U3393 , U3394;
wire U3395 , U3396 , U3397 , U3398 , U3399 , U3400 , U3401 , U3402 , U3403 , U3404;
wire U3405 , U3406 , U3407 , U3408 , U3409 , U3410 , U3411 , U3412 , U3413 , U3414;
wire U3415 , U3416 , U3417 , U3418 , U3419 , U3420 , U3421 , U3422 , U3423 , U3424;
wire U3425 , U3426 , U3427 , U3428 , U3429 , U3430 , U3431 , U3432 , U3433 , U3434;
wire U3435 , U3436 , U3437 , U3438 , U3439 , U3440 , U3441 , U3442 , U3443 , U3444;
wire U3449 , U3450 , U3454 , U3457 , U3458 , U3466 , U3467 , U3475 , U3476 , U3477;
wire U3478 , U3479 , U3480 , U3481 , U3482 , U3483 , U3484 , U3485 , U3486 , U3487;
wire U3488 , U3489 , U3490 , U3491 , U3492 , U3493 , U3494 , U3495 , U3496 , U3497;
wire U3498 , U3499 , U3500 , U3501 , U3502 , U3503 , U3504 , U3505 , U3506 , U3507;
wire U3508 , U3509 , U3510 , U3511 , U3512 , U3513 , U3514 , U3515 , U3516 , U3517;
wire U3518 , U3519 , U3520 , U3521 , U3522 , U3523 , U3524 , U3525 , U3526 , U3527;
wire U3528 , U3529 , U3530 , U3531 , U3532 , U3533 , U3534 , U3535 , U3536 , U3537;
wire U3538 , U3539 , U3540 , U3541 , U3542 , U3543 , U3544 , U3545 , U3546 , U3547;
wire U3548 , U3549 , U3550 , U3551 , U3552 , U3553 , U3554 , U3555 , U3556 , U3557;
wire U3558 , U3559 , U3560 , U3561 , U3562 , U3563 , U3564 , U3565 , U3566 , U3567;
wire U3568 , U3569 , U3570 , U3571 , U3572 , U3573 , U3574 , U3575 , U3576 , U3577;
wire U3578 , U3579 , U3580 , U3581 , U3582 , U3583 , U3584 , U3585 , U3586 , U3587;
wire U3588 , U3589 , U3590 , U3591 , U3592 , U3593 , U3594 , U3595 , U3596 , U3597;
wire U3598 , U3599 , U3600 , U3601 , U3602 , U3603 , U3604 , U3605 , U3606 , U3607;
wire U3608 , U3609 , U3610 , U3611 , U3612 , U3613 , U3614 , U3615 , U3616 , U3617;
wire U3618 , U3619 , U3620 , U3621 , U3622 , U3623 , U3624 , U3625 , U3626 , U3627;
wire U3628 , U3629 , U3630 , U3631 , U3632 , U3633 , U3634 , U3635 , U3636 , U3637;
wire U3638 , U3639 , U3640 , U3641 , U3642 , U3643 , U3644 , U3645 , U3646 , U3647;
wire U3648 , U3649 , U3650 , U3651 , U3652 , U3653 , U3654 , U3655 , U3656 , U3657;
wire U3658 , U3659 , U3660 , U3661 , U3662 , U3663 , U3664 , U3665 , U3666 , U3667;
wire U3668 , U3669 , U3670 , U3671 , U3672 , U3673 , U3674 , U3675 , U3676 , U3677;
wire U3678 , U3679 , U3680 , U3681 , U3682 , U3683 , U3684 , U3685 , U3686 , U3687;
wire U3688 , U3689 , U3690 , U3691 , U3692 , U3693 , U3694 , U3695 , U3696 , U3697;
wire U3698 , U3699 , U3700 , U3701 , U3702 , U3703 , U3704 , U3705 , U3706 , U3707;
wire U3708 , U3709 , U3710 , U3711 , U3712 , U3713 , U3714 , U3715 , U3716 , U3717;
wire U3718 , U3719 , U3720 , U3721 , U3722 , U3723 , U3724 , U3725 , U3726 , U3727;
wire U3728 , U3729 , U3730 , U3731 , U3732 , U3733 , U3734 , U3735 , U3736 , U3737;
wire U3738 , U3739 , U3740 , U3741 , U3742 , U3743 , U3744 , U3745 , U3746 , U3747;
wire U3748 , U3749 , U3750 , U3751 , U3752 , U3753 , U3754 , U3755 , U3756 , U3757;
wire U3758 , U3759 , U3760 , U3761 , U3762 , U3763 , U3764 , U3765 , U3766 , U3767;
wire U3768 , U3769 , U3770 , U3771 , U3772 , U3773 , U3774 , U3775 , U3776 , U3777;
wire U3778 , U3779 , U3780 , U3781 , U3782 , U3783 , U3784 , U3785 , U3786 , U3787;
wire U3788 , U3789 , U3790 , U3791 , U3792 , U3793 , U3794 , U3795 , U3796 , U3797;
wire U3798 , U3799 , U3800 , U3801 , U3802 , U3803 , U3804 , U3805 , U3806 , U3807;
wire U3808 , U3809 , U3810 , U3811 , U3812 , U3813 , U3814 , U3815 , U3816 , U3817;
wire U3818 , U3819 , U3820 , U3821 , U3822 , U3823 , U3824 , U3825 , U3826 , U3827;
wire U3828 , U3829 , U3830 , U3831 , U3832 , U3833 , U3834 , U3835 , U3836 , U3837;
wire U3838 , U3839 , U3840 , U3841 , U3842 , U3843 , U3844 , U3845 , U3846 , U3847;
wire U3848 , U3849 , U3850 , U3851 , U3852 , U3853 , U3854 , U3855 , U3856 , U3857;
wire U3858 , U3859 , U3860 , U3861 , U3862 , U3863 , U3864 , U3865 , U3866 , U3867;
wire U3868 , U3869 , U3870 , U3871 , U3872 , U3873 , U3874 , U3875 , U3876 , U3877;
wire U3878 , U3879 , U3880 , U3881 , U3882 , U3883 , U3884 , U3885 , U3886 , U3887;
wire U3888 , U3889 , U3890 , U3891 , U3892 , U3893 , U3894 , U3895 , U3896 , U3897;
wire U3898 , U3899 , U3900 , U3901 , U3902 , U3903 , U3904 , U3905 , U3906 , U3907;
wire U3908 , U3909 , U3910 , U3911 , U3912 , U3913 , U3914 , U3915 , U3916 , U3917;
wire U3918 , U3919 , U3920 , U3921 , U3922 , U3923 , U3924 , U3925 , U3926 , U3927;
wire U3928 , U3929 , U3930 , U3931 , U3932 , U3933 , U3934 , U3935 , U3936 , U3937;
wire U3938 , U3939 , U3940 , U3941 , U3942 , U3943 , U3944 , U3945 , U3946 , U3947;
wire U3948 , U3949 , U3950 , U3951 , U3952 , U3953 , U3954 , U3955 , U3956 , U3957;
wire U3958 , U3959 , U3960 , U3961 , U3962 , U3963 , U3964 , U3965 , U3966 , U3967;
wire U3968 , U3969 , U3970 , U3971 , U3972 , U3973 , U3974 , U3975 , U3976 , U3977;
wire U3978 , U3979 , U3980 , U3981 , U3982 , U3983 , U3984 , U3985 , U3986 , U3987;
wire U3988 , U3989 , U3990 , U3991 , U3992 , U3993 , U3994 , U3995 , U3996 , U3997;
wire U3998 , U3999 , U4000 , U4001 , U4002 , U4003 , U4004 , U4005 , U4006 , U4007;
wire U4008 , U4009 , U4010 , U4011 , U4012 , U4013 , U4014 , U4015 , U4016 , U4017;
wire U4018 , U4019 , U4020 , U4021 , U4022 , U4023 , U4024 , U4025 , U4026 , U4027;
wire U4028 , U4029 , U4030 , U4031 , U4032 , U4033 , U4034 , U4035 , U4036 , U4037;
wire U4038 , U4039 , U4040 , U4041 , U4042 , U4043 , U4044 , U4045 , U4046 , U4047;
wire U4048 , U4049 , U4050 , U4051 , U4052 , U4053 , U4054 , U4055 , U4056 , U4057;
wire U4058 , U4059 , U4060 , U4061 , U4062 , U4063 , U4064 , U4065 , U4066 , U4067;
wire U4068 , U4069 , U4070 , U4071 , U4072 , U4073 , U4074 , U4075 , U4076 , U4077;
wire U4078 , U4079 , U4080 , U4081 , U4082 , U4083 , U4084 , U4085 , U4086 , U4087;
wire U4088 , U4089 , U4090 , U4091 , U4092 , U4093 , U4094 , U4095 , U4096 , U4097;
wire U4098 , U4099 , U4100 , U4101 , U4102 , U4103 , U4104 , U4105 , U4106 , U4107;
wire U4108 , U4109 , U4110 , U4111 , U4112 , U4113 , U4114 , U4115 , U4116 , U4117;
wire U4118 , U4119 , U4120 , U4121 , U4122 , U4123 , U4124 , U4125 , U4126 , U4127;
wire U4128 , U4129 , U4130 , U4131 , U4132 , U4133 , U4134 , U4135 , U4136 , U4137;
wire U4138 , U4139 , U4140 , U4141 , U4142 , U4143 , U4144 , U4145 , U4146 , U4147;
wire U4148 , U4149 , U4150 , U4151 , U4152 , U4153 , U4154 , U4155 , U4156 , U4157;
wire U4158 , U4159 , U4160 , U4161 , U4162 , U4163 , U4164 , U4165 , U4166 , U4167;
wire U4168 , U4169 , U4170 , U4171 , U4172 , U4173 , U4174 , U4175 , U4176 , U4177;
wire U4178 , U4179 , U4180 , U4181 , U4182 , U4183 , U4184 , U4185 , U4186 , U4187;
wire U4188 , U4189 , U4190 , U4191 , U4192 , U4193 , U4194 , U4195 , U4196 , U4197;
wire U4198 , U4199 , U4200 , U4201 , U4202 , U4203 , U4204 , U4205 , U4206 , U4207;
wire U4208 , U4209 , U4210 , U4211 , U4212 , U4213 , U4214 , U4215 , U4216 , U4217;
wire U4218 , U4219 , U4220 , U4221 , U4222 , U4223 , U4224 , U4225 , U4226 , U4227;
wire U4228 , U4229 , U4230 , U4231 , U4232 , U4233 , U4234 , U4235 , U4236 , U4237;
wire U4238 , U4239 , U4240 , U4241 , U4242 , U4243 , U4244 , U4245 , U4246 , U4247;
wire U4248 , U4249 , U4250 , U4251 , U4252 , U4253 , U4254 , U4255 , U4256 , U4257;
wire U4258 , U4259 , U4260 , U4261 , U4262 , U4263 , U4264 , U4265 , U4266 , U4267;
wire U4268 , U4269 , U4270 , U4271 , U4272 , U4273 , U4274 , U4275 , U4276 , U4277;
wire U4278 , U4279 , U4280 , U4281 , U4282 , U4283 , U4284 , U4285 , U4286 , U4287;
wire U4288 , U4289 , U4290 , U4291 , U4292 , U4293 , U4294 , U4295 , U4296 , U4297;
wire U4298 , U4299 , U4300 , U4301 , U4302 , U4303 , U4304 , U4305 , U4306 , U4307;
wire U4308 , U4309 , U4310 , U4311 , U4312 , U4313 , U4314 , U4315 , U4316 , U4317;
wire U4318 , U4319 , U4320 , U4321 , U4322 , U4323 , U4324 , U4325 , U4326 , U4327;
wire U4328 , U4329 , U4330 , U4331 , U4332 , U4333 , U4334 , U4335 , U4336 , U4337;
wire U4338 , U4339 , U4340 , U4341 , U4342 , U4343 , U4344 , U4345 , U4346 , U4347;
wire U4348 , U4349 , U4350 , U4351 , U4352 , U4353 , U4354 , U4355 , U4356 , U4357;
wire U4358 , U4359 , U4360 , U4361 , U4362 , U4363 , U4364 , U4365 , U4366 , U4367;
wire U4368 , U4369 , U4370 , U4371 , U4372 , U4373 , U4374 , U4375 , U4376 , U4377;
wire U4378 , U4379 , U4380 , U4381 , U4382 , U4383 , U4384 , U4385 , U4386 , U4387;
wire U4388 , U4389 , U4390 , U4391 , U4392 , U4393 , U4394 , U4395 , U4396 , U4397;
wire U4398 , U4399 , U4400 , U4401 , U4402 , U4403 , U4404 , U4405 , U4406 , U4407;
wire U4408 , U4409 , U4410 , U4411 , U4412 , U4413 , U4414 , U4415 , U4416 , U4417;
wire U4418 , U4419 , U4420 , U4421 , U4422 , U4423 , U4424 , U4425 , U4426 , U4427;
wire U4428 , U4429 , U4430 , U4431 , U4432 , U4433 , U4434 , U4435 , U4436 , U4437;
wire U4438 , U4439 , U4440 , U4441 , U4442 , U4443 , U4444 , U4445 , U4446 , U4447;
wire U4448 , U4449 , U4450 , U4451 , U4452 , U4453 , U4454 , U4455 , U4456 , U4457;
wire U4458 , U4459 , U4460 , U4461 , U4462 , U4463 , U4464 , U4465 , U4466 , U4467;
wire U4468 , U4469 , U4470 , U4471 , U4472 , U4473 , U4474 , U4475 , U4476 , U4477;
wire U4478 , U4479 , U4480 , U4481 , U4482 , U4483 , U4484 , U4485 , U4486 , U4487;
wire U4488 , U4489 , U4490 , U4491 , U4492 , U4493 , U4494 , U4495 , U4496 , U4497;
wire U4498 , U4499 , U4500 , U4501 , U4502 , U4503 , U4504 , U4505 , U4506 , U4507;
wire U4508 , U4509 , U4510 , U4511 , U4512 , U4513 , U4514 , U4515 , U4516 , U4517;
wire U4518 , U4519 , U4520 , U4521 , U4522 , U4523 , U4524 , U4525 , U4526 , U4527;
wire U4528 , U4529 , U4530 , U4531 , U4532 , U4533 , U4534 , U4535 , U4536 , U4537;
wire U4538 , U4539 , U4540 , U4541 , U4542 , U4543 , U4544 , U4545 , U4546 , U4547;
wire U4548 , U4549 , U4550 , U4551 , U4552 , U4553 , U4554 , U4555 , U4556 , U4557;
wire U4558 , U4559 , U4560 , U4561 , U4562 , U4563 , U4564 , U4565 , U4566 , U4567;
wire U4568 , U4569 , U4570 , U4571 , U4572 , U4573 , U4574 , U4575 , U4576 , U4577;
wire U4578 , U4579 , U4580 , U4581 , U4582 , U4583 , U4584 , U4585 , U4586 , U4587;
wire U4588 , U4589 , U4590 , U4591 , U4592 , U4593 , U4594 , U4595 , U4596 , U4597;
wire U4598 , U4599 , U4600 , U4601 , U4602 , U4603 , U4604 , U4605 , U4606 , U4607;
wire U4608 , U4609 , U4610 , U4611 , U4612 , U4613 , U4614 , U4615 , U4616 , U4617;
wire U4618 , U4619 , U4620 , U4621 , U4622 , U4623 , U4624 , U4625 , U4626 , U4627;
wire U4628 , U4629 , U4630 , U4631 , U4632 , U4633 , U4634 , U4635 , U4636 , U4637;
wire U4638 , U4639 , U4640 , U4641 , U4642 , U4643 , U4644 , U4645 , U4646 , U4647;
wire U4648 , U4649 , U4650 , U4651 , U4652 , U4653 , U4654 , U4655 , U4656 , U4657;
wire U4658 , U4659 , U4660 , U4661 , U4662 , U4663 , U4664 , U4665 , U4666 , U4667;
wire U4668 , U4669 , U4670 , U4671 , U4672 , U4673 , U4674 , U4675 , U4676 , U4677;
wire U4678 , U4679 , U4680 , U4681 , U4682 , U4683 , U4684 , U4685 , U4686 , U4687;
wire U4688 , U4689 , U4690 , U4691 , U4692 , U4693 , U4694 , U4695 , U4696 , U4697;
wire U4698 , U4699 , U4700 , U4701 , U4702 , U4703 , U4704 , U4705 , U4706 , U4707;
wire U4708 , U4709 , U4710 , U4711 , U4712 , U4713 , U4714 , U4715 , U4716 , U4717;
wire U4718 , U4719 , U4720 , U4721 , U4722 , U4723 , U4724 , U4725 , U4726 , U4727;
wire U4728 , U4729 , U4730 , U4731 , U4732 , U4733 , U4734 , U4735 , U4736 , U4737;
wire U4738 , U4739 , U4740 , U4741 , U4742 , U4743 , U4744 , U4745 , U4746 , U4747;
wire U4748 , U4749 , U4750 , U4751 , U4752 , U4753 , U4754 , U4755 , U4756 , U4757;
wire U4758 , U4759 , U4760 , U4761 , U4762 , U4763 , U4764 , U4765 , U4766 , U4767;
wire U4768 , U4769 , U4770 , U4771 , U4772 , U4773 , U4774 , U4775 , U4776 , U4777;
wire U4778 , U4779 , U4780 , U4781 , U4782 , U4783 , U4784 , U4785 , U4786 , U4787;
wire U4788 , U4789 , U4790 , U4791 , U4792 , U4793 , U4794 , U4795 , U4796 , U4797;
wire U4798 , U4799 , U4800 , U4801 , U4802 , U4803 , U4804 , U4805 , U4806 , U4807;
wire U4808 , U4809 , U4810 , U4811 , U4812 , U4813 , U4814 , U4815 , U4816 , U4817;
wire U4818 , U4819 , U4820 , U4821 , U4822 , U4823 , U4824 , U4825 , U4826 , U4827;
wire U4828 , U4829 , U4830 , U4831 , U4832 , U4833 , U4834 , U4835 , U4836 , U4837;
wire U4838 , U4839 , U4840 , U4841 , U4842 , U4843 , U4844 , U4845 , U4846 , U4847;
wire U4848 , U4849 , U4850 , U4851 , U4852 , U4853 , U4854 , U4855 , U4856 , U4857;
wire U4858 , U4859 , U4860 , U4861 , U4862 , U4863 , U4864 , U4865 , U4866 , U4867;
wire U4868 , U4869 , U4870 , U4871 , U4872 , U4873 , U4874 , U4875 , U4876 , U4877;
wire U4878 , U4879 , U4880 , U4881 , U4882 , U4883 , U4884 , U4885 , U4886 , U4887;
wire U4888 , U4889 , U4890 , U4891 , U4892 , U4893 , U4894 , U4895 , U4896 , U4897;
wire U4898 , U4899 , U4900 , U4901 , U4902 , U4903 , U4904 , U4905 , U4906 , U4907;
wire U4908 , U4909 , U4910 , U4911 , U4912 , U4913 , U4914 , U4915 , U4916 , U4917;
wire U4918 , U4919 , U4920 , U4921 , U4922 , U4923 , U4924 , U4925 , U4926 , U4927;
wire U4928 , U4929 , U4930 , U4931 , U4932 , U4933 , U4934 , U4935 , U4936 , U4937;
wire U4938 , U4939 , U4940 , U4941 , U4942 , U4943 , U4944 , U4945 , U4946 , U4947;
wire U4948 , U4949 , U4950 , U4951 , U4952 , U4953 , U4954 , U4955 , U4956 , U4957;
wire U4958 , U4959 , U4960 , U4961 , U4962 , U4963 , U4964 , U4965 , U4966 , U4967;
wire U4968 , U4969 , U4970 , U4971 , U4972 , U4973 , U4974 , U4975 , U4976 , U4977;
wire U4978 , U4979 , U4980 , U4981 , U4982 , U4983 , U4984 , U4985 , U4986 , U4987;
wire U4988 , U4989 , U4990 , U4991 , U4992 , U4993 , U4994 , U4995 , U4996 , U4997;
wire U4998 , U4999 , U5000 , U5001 , U5002 , U5003 , U5004 , U5005 , U5006 , U5007;
wire U5008 , U5009 , U5010 , U5011 , U5012 , U5013 , U5014 , U5015 , U5016 , U5017;
wire U5018 , U5019 , U5020 , U5021 , U5022 , U5023 , U5024 , U5025 , U5026 , U5027;
wire U5028 , U5029 , U5030 , U5031 , U5032 , U5033 , U5034 , U5035 , U5036 , U5037;
wire U5038 , U5039 , U5040 , U5041 , U5042 , U5043 , U5044 , U5045 , U5046 , U5047;
wire U5048 , U5049 , U5050 , U5051 , U5052 , U5053 , U5054 , U5055 , U5056 , U5057;
wire U5058 , U5059 , U5060 , U5061 , U5062 , U5063 , U5064 , U5065 , U5066 , U5067;
wire U5068 , U5069 , U5070 , U5071 , U5072 , U5073 , U5074 , U5075 , U5076 , U5077;
wire U5078 , U5079 , U5080 , U5081 , U5082 , U5083 , U5084 , U5085 , U5086 , U5087;
wire U5088 , U5089 , U5090 , U5091 , U5092 , U5093 , U5094 , U5095 , U5096 , U5097;
wire U5098 , U5099 , U5100 , U5101 , U5102 , U5103 , U5104 , U5105 , U5106 , U5107;
wire U5108 , U5109 , U5110 , U5111 , U5112 , U5113 , U5114 , U5115 , U5116 , U5117;
wire U5118 , U5119 , U5120 , U5121 , U5122 , U5123 , U5124 , U5125 , U5126 , U5127;
wire U5128 , U5129 , U5130 , U5131 , U5132 , U5133 , U5134 , U5135 , U5136 , U5137;
wire U5138 , U5139 , U5140 , U5141 , U5142 , U5143 , U5144 , U5145 , U5146 , U5147;
wire U5148 , U5149 , U5150 , U5151 , U5152 , U5153 , U5154 , U5155 , U5156 , U5157;
wire U5158 , U5159 , U5160 , U5161 , U5162 , U5163 , U5164 , U5165 , U5166 , U5167;
wire U5168 , U5169 , U5170 , U5171 , U5172 , U5173 , U5174 , U5175 , U5176 , U5177;
wire U5178 , U5179 , U5180 , U5181 , U5182 , U5183 , U5184 , U5185 , U5186 , U5187;
wire U5188 , U5189 , U5190 , U5191 , U5192 , U5193 , U5194 , U5195 , U5196 , U5197;
wire U5198 , U5199 , U5200 , U5201 , U5202 , U5203 , U5204 , U5205 , U5206 , U5207;
wire U5208 , U5209 , U5210 , U5211 , U5212 , U5213 , U5214 , U5215 , U5216 , U5217;
wire U5218 , U5219 , U5220 , U5221 , U5222 , U5223 , U5224 , U5225 , U5226 , U5227;
wire U5228 , U5229 , U5230 , U5231 , U5232 , U5233 , U5234 , U5235 , U5236 , U5237;
wire U5238 , U5239 , U5240 , U5241 , U5242 , U5243 , U5244 , U5245 , U5246 , U5247;
wire U5248 , U5249 , U5250 , U5251 , U5252 , U5253 , U5254 , U5255 , U5256 , U5257;
wire U5258 , U5259 , U5260 , U5261 , U5262 , U5263 , U5264 , U5265 , U5266 , U5267;
wire U5268 , U5269 , U5270 , U5271 , U5272 , U5273 , U5274 , U5275 , U5276 , U5277;
wire U5278 , U5279 , U5280 , U5281 , U5282 , U5283 , U5284 , U5285 , U5286 , U5287;
wire U5288 , U5289 , U5290 , U5291 , U5292 , U5293 , U5294 , U5295 , U5296 , U5297;
wire U5298 , U5299 , U5300 , U5301 , U5302 , U5303 , U5304 , U5305 , U5306 , U5307;
wire U5308 , U5309 , U5310 , U5311 , U5312 , U5313 , U5314 , U5315 , U5316 , U5317;
wire U5318 , U5319 , U5320 , U5321 , U5322 , U5323 , U5324 , U5325 , U5326 , U5327;
wire U5328 , U5329 , U5330 , U5331 , U5332 , U5333 , U5334 , U5335 , U5336 , U5337;
wire U5338 , U5339 , U5340 , U5341 , U5342 , U5343 , U5344 , U5345 , U5346 , U5347;
wire U5348 , U5349 , U5350 , U5351 , U5352 , U5353 , U5354 , U5355 , U5356 , U5357;
wire U5358 , U5359 , U5360 , U5361 , U5362 , U5363 , U5364 , U5365 , U5366 , U5367;
wire U5368 , U5369 , U5370 , U5371 , U5372 , U5373 , U5374 , U5375 , U5376 , U5377;
wire U5378 , U5379 , U5380 , U5381 , U5382 , U5383 , U5384 , U5385 , U5386 , U5387;
wire U5388 , U5389 , U5390 , U5391 , U5392 , U5393 , U5394 , U5395 , U5396 , U5397;
wire U5398 , U5399 , U5400 , U5401 , U5402 , U5403 , U5404 , U5405 , U5406 , U5407;
wire U5408 , U5409 , U5410 , U5411 , U5412 , U5413 , U5414 , U5415 , U5416 , U5417;
wire U5418 , U5419 , U5420 , U5421 , U5422 , U5423 , U5424 , U5425 , U5426 , U5427;
wire U5428 , U5429 , U5430 , U5431 , U5432 , U5433 , U5434 , U5435 , U5436 , U5437;
wire U5438 , U5439 , U5440 , U5441 , U5442 , U5443 , U5444 , U5445 , U5446 , U5447;
wire U5448 , U5449 , U5450 , U5451 , U5452 , U5453 , U5454 , U5455 , U5456 , U5457;
wire U5458 , U5459 , U5460 , U5461 , U5462 , U5463 , U5464 , U5465 , U5466 , U5467;
wire U5468 , U5469 , U5470 , U5471 , U5472 , U5473 , U5474 , U5475 , U5476 , U5477;
wire U5478 , U5479 , U5480 , U5481 , U5482 , U5483 , U5484 , U5485 , U5486 , U5487;
wire U5488 , U5489 , U5490 , U5491 , U5492 , U5493 , U5494 , U5495 , U5496 , U5497;
wire U5498 , U5499 , U5500 , U5501 , U5502 , U5503 , U5504 , U5505 , U5506 , U5507;
wire U5508 , U5509 , U5510 , U5511 , U5512 , U5513 , U5514 , U5515 , U5516 , U5517;
wire U5518 , U5519 , U5520 , U5521 , U5522 , U5523 , U5524 , U5525 , U5526 , U5527;
wire U5528 , U5529 , U5530 , U5531 , U5532 , U5533 , U5534 , U5535 , U5536 , U5537;
wire U5538 , U5539 , U5540 , U5541 , U5542 , U5543 , U5544 , U5545 , U5546 , U5547;
wire U5548 , U5549 , U5550 , U5551 , U5552 , U5553 , U5554 , U5555 , U5556 , U5557;
wire U5558 , U5559 , U5560 , U5561 , U5562 , U5563 , U5564 , U5565 , U5566 , U5567;
wire U5568 , U5569 , U5570 , U5571 , U5572 , U5573 , U5574 , U5575 , U5576 , U5577;
wire U5578 , U5579 , U5580 , U5581 , U5582 , U5583 , U5584 , U5585 , U5586 , U5587;
wire U5588 , U5589 , U5590 , U5591 , U5592 , U5593 , U5594 , U5595 , U5596 , U5597;
wire U5598 , U5599 , U5600 , U5601 , U5602 , U5603 , U5604 , U5605 , U5606 , U5607;
wire U5608 , U5609 , U5610 , U5611 , U5612 , U5613 , U5614 , U5615 , U5616 , U5617;
wire U5618 , U5619 , U5620 , U5621 , U5622 , U5623 , U5624 , U5625 , U5626 , U5627;
wire U5628 , U5629 , U5630 , U5631 , U5632 , U5633 , U5634 , U5635 , U5636 , U5637;
wire U5638 , U5639 , U5640 , U5641 , U5642 , U5643 , U5644 , U5645 , U5646 , U5647;
wire U5648 , U5649 , U5650 , U5651 , U5652 , U5653 , U5654 , U5655 , U5656 , U5657;
wire U5658 , U5659 , U5660 , U5661 , U5662 , U5663 , U5664 , U5665 , U5666 , U5667;
wire U5668 , U5669 , U5670 , U5671 , U5672 , U5673 , U5674 , U5675 , U5676 , U5677;
wire U5678 , U5679 , U5680 , U5681 , U5682 , U5683 , U5684 , U5685 , U5686 , U5687;
wire U5688 , U5689 , U5690 , U5691 , U5692 , U5693 , U5694 , U5695 , U5696 , U5697;
wire U5698 , U5699 , U5700 , U5701 , U5702 , U5703 , U5704 , U5705 , U5706 , U5707;
wire U5708 , U5709 , U5710 , U5711 , U5712 , U5713 , U5714 , U5715 , U5716 , U5717;
wire U5718 , U5719 , U5720 , U5721 , U5722 , U5723 , U5724 , U5725 , U5726 , U5727;
wire U5728 , U5729 , U5730 , U5731 , U5732 , U5733 , U5734 , U5735 , U5736 , U5737;
wire U5738 , U5739 , U5740 , U5741 , U5742 , U5743 , U5744 , U5745 , U5746 , U5747;
wire U5748 , U5749 , U5750 , U5751 , U5752 , U5753 , U5754 , U5755 , U5756 , U5757;
wire U5758 , U5759 , U5760 , U5761 , U5762 , U5763 , U5764 , U5765 , U5766 , U5767;
wire U5768 , U5769 , U5770 , U5771 , U5772 , U5773 , U5774 , U5775 , U5776 , U5777;
wire U5778 , U5779 , U5780 , U5781 , U5782 , U5783 , U5784 , U5785 , U5786 , U5787;
wire U5788 , U5789 , U5790 , U5791 , U5792 , U5793 , U5794 , U5795 , U5796 , U5797;
wire U5798 , U5799 , U5800 , U5801 , U5802 , U5803 , U5804 , U5805 , U5806 , U5807;
wire U5808 , U5809 , U5810 , U5811 , U5812 , U5813 , U5814 , U5815 , U5816 , U5817;
wire U5818 , U5819 , U5820 , U5821 , U5822 , U5823 , U5824 , U5825 , U5826 , U5827;
wire U5828 , U5829 , U5830 , U5831 , U5832 , U5833 , U5834 , U5835 , U5836 , U5837;
wire U5838 , U5839 , U5840 , U5841 , U5842 , U5843 , U5844 , U5845 , U5846 , U5847;
wire U5848 , U5849 , U5850 , U5851 , U5852 , U5853 , U5854 , U5855 , U5856 , U5857;
wire U5858 , U5859 , U5860 , U5861 , U5862 , U5863 , U5864 , U5865 , U5866 , U5867;
wire U5868 , U5869 , U5870 , U5871 , U5872 , U5873 , U5874 , U5875 , U5876 , U5877;
wire U5878 , U5879 , U5880 , U5881 , U5882 , U5883 , U5884 , U5885 , U5886 , U5887;
wire U5888 , U5889 , U5890 , U5891 , U5892 , U5893 , U5894 , U5895 , U5896 , U5897;
wire U5898 , U5899 , U5900 , U5901 , U5902 , U5903 , U5904 , U5905 , U5906 , U5907;
wire U5908 , U5909 , U5910 , U5911 , U5912 , U5913 , U5914 , U5915 , U5916 , U5917;
wire U5918 , U5919 , U5920 , U5921 , U5922 , U5923 , U5924 , U5925 , U5926 , U5927;
wire U5928 , U5929 , U5930 , U5931 , U5932 , U5933 , U5934 , U5935 , U5936 , U5937;
wire U5938 , U5939 , U5940 , U5941 , U5942 , U5943 , U5944 , U5945 , U5946 , U5947;
wire U5948 , U5949 , U5950 , U5951 , U5952 , U5953 , U5954 , U5955 , U5956 , U5957;
wire U5958 , U5959 , U5960 , U5961 , U5962 , U5963 , U5964 , U5965 , U5966 , U5967;
wire U5968 , U5969 , U5970 , U5971 , U5972 , U5973 , U5974 , U5975 , U5976 , U5977;
wire U5978 , U5979 , U5980 , U5981 , U5982 , U5983 , U5984 , U5985 , U5986 , U5987;
wire U5988 , U5989 , U5990 , U5991 , U5992 , U5993 , U5994 , U5995 , U5996 , U5997;
wire U5998 , U5999 , U6000 , U6001 , U6002 , U6003 , U6004 , U6005 , U6006 , U6007;
wire U6008 , U6009 , U6010 , U6011 , U6012 , U6013 , U6014 , U6015 , U6016 , U6017;
wire U6018 , U6019 , U6020 , U6021 , U6022 , U6023 , U6024 , U6025 , U6026 , U6027;
wire U6028 , U6029 , U6030 , U6031 , U6032 , U6033 , U6034 , U6035 , U6036 , U6037;
wire U6038 , U6039 , U6040 , U6041 , U6042 , U6043 , U6044 , U6045 , U6046 , U6047;
wire U6048 , U6049 , U6050 , U6051 , U6052 , U6053 , U6054 , U6055 , U6056 , U6057;
wire U6058 , U6059 , U6060 , U6061 , U6062 , U6063 , U6064 , U6065 , U6066 , U6067;
wire U6068 , U6069 , U6070 , U6071 , U6072 , U6073 , U6074 , U6075 , U6076 , U6077;
wire U6078 , U6079 , U6080 , U6081 , U6082 , U6083 , U6084 , U6085 , U6086 , U6087;
wire U6088 , U6089 , U6090 , U6091 , U6092 , U6093 , U6094 , U6095 , U6096 , U6097;
wire U6098 , U6099 , U6100 , U6101 , U6102 , U6103 , U6104 , U6105 , U6106 , U6107;
wire U6108 , U6109 , U6110 , U6111 , U6112 , U6113 , U6114 , U6115 , U6116 , U6117;
wire U6118 , U6119 , U6120 , U6121 , U6122 , U6123 , U6124 , U6125 , U6126 , U6127;
wire U6128 , U6129 , U6130 , U6131 , U6132 , U6133 , U6134 , U6135 , U6136 , U6137;
wire U6138 , U6139 , U6140 , U6141 , U6142 , U6143 , U6144 , U6145 , U6146 , U6147;
wire U6148 , U6149 , U6150 , U6151 , U6152 , U6153 , U6154 , U6155 , U6156 , U6157;
wire U6158 , U6159 , U6160 , U6161 , U6162 , U6163 , U6164 , U6165 , U6166 , U6167;
wire U6168 , U6169 , U6170 , U6171 , U6172 , U6173 , U6174 , U6175 , U6176 , U6177;
wire U6178 , U6179 , U6180 , U6181 , U6182 , U6183 , U6184 , U6185 , U6186 , U6187;
wire U6188 , U6189 , U6190 , U6191 , U6192 , U6193 , U6194 , U6195 , U6196 , U6197;
wire U6198 , U6199 , U6200 , U6201 , U6202 , U6203 , U6204 , U6205 , U6206 , U6207;
wire U6208 , U6209 , U6210 , U6211 , U6212 , U6213 , U6214 , U6215 , U6216 , U6217;
wire U6218 , U6219 , U6220 , U6221 , U6222 , U6223 , U6224 , U6225 , U6226 , U6227;
wire U6228 , U6229 , U6230 , U6231 , U6232 , U6233 , U6234 , U6235 , U6236 , U6237;
wire U6238 , U6239 , U6240 , U6241 , U6242 , U6243 , U6244 , U6245 , U6246 , U6247;
wire U6248 , U6249 , U6250 , U6251 , U6252 , U6253 , U6254 , U6255 , U6256 , U6257;
wire U6258 , U6259 , U6260 , U6261 , U6262 , U6263 , U6264 , U6265 , U6266 , U6267;
wire U6268 , U6269 , U6270 , U6271 , U6272 , U6273 , U6274 , U6275 , U6276 , U6277;
wire U6278 , U6279 , U6280 , U6281 , U6282 , U6283 , U6284 , U6285 , U6286 , U6287;
wire U6288 , U6289 , U6290 , U6291 , U6292 , U6293 , U6294 , U6295 , U6296 , U6297;
wire U6298 , U6299 , U6300 , U6301 , U6302 , U6303 , U6304 , U6305 , U6306 , U6307;
wire U6308 , U6309 , U6310 , U6311 , U6312 , U6313 , U6314 , U6315 , U6316 , U6317;
wire U6318 , U6319 , U6320 , U6321 , U6322 , U6323 , U6324 , U6325 , U6326 , U6327;
wire U6328 , U6329 , U6330 , U6331 , U6332 , U6333 , U6334 , U6335 , U6336 , U6337;
wire U6338 , U6339 , U6340 , U6341 , U6342 , U6343 , U6344 , U6345 , U6346 , U6347;
wire U6348 , U6349 , U6350 , U6351 , U6352 , U6353 , U6354 , U6355 , U6356 , U6357;
wire U6358 , U6359 , U6360 , U6361 , U6362 , U6363 , U6364 , U6365 , U6366 , U6367;
wire U6368 , U6369 , U6370 , U6371 , U6372 , U6373 , U6374 , U6375 , U6376 , U6377;
wire U6378 , U6379 , U6380 , U6381 , U6382 , U6383 , U6384 , U6385 , U6386 , U6387;
wire U6388 , U6389 , U6390 , U6391 , U6392 , U6393 , U6394 , U6395 , U6396 , U6397;
wire U6398 , U6399 , U6400 , U6401 , U6402 , U6403 , U6404 , U6405 , U6406 , U6407;
wire U6408 , U6409 , U6410 , U6411 , U6412 , U6413 , U6414 , U6415 , U6416 , U6417;
wire U6418 , U6419 , U6420 , U6421 , U6422 , U6423 , U6424 , U6425 , U6426 , U6427;
wire U6428 , U6429 , U6430 , U6431 , U6432 , U6433 , U6434 , U6435 , U6436 , U6437;
wire U6438 , U6439 , U6440 , U6441 , U6442 , U6443 , U6444 , U6445 , U6446 , U6447;
wire U6448 , U6449 , U6450 , U6451 , U6452 , U6453 , U6454 , U6455 , U6456 , U6457;
wire U6458 , U6459 , U6460 , U6461 , U6462 , U6463 , U6464 , U6465 , U6466 , U6467;
wire U6468 , U6469 , U6470 , U6471 , U6472 , U6473 , U6474 , U6475 , U6476 , U6477;
wire U6478 , U6479 , U6480 , U6481 , U6482 , U6483 , U6484 , U6485 , U6486 , U6487;
wire U6488 , U6489 , U6490 , U6491 , U6492 , U6493 , U6494 , U6495 , U6496 , U6497;
wire U6498 , U6499 , U6500 , U6501 , U6502 , U6503 , U6504 , U6505 , U6506 , U6507;
wire U6508 , U6509 , U6510 , U6511 , U6512 , U6513 , U6514 , U6515 , U6516 , U6517;
wire U6518 , U6519 , U6520 , U6521 , U6522 , U6523 , U6524 , U6525 , U6526 , U6527;
wire U6528 , U6529 , U6530 , U6531 , U6532 , U6533 , U6534 , U6535 , U6536 , U6537;
wire U6538 , U6539 , U6540 , U6541 , U6542 , U6543 , U6544 , U6545 , U6546 , U6547;
wire U6548 , U6549 , U6550 , U6551 , U6552 , U6553 , U6554 , U6555 , U6556 , U6557;
wire U6558 , U6559 , U6560 , U6561 , U6562 , U6563 , U6564 , U6565 , U6566 , U6567;
wire U6568 , U6569 , U6570 , U6571 , U6572 , U6573 , U6574 , U6575 , U6576 , U6577;
wire U6578 , U6579 , U6580 , U6581 , U6582 , U6583 , U6584 , U6585 , U6586 , U6587;
wire U6588 , U6589 , U6590 , U6591 , U6592 , U6593 , U6594 , U6595 , U6596 , U6597;
wire U6598 , U6599 , U6600 , U6601 , U6602 , U6603 , U6604 , U6605 , U6606 , U6607;
wire U6608 , U6609 , U6610 , U6611 , U6612 , U6613 , U6614 , U6615 , U6616 , U6617;
wire U6618 , U6619 , U6620 , U6621 , U6622 , U6623 , U6624 , U6625 , U6626 , U6627;
wire U6628 , U6629 , U6630 , U6631 , U6632 , U6633 , U6634 , U6635 , U6636 , U6637;
wire U6638 , U6639 , U6640 , U6641 , U6642 , U6643 , U6644 , U6645 , U6646 , U6647;
wire U6648 , U6649 , U6650 , U6651 , U6652 , U6653 , U6654 , U6655 , U6656 , U6657;
wire U6658 , U6659 , U6660 , U6661 , U6662 , U6663 , U6664 , U6665 , U6666 , U6667;
wire U6668 , U6669 , U6670 , U6671 , U6672 , U6673 , U6674 , U6675 , U6676 , U6677;
wire U6678 , U6679 , U6680 , U6681 , U6682 , U6683 , U6684 , U6685 , U6686 , U6687;
wire U6688 , U6689 , U6690 , U6691 , U6692 , U6693 , U6694 , U6695 , U6696 , U6697;
wire U6698 , U6699 , U6700 , U6701 , U6702 , U6703 , U6704 , U6705 , U6706 , U6707;
wire U6708 , U6709 , U6710 , U6711 , U6712 , U6713 , U6714 , U6715 , U6716 , U6717;
wire U6718 , U6719 , U6720 , U6721 , U6722 , U6723 , U6724 , U6725 , U6726 , U6727;
wire U6728 , U6729 , U6730 , U6731 , U6732 , U6733 , U6734 , U6735 , U6736 , U6737;
wire U6738 , U6739 , U6740 , U6741 , U6742 , U6743 , U6744 , U6745 , U6746 , U6747;
wire U6748 , U6749 , U6750 , U6751 , U6752 , U6753 , U6754 , U6755 , U6756 , U6757;
wire U6758 , U6759 , U6760 , U6761 , U6762 , U6763 , U6764 , U6765 , U6766 , U6767;
wire U6768 , U6769 , U6770 , U6771 , U6772 , U6773 , U6774 , U6775 , U6776 , U6777;
wire U6778 , U6779 , U6780 , U6781 , U6782 , U6783 , U6784 , U6785 , U6786 , U6787;
wire U6788 , U6789 , U6790 , U6791 , U6792 , U6793 , U6794 , U6795 , U6796 , U6797;
wire U6798 , U6799 , U6800 , U6801 , U6802 , U6803 , U6804 , U6805 , U6806 , U6807;
wire U6808 , U6809 , U6810 , U6811 , U6812 , U6813 , U6814 , U6815 , U6816 , U6817;
wire U6818 , U6819 , U6820 , U6821 , U6822 , U6823 , U6824 , U6825 , U6826 , U6827;
wire U6828 , U6829 , U6830 , U6831 , U6832 , U6833 , U6834 , U6835 , U6836 , U6837;
wire U6838 , U6839 , U6840 , U6841 , U6842 , U6843 , U6844 , U6845 , U6846 , U6847;
wire U6848 , U6849 , U6850 , U6851 , U6852 , U6853 , U6854 , U6855 , U6856 , U6857;
wire U6858 , U6859 , U6860 , U6861 , U6862 , U6863 , U6864 , U6865 , U6866 , U6867;
wire U6868 , U6869 , U6870 , U6871 , U6872 , U6873 , U6874 , U6875 , U6876 , U6877;
wire U6878 , U6879 , U6880 , U6881 , U6882 , U6883 , U6884 , U6885 , U6886 , U6887;
wire U6888 , U6889 , U6890 , U6891 , U6892 , U6893 , U6894 , U6895 , U6896 , U6897;
wire U6898 , U6899 , U6900 , U6901 , U6902 , U6903 , U6904 , U6905 , U6906 , U6907;
wire U6908 , U6909 , U6910 , U6911 , U6912 , U6913 , U6914 , U6915 , U6916 , U6917;
wire U6918 , U6919 , U6920 , U6921 , U6922 , U6923 , U6924 , U6925 , U6926 , U6927;
wire U6928 , U6929 , U6930 , U6931 , U6932 , U6933 , U6934 , U6935 , U6936 , U6937;
wire U6938 , U6939 , U6940 , U6941 , U6942 , U6943 , U6944 , U6945 , U6946 , U6947;
wire U6948 , U6949 , U6950 , U6951 , U6952 , U6953 , U6954 , U6955 , U6956 , U6957;
wire U6958 , U6959 , U6960 , U6961 , U6962 , U6963 , U6964 , U6965 , U6966 , U6967;
wire U6968 , U6969 , U6970 , U6971 , U6972 , U6973 , U6974 , U6975 , U6976 , U6977;
wire U6978 , U6979 , U6980 , U6981 , U6982 , U6983 , U6984 , U6985 , U6986 , U6987;
wire U6988 , U6989 , U6990 , U6991 , U6992 , U6993 , U6994 , U6995 , U6996 , U6997;
wire U6998 , U6999 , U7000 , U7001 , U7002 , U7003 , U7004 , U7005 , U7006 , U7007;
wire U7008 , U7009 , U7010 , U7011 , U7012 , U7013 , U7014 , U7015 , U7016 , U7017;
wire U7018 , U7019 , U7020 , U7021 , U7022 , U7023 , U7024 , U7025 , U7026 , U7027;
wire U7028 , U7029 , U7030 , U7031 , U7032 , U7033 , U7034 , U7035 , U7036 , U7037;
wire U7038 , U7039 , U7040 , U7041 , U7042 , U7043 , U7044 , U7045 , U7046 , U7047;
wire U7048 , U7049 , U7050 , U7051 , U7052 , U7053 , U7054 , U7055 , U7056 , U7057;
wire U7058 , U7059 , U7060 , U7061 , U7062 , U7063 , U7064 , U7065 , U7066 , U7067;
wire U7068 , U7069 , U7070 , U7071 , U7072 , U7073 , U7074 , U7075 , U7076 , U7077;
wire U7078 , U7079 , U7080 , U7081 , U7082 , U7083 , U7084 , U7085 , U7086 , U7087;
wire U7088 , U7089 , U7090 , U7091 , U7092 , U7093 , U7094 , U7095 , U7096 , U7097;
wire U7098 , U7099 , U7100 , U7101 , U7102 , U7103 , U7104 , U7105 , U7106 , U7107;
wire U7108 , U7109 , U7110 , U7111 , U7112 , U7113 , U7114 , U7115 , U7116 , U7117;
wire U7118 , U7119 , U7120 , U7121 , U7122 , U7123 , U7124 , U7125 , U7126 , U7127;
wire U7128 , U7129 , U7130 , U7131 , U7132 , U7133 , U7134 , U7135 , U7136 , U7137;
wire U7138 , U7139 , U7140 , U7141 , U7142 , U7143 , U7144 , U7145 , U7146 , U7147;
wire U7148 , U7149 , U7150 , U7151 , U7152 , U7153 , U7154 , U7155 , U7156 , U7157;
wire U7158 , U7159 , U7160 , U7161 , U7162 , U7163 , U7164 , U7165 , U7166 , U7167;
wire U7168 , U7169 , U7170 , U7171 , U7172 , U7173 , U7174 , U7175 , U7176 , U7177;
wire U7178 , U7179 , U7180 , U7181 , U7182 , U7183 , U7184 , U7185 , U7186 , U7187;
wire U7188 , U7189 , U7190 , U7191 , U7192 , U7193 , U7194 , U7195 , U7196 , U7197;
wire U7198 , U7199 , U7200 , U7201 , U7202 , U7203 , U7204 , U7205 , U7206 , U7207;
wire U7208 , U7209 , U7210 , U7211 , U7212 , U7213 , U7214 , U7215 , U7216 , U7217;
wire U7218 , U7219 , U7220 , U7221 , U7222 , U7223 , U7224 , U7225 , U7226 , U7227;
wire U7228 , U7229 , U7230 , U7231 , U7232 , U7233 , U7234 , U7235 , U7236 , U7237;
wire U7238 , U7239 , U7240 , U7241 , U7242 , U7243 , U7244 , U7245 , U7246 , U7247;
wire U7248 , U7249 , U7250 , U7251 , U7252 , U7253 , U7254 , U7255 , U7256 , U7257;
wire U7258 , U7259 , U7260 , U7261 , U7262 , U7263 , U7264 , U7265 , U7266 , U7267;
wire U7268 , U7269 , U7270 , U7271 , U7272 , U7273 , U7274 , U7275 , U7276 , U7277;
wire U7278 , U7279 , U7280 , U7281 , U7282 , U7283 , U7284 , U7285 , U7286 , U7287;
wire U7288 , U7289 , U7290 , U7291 , U7292 , U7293 , U7294 , U7295 , U7296 , U7297;
wire U7298 , U7299 , U7300 , U7301 , U7302 , U7303 , U7304 , U7305 , U7306 , U7307;
wire U7308 , U7309 , U7310 , U7311 , U7312 , U7313 , U7314 , U7315 , U7316 , U7317;
wire U7318 , U7319 , U7320 , U7321 , U7322 , U7323 , U7324 , U7325 , U7326 , U7327;
wire U7328 , U7329 , U7330 , U7331 , U7332 , U7333 , U7334 , U7335 , U7336 , U7337;
wire U7338 , U7339 , U7340 , U7341 , U7342 , U7343 , U7344 , U7345 , U7346 , U7347;
wire U7348 , U7349 , U7350 , U7351 , U7352 , U7353 , U7354 , U7355 , U7356 , U7357;
wire U7358 , U7359 , U7360 , U7361 , U7362 , U7363 , U7364 , U7365 , U7366 , U7367;
wire U7368 , U7369 , U7370 , U7371 , U7372 , U7373 , U7374 , U7375 , U7376 , U7377;
wire U7378 , U7379 , U7380 , U7381 , U7382 , U7383 , U7384 , U7385 , U7386 , U7387;
wire U7388 , U7389 , U7390 , U7391 , U7392 , U7393 , U7394 , U7395 , U7396 , U7397;
wire U7398 , U7399 , U7400 , U7401 , U7402 , U7403 , U7404 , U7405 , U7406 , U7407;
wire U7408 , U7409 , U7410 , U7411 , U7412 , U7413 , U7414 , U7415 , U7416 , U7417;
wire U7418 , U7419 , U7420 , U7421 , U7422 , U7423 , U7424 , U7425 , U7426 , U7427;
wire U7428 , U7429 , U7430 , U7431 , U7432 , U7433 , U7434 , U7435 , U7436 , U7437;
wire U7438 , U7439 , U7440 , U7441 , U7442 , U7443 , U7444 , U7445 , U7446 , U7447;
wire U7448 , U7449 , U7450 , U7451 , U7452 , U7453 , U7454 , U7455 , U7456 , U7457;
wire U7458 , U7459 , U7460 , U7461 , U7462 , U7463 , U7464 , U7465 , U7466 , U7467;
wire U7468 , U7469 , U7470 , U7471 , U7472 , U7473 , U7474 , U7475 , U7476 , U7477;
wire U7478 , U7479 , U7480 , U7481 , U7482 , U7483 , U7484 , U7485 , U7486 , U7487;
wire U7488 , U7489 , U7490 , U7491 , U7492 , U7493 , U7494 , U7495 , U7496 , U7497;
wire U7498 , U7499 , U7500 , U7501 , U7502 , U7503 , U7504 , U7505 , U7506 , U7507;
wire U7508 , U7509 , U7510 , U7511 , U7512 , U7513 , U7514 , U7515 , U7516 , U7517;
wire U7518 , U7519 , U7520 , U7521 , U7522 , U7523 , U7524 , U7525 , U7526 , U7527;
wire U7528 , U7529 , U7530 , U7531 , U7532 , U7533 , U7534 , U7535 , U7536 , U7537;
wire U7538 , U7539 , U7540 , U7541 , U7542 , U7543 , U7544 , U7545 , U7546 , U7547;
wire U7548 , U7549 , U7550 , U7551 , U7552 , U7553 , U7554 , U7555 , U7556 , U7557;
wire U7558 , U7559 , U7560 , U7561 , U7562 , U7563 , U7564 , U7565 , U7566 , U7567;
wire U7568 , U7569 , U7570 , U7571 , U7572 , U7573 , U7574 , U7575 , U7576 , U7577;
wire U7578 , U7579 , U7580 , U7581 , U7582 , U7583 , U7584 , U7585 , U7586 , U7587;
wire U7588 , U7589 , U7590 , U7591 , U7592 , U7593 , U7594 , U7595 , U7596 , U7597;
wire U7598 , U7599 , U7600 , U7601 , U7602 , U7603 , U7604 , U7605 , U7606 , U7607;
wire U7608 , U7609 , U7610 , U7611 , U7612 , U7613 , U7614 , U7615 , U7616 , U7617;
wire U7618 , U7619 , U7620 , U7621 , U7622 , U7623 , U7624 , U7625 , U7626 , U7627;
wire U7628 , U7629 , U7630 , U7631 , U7632 , U7633 , U7634 , U7635 , U7636 , U7637;
wire U7638 , U7639 , U7640 , U7641 , U7642 , U7643 , U7644 , U7645 , U7646 , U7647;
wire U7648 , U7649 , U7650 , U7651 , U7652 , U7653 , U7654 , U7655 , U7656 , U7657;
wire U7658 , U7659 , U7660 , U7661 , U7662 , U7663 , U7664 , U7665 , U7666 , U7667;
wire U7668 , U7669 , U7670 , U7671 , U7672 , U7673 , U7674 , U7675 , U7676 , U7677;
wire U7678 , U7679 , U7680 , U7681 , U7682 , U7683 , U7684 , U7685 , U7686 , U7687;
wire U7688 , U7689 , U7690 , U7691 , U7692 , U7693 , U7694 , U7695 , U7696 , U7697;
wire U7698 , U7699 , U7700 , U7701 , U7702 , U7703 , U7704 , U7705 , U7706 , U7707;
wire U7708 , U7709 , U7710 , U7711 , U7712 , U7713 , U7714 , U7715 , U7716 , U7717;
wire U7718 , U7719 , U7720 , U7721 , U7722 , U7723 , U7724 , U7725 , U7726 , U7727;
wire U7728 , U7729 , U7730 , U7731 , U7732 , U7733 , U7734 , U7735 , U7736 , U7737;
wire U7738 , U7739 , U7740 , U7741 , U7742 , U7743 , U7744 , U7745 , U7746 , U7747;
wire U7748 , U7749 , U7750 , U7751 , U7752 , U7753 , U7754 , U7755 , U7756 , U7757;
wire U7758 , U7759 , U7760 , U7761 , U7762 , U7763 , U7764 , U7765 , U7766 , U7767;
wire U7768 , U7769 , U7770 , U7771 , U7772 , U7773 , U7774 , U7775 , U7776 , U7777;
wire U7778 , U7779 , U7780 , U7781 , U7782 , ADD_515_U178 , ADD_515_U177 , ADD_515_U176 , ADD_515_U175 , ADD_515_U174;
wire ADD_515_U173 , ADD_515_U172 , ADD_515_U171 , ADD_515_U170 , ADD_515_U169 , ADD_515_U168 , ADD_515_U167 , ADD_515_U166 , ADD_515_U165 , ADD_515_U164;
wire ADD_515_U163 , ADD_515_U162 , ADD_515_U161 , ADD_515_U160 , ADD_515_U159 , ADD_515_U158 , ADD_515_U157 , ADD_515_U156 , ADD_515_U155 , ADD_515_U154;
wire ADD_515_U153 , ADD_515_U152 , R2027_U5 , R2027_U6 , R2027_U7 , R2027_U8 , R2027_U9 , R2027_U10 , R2027_U11 , R2027_U12;
wire R2027_U13 , R2027_U14 , R2027_U15 , R2027_U16 , R2027_U17 , R2027_U18 , R2027_U19 , R2027_U20 , R2027_U21 , R2027_U22;
wire R2027_U23 , R2027_U24 , R2027_U25 , R2027_U26 , R2027_U27 , R2027_U28 , R2027_U29 , R2027_U30 , R2027_U31 , R2027_U32;
wire R2027_U33 , R2027_U34 , R2027_U35 , R2027_U36 , R2027_U37 , R2027_U38 , R2027_U39 , R2027_U40 , R2027_U41 , R2027_U42;
wire R2027_U43 , R2027_U44 , R2027_U45 , R2027_U46 , R2027_U47 , R2027_U48 , R2027_U49 , R2027_U50 , R2027_U51 , R2027_U52;
wire R2027_U53 , R2027_U54 , R2027_U55 , R2027_U56 , R2027_U57 , R2027_U58 , R2027_U59 , R2027_U60 , R2027_U61 , R2027_U62;
wire R2027_U63 , R2027_U64 , R2027_U65 , R2027_U66 , R2027_U67 , R2027_U68 , R2027_U69 , R2027_U70 , R2027_U71 , R2027_U72;
wire R2027_U73 , R2027_U74 , R2027_U75 , R2027_U76 , R2027_U77 , R2027_U78 , R2027_U79 , R2027_U80 , R2027_U81 , R2027_U82;
wire R2027_U83 , R2027_U84 , R2027_U85 , R2027_U86 , R2027_U87 , R2027_U88 , R2027_U89 , R2027_U90 , R2027_U91 , R2027_U92;
wire R2027_U93 , R2027_U94 , R2027_U95 , R2027_U96 , R2027_U97 , R2027_U98 , R2027_U99 , R2027_U100 , R2027_U101 , R2027_U102;
wire R2027_U103 , R2027_U104 , R2027_U105 , R2027_U106 , R2027_U107 , R2027_U108 , R2027_U109 , R2027_U110 , R2027_U111 , R2027_U112;
wire R2027_U113 , R2027_U114 , R2027_U115 , R2027_U116 , R2027_U117 , R2027_U118 , R2027_U119 , R2027_U120 , R2027_U121 , R2027_U122;
wire R2027_U123 , R2027_U124 , R2027_U125 , R2027_U126 , R2027_U127 , R2027_U128 , R2027_U129 , R2027_U130 , R2027_U131 , R2027_U132;
wire R2027_U133 , R2027_U134 , R2027_U135 , R2027_U136 , R2027_U137 , R2027_U138 , R2027_U139 , R2027_U140 , R2027_U141 , R2027_U142;
wire R2027_U143 , R2027_U144 , R2027_U145 , R2027_U146 , R2027_U147 , R2027_U148 , R2027_U149 , R2027_U150 , R2027_U151 , R2027_U152;
wire R2027_U153 , R2027_U154 , R2027_U155 , R2027_U156 , R2027_U157 , R2027_U158 , R2027_U159 , R2027_U160 , R2027_U161 , R2027_U162;
wire R2027_U163 , R2027_U164 , R2027_U165 , R2027_U166 , R2027_U167 , R2027_U168 , R2027_U169 , R2027_U170 , R2027_U171 , R2027_U172;
wire R2027_U173 , R2027_U174 , R2027_U175 , R2027_U176 , R2027_U177 , R2027_U178 , R2027_U179 , R2027_U180 , R2027_U181 , R2027_U182;
wire R2027_U183 , R2027_U184 , R2027_U185 , R2027_U186 , R2027_U187 , R2027_U188 , R2027_U189 , R2027_U190 , R2027_U191 , R2027_U192;
wire R2027_U193 , R2027_U194 , R2027_U195 , R2027_U196 , R2027_U197 , R2027_U198 , R2027_U199 , R2027_U200 , R2027_U201 , R2027_U202;
wire R2278_U5 , R2278_U6 , R2278_U7 , R2278_U8 , R2278_U9 , R2278_U10 , R2278_U11 , R2278_U12 , R2278_U13 , R2278_U14;
wire R2278_U15 , R2278_U16 , R2278_U17 , R2278_U18 , R2278_U19 , R2278_U20 , R2278_U21 , R2278_U22 , R2278_U23 , R2278_U24;
wire R2278_U25 , R2278_U26 , R2278_U27 , R2278_U28 , R2278_U29 , R2278_U30 , R2278_U31 , R2278_U32 , R2278_U33 , R2278_U34;
wire R2278_U35 , R2278_U36 , R2278_U37 , R2278_U38 , R2278_U39 , R2278_U40 , R2278_U41 , R2278_U42 , R2278_U43 , R2278_U44;
wire R2278_U45 , R2278_U46 , R2278_U47 , R2278_U48 , R2278_U49 , R2278_U50 , R2278_U51 , R2278_U52 , R2278_U53 , R2278_U54;
wire R2278_U55 , R2278_U56 , R2278_U57 , R2278_U58 , R2278_U59 , R2278_U60 , R2278_U61 , R2278_U62 , R2278_U63 , R2278_U64;
wire R2278_U65 , R2278_U66 , R2278_U67 , R2278_U68 , R2278_U69 , R2278_U70 , R2278_U71 , R2278_U72 , R2278_U73 , R2278_U74;
wire R2278_U75 , R2278_U76 , R2278_U77 , R2278_U78 , R2278_U79 , R2278_U80 , R2278_U81 , R2278_U82 , R2278_U83 , R2278_U84;
wire R2278_U85 , R2278_U86 , R2278_U87 , R2278_U88 , R2278_U89 , R2278_U90 , R2278_U91 , R2278_U92 , R2278_U93 , R2278_U94;
wire R2278_U95 , R2278_U96 , R2278_U97 , R2278_U98 , R2278_U99 , R2278_U100 , R2278_U101 , R2278_U102 , R2278_U103 , R2278_U104;
wire R2278_U105 , R2278_U106 , R2278_U107 , R2278_U108 , R2278_U109 , R2278_U110 , R2278_U111 , R2278_U112 , R2278_U113 , R2278_U114;
wire R2278_U115 , R2278_U116 , R2278_U117 , R2278_U118 , R2278_U119 , R2278_U120 , R2278_U121 , R2278_U122 , R2278_U123 , R2278_U124;
wire R2278_U125 , R2278_U126 , R2278_U127 , R2278_U128 , R2278_U129 , R2278_U130 , R2278_U131 , R2278_U132 , R2278_U133 , R2278_U134;
wire R2278_U135 , R2278_U136 , R2278_U137 , R2278_U138 , R2278_U139 , R2278_U140 , R2278_U141 , R2278_U142 , R2278_U143 , R2278_U144;
wire R2278_U145 , R2278_U146 , R2278_U147 , R2278_U148 , R2278_U149 , R2278_U150 , R2278_U151 , R2278_U152 , R2278_U153 , R2278_U154;
wire R2278_U155 , R2278_U156 , R2278_U157 , R2278_U158 , R2278_U159 , R2278_U160 , R2278_U161 , R2278_U162 , R2278_U163 , R2278_U164;
wire R2278_U165 , R2278_U166 , R2278_U167 , R2278_U168 , R2278_U169 , R2278_U170 , R2278_U171 , R2278_U172 , R2278_U173 , R2278_U174;
wire R2278_U175 , R2278_U176 , R2278_U177 , R2278_U178 , R2278_U179 , R2278_U180 , R2278_U181 , R2278_U182 , R2278_U183 , R2278_U184;
wire R2278_U185 , R2278_U186 , R2278_U187 , R2278_U188 , R2278_U189 , R2278_U190 , R2278_U191 , R2278_U192 , R2278_U193 , R2278_U194;
wire R2278_U195 , R2278_U196 , R2278_U197 , R2278_U198 , R2278_U199 , R2278_U200 , R2278_U201 , R2278_U202 , R2278_U203 , R2278_U204;
wire R2278_U205 , R2278_U206 , R2278_U207 , R2278_U208 , R2278_U209 , R2278_U210 , R2278_U211 , R2278_U212 , R2278_U213 , R2278_U214;
wire R2278_U215 , R2278_U216 , R2278_U217 , R2278_U218 , R2278_U219 , R2278_U220 , R2278_U221 , R2278_U222 , R2278_U223 , R2278_U224;
wire R2278_U225 , R2278_U226 , R2278_U227 , R2278_U228 , R2278_U229 , R2278_U230 , R2278_U231 , R2278_U232 , R2278_U233 , R2278_U234;
wire R2278_U235 , R2278_U236 , R2278_U237 , R2278_U238 , R2278_U239 , R2278_U240 , R2278_U241 , R2278_U242 , R2278_U243 , R2278_U244;
wire R2278_U245 , R2278_U246 , R2278_U247 , R2278_U248 , R2278_U249 , R2278_U250 , R2278_U251 , R2278_U252 , R2278_U253 , R2278_U254;
wire R2278_U255 , R2278_U256 , R2278_U257 , R2278_U258 , R2278_U259 , R2278_U260 , R2278_U261 , R2278_U262 , R2278_U263 , R2278_U264;
wire R2278_U265 , R2278_U266 , R2278_U267 , R2278_U268 , R2278_U269 , R2278_U270 , R2278_U271 , R2278_U272 , R2278_U273 , R2278_U274;
wire R2278_U275 , R2278_U276 , R2278_U277 , R2278_U278 , R2278_U279 , R2278_U280 , R2278_U281 , R2278_U282 , R2278_U283 , R2278_U284;
wire R2278_U285 , R2278_U286 , R2278_U287 , R2278_U288 , R2278_U289 , R2278_U290 , R2278_U291 , R2278_U292 , R2278_U293 , R2278_U294;
wire R2278_U295 , R2278_U296 , R2278_U297 , R2278_U298 , R2278_U299 , R2278_U300 , R2278_U301 , R2278_U302 , R2278_U303 , R2278_U304;
wire R2278_U305 , R2278_U306 , R2278_U307 , R2278_U308 , R2278_U309 , R2278_U310 , R2278_U311 , R2278_U312 , R2278_U313 , R2278_U314;
wire R2278_U315 , R2278_U316 , R2278_U317 , R2278_U318 , R2278_U319 , R2278_U320 , R2278_U321 , R2278_U322 , R2278_U323 , R2278_U324;
wire R2278_U325 , R2278_U326 , R2278_U327 , R2278_U328 , R2278_U329 , R2278_U330 , R2278_U331 , R2278_U332 , R2278_U333 , R2278_U334;
wire R2278_U335 , R2278_U336 , R2278_U337 , R2278_U338 , R2278_U339 , R2278_U340 , R2278_U341 , R2278_U342 , R2278_U343 , R2278_U344;
wire R2278_U345 , R2278_U346 , R2278_U347 , R2278_U348 , R2278_U349 , R2278_U350 , R2278_U351 , R2278_U352 , R2278_U353 , R2278_U354;
wire R2278_U355 , R2278_U356 , R2278_U357 , R2278_U358 , R2278_U359 , R2278_U360 , R2278_U361 , R2278_U362 , R2278_U363 , R2278_U364;
wire R2278_U365 , R2278_U366 , R2278_U367 , R2278_U368 , R2278_U369 , R2278_U370 , R2278_U371 , R2278_U372 , R2278_U373 , R2278_U374;
wire R2278_U375 , R2278_U376 , R2278_U377 , R2278_U378 , R2278_U379 , R2278_U380 , R2278_U381 , R2278_U382 , R2278_U383 , R2278_U384;
wire R2278_U385 , R2278_U386 , R2278_U387 , R2278_U388 , R2278_U389 , R2278_U390 , R2278_U391 , R2278_U392 , R2278_U393 , R2278_U394;
wire R2278_U395 , R2278_U396 , R2278_U397 , R2278_U398 , R2278_U399 , R2278_U400 , R2278_U401 , R2278_U402 , R2278_U403 , R2278_U404;
wire R2278_U405 , R2278_U406 , R2278_U407 , R2278_U408 , R2278_U409 , R2278_U410 , R2278_U411 , R2278_U412 , R2278_U413 , R2278_U414;
wire R2278_U415 , R2278_U416 , R2278_U417 , R2278_U418 , R2278_U419 , R2278_U420 , R2278_U421 , R2278_U422 , R2358_U5 , R2358_U6;
wire R2358_U7 , R2358_U8 , R2358_U9 , R2358_U10 , R2358_U11 , R2358_U12 , R2358_U13 , R2358_U14 , R2358_U15 , R2358_U16;
wire R2358_U17 , R2358_U18 , R2358_U19 , R2358_U20 , R2358_U21 , R2358_U22 , R2358_U23 , R2358_U24 , R2358_U25 , R2358_U26;
wire R2358_U27 , R2358_U28 , R2358_U29 , R2358_U30 , R2358_U31 , R2358_U32 , R2358_U33 , R2358_U34 , R2358_U35 , R2358_U36;
wire R2358_U37 , R2358_U38 , R2358_U39 , R2358_U40 , R2358_U41 , R2358_U42 , R2358_U43 , R2358_U44 , R2358_U45 , R2358_U46;
wire R2358_U47 , R2358_U48 , R2358_U49 , R2358_U50 , R2358_U51 , R2358_U52 , R2358_U53 , R2358_U54 , R2358_U55 , R2358_U56;
wire R2358_U57 , R2358_U58 , R2358_U59 , R2358_U60 , R2358_U61 , R2358_U62 , R2358_U63 , R2358_U64 , R2358_U65 , R2358_U66;
wire R2358_U67 , R2358_U68 , R2358_U69 , R2358_U70 , R2358_U71 , R2358_U72 , R2358_U73 , R2358_U74 , R2358_U75 , R2358_U76;
wire R2358_U77 , R2358_U78 , R2358_U79 , R2358_U80 , R2358_U81 , R2358_U82 , R2358_U83 , R2358_U84 , R2358_U85 , R2358_U86;
wire R2358_U87 , R2358_U88 , R2358_U89 , R2358_U90 , R2358_U91 , R2358_U92 , R2358_U93 , R2358_U94 , R2358_U95 , R2358_U96;
wire R2358_U97 , R2358_U98 , R2358_U99 , R2358_U100 , R2358_U101 , R2358_U102 , R2358_U103 , R2358_U104 , R2358_U105 , R2358_U106;
wire R2358_U107 , R2358_U108 , R2358_U109 , R2358_U110 , R2358_U111 , R2358_U112 , R2358_U113 , R2358_U114 , R2358_U115 , R2358_U116;
wire R2358_U117 , R2358_U118 , R2358_U119 , R2358_U120 , R2358_U121 , R2358_U122 , R2358_U123 , R2358_U124 , R2358_U125 , R2358_U126;
wire R2358_U127 , R2358_U128 , R2358_U129 , R2358_U130 , R2358_U131 , R2358_U132 , R2358_U133 , R2358_U134 , R2358_U135 , R2358_U136;
wire R2358_U137 , R2358_U138 , R2358_U139 , R2358_U140 , R2358_U141 , R2358_U142 , R2358_U143 , R2358_U144 , R2358_U145 , R2358_U146;
wire R2358_U147 , R2358_U148 , R2358_U149 , R2358_U150 , R2358_U151 , R2358_U152 , R2358_U153 , R2358_U154 , R2358_U155 , R2358_U156;
wire R2358_U157 , R2358_U158 , R2358_U159 , R2358_U160 , R2358_U161 , R2358_U162 , R2358_U163 , R2358_U164 , R2358_U165 , R2358_U166;
wire R2358_U167 , R2358_U168 , R2358_U169 , R2358_U170 , R2358_U171 , R2358_U172 , R2358_U173 , R2358_U174 , R2358_U175 , R2358_U176;
wire R2358_U177 , R2358_U178 , R2358_U179 , R2358_U180 , R2358_U181 , R2358_U182 , R2358_U183 , R2358_U184 , R2358_U185 , R2358_U186;
wire R2358_U187 , R2358_U188 , R2358_U189 , R2358_U190 , R2358_U191 , R2358_U192 , R2358_U193 , R2358_U194 , R2358_U195 , R2358_U196;
wire R2358_U197 , R2358_U198 , R2358_U199 , R2358_U200 , R2358_U201 , R2358_U202 , R2358_U203 , R2358_U204 , R2358_U205 , R2358_U206;
wire R2358_U207 , R2358_U208 , R2358_U209 , R2358_U210 , R2358_U211 , R2358_U212 , R2358_U213 , R2358_U214 , R2358_U215 , R2358_U216;
wire R2358_U217 , R2358_U218 , R2358_U219 , R2358_U220 , R2358_U221 , R2358_U222 , R2358_U223 , R2358_U224 , R2358_U225 , R2358_U226;
wire R2358_U227 , R2358_U228 , R2358_U229 , R2358_U230 , R2358_U231 , R2358_U232 , R2358_U233 , R2358_U234 , R2358_U235 , R2358_U236;
wire R2358_U237 , R2358_U238 , R2358_U239 , R2358_U240 , R2358_U241 , R2358_U242 , R2358_U243 , R2358_U244 , R2358_U245 , R2358_U246;
wire R2358_U247 , R2358_U248 , R2358_U249 , R2358_U250 , R2358_U251 , R2358_U252 , R2358_U253 , R2358_U254 , R2358_U255 , R2358_U256;
wire R2358_U257 , R2358_U258 , R2358_U259 , R2358_U260 , R2358_U261 , R2358_U262 , R2358_U263 , R2358_U264 , R2358_U265 , R2358_U266;
wire R2358_U267 , R2358_U268 , R2358_U269 , R2358_U270 , R2358_U271 , R2358_U272 , R2358_U273 , R2358_U274 , R2358_U275 , R2358_U276;
wire R2358_U277 , R2358_U278 , R2358_U279 , R2358_U280 , R2358_U281 , R2358_U282 , R2358_U283 , R2358_U284 , R2358_U285 , R2358_U286;
wire R2358_U287 , R2358_U288 , R2358_U289 , R2358_U290 , R2358_U291 , R2358_U292 , R2358_U293 , R2358_U294 , R2358_U295 , R2358_U296;
wire R2358_U297 , R2358_U298 , R2358_U299 , R2358_U300 , R2358_U301 , R2358_U302 , R2358_U303 , R2358_U304 , R2358_U305 , R2358_U306;
wire R2358_U307 , R2358_U308 , R2358_U309 , R2358_U310 , R2358_U311 , R2358_U312 , R2358_U313 , R2358_U314 , R2358_U315 , R2358_U316;
wire R2358_U317 , R2358_U318 , R2358_U319 , R2358_U320 , R2358_U321 , R2358_U322 , R2358_U323 , R2358_U324 , R2358_U325 , R2358_U326;
wire R2358_U327 , R2358_U328 , R2358_U329 , R2358_U330 , R2358_U331 , R2358_U332 , R2358_U333 , R2358_U334 , R2358_U335 , R2358_U336;
wire R2358_U337 , R2358_U338 , R2358_U339 , R2358_U340 , R2358_U341 , R2358_U342 , R2358_U343 , R2358_U344 , R2358_U345 , R2358_U346;
wire R2358_U347 , R2358_U348 , R2358_U349 , R2358_U350 , R2358_U351 , R2358_U352 , R2358_U353 , R2358_U354 , R2358_U355 , R2358_U356;
wire R2358_U357 , R2358_U358 , R2358_U359 , R2358_U360 , R2358_U361 , R2358_U362 , R2358_U363 , R2358_U364 , R2358_U365 , R2358_U366;
wire R2358_U367 , R2358_U368 , R2358_U369 , R2358_U370 , R2358_U371 , R2358_U372 , R2358_U373 , R2358_U374 , R2358_U375 , R2358_U376;
wire R2358_U377 , R2358_U378 , R2358_U379 , R2358_U380 , R2358_U381 , R2358_U382 , R2358_U383 , R2358_U384 , R2358_U385 , R2358_U386;
wire R2358_U387 , R2358_U388 , R2358_U389 , R2358_U390 , R2358_U391 , R2358_U392 , R2358_U393 , R2358_U394 , R2358_U395 , R2358_U396;
wire R2358_U397 , R2358_U398 , R2358_U399 , R2358_U400 , R2358_U401 , R2358_U402 , R2358_U403 , R2358_U404 , R2358_U405 , R2358_U406;
wire R2358_U407 , R2358_U408 , R2358_U409 , R2358_U410 , R2358_U411 , R2358_U412 , R2358_U413 , R2358_U414 , R2358_U415 , R2358_U416;
wire R2358_U417 , R2358_U418 , R2358_U419 , R2358_U420 , R2358_U421 , R2358_U422 , R2358_U423 , R2358_U424 , R2358_U425 , R2358_U426;
wire R2358_U427 , R2358_U428 , R2358_U429 , R2358_U430 , R2358_U431 , R2358_U432 , R2358_U433 , R2358_U434 , R2358_U435 , R2358_U436;
wire R2358_U437 , R2358_U438 , R2358_U439 , R2358_U440 , R2358_U441 , R2358_U442 , R2358_U443 , R2358_U444 , R2358_U445 , R2358_U446;
wire R2358_U447 , R2358_U448 , R2358_U449 , R2358_U450 , R2358_U451 , R2358_U452 , R2358_U453 , R2358_U454 , R2358_U455 , R2358_U456;
wire R2358_U457 , R2358_U458 , R2358_U459 , R2358_U460 , R2358_U461 , R2358_U462 , R2358_U463 , R2358_U464 , R2358_U465 , R2358_U466;
wire R2358_U467 , R2358_U468 , R2358_U469 , R2358_U470 , R2358_U471 , R2358_U472 , R2358_U473 , R2358_U474 , R2358_U475 , R2358_U476;
wire R2358_U477 , R2358_U478 , R2358_U479 , R2358_U480 , R2358_U481 , R2358_U482 , R2358_U483 , R2358_U484 , R2358_U485 , R2358_U486;
wire R2358_U487 , R2358_U488 , R2358_U489 , R2358_U490 , R2358_U491 , R2358_U492 , R2358_U493 , R2358_U494 , R2358_U495 , R2358_U496;
wire R2358_U497 , R2358_U498 , R2358_U499 , R2358_U500 , R2358_U501 , R2358_U502 , R2358_U503 , R2358_U504 , R2358_U505 , R2358_U506;
wire R2358_U507 , R2358_U508 , R2358_U509 , R2358_U510 , R2358_U511 , R2358_U512 , R2358_U513 , R2358_U514 , R2358_U515 , R2358_U516;
wire R2358_U517 , R2358_U518 , R2358_U519 , R2358_U520 , R2358_U521 , R2358_U522 , R2358_U523 , R2358_U524 , R2358_U525 , R2358_U526;
wire R2358_U527 , R2358_U528 , R2358_U529 , R2358_U530 , R2358_U531 , R2358_U532 , R2358_U533 , R2358_U534 , R2358_U535 , R2358_U536;
wire R2358_U537 , R2358_U538 , R2358_U539 , R2358_U540 , R2358_U541 , R2358_U542 , R2358_U543 , R2358_U544 , R2358_U545 , R2358_U546;
wire R2358_U547 , R2358_U548 , R2358_U549 , R2358_U550 , R2358_U551 , R2358_U552 , R2358_U553 , R2358_U554 , R2358_U555 , R2358_U556;
wire R2358_U557 , R2358_U558 , R2358_U559 , R2358_U560 , R2358_U561 , R2358_U562 , R2358_U563 , R2358_U564 , R2358_U565 , R2358_U566;
wire R2358_U567 , R2358_U568 , R2358_U569 , R2358_U570 , R2358_U571 , R2358_U572 , R2358_U573 , R2358_U574 , R2358_U575 , R2358_U576;
wire R2358_U577 , R2358_U578 , R2358_U579 , R2358_U580 , R2358_U581 , R2358_U582 , R2358_U583 , R2358_U584 , R2358_U585 , R2358_U586;
wire R2358_U587 , R2358_U588 , R2358_U589 , R2358_U590 , R2358_U591 , R2358_U592 , R2358_U593 , R2358_U594 , R2358_U595 , R2358_U596;
wire R2358_U597 , R2358_U598 , R2358_U599 , R2358_U600 , R2358_U601 , R2358_U602 , R2358_U603 , R2358_U604 , R2358_U605 , R2358_U606;
wire R2358_U607 , R2358_U608 , R2358_U609 , R2358_U610 , R2358_U611 , R2358_U612 , R2358_U613 , R2358_U614 , R2358_U615 , R2358_U616;
wire R2358_U617 , R2358_U618 , R2358_U619 , R2358_U620 , R2358_U621 , R2358_U622 , R2358_U623 , R2358_U624 , R2358_U625 , R2358_U626;
wire R2358_U627 , R2358_U628 , R2358_U629 , R2358_U630 , R2358_U631 , R2358_U632 , R2358_U633 , R2358_U634 , R2358_U635 , R2358_U636;
wire R2358_U637 , R2358_U638 , R2358_U639 , R2358_U640 , R2358_U641 , R2358_U642 , R2358_U643 , R2358_U644 , R2358_U645 , R2358_U646;
wire R2358_U647 , R2358_U648 , R2358_U649 , R2358_U650 , R2358_U651 , R2358_U652 , R2358_U653 , R2358_U654 , R2337_U5 , R2337_U6;
wire R2337_U7 , R2337_U8 , R2337_U9 , R2337_U10 , R2337_U11 , R2337_U12 , R2337_U13 , R2337_U14 , R2337_U15 , R2337_U16;
wire R2337_U17 , R2337_U18 , R2337_U19 , R2337_U20 , R2337_U21 , R2337_U22 , R2337_U23 , R2337_U24 , R2337_U25 , R2337_U26;
wire R2337_U27 , R2337_U28 , R2337_U29 , R2337_U30 , R2337_U31 , R2337_U32 , R2337_U33 , R2337_U34 , R2337_U35 , R2337_U36;
wire R2337_U37 , R2337_U38 , R2337_U39 , R2337_U40 , R2337_U41 , R2337_U42 , R2337_U43 , R2337_U44 , R2337_U45 , R2337_U46;
wire R2337_U47 , R2337_U48 , R2337_U49 , R2337_U50 , R2337_U51 , R2337_U52 , R2337_U53 , R2337_U54 , R2337_U55 , R2337_U56;
wire R2337_U57 , R2337_U58 , R2337_U59 , R2337_U60 , R2337_U61 , R2337_U62 , R2337_U63 , R2337_U64 , R2337_U65 , R2337_U66;
wire R2337_U67 , R2337_U68 , R2337_U69 , R2337_U70 , R2337_U71 , R2337_U72 , R2337_U73 , R2337_U74 , R2337_U75 , R2337_U76;
wire R2337_U77 , R2337_U78 , R2337_U79 , R2337_U80 , R2337_U81 , R2337_U82 , R2337_U83 , R2337_U84 , R2337_U85 , R2337_U86;
wire R2337_U87 , R2337_U88 , R2337_U89 , R2337_U90 , R2337_U91 , R2337_U92 , R2337_U93 , R2337_U94 , R2337_U95 , R2337_U96;
wire R2337_U97 , R2337_U98 , R2337_U99 , R2337_U100 , R2337_U101 , R2337_U102 , R2337_U103 , R2337_U104 , R2337_U105 , R2337_U106;
wire R2337_U107 , R2337_U108 , R2337_U109 , R2337_U110 , R2337_U111 , R2337_U112 , R2337_U113 , R2337_U114 , R2337_U115 , R2337_U116;
wire R2337_U117 , R2337_U118 , R2337_U119 , R2337_U120 , R2337_U121 , R2337_U122 , R2337_U123 , R2337_U124 , R2337_U125 , R2337_U126;
wire R2337_U127 , R2337_U128 , R2337_U129 , R2337_U130 , R2337_U131 , R2337_U132 , R2337_U133 , R2337_U134 , R2337_U135 , R2337_U136;
wire R2337_U137 , R2337_U138 , R2337_U139 , R2337_U140 , R2337_U141 , R2337_U142 , R2337_U143 , R2337_U144 , R2337_U145 , R2337_U146;
wire R2337_U147 , R2337_U148 , R2337_U149 , R2337_U150 , R2337_U151 , R2337_U152 , R2337_U153 , R2337_U154 , R2337_U155 , R2337_U156;
wire R2337_U157 , R2337_U158 , R2337_U159 , R2337_U160 , R2337_U161 , R2337_U162 , R2337_U163 , R2337_U164 , R2337_U165 , R2337_U166;
wire R2337_U167 , R2337_U168 , R2337_U169 , R2337_U170 , R2337_U171 , R2337_U172 , R2337_U173 , R2337_U174 , R2337_U175 , R2337_U176;
wire R2337_U177 , R2337_U178 , R2337_U179 , R2337_U180 , R2337_U181 , R2337_U182 , R2337_U183 , R2337_U184 , R2337_U185 , R2337_U186;
wire R2337_U187 , R2337_U188 , R2337_U189 , R2337_U190 , R2337_U191 , R2337_U192 , R2337_U193 , R2182_U5 , R2182_U6 , R2182_U7;
wire R2182_U8 , R2182_U9 , R2182_U10 , R2182_U11 , R2182_U12 , R2182_U13 , R2182_U14 , R2182_U15 , R2182_U16 , R2182_U17;
wire R2182_U18 , R2182_U19 , R2182_U20 , R2182_U21 , R2182_U22 , R2182_U23 , R2182_U24 , R2182_U25 , R2182_U26 , R2182_U27;
wire R2182_U28 , R2182_U29 , R2182_U30 , R2182_U31 , R2182_U32 , R2182_U33 , R2182_U34 , R2182_U35 , R2182_U36 , R2182_U37;
wire R2182_U38 , R2182_U39 , R2182_U40 , R2182_U41 , R2182_U42 , R2182_U43 , R2182_U44 , R2182_U45 , R2182_U46 , R2182_U47;
wire R2182_U48 , R2182_U49 , R2182_U50 , R2182_U51 , R2182_U52 , R2182_U53 , R2182_U54 , R2182_U55 , R2182_U56 , R2182_U57;
wire R2182_U58 , R2182_U59 , R2182_U60 , R2182_U61 , R2182_U62 , R2182_U63 , R2182_U64 , R2182_U65 , R2182_U66 , R2182_U67;
wire R2182_U68 , R2182_U69 , R2182_U70 , R2182_U71 , R2182_U72 , R2182_U73 , R2182_U74 , R2182_U75 , R2182_U76 , R2182_U77;
wire R2182_U78 , R2182_U79 , R2182_U80 , R2182_U81 , R2182_U82 , R2182_U83 , R2182_U84 , R2182_U85 , R2182_U86 , R2144_U5;
wire R2144_U6 , R2144_U7 , R2144_U8 , R2144_U9 , R2144_U10 , R2144_U11 , R2144_U12 , R2144_U13 , R2144_U14 , R2144_U15;
wire R2144_U16 , R2144_U17 , R2144_U18 , R2144_U19 , R2144_U20 , R2144_U21 , R2144_U22 , R2144_U23 , R2144_U24 , R2144_U25;
wire R2144_U26 , R2144_U27 , R2144_U28 , R2144_U29 , R2144_U30 , R2144_U31 , R2144_U32 , R2144_U33 , R2144_U34 , R2144_U35;
wire R2144_U36 , R2144_U37 , R2144_U38 , R2144_U39 , R2144_U40 , R2144_U41 , R2144_U42 , R2144_U43 , R2144_U44 , R2144_U45;
wire R2144_U46 , R2144_U47 , R2144_U48 , R2144_U49 , R2144_U50 , R2144_U51 , R2144_U52 , R2144_U53 , R2144_U54 , R2144_U55;
wire R2144_U56 , R2144_U57 , R2144_U58 , R2144_U59 , R2144_U60 , R2144_U61 , R2144_U62 , R2144_U63 , R2144_U64 , R2144_U65;
wire R2144_U66 , R2144_U67 , R2144_U68 , R2144_U69 , R2144_U70 , R2144_U71 , R2144_U72 , R2144_U73 , R2144_U74 , R2144_U75;
wire R2144_U76 , R2144_U77 , R2144_U78 , R2144_U79 , R2144_U80 , R2144_U81 , R2144_U82 , R2144_U83 , R2144_U84 , R2144_U85;
wire R2144_U86 , R2144_U87 , R2144_U88 , R2144_U89 , R2144_U90 , R2144_U91 , R2144_U92 , R2144_U93 , R2144_U94 , R2144_U95;
wire R2144_U96 , R2144_U97 , R2144_U98 , R2144_U99 , R2144_U100 , R2144_U101 , R2144_U102 , R2144_U103 , R2144_U104 , R2144_U105;
wire R2144_U106 , R2144_U107 , R2144_U108 , R2144_U109 , R2144_U110 , R2144_U111 , R2144_U112 , R2144_U113 , R2144_U114 , R2144_U115;
wire R2144_U116 , R2144_U117 , R2144_U118 , R2144_U119 , R2144_U120 , R2144_U121 , R2144_U122 , R2144_U123 , R2144_U124 , R2144_U125;
wire R2144_U126 , R2144_U127 , R2144_U128 , R2144_U129 , R2144_U130 , R2144_U131 , R2144_U132 , R2144_U133 , R2144_U134 , R2144_U135;
wire R2144_U136 , R2144_U137 , R2144_U138 , R2144_U139 , R2144_U140 , R2144_U141 , R2144_U142 , R2144_U143 , R2144_U144 , R2144_U145;
wire R2144_U146 , R2144_U147 , R2144_U148 , R2144_U149 , R2144_U150 , R2144_U151 , R2144_U152 , R2144_U153 , R2144_U154 , R2144_U155;
wire R2144_U156 , R2144_U157 , R2144_U158 , R2144_U159 , R2144_U160 , R2144_U161 , R2144_U162 , R2144_U163 , R2144_U164 , R2144_U165;
wire R2144_U166 , R2144_U167 , R2144_U168 , R2144_U169 , R2144_U170 , R2144_U171 , R2144_U172 , R2144_U173 , R2144_U174 , R2144_U175;
wire R2144_U176 , R2144_U177 , R2144_U178 , R2144_U179 , R2144_U180 , R2144_U181 , R2144_U182 , R2144_U183 , R2144_U184 , R2144_U185;
wire R2144_U186 , R2144_U187 , R2144_U188 , R2144_U189 , R2144_U190 , R2144_U191 , R2144_U192 , R2144_U193 , R2144_U194 , R2144_U195;
wire R2144_U196 , R2144_U197 , R2144_U198 , R2144_U199 , R2144_U200 , R2144_U201 , R2144_U202 , R2144_U203 , R2144_U204 , R2144_U205;
wire R2144_U206 , R2144_U207 , R2144_U208 , R2144_U209 , R2144_U210 , R2144_U211 , R2144_U212 , R2144_U213 , R2144_U214 , R2144_U215;
wire R2144_U216 , R2144_U217 , R2144_U218 , R2144_U219 , R2144_U220 , R2144_U221 , R2144_U222 , R2144_U223 , R2144_U224 , R2144_U225;
wire R2144_U226 , R2144_U227 , R2144_U228 , R2144_U229 , R2144_U230 , R2144_U231 , R2144_U232 , R2144_U233 , R2144_U234 , R2144_U235;
wire R2144_U236 , R2144_U237 , R2144_U238 , R2144_U239 , R2144_U240 , R2144_U241 , R2144_U242 , R2144_U243 , R2144_U244 , R2144_U245;
wire R2144_U246 , R2144_U247 , R2144_U248 , R2144_U249 , R2144_U250 , R2144_U251 , R2144_U252 , R2144_U253 , R2144_U254 , R2144_U255;
wire R2144_U256 , R2144_U257 , R2144_U258 , R2144_U259 , R2144_U260 , LT_589_U6 , LT_589_U7 , LT_589_U8 , R584_U6 , R584_U7;
wire R584_U8 , R584_U9 , R2099_U4 , R2099_U5 , R2099_U6 , R2099_U7 , R2099_U8 , R2099_U9 , R2099_U10 , R2099_U11;
wire R2099_U12 , R2099_U13 , R2099_U14 , R2099_U15 , R2099_U16 , R2099_U17 , R2099_U18 , R2099_U19 , R2099_U20 , R2099_U21;
wire R2099_U22 , R2099_U23 , R2099_U24 , R2099_U25 , R2099_U26 , R2099_U27 , R2099_U28 , R2099_U29 , R2099_U30 , R2099_U31;
wire R2099_U32 , R2099_U33 , R2099_U34 , R2099_U35 , R2099_U36 , R2099_U37 , R2099_U38 , R2099_U39 , R2099_U40 , R2099_U41;
wire R2099_U42 , R2099_U43 , R2099_U44 , R2099_U45 , R2099_U46 , R2099_U47 , R2099_U48 , R2099_U49 , R2099_U50 , R2099_U51;
wire R2099_U52 , R2099_U53 , R2099_U54 , R2099_U55 , R2099_U56 , R2099_U57 , R2099_U58 , R2099_U59 , R2099_U60 , R2099_U61;
wire R2099_U62 , R2099_U63 , R2099_U64 , R2099_U65 , R2099_U66 , R2099_U67 , R2099_U68 , R2099_U69 , R2099_U70 , R2099_U71;
wire R2099_U72 , R2099_U73 , R2099_U74 , R2099_U75 , R2099_U76 , R2099_U77 , R2099_U78 , R2099_U79 , R2099_U80 , R2099_U81;
wire R2099_U82 , R2099_U83 , R2099_U84 , R2099_U85 , R2099_U86 , R2099_U87 , R2099_U88 , R2099_U89 , R2099_U90 , R2099_U91;
wire R2099_U92 , R2099_U93 , R2099_U94 , R2099_U95 , R2099_U96 , R2099_U97 , R2099_U98 , R2099_U99 , R2099_U100 , R2099_U101;
wire R2099_U102 , R2099_U103 , R2099_U104 , R2099_U105 , R2099_U106 , R2099_U107 , R2099_U108 , R2099_U109 , R2099_U110 , R2099_U111;
wire R2099_U112 , R2099_U113 , R2099_U114 , R2099_U115 , R2099_U116 , R2099_U117 , R2099_U118 , R2099_U119 , R2099_U120 , R2099_U121;
wire R2099_U122 , R2099_U123 , R2099_U124 , R2099_U125 , R2099_U126 , R2099_U127 , R2099_U128 , R2099_U129 , R2099_U130 , R2099_U131;
wire R2099_U132 , R2099_U133 , R2099_U134 , R2099_U135 , R2099_U136 , R2099_U137 , R2099_U138 , R2099_U139 , R2099_U140 , R2099_U141;
wire R2099_U142 , R2099_U143 , R2099_U144 , R2099_U145 , R2099_U146 , R2099_U147 , R2099_U148 , R2099_U149 , R2099_U150 , R2099_U151;
wire R2099_U152 , R2099_U153 , R2099_U154 , R2099_U155 , R2099_U156 , R2099_U157 , R2099_U158 , R2099_U159 , R2099_U160 , R2099_U161;
wire R2099_U162 , R2099_U163 , R2099_U164 , R2099_U165 , R2099_U166 , R2099_U167 , R2099_U168 , R2099_U169 , R2099_U170 , R2099_U171;
wire R2099_U172 , R2099_U173 , R2099_U174 , R2099_U175 , R2099_U176 , R2099_U177 , R2099_U178 , R2099_U179 , R2099_U180 , R2099_U181;
wire R2099_U182 , R2099_U183 , R2099_U184 , R2099_U185 , R2099_U186 , R2099_U187 , R2099_U188 , R2099_U189 , R2099_U190 , R2099_U191;
wire R2099_U192 , R2099_U193 , R2099_U194 , R2099_U195 , R2099_U196 , R2099_U197 , R2099_U198 , R2099_U199 , R2099_U200 , R2099_U201;
wire R2099_U202 , R2099_U203 , R2099_U204 , R2099_U205 , R2099_U206 , R2099_U207 , R2099_U208 , R2099_U209 , R2099_U210 , R2099_U211;
wire R2099_U212 , R2099_U213 , R2099_U214 , R2099_U215 , R2099_U216 , R2099_U217 , R2099_U218 , R2099_U219 , R2099_U220 , R2099_U221;
wire R2099_U222 , R2099_U223 , R2099_U224 , R2099_U225 , R2099_U226 , R2099_U227 , R2099_U228 , R2099_U229 , R2099_U230 , R2099_U231;
wire R2099_U232 , R2099_U233 , R2099_U234 , R2099_U235 , R2099_U236 , R2099_U237 , R2099_U238 , R2099_U239 , R2099_U240 , R2099_U241;
wire R2099_U242 , R2099_U243 , R2099_U244 , R2099_U245 , R2099_U246 , R2099_U247 , R2099_U248 , R2099_U249 , R2099_U250 , R2099_U251;
wire R2099_U252 , R2099_U253 , R2099_U254 , R2099_U255 , R2099_U256 , R2099_U257 , R2099_U258 , R2099_U259 , R2099_U260 , R2099_U261;
wire R2099_U262 , R2099_U263 , R2099_U264 , R2099_U265 , R2099_U266 , R2099_U267 , R2099_U268 , R2099_U269 , R2099_U270 , R2099_U271;
wire R2099_U272 , R2099_U273 , R2099_U274 , R2099_U275 , R2099_U276 , R2099_U277 , R2099_U278 , R2099_U279 , R2099_U280 , R2099_U281;
wire R2099_U282 , R2099_U283 , R2099_U284 , R2099_U285 , R2099_U286 , R2099_U287 , R2099_U288 , R2099_U289 , R2099_U290 , R2099_U291;
wire R2099_U292 , R2099_U293 , R2099_U294 , R2099_U295 , R2099_U296 , R2099_U297 , R2099_U298 , R2099_U299 , R2099_U300 , R2099_U301;
wire R2099_U302 , R2099_U303 , R2099_U304 , R2099_U305 , R2099_U306 , R2099_U307 , R2099_U308 , R2099_U309 , R2099_U310 , R2099_U311;
wire R2099_U312 , R2099_U313 , R2099_U314 , R2099_U315 , R2099_U316 , R2099_U317 , R2099_U318 , R2099_U319 , R2099_U320 , R2099_U321;
wire R2099_U322 , R2099_U323 , R2099_U324 , R2099_U325 , R2099_U326 , R2099_U327 , R2099_U328 , R2099_U329 , R2099_U330 , R2099_U331;
wire R2099_U332 , R2099_U333 , R2099_U334 , R2099_U335 , R2099_U336 , R2099_U337 , R2099_U338 , R2099_U339 , R2099_U340 , R2099_U341;
wire R2099_U342 , R2099_U343 , R2099_U344 , R2099_U345 , R2099_U346 , R2099_U347 , R2099_U348 , R2099_U349 , R2167_U6 , R2167_U7;
wire R2167_U8 , R2167_U9 , R2167_U10 , R2167_U11 , R2167_U12 , R2167_U13 , R2167_U14 , R2167_U15 , R2167_U16 , R2167_U17;
wire R2167_U18 , R2167_U19 , R2167_U20 , R2167_U21 , R2167_U22 , R2167_U23 , R2167_U24 , R2167_U25 , R2167_U26 , R2167_U27;
wire R2167_U28 , R2167_U29 , R2167_U30 , R2167_U31 , R2167_U32 , R2167_U33 , R2167_U34 , R2167_U35 , R2167_U36 , R2167_U37;
wire R2167_U38 , R2167_U39 , R2167_U40 , R2167_U41 , R2167_U42 , R2167_U43 , R2167_U44 , R2167_U45 , R2167_U46 , R2167_U47;
wire R2167_U48 , R2167_U49 , R2167_U50 , SUB_357_U6 , SUB_357_U7 , SUB_357_U8 , SUB_357_U9 , SUB_357_U10 , SUB_357_U11 , SUB_357_U12;
wire SUB_357_U13 , LT_563_1260_U6 , LT_563_1260_U7 , LT_563_1260_U8 , LT_563_1260_U9 , SUB_580_U6 , SUB_580_U7 , SUB_580_U8 , SUB_580_U9 , SUB_580_U10;
wire R2096_U4 , R2096_U5 , R2096_U6 , R2096_U7 , R2096_U8 , R2096_U9 , R2096_U10 , R2096_U11 , R2096_U12 , R2096_U13;
wire R2096_U14 , R2096_U15 , R2096_U16 , R2096_U17 , R2096_U18 , R2096_U19 , R2096_U20 , R2096_U21 , R2096_U22 , R2096_U23;
wire R2096_U24 , R2096_U25 , R2096_U26 , R2096_U27 , R2096_U28 , R2096_U29 , R2096_U30 , R2096_U31 , R2096_U32 , R2096_U33;
wire R2096_U34 , R2096_U35 , R2096_U36 , R2096_U37 , R2096_U38 , R2096_U39 , R2096_U40 , R2096_U41 , R2096_U42 , R2096_U43;
wire R2096_U44 , R2096_U45 , R2096_U46 , R2096_U47 , R2096_U48 , R2096_U49 , R2096_U50 , R2096_U51 , R2096_U52 , R2096_U53;
wire R2096_U54 , R2096_U55 , R2096_U56 , R2096_U57 , R2096_U58 , R2096_U59 , R2096_U60 , R2096_U61 , R2096_U62 , R2096_U63;
wire R2096_U64 , R2096_U65 , R2096_U66 , R2096_U67 , R2096_U68 , R2096_U69 , R2096_U70 , R2096_U71 , R2096_U72 , R2096_U73;
wire R2096_U74 , R2096_U75 , R2096_U76 , R2096_U77 , R2096_U78 , R2096_U79 , R2096_U80 , R2096_U81 , R2096_U82 , R2096_U83;
wire R2096_U84 , R2096_U85 , R2096_U86 , R2096_U87 , R2096_U88 , R2096_U89 , R2096_U90 , R2096_U91 , R2096_U92 , R2096_U93;
wire R2096_U94 , R2096_U95 , R2096_U96 , R2096_U97 , R2096_U98 , R2096_U99 , R2096_U100 , R2096_U101 , R2096_U102 , R2096_U103;
wire R2096_U104 , R2096_U105 , R2096_U106 , R2096_U107 , R2096_U108 , R2096_U109 , R2096_U110 , R2096_U111 , R2096_U112 , R2096_U113;
wire R2096_U114 , R2096_U115 , R2096_U116 , R2096_U117 , R2096_U118 , R2096_U119 , R2096_U120 , R2096_U121 , R2096_U122 , R2096_U123;
wire R2096_U124 , R2096_U125 , R2096_U126 , R2096_U127 , R2096_U128 , R2096_U129 , R2096_U130 , R2096_U131 , R2096_U132 , R2096_U133;
wire R2096_U134 , R2096_U135 , R2096_U136 , R2096_U137 , R2096_U138 , R2096_U139 , R2096_U140 , R2096_U141 , R2096_U142 , R2096_U143;
wire R2096_U144 , R2096_U145 , R2096_U146 , R2096_U147 , R2096_U148 , R2096_U149 , R2096_U150 , R2096_U151 , R2096_U152 , R2096_U153;
wire R2096_U154 , R2096_U155 , R2096_U156 , R2096_U157 , R2096_U158 , R2096_U159 , R2096_U160 , R2096_U161 , R2096_U162 , R2096_U163;
wire R2096_U164 , R2096_U165 , R2096_U166 , R2096_U167 , R2096_U168 , R2096_U169 , R2096_U170 , R2096_U171 , R2096_U172 , R2096_U173;
wire R2096_U174 , R2096_U175 , R2096_U176 , R2096_U177 , R2096_U178 , R2096_U179 , R2096_U180 , R2096_U181 , R2096_U182 , LT_563_U6;
wire LT_563_U7 , LT_563_U8 , LT_563_U9 , LT_563_U10 , LT_563_U11 , LT_563_U12 , LT_563_U13 , LT_563_U14 , LT_563_U15 , LT_563_U16;
wire LT_563_U17 , LT_563_U18 , LT_563_U19 , LT_563_U20 , LT_563_U21 , LT_563_U22 , LT_563_U23 , LT_563_U24 , LT_563_U25 , LT_563_U26;
wire LT_563_U27 , LT_563_U28 , R2238_U6 , R2238_U7 , R2238_U8 , R2238_U9 , R2238_U10 , R2238_U11 , R2238_U12 , R2238_U13;
wire R2238_U14 , R2238_U15 , R2238_U16 , R2238_U17 , R2238_U18 , R2238_U19 , R2238_U20 , R2238_U21 , R2238_U22 , R2238_U23;
wire R2238_U24 , R2238_U25 , R2238_U26 , R2238_U27 , R2238_U28 , R2238_U29 , R2238_U30 , R2238_U31 , R2238_U32 , R2238_U33;
wire R2238_U34 , R2238_U35 , R2238_U36 , R2238_U37 , R2238_U38 , R2238_U39 , R2238_U40 , R2238_U41 , R2238_U42 , R2238_U43;
wire R2238_U44 , R2238_U45 , R2238_U46 , R2238_U47 , R2238_U48 , R2238_U49 , R2238_U50 , R2238_U51 , R2238_U52 , R2238_U53;
wire R2238_U54 , R2238_U55 , R2238_U56 , R2238_U57 , R2238_U58 , R2238_U59 , R2238_U60 , R2238_U61 , R2238_U62 , R2238_U63;
wire R2238_U64 , R2238_U65 , R2238_U66 , SUB_450_U6 , SUB_450_U7 , SUB_450_U8 , SUB_450_U9 , SUB_450_U10 , SUB_450_U11 , SUB_450_U12;
wire SUB_450_U13 , SUB_450_U14 , SUB_450_U15 , SUB_450_U16 , SUB_450_U17 , SUB_450_U18 , SUB_450_U19 , SUB_450_U20 , SUB_450_U21 , SUB_450_U22;
wire SUB_450_U23 , SUB_450_U24 , SUB_450_U25 , SUB_450_U26 , SUB_450_U27 , SUB_450_U28 , SUB_450_U29 , SUB_450_U30 , SUB_450_U31 , SUB_450_U32;
wire SUB_450_U33 , SUB_450_U34 , SUB_450_U35 , SUB_450_U36 , SUB_450_U37 , SUB_450_U38 , SUB_450_U39 , SUB_450_U40 , SUB_450_U41 , SUB_450_U42;
wire SUB_450_U43 , SUB_450_U44 , SUB_450_U45 , SUB_450_U46 , SUB_450_U47 , SUB_450_U48 , SUB_450_U49 , SUB_450_U50 , SUB_450_U51 , SUB_450_U52;
wire SUB_450_U53 , SUB_450_U54 , SUB_450_U55 , SUB_450_U56 , SUB_450_U57 , SUB_450_U58 , SUB_450_U59 , SUB_450_U60 , SUB_450_U61 , SUB_450_U62;
wire SUB_450_U63 , SUB_450_U64 , SUB_450_U65 , SUB_450_U66 , ADD_371_U4 , ADD_371_U5 , ADD_371_U6 , ADD_371_U7 , ADD_371_U8 , ADD_371_U9;
wire ADD_371_U10 , ADD_371_U11 , ADD_371_U12 , ADD_371_U13 , ADD_371_U14 , ADD_371_U15 , ADD_371_U16 , ADD_371_U17 , ADD_371_U18 , ADD_371_U19;
wire ADD_371_U20 , ADD_371_U21 , ADD_371_U22 , ADD_371_U23 , ADD_371_U24 , ADD_371_U25 , ADD_371_U26 , ADD_371_U27 , ADD_371_U28 , ADD_371_U29;
wire ADD_371_U30 , ADD_371_U31 , ADD_371_U32 , ADD_371_U33 , ADD_371_U34 , ADD_371_U35 , ADD_371_U36 , ADD_371_U37 , ADD_371_U38 , ADD_371_U39;
wire ADD_371_U40 , ADD_371_U41 , ADD_371_U42 , ADD_371_U43 , ADD_371_U44 , ADD_405_U4 , ADD_405_U5 , ADD_405_U6 , ADD_405_U7 , ADD_405_U8;
wire ADD_405_U9 , ADD_405_U10 , ADD_405_U11 , ADD_405_U12 , ADD_405_U13 , ADD_405_U14 , ADD_405_U15 , ADD_405_U16 , ADD_405_U17 , ADD_405_U18;
wire ADD_405_U19 , ADD_405_U20 , ADD_405_U21 , ADD_405_U22 , ADD_405_U23 , ADD_405_U24 , ADD_405_U25 , ADD_405_U26 , ADD_405_U27 , ADD_405_U28;
wire ADD_405_U29 , ADD_405_U30 , ADD_405_U31 , ADD_405_U32 , ADD_405_U33 , ADD_405_U34 , ADD_405_U35 , ADD_405_U36 , ADD_405_U37 , ADD_405_U38;
wire ADD_405_U39 , ADD_405_U40 , ADD_405_U41 , ADD_405_U42 , ADD_405_U43 , ADD_405_U44 , ADD_405_U45 , ADD_405_U46 , ADD_405_U47 , ADD_405_U48;
wire ADD_405_U49 , ADD_405_U50 , ADD_405_U51 , ADD_405_U52 , ADD_405_U53 , ADD_405_U54 , ADD_405_U55 , ADD_405_U56 , ADD_405_U57 , ADD_405_U58;
wire ADD_405_U59 , ADD_405_U60 , ADD_405_U61 , ADD_405_U62 , ADD_405_U63 , ADD_405_U64 , ADD_405_U65 , ADD_405_U66 , ADD_405_U67 , ADD_405_U68;
wire ADD_405_U69 , ADD_405_U70 , ADD_405_U71 , ADD_405_U72 , ADD_405_U73 , ADD_405_U74 , ADD_405_U75 , ADD_405_U76 , ADD_405_U77 , ADD_405_U78;
wire ADD_405_U79 , ADD_405_U80 , ADD_405_U81 , ADD_405_U82 , ADD_405_U83 , ADD_405_U84 , ADD_405_U85 , ADD_405_U86 , ADD_405_U87 , ADD_405_U88;
wire ADD_405_U89 , ADD_405_U90 , ADD_405_U91 , ADD_405_U92 , ADD_405_U93 , ADD_405_U94 , ADD_405_U95 , ADD_405_U96 , ADD_405_U97 , ADD_405_U98;
wire ADD_405_U99 , ADD_405_U100 , ADD_405_U101 , ADD_405_U102 , ADD_405_U103 , ADD_405_U104 , ADD_405_U105 , ADD_405_U106 , ADD_405_U107 , ADD_405_U108;
wire ADD_405_U109 , ADD_405_U110 , ADD_405_U111 , ADD_405_U112 , ADD_405_U113 , ADD_405_U114 , ADD_405_U115 , ADD_405_U116 , ADD_405_U117 , ADD_405_U118;
wire ADD_405_U119 , ADD_405_U120 , ADD_405_U121 , ADD_405_U122 , ADD_405_U123 , ADD_405_U124 , ADD_405_U125 , ADD_405_U126 , ADD_405_U127 , ADD_405_U128;
wire ADD_405_U129 , ADD_405_U130 , ADD_405_U131 , ADD_405_U132 , ADD_405_U133 , ADD_405_U134 , ADD_405_U135 , ADD_405_U136 , ADD_405_U137 , ADD_405_U138;
wire ADD_405_U139 , ADD_405_U140 , ADD_405_U141 , ADD_405_U142 , ADD_405_U143 , ADD_405_U144 , ADD_405_U145 , ADD_405_U146 , ADD_405_U147 , ADD_405_U148;
wire ADD_405_U149 , ADD_405_U150 , ADD_405_U151 , ADD_405_U152 , ADD_405_U153 , ADD_405_U154 , ADD_405_U155 , ADD_405_U156 , ADD_405_U157 , ADD_405_U158;
wire ADD_405_U159 , ADD_405_U160 , ADD_405_U161 , ADD_405_U162 , ADD_405_U163 , ADD_405_U164 , ADD_405_U165 , ADD_405_U166 , ADD_405_U167 , ADD_405_U168;
wire ADD_405_U169 , ADD_405_U170 , ADD_405_U171 , ADD_405_U172 , ADD_405_U173 , ADD_405_U174 , ADD_405_U175 , ADD_405_U176 , ADD_405_U177 , ADD_405_U178;
wire ADD_405_U179 , ADD_405_U180 , ADD_405_U181 , ADD_405_U182 , ADD_405_U183 , ADD_405_U184 , ADD_405_U185 , ADD_405_U186 , GTE_485_U6 , GTE_485_U7;
wire ADD_515_U4 , ADD_515_U5 , ADD_515_U6 , ADD_515_U7 , ADD_515_U8 , ADD_515_U9 , ADD_515_U10 , ADD_515_U11 , ADD_515_U12 , ADD_515_U13;
wire ADD_515_U14 , ADD_515_U15 , ADD_515_U16 , ADD_515_U17 , ADD_515_U18 , ADD_515_U19 , ADD_515_U20 , ADD_515_U21 , ADD_515_U22 , ADD_515_U23;
wire ADD_515_U24 , ADD_515_U25 , ADD_515_U26 , ADD_515_U27 , ADD_515_U28 , ADD_515_U29 , ADD_515_U30 , ADD_515_U31 , ADD_515_U32 , ADD_515_U33;
wire ADD_515_U34 , ADD_515_U35 , ADD_515_U36 , ADD_515_U37 , ADD_515_U38 , ADD_515_U39 , ADD_515_U40 , ADD_515_U41 , ADD_515_U42 , ADD_515_U43;
wire ADD_515_U44 , ADD_515_U45 , ADD_515_U46 , ADD_515_U47 , ADD_515_U48 , ADD_515_U49 , ADD_515_U50 , ADD_515_U51 , ADD_515_U52 , ADD_515_U53;
wire ADD_515_U54 , ADD_515_U55 , ADD_515_U56 , ADD_515_U57 , ADD_515_U58 , ADD_515_U59 , ADD_515_U60 , ADD_515_U61 , ADD_515_U62 , ADD_515_U63;
wire ADD_515_U64 , ADD_515_U65 , ADD_515_U66 , ADD_515_U67 , ADD_515_U68 , ADD_515_U69 , ADD_515_U70 , ADD_515_U71 , ADD_515_U72 , ADD_515_U73;
wire ADD_515_U74 , ADD_515_U75 , ADD_515_U76 , ADD_515_U77 , ADD_515_U78 , ADD_515_U79 , ADD_515_U80 , ADD_515_U81 , ADD_515_U82 , ADD_515_U83;
wire ADD_515_U84 , ADD_515_U85 , ADD_515_U86 , ADD_515_U87 , ADD_515_U88 , ADD_515_U89 , ADD_515_U90 , ADD_515_U91 , ADD_515_U92 , ADD_515_U93;
wire ADD_515_U94 , ADD_515_U95 , ADD_515_U96 , ADD_515_U97 , ADD_515_U98 , ADD_515_U99 , ADD_515_U100 , ADD_515_U101 , ADD_515_U102 , ADD_515_U103;
wire ADD_515_U104 , ADD_515_U105 , ADD_515_U106 , ADD_515_U107 , ADD_515_U108 , ADD_515_U109 , ADD_515_U110 , ADD_515_U111 , ADD_515_U112 , ADD_515_U113;
wire ADD_515_U114 , ADD_515_U115 , ADD_515_U116 , ADD_515_U117 , ADD_515_U118 , ADD_515_U119 , ADD_515_U120 , ADD_515_U121 , ADD_515_U122 , ADD_515_U123;
wire ADD_515_U124 , ADD_515_U125 , ADD_515_U126 , ADD_515_U127 , ADD_515_U128 , ADD_515_U129 , ADD_515_U130 , ADD_515_U131 , ADD_515_U132 , ADD_515_U133;
wire ADD_515_U134 , ADD_515_U135 , ADD_515_U136 , ADD_515_U137 , ADD_515_U138 , ADD_515_U139 , ADD_515_U140 , ADD_515_U141 , ADD_515_U142 , ADD_515_U143;
wire ADD_515_U144 , ADD_515_U145 , ADD_515_U146 , ADD_515_U147 , ADD_515_U148 , ADD_515_U149 , ADD_515_U150 , ADD_515_U151;


nand NAND2_1 ( ADD_515_U182 , ADD_515_U101 , ADD_515_U21 );
nand NAND2_2 ( ADD_515_U181 , INSTADDRPOINTER_REG_10_ , ADD_515_U20 );
nand NAND2_3 ( ADD_515_U180 , ADD_515_U102 , ADD_515_U23 );
nor nor_4 ( U2352 , STATEBS16_REG , STATE2_REG_2_ );
and AND2_5 ( U2353 , U4219 , STATE2_REG_2_ );
and AND2_6 ( U2354 , U4253 , U4465 );
and AND2_7 ( U2355 , U3221 , U2450 );
and AND2_8 ( U2356 , R2238_U6 , U4180 );
and AND3_9 ( U2357 , U5947 , U3853 , R2167_U17 );
and AND2_10 ( U2358 , U2388 , U4212 );
and AND2_11 ( U2359 , STATE2_REG_2_ , U3418 );
and AND2_12 ( U2360 , STATE2_REG_2_ , U3401 );
and AND2_13 ( U2361 , U4212 , STATE2_REG_3_ );
and AND2_14 ( U2362 , U2359 , U4196 );
and AND2_15 ( U2363 , U2359 , U4198 );
and AND2_16 ( U2364 , U3852 , U3403 );
and AND2_17 ( U2365 , U4249 , U3403 );
and AND3_18 ( U2366 , U3418 , STATE2_REG_1_ , U3417 );
and AND3_19 ( U2367 , STATE2_REG_1_ , U3418 , R2337_U58 );
and AND2_20 ( U2368 , U4223 , STATE2_REG_0_ );
and AND2_21 ( U2369 , U2362 , U4485 );
and AND2_22 ( U2370 , U3401 , U3250 );
and AND2_23 ( U2371 , U4210 , U4437 );
and AND2_24 ( U2372 , STATE2_REG_0_ , U3403 );
and AND2_25 ( U2373 , STATE2_REG_3_ , U3418 );
and AND2_26 ( U2374 , U2360 , U4202 );
and AND2_27 ( U2375 , U2360 , U4204 );
and AND2_28 ( U2376 , U5786 , U3403 );
and AND2_29 ( U2377 , U3750 , U3401 );
and AND2_30 ( U2378 , U2360 , U5557 );
and AND2_31 ( U2379 , U2363 , U3267 );
and AND2_32 ( U2380 , U2360 , U7596 );
and AND2_33 ( U2381 , U2357 , U3258 );
and AND2_34 ( U2382 , U2357 , U4465 );
and AND2_35 ( U2383 , U4210 , U3378 );
and AND2_36 ( U2384 , STATE2_REG_0_ , U3404 );
and AND2_37 ( U2385 , U3404 , U3281 );
and AND2_38 ( U2386 , U4211 , U3410 );
and AND2_39 ( U2387 , U3872 , U4211 );
and AND2_40 ( U2388 , STATEBS16_REG , U4197 );
and AND2_41 ( U2389 , U2452 , U7482 );
and AND2_42 ( U2390 , DATAI_0_ , U4212 );
and AND2_43 ( U2391 , DATAI_1_ , U4212 );
and AND2_44 ( U2392 , DATAI_2_ , U4212 );
and AND2_45 ( U2393 , DATAI_3_ , U4212 );
and AND2_46 ( U2394 , DATAI_4_ , U4212 );
and AND2_47 ( U2395 , DATAI_5_ , U4212 );
and AND2_48 ( U2396 , DATAI_6_ , U4212 );
and AND2_49 ( U2397 , DATAI_7_ , U4212 );
and AND2_50 ( U2398 , DATAI_24_ , U2358 );
and AND2_51 ( U2399 , DATAI_16_ , U2358 );
and AND2_52 ( U2400 , DATAI_25_ , U2358 );
and AND2_53 ( U2401 , DATAI_17_ , U2358 );
and AND2_54 ( U2402 , DATAI_26_ , U2358 );
and AND2_55 ( U2403 , DATAI_18_ , U2358 );
and AND2_56 ( U2404 , DATAI_27_ , U2358 );
and AND2_57 ( U2405 , DATAI_19_ , U2358 );
and AND2_58 ( U2406 , DATAI_28_ , U2358 );
and AND2_59 ( U2407 , DATAI_20_ , U2358 );
and AND2_60 ( U2408 , DATAI_29_ , U2358 );
and AND2_61 ( U2409 , DATAI_21_ , U2358 );
and AND2_62 ( U2410 , DATAI_30_ , U2358 );
and AND2_63 ( U2411 , DATAI_22_ , U2358 );
and AND2_64 ( U2412 , DATAI_31_ , U2358 );
and AND2_65 ( U2413 , DATAI_23_ , U2358 );
and AND2_66 ( U2414 , U2361 , U3258 );
and AND2_67 ( U2415 , U2361 , U3378 );
and AND2_68 ( U2416 , U2361 , U3264 );
and AND2_69 ( U2417 , U2361 , U3271 );
and AND2_70 ( U2418 , U2361 , U3270 );
and AND2_71 ( U2419 , U2361 , U3265 );
and AND2_72 ( U2420 , U2361 , U4161 );
and AND2_73 ( U2421 , U2361 , U4159 );
and AND2_74 ( U2422 , U4211 , U5449 );
and AND2_75 ( U2423 , U4211 , U4219 );
and AND2_76 ( U2424 , U2384 , U3271 );
and AND2_77 ( U2425 , U2368 , U2448 );
and AND2_78 ( U2426 , U3877 , U3418 );
nor nor_79 ( U2427 , STATE2_REG_1_ , STATE2_REG_3_ );
and AND2_80 ( U2428 , STATE2_REG_2_ , STATE2_REG_1_ );
and AND2_81 ( U2429 , U6354 , U3418 );
and AND2_82 ( U2430 , STATE2_REG_1_ , U3374 );
and AND2_83 ( U2431 , U4187 , U7482 );
and AND2_84 ( U2432 , U3442 , U3347 );
and AND2_85 ( U2433 , U4528 , U3442 );
and AND2_86 ( U2434 , U7684 , U3347 );
and AND2_87 ( U2435 , U4528 , U7684 );
and AND2_88 ( U2436 , U3222 , U3288 );
and AND2_89 ( U2437 , U4531 , U3288 );
and AND2_90 ( U2438 , R2182_U42 , R2182_U25 );
and AND2_91 ( U2439 , R2182_U42 , U3303 );
and AND2_92 ( U2440 , R2182_U25 , U3304 );
nor nor_93 ( U2441 , R2182_U42 , R2182_U25 );
and AND2_94 ( U2442 , R2182_U33 , R2182_U34 );
and AND2_95 ( U2443 , R2182_U33 , U3305 );
and AND2_96 ( U2444 , R2182_U34 , U3306 );
nor nor_97 ( U2445 , R2182_U33 , R2182_U34 );
and AND2_98 ( U2446 , STATE2_REG_1_ , U3458 );
and AND2_99 ( U2447 , U3565 , U2452 );
and AND2_100 ( U2448 , R2167_U17 , U3271 );
and AND2_101 ( U2449 , U4482 , U3258 );
and AND2_102 ( U2450 , STATE2_REG_0_ , U4388 );
and AND2_103 ( U2451 , U4239 , STATE2_REG_0_ );
and AND4_104 ( U2452 , U4388 , U3264 , U3378 , U4161 );
and AND4_105 ( U2453 , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ );
and AND2_106 ( U2454 , INSTQUEUERD_ADDR_REG_1_ , U3253 );
and AND4_107 ( U2455 , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ , U3253 );
and AND2_108 ( U2456 , INSTQUEUERD_ADDR_REG_0_ , U3252 );
and AND4_109 ( U2457 , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_2_ , U3252 );
and AND2_110 ( U2458 , U3495 , U4366 );
and AND4_111 ( U2459 , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ , U3251 );
and AND3_112 ( U2460 , U3251 , U3253 , INSTQUEUERD_ADDR_REG_1_ );
and AND2_113 ( U2461 , U3494 , U3493 );
and AND3_114 ( U2462 , U3251 , U3252 , INSTQUEUERD_ADDR_REG_0_ );
and AND2_115 ( U2463 , U3492 , U3491 );
and AND2_116 ( U2464 , INSTQUEUERD_ADDR_REG_3_ , U4368 );
and AND2_117 ( U2465 , U3490 , U3489 );
and AND2_118 ( U2466 , U3488 , U3487 );
and AND3_119 ( U2467 , INSTQUEUERD_ADDR_REG_2_ , U3257 , U4366 );
and AND2_120 ( U2468 , U3486 , U3485 );
nor nor_121 ( U2469 , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_2_ );
and AND3_122 ( U2470 , INSTQUEUERD_ADDR_REG_1_ , U3253 , U2469 );
and AND3_123 ( U2471 , INSTQUEUERD_ADDR_REG_0_ , U3252 , U2469 );
and AND2_124 ( U2472 , U4368 , U3257 );
and AND3_125 ( U2473 , U7668 , U7667 , U3393 );
and AND2_126 ( U2474 , R2144_U49 , U3299 );
and AND2_127 ( U2475 , U3441 , U3345 );
and AND2_128 ( U2476 , R2144_U8 , R2144_U49 );
and AND2_129 ( U2477 , U4516 , U2476 );
and AND2_130 ( U2478 , INSTQUEUEWR_ADDR_REG_2_ , INSTQUEUEWR_ADDR_REG_3_ );
and AND2_131 ( U2479 , INSTQUEUEWR_ADDR_REG_2_ , U3290 );
and AND2_132 ( U2480 , U3302 , U4536 );
and AND2_133 ( U2481 , U4512 , U2476 );
and AND2_134 ( U2482 , U3314 , U4594 );
and AND2_135 ( U2483 , U4513 , U2476 );
and AND2_136 ( U2484 , U3321 , U4653 );
and AND2_137 ( U2485 , U4514 , R2144_U43 );
nor nor_138 ( U2486 , R2144_U43 , R2144_U50 );
and AND2_139 ( U2487 , U2486 , U2476 );
nor nor_140 ( U2488 , INSTQUEUEWR_ADDR_REG_0_ , INSTQUEUEWR_ADDR_REG_1_ );
and AND2_141 ( U2489 , U3325 , U4710 );
and AND2_142 ( U2490 , U7681 , U3345 );
and AND2_143 ( U2491 , U4517 , U4516 );
and AND2_144 ( U2492 , U3330 , U4768 );
and AND2_145 ( U2493 , U4517 , U4512 );
and AND2_146 ( U2494 , U3334 , U4825 );
and AND2_147 ( U2495 , U4517 , U4513 );
and AND2_148 ( U2496 , U3337 , U4883 );
and AND2_149 ( U2497 , U4517 , U2486 );
and AND2_150 ( U2498 , U3341 , U4940 );
and AND2_151 ( U2499 , U4519 , U3441 );
and AND2_152 ( U2500 , U3346 , U3344 );
and AND2_153 ( U2501 , U4512 , U2474 );
and AND2_154 ( U2502 , U3351 , U5053 );
and AND2_155 ( U2503 , U4513 , U2474 );
and AND2_156 ( U2504 , U3354 , U5111 );
and AND2_157 ( U2505 , U2486 , U2474 );
and AND2_158 ( U2506 , U3358 , U5168 );
and AND2_159 ( U2507 , U4519 , U7681 );
nor nor_160 ( U2508 , R2144_U49 , R2144_U8 );
and AND2_161 ( U2509 , U2508 , U4516 );
nor nor_162 ( U2510 , INSTQUEUEWR_ADDR_REG_3_ , INSTQUEUEWR_ADDR_REG_2_ );
and AND2_163 ( U2511 , U3361 , U5226 );
and AND2_164 ( U2512 , U2508 , U4512 );
and AND2_165 ( U2513 , U3365 , U5283 );
and AND2_166 ( U2514 , U2508 , U4513 );
and AND2_167 ( U2515 , U3368 , U5341 );
and AND2_168 ( U2516 , U2508 , U2486 );
and AND2_169 ( U2517 , U3372 , U5398 );
and AND3_170 ( U2518 , U7688 , U7687 , U5456 );
and AND2_171 ( U2519 , U3732 , U5487 );
and AND2_172 ( U2520 , U4207 , U3433 );
and AND2_173 ( U2521 , INSTQUEUERD_ADDR_REG_0_ , U3389 );
and AND2_174 ( U2522 , U5471 , U5499 );
and AND2_175 ( U2523 , U2522 , U2521 );
and AND2_176 ( U2524 , U3253 , U3389 );
and AND2_177 ( U2525 , U2522 , U2524 );
and AND2_178 ( U2526 , U5507 , INSTQUEUERD_ADDR_REG_0_ );
and AND2_179 ( U2527 , U2522 , U2526 );
and AND2_180 ( U2528 , U5507 , U3253 );
and AND2_181 ( U2529 , U2522 , U2528 );
and AND2_182 ( U2530 , U5471 , U3388 );
and AND2_183 ( U2531 , U2530 , U2521 );
and AND2_184 ( U2532 , U2530 , U2524 );
and AND2_185 ( U2533 , U2530 , U2526 );
and AND2_186 ( U2534 , U2530 , U2528 );
and AND2_187 ( U2535 , U5499 , U3425 );
and AND2_188 ( U2536 , U2535 , U2521 );
and AND2_189 ( U2537 , U2535 , U2524 );
and AND2_190 ( U2538 , U2535 , U2526 );
and AND2_191 ( U2539 , U2535 , U2528 );
and AND2_192 ( U2540 , U3425 , U3388 );
and AND2_193 ( U2541 , U2521 , U2540 );
and AND2_194 ( U2542 , U2524 , U2540 );
and AND2_195 ( U2543 , U2526 , U2540 );
and AND2_196 ( U2544 , U2528 , U2540 );
and AND2_197 ( U2545 , U5468 , U7708 );
and AND2_198 ( U2546 , U2545 , U2454 );
and AND2_199 ( U2547 , U2545 , U3486 );
and AND2_200 ( U2548 , U2545 , U4366 );
and AND2_201 ( U2549 , U2545 , U2456 );
and AND2_202 ( U2550 , U5468 , U3443 );
and AND2_203 ( U2551 , U2550 , U2454 );
and AND2_204 ( U2552 , U2550 , U3486 );
and AND2_205 ( U2553 , U2550 , U4366 );
and AND2_206 ( U2554 , U2550 , U2456 );
and AND2_207 ( U2555 , U7708 , U3429 );
and AND2_208 ( U2556 , U2555 , U2454 );
and AND2_209 ( U2557 , U2555 , U3486 );
and AND2_210 ( U2558 , U2555 , U4366 );
and AND2_211 ( U2559 , U2555 , U2456 );
and AND2_212 ( U2560 , U3443 , U3429 );
and AND2_213 ( U2561 , U2560 , U2454 );
and AND2_214 ( U2562 , U2560 , U3486 );
and AND2_215 ( U2563 , U2560 , U4366 );
and AND2_216 ( U2564 , U2560 , U2456 );
and AND2_217 ( U2565 , U7053 , U4367 );
and AND2_218 ( U2566 , U7053 , U2460 );
and AND2_219 ( U2567 , U7053 , U2462 );
and AND2_220 ( U2568 , U7053 , U4368 );
and AND2_221 ( U2569 , U7053 , INSTQUEUERD_ADDR_REG_2_ );
and AND2_222 ( U2570 , U2569 , U3486 );
and AND2_223 ( U2571 , U2569 , U2454 );
and AND2_224 ( U2572 , U2569 , U2456 );
and AND2_225 ( U2573 , U2569 , U4366 );
and AND2_226 ( U2574 , U4367 , U3432 );
and AND2_227 ( U2575 , U2460 , U3432 );
and AND2_228 ( U2576 , U2462 , U3432 );
and AND2_229 ( U2577 , U4368 , U3432 );
and AND2_230 ( U2578 , INSTQUEUERD_ADDR_REG_2_ , U3432 );
and AND2_231 ( U2579 , U2578 , U3486 );
and AND2_232 ( U2580 , U2578 , U2454 );
and AND2_233 ( U2581 , U2578 , U2456 );
and AND2_234 ( U2582 , U2578 , U4366 );
and AND2_235 ( U2583 , U7778 , U4172 );
and AND2_236 ( U2584 , U2583 , U2524 );
and AND2_237 ( U2585 , U2583 , U2521 );
and AND2_238 ( U2586 , U2583 , U2528 );
and AND2_239 ( U2587 , U2583 , U2526 );
and AND2_240 ( U2588 , U7778 , U3439 );
and AND2_241 ( U2589 , U2588 , U2524 );
and AND2_242 ( U2590 , U2588 , U2521 );
and AND2_243 ( U2591 , U2588 , U2528 );
and AND2_244 ( U2592 , U2588 , U2526 );
and AND2_245 ( U2593 , U4172 , U3444 );
and AND2_246 ( U2594 , U2593 , U2524 );
and AND2_247 ( U2595 , U2593 , U2521 );
and AND2_248 ( U2596 , U2593 , U2528 );
and AND2_249 ( U2597 , U2593 , U2526 );
and AND2_250 ( U2598 , U3444 , U3439 );
and AND2_251 ( U2599 , U2598 , U2524 );
and AND2_252 ( U2600 , U2598 , U2521 );
and AND2_253 ( U2601 , U2598 , U2528 );
and AND2_254 ( U2602 , U2598 , U2526 );
and AND2_255 ( U2603 , STATE2_REG_0_ , U3376 );
and AND2_256 ( U2604 , EBX_REG_31_ , U2379 );
and AND5_257 ( U2605 , U3521 , U2607 , U3520 , U3519 , U3518 );
and AND2_258 ( U2606 , U7492 , U3414 );
and AND2_259 ( U2607 , U7660 , U7659 );
and AND2_260 ( U2608 , U7775 , U7774 );
nand NAND2_261 ( U2609 , U6744 , U3993 );
nand NAND2_262 ( U2610 , U6741 , U3992 );
nand NAND2_263 ( U2611 , U6738 , U3991 );
nand NAND2_264 ( U2612 , U6735 , U3990 );
nand NAND2_265 ( U2613 , U6844 , U4014 );
nand NAND3_266 ( U2614 , U6841 , U6842 , U6843 );
nand NAND3_267 ( U2615 , U6838 , U6839 , U6840 );
nand NAND3_268 ( U2616 , U6835 , U6836 , U6837 );
nand NAND3_269 ( U2617 , U6832 , U6833 , U6834 );
nand NAND3_270 ( U2618 , U6829 , U6830 , U6831 );
nand NAND2_271 ( ADD_515_U179 , INSTADDRPOINTER_REG_11_ , ADD_515_U22 );
and AND2_272 ( U2620 , R2144_U145 , U6734 );
and AND2_273 ( U2621 , R2144_U145 , U6734 );
and AND2_274 ( U2622 , R2144_U145 , U6734 );
and AND2_275 ( U2623 , R2144_U145 , U6734 );
and AND2_276 ( U2624 , R2144_U145 , U6734 );
and AND2_277 ( U2625 , R2144_U145 , U6734 );
and AND2_278 ( U2626 , R2144_U145 , U6734 );
and AND2_279 ( U2627 , R2144_U145 , U6734 );
and AND2_280 ( U2628 , R2144_U145 , U6734 );
and AND2_281 ( U2629 , R2144_U145 , U6734 );
and AND2_282 ( U2630 , R2144_U145 , U6734 );
and AND2_283 ( U2631 , R2144_U145 , U6734 );
and AND2_284 ( U2632 , R2144_U145 , U6734 );
and AND2_285 ( U2633 , R2144_U145 , U6734 );
and AND2_286 ( U2634 , R2144_U11 , U6734 );
and AND2_287 ( U2635 , R2144_U37 , U6734 );
and AND2_288 ( U2636 , R2144_U38 , U6734 );
and AND2_289 ( U2637 , R2144_U39 , U6734 );
and AND2_290 ( U2638 , R2144_U40 , U6734 );
and AND2_291 ( U2639 , R2144_U41 , U6734 );
and AND2_292 ( U2640 , R2144_U42 , U6734 );
and AND2_293 ( U2641 , R2144_U30 , U6734 );
and AND2_294 ( U2642 , R2144_U80 , U6734 );
and AND2_295 ( U2643 , R2144_U10 , U6734 );
and AND2_296 ( U2644 , R2144_U9 , U6734 );
and AND2_297 ( U2645 , R2144_U45 , U6734 );
and AND2_298 ( U2646 , R2144_U47 , U6734 );
and AND2_299 ( U2647 , R2144_U8 , U6734 );
nand NAND2_300 ( U2648 , U3427 , U6857 );
and AND2_301 ( U2649 , R2144_U50 , U6734 );
and AND2_302 ( U2650 , STATE2_REG_2_ , U6858 );
nand NAND3_303 ( U2651 , U6757 , U6756 , U6758 );
nand NAND2_304 ( U2652 , U6759 , U3997 );
nand NAND2_305 ( U2653 , U6768 , U3999 );
nand NAND2_306 ( U2654 , U6772 , U4000 );
nand NAND2_307 ( U2655 , U6776 , U4001 );
nand NAND2_308 ( U2656 , U6780 , U4002 );
nand NAND2_309 ( U2657 , U6784 , U4003 );
nand NAND2_310 ( U2658 , U6788 , U4004 );
nand NAND2_311 ( U2659 , U6792 , U4005 );
nand NAND2_312 ( U2660 , U6796 , U4006 );
nand NAND2_313 ( U2661 , U6800 , U4007 );
nand NAND2_314 ( U2662 , U6804 , U4008 );
nand NAND2_315 ( U2663 , U6813 , U4010 );
nand NAND2_316 ( U2664 , U6817 , U4011 );
nand NAND2_317 ( U2665 , U6821 , U4012 );
nand NAND2_318 ( U2666 , U6825 , U4013 );
nand NAND2_319 ( U2667 , U6747 , U3994 );
nand NAND4_320 ( U2668 , U6755 , U6754 , U3996 , U6751 );
nand NAND4_321 ( U2669 , U6767 , U6766 , U3998 , U6763 );
nand NAND4_322 ( U2670 , U6812 , U6811 , U4009 , U6808 );
nand NAND4_323 ( U2671 , U6851 , U6850 , U4015 , U6847 );
nand NAND5_324 ( U2672 , U6854 , U6852 , U6853 , U6856 , U6855 );
nand NAND2_325 ( U2673 , U7446 , U7445 );
nand NAND2_326 ( U2674 , U7448 , U7447 );
nand NAND2_327 ( U2675 , U4156 , U7451 );
nand NAND2_328 ( U2676 , U4157 , U7454 );
nand NAND3_329 ( U2677 , U7782 , U7781 , U7455 );
nand NAND2_330 ( U2678 , U7444 , U3271 );
nand NAND2_331 ( U2679 , U7393 , U7392 );
nand NAND2_332 ( U2680 , U7395 , U7394 );
nand NAND2_333 ( U2681 , U7399 , U7398 );
nand NAND2_334 ( U2682 , U7401 , U7400 );
nand NAND2_335 ( U2683 , U7403 , U7402 );
nand NAND2_336 ( U2684 , U7405 , U7404 );
nand NAND2_337 ( U2685 , U7407 , U7406 );
nand NAND2_338 ( U2686 , U7409 , U7408 );
nand NAND2_339 ( U2687 , U7411 , U7410 );
nand NAND2_340 ( U2688 , U7413 , U7412 );
nand NAND2_341 ( U2689 , U7415 , U7414 );
nand NAND2_342 ( U2690 , U7417 , U7416 );
nand NAND2_343 ( U2691 , U7421 , U7420 );
nand NAND2_344 ( U2692 , U7423 , U7422 );
nand NAND2_345 ( U2693 , U7425 , U7424 );
nand NAND2_346 ( U2694 , U7427 , U7426 );
nand NAND2_347 ( U2695 , U7429 , U7428 );
nand NAND2_348 ( U2696 , U7431 , U7430 );
nand NAND2_349 ( U2697 , U7433 , U7432 );
nand NAND2_350 ( U2698 , U7435 , U7434 );
nand NAND2_351 ( U2699 , U7437 , U7436 );
nand NAND2_352 ( U2700 , U7439 , U7438 );
nand NAND2_353 ( U2701 , U7381 , U7380 );
nand NAND2_354 ( U2702 , U7383 , U7382 );
nand NAND2_355 ( U2703 , U7385 , U7384 );
nand NAND2_356 ( U2704 , U7387 , U7386 );
nand NAND2_357 ( U2705 , U7389 , U7388 );
nand NAND2_358 ( U2706 , U7391 , U7390 );
nand NAND2_359 ( U2707 , U7397 , U7396 );
nand NAND2_360 ( U2708 , U7419 , U7418 );
nand NAND2_361 ( U2709 , U7441 , U7440 );
nand NAND2_362 ( U2710 , U7443 , U7442 );
nand NAND2_363 ( U2711 , U7365 , U7364 );
nand NAND2_364 ( U2712 , U7367 , U7366 );
nand NAND2_365 ( U2713 , U4153 , U4227 );
nand NAND4_366 ( U2714 , U7374 , U7373 , U4154 , U3421 );
nand NAND2_367 ( U2715 , U4227 , U4155 );
nand NAND2_368 ( U2716 , U7353 , U7352 );
nand NAND2_369 ( U2717 , U7355 , U7354 );
nand NAND2_370 ( U2718 , U4149 , U7356 );
nand NAND2_371 ( U2719 , U4150 , U7358 );
nand NAND2_372 ( U2720 , U4151 , U7360 );
nand NAND2_373 ( U2721 , U4152 , U7362 );
nand NAND2_374 ( U2722 , U4147 , U4180 );
and AND2_375 ( U2723 , U7224 , U7071 );
and AND2_376 ( U2724 , U7241 , U7071 );
and AND2_377 ( U2725 , U7258 , U7071 );
and AND2_378 ( U2726 , U7608 , U7071 );
and AND2_379 ( U2727 , U7290 , U7071 );
and AND2_380 ( U2728 , U7307 , U7071 );
and AND2_381 ( U2729 , U7324 , U7071 );
and AND2_382 ( U2730 , U7341 , U7071 );
nand NAND2_383 ( U2731 , U2606 , U7342 );
and AND2_384 ( U2732 , U7071 , U7070 );
and AND2_385 ( U2733 , U7102 , U7071 );
and AND2_386 ( U2734 , U7119 , U7071 );
and AND2_387 ( U2735 , U7606 , U7071 );
and AND2_388 ( U2736 , U7151 , U7071 );
and AND2_389 ( U2737 , U7168 , U7071 );
and AND2_390 ( U2738 , U7185 , U7071 );
and AND2_391 ( U2739 , U7202 , U7071 );
and AND2_392 ( U2740 , INSTQUEUERD_ADDR_REG_4_ , U7051 );
nand NAND2_393 ( U2741 , U4066 , U7084 );
and AND2_394 ( U2742 , U7480 , U7479 );
and AND2_395 ( U2743 , U7494 , U7458 );
and AND2_396 ( U2744 , U7467 , U7466 );
nand NAND2_397 ( U2745 , U7036 , U7035 );
nand NAND2_398 ( U2746 , U7038 , U7037 );
nand NAND2_399 ( U2747 , U7040 , U7039 );
nand NAND2_400 ( U2748 , U7604 , U7041 );
nand NAND2_401 ( U2749 , U7043 , U7042 );
nand NAND2_402 ( U2750 , U7045 , U7044 );
nand NAND2_403 ( U2751 , U4049 , U7046 );
nand NAND3_404 ( U2752 , U4050 , U7048 , U7049 );
and AND2_405 ( U2753 , U6945 , U6897 );
and AND2_406 ( U2754 , U6962 , U6897 );
and AND2_407 ( U2755 , U6979 , U6897 );
and AND2_408 ( U2756 , U7603 , U6897 );
and AND2_409 ( U2757 , U7011 , U6897 );
and AND2_410 ( U2758 , U7028 , U6897 );
and AND2_411 ( U2759 , U6897 , U6896 );
and AND2_412 ( U2760 , U6914 , U6897 );
nand NAND2_413 ( U2761 , U6916 , U6915 );
nand NAND2_414 ( U2762 , U6918 , U6917 );
nand NAND2_415 ( U2763 , U6920 , U6919 );
nand NAND2_416 ( U2764 , U6922 , U6921 );
nand NAND3_417 ( U2765 , U6924 , U6923 , U6925 );
nand NAND3_418 ( U2766 , U6927 , U6926 , U6928 );
nand NAND3_419 ( U2767 , U7031 , U7029 , U7030 );
nand NAND3_420 ( U2768 , U7034 , U7032 , U7033 );
and AND2_421 ( U2769 , R2144_U145 , U4147 );
and AND2_422 ( U2770 , U4147 , R2144_U145 );
and AND2_423 ( U2771 , U4147 , R2144_U11 );
and AND2_424 ( U2772 , U4147 , R2144_U37 );
and AND2_425 ( U2773 , U4147 , R2144_U38 );
and AND2_426 ( U2774 , U4147 , R2144_U39 );
and AND2_427 ( U2775 , U4147 , R2144_U40 );
and AND2_428 ( U2776 , U4147 , R2144_U41 );
and AND2_429 ( U2777 , U4147 , R2144_U42 );
and AND2_430 ( U2778 , U4147 , R2144_U30 );
nand NAND2_431 ( U2779 , U6860 , U6859 );
nand NAND2_432 ( U2780 , U6862 , U6861 );
nand NAND2_433 ( U2781 , U6864 , U6863 );
nand NAND2_434 ( U2782 , U6866 , U6865 );
nand NAND2_435 ( U2783 , U6868 , U6867 );
nand NAND2_436 ( U2784 , U6870 , U6869 );
nand NAND3_437 ( U2785 , U6872 , U6873 , U6871 );
nand NAND3_438 ( U2786 , U4016 , U6875 , U6874 );
nand NAND3_439 ( U2787 , U6878 , U6879 , U6877 );
nand NAND3_440 ( U2788 , U6605 , U3419 , U7486 );
nand NAND2_441 ( U2789 , U7638 , U6601 );
nand NAND2_442 ( U2790 , U6600 , U6599 );
nand NAND3_443 ( U2791 , U7757 , U7756 , U4231 );
nand NAND3_444 ( U2792 , U7753 , U7752 , U4231 );
nand NAND2_445 ( U2793 , U6589 , U4236 );
nand NAND3_446 ( U2794 , U7745 , U7744 , U4228 );
nand NAND3_447 ( U2795 , U7735 , U7734 , U4228 );
nand NAND5_448 ( U2796 , U6581 , U3936 , U3937 , U6579 , U6583 );
nand NAND5_449 ( U2797 , U6574 , U3934 , U3935 , U6572 , U6576 );
nand NAND5_450 ( U2798 , U6567 , U3932 , U3933 , U6565 , U6569 );
nand NAND5_451 ( U2799 , U6560 , U3930 , U3931 , U6558 , U6562 );
nand NAND5_452 ( U2800 , U6553 , U3928 , U3929 , U6551 , U6555 );
nand NAND5_453 ( U2801 , U6546 , U3926 , U3927 , U6544 , U6548 );
nand NAND5_454 ( U2802 , U6539 , U3924 , U3925 , U6537 , U6541 );
nand NAND5_455 ( U2803 , U6532 , U3922 , U3923 , U6530 , U6534 );
nand NAND5_456 ( U2804 , U6525 , U3920 , U3921 , U6523 , U6527 );
nand NAND5_457 ( U2805 , U6518 , U3918 , U3919 , U6516 , U6520 );
nand NAND5_458 ( U2806 , U6511 , U3916 , U3917 , U6509 , U6513 );
nand NAND5_459 ( U2807 , U6504 , U3914 , U3915 , U6502 , U6506 );
nand NAND5_460 ( U2808 , U3912 , U6497 , U3913 , U6495 , U6499 );
nand NAND5_461 ( U2809 , U3910 , U6490 , U3911 , U6488 , U6492 );
nand NAND5_462 ( U2810 , U3908 , U6483 , U3909 , U6481 , U6485 );
nand NAND5_463 ( U2811 , U6476 , U6475 , U3907 , U3906 , U6478 );
nand NAND5_464 ( U2812 , U6469 , U6468 , U3905 , U3904 , U6471 );
nand NAND5_465 ( U2813 , U3903 , U6462 , U3902 , U6461 , U6464 );
nand NAND5_466 ( U2814 , U3901 , U6455 , U3900 , U6454 , U6457 );
nand NAND5_467 ( U2815 , U3899 , U6448 , U3898 , U6447 , U6450 );
nand NAND5_468 ( U2816 , U3897 , U6441 , U3896 , U6440 , U6443 );
nand NAND5_469 ( U2817 , U3895 , U6434 , U3894 , U6433 , U6436 );
nand NAND5_470 ( U2818 , U3893 , U6427 , U3892 , U6426 , U6429 );
nand NAND5_471 ( U2819 , U3891 , U6420 , U3890 , U6419 , U6422 );
nand NAND5_472 ( U2820 , U3889 , U6413 , U3888 , U6412 , U6415 );
nand NAND5_473 ( U2821 , U3887 , U6406 , U3886 , U6405 , U6408 );
nand NAND4_474 ( U2822 , U3884 , U6397 , U6398 , U3885 );
nand NAND5_475 ( U2823 , U3882 , U6389 , U3883 , U6391 , U6390 );
nand NAND4_476 ( U2824 , U6381 , U6380 , U6382 , U3881 );
nand NAND4_477 ( U2825 , U6373 , U6372 , U6374 , U3880 );
nand NAND4_478 ( U2826 , U6365 , U6364 , U6366 , U3879 );
nand NAND4_479 ( U2827 , U6357 , U6356 , U6358 , U3878 );
nand NAND2_480 ( U2828 , U6347 , U6346 );
nand NAND3_481 ( U2829 , U6344 , U6345 , U6343 );
nand NAND3_482 ( U2830 , U6341 , U6342 , U6340 );
nand NAND3_483 ( U2831 , U6338 , U6339 , U6337 );
nand NAND3_484 ( U2832 , U6335 , U6336 , U6334 );
nand NAND3_485 ( U2833 , U6332 , U6333 , U6331 );
nand NAND3_486 ( U2834 , U6329 , U6330 , U6328 );
nand NAND3_487 ( U2835 , U6326 , U6327 , U6325 );
nand NAND3_488 ( U2836 , U6323 , U6324 , U6322 );
nand NAND3_489 ( U2837 , U6320 , U6321 , U6319 );
nand NAND3_490 ( U2838 , U6317 , U6318 , U6316 );
nand NAND3_491 ( U2839 , U6314 , U6315 , U6313 );
nand NAND3_492 ( U2840 , U6311 , U6312 , U6310 );
nand NAND3_493 ( U2841 , U6308 , U6309 , U6307 );
nand NAND3_494 ( U2842 , U6305 , U6306 , U6304 );
nand NAND3_495 ( U2843 , U6302 , U6303 , U6301 );
nand NAND3_496 ( U2844 , U6299 , U6300 , U6298 );
nand NAND3_497 ( U2845 , U6296 , U6297 , U6295 );
nand NAND3_498 ( U2846 , U6293 , U6294 , U6292 );
nand NAND3_499 ( U2847 , U6290 , U6291 , U6289 );
nand NAND3_500 ( U2848 , U6287 , U6288 , U6286 );
nand NAND3_501 ( U2849 , U6284 , U6285 , U6283 );
nand NAND3_502 ( U2850 , U6281 , U6282 , U6280 );
nand NAND3_503 ( U2851 , U6278 , U6279 , U6277 );
nand NAND3_504 ( U2852 , U6275 , U6276 , U6274 );
nand NAND3_505 ( U2853 , U6272 , U6273 , U6271 );
nand NAND3_506 ( U2854 , U6269 , U6270 , U6268 );
nand NAND3_507 ( U2855 , U6266 , U6267 , U6265 );
nand NAND3_508 ( U2856 , U6263 , U6264 , U6262 );
nand NAND3_509 ( U2857 , U6260 , U6261 , U6259 );
nand NAND3_510 ( U2858 , U6257 , U6258 , U6256 );
nand NAND3_511 ( U2859 , U6254 , U6253 , U6255 );
nand NAND2_512 ( U2860 , U4164 , U6250 );
nand NAND4_513 ( U2861 , U6247 , U6246 , U6249 , U6248 );
nand NAND4_514 ( U2862 , U6243 , U6242 , U6245 , U6244 );
nand NAND4_515 ( U2863 , U6239 , U6238 , U6241 , U6240 );
nand NAND4_516 ( U2864 , U6235 , U6234 , U6237 , U6236 );
nand NAND4_517 ( U2865 , U6231 , U6230 , U6233 , U6232 );
nand NAND4_518 ( U2866 , U6227 , U6226 , U6229 , U6228 );
nand NAND4_519 ( U2867 , U6223 , U6222 , U6225 , U6224 );
nand NAND4_520 ( U2868 , U6219 , U6218 , U6221 , U6220 );
nand NAND4_521 ( U2869 , U6215 , U6214 , U6217 , U6216 );
nand NAND4_522 ( U2870 , U6211 , U6210 , U6213 , U6212 );
nand NAND4_523 ( U2871 , U6207 , U6206 , U6209 , U6208 );
nand NAND4_524 ( U2872 , U6203 , U6202 , U6205 , U6204 );
nand NAND4_525 ( U2873 , U6199 , U6198 , U6201 , U6200 );
nand NAND4_526 ( U2874 , U6195 , U6194 , U6197 , U6196 );
nand NAND4_527 ( U2875 , U6191 , U6190 , U6193 , U6192 );
nand NAND3_528 ( U2876 , U6189 , U6187 , U6188 );
nand NAND3_529 ( U2877 , U6186 , U6184 , U6185 );
nand NAND3_530 ( U2878 , U6183 , U6181 , U6182 );
nand NAND3_531 ( U2879 , U6180 , U6178 , U6179 );
nand NAND3_532 ( U2880 , U6177 , U6175 , U6176 );
nand NAND3_533 ( U2881 , U6174 , U6172 , U6173 );
nand NAND3_534 ( U2882 , U6171 , U6169 , U6170 );
nand NAND3_535 ( U2883 , U6168 , U6166 , U6167 );
nand NAND3_536 ( U2884 , U6165 , U6163 , U6164 );
nand NAND3_537 ( U2885 , U6162 , U6160 , U6161 );
nand NAND3_538 ( U2886 , U6159 , U6157 , U6158 );
nand NAND3_539 ( U2887 , U6156 , U6154 , U6155 );
nand NAND3_540 ( U2888 , U6153 , U6151 , U6152 );
nand NAND3_541 ( U2889 , U6150 , U6148 , U6149 );
nand NAND3_542 ( U2890 , U6146 , U6145 , U6147 );
nand NAND3_543 ( U2891 , U6143 , U6142 , U6144 );
and AND2_544 ( U2892 , DATAO_REG_31_ , U6043 );
nand NAND2_545 ( U2893 , U3870 , U6134 );
nand NAND2_546 ( U2894 , U3869 , U6131 );
nand NAND2_547 ( U2895 , U3868 , U6128 );
nand NAND2_548 ( U2896 , U3867 , U6125 );
nand NAND2_549 ( U2897 , U3866 , U6122 );
nand NAND2_550 ( U2898 , U3865 , U6119 );
nand NAND2_551 ( U2899 , U3864 , U6116 );
nand NAND2_552 ( U2900 , U3863 , U6113 );
nand NAND2_553 ( U2901 , U3862 , U6110 );
nand NAND2_554 ( U2902 , U3861 , U6107 );
nand NAND2_555 ( U2903 , U3860 , U6104 );
nand NAND2_556 ( U2904 , U3859 , U6101 );
nand NAND2_557 ( U2905 , U3858 , U6098 );
nand NAND2_558 ( U2906 , U3857 , U6095 );
nand NAND2_559 ( U2907 , U3856 , U6092 );
nand NAND3_560 ( U2908 , U6090 , U6089 , U6091 );
nand NAND3_561 ( U2909 , U6087 , U6086 , U6088 );
nand NAND3_562 ( U2910 , U6084 , U6083 , U6085 );
nand NAND3_563 ( U2911 , U6081 , U6080 , U6082 );
nand NAND3_564 ( U2912 , U6078 , U6077 , U6079 );
nand NAND3_565 ( U2913 , U6075 , U6074 , U6076 );
nand NAND3_566 ( U2914 , U6072 , U6071 , U6073 );
nand NAND3_567 ( U2915 , U6069 , U6068 , U6070 );
nand NAND3_568 ( U2916 , U6066 , U6065 , U6067 );
nand NAND3_569 ( U2917 , U6063 , U6062 , U6064 );
nand NAND3_570 ( U2918 , U6060 , U6059 , U6061 );
nand NAND3_571 ( U2919 , U6057 , U6056 , U6058 );
nand NAND3_572 ( U2920 , U6054 , U6053 , U6055 );
nand NAND3_573 ( U2921 , U6051 , U6050 , U6052 );
nand NAND3_574 ( U2922 , U6048 , U6047 , U6049 );
nand NAND3_575 ( U2923 , U6045 , U6044 , U6046 );
nand NAND2_576 ( U2924 , U7528 , U7530 );
nand NAND2_577 ( U2925 , U7527 , U7532 );
nand NAND2_578 ( U2926 , U7526 , U7534 );
nand NAND2_579 ( U2927 , U7525 , U7536 );
nand NAND2_580 ( U2928 , U7524 , U7538 );
nand NAND2_581 ( U2929 , U7523 , U7540 );
nand NAND2_582 ( U2930 , U7522 , U7542 );
nand NAND2_583 ( U2931 , U7521 , U7544 );
nand NAND2_584 ( U2932 , U7520 , U7546 );
nand NAND2_585 ( U2933 , U7519 , U7548 );
nand NAND2_586 ( U2934 , U7518 , U7550 );
nand NAND2_587 ( U2935 , U7517 , U7552 );
nand NAND2_588 ( U2936 , U7516 , U7554 );
nand NAND2_589 ( U2937 , U7515 , U7556 );
nand NAND2_590 ( U2938 , U7514 , U7558 );
nand NAND2_591 ( U2939 , U7513 , U7560 );
nand NAND2_592 ( U2940 , U7512 , U7562 );
nand NAND2_593 ( U2941 , U7511 , U7564 );
nand NAND2_594 ( U2942 , U7510 , U7566 );
nand NAND2_595 ( U2943 , U7509 , U7568 );
nand NAND2_596 ( U2944 , U7508 , U7570 );
nand NAND2_597 ( U2945 , U7507 , U7572 );
nand NAND2_598 ( U2946 , U7506 , U7574 );
nand NAND2_599 ( U2947 , U7505 , U7576 );
nand NAND2_600 ( U2948 , U7504 , U7578 );
nand NAND2_601 ( U2949 , U7503 , U7580 );
nand NAND2_602 ( U2950 , U7502 , U7582 );
nand NAND2_603 ( U2951 , U7501 , U7584 );
nand NAND2_604 ( U2952 , U7500 , U7586 );
nand NAND2_605 ( U2953 , U7499 , U7588 );
nand NAND2_606 ( U2954 , U7498 , U7590 );
nand NAND5_607 ( U2955 , U5944 , U5942 , U5946 , U5943 , U5945 );
nand NAND5_608 ( U2956 , U5939 , U5937 , U5941 , U5938 , U5940 );
nand NAND5_609 ( U2957 , U5934 , U5932 , U5936 , U5933 , U5935 );
nand NAND5_610 ( U2958 , U5929 , U5927 , U5931 , U5928 , U5930 );
nand NAND5_611 ( U2959 , U5924 , U5922 , U5926 , U5923 , U5925 );
nand NAND5_612 ( U2960 , U5919 , U5917 , U5921 , U5918 , U5920 );
nand NAND5_613 ( U2961 , U5914 , U5912 , U5916 , U5913 , U5915 );
nand NAND5_614 ( U2962 , U5909 , U5907 , U5911 , U5908 , U5910 );
nand NAND5_615 ( U2963 , U5904 , U5902 , U5906 , U5903 , U5905 );
nand NAND5_616 ( U2964 , U5899 , U5897 , U5901 , U5898 , U5900 );
nand NAND5_617 ( U2965 , U5894 , U5892 , U5896 , U5893 , U5895 );
nand NAND5_618 ( U2966 , U5889 , U5887 , U5891 , U5888 , U5890 );
nand NAND5_619 ( U2967 , U5884 , U5882 , U5886 , U5883 , U5885 );
nand NAND5_620 ( U2968 , U5879 , U5877 , U5881 , U5878 , U5880 );
nand NAND5_621 ( U2969 , U5874 , U5872 , U5876 , U5873 , U5875 );
nand NAND5_622 ( U2970 , U5869 , U5867 , U5871 , U5868 , U5870 );
nand NAND5_623 ( U2971 , U5864 , U5862 , U5866 , U5863 , U5865 );
nand NAND5_624 ( U2972 , U5859 , U5857 , U5861 , U5858 , U5860 );
nand NAND5_625 ( U2973 , U5854 , U5852 , U5856 , U5853 , U5855 );
nand NAND5_626 ( U2974 , U5849 , U5847 , U5851 , U5848 , U5850 );
nand NAND5_627 ( U2975 , U5844 , U5842 , U5846 , U5843 , U5845 );
nand NAND5_628 ( U2976 , U5839 , U5837 , U5841 , U5838 , U5840 );
nand NAND5_629 ( U2977 , U5834 , U5832 , U5836 , U5833 , U5835 );
nand NAND5_630 ( U2978 , U5829 , U5827 , U5831 , U5828 , U5830 );
nand NAND5_631 ( U2979 , U5824 , U5822 , U5823 , U5826 , U5825 );
nand NAND5_632 ( U2980 , U5819 , U5817 , U5818 , U5821 , U5820 );
nand NAND5_633 ( U2981 , U5814 , U5812 , U5813 , U5816 , U5815 );
nand NAND5_634 ( U2982 , U5809 , U5807 , U5808 , U5811 , U5810 );
nand NAND5_635 ( U2983 , U5804 , U5802 , U5803 , U5806 , U5805 );
nand NAND5_636 ( U2984 , U5799 , U5797 , U5798 , U5801 , U5800 );
nand NAND5_637 ( U2985 , U5793 , U5792 , U5794 , U5796 , U5795 );
nand NAND5_638 ( U2986 , U5788 , U5787 , U5789 , U5791 , U5790 );
nand NAND4_639 ( U2987 , U3849 , U3847 , U5775 , U5777 );
nand NAND4_640 ( U2988 , U3846 , U3844 , U5768 , U5770 );
nand NAND4_641 ( U2989 , U3843 , U3841 , U5761 , U5763 );
nand NAND4_642 ( U2990 , U3840 , U3838 , U5754 , U5756 );
nand NAND4_643 ( U2991 , U3837 , U3835 , U5747 , U5749 );
nand NAND4_644 ( U2992 , U3834 , U3832 , U5740 , U5742 );
nand NAND4_645 ( U2993 , U3831 , U3829 , U5733 , U5735 );
nand NAND4_646 ( U2994 , U3828 , U3826 , U5726 , U5728 );
nand NAND4_647 ( U2995 , U3825 , U3823 , U5719 , U5721 );
nand NAND4_648 ( U2996 , U3822 , U3820 , U5712 , U5714 );
nand NAND4_649 ( U2997 , U3819 , U3817 , U5705 , U5707 );
nand NAND4_650 ( U2998 , U3816 , U3814 , U5698 , U5700 );
nand NAND4_651 ( U2999 , U3813 , U3811 , U5691 , U5693 );
nand NAND4_652 ( U3000 , U3810 , U3808 , U5684 , U5686 );
nand NAND4_653 ( U3001 , U3807 , U3805 , U5677 , U5679 );
nand NAND4_654 ( U3002 , U3804 , U3802 , U5670 , U5672 );
nand NAND4_655 ( U3003 , U3801 , U3799 , U5663 , U5665 );
nand NAND4_656 ( U3004 , U3798 , U3796 , U5656 , U5658 );
nand NAND4_657 ( U3005 , U3795 , U3793 , U5649 , U5651 );
nand NAND3_658 ( U3006 , U3790 , U3792 , U5644 );
nand NAND3_659 ( U3007 , U3787 , U3789 , U5637 );
nand NAND3_660 ( U3008 , U3784 , U3786 , U5630 );
nand NAND3_661 ( U3009 , U3781 , U3783 , U5623 );
nand NAND3_662 ( U3010 , U3778 , U3780 , U5616 );
nand NAND3_663 ( U3011 , U3775 , U3777 , U5609 );
nand NAND3_664 ( U3012 , U3772 , U3774 , U5602 );
nand NAND3_665 ( U3013 , U3769 , U3771 , U5595 );
nand NAND3_666 ( U3014 , U3766 , U3768 , U5588 );
nand NAND2_667 ( U3015 , U3763 , U3764 );
nand NAND3_668 ( U3016 , U3760 , U3759 , U3762 );
nand NAND3_669 ( U3017 , U3756 , U3755 , U3758 );
nand NAND3_670 ( U3018 , U3752 , U3751 , U3754 );
and AND2_671 ( U3019 , INSTQUEUEWR_ADDR_REG_4_ , U5525 );
nand NAND3_672 ( U3020 , U5448 , U5447 , U3718 );
nand NAND3_673 ( U3021 , U5443 , U5442 , U3717 );
nand NAND3_674 ( U3022 , U5438 , U5437 , U3716 );
nand NAND3_675 ( U3023 , U5433 , U5432 , U3715 );
nand NAND3_676 ( U3024 , U7600 , U5428 , U3714 );
nand NAND3_677 ( U3025 , U5424 , U5423 , U3713 );
nand NAND3_678 ( U3026 , U5419 , U5418 , U3712 );
nand NAND3_679 ( U3027 , U5414 , U5413 , U3711 );
nand NAND3_680 ( U3028 , U5392 , U5391 , U3709 );
nand NAND3_681 ( U3029 , U5387 , U5386 , U3708 );
nand NAND3_682 ( U3030 , U5382 , U5381 , U3707 );
nand NAND3_683 ( U3031 , U5377 , U5376 , U3706 );
nand NAND3_684 ( U3032 , U5372 , U5371 , U3705 );
nand NAND3_685 ( U3033 , U5367 , U5366 , U3704 );
nand NAND3_686 ( U3034 , U5362 , U5361 , U3703 );
nand NAND3_687 ( U3035 , U5357 , U5356 , U3702 );
nand NAND3_688 ( U3036 , U5334 , U5333 , U3700 );
nand NAND3_689 ( U3037 , U5329 , U5328 , U3699 );
nand NAND3_690 ( U3038 , U5324 , U5323 , U3698 );
nand NAND3_691 ( U3039 , U5319 , U5318 , U3697 );
nand NAND3_692 ( U3040 , U5314 , U5313 , U3696 );
nand NAND3_693 ( U3041 , U5309 , U5308 , U3695 );
nand NAND3_694 ( U3042 , U5304 , U5303 , U3694 );
nand NAND3_695 ( U3043 , U5299 , U5298 , U3693 );
nand NAND3_696 ( U3044 , U5277 , U5276 , U3691 );
nand NAND3_697 ( U3045 , U5272 , U5271 , U3690 );
nand NAND3_698 ( U3046 , U5267 , U5266 , U3689 );
nand NAND3_699 ( U3047 , U5262 , U5261 , U3688 );
nand NAND3_700 ( U3048 , U5257 , U5256 , U3687 );
nand NAND3_701 ( U3049 , U5252 , U5251 , U3686 );
nand NAND3_702 ( U3050 , U5247 , U5246 , U3685 );
nand NAND3_703 ( U3051 , U5242 , U5241 , U3684 );
nand NAND3_704 ( U3052 , U5219 , U5218 , U3682 );
nand NAND3_705 ( U3053 , U5214 , U5213 , U3681 );
nand NAND3_706 ( U3054 , U5209 , U5208 , U3680 );
nand NAND3_707 ( U3055 , U5204 , U5203 , U3679 );
nand NAND3_708 ( U3056 , U5199 , U5198 , U3678 );
nand NAND3_709 ( U3057 , U5194 , U5193 , U3677 );
nand NAND3_710 ( U3058 , U5189 , U5188 , U3676 );
nand NAND3_711 ( U3059 , U5184 , U5183 , U3675 );
nand NAND3_712 ( U3060 , U5162 , U5161 , U3673 );
nand NAND3_713 ( U3061 , U5157 , U5156 , U3672 );
nand NAND3_714 ( U3062 , U5152 , U5151 , U3671 );
nand NAND3_715 ( U3063 , U5147 , U5146 , U3670 );
nand NAND3_716 ( U3064 , U5142 , U5141 , U3669 );
nand NAND3_717 ( U3065 , U5137 , U5136 , U3668 );
nand NAND3_718 ( U3066 , U5132 , U5131 , U3667 );
nand NAND3_719 ( U3067 , U5127 , U5126 , U3666 );
nand NAND3_720 ( U3068 , U5104 , U5103 , U3664 );
nand NAND3_721 ( U3069 , U5099 , U5098 , U3663 );
nand NAND3_722 ( U3070 , U5094 , U5093 , U3662 );
nand NAND3_723 ( U3071 , U5089 , U5088 , U3661 );
nand NAND3_724 ( U3072 , U5084 , U5083 , U3660 );
nand NAND3_725 ( U3073 , U5079 , U5078 , U3659 );
nand NAND3_726 ( U3074 , U5074 , U5073 , U3658 );
nand NAND3_727 ( U3075 , U5069 , U5068 , U3657 );
nand NAND3_728 ( U3076 , U5047 , U5046 , U3655 );
nand NAND3_729 ( U3077 , U5042 , U5041 , U3654 );
nand NAND3_730 ( U3078 , U5037 , U5036 , U3653 );
nand NAND3_731 ( U3079 , U5032 , U5031 , U3652 );
nand NAND3_732 ( U3080 , U5027 , U5026 , U3651 );
nand NAND3_733 ( U3081 , U5022 , U5021 , U3650 );
nand NAND3_734 ( U3082 , U5017 , U5016 , U3649 );
nand NAND3_735 ( U3083 , U5012 , U5011 , U3648 );
nand NAND3_736 ( U3084 , U4991 , U4990 , U3646 );
nand NAND3_737 ( U3085 , U4986 , U4985 , U3645 );
nand NAND3_738 ( U3086 , U4981 , U4980 , U3644 );
nand NAND3_739 ( U3087 , U4976 , U4975 , U3643 );
nand NAND3_740 ( U3088 , U4971 , U4970 , U3642 );
nand NAND3_741 ( U3089 , U4966 , U4965 , U3641 );
nand NAND3_742 ( U3090 , U4961 , U4960 , U3640 );
nand NAND3_743 ( U3091 , U4956 , U4955 , U3639 );
nand NAND3_744 ( U3092 , U4934 , U4933 , U3637 );
nand NAND3_745 ( U3093 , U4929 , U4928 , U3636 );
nand NAND3_746 ( U3094 , U4924 , U4923 , U3635 );
nand NAND3_747 ( U3095 , U4919 , U4918 , U3634 );
nand NAND3_748 ( U3096 , U4914 , U4913 , U3633 );
nand NAND3_749 ( U3097 , U4909 , U4908 , U3632 );
nand NAND3_750 ( U3098 , U4904 , U4903 , U3631 );
nand NAND3_751 ( U3099 , U4899 , U4898 , U3630 );
nand NAND3_752 ( U3100 , U4876 , U4875 , U3628 );
nand NAND3_753 ( U3101 , U4871 , U4870 , U3627 );
nand NAND3_754 ( U3102 , U4866 , U4865 , U3626 );
nand NAND3_755 ( U3103 , U4861 , U4860 , U3625 );
nand NAND3_756 ( U3104 , U4856 , U4855 , U3624 );
nand NAND3_757 ( U3105 , U4851 , U4850 , U3623 );
nand NAND3_758 ( U3106 , U4846 , U4845 , U3622 );
nand NAND3_759 ( U3107 , U4841 , U4840 , U3621 );
nand NAND3_760 ( U3108 , U4819 , U4818 , U3619 );
nand NAND3_761 ( U3109 , U4814 , U4813 , U3618 );
nand NAND3_762 ( U3110 , U4809 , U4808 , U3617 );
nand NAND3_763 ( U3111 , U4804 , U4803 , U3616 );
nand NAND3_764 ( U3112 , U4799 , U4798 , U3615 );
nand NAND3_765 ( U3113 , U4794 , U4793 , U3614 );
nand NAND3_766 ( U3114 , U4789 , U4788 , U3613 );
nand NAND3_767 ( U3115 , U4784 , U4783 , U3612 );
nand NAND3_768 ( U3116 , U4761 , U4760 , U3610 );
nand NAND3_769 ( U3117 , U4756 , U4755 , U3609 );
nand NAND3_770 ( U3118 , U4751 , U4750 , U3608 );
nand NAND3_771 ( U3119 , U4746 , U4745 , U3607 );
nand NAND3_772 ( U3120 , U4741 , U4740 , U3606 );
nand NAND3_773 ( U3121 , U4736 , U4735 , U3605 );
nand NAND3_774 ( U3122 , U4731 , U4730 , U3604 );
nand NAND3_775 ( U3123 , U4726 , U4725 , U3603 );
nand NAND3_776 ( U3124 , U4704 , U4703 , U3601 );
nand NAND3_777 ( U3125 , U4699 , U4698 , U3600 );
nand NAND3_778 ( U3126 , U4694 , U4693 , U3599 );
nand NAND3_779 ( U3127 , U4689 , U4688 , U3598 );
nand NAND3_780 ( U3128 , U4684 , U4683 , U3597 );
nand NAND3_781 ( U3129 , U4679 , U4678 , U3596 );
nand NAND3_782 ( U3130 , U4674 , U4673 , U3595 );
nand NAND3_783 ( U3131 , U4669 , U4668 , U3594 );
nand NAND3_784 ( U3132 , U4645 , U4644 , U3592 );
nand NAND3_785 ( U3133 , U4640 , U4639 , U3591 );
nand NAND3_786 ( U3134 , U4635 , U4634 , U3590 );
nand NAND3_787 ( U3135 , U4630 , U4629 , U3589 );
nand NAND3_788 ( U3136 , U4625 , U4624 , U3588 );
nand NAND3_789 ( U3137 , U4620 , U4619 , U3587 );
nand NAND3_790 ( U3138 , U4615 , U4614 , U3586 );
nand NAND3_791 ( U3139 , U4610 , U4609 , U3585 );
nand NAND3_792 ( U3140 , U4587 , U4586 , U3583 );
nand NAND3_793 ( U3141 , U4582 , U4581 , U3582 );
nand NAND3_794 ( U3142 , U4577 , U4576 , U3581 );
nand NAND3_795 ( U3143 , U4572 , U4571 , U3580 );
nand NAND3_796 ( U3144 , U4567 , U4566 , U3579 );
nand NAND3_797 ( U3145 , U4562 , U4561 , U3578 );
nand NAND3_798 ( U3146 , U4557 , U4556 , U3577 );
nand NAND3_799 ( U3147 , U4552 , U4551 , U3576 );
nand NAND3_800 ( U3148 , U7678 , U7677 , U3574 );
nand NAND4_801 ( U3149 , U4508 , U4507 , U4506 , U4232 );
nand NAND2_802 ( U3150 , U3570 , U4504 );
and AND2_803 ( U3151 , DATAWIDTH_REG_31_ , U7638 );
and AND2_804 ( U3152 , DATAWIDTH_REG_30_ , U7638 );
and AND2_805 ( U3153 , DATAWIDTH_REG_29_ , U7638 );
and AND2_806 ( U3154 , DATAWIDTH_REG_28_ , U7638 );
and AND2_807 ( U3155 , DATAWIDTH_REG_27_ , U7638 );
and AND2_808 ( U3156 , DATAWIDTH_REG_26_ , U7638 );
and AND2_809 ( U3157 , DATAWIDTH_REG_25_ , U7638 );
and AND2_810 ( U3158 , DATAWIDTH_REG_24_ , U7638 );
and AND2_811 ( U3159 , DATAWIDTH_REG_23_ , U7638 );
and AND2_812 ( U3160 , DATAWIDTH_REG_22_ , U7638 );
and AND2_813 ( U3161 , DATAWIDTH_REG_21_ , U7638 );
and AND2_814 ( U3162 , DATAWIDTH_REG_20_ , U7638 );
and AND2_815 ( U3163 , DATAWIDTH_REG_19_ , U7638 );
and AND2_816 ( U3164 , DATAWIDTH_REG_18_ , U7638 );
and AND2_817 ( U3165 , DATAWIDTH_REG_17_ , U7638 );
and AND2_818 ( U3166 , DATAWIDTH_REG_16_ , U7638 );
and AND2_819 ( U3167 , DATAWIDTH_REG_15_ , U7638 );
and AND2_820 ( U3168 , DATAWIDTH_REG_14_ , U7638 );
and AND2_821 ( U3169 , DATAWIDTH_REG_13_ , U7638 );
and AND2_822 ( U3170 , DATAWIDTH_REG_12_ , U7638 );
and AND2_823 ( U3171 , DATAWIDTH_REG_11_ , U7638 );
and AND2_824 ( U3172 , DATAWIDTH_REG_10_ , U7638 );
and AND2_825 ( U3173 , DATAWIDTH_REG_9_ , U7638 );
and AND2_826 ( U3174 , DATAWIDTH_REG_8_ , U7638 );
and AND2_827 ( U3175 , DATAWIDTH_REG_7_ , U7638 );
and AND2_828 ( U3176 , DATAWIDTH_REG_6_ , U7638 );
and AND2_829 ( U3177 , DATAWIDTH_REG_5_ , U7638 );
and AND2_830 ( U3178 , DATAWIDTH_REG_4_ , U7638 );
and AND2_831 ( U3179 , DATAWIDTH_REG_3_ , U7638 );
and AND2_832 ( U3180 , DATAWIDTH_REG_2_ , U7638 );
nand NAND3_833 ( U3181 , U7635 , U7634 , U4363 );
nand NAND3_834 ( U3182 , U7633 , U7632 , U3483 );
nand NAND2_835 ( U3183 , U3482 , U4357 );
nand NAND3_836 ( U3184 , U4343 , U4342 , U4344 );
nand NAND3_837 ( U3185 , U4340 , U4339 , U4341 );
nand NAND3_838 ( U3186 , U4337 , U4336 , U4338 );
nand NAND3_839 ( U3187 , U4334 , U4333 , U4335 );
nand NAND3_840 ( U3188 , U4331 , U4330 , U4332 );
nand NAND3_841 ( U3189 , U4328 , U4327 , U4329 );
nand NAND3_842 ( U3190 , U4325 , U4324 , U4326 );
nand NAND3_843 ( U3191 , U4322 , U4321 , U4323 );
nand NAND3_844 ( U3192 , U4319 , U4318 , U4320 );
nand NAND3_845 ( U3193 , U4316 , U4315 , U4317 );
nand NAND3_846 ( U3194 , U4313 , U4312 , U4314 );
nand NAND3_847 ( U3195 , U4310 , U4309 , U4311 );
nand NAND3_848 ( U3196 , U4307 , U4306 , U4308 );
nand NAND3_849 ( U3197 , U4304 , U4303 , U4305 );
nand NAND3_850 ( U3198 , U4301 , U4300 , U4302 );
nand NAND3_851 ( U3199 , U4298 , U4297 , U4299 );
nand NAND3_852 ( U3200 , U4295 , U4294 , U4296 );
nand NAND3_853 ( U3201 , U4292 , U4291 , U4293 );
nand NAND3_854 ( U3202 , U4289 , U4288 , U4290 );
nand NAND3_855 ( U3203 , U4286 , U4285 , U4287 );
nand NAND3_856 ( U3204 , U4283 , U4282 , U4284 );
nand NAND3_857 ( U3205 , U4280 , U4279 , U4281 );
nand NAND3_858 ( U3206 , U4277 , U4276 , U4278 );
nand NAND3_859 ( U3207 , U4274 , U4273 , U4275 );
nand NAND3_860 ( U3208 , U4271 , U4270 , U4272 );
nand NAND3_861 ( U3209 , U4268 , U4267 , U4269 );
nand NAND3_862 ( U3210 , U4265 , U4264 , U4266 );
nand NAND3_863 ( U3211 , U4262 , U4261 , U4263 );
nand NAND3_864 ( U3212 , U4259 , U4258 , U4260 );
nand NAND3_865 ( U3213 , U4256 , U4255 , U4257 );
nand NAND4_866 ( U3214 , U3989 , U3988 , U3987 , U3986 );
nand NAND4_867 ( U3215 , U3985 , U3984 , U3983 , U3982 );
nand NAND4_868 ( U3216 , U3981 , U3980 , U3979 , U3978 );
nand NAND4_869 ( U3217 , U3977 , U3976 , U3975 , U3974 );
nand NAND4_870 ( U3218 , U3973 , U3972 , U3971 , U3970 );
nand NAND4_871 ( U3219 , U3969 , U3968 , U3967 , U3966 );
nand NAND4_872 ( U3220 , U3965 , U3964 , U3963 , U3962 );
nand NAND4_873 ( U3221 , U3961 , U3960 , U3959 , U3958 );
nand NAND2_874 ( U3222 , U3316 , U3310 );
nand NAND2_875 ( U3223 , U2432 , U3222 );
nand NAND2_876 ( U3224 , U2432 , U4531 );
nand NAND2_877 ( U3225 , U2434 , U3222 );
nand NAND2_878 ( U3226 , U2434 , U4531 );
nand NAND2_879 ( U3227 , U2433 , U3222 );
nand NAND2_880 ( U3228 , U2433 , U4531 );
nand NAND2_881 ( U3229 , U2435 , U3222 );
nand NAND2_882 ( U3230 , U2435 , U4531 );
nand NAND3_883 ( U3231 , U3378 , U3381 , U5451 );
nand NAND2_884 ( U3232 , U7074 , U5452 );
nand NAND4_885 ( U3233 , U7780 , U7779 , U4146 , U4144 );
not NOT1_886 ( U3234 , REQUESTPENDING_REG );
not NOT1_887 ( U3235 , STATE_REG_1_ );
nand NAND2_888 ( U3236 , STATE_REG_1_ , U3245 );
nand NAND2_889 ( U3237 , U4209 , U3238 );
not NOT1_890 ( U3238 , STATE_REG_2_ );
nand NAND2_891 ( U3239 , STATE_REG_2_ , U4209 );
not NOT1_892 ( U3240 , REIP_REG_1_ );
nand NAND2_893 ( U3241 , STATE_REG_1_ , U3238 );
or OR2_894 ( U3242 , STATE_REG_1_ , STATE_REG_2_ );
not NOT1_895 ( U3243 , HOLD );
not NOT1_896 ( U3244 , READY_N );
not NOT1_897 ( U3245 , STATE_REG_0_ );
nand NAND2_898 ( U3246 , STATE_REG_0_ , U3247 );
nand NAND2_899 ( U3247 , REQUESTPENDING_REG , U3243 );
or OR2_900 ( U3248 , HOLD , REQUESTPENDING_REG );
not NOT1_901 ( U3249 , STATE2_REG_1_ );
not NOT1_902 ( U3250 , STATE2_REG_2_ );
not NOT1_903 ( U3251 , INSTQUEUERD_ADDR_REG_2_ );
not NOT1_904 ( U3252 , INSTQUEUERD_ADDR_REG_1_ );
not NOT1_905 ( U3253 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND4_906 ( U3254 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ , U3257 );
or OR3_907 ( U3255 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ );
or OR2_908 ( U3256 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_0_ );
not NOT1_909 ( U3257 , INSTQUEUERD_ADDR_REG_3_ );
nand NAND4_910 ( U3258 , U3555 , U3554 , U3553 , U3552 );
nand NAND2_911 ( U3259 , U4484 , U3245 );
not NOT1_912 ( U3260 , R2167_U17 );
nand NAND2_913 ( U3261 , INSTQUEUERD_ADDR_REG_2_ , U3257 );
nand NAND2_914 ( U3262 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ );
nand NAND4_915 ( U3263 , U3507 , U3506 , U3505 , U3504 );
nand NAND5_916 ( U3264 , U3527 , U4158 , U3526 , U3525 , U3524 );
nand NAND4_917 ( U3265 , U3545 , U3544 , U3543 , U3542 );
nand NAND2_918 ( U3266 , U3547 , U3546 );
or OR2_919 ( U3267 , STATEBS16_REG , READY_N );
nand NAND2_920 ( U3268 , R2167_U17 , U4485 );
nand NAND2_921 ( U3269 , U4465 , U3271 );
nand NAND4_922 ( U3270 , U3499 , U3498 , U3497 , U3496 );
nand NAND4_923 ( U3271 , U3551 , U3550 , U3549 , U3548 );
nand NAND2_924 ( U3272 , U2473 , U4489 );
nand NAND2_925 ( U3273 , U2389 , U3270 );
nand NAND2_926 ( U3274 , U4482 , U4465 );
nand NAND2_927 ( U3275 , U4237 , U2447 );
nand NAND4_928 ( U3276 , U4448 , U3378 , U4161 , U3265 );
nand NAND2_929 ( U3277 , U3258 , U3270 );
nand NAND2_930 ( U3278 , U4178 , U3271 );
nand NAND2_931 ( U3279 , U4244 , U2431 );
nand NAND5_932 ( U3280 , U4166 , U4497 , U7614 , U4213 , LT_563_U6 );
not NOT1_933 ( U3281 , STATE2_REG_0_ );
nand NAND2_934 ( U3282 , STATE2_REG_0_ , U7592 );
not NOT1_935 ( U3283 , STATE2_REG_3_ );
nand NAND2_936 ( U3284 , STATE2_REG_2_ , U3249 );
or OR2_937 ( U3285 , STATE2_REG_2_ , STATE2_REG_1_ );
nand NAND2_938 ( U3286 , STATE2_REG_3_ , R2167_U17 );
nand NAND2_939 ( U3287 , U4535 , U3281 );
not NOT1_940 ( U3288 , INSTQUEUEWR_ADDR_REG_0_ );
not NOT1_941 ( U3289 , INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_942 ( U3290 , INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_943 ( U3291 , INSTQUEUEWR_ADDR_REG_2_ );
nand NAND2_944 ( U3292 , INSTQUEUEWR_ADDR_REG_1_ , INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_945 ( U3293 , U4521 , U2478 );
or OR2_946 ( U3294 , STATE2_REG_2_ , STATE2_REG_3_ );
not NOT1_947 ( U3295 , STATEBS16_REG );
not NOT1_948 ( U3296 , R2144_U43 );
not NOT1_949 ( U3297 , R2144_U50 );
not NOT1_950 ( U3298 , R2144_U49 );
not NOT1_951 ( U3299 , R2144_U8 );
nand NAND2_952 ( U3300 , R2144_U50 , R2144_U43 );
nand NAND2_953 ( U3301 , U3319 , U3296 );
nand NAND2_954 ( U3302 , U4515 , U2475 );
not NOT1_955 ( U3303 , R2182_U25 );
not NOT1_956 ( U3304 , R2182_U42 );
not NOT1_957 ( U3305 , R2182_U34 );
not NOT1_958 ( U3306 , R2182_U33 );
nand NAND2_959 ( U3307 , U4197 , U3295 );
nand NAND2_960 ( U3308 , U3293 , U4523 );
nand NAND2_961 ( U3309 , U3293 , U4532 );
nand NAND2_962 ( U3310 , INSTQUEUEWR_ADDR_REG_1_ , U3288 );
nand NAND2_963 ( U3311 , U4530 , U2478 );
nand NAND2_964 ( U3312 , R2144_U50 , U3296 );
nand NAND2_965 ( U3313 , R2144_U43 , U3319 );
nand NAND2_966 ( U3314 , U4588 , U2475 );
nand NAND2_967 ( U3315 , U3311 , U4591 );
nand NAND2_968 ( U3316 , INSTQUEUEWR_ADDR_REG_0_ , U3289 );
nand NAND2_969 ( U3317 , U4529 , U2478 );
nand NAND2_970 ( U3318 , R2144_U43 , U3297 );
nand NAND2_971 ( U3319 , U3312 , U3318 );
nand NAND2_972 ( U3320 , U4514 , U3296 );
nand NAND2_973 ( U3321 , U4646 , U2475 );
nand NAND2_974 ( U3322 , U3317 , U4649 );
nand NAND2_975 ( U3323 , U3317 , U4651 );
nand NAND2_976 ( U3324 , U2488 , U2478 );
nand NAND2_977 ( U3325 , U2485 , U2475 );
nand NAND2_978 ( U3326 , U3324 , U4707 );
nand NAND2_979 ( U3327 , INSTQUEUEWR_ADDR_REG_3_ , U3291 );
nand NAND2_980 ( U3328 , U4526 , U4521 );
nand NAND2_981 ( U3329 , R2144_U8 , U3298 );
nand NAND2_982 ( U3330 , U2490 , U4515 );
nand NAND2_983 ( U3331 , U3328 , U4764 );
nand NAND2_984 ( U3332 , U3328 , U4766 );
nand NAND2_985 ( U3333 , U4526 , U4530 );
nand NAND2_986 ( U3334 , U2490 , U4588 );
nand NAND2_987 ( U3335 , U3333 , U4822 );
nand NAND2_988 ( U3336 , U4526 , U4529 );
nand NAND2_989 ( U3337 , U2490 , U4646 );
nand NAND2_990 ( U3338 , U3336 , U4879 );
nand NAND2_991 ( U3339 , U3336 , U4881 );
nand NAND2_992 ( U3340 , U4526 , U2488 );
nand NAND2_993 ( U3341 , U2490 , U2485 );
nand NAND2_994 ( U3342 , U3340 , U4937 );
nand NAND2_995 ( U3343 , U2479 , U4521 );
nand NAND2_996 ( U3344 , U2474 , U4516 );
nand NAND3_997 ( U3345 , U3329 , U4518 , U3344 );
nand NAND2_998 ( U3346 , U2499 , U4515 );
nand NAND3_999 ( U3347 , U3327 , U4527 , U3343 );
nand NAND2_1000 ( U3348 , U3343 , U4993 );
nand NAND2_1001 ( U3349 , U3343 , U4995 );
nand NAND2_1002 ( U3350 , U4530 , U2479 );
nand NAND2_1003 ( U3351 , U2499 , U4588 );
nand NAND2_1004 ( U3352 , U3350 , U5050 );
nand NAND2_1005 ( U3353 , U4529 , U2479 );
nand NAND2_1006 ( U3354 , U2499 , U4646 );
nand NAND2_1007 ( U3355 , U3353 , U5107 );
nand NAND2_1008 ( U3356 , U3353 , U5109 );
nand NAND2_1009 ( U3357 , U2488 , U2479 );
nand NAND2_1010 ( U3358 , U2499 , U2485 );
nand NAND2_1011 ( U3359 , U3357 , U5165 );
nand NAND2_1012 ( U3360 , U2510 , U4521 );
nand NAND2_1013 ( U3361 , U2507 , U4515 );
nand NAND2_1014 ( U3362 , U3360 , U5222 );
nand NAND2_1015 ( U3363 , U3360 , U5224 );
nand NAND2_1016 ( U3364 , U2510 , U4530 );
nand NAND2_1017 ( U3365 , U2507 , U4588 );
nand NAND2_1018 ( U3366 , U3364 , U5280 );
nand NAND2_1019 ( U3367 , U2510 , U4529 );
nand NAND2_1020 ( U3368 , U2507 , U4646 );
nand NAND2_1021 ( U3369 , U3367 , U5337 );
nand NAND2_1022 ( U3370 , U3367 , U5339 );
nand NAND2_1023 ( U3371 , U2510 , U2488 );
nand NAND2_1024 ( U3372 , U2507 , U2485 );
nand NAND2_1025 ( U3373 , U3371 , U5395 );
not NOT1_1026 ( U3374 , FLUSH_REG );
not NOT1_1027 ( U3375 , GTE_485_U6 );
nand NAND2_1028 ( U3376 , U3271 , U3265 );
nand NAND2_1029 ( U3377 , U3271 , U3258 );
nand NAND4_1030 ( U3378 , U3503 , U3502 , U3501 , U3500 );
nand NAND3_1031 ( U3379 , U5478 , U5477 , U7616 );
nand NAND2_1032 ( U3380 , U4387 , U3271 );
nand NAND2_1033 ( U3381 , U2605 , U3264 );
nand NAND3_1034 ( U3382 , U4387 , U7482 , U4482 );
nand NAND2_1035 ( U3383 , U3729 , U4235 );
nand NAND5_1036 ( U3384 , U7482 , U4465 , U2605 , U4482 , U4387 );
nand NAND5_1037 ( U3385 , U2605 , U4448 , U4159 , U4437 , U4388 );
nand NAND3_1038 ( U3386 , U4187 , U4465 , U4222 );
nand NAND2_1039 ( U3387 , U2449 , U2447 );
nand NAND2_1040 ( U3388 , U3431 , U5498 );
nand NAND2_1041 ( U3389 , U3256 , U3262 );
not NOT1_1042 ( U3390 , LT_589_U6 );
nand NAND3_1043 ( U3391 , U4230 , U3287 , U5524 );
nand NAND3_1044 ( U3392 , STATE2_REG_0_ , U3265 , U3271 );
nand NAND2_1045 ( U3393 , U3258 , U3260 );
nand NAND2_1046 ( U3394 , U3264 , U3378 );
nand NAND2_1047 ( U3395 , U2427 , U3281 );
nand NAND2_1048 ( U3396 , U4448 , U3378 );
nand NAND2_1049 ( U3397 , U4241 , U3265 );
nand NAND2_1050 ( U3398 , U4178 , U2452 );
nand NAND2_1051 ( U3399 , STATE2_REG_2_ , U3258 );
not NOT1_1052 ( U3400 , REIP_REG_0_ );
nand NAND2_1053 ( U3401 , U3744 , U5550 );
nand NAND2_1054 ( U3402 , U4388 , U4161 );
nand NAND2_1055 ( U3403 , U3851 , U4236 );
nand NAND2_1056 ( U3404 , U6042 , U6041 );
nand NAND2_1057 ( U3405 , STATE2_REG_0_ , U4482 );
nand NAND2_1058 ( U3406 , U4387 , U7482 );
nand NAND2_1059 ( U3407 , U4194 , U4465 );
nand NAND2_1060 ( U3408 , U4182 , U2431 );
nand NAND2_1061 ( U3409 , U4198 , STATE2_REG_0_ );
nand NAND2_1062 ( U3410 , U4491 , U3378 );
nand NAND2_1063 ( U3411 , U4223 , U6141 );
nand NAND2_1064 ( U3412 , STATE2_REG_0_ , U4204 );
nand NAND2_1065 ( U3413 , U4223 , U6252 );
nand NAND4_1066 ( U3414 , STATE2_REG_0_ , U4237 , U3874 , U2452 );
nand NAND2_1067 ( U3415 , U3854 , U2447 );
not NOT1_1068 ( U3416 , EBX_REG_31_ );
not NOT1_1069 ( U3417 , R2337_U58 );
nand NAND2_1070 ( U3418 , U4216 , U3875 );
nand NAND2_1071 ( U3419 , U4197 , U3249 );
nand NAND4_1072 ( U3420 , U3950 , U3946 , U3943 , U3940 );
nand NAND2_1073 ( U3421 , U4194 , U3258 );
not NOT1_1074 ( U3422 , CODEFETCH_REG );
not NOT1_1075 ( U3423 , READREQUEST_REG );
nand NAND2_1076 ( U3424 , U2447 , U4486 );
nand NAND2_1077 ( U3425 , U3254 , U5470 );
nand NAND2_1078 ( U3426 , U4437 , STATE2_REG_2_ );
nand NAND2_1079 ( U3427 , STATEBS16_REG , U3250 );
not NOT1_1080 ( U3428 , U3221 );
nand NAND2_1081 ( U3429 , U5467 , U5466 );
nand NAND2_1082 ( U3430 , U2450 , U3428 );
nand NAND3_1083 ( U3431 , INSTQUEUERD_ADDR_REG_1_ , U3251 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_1084 ( U3432 , U3261 , U7052 );
nand NAND2_1085 ( U3433 , U4185 , U4222 );
nand NAND3_1086 ( U3434 , U4219 , U4388 , U4238 );
nand NAND3_1087 ( U3435 , U4219 , U3265 , U4238 );
nand NAND2_1088 ( U3436 , U4465 , U4484 );
nand NAND4_1089 ( U3437 , U4062 , U7081 , U4063 , U4065 );
nand NAND2_1090 ( U3438 , U4242 , U4254 );
nand NAND2_1091 ( U3439 , U4171 , U3255 );
nand NAND2_1092 ( U3440 , STATE2_REG_0_ , U2605 );
nand NAND2_1093 ( U3441 , U7680 , U7679 );
nand NAND2_1094 ( U3442 , U7683 , U7682 );
nand NAND2_1095 ( U3443 , U7707 , U7706 );
nand NAND2_1096 ( U3444 , U7777 , U7776 );
nand NAND2_1097 ( U3445 , U7622 , U7621 );
nand NAND2_1098 ( U3446 , U7624 , U7623 );
nand NAND2_1099 ( U3447 , U7626 , U7625 );
nand NAND2_1100 ( U3448 , U7628 , U7627 );
nand NAND2_1101 ( U3449 , U7637 , U7636 );
and AND2_1102 ( U3450 , U3242 , U4167 );
nand NAND2_1103 ( U3451 , U7640 , U7639 );
nand NAND2_1104 ( U3452 , U7642 , U7641 );
nand NAND2_1105 ( U3453 , U7674 , U7673 );
and AND3_1106 ( U3454 , U2427 , U4203 , R2182_U24 );
nand NAND2_1107 ( U3455 , U7690 , U7689 );
nand NAND2_1108 ( U3456 , U7697 , U7696 );
nand NAND2_1109 ( U3457 , U7699 , U7698 );
nand NAND2_1110 ( U3458 , U7702 , U7701 );
nand NAND2_1111 ( U3459 , U7710 , U7709 );
nand NAND2_1112 ( U3460 , U7712 , U7711 );
nand NAND2_1113 ( U3461 , U7716 , U7715 );
nand NAND2_1114 ( U3462 , U7718 , U7717 );
nand NAND2_1115 ( U3463 , U7723 , U7722 );
nand NAND2_1116 ( U3464 , U7725 , U7724 );
nand NAND2_1117 ( U3465 , U7727 , U7726 );
and AND2_1118 ( U3466 , R2358_U91 , U4437 );
nor nor_1119 ( U3467 , DATAWIDTH_REG_1_ , REIP_REG_1_ );
nand NAND2_1120 ( U3468 , U7743 , U7742 );
nand NAND2_1121 ( U3469 , U7747 , U7746 );
nand NAND2_1122 ( U3470 , U7749 , U7748 );
nand NAND2_1123 ( U3471 , U7751 , U7750 );
nand NAND2_1124 ( U3472 , U7755 , U7754 );
nand NAND2_1125 ( U3473 , U7759 , U7758 );
nand NAND2_1126 ( U3474 , U7761 , U7760 );
and AND2_1127 ( U3475 , R2182_U24 , U4203 );
nand NAND2_1128 ( U3476 , U7763 , U7762 );
nand NAND2_1129 ( U3477 , U7765 , U7764 );
nand NAND2_1130 ( U3478 , U7767 , U7766 );
nand NAND2_1131 ( U3479 , U7769 , U7768 );
nand NAND2_1132 ( U3480 , U7771 , U7770 );
and AND2_1133 ( U3481 , STATE_REG_1_ , READY_N );
and AND2_1134 ( U3482 , U4356 , U3239 );
and AND2_1135 ( U3483 , U4358 , U3237 );
and AND2_1136 ( U3484 , REQUESTPENDING_REG , STATE_REG_0_ );
nor nor_1137 ( U3485 , INSTQUEUERD_ADDR_REG_2_ , INSTQUEUERD_ADDR_REG_3_ );
and AND2_1138 ( U3486 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ );
nor nor_1139 ( U3487 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_3_ );
and AND2_1140 ( U3488 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_2_ );
nor nor_1141 ( U3489 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_3_ );
and AND2_1142 ( U3490 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ );
nor nor_1143 ( U3491 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ );
and AND2_1144 ( U3492 , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_0_ );
nor nor_1145 ( U3493 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_2_ );
and AND2_1146 ( U3494 , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_1_ );
and AND2_1147 ( U3495 , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_2_ );
and AND4_1148 ( U3496 , U4374 , U4373 , U4372 , U4371 );
and AND4_1149 ( U3497 , U4378 , U4377 , U4376 , U4375 );
and AND4_1150 ( U3498 , U4382 , U4381 , U4380 , U4379 );
and AND4_1151 ( U3499 , U4386 , U4385 , U4384 , U4383 );
and AND4_1152 ( U3500 , U4424 , U4423 , U4422 , U4421 );
and AND4_1153 ( U3501 , U4428 , U4427 , U4426 , U4425 );
and AND4_1154 ( U3502 , U4432 , U4431 , U4430 , U4429 );
and AND4_1155 ( U3503 , U4436 , U4435 , U4434 , U4433 );
and AND4_1156 ( U3504 , U4407 , U4406 , U4405 , U4404 );
and AND4_1157 ( U3505 , U4411 , U4410 , U4409 , U4408 );
and AND4_1158 ( U3506 , U4415 , U4414 , U4413 , U4412 );
and AND4_1159 ( U3507 , U4419 , U4418 , U4417 , U4416 );
nor nor_1160 ( U3508 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_3_ );
and AND2_1161 ( U3509 , INSTQUEUE_REG_5__5_ , INSTQUEUERD_ADDR_REG_0_ );
nor nor_1162 ( U3510 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_3_ );
and AND2_1163 ( U3511 , INSTQUEUE_REG_6__5_ , INSTQUEUERD_ADDR_REG_1_ );
and AND2_1164 ( U3512 , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUE_REG_8__5_ );
nor nor_1165 ( U3513 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_2_ );
and AND2_1166 ( U3514 , INSTQUEUE_REG_10__5_ , INSTQUEUERD_ADDR_REG_3_ );
and AND2_1167 ( U3515 , INSTQUEUE_REG_12__5_ , INSTQUEUERD_ADDR_REG_3_ );
nor nor_1168 ( U3516 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ );
and AND2_1169 ( U3517 , INSTQUEUE_REG_9__5_ , INSTQUEUERD_ADDR_REG_0_ );
and AND4_1170 ( U3518 , U4392 , U4391 , U4390 , U4389 );
and AND4_1171 ( U3519 , U4396 , U4395 , U4394 , U4393 );
and AND4_1172 ( U3520 , U4400 , U4399 , U4398 , U4397 );
and AND2_1173 ( U3521 , U4402 , U4401 );
nor nor_1174 ( U3522 , INSTQUEUERD_ADDR_REG_2_ , INSTQUEUERD_ADDR_REG_3_ );
and AND2_1175 ( U3523 , INSTQUEUE_REG_3__6_ , INSTQUEUERD_ADDR_REG_0_ );
and AND4_1176 ( U3524 , U4441 , U4440 , U4439 , U4438 );
and AND3_1177 ( U3525 , U4443 , U4442 , U4444 );
and AND3_1178 ( U3526 , U4446 , U4445 , U4447 );
and AND4_1179 ( U3527 , U7666 , U7665 , U7664 , U7663 );
nor nor_1180 ( U3528 , INSTQUEUERD_ADDR_REG_2_ , INSTQUEUERD_ADDR_REG_3_ );
and AND2_1181 ( U3529 , INSTQUEUE_REG_1__4_ , INSTQUEUERD_ADDR_REG_0_ );
nor nor_1182 ( U3530 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ );
and AND2_1183 ( U3531 , INSTQUEUE_REG_4__4_ , INSTQUEUERD_ADDR_REG_2_ );
nor nor_1184 ( U3532 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ );
and AND2_1185 ( U3533 , INSTQUEUE_REG_12__4_ , INSTQUEUERD_ADDR_REG_2_ );
and AND2_1186 ( U3534 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_2_ );
and AND2_1187 ( U3535 , INSTQUEUE_REG_13__4_ , INSTQUEUERD_ADDR_REG_3_ );
nor nor_1188 ( U3536 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_3_ );
and AND2_1189 ( U3537 , INSTQUEUE_REG_6__4_ , INSTQUEUERD_ADDR_REG_2_ );
and AND2_1190 ( U3538 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ );
and AND2_1191 ( U3539 , INSTQUEUE_REG_14__4_ , INSTQUEUERD_ADDR_REG_3_ );
nor nor_1192 ( U3540 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ );
and AND2_1193 ( U3541 , INSTQUEUE_REG_9__4_ , INSTQUEUERD_ADDR_REG_3_ );
and AND4_1194 ( U3542 , U7646 , U7645 , U7644 , U7643 );
and AND4_1195 ( U3543 , U7650 , U7649 , U7648 , U7647 );
and AND4_1196 ( U3544 , U7654 , U7653 , U7652 , U7651 );
and AND4_1197 ( U3545 , U7658 , U7657 , U7656 , U7655 );
and AND3_1198 ( U3546 , U3378 , U3270 , U7482 );
and AND3_1199 ( U3547 , U4448 , U2605 , U4388 );
and AND4_1200 ( U3548 , U4469 , U4468 , U4467 , U4466 );
and AND4_1201 ( U3549 , U4473 , U4472 , U4471 , U4470 );
and AND4_1202 ( U3550 , U4477 , U4476 , U4475 , U4474 );
and AND4_1203 ( U3551 , U4481 , U4480 , U4479 , U4478 );
and AND4_1204 ( U3552 , U4452 , U4451 , U4450 , U4449 );
and AND4_1205 ( U3553 , U4456 , U4455 , U4454 , U4453 );
and AND4_1206 ( U3554 , U4460 , U4459 , U4458 , U4457 );
and AND4_1207 ( U3555 , U4464 , U4463 , U4462 , U4461 );
and AND2_1208 ( U3556 , U4365 , U4196 );
and AND4_1209 ( U3557 , U4407 , U4406 , U4405 , U4404 );
and AND4_1210 ( U3558 , U4411 , U4410 , U4409 , U4408 );
and AND4_1211 ( U3559 , U4415 , U4414 , U4413 , U4412 );
and AND4_1212 ( U3560 , U4419 , U4418 , U4417 , U4416 );
and AND4_1213 ( U3561 , U4392 , U4391 , U4390 , U4389 );
and AND4_1214 ( U3562 , U4396 , U4395 , U4394 , U4393 );
and AND4_1215 ( U3563 , U4400 , U4399 , U4398 , U4397 );
and AND2_1216 ( U3564 , U4402 , U4401 );
and AND2_1217 ( U3565 , U4387 , U4159 );
and AND2_1218 ( U3566 , U4237 , U3270 );
and AND4_1219 ( U3567 , U3271 , U3270 , U4388 , U7482 );
and AND2_1220 ( U3568 , U4205 , U3387 );
and AND2_1221 ( U3569 , STATE2_REG_2_ , U7591 );
and AND2_1222 ( U3570 , U4503 , U3284 );
and AND2_1223 ( U3571 , U2427 , U3244 );
and AND2_1224 ( U3572 , STATE2_REG_3_ , STATE2_REG_0_ );
and AND2_1225 ( U3573 , U4234 , U4229 );
and AND2_1226 ( U3574 , U3573 , U4511 );
and AND3_1227 ( U3575 , U4540 , U4541 , U4212 );
and AND3_1228 ( U3576 , U4549 , U4548 , U4550 );
and AND3_1229 ( U3577 , U4554 , U4553 , U4555 );
and AND3_1230 ( U3578 , U4559 , U4558 , U4560 );
and AND3_1231 ( U3579 , U4564 , U4563 , U4565 );
and AND3_1232 ( U3580 , U4569 , U4568 , U4570 );
and AND3_1233 ( U3581 , U4574 , U4573 , U4575 );
and AND3_1234 ( U3582 , U4579 , U4578 , U4580 );
and AND3_1235 ( U3583 , U4584 , U4583 , U4585 );
and AND3_1236 ( U3584 , U4598 , U4599 , U4212 );
and AND3_1237 ( U3585 , U4607 , U4606 , U4608 );
and AND3_1238 ( U3586 , U4612 , U4611 , U4613 );
and AND3_1239 ( U3587 , U4617 , U4616 , U4618 );
and AND3_1240 ( U3588 , U4622 , U4621 , U4623 );
and AND3_1241 ( U3589 , U4627 , U4626 , U4628 );
and AND3_1242 ( U3590 , U4632 , U4631 , U4633 );
and AND3_1243 ( U3591 , U4637 , U4636 , U4638 );
and AND3_1244 ( U3592 , U4642 , U4641 , U4643 );
and AND3_1245 ( U3593 , U4657 , U4658 , U4212 );
and AND3_1246 ( U3594 , U4666 , U4665 , U4667 );
and AND3_1247 ( U3595 , U4671 , U4670 , U4672 );
and AND3_1248 ( U3596 , U4676 , U4675 , U4677 );
and AND3_1249 ( U3597 , U4681 , U4680 , U4682 );
and AND3_1250 ( U3598 , U4686 , U4685 , U4687 );
and AND3_1251 ( U3599 , U4691 , U4690 , U4692 );
and AND3_1252 ( U3600 , U4696 , U4695 , U4697 );
and AND3_1253 ( U3601 , U4701 , U4700 , U4702 );
and AND3_1254 ( U3602 , U4714 , U4715 , U4212 );
and AND3_1255 ( U3603 , U4723 , U4722 , U4724 );
and AND3_1256 ( U3604 , U4728 , U4727 , U4729 );
and AND3_1257 ( U3605 , U4733 , U4732 , U4734 );
and AND3_1258 ( U3606 , U4738 , U4737 , U4739 );
and AND3_1259 ( U3607 , U4743 , U4742 , U4744 );
and AND3_1260 ( U3608 , U4748 , U4747 , U4749 );
and AND3_1261 ( U3609 , U4753 , U4752 , U4754 );
and AND3_1262 ( U3610 , U4758 , U4757 , U4759 );
and AND3_1263 ( U3611 , U4772 , U4773 , U4212 );
and AND3_1264 ( U3612 , U4781 , U4780 , U4782 );
and AND3_1265 ( U3613 , U4786 , U4785 , U4787 );
and AND3_1266 ( U3614 , U4791 , U4790 , U4792 );
and AND3_1267 ( U3615 , U4796 , U4795 , U4797 );
and AND3_1268 ( U3616 , U4801 , U4800 , U4802 );
and AND3_1269 ( U3617 , U4806 , U4805 , U4807 );
and AND3_1270 ( U3618 , U4811 , U4810 , U4812 );
and AND3_1271 ( U3619 , U4816 , U4815 , U4817 );
and AND3_1272 ( U3620 , U4829 , U4830 , U4212 );
and AND3_1273 ( U3621 , U4838 , U4837 , U4839 );
and AND3_1274 ( U3622 , U4843 , U4842 , U4844 );
and AND3_1275 ( U3623 , U4848 , U4847 , U4849 );
and AND3_1276 ( U3624 , U4853 , U4852 , U4854 );
and AND3_1277 ( U3625 , U4858 , U4857 , U4859 );
and AND3_1278 ( U3626 , U4863 , U4862 , U4864 );
and AND3_1279 ( U3627 , U4868 , U4867 , U4869 );
and AND3_1280 ( U3628 , U4873 , U4872 , U4874 );
and AND3_1281 ( U3629 , U4887 , U4888 , U4212 );
and AND3_1282 ( U3630 , U4896 , U4895 , U4897 );
and AND3_1283 ( U3631 , U4901 , U4900 , U4902 );
and AND3_1284 ( U3632 , U4906 , U4905 , U4907 );
and AND3_1285 ( U3633 , U4911 , U4910 , U4912 );
and AND3_1286 ( U3634 , U4916 , U4915 , U4917 );
and AND3_1287 ( U3635 , U4921 , U4920 , U4922 );
and AND3_1288 ( U3636 , U4926 , U4925 , U4927 );
and AND3_1289 ( U3637 , U4931 , U4930 , U4932 );
and AND3_1290 ( U3638 , U4944 , U4945 , U4212 );
and AND3_1291 ( U3639 , U4953 , U4952 , U4954 );
and AND3_1292 ( U3640 , U4958 , U4957 , U4959 );
and AND3_1293 ( U3641 , U4963 , U4962 , U4964 );
and AND3_1294 ( U3642 , U4968 , U4967 , U4969 );
and AND3_1295 ( U3643 , U4973 , U4972 , U4974 );
and AND3_1296 ( U3644 , U4978 , U4977 , U4979 );
and AND3_1297 ( U3645 , U4983 , U4982 , U4984 );
and AND3_1298 ( U3646 , U4988 , U4987 , U4989 );
and AND3_1299 ( U3647 , U5000 , U5001 , U4212 );
and AND3_1300 ( U3648 , U5009 , U5008 , U5010 );
and AND3_1301 ( U3649 , U5014 , U5013 , U5015 );
and AND3_1302 ( U3650 , U5019 , U5018 , U5020 );
and AND3_1303 ( U3651 , U5024 , U5023 , U5025 );
and AND3_1304 ( U3652 , U5029 , U5028 , U5030 );
and AND3_1305 ( U3653 , U5034 , U5033 , U5035 );
and AND3_1306 ( U3654 , U5039 , U5038 , U5040 );
and AND3_1307 ( U3655 , U5044 , U5043 , U5045 );
and AND3_1308 ( U3656 , U5057 , U5058 , U4212 );
and AND3_1309 ( U3657 , U5066 , U5065 , U5067 );
and AND3_1310 ( U3658 , U5071 , U5070 , U5072 );
and AND3_1311 ( U3659 , U5076 , U5075 , U5077 );
and AND3_1312 ( U3660 , U5081 , U5080 , U5082 );
and AND3_1313 ( U3661 , U5086 , U5085 , U5087 );
and AND3_1314 ( U3662 , U5091 , U5090 , U5092 );
and AND3_1315 ( U3663 , U5096 , U5095 , U5097 );
and AND3_1316 ( U3664 , U5101 , U5100 , U5102 );
and AND3_1317 ( U3665 , U5115 , U5116 , U4212 );
and AND3_1318 ( U3666 , U5124 , U5123 , U5125 );
and AND3_1319 ( U3667 , U5129 , U5128 , U5130 );
and AND3_1320 ( U3668 , U5134 , U5133 , U5135 );
and AND3_1321 ( U3669 , U5139 , U5138 , U5140 );
and AND3_1322 ( U3670 , U5144 , U5143 , U5145 );
and AND3_1323 ( U3671 , U5149 , U5148 , U5150 );
and AND3_1324 ( U3672 , U5154 , U5153 , U5155 );
and AND3_1325 ( U3673 , U5159 , U5158 , U5160 );
and AND3_1326 ( U3674 , U5172 , U5173 , U4212 );
and AND3_1327 ( U3675 , U5181 , U5180 , U5182 );
and AND3_1328 ( U3676 , U5186 , U5185 , U5187 );
and AND3_1329 ( U3677 , U5191 , U5190 , U5192 );
and AND3_1330 ( U3678 , U5196 , U5195 , U5197 );
and AND3_1331 ( U3679 , U5201 , U5200 , U5202 );
and AND3_1332 ( U3680 , U5206 , U5205 , U5207 );
and AND3_1333 ( U3681 , U5211 , U5210 , U5212 );
and AND3_1334 ( U3682 , U5216 , U5215 , U5217 );
and AND3_1335 ( U3683 , U5230 , U5231 , U4212 );
and AND3_1336 ( U3684 , U5239 , U5238 , U5240 );
and AND3_1337 ( U3685 , U5244 , U5243 , U5245 );
and AND3_1338 ( U3686 , U5249 , U5248 , U5250 );
and AND3_1339 ( U3687 , U5254 , U5253 , U5255 );
and AND3_1340 ( U3688 , U5259 , U5258 , U5260 );
and AND3_1341 ( U3689 , U5264 , U5263 , U5265 );
and AND3_1342 ( U3690 , U5269 , U5268 , U5270 );
and AND3_1343 ( U3691 , U5274 , U5273 , U5275 );
and AND3_1344 ( U3692 , U5287 , U5288 , U4212 );
and AND3_1345 ( U3693 , U5296 , U5295 , U5297 );
and AND3_1346 ( U3694 , U5301 , U5300 , U5302 );
and AND3_1347 ( U3695 , U5306 , U5305 , U5307 );
and AND3_1348 ( U3696 , U5311 , U5310 , U5312 );
and AND3_1349 ( U3697 , U5316 , U5315 , U5317 );
and AND3_1350 ( U3698 , U5321 , U5320 , U5322 );
and AND3_1351 ( U3699 , U5326 , U5325 , U5327 );
and AND3_1352 ( U3700 , U5331 , U5330 , U5332 );
and AND3_1353 ( U3701 , U5345 , U5346 , U4212 );
and AND3_1354 ( U3702 , U5354 , U5353 , U5355 );
and AND3_1355 ( U3703 , U5359 , U5358 , U5360 );
and AND3_1356 ( U3704 , U5364 , U5363 , U5365 );
and AND3_1357 ( U3705 , U5369 , U5368 , U5370 );
and AND3_1358 ( U3706 , U5374 , U5373 , U5375 );
and AND3_1359 ( U3707 , U5379 , U5378 , U5380 );
and AND3_1360 ( U3708 , U5384 , U5383 , U5385 );
and AND3_1361 ( U3709 , U5389 , U5388 , U5390 );
and AND3_1362 ( U3710 , U5402 , U5403 , U4212 );
and AND3_1363 ( U3711 , U5411 , U5410 , U5412 );
and AND3_1364 ( U3712 , U5416 , U5415 , U5417 );
and AND3_1365 ( U3713 , U5421 , U5420 , U5422 );
and AND3_1366 ( U3714 , U5426 , U5425 , U5427 );
and AND3_1367 ( U3715 , U5430 , U5429 , U5431 );
and AND3_1368 ( U3716 , U5435 , U5434 , U5436 );
and AND3_1369 ( U3717 , U5440 , U5439 , U5441 );
and AND3_1370 ( U3718 , U5445 , U5444 , U5446 );
and AND2_1371 ( U3719 , FLUSH_REG , STATE2_REG_0_ );
and AND2_1372 ( U3720 , U4482 , U4387 );
and AND2_1373 ( U3721 , U4485 , U3244 );
and AND2_1374 ( U3722 , U4198 , U3244 );
and AND2_1375 ( U3723 , U7484 , U4205 );
and AND2_1376 ( U3724 , U5459 , U5460 );
and AND2_1377 ( U3725 , U3724 , U5458 );
and AND2_1378 ( U3726 , U3725 , U2518 );
and AND2_1379 ( U3727 , U5463 , U4230 );
and AND2_1380 ( U3728 , U5474 , U5473 );
and AND2_1381 ( U3729 , U4437 , U4388 );
and AND2_1382 ( U3730 , U5484 , U3380 );
and AND2_1383 ( U3731 , U5486 , U5485 );
and AND4_1384 ( U3732 , U5488 , U7615 , U3730 , U3731 );
and AND2_1385 ( U3733 , U4251 , U3384 );
and AND5_1386 ( U3734 , U3398 , U3275 , U3733 , U2520 , U3266 );
and AND2_1387 ( U3735 , U3736 , U5490 );
and AND2_1388 ( U3736 , U5493 , U5492 );
and AND3_1389 ( U3737 , U7705 , U7704 , U5501 );
and AND2_1390 ( U3738 , U5512 , U5510 );
and AND2_1391 ( U3739 , U5531 , U5532 );
and AND2_1392 ( U3740 , U5535 , U5536 );
and AND2_1393 ( U3741 , U5540 , U5541 );
and AND2_1394 ( U3742 , U5546 , U3244 );
and AND2_1395 ( U3743 , U3271 , U3394 );
and AND2_1396 ( U3744 , U5551 , U5549 );
and AND3_1397 ( U3745 , U3385 , U3386 , U5555 );
and AND3_1398 ( U3746 , U2520 , U5556 , U3745 );
and AND2_1399 ( U3747 , U4174 , U3271 );
and AND3_1400 ( U3748 , U3275 , U4205 , U3435 );
and AND2_1401 ( U3749 , U5554 , U7495 );
and AND2_1402 ( U3750 , U7496 , STATE2_REG_2_ );
and AND2_1403 ( U3751 , U5559 , U5558 );
and AND2_1404 ( U3752 , U5561 , U5560 );
and AND2_1405 ( U3753 , U5563 , U5564 );
and AND2_1406 ( U3754 , U3753 , U5562 );
and AND2_1407 ( U3755 , U5566 , U5565 );
and AND2_1408 ( U3756 , U5568 , U5567 );
and AND2_1409 ( U3757 , U5570 , U5571 );
and AND2_1410 ( U3758 , U3757 , U5569 );
and AND2_1411 ( U3759 , U5573 , U5572 );
and AND2_1412 ( U3760 , U5575 , U5574 );
and AND2_1413 ( U3761 , U5577 , U5578 );
and AND2_1414 ( U3762 , U3761 , U5576 );
and AND3_1415 ( U3763 , U5580 , U5579 , U5582 );
and AND3_1416 ( U3764 , U3765 , U5583 , U5581 );
and AND2_1417 ( U3765 , U5584 , U5585 );
and AND3_1418 ( U3766 , U5587 , U5586 , U5589 );
and AND2_1419 ( U3767 , U5591 , U5592 );
and AND2_1420 ( U3768 , U3767 , U5590 );
and AND3_1421 ( U3769 , U5594 , U5593 , U5596 );
and AND2_1422 ( U3770 , U5598 , U5599 );
and AND2_1423 ( U3771 , U3770 , U5597 );
and AND3_1424 ( U3772 , U5601 , U5600 , U5603 );
and AND2_1425 ( U3773 , U5605 , U5606 );
and AND2_1426 ( U3774 , U3773 , U5604 );
and AND3_1427 ( U3775 , U5608 , U5607 , U5610 );
and AND2_1428 ( U3776 , U5612 , U5613 );
and AND2_1429 ( U3777 , U3776 , U5611 );
and AND3_1430 ( U3778 , U5615 , U5614 , U5617 );
and AND2_1431 ( U3779 , U5619 , U5620 );
and AND2_1432 ( U3780 , U3779 , U5618 );
and AND3_1433 ( U3781 , U5622 , U5621 , U5624 );
and AND2_1434 ( U3782 , U5626 , U5627 );
and AND2_1435 ( U3783 , U3782 , U5625 );
and AND3_1436 ( U3784 , U5629 , U5628 , U5631 );
and AND2_1437 ( U3785 , U5633 , U5634 );
and AND2_1438 ( U3786 , U3785 , U5632 );
and AND3_1439 ( U3787 , U5636 , U5635 , U5638 );
and AND2_1440 ( U3788 , U5640 , U5641 );
and AND2_1441 ( U3789 , U3788 , U5639 );
and AND3_1442 ( U3790 , U5643 , U5642 , U5645 );
and AND2_1443 ( U3791 , U5647 , U5648 );
and AND2_1444 ( U3792 , U3791 , U5646 );
and AND2_1445 ( U3793 , U5650 , U5652 );
and AND2_1446 ( U3794 , U5654 , U5655 );
and AND2_1447 ( U3795 , U3794 , U5653 );
and AND2_1448 ( U3796 , U5657 , U5659 );
and AND2_1449 ( U3797 , U5661 , U5662 );
and AND2_1450 ( U3798 , U3797 , U5660 );
and AND2_1451 ( U3799 , U5664 , U5666 );
and AND2_1452 ( U3800 , U5668 , U5669 );
and AND2_1453 ( U3801 , U3800 , U5667 );
and AND2_1454 ( U3802 , U5671 , U5673 );
and AND2_1455 ( U3803 , U5675 , U5676 );
and AND2_1456 ( U3804 , U3803 , U5674 );
and AND2_1457 ( U3805 , U5678 , U5680 );
and AND2_1458 ( U3806 , U5682 , U5683 );
and AND2_1459 ( U3807 , U3806 , U5681 );
and AND2_1460 ( U3808 , U5685 , U5687 );
and AND2_1461 ( U3809 , U5689 , U5690 );
and AND2_1462 ( U3810 , U3809 , U5688 );
and AND2_1463 ( U3811 , U5692 , U5694 );
and AND2_1464 ( U3812 , U5696 , U5697 );
and AND2_1465 ( U3813 , U3812 , U5695 );
and AND2_1466 ( U3814 , U5699 , U5701 );
and AND2_1467 ( U3815 , U5703 , U5704 );
and AND2_1468 ( U3816 , U3815 , U5702 );
and AND2_1469 ( U3817 , U5706 , U5708 );
and AND2_1470 ( U3818 , U5710 , U5711 );
and AND2_1471 ( U3819 , U3818 , U5709 );
and AND2_1472 ( U3820 , U5713 , U5715 );
and AND2_1473 ( U3821 , U5717 , U5718 );
and AND2_1474 ( U3822 , U3821 , U5716 );
and AND2_1475 ( U3823 , U5720 , U5722 );
and AND2_1476 ( U3824 , U5724 , U5725 );
and AND2_1477 ( U3825 , U3824 , U5723 );
and AND2_1478 ( U3826 , U5727 , U5729 );
and AND2_1479 ( U3827 , U5731 , U5732 );
and AND2_1480 ( U3828 , U3827 , U5730 );
and AND2_1481 ( U3829 , U5734 , U5736 );
and AND2_1482 ( U3830 , U5738 , U5739 );
and AND2_1483 ( U3831 , U3830 , U5737 );
and AND2_1484 ( U3832 , U5741 , U5743 );
and AND2_1485 ( U3833 , U5745 , U5746 );
and AND2_1486 ( U3834 , U3833 , U5744 );
and AND2_1487 ( U3835 , U5748 , U5750 );
and AND2_1488 ( U3836 , U5752 , U5753 );
and AND2_1489 ( U3837 , U3836 , U5751 );
and AND2_1490 ( U3838 , U5755 , U5757 );
and AND2_1491 ( U3839 , U5759 , U5760 );
and AND2_1492 ( U3840 , U3839 , U5758 );
and AND2_1493 ( U3841 , U5762 , U5764 );
and AND2_1494 ( U3842 , U5766 , U5767 );
and AND2_1495 ( U3843 , U3842 , U5765 );
and AND2_1496 ( U3844 , U5769 , U5771 );
and AND2_1497 ( U3845 , U5773 , U5774 );
and AND2_1498 ( U3846 , U3845 , U5772 );
and AND2_1499 ( U3847 , U5776 , U5778 );
and AND2_1500 ( U3848 , U5780 , U5781 );
and AND2_1501 ( U3849 , U3848 , U5779 );
and AND3_1502 ( U3850 , U3270 , U3249 , U7482 );
and AND2_1503 ( U3851 , U5782 , U3395 );
and AND2_1504 ( U3852 , STATE2_REG_1_ , STATEBS16_REG );
and AND2_1505 ( U3853 , U2368 , U3271 );
and AND2_1506 ( U3854 , U2449 , STATE2_REG_0_ );
and AND2_1507 ( U3855 , U4196 , U2368 );
and AND2_1508 ( U3856 , U6093 , U6094 );
and AND2_1509 ( U3857 , U6096 , U6097 );
and AND2_1510 ( U3858 , U6099 , U6100 );
and AND2_1511 ( U3859 , U6102 , U6103 );
and AND2_1512 ( U3860 , U6105 , U6106 );
and AND2_1513 ( U3861 , U6108 , U6109 );
and AND2_1514 ( U3862 , U6111 , U6112 );
and AND2_1515 ( U3863 , U6114 , U6115 );
and AND2_1516 ( U3864 , U6117 , U6118 );
and AND2_1517 ( U3865 , U6120 , U6121 );
and AND2_1518 ( U3866 , U6123 , U6124 );
and AND2_1519 ( U3867 , U6126 , U6127 );
and AND2_1520 ( U3868 , U6129 , U6130 );
and AND2_1521 ( U3869 , U6132 , U6133 );
and AND2_1522 ( U3870 , U6135 , U6136 );
and AND2_1523 ( U3871 , U6139 , U6138 );
and AND2_1524 ( U3872 , U2605 , U3378 );
and AND3_1525 ( U3873 , STATE2_REG_0_ , U3258 , U7482 );
and AND2_1526 ( U3874 , U4387 , U4159 );
and AND3_1527 ( U3875 , U4229 , U4232 , U6350 );
nor nor_1528 ( U3876 , READY_N , STATEBS16_REG );
and AND2_1529 ( U3877 , U4482 , U4174 );
and AND5_1530 ( U3878 , U6361 , U6360 , U6363 , U6362 , U6359 );
and AND5_1531 ( U3879 , U6369 , U6368 , U6371 , U6370 , U6367 );
and AND5_1532 ( U3880 , U6377 , U6376 , U6379 , U6378 , U6375 );
and AND5_1533 ( U3881 , U6385 , U6384 , U6387 , U6386 , U6383 );
and AND2_1534 ( U3882 , U6388 , U4215 );
and AND4_1535 ( U3883 , U6393 , U6392 , U6395 , U6394 );
and AND2_1536 ( U3884 , U6396 , U4215 );
and AND5_1537 ( U3885 , U6401 , U6400 , U6403 , U6402 , U6399 );
and AND2_1538 ( U3886 , U6404 , U4215 );
and AND3_1539 ( U3887 , U6410 , U6407 , U6409 );
and AND2_1540 ( U3888 , U6411 , U4215 );
and AND3_1541 ( U3889 , U6417 , U6414 , U6416 );
and AND2_1542 ( U3890 , U6418 , U4215 );
and AND3_1543 ( U3891 , U6424 , U6421 , U6423 );
and AND2_1544 ( U3892 , U6425 , U4215 );
and AND3_1545 ( U3893 , U6431 , U6428 , U6430 );
and AND2_1546 ( U3894 , U6432 , U4215 );
and AND3_1547 ( U3895 , U6438 , U6435 , U6437 );
and AND2_1548 ( U3896 , U6439 , U4215 );
and AND3_1549 ( U3897 , U6445 , U6442 , U6444 );
and AND2_1550 ( U3898 , U6446 , U4215 );
and AND3_1551 ( U3899 , U6452 , U6449 , U6451 );
and AND2_1552 ( U3900 , U6453 , U4215 );
and AND3_1553 ( U3901 , U6459 , U6456 , U6458 );
and AND2_1554 ( U3902 , U6460 , U4215 );
and AND3_1555 ( U3903 , U6466 , U6463 , U6465 );
and AND2_1556 ( U3904 , U6467 , U4215 );
and AND3_1557 ( U3905 , U6473 , U6470 , U6472 );
and AND2_1558 ( U3906 , U6474 , U4215 );
and AND3_1559 ( U3907 , U6480 , U6477 , U6479 );
and AND2_1560 ( U3908 , U4215 , U6482 );
and AND3_1561 ( U3909 , U6487 , U6484 , U6486 );
and AND2_1562 ( U3910 , U4215 , U6489 );
and AND3_1563 ( U3911 , U6494 , U6491 , U6493 );
and AND2_1564 ( U3912 , U4215 , U6496 );
and AND3_1565 ( U3913 , U6501 , U6498 , U6500 );
and AND2_1566 ( U3914 , U6505 , U6503 );
and AND2_1567 ( U3915 , U6507 , U6508 );
and AND2_1568 ( U3916 , U6512 , U6510 );
and AND2_1569 ( U3917 , U6514 , U6515 );
and AND2_1570 ( U3918 , U6519 , U6517 );
and AND2_1571 ( U3919 , U6521 , U6522 );
and AND2_1572 ( U3920 , U6526 , U6524 );
and AND2_1573 ( U3921 , U6528 , U6529 );
and AND2_1574 ( U3922 , U6533 , U6531 );
and AND2_1575 ( U3923 , U6535 , U6536 );
and AND2_1576 ( U3924 , U6540 , U6538 );
and AND2_1577 ( U3925 , U6542 , U6543 );
and AND2_1578 ( U3926 , U6547 , U6545 );
and AND2_1579 ( U3927 , U6549 , U6550 );
and AND2_1580 ( U3928 , U6554 , U6552 );
and AND2_1581 ( U3929 , U6556 , U6557 );
and AND2_1582 ( U3930 , U6561 , U6559 );
and AND2_1583 ( U3931 , U6563 , U6564 );
and AND2_1584 ( U3932 , U6568 , U6566 );
and AND2_1585 ( U3933 , U6570 , U6571 );
and AND2_1586 ( U3934 , U6575 , U6573 );
and AND2_1587 ( U3935 , U6577 , U6578 );
and AND2_1588 ( U3936 , U6582 , U6580 );
and AND2_1589 ( U3937 , U6584 , U6585 );
nor nor_1590 ( U3938 , DATAWIDTH_REG_2_ , DATAWIDTH_REG_3_ , DATAWIDTH_REG_4_ , DATAWIDTH_REG_5_ );
nor nor_1591 ( U3939 , DATAWIDTH_REG_6_ , DATAWIDTH_REG_7_ , DATAWIDTH_REG_8_ , DATAWIDTH_REG_9_ );
and AND2_1592 ( U3940 , U3939 , U3938 );
nor nor_1593 ( U3941 , DATAWIDTH_REG_10_ , DATAWIDTH_REG_11_ , DATAWIDTH_REG_12_ , DATAWIDTH_REG_13_ );
nor nor_1594 ( U3942 , DATAWIDTH_REG_14_ , DATAWIDTH_REG_15_ , DATAWIDTH_REG_16_ , DATAWIDTH_REG_17_ );
and AND2_1595 ( U3943 , U3942 , U3941 );
nor nor_1596 ( U3944 , DATAWIDTH_REG_18_ , DATAWIDTH_REG_19_ , DATAWIDTH_REG_20_ , DATAWIDTH_REG_21_ );
nor nor_1597 ( U3945 , DATAWIDTH_REG_22_ , DATAWIDTH_REG_23_ , DATAWIDTH_REG_24_ , DATAWIDTH_REG_25_ );
and AND2_1598 ( U3946 , U3945 , U3944 );
nor nor_1599 ( U3947 , DATAWIDTH_REG_26_ , DATAWIDTH_REG_27_ );
nor nor_1600 ( U3948 , DATAWIDTH_REG_28_ , DATAWIDTH_REG_29_ );
nor nor_1601 ( U3949 , DATAWIDTH_REG_30_ , DATAWIDTH_REG_31_ );
and AND4_1602 ( U3950 , U3949 , U6586 , U3948 , U3947 );
nor nor_1603 ( U3951 , REIP_REG_0_ , DATAWIDTH_REG_0_ , DATAWIDTH_REG_1_ );
and AND2_1604 ( U3952 , STATE2_REG_2_ , U3244 );
and AND2_1605 ( U3953 , U6596 , U3285 );
nor nor_1606 ( U3954 , READY_N , STATE2_REG_0_ );
and AND3_1607 ( U3955 , U3294 , U3395 , U6590 );
and AND2_1608 ( U3956 , STATE2_REG_2_ , U3274 );
and AND2_1609 ( U3957 , U4223 , U4194 );
and AND4_1610 ( U3958 , U6609 , U6608 , U6607 , U6606 );
and AND4_1611 ( U3959 , U6613 , U6612 , U6611 , U6610 );
and AND4_1612 ( U3960 , U6617 , U6616 , U6615 , U6614 );
and AND4_1613 ( U3961 , U6621 , U6620 , U6619 , U6618 );
and AND4_1614 ( U3962 , U6625 , U6624 , U6623 , U6622 );
and AND4_1615 ( U3963 , U6629 , U6628 , U6627 , U6626 );
and AND4_1616 ( U3964 , U6633 , U6632 , U6631 , U6630 );
and AND4_1617 ( U3965 , U6637 , U6636 , U6635 , U6634 );
and AND4_1618 ( U3966 , U6641 , U6640 , U6639 , U6638 );
and AND4_1619 ( U3967 , U6645 , U6644 , U6643 , U6642 );
and AND4_1620 ( U3968 , U6649 , U6648 , U6647 , U6646 );
and AND4_1621 ( U3969 , U6653 , U6652 , U6651 , U6650 );
and AND4_1622 ( U3970 , U6657 , U6656 , U6655 , U6654 );
and AND4_1623 ( U3971 , U6661 , U6660 , U6659 , U6658 );
and AND4_1624 ( U3972 , U6665 , U6664 , U6663 , U6662 );
and AND4_1625 ( U3973 , U7601 , U6668 , U6667 , U6666 );
and AND4_1626 ( U3974 , U6672 , U6671 , U6670 , U6669 );
and AND4_1627 ( U3975 , U6676 , U6675 , U6674 , U6673 );
and AND4_1628 ( U3976 , U6680 , U6679 , U6678 , U6677 );
and AND4_1629 ( U3977 , U6684 , U6683 , U6682 , U6681 );
and AND4_1630 ( U3978 , U6688 , U6687 , U6686 , U6685 );
and AND4_1631 ( U3979 , U6692 , U6691 , U6690 , U6689 );
and AND4_1632 ( U3980 , U6696 , U6695 , U6694 , U6693 );
and AND4_1633 ( U3981 , U6700 , U6699 , U6698 , U6697 );
and AND4_1634 ( U3982 , U6704 , U6703 , U6702 , U6701 );
and AND4_1635 ( U3983 , U6708 , U6707 , U6706 , U6705 );
and AND4_1636 ( U3984 , U6712 , U6711 , U6710 , U6709 );
and AND4_1637 ( U3985 , U6716 , U6715 , U6714 , U6713 );
and AND4_1638 ( U3986 , U6720 , U6719 , U6718 , U6717 );
and AND4_1639 ( U3987 , U6724 , U6723 , U6722 , U6721 );
and AND4_1640 ( U3988 , U6728 , U6727 , U6726 , U6725 );
and AND4_1641 ( U3989 , U6732 , U6731 , U6730 , U6729 );
and AND2_1642 ( U3990 , U6737 , U6736 );
and AND2_1643 ( U3991 , U6740 , U6739 );
and AND2_1644 ( U3992 , U6743 , U6742 );
and AND2_1645 ( U3993 , U6746 , U6745 );
and AND2_1646 ( U3994 , U6748 , U3995 );
and AND2_1647 ( U3995 , U6750 , U6749 );
and AND2_1648 ( U3996 , U6752 , U6753 );
and AND3_1649 ( U3997 , U6760 , U6761 , U6762 );
and AND2_1650 ( U3998 , U6764 , U6765 );
and AND3_1651 ( U3999 , U6769 , U6770 , U6771 );
and AND3_1652 ( U4000 , U6773 , U6774 , U6775 );
and AND3_1653 ( U4001 , U6777 , U6778 , U6779 );
and AND3_1654 ( U4002 , U6781 , U6782 , U6783 );
and AND3_1655 ( U4003 , U6785 , U6786 , U6787 );
and AND3_1656 ( U4004 , U6789 , U6790 , U6791 );
and AND3_1657 ( U4005 , U6793 , U6794 , U6795 );
and AND3_1658 ( U4006 , U6797 , U6798 , U6799 );
and AND3_1659 ( U4007 , U6801 , U6802 , U6803 );
and AND3_1660 ( U4008 , U6805 , U6806 , U6807 );
and AND2_1661 ( U4009 , U6809 , U6810 );
and AND3_1662 ( U4010 , U6814 , U6815 , U6816 );
and AND3_1663 ( U4011 , U6818 , U6819 , U6820 );
and AND3_1664 ( U4012 , U6822 , U6823 , U6824 );
and AND3_1665 ( U4013 , U6826 , U6827 , U6828 );
and AND2_1666 ( U4014 , U6846 , U6845 );
and AND2_1667 ( U4015 , U6848 , U6849 );
and AND3_1668 ( U4016 , U7482 , U6876 , U3270 );
and AND4_1669 ( U4017 , U6883 , U6882 , U6881 , U6880 );
and AND4_1670 ( U4018 , U6887 , U6886 , U6885 , U6884 );
and AND4_1671 ( U4019 , U6891 , U6890 , U6889 , U6888 );
and AND4_1672 ( U4020 , U6895 , U6894 , U6893 , U6892 );
and AND4_1673 ( U4021 , U6901 , U6900 , U6899 , U6898 );
and AND4_1674 ( U4022 , U6905 , U6904 , U6903 , U6902 );
and AND4_1675 ( U4023 , U6909 , U6908 , U6907 , U6906 );
and AND4_1676 ( U4024 , U6913 , U6912 , U6911 , U6910 );
and AND4_1677 ( U4025 , U6932 , U6931 , U6930 , U6929 );
and AND4_1678 ( U4026 , U6936 , U6935 , U6934 , U6933 );
and AND4_1679 ( U4027 , U6940 , U6939 , U6938 , U6937 );
and AND4_1680 ( U4028 , U6944 , U6943 , U6942 , U6941 );
and AND4_1681 ( U4029 , U6949 , U6948 , U6947 , U6946 );
and AND4_1682 ( U4030 , U6953 , U6952 , U6951 , U6950 );
and AND4_1683 ( U4031 , U6957 , U6956 , U6955 , U6954 );
and AND4_1684 ( U4032 , U6961 , U6960 , U6959 , U6958 );
and AND4_1685 ( U4033 , U6966 , U6965 , U6964 , U6963 );
and AND4_1686 ( U4034 , U6970 , U6969 , U6968 , U6967 );
and AND4_1687 ( U4035 , U6974 , U6973 , U6972 , U6971 );
and AND4_1688 ( U4036 , U6978 , U6977 , U6976 , U6975 );
and AND4_1689 ( U4037 , U6983 , U6982 , U6981 , U6980 );
and AND4_1690 ( U4038 , U6987 , U6986 , U6985 , U6984 );
and AND4_1691 ( U4039 , U6991 , U6990 , U6989 , U6988 );
and AND4_1692 ( U4040 , U7602 , U6994 , U6993 , U6992 );
and AND4_1693 ( U4041 , U6998 , U6997 , U6996 , U6995 );
and AND4_1694 ( U4042 , U7002 , U7001 , U7000 , U6999 );
and AND4_1695 ( U4043 , U7006 , U7005 , U7004 , U7003 );
and AND4_1696 ( U4044 , U7010 , U7009 , U7008 , U7007 );
and AND4_1697 ( U4045 , U7015 , U7014 , U7013 , U7012 );
and AND4_1698 ( U4046 , U7019 , U7018 , U7017 , U7016 );
and AND4_1699 ( U4047 , U7023 , U7022 , U7021 , U7020 );
and AND4_1700 ( U4048 , U7027 , U7026 , U7025 , U7024 );
and AND2_1701 ( U4049 , U7047 , U3430 );
and AND2_1702 ( U4050 , STATE2_REG_0_ , U7050 );
and AND4_1703 ( U4051 , U7057 , U7056 , U7055 , U7054 );
and AND4_1704 ( U4052 , U7061 , U7060 , U7059 , U7058 );
and AND4_1705 ( U4053 , U7065 , U7064 , U7063 , U7062 );
and AND4_1706 ( U4054 , U7069 , U7068 , U7067 , U7066 );
and AND2_1707 ( U4055 , U4244 , STATE2_REG_0_ );
and AND4_1708 ( U4056 , U4393 , U4392 , U4391 , U4389 );
and AND3_1709 ( U4057 , U4395 , U4394 , U4396 );
and AND4_1710 ( U4058 , U4400 , U4399 , U4398 , U4397 );
and AND2_1711 ( U4059 , U4402 , U4401 );
and AND2_1712 ( U4060 , U4388 , U3378 );
and AND2_1713 ( U4061 , STATE2_REG_0_ , U3271 );
and AND2_1714 ( U4062 , U7078 , U7077 );
and AND3_1715 ( U4063 , U7460 , U3421 , U7461 );
and AND3_1716 ( U4064 , U7463 , U7464 , U7462 );
and AND3_1717 ( U4065 , U2606 , U7465 , U4064 );
and AND2_1718 ( U4066 , U7085 , U7083 );
and AND4_1719 ( U4067 , U7089 , U7088 , U7087 , U7086 );
and AND4_1720 ( U4068 , U7093 , U7092 , U7091 , U7090 );
and AND4_1721 ( U4069 , U7097 , U7096 , U7095 , U7094 );
and AND4_1722 ( U4070 , U7101 , U7100 , U7099 , U7098 );
and AND4_1723 ( U4071 , U7106 , U7105 , U7104 , U7103 );
and AND4_1724 ( U4072 , U7110 , U7109 , U7108 , U7107 );
and AND4_1725 ( U4073 , U7114 , U7113 , U7112 , U7111 );
and AND4_1726 ( U4074 , U7118 , U7117 , U7116 , U7115 );
and AND4_1727 ( U4075 , U7123 , U7122 , U7121 , U7120 );
and AND4_1728 ( U4076 , U7127 , U7126 , U7125 , U7124 );
and AND4_1729 ( U4077 , U7131 , U7130 , U7129 , U7128 );
and AND2_1730 ( U4078 , U7133 , U7132 );
and AND3_1731 ( U4079 , U7605 , U7134 , U4078 );
and AND4_1732 ( U4080 , U7138 , U7137 , U7136 , U7135 );
and AND4_1733 ( U4081 , U7142 , U7141 , U7140 , U7139 );
and AND4_1734 ( U4082 , U7146 , U7145 , U7144 , U7143 );
and AND4_1735 ( U4083 , U7150 , U7149 , U7148 , U7147 );
and AND4_1736 ( U4084 , U7155 , U7154 , U7153 , U7152 );
and AND4_1737 ( U4085 , U7159 , U7158 , U7157 , U7156 );
and AND4_1738 ( U4086 , U7163 , U7162 , U7161 , U7160 );
and AND4_1739 ( U4087 , U7167 , U7166 , U7165 , U7164 );
and AND4_1740 ( U4088 , U7172 , U7171 , U7170 , U7169 );
and AND4_1741 ( U4089 , U7176 , U7175 , U7174 , U7173 );
and AND4_1742 ( U4090 , U7180 , U7179 , U7178 , U7177 );
and AND4_1743 ( U4091 , U7184 , U7183 , U7182 , U7181 );
and AND4_1744 ( U4092 , U7189 , U7188 , U7187 , U7186 );
and AND4_1745 ( U4093 , U7193 , U7192 , U7191 , U7190 );
and AND4_1746 ( U4094 , U7197 , U7196 , U7195 , U7194 );
and AND4_1747 ( U4095 , U7201 , U7200 , U7199 , U7198 );
and AND2_1748 ( U4096 , U7203 , U3251 );
and AND2_1749 ( U4097 , U7204 , U7203 );
and AND2_1750 ( U4098 , U7205 , U3252 );
and AND2_1751 ( U4099 , U7077 , U3414 );
and AND2_1752 ( U4100 , U7206 , U7205 );
and AND3_1753 ( U4101 , U4100 , U7460 , U7461 );
and AND4_1754 ( U4102 , U7078 , U3421 , U4099 , U4101 );
and AND4_1755 ( U4103 , U7474 , U7468 , U7464 , U7462 );
and AND4_1756 ( U4104 , U7493 , U7477 , U7476 , U7475 );
and AND2_1757 ( U4105 , U7078 , U7077 );
and AND3_1758 ( U4106 , U7460 , U3421 , U7461 );
and AND3_1759 ( U4107 , U7463 , U7464 , U7462 );
and AND4_1760 ( U4108 , U2608 , U7465 , U2606 , U4107 );
and AND4_1761 ( U4109 , U7211 , U7210 , U7209 , U7208 );
and AND4_1762 ( U4110 , U7215 , U7214 , U7213 , U7212 );
and AND4_1763 ( U4111 , U7219 , U7218 , U7217 , U7216 );
and AND4_1764 ( U4112 , U7223 , U7222 , U7221 , U7220 );
and AND4_1765 ( U4113 , U7228 , U7227 , U7226 , U7225 );
and AND4_1766 ( U4114 , U7232 , U7231 , U7230 , U7229 );
and AND4_1767 ( U4115 , U7236 , U7235 , U7234 , U7233 );
and AND4_1768 ( U4116 , U7240 , U7239 , U7238 , U7237 );
and AND4_1769 ( U4117 , U7245 , U7244 , U7243 , U7242 );
and AND4_1770 ( U4118 , U7249 , U7248 , U7247 , U7246 );
and AND4_1771 ( U4119 , U7253 , U7252 , U7251 , U7250 );
and AND4_1772 ( U4120 , U7257 , U7256 , U7255 , U7254 );
and AND4_1773 ( U4121 , U7262 , U7261 , U7260 , U7259 );
and AND4_1774 ( U4122 , U7266 , U7265 , U7264 , U7263 );
and AND4_1775 ( U4123 , U7270 , U7269 , U7268 , U7267 );
and AND4_1776 ( U4124 , U7607 , U7273 , U7272 , U7271 );
and AND4_1777 ( U4125 , U7277 , U7276 , U7275 , U7274 );
and AND4_1778 ( U4126 , U7281 , U7280 , U7279 , U7278 );
and AND4_1779 ( U4127 , U7285 , U7284 , U7283 , U7282 );
and AND4_1780 ( U4128 , U7289 , U7288 , U7287 , U7286 );
and AND4_1781 ( U4129 , U7294 , U7293 , U7292 , U7291 );
and AND4_1782 ( U4130 , U7298 , U7297 , U7296 , U7295 );
and AND4_1783 ( U4131 , U7302 , U7301 , U7300 , U7299 );
and AND4_1784 ( U4132 , U7306 , U7305 , U7304 , U7303 );
and AND4_1785 ( U4133 , U7311 , U7310 , U7309 , U7308 );
and AND4_1786 ( U4134 , U7315 , U7314 , U7313 , U7312 );
and AND4_1787 ( U4135 , U7319 , U7318 , U7317 , U7316 );
and AND4_1788 ( U4136 , U7323 , U7322 , U7321 , U7320 );
and AND4_1789 ( U4137 , U7328 , U7327 , U7326 , U7325 );
and AND4_1790 ( U4138 , U7332 , U7331 , U7330 , U7329 );
and AND4_1791 ( U4139 , U7336 , U7335 , U7334 , U7333 );
and AND4_1792 ( U4140 , U7340 , U7339 , U7338 , U7337 );
and AND2_1793 ( U4141 , U3271 , U3406 );
and AND2_1794 ( U4142 , U3270 , U3378 );
and AND3_1795 ( U4143 , U7345 , U7346 , U4251 );
and AND2_1796 ( U4144 , U4143 , U7347 );
and AND2_1797 ( U4145 , STATE2_REG_0_ , U2427 );
and AND2_1798 ( U4146 , U4145 , U7348 );
and AND2_1799 ( U4147 , U3258 , U4161 );
and AND2_1800 ( U4148 , STATE2_REG_0_ , U4161 );
and AND2_1801 ( U4149 , U7357 , STATE2_REG_0_ );
and AND2_1802 ( U4150 , U7359 , U2603 );
and AND2_1803 ( U4151 , U7361 , STATE2_REG_0_ );
and AND2_1804 ( U4152 , U7363 , U2603 );
and AND2_1805 ( U4153 , U7370 , U7371 );
and AND2_1806 ( U4154 , U3440 , U7372 );
and AND3_1807 ( U4155 , U7377 , U7376 , U7375 );
and AND2_1808 ( U4156 , U7450 , U7449 );
and AND2_1809 ( U4157 , U7453 , U7452 );
and AND2_1810 ( U4158 , U7662 , U7661 );
nand NAND4_1811 ( U4159 , U3560 , U3559 , U3558 , U3557 );
nand NAND2_1812 ( U4160 , U3727 , U5462 );
nand NAND5_1813 ( U4161 , U3564 , U2607 , U3563 , U3562 , U3561 );
not NOT1_1814 ( U4162 , INSTADDRPOINTER_REG_31_ );
and AND2_1815 ( U4163 , U7714 , U7713 );
and AND2_1816 ( U4164 , U7733 , U7732 );
nand NAND2_1817 ( U4165 , U2368 , U3272 );
nand NAND2_1818 ( U4166 , U4496 , U3378 );
not NOT1_1819 ( U4167 , BS16_N );
nand NAND2_1820 ( U4168 , U3955 , U4216 );
nand NAND2_1821 ( U4169 , U4216 , U3419 );
nand NAND3_1822 ( U4170 , U7686 , U7685 , U3726 );
nand NAND2_1823 ( U4171 , INSTQUEUERD_ADDR_REG_2_ , U3256 );
not NOT1_1824 ( U4172 , U3439 );
nand NAND2_1825 ( U4173 , HOLD , U3244 );
not NOT1_1826 ( U4174 , U3399 );
not NOT1_1827 ( U4175 , U3427 );
not NOT1_1828 ( U4176 , U3426 );
not NOT1_1829 ( U4177 , U3380 );
not NOT1_1830 ( U4178 , U3277 );
not NOT1_1831 ( U4179 , U3436 );
not NOT1_1832 ( U4180 , U3392 );
not NOT1_1833 ( U4181 , U3421 );
not NOT1_1834 ( U4182 , U3407 );
nand NAND2_1835 ( U4183 , U4253 , U3258 );
nand NAND2_1836 ( U4184 , U4448 , U2605 );
not NOT1_1837 ( U4185 , U3383 );
not NOT1_1838 ( U4186 , U3412 );
not NOT1_1839 ( U4187 , U3276 );
not NOT1_1840 ( U4188 , U3408 );
not NOT1_1841 ( U4189 , U3409 );
not NOT1_1842 ( U4190 , U3415 );
not NOT1_1843 ( U4191 , U3395 );
not NOT1_1844 ( U4192 , U3414 );
nand NAND3_1845 ( U4193 , U3873 , U4177 , U4185 );
not NOT1_1846 ( U4194 , U3405 );
not NOT1_1847 ( U4195 , U3430 );
not NOT1_1848 ( U4196 , U3269 );
not NOT1_1849 ( U4197 , U3294 );
not NOT1_1850 ( U4198 , U3377 );
not NOT1_1851 ( U4199 , U3433 );
not NOT1_1852 ( U4200 , U3434 );
not NOT1_1853 ( U4201 , U3435 );
not NOT1_1854 ( U4202 , U3387 );
not NOT1_1855 ( U4203 , U3275 );
not NOT1_1856 ( U4204 , U3279 );
nand NAND2_1857 ( U4205 , U3566 , U2431 );
not NOT1_1858 ( U4206 , U3386 );
nand NAND2_1859 ( U4207 , U4437 , U3258 );
not NOT1_1860 ( U4208 , U3420 );
not NOT1_1861 ( U4209 , U3236 );
not NOT1_1862 ( U4210 , U3413 );
not NOT1_1863 ( U4211 , U3411 );
not NOT1_1864 ( U4212 , U3287 );
not NOT1_1865 ( U4213 , LT_563_1260_U6 );
not NOT1_1866 ( U4214 , U3307 );
nand NAND2_1867 ( U4215 , U4243 , U3418 );
nand NAND2_1868 ( U4216 , U4223 , U7488 );
nand NAND2_1869 ( U4217 , U2362 , U3259 );
nand NAND2_1870 ( U4218 , U2363 , U4365 );
not NOT1_1871 ( U4219 , U3394 );
not NOT1_1872 ( U4220 , U3239 );
not NOT1_1873 ( U4221 , U3237 );
not NOT1_1874 ( U4222 , U3382 );
not NOT1_1875 ( U4223 , U3284 );
not NOT1_1876 ( U4224 , U3385 );
not NOT1_1877 ( U4225 , U4166 );
not NOT1_1878 ( U4226 , U3344 );
nand NAND2_1879 ( U4227 , U4465 , U7369 );
nand NAND2_1880 ( U4228 , U3951 , U4208 );
nand NAND2_1881 ( U4229 , U3572 , U4249 );
nand NAND2_1882 ( U4230 , U3719 , U2428 );
nand NAND2_1883 ( U4231 , U4352 , U3245 );
nand NAND3_1884 ( U4232 , STATE2_REG_1_ , U3281 , U2352 );
nand NAND2_1885 ( U4233 , U2428 , U3390 );
nand NAND3_1886 ( U4234 , READY_N , U3250 , STATE2_REG_0_ );
not NOT1_1887 ( U4235 , U3381 );
nand NAND4_1888 ( U4236 , U2451 , U2353 , U3850 , U2448 );
not NOT1_1889 ( U4237 , U3274 );
not NOT1_1890 ( U4238 , U3384 );
not NOT1_1891 ( U4239 , U3402 );
not NOT1_1892 ( U4240 , U3286 );
not NOT1_1893 ( U4241 , U3396 );
not NOT1_1894 ( U4242 , U3406 );
not NOT1_1895 ( U4243 , U3419 );
not NOT1_1896 ( U4244 , U3278 );
not NOT1_1897 ( U4245 , U3376 );
not NOT1_1898 ( U4246 , U3241 );
not NOT1_1899 ( U4247 , U3268 );
not NOT1_1900 ( U4248 , U3393 );
not NOT1_1901 ( U4249 , U3285 );
not NOT1_1902 ( U4250 , U3273 );
nand NAND2_1903 ( U4251 , U4224 , U4387 );
not NOT1_1904 ( U4252 , U3398 );
not NOT1_1905 ( U4253 , U3440 );
not NOT1_1906 ( U4254 , U3397 );
nand NAND2_1907 ( U4255 , REIP_REG_31_ , U4221 );
nand NAND2_1908 ( U4256 , REIP_REG_30_ , U4220 );
nand NAND2_1909 ( U4257 , ADDRESS_REG_29_ , U3236 );
nand NAND2_1910 ( U4258 , REIP_REG_30_ , U4221 );
nand NAND2_1911 ( U4259 , REIP_REG_29_ , U4220 );
nand NAND2_1912 ( U4260 , ADDRESS_REG_28_ , U3236 );
nand NAND2_1913 ( U4261 , REIP_REG_29_ , U4221 );
nand NAND2_1914 ( U4262 , REIP_REG_28_ , U4220 );
nand NAND2_1915 ( U4263 , ADDRESS_REG_27_ , U3236 );
nand NAND2_1916 ( U4264 , REIP_REG_28_ , U4221 );
nand NAND2_1917 ( U4265 , REIP_REG_27_ , U4220 );
nand NAND2_1918 ( U4266 , ADDRESS_REG_26_ , U3236 );
nand NAND2_1919 ( U4267 , REIP_REG_27_ , U4221 );
nand NAND2_1920 ( U4268 , REIP_REG_26_ , U4220 );
nand NAND2_1921 ( U4269 , ADDRESS_REG_25_ , U3236 );
nand NAND2_1922 ( U4270 , REIP_REG_26_ , U4221 );
nand NAND2_1923 ( U4271 , REIP_REG_25_ , U4220 );
nand NAND2_1924 ( U4272 , ADDRESS_REG_24_ , U3236 );
nand NAND2_1925 ( U4273 , REIP_REG_25_ , U4221 );
nand NAND2_1926 ( U4274 , REIP_REG_24_ , U4220 );
nand NAND2_1927 ( U4275 , ADDRESS_REG_23_ , U3236 );
nand NAND2_1928 ( U4276 , REIP_REG_24_ , U4221 );
nand NAND2_1929 ( U4277 , REIP_REG_23_ , U4220 );
nand NAND2_1930 ( U4278 , ADDRESS_REG_22_ , U3236 );
nand NAND2_1931 ( U4279 , REIP_REG_23_ , U4221 );
nand NAND2_1932 ( U4280 , REIP_REG_22_ , U4220 );
nand NAND2_1933 ( U4281 , ADDRESS_REG_21_ , U3236 );
nand NAND2_1934 ( U4282 , REIP_REG_22_ , U4221 );
nand NAND2_1935 ( U4283 , REIP_REG_21_ , U4220 );
nand NAND2_1936 ( U4284 , ADDRESS_REG_20_ , U3236 );
nand NAND2_1937 ( U4285 , REIP_REG_21_ , U4221 );
nand NAND2_1938 ( U4286 , REIP_REG_20_ , U4220 );
nand NAND2_1939 ( U4287 , ADDRESS_REG_19_ , U3236 );
nand NAND2_1940 ( U4288 , REIP_REG_20_ , U4221 );
nand NAND2_1941 ( U4289 , REIP_REG_19_ , U4220 );
nand NAND2_1942 ( U4290 , ADDRESS_REG_18_ , U3236 );
nand NAND2_1943 ( U4291 , REIP_REG_19_ , U4221 );
nand NAND2_1944 ( U4292 , REIP_REG_18_ , U4220 );
nand NAND2_1945 ( U4293 , ADDRESS_REG_17_ , U3236 );
nand NAND2_1946 ( U4294 , REIP_REG_18_ , U4221 );
nand NAND2_1947 ( U4295 , REIP_REG_17_ , U4220 );
nand NAND2_1948 ( U4296 , ADDRESS_REG_16_ , U3236 );
nand NAND2_1949 ( U4297 , REIP_REG_17_ , U4221 );
nand NAND2_1950 ( U4298 , REIP_REG_16_ , U4220 );
nand NAND2_1951 ( U4299 , ADDRESS_REG_15_ , U3236 );
nand NAND2_1952 ( U4300 , REIP_REG_16_ , U4221 );
nand NAND2_1953 ( U4301 , REIP_REG_15_ , U4220 );
nand NAND2_1954 ( U4302 , ADDRESS_REG_14_ , U3236 );
nand NAND2_1955 ( U4303 , REIP_REG_15_ , U4221 );
nand NAND2_1956 ( U4304 , REIP_REG_14_ , U4220 );
nand NAND2_1957 ( U4305 , ADDRESS_REG_13_ , U3236 );
nand NAND2_1958 ( U4306 , REIP_REG_14_ , U4221 );
nand NAND2_1959 ( U4307 , REIP_REG_13_ , U4220 );
nand NAND2_1960 ( U4308 , ADDRESS_REG_12_ , U3236 );
nand NAND2_1961 ( U4309 , REIP_REG_13_ , U4221 );
nand NAND2_1962 ( U4310 , REIP_REG_12_ , U4220 );
nand NAND2_1963 ( U4311 , ADDRESS_REG_11_ , U3236 );
nand NAND2_1964 ( U4312 , REIP_REG_12_ , U4221 );
nand NAND2_1965 ( U4313 , REIP_REG_11_ , U4220 );
nand NAND2_1966 ( U4314 , ADDRESS_REG_10_ , U3236 );
nand NAND2_1967 ( U4315 , REIP_REG_11_ , U4221 );
nand NAND2_1968 ( U4316 , REIP_REG_10_ , U4220 );
nand NAND2_1969 ( U4317 , ADDRESS_REG_9_ , U3236 );
nand NAND2_1970 ( U4318 , REIP_REG_10_ , U4221 );
nand NAND2_1971 ( U4319 , REIP_REG_9_ , U4220 );
nand NAND2_1972 ( U4320 , ADDRESS_REG_8_ , U3236 );
nand NAND2_1973 ( U4321 , REIP_REG_9_ , U4221 );
nand NAND2_1974 ( U4322 , REIP_REG_8_ , U4220 );
nand NAND2_1975 ( U4323 , ADDRESS_REG_7_ , U3236 );
nand NAND2_1976 ( U4324 , REIP_REG_8_ , U4221 );
nand NAND2_1977 ( U4325 , REIP_REG_7_ , U4220 );
nand NAND2_1978 ( U4326 , ADDRESS_REG_6_ , U3236 );
nand NAND2_1979 ( U4327 , REIP_REG_7_ , U4221 );
nand NAND2_1980 ( U4328 , REIP_REG_6_ , U4220 );
nand NAND2_1981 ( U4329 , ADDRESS_REG_5_ , U3236 );
nand NAND2_1982 ( U4330 , REIP_REG_6_ , U4221 );
nand NAND2_1983 ( U4331 , REIP_REG_5_ , U4220 );
nand NAND2_1984 ( U4332 , ADDRESS_REG_4_ , U3236 );
nand NAND2_1985 ( U4333 , REIP_REG_5_ , U4221 );
nand NAND2_1986 ( U4334 , REIP_REG_4_ , U4220 );
nand NAND2_1987 ( U4335 , ADDRESS_REG_3_ , U3236 );
nand NAND2_1988 ( U4336 , REIP_REG_4_ , U4221 );
nand NAND2_1989 ( U4337 , REIP_REG_3_ , U4220 );
nand NAND2_1990 ( U4338 , ADDRESS_REG_2_ , U3236 );
nand NAND2_1991 ( U4339 , REIP_REG_3_ , U4221 );
nand NAND2_1992 ( U4340 , REIP_REG_2_ , U4220 );
nand NAND2_1993 ( U4341 , ADDRESS_REG_1_ , U3236 );
nand NAND2_1994 ( U4342 , REIP_REG_2_ , U4221 );
nand NAND2_1995 ( U4343 , REIP_REG_1_ , U4220 );
nand NAND2_1996 ( U4344 , ADDRESS_REG_0_ , U3236 );
not NOT1_1997 ( U4345 , U3247 );
nand NAND2_1998 ( U4346 , U4345 , U3244 );
nand NAND2_1999 ( U4347 , NA_N , U4246 );
not NOT1_2000 ( U4348 , U3248 );
nand NAND2_2001 ( U4349 , U4348 , U3244 );
or OR2_2002 ( U4350 , STATE_REG_0_ , NA_N );
nand NAND3_2003 ( U4351 , U7610 , U4350 , U7611 );
not NOT1_2004 ( U4352 , U3242 );
nand NAND3_2005 ( U4353 , HOLD , U3234 , U4352 );
nand NAND2_2006 ( U4354 , U3481 , U3248 );
nand NAND2_2007 ( U4355 , U4354 , U4353 );
nand NAND3_2008 ( U4356 , STATE_REG_0_ , U4347 , U4355 );
nand NAND2_2009 ( U4357 , STATE_REG_2_ , U4351 );
nand NAND2_2010 ( U4358 , READY_N , U4209 );
nand NAND2_2011 ( U4359 , U3484 , U7613 );
nand NAND2_2012 ( U4360 , STATE_REG_2_ , U3247 );
nand NAND2_2013 ( U4361 , NA_N , U3245 );
nand NAND2_2014 ( U4362 , U4361 , U4360 );
nand NAND2_2015 ( U4363 , U4362 , U3235 );
nand NAND2_2016 ( U4364 , U4167 , U3242 );
not NOT1_2017 ( U4365 , U3267 );
not NOT1_2018 ( U4366 , U3256 );
not NOT1_2019 ( U4367 , U3431 );
not NOT1_2020 ( U4368 , U3255 );
not NOT1_2021 ( U4369 , U3261 );
not NOT1_2022 ( U4370 , U3254 );
nand NAND2_2023 ( U4371 , INSTQUEUE_REG_7__3_ , U4370 );
nand NAND2_2024 ( U4372 , INSTQUEUE_REG_0__3_ , U2472 );
nand NAND2_2025 ( U4373 , INSTQUEUE_REG_1__3_ , U2471 );
nand NAND2_2026 ( U4374 , INSTQUEUE_REG_2__3_ , U2470 );
nand NAND2_2027 ( U4375 , INSTQUEUE_REG_3__3_ , U2468 );
nand NAND2_2028 ( U4376 , INSTQUEUE_REG_4__3_ , U2467 );
nand NAND2_2029 ( U4377 , INSTQUEUE_REG_5__3_ , U2466 );
nand NAND2_2030 ( U4378 , INSTQUEUE_REG_6__3_ , U2465 );
nand NAND2_2031 ( U4379 , INSTQUEUE_REG_8__3_ , U2464 );
nand NAND2_2032 ( U4380 , INSTQUEUE_REG_9__3_ , U2463 );
nand NAND2_2033 ( U4381 , INSTQUEUE_REG_10__3_ , U2461 );
nand NAND2_2034 ( U4382 , INSTQUEUE_REG_11__3_ , U2459 );
nand NAND2_2035 ( U4383 , INSTQUEUE_REG_12__3_ , U2458 );
nand NAND2_2036 ( U4384 , INSTQUEUE_REG_13__3_ , U2457 );
nand NAND2_2037 ( U4385 , INSTQUEUE_REG_14__3_ , U2455 );
nand NAND2_2038 ( U4386 , INSTQUEUE_REG_15__3_ , U2453 );
not NOT1_2039 ( U4387 , U3270 );
not NOT1_2040 ( U4388 , U3265 );
nand NAND5_2041 ( U4389 , INSTQUEUERD_ADDR_REG_2_ , U3257 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUE_REG_7__5_ , INSTQUEUERD_ADDR_REG_0_ );
nand NAND3_2042 ( U4390 , INSTQUEUE_REG_0__5_ , U3257 , U4368 );
nand NAND4_2043 ( U4391 , INSTQUEUE_REG_1__5_ , U2469 , INSTQUEUERD_ADDR_REG_0_ , U3252 );
nand NAND4_2044 ( U4392 , INSTQUEUE_REG_2__5_ , U2469 , INSTQUEUERD_ADDR_REG_1_ , U3253 );
nand NAND4_2045 ( U4393 , INSTQUEUE_REG_4__5_ , U4366 , INSTQUEUERD_ADDR_REG_2_ , U3257 );
nand NAND3_2046 ( U4394 , U3508 , INSTQUEUERD_ADDR_REG_2_ , U3509 );
nand NAND3_2047 ( U4395 , U3510 , INSTQUEUERD_ADDR_REG_2_ , U3511 );
nand NAND2_2048 ( U4396 , U3512 , U4368 );
nand NAND3_2049 ( U4397 , U3513 , INSTQUEUERD_ADDR_REG_1_ , U3514 );
nand NAND5_2050 ( U4398 , INSTQUEUERD_ADDR_REG_1_ , U3251 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUE_REG_11__5_ , INSTQUEUERD_ADDR_REG_3_ );
nand NAND3_2051 ( U4399 , U4366 , INSTQUEUERD_ADDR_REG_2_ , U3515 );
nand NAND5_2052 ( U4400 , INSTQUEUERD_ADDR_REG_2_ , U3252 , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUE_REG_13__5_ , INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_2053 ( U4401 , INSTQUEUERD_ADDR_REG_2_ , U3253 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUE_REG_14__5_ , INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_2054 ( U4402 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUE_REG_15__5_ , INSTQUEUERD_ADDR_REG_3_ );
not NOT1_2055 ( U4403 , U4161 );
nand NAND2_2056 ( U4404 , INSTQUEUE_REG_7__2_ , U4370 );
nand NAND2_2057 ( U4405 , INSTQUEUE_REG_0__2_ , U2472 );
nand NAND2_2058 ( U4406 , INSTQUEUE_REG_1__2_ , U2471 );
nand NAND2_2059 ( U4407 , INSTQUEUE_REG_2__2_ , U2470 );
nand NAND2_2060 ( U4408 , INSTQUEUE_REG_3__2_ , U2468 );
nand NAND2_2061 ( U4409 , INSTQUEUE_REG_4__2_ , U2467 );
nand NAND2_2062 ( U4410 , INSTQUEUE_REG_5__2_ , U2466 );
nand NAND2_2063 ( U4411 , INSTQUEUE_REG_6__2_ , U2465 );
nand NAND2_2064 ( U4412 , INSTQUEUE_REG_8__2_ , U2464 );
nand NAND2_2065 ( U4413 , INSTQUEUE_REG_9__2_ , U2463 );
nand NAND2_2066 ( U4414 , INSTQUEUE_REG_10__2_ , U2461 );
nand NAND2_2067 ( U4415 , INSTQUEUE_REG_11__2_ , U2459 );
nand NAND2_2068 ( U4416 , INSTQUEUE_REG_12__2_ , U2458 );
nand NAND2_2069 ( U4417 , INSTQUEUE_REG_13__2_ , U2457 );
nand NAND2_2070 ( U4418 , INSTQUEUE_REG_14__2_ , U2455 );
nand NAND2_2071 ( U4419 , INSTQUEUE_REG_15__2_ , U2453 );
not NOT1_2072 ( U4420 , U4159 );
nand NAND2_2073 ( U4421 , INSTQUEUE_REG_7__7_ , U4370 );
nand NAND2_2074 ( U4422 , INSTQUEUE_REG_0__7_ , U2472 );
nand NAND2_2075 ( U4423 , INSTQUEUE_REG_1__7_ , U2471 );
nand NAND2_2076 ( U4424 , INSTQUEUE_REG_2__7_ , U2470 );
nand NAND2_2077 ( U4425 , INSTQUEUE_REG_3__7_ , U2468 );
nand NAND2_2078 ( U4426 , INSTQUEUE_REG_4__7_ , U2467 );
nand NAND2_2079 ( U4427 , INSTQUEUE_REG_5__7_ , U2466 );
nand NAND2_2080 ( U4428 , INSTQUEUE_REG_6__7_ , U2465 );
nand NAND2_2081 ( U4429 , INSTQUEUE_REG_8__7_ , U2464 );
nand NAND2_2082 ( U4430 , INSTQUEUE_REG_9__7_ , U2463 );
nand NAND2_2083 ( U4431 , INSTQUEUE_REG_10__7_ , U2461 );
nand NAND2_2084 ( U4432 , INSTQUEUE_REG_11__7_ , U2459 );
nand NAND2_2085 ( U4433 , INSTQUEUE_REG_12__7_ , U2458 );
nand NAND2_2086 ( U4434 , INSTQUEUE_REG_13__7_ , U2457 );
nand NAND2_2087 ( U4435 , INSTQUEUE_REG_14__7_ , U2455 );
nand NAND2_2088 ( U4436 , INSTQUEUE_REG_15__7_ , U2453 );
not NOT1_2089 ( U4437 , U3378 );
nand NAND3_2090 ( U4438 , U3486 , U4369 , INSTQUEUE_REG_7__6_ );
nand NAND3_2091 ( U4439 , INSTQUEUE_REG_1__6_ , U2469 , U2456 );
nand NAND3_2092 ( U4440 , INSTQUEUE_REG_2__6_ , U2469 , U2454 );
nand NAND3_2093 ( U4441 , INSTQUEUE_REG_4__6_ , U4366 , U4369 );
nand NAND3_2094 ( U4442 , U2456 , U4369 , INSTQUEUE_REG_5__6_ );
nand NAND3_2095 ( U4443 , U2454 , U4369 , INSTQUEUE_REG_6__6_ );
nand NAND3_2096 ( U4444 , INSTQUEUE_REG_12__6_ , U4366 , U3495 );
nand NAND3_2097 ( U4445 , U3495 , U2456 , INSTQUEUE_REG_13__6_ );
nand NAND3_2098 ( U4446 , U3495 , U2454 , INSTQUEUE_REG_14__6_ );
nand NAND3_2099 ( U4447 , U3495 , U3486 , INSTQUEUE_REG_15__6_ );
not NOT1_2100 ( U4448 , U3264 );
nand NAND2_2101 ( U4449 , INSTQUEUE_REG_7__1_ , U4370 );
nand NAND2_2102 ( U4450 , INSTQUEUE_REG_0__1_ , U2472 );
nand NAND2_2103 ( U4451 , INSTQUEUE_REG_1__1_ , U2471 );
nand NAND2_2104 ( U4452 , INSTQUEUE_REG_2__1_ , U2470 );
nand NAND2_2105 ( U4453 , INSTQUEUE_REG_3__1_ , U2468 );
nand NAND2_2106 ( U4454 , INSTQUEUE_REG_4__1_ , U2467 );
nand NAND2_2107 ( U4455 , INSTQUEUE_REG_5__1_ , U2466 );
nand NAND2_2108 ( U4456 , INSTQUEUE_REG_6__1_ , U2465 );
nand NAND2_2109 ( U4457 , INSTQUEUE_REG_8__1_ , U2464 );
nand NAND2_2110 ( U4458 , INSTQUEUE_REG_9__1_ , U2463 );
nand NAND2_2111 ( U4459 , INSTQUEUE_REG_10__1_ , U2461 );
nand NAND2_2112 ( U4460 , INSTQUEUE_REG_11__1_ , U2459 );
nand NAND2_2113 ( U4461 , INSTQUEUE_REG_12__1_ , U2458 );
nand NAND2_2114 ( U4462 , INSTQUEUE_REG_13__1_ , U2457 );
nand NAND2_2115 ( U4463 , INSTQUEUE_REG_14__1_ , U2455 );
nand NAND2_2116 ( U4464 , INSTQUEUE_REG_15__1_ , U2453 );
not NOT1_2117 ( U4465 , U3258 );
nand NAND2_2118 ( U4466 , INSTQUEUE_REG_7__0_ , U4370 );
nand NAND2_2119 ( U4467 , INSTQUEUE_REG_0__0_ , U2472 );
nand NAND2_2120 ( U4468 , INSTQUEUE_REG_1__0_ , U2471 );
nand NAND2_2121 ( U4469 , INSTQUEUE_REG_2__0_ , U2470 );
nand NAND2_2122 ( U4470 , INSTQUEUE_REG_3__0_ , U2468 );
nand NAND2_2123 ( U4471 , INSTQUEUE_REG_4__0_ , U2467 );
nand NAND2_2124 ( U4472 , INSTQUEUE_REG_5__0_ , U2466 );
nand NAND2_2125 ( U4473 , INSTQUEUE_REG_6__0_ , U2465 );
nand NAND2_2126 ( U4474 , INSTQUEUE_REG_8__0_ , U2464 );
nand NAND2_2127 ( U4475 , INSTQUEUE_REG_9__0_ , U2463 );
nand NAND2_2128 ( U4476 , INSTQUEUE_REG_10__0_ , U2461 );
nand NAND2_2129 ( U4477 , INSTQUEUE_REG_11__0_ , U2459 );
nand NAND2_2130 ( U4478 , INSTQUEUE_REG_12__0_ , U2458 );
nand NAND2_2131 ( U4479 , INSTQUEUE_REG_13__0_ , U2457 );
nand NAND2_2132 ( U4480 , INSTQUEUE_REG_14__0_ , U2455 );
nand NAND2_2133 ( U4481 , INSTQUEUE_REG_15__0_ , U2453 );
not NOT1_2134 ( U4482 , U3271 );
nand NAND2_2135 ( U4483 , STATE_REG_2_ , U3235 );
nand NAND2_2136 ( U4484 , U3241 , U4483 );
not NOT1_2137 ( U4485 , U3259 );
nand NAND2_2138 ( U4486 , U4465 , U3375 );
not NOT1_2139 ( U4487 , U3424 );
nand NAND3_2140 ( U4488 , U3259 , U3377 , U3274 );
nand NAND2_2141 ( U4489 , U4488 , U3244 );
not NOT1_2142 ( U4490 , U3272 );
nand NAND2_2143 ( U4491 , U4448 , U4161 );
nand NAND2_2144 ( U4492 , U4184 , U3273 );
nand NAND2_2145 ( U4493 , U4492 , U3567 );
nand NAND2_2146 ( U4494 , U3568 , U4493 );
nand NAND2_2147 ( U4495 , U4203 , U3375 );
nand NAND3_2148 ( U4496 , U7670 , U7669 , U4495 );
nand NAND2_2149 ( U4497 , U2448 , U4250 );
or OR2_2150 ( U4498 , MORE_REG , FLUSH_REG );
not NOT1_2151 ( U4499 , U3280 );
nand NAND2_2152 ( U4500 , U4499 , U3249 );
nand NAND2_2153 ( U4501 , STATE2_REG_1_ , READY_N );
not NOT1_2154 ( U4502 , U3282 );
nand NAND3_2155 ( U4503 , U7676 , U7675 , STATE2_REG_1_ );
nand NAND2_2156 ( U4504 , STATE2_REG_2_ , U3282 );
nand NAND2_2157 ( U4505 , U7592 , U4234 );
nand NAND2_2158 ( U4506 , U3571 , U4502 );
nand NAND2_2159 ( U4507 , STATE2_REG_1_ , U4505 );
nand NAND2_2160 ( U4508 , U2368 , U7592 );
nand NAND2_2161 ( U4509 , U4240 , U4249 );
nand NAND2_2162 ( U4510 , U7592 , U4233 );
nand NAND2_2163 ( U4511 , U2368 , U3280 );
not NOT1_2164 ( U4512 , U3312 );
not NOT1_2165 ( U4513 , U3318 );
not NOT1_2166 ( U4514 , U3319 );
not NOT1_2167 ( U4515 , U3301 );
not NOT1_2168 ( U4516 , U3300 );
not NOT1_2169 ( U4517 , U3329 );
nand NAND2_2170 ( U4518 , R2144_U8 , U3300 );
not NOT1_2171 ( U4519 , U3345 );
not NOT1_2172 ( U4520 , U3302 );
not NOT1_2173 ( U4521 , U3292 );
not NOT1_2174 ( U4522 , U3293 );
nand NAND2_2175 ( U4523 , U2438 , U2442 );
not NOT1_2176 ( U4524 , U3308 );
not NOT1_2177 ( U4525 , U3343 );
not NOT1_2178 ( U4526 , U3327 );
nand NAND2_2179 ( U4527 , INSTQUEUEWR_ADDR_REG_3_ , U3292 );
not NOT1_2180 ( U4528 , U3347 );
not NOT1_2181 ( U4529 , U3316 );
not NOT1_2182 ( U4530 , U3310 );
not NOT1_2183 ( U4531 , U3222 );
nand NAND2_2184 ( U4532 , U2432 , U2436 );
not NOT1_2185 ( U4533 , U3309 );
nand NAND2_2186 ( U4534 , STATE2_REG_1_ , U3250 );
nand NAND3_2187 ( U4535 , U4534 , U3284 , U3286 );
nand NAND2_2188 ( U4536 , U4516 , U2476 );
nand NAND2_2189 ( U4537 , U2480 , U2358 );
nand NAND2_2190 ( U4538 , U3307 , U4537 );
nand NAND2_2191 ( U4539 , U4524 , U4538 );
nand NAND2_2192 ( U4540 , STATE2_REG_3_ , U3293 );
nand NAND2_2193 ( U4541 , U4533 , STATE2_REG_2_ );
nand NAND2_2194 ( U4542 , U4539 , U3575 );
nand NAND2_2195 ( U4543 , U2480 , U2388 );
nand NAND2_2196 ( U4544 , U3307 , U4543 );
nand NAND2_2197 ( U4545 , U4544 , U3308 );
nand NAND2_2198 ( U4546 , STATE2_REG_2_ , U3309 );
nand NAND2_2199 ( U4547 , U4546 , U4545 );
nand NAND2_2200 ( U4548 , U2415 , U4522 );
nand NAND2_2201 ( U4549 , U2413 , U2477 );
nand NAND2_2202 ( U4550 , U2412 , U4520 );
nand NAND2_2203 ( U4551 , U2397 , U4547 );
nand NAND2_2204 ( U4552 , INSTQUEUE_REG_15__7_ , U4542 );
nand NAND2_2205 ( U4553 , U2416 , U4522 );
nand NAND2_2206 ( U4554 , U2411 , U2477 );
nand NAND2_2207 ( U4555 , U2410 , U4520 );
nand NAND2_2208 ( U4556 , U2396 , U4547 );
nand NAND2_2209 ( U4557 , INSTQUEUE_REG_15__6_ , U4542 );
nand NAND2_2210 ( U4558 , U2420 , U4522 );
nand NAND2_2211 ( U4559 , U2409 , U2477 );
nand NAND2_2212 ( U4560 , U2408 , U4520 );
nand NAND2_2213 ( U4561 , U2395 , U4547 );
nand NAND2_2214 ( U4562 , INSTQUEUE_REG_15__5_ , U4542 );
nand NAND2_2215 ( U4563 , U2419 , U4522 );
nand NAND2_2216 ( U4564 , U2407 , U2477 );
nand NAND2_2217 ( U4565 , U2406 , U4520 );
nand NAND2_2218 ( U4566 , U2394 , U4547 );
nand NAND2_2219 ( U4567 , INSTQUEUE_REG_15__4_ , U4542 );
nand NAND2_2220 ( U4568 , U2418 , U4522 );
nand NAND2_2221 ( U4569 , U2405 , U2477 );
nand NAND2_2222 ( U4570 , U2404 , U4520 );
nand NAND2_2223 ( U4571 , U2393 , U4547 );
nand NAND2_2224 ( U4572 , INSTQUEUE_REG_15__3_ , U4542 );
nand NAND2_2225 ( U4573 , U2421 , U4522 );
nand NAND2_2226 ( U4574 , U2403 , U2477 );
nand NAND2_2227 ( U4575 , U2402 , U4520 );
nand NAND2_2228 ( U4576 , U2392 , U4547 );
nand NAND2_2229 ( U4577 , INSTQUEUE_REG_15__2_ , U4542 );
nand NAND2_2230 ( U4578 , U2414 , U4522 );
nand NAND2_2231 ( U4579 , U2401 , U2477 );
nand NAND2_2232 ( U4580 , U2400 , U4520 );
nand NAND2_2233 ( U4581 , U2391 , U4547 );
nand NAND2_2234 ( U4582 , INSTQUEUE_REG_15__1_ , U4542 );
nand NAND2_2235 ( U4583 , U2417 , U4522 );
nand NAND2_2236 ( U4584 , U2399 , U2477 );
nand NAND2_2237 ( U4585 , U2398 , U4520 );
nand NAND2_2238 ( U4586 , U2390 , U4547 );
nand NAND2_2239 ( U4587 , INSTQUEUE_REG_15__0_ , U4542 );
not NOT1_2240 ( U4588 , U3313 );
not NOT1_2241 ( U4589 , U3314 );
not NOT1_2242 ( U4590 , U3311 );
nand NAND2_2243 ( U4591 , U2443 , U2438 );
not NOT1_2244 ( U4592 , U3315 );
not NOT1_2245 ( U4593 , U3223 );
nand NAND2_2246 ( U4594 , U4512 , U2476 );
nand NAND2_2247 ( U4595 , U2482 , U2358 );
nand NAND2_2248 ( U4596 , U3307 , U4595 );
nand NAND2_2249 ( U4597 , U4592 , U4596 );
nand NAND2_2250 ( U4598 , STATE2_REG_3_ , U3311 );
nand NAND2_2251 ( U4599 , STATE2_REG_2_ , U3223 );
nand NAND2_2252 ( U4600 , U4597 , U3584 );
nand NAND2_2253 ( U4601 , U2482 , U2388 );
nand NAND2_2254 ( U4602 , U3307 , U4601 );
nand NAND2_2255 ( U4603 , U4602 , U3315 );
nand NAND2_2256 ( U4604 , STATE2_REG_2_ , U4593 );
nand NAND2_2257 ( U4605 , U4604 , U4603 );
nand NAND2_2258 ( U4606 , U4590 , U2415 );
nand NAND2_2259 ( U4607 , U2481 , U2413 );
nand NAND2_2260 ( U4608 , U4589 , U2412 );
nand NAND2_2261 ( U4609 , U2397 , U4605 );
nand NAND2_2262 ( U4610 , INSTQUEUE_REG_14__7_ , U4600 );
nand NAND2_2263 ( U4611 , U4590 , U2416 );
nand NAND2_2264 ( U4612 , U2481 , U2411 );
nand NAND2_2265 ( U4613 , U4589 , U2410 );
nand NAND2_2266 ( U4614 , U2396 , U4605 );
nand NAND2_2267 ( U4615 , INSTQUEUE_REG_14__6_ , U4600 );
nand NAND2_2268 ( U4616 , U4590 , U2420 );
nand NAND2_2269 ( U4617 , U2481 , U2409 );
nand NAND2_2270 ( U4618 , U4589 , U2408 );
nand NAND2_2271 ( U4619 , U2395 , U4605 );
nand NAND2_2272 ( U4620 , INSTQUEUE_REG_14__5_ , U4600 );
nand NAND2_2273 ( U4621 , U4590 , U2419 );
nand NAND2_2274 ( U4622 , U2481 , U2407 );
nand NAND2_2275 ( U4623 , U4589 , U2406 );
nand NAND2_2276 ( U4624 , U2394 , U4605 );
nand NAND2_2277 ( U4625 , INSTQUEUE_REG_14__4_ , U4600 );
nand NAND2_2278 ( U4626 , U4590 , U2418 );
nand NAND2_2279 ( U4627 , U2481 , U2405 );
nand NAND2_2280 ( U4628 , U4589 , U2404 );
nand NAND2_2281 ( U4629 , U2393 , U4605 );
nand NAND2_2282 ( U4630 , INSTQUEUE_REG_14__3_ , U4600 );
nand NAND2_2283 ( U4631 , U4590 , U2421 );
nand NAND2_2284 ( U4632 , U2481 , U2403 );
nand NAND2_2285 ( U4633 , U4589 , U2402 );
nand NAND2_2286 ( U4634 , U2392 , U4605 );
nand NAND2_2287 ( U4635 , INSTQUEUE_REG_14__2_ , U4600 );
nand NAND2_2288 ( U4636 , U4590 , U2414 );
nand NAND2_2289 ( U4637 , U2481 , U2401 );
nand NAND2_2290 ( U4638 , U4589 , U2400 );
nand NAND2_2291 ( U4639 , U2391 , U4605 );
nand NAND2_2292 ( U4640 , INSTQUEUE_REG_14__1_ , U4600 );
nand NAND2_2293 ( U4641 , U4590 , U2417 );
nand NAND2_2294 ( U4642 , U2481 , U2399 );
nand NAND2_2295 ( U4643 , U4589 , U2398 );
nand NAND2_2296 ( U4644 , U2390 , U4605 );
nand NAND2_2297 ( U4645 , INSTQUEUE_REG_14__0_ , U4600 );
not NOT1_2298 ( U4646 , U3320 );
not NOT1_2299 ( U4647 , U3321 );
not NOT1_2300 ( U4648 , U3317 );
nand NAND2_2301 ( U4649 , U2444 , U2438 );
not NOT1_2302 ( U4650 , U3322 );
nand NAND2_2303 ( U4651 , U2437 , U2432 );
not NOT1_2304 ( U4652 , U3323 );
nand NAND2_2305 ( U4653 , U4513 , U2476 );
nand NAND2_2306 ( U4654 , U2484 , U2358 );
nand NAND2_2307 ( U4655 , U3307 , U4654 );
nand NAND2_2308 ( U4656 , U4650 , U4655 );
nand NAND2_2309 ( U4657 , STATE2_REG_3_ , U3317 );
nand NAND2_2310 ( U4658 , U4652 , STATE2_REG_2_ );
nand NAND2_2311 ( U4659 , U4656 , U3593 );
nand NAND2_2312 ( U4660 , U2484 , U2388 );
nand NAND2_2313 ( U4661 , U3307 , U4660 );
nand NAND2_2314 ( U4662 , U4661 , U3322 );
nand NAND2_2315 ( U4663 , STATE2_REG_2_ , U3323 );
nand NAND2_2316 ( U4664 , U4663 , U4662 );
nand NAND2_2317 ( U4665 , U4648 , U2415 );
nand NAND2_2318 ( U4666 , U2483 , U2413 );
nand NAND2_2319 ( U4667 , U4647 , U2412 );
nand NAND2_2320 ( U4668 , U2397 , U4664 );
nand NAND2_2321 ( U4669 , INSTQUEUE_REG_13__7_ , U4659 );
nand NAND2_2322 ( U4670 , U4648 , U2416 );
nand NAND2_2323 ( U4671 , U2483 , U2411 );
nand NAND2_2324 ( U4672 , U4647 , U2410 );
nand NAND2_2325 ( U4673 , U2396 , U4664 );
nand NAND2_2326 ( U4674 , INSTQUEUE_REG_13__6_ , U4659 );
nand NAND2_2327 ( U4675 , U4648 , U2420 );
nand NAND2_2328 ( U4676 , U2483 , U2409 );
nand NAND2_2329 ( U4677 , U4647 , U2408 );
nand NAND2_2330 ( U4678 , U2395 , U4664 );
nand NAND2_2331 ( U4679 , INSTQUEUE_REG_13__5_ , U4659 );
nand NAND2_2332 ( U4680 , U4648 , U2419 );
nand NAND2_2333 ( U4681 , U2483 , U2407 );
nand NAND2_2334 ( U4682 , U4647 , U2406 );
nand NAND2_2335 ( U4683 , U2394 , U4664 );
nand NAND2_2336 ( U4684 , INSTQUEUE_REG_13__4_ , U4659 );
nand NAND2_2337 ( U4685 , U4648 , U2418 );
nand NAND2_2338 ( U4686 , U2483 , U2405 );
nand NAND2_2339 ( U4687 , U4647 , U2404 );
nand NAND2_2340 ( U4688 , U2393 , U4664 );
nand NAND2_2341 ( U4689 , INSTQUEUE_REG_13__3_ , U4659 );
nand NAND2_2342 ( U4690 , U4648 , U2421 );
nand NAND2_2343 ( U4691 , U2483 , U2403 );
nand NAND2_2344 ( U4692 , U4647 , U2402 );
nand NAND2_2345 ( U4693 , U2392 , U4664 );
nand NAND2_2346 ( U4694 , INSTQUEUE_REG_13__2_ , U4659 );
nand NAND2_2347 ( U4695 , U4648 , U2414 );
nand NAND2_2348 ( U4696 , U2483 , U2401 );
nand NAND2_2349 ( U4697 , U4647 , U2400 );
nand NAND2_2350 ( U4698 , U2391 , U4664 );
nand NAND2_2351 ( U4699 , INSTQUEUE_REG_13__1_ , U4659 );
nand NAND2_2352 ( U4700 , U4648 , U2417 );
nand NAND2_2353 ( U4701 , U2483 , U2399 );
nand NAND2_2354 ( U4702 , U4647 , U2398 );
nand NAND2_2355 ( U4703 , U2390 , U4664 );
nand NAND2_2356 ( U4704 , INSTQUEUE_REG_13__0_ , U4659 );
not NOT1_2357 ( U4705 , U3325 );
not NOT1_2358 ( U4706 , U3324 );
nand NAND2_2359 ( U4707 , U2445 , U2438 );
not NOT1_2360 ( U4708 , U3326 );
not NOT1_2361 ( U4709 , U3224 );
nand NAND2_2362 ( U4710 , U2486 , U2476 );
nand NAND2_2363 ( U4711 , U2489 , U2358 );
nand NAND2_2364 ( U4712 , U3307 , U4711 );
nand NAND2_2365 ( U4713 , U4708 , U4712 );
nand NAND2_2366 ( U4714 , STATE2_REG_3_ , U3324 );
nand NAND2_2367 ( U4715 , STATE2_REG_2_ , U3224 );
nand NAND2_2368 ( U4716 , U4713 , U3602 );
nand NAND2_2369 ( U4717 , U2489 , U2388 );
nand NAND2_2370 ( U4718 , U3307 , U4717 );
nand NAND2_2371 ( U4719 , U4718 , U3326 );
nand NAND2_2372 ( U4720 , STATE2_REG_2_ , U4709 );
nand NAND2_2373 ( U4721 , U4720 , U4719 );
nand NAND2_2374 ( U4722 , U4706 , U2415 );
nand NAND2_2375 ( U4723 , U2487 , U2413 );
nand NAND2_2376 ( U4724 , U4705 , U2412 );
nand NAND2_2377 ( U4725 , U2397 , U4721 );
nand NAND2_2378 ( U4726 , INSTQUEUE_REG_12__7_ , U4716 );
nand NAND2_2379 ( U4727 , U4706 , U2416 );
nand NAND2_2380 ( U4728 , U2487 , U2411 );
nand NAND2_2381 ( U4729 , U4705 , U2410 );
nand NAND2_2382 ( U4730 , U2396 , U4721 );
nand NAND2_2383 ( U4731 , INSTQUEUE_REG_12__6_ , U4716 );
nand NAND2_2384 ( U4732 , U4706 , U2420 );
nand NAND2_2385 ( U4733 , U2487 , U2409 );
nand NAND2_2386 ( U4734 , U4705 , U2408 );
nand NAND2_2387 ( U4735 , U2395 , U4721 );
nand NAND2_2388 ( U4736 , INSTQUEUE_REG_12__5_ , U4716 );
nand NAND2_2389 ( U4737 , U4706 , U2419 );
nand NAND2_2390 ( U4738 , U2487 , U2407 );
nand NAND2_2391 ( U4739 , U4705 , U2406 );
nand NAND2_2392 ( U4740 , U2394 , U4721 );
nand NAND2_2393 ( U4741 , INSTQUEUE_REG_12__4_ , U4716 );
nand NAND2_2394 ( U4742 , U4706 , U2418 );
nand NAND2_2395 ( U4743 , U2487 , U2405 );
nand NAND2_2396 ( U4744 , U4705 , U2404 );
nand NAND2_2397 ( U4745 , U2393 , U4721 );
nand NAND2_2398 ( U4746 , INSTQUEUE_REG_12__3_ , U4716 );
nand NAND2_2399 ( U4747 , U4706 , U2421 );
nand NAND2_2400 ( U4748 , U2487 , U2403 );
nand NAND2_2401 ( U4749 , U4705 , U2402 );
nand NAND2_2402 ( U4750 , U2392 , U4721 );
nand NAND2_2403 ( U4751 , INSTQUEUE_REG_12__2_ , U4716 );
nand NAND2_2404 ( U4752 , U4706 , U2414 );
nand NAND2_2405 ( U4753 , U2487 , U2401 );
nand NAND2_2406 ( U4754 , U4705 , U2400 );
nand NAND2_2407 ( U4755 , U2391 , U4721 );
nand NAND2_2408 ( U4756 , INSTQUEUE_REG_12__1_ , U4716 );
nand NAND2_2409 ( U4757 , U4706 , U2417 );
nand NAND2_2410 ( U4758 , U2487 , U2399 );
nand NAND2_2411 ( U4759 , U4705 , U2398 );
nand NAND2_2412 ( U4760 , U2390 , U4721 );
nand NAND2_2413 ( U4761 , INSTQUEUE_REG_12__0_ , U4716 );
not NOT1_2414 ( U4762 , U3330 );
not NOT1_2415 ( U4763 , U3328 );
nand NAND2_2416 ( U4764 , U2440 , U2442 );
not NOT1_2417 ( U4765 , U3331 );
nand NAND2_2418 ( U4766 , U2434 , U2436 );
not NOT1_2419 ( U4767 , U3332 );
nand NAND2_2420 ( U4768 , U4517 , U4516 );
nand NAND2_2421 ( U4769 , U2492 , U2358 );
nand NAND2_2422 ( U4770 , U3307 , U4769 );
nand NAND2_2423 ( U4771 , U4765 , U4770 );
nand NAND2_2424 ( U4772 , STATE2_REG_3_ , U3328 );
nand NAND2_2425 ( U4773 , U4767 , STATE2_REG_2_ );
nand NAND2_2426 ( U4774 , U4771 , U3611 );
nand NAND2_2427 ( U4775 , U2492 , U2388 );
nand NAND2_2428 ( U4776 , U3307 , U4775 );
nand NAND2_2429 ( U4777 , U4776 , U3331 );
nand NAND2_2430 ( U4778 , STATE2_REG_2_ , U3332 );
nand NAND2_2431 ( U4779 , U4778 , U4777 );
nand NAND2_2432 ( U4780 , U4763 , U2415 );
nand NAND2_2433 ( U4781 , U2491 , U2413 );
nand NAND2_2434 ( U4782 , U4762 , U2412 );
nand NAND2_2435 ( U4783 , U2397 , U4779 );
nand NAND2_2436 ( U4784 , INSTQUEUE_REG_11__7_ , U4774 );
nand NAND2_2437 ( U4785 , U4763 , U2416 );
nand NAND2_2438 ( U4786 , U2491 , U2411 );
nand NAND2_2439 ( U4787 , U4762 , U2410 );
nand NAND2_2440 ( U4788 , U2396 , U4779 );
nand NAND2_2441 ( U4789 , INSTQUEUE_REG_11__6_ , U4774 );
nand NAND2_2442 ( U4790 , U4763 , U2420 );
nand NAND2_2443 ( U4791 , U2491 , U2409 );
nand NAND2_2444 ( U4792 , U4762 , U2408 );
nand NAND2_2445 ( U4793 , U2395 , U4779 );
nand NAND2_2446 ( U4794 , INSTQUEUE_REG_11__5_ , U4774 );
nand NAND2_2447 ( U4795 , U4763 , U2419 );
nand NAND2_2448 ( U4796 , U2491 , U2407 );
nand NAND2_2449 ( U4797 , U4762 , U2406 );
nand NAND2_2450 ( U4798 , U2394 , U4779 );
nand NAND2_2451 ( U4799 , INSTQUEUE_REG_11__4_ , U4774 );
nand NAND2_2452 ( U4800 , U4763 , U2418 );
nand NAND2_2453 ( U4801 , U2491 , U2405 );
nand NAND2_2454 ( U4802 , U4762 , U2404 );
nand NAND2_2455 ( U4803 , U2393 , U4779 );
nand NAND2_2456 ( U4804 , INSTQUEUE_REG_11__3_ , U4774 );
nand NAND2_2457 ( U4805 , U4763 , U2421 );
nand NAND2_2458 ( U4806 , U2491 , U2403 );
nand NAND2_2459 ( U4807 , U4762 , U2402 );
nand NAND2_2460 ( U4808 , U2392 , U4779 );
nand NAND2_2461 ( U4809 , INSTQUEUE_REG_11__2_ , U4774 );
nand NAND2_2462 ( U4810 , U4763 , U2414 );
nand NAND2_2463 ( U4811 , U2491 , U2401 );
nand NAND2_2464 ( U4812 , U4762 , U2400 );
nand NAND2_2465 ( U4813 , U2391 , U4779 );
nand NAND2_2466 ( U4814 , INSTQUEUE_REG_11__1_ , U4774 );
nand NAND2_2467 ( U4815 , U4763 , U2417 );
nand NAND2_2468 ( U4816 , U2491 , U2399 );
nand NAND2_2469 ( U4817 , U4762 , U2398 );
nand NAND2_2470 ( U4818 , U2390 , U4779 );
nand NAND2_2471 ( U4819 , INSTQUEUE_REG_11__0_ , U4774 );
not NOT1_2472 ( U4820 , U3334 );
not NOT1_2473 ( U4821 , U3333 );
nand NAND2_2474 ( U4822 , U2440 , U2443 );
not NOT1_2475 ( U4823 , U3335 );
not NOT1_2476 ( U4824 , U3225 );
nand NAND2_2477 ( U4825 , U4517 , U4512 );
nand NAND2_2478 ( U4826 , U2494 , U2358 );
nand NAND2_2479 ( U4827 , U3307 , U4826 );
nand NAND2_2480 ( U4828 , U4823 , U4827 );
nand NAND2_2481 ( U4829 , STATE2_REG_3_ , U3333 );
nand NAND2_2482 ( U4830 , STATE2_REG_2_ , U3225 );
nand NAND2_2483 ( U4831 , U4828 , U3620 );
nand NAND2_2484 ( U4832 , U2494 , U2388 );
nand NAND2_2485 ( U4833 , U3307 , U4832 );
nand NAND2_2486 ( U4834 , U4833 , U3335 );
nand NAND2_2487 ( U4835 , STATE2_REG_2_ , U4824 );
nand NAND2_2488 ( U4836 , U4835 , U4834 );
nand NAND2_2489 ( U4837 , U4821 , U2415 );
nand NAND2_2490 ( U4838 , U2493 , U2413 );
nand NAND2_2491 ( U4839 , U4820 , U2412 );
nand NAND2_2492 ( U4840 , U2397 , U4836 );
nand NAND2_2493 ( U4841 , INSTQUEUE_REG_10__7_ , U4831 );
nand NAND2_2494 ( U4842 , U4821 , U2416 );
nand NAND2_2495 ( U4843 , U2493 , U2411 );
nand NAND2_2496 ( U4844 , U4820 , U2410 );
nand NAND2_2497 ( U4845 , U2396 , U4836 );
nand NAND2_2498 ( U4846 , INSTQUEUE_REG_10__6_ , U4831 );
nand NAND2_2499 ( U4847 , U4821 , U2420 );
nand NAND2_2500 ( U4848 , U2493 , U2409 );
nand NAND2_2501 ( U4849 , U4820 , U2408 );
nand NAND2_2502 ( U4850 , U2395 , U4836 );
nand NAND2_2503 ( U4851 , INSTQUEUE_REG_10__5_ , U4831 );
nand NAND2_2504 ( U4852 , U4821 , U2419 );
nand NAND2_2505 ( U4853 , U2493 , U2407 );
nand NAND2_2506 ( U4854 , U4820 , U2406 );
nand NAND2_2507 ( U4855 , U2394 , U4836 );
nand NAND2_2508 ( U4856 , INSTQUEUE_REG_10__4_ , U4831 );
nand NAND2_2509 ( U4857 , U4821 , U2418 );
nand NAND2_2510 ( U4858 , U2493 , U2405 );
nand NAND2_2511 ( U4859 , U4820 , U2404 );
nand NAND2_2512 ( U4860 , U2393 , U4836 );
nand NAND2_2513 ( U4861 , INSTQUEUE_REG_10__3_ , U4831 );
nand NAND2_2514 ( U4862 , U4821 , U2421 );
nand NAND2_2515 ( U4863 , U2493 , U2403 );
nand NAND2_2516 ( U4864 , U4820 , U2402 );
nand NAND2_2517 ( U4865 , U2392 , U4836 );
nand NAND2_2518 ( U4866 , INSTQUEUE_REG_10__2_ , U4831 );
nand NAND2_2519 ( U4867 , U4821 , U2414 );
nand NAND2_2520 ( U4868 , U2493 , U2401 );
nand NAND2_2521 ( U4869 , U4820 , U2400 );
nand NAND2_2522 ( U4870 , U2391 , U4836 );
nand NAND2_2523 ( U4871 , INSTQUEUE_REG_10__1_ , U4831 );
nand NAND2_2524 ( U4872 , U4821 , U2417 );
nand NAND2_2525 ( U4873 , U2493 , U2399 );
nand NAND2_2526 ( U4874 , U4820 , U2398 );
nand NAND2_2527 ( U4875 , U2390 , U4836 );
nand NAND2_2528 ( U4876 , INSTQUEUE_REG_10__0_ , U4831 );
not NOT1_2529 ( U4877 , U3337 );
not NOT1_2530 ( U4878 , U3336 );
nand NAND2_2531 ( U4879 , U2440 , U2444 );
not NOT1_2532 ( U4880 , U3338 );
nand NAND2_2533 ( U4881 , U2434 , U2437 );
not NOT1_2534 ( U4882 , U3339 );
nand NAND2_2535 ( U4883 , U4517 , U4513 );
nand NAND2_2536 ( U4884 , U2496 , U2358 );
nand NAND2_2537 ( U4885 , U3307 , U4884 );
nand NAND2_2538 ( U4886 , U4880 , U4885 );
nand NAND2_2539 ( U4887 , STATE2_REG_3_ , U3336 );
nand NAND2_2540 ( U4888 , U4882 , STATE2_REG_2_ );
nand NAND2_2541 ( U4889 , U4886 , U3629 );
nand NAND2_2542 ( U4890 , U2496 , U2388 );
nand NAND2_2543 ( U4891 , U3307 , U4890 );
nand NAND2_2544 ( U4892 , U4891 , U3338 );
nand NAND2_2545 ( U4893 , STATE2_REG_2_ , U3339 );
nand NAND2_2546 ( U4894 , U4893 , U4892 );
nand NAND2_2547 ( U4895 , U4878 , U2415 );
nand NAND2_2548 ( U4896 , U2495 , U2413 );
nand NAND2_2549 ( U4897 , U4877 , U2412 );
nand NAND2_2550 ( U4898 , U2397 , U4894 );
nand NAND2_2551 ( U4899 , INSTQUEUE_REG_9__7_ , U4889 );
nand NAND2_2552 ( U4900 , U4878 , U2416 );
nand NAND2_2553 ( U4901 , U2495 , U2411 );
nand NAND2_2554 ( U4902 , U4877 , U2410 );
nand NAND2_2555 ( U4903 , U2396 , U4894 );
nand NAND2_2556 ( U4904 , INSTQUEUE_REG_9__6_ , U4889 );
nand NAND2_2557 ( U4905 , U4878 , U2420 );
nand NAND2_2558 ( U4906 , U2495 , U2409 );
nand NAND2_2559 ( U4907 , U4877 , U2408 );
nand NAND2_2560 ( U4908 , U2395 , U4894 );
nand NAND2_2561 ( U4909 , INSTQUEUE_REG_9__5_ , U4889 );
nand NAND2_2562 ( U4910 , U4878 , U2419 );
nand NAND2_2563 ( U4911 , U2495 , U2407 );
nand NAND2_2564 ( U4912 , U4877 , U2406 );
nand NAND2_2565 ( U4913 , U2394 , U4894 );
nand NAND2_2566 ( U4914 , INSTQUEUE_REG_9__4_ , U4889 );
nand NAND2_2567 ( U4915 , U4878 , U2418 );
nand NAND2_2568 ( U4916 , U2495 , U2405 );
nand NAND2_2569 ( U4917 , U4877 , U2404 );
nand NAND2_2570 ( U4918 , U2393 , U4894 );
nand NAND2_2571 ( U4919 , INSTQUEUE_REG_9__3_ , U4889 );
nand NAND2_2572 ( U4920 , U4878 , U2421 );
nand NAND2_2573 ( U4921 , U2495 , U2403 );
nand NAND2_2574 ( U4922 , U4877 , U2402 );
nand NAND2_2575 ( U4923 , U2392 , U4894 );
nand NAND2_2576 ( U4924 , INSTQUEUE_REG_9__2_ , U4889 );
nand NAND2_2577 ( U4925 , U4878 , U2414 );
nand NAND2_2578 ( U4926 , U2495 , U2401 );
nand NAND2_2579 ( U4927 , U4877 , U2400 );
nand NAND2_2580 ( U4928 , U2391 , U4894 );
nand NAND2_2581 ( U4929 , INSTQUEUE_REG_9__1_ , U4889 );
nand NAND2_2582 ( U4930 , U4878 , U2417 );
nand NAND2_2583 ( U4931 , U2495 , U2399 );
nand NAND2_2584 ( U4932 , U4877 , U2398 );
nand NAND2_2585 ( U4933 , U2390 , U4894 );
nand NAND2_2586 ( U4934 , INSTQUEUE_REG_9__0_ , U4889 );
not NOT1_2587 ( U4935 , U3341 );
not NOT1_2588 ( U4936 , U3340 );
nand NAND2_2589 ( U4937 , U2440 , U2445 );
not NOT1_2590 ( U4938 , U3342 );
not NOT1_2591 ( U4939 , U3226 );
nand NAND2_2592 ( U4940 , U4517 , U2486 );
nand NAND2_2593 ( U4941 , U2498 , U2358 );
nand NAND2_2594 ( U4942 , U3307 , U4941 );
nand NAND2_2595 ( U4943 , U4938 , U4942 );
nand NAND2_2596 ( U4944 , STATE2_REG_3_ , U3340 );
nand NAND2_2597 ( U4945 , STATE2_REG_2_ , U3226 );
nand NAND2_2598 ( U4946 , U4943 , U3638 );
nand NAND2_2599 ( U4947 , U2498 , U2388 );
nand NAND2_2600 ( U4948 , U3307 , U4947 );
nand NAND2_2601 ( U4949 , U4948 , U3342 );
nand NAND2_2602 ( U4950 , STATE2_REG_2_ , U4939 );
nand NAND2_2603 ( U4951 , U4950 , U4949 );
nand NAND2_2604 ( U4952 , U4936 , U2415 );
nand NAND2_2605 ( U4953 , U2497 , U2413 );
nand NAND2_2606 ( U4954 , U4935 , U2412 );
nand NAND2_2607 ( U4955 , U2397 , U4951 );
nand NAND2_2608 ( U4956 , INSTQUEUE_REG_8__7_ , U4946 );
nand NAND2_2609 ( U4957 , U4936 , U2416 );
nand NAND2_2610 ( U4958 , U2497 , U2411 );
nand NAND2_2611 ( U4959 , U4935 , U2410 );
nand NAND2_2612 ( U4960 , U2396 , U4951 );
nand NAND2_2613 ( U4961 , INSTQUEUE_REG_8__6_ , U4946 );
nand NAND2_2614 ( U4962 , U4936 , U2420 );
nand NAND2_2615 ( U4963 , U2497 , U2409 );
nand NAND2_2616 ( U4964 , U4935 , U2408 );
nand NAND2_2617 ( U4965 , U2395 , U4951 );
nand NAND2_2618 ( U4966 , INSTQUEUE_REG_8__5_ , U4946 );
nand NAND2_2619 ( U4967 , U4936 , U2419 );
nand NAND2_2620 ( U4968 , U2497 , U2407 );
nand NAND2_2621 ( U4969 , U4935 , U2406 );
nand NAND2_2622 ( U4970 , U2394 , U4951 );
nand NAND2_2623 ( U4971 , INSTQUEUE_REG_8__4_ , U4946 );
nand NAND2_2624 ( U4972 , U4936 , U2418 );
nand NAND2_2625 ( U4973 , U2497 , U2405 );
nand NAND2_2626 ( U4974 , U4935 , U2404 );
nand NAND2_2627 ( U4975 , U2393 , U4951 );
nand NAND2_2628 ( U4976 , INSTQUEUE_REG_8__3_ , U4946 );
nand NAND2_2629 ( U4977 , U4936 , U2421 );
nand NAND2_2630 ( U4978 , U2497 , U2403 );
nand NAND2_2631 ( U4979 , U4935 , U2402 );
nand NAND2_2632 ( U4980 , U2392 , U4951 );
nand NAND2_2633 ( U4981 , INSTQUEUE_REG_8__2_ , U4946 );
nand NAND2_2634 ( U4982 , U4936 , U2414 );
nand NAND2_2635 ( U4983 , U2497 , U2401 );
nand NAND2_2636 ( U4984 , U4935 , U2400 );
nand NAND2_2637 ( U4985 , U2391 , U4951 );
nand NAND2_2638 ( U4986 , INSTQUEUE_REG_8__1_ , U4946 );
nand NAND2_2639 ( U4987 , U4936 , U2417 );
nand NAND2_2640 ( U4988 , U2497 , U2399 );
nand NAND2_2641 ( U4989 , U4935 , U2398 );
nand NAND2_2642 ( U4990 , U2390 , U4951 );
nand NAND2_2643 ( U4991 , INSTQUEUE_REG_8__0_ , U4946 );
not NOT1_2644 ( U4992 , U3346 );
nand NAND2_2645 ( U4993 , U2439 , U2442 );
not NOT1_2646 ( U4994 , U3348 );
nand NAND2_2647 ( U4995 , U2433 , U2436 );
not NOT1_2648 ( U4996 , U3349 );
nand NAND2_2649 ( U4997 , U2500 , U2358 );
nand NAND2_2650 ( U4998 , U3307 , U4997 );
nand NAND2_2651 ( U4999 , U4994 , U4998 );
nand NAND2_2652 ( U5000 , STATE2_REG_3_ , U3343 );
nand NAND2_2653 ( U5001 , U4996 , STATE2_REG_2_ );
nand NAND2_2654 ( U5002 , U4999 , U3647 );
nand NAND2_2655 ( U5003 , U2500 , U2388 );
nand NAND2_2656 ( U5004 , U3307 , U5003 );
nand NAND2_2657 ( U5005 , U5004 , U3348 );
nand NAND2_2658 ( U5006 , STATE2_REG_2_ , U3349 );
nand NAND2_2659 ( U5007 , U5006 , U5005 );
nand NAND2_2660 ( U5008 , U4525 , U2415 );
nand NAND2_2661 ( U5009 , U4226 , U2413 );
nand NAND2_2662 ( U5010 , U4992 , U2412 );
nand NAND2_2663 ( U5011 , U2397 , U5007 );
nand NAND2_2664 ( U5012 , INSTQUEUE_REG_7__7_ , U5002 );
nand NAND2_2665 ( U5013 , U4525 , U2416 );
nand NAND2_2666 ( U5014 , U4226 , U2411 );
nand NAND2_2667 ( U5015 , U4992 , U2410 );
nand NAND2_2668 ( U5016 , U2396 , U5007 );
nand NAND2_2669 ( U5017 , INSTQUEUE_REG_7__6_ , U5002 );
nand NAND2_2670 ( U5018 , U4525 , U2420 );
nand NAND2_2671 ( U5019 , U4226 , U2409 );
nand NAND2_2672 ( U5020 , U4992 , U2408 );
nand NAND2_2673 ( U5021 , U2395 , U5007 );
nand NAND2_2674 ( U5022 , INSTQUEUE_REG_7__5_ , U5002 );
nand NAND2_2675 ( U5023 , U4525 , U2419 );
nand NAND2_2676 ( U5024 , U4226 , U2407 );
nand NAND2_2677 ( U5025 , U4992 , U2406 );
nand NAND2_2678 ( U5026 , U2394 , U5007 );
nand NAND2_2679 ( U5027 , INSTQUEUE_REG_7__4_ , U5002 );
nand NAND2_2680 ( U5028 , U4525 , U2418 );
nand NAND2_2681 ( U5029 , U4226 , U2405 );
nand NAND2_2682 ( U5030 , U4992 , U2404 );
nand NAND2_2683 ( U5031 , U2393 , U5007 );
nand NAND2_2684 ( U5032 , INSTQUEUE_REG_7__3_ , U5002 );
nand NAND2_2685 ( U5033 , U4525 , U2421 );
nand NAND2_2686 ( U5034 , U4226 , U2403 );
nand NAND2_2687 ( U5035 , U4992 , U2402 );
nand NAND2_2688 ( U5036 , U2392 , U5007 );
nand NAND2_2689 ( U5037 , INSTQUEUE_REG_7__2_ , U5002 );
nand NAND2_2690 ( U5038 , U4525 , U2414 );
nand NAND2_2691 ( U5039 , U4226 , U2401 );
nand NAND2_2692 ( U5040 , U4992 , U2400 );
nand NAND2_2693 ( U5041 , U2391 , U5007 );
nand NAND2_2694 ( U5042 , INSTQUEUE_REG_7__1_ , U5002 );
nand NAND2_2695 ( U5043 , U4525 , U2417 );
nand NAND2_2696 ( U5044 , U4226 , U2399 );
nand NAND2_2697 ( U5045 , U4992 , U2398 );
nand NAND2_2698 ( U5046 , U2390 , U5007 );
nand NAND2_2699 ( U5047 , INSTQUEUE_REG_7__0_ , U5002 );
not NOT1_2700 ( U5048 , U3351 );
not NOT1_2701 ( U5049 , U3350 );
nand NAND2_2702 ( U5050 , U2439 , U2443 );
not NOT1_2703 ( U5051 , U3352 );
not NOT1_2704 ( U5052 , U3227 );
nand NAND2_2705 ( U5053 , U4512 , U2474 );
nand NAND2_2706 ( U5054 , U2502 , U2358 );
nand NAND2_2707 ( U5055 , U3307 , U5054 );
nand NAND2_2708 ( U5056 , U5051 , U5055 );
nand NAND2_2709 ( U5057 , STATE2_REG_3_ , U3350 );
nand NAND2_2710 ( U5058 , STATE2_REG_2_ , U3227 );
nand NAND2_2711 ( U5059 , U5056 , U3656 );
nand NAND2_2712 ( U5060 , U2502 , U2388 );
nand NAND2_2713 ( U5061 , U3307 , U5060 );
nand NAND2_2714 ( U5062 , U5061 , U3352 );
nand NAND2_2715 ( U5063 , STATE2_REG_2_ , U5052 );
nand NAND2_2716 ( U5064 , U5063 , U5062 );
nand NAND2_2717 ( U5065 , U5049 , U2415 );
nand NAND2_2718 ( U5066 , U2501 , U2413 );
nand NAND2_2719 ( U5067 , U5048 , U2412 );
nand NAND2_2720 ( U5068 , U2397 , U5064 );
nand NAND2_2721 ( U5069 , INSTQUEUE_REG_6__7_ , U5059 );
nand NAND2_2722 ( U5070 , U5049 , U2416 );
nand NAND2_2723 ( U5071 , U2501 , U2411 );
nand NAND2_2724 ( U5072 , U5048 , U2410 );
nand NAND2_2725 ( U5073 , U2396 , U5064 );
nand NAND2_2726 ( U5074 , INSTQUEUE_REG_6__6_ , U5059 );
nand NAND2_2727 ( U5075 , U5049 , U2420 );
nand NAND2_2728 ( U5076 , U2501 , U2409 );
nand NAND2_2729 ( U5077 , U5048 , U2408 );
nand NAND2_2730 ( U5078 , U2395 , U5064 );
nand NAND2_2731 ( U5079 , INSTQUEUE_REG_6__5_ , U5059 );
nand NAND2_2732 ( U5080 , U5049 , U2419 );
nand NAND2_2733 ( U5081 , U2501 , U2407 );
nand NAND2_2734 ( U5082 , U5048 , U2406 );
nand NAND2_2735 ( U5083 , U2394 , U5064 );
nand NAND2_2736 ( U5084 , INSTQUEUE_REG_6__4_ , U5059 );
nand NAND2_2737 ( U5085 , U5049 , U2418 );
nand NAND2_2738 ( U5086 , U2501 , U2405 );
nand NAND2_2739 ( U5087 , U5048 , U2404 );
nand NAND2_2740 ( U5088 , U2393 , U5064 );
nand NAND2_2741 ( U5089 , INSTQUEUE_REG_6__3_ , U5059 );
nand NAND2_2742 ( U5090 , U5049 , U2421 );
nand NAND2_2743 ( U5091 , U2501 , U2403 );
nand NAND2_2744 ( U5092 , U5048 , U2402 );
nand NAND2_2745 ( U5093 , U2392 , U5064 );
nand NAND2_2746 ( U5094 , INSTQUEUE_REG_6__2_ , U5059 );
nand NAND2_2747 ( U5095 , U5049 , U2414 );
nand NAND2_2748 ( U5096 , U2501 , U2401 );
nand NAND2_2749 ( U5097 , U5048 , U2400 );
nand NAND2_2750 ( U5098 , U2391 , U5064 );
nand NAND2_2751 ( U5099 , INSTQUEUE_REG_6__1_ , U5059 );
nand NAND2_2752 ( U5100 , U5049 , U2417 );
nand NAND2_2753 ( U5101 , U2501 , U2399 );
nand NAND2_2754 ( U5102 , U5048 , U2398 );
nand NAND2_2755 ( U5103 , U2390 , U5064 );
nand NAND2_2756 ( U5104 , INSTQUEUE_REG_6__0_ , U5059 );
not NOT1_2757 ( U5105 , U3354 );
not NOT1_2758 ( U5106 , U3353 );
nand NAND2_2759 ( U5107 , U2439 , U2444 );
not NOT1_2760 ( U5108 , U3355 );
nand NAND2_2761 ( U5109 , U2433 , U2437 );
not NOT1_2762 ( U5110 , U3356 );
nand NAND2_2763 ( U5111 , U4513 , U2474 );
nand NAND2_2764 ( U5112 , U2504 , U2358 );
nand NAND2_2765 ( U5113 , U3307 , U5112 );
nand NAND2_2766 ( U5114 , U5108 , U5113 );
nand NAND2_2767 ( U5115 , STATE2_REG_3_ , U3353 );
nand NAND2_2768 ( U5116 , U5110 , STATE2_REG_2_ );
nand NAND2_2769 ( U5117 , U5114 , U3665 );
nand NAND2_2770 ( U5118 , U2504 , U2388 );
nand NAND2_2771 ( U5119 , U3307 , U5118 );
nand NAND2_2772 ( U5120 , U5119 , U3355 );
nand NAND2_2773 ( U5121 , STATE2_REG_2_ , U3356 );
nand NAND2_2774 ( U5122 , U5121 , U5120 );
nand NAND2_2775 ( U5123 , U5106 , U2415 );
nand NAND2_2776 ( U5124 , U2503 , U2413 );
nand NAND2_2777 ( U5125 , U5105 , U2412 );
nand NAND2_2778 ( U5126 , U2397 , U5122 );
nand NAND2_2779 ( U5127 , INSTQUEUE_REG_5__7_ , U5117 );
nand NAND2_2780 ( U5128 , U5106 , U2416 );
nand NAND2_2781 ( U5129 , U2503 , U2411 );
nand NAND2_2782 ( U5130 , U5105 , U2410 );
nand NAND2_2783 ( U5131 , U2396 , U5122 );
nand NAND2_2784 ( U5132 , INSTQUEUE_REG_5__6_ , U5117 );
nand NAND2_2785 ( U5133 , U5106 , U2420 );
nand NAND2_2786 ( U5134 , U2503 , U2409 );
nand NAND2_2787 ( U5135 , U5105 , U2408 );
nand NAND2_2788 ( U5136 , U2395 , U5122 );
nand NAND2_2789 ( U5137 , INSTQUEUE_REG_5__5_ , U5117 );
nand NAND2_2790 ( U5138 , U5106 , U2419 );
nand NAND2_2791 ( U5139 , U2503 , U2407 );
nand NAND2_2792 ( U5140 , U5105 , U2406 );
nand NAND2_2793 ( U5141 , U2394 , U5122 );
nand NAND2_2794 ( U5142 , INSTQUEUE_REG_5__4_ , U5117 );
nand NAND2_2795 ( U5143 , U5106 , U2418 );
nand NAND2_2796 ( U5144 , U2503 , U2405 );
nand NAND2_2797 ( U5145 , U5105 , U2404 );
nand NAND2_2798 ( U5146 , U2393 , U5122 );
nand NAND2_2799 ( U5147 , INSTQUEUE_REG_5__3_ , U5117 );
nand NAND2_2800 ( U5148 , U5106 , U2421 );
nand NAND2_2801 ( U5149 , U2503 , U2403 );
nand NAND2_2802 ( U5150 , U5105 , U2402 );
nand NAND2_2803 ( U5151 , U2392 , U5122 );
nand NAND2_2804 ( U5152 , INSTQUEUE_REG_5__2_ , U5117 );
nand NAND2_2805 ( U5153 , U5106 , U2414 );
nand NAND2_2806 ( U5154 , U2503 , U2401 );
nand NAND2_2807 ( U5155 , U5105 , U2400 );
nand NAND2_2808 ( U5156 , U2391 , U5122 );
nand NAND2_2809 ( U5157 , INSTQUEUE_REG_5__1_ , U5117 );
nand NAND2_2810 ( U5158 , U5106 , U2417 );
nand NAND2_2811 ( U5159 , U2503 , U2399 );
nand NAND2_2812 ( U5160 , U5105 , U2398 );
nand NAND2_2813 ( U5161 , U2390 , U5122 );
nand NAND2_2814 ( U5162 , INSTQUEUE_REG_5__0_ , U5117 );
not NOT1_2815 ( U5163 , U3358 );
not NOT1_2816 ( U5164 , U3357 );
nand NAND2_2817 ( U5165 , U2439 , U2445 );
not NOT1_2818 ( U5166 , U3359 );
not NOT1_2819 ( U5167 , U3228 );
nand NAND2_2820 ( U5168 , U2486 , U2474 );
nand NAND2_2821 ( U5169 , U2506 , U2358 );
nand NAND2_2822 ( U5170 , U3307 , U5169 );
nand NAND2_2823 ( U5171 , U5166 , U5170 );
nand NAND2_2824 ( U5172 , STATE2_REG_3_ , U3357 );
nand NAND2_2825 ( U5173 , STATE2_REG_2_ , U3228 );
nand NAND2_2826 ( U5174 , U5171 , U3674 );
nand NAND2_2827 ( U5175 , U2506 , U2388 );
nand NAND2_2828 ( U5176 , U3307 , U5175 );
nand NAND2_2829 ( U5177 , U5176 , U3359 );
nand NAND2_2830 ( U5178 , STATE2_REG_2_ , U5167 );
nand NAND2_2831 ( U5179 , U5178 , U5177 );
nand NAND2_2832 ( U5180 , U5164 , U2415 );
nand NAND2_2833 ( U5181 , U2505 , U2413 );
nand NAND2_2834 ( U5182 , U5163 , U2412 );
nand NAND2_2835 ( U5183 , U2397 , U5179 );
nand NAND2_2836 ( U5184 , INSTQUEUE_REG_4__7_ , U5174 );
nand NAND2_2837 ( U5185 , U5164 , U2416 );
nand NAND2_2838 ( U5186 , U2505 , U2411 );
nand NAND2_2839 ( U5187 , U5163 , U2410 );
nand NAND2_2840 ( U5188 , U2396 , U5179 );
nand NAND2_2841 ( U5189 , INSTQUEUE_REG_4__6_ , U5174 );
nand NAND2_2842 ( U5190 , U5164 , U2420 );
nand NAND2_2843 ( U5191 , U2505 , U2409 );
nand NAND2_2844 ( U5192 , U5163 , U2408 );
nand NAND2_2845 ( U5193 , U2395 , U5179 );
nand NAND2_2846 ( U5194 , INSTQUEUE_REG_4__5_ , U5174 );
nand NAND2_2847 ( U5195 , U5164 , U2419 );
nand NAND2_2848 ( U5196 , U2505 , U2407 );
nand NAND2_2849 ( U5197 , U5163 , U2406 );
nand NAND2_2850 ( U5198 , U2394 , U5179 );
nand NAND2_2851 ( U5199 , INSTQUEUE_REG_4__4_ , U5174 );
nand NAND2_2852 ( U5200 , U5164 , U2418 );
nand NAND2_2853 ( U5201 , U2505 , U2405 );
nand NAND2_2854 ( U5202 , U5163 , U2404 );
nand NAND2_2855 ( U5203 , U2393 , U5179 );
nand NAND2_2856 ( U5204 , INSTQUEUE_REG_4__3_ , U5174 );
nand NAND2_2857 ( U5205 , U5164 , U2421 );
nand NAND2_2858 ( U5206 , U2505 , U2403 );
nand NAND2_2859 ( U5207 , U5163 , U2402 );
nand NAND2_2860 ( U5208 , U2392 , U5179 );
nand NAND2_2861 ( U5209 , INSTQUEUE_REG_4__2_ , U5174 );
nand NAND2_2862 ( U5210 , U5164 , U2414 );
nand NAND2_2863 ( U5211 , U2505 , U2401 );
nand NAND2_2864 ( U5212 , U5163 , U2400 );
nand NAND2_2865 ( U5213 , U2391 , U5179 );
nand NAND2_2866 ( U5214 , INSTQUEUE_REG_4__1_ , U5174 );
nand NAND2_2867 ( U5215 , U5164 , U2417 );
nand NAND2_2868 ( U5216 , U2505 , U2399 );
nand NAND2_2869 ( U5217 , U5163 , U2398 );
nand NAND2_2870 ( U5218 , U2390 , U5179 );
nand NAND2_2871 ( U5219 , INSTQUEUE_REG_4__0_ , U5174 );
not NOT1_2872 ( U5220 , U3361 );
not NOT1_2873 ( U5221 , U3360 );
nand NAND2_2874 ( U5222 , U2441 , U2442 );
not NOT1_2875 ( U5223 , U3362 );
nand NAND2_2876 ( U5224 , U2435 , U2436 );
not NOT1_2877 ( U5225 , U3363 );
nand NAND2_2878 ( U5226 , U2508 , U4516 );
nand NAND2_2879 ( U5227 , U2511 , U2358 );
nand NAND2_2880 ( U5228 , U3307 , U5227 );
nand NAND2_2881 ( U5229 , U5223 , U5228 );
nand NAND2_2882 ( U5230 , STATE2_REG_3_ , U3360 );
nand NAND2_2883 ( U5231 , U5225 , STATE2_REG_2_ );
nand NAND2_2884 ( U5232 , U5229 , U3683 );
nand NAND2_2885 ( U5233 , U2511 , U2388 );
nand NAND2_2886 ( U5234 , U3307 , U5233 );
nand NAND2_2887 ( U5235 , U5234 , U3362 );
nand NAND2_2888 ( U5236 , STATE2_REG_2_ , U3363 );
nand NAND2_2889 ( U5237 , U5236 , U5235 );
nand NAND2_2890 ( U5238 , U5221 , U2415 );
nand NAND2_2891 ( U5239 , U2509 , U2413 );
nand NAND2_2892 ( U5240 , U5220 , U2412 );
nand NAND2_2893 ( U5241 , U2397 , U5237 );
nand NAND2_2894 ( U5242 , INSTQUEUE_REG_3__7_ , U5232 );
nand NAND2_2895 ( U5243 , U5221 , U2416 );
nand NAND2_2896 ( U5244 , U2509 , U2411 );
nand NAND2_2897 ( U5245 , U5220 , U2410 );
nand NAND2_2898 ( U5246 , U2396 , U5237 );
nand NAND2_2899 ( U5247 , INSTQUEUE_REG_3__6_ , U5232 );
nand NAND2_2900 ( U5248 , U5221 , U2420 );
nand NAND2_2901 ( U5249 , U2509 , U2409 );
nand NAND2_2902 ( U5250 , U5220 , U2408 );
nand NAND2_2903 ( U5251 , U2395 , U5237 );
nand NAND2_2904 ( U5252 , INSTQUEUE_REG_3__5_ , U5232 );
nand NAND2_2905 ( U5253 , U5221 , U2419 );
nand NAND2_2906 ( U5254 , U2509 , U2407 );
nand NAND2_2907 ( U5255 , U5220 , U2406 );
nand NAND2_2908 ( U5256 , U2394 , U5237 );
nand NAND2_2909 ( U5257 , INSTQUEUE_REG_3__4_ , U5232 );
nand NAND2_2910 ( U5258 , U5221 , U2418 );
nand NAND2_2911 ( U5259 , U2509 , U2405 );
nand NAND2_2912 ( U5260 , U5220 , U2404 );
nand NAND2_2913 ( U5261 , U2393 , U5237 );
nand NAND2_2914 ( U5262 , INSTQUEUE_REG_3__3_ , U5232 );
nand NAND2_2915 ( U5263 , U5221 , U2421 );
nand NAND2_2916 ( U5264 , U2509 , U2403 );
nand NAND2_2917 ( U5265 , U5220 , U2402 );
nand NAND2_2918 ( U5266 , U2392 , U5237 );
nand NAND2_2919 ( U5267 , INSTQUEUE_REG_3__2_ , U5232 );
nand NAND2_2920 ( U5268 , U5221 , U2414 );
nand NAND2_2921 ( U5269 , U2509 , U2401 );
nand NAND2_2922 ( U5270 , U5220 , U2400 );
nand NAND2_2923 ( U5271 , U2391 , U5237 );
nand NAND2_2924 ( U5272 , INSTQUEUE_REG_3__1_ , U5232 );
nand NAND2_2925 ( U5273 , U5221 , U2417 );
nand NAND2_2926 ( U5274 , U2509 , U2399 );
nand NAND2_2927 ( U5275 , U5220 , U2398 );
nand NAND2_2928 ( U5276 , U2390 , U5237 );
nand NAND2_2929 ( U5277 , INSTQUEUE_REG_3__0_ , U5232 );
not NOT1_2930 ( U5278 , U3365 );
not NOT1_2931 ( U5279 , U3364 );
nand NAND2_2932 ( U5280 , U2441 , U2443 );
not NOT1_2933 ( U5281 , U3366 );
not NOT1_2934 ( U5282 , U3229 );
nand NAND2_2935 ( U5283 , U2508 , U4512 );
nand NAND2_2936 ( U5284 , U2513 , U2358 );
nand NAND2_2937 ( U5285 , U3307 , U5284 );
nand NAND2_2938 ( U5286 , U5281 , U5285 );
nand NAND2_2939 ( U5287 , STATE2_REG_3_ , U3364 );
nand NAND2_2940 ( U5288 , STATE2_REG_2_ , U3229 );
nand NAND2_2941 ( U5289 , U5286 , U3692 );
nand NAND2_2942 ( U5290 , U2513 , U2388 );
nand NAND2_2943 ( U5291 , U3307 , U5290 );
nand NAND2_2944 ( U5292 , U5291 , U3366 );
nand NAND2_2945 ( U5293 , STATE2_REG_2_ , U5282 );
nand NAND2_2946 ( U5294 , U5293 , U5292 );
nand NAND2_2947 ( U5295 , U5279 , U2415 );
nand NAND2_2948 ( U5296 , U2512 , U2413 );
nand NAND2_2949 ( U5297 , U5278 , U2412 );
nand NAND2_2950 ( U5298 , U2397 , U5294 );
nand NAND2_2951 ( U5299 , INSTQUEUE_REG_2__7_ , U5289 );
nand NAND2_2952 ( U5300 , U5279 , U2416 );
nand NAND2_2953 ( U5301 , U2512 , U2411 );
nand NAND2_2954 ( U5302 , U5278 , U2410 );
nand NAND2_2955 ( U5303 , U2396 , U5294 );
nand NAND2_2956 ( U5304 , INSTQUEUE_REG_2__6_ , U5289 );
nand NAND2_2957 ( U5305 , U5279 , U2420 );
nand NAND2_2958 ( U5306 , U2512 , U2409 );
nand NAND2_2959 ( U5307 , U5278 , U2408 );
nand NAND2_2960 ( U5308 , U2395 , U5294 );
nand NAND2_2961 ( U5309 , INSTQUEUE_REG_2__5_ , U5289 );
nand NAND2_2962 ( U5310 , U5279 , U2419 );
nand NAND2_2963 ( U5311 , U2512 , U2407 );
nand NAND2_2964 ( U5312 , U5278 , U2406 );
nand NAND2_2965 ( U5313 , U2394 , U5294 );
nand NAND2_2966 ( U5314 , INSTQUEUE_REG_2__4_ , U5289 );
nand NAND2_2967 ( U5315 , U5279 , U2418 );
nand NAND2_2968 ( U5316 , U2512 , U2405 );
nand NAND2_2969 ( U5317 , U5278 , U2404 );
nand NAND2_2970 ( U5318 , U2393 , U5294 );
nand NAND2_2971 ( U5319 , INSTQUEUE_REG_2__3_ , U5289 );
nand NAND2_2972 ( U5320 , U5279 , U2421 );
nand NAND2_2973 ( U5321 , U2512 , U2403 );
nand NAND2_2974 ( U5322 , U5278 , U2402 );
nand NAND2_2975 ( U5323 , U2392 , U5294 );
nand NAND2_2976 ( U5324 , INSTQUEUE_REG_2__2_ , U5289 );
nand NAND2_2977 ( U5325 , U5279 , U2414 );
nand NAND2_2978 ( U5326 , U2512 , U2401 );
nand NAND2_2979 ( U5327 , U5278 , U2400 );
nand NAND2_2980 ( U5328 , U2391 , U5294 );
nand NAND2_2981 ( U5329 , INSTQUEUE_REG_2__1_ , U5289 );
nand NAND2_2982 ( U5330 , U5279 , U2417 );
nand NAND2_2983 ( U5331 , U2512 , U2399 );
nand NAND2_2984 ( U5332 , U5278 , U2398 );
nand NAND2_2985 ( U5333 , U2390 , U5294 );
nand NAND2_2986 ( U5334 , INSTQUEUE_REG_2__0_ , U5289 );
not NOT1_2987 ( U5335 , U3368 );
not NOT1_2988 ( U5336 , U3367 );
nand NAND2_2989 ( U5337 , U2441 , U2444 );
not NOT1_2990 ( U5338 , U3369 );
nand NAND2_2991 ( U5339 , U2435 , U2437 );
not NOT1_2992 ( U5340 , U3370 );
nand NAND2_2993 ( U5341 , U2508 , U4513 );
nand NAND2_2994 ( U5342 , U2515 , U2358 );
nand NAND2_2995 ( U5343 , U3307 , U5342 );
nand NAND2_2996 ( U5344 , U5338 , U5343 );
nand NAND2_2997 ( U5345 , STATE2_REG_3_ , U3367 );
nand NAND2_2998 ( U5346 , U5340 , STATE2_REG_2_ );
nand NAND2_2999 ( U5347 , U5344 , U3701 );
nand NAND2_3000 ( U5348 , U2515 , U2388 );
nand NAND2_3001 ( U5349 , U3307 , U5348 );
nand NAND2_3002 ( U5350 , U5349 , U3369 );
nand NAND2_3003 ( U5351 , STATE2_REG_2_ , U3370 );
nand NAND2_3004 ( U5352 , U5351 , U5350 );
nand NAND2_3005 ( U5353 , U5336 , U2415 );
nand NAND2_3006 ( U5354 , U2514 , U2413 );
nand NAND2_3007 ( U5355 , U5335 , U2412 );
nand NAND2_3008 ( U5356 , U2397 , U5352 );
nand NAND2_3009 ( U5357 , INSTQUEUE_REG_1__7_ , U5347 );
nand NAND2_3010 ( U5358 , U5336 , U2416 );
nand NAND2_3011 ( U5359 , U2514 , U2411 );
nand NAND2_3012 ( U5360 , U5335 , U2410 );
nand NAND2_3013 ( U5361 , U2396 , U5352 );
nand NAND2_3014 ( U5362 , INSTQUEUE_REG_1__6_ , U5347 );
nand NAND2_3015 ( U5363 , U5336 , U2420 );
nand NAND2_3016 ( U5364 , U2514 , U2409 );
nand NAND2_3017 ( U5365 , U5335 , U2408 );
nand NAND2_3018 ( U5366 , U2395 , U5352 );
nand NAND2_3019 ( U5367 , INSTQUEUE_REG_1__5_ , U5347 );
nand NAND2_3020 ( U5368 , U5336 , U2419 );
nand NAND2_3021 ( U5369 , U2514 , U2407 );
nand NAND2_3022 ( U5370 , U5335 , U2406 );
nand NAND2_3023 ( U5371 , U2394 , U5352 );
nand NAND2_3024 ( U5372 , INSTQUEUE_REG_1__4_ , U5347 );
nand NAND2_3025 ( U5373 , U5336 , U2418 );
nand NAND2_3026 ( U5374 , U2514 , U2405 );
nand NAND2_3027 ( U5375 , U5335 , U2404 );
nand NAND2_3028 ( U5376 , U2393 , U5352 );
nand NAND2_3029 ( U5377 , INSTQUEUE_REG_1__3_ , U5347 );
nand NAND2_3030 ( U5378 , U5336 , U2421 );
nand NAND2_3031 ( U5379 , U2514 , U2403 );
nand NAND2_3032 ( U5380 , U5335 , U2402 );
nand NAND2_3033 ( U5381 , U2392 , U5352 );
nand NAND2_3034 ( U5382 , INSTQUEUE_REG_1__2_ , U5347 );
nand NAND2_3035 ( U5383 , U5336 , U2414 );
nand NAND2_3036 ( U5384 , U2514 , U2401 );
nand NAND2_3037 ( U5385 , U5335 , U2400 );
nand NAND2_3038 ( U5386 , U2391 , U5352 );
nand NAND2_3039 ( U5387 , INSTQUEUE_REG_1__1_ , U5347 );
nand NAND2_3040 ( U5388 , U5336 , U2417 );
nand NAND2_3041 ( U5389 , U2514 , U2399 );
nand NAND2_3042 ( U5390 , U5335 , U2398 );
nand NAND2_3043 ( U5391 , U2390 , U5352 );
nand NAND2_3044 ( U5392 , INSTQUEUE_REG_1__0_ , U5347 );
not NOT1_3045 ( U5393 , U3372 );
not NOT1_3046 ( U5394 , U3371 );
nand NAND2_3047 ( U5395 , U2441 , U2445 );
not NOT1_3048 ( U5396 , U3373 );
not NOT1_3049 ( U5397 , U3230 );
nand NAND2_3050 ( U5398 , U2508 , U2486 );
nand NAND2_3051 ( U5399 , U2517 , U2358 );
nand NAND2_3052 ( U5400 , U3307 , U5399 );
nand NAND2_3053 ( U5401 , U5396 , U5400 );
nand NAND2_3054 ( U5402 , STATE2_REG_3_ , U3371 );
nand NAND2_3055 ( U5403 , STATE2_REG_2_ , U3230 );
nand NAND2_3056 ( U5404 , U5401 , U3710 );
nand NAND2_3057 ( U5405 , U2517 , U2388 );
nand NAND2_3058 ( U5406 , U3307 , U5405 );
nand NAND2_3059 ( U5407 , U5406 , U3373 );
nand NAND2_3060 ( U5408 , STATE2_REG_2_ , U5397 );
nand NAND2_3061 ( U5409 , U5408 , U5407 );
nand NAND2_3062 ( U5410 , U5394 , U2415 );
nand NAND2_3063 ( U5411 , U2516 , U2413 );
nand NAND2_3064 ( U5412 , U5393 , U2412 );
nand NAND2_3065 ( U5413 , U2397 , U5409 );
nand NAND2_3066 ( U5414 , INSTQUEUE_REG_0__7_ , U5404 );
nand NAND2_3067 ( U5415 , U5394 , U2416 );
nand NAND2_3068 ( U5416 , U2516 , U2411 );
nand NAND2_3069 ( U5417 , U5393 , U2410 );
nand NAND2_3070 ( U5418 , U2396 , U5409 );
nand NAND2_3071 ( U5419 , INSTQUEUE_REG_0__6_ , U5404 );
nand NAND2_3072 ( U5420 , U5394 , U2420 );
nand NAND2_3073 ( U5421 , U2516 , U2409 );
nand NAND2_3074 ( U5422 , U5393 , U2408 );
nand NAND2_3075 ( U5423 , U2395 , U5409 );
nand NAND2_3076 ( U5424 , INSTQUEUE_REG_0__5_ , U5404 );
nand NAND2_3077 ( U5425 , U5394 , U2419 );
nand NAND2_3078 ( U5426 , U2516 , U2407 );
nand NAND2_3079 ( U5427 , U5393 , U2406 );
nand NAND2_3080 ( U5428 , U2394 , U5409 );
nand NAND2_3081 ( U5429 , U5394 , U2418 );
nand NAND2_3082 ( U5430 , U2516 , U2405 );
nand NAND2_3083 ( U5431 , U5393 , U2404 );
nand NAND2_3084 ( U5432 , U2393 , U5409 );
nand NAND2_3085 ( U5433 , INSTQUEUE_REG_0__3_ , U5404 );
nand NAND2_3086 ( U5434 , U5394 , U2421 );
nand NAND2_3087 ( U5435 , U2516 , U2403 );
nand NAND2_3088 ( U5436 , U5393 , U2402 );
nand NAND2_3089 ( U5437 , U2392 , U5409 );
nand NAND2_3090 ( U5438 , INSTQUEUE_REG_0__2_ , U5404 );
nand NAND2_3091 ( U5439 , U5394 , U2414 );
nand NAND2_3092 ( U5440 , U2516 , U2401 );
nand NAND2_3093 ( U5441 , U5393 , U2400 );
nand NAND2_3094 ( U5442 , U2391 , U5409 );
nand NAND2_3095 ( U5443 , INSTQUEUE_REG_0__1_ , U5404 );
nand NAND2_3096 ( U5444 , U5394 , U2417 );
nand NAND2_3097 ( U5445 , U2516 , U2399 );
nand NAND2_3098 ( U5446 , U5393 , U2398 );
nand NAND2_3099 ( U5447 , U2390 , U5409 );
nand NAND2_3100 ( U5448 , INSTQUEUE_REG_0__0_ , U5404 );
not NOT1_3101 ( U5449 , U3410 );
nand NAND3_3102 ( U5450 , U3378 , U3381 , U4491 );
nand NAND3_3103 ( U5451 , U4388 , U4161 , U4448 );
not NOT1_3104 ( U5452 , U3231 );
nand NAND2_3105 ( U5453 , U4482 , U3276 );
nand NAND3_3106 ( U5454 , U5453 , U3270 , U5452 );
nand NAND2_3107 ( U5455 , U3720 , U2452 );
nand NAND2_3108 ( U5456 , U4196 , U5450 );
nand NAND2_3109 ( U5457 , U3721 , U7597 );
nand NAND3_3110 ( U5458 , U4203 , U3244 , GTE_485_U6 );
nand NAND2_3111 ( U5459 , U2449 , U7482 );
nand NAND2_3112 ( U5460 , U4245 , U4491 );
not NOT1_3113 ( U5461 , U4170 );
nand NAND2_3114 ( U5462 , U2368 , U4170 );
nand NAND2_3115 ( U5463 , STATE2_REG_3_ , U3281 );
not NOT1_3116 ( U5464 , U4160 );
nand NAND2_3117 ( U5465 , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_3118 ( U5466 , INSTQUEUERD_ADDR_REG_3_ , U5465 );
nand NAND2_3119 ( U5467 , U4369 , INSTQUEUERD_ADDR_REG_1_ );
not NOT1_3120 ( U5468 , U3429 );
nand NAND2_3121 ( U5469 , U3486 , INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_3122 ( U5470 , INSTQUEUERD_ADDR_REG_3_ , U5469 );
not NOT1_3123 ( U5471 , U3425 );
nand NAND2_3124 ( U5472 , U3262 , U3251 );
nand NAND2_3125 ( U5473 , INSTQUEUERD_ADDR_REG_3_ , U5472 );
nand NAND2_3126 ( U5474 , U2469 , U3262 );
nand NAND2_3127 ( U5475 , U4482 , U3277 );
nand NAND2_3128 ( U5476 , U4388 , U2605 );
nand NAND3_3129 ( U5477 , U7692 , U7691 , U7482 );
nand NAND2_3130 ( U5478 , U4437 , U5476 );
nand NAND3_3131 ( U5479 , U4388 , U3381 , U3396 );
nand NAND2_3132 ( U5480 , U5479 , U4159 );
nand NAND2_3133 ( U5481 , U7617 , U5480 );
nand NAND2_3134 ( U5482 , U4448 , U4159 );
nand NAND2_3135 ( U5483 , U3382 , U5482 );
nand NAND2_3136 ( U5484 , U4196 , U5450 );
nand NAND2_3137 ( U5485 , U4245 , U4491 );
nand NAND2_3138 ( U5486 , U5483 , U3258 );
nand NAND2_3139 ( U5487 , U4482 , U7695 );
nand NAND2_3140 ( U5488 , U4178 , U3231 );
nand NAND2_3141 ( U5489 , U3279 , U4205 );
nand NAND2_3142 ( U5490 , U3728 , U5489 );
nand NAND2_3143 ( U5491 , R2182_U25 , U7497 );
nand NAND2_3144 ( U5492 , U4206 , U3425 );
nand NAND2_3145 ( U5493 , U4202 , U3429 );
nand NAND2_3146 ( U5494 , U5491 , U3735 );
nand NAND2_3147 ( U5495 , U4240 , U3425 );
nand NAND2_3148 ( U5496 , U2427 , U5494 );
nand NAND2_3149 ( U5497 , U5496 , U5495 );
nand NAND2_3150 ( U5498 , INSTQUEUERD_ADDR_REG_2_ , U3262 );
not NOT1_3151 ( U5499 , U3388 );
nand NAND2_3152 ( U5500 , R2182_U42 , U7497 );
nand NAND2_3153 ( U5501 , U4202 , U3443 );
nand NAND2_3154 ( U5502 , U3737 , U5500 );
nand NAND2_3155 ( U5503 , U2446 , U3457 );
nand NAND2_3156 ( U5504 , U4240 , U3388 );
nand NAND2_3157 ( U5505 , U2427 , U5502 );
nand NAND3_3158 ( U5506 , U5505 , U5503 , U5504 );
not NOT1_3159 ( U5507 , U3389 );
nand NAND2_3160 ( U5508 , U2431 , U4237 );
nand NAND2_3161 ( U5509 , U3279 , U5508 );
nand NAND2_3162 ( U5510 , U5507 , U5509 );
nand NAND2_3163 ( U5511 , R2182_U33 , U7497 );
nand NAND2_3164 ( U5512 , U4202 , U3252 );
nand NAND2_3165 ( U5513 , U3738 , U5511 );
nand NAND2_3166 ( U5514 , U7700 , U2446 );
nand NAND2_3167 ( U5515 , U5507 , U4240 );
nand NAND2_3168 ( U5516 , U2427 , U5513 );
nand NAND3_3169 ( U5517 , U5516 , U5514 , U5515 );
nand NAND2_3170 ( U5518 , R2182_U34 , U7497 );
nand NAND2_3171 ( U5519 , U4163 , U5518 );
nand NAND2_3172 ( U5520 , U4240 , U3253 );
nand NAND2_3173 ( U5521 , U2427 , U5519 );
nand NAND2_3174 ( U5522 , U7703 , STATE2_REG_1_ );
nand NAND3_3175 ( U5523 , U5521 , U5522 , U5520 );
nand NAND3_3176 ( U5524 , U2428 , STATE2_REG_0_ , LT_589_U6 );
not NOT1_3177 ( U5525 , U3391 );
nand NAND2_3178 ( U5526 , STATE2_REG_1_ , U3283 );
nand NAND2_3179 ( U5527 , U4515 , U3441 );
nand NAND2_3180 ( U5528 , U3345 , U5527 );
nand NAND2_3181 ( U5529 , U3346 , U5528 );
nand NAND2_3182 ( U5530 , U2388 , U5529 );
nand NAND2_3183 ( U5531 , R2182_U25 , U5526 );
nand NAND2_3184 ( U5532 , U4214 , R2144_U8 );
nand NAND2_3185 ( U5533 , U3739 , U5530 );
nand NAND2_3186 ( U5534 , U2388 , U7721 );
nand NAND2_3187 ( U5535 , R2182_U42 , U5526 );
nand NAND2_3188 ( U5536 , U4214 , R2144_U49 );
nand NAND2_3189 ( U5537 , U3740 , U5534 );
nand NAND2_3190 ( U5538 , U3313 , U3320 );
nand NAND2_3191 ( U5539 , U2388 , U5538 );
nand NAND2_3192 ( U5540 , R2182_U33 , U5526 );
nand NAND2_3193 ( U5541 , U4214 , R2144_U50 );
nand NAND2_3194 ( U5542 , U3741 , U5539 );
nand NAND2_3195 ( U5543 , R2182_U34 , U5526 );
nand NAND2_3196 ( U5544 , R2144_U43 , U4197 );
nand NAND3_3197 ( U5545 , U5543 , U5544 , U4233 );
nand NAND2_3198 ( U5546 , U4465 , U3259 );
nand NAND2_3199 ( U5547 , U4248 , U2431 );
nand NAND4_3200 ( U5548 , U2518 , U5547 , U7731 , U7730 );
nand NAND3_3201 ( U5549 , U4223 , U4491 , U4180 );
nand NAND2_3202 ( U5550 , U2368 , U5548 );
nand NAND2_3203 ( U5551 , U4191 , U3250 );
not NOT1_3204 ( U5552 , U3401 );
nand NAND2_3205 ( U5553 , U4250 , U4196 );
nand NAND2_3206 ( U5554 , U4244 , U2389 );
nand NAND2_3207 ( U5555 , U4254 , U4238 );
nand NAND2_3208 ( U5556 , U4252 , U4482 );
nand NAND2_3209 ( U5557 , U3746 , U2519 );
nand NAND2_3210 ( U5558 , R2099_U86 , U2380 );
nand NAND2_3211 ( U5559 , R2027_U5 , U2378 );
nand NAND2_3212 ( U5560 , R2278_U17 , U2377 );
nand NAND2_3213 ( U5561 , ADD_405_U4 , U2375 );
nand NAND2_3214 ( U5562 , INSTADDRPOINTER_REG_0_ , U2374 );
nand NAND2_3215 ( U5563 , REIP_REG_0_ , U2370 );
nand NAND2_3216 ( U5564 , U5552 , INSTADDRPOINTER_REG_0_ );
nand NAND2_3217 ( U5565 , R2099_U87 , U2380 );
nand NAND2_3218 ( U5566 , R2027_U71 , U2378 );
nand NAND2_3219 ( U5567 , R2278_U42 , U2377 );
nand NAND2_3220 ( U5568 , ADD_405_U81 , U2375 );
nand NAND2_3221 ( U5569 , ADD_515_U4 , U2374 );
nand NAND2_3222 ( U5570 , U2370 , REIP_REG_1_ );
nand NAND2_3223 ( U5571 , U5552 , INSTADDRPOINTER_REG_1_ );
nand NAND2_3224 ( U5572 , R2099_U138 , U2380 );
nand NAND2_3225 ( U5573 , R2027_U60 , U2378 );
nand NAND2_3226 ( U5574 , R2278_U101 , U2377 );
nand NAND2_3227 ( U5575 , ADD_405_U5 , U2375 );
nand NAND2_3228 ( U5576 , ADD_515_U71 , U2374 );
nand NAND2_3229 ( U5577 , U2370 , REIP_REG_2_ );
nand NAND2_3230 ( U5578 , INSTADDRPOINTER_REG_2_ , U5552 );
nand NAND2_3231 ( U5579 , R2099_U42 , U2380 );
nand NAND2_3232 ( U5580 , R2027_U57 , U2378 );
nand NAND2_3233 ( U5581 , R2278_U92 , U2377 );
nand NAND2_3234 ( U5582 , ADD_405_U93 , U2375 );
nand NAND2_3235 ( U5583 , ADD_515_U68 , U2374 );
nand NAND2_3236 ( U5584 , U2370 , REIP_REG_3_ );
nand NAND2_3237 ( U5585 , INSTADDRPOINTER_REG_3_ , U5552 );
nand NAND2_3238 ( U5586 , R2099_U41 , U2380 );
nand NAND2_3239 ( U5587 , R2027_U56 , U2378 );
nand NAND2_3240 ( U5588 , R2278_U89 , U2377 );
nand NAND2_3241 ( U5589 , ADD_405_U68 , U2375 );
nand NAND2_3242 ( U5590 , ADD_515_U67 , U2374 );
nand NAND2_3243 ( U5591 , U2370 , REIP_REG_4_ );
nand NAND2_3244 ( U5592 , INSTADDRPOINTER_REG_4_ , U5552 );
nand NAND2_3245 ( U5593 , R2099_U40 , U2380 );
nand NAND2_3246 ( U5594 , R2027_U55 , U2378 );
nand NAND2_3247 ( U5595 , R2278_U86 , U2377 );
nand NAND2_3248 ( U5596 , ADD_405_U67 , U2375 );
nand NAND2_3249 ( U5597 , ADD_515_U66 , U2374 );
nand NAND2_3250 ( U5598 , U2370 , REIP_REG_5_ );
nand NAND2_3251 ( U5599 , INSTADDRPOINTER_REG_5_ , U5552 );
nand NAND2_3252 ( U5600 , R2099_U39 , U2380 );
nand NAND2_3253 ( U5601 , R2027_U54 , U2378 );
nand NAND2_3254 ( U5602 , R2278_U83 , U2377 );
nand NAND2_3255 ( U5603 , ADD_405_U66 , U2375 );
nand NAND2_3256 ( U5604 , ADD_515_U65 , U2374 );
nand NAND2_3257 ( U5605 , U2370 , REIP_REG_6_ );
nand NAND2_3258 ( U5606 , INSTADDRPOINTER_REG_6_ , U5552 );
nand NAND2_3259 ( U5607 , R2099_U38 , U2380 );
nand NAND2_3260 ( U5608 , R2027_U53 , U2378 );
nand NAND2_3261 ( U5609 , R2278_U80 , U2377 );
nand NAND2_3262 ( U5610 , ADD_405_U65 , U2375 );
nand NAND2_3263 ( U5611 , ADD_515_U64 , U2374 );
nand NAND2_3264 ( U5612 , U2370 , REIP_REG_7_ );
nand NAND2_3265 ( U5613 , INSTADDRPOINTER_REG_7_ , U5552 );
nand NAND2_3266 ( U5614 , R2099_U37 , U2380 );
nand NAND2_3267 ( U5615 , R2027_U52 , U2378 );
nand NAND2_3268 ( U5616 , R2278_U77 , U2377 );
nand NAND2_3269 ( U5617 , ADD_405_U64 , U2375 );
nand NAND2_3270 ( U5618 , ADD_515_U63 , U2374 );
nand NAND2_3271 ( U5619 , U2370 , REIP_REG_8_ );
nand NAND2_3272 ( U5620 , INSTADDRPOINTER_REG_8_ , U5552 );
nand NAND2_3273 ( U5621 , R2099_U36 , U2380 );
nand NAND2_3274 ( U5622 , R2027_U51 , U2378 );
nand NAND2_3275 ( U5623 , R2278_U74 , U2377 );
nand NAND2_3276 ( U5624 , ADD_405_U63 , U2375 );
nand NAND2_3277 ( U5625 , ADD_515_U62 , U2374 );
nand NAND2_3278 ( U5626 , U2370 , REIP_REG_9_ );
nand NAND2_3279 ( U5627 , INSTADDRPOINTER_REG_9_ , U5552 );
nand NAND2_3280 ( U5628 , R2099_U85 , U2380 );
nand NAND2_3281 ( U5629 , R2027_U81 , U2378 );
nand NAND2_3282 ( U5630 , R2278_U160 , U2377 );
nand NAND2_3283 ( U5631 , ADD_405_U91 , U2375 );
nand NAND2_3284 ( U5632 , ADD_515_U91 , U2374 );
nand NAND2_3285 ( U5633 , U2370 , REIP_REG_10_ );
nand NAND2_3286 ( U5634 , INSTADDRPOINTER_REG_10_ , U5552 );
nand NAND2_3287 ( U5635 , R2099_U84 , U2380 );
nand NAND2_3288 ( U5636 , R2027_U80 , U2378 );
nand NAND2_3289 ( U5637 , R2278_U157 , U2377 );
nand NAND2_3290 ( U5638 , ADD_405_U90 , U2375 );
nand NAND2_3291 ( U5639 , ADD_515_U90 , U2374 );
nand NAND2_3292 ( U5640 , U2370 , REIP_REG_11_ );
nand NAND2_3293 ( U5641 , INSTADDRPOINTER_REG_11_ , U5552 );
nand NAND2_3294 ( U5642 , R2099_U83 , U2380 );
nand NAND2_3295 ( U5643 , R2027_U79 , U2378 );
nand NAND2_3296 ( U5644 , R2278_U154 , U2377 );
nand NAND2_3297 ( U5645 , ADD_405_U89 , U2375 );
nand NAND2_3298 ( U5646 , ADD_515_U89 , U2374 );
nand NAND2_3299 ( U5647 , U2370 , REIP_REG_12_ );
nand NAND2_3300 ( U5648 , INSTADDRPOINTER_REG_12_ , U5552 );
nand NAND2_3301 ( U5649 , R2099_U82 , U2380 );
nand NAND2_3302 ( U5650 , R2027_U78 , U2378 );
nand NAND2_3303 ( U5651 , R2278_U151 , U2377 );
nand NAND2_3304 ( U5652 , ADD_405_U88 , U2375 );
nand NAND2_3305 ( U5653 , ADD_515_U88 , U2374 );
nand NAND2_3306 ( U5654 , U2370 , REIP_REG_13_ );
nand NAND2_3307 ( U5655 , INSTADDRPOINTER_REG_13_ , U5552 );
nand NAND2_3308 ( U5656 , R2099_U81 , U2380 );
nand NAND2_3309 ( U5657 , R2027_U77 , U2378 );
nand NAND2_3310 ( U5658 , R2278_U148 , U2377 );
nand NAND2_3311 ( U5659 , ADD_405_U87 , U2375 );
nand NAND2_3312 ( U5660 , ADD_515_U87 , U2374 );
nand NAND2_3313 ( U5661 , U2370 , REIP_REG_14_ );
nand NAND2_3314 ( U5662 , INSTADDRPOINTER_REG_14_ , U5552 );
nand NAND2_3315 ( U5663 , R2099_U80 , U2380 );
nand NAND2_3316 ( U5664 , R2027_U76 , U2378 );
nand NAND2_3317 ( U5665 , R2278_U145 , U2377 );
nand NAND2_3318 ( U5666 , ADD_405_U86 , U2375 );
nand NAND2_3319 ( U5667 , ADD_515_U86 , U2374 );
nand NAND2_3320 ( U5668 , U2370 , REIP_REG_15_ );
nand NAND2_3321 ( U5669 , INSTADDRPOINTER_REG_15_ , U5552 );
nand NAND2_3322 ( U5670 , R2099_U79 , U2380 );
nand NAND2_3323 ( U5671 , R2027_U75 , U2378 );
nand NAND2_3324 ( U5672 , R2278_U142 , U2377 );
nand NAND2_3325 ( U5673 , ADD_405_U85 , U2375 );
nand NAND2_3326 ( U5674 , ADD_515_U85 , U2374 );
nand NAND2_3327 ( U5675 , U2370 , REIP_REG_16_ );
nand NAND2_3328 ( U5676 , INSTADDRPOINTER_REG_16_ , U5552 );
nand NAND2_3329 ( U5677 , R2099_U78 , U2380 );
nand NAND2_3330 ( U5678 , R2027_U74 , U2378 );
nand NAND2_3331 ( U5679 , R2278_U139 , U2377 );
nand NAND2_3332 ( U5680 , ADD_405_U84 , U2375 );
nand NAND2_3333 ( U5681 , ADD_515_U84 , U2374 );
nand NAND2_3334 ( U5682 , U2370 , REIP_REG_17_ );
nand NAND2_3335 ( U5683 , INSTADDRPOINTER_REG_17_ , U5552 );
nand NAND2_3336 ( U5684 , R2099_U77 , U2380 );
nand NAND2_3337 ( U5685 , R2027_U73 , U2378 );
nand NAND2_3338 ( U5686 , R2278_U136 , U2377 );
nand NAND2_3339 ( U5687 , ADD_405_U83 , U2375 );
nand NAND2_3340 ( U5688 , ADD_515_U83 , U2374 );
nand NAND2_3341 ( U5689 , U2370 , REIP_REG_18_ );
nand NAND2_3342 ( U5690 , INSTADDRPOINTER_REG_18_ , U5552 );
nand NAND2_3343 ( U5691 , R2099_U76 , U2380 );
nand NAND2_3344 ( U5692 , R2027_U72 , U2378 );
nand NAND2_3345 ( U5693 , R2278_U133 , U2377 );
nand NAND2_3346 ( U5694 , ADD_405_U82 , U2375 );
nand NAND2_3347 ( U5695 , ADD_515_U82 , U2374 );
nand NAND2_3348 ( U5696 , U2370 , REIP_REG_19_ );
nand NAND2_3349 ( U5697 , INSTADDRPOINTER_REG_19_ , U5552 );
nand NAND2_3350 ( U5698 , R2099_U75 , U2380 );
nand NAND2_3351 ( U5699 , R2027_U70 , U2378 );
nand NAND2_3352 ( U5700 , R2278_U129 , U2377 );
nand NAND2_3353 ( U5701 , ADD_405_U80 , U2375 );
nand NAND2_3354 ( U5702 , ADD_515_U81 , U2374 );
nand NAND2_3355 ( U5703 , U2370 , REIP_REG_20_ );
nand NAND2_3356 ( U5704 , INSTADDRPOINTER_REG_20_ , U5552 );
nand NAND2_3357 ( U5705 , R2099_U74 , U2380 );
nand NAND2_3358 ( U5706 , R2027_U69 , U2378 );
nand NAND2_3359 ( U5707 , R2278_U126 , U2377 );
nand NAND2_3360 ( U5708 , ADD_405_U79 , U2375 );
nand NAND2_3361 ( U5709 , ADD_515_U80 , U2374 );
nand NAND2_3362 ( U5710 , U2370 , REIP_REG_21_ );
nand NAND2_3363 ( U5711 , INSTADDRPOINTER_REG_21_ , U5552 );
nand NAND2_3364 ( U5712 , R2099_U73 , U2380 );
nand NAND2_3365 ( U5713 , R2027_U68 , U2378 );
nand NAND2_3366 ( U5714 , R2278_U123 , U2377 );
nand NAND2_3367 ( U5715 , ADD_405_U78 , U2375 );
nand NAND2_3368 ( U5716 , ADD_515_U79 , U2374 );
nand NAND2_3369 ( U5717 , U2370 , REIP_REG_22_ );
nand NAND2_3370 ( U5718 , INSTADDRPOINTER_REG_22_ , U5552 );
nand NAND2_3371 ( U5719 , R2099_U72 , U2380 );
nand NAND2_3372 ( U5720 , R2027_U67 , U2378 );
nand NAND2_3373 ( U5721 , R2278_U120 , U2377 );
nand NAND2_3374 ( U5722 , ADD_405_U77 , U2375 );
nand NAND2_3375 ( U5723 , ADD_515_U78 , U2374 );
nand NAND2_3376 ( U5724 , U2370 , REIP_REG_23_ );
nand NAND2_3377 ( U5725 , INSTADDRPOINTER_REG_23_ , U5552 );
nand NAND2_3378 ( U5726 , R2099_U71 , U2380 );
nand NAND2_3379 ( U5727 , R2027_U66 , U2378 );
nand NAND2_3380 ( U5728 , R2278_U117 , U2377 );
nand NAND2_3381 ( U5729 , ADD_405_U76 , U2375 );
nand NAND2_3382 ( U5730 , ADD_515_U77 , U2374 );
nand NAND2_3383 ( U5731 , U2370 , REIP_REG_24_ );
nand NAND2_3384 ( U5732 , INSTADDRPOINTER_REG_24_ , U5552 );
nand NAND2_3385 ( U5733 , R2099_U70 , U2380 );
nand NAND2_3386 ( U5734 , R2027_U65 , U2378 );
nand NAND2_3387 ( U5735 , R2278_U114 , U2377 );
nand NAND2_3388 ( U5736 , ADD_405_U75 , U2375 );
nand NAND2_3389 ( U5737 , ADD_515_U76 , U2374 );
nand NAND2_3390 ( U5738 , U2370 , REIP_REG_25_ );
nand NAND2_3391 ( U5739 , INSTADDRPOINTER_REG_25_ , U5552 );
nand NAND2_3392 ( U5740 , R2099_U69 , U2380 );
nand NAND2_3393 ( U5741 , R2027_U64 , U2378 );
nand NAND2_3394 ( U5742 , R2278_U111 , U2377 );
nand NAND2_3395 ( U5743 , ADD_405_U74 , U2375 );
nand NAND2_3396 ( U5744 , ADD_515_U75 , U2374 );
nand NAND2_3397 ( U5745 , U2370 , REIP_REG_26_ );
nand NAND2_3398 ( U5746 , INSTADDRPOINTER_REG_26_ , U5552 );
nand NAND2_3399 ( U5747 , R2099_U68 , U2380 );
nand NAND2_3400 ( U5748 , R2027_U63 , U2378 );
nand NAND2_3401 ( U5749 , R2278_U108 , U2377 );
nand NAND2_3402 ( U5750 , ADD_405_U73 , U2375 );
nand NAND2_3403 ( U5751 , ADD_515_U74 , U2374 );
nand NAND2_3404 ( U5752 , U2370 , REIP_REG_27_ );
nand NAND2_3405 ( U5753 , INSTADDRPOINTER_REG_27_ , U5552 );
nand NAND2_3406 ( U5754 , R2099_U67 , U2380 );
nand NAND2_3407 ( U5755 , R2027_U62 , U2378 );
nand NAND2_3408 ( U5756 , R2278_U105 , U2377 );
nand NAND2_3409 ( U5757 , ADD_405_U72 , U2375 );
nand NAND2_3410 ( U5758 , ADD_515_U73 , U2374 );
nand NAND2_3411 ( U5759 , U2370 , REIP_REG_28_ );
nand NAND2_3412 ( U5760 , INSTADDRPOINTER_REG_28_ , U5552 );
nand NAND2_3413 ( U5761 , R2099_U66 , U2380 );
nand NAND2_3414 ( U5762 , R2027_U61 , U2378 );
nand NAND2_3415 ( U5763 , R2278_U103 , U2377 );
nand NAND2_3416 ( U5764 , ADD_405_U71 , U2375 );
nand NAND2_3417 ( U5765 , ADD_515_U72 , U2374 );
nand NAND2_3418 ( U5766 , U2370 , REIP_REG_29_ );
nand NAND2_3419 ( U5767 , INSTADDRPOINTER_REG_29_ , U5552 );
nand NAND2_3420 ( U5768 , R2099_U65 , U2380 );
nand NAND2_3421 ( U5769 , R2027_U59 , U2378 );
nand NAND2_3422 ( U5770 , R2278_U98 , U2377 );
nand NAND2_3423 ( U5771 , ADD_405_U70 , U2375 );
nand NAND2_3424 ( U5772 , ADD_515_U70 , U2374 );
nand NAND2_3425 ( U5773 , U2370 , REIP_REG_30_ );
nand NAND2_3426 ( U5774 , INSTADDRPOINTER_REG_30_ , U5552 );
nand NAND2_3427 ( U5775 , R2099_U64 , U2380 );
nand NAND2_3428 ( U5776 , R2027_U58 , U2378 );
nand NAND2_3429 ( U5777 , R2278_U96 , U2377 );
nand NAND2_3430 ( U5778 , ADD_405_U69 , U2375 );
nand NAND2_3431 ( U5779 , ADD_515_U69 , U2374 );
nand NAND2_3432 ( U5780 , U2370 , REIP_REG_31_ );
nand NAND2_3433 ( U5781 , INSTADDRPOINTER_REG_31_ , U5552 );
nand NAND2_3434 ( U5782 , U4197 , U3281 );
not NOT1_3435 ( U5783 , U3403 );
nand NAND2_3436 ( U5784 , STATE2_REG_2_ , U3281 );
nand NAND2_3437 ( U5785 , STATE2_REG_1_ , U3295 );
nand NAND2_3438 ( U5786 , U5785 , U5784 );
nand NAND2_3439 ( U5787 , PHYADDRPOINTER_REG_0_ , U2376 );
nand NAND2_3440 ( U5788 , U2372 , R2278_U17 );
nand NAND2_3441 ( U5789 , U2365 , REIP_REG_0_ );
nand NAND2_3442 ( U5790 , R2358_U82 , U2364 );
nand NAND2_3443 ( U5791 , PHYADDRPOINTER_REG_0_ , U5783 );
nand NAND2_3444 ( U5792 , R2337_U5 , U2376 );
nand NAND2_3445 ( U5793 , U2372 , R2278_U42 );
nand NAND2_3446 ( U5794 , U2365 , REIP_REG_1_ );
nand NAND2_3447 ( U5795 , R2358_U112 , U2364 );
nand NAND2_3448 ( U5796 , PHYADDRPOINTER_REG_1_ , U5783 );
nand NAND2_3449 ( U5797 , R2337_U60 , U2376 );
nand NAND2_3450 ( U5798 , U2372 , R2278_U101 );
nand NAND2_3451 ( U5799 , U2365 , REIP_REG_2_ );
nand NAND2_3452 ( U5800 , R2358_U19 , U2364 );
nand NAND2_3453 ( U5801 , PHYADDRPOINTER_REG_2_ , U5783 );
nand NAND2_3454 ( U5802 , R2337_U57 , U2376 );
nand NAND2_3455 ( U5803 , U2372 , R2278_U92 );
nand NAND2_3456 ( U5804 , U2365 , REIP_REG_3_ );
nand NAND2_3457 ( U5805 , R2358_U20 , U2364 );
nand NAND2_3458 ( U5806 , PHYADDRPOINTER_REG_3_ , U5783 );
nand NAND2_3459 ( U5807 , R2337_U56 , U2376 );
nand NAND2_3460 ( U5808 , U2372 , R2278_U89 );
nand NAND2_3461 ( U5809 , U2365 , REIP_REG_4_ );
nand NAND2_3462 ( U5810 , R2358_U90 , U2364 );
nand NAND2_3463 ( U5811 , PHYADDRPOINTER_REG_4_ , U5783 );
nand NAND2_3464 ( U5812 , R2337_U55 , U2376 );
nand NAND2_3465 ( U5813 , U2372 , R2278_U86 );
nand NAND2_3466 ( U5814 , U2365 , REIP_REG_5_ );
nand NAND2_3467 ( U5815 , R2358_U88 , U2364 );
nand NAND2_3468 ( U5816 , PHYADDRPOINTER_REG_5_ , U5783 );
nand NAND2_3469 ( U5817 , R2337_U54 , U2376 );
nand NAND2_3470 ( U5818 , U2372 , R2278_U83 );
nand NAND2_3471 ( U5819 , U2365 , REIP_REG_6_ );
nand NAND2_3472 ( U5820 , R2358_U86 , U2364 );
nand NAND2_3473 ( U5821 , PHYADDRPOINTER_REG_6_ , U5783 );
nand NAND2_3474 ( U5822 , R2337_U53 , U2376 );
nand NAND2_3475 ( U5823 , U2372 , R2278_U80 );
nand NAND2_3476 ( U5824 , U2365 , REIP_REG_7_ );
nand NAND2_3477 ( U5825 , R2358_U21 , U2364 );
nand NAND2_3478 ( U5826 , PHYADDRPOINTER_REG_7_ , U5783 );
nand NAND2_3479 ( U5827 , R2337_U52 , U2376 );
nand NAND2_3480 ( U5828 , U2372 , R2278_U77 );
nand NAND2_3481 ( U5829 , U2365 , REIP_REG_8_ );
nand NAND2_3482 ( U5830 , R2358_U85 , U2364 );
nand NAND2_3483 ( U5831 , PHYADDRPOINTER_REG_8_ , U5783 );
nand NAND2_3484 ( U5832 , R2337_U51 , U2376 );
nand NAND2_3485 ( U5833 , U2372 , R2278_U74 );
nand NAND2_3486 ( U5834 , U2365 , REIP_REG_9_ );
nand NAND2_3487 ( U5835 , R2358_U83 , U2364 );
nand NAND2_3488 ( U5836 , PHYADDRPOINTER_REG_9_ , U5783 );
nand NAND2_3489 ( U5837 , R2337_U80 , U2376 );
nand NAND2_3490 ( U5838 , U2372 , R2278_U160 );
nand NAND2_3491 ( U5839 , U2365 , REIP_REG_10_ );
nand NAND2_3492 ( U5840 , R2358_U14 , U2364 );
nand NAND2_3493 ( U5841 , PHYADDRPOINTER_REG_10_ , U5783 );
nand NAND2_3494 ( U5842 , R2337_U79 , U2376 );
nand NAND2_3495 ( U5843 , U2372 , R2278_U157 );
nand NAND2_3496 ( U5844 , U2365 , REIP_REG_11_ );
nand NAND2_3497 ( U5845 , R2358_U15 , U2364 );
nand NAND2_3498 ( U5846 , PHYADDRPOINTER_REG_11_ , U5783 );
nand NAND2_3499 ( U5847 , R2337_U78 , U2376 );
nand NAND2_3500 ( U5848 , U2372 , R2278_U154 );
nand NAND2_3501 ( U5849 , U2365 , REIP_REG_12_ );
nand NAND2_3502 ( U5850 , R2358_U122 , U2364 );
nand NAND2_3503 ( U5851 , PHYADDRPOINTER_REG_12_ , U5783 );
nand NAND2_3504 ( U5852 , R2337_U77 , U2376 );
nand NAND2_3505 ( U5853 , U2372 , R2278_U151 );
nand NAND2_3506 ( U5854 , U2365 , REIP_REG_13_ );
nand NAND2_3507 ( U5855 , R2358_U120 , U2364 );
nand NAND2_3508 ( U5856 , PHYADDRPOINTER_REG_13_ , U5783 );
nand NAND2_3509 ( U5857 , R2337_U76 , U2376 );
nand NAND2_3510 ( U5858 , U2372 , R2278_U148 );
nand NAND2_3511 ( U5859 , U2365 , REIP_REG_14_ );
nand NAND2_3512 ( U5860 , R2358_U119 , U2364 );
nand NAND2_3513 ( U5861 , PHYADDRPOINTER_REG_14_ , U5783 );
nand NAND2_3514 ( U5862 , R2337_U75 , U2376 );
nand NAND2_3515 ( U5863 , U2372 , R2278_U145 );
nand NAND2_3516 ( U5864 , U2365 , REIP_REG_15_ );
nand NAND2_3517 ( U5865 , R2358_U16 , U2364 );
nand NAND2_3518 ( U5866 , PHYADDRPOINTER_REG_15_ , U5783 );
nand NAND2_3519 ( U5867 , R2337_U74 , U2376 );
nand NAND2_3520 ( U5868 , U2372 , R2278_U142 );
nand NAND2_3521 ( U5869 , U2365 , REIP_REG_16_ );
nand NAND2_3522 ( U5870 , R2358_U17 , U2364 );
nand NAND2_3523 ( U5871 , PHYADDRPOINTER_REG_16_ , U5783 );
nand NAND2_3524 ( U5872 , R2337_U73 , U2376 );
nand NAND2_3525 ( U5873 , U2372 , R2278_U139 );
nand NAND2_3526 ( U5874 , U2365 , REIP_REG_17_ );
nand NAND2_3527 ( U5875 , R2358_U118 , U2364 );
nand NAND2_3528 ( U5876 , PHYADDRPOINTER_REG_17_ , U5783 );
nand NAND2_3529 ( U5877 , R2337_U72 , U2376 );
nand NAND2_3530 ( U5878 , U2372 , R2278_U136 );
nand NAND2_3531 ( U5879 , U2365 , REIP_REG_18_ );
nand NAND2_3532 ( U5880 , R2358_U116 , U2364 );
nand NAND2_3533 ( U5881 , PHYADDRPOINTER_REG_18_ , U5783 );
nand NAND2_3534 ( U5882 , R2337_U71 , U2376 );
nand NAND2_3535 ( U5883 , U2372 , R2278_U133 );
nand NAND2_3536 ( U5884 , U2365 , REIP_REG_19_ );
nand NAND2_3537 ( U5885 , R2358_U114 , U2364 );
nand NAND2_3538 ( U5886 , PHYADDRPOINTER_REG_19_ , U5783 );
nand NAND2_3539 ( U5887 , R2337_U70 , U2376 );
nand NAND2_3540 ( U5888 , U2372 , R2278_U129 );
nand NAND2_3541 ( U5889 , U2365 , REIP_REG_20_ );
nand NAND2_3542 ( U5890 , R2358_U110 , U2364 );
nand NAND2_3543 ( U5891 , PHYADDRPOINTER_REG_20_ , U5783 );
nand NAND2_3544 ( U5892 , R2337_U69 , U2376 );
nand NAND2_3545 ( U5893 , U2372 , R2278_U126 );
nand NAND2_3546 ( U5894 , U2365 , REIP_REG_21_ );
nand NAND2_3547 ( U5895 , R2358_U18 , U2364 );
nand NAND2_3548 ( U5896 , PHYADDRPOINTER_REG_21_ , U5783 );
nand NAND2_3549 ( U5897 , R2337_U68 , U2376 );
nand NAND2_3550 ( U5898 , U2372 , R2278_U123 );
nand NAND2_3551 ( U5899 , U2365 , REIP_REG_22_ );
nand NAND2_3552 ( U5900 , R2358_U109 , U2364 );
nand NAND2_3553 ( U5901 , PHYADDRPOINTER_REG_22_ , U5783 );
nand NAND2_3554 ( U5902 , R2337_U67 , U2376 );
nand NAND2_3555 ( U5903 , U2372 , R2278_U120 );
nand NAND2_3556 ( U5904 , U2365 , REIP_REG_23_ );
nand NAND2_3557 ( U5905 , R2358_U107 , U2364 );
nand NAND2_3558 ( U5906 , PHYADDRPOINTER_REG_23_ , U5783 );
nand NAND2_3559 ( U5907 , R2337_U66 , U2376 );
nand NAND2_3560 ( U5908 , U2372 , R2278_U117 );
nand NAND2_3561 ( U5909 , U2365 , REIP_REG_24_ );
nand NAND2_3562 ( U5910 , R2358_U105 , U2364 );
nand NAND2_3563 ( U5911 , PHYADDRPOINTER_REG_24_ , U5783 );
nand NAND2_3564 ( U5912 , R2337_U65 , U2376 );
nand NAND2_3565 ( U5913 , U2372 , R2278_U114 );
nand NAND2_3566 ( U5914 , U2365 , REIP_REG_25_ );
nand NAND2_3567 ( U5915 , R2358_U103 , U2364 );
nand NAND2_3568 ( U5916 , PHYADDRPOINTER_REG_25_ , U5783 );
nand NAND2_3569 ( U5917 , R2337_U64 , U2376 );
nand NAND2_3570 ( U5918 , U2372 , R2278_U111 );
nand NAND2_3571 ( U5919 , U2365 , REIP_REG_26_ );
nand NAND2_3572 ( U5920 , R2358_U101 , U2364 );
nand NAND2_3573 ( U5921 , PHYADDRPOINTER_REG_26_ , U5783 );
nand NAND2_3574 ( U5922 , R2337_U63 , U2376 );
nand NAND2_3575 ( U5923 , U2372 , R2278_U108 );
nand NAND2_3576 ( U5924 , U2365 , REIP_REG_27_ );
nand NAND2_3577 ( U5925 , R2358_U99 , U2364 );
nand NAND2_3578 ( U5926 , PHYADDRPOINTER_REG_27_ , U5783 );
nand NAND2_3579 ( U5927 , R2337_U62 , U2376 );
nand NAND2_3580 ( U5928 , U2372 , R2278_U105 );
nand NAND2_3581 ( U5929 , U2365 , REIP_REG_28_ );
nand NAND2_3582 ( U5930 , R2358_U97 , U2364 );
nand NAND2_3583 ( U5931 , PHYADDRPOINTER_REG_28_ , U5783 );
nand NAND2_3584 ( U5932 , R2337_U61 , U2376 );
nand NAND2_3585 ( U5933 , U2372 , R2278_U103 );
nand NAND2_3586 ( U5934 , U2365 , REIP_REG_29_ );
nand NAND2_3587 ( U5935 , R2358_U95 , U2364 );
nand NAND2_3588 ( U5936 , PHYADDRPOINTER_REG_29_ , U5783 );
nand NAND2_3589 ( U5937 , R2337_U59 , U2376 );
nand NAND2_3590 ( U5938 , U2372 , R2278_U98 );
nand NAND2_3591 ( U5939 , U2365 , REIP_REG_30_ );
nand NAND2_3592 ( U5940 , R2358_U93 , U2364 );
nand NAND2_3593 ( U5941 , PHYADDRPOINTER_REG_30_ , U5783 );
nand NAND2_3594 ( U5942 , R2337_U58 , U2376 );
nand NAND2_3595 ( U5943 , U2372 , R2278_U96 );
nand NAND2_3596 ( U5944 , U2365 , REIP_REG_31_ );
nand NAND2_3597 ( U5945 , R2358_U91 , U2364 );
nand NAND2_3598 ( U5946 , PHYADDRPOINTER_REG_31_ , U5783 );
nand NAND2_3599 ( U5947 , READY_N , U3269 );
nand NAND2_3600 ( U5948 , EAX_REG_15_ , U2382 );
nand NAND2_3601 ( U5949 , DATAI_15_ , U2381 );
nand NAND2_3602 ( U5950 , U5949 , U5948 );
nand NAND2_3603 ( U5951 , EAX_REG_14_ , U2382 );
nand NAND2_3604 ( U5952 , DATAI_14_ , U2381 );
nand NAND2_3605 ( U5953 , U5952 , U5951 );
nand NAND2_3606 ( U5954 , EAX_REG_13_ , U2382 );
nand NAND2_3607 ( U5955 , DATAI_13_ , U2381 );
nand NAND2_3608 ( U5956 , U5955 , U5954 );
nand NAND2_3609 ( U5957 , EAX_REG_12_ , U2382 );
nand NAND2_3610 ( U5958 , DATAI_12_ , U2381 );
nand NAND2_3611 ( U5959 , U5958 , U5957 );
nand NAND2_3612 ( U5960 , EAX_REG_11_ , U2382 );
nand NAND2_3613 ( U5961 , DATAI_11_ , U2381 );
nand NAND2_3614 ( U5962 , U5961 , U5960 );
nand NAND2_3615 ( U5963 , EAX_REG_10_ , U2382 );
nand NAND2_3616 ( U5964 , DATAI_10_ , U2381 );
nand NAND2_3617 ( U5965 , U5964 , U5963 );
nand NAND2_3618 ( U5966 , EAX_REG_9_ , U2382 );
nand NAND2_3619 ( U5967 , DATAI_9_ , U2381 );
nand NAND2_3620 ( U5968 , U5967 , U5966 );
nand NAND2_3621 ( U5969 , EAX_REG_8_ , U2382 );
nand NAND2_3622 ( U5970 , DATAI_8_ , U2381 );
nand NAND2_3623 ( U5971 , U5970 , U5969 );
nand NAND2_3624 ( U5972 , EAX_REG_7_ , U2382 );
nand NAND2_3625 ( U5973 , U2381 , DATAI_7_ );
nand NAND2_3626 ( U5974 , U5973 , U5972 );
nand NAND2_3627 ( U5975 , EAX_REG_6_ , U2382 );
nand NAND2_3628 ( U5976 , U2381 , DATAI_6_ );
nand NAND2_3629 ( U5977 , U5976 , U5975 );
nand NAND2_3630 ( U5978 , EAX_REG_5_ , U2382 );
nand NAND2_3631 ( U5979 , U2381 , DATAI_5_ );
nand NAND2_3632 ( U5980 , U5979 , U5978 );
nand NAND2_3633 ( U5981 , EAX_REG_4_ , U2382 );
nand NAND2_3634 ( U5982 , U2381 , DATAI_4_ );
nand NAND2_3635 ( U5983 , U5982 , U5981 );
nand NAND2_3636 ( U5984 , EAX_REG_3_ , U2382 );
nand NAND2_3637 ( U5985 , U2381 , DATAI_3_ );
nand NAND2_3638 ( U5986 , U5985 , U5984 );
nand NAND2_3639 ( U5987 , EAX_REG_2_ , U2382 );
nand NAND2_3640 ( U5988 , U2381 , DATAI_2_ );
nand NAND2_3641 ( U5989 , U5988 , U5987 );
nand NAND2_3642 ( U5990 , EAX_REG_1_ , U2382 );
nand NAND2_3643 ( U5991 , U2381 , DATAI_1_ );
nand NAND2_3644 ( U5992 , U5991 , U5990 );
nand NAND2_3645 ( U5993 , EAX_REG_0_ , U2382 );
nand NAND2_3646 ( U5994 , U2381 , DATAI_0_ );
nand NAND2_3647 ( U5995 , U5994 , U5993 );
nand NAND2_3648 ( U5996 , EAX_REG_30_ , U2382 );
nand NAND2_3649 ( U5997 , DATAI_14_ , U2381 );
nand NAND2_3650 ( U5998 , U5997 , U5996 );
nand NAND2_3651 ( U5999 , EAX_REG_29_ , U2382 );
nand NAND2_3652 ( U6000 , DATAI_13_ , U2381 );
nand NAND2_3653 ( U6001 , U6000 , U5999 );
nand NAND2_3654 ( U6002 , EAX_REG_28_ , U2382 );
nand NAND2_3655 ( U6003 , DATAI_12_ , U2381 );
nand NAND2_3656 ( U6004 , U6003 , U6002 );
nand NAND2_3657 ( U6005 , EAX_REG_27_ , U2382 );
nand NAND2_3658 ( U6006 , DATAI_11_ , U2381 );
nand NAND2_3659 ( U6007 , U6006 , U6005 );
nand NAND2_3660 ( U6008 , EAX_REG_26_ , U2382 );
nand NAND2_3661 ( U6009 , DATAI_10_ , U2381 );
nand NAND2_3662 ( U6010 , U6009 , U6008 );
nand NAND2_3663 ( U6011 , EAX_REG_25_ , U2382 );
nand NAND2_3664 ( U6012 , DATAI_9_ , U2381 );
nand NAND2_3665 ( U6013 , U6012 , U6011 );
nand NAND2_3666 ( U6014 , EAX_REG_24_ , U2382 );
nand NAND2_3667 ( U6015 , DATAI_8_ , U2381 );
nand NAND2_3668 ( U6016 , U6015 , U6014 );
nand NAND2_3669 ( U6017 , EAX_REG_23_ , U2382 );
nand NAND2_3670 ( U6018 , U2381 , DATAI_7_ );
nand NAND2_3671 ( U6019 , U6018 , U6017 );
nand NAND2_3672 ( U6020 , EAX_REG_22_ , U2382 );
nand NAND2_3673 ( U6021 , U2381 , DATAI_6_ );
nand NAND2_3674 ( U6022 , U6021 , U6020 );
nand NAND2_3675 ( U6023 , EAX_REG_21_ , U2382 );
nand NAND2_3676 ( U6024 , U2381 , DATAI_5_ );
nand NAND2_3677 ( U6025 , U6024 , U6023 );
nand NAND2_3678 ( U6026 , EAX_REG_20_ , U2382 );
nand NAND2_3679 ( U6027 , U2381 , DATAI_4_ );
nand NAND2_3680 ( U6028 , U6027 , U6026 );
nand NAND2_3681 ( U6029 , EAX_REG_19_ , U2382 );
nand NAND2_3682 ( U6030 , U2381 , DATAI_3_ );
nand NAND2_3683 ( U6031 , U6030 , U6029 );
nand NAND2_3684 ( U6032 , EAX_REG_18_ , U2382 );
nand NAND2_3685 ( U6033 , U2381 , DATAI_2_ );
nand NAND2_3686 ( U6034 , U6033 , U6032 );
nand NAND2_3687 ( U6035 , EAX_REG_17_ , U2382 );
nand NAND2_3688 ( U6036 , U2381 , DATAI_1_ );
nand NAND2_3689 ( U6037 , U6036 , U6035 );
nand NAND2_3690 ( U6038 , EAX_REG_16_ , U2382 );
nand NAND2_3691 ( U6039 , U2381 , DATAI_0_ );
nand NAND2_3692 ( U6040 , U6039 , U6038 );
nand NAND3_3693 ( U6041 , U4223 , U7594 , U4247 );
nand NAND2_3694 ( U6042 , U2428 , U3281 );
not NOT1_3695 ( U6043 , U3404 );
nand NAND2_3696 ( U6044 , U2385 , LWORD_REG_0_ );
nand NAND2_3697 ( U6045 , U2384 , EAX_REG_0_ );
nand NAND2_3698 ( U6046 , DATAO_REG_0_ , U6043 );
nand NAND2_3699 ( U6047 , U2385 , LWORD_REG_1_ );
nand NAND2_3700 ( U6048 , U2384 , EAX_REG_1_ );
nand NAND2_3701 ( U6049 , DATAO_REG_1_ , U6043 );
nand NAND2_3702 ( U6050 , U2385 , LWORD_REG_2_ );
nand NAND2_3703 ( U6051 , U2384 , EAX_REG_2_ );
nand NAND2_3704 ( U6052 , DATAO_REG_2_ , U6043 );
nand NAND2_3705 ( U6053 , U2385 , LWORD_REG_3_ );
nand NAND2_3706 ( U6054 , U2384 , EAX_REG_3_ );
nand NAND2_3707 ( U6055 , DATAO_REG_3_ , U6043 );
nand NAND2_3708 ( U6056 , U2385 , LWORD_REG_4_ );
nand NAND2_3709 ( U6057 , U2384 , EAX_REG_4_ );
nand NAND2_3710 ( U6058 , DATAO_REG_4_ , U6043 );
nand NAND2_3711 ( U6059 , U2385 , LWORD_REG_5_ );
nand NAND2_3712 ( U6060 , U2384 , EAX_REG_5_ );
nand NAND2_3713 ( U6061 , DATAO_REG_5_ , U6043 );
nand NAND2_3714 ( U6062 , U2385 , LWORD_REG_6_ );
nand NAND2_3715 ( U6063 , U2384 , EAX_REG_6_ );
nand NAND2_3716 ( U6064 , DATAO_REG_6_ , U6043 );
nand NAND2_3717 ( U6065 , U2385 , LWORD_REG_7_ );
nand NAND2_3718 ( U6066 , U2384 , EAX_REG_7_ );
nand NAND2_3719 ( U6067 , DATAO_REG_7_ , U6043 );
nand NAND2_3720 ( U6068 , U2385 , LWORD_REG_8_ );
nand NAND2_3721 ( U6069 , U2384 , EAX_REG_8_ );
nand NAND2_3722 ( U6070 , DATAO_REG_8_ , U6043 );
nand NAND2_3723 ( U6071 , U2385 , LWORD_REG_9_ );
nand NAND2_3724 ( U6072 , U2384 , EAX_REG_9_ );
nand NAND2_3725 ( U6073 , DATAO_REG_9_ , U6043 );
nand NAND2_3726 ( U6074 , U2385 , LWORD_REG_10_ );
nand NAND2_3727 ( U6075 , U2384 , EAX_REG_10_ );
nand NAND2_3728 ( U6076 , DATAO_REG_10_ , U6043 );
nand NAND2_3729 ( U6077 , U2385 , LWORD_REG_11_ );
nand NAND2_3730 ( U6078 , U2384 , EAX_REG_11_ );
nand NAND2_3731 ( U6079 , DATAO_REG_11_ , U6043 );
nand NAND2_3732 ( U6080 , U2385 , LWORD_REG_12_ );
nand NAND2_3733 ( U6081 , U2384 , EAX_REG_12_ );
nand NAND2_3734 ( U6082 , DATAO_REG_12_ , U6043 );
nand NAND2_3735 ( U6083 , U2385 , LWORD_REG_13_ );
nand NAND2_3736 ( U6084 , U2384 , EAX_REG_13_ );
nand NAND2_3737 ( U6085 , DATAO_REG_13_ , U6043 );
nand NAND2_3738 ( U6086 , U2385 , LWORD_REG_14_ );
nand NAND2_3739 ( U6087 , U2384 , EAX_REG_14_ );
nand NAND2_3740 ( U6088 , DATAO_REG_14_ , U6043 );
nand NAND2_3741 ( U6089 , U2385 , LWORD_REG_15_ );
nand NAND2_3742 ( U6090 , U2384 , EAX_REG_15_ );
nand NAND2_3743 ( U6091 , DATAO_REG_15_ , U6043 );
nand NAND2_3744 ( U6092 , U2424 , EAX_REG_16_ );
nand NAND2_3745 ( U6093 , U2385 , UWORD_REG_0_ );
nand NAND2_3746 ( U6094 , DATAO_REG_16_ , U6043 );
nand NAND2_3747 ( U6095 , U2424 , EAX_REG_17_ );
nand NAND2_3748 ( U6096 , U2385 , UWORD_REG_1_ );
nand NAND2_3749 ( U6097 , DATAO_REG_17_ , U6043 );
nand NAND2_3750 ( U6098 , U2424 , EAX_REG_18_ );
nand NAND2_3751 ( U6099 , U2385 , UWORD_REG_2_ );
nand NAND2_3752 ( U6100 , DATAO_REG_18_ , U6043 );
nand NAND2_3753 ( U6101 , U2424 , EAX_REG_19_ );
nand NAND2_3754 ( U6102 , U2385 , UWORD_REG_3_ );
nand NAND2_3755 ( U6103 , DATAO_REG_19_ , U6043 );
nand NAND2_3756 ( U6104 , U2424 , EAX_REG_20_ );
nand NAND2_3757 ( U6105 , U2385 , UWORD_REG_4_ );
nand NAND2_3758 ( U6106 , DATAO_REG_20_ , U6043 );
nand NAND2_3759 ( U6107 , U2424 , EAX_REG_21_ );
nand NAND2_3760 ( U6108 , U2385 , UWORD_REG_5_ );
nand NAND2_3761 ( U6109 , DATAO_REG_21_ , U6043 );
nand NAND2_3762 ( U6110 , U2424 , EAX_REG_22_ );
nand NAND2_3763 ( U6111 , U2385 , UWORD_REG_6_ );
nand NAND2_3764 ( U6112 , DATAO_REG_22_ , U6043 );
nand NAND2_3765 ( U6113 , U2424 , EAX_REG_23_ );
nand NAND2_3766 ( U6114 , U2385 , UWORD_REG_7_ );
nand NAND2_3767 ( U6115 , DATAO_REG_23_ , U6043 );
nand NAND2_3768 ( U6116 , U2424 , EAX_REG_24_ );
nand NAND2_3769 ( U6117 , U2385 , UWORD_REG_8_ );
nand NAND2_3770 ( U6118 , DATAO_REG_24_ , U6043 );
nand NAND2_3771 ( U6119 , U2424 , EAX_REG_25_ );
nand NAND2_3772 ( U6120 , U2385 , UWORD_REG_9_ );
nand NAND2_3773 ( U6121 , DATAO_REG_25_ , U6043 );
nand NAND2_3774 ( U6122 , U2424 , EAX_REG_26_ );
nand NAND2_3775 ( U6123 , U2385 , UWORD_REG_10_ );
nand NAND2_3776 ( U6124 , DATAO_REG_26_ , U6043 );
nand NAND2_3777 ( U6125 , U2424 , EAX_REG_27_ );
nand NAND2_3778 ( U6126 , U2385 , UWORD_REG_11_ );
nand NAND2_3779 ( U6127 , DATAO_REG_27_ , U6043 );
nand NAND2_3780 ( U6128 , U2424 , EAX_REG_28_ );
nand NAND2_3781 ( U6129 , U2385 , UWORD_REG_12_ );
nand NAND2_3782 ( U6130 , DATAO_REG_28_ , U6043 );
nand NAND2_3783 ( U6131 , U2424 , EAX_REG_29_ );
nand NAND2_3784 ( U6132 , U2385 , UWORD_REG_13_ );
nand NAND2_3785 ( U6133 , DATAO_REG_29_ , U6043 );
nand NAND2_3786 ( U6134 , U2424 , EAX_REG_30_ );
nand NAND2_3787 ( U6135 , U2385 , UWORD_REG_14_ );
nand NAND2_3788 ( U6136 , DATAO_REG_30_ , U6043 );
nand NAND3_3789 ( U6137 , U4182 , U2447 , GTE_485_U6 );
nand NAND3_3790 ( U6138 , U4242 , U4185 , U4182 );
nand NAND3_3791 ( U6139 , U4188 , U3270 , R2167_U17 );
nand NAND2_3792 ( U6140 , U7491 , U3244 );
nand NAND2_3793 ( U6141 , U3871 , U6140 );
nand NAND2_3794 ( U6142 , U2422 , DATAI_0_ );
nand NAND2_3795 ( U6143 , U2386 , R2358_U82 );
nand NAND2_3796 ( U6144 , EAX_REG_0_ , U3411 );
nand NAND2_3797 ( U6145 , U2422 , DATAI_1_ );
nand NAND2_3798 ( U6146 , U2386 , R2358_U112 );
nand NAND2_3799 ( U6147 , EAX_REG_1_ , U3411 );
nand NAND2_3800 ( U6148 , U2422 , DATAI_2_ );
nand NAND2_3801 ( U6149 , U2386 , R2358_U19 );
nand NAND2_3802 ( U6150 , EAX_REG_2_ , U3411 );
nand NAND2_3803 ( U6151 , U2422 , DATAI_3_ );
nand NAND2_3804 ( U6152 , U2386 , R2358_U20 );
nand NAND2_3805 ( U6153 , EAX_REG_3_ , U3411 );
nand NAND2_3806 ( U6154 , U2422 , DATAI_4_ );
nand NAND2_3807 ( U6155 , U2386 , R2358_U90 );
nand NAND2_3808 ( U6156 , EAX_REG_4_ , U3411 );
nand NAND2_3809 ( U6157 , U2422 , DATAI_5_ );
nand NAND2_3810 ( U6158 , U2386 , R2358_U88 );
nand NAND2_3811 ( U6159 , EAX_REG_5_ , U3411 );
nand NAND2_3812 ( U6160 , U2422 , DATAI_6_ );
nand NAND2_3813 ( U6161 , U2386 , R2358_U86 );
nand NAND2_3814 ( U6162 , EAX_REG_6_ , U3411 );
nand NAND2_3815 ( U6163 , U2422 , DATAI_7_ );
nand NAND2_3816 ( U6164 , U2386 , R2358_U21 );
nand NAND2_3817 ( U6165 , EAX_REG_7_ , U3411 );
nand NAND2_3818 ( U6166 , U2422 , DATAI_8_ );
nand NAND2_3819 ( U6167 , U2386 , R2358_U85 );
nand NAND2_3820 ( U6168 , EAX_REG_8_ , U3411 );
nand NAND2_3821 ( U6169 , U2422 , DATAI_9_ );
nand NAND2_3822 ( U6170 , U2386 , R2358_U83 );
nand NAND2_3823 ( U6171 , EAX_REG_9_ , U3411 );
nand NAND2_3824 ( U6172 , U2422 , DATAI_10_ );
nand NAND2_3825 ( U6173 , U2386 , R2358_U14 );
nand NAND2_3826 ( U6174 , EAX_REG_10_ , U3411 );
nand NAND2_3827 ( U6175 , U2422 , DATAI_11_ );
nand NAND2_3828 ( U6176 , U2386 , R2358_U15 );
nand NAND2_3829 ( U6177 , EAX_REG_11_ , U3411 );
nand NAND2_3830 ( U6178 , U2422 , DATAI_12_ );
nand NAND2_3831 ( U6179 , U2386 , R2358_U122 );
nand NAND2_3832 ( U6180 , EAX_REG_12_ , U3411 );
nand NAND2_3833 ( U6181 , U2422 , DATAI_13_ );
nand NAND2_3834 ( U6182 , U2386 , R2358_U120 );
nand NAND2_3835 ( U6183 , EAX_REG_13_ , U3411 );
nand NAND2_3836 ( U6184 , U2422 , DATAI_14_ );
nand NAND2_3837 ( U6185 , U2386 , R2358_U119 );
nand NAND2_3838 ( U6186 , EAX_REG_14_ , U3411 );
nand NAND2_3839 ( U6187 , U2422 , DATAI_15_ );
nand NAND2_3840 ( U6188 , U2386 , R2358_U16 );
nand NAND2_3841 ( U6189 , EAX_REG_15_ , U3411 );
nand NAND2_3842 ( U6190 , U2423 , DATAI_16_ );
nand NAND2_3843 ( U6191 , U2387 , DATAI_0_ );
nand NAND2_3844 ( U6192 , U2386 , R2358_U17 );
nand NAND2_3845 ( U6193 , EAX_REG_16_ , U3411 );
nand NAND2_3846 ( U6194 , U2423 , DATAI_17_ );
nand NAND2_3847 ( U6195 , U2387 , DATAI_1_ );
nand NAND2_3848 ( U6196 , U2386 , R2358_U118 );
nand NAND2_3849 ( U6197 , EAX_REG_17_ , U3411 );
nand NAND2_3850 ( U6198 , U2423 , DATAI_18_ );
nand NAND2_3851 ( U6199 , U2387 , DATAI_2_ );
nand NAND2_3852 ( U6200 , U2386 , R2358_U116 );
nand NAND2_3853 ( U6201 , EAX_REG_18_ , U3411 );
nand NAND2_3854 ( U6202 , U2423 , DATAI_19_ );
nand NAND2_3855 ( U6203 , U2387 , DATAI_3_ );
nand NAND2_3856 ( U6204 , U2386 , R2358_U114 );
nand NAND2_3857 ( U6205 , EAX_REG_19_ , U3411 );
nand NAND2_3858 ( U6206 , U2423 , DATAI_20_ );
nand NAND2_3859 ( U6207 , U2387 , DATAI_4_ );
nand NAND2_3860 ( U6208 , U2386 , R2358_U110 );
nand NAND2_3861 ( U6209 , EAX_REG_20_ , U3411 );
nand NAND2_3862 ( U6210 , U2423 , DATAI_21_ );
nand NAND2_3863 ( U6211 , U2387 , DATAI_5_ );
nand NAND2_3864 ( U6212 , U2386 , R2358_U18 );
nand NAND2_3865 ( U6213 , EAX_REG_21_ , U3411 );
nand NAND2_3866 ( U6214 , U2423 , DATAI_22_ );
nand NAND2_3867 ( U6215 , U2387 , DATAI_6_ );
nand NAND2_3868 ( U6216 , U2386 , R2358_U109 );
nand NAND2_3869 ( U6217 , EAX_REG_22_ , U3411 );
nand NAND2_3870 ( U6218 , U2423 , DATAI_23_ );
nand NAND2_3871 ( U6219 , U2387 , DATAI_7_ );
nand NAND2_3872 ( U6220 , U2386 , R2358_U107 );
nand NAND2_3873 ( U6221 , EAX_REG_23_ , U3411 );
nand NAND2_3874 ( U6222 , U2423 , DATAI_24_ );
nand NAND2_3875 ( U6223 , U2387 , DATAI_8_ );
nand NAND2_3876 ( U6224 , U2386 , R2358_U105 );
nand NAND2_3877 ( U6225 , EAX_REG_24_ , U3411 );
nand NAND2_3878 ( U6226 , U2423 , DATAI_25_ );
nand NAND2_3879 ( U6227 , U2387 , DATAI_9_ );
nand NAND2_3880 ( U6228 , U2386 , R2358_U103 );
nand NAND2_3881 ( U6229 , EAX_REG_25_ , U3411 );
nand NAND2_3882 ( U6230 , U2423 , DATAI_26_ );
nand NAND2_3883 ( U6231 , U2387 , DATAI_10_ );
nand NAND2_3884 ( U6232 , U2386 , R2358_U101 );
nand NAND2_3885 ( U6233 , EAX_REG_26_ , U3411 );
nand NAND2_3886 ( U6234 , U2423 , DATAI_27_ );
nand NAND2_3887 ( U6235 , U2387 , DATAI_11_ );
nand NAND2_3888 ( U6236 , U2386 , R2358_U99 );
nand NAND2_3889 ( U6237 , EAX_REG_27_ , U3411 );
nand NAND2_3890 ( U6238 , U2423 , DATAI_28_ );
nand NAND2_3891 ( U6239 , U2387 , DATAI_12_ );
nand NAND2_3892 ( U6240 , U2386 , R2358_U97 );
nand NAND2_3893 ( U6241 , EAX_REG_28_ , U3411 );
nand NAND2_3894 ( U6242 , U2423 , DATAI_29_ );
nand NAND2_3895 ( U6243 , U2387 , DATAI_13_ );
nand NAND2_3896 ( U6244 , U2386 , R2358_U95 );
nand NAND2_3897 ( U6245 , EAX_REG_29_ , U3411 );
nand NAND2_3898 ( U6246 , U2423 , DATAI_30_ );
nand NAND2_3899 ( U6247 , U2387 , DATAI_14_ );
nand NAND2_3900 ( U6248 , U2386 , R2358_U93 );
nand NAND2_3901 ( U6249 , EAX_REG_30_ , U3411 );
nand NAND2_3902 ( U6250 , U2423 , DATAI_31_ );
nand NAND2_3903 ( U6251 , U4186 , U3260 );
nand NAND2_3904 ( U6252 , U4193 , U6251 );
nand NAND2_3905 ( U6253 , U2383 , R2358_U82 );
nand NAND2_3906 ( U6254 , U2371 , R2099_U86 );
nand NAND2_3907 ( U6255 , EBX_REG_0_ , U3413 );
nand NAND2_3908 ( U6256 , U2383 , R2358_U112 );
nand NAND2_3909 ( U6257 , U2371 , R2099_U87 );
nand NAND2_3910 ( U6258 , EBX_REG_1_ , U3413 );
nand NAND2_3911 ( U6259 , U2383 , R2358_U19 );
nand NAND2_3912 ( U6260 , U2371 , R2099_U138 );
nand NAND2_3913 ( U6261 , EBX_REG_2_ , U3413 );
nand NAND2_3914 ( U6262 , U2383 , R2358_U20 );
nand NAND2_3915 ( U6263 , U2371 , R2099_U42 );
nand NAND2_3916 ( U6264 , EBX_REG_3_ , U3413 );
nand NAND2_3917 ( U6265 , U2383 , R2358_U90 );
nand NAND2_3918 ( U6266 , U2371 , R2099_U41 );
nand NAND2_3919 ( U6267 , EBX_REG_4_ , U3413 );
nand NAND2_3920 ( U6268 , U2383 , R2358_U88 );
nand NAND2_3921 ( U6269 , U2371 , R2099_U40 );
nand NAND2_3922 ( U6270 , EBX_REG_5_ , U3413 );
nand NAND2_3923 ( U6271 , U2383 , R2358_U86 );
nand NAND2_3924 ( U6272 , U2371 , R2099_U39 );
nand NAND2_3925 ( U6273 , EBX_REG_6_ , U3413 );
nand NAND2_3926 ( U6274 , U2383 , R2358_U21 );
nand NAND2_3927 ( U6275 , U2371 , R2099_U38 );
nand NAND2_3928 ( U6276 , EBX_REG_7_ , U3413 );
nand NAND2_3929 ( U6277 , U2383 , R2358_U85 );
nand NAND2_3930 ( U6278 , U2371 , R2099_U37 );
nand NAND2_3931 ( U6279 , EBX_REG_8_ , U3413 );
nand NAND2_3932 ( U6280 , U2383 , R2358_U83 );
nand NAND2_3933 ( U6281 , U2371 , R2099_U36 );
nand NAND2_3934 ( U6282 , EBX_REG_9_ , U3413 );
nand NAND2_3935 ( U6283 , U2383 , R2358_U14 );
nand NAND2_3936 ( U6284 , U2371 , R2099_U85 );
nand NAND2_3937 ( U6285 , EBX_REG_10_ , U3413 );
nand NAND2_3938 ( U6286 , U2383 , R2358_U15 );
nand NAND2_3939 ( U6287 , U2371 , R2099_U84 );
nand NAND2_3940 ( U6288 , EBX_REG_11_ , U3413 );
nand NAND2_3941 ( U6289 , U2383 , R2358_U122 );
nand NAND2_3942 ( U6290 , U2371 , R2099_U83 );
nand NAND2_3943 ( U6291 , EBX_REG_12_ , U3413 );
nand NAND2_3944 ( U6292 , U2383 , R2358_U120 );
nand NAND2_3945 ( U6293 , U2371 , R2099_U82 );
nand NAND2_3946 ( U6294 , EBX_REG_13_ , U3413 );
nand NAND2_3947 ( U6295 , U2383 , R2358_U119 );
nand NAND2_3948 ( U6296 , U2371 , R2099_U81 );
nand NAND2_3949 ( U6297 , EBX_REG_14_ , U3413 );
nand NAND2_3950 ( U6298 , U2383 , R2358_U16 );
nand NAND2_3951 ( U6299 , U2371 , R2099_U80 );
nand NAND2_3952 ( U6300 , EBX_REG_15_ , U3413 );
nand NAND2_3953 ( U6301 , U2383 , R2358_U17 );
nand NAND2_3954 ( U6302 , U2371 , R2099_U79 );
nand NAND2_3955 ( U6303 , EBX_REG_16_ , U3413 );
nand NAND2_3956 ( U6304 , U2383 , R2358_U118 );
nand NAND2_3957 ( U6305 , U2371 , R2099_U78 );
nand NAND2_3958 ( U6306 , EBX_REG_17_ , U3413 );
nand NAND2_3959 ( U6307 , U2383 , R2358_U116 );
nand NAND2_3960 ( U6308 , U2371 , R2099_U77 );
nand NAND2_3961 ( U6309 , EBX_REG_18_ , U3413 );
nand NAND2_3962 ( U6310 , U2383 , R2358_U114 );
nand NAND2_3963 ( U6311 , U2371 , R2099_U76 );
nand NAND2_3964 ( U6312 , EBX_REG_19_ , U3413 );
nand NAND2_3965 ( U6313 , U2383 , R2358_U110 );
nand NAND2_3966 ( U6314 , U2371 , R2099_U75 );
nand NAND2_3967 ( U6315 , EBX_REG_20_ , U3413 );
nand NAND2_3968 ( U6316 , U2383 , R2358_U18 );
nand NAND2_3969 ( U6317 , U2371 , R2099_U74 );
nand NAND2_3970 ( U6318 , EBX_REG_21_ , U3413 );
nand NAND2_3971 ( U6319 , U2383 , R2358_U109 );
nand NAND2_3972 ( U6320 , U2371 , R2099_U73 );
nand NAND2_3973 ( U6321 , EBX_REG_22_ , U3413 );
nand NAND2_3974 ( U6322 , U2383 , R2358_U107 );
nand NAND2_3975 ( U6323 , U2371 , R2099_U72 );
nand NAND2_3976 ( U6324 , EBX_REG_23_ , U3413 );
nand NAND2_3977 ( U6325 , U2383 , R2358_U105 );
nand NAND2_3978 ( U6326 , U2371 , R2099_U71 );
nand NAND2_3979 ( U6327 , EBX_REG_24_ , U3413 );
nand NAND2_3980 ( U6328 , U2383 , R2358_U103 );
nand NAND2_3981 ( U6329 , U2371 , R2099_U70 );
nand NAND2_3982 ( U6330 , EBX_REG_25_ , U3413 );
nand NAND2_3983 ( U6331 , U2383 , R2358_U101 );
nand NAND2_3984 ( U6332 , U2371 , R2099_U69 );
nand NAND2_3985 ( U6333 , EBX_REG_26_ , U3413 );
nand NAND2_3986 ( U6334 , U2383 , R2358_U99 );
nand NAND2_3987 ( U6335 , U2371 , R2099_U68 );
nand NAND2_3988 ( U6336 , EBX_REG_27_ , U3413 );
nand NAND2_3989 ( U6337 , U2383 , R2358_U97 );
nand NAND2_3990 ( U6338 , U2371 , R2099_U67 );
nand NAND2_3991 ( U6339 , EBX_REG_28_ , U3413 );
nand NAND2_3992 ( U6340 , U2383 , R2358_U95 );
nand NAND2_3993 ( U6341 , U2371 , R2099_U66 );
nand NAND2_3994 ( U6342 , EBX_REG_29_ , U3413 );
nand NAND2_3995 ( U6343 , U2383 , R2358_U93 );
nand NAND2_3996 ( U6344 , U2371 , R2099_U65 );
nand NAND2_3997 ( U6345 , EBX_REG_30_ , U3413 );
nand NAND2_3998 ( U6346 , U2371 , R2099_U64 );
nand NAND2_3999 ( U6347 , EBX_REG_31_ , U3413 );
nand NAND2_4000 ( U6348 , U4192 , GTE_485_U6 );
nand NAND2_4001 ( U6349 , U4190 , R2167_U17 );
nand NAND2_4002 ( U6350 , U4191 , U3250 );
not NOT1_4003 ( U6351 , U3418 );
nand NAND2_4004 ( U6352 , U4237 , STATE2_REG_2_ );
nand NAND2_4005 ( U6353 , R2337_U58 , STATE2_REG_1_ );
nand NAND2_4006 ( U6354 , U6353 , U6352 );
or OR2_4007 ( U6355 , STATEBS16_REG , READY_N );
nand NAND2_4008 ( U6356 , U2604 , R2099_U86 );
nand NAND2_4009 ( U6357 , REIP_REG_0_ , U7473 );
nand NAND2_4010 ( U6358 , EBX_REG_0_ , U7472 );
nand NAND2_4011 ( U6359 , U2429 , R2358_U82 );
nand NAND2_4012 ( U6360 , U2426 , R2182_U34 );
nand NAND2_4013 ( U6361 , U2373 , PHYADDRPOINTER_REG_0_ );
nand NAND2_4014 ( U6362 , U2366 , PHYADDRPOINTER_REG_0_ );
nand NAND2_4015 ( U6363 , U6351 , REIP_REG_0_ );
nand NAND2_4016 ( U6364 , U2604 , R2099_U87 );
nand NAND2_4017 ( U6365 , R2096_U4 , U7473 );
nand NAND2_4018 ( U6366 , EBX_REG_1_ , U7472 );
nand NAND2_4019 ( U6367 , U2429 , R2358_U112 );
nand NAND2_4020 ( U6368 , U2426 , R2182_U33 );
nand NAND2_4021 ( U6369 , U2373 , PHYADDRPOINTER_REG_1_ );
nand NAND2_4022 ( U6370 , U2366 , R2337_U5 );
nand NAND2_4023 ( U6371 , U6351 , REIP_REG_1_ );
nand NAND2_4024 ( U6372 , U2604 , R2099_U138 );
nand NAND2_4025 ( U6373 , R2096_U71 , U7473 );
nand NAND2_4026 ( U6374 , EBX_REG_2_ , U7472 );
nand NAND2_4027 ( U6375 , U2429 , R2358_U19 );
nand NAND2_4028 ( U6376 , U2426 , R2182_U42 );
nand NAND2_4029 ( U6377 , U2373 , PHYADDRPOINTER_REG_2_ );
nand NAND2_4030 ( U6378 , U2366 , R2337_U60 );
nand NAND2_4031 ( U6379 , U6351 , REIP_REG_2_ );
nand NAND2_4032 ( U6380 , U2604 , R2099_U42 );
nand NAND2_4033 ( U6381 , R2096_U68 , U7473 );
nand NAND2_4034 ( U6382 , EBX_REG_3_ , U7472 );
nand NAND2_4035 ( U6383 , U2429 , R2358_U20 );
nand NAND2_4036 ( U6384 , U2426 , R2182_U25 );
nand NAND2_4037 ( U6385 , U2373 , PHYADDRPOINTER_REG_3_ );
nand NAND2_4038 ( U6386 , U2366 , R2337_U57 );
nand NAND2_4039 ( U6387 , U6351 , REIP_REG_3_ );
nand NAND2_4040 ( U6388 , U2604 , R2099_U41 );
nand NAND2_4041 ( U6389 , R2096_U67 , U7473 );
nand NAND2_4042 ( U6390 , EBX_REG_4_ , U7472 );
nand NAND2_4043 ( U6391 , U2429 , R2358_U90 );
nand NAND2_4044 ( U6392 , U2426 , R2182_U24 );
nand NAND2_4045 ( U6393 , U2373 , PHYADDRPOINTER_REG_4_ );
nand NAND2_4046 ( U6394 , U2366 , R2337_U56 );
nand NAND2_4047 ( U6395 , U6351 , REIP_REG_4_ );
nand NAND2_4048 ( U6396 , U2604 , R2099_U40 );
nand NAND2_4049 ( U6397 , R2096_U66 , U7473 );
nand NAND2_4050 ( U6398 , EBX_REG_5_ , U7472 );
nand NAND2_4051 ( U6399 , U2429 , R2358_U88 );
nand NAND2_4052 ( U6400 , R2182_U5 , U2426 );
nand NAND2_4053 ( U6401 , U2373 , PHYADDRPOINTER_REG_5_ );
nand NAND2_4054 ( U6402 , U2366 , R2337_U55 );
nand NAND2_4055 ( U6403 , U6351 , REIP_REG_5_ );
nand NAND2_4056 ( U6404 , U2604 , R2099_U39 );
nand NAND2_4057 ( U6405 , R2096_U65 , U7473 );
nand NAND2_4058 ( U6406 , EBX_REG_6_ , U7472 );
nand NAND2_4059 ( U6407 , U2373 , PHYADDRPOINTER_REG_6_ );
nand NAND2_4060 ( U6408 , U2367 , R2358_U86 );
nand NAND2_4061 ( U6409 , U2366 , R2337_U54 );
nand NAND2_4062 ( U6410 , U6351 , REIP_REG_6_ );
nand NAND2_4063 ( U6411 , U2604 , R2099_U38 );
nand NAND2_4064 ( U6412 , R2096_U64 , U7473 );
nand NAND2_4065 ( U6413 , EBX_REG_7_ , U7472 );
nand NAND2_4066 ( U6414 , U2373 , PHYADDRPOINTER_REG_7_ );
nand NAND2_4067 ( U6415 , U2367 , R2358_U21 );
nand NAND2_4068 ( U6416 , U2366 , R2337_U53 );
nand NAND2_4069 ( U6417 , U6351 , REIP_REG_7_ );
nand NAND2_4070 ( U6418 , U2604 , R2099_U37 );
nand NAND2_4071 ( U6419 , R2096_U63 , U7473 );
nand NAND2_4072 ( U6420 , EBX_REG_8_ , U7472 );
nand NAND2_4073 ( U6421 , U2373 , PHYADDRPOINTER_REG_8_ );
nand NAND2_4074 ( U6422 , U2367 , R2358_U85 );
nand NAND2_4075 ( U6423 , U2366 , R2337_U52 );
nand NAND2_4076 ( U6424 , U6351 , REIP_REG_8_ );
nand NAND2_4077 ( U6425 , U2604 , R2099_U36 );
nand NAND2_4078 ( U6426 , R2096_U62 , U7473 );
nand NAND2_4079 ( U6427 , EBX_REG_9_ , U7472 );
nand NAND2_4080 ( U6428 , U2373 , PHYADDRPOINTER_REG_9_ );
nand NAND2_4081 ( U6429 , U2367 , R2358_U83 );
nand NAND2_4082 ( U6430 , U2366 , R2337_U51 );
nand NAND2_4083 ( U6431 , U6351 , REIP_REG_9_ );
nand NAND2_4084 ( U6432 , U2604 , R2099_U85 );
nand NAND2_4085 ( U6433 , R2096_U91 , U7473 );
nand NAND2_4086 ( U6434 , EBX_REG_10_ , U7472 );
nand NAND2_4087 ( U6435 , U2373 , PHYADDRPOINTER_REG_10_ );
nand NAND2_4088 ( U6436 , U2367 , R2358_U14 );
nand NAND2_4089 ( U6437 , U2366 , R2337_U80 );
nand NAND2_4090 ( U6438 , U6351 , REIP_REG_10_ );
nand NAND2_4091 ( U6439 , U2604 , R2099_U84 );
nand NAND2_4092 ( U6440 , R2096_U90 , U7473 );
nand NAND2_4093 ( U6441 , EBX_REG_11_ , U7472 );
nand NAND2_4094 ( U6442 , U2373 , PHYADDRPOINTER_REG_11_ );
nand NAND2_4095 ( U6443 , U2367 , R2358_U15 );
nand NAND2_4096 ( U6444 , U2366 , R2337_U79 );
nand NAND2_4097 ( U6445 , U6351 , REIP_REG_11_ );
nand NAND2_4098 ( U6446 , U2604 , R2099_U83 );
nand NAND2_4099 ( U6447 , R2096_U89 , U7473 );
nand NAND2_4100 ( U6448 , EBX_REG_12_ , U7472 );
nand NAND2_4101 ( U6449 , U2373 , PHYADDRPOINTER_REG_12_ );
nand NAND2_4102 ( U6450 , U2367 , R2358_U122 );
nand NAND2_4103 ( U6451 , U2366 , R2337_U78 );
nand NAND2_4104 ( U6452 , U6351 , REIP_REG_12_ );
nand NAND2_4105 ( U6453 , U2604 , R2099_U82 );
nand NAND2_4106 ( U6454 , R2096_U88 , U7473 );
nand NAND2_4107 ( U6455 , EBX_REG_13_ , U7472 );
nand NAND2_4108 ( U6456 , U2373 , PHYADDRPOINTER_REG_13_ );
nand NAND2_4109 ( U6457 , U2367 , R2358_U120 );
nand NAND2_4110 ( U6458 , U2366 , R2337_U77 );
nand NAND2_4111 ( U6459 , U6351 , REIP_REG_13_ );
nand NAND2_4112 ( U6460 , U2604 , R2099_U81 );
nand NAND2_4113 ( U6461 , R2096_U87 , U7473 );
nand NAND2_4114 ( U6462 , EBX_REG_14_ , U7472 );
nand NAND2_4115 ( U6463 , U2373 , PHYADDRPOINTER_REG_14_ );
nand NAND2_4116 ( U6464 , U2367 , R2358_U119 );
nand NAND2_4117 ( U6465 , U2366 , R2337_U76 );
nand NAND2_4118 ( U6466 , U6351 , REIP_REG_14_ );
nand NAND2_4119 ( U6467 , U2604 , R2099_U80 );
nand NAND2_4120 ( U6468 , R2096_U86 , U7473 );
nand NAND2_4121 ( U6469 , EBX_REG_15_ , U7472 );
nand NAND2_4122 ( U6470 , U2373 , PHYADDRPOINTER_REG_15_ );
nand NAND2_4123 ( U6471 , U2367 , R2358_U16 );
nand NAND2_4124 ( U6472 , U2366 , R2337_U75 );
nand NAND2_4125 ( U6473 , U6351 , REIP_REG_15_ );
nand NAND2_4126 ( U6474 , U2604 , R2099_U79 );
nand NAND2_4127 ( U6475 , R2096_U85 , U7473 );
nand NAND2_4128 ( U6476 , EBX_REG_16_ , U7472 );
nand NAND2_4129 ( U6477 , U2373 , PHYADDRPOINTER_REG_16_ );
nand NAND2_4130 ( U6478 , U2367 , R2358_U17 );
nand NAND2_4131 ( U6479 , U2366 , R2337_U74 );
nand NAND2_4132 ( U6480 , U6351 , REIP_REG_16_ );
nand NAND2_4133 ( U6481 , U2604 , R2099_U78 );
nand NAND2_4134 ( U6482 , R2096_U84 , U7473 );
nand NAND2_4135 ( U6483 , EBX_REG_17_ , U7472 );
nand NAND2_4136 ( U6484 , U2373 , PHYADDRPOINTER_REG_17_ );
nand NAND2_4137 ( U6485 , U2367 , R2358_U118 );
nand NAND2_4138 ( U6486 , U2366 , R2337_U73 );
nand NAND2_4139 ( U6487 , U6351 , REIP_REG_17_ );
nand NAND2_4140 ( U6488 , U2604 , R2099_U77 );
nand NAND2_4141 ( U6489 , R2096_U83 , U7473 );
nand NAND2_4142 ( U6490 , EBX_REG_18_ , U7472 );
nand NAND2_4143 ( U6491 , U2373 , PHYADDRPOINTER_REG_18_ );
nand NAND2_4144 ( U6492 , U2367 , R2358_U116 );
nand NAND2_4145 ( U6493 , U2366 , R2337_U72 );
nand NAND2_4146 ( U6494 , U6351 , REIP_REG_18_ );
nand NAND2_4147 ( U6495 , U2604 , R2099_U76 );
nand NAND2_4148 ( U6496 , R2096_U82 , U7473 );
nand NAND2_4149 ( U6497 , EBX_REG_19_ , U7472 );
nand NAND2_4150 ( U6498 , U2373 , PHYADDRPOINTER_REG_19_ );
nand NAND2_4151 ( U6499 , U2367 , R2358_U114 );
nand NAND2_4152 ( U6500 , U2366 , R2337_U71 );
nand NAND2_4153 ( U6501 , U6351 , REIP_REG_19_ );
nand NAND2_4154 ( U6502 , U2604 , R2099_U75 );
nand NAND2_4155 ( U6503 , R2096_U81 , U7473 );
nand NAND2_4156 ( U6504 , EBX_REG_20_ , U7472 );
nand NAND2_4157 ( U6505 , U2373 , PHYADDRPOINTER_REG_20_ );
nand NAND2_4158 ( U6506 , U2367 , R2358_U110 );
nand NAND2_4159 ( U6507 , U2366 , R2337_U70 );
nand NAND2_4160 ( U6508 , U6351 , REIP_REG_20_ );
nand NAND2_4161 ( U6509 , U2604 , R2099_U74 );
nand NAND2_4162 ( U6510 , R2096_U80 , U7473 );
nand NAND2_4163 ( U6511 , EBX_REG_21_ , U7472 );
nand NAND2_4164 ( U6512 , U2373 , PHYADDRPOINTER_REG_21_ );
nand NAND2_4165 ( U6513 , U2367 , R2358_U18 );
nand NAND2_4166 ( U6514 , U2366 , R2337_U69 );
nand NAND2_4167 ( U6515 , U6351 , REIP_REG_21_ );
nand NAND2_4168 ( U6516 , U2604 , R2099_U73 );
nand NAND2_4169 ( U6517 , R2096_U79 , U7473 );
nand NAND2_4170 ( U6518 , EBX_REG_22_ , U7472 );
nand NAND2_4171 ( U6519 , U2373 , PHYADDRPOINTER_REG_22_ );
nand NAND2_4172 ( U6520 , U2367 , R2358_U109 );
nand NAND2_4173 ( U6521 , U2366 , R2337_U68 );
nand NAND2_4174 ( U6522 , U6351 , REIP_REG_22_ );
nand NAND2_4175 ( U6523 , U2604 , R2099_U72 );
nand NAND2_4176 ( U6524 , R2096_U78 , U7473 );
nand NAND2_4177 ( U6525 , EBX_REG_23_ , U7472 );
nand NAND2_4178 ( U6526 , U2373 , PHYADDRPOINTER_REG_23_ );
nand NAND2_4179 ( U6527 , U2367 , R2358_U107 );
nand NAND2_4180 ( U6528 , U2366 , R2337_U67 );
nand NAND2_4181 ( U6529 , U6351 , REIP_REG_23_ );
nand NAND2_4182 ( U6530 , U2604 , R2099_U71 );
nand NAND2_4183 ( U6531 , R2096_U77 , U7473 );
nand NAND2_4184 ( U6532 , EBX_REG_24_ , U7472 );
nand NAND2_4185 ( U6533 , U2373 , PHYADDRPOINTER_REG_24_ );
nand NAND2_4186 ( U6534 , U2367 , R2358_U105 );
nand NAND2_4187 ( U6535 , U2366 , R2337_U66 );
nand NAND2_4188 ( U6536 , U6351 , REIP_REG_24_ );
nand NAND2_4189 ( U6537 , U2604 , R2099_U70 );
nand NAND2_4190 ( U6538 , R2096_U76 , U7473 );
nand NAND2_4191 ( U6539 , EBX_REG_25_ , U7472 );
nand NAND2_4192 ( U6540 , U2373 , PHYADDRPOINTER_REG_25_ );
nand NAND2_4193 ( U6541 , U2367 , R2358_U103 );
nand NAND2_4194 ( U6542 , U2366 , R2337_U65 );
nand NAND2_4195 ( U6543 , U6351 , REIP_REG_25_ );
nand NAND2_4196 ( U6544 , U2604 , R2099_U69 );
nand NAND2_4197 ( U6545 , R2096_U75 , U7473 );
nand NAND2_4198 ( U6546 , EBX_REG_26_ , U7472 );
nand NAND2_4199 ( U6547 , U2373 , PHYADDRPOINTER_REG_26_ );
nand NAND2_4200 ( U6548 , U2367 , R2358_U101 );
nand NAND2_4201 ( U6549 , U2366 , R2337_U64 );
nand NAND2_4202 ( U6550 , U6351 , REIP_REG_26_ );
nand NAND2_4203 ( U6551 , U2604 , R2099_U68 );
nand NAND2_4204 ( U6552 , R2096_U74 , U7473 );
nand NAND2_4205 ( U6553 , EBX_REG_27_ , U7472 );
nand NAND2_4206 ( U6554 , U2373 , PHYADDRPOINTER_REG_27_ );
nand NAND2_4207 ( U6555 , U2367 , R2358_U99 );
nand NAND2_4208 ( U6556 , U2366 , R2337_U63 );
nand NAND2_4209 ( U6557 , U6351 , REIP_REG_27_ );
nand NAND2_4210 ( U6558 , U2604 , R2099_U67 );
nand NAND2_4211 ( U6559 , R2096_U73 , U7473 );
nand NAND2_4212 ( U6560 , EBX_REG_28_ , U7472 );
nand NAND2_4213 ( U6561 , U2373 , PHYADDRPOINTER_REG_28_ );
nand NAND2_4214 ( U6562 , U2367 , R2358_U97 );
nand NAND2_4215 ( U6563 , U2366 , R2337_U62 );
nand NAND2_4216 ( U6564 , U6351 , REIP_REG_28_ );
nand NAND2_4217 ( U6565 , U2604 , R2099_U66 );
nand NAND2_4218 ( U6566 , R2096_U72 , U7473 );
nand NAND2_4219 ( U6567 , EBX_REG_29_ , U7472 );
nand NAND2_4220 ( U6568 , U2373 , PHYADDRPOINTER_REG_29_ );
nand NAND2_4221 ( U6569 , U2367 , R2358_U95 );
nand NAND2_4222 ( U6570 , U2366 , R2337_U61 );
nand NAND2_4223 ( U6571 , U6351 , REIP_REG_29_ );
nand NAND2_4224 ( U6572 , U2604 , R2099_U65 );
nand NAND2_4225 ( U6573 , R2096_U70 , U7473 );
nand NAND2_4226 ( U6574 , EBX_REG_30_ , U7472 );
nand NAND2_4227 ( U6575 , U2373 , PHYADDRPOINTER_REG_30_ );
nand NAND2_4228 ( U6576 , U2367 , R2358_U93 );
nand NAND2_4229 ( U6577 , U2366 , R2337_U59 );
nand NAND2_4230 ( U6578 , U6351 , REIP_REG_30_ );
nand NAND2_4231 ( U6579 , U2604 , R2099_U64 );
nand NAND2_4232 ( U6580 , R2096_U69 , U7473 );
nand NAND2_4233 ( U6581 , EBX_REG_31_ , U7472 );
nand NAND2_4234 ( U6582 , U2373 , PHYADDRPOINTER_REG_31_ );
nand NAND2_4235 ( U6583 , U2367 , R2358_U91 );
nand NAND2_4236 ( U6584 , U2366 , R2337_U58 );
nand NAND2_4237 ( U6585 , U6351 , REIP_REG_31_ );
nand NAND2_4238 ( U6586 , DATAWIDTH_REG_1_ , DATAWIDTH_REG_0_ );
or OR2_4239 ( U6587 , REIP_REG_1_ , REIP_REG_0_ );
not NOT1_4240 ( U6588 , U4165 );
nand NAND2_4241 ( U6589 , FLUSH_REG , U4165 );
nand NAND2_4242 ( U6590 , U3954 , U2428 );
not NOT1_4243 ( U6591 , U4168 );
nand NAND2_4244 ( U6592 , STATEBS16_REG , U4485 );
nand NAND2_4245 ( U6593 , U4196 , U6592 );
nand NAND2_4246 ( U6594 , U3952 , U6593 );
nand NAND2_4247 ( U6595 , STATE2_REG_0_ , U6594 );
nand NAND2_4248 ( U6596 , U4181 , U3259 );
nand NAND2_4249 ( U6597 , U3953 , U6595 );
nand NAND2_4250 ( U6598 , U2368 , U2473 );
nand NAND2_4251 ( U6599 , CODEFETCH_REG , U6598 );
nand NAND2_4252 ( U6600 , U4243 , STATE2_REG_0_ );
nand NAND2_4253 ( U6601 , ADS_N_REG , STATE_REG_0_ );
not NOT1_4254 ( U6602 , U4169 );
nand NAND2_4255 ( U6603 , U3956 , U3278 );
nand NAND3_4256 ( U6604 , U4487 , U3957 , U3393 );
nand NAND2_4257 ( U6605 , MEMORYFETCH_REG , U6604 );
nand NAND2_4258 ( U6606 , U2544 , INSTQUEUE_REG_15__7_ );
nand NAND2_4259 ( U6607 , U2543 , INSTQUEUE_REG_14__7_ );
nand NAND2_4260 ( U6608 , U2542 , INSTQUEUE_REG_13__7_ );
nand NAND2_4261 ( U6609 , U2541 , INSTQUEUE_REG_12__7_ );
nand NAND2_4262 ( U6610 , U2539 , INSTQUEUE_REG_11__7_ );
nand NAND2_4263 ( U6611 , U2538 , INSTQUEUE_REG_10__7_ );
nand NAND2_4264 ( U6612 , U2537 , INSTQUEUE_REG_9__7_ );
nand NAND2_4265 ( U6613 , U2536 , INSTQUEUE_REG_8__7_ );
nand NAND2_4266 ( U6614 , U2534 , INSTQUEUE_REG_7__7_ );
nand NAND2_4267 ( U6615 , U2533 , INSTQUEUE_REG_6__7_ );
nand NAND2_4268 ( U6616 , U2532 , INSTQUEUE_REG_5__7_ );
nand NAND2_4269 ( U6617 , U2531 , INSTQUEUE_REG_4__7_ );
nand NAND2_4270 ( U6618 , U2529 , INSTQUEUE_REG_3__7_ );
nand NAND2_4271 ( U6619 , U2527 , INSTQUEUE_REG_2__7_ );
nand NAND2_4272 ( U6620 , U2525 , INSTQUEUE_REG_1__7_ );
nand NAND2_4273 ( U6621 , U2523 , INSTQUEUE_REG_0__7_ );
nand NAND2_4274 ( U6622 , U2544 , INSTQUEUE_REG_15__6_ );
nand NAND2_4275 ( U6623 , U2543 , INSTQUEUE_REG_14__6_ );
nand NAND2_4276 ( U6624 , U2542 , INSTQUEUE_REG_13__6_ );
nand NAND2_4277 ( U6625 , U2541 , INSTQUEUE_REG_12__6_ );
nand NAND2_4278 ( U6626 , U2539 , INSTQUEUE_REG_11__6_ );
nand NAND2_4279 ( U6627 , U2538 , INSTQUEUE_REG_10__6_ );
nand NAND2_4280 ( U6628 , U2537 , INSTQUEUE_REG_9__6_ );
nand NAND2_4281 ( U6629 , U2536 , INSTQUEUE_REG_8__6_ );
nand NAND2_4282 ( U6630 , U2534 , INSTQUEUE_REG_7__6_ );
nand NAND2_4283 ( U6631 , U2533 , INSTQUEUE_REG_6__6_ );
nand NAND2_4284 ( U6632 , U2532 , INSTQUEUE_REG_5__6_ );
nand NAND2_4285 ( U6633 , U2531 , INSTQUEUE_REG_4__6_ );
nand NAND2_4286 ( U6634 , U2529 , INSTQUEUE_REG_3__6_ );
nand NAND2_4287 ( U6635 , U2527 , INSTQUEUE_REG_2__6_ );
nand NAND2_4288 ( U6636 , U2525 , INSTQUEUE_REG_1__6_ );
nand NAND2_4289 ( U6637 , U2523 , INSTQUEUE_REG_0__6_ );
nand NAND2_4290 ( U6638 , U2544 , INSTQUEUE_REG_15__5_ );
nand NAND2_4291 ( U6639 , U2543 , INSTQUEUE_REG_14__5_ );
nand NAND2_4292 ( U6640 , U2542 , INSTQUEUE_REG_13__5_ );
nand NAND2_4293 ( U6641 , U2541 , INSTQUEUE_REG_12__5_ );
nand NAND2_4294 ( U6642 , U2539 , INSTQUEUE_REG_11__5_ );
nand NAND2_4295 ( U6643 , U2538 , INSTQUEUE_REG_10__5_ );
nand NAND2_4296 ( U6644 , U2537 , INSTQUEUE_REG_9__5_ );
nand NAND2_4297 ( U6645 , U2536 , INSTQUEUE_REG_8__5_ );
nand NAND2_4298 ( U6646 , U2534 , INSTQUEUE_REG_7__5_ );
nand NAND2_4299 ( U6647 , U2533 , INSTQUEUE_REG_6__5_ );
nand NAND2_4300 ( U6648 , U2532 , INSTQUEUE_REG_5__5_ );
nand NAND2_4301 ( U6649 , U2531 , INSTQUEUE_REG_4__5_ );
nand NAND2_4302 ( U6650 , U2529 , INSTQUEUE_REG_3__5_ );
nand NAND2_4303 ( U6651 , U2527 , INSTQUEUE_REG_2__5_ );
nand NAND2_4304 ( U6652 , U2525 , INSTQUEUE_REG_1__5_ );
nand NAND2_4305 ( U6653 , U2523 , INSTQUEUE_REG_0__5_ );
nand NAND2_4306 ( U6654 , U2544 , INSTQUEUE_REG_15__4_ );
nand NAND2_4307 ( U6655 , U2543 , INSTQUEUE_REG_14__4_ );
nand NAND2_4308 ( U6656 , U2542 , INSTQUEUE_REG_13__4_ );
nand NAND2_4309 ( U6657 , U2541 , INSTQUEUE_REG_12__4_ );
nand NAND2_4310 ( U6658 , U2539 , INSTQUEUE_REG_11__4_ );
nand NAND2_4311 ( U6659 , U2538 , INSTQUEUE_REG_10__4_ );
nand NAND2_4312 ( U6660 , U2537 , INSTQUEUE_REG_9__4_ );
nand NAND2_4313 ( U6661 , U2536 , INSTQUEUE_REG_8__4_ );
nand NAND2_4314 ( U6662 , U2534 , INSTQUEUE_REG_7__4_ );
nand NAND2_4315 ( U6663 , U2533 , INSTQUEUE_REG_6__4_ );
nand NAND2_4316 ( U6664 , U2532 , INSTQUEUE_REG_5__4_ );
nand NAND2_4317 ( U6665 , U2531 , INSTQUEUE_REG_4__4_ );
nand NAND2_4318 ( U6666 , U2529 , INSTQUEUE_REG_3__4_ );
nand NAND2_4319 ( U6667 , U2527 , INSTQUEUE_REG_2__4_ );
nand NAND2_4320 ( U6668 , U2525 , INSTQUEUE_REG_1__4_ );
nand NAND2_4321 ( U6669 , U2544 , INSTQUEUE_REG_15__3_ );
nand NAND2_4322 ( U6670 , U2543 , INSTQUEUE_REG_14__3_ );
nand NAND2_4323 ( U6671 , U2542 , INSTQUEUE_REG_13__3_ );
nand NAND2_4324 ( U6672 , U2541 , INSTQUEUE_REG_12__3_ );
nand NAND2_4325 ( U6673 , U2539 , INSTQUEUE_REG_11__3_ );
nand NAND2_4326 ( U6674 , U2538 , INSTQUEUE_REG_10__3_ );
nand NAND2_4327 ( U6675 , U2537 , INSTQUEUE_REG_9__3_ );
nand NAND2_4328 ( U6676 , U2536 , INSTQUEUE_REG_8__3_ );
nand NAND2_4329 ( U6677 , U2534 , INSTQUEUE_REG_7__3_ );
nand NAND2_4330 ( U6678 , U2533 , INSTQUEUE_REG_6__3_ );
nand NAND2_4331 ( U6679 , U2532 , INSTQUEUE_REG_5__3_ );
nand NAND2_4332 ( U6680 , U2531 , INSTQUEUE_REG_4__3_ );
nand NAND2_4333 ( U6681 , U2529 , INSTQUEUE_REG_3__3_ );
nand NAND2_4334 ( U6682 , U2527 , INSTQUEUE_REG_2__3_ );
nand NAND2_4335 ( U6683 , U2525 , INSTQUEUE_REG_1__3_ );
nand NAND2_4336 ( U6684 , U2523 , INSTQUEUE_REG_0__3_ );
nand NAND2_4337 ( U6685 , U2544 , INSTQUEUE_REG_15__2_ );
nand NAND2_4338 ( U6686 , U2543 , INSTQUEUE_REG_14__2_ );
nand NAND2_4339 ( U6687 , U2542 , INSTQUEUE_REG_13__2_ );
nand NAND2_4340 ( U6688 , U2541 , INSTQUEUE_REG_12__2_ );
nand NAND2_4341 ( U6689 , U2539 , INSTQUEUE_REG_11__2_ );
nand NAND2_4342 ( U6690 , U2538 , INSTQUEUE_REG_10__2_ );
nand NAND2_4343 ( U6691 , U2537 , INSTQUEUE_REG_9__2_ );
nand NAND2_4344 ( U6692 , U2536 , INSTQUEUE_REG_8__2_ );
nand NAND2_4345 ( U6693 , U2534 , INSTQUEUE_REG_7__2_ );
nand NAND2_4346 ( U6694 , U2533 , INSTQUEUE_REG_6__2_ );
nand NAND2_4347 ( U6695 , U2532 , INSTQUEUE_REG_5__2_ );
nand NAND2_4348 ( U6696 , U2531 , INSTQUEUE_REG_4__2_ );
nand NAND2_4349 ( U6697 , U2529 , INSTQUEUE_REG_3__2_ );
nand NAND2_4350 ( U6698 , U2527 , INSTQUEUE_REG_2__2_ );
nand NAND2_4351 ( U6699 , U2525 , INSTQUEUE_REG_1__2_ );
nand NAND2_4352 ( U6700 , U2523 , INSTQUEUE_REG_0__2_ );
nand NAND2_4353 ( U6701 , U2544 , INSTQUEUE_REG_15__1_ );
nand NAND2_4354 ( U6702 , U2543 , INSTQUEUE_REG_14__1_ );
nand NAND2_4355 ( U6703 , U2542 , INSTQUEUE_REG_13__1_ );
nand NAND2_4356 ( U6704 , U2541 , INSTQUEUE_REG_12__1_ );
nand NAND2_4357 ( U6705 , U2539 , INSTQUEUE_REG_11__1_ );
nand NAND2_4358 ( U6706 , U2538 , INSTQUEUE_REG_10__1_ );
nand NAND2_4359 ( U6707 , U2537 , INSTQUEUE_REG_9__1_ );
nand NAND2_4360 ( U6708 , U2536 , INSTQUEUE_REG_8__1_ );
nand NAND2_4361 ( U6709 , U2534 , INSTQUEUE_REG_7__1_ );
nand NAND2_4362 ( U6710 , U2533 , INSTQUEUE_REG_6__1_ );
nand NAND2_4363 ( U6711 , U2532 , INSTQUEUE_REG_5__1_ );
nand NAND2_4364 ( U6712 , U2531 , INSTQUEUE_REG_4__1_ );
nand NAND2_4365 ( U6713 , U2529 , INSTQUEUE_REG_3__1_ );
nand NAND2_4366 ( U6714 , U2527 , INSTQUEUE_REG_2__1_ );
nand NAND2_4367 ( U6715 , U2525 , INSTQUEUE_REG_1__1_ );
nand NAND2_4368 ( U6716 , U2523 , INSTQUEUE_REG_0__1_ );
nand NAND2_4369 ( U6717 , U2544 , INSTQUEUE_REG_15__0_ );
nand NAND2_4370 ( U6718 , U2543 , INSTQUEUE_REG_14__0_ );
nand NAND2_4371 ( U6719 , U2542 , INSTQUEUE_REG_13__0_ );
nand NAND2_4372 ( U6720 , U2541 , INSTQUEUE_REG_12__0_ );
nand NAND2_4373 ( U6721 , U2539 , INSTQUEUE_REG_11__0_ );
nand NAND2_4374 ( U6722 , U2538 , INSTQUEUE_REG_10__0_ );
nand NAND2_4375 ( U6723 , U2537 , INSTQUEUE_REG_9__0_ );
nand NAND2_4376 ( U6724 , U2536 , INSTQUEUE_REG_8__0_ );
nand NAND2_4377 ( U6725 , U2534 , INSTQUEUE_REG_7__0_ );
nand NAND2_4378 ( U6726 , U2533 , INSTQUEUE_REG_6__0_ );
nand NAND2_4379 ( U6727 , U2532 , INSTQUEUE_REG_5__0_ );
nand NAND2_4380 ( U6728 , U2531 , INSTQUEUE_REG_4__0_ );
nand NAND2_4381 ( U6729 , U2529 , INSTQUEUE_REG_3__0_ );
nand NAND2_4382 ( U6730 , U2527 , INSTQUEUE_REG_2__0_ );
nand NAND2_4383 ( U6731 , U2525 , INSTQUEUE_REG_1__0_ );
nand NAND2_4384 ( U6732 , U2523 , INSTQUEUE_REG_0__0_ );
nand NAND2_4385 ( U6733 , U4448 , STATE2_REG_2_ );
nand NAND2_4386 ( U6734 , U3399 , U6733 );
nand NAND2_4387 ( U6735 , U4176 , EAX_REG_9_ );
nand NAND2_4388 ( U6736 , U4175 , PHYADDRPOINTER_REG_9_ );
nand NAND2_4389 ( U6737 , R2337_U51 , U2352 );
nand NAND2_4390 ( U6738 , U4176 , EAX_REG_8_ );
nand NAND2_4391 ( U6739 , U4175 , PHYADDRPOINTER_REG_8_ );
nand NAND2_4392 ( U6740 , R2337_U52 , U2352 );
nand NAND2_4393 ( U6741 , U4176 , EAX_REG_7_ );
nand NAND2_4394 ( U6742 , U4175 , PHYADDRPOINTER_REG_7_ );
nand NAND2_4395 ( U6743 , R2337_U53 , U2352 );
nand NAND2_4396 ( U6744 , U4176 , EAX_REG_6_ );
nand NAND2_4397 ( U6745 , U4175 , PHYADDRPOINTER_REG_6_ );
nand NAND2_4398 ( U6746 , R2337_U54 , U2352 );
nand NAND2_4399 ( U6747 , R2182_U5 , U6734 );
nand NAND2_4400 ( U6748 , U4176 , EAX_REG_5_ );
nand NAND2_4401 ( U6749 , U4175 , PHYADDRPOINTER_REG_5_ );
nand NAND2_4402 ( U6750 , R2337_U55 , U2352 );
nand NAND2_4403 ( U6751 , R2182_U24 , U6734 );
nand NAND2_4404 ( U6752 , U4176 , EAX_REG_4_ );
nand NAND2_4405 ( U6753 , U4175 , PHYADDRPOINTER_REG_4_ );
nand NAND2_4406 ( U6754 , R2337_U56 , U2352 );
nand NAND2_4407 ( U6755 , U2353 , INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_4408 ( U6756 , U4176 , EAX_REG_31_ );
nand NAND2_4409 ( U6757 , U4175 , PHYADDRPOINTER_REG_31_ );
nand NAND2_4410 ( U6758 , R2337_U58 , U2352 );
nand NAND2_4411 ( U6759 , R2182_U26 , U6734 );
nand NAND2_4412 ( U6760 , U4176 , EAX_REG_30_ );
nand NAND2_4413 ( U6761 , U4175 , PHYADDRPOINTER_REG_30_ );
nand NAND2_4414 ( U6762 , R2337_U59 , U2352 );
nand NAND2_4415 ( U6763 , R2182_U25 , U6734 );
nand NAND2_4416 ( U6764 , U4176 , EAX_REG_3_ );
nand NAND2_4417 ( U6765 , U4175 , PHYADDRPOINTER_REG_3_ );
nand NAND2_4418 ( U6766 , R2337_U57 , U2352 );
nand NAND2_4419 ( U6767 , U2353 , INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_4420 ( U6768 , R2182_U27 , U6734 );
nand NAND2_4421 ( U6769 , U4176 , EAX_REG_29_ );
nand NAND2_4422 ( U6770 , U4175 , PHYADDRPOINTER_REG_29_ );
nand NAND2_4423 ( U6771 , R2337_U61 , U2352 );
nand NAND2_4424 ( U6772 , R2182_U28 , U6734 );
nand NAND2_4425 ( U6773 , U4176 , EAX_REG_28_ );
nand NAND2_4426 ( U6774 , U4175 , PHYADDRPOINTER_REG_28_ );
nand NAND2_4427 ( U6775 , R2337_U62 , U2352 );
nand NAND2_4428 ( U6776 , R2182_U29 , U6734 );
nand NAND2_4429 ( U6777 , U4176 , EAX_REG_27_ );
nand NAND2_4430 ( U6778 , U4175 , PHYADDRPOINTER_REG_27_ );
nand NAND2_4431 ( U6779 , R2337_U63 , U2352 );
nand NAND2_4432 ( U6780 , R2182_U30 , U6734 );
nand NAND2_4433 ( U6781 , U4176 , EAX_REG_26_ );
nand NAND2_4434 ( U6782 , U4175 , PHYADDRPOINTER_REG_26_ );
nand NAND2_4435 ( U6783 , R2337_U64 , U2352 );
nand NAND2_4436 ( U6784 , R2182_U31 , U6734 );
nand NAND2_4437 ( U6785 , U4176 , EAX_REG_25_ );
nand NAND2_4438 ( U6786 , U4175 , PHYADDRPOINTER_REG_25_ );
nand NAND2_4439 ( U6787 , R2337_U65 , U2352 );
nand NAND2_4440 ( U6788 , R2182_U32 , U6734 );
nand NAND2_4441 ( U6789 , U4176 , EAX_REG_24_ );
nand NAND2_4442 ( U6790 , U4175 , PHYADDRPOINTER_REG_24_ );
nand NAND2_4443 ( U6791 , R2337_U66 , U2352 );
nand NAND2_4444 ( U6792 , R2182_U6 , U6734 );
nand NAND2_4445 ( U6793 , U4176 , EAX_REG_23_ );
nand NAND2_4446 ( U6794 , U4175 , PHYADDRPOINTER_REG_23_ );
nand NAND2_4447 ( U6795 , R2337_U67 , U2352 );
nand NAND2_4448 ( U6796 , U2724 , U6734 );
nand NAND2_4449 ( U6797 , U4176 , EAX_REG_22_ );
nand NAND2_4450 ( U6798 , U4175 , PHYADDRPOINTER_REG_22_ );
nand NAND2_4451 ( U6799 , R2337_U68 , U2352 );
nand NAND2_4452 ( U6800 , U2725 , U6734 );
nand NAND2_4453 ( U6801 , U4176 , EAX_REG_21_ );
nand NAND2_4454 ( U6802 , U4175 , PHYADDRPOINTER_REG_21_ );
nand NAND2_4455 ( U6803 , R2337_U69 , U2352 );
nand NAND2_4456 ( U6804 , U2726 , U6734 );
nand NAND2_4457 ( U6805 , U4176 , EAX_REG_20_ );
nand NAND2_4458 ( U6806 , U4175 , PHYADDRPOINTER_REG_20_ );
nand NAND2_4459 ( U6807 , R2337_U70 , U2352 );
nand NAND2_4460 ( U6808 , R2182_U42 , U6734 );
nand NAND2_4461 ( U6809 , U4176 , EAX_REG_2_ );
nand NAND2_4462 ( U6810 , U4175 , PHYADDRPOINTER_REG_2_ );
nand NAND2_4463 ( U6811 , R2337_U60 , U2352 );
nand NAND2_4464 ( U6812 , U2353 , INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_4465 ( U6813 , U2727 , U6734 );
nand NAND2_4466 ( U6814 , U4176 , EAX_REG_19_ );
nand NAND2_4467 ( U6815 , U4175 , PHYADDRPOINTER_REG_19_ );
nand NAND2_4468 ( U6816 , R2337_U71 , U2352 );
nand NAND2_4469 ( U6817 , U2728 , U6734 );
nand NAND2_4470 ( U6818 , U4176 , EAX_REG_18_ );
nand NAND2_4471 ( U6819 , U4175 , PHYADDRPOINTER_REG_18_ );
nand NAND2_4472 ( U6820 , R2337_U72 , U2352 );
nand NAND2_4473 ( U6821 , U2729 , U6734 );
nand NAND2_4474 ( U6822 , U4176 , EAX_REG_17_ );
nand NAND2_4475 ( U6823 , U4175 , PHYADDRPOINTER_REG_17_ );
nand NAND2_4476 ( U6824 , R2337_U73 , U2352 );
nand NAND2_4477 ( U6825 , U2730 , U6734 );
nand NAND2_4478 ( U6826 , U4176 , EAX_REG_16_ );
nand NAND2_4479 ( U6827 , U4175 , PHYADDRPOINTER_REG_16_ );
nand NAND2_4480 ( U6828 , R2337_U74 , U2352 );
nand NAND2_4481 ( U6829 , U4176 , EAX_REG_15_ );
nand NAND2_4482 ( U6830 , U4175 , PHYADDRPOINTER_REG_15_ );
nand NAND2_4483 ( U6831 , R2337_U75 , U2352 );
nand NAND2_4484 ( U6832 , U4176 , EAX_REG_14_ );
nand NAND2_4485 ( U6833 , U4175 , PHYADDRPOINTER_REG_14_ );
nand NAND2_4486 ( U6834 , R2337_U76 , U2352 );
nand NAND2_4487 ( U6835 , U4176 , EAX_REG_13_ );
nand NAND2_4488 ( U6836 , U4175 , PHYADDRPOINTER_REG_13_ );
nand NAND2_4489 ( U6837 , R2337_U77 , U2352 );
nand NAND2_4490 ( U6838 , U4176 , EAX_REG_12_ );
nand NAND2_4491 ( U6839 , U4175 , PHYADDRPOINTER_REG_12_ );
nand NAND2_4492 ( U6840 , R2337_U78 , U2352 );
nand NAND2_4493 ( U6841 , U4176 , EAX_REG_11_ );
nand NAND2_4494 ( U6842 , U4175 , PHYADDRPOINTER_REG_11_ );
nand NAND2_4495 ( U6843 , R2337_U79 , U2352 );
nand NAND2_4496 ( U6844 , U4176 , EAX_REG_10_ );
nand NAND2_4497 ( U6845 , U4175 , PHYADDRPOINTER_REG_10_ );
nand NAND2_4498 ( U6846 , R2337_U80 , U2352 );
nand NAND2_4499 ( U6847 , R2182_U33 , U6734 );
nand NAND2_4500 ( U6848 , U4176 , EAX_REG_1_ );
nand NAND2_4501 ( U6849 , U4175 , PHYADDRPOINTER_REG_1_ );
nand NAND2_4502 ( U6850 , R2337_U5 , U2352 );
nand NAND2_4503 ( U6851 , U2353 , INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_4504 ( U6852 , R2182_U34 , U6734 );
nand NAND2_4505 ( U6853 , U4176 , EAX_REG_0_ );
nand NAND2_4506 ( U6854 , U4175 , PHYADDRPOINTER_REG_0_ );
nand NAND2_4507 ( U6855 , PHYADDRPOINTER_REG_0_ , U2352 );
nand NAND2_4508 ( U6856 , U2353 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_4509 ( U6857 , R2144_U49 , U6734 );
nand NAND3_4510 ( U6858 , U3426 , U4448 , U3296 );
nand NAND2_4511 ( U6859 , U4147 , R2144_U80 );
nand NAND2_4512 ( U6860 , ADD_371_U6 , U4196 );
nand NAND2_4513 ( U6861 , U4147 , R2144_U10 );
nand NAND2_4514 ( U6862 , ADD_371_U17 , U4196 );
nand NAND2_4515 ( U6863 , U4147 , R2144_U9 );
nand NAND2_4516 ( U6864 , ADD_371_U18 , U4196 );
nand NAND2_4517 ( U6865 , U4147 , R2144_U45 );
nand NAND2_4518 ( U6866 , ADD_371_U19 , U4196 );
nand NAND2_4519 ( U6867 , U4147 , R2144_U47 );
nand NAND2_4520 ( U6868 , ADD_371_U20 , U4196 );
nand NAND2_4521 ( U6869 , U4147 , R2144_U8 );
nand NAND2_4522 ( U6870 , ADD_371_U25 , U4196 );
nand NAND2_4523 ( U6871 , U4147 , R2144_U49 );
nand NAND2_4524 ( U6872 , ADD_371_U5 , U4196 );
nand NAND2_4525 ( U6873 , U4482 , U3270 );
nand NAND2_4526 ( U6874 , U4147 , R2144_U50 );
nand NAND2_4527 ( U6875 , ADD_371_U21 , U4196 );
nand NAND2_4528 ( U6876 , U2605 , U3271 );
nand NAND2_4529 ( U6877 , U4147 , R2144_U43 );
nand NAND2_4530 ( U6878 , ADD_371_U4 , U4196 );
nand NAND2_4531 ( U6879 , U4482 , U3270 );
nand NAND2_4532 ( U6880 , U2564 , INSTQUEUE_REG_15__1_ );
nand NAND2_4533 ( U6881 , U2563 , INSTQUEUE_REG_14__1_ );
nand NAND2_4534 ( U6882 , U2562 , INSTQUEUE_REG_13__1_ );
nand NAND2_4535 ( U6883 , U2561 , INSTQUEUE_REG_12__1_ );
nand NAND2_4536 ( U6884 , U2559 , INSTQUEUE_REG_11__1_ );
nand NAND2_4537 ( U6885 , U2558 , INSTQUEUE_REG_10__1_ );
nand NAND2_4538 ( U6886 , U2557 , INSTQUEUE_REG_9__1_ );
nand NAND2_4539 ( U6887 , U2556 , INSTQUEUE_REG_8__1_ );
nand NAND2_4540 ( U6888 , U2554 , INSTQUEUE_REG_7__1_ );
nand NAND2_4541 ( U6889 , U2553 , INSTQUEUE_REG_6__1_ );
nand NAND2_4542 ( U6890 , U2552 , INSTQUEUE_REG_5__1_ );
nand NAND2_4543 ( U6891 , U2551 , INSTQUEUE_REG_4__1_ );
nand NAND2_4544 ( U6892 , U2549 , INSTQUEUE_REG_3__1_ );
nand NAND2_4545 ( U6893 , U2548 , INSTQUEUE_REG_2__1_ );
nand NAND2_4546 ( U6894 , U2547 , INSTQUEUE_REG_1__1_ );
nand NAND2_4547 ( U6895 , U2546 , INSTQUEUE_REG_0__1_ );
nand NAND4_4548 ( U6896 , U4020 , U4019 , U4018 , U4017 );
nand NAND2_4549 ( U6897 , U3392 , U3405 );
nand NAND2_4550 ( U6898 , U2564 , INSTQUEUE_REG_15__0_ );
nand NAND2_4551 ( U6899 , U2563 , INSTQUEUE_REG_14__0_ );
nand NAND2_4552 ( U6900 , U2562 , INSTQUEUE_REG_13__0_ );
nand NAND2_4553 ( U6901 , U2561 , INSTQUEUE_REG_12__0_ );
nand NAND2_4554 ( U6902 , U2559 , INSTQUEUE_REG_11__0_ );
nand NAND2_4555 ( U6903 , U2558 , INSTQUEUE_REG_10__0_ );
nand NAND2_4556 ( U6904 , U2557 , INSTQUEUE_REG_9__0_ );
nand NAND2_4557 ( U6905 , U2556 , INSTQUEUE_REG_8__0_ );
nand NAND2_4558 ( U6906 , U2554 , INSTQUEUE_REG_7__0_ );
nand NAND2_4559 ( U6907 , U2553 , INSTQUEUE_REG_6__0_ );
nand NAND2_4560 ( U6908 , U2552 , INSTQUEUE_REG_5__0_ );
nand NAND2_4561 ( U6909 , U2551 , INSTQUEUE_REG_4__0_ );
nand NAND2_4562 ( U6910 , U2549 , INSTQUEUE_REG_3__0_ );
nand NAND2_4563 ( U6911 , U2548 , INSTQUEUE_REG_2__0_ );
nand NAND2_4564 ( U6912 , U2547 , INSTQUEUE_REG_1__0_ );
nand NAND2_4565 ( U6913 , U2546 , INSTQUEUE_REG_0__0_ );
nand NAND4_4566 ( U6914 , U4024 , U4023 , U4022 , U4021 );
nand NAND2_4567 ( U6915 , U4195 , U3221 );
nand NAND2_4568 ( U6916 , U2355 , SUB_357_U8 );
nand NAND2_4569 ( U6917 , U4195 , U3220 );
nand NAND2_4570 ( U6918 , SUB_357_U6 , U2355 );
nand NAND2_4571 ( U6919 , U4195 , U3219 );
nand NAND2_4572 ( U6920 , SUB_357_U9 , U2355 );
nand NAND2_4573 ( U6921 , U4195 , U3218 );
nand NAND2_4574 ( U6922 , SUB_357_U13 , U2355 );
nand NAND2_4575 ( U6923 , U4195 , U3217 );
nand NAND2_4576 ( U6924 , SUB_357_U11 , U2355 );
nand NAND2_4577 ( U6925 , R2182_U25 , U3281 );
nand NAND2_4578 ( U6926 , U4195 , U3216 );
nand NAND2_4579 ( U6927 , SUB_357_U12 , U2355 );
nand NAND2_4580 ( U6928 , R2182_U42 , U3281 );
nand NAND2_4581 ( U6929 , U2564 , INSTQUEUE_REG_15__7_ );
nand NAND2_4582 ( U6930 , U2563 , INSTQUEUE_REG_14__7_ );
nand NAND2_4583 ( U6931 , U2562 , INSTQUEUE_REG_13__7_ );
nand NAND2_4584 ( U6932 , U2561 , INSTQUEUE_REG_12__7_ );
nand NAND2_4585 ( U6933 , U2559 , INSTQUEUE_REG_11__7_ );
nand NAND2_4586 ( U6934 , U2558 , INSTQUEUE_REG_10__7_ );
nand NAND2_4587 ( U6935 , U2557 , INSTQUEUE_REG_9__7_ );
nand NAND2_4588 ( U6936 , U2556 , INSTQUEUE_REG_8__7_ );
nand NAND2_4589 ( U6937 , U2554 , INSTQUEUE_REG_7__7_ );
nand NAND2_4590 ( U6938 , U2553 , INSTQUEUE_REG_6__7_ );
nand NAND2_4591 ( U6939 , U2552 , INSTQUEUE_REG_5__7_ );
nand NAND2_4592 ( U6940 , U2551 , INSTQUEUE_REG_4__7_ );
nand NAND2_4593 ( U6941 , U2549 , INSTQUEUE_REG_3__7_ );
nand NAND2_4594 ( U6942 , U2548 , INSTQUEUE_REG_2__7_ );
nand NAND2_4595 ( U6943 , U2547 , INSTQUEUE_REG_1__7_ );
nand NAND2_4596 ( U6944 , U2546 , INSTQUEUE_REG_0__7_ );
nand NAND4_4597 ( U6945 , U4028 , U4027 , U4026 , U4025 );
nand NAND2_4598 ( U6946 , U2564 , INSTQUEUE_REG_15__6_ );
nand NAND2_4599 ( U6947 , U2563 , INSTQUEUE_REG_14__6_ );
nand NAND2_4600 ( U6948 , U2562 , INSTQUEUE_REG_13__6_ );
nand NAND2_4601 ( U6949 , U2561 , INSTQUEUE_REG_12__6_ );
nand NAND2_4602 ( U6950 , U2559 , INSTQUEUE_REG_11__6_ );
nand NAND2_4603 ( U6951 , U2558 , INSTQUEUE_REG_10__6_ );
nand NAND2_4604 ( U6952 , U2557 , INSTQUEUE_REG_9__6_ );
nand NAND2_4605 ( U6953 , U2556 , INSTQUEUE_REG_8__6_ );
nand NAND2_4606 ( U6954 , U2554 , INSTQUEUE_REG_7__6_ );
nand NAND2_4607 ( U6955 , U2553 , INSTQUEUE_REG_6__6_ );
nand NAND2_4608 ( U6956 , U2552 , INSTQUEUE_REG_5__6_ );
nand NAND2_4609 ( U6957 , U2551 , INSTQUEUE_REG_4__6_ );
nand NAND2_4610 ( U6958 , U2549 , INSTQUEUE_REG_3__6_ );
nand NAND2_4611 ( U6959 , U2548 , INSTQUEUE_REG_2__6_ );
nand NAND2_4612 ( U6960 , U2547 , INSTQUEUE_REG_1__6_ );
nand NAND2_4613 ( U6961 , U2546 , INSTQUEUE_REG_0__6_ );
nand NAND4_4614 ( U6962 , U4032 , U4031 , U4030 , U4029 );
nand NAND2_4615 ( U6963 , U2564 , INSTQUEUE_REG_15__5_ );
nand NAND2_4616 ( U6964 , U2563 , INSTQUEUE_REG_14__5_ );
nand NAND2_4617 ( U6965 , U2562 , INSTQUEUE_REG_13__5_ );
nand NAND2_4618 ( U6966 , U2561 , INSTQUEUE_REG_12__5_ );
nand NAND2_4619 ( U6967 , U2559 , INSTQUEUE_REG_11__5_ );
nand NAND2_4620 ( U6968 , U2558 , INSTQUEUE_REG_10__5_ );
nand NAND2_4621 ( U6969 , U2557 , INSTQUEUE_REG_9__5_ );
nand NAND2_4622 ( U6970 , U2556 , INSTQUEUE_REG_8__5_ );
nand NAND2_4623 ( U6971 , U2554 , INSTQUEUE_REG_7__5_ );
nand NAND2_4624 ( U6972 , U2553 , INSTQUEUE_REG_6__5_ );
nand NAND2_4625 ( U6973 , U2552 , INSTQUEUE_REG_5__5_ );
nand NAND2_4626 ( U6974 , U2551 , INSTQUEUE_REG_4__5_ );
nand NAND2_4627 ( U6975 , U2549 , INSTQUEUE_REG_3__5_ );
nand NAND2_4628 ( U6976 , U2548 , INSTQUEUE_REG_2__5_ );
nand NAND2_4629 ( U6977 , U2547 , INSTQUEUE_REG_1__5_ );
nand NAND2_4630 ( U6978 , U2546 , INSTQUEUE_REG_0__5_ );
nand NAND4_4631 ( U6979 , U4036 , U4035 , U4034 , U4033 );
nand NAND2_4632 ( U6980 , U2564 , INSTQUEUE_REG_15__4_ );
nand NAND2_4633 ( U6981 , U2563 , INSTQUEUE_REG_14__4_ );
nand NAND2_4634 ( U6982 , U2562 , INSTQUEUE_REG_13__4_ );
nand NAND2_4635 ( U6983 , U2561 , INSTQUEUE_REG_12__4_ );
nand NAND2_4636 ( U6984 , U2559 , INSTQUEUE_REG_11__4_ );
nand NAND2_4637 ( U6985 , U2558 , INSTQUEUE_REG_10__4_ );
nand NAND2_4638 ( U6986 , U2557 , INSTQUEUE_REG_9__4_ );
nand NAND2_4639 ( U6987 , U2556 , INSTQUEUE_REG_8__4_ );
nand NAND2_4640 ( U6988 , U2554 , INSTQUEUE_REG_7__4_ );
nand NAND2_4641 ( U6989 , U2553 , INSTQUEUE_REG_6__4_ );
nand NAND2_4642 ( U6990 , U2552 , INSTQUEUE_REG_5__4_ );
nand NAND2_4643 ( U6991 , U2551 , INSTQUEUE_REG_4__4_ );
nand NAND2_4644 ( U6992 , U2549 , INSTQUEUE_REG_3__4_ );
nand NAND2_4645 ( U6993 , U2548 , INSTQUEUE_REG_2__4_ );
nand NAND2_4646 ( U6994 , U2547 , INSTQUEUE_REG_1__4_ );
nand NAND2_4647 ( U6995 , U2564 , INSTQUEUE_REG_15__3_ );
nand NAND2_4648 ( U6996 , U2563 , INSTQUEUE_REG_14__3_ );
nand NAND2_4649 ( U6997 , U2562 , INSTQUEUE_REG_13__3_ );
nand NAND2_4650 ( U6998 , U2561 , INSTQUEUE_REG_12__3_ );
nand NAND2_4651 ( U6999 , U2559 , INSTQUEUE_REG_11__3_ );
nand NAND2_4652 ( U7000 , U2558 , INSTQUEUE_REG_10__3_ );
nand NAND2_4653 ( U7001 , U2557 , INSTQUEUE_REG_9__3_ );
nand NAND2_4654 ( U7002 , U2556 , INSTQUEUE_REG_8__3_ );
nand NAND2_4655 ( U7003 , U2554 , INSTQUEUE_REG_7__3_ );
nand NAND2_4656 ( U7004 , U2553 , INSTQUEUE_REG_6__3_ );
nand NAND2_4657 ( U7005 , U2552 , INSTQUEUE_REG_5__3_ );
nand NAND2_4658 ( U7006 , U2551 , INSTQUEUE_REG_4__3_ );
nand NAND2_4659 ( U7007 , U2549 , INSTQUEUE_REG_3__3_ );
nand NAND2_4660 ( U7008 , U2548 , INSTQUEUE_REG_2__3_ );
nand NAND2_4661 ( U7009 , U2547 , INSTQUEUE_REG_1__3_ );
nand NAND2_4662 ( U7010 , U2546 , INSTQUEUE_REG_0__3_ );
nand NAND4_4663 ( U7011 , U4044 , U4043 , U4042 , U4041 );
nand NAND2_4664 ( U7012 , U2564 , INSTQUEUE_REG_15__2_ );
nand NAND2_4665 ( U7013 , U2563 , INSTQUEUE_REG_14__2_ );
nand NAND2_4666 ( U7014 , U2562 , INSTQUEUE_REG_13__2_ );
nand NAND2_4667 ( U7015 , U2561 , INSTQUEUE_REG_12__2_ );
nand NAND2_4668 ( U7016 , U2559 , INSTQUEUE_REG_11__2_ );
nand NAND2_4669 ( U7017 , U2558 , INSTQUEUE_REG_10__2_ );
nand NAND2_4670 ( U7018 , U2557 , INSTQUEUE_REG_9__2_ );
nand NAND2_4671 ( U7019 , U2556 , INSTQUEUE_REG_8__2_ );
nand NAND2_4672 ( U7020 , U2554 , INSTQUEUE_REG_7__2_ );
nand NAND2_4673 ( U7021 , U2553 , INSTQUEUE_REG_6__2_ );
nand NAND2_4674 ( U7022 , U2552 , INSTQUEUE_REG_5__2_ );
nand NAND2_4675 ( U7023 , U2551 , INSTQUEUE_REG_4__2_ );
nand NAND2_4676 ( U7024 , U2549 , INSTQUEUE_REG_3__2_ );
nand NAND2_4677 ( U7025 , U2548 , INSTQUEUE_REG_2__2_ );
nand NAND2_4678 ( U7026 , U2547 , INSTQUEUE_REG_1__2_ );
nand NAND2_4679 ( U7027 , U2546 , INSTQUEUE_REG_0__2_ );
nand NAND4_4680 ( U7028 , U4048 , U4047 , U4046 , U4045 );
nand NAND2_4681 ( U7029 , U4195 , U3215 );
nand NAND2_4682 ( U7030 , SUB_357_U7 , U2355 );
nand NAND2_4683 ( U7031 , R2182_U33 , U3281 );
nand NAND2_4684 ( U7032 , U4195 , U3214 );
nand NAND2_4685 ( U7033 , SUB_357_U10 , U2355 );
nand NAND2_4686 ( U7034 , R2182_U34 , U3281 );
nand NAND2_4687 ( U7035 , U4194 , U3221 );
nand NAND2_4688 ( U7036 , U4180 , INSTQUEUE_REG_0__7_ );
nand NAND2_4689 ( U7037 , U4194 , U3220 );
nand NAND2_4690 ( U7038 , U4180 , INSTQUEUE_REG_0__6_ );
nand NAND2_4691 ( U7039 , U4194 , U3219 );
nand NAND2_4692 ( U7040 , U4180 , INSTQUEUE_REG_0__5_ );
nand NAND2_4693 ( U7041 , U4194 , U3218 );
nand NAND2_4694 ( U7042 , U4194 , U3217 );
nand NAND2_4695 ( U7043 , U4180 , INSTQUEUE_REG_0__3_ );
nand NAND2_4696 ( U7044 , U4194 , U3216 );
nand NAND2_4697 ( U7045 , U4180 , INSTQUEUE_REG_0__2_ );
nand NAND2_4698 ( U7046 , U4194 , U3215 );
nand NAND2_4699 ( U7047 , U4180 , INSTQUEUE_REG_0__1_ );
nand NAND2_4700 ( U7048 , U4194 , U3214 );
nand NAND2_4701 ( U7049 , U3221 , U4388 );
nand NAND2_4702 ( U7050 , U4180 , INSTQUEUE_REG_0__0_ );
nand NAND2_4703 ( U7051 , U3415 , U3414 );
nand NAND2_4704 ( U7052 , INSTQUEUERD_ADDR_REG_3_ , U3251 );
not NOT1_4705 ( U7053 , U3432 );
nand NAND2_4706 ( U7054 , U2582 , INSTQUEUE_REG_8__7_ );
nand NAND2_4707 ( U7055 , U2581 , INSTQUEUE_REG_9__7_ );
nand NAND2_4708 ( U7056 , U2580 , INSTQUEUE_REG_10__7_ );
nand NAND2_4709 ( U7057 , U2579 , INSTQUEUE_REG_11__7_ );
nand NAND2_4710 ( U7058 , U2577 , INSTQUEUE_REG_12__7_ );
nand NAND2_4711 ( U7059 , U2576 , INSTQUEUE_REG_13__7_ );
nand NAND2_4712 ( U7060 , U2575 , INSTQUEUE_REG_14__7_ );
nand NAND2_4713 ( U7061 , U2574 , INSTQUEUE_REG_15__7_ );
nand NAND2_4714 ( U7062 , U2573 , INSTQUEUE_REG_0__7_ );
nand NAND2_4715 ( U7063 , U2572 , INSTQUEUE_REG_1__7_ );
nand NAND2_4716 ( U7064 , U2571 , INSTQUEUE_REG_2__7_ );
nand NAND2_4717 ( U7065 , U2570 , INSTQUEUE_REG_3__7_ );
nand NAND2_4718 ( U7066 , U2568 , INSTQUEUE_REG_4__7_ );
nand NAND2_4719 ( U7067 , U2567 , INSTQUEUE_REG_5__7_ );
nand NAND2_4720 ( U7068 , U2566 , INSTQUEUE_REG_6__7_ );
nand NAND2_4721 ( U7069 , U2565 , INSTQUEUE_REG_7__7_ );
nand NAND4_4722 ( U7070 , U4054 , U4053 , U4052 , U4051 );
nand NAND2_4723 ( U7071 , U3412 , U3408 );
nand NAND2_4724 ( U7072 , U4061 , U4179 );
nand NAND2_4725 ( U7073 , U7072 , U3409 );
nand NAND2_4726 ( U7074 , U4491 , U3265 );
not NOT1_4727 ( U7075 , U3232 );
nand NAND4_4728 ( U7076 , U4388 , U4491 , U4142 , U3381 );
nand NAND2_4729 ( U7077 , U4177 , STATE2_REG_0_ );
nand NAND2_4730 ( U7078 , U4055 , U3232 );
not NOT1_4731 ( U7079 , U3438 );
nand NAND3_4732 ( U7080 , U3438 , U5480 , U7617 );
nand NAND2_4733 ( U7081 , U4182 , U7080 );
not NOT1_4734 ( U7082 , U3437 );
nand NAND2_4735 ( U7083 , INSTQUEUEWR_ADDR_REG_3_ , U3284 );
nand NAND2_4736 ( U7084 , INSTQUEUERD_ADDR_REG_3_ , U3437 );
nand NAND2_4737 ( U7085 , U4191 , U3347 );
nand NAND2_4738 ( U7086 , U2582 , INSTQUEUE_REG_8__6_ );
nand NAND2_4739 ( U7087 , U2581 , INSTQUEUE_REG_9__6_ );
nand NAND2_4740 ( U7088 , U2580 , INSTQUEUE_REG_10__6_ );
nand NAND2_4741 ( U7089 , U2579 , INSTQUEUE_REG_11__6_ );
nand NAND2_4742 ( U7090 , U2577 , INSTQUEUE_REG_12__6_ );
nand NAND2_4743 ( U7091 , U2576 , INSTQUEUE_REG_13__6_ );
nand NAND2_4744 ( U7092 , U2575 , INSTQUEUE_REG_14__6_ );
nand NAND2_4745 ( U7093 , U2574 , INSTQUEUE_REG_15__6_ );
nand NAND2_4746 ( U7094 , U2573 , INSTQUEUE_REG_0__6_ );
nand NAND2_4747 ( U7095 , U2572 , INSTQUEUE_REG_1__6_ );
nand NAND2_4748 ( U7096 , U2571 , INSTQUEUE_REG_2__6_ );
nand NAND2_4749 ( U7097 , U2570 , INSTQUEUE_REG_3__6_ );
nand NAND2_4750 ( U7098 , U2568 , INSTQUEUE_REG_4__6_ );
nand NAND2_4751 ( U7099 , U2567 , INSTQUEUE_REG_5__6_ );
nand NAND2_4752 ( U7100 , U2566 , INSTQUEUE_REG_6__6_ );
nand NAND2_4753 ( U7101 , U2565 , INSTQUEUE_REG_7__6_ );
nand NAND4_4754 ( U7102 , U4070 , U4069 , U4068 , U4067 );
nand NAND2_4755 ( U7103 , U2582 , INSTQUEUE_REG_8__5_ );
nand NAND2_4756 ( U7104 , U2581 , INSTQUEUE_REG_9__5_ );
nand NAND2_4757 ( U7105 , U2580 , INSTQUEUE_REG_10__5_ );
nand NAND2_4758 ( U7106 , U2579 , INSTQUEUE_REG_11__5_ );
nand NAND2_4759 ( U7107 , U2577 , INSTQUEUE_REG_12__5_ );
nand NAND2_4760 ( U7108 , U2576 , INSTQUEUE_REG_13__5_ );
nand NAND2_4761 ( U7109 , U2575 , INSTQUEUE_REG_14__5_ );
nand NAND2_4762 ( U7110 , U2574 , INSTQUEUE_REG_15__5_ );
nand NAND2_4763 ( U7111 , U2573 , INSTQUEUE_REG_0__5_ );
nand NAND2_4764 ( U7112 , U2572 , INSTQUEUE_REG_1__5_ );
nand NAND2_4765 ( U7113 , U2571 , INSTQUEUE_REG_2__5_ );
nand NAND2_4766 ( U7114 , U2570 , INSTQUEUE_REG_3__5_ );
nand NAND2_4767 ( U7115 , U2568 , INSTQUEUE_REG_4__5_ );
nand NAND2_4768 ( U7116 , U2567 , INSTQUEUE_REG_5__5_ );
nand NAND2_4769 ( U7117 , U2566 , INSTQUEUE_REG_6__5_ );
nand NAND2_4770 ( U7118 , U2565 , INSTQUEUE_REG_7__5_ );
nand NAND4_4771 ( U7119 , U4074 , U4073 , U4072 , U4071 );
nand NAND2_4772 ( U7120 , U2582 , INSTQUEUE_REG_8__4_ );
nand NAND2_4773 ( U7121 , U2581 , INSTQUEUE_REG_9__4_ );
nand NAND2_4774 ( U7122 , U2580 , INSTQUEUE_REG_10__4_ );
nand NAND2_4775 ( U7123 , U2579 , INSTQUEUE_REG_11__4_ );
nand NAND2_4776 ( U7124 , U2577 , INSTQUEUE_REG_12__4_ );
nand NAND2_4777 ( U7125 , U2576 , INSTQUEUE_REG_13__4_ );
nand NAND2_4778 ( U7126 , U2575 , INSTQUEUE_REG_14__4_ );
nand NAND2_4779 ( U7127 , U2574 , INSTQUEUE_REG_15__4_ );
nand NAND2_4780 ( U7128 , U2572 , INSTQUEUE_REG_1__4_ );
nand NAND2_4781 ( U7129 , U2571 , INSTQUEUE_REG_2__4_ );
nand NAND2_4782 ( U7130 , U2570 , INSTQUEUE_REG_3__4_ );
nand NAND2_4783 ( U7131 , U2568 , INSTQUEUE_REG_4__4_ );
nand NAND2_4784 ( U7132 , U2567 , INSTQUEUE_REG_5__4_ );
nand NAND2_4785 ( U7133 , U2566 , INSTQUEUE_REG_6__4_ );
nand NAND2_4786 ( U7134 , U2565 , INSTQUEUE_REG_7__4_ );
nand NAND2_4787 ( U7135 , U2582 , INSTQUEUE_REG_8__3_ );
nand NAND2_4788 ( U7136 , U2581 , INSTQUEUE_REG_9__3_ );
nand NAND2_4789 ( U7137 , U2580 , INSTQUEUE_REG_10__3_ );
nand NAND2_4790 ( U7138 , U2579 , INSTQUEUE_REG_11__3_ );
nand NAND2_4791 ( U7139 , U2577 , INSTQUEUE_REG_12__3_ );
nand NAND2_4792 ( U7140 , U2576 , INSTQUEUE_REG_13__3_ );
nand NAND2_4793 ( U7141 , U2575 , INSTQUEUE_REG_14__3_ );
nand NAND2_4794 ( U7142 , U2574 , INSTQUEUE_REG_15__3_ );
nand NAND2_4795 ( U7143 , U2573 , INSTQUEUE_REG_0__3_ );
nand NAND2_4796 ( U7144 , U2572 , INSTQUEUE_REG_1__3_ );
nand NAND2_4797 ( U7145 , U2571 , INSTQUEUE_REG_2__3_ );
nand NAND2_4798 ( U7146 , U2570 , INSTQUEUE_REG_3__3_ );
nand NAND2_4799 ( U7147 , U2568 , INSTQUEUE_REG_4__3_ );
nand NAND2_4800 ( U7148 , U2567 , INSTQUEUE_REG_5__3_ );
nand NAND2_4801 ( U7149 , U2566 , INSTQUEUE_REG_6__3_ );
nand NAND2_4802 ( U7150 , U2565 , INSTQUEUE_REG_7__3_ );
nand NAND4_4803 ( U7151 , U4083 , U4082 , U4081 , U4080 );
nand NAND2_4804 ( U7152 , U2582 , INSTQUEUE_REG_8__2_ );
nand NAND2_4805 ( U7153 , U2581 , INSTQUEUE_REG_9__2_ );
nand NAND2_4806 ( U7154 , U2580 , INSTQUEUE_REG_10__2_ );
nand NAND2_4807 ( U7155 , U2579 , INSTQUEUE_REG_11__2_ );
nand NAND2_4808 ( U7156 , U2577 , INSTQUEUE_REG_12__2_ );
nand NAND2_4809 ( U7157 , U2576 , INSTQUEUE_REG_13__2_ );
nand NAND2_4810 ( U7158 , U2575 , INSTQUEUE_REG_14__2_ );
nand NAND2_4811 ( U7159 , U2574 , INSTQUEUE_REG_15__2_ );
nand NAND2_4812 ( U7160 , U2573 , INSTQUEUE_REG_0__2_ );
nand NAND2_4813 ( U7161 , U2572 , INSTQUEUE_REG_1__2_ );
nand NAND2_4814 ( U7162 , U2571 , INSTQUEUE_REG_2__2_ );
nand NAND2_4815 ( U7163 , U2570 , INSTQUEUE_REG_3__2_ );
nand NAND2_4816 ( U7164 , U2568 , INSTQUEUE_REG_4__2_ );
nand NAND2_4817 ( U7165 , U2567 , INSTQUEUE_REG_5__2_ );
nand NAND2_4818 ( U7166 , U2566 , INSTQUEUE_REG_6__2_ );
nand NAND2_4819 ( U7167 , U2565 , INSTQUEUE_REG_7__2_ );
nand NAND4_4820 ( U7168 , U4087 , U4086 , U4085 , U4084 );
nand NAND2_4821 ( U7169 , U2582 , INSTQUEUE_REG_8__1_ );
nand NAND2_4822 ( U7170 , U2581 , INSTQUEUE_REG_9__1_ );
nand NAND2_4823 ( U7171 , U2580 , INSTQUEUE_REG_10__1_ );
nand NAND2_4824 ( U7172 , U2579 , INSTQUEUE_REG_11__1_ );
nand NAND2_4825 ( U7173 , U2577 , INSTQUEUE_REG_12__1_ );
nand NAND2_4826 ( U7174 , U2576 , INSTQUEUE_REG_13__1_ );
nand NAND2_4827 ( U7175 , U2575 , INSTQUEUE_REG_14__1_ );
nand NAND2_4828 ( U7176 , U2574 , INSTQUEUE_REG_15__1_ );
nand NAND2_4829 ( U7177 , U2573 , INSTQUEUE_REG_0__1_ );
nand NAND2_4830 ( U7178 , U2572 , INSTQUEUE_REG_1__1_ );
nand NAND2_4831 ( U7179 , U2571 , INSTQUEUE_REG_2__1_ );
nand NAND2_4832 ( U7180 , U2570 , INSTQUEUE_REG_3__1_ );
nand NAND2_4833 ( U7181 , U2568 , INSTQUEUE_REG_4__1_ );
nand NAND2_4834 ( U7182 , U2567 , INSTQUEUE_REG_5__1_ );
nand NAND2_4835 ( U7183 , U2566 , INSTQUEUE_REG_6__1_ );
nand NAND2_4836 ( U7184 , U2565 , INSTQUEUE_REG_7__1_ );
nand NAND4_4837 ( U7185 , U4091 , U4090 , U4089 , U4088 );
nand NAND2_4838 ( U7186 , U2582 , INSTQUEUE_REG_8__0_ );
nand NAND2_4839 ( U7187 , U2581 , INSTQUEUE_REG_9__0_ );
nand NAND2_4840 ( U7188 , U2580 , INSTQUEUE_REG_10__0_ );
nand NAND2_4841 ( U7189 , U2579 , INSTQUEUE_REG_11__0_ );
nand NAND2_4842 ( U7190 , U2577 , INSTQUEUE_REG_12__0_ );
nand NAND2_4843 ( U7191 , U2576 , INSTQUEUE_REG_13__0_ );
nand NAND2_4844 ( U7192 , U2575 , INSTQUEUE_REG_14__0_ );
nand NAND2_4845 ( U7193 , U2574 , INSTQUEUE_REG_15__0_ );
nand NAND2_4846 ( U7194 , U2573 , INSTQUEUE_REG_0__0_ );
nand NAND2_4847 ( U7195 , U2572 , INSTQUEUE_REG_1__0_ );
nand NAND2_4848 ( U7196 , U2571 , INSTQUEUE_REG_2__0_ );
nand NAND2_4849 ( U7197 , U2570 , INSTQUEUE_REG_3__0_ );
nand NAND2_4850 ( U7198 , U2568 , INSTQUEUE_REG_4__0_ );
nand NAND2_4851 ( U7199 , U2567 , INSTQUEUE_REG_5__0_ );
nand NAND2_4852 ( U7200 , U2566 , INSTQUEUE_REG_6__0_ );
nand NAND2_4853 ( U7201 , U2565 , INSTQUEUE_REG_7__0_ );
nand NAND4_4854 ( U7202 , U4095 , U4094 , U4093 , U4092 );
nand NAND2_4855 ( U7203 , INSTQUEUEWR_ADDR_REG_2_ , U3284 );
nand NAND2_4856 ( U7204 , U4191 , U3442 );
nand NAND2_4857 ( U7205 , INSTQUEUEWR_ADDR_REG_1_ , U3284 );
nand NAND2_4858 ( U7206 , U4191 , U3222 );
not NOT1_4859 ( U7207 , U4171 );
nand NAND2_4860 ( U7208 , U2602 , INSTQUEUE_REG_8__7_ );
nand NAND2_4861 ( U7209 , U2601 , INSTQUEUE_REG_9__7_ );
nand NAND2_4862 ( U7210 , U2600 , INSTQUEUE_REG_10__7_ );
nand NAND2_4863 ( U7211 , U2599 , INSTQUEUE_REG_11__7_ );
nand NAND2_4864 ( U7212 , U2597 , INSTQUEUE_REG_12__7_ );
nand NAND2_4865 ( U7213 , U2596 , INSTQUEUE_REG_13__7_ );
nand NAND2_4866 ( U7214 , U2595 , INSTQUEUE_REG_14__7_ );
nand NAND2_4867 ( U7215 , U2594 , INSTQUEUE_REG_15__7_ );
nand NAND2_4868 ( U7216 , U2592 , INSTQUEUE_REG_0__7_ );
nand NAND2_4869 ( U7217 , U2591 , INSTQUEUE_REG_1__7_ );
nand NAND2_4870 ( U7218 , U2590 , INSTQUEUE_REG_2__7_ );
nand NAND2_4871 ( U7219 , U2589 , INSTQUEUE_REG_3__7_ );
nand NAND2_4872 ( U7220 , U2587 , INSTQUEUE_REG_4__7_ );
nand NAND2_4873 ( U7221 , U2586 , INSTQUEUE_REG_5__7_ );
nand NAND2_4874 ( U7222 , U2585 , INSTQUEUE_REG_6__7_ );
nand NAND2_4875 ( U7223 , U2584 , INSTQUEUE_REG_7__7_ );
nand NAND4_4876 ( U7224 , U4112 , U4111 , U4110 , U4109 );
nand NAND2_4877 ( U7225 , U2602 , INSTQUEUE_REG_8__6_ );
nand NAND2_4878 ( U7226 , U2601 , INSTQUEUE_REG_9__6_ );
nand NAND2_4879 ( U7227 , U2600 , INSTQUEUE_REG_10__6_ );
nand NAND2_4880 ( U7228 , U2599 , INSTQUEUE_REG_11__6_ );
nand NAND2_4881 ( U7229 , U2597 , INSTQUEUE_REG_12__6_ );
nand NAND2_4882 ( U7230 , U2596 , INSTQUEUE_REG_13__6_ );
nand NAND2_4883 ( U7231 , U2595 , INSTQUEUE_REG_14__6_ );
nand NAND2_4884 ( U7232 , U2594 , INSTQUEUE_REG_15__6_ );
nand NAND2_4885 ( U7233 , U2592 , INSTQUEUE_REG_0__6_ );
nand NAND2_4886 ( U7234 , U2591 , INSTQUEUE_REG_1__6_ );
nand NAND2_4887 ( U7235 , U2590 , INSTQUEUE_REG_2__6_ );
nand NAND2_4888 ( U7236 , U2589 , INSTQUEUE_REG_3__6_ );
nand NAND2_4889 ( U7237 , U2587 , INSTQUEUE_REG_4__6_ );
nand NAND2_4890 ( U7238 , U2586 , INSTQUEUE_REG_5__6_ );
nand NAND2_4891 ( U7239 , U2585 , INSTQUEUE_REG_6__6_ );
nand NAND2_4892 ( U7240 , U2584 , INSTQUEUE_REG_7__6_ );
nand NAND4_4893 ( U7241 , U4116 , U4115 , U4114 , U4113 );
nand NAND2_4894 ( U7242 , U2602 , INSTQUEUE_REG_8__5_ );
nand NAND2_4895 ( U7243 , U2601 , INSTQUEUE_REG_9__5_ );
nand NAND2_4896 ( U7244 , U2600 , INSTQUEUE_REG_10__5_ );
nand NAND2_4897 ( U7245 , U2599 , INSTQUEUE_REG_11__5_ );
nand NAND2_4898 ( U7246 , U2597 , INSTQUEUE_REG_12__5_ );
nand NAND2_4899 ( U7247 , U2596 , INSTQUEUE_REG_13__5_ );
nand NAND2_4900 ( U7248 , U2595 , INSTQUEUE_REG_14__5_ );
nand NAND2_4901 ( U7249 , U2594 , INSTQUEUE_REG_15__5_ );
nand NAND2_4902 ( U7250 , U2592 , INSTQUEUE_REG_0__5_ );
nand NAND2_4903 ( U7251 , U2591 , INSTQUEUE_REG_1__5_ );
nand NAND2_4904 ( U7252 , U2590 , INSTQUEUE_REG_2__5_ );
nand NAND2_4905 ( U7253 , U2589 , INSTQUEUE_REG_3__5_ );
nand NAND2_4906 ( U7254 , U2587 , INSTQUEUE_REG_4__5_ );
nand NAND2_4907 ( U7255 , U2586 , INSTQUEUE_REG_5__5_ );
nand NAND2_4908 ( U7256 , U2585 , INSTQUEUE_REG_6__5_ );
nand NAND2_4909 ( U7257 , U2584 , INSTQUEUE_REG_7__5_ );
nand NAND4_4910 ( U7258 , U4120 , U4119 , U4118 , U4117 );
nand NAND2_4911 ( U7259 , U2602 , INSTQUEUE_REG_8__4_ );
nand NAND2_4912 ( U7260 , U2601 , INSTQUEUE_REG_9__4_ );
nand NAND2_4913 ( U7261 , U2600 , INSTQUEUE_REG_10__4_ );
nand NAND2_4914 ( U7262 , U2599 , INSTQUEUE_REG_11__4_ );
nand NAND2_4915 ( U7263 , U2597 , INSTQUEUE_REG_12__4_ );
nand NAND2_4916 ( U7264 , U2596 , INSTQUEUE_REG_13__4_ );
nand NAND2_4917 ( U7265 , U2595 , INSTQUEUE_REG_14__4_ );
nand NAND2_4918 ( U7266 , U2594 , INSTQUEUE_REG_15__4_ );
nand NAND2_4919 ( U7267 , U2591 , INSTQUEUE_REG_1__4_ );
nand NAND2_4920 ( U7268 , U2590 , INSTQUEUE_REG_2__4_ );
nand NAND2_4921 ( U7269 , U2589 , INSTQUEUE_REG_3__4_ );
nand NAND2_4922 ( U7270 , U2587 , INSTQUEUE_REG_4__4_ );
nand NAND2_4923 ( U7271 , U2586 , INSTQUEUE_REG_5__4_ );
nand NAND2_4924 ( U7272 , U2585 , INSTQUEUE_REG_6__4_ );
nand NAND2_4925 ( U7273 , U2584 , INSTQUEUE_REG_7__4_ );
nand NAND2_4926 ( U7274 , U2602 , INSTQUEUE_REG_8__3_ );
nand NAND2_4927 ( U7275 , U2601 , INSTQUEUE_REG_9__3_ );
nand NAND2_4928 ( U7276 , U2600 , INSTQUEUE_REG_10__3_ );
nand NAND2_4929 ( U7277 , U2599 , INSTQUEUE_REG_11__3_ );
nand NAND2_4930 ( U7278 , U2597 , INSTQUEUE_REG_12__3_ );
nand NAND2_4931 ( U7279 , U2596 , INSTQUEUE_REG_13__3_ );
nand NAND2_4932 ( U7280 , U2595 , INSTQUEUE_REG_14__3_ );
nand NAND2_4933 ( U7281 , U2594 , INSTQUEUE_REG_15__3_ );
nand NAND2_4934 ( U7282 , U2592 , INSTQUEUE_REG_0__3_ );
nand NAND2_4935 ( U7283 , U2591 , INSTQUEUE_REG_1__3_ );
nand NAND2_4936 ( U7284 , U2590 , INSTQUEUE_REG_2__3_ );
nand NAND2_4937 ( U7285 , U2589 , INSTQUEUE_REG_3__3_ );
nand NAND2_4938 ( U7286 , U2587 , INSTQUEUE_REG_4__3_ );
nand NAND2_4939 ( U7287 , U2586 , INSTQUEUE_REG_5__3_ );
nand NAND2_4940 ( U7288 , U2585 , INSTQUEUE_REG_6__3_ );
nand NAND2_4941 ( U7289 , U2584 , INSTQUEUE_REG_7__3_ );
nand NAND4_4942 ( U7290 , U4128 , U4127 , U4126 , U4125 );
nand NAND2_4943 ( U7291 , U2602 , INSTQUEUE_REG_8__2_ );
nand NAND2_4944 ( U7292 , U2601 , INSTQUEUE_REG_9__2_ );
nand NAND2_4945 ( U7293 , U2600 , INSTQUEUE_REG_10__2_ );
nand NAND2_4946 ( U7294 , U2599 , INSTQUEUE_REG_11__2_ );
nand NAND2_4947 ( U7295 , U2597 , INSTQUEUE_REG_12__2_ );
nand NAND2_4948 ( U7296 , U2596 , INSTQUEUE_REG_13__2_ );
nand NAND2_4949 ( U7297 , U2595 , INSTQUEUE_REG_14__2_ );
nand NAND2_4950 ( U7298 , U2594 , INSTQUEUE_REG_15__2_ );
nand NAND2_4951 ( U7299 , U2592 , INSTQUEUE_REG_0__2_ );
nand NAND2_4952 ( U7300 , U2591 , INSTQUEUE_REG_1__2_ );
nand NAND2_4953 ( U7301 , U2590 , INSTQUEUE_REG_2__2_ );
nand NAND2_4954 ( U7302 , U2589 , INSTQUEUE_REG_3__2_ );
nand NAND2_4955 ( U7303 , U2587 , INSTQUEUE_REG_4__2_ );
nand NAND2_4956 ( U7304 , U2586 , INSTQUEUE_REG_5__2_ );
nand NAND2_4957 ( U7305 , U2585 , INSTQUEUE_REG_6__2_ );
nand NAND2_4958 ( U7306 , U2584 , INSTQUEUE_REG_7__2_ );
nand NAND4_4959 ( U7307 , U4132 , U4131 , U4130 , U4129 );
nand NAND2_4960 ( U7308 , U2602 , INSTQUEUE_REG_8__1_ );
nand NAND2_4961 ( U7309 , U2601 , INSTQUEUE_REG_9__1_ );
nand NAND2_4962 ( U7310 , U2600 , INSTQUEUE_REG_10__1_ );
nand NAND2_4963 ( U7311 , U2599 , INSTQUEUE_REG_11__1_ );
nand NAND2_4964 ( U7312 , U2597 , INSTQUEUE_REG_12__1_ );
nand NAND2_4965 ( U7313 , U2596 , INSTQUEUE_REG_13__1_ );
nand NAND2_4966 ( U7314 , U2595 , INSTQUEUE_REG_14__1_ );
nand NAND2_4967 ( U7315 , U2594 , INSTQUEUE_REG_15__1_ );
nand NAND2_4968 ( U7316 , U2592 , INSTQUEUE_REG_0__1_ );
nand NAND2_4969 ( U7317 , U2591 , INSTQUEUE_REG_1__1_ );
nand NAND2_4970 ( U7318 , U2590 , INSTQUEUE_REG_2__1_ );
nand NAND2_4971 ( U7319 , U2589 , INSTQUEUE_REG_3__1_ );
nand NAND2_4972 ( U7320 , U2587 , INSTQUEUE_REG_4__1_ );
nand NAND2_4973 ( U7321 , U2586 , INSTQUEUE_REG_5__1_ );
nand NAND2_4974 ( U7322 , U2585 , INSTQUEUE_REG_6__1_ );
nand NAND2_4975 ( U7323 , U2584 , INSTQUEUE_REG_7__1_ );
nand NAND4_4976 ( U7324 , U4136 , U4135 , U4134 , U4133 );
nand NAND2_4977 ( U7325 , U2602 , INSTQUEUE_REG_8__0_ );
nand NAND2_4978 ( U7326 , U2601 , INSTQUEUE_REG_9__0_ );
nand NAND2_4979 ( U7327 , U2600 , INSTQUEUE_REG_10__0_ );
nand NAND2_4980 ( U7328 , U2599 , INSTQUEUE_REG_11__0_ );
nand NAND2_4981 ( U7329 , U2597 , INSTQUEUE_REG_12__0_ );
nand NAND2_4982 ( U7330 , U2596 , INSTQUEUE_REG_13__0_ );
nand NAND2_4983 ( U7331 , U2595 , INSTQUEUE_REG_14__0_ );
nand NAND2_4984 ( U7332 , U2594 , INSTQUEUE_REG_15__0_ );
nand NAND2_4985 ( U7333 , U2592 , INSTQUEUE_REG_0__0_ );
nand NAND2_4986 ( U7334 , U2591 , INSTQUEUE_REG_1__0_ );
nand NAND2_4987 ( U7335 , U2590 , INSTQUEUE_REG_2__0_ );
nand NAND2_4988 ( U7336 , U2589 , INSTQUEUE_REG_3__0_ );
nand NAND2_4989 ( U7337 , U2587 , INSTQUEUE_REG_4__0_ );
nand NAND2_4990 ( U7338 , U2586 , INSTQUEUE_REG_5__0_ );
nand NAND2_4991 ( U7339 , U2585 , INSTQUEUE_REG_6__0_ );
nand NAND2_4992 ( U7340 , U2584 , INSTQUEUE_REG_7__0_ );
nand NAND4_4993 ( U7341 , U4140 , U4139 , U4138 , U4137 );
nand NAND3_4994 ( U7342 , U4219 , U2354 , U4222 );
nand NAND2_4995 ( U7343 , U4141 , U7075 );
nand NAND2_4996 ( U7344 , U3383 , U3397 );
nand NAND2_4997 ( U7345 , U4222 , U7344 );
nand NAND2_4998 ( U7346 , U4178 , U2452 );
nand NAND2_4999 ( U7347 , U7343 , U3258 );
nand NAND2_5000 ( U7348 , U4196 , U7076 );
nand NAND2_5001 ( U7349 , U4148 , U4196 );
nand NAND2_5002 ( U7350 , U2451 , U4198 );
nand NAND5_5003 ( U7351 , U3407 , U3421 , U4183 , U7350 , U7349 );
nand NAND2_5004 ( U7352 , R2238_U6 , U7351 );
nand NAND2_5005 ( U7353 , SUB_450_U6 , U2354 );
nand NAND2_5006 ( U7354 , R2238_U19 , U7351 );
nand NAND2_5007 ( U7355 , SUB_450_U19 , U2354 );
nand NAND2_5008 ( U7356 , R2238_U20 , U7351 );
nand NAND2_5009 ( U7357 , SUB_450_U20 , U2354 );
nand NAND2_5010 ( U7358 , R2238_U21 , U7351 );
nand NAND2_5011 ( U7359 , SUB_450_U21 , U2354 );
nand NAND2_5012 ( U7360 , R2238_U22 , U7351 );
nand NAND2_5013 ( U7361 , SUB_450_U22 , U2354 );
nand NAND2_5014 ( U7362 , R2238_U7 , U7351 );
nand NAND2_5015 ( U7363 , SUB_450_U7 , U2354 );
nand NAND2_5016 ( U7364 , R2238_U19 , U4180 );
nand NAND2_5017 ( U7365 , INSTQUEUERD_ADDR_REG_4_ , U3281 );
nand NAND2_5018 ( U7366 , R2238_U20 , U4180 );
nand NAND2_5019 ( U7367 , INSTQUEUERD_ADDR_REG_3_ , U3281 );
nand NAND2_5020 ( U7368 , STATE2_REG_0_ , U4161 );
nand NAND2_5021 ( U7369 , U3407 , U7368 );
nand NAND2_5022 ( U7370 , R2238_U21 , U4180 );
nand NAND2_5023 ( U7371 , INSTQUEUERD_ADDR_REG_2_ , U3281 );
nand NAND2_5024 ( U7372 , U2450 , U3258 );
nand NAND2_5025 ( U7373 , R2238_U22 , U4180 );
nand NAND2_5026 ( U7374 , INSTQUEUERD_ADDR_REG_1_ , U3281 );
nand NAND2_5027 ( U7375 , U2451 , U3271 );
nand NAND2_5028 ( U7376 , R2238_U7 , U4180 );
nand NAND2_5029 ( U7377 , INSTQUEUERD_ADDR_REG_0_ , U3281 );
nand NAND2_5030 ( U7378 , U3380 , U3277 );
nand NAND2_5031 ( U7379 , U3271 , U3436 );
nand NAND2_5032 ( U7380 , INSTADDRPOINTER_REG_9_ , U7379 );
nand NAND2_5033 ( U7381 , EBX_REG_9_ , U7378 );
nand NAND2_5034 ( U7382 , INSTADDRPOINTER_REG_8_ , U7379 );
nand NAND2_5035 ( U7383 , EBX_REG_8_ , U7378 );
nand NAND2_5036 ( U7384 , INSTADDRPOINTER_REG_7_ , U7379 );
nand NAND2_5037 ( U7385 , EBX_REG_7_ , U7378 );
nand NAND2_5038 ( U7386 , INSTADDRPOINTER_REG_6_ , U7379 );
nand NAND2_5039 ( U7387 , EBX_REG_6_ , U7378 );
nand NAND2_5040 ( U7388 , INSTADDRPOINTER_REG_5_ , U7379 );
nand NAND2_5041 ( U7389 , EBX_REG_5_ , U7378 );
nand NAND2_5042 ( U7390 , INSTADDRPOINTER_REG_4_ , U7379 );
nand NAND2_5043 ( U7391 , EBX_REG_4_ , U7378 );
nand NAND2_5044 ( U7392 , INSTADDRPOINTER_REG_31_ , U7379 );
nand NAND2_5045 ( U7393 , EBX_REG_31_ , U7378 );
nand NAND2_5046 ( U7394 , INSTADDRPOINTER_REG_30_ , U7379 );
nand NAND2_5047 ( U7395 , EBX_REG_30_ , U7378 );
nand NAND2_5048 ( U7396 , INSTADDRPOINTER_REG_3_ , U7379 );
nand NAND2_5049 ( U7397 , EBX_REG_3_ , U7378 );
nand NAND2_5050 ( U7398 , INSTADDRPOINTER_REG_29_ , U7379 );
nand NAND2_5051 ( U7399 , EBX_REG_29_ , U7378 );
nand NAND2_5052 ( U7400 , INSTADDRPOINTER_REG_28_ , U7379 );
nand NAND2_5053 ( U7401 , EBX_REG_28_ , U7378 );
nand NAND2_5054 ( U7402 , INSTADDRPOINTER_REG_27_ , U7379 );
nand NAND2_5055 ( U7403 , EBX_REG_27_ , U7378 );
nand NAND2_5056 ( U7404 , INSTADDRPOINTER_REG_26_ , U7379 );
nand NAND2_5057 ( U7405 , EBX_REG_26_ , U7378 );
nand NAND2_5058 ( U7406 , INSTADDRPOINTER_REG_25_ , U7379 );
nand NAND2_5059 ( U7407 , EBX_REG_25_ , U7378 );
nand NAND2_5060 ( U7408 , INSTADDRPOINTER_REG_24_ , U7379 );
nand NAND2_5061 ( U7409 , EBX_REG_24_ , U7378 );
nand NAND2_5062 ( U7410 , INSTADDRPOINTER_REG_23_ , U7379 );
nand NAND2_5063 ( U7411 , EBX_REG_23_ , U7378 );
nand NAND2_5064 ( U7412 , INSTADDRPOINTER_REG_22_ , U7379 );
nand NAND2_5065 ( U7413 , EBX_REG_22_ , U7378 );
nand NAND2_5066 ( U7414 , INSTADDRPOINTER_REG_21_ , U7379 );
nand NAND2_5067 ( U7415 , EBX_REG_21_ , U7378 );
nand NAND2_5068 ( U7416 , INSTADDRPOINTER_REG_20_ , U7379 );
nand NAND2_5069 ( U7417 , EBX_REG_20_ , U7378 );
nand NAND2_5070 ( U7418 , INSTADDRPOINTER_REG_2_ , U7379 );
nand NAND2_5071 ( U7419 , EBX_REG_2_ , U7378 );
nand NAND2_5072 ( U7420 , INSTADDRPOINTER_REG_19_ , U7379 );
nand NAND2_5073 ( U7421 , EBX_REG_19_ , U7378 );
nand NAND2_5074 ( U7422 , INSTADDRPOINTER_REG_18_ , U7379 );
nand NAND2_5075 ( U7423 , EBX_REG_18_ , U7378 );
nand NAND2_5076 ( U7424 , INSTADDRPOINTER_REG_17_ , U7379 );
nand NAND2_5077 ( U7425 , EBX_REG_17_ , U7378 );
nand NAND2_5078 ( U7426 , INSTADDRPOINTER_REG_16_ , U7379 );
nand NAND2_5079 ( U7427 , EBX_REG_16_ , U7378 );
nand NAND2_5080 ( U7428 , INSTADDRPOINTER_REG_15_ , U7379 );
nand NAND2_5081 ( U7429 , EBX_REG_15_ , U7378 );
nand NAND2_5082 ( U7430 , INSTADDRPOINTER_REG_14_ , U7379 );
nand NAND2_5083 ( U7431 , EBX_REG_14_ , U7378 );
nand NAND2_5084 ( U7432 , INSTADDRPOINTER_REG_13_ , U7379 );
nand NAND2_5085 ( U7433 , EBX_REG_13_ , U7378 );
nand NAND2_5086 ( U7434 , INSTADDRPOINTER_REG_12_ , U7379 );
nand NAND2_5087 ( U7435 , EBX_REG_12_ , U7378 );
nand NAND2_5088 ( U7436 , INSTADDRPOINTER_REG_11_ , U7379 );
nand NAND2_5089 ( U7437 , EBX_REG_11_ , U7378 );
nand NAND2_5090 ( U7438 , INSTADDRPOINTER_REG_10_ , U7379 );
nand NAND2_5091 ( U7439 , EBX_REG_10_ , U7378 );
nand NAND2_5092 ( U7440 , INSTADDRPOINTER_REG_1_ , U7379 );
nand NAND2_5093 ( U7441 , EBX_REG_1_ , U7378 );
nand NAND2_5094 ( U7442 , INSTADDRPOINTER_REG_0_ , U7379 );
nand NAND2_5095 ( U7443 , EBX_REG_0_ , U7378 );
nand NAND2_5096 ( U7444 , U4465 , U4484 );
nand NAND2_5097 ( U7445 , U2430 , INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_5098 ( U7446 , U3476 , U3249 );
nand NAND2_5099 ( U7447 , U2430 , INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_5100 ( U7448 , U3477 , U3249 );
nand NAND3_5101 ( U7449 , FLUSH_REG , U2446 , U3457 );
nand NAND2_5102 ( U7450 , U2430 , INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_5103 ( U7451 , U3478 , U3249 );
nand NAND3_5104 ( U7452 , U2446 , FLUSH_REG , U7700 );
nand NAND2_5105 ( U7453 , U2430 , INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_5106 ( U7454 , U3479 , U3249 );
nand NAND2_5107 ( U7455 , U2430 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_5108 ( U7456 , STATE_REG_0_ , U4173 );
or OR2_5109 ( U7457 , READY_N , STATE2_REG_2_ );
nand NAND2_5110 ( U7458 , U4098 , U7206 );
nand NAND2_5111 ( U7459 , U7072 , U3409 );
nand NAND2_5112 ( U7460 , U4199 , STATE2_REG_0_ );
nand NAND2_5113 ( U7461 , U4200 , STATE2_REG_0_ );
nand NAND2_5114 ( U7462 , U4201 , STATE2_REG_0_ );
nand NAND2_5115 ( U7463 , U4224 , STATE2_REG_0_ );
nand NAND2_5116 ( U7464 , U4252 , STATE2_REG_0_ );
nand NAND2_5117 ( U7465 , STATE2_REG_0_ , U7620 );
nand NAND2_5118 ( U7466 , U2608 , U3253 );
nand NAND4_5119 ( U7467 , U4105 , U7081 , U4106 , U4108 );
nand NAND2_5120 ( U7468 , STATE2_REG_0_ , U7620 );
nand NAND2_5121 ( U7469 , U2379 , U3416 );
nand NAND2_5122 ( U7470 , U2369 , U6355 );
nand NAND2_5123 ( U7471 , U3876 , U2369 );
nand NAND3_5124 ( U7472 , U7469 , U4217 , U7470 );
nand NAND2_5125 ( U7473 , U7471 , U4218 );
nand NAND3_5126 ( U7474 , U5479 , U4159 , U4182 );
nand NAND2_5127 ( U7475 , U7079 , U4182 );
nand NAND2_5128 ( U7476 , U4182 , U3379 );
nand NAND2_5129 ( U7477 , U4224 , STATE2_REG_0_ );
nand NAND3_5130 ( U7478 , U7773 , U7772 , U4060 );
nand NAND2_5131 ( U7479 , U4096 , U7204 );
nand NAND2_5132 ( U7480 , U4097 , U7082 );
not NOT1_5133 ( U7481 , U3266 );
not NOT1_5134 ( U7482 , U3263 );
nand NAND5_5135 ( U7483 , U4059 , U2607 , U4058 , U4057 , U4056 );
nand NAND2_5136 ( U7484 , U3722 , U7481 );
nand NAND2_5137 ( U7485 , U3723 , U5457 );
nand NAND2_5138 ( U7486 , U2425 , U7481 );
nand NAND2_5139 ( U7487 , U2425 , U7481 );
nand NAND3_5140 ( U7488 , U6349 , U6348 , U7487 );
nand NAND2_5141 ( U7489 , U7481 , R2167_U17 );
nand NAND3_5142 ( U7490 , U7481 , U4189 , R2167_U17 );
nand NAND2_5143 ( U7491 , U7490 , U6137 );
nand NAND2_5144 ( U7492 , U7481 , U7073 );
nand NAND2_5145 ( U7493 , U7481 , U7459 );
nand NAND3_5146 ( U7494 , U4104 , U4103 , U4102 );
nand NAND2_5147 ( U7495 , U3747 , U7481 );
nand NAND3_5148 ( U7496 , U3749 , U5553 , U3748 );
nand NAND2_5149 ( U7497 , U3734 , U2519 );
nand NAND2_5150 ( U7498 , U7481 , U5950 );
nand NAND2_5151 ( U7499 , U7481 , U5953 );
nand NAND2_5152 ( U7500 , U7481 , U5956 );
nand NAND2_5153 ( U7501 , U7481 , U5959 );
nand NAND2_5154 ( U7502 , U7481 , U5962 );
nand NAND2_5155 ( U7503 , U7481 , U5965 );
nand NAND2_5156 ( U7504 , U7481 , U5968 );
nand NAND2_5157 ( U7505 , U7481 , U5971 );
nand NAND2_5158 ( U7506 , U7481 , U5974 );
nand NAND2_5159 ( U7507 , U7481 , U5977 );
nand NAND2_5160 ( U7508 , U7481 , U5980 );
nand NAND2_5161 ( U7509 , U7481 , U5983 );
nand NAND2_5162 ( U7510 , U7481 , U5986 );
nand NAND2_5163 ( U7511 , U7481 , U5989 );
nand NAND2_5164 ( U7512 , U7481 , U5992 );
nand NAND2_5165 ( U7513 , U7481 , U5995 );
nand NAND2_5166 ( U7514 , U7481 , U5998 );
nand NAND2_5167 ( U7515 , U7481 , U6001 );
nand NAND2_5168 ( U7516 , U7481 , U6004 );
nand NAND2_5169 ( U7517 , U7481 , U6007 );
nand NAND2_5170 ( U7518 , U7481 , U6010 );
nand NAND2_5171 ( U7519 , U7481 , U6013 );
nand NAND2_5172 ( U7520 , U7481 , U6016 );
nand NAND2_5173 ( U7521 , U7481 , U6019 );
nand NAND2_5174 ( U7522 , U7481 , U6022 );
nand NAND2_5175 ( U7523 , U7481 , U6025 );
nand NAND2_5176 ( U7524 , U7481 , U6028 );
nand NAND2_5177 ( U7525 , U7481 , U6031 );
nand NAND2_5178 ( U7526 , U7481 , U6034 );
nand NAND2_5179 ( U7527 , U7481 , U6037 );
nand NAND2_5180 ( U7528 , U7481 , U6040 );
nand NAND2_5181 ( U7529 , U2357 , U7481 );
nand NAND2_5182 ( U7530 , UWORD_REG_0_ , U7529 );
nand NAND2_5183 ( U7531 , U2357 , U7481 );
nand NAND2_5184 ( U7532 , UWORD_REG_1_ , U7531 );
nand NAND2_5185 ( U7533 , U2357 , U7481 );
nand NAND2_5186 ( U7534 , UWORD_REG_2_ , U7533 );
nand NAND2_5187 ( U7535 , U2357 , U7481 );
nand NAND2_5188 ( U7536 , UWORD_REG_3_ , U7535 );
nand NAND2_5189 ( U7537 , U2357 , U7481 );
nand NAND2_5190 ( U7538 , UWORD_REG_4_ , U7537 );
nand NAND2_5191 ( U7539 , U2357 , U7481 );
nand NAND2_5192 ( U7540 , UWORD_REG_5_ , U7539 );
nand NAND2_5193 ( U7541 , U2357 , U7481 );
nand NAND2_5194 ( U7542 , UWORD_REG_6_ , U7541 );
nand NAND2_5195 ( U7543 , U2357 , U7481 );
nand NAND2_5196 ( U7544 , UWORD_REG_7_ , U7543 );
nand NAND2_5197 ( U7545 , U2357 , U7481 );
nand NAND2_5198 ( U7546 , UWORD_REG_8_ , U7545 );
nand NAND2_5199 ( U7547 , U2357 , U7481 );
nand NAND2_5200 ( U7548 , UWORD_REG_9_ , U7547 );
nand NAND2_5201 ( U7549 , U2357 , U7481 );
nand NAND2_5202 ( U7550 , UWORD_REG_10_ , U7549 );
nand NAND2_5203 ( U7551 , U2357 , U7481 );
nand NAND2_5204 ( U7552 , UWORD_REG_11_ , U7551 );
nand NAND2_5205 ( U7553 , U2357 , U7481 );
nand NAND2_5206 ( U7554 , UWORD_REG_12_ , U7553 );
nand NAND2_5207 ( U7555 , U2357 , U7481 );
nand NAND2_5208 ( U7556 , UWORD_REG_13_ , U7555 );
nand NAND2_5209 ( U7557 , U2357 , U7481 );
nand NAND2_5210 ( U7558 , UWORD_REG_14_ , U7557 );
nand NAND2_5211 ( U7559 , U2357 , U7481 );
nand NAND2_5212 ( U7560 , LWORD_REG_0_ , U7559 );
nand NAND2_5213 ( U7561 , U2357 , U7481 );
nand NAND2_5214 ( U7562 , LWORD_REG_1_ , U7561 );
nand NAND2_5215 ( U7563 , U2357 , U7481 );
nand NAND2_5216 ( U7564 , LWORD_REG_2_ , U7563 );
nand NAND2_5217 ( U7565 , U2357 , U7481 );
nand NAND2_5218 ( U7566 , LWORD_REG_3_ , U7565 );
nand NAND2_5219 ( U7567 , U2357 , U7481 );
nand NAND2_5220 ( U7568 , LWORD_REG_4_ , U7567 );
nand NAND2_5221 ( U7569 , U2357 , U7481 );
nand NAND2_5222 ( U7570 , LWORD_REG_5_ , U7569 );
nand NAND2_5223 ( U7571 , U2357 , U7481 );
nand NAND2_5224 ( U7572 , LWORD_REG_6_ , U7571 );
nand NAND2_5225 ( U7573 , U2357 , U7481 );
nand NAND2_5226 ( U7574 , LWORD_REG_7_ , U7573 );
nand NAND2_5227 ( U7575 , U2357 , U7481 );
nand NAND2_5228 ( U7576 , LWORD_REG_8_ , U7575 );
nand NAND2_5229 ( U7577 , U2357 , U7481 );
nand NAND2_5230 ( U7578 , LWORD_REG_9_ , U7577 );
nand NAND2_5231 ( U7579 , U2357 , U7481 );
nand NAND2_5232 ( U7580 , LWORD_REG_10_ , U7579 );
nand NAND2_5233 ( U7581 , U2357 , U7481 );
nand NAND2_5234 ( U7582 , LWORD_REG_11_ , U7581 );
nand NAND2_5235 ( U7583 , U2357 , U7481 );
nand NAND2_5236 ( U7584 , LWORD_REG_12_ , U7583 );
nand NAND2_5237 ( U7585 , U2357 , U7481 );
nand NAND2_5238 ( U7586 , LWORD_REG_13_ , U7585 );
nand NAND2_5239 ( U7587 , U2357 , U7481 );
nand NAND2_5240 ( U7588 , LWORD_REG_14_ , U7587 );
nand NAND2_5241 ( U7589 , U2357 , U7481 );
nand NAND2_5242 ( U7590 , LWORD_REG_15_ , U7589 );
nand NAND3_5243 ( U7591 , U7481 , U3556 , U4247 );
nand NAND3_5244 ( U7592 , U7672 , U7671 , U3569 );
nand NAND2_5245 ( U7593 , U3855 , U7481 );
nand NAND2_5246 ( U7594 , U7593 , U3415 );
nand NAND2_5247 ( U7595 , U4196 , U7481 );
nand NAND2_5248 ( U7596 , U7595 , U3434 );
nand NAND2_5249 ( U7597 , U3266 , U3387 );
nand NAND2_5250 ( U7598 , U3742 , U7481 );
nand NAND2_5251 ( U7599 , U3743 , U7598 );
nand NAND2_5252 ( U7600 , INSTQUEUE_REG_0__4_ , U5404 );
nand NAND2_5253 ( U7601 , U2523 , INSTQUEUE_REG_0__4_ );
nand NAND2_5254 ( U7602 , U2546 , INSTQUEUE_REG_0__4_ );
nand NAND4_5255 ( U7603 , U4040 , U4039 , U4038 , U4037 );
nand NAND2_5256 ( U7604 , U4180 , INSTQUEUE_REG_0__4_ );
nand NAND2_5257 ( U7605 , U2573 , INSTQUEUE_REG_0__4_ );
nand NAND4_5258 ( U7606 , U4079 , U4077 , U4076 , U4075 );
nand NAND2_5259 ( U7607 , U2592 , INSTQUEUE_REG_0__4_ );
nand NAND4_5260 ( U7608 , U4124 , U4123 , U4122 , U4121 );
not NOT1_5261 ( U7609 , U3246 );
nand NAND2_5262 ( U7610 , U7609 , U3248 );
nand NAND3_5263 ( U7611 , U4349 , STATE_REG_1_ , U4346 );
nand NAND2_5264 ( U7612 , STATE_REG_2_ , U7456 );
nand NAND2_5265 ( U7613 , STATE_REG_1_ , U4346 );
nand NAND2_5266 ( U7614 , U4490 , U4498 );
nand NAND2_5267 ( U7615 , U5475 , U4159 );
nand NAND2_5268 ( U7616 , U3270 , U3276 );
not NOT1_5269 ( U7617 , U3379 );
nand NAND2_5270 ( U7618 , U4196 , U7478 );
nand NAND2_5271 ( U7619 , U5475 , U4159 );
nand NAND2_5272 ( U7620 , U7619 , U7618 );
nand NAND2_5273 ( U7621 , BE_N_REG_3_ , U3236 );
nand NAND2_5274 ( U7622 , BYTEENABLE_REG_3_ , U4209 );
nand NAND2_5275 ( U7623 , BE_N_REG_2_ , U3236 );
nand NAND2_5276 ( U7624 , BYTEENABLE_REG_2_ , U4209 );
nand NAND2_5277 ( U7625 , BE_N_REG_1_ , U3236 );
nand NAND2_5278 ( U7626 , BYTEENABLE_REG_1_ , U4209 );
nand NAND2_5279 ( U7627 , BE_N_REG_0_ , U3236 );
nand NAND2_5280 ( U7628 , BYTEENABLE_REG_0_ , U4209 );
nand NAND3_5281 ( U7629 , STATE_REG_0_ , REQUESTPENDING_REG , U3238 );
nand NAND2_5282 ( U7630 , STATE_REG_2_ , U3246 );
nand NAND2_5283 ( U7631 , U7630 , U7629 );
nand NAND3_5284 ( U7632 , U7612 , U4349 , STATE_REG_1_ );
nand NAND2_5285 ( U7633 , U7631 , U3235 );
nand NAND3_5286 ( U7634 , STATE_REG_0_ , U3247 , STATE_REG_2_ );
nand NAND2_5287 ( U7635 , U4359 , U3238 );
or OR2_5288 ( U7636 , STATE_REG_0_ , STATE_REG_1_ );
nand NAND2_5289 ( U7637 , STATE_REG_0_ , U4246 );
not NOT1_5290 ( U7638 , U3449 );
nand NAND2_5291 ( U7639 , U7638 , DATAWIDTH_REG_0_ );
nand NAND2_5292 ( U7640 , U3450 , U3449 );
nand NAND2_5293 ( U7641 , U3449 , U4364 );
nand NAND2_5294 ( U7642 , U7638 , DATAWIDTH_REG_1_ );
nand NAND3_5295 ( U7643 , U3529 , U3528 , U3252 );
nand NAND5_5296 ( U7644 , INSTQUEUE_REG_7__4_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_2_ , U3257 , INSTQUEUERD_ADDR_REG_1_ );
nand NAND5_5297 ( U7645 , INSTQUEUE_REG_5__4_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_2_ , U3257 , U3252 );
nand NAND5_5298 ( U7646 , INSTQUEUE_REG_2__4_ , U3257 , U3251 , U3253 , INSTQUEUERD_ADDR_REG_1_ );
nand NAND3_5299 ( U7647 , U3531 , U3530 , U3257 );
nand NAND3_5300 ( U7648 , U3533 , U3532 , INSTQUEUERD_ADDR_REG_3_ );
nand NAND3_5301 ( U7649 , U3535 , U3534 , U3252 );
nand NAND3_5302 ( U7650 , U3537 , U3536 , INSTQUEUERD_ADDR_REG_1_ );
nand NAND3_5303 ( U7651 , U3539 , U3538 , U3253 );
nand NAND5_5304 ( U7652 , INSTQUEUE_REG_15__4_ , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_1_ , INSTQUEUERD_ADDR_REG_2_ , INSTQUEUERD_ADDR_REG_0_ );
nand NAND5_5305 ( U7653 , INSTQUEUE_REG_0__4_ , U3251 , U3252 , U3253 , U3257 );
nand NAND5_5306 ( U7654 , INSTQUEUE_REG_8__4_ , U3251 , U3252 , U3253 , INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_5307 ( U7655 , INSTQUEUE_REG_10__4_ , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_1_ , U3251 , U3253 );
nand NAND3_5308 ( U7656 , U3541 , U3540 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND5_5309 ( U7657 , INSTQUEUE_REG_3__4_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ , U3251 , U3257 );
nand NAND5_5310 ( U7658 , INSTQUEUE_REG_11__4_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ , U3251 , INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_5311 ( U7659 , INSTQUEUE_REG_3__5_ , INSTQUEUERD_ADDR_REG_0_ , INSTQUEUERD_ADDR_REG_1_ , U3251 , U3257 );
nand NAND3_5312 ( U7660 , U3517 , U3516 , INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_5313 ( U7661 , INSTQUEUE_REG_9__6_ , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_0_ , U3251 , U3252 );
nand NAND3_5314 ( U7662 , U3523 , U3522 , INSTQUEUERD_ADDR_REG_1_ );
nand NAND5_5315 ( U7663 , INSTQUEUE_REG_10__6_ , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_1_ , U3251 , U3253 );
nand NAND5_5316 ( U7664 , INSTQUEUE_REG_11__6_ , INSTQUEUERD_ADDR_REG_3_ , INSTQUEUERD_ADDR_REG_1_ , U3251 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND5_5317 ( U7665 , INSTQUEUE_REG_0__6_ , U3251 , U3252 , U3253 , U3257 );
nand NAND5_5318 ( U7666 , INSTQUEUE_REG_8__6_ , U3251 , U3252 , U3253 , INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_5319 ( U7667 , U4482 , U3424 );
nand NAND2_5320 ( U7668 , U7489 , U3271 );
nand NAND2_5321 ( U7669 , U4204 , R2167_U17 );
nand NAND2_5322 ( U7670 , U4494 , U3260 );
nand NAND2_5323 ( U7671 , STATE2_REG_0_ , U4500 );
nand NAND2_5324 ( U7672 , U4501 , U3281 );
nand NAND2_5325 ( U7673 , STATE2_REG_3_ , U3282 );
nand NAND2_5326 ( U7674 , U2428 , U4502 );
or OR2_5327 ( U7675 , STATEBS16_REG , STATE2_REG_0_ );
nand NAND2_5328 ( U7676 , STATE2_REG_0_ , U7457 );
nand NAND2_5329 ( U7677 , STATE2_REG_0_ , U4510 );
nand NAND3_5330 ( U7678 , U7592 , U4509 , U3281 );
nand NAND2_5331 ( U7679 , R2144_U49 , U3300 );
nand NAND2_5332 ( U7680 , U4516 , U3298 );
not NOT1_5333 ( U7681 , U3441 );
nand NAND2_5334 ( U7682 , INSTQUEUEWR_ADDR_REG_2_ , U3292 );
nand NAND2_5335 ( U7683 , U4521 , U3291 );
not NOT1_5336 ( U7684 , U3442 );
nand NAND2_5337 ( U7685 , U4204 , U3260 );
nand NAND2_5338 ( U7686 , R2167_U17 , U7485 );
nand NAND2_5339 ( U7687 , U4420 , U5454 );
nand NAND2_5340 ( U7688 , U5455 , U4159 );
nand NAND2_5341 ( U7689 , U3454 , U4160 );
nand NAND2_5342 ( U7690 , U5464 , INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_5343 ( U7691 , U4448 , U3265 );
nand NAND2_5344 ( U7692 , U4403 , U3264 );
nand NAND2_5345 ( U7693 , U3258 , U3402 );
nand NAND2_5346 ( U7694 , U4465 , U5481 );
nand NAND2_5347 ( U7695 , U7694 , U7693 );
nand NAND2_5348 ( U7696 , U5464 , INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_5349 ( U7697 , U5497 , U4160 );
nand NAND2_5350 ( U7698 , INSTADDRPOINTER_REG_1_ , U4162 );
nand NAND2_5351 ( U7699 , SUB_580_U6 , INSTADDRPOINTER_REG_31_ );
not NOT1_5352 ( U7700 , U3457 );
nand NAND2_5353 ( U7701 , INSTADDRPOINTER_REG_0_ , U4162 );
nand NAND2_5354 ( U7702 , INSTADDRPOINTER_REG_0_ , INSTADDRPOINTER_REG_31_ );
not NOT1_5355 ( U7703 , U3458 );
nand NAND2_5356 ( U7704 , U5499 , U5489 );
nand NAND2_5357 ( U7705 , U4206 , U3388 );
nand NAND2_5358 ( U7706 , INSTQUEUERD_ADDR_REG_1_ , U3251 );
nand NAND2_5359 ( U7707 , INSTQUEUERD_ADDR_REG_2_ , U3252 );
not NOT1_5360 ( U7708 , U3443 );
nand NAND2_5361 ( U7709 , U5464 , INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_5362 ( U7710 , U5506 , U4160 );
nand NAND2_5363 ( U7711 , U5464 , INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_5364 ( U7712 , U5517 , U4160 );
nand NAND2_5365 ( U7713 , U4202 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_5366 ( U7714 , U5509 , U3253 );
nand NAND2_5367 ( U7715 , U5464 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_5368 ( U7716 , U5523 , U4160 );
nand NAND2_5369 ( U7717 , U5525 , INSTQUEUEWR_ADDR_REG_3_ );
nand NAND2_5370 ( U7718 , U5533 , U3391 );
nand NAND2_5371 ( U7719 , U7681 , U4515 );
nand NAND2_5372 ( U7720 , U3441 , U3301 );
nand NAND2_5373 ( U7721 , U7720 , U7719 );
nand NAND2_5374 ( U7722 , U5525 , INSTQUEUEWR_ADDR_REG_2_ );
nand NAND2_5375 ( U7723 , U5537 , U3391 );
nand NAND2_5376 ( U7724 , U5525 , INSTQUEUEWR_ADDR_REG_1_ );
nand NAND2_5377 ( U7725 , U5542 , U3391 );
nand NAND2_5378 ( U7726 , U5525 , INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_5379 ( U7727 , U5545 , U3391 );
nand NAND2_5380 ( U7728 , U4465 , U3375 );
nand NAND2_5381 ( U7729 , U3258 , U3268 );
nand NAND4_5382 ( U7730 , U7729 , U7728 , U3244 , U4159 );
nand NAND3_5383 ( U7731 , R2167_U17 , U7599 , U4420 );
nand NAND2_5384 ( U7732 , EAX_REG_31_ , U3411 );
nand NAND2_5385 ( U7733 , U3466 , U4211 );
nand NAND2_5386 ( U7734 , BYTEENABLE_REG_3_ , U3420 );
nand NAND2_5387 ( U7735 , U3467 , U4208 );
or OR2_5388 ( U7736 , DATAWIDTH_REG_0_ , DATAWIDTH_REG_1_ );
nand NAND2_5389 ( U7737 , DATAWIDTH_REG_0_ , U3400 );
nand NAND2_5390 ( U7738 , U7737 , U7736 );
nand NAND2_5391 ( U7739 , U7738 , U3240 );
nand NAND2_5392 ( U7740 , REIP_REG_0_ , REIP_REG_1_ );
nand NAND2_5393 ( U7741 , U7740 , U7739 );
nand NAND2_5394 ( U7742 , BYTEENABLE_REG_2_ , U3420 );
nand NAND2_5395 ( U7743 , U7741 , U4208 );
nand NAND2_5396 ( U7744 , BYTEENABLE_REG_1_ , U3420 );
nand NAND2_5397 ( U7745 , U4208 , REIP_REG_1_ );
nand NAND2_5398 ( U7746 , BYTEENABLE_REG_0_ , U3420 );
nand NAND2_5399 ( U7747 , U4208 , U6587 );
nand NAND2_5400 ( U7748 , U4209 , U3423 );
nand NAND2_5401 ( U7749 , W_R_N_REG , U3236 );
nand NAND2_5402 ( U7750 , MORE_REG , U4165 );
nand NAND2_5403 ( U7751 , U4225 , U6588 );
nand NAND2_5404 ( U7752 , U7638 , STATEBS16_REG );
nand NAND2_5405 ( U7753 , BS16_N , U3449 );
nand NAND2_5406 ( U7754 , U6591 , REQUESTPENDING_REG );
nand NAND2_5407 ( U7755 , U6597 , U4168 );
nand NAND2_5408 ( U7756 , U4209 , U3422 );
nand NAND2_5409 ( U7757 , D_C_N_REG , U3236 );
nand NAND2_5410 ( U7758 , M_IO_N_REG , U3236 );
nand NAND2_5411 ( U7759 , MEMORYFETCH_REG , U4209 );
nand NAND2_5412 ( U7760 , U6602 , READREQUEST_REG );
nand NAND2_5413 ( U7761 , U6603 , U4169 );
nand NAND2_5414 ( U7762 , U3475 , U4170 );
nand NAND2_5415 ( U7763 , U5461 , INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_5416 ( U7764 , U5461 , INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_5417 ( U7765 , U5494 , U4170 );
nand NAND2_5418 ( U7766 , U5461 , INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_5419 ( U7767 , U5502 , U4170 );
nand NAND2_5420 ( U7768 , U5461 , INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_5421 ( U7769 , U5513 , U4170 );
nand NAND2_5422 ( U7770 , U5461 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_5423 ( U7771 , U5519 , U4170 );
nand NAND2_5424 ( U7772 , U2605 , U3264 );
nand NAND2_5425 ( U7773 , U4448 , U7483 );
nand NAND2_5426 ( U7774 , U4191 , U3288 );
nand NAND2_5427 ( U7775 , INSTQUEUEWR_ADDR_REG_0_ , U3284 );
nand NAND2_5428 ( U7776 , INSTQUEUERD_ADDR_REG_3_ , U4171 );
nand NAND2_5429 ( U7777 , U7207 , U3257 );
not NOT1_5430 ( U7778 , U3444 );
nand NAND2_5431 ( U7779 , U3263 , U3271 );
nand NAND2_5432 ( U7780 , U7695 , U4482 );
nand NAND2_5433 ( U7781 , U3480 , U3249 );
nand NAND3_5434 ( U7782 , FLUSH_REG , U7703 , STATE2_REG_1_ );
nand NAND2_5435 ( ADD_515_U178 , ADD_515_U103 , ADD_515_U25 );
nand NAND2_5436 ( ADD_515_U177 , INSTADDRPOINTER_REG_12_ , ADD_515_U24 );
nand NAND2_5437 ( ADD_515_U176 , ADD_515_U104 , ADD_515_U27 );
nand NAND2_5438 ( ADD_515_U175 , INSTADDRPOINTER_REG_13_ , ADD_515_U26 );
nand NAND2_5439 ( ADD_515_U174 , ADD_515_U105 , ADD_515_U29 );
nand NAND2_5440 ( ADD_515_U173 , INSTADDRPOINTER_REG_14_ , ADD_515_U28 );
nand NAND2_5441 ( ADD_515_U172 , ADD_515_U106 , ADD_515_U31 );
nand NAND2_5442 ( ADD_515_U171 , INSTADDRPOINTER_REG_15_ , ADD_515_U30 );
nand NAND2_5443 ( ADD_515_U170 , ADD_515_U107 , ADD_515_U33 );
nand NAND2_5444 ( ADD_515_U169 , INSTADDRPOINTER_REG_16_ , ADD_515_U32 );
nand NAND2_5445 ( ADD_515_U168 , ADD_515_U108 , ADD_515_U35 );
nand NAND2_5446 ( ADD_515_U167 , INSTADDRPOINTER_REG_17_ , ADD_515_U34 );
nand NAND2_5447 ( ADD_515_U166 , ADD_515_U109 , ADD_515_U37 );
nand NAND2_5448 ( ADD_515_U165 , INSTADDRPOINTER_REG_18_ , ADD_515_U36 );
nand NAND2_5449 ( ADD_515_U164 , ADD_515_U110 , ADD_515_U39 );
nand NAND2_5450 ( ADD_515_U163 , INSTADDRPOINTER_REG_19_ , ADD_515_U38 );
nand NAND2_5451 ( ADD_515_U162 , ADD_515_U111 , ADD_515_U41 );
nand NAND2_5452 ( ADD_515_U161 , INSTADDRPOINTER_REG_20_ , ADD_515_U40 );
nand NAND2_5453 ( ADD_515_U160 , ADD_515_U112 , ADD_515_U43 );
nand NAND2_5454 ( ADD_515_U159 , INSTADDRPOINTER_REG_21_ , ADD_515_U42 );
nand NAND2_5455 ( ADD_515_U158 , ADD_515_U113 , ADD_515_U45 );
nand NAND2_5456 ( ADD_515_U157 , INSTADDRPOINTER_REG_22_ , ADD_515_U44 );
nand NAND2_5457 ( ADD_515_U156 , ADD_515_U114 , ADD_515_U47 );
nand NAND2_5458 ( ADD_515_U155 , INSTADDRPOINTER_REG_23_ , ADD_515_U46 );
nand NAND2_5459 ( ADD_515_U154 , ADD_515_U115 , ADD_515_U49 );
nand NAND2_5460 ( ADD_515_U153 , INSTADDRPOINTER_REG_24_ , ADD_515_U48 );
nand NAND2_5461 ( ADD_515_U152 , ADD_515_U116 , ADD_515_U51 );
not NOT1_5462 ( R2027_U5 , INSTADDRPOINTER_REG_0_ );
not NOT1_5463 ( R2027_U6 , INSTADDRPOINTER_REG_2_ );
not NOT1_5464 ( R2027_U7 , INSTADDRPOINTER_REG_1_ );
not NOT1_5465 ( R2027_U8 , INSTADDRPOINTER_REG_4_ );
not NOT1_5466 ( R2027_U9 , INSTADDRPOINTER_REG_3_ );
nand NAND3_5467 ( R2027_U10 , INSTADDRPOINTER_REG_2_ , INSTADDRPOINTER_REG_0_ , INSTADDRPOINTER_REG_1_ );
not NOT1_5468 ( R2027_U11 , INSTADDRPOINTER_REG_6_ );
not NOT1_5469 ( R2027_U12 , INSTADDRPOINTER_REG_5_ );
nand NAND2_5470 ( R2027_U13 , R2027_U82 , R2027_U111 );
not NOT1_5471 ( R2027_U14 , INSTADDRPOINTER_REG_8_ );
not NOT1_5472 ( R2027_U15 , INSTADDRPOINTER_REG_7_ );
nand NAND2_5473 ( R2027_U16 , R2027_U83 , R2027_U112 );
nand NAND2_5474 ( R2027_U17 , R2027_U84 , R2027_U118 );
not NOT1_5475 ( R2027_U18 , INSTADDRPOINTER_REG_9_ );
not NOT1_5476 ( R2027_U19 , INSTADDRPOINTER_REG_10_ );
not NOT1_5477 ( R2027_U20 , INSTADDRPOINTER_REG_12_ );
not NOT1_5478 ( R2027_U21 , INSTADDRPOINTER_REG_11_ );
nand NAND2_5479 ( R2027_U22 , R2027_U85 , R2027_U120 );
not NOT1_5480 ( R2027_U23 , INSTADDRPOINTER_REG_14_ );
not NOT1_5481 ( R2027_U24 , INSTADDRPOINTER_REG_13_ );
nand NAND2_5482 ( R2027_U25 , R2027_U86 , R2027_U113 );
not NOT1_5483 ( R2027_U26 , INSTADDRPOINTER_REG_15_ );
nand NAND2_5484 ( R2027_U27 , R2027_U87 , R2027_U119 );
not NOT1_5485 ( R2027_U28 , INSTADDRPOINTER_REG_16_ );
not NOT1_5486 ( R2027_U29 , INSTADDRPOINTER_REG_18_ );
not NOT1_5487 ( R2027_U30 , INSTADDRPOINTER_REG_17_ );
nand NAND2_5488 ( R2027_U31 , R2027_U88 , R2027_U124 );
not NOT1_5489 ( R2027_U32 , INSTADDRPOINTER_REG_20_ );
not NOT1_5490 ( R2027_U33 , INSTADDRPOINTER_REG_19_ );
nand NAND2_5491 ( R2027_U34 , R2027_U89 , R2027_U117 );
not NOT1_5492 ( R2027_U35 , INSTADDRPOINTER_REG_21_ );
nand NAND2_5493 ( R2027_U36 , R2027_U90 , R2027_U114 );
not NOT1_5494 ( R2027_U37 , INSTADDRPOINTER_REG_22_ );
not NOT1_5495 ( R2027_U38 , INSTADDRPOINTER_REG_24_ );
not NOT1_5496 ( R2027_U39 , INSTADDRPOINTER_REG_23_ );
nand NAND2_5497 ( R2027_U40 , R2027_U91 , R2027_U121 );
not NOT1_5498 ( R2027_U41 , INSTADDRPOINTER_REG_26_ );
not NOT1_5499 ( R2027_U42 , INSTADDRPOINTER_REG_25_ );
nand NAND2_5500 ( R2027_U43 , R2027_U92 , R2027_U115 );
not NOT1_5501 ( R2027_U44 , INSTADDRPOINTER_REG_27_ );
not NOT1_5502 ( R2027_U45 , INSTADDRPOINTER_REG_28_ );
nand NAND2_5503 ( R2027_U46 , R2027_U93 , R2027_U116 );
not NOT1_5504 ( R2027_U47 , INSTADDRPOINTER_REG_29_ );
nand NAND2_5505 ( R2027_U48 , R2027_U94 , R2027_U122 );
nand NAND2_5506 ( R2027_U49 , R2027_U123 , INSTADDRPOINTER_REG_29_ );
not NOT1_5507 ( R2027_U50 , INSTADDRPOINTER_REG_30_ );
nand NAND2_5508 ( R2027_U51 , R2027_U142 , R2027_U141 );
nand NAND2_5509 ( R2027_U52 , R2027_U144 , R2027_U143 );
nand NAND2_5510 ( R2027_U53 , R2027_U146 , R2027_U145 );
nand NAND2_5511 ( R2027_U54 , R2027_U148 , R2027_U147 );
nand NAND2_5512 ( R2027_U55 , R2027_U150 , R2027_U149 );
nand NAND2_5513 ( R2027_U56 , R2027_U152 , R2027_U151 );
nand NAND2_5514 ( R2027_U57 , R2027_U154 , R2027_U153 );
nand NAND2_5515 ( R2027_U58 , R2027_U156 , R2027_U155 );
nand NAND2_5516 ( R2027_U59 , R2027_U158 , R2027_U157 );
nand NAND2_5517 ( R2027_U60 , R2027_U160 , R2027_U159 );
nand NAND2_5518 ( R2027_U61 , R2027_U162 , R2027_U161 );
nand NAND2_5519 ( R2027_U62 , R2027_U164 , R2027_U163 );
nand NAND2_5520 ( R2027_U63 , R2027_U166 , R2027_U165 );
nand NAND2_5521 ( R2027_U64 , R2027_U168 , R2027_U167 );
nand NAND2_5522 ( R2027_U65 , R2027_U170 , R2027_U169 );
nand NAND2_5523 ( R2027_U66 , R2027_U172 , R2027_U171 );
nand NAND2_5524 ( R2027_U67 , R2027_U174 , R2027_U173 );
nand NAND2_5525 ( R2027_U68 , R2027_U176 , R2027_U175 );
nand NAND2_5526 ( R2027_U69 , R2027_U178 , R2027_U177 );
nand NAND2_5527 ( R2027_U70 , R2027_U180 , R2027_U179 );
nand NAND2_5528 ( R2027_U71 , R2027_U182 , R2027_U181 );
nand NAND2_5529 ( R2027_U72 , R2027_U184 , R2027_U183 );
nand NAND2_5530 ( R2027_U73 , R2027_U186 , R2027_U185 );
nand NAND2_5531 ( R2027_U74 , R2027_U188 , R2027_U187 );
nand NAND2_5532 ( R2027_U75 , R2027_U190 , R2027_U189 );
nand NAND2_5533 ( R2027_U76 , R2027_U192 , R2027_U191 );
nand NAND2_5534 ( R2027_U77 , R2027_U194 , R2027_U193 );
nand NAND2_5535 ( R2027_U78 , R2027_U196 , R2027_U195 );
nand NAND2_5536 ( R2027_U79 , R2027_U198 , R2027_U197 );
nand NAND2_5537 ( R2027_U80 , R2027_U200 , R2027_U199 );
nand NAND2_5538 ( R2027_U81 , R2027_U202 , R2027_U201 );
and AND2_5539 ( R2027_U82 , INSTADDRPOINTER_REG_3_ , INSTADDRPOINTER_REG_4_ );
and AND2_5540 ( R2027_U83 , INSTADDRPOINTER_REG_5_ , INSTADDRPOINTER_REG_6_ );
and AND2_5541 ( R2027_U84 , INSTADDRPOINTER_REG_7_ , INSTADDRPOINTER_REG_8_ );
and AND2_5542 ( R2027_U85 , INSTADDRPOINTER_REG_9_ , INSTADDRPOINTER_REG_10_ );
and AND2_5543 ( R2027_U86 , INSTADDRPOINTER_REG_11_ , INSTADDRPOINTER_REG_12_ );
and AND2_5544 ( R2027_U87 , INSTADDRPOINTER_REG_13_ , INSTADDRPOINTER_REG_14_ );
and AND2_5545 ( R2027_U88 , INSTADDRPOINTER_REG_16_ , INSTADDRPOINTER_REG_15_ );
and AND2_5546 ( R2027_U89 , INSTADDRPOINTER_REG_17_ , INSTADDRPOINTER_REG_18_ );
and AND2_5547 ( R2027_U90 , INSTADDRPOINTER_REG_19_ , INSTADDRPOINTER_REG_20_ );
and AND2_5548 ( R2027_U91 , INSTADDRPOINTER_REG_22_ , INSTADDRPOINTER_REG_21_ );
and AND2_5549 ( R2027_U92 , INSTADDRPOINTER_REG_23_ , INSTADDRPOINTER_REG_24_ );
and AND2_5550 ( R2027_U93 , INSTADDRPOINTER_REG_25_ , INSTADDRPOINTER_REG_26_ );
and AND2_5551 ( R2027_U94 , INSTADDRPOINTER_REG_28_ , INSTADDRPOINTER_REG_27_ );
nand NAND2_5552 ( R2027_U95 , R2027_U118 , INSTADDRPOINTER_REG_7_ );
nand NAND2_5553 ( R2027_U96 , R2027_U112 , INSTADDRPOINTER_REG_5_ );
nand NAND2_5554 ( R2027_U97 , R2027_U111 , INSTADDRPOINTER_REG_3_ );
not NOT1_5555 ( R2027_U98 , INSTADDRPOINTER_REG_31_ );
nand NAND2_5556 ( R2027_U99 , INSTADDRPOINTER_REG_30_ , R2027_U128 );
nand NAND2_5557 ( R2027_U100 , INSTADDRPOINTER_REG_1_ , INSTADDRPOINTER_REG_0_ );
nand NAND2_5558 ( R2027_U101 , R2027_U122 , INSTADDRPOINTER_REG_27_ );
nand NAND2_5559 ( R2027_U102 , R2027_U116 , INSTADDRPOINTER_REG_25_ );
nand NAND2_5560 ( R2027_U103 , R2027_U115 , INSTADDRPOINTER_REG_23_ );
nand NAND2_5561 ( R2027_U104 , R2027_U121 , INSTADDRPOINTER_REG_21_ );
nand NAND2_5562 ( R2027_U105 , R2027_U114 , INSTADDRPOINTER_REG_19_ );
nand NAND2_5563 ( R2027_U106 , R2027_U117 , INSTADDRPOINTER_REG_17_ );
nand NAND2_5564 ( R2027_U107 , R2027_U124 , INSTADDRPOINTER_REG_15_ );
nand NAND2_5565 ( R2027_U108 , R2027_U119 , INSTADDRPOINTER_REG_13_ );
nand NAND2_5566 ( R2027_U109 , R2027_U113 , INSTADDRPOINTER_REG_11_ );
nand NAND2_5567 ( R2027_U110 , INSTADDRPOINTER_REG_9_ , R2027_U120 );
not NOT1_5568 ( R2027_U111 , R2027_U10 );
not NOT1_5569 ( R2027_U112 , R2027_U13 );
not NOT1_5570 ( R2027_U113 , R2027_U22 );
not NOT1_5571 ( R2027_U114 , R2027_U34 );
not NOT1_5572 ( R2027_U115 , R2027_U40 );
not NOT1_5573 ( R2027_U116 , R2027_U43 );
not NOT1_5574 ( R2027_U117 , R2027_U31 );
not NOT1_5575 ( R2027_U118 , R2027_U16 );
not NOT1_5576 ( R2027_U119 , R2027_U25 );
not NOT1_5577 ( R2027_U120 , R2027_U17 );
not NOT1_5578 ( R2027_U121 , R2027_U36 );
not NOT1_5579 ( R2027_U122 , R2027_U46 );
not NOT1_5580 ( R2027_U123 , R2027_U48 );
not NOT1_5581 ( R2027_U124 , R2027_U27 );
not NOT1_5582 ( R2027_U125 , R2027_U95 );
not NOT1_5583 ( R2027_U126 , R2027_U96 );
not NOT1_5584 ( R2027_U127 , R2027_U97 );
not NOT1_5585 ( R2027_U128 , R2027_U49 );
not NOT1_5586 ( R2027_U129 , R2027_U99 );
not NOT1_5587 ( R2027_U130 , R2027_U100 );
not NOT1_5588 ( R2027_U131 , R2027_U101 );
not NOT1_5589 ( R2027_U132 , R2027_U102 );
not NOT1_5590 ( R2027_U133 , R2027_U103 );
not NOT1_5591 ( R2027_U134 , R2027_U104 );
not NOT1_5592 ( R2027_U135 , R2027_U105 );
not NOT1_5593 ( R2027_U136 , R2027_U106 );
not NOT1_5594 ( R2027_U137 , R2027_U107 );
not NOT1_5595 ( R2027_U138 , R2027_U108 );
not NOT1_5596 ( R2027_U139 , R2027_U109 );
not NOT1_5597 ( R2027_U140 , R2027_U110 );
nand NAND2_5598 ( R2027_U141 , R2027_U120 , R2027_U18 );
nand NAND2_5599 ( R2027_U142 , INSTADDRPOINTER_REG_9_ , R2027_U17 );
nand NAND2_5600 ( R2027_U143 , INSTADDRPOINTER_REG_8_ , R2027_U95 );
nand NAND2_5601 ( R2027_U144 , R2027_U125 , R2027_U14 );
nand NAND2_5602 ( R2027_U145 , R2027_U118 , R2027_U15 );
nand NAND2_5603 ( R2027_U146 , INSTADDRPOINTER_REG_7_ , R2027_U16 );
nand NAND2_5604 ( R2027_U147 , INSTADDRPOINTER_REG_6_ , R2027_U96 );
nand NAND2_5605 ( R2027_U148 , R2027_U126 , R2027_U11 );
nand NAND2_5606 ( R2027_U149 , R2027_U112 , R2027_U12 );
nand NAND2_5607 ( R2027_U150 , INSTADDRPOINTER_REG_5_ , R2027_U13 );
nand NAND2_5608 ( R2027_U151 , INSTADDRPOINTER_REG_4_ , R2027_U97 );
nand NAND2_5609 ( R2027_U152 , R2027_U127 , R2027_U8 );
nand NAND2_5610 ( R2027_U153 , R2027_U111 , R2027_U9 );
nand NAND2_5611 ( R2027_U154 , INSTADDRPOINTER_REG_3_ , R2027_U10 );
nand NAND2_5612 ( R2027_U155 , INSTADDRPOINTER_REG_31_ , R2027_U99 );
nand NAND2_5613 ( R2027_U156 , R2027_U129 , R2027_U98 );
nand NAND2_5614 ( R2027_U157 , INSTADDRPOINTER_REG_30_ , R2027_U49 );
nand NAND2_5615 ( R2027_U158 , R2027_U128 , R2027_U50 );
nand NAND2_5616 ( R2027_U159 , INSTADDRPOINTER_REG_2_ , R2027_U100 );
nand NAND2_5617 ( R2027_U160 , R2027_U130 , R2027_U6 );
nand NAND2_5618 ( R2027_U161 , R2027_U123 , R2027_U47 );
nand NAND2_5619 ( R2027_U162 , INSTADDRPOINTER_REG_29_ , R2027_U48 );
nand NAND2_5620 ( R2027_U163 , INSTADDRPOINTER_REG_28_ , R2027_U101 );
nand NAND2_5621 ( R2027_U164 , R2027_U131 , R2027_U45 );
nand NAND2_5622 ( R2027_U165 , R2027_U122 , R2027_U44 );
nand NAND2_5623 ( R2027_U166 , INSTADDRPOINTER_REG_27_ , R2027_U46 );
nand NAND2_5624 ( R2027_U167 , INSTADDRPOINTER_REG_26_ , R2027_U102 );
nand NAND2_5625 ( R2027_U168 , R2027_U132 , R2027_U41 );
nand NAND2_5626 ( R2027_U169 , R2027_U116 , R2027_U42 );
nand NAND2_5627 ( R2027_U170 , INSTADDRPOINTER_REG_25_ , R2027_U43 );
nand NAND2_5628 ( R2027_U171 , INSTADDRPOINTER_REG_24_ , R2027_U103 );
nand NAND2_5629 ( R2027_U172 , R2027_U133 , R2027_U38 );
nand NAND2_5630 ( R2027_U173 , R2027_U115 , R2027_U39 );
nand NAND2_5631 ( R2027_U174 , INSTADDRPOINTER_REG_23_ , R2027_U40 );
nand NAND2_5632 ( R2027_U175 , INSTADDRPOINTER_REG_22_ , R2027_U104 );
nand NAND2_5633 ( R2027_U176 , R2027_U134 , R2027_U37 );
nand NAND2_5634 ( R2027_U177 , R2027_U121 , R2027_U35 );
nand NAND2_5635 ( R2027_U178 , INSTADDRPOINTER_REG_21_ , R2027_U36 );
nand NAND2_5636 ( R2027_U179 , INSTADDRPOINTER_REG_20_ , R2027_U105 );
nand NAND2_5637 ( R2027_U180 , R2027_U135 , R2027_U32 );
nand NAND2_5638 ( R2027_U181 , INSTADDRPOINTER_REG_0_ , R2027_U7 );
nand NAND2_5639 ( R2027_U182 , INSTADDRPOINTER_REG_1_ , R2027_U5 );
nand NAND2_5640 ( R2027_U183 , R2027_U114 , R2027_U33 );
nand NAND2_5641 ( R2027_U184 , INSTADDRPOINTER_REG_19_ , R2027_U34 );
nand NAND2_5642 ( R2027_U185 , INSTADDRPOINTER_REG_18_ , R2027_U106 );
nand NAND2_5643 ( R2027_U186 , R2027_U136 , R2027_U29 );
nand NAND2_5644 ( R2027_U187 , R2027_U117 , R2027_U30 );
nand NAND2_5645 ( R2027_U188 , INSTADDRPOINTER_REG_17_ , R2027_U31 );
nand NAND2_5646 ( R2027_U189 , INSTADDRPOINTER_REG_16_ , R2027_U107 );
nand NAND2_5647 ( R2027_U190 , R2027_U137 , R2027_U28 );
nand NAND2_5648 ( R2027_U191 , R2027_U124 , R2027_U26 );
nand NAND2_5649 ( R2027_U192 , INSTADDRPOINTER_REG_15_ , R2027_U27 );
nand NAND2_5650 ( R2027_U193 , INSTADDRPOINTER_REG_14_ , R2027_U108 );
nand NAND2_5651 ( R2027_U194 , R2027_U138 , R2027_U23 );
nand NAND2_5652 ( R2027_U195 , R2027_U119 , R2027_U24 );
nand NAND2_5653 ( R2027_U196 , INSTADDRPOINTER_REG_13_ , R2027_U25 );
nand NAND2_5654 ( R2027_U197 , INSTADDRPOINTER_REG_12_ , R2027_U109 );
nand NAND2_5655 ( R2027_U198 , R2027_U139 , R2027_U20 );
nand NAND2_5656 ( R2027_U199 , R2027_U113 , R2027_U21 );
nand NAND2_5657 ( R2027_U200 , INSTADDRPOINTER_REG_11_ , R2027_U22 );
nand NAND2_5658 ( R2027_U201 , INSTADDRPOINTER_REG_10_ , R2027_U110 );
nand NAND2_5659 ( R2027_U202 , R2027_U140 , R2027_U19 );
and AND2_5660 ( R2278_U5 , R2278_U217 , R2278_U215 );
and AND2_5661 ( R2278_U6 , R2278_U227 , R2278_U225 );
and AND2_5662 ( R2278_U7 , R2278_U6 , R2278_U208 );
and AND2_5663 ( R2278_U8 , R2278_U7 , R2278_U207 );
and AND2_5664 ( R2278_U9 , R2278_U235 , R2278_U231 );
and AND2_5665 ( R2278_U10 , R2278_U9 , R2278_U206 );
and AND2_5666 ( R2278_U11 , R2278_U10 , R2278_U205 );
and AND2_5667 ( R2278_U12 , R2278_U11 , R2278_U242 );
and AND2_5668 ( R2278_U13 , R2278_U12 , R2278_U204 );
and AND2_5669 ( R2278_U14 , R2278_U250 , R2278_U246 );
and AND2_5670 ( R2278_U15 , R2278_U14 , R2278_U253 );
and AND2_5671 ( R2278_U16 , R2278_U15 , R2278_U256 );
and AND2_5672 ( R2278_U17 , R2278_U292 , R2278_U19 );
nand NAND2_5673 ( R2278_U18 , U2783 , INSTADDRPOINTER_REG_4_ );
nand NAND2_5674 ( R2278_U19 , U2787 , INSTADDRPOINTER_REG_0_ );
nand NAND2_5675 ( R2278_U20 , U2782 , INSTADDRPOINTER_REG_5_ );
not NOT1_5676 ( R2278_U21 , INSTADDRPOINTER_REG_30_ );
not NOT1_5677 ( R2278_U22 , U2770 );
nand NAND2_5678 ( R2278_U23 , U2770 , INSTADDRPOINTER_REG_19_ );
nand NAND2_5679 ( R2278_U24 , U2771 , INSTADDRPOINTER_REG_16_ );
nand NAND2_5680 ( R2278_U25 , R2278_U40 , R2278_U207 );
nand NAND2_5681 ( R2278_U26 , U2779 , INSTADDRPOINTER_REG_8_ );
nand NAND2_5682 ( R2278_U27 , U2778 , INSTADDRPOINTER_REG_9_ );
nand NAND2_5683 ( R2278_U28 , U2777 , INSTADDRPOINTER_REG_10_ );
nand NAND2_5684 ( R2278_U29 , U2775 , INSTADDRPOINTER_REG_12_ );
nand NAND2_5685 ( R2278_U30 , U2773 , INSTADDRPOINTER_REG_14_ );
nand NAND2_5686 ( R2278_U31 , U2774 , INSTADDRPOINTER_REG_13_ );
not NOT1_5687 ( R2278_U32 , INSTADDRPOINTER_REG_29_ );
not NOT1_5688 ( R2278_U33 , U2770 );
not NOT1_5689 ( R2278_U34 , INSTADDRPOINTER_REG_28_ );
not NOT1_5690 ( R2278_U35 , U2770 );
nand NAND2_5691 ( R2278_U36 , U2770 , INSTADDRPOINTER_REG_26_ );
nand NAND2_5692 ( R2278_U37 , R2278_U328 , R2278_U257 );
nand NAND2_5693 ( R2278_U38 , R2278_U325 , R2278_U254 );
nand NAND2_5694 ( R2278_U39 , R2278_U322 , R2278_U251 );
nand NAND2_5695 ( R2278_U40 , R2278_U306 , R2278_U229 );
nand NAND2_5696 ( R2278_U41 , R2278_U304 , R2278_U228 );
nand NAND2_5697 ( R2278_U42 , R2278_U402 , R2278_U401 );
and AND2_5698 ( R2278_U43 , R2278_U178 , R2278_U162 );
and AND2_5699 ( R2278_U44 , R2278_U303 , R2278_U179 );
and AND2_5700 ( R2278_U45 , R2278_U182 , R2278_U163 );
and AND2_5701 ( R2278_U46 , R2278_U302 , R2278_U301 );
and AND2_5702 ( R2278_U47 , INSTADDRPOINTER_REG_20_ , U2770 );
and AND2_5703 ( R2278_U48 , R2278_U178 , R2278_U162 );
and AND2_5704 ( R2278_U49 , R2278_U337 , R2278_U179 );
and AND3_5705 ( R2278_U50 , R2278_U301 , R2278_U163 , R2278_U182 );
and AND2_5706 ( R2278_U51 , R2278_U189 , R2278_U185 );
and AND2_5707 ( R2278_U52 , R2278_U5 , R2278_U51 );
and AND2_5708 ( R2278_U53 , R2278_U186 , R2278_U189 );
and AND4_5709 ( R2278_U54 , R2278_U293 , R2278_U216 , R2278_U296 , R2278_U295 );
and AND4_5710 ( R2278_U55 , R2278_U211 , R2278_U213 , R2278_U221 , R2278_U209 );
and AND4_5711 ( R2278_U56 , R2278_U294 , R2278_U210 , R2278_U298 , R2278_U297 );
and AND2_5712 ( R2278_U57 , R2278_U13 , R2278_U8 );
and AND2_5713 ( R2278_U58 , R2278_U332 , R2278_U245 );
and AND3_5714 ( R2278_U59 , R2278_U333 , R2278_U320 , R2278_U58 );
and AND2_5715 ( R2278_U60 , R2278_U16 , R2278_U259 );
and AND2_5716 ( R2278_U61 , R2278_U331 , R2278_U260 );
nand NAND2_5717 ( R2278_U62 , R2278_U364 , R2278_U363 );
nand NAND2_5718 ( R2278_U63 , R2278_U369 , R2278_U368 );
nand NAND2_5719 ( R2278_U64 , R2278_U376 , R2278_U375 );
nand NAND2_5720 ( R2278_U65 , R2278_U381 , R2278_U380 );
and AND2_5721 ( R2278_U66 , R2278_U25 , R2278_U23 );
and AND2_5722 ( R2278_U67 , R2278_U318 , R2278_U243 );
and AND2_5723 ( R2278_U68 , R2278_U315 , R2278_U240 );
and AND2_5724 ( R2278_U69 , R2278_U312 , R2278_U238 );
and AND2_5725 ( R2278_U70 , R2278_U310 , R2278_U236 );
and AND4_5726 ( R2278_U71 , R2278_U293 , R2278_U216 , R2278_U296 , R2278_U295 );
nand NAND2_5727 ( R2278_U72 , R2278_U26 , R2278_U187 );
nand NAND2_5728 ( R2278_U73 , R2278_U189 , R2278_U27 );
and AND2_5729 ( R2278_U74 , R2278_U350 , R2278_U349 );
nand NAND3_5730 ( R2278_U75 , R2278_U46 , R2278_U183 , R2278_U45 );
nand NAND2_5731 ( R2278_U76 , R2278_U185 , R2278_U26 );
and AND2_5732 ( R2278_U77 , R2278_U352 , R2278_U351 );
nand NAND2_5733 ( R2278_U78 , R2278_U197 , R2278_U165 );
nand NAND2_5734 ( R2278_U79 , R2278_U162 , R2278_U163 );
and AND2_5735 ( R2278_U80 , R2278_U354 , R2278_U353 );
nand NAND2_5736 ( R2278_U81 , R2278_U20 , R2278_U195 );
nand NAND2_5737 ( R2278_U82 , R2278_U165 , R2278_U164 );
and AND2_5738 ( R2278_U83 , R2278_U356 , R2278_U355 );
nand NAND2_5739 ( R2278_U84 , R2278_U18 , R2278_U193 );
nand NAND2_5740 ( R2278_U85 , R2278_U179 , R2278_U20 );
and AND2_5741 ( R2278_U86 , R2278_U358 , R2278_U357 );
nand NAND2_5742 ( R2278_U87 , R2278_U175 , R2278_U176 );
nand NAND2_5743 ( R2278_U88 , R2278_U178 , R2278_U18 );
and AND2_5744 ( R2278_U89 , R2278_U360 , R2278_U359 );
nand NAND2_5745 ( R2278_U90 , R2278_U172 , R2278_U173 );
nand NAND2_5746 ( R2278_U91 , R2278_U166 , R2278_U175 );
and AND2_5747 ( R2278_U92 , R2278_U362 , R2278_U361 );
not NOT1_5748 ( R2278_U93 , U2769 );
not NOT1_5749 ( R2278_U94 , INSTADDRPOINTER_REG_31_ );
nand NAND2_5750 ( R2278_U95 , R2278_U61 , R2278_U330 );
and AND2_5751 ( R2278_U96 , R2278_U367 , R2278_U366 );
nand NAND2_5752 ( R2278_U97 , R2278_U329 , R2278_U327 );
and AND2_5753 ( R2278_U98 , R2278_U372 , R2278_U371 );
nand NAND2_5754 ( R2278_U99 , R2278_U169 , R2278_U170 );
nand NAND2_5755 ( R2278_U100 , R2278_U167 , R2278_U172 );
and AND2_5756 ( R2278_U101 , R2278_U374 , R2278_U373 );
nand NAND2_5757 ( R2278_U102 , R2278_U326 , R2278_U324 );
and AND2_5758 ( R2278_U103 , R2278_U379 , R2278_U378 );
nand NAND2_5759 ( R2278_U104 , R2278_U323 , R2278_U321 );
and AND2_5760 ( R2278_U105 , R2278_U384 , R2278_U383 );
nand NAND2_5761 ( R2278_U106 , R2278_U36 , R2278_U248 );
nand NAND2_5762 ( R2278_U107 , R2278_U250 , R2278_U251 );
and AND2_5763 ( R2278_U108 , R2278_U386 , R2278_U385 );
nand NAND2_5764 ( R2278_U109 , R2278_U246 , R2278_U36 );
nand NAND2_5765 ( R2278_U110 , R2278_U59 , R2278_U347 );
and AND2_5766 ( R2278_U111 , R2278_U388 , R2278_U387 );
nand NAND2_5767 ( R2278_U112 , R2278_U67 , R2278_U316 );
nand NAND2_5768 ( R2278_U113 , R2278_U204 , R2278_U245 );
and AND2_5769 ( R2278_U114 , R2278_U390 , R2278_U389 );
nand NAND2_5770 ( R2278_U115 , R2278_U68 , R2278_U313 );
nand NAND2_5771 ( R2278_U116 , R2278_U243 , R2278_U242 );
and AND2_5772 ( R2278_U117 , R2278_U392 , R2278_U391 );
nand NAND2_5773 ( R2278_U118 , R2278_U69 , R2278_U311 );
nand NAND2_5774 ( R2278_U119 , R2278_U240 , R2278_U205 );
and AND2_5775 ( R2278_U120 , R2278_U394 , R2278_U393 );
nand NAND2_5776 ( R2278_U121 , R2278_U70 , R2278_U309 );
nand NAND2_5777 ( R2278_U122 , R2278_U238 , R2278_U206 );
and AND2_5778 ( R2278_U123 , R2278_U396 , R2278_U395 );
nand NAND2_5779 ( R2278_U124 , R2278_U232 , R2278_U233 );
nand NAND2_5780 ( R2278_U125 , R2278_U236 , R2278_U235 );
and AND2_5781 ( R2278_U126 , R2278_U398 , R2278_U397 );
nand NAND2_5782 ( R2278_U127 , R2278_U231 , R2278_U232 );
nand NAND2_5783 ( R2278_U128 , R2278_U66 , R2278_U345 );
and AND2_5784 ( R2278_U129 , R2278_U400 , R2278_U399 );
nand NAND2_5785 ( R2278_U130 , R2278_U168 , R2278_U169 );
nand NAND2_5786 ( R2278_U131 , R2278_U207 , R2278_U23 );
nand NAND2_5787 ( R2278_U132 , R2278_U307 , R2278_U343 );
and AND2_5788 ( R2278_U133 , R2278_U404 , R2278_U403 );
nand NAND2_5789 ( R2278_U134 , R2278_U208 , R2278_U229 );
nand NAND2_5790 ( R2278_U135 , R2278_U305 , R2278_U341 );
and AND2_5791 ( R2278_U136 , R2278_U406 , R2278_U405 );
nand NAND2_5792 ( R2278_U137 , R2278_U227 , R2278_U228 );
nand NAND2_5793 ( R2278_U138 , R2278_U339 , R2278_U24 );
and AND2_5794 ( R2278_U139 , R2278_U408 , R2278_U407 );
nand NAND2_5795 ( R2278_U140 , R2278_U223 , R2278_U56 );
nand NAND2_5796 ( R2278_U141 , R2278_U225 , R2278_U24 );
and AND2_5797 ( R2278_U142 , R2278_U410 , R2278_U409 );
nand NAND2_5798 ( R2278_U143 , R2278_U280 , R2278_U30 );
nand NAND2_5799 ( R2278_U144 , R2278_U209 , R2278_U210 );
and AND2_5800 ( R2278_U145 , R2278_U412 , R2278_U411 );
nand NAND2_5801 ( R2278_U146 , R2278_U31 , R2278_U278 );
nand NAND2_5802 ( R2278_U147 , R2278_U30 , R2278_U211 );
and AND2_5803 ( R2278_U148 , R2278_U414 , R2278_U413 );
nand NAND2_5804 ( R2278_U149 , R2278_U29 , R2278_U276 );
nand NAND2_5805 ( R2278_U150 , R2278_U213 , R2278_U31 );
and AND2_5806 ( R2278_U151 , R2278_U416 , R2278_U415 );
nand NAND2_5807 ( R2278_U152 , R2278_U219 , R2278_U71 );
nand NAND2_5808 ( R2278_U153 , R2278_U221 , R2278_U29 );
and AND2_5809 ( R2278_U154 , R2278_U418 , R2278_U417 );
nand NAND2_5810 ( R2278_U155 , R2278_U288 , R2278_U28 );
nand NAND2_5811 ( R2278_U156 , R2278_U215 , R2278_U216 );
and AND2_5812 ( R2278_U157 , R2278_U420 , R2278_U419 );
nand NAND2_5813 ( R2278_U158 , R2278_U27 , R2278_U286 );
nand NAND2_5814 ( R2278_U159 , R2278_U28 , R2278_U217 );
and AND2_5815 ( R2278_U160 , R2278_U422 , R2278_U421 );
not NOT1_5816 ( R2278_U161 , R2278_U19 );
or OR2_5817 ( R2278_U162 , INSTADDRPOINTER_REG_7_ , U2780 );
nand NAND2_5818 ( R2278_U163 , U2780 , INSTADDRPOINTER_REG_7_ );
or OR2_5819 ( R2278_U164 , INSTADDRPOINTER_REG_6_ , U2781 );
nand NAND2_5820 ( R2278_U165 , U2781 , INSTADDRPOINTER_REG_6_ );
or OR2_5821 ( R2278_U166 , INSTADDRPOINTER_REG_3_ , U2784 );
or OR2_5822 ( R2278_U167 , INSTADDRPOINTER_REG_2_ , U2785 );
or OR2_5823 ( R2278_U168 , INSTADDRPOINTER_REG_1_ , U2786 );
nand NAND2_5824 ( R2278_U169 , U2786 , INSTADDRPOINTER_REG_1_ );
nand NAND2_5825 ( R2278_U170 , R2278_U161 , R2278_U168 );
not NOT1_5826 ( R2278_U171 , R2278_U99 );
nand NAND2_5827 ( R2278_U172 , U2785 , INSTADDRPOINTER_REG_2_ );
nand NAND2_5828 ( R2278_U173 , R2278_U99 , R2278_U299 );
not NOT1_5829 ( R2278_U174 , R2278_U90 );
nand NAND2_5830 ( R2278_U175 , U2784 , INSTADDRPOINTER_REG_3_ );
nand NAND2_5831 ( R2278_U176 , R2278_U300 , R2278_U166 );
not NOT1_5832 ( R2278_U177 , R2278_U87 );
or OR2_5833 ( R2278_U178 , INSTADDRPOINTER_REG_4_ , U2783 );
or OR2_5834 ( R2278_U179 , INSTADDRPOINTER_REG_5_ , U2782 );
not NOT1_5835 ( R2278_U180 , R2278_U20 );
not NOT1_5836 ( R2278_U181 , R2278_U18 );
nand NAND4_5837 ( R2278_U182 , R2278_U181 , R2278_U179 , R2278_U164 , R2278_U162 );
nand NAND3_5838 ( R2278_U183 , R2278_U43 , R2278_U87 , R2278_U44 );
not NOT1_5839 ( R2278_U184 , R2278_U75 );
or OR2_5840 ( R2278_U185 , INSTADDRPOINTER_REG_8_ , U2779 );
not NOT1_5841 ( R2278_U186 , R2278_U26 );
nand NAND2_5842 ( R2278_U187 , R2278_U185 , R2278_U75 );
not NOT1_5843 ( R2278_U188 , R2278_U72 );
or OR2_5844 ( R2278_U189 , INSTADDRPOINTER_REG_9_ , U2778 );
not NOT1_5845 ( R2278_U190 , R2278_U27 );
not NOT1_5846 ( R2278_U191 , R2278_U73 );
not NOT1_5847 ( R2278_U192 , R2278_U76 );
nand NAND2_5848 ( R2278_U193 , R2278_U178 , R2278_U87 );
not NOT1_5849 ( R2278_U194 , R2278_U84 );
nand NAND2_5850 ( R2278_U195 , R2278_U84 , R2278_U179 );
not NOT1_5851 ( R2278_U196 , R2278_U81 );
nand NAND2_5852 ( R2278_U197 , R2278_U81 , R2278_U164 );
not NOT1_5853 ( R2278_U198 , R2278_U78 );
not NOT1_5854 ( R2278_U199 , R2278_U79 );
not NOT1_5855 ( R2278_U200 , R2278_U82 );
not NOT1_5856 ( R2278_U201 , R2278_U85 );
not NOT1_5857 ( R2278_U202 , R2278_U88 );
not NOT1_5858 ( R2278_U203 , R2278_U91 );
or OR2_5859 ( R2278_U204 , INSTADDRPOINTER_REG_25_ , U2770 );
or OR2_5860 ( R2278_U205 , INSTADDRPOINTER_REG_23_ , U2770 );
or OR2_5861 ( R2278_U206 , INSTADDRPOINTER_REG_22_ , U2770 );
or OR2_5862 ( R2278_U207 , INSTADDRPOINTER_REG_19_ , U2770 );
or OR2_5863 ( R2278_U208 , INSTADDRPOINTER_REG_18_ , U2770 );
or OR2_5864 ( R2278_U209 , INSTADDRPOINTER_REG_15_ , U2772 );
nand NAND2_5865 ( R2278_U210 , U2772 , INSTADDRPOINTER_REG_15_ );
or OR2_5866 ( R2278_U211 , INSTADDRPOINTER_REG_14_ , U2773 );
not NOT1_5867 ( R2278_U212 , R2278_U30 );
or OR2_5868 ( R2278_U213 , INSTADDRPOINTER_REG_13_ , U2774 );
not NOT1_5869 ( R2278_U214 , R2278_U31 );
or OR2_5870 ( R2278_U215 , INSTADDRPOINTER_REG_11_ , U2776 );
nand NAND2_5871 ( R2278_U216 , U2776 , INSTADDRPOINTER_REG_11_ );
or OR2_5872 ( R2278_U217 , INSTADDRPOINTER_REG_10_ , U2777 );
not NOT1_5873 ( R2278_U218 , R2278_U28 );
nand NAND2_5874 ( R2278_U219 , R2278_U52 , R2278_U335 );
not NOT1_5875 ( R2278_U220 , R2278_U152 );
or OR2_5876 ( R2278_U221 , INSTADDRPOINTER_REG_12_ , U2775 );
not NOT1_5877 ( R2278_U222 , R2278_U29 );
nand NAND2_5878 ( R2278_U223 , R2278_U55 , R2278_U338 );
not NOT1_5879 ( R2278_U224 , R2278_U140 );
or OR2_5880 ( R2278_U225 , INSTADDRPOINTER_REG_16_ , U2771 );
not NOT1_5881 ( R2278_U226 , R2278_U24 );
or OR2_5882 ( R2278_U227 , INSTADDRPOINTER_REG_17_ , U2770 );
nand NAND2_5883 ( R2278_U228 , U2770 , INSTADDRPOINTER_REG_17_ );
nand NAND2_5884 ( R2278_U229 , U2770 , INSTADDRPOINTER_REG_18_ );
not NOT1_5885 ( R2278_U230 , R2278_U23 );
or OR2_5886 ( R2278_U231 , INSTADDRPOINTER_REG_20_ , U2770 );
nand NAND2_5887 ( R2278_U232 , U2770 , INSTADDRPOINTER_REG_20_ );
nand NAND2_5888 ( R2278_U233 , R2278_U231 , R2278_U128 );
not NOT1_5889 ( R2278_U234 , R2278_U124 );
or OR2_5890 ( R2278_U235 , INSTADDRPOINTER_REG_21_ , U2770 );
nand NAND2_5891 ( R2278_U236 , U2770 , INSTADDRPOINTER_REG_21_ );
not NOT1_5892 ( R2278_U237 , R2278_U121 );
nand NAND2_5893 ( R2278_U238 , U2770 , INSTADDRPOINTER_REG_22_ );
not NOT1_5894 ( R2278_U239 , R2278_U118 );
nand NAND2_5895 ( R2278_U240 , U2770 , INSTADDRPOINTER_REG_23_ );
not NOT1_5896 ( R2278_U241 , R2278_U115 );
or OR2_5897 ( R2278_U242 , INSTADDRPOINTER_REG_24_ , U2770 );
nand NAND2_5898 ( R2278_U243 , U2770 , INSTADDRPOINTER_REG_24_ );
not NOT1_5899 ( R2278_U244 , R2278_U112 );
nand NAND2_5900 ( R2278_U245 , U2770 , INSTADDRPOINTER_REG_25_ );
or OR2_5901 ( R2278_U246 , INSTADDRPOINTER_REG_26_ , U2770 );
not NOT1_5902 ( R2278_U247 , R2278_U36 );
nand NAND2_5903 ( R2278_U248 , R2278_U246 , R2278_U110 );
not NOT1_5904 ( R2278_U249 , R2278_U106 );
or OR2_5905 ( R2278_U250 , INSTADDRPOINTER_REG_27_ , U2770 );
nand NAND2_5906 ( R2278_U251 , U2770 , INSTADDRPOINTER_REG_27_ );
not NOT1_5907 ( R2278_U252 , R2278_U104 );
or OR2_5908 ( R2278_U253 , INSTADDRPOINTER_REG_28_ , U2770 );
nand NAND2_5909 ( R2278_U254 , U2770 , INSTADDRPOINTER_REG_28_ );
not NOT1_5910 ( R2278_U255 , R2278_U102 );
or OR2_5911 ( R2278_U256 , INSTADDRPOINTER_REG_29_ , U2770 );
nand NAND2_5912 ( R2278_U257 , U2770 , INSTADDRPOINTER_REG_29_ );
not NOT1_5913 ( R2278_U258 , R2278_U97 );
or OR2_5914 ( R2278_U259 , INSTADDRPOINTER_REG_30_ , U2770 );
nand NAND2_5915 ( R2278_U260 , U2770 , INSTADDRPOINTER_REG_30_ );
not NOT1_5916 ( R2278_U261 , R2278_U95 );
not NOT1_5917 ( R2278_U262 , R2278_U100 );
not NOT1_5918 ( R2278_U263 , R2278_U107 );
not NOT1_5919 ( R2278_U264 , R2278_U109 );
not NOT1_5920 ( R2278_U265 , R2278_U113 );
not NOT1_5921 ( R2278_U266 , R2278_U116 );
not NOT1_5922 ( R2278_U267 , R2278_U119 );
not NOT1_5923 ( R2278_U268 , R2278_U122 );
not NOT1_5924 ( R2278_U269 , R2278_U125 );
not NOT1_5925 ( R2278_U270 , R2278_U127 );
not NOT1_5926 ( R2278_U271 , R2278_U130 );
not NOT1_5927 ( R2278_U272 , R2278_U131 );
not NOT1_5928 ( R2278_U273 , R2278_U134 );
not NOT1_5929 ( R2278_U274 , R2278_U137 );
not NOT1_5930 ( R2278_U275 , R2278_U141 );
nand NAND2_5931 ( R2278_U276 , R2278_U221 , R2278_U152 );
not NOT1_5932 ( R2278_U277 , R2278_U149 );
nand NAND2_5933 ( R2278_U278 , R2278_U149 , R2278_U213 );
not NOT1_5934 ( R2278_U279 , R2278_U146 );
nand NAND2_5935 ( R2278_U280 , R2278_U146 , R2278_U211 );
not NOT1_5936 ( R2278_U281 , R2278_U143 );
not NOT1_5937 ( R2278_U282 , R2278_U144 );
not NOT1_5938 ( R2278_U283 , R2278_U147 );
not NOT1_5939 ( R2278_U284 , R2278_U150 );
not NOT1_5940 ( R2278_U285 , R2278_U153 );
nand NAND2_5941 ( R2278_U286 , R2278_U189 , R2278_U72 );
not NOT1_5942 ( R2278_U287 , R2278_U158 );
nand NAND2_5943 ( R2278_U288 , R2278_U158 , R2278_U217 );
not NOT1_5944 ( R2278_U289 , R2278_U155 );
not NOT1_5945 ( R2278_U290 , R2278_U156 );
not NOT1_5946 ( R2278_U291 , R2278_U159 );
or OR2_5947 ( R2278_U292 , INSTADDRPOINTER_REG_0_ , U2787 );
nand NAND2_5948 ( R2278_U293 , R2278_U53 , R2278_U5 );
nand NAND4_5949 ( R2278_U294 , R2278_U222 , R2278_U213 , R2278_U211 , R2278_U209 );
nand NAND2_5950 ( R2278_U295 , R2278_U190 , R2278_U5 );
nand NAND2_5951 ( R2278_U296 , R2278_U218 , R2278_U5 );
nand NAND2_5952 ( R2278_U297 , R2278_U212 , R2278_U209 );
nand NAND3_5953 ( R2278_U298 , R2278_U211 , R2278_U214 , R2278_U209 );
or OR2_5954 ( R2278_U299 , INSTADDRPOINTER_REG_2_ , U2785 );
nand NAND2_5955 ( R2278_U300 , R2278_U172 , R2278_U173 );
nand NAND3_5956 ( R2278_U301 , INSTADDRPOINTER_REG_6_ , R2278_U162 , U2781 );
nand NAND3_5957 ( R2278_U302 , R2278_U180 , R2278_U162 , R2278_U164 );
or OR2_5958 ( R2278_U303 , INSTADDRPOINTER_REG_6_ , U2781 );
nand NAND2_5959 ( R2278_U304 , R2278_U226 , R2278_U227 );
not NOT1_5960 ( R2278_U305 , R2278_U41 );
nand NAND2_5961 ( R2278_U306 , R2278_U41 , R2278_U208 );
not NOT1_5962 ( R2278_U307 , R2278_U40 );
not NOT1_5963 ( R2278_U308 , R2278_U25 );
nand NAND2_5964 ( R2278_U309 , R2278_U9 , R2278_U128 );
nand NAND2_5965 ( R2278_U310 , R2278_U47 , R2278_U235 );
nand NAND2_5966 ( R2278_U311 , R2278_U10 , R2278_U128 );
nand NAND2_5967 ( R2278_U312 , R2278_U334 , R2278_U206 );
nand NAND2_5968 ( R2278_U313 , R2278_U11 , R2278_U128 );
nand NAND2_5969 ( R2278_U314 , R2278_U312 , R2278_U238 );
nand NAND2_5970 ( R2278_U315 , R2278_U314 , R2278_U205 );
nand NAND2_5971 ( R2278_U316 , R2278_U12 , R2278_U128 );
nand NAND2_5972 ( R2278_U317 , R2278_U315 , R2278_U240 );
nand NAND2_5973 ( R2278_U318 , R2278_U317 , R2278_U242 );
nand NAND2_5974 ( R2278_U319 , R2278_U318 , R2278_U243 );
nand NAND2_5975 ( R2278_U320 , R2278_U319 , R2278_U204 );
nand NAND2_5976 ( R2278_U321 , R2278_U14 , R2278_U110 );
nand NAND2_5977 ( R2278_U322 , R2278_U247 , R2278_U250 );
not NOT1_5978 ( R2278_U323 , R2278_U39 );
nand NAND2_5979 ( R2278_U324 , R2278_U15 , R2278_U110 );
nand NAND2_5980 ( R2278_U325 , R2278_U39 , R2278_U253 );
not NOT1_5981 ( R2278_U326 , R2278_U38 );
nand NAND2_5982 ( R2278_U327 , R2278_U16 , R2278_U110 );
nand NAND2_5983 ( R2278_U328 , R2278_U38 , R2278_U256 );
not NOT1_5984 ( R2278_U329 , R2278_U37 );
nand NAND2_5985 ( R2278_U330 , R2278_U60 , R2278_U110 );
nand NAND2_5986 ( R2278_U331 , R2278_U37 , R2278_U259 );
nand NAND2_5987 ( R2278_U332 , R2278_U230 , R2278_U13 );
nand NAND2_5988 ( R2278_U333 , R2278_U308 , R2278_U13 );
nand NAND2_5989 ( R2278_U334 , R2278_U310 , R2278_U236 );
nand NAND3_5990 ( R2278_U335 , R2278_U336 , R2278_U302 , R2278_U50 );
nand NAND3_5991 ( R2278_U336 , R2278_U48 , R2278_U87 , R2278_U49 );
or OR2_5992 ( R2278_U337 , INSTADDRPOINTER_REG_6_ , U2781 );
nand NAND2_5993 ( R2278_U338 , R2278_U219 , R2278_U54 );
nand NAND2_5994 ( R2278_U339 , R2278_U225 , R2278_U140 );
not NOT1_5995 ( R2278_U340 , R2278_U138 );
nand NAND2_5996 ( R2278_U341 , R2278_U6 , R2278_U140 );
not NOT1_5997 ( R2278_U342 , R2278_U135 );
nand NAND2_5998 ( R2278_U343 , R2278_U7 , R2278_U140 );
not NOT1_5999 ( R2278_U344 , R2278_U132 );
nand NAND2_6000 ( R2278_U345 , R2278_U8 , R2278_U140 );
not NOT1_6001 ( R2278_U346 , R2278_U128 );
nand NAND2_6002 ( R2278_U347 , R2278_U57 , R2278_U140 );
not NOT1_6003 ( R2278_U348 , R2278_U110 );
nand NAND2_6004 ( R2278_U349 , R2278_U188 , R2278_U73 );
nand NAND2_6005 ( R2278_U350 , R2278_U191 , R2278_U72 );
nand NAND2_6006 ( R2278_U351 , R2278_U184 , R2278_U76 );
nand NAND2_6007 ( R2278_U352 , R2278_U192 , R2278_U75 );
nand NAND2_6008 ( R2278_U353 , R2278_U198 , R2278_U79 );
nand NAND2_6009 ( R2278_U354 , R2278_U199 , R2278_U78 );
nand NAND2_6010 ( R2278_U355 , R2278_U196 , R2278_U82 );
nand NAND2_6011 ( R2278_U356 , R2278_U200 , R2278_U81 );
nand NAND2_6012 ( R2278_U357 , R2278_U194 , R2278_U85 );
nand NAND2_6013 ( R2278_U358 , R2278_U201 , R2278_U84 );
nand NAND2_6014 ( R2278_U359 , R2278_U177 , R2278_U88 );
nand NAND2_6015 ( R2278_U360 , R2278_U202 , R2278_U87 );
nand NAND2_6016 ( R2278_U361 , R2278_U174 , R2278_U91 );
nand NAND2_6017 ( R2278_U362 , R2278_U203 , R2278_U90 );
nand NAND2_6018 ( R2278_U363 , U2769 , R2278_U94 );
nand NAND2_6019 ( R2278_U364 , INSTADDRPOINTER_REG_31_ , R2278_U93 );
not NOT1_6020 ( R2278_U365 , R2278_U62 );
nand NAND2_6021 ( R2278_U366 , R2278_U261 , R2278_U365 );
nand NAND2_6022 ( R2278_U367 , R2278_U62 , R2278_U95 );
nand NAND2_6023 ( R2278_U368 , U2770 , R2278_U21 );
nand NAND2_6024 ( R2278_U369 , INSTADDRPOINTER_REG_30_ , R2278_U22 );
not NOT1_6025 ( R2278_U370 , R2278_U63 );
nand NAND2_6026 ( R2278_U371 , R2278_U258 , R2278_U370 );
nand NAND2_6027 ( R2278_U372 , R2278_U63 , R2278_U97 );
nand NAND2_6028 ( R2278_U373 , R2278_U171 , R2278_U100 );
nand NAND2_6029 ( R2278_U374 , R2278_U262 , R2278_U99 );
nand NAND2_6030 ( R2278_U375 , U2770 , R2278_U32 );
nand NAND2_6031 ( R2278_U376 , INSTADDRPOINTER_REG_29_ , R2278_U33 );
not NOT1_6032 ( R2278_U377 , R2278_U64 );
nand NAND2_6033 ( R2278_U378 , R2278_U255 , R2278_U377 );
nand NAND2_6034 ( R2278_U379 , R2278_U64 , R2278_U102 );
nand NAND2_6035 ( R2278_U380 , U2770 , R2278_U34 );
nand NAND2_6036 ( R2278_U381 , INSTADDRPOINTER_REG_28_ , R2278_U35 );
not NOT1_6037 ( R2278_U382 , R2278_U65 );
nand NAND2_6038 ( R2278_U383 , R2278_U252 , R2278_U382 );
nand NAND2_6039 ( R2278_U384 , R2278_U65 , R2278_U104 );
nand NAND2_6040 ( R2278_U385 , R2278_U249 , R2278_U107 );
nand NAND2_6041 ( R2278_U386 , R2278_U263 , R2278_U106 );
nand NAND2_6042 ( R2278_U387 , R2278_U264 , R2278_U110 );
nand NAND2_6043 ( R2278_U388 , R2278_U348 , R2278_U109 );
nand NAND2_6044 ( R2278_U389 , R2278_U244 , R2278_U113 );
nand NAND2_6045 ( R2278_U390 , R2278_U265 , R2278_U112 );
nand NAND2_6046 ( R2278_U391 , R2278_U241 , R2278_U116 );
nand NAND2_6047 ( R2278_U392 , R2278_U266 , R2278_U115 );
nand NAND2_6048 ( R2278_U393 , R2278_U239 , R2278_U119 );
nand NAND2_6049 ( R2278_U394 , R2278_U267 , R2278_U118 );
nand NAND2_6050 ( R2278_U395 , R2278_U237 , R2278_U122 );
nand NAND2_6051 ( R2278_U396 , R2278_U268 , R2278_U121 );
nand NAND2_6052 ( R2278_U397 , R2278_U234 , R2278_U125 );
nand NAND2_6053 ( R2278_U398 , R2278_U269 , R2278_U124 );
nand NAND2_6054 ( R2278_U399 , R2278_U270 , R2278_U128 );
nand NAND2_6055 ( R2278_U400 , R2278_U346 , R2278_U127 );
nand NAND2_6056 ( R2278_U401 , R2278_U161 , R2278_U130 );
nand NAND2_6057 ( R2278_U402 , R2278_U271 , R2278_U19 );
nand NAND2_6058 ( R2278_U403 , R2278_U272 , R2278_U132 );
nand NAND2_6059 ( R2278_U404 , R2278_U344 , R2278_U131 );
nand NAND2_6060 ( R2278_U405 , R2278_U273 , R2278_U135 );
nand NAND2_6061 ( R2278_U406 , R2278_U342 , R2278_U134 );
nand NAND2_6062 ( R2278_U407 , R2278_U274 , R2278_U138 );
nand NAND2_6063 ( R2278_U408 , R2278_U340 , R2278_U137 );
nand NAND2_6064 ( R2278_U409 , R2278_U224 , R2278_U141 );
nand NAND2_6065 ( R2278_U410 , R2278_U275 , R2278_U140 );
nand NAND2_6066 ( R2278_U411 , R2278_U281 , R2278_U144 );
nand NAND2_6067 ( R2278_U412 , R2278_U282 , R2278_U143 );
nand NAND2_6068 ( R2278_U413 , R2278_U279 , R2278_U147 );
nand NAND2_6069 ( R2278_U414 , R2278_U283 , R2278_U146 );
nand NAND2_6070 ( R2278_U415 , R2278_U277 , R2278_U150 );
nand NAND2_6071 ( R2278_U416 , R2278_U284 , R2278_U149 );
nand NAND2_6072 ( R2278_U417 , R2278_U220 , R2278_U153 );
nand NAND2_6073 ( R2278_U418 , R2278_U285 , R2278_U152 );
nand NAND2_6074 ( R2278_U419 , R2278_U289 , R2278_U156 );
nand NAND2_6075 ( R2278_U420 , R2278_U290 , R2278_U155 );
nand NAND2_6076 ( R2278_U421 , R2278_U287 , R2278_U159 );
nand NAND2_6077 ( R2278_U422 , R2278_U291 , R2278_U158 );
and AND4_6078 ( R2358_U5 , R2358_U293 , R2358_U285 , R2358_U282 , R2358_U281 );
and AND2_6079 ( R2358_U6 , R2358_U329 , R2358_U325 );
and AND3_6080 ( R2358_U7 , R2358_U6 , R2358_U324 , R2358_U141 );
and AND2_6081 ( R2358_U8 , R2358_U135 , R2358_U5 );
and AND2_6082 ( R2358_U9 , R2358_U296 , R2358_U294 );
and AND2_6083 ( R2358_U10 , R2358_U304 , R2358_U253 );
and AND2_6084 ( R2358_U11 , R2358_U303 , R2358_U301 );
and AND2_6085 ( R2358_U12 , R2358_U8 , R2358_U7 );
and AND2_6086 ( R2358_U13 , R2358_U528 , R2358_U527 );
and AND2_6087 ( R2358_U14 , R2358_U379 , R2358_U378 );
and AND2_6088 ( R2358_U15 , R2358_U376 , R2358_U374 );
and AND2_6089 ( R2358_U16 , R2358_U370 , R2358_U367 );
and AND2_6090 ( R2358_U17 , R2358_U360 , R2358_U359 );
and AND2_6091 ( R2358_U18 , R2358_U354 , R2358_U352 );
and AND2_6092 ( R2358_U19 , R2358_U336 , R2358_U335 );
and AND2_6093 ( R2358_U20 , R2358_U276 , R2358_U274 );
and AND2_6094 ( R2358_U21 , R2358_U266 , R2358_U262 );
not NOT1_6095 ( R2358_U22 , U2352 );
not NOT1_6096 ( R2358_U23 , U2643 );
not NOT1_6097 ( R2358_U24 , U2644 );
not NOT1_6098 ( R2358_U25 , U2645 );
not NOT1_6099 ( R2358_U26 , U2646 );
not NOT1_6100 ( R2358_U27 , U2649 );
not NOT1_6101 ( R2358_U28 , U2648 );
not NOT1_6102 ( R2358_U29 , U2650 );
not NOT1_6103 ( R2358_U30 , U2647 );
nand NAND2_6104 ( R2358_U31 , U2644 , R2358_U77 );
not NOT1_6105 ( R2358_U32 , U2642 );
not NOT1_6106 ( R2358_U33 , U2641 );
nand NAND2_6107 ( R2358_U34 , R2358_U246 , R2358_U259 );
not NOT1_6108 ( R2358_U35 , U2620 );
not NOT1_6109 ( R2358_U36 , U2625 );
not NOT1_6110 ( R2358_U37 , U2624 );
not NOT1_6111 ( R2358_U38 , U2622 );
not NOT1_6112 ( R2358_U39 , U2623 );
not NOT1_6113 ( R2358_U40 , U2621 );
not NOT1_6114 ( R2358_U41 , U2626 );
not NOT1_6115 ( R2358_U42 , U2627 );
not NOT1_6116 ( R2358_U43 , U2628 );
not NOT1_6117 ( R2358_U44 , U2629 );
not NOT1_6118 ( R2358_U45 , U2630 );
nand NAND2_6119 ( R2358_U46 , U2630 , R2358_U78 );
not NOT1_6120 ( R2358_U47 , U2639 );
not NOT1_6121 ( R2358_U48 , U2640 );
nand NAND2_6122 ( R2358_U49 , U2642 , R2358_U490 );
not NOT1_6123 ( R2358_U50 , U2637 );
nand NAND2_6124 ( R2358_U51 , U2637 , R2358_U80 );
not NOT1_6125 ( R2358_U52 , U2638 );
nand NAND2_6126 ( R2358_U53 , U2638 , R2358_U531 );
not NOT1_6127 ( R2358_U54 , U2636 );
nand NAND2_6128 ( R2358_U55 , R2358_U142 , R2358_U9 );
not NOT1_6129 ( R2358_U56 , U2631 );
not NOT1_6130 ( R2358_U57 , U2632 );
not NOT1_6131 ( R2358_U58 , U2633 );
nand NAND2_6132 ( R2358_U59 , U2633 , R2358_U607 );
not NOT1_6133 ( R2358_U60 , U2634 );
nand NAND2_6134 ( R2358_U61 , U2634 , R2358_U601 );
nand NAND2_6135 ( R2358_U62 , R2358_U438 , R2358_U320 );
nand NAND2_6136 ( R2358_U63 , R2358_U280 , R2358_U291 );
nand NAND2_6137 ( R2358_U64 , R2358_U233 , R2358_U270 );
nand NAND2_6138 ( R2358_U65 , R2358_U64 , R2358_U229 );
nand NAND2_6139 ( R2358_U66 , R2358_U417 , R2358_U316 );
nand NAND3_6140 ( R2358_U67 , R2358_U410 , R2358_U219 , R2358_U146 );
nand NAND2_6141 ( R2358_U68 , R2358_U418 , R2358_U416 );
nand NAND3_6142 ( R2358_U69 , R2358_U407 , R2358_U295 , R2358_U408 );
nand NAND2_6143 ( R2358_U70 , R2358_U313 , R2358_U67 );
not NOT1_6144 ( R2358_U71 , U2635 );
nand NAND2_6145 ( R2358_U72 , R2358_U51 , R2358_U364 );
nand NAND2_6146 ( R2358_U73 , R2358_U414 , R2358_U305 );
nand NAND2_6147 ( R2358_U74 , R2358_U423 , R2358_U413 );
nand NAND2_6148 ( R2358_U75 , R2358_U74 , R2358_U301 );
nand NAND2_6149 ( R2358_U76 , R2358_U441 , R2358_U440 );
nand NAND2_6150 ( R2358_U77 , R2358_U454 , R2358_U453 );
nand NAND2_6151 ( R2358_U78 , R2358_U552 , R2358_U551 );
nand NAND2_6152 ( R2358_U79 , R2358_U520 , R2358_U519 );
nand NAND2_6153 ( R2358_U80 , R2358_U525 , R2358_U524 );
nand NAND2_6154 ( R2358_U81 , R2358_U533 , R2358_U532 );
nand NAND2_6155 ( R2358_U82 , R2358_U654 , R2358_U653 );
nand NAND2_6156 ( R2358_U83 , R2358_U492 , R2358_U491 );
and AND2_6157 ( R2358_U84 , R2358_U49 , R2358_U253 );
nand NAND2_6158 ( R2358_U85 , R2358_U494 , R2358_U493 );
nand NAND2_6159 ( R2358_U86 , R2358_U499 , R2358_U498 );
and AND2_6160 ( R2358_U87 , R2358_U246 , R2358_U243 );
nand NAND2_6161 ( R2358_U88 , R2358_U501 , R2358_U500 );
and AND2_6162 ( R2358_U89 , R2358_U247 , R2358_U244 );
nand NAND2_6163 ( R2358_U90 , R2358_U503 , R2358_U502 );
nand NAND2_6164 ( R2358_U91 , R2358_U609 , R2358_U608 );
and AND2_6165 ( R2358_U92 , R2358_U278 , R2358_U277 );
nand NAND2_6166 ( R2358_U93 , R2358_U611 , R2358_U610 );
and AND2_6167 ( R2358_U94 , R2358_U280 , R2358_U279 );
nand NAND2_6168 ( R2358_U95 , R2358_U613 , R2358_U612 );
and AND2_6169 ( R2358_U96 , R2358_U288 , R2358_U281 );
nand NAND2_6170 ( R2358_U97 , R2358_U615 , R2358_U614 );
and AND2_6171 ( R2358_U98 , R2358_U289 , R2358_U282 );
nand NAND2_6172 ( R2358_U99 , R2358_U617 , R2358_U616 );
and AND2_6173 ( R2358_U100 , R2358_U285 , R2358_U284 );
nand NAND2_6174 ( R2358_U101 , R2358_U619 , R2358_U618 );
and AND2_6175 ( R2358_U102 , R2358_U293 , R2358_U283 );
nand NAND2_6176 ( R2358_U103 , R2358_U621 , R2358_U620 );
and AND2_6177 ( R2358_U104 , R2358_U320 , R2358_U319 );
nand NAND2_6178 ( R2358_U105 , R2358_U623 , R2358_U622 );
and AND2_6179 ( R2358_U106 , R2358_U322 , R2358_U321 );
nand NAND2_6180 ( R2358_U107 , R2358_U625 , R2358_U624 );
and AND2_6181 ( R2358_U108 , R2358_U324 , R2358_U323 );
nand NAND2_6182 ( R2358_U109 , R2358_U627 , R2358_U626 );
nand NAND2_6183 ( R2358_U110 , R2358_U632 , R2358_U631 );
and AND2_6184 ( R2358_U111 , R2358_U233 , R2358_U232 );
nand NAND2_6185 ( R2358_U112 , R2358_U634 , R2358_U633 );
and AND2_6186 ( R2358_U113 , R2358_U317 , R2358_U316 );
nand NAND2_6187 ( R2358_U114 , R2358_U636 , R2358_U635 );
and AND2_6188 ( R2358_U115 , R2358_U295 , R2358_U294 );
nand NAND2_6189 ( R2358_U116 , R2358_U638 , R2358_U637 );
and AND2_6190 ( R2358_U117 , R2358_U59 , R2358_U296 );
nand NAND2_6191 ( R2358_U118 , R2358_U640 , R2358_U639 );
nand NAND2_6192 ( R2358_U119 , R2358_U645 , R2358_U644 );
nand NAND2_6193 ( R2358_U120 , R2358_U650 , R2358_U649 );
and AND2_6194 ( R2358_U121 , R2358_U310 , R2358_U53 );
nand NAND2_6195 ( R2358_U122 , R2358_U652 , R2358_U651 );
and AND2_6196 ( R2358_U123 , R2358_U235 , R2358_U232 );
and AND2_6197 ( R2358_U124 , R2358_U231 , R2358_U229 );
and AND2_6198 ( R2358_U125 , R2358_U244 , R2358_U243 );
and AND2_6199 ( R2358_U126 , R2358_U249 , R2358_U245 );
and AND2_6200 ( R2358_U127 , R2358_U245 , R2358_U222 );
and AND2_6201 ( R2358_U128 , R2358_U265 , R2358_U31 );
and AND2_6202 ( R2358_U129 , R2358_U231 , R2358_U230 );
and AND2_6203 ( R2358_U130 , R2358_U285 , R2358_U282 );
and AND2_6204 ( R2358_U131 , R2358_U288 , R2358_U289 );
and AND2_6205 ( R2358_U132 , R2358_U281 , R2358_U279 );
and AND2_6206 ( R2358_U133 , R2358_U326 , R2358_U323 );
and AND2_6207 ( R2358_U134 , R2358_U322 , R2358_U319 );
and AND2_6208 ( R2358_U135 , R2358_U279 , R2358_U277 );
and AND2_6209 ( R2358_U136 , R2358_U11 , R2358_U10 );
and AND2_6210 ( R2358_U137 , R2358_U432 , R2358_U425 );
and AND2_6211 ( R2358_U138 , R2358_U310 , R2358_U224 );
and AND2_6212 ( R2358_U139 , R2358_U415 , R2358_U311 );
and AND2_6213 ( R2358_U140 , R2358_U420 , R2358_U411 );
and AND2_6214 ( R2358_U141 , R2358_U322 , R2358_U319 );
and AND2_6215 ( R2358_U142 , R2358_U317 , R2358_U313 );
and AND2_6216 ( R2358_U143 , R2358_U12 , R2358_U426 );
and AND2_6217 ( R2358_U144 , R2358_U402 , R2358_U278 );
and AND3_6218 ( R2358_U145 , R2358_U144 , R2358_U406 , R2358_U430 );
and AND2_6219 ( R2358_U146 , R2358_U420 , R2358_U411 );
and AND2_6220 ( R2358_U147 , R2358_U313 , R2358_U317 );
and AND2_6221 ( R2358_U148 , R2358_U7 , R2358_U149 );
and AND2_6222 ( R2358_U149 , R2358_U9 , R2358_U147 );
and AND2_6223 ( R2358_U150 , R2358_U422 , R2358_U439 );
and AND2_6224 ( R2358_U151 , R2358_U5 , R2358_U279 );
and AND3_6225 ( R2358_U152 , R2358_U285 , R2358_U282 , R2358_U293 );
and AND2_6226 ( R2358_U153 , R2358_U289 , R2358_U287 );
and AND2_6227 ( R2358_U154 , R2358_U284 , R2358_U283 );
and AND2_6228 ( R2358_U155 , R2358_U156 , R2358_U434 );
and AND2_6229 ( R2358_U156 , R2358_U6 , R2358_U324 );
and AND2_6230 ( R2358_U157 , R2358_U418 , R2358_U46 );
and AND2_6231 ( R2358_U158 , R2358_U6 , R2358_U326 );
and AND2_6232 ( R2358_U159 , R2358_U313 , R2358_U9 );
and AND3_6233 ( R2358_U160 , R2358_U299 , R2358_U224 , R2358_U300 );
and AND2_6234 ( R2358_U161 , R2358_U369 , R2358_U227 );
and AND2_6235 ( R2358_U162 , R2358_U303 , R2358_U302 );
and AND2_6236 ( R2358_U163 , R2358_U375 , R2358_U307 );
not NOT1_6237 ( R2358_U164 , U2612 );
and AND2_6238 ( R2358_U165 , R2358_U444 , R2358_U443 );
not NOT1_6239 ( R2358_U166 , U2610 );
not NOT1_6240 ( R2358_U167 , U2609 );
not NOT1_6241 ( R2358_U168 , U2667 );
not NOT1_6242 ( R2358_U169 , U2668 );
not NOT1_6243 ( R2358_U170 , U2670 );
not NOT1_6244 ( R2358_U171 , U2671 );
not NOT1_6245 ( R2358_U172 , U2672 );
not NOT1_6246 ( R2358_U173 , U2669 );
not NOT1_6247 ( R2358_U174 , U2611 );
nand NAND2_6248 ( R2358_U175 , R2358_U49 , R2358_U255 );
nand NAND3_6249 ( R2358_U176 , R2358_U251 , R2358_U250 , R2358_U126 );
nand NAND2_6250 ( R2358_U177 , R2358_U247 , R2358_U257 );
nand NAND2_6251 ( R2358_U178 , R2358_U230 , R2358_U240 );
not NOT1_6252 ( R2358_U179 , U2651 );
and AND2_6253 ( R2358_U180 , R2358_U505 , R2358_U504 );
not NOT1_6254 ( R2358_U181 , U2613 );
not NOT1_6255 ( R2358_U182 , U2614 );
not NOT1_6256 ( R2358_U183 , U2617 );
not NOT1_6257 ( R2358_U184 , U2615 );
not NOT1_6258 ( R2358_U185 , U2616 );
not NOT1_6259 ( R2358_U186 , U2618 );
not NOT1_6260 ( R2358_U187 , U2664 );
not NOT1_6261 ( R2358_U188 , U2665 );
not NOT1_6262 ( R2358_U189 , U2666 );
not NOT1_6263 ( R2358_U190 , U2663 );
not NOT1_6264 ( R2358_U191 , U2658 );
not NOT1_6265 ( R2358_U192 , U2659 );
not NOT1_6266 ( R2358_U193 , U2660 );
not NOT1_6267 ( R2358_U194 , U2661 );
not NOT1_6268 ( R2358_U195 , U2662 );
not NOT1_6269 ( R2358_U196 , U2654 );
not NOT1_6270 ( R2358_U197 , U2655 );
not NOT1_6271 ( R2358_U198 , U2656 );
not NOT1_6272 ( R2358_U199 , U2657 );
not NOT1_6273 ( R2358_U200 , U2652 );
not NOT1_6274 ( R2358_U201 , U2653 );
nand NAND2_6275 ( R2358_U202 , R2358_U145 , R2358_U429 );
nand NAND2_6276 ( R2358_U203 , R2358_U292 , R2358_U332 );
nand NAND2_6277 ( R2358_U204 , R2358_U338 , R2358_U337 );
nand NAND2_6278 ( R2358_U205 , R2358_U153 , R2358_U340 );
nand NAND2_6279 ( R2358_U206 , R2358_U344 , R2358_U285 );
nand NAND2_6280 ( R2358_U207 , R2358_U283 , R2358_U342 );
nand NAND2_6281 ( R2358_U208 , R2358_U150 , R2358_U421 );
nand NAND2_6282 ( R2358_U209 , R2358_U321 , R2358_U347 );
nand NAND2_6283 ( R2358_U210 , R2358_U345 , R2358_U437 );
nand NAND2_6284 ( R2358_U211 , R2358_U350 , R2358_U325 );
nand NAND2_6285 ( R2358_U212 , R2358_U236 , R2358_U268 );
nand NAND2_6286 ( R2358_U213 , R2358_U412 , R2358_U409 );
nand NAND2_6287 ( R2358_U214 , R2358_U356 , R2358_U59 );
nand NAND2_6288 ( R2358_U215 , R2358_U61 , R2358_U70 );
nand NAND2_6289 ( R2358_U216 , R2358_U53 , R2358_U361 );
nand NAND2_6290 ( R2358_U217 , R2358_U137 , R2358_U431 );
nand NAND2_6291 ( R2358_U218 , R2358_U236 , R2358_U235 );
nand NAND3_6292 ( R2358_U219 , R2358_U138 , R2358_U217 , R2358_U139 );
not NOT1_6293 ( R2358_U220 , R2358_U211 );
not NOT1_6294 ( R2358_U221 , R2358_U206 );
nand NAND2_6295 ( R2358_U222 , R2358_U404 , R2358_U403 );
not NOT1_6296 ( R2358_U223 , R2358_U51 );
nand NAND2_6297 ( R2358_U224 , R2358_U521 , R2358_U54 );
not NOT1_6298 ( R2358_U225 , R2358_U46 );
nand NAND2_6299 ( R2358_U226 , R2358_U349 , R2358_U329 );
nand NAND2_6300 ( R2358_U227 , U2636 , R2358_U79 );
not NOT1_6301 ( R2358_U228 , R2358_U31 );
nand NAND3_6302 ( R2358_U229 , R2358_U480 , R2358_U479 , R2358_U28 );
nand NAND2_6303 ( R2358_U230 , U2647 , R2358_U485 );
nand NAND3_6304 ( R2358_U231 , R2358_U482 , R2358_U481 , R2358_U30 );
nand NAND3_6305 ( R2358_U232 , R2358_U476 , R2358_U475 , R2358_U27 );
nand NAND2_6306 ( R2358_U233 , U2649 , R2358_U471 );
nand NAND2_6307 ( R2358_U234 , U2648 , R2358_U468 );
nand NAND3_6308 ( R2358_U235 , R2358_U478 , R2358_U477 , R2358_U29 );
nand NAND2_6309 ( R2358_U236 , U2650 , R2358_U474 );
nand NAND2_6310 ( R2358_U237 , R2358_U236 , R2358_U22 );
nand NAND2_6311 ( R2358_U238 , R2358_U123 , R2358_U237 );
nand NAND3_6312 ( R2358_U239 , R2358_U238 , R2358_U233 , R2358_U234 );
nand NAND2_6313 ( R2358_U240 , R2358_U124 , R2358_U239 );
not NOT1_6314 ( R2358_U241 , R2358_U178 );
nand NAND3_6315 ( R2358_U242 , R2358_U452 , R2358_U451 , R2358_U23 );
nand NAND3_6316 ( R2358_U243 , R2358_U463 , R2358_U462 , R2358_U25 );
nand NAND3_6317 ( R2358_U244 , R2358_U465 , R2358_U464 , R2358_U26 );
nand NAND2_6318 ( R2358_U245 , U2643 , R2358_U450 );
nand NAND2_6319 ( R2358_U246 , U2645 , R2358_U458 );
nand NAND2_6320 ( R2358_U247 , U2646 , R2358_U461 );
nand NAND2_6321 ( R2358_U248 , R2358_U247 , R2358_U246 );
nand NAND3_6322 ( R2358_U249 , R2358_U243 , R2358_U248 , R2358_U222 );
nand NAND3_6323 ( R2358_U250 , R2358_U178 , R2358_U125 , R2358_U222 );
nand NAND2_6324 ( R2358_U251 , R2358_U228 , R2358_U242 );
not NOT1_6325 ( R2358_U252 , R2358_U176 );
nand NAND3_6326 ( R2358_U253 , R2358_U487 , R2358_U486 , R2358_U32 );
not NOT1_6327 ( R2358_U254 , R2358_U49 );
nand NAND2_6328 ( R2358_U255 , R2358_U253 , R2358_U176 );
not NOT1_6329 ( R2358_U256 , R2358_U175 );
nand NAND2_6330 ( R2358_U257 , R2358_U244 , R2358_U178 );
not NOT1_6331 ( R2358_U258 , R2358_U177 );
nand NAND2_6332 ( R2358_U259 , R2358_U177 , R2358_U243 );
not NOT1_6333 ( R2358_U260 , R2358_U34 );
nand NAND2_6334 ( R2358_U261 , R2358_U260 , R2358_U31 );
nand NAND2_6335 ( R2358_U262 , R2358_U127 , R2358_U261 );
nand NAND2_6336 ( R2358_U263 , R2358_U455 , R2358_U24 );
nand NAND2_6337 ( R2358_U264 , R2358_U263 , R2358_U34 );
nand NAND2_6338 ( R2358_U265 , R2358_U245 , R2358_U242 );
nand NAND2_6339 ( R2358_U266 , R2358_U128 , R2358_U264 );
nand NAND2_6340 ( R2358_U267 , R2358_U455 , R2358_U24 );
nand NAND2_6341 ( R2358_U268 , U2352 , R2358_U235 );
not NOT1_6342 ( R2358_U269 , R2358_U212 );
nand NAND2_6343 ( R2358_U270 , R2358_U212 , R2358_U232 );
not NOT1_6344 ( R2358_U271 , R2358_U64 );
not NOT1_6345 ( R2358_U272 , R2358_U65 );
nand NAND2_6346 ( R2358_U273 , R2358_U65 , R2358_U234 );
nand NAND2_6347 ( R2358_U274 , R2358_U129 , R2358_U273 );
nand NAND2_6348 ( R2358_U275 , R2358_U231 , R2358_U230 );
nand NAND3_6349 ( R2358_U276 , R2358_U65 , R2358_U234 , R2358_U275 );
nand NAND3_6350 ( R2358_U277 , R2358_U563 , R2358_U562 , R2358_U35 );
nand NAND2_6351 ( R2358_U278 , U2620 , R2358_U580 );
nand NAND3_6352 ( R2358_U279 , R2358_U565 , R2358_U564 , R2358_U40 );
nand NAND2_6353 ( R2358_U280 , U2621 , R2358_U595 );
nand NAND3_6354 ( R2358_U281 , R2358_U555 , R2358_U554 , R2358_U38 );
nand NAND3_6355 ( R2358_U282 , R2358_U557 , R2358_U556 , R2358_U39 );
nand NAND2_6356 ( R2358_U283 , U2625 , R2358_U583 );
nand NAND2_6357 ( R2358_U284 , U2624 , R2358_U586 );
nand NAND3_6358 ( R2358_U285 , R2358_U559 , R2358_U558 , R2358_U37 );
nand NAND2_6359 ( R2358_U286 , R2358_U284 , R2358_U283 );
nand NAND2_6360 ( R2358_U287 , R2358_U130 , R2358_U286 );
nand NAND2_6361 ( R2358_U288 , U2622 , R2358_U592 );
nand NAND2_6362 ( R2358_U289 , U2623 , R2358_U589 );
nand NAND2_6363 ( R2358_U290 , R2358_U131 , R2358_U287 );
nand NAND2_6364 ( R2358_U291 , R2358_U132 , R2358_U290 );
not NOT1_6365 ( R2358_U292 , R2358_U63 );
nand NAND3_6366 ( R2358_U293 , R2358_U561 , R2358_U560 , R2358_U36 );
nand NAND3_6367 ( R2358_U294 , R2358_U536 , R2358_U535 , R2358_U57 );
nand NAND2_6368 ( R2358_U295 , U2632 , R2358_U604 );
nand NAND3_6369 ( R2358_U296 , R2358_U538 , R2358_U537 , R2358_U58 );
not NOT1_6370 ( R2358_U297 , R2358_U59 );
not NOT1_6371 ( R2358_U298 , R2358_U61 );
nand NAND2_6372 ( R2358_U299 , R2358_U13 , R2358_U71 );
nand NAND2_6373 ( R2358_U300 , U2635 , R2358_U81 );
nand NAND3_6374 ( R2358_U301 , R2358_U510 , R2358_U509 , R2358_U48 );
nand NAND2_6375 ( R2358_U302 , U2639 , R2358_U515 );
nand NAND3_6376 ( R2358_U303 , R2358_U512 , R2358_U511 , R2358_U47 );
nand NAND2_6377 ( R2358_U304 , R2358_U442 , R2358_U33 );
nand NAND2_6378 ( R2358_U305 , U2641 , R2358_U76 );
not NOT1_6379 ( R2358_U306 , R2358_U74 );
nand NAND2_6380 ( R2358_U307 , U2640 , R2358_U518 );
not NOT1_6381 ( R2358_U308 , R2358_U217 );
not NOT1_6382 ( R2358_U309 , R2358_U53 );
nand NAND3_6383 ( R2358_U310 , R2358_U523 , R2358_U522 , R2358_U52 );
nand NAND2_6384 ( R2358_U311 , R2358_U526 , R2358_U50 );
not NOT1_6385 ( R2358_U312 , R2358_U67 );
nand NAND3_6386 ( R2358_U313 , R2358_U540 , R2358_U539 , R2358_U60 );
not NOT1_6387 ( R2358_U314 , R2358_U70 );
not NOT1_6388 ( R2358_U315 , R2358_U213 );
nand NAND2_6389 ( R2358_U316 , U2631 , R2358_U598 );
nand NAND3_6390 ( R2358_U317 , R2358_U542 , R2358_U541 , R2358_U56 );
not NOT1_6391 ( R2358_U318 , R2358_U68 );
nand NAND3_6392 ( R2358_U319 , R2358_U544 , R2358_U543 , R2358_U41 );
nand NAND2_6393 ( R2358_U320 , U2626 , R2358_U568 );
nand NAND2_6394 ( R2358_U321 , U2627 , R2358_U571 );
nand NAND3_6395 ( R2358_U322 , R2358_U546 , R2358_U545 , R2358_U42 );
nand NAND2_6396 ( R2358_U323 , U2628 , R2358_U574 );
nand NAND3_6397 ( R2358_U324 , R2358_U548 , R2358_U547 , R2358_U43 );
nand NAND3_6398 ( R2358_U325 , R2358_U550 , R2358_U549 , R2358_U44 );
nand NAND2_6399 ( R2358_U326 , U2629 , R2358_U577 );
nand NAND2_6400 ( R2358_U327 , R2358_U225 , R2358_U325 );
nand NAND2_6401 ( R2358_U328 , R2358_U437 , R2358_U321 );
nand NAND2_6402 ( R2358_U329 , R2358_U553 , R2358_U45 );
not NOT1_6403 ( R2358_U330 , R2358_U202 );
not NOT1_6404 ( R2358_U331 , R2358_U208 );
nand NAND2_6405 ( R2358_U332 , R2358_U151 , R2358_U208 );
not NOT1_6406 ( R2358_U333 , R2358_U203 );
nand NAND2_6407 ( R2358_U334 , R2358_U234 , R2358_U229 );
nand NAND2_6408 ( R2358_U335 , R2358_U271 , R2358_U334 );
nand NAND2_6409 ( R2358_U336 , R2358_U272 , R2358_U234 );
nand NAND2_6410 ( R2358_U337 , R2358_U290 , R2358_U281 );
nand NAND2_6411 ( R2358_U338 , R2358_U5 , R2358_U208 );
not NOT1_6412 ( R2358_U339 , R2358_U204 );
nand NAND2_6413 ( R2358_U340 , R2358_U152 , R2358_U208 );
not NOT1_6414 ( R2358_U341 , R2358_U205 );
nand NAND2_6415 ( R2358_U342 , R2358_U208 , R2358_U293 );
not NOT1_6416 ( R2358_U343 , R2358_U207 );
nand NAND2_6417 ( R2358_U344 , R2358_U154 , R2358_U342 );
nand NAND2_6418 ( R2358_U345 , R2358_U433 , R2358_U155 );
not NOT1_6419 ( R2358_U346 , R2358_U210 );
nand NAND2_6420 ( R2358_U347 , R2358_U210 , R2358_U322 );
not NOT1_6421 ( R2358_U348 , R2358_U209 );
nand NAND2_6422 ( R2358_U349 , R2358_U157 , R2358_U416 );
nand NAND2_6423 ( R2358_U350 , R2358_U326 , R2358_U226 );
nand NAND2_6424 ( R2358_U351 , R2358_U318 , R2358_U46 );
nand NAND2_6425 ( R2358_U352 , R2358_U158 , R2358_U351 );
nand NAND2_6426 ( R2358_U353 , R2358_U326 , R2358_U325 );
nand NAND2_6427 ( R2358_U354 , R2358_U226 , R2358_U353 );
not NOT1_6428 ( R2358_U355 , R2358_U215 );
nand NAND2_6429 ( R2358_U356 , R2358_U215 , R2358_U296 );
not NOT1_6430 ( R2358_U357 , R2358_U214 );
nand NAND2_6431 ( R2358_U358 , R2358_U313 , R2358_U61 );
nand NAND2_6432 ( R2358_U359 , R2358_U312 , R2358_U358 );
nand NAND2_6433 ( R2358_U360 , R2358_U314 , R2358_U61 );
nand NAND2_6434 ( R2358_U361 , R2358_U310 , R2358_U217 );
not NOT1_6435 ( R2358_U362 , R2358_U216 );
nand NAND2_6436 ( R2358_U363 , R2358_U526 , R2358_U50 );
nand NAND2_6437 ( R2358_U364 , R2358_U363 , R2358_U216 );
not NOT1_6438 ( R2358_U365 , R2358_U72 );
nand NAND2_6439 ( R2358_U366 , R2358_U365 , R2358_U227 );
nand NAND2_6440 ( R2358_U367 , R2358_U160 , R2358_U366 );
nand NAND2_6441 ( R2358_U368 , R2358_U72 , R2358_U224 );
nand NAND2_6442 ( R2358_U369 , R2358_U300 , R2358_U299 );
nand NAND2_6443 ( R2358_U370 , R2358_U161 , R2358_U368 );
nand NAND2_6444 ( R2358_U371 , R2358_U526 , R2358_U50 );
not NOT1_6445 ( R2358_U372 , R2358_U75 );
nand NAND2_6446 ( R2358_U373 , R2358_U75 , R2358_U307 );
nand NAND2_6447 ( R2358_U374 , R2358_U162 , R2358_U373 );
nand NAND2_6448 ( R2358_U375 , R2358_U303 , R2358_U302 );
nand NAND2_6449 ( R2358_U376 , R2358_U163 , R2358_U75 );
nand NAND2_6450 ( R2358_U377 , R2358_U307 , R2358_U301 );
nand NAND2_6451 ( R2358_U378 , R2358_U306 , R2358_U377 );
nand NAND2_6452 ( R2358_U379 , R2358_U372 , R2358_U307 );
not NOT1_6453 ( R2358_U380 , R2358_U218 );
nand NAND2_6454 ( R2358_U381 , R2358_U49 , R2358_U253 );
nand NAND2_6455 ( R2358_U382 , R2358_U267 , R2358_U31 );
nand NAND2_6456 ( R2358_U383 , R2358_U246 , R2358_U243 );
nand NAND2_6457 ( R2358_U384 , R2358_U247 , R2358_U244 );
nand NAND2_6458 ( R2358_U385 , R2358_U278 , R2358_U277 );
nand NAND2_6459 ( R2358_U386 , R2358_U280 , R2358_U279 );
nand NAND2_6460 ( R2358_U387 , R2358_U288 , R2358_U281 );
nand NAND2_6461 ( R2358_U388 , R2358_U289 , R2358_U282 );
nand NAND2_6462 ( R2358_U389 , R2358_U285 , R2358_U284 );
nand NAND2_6463 ( R2358_U390 , R2358_U293 , R2358_U283 );
nand NAND2_6464 ( R2358_U391 , R2358_U320 , R2358_U319 );
nand NAND2_6465 ( R2358_U392 , R2358_U322 , R2358_U321 );
nand NAND2_6466 ( R2358_U393 , R2358_U324 , R2358_U323 );
nand NAND2_6467 ( R2358_U394 , R2358_U329 , R2358_U46 );
nand NAND2_6468 ( R2358_U395 , R2358_U233 , R2358_U232 );
nand NAND2_6469 ( R2358_U396 , R2358_U317 , R2358_U316 );
nand NAND2_6470 ( R2358_U397 , R2358_U295 , R2358_U294 );
nand NAND2_6471 ( R2358_U398 , R2358_U59 , R2358_U296 );
nand NAND2_6472 ( R2358_U399 , R2358_U227 , R2358_U224 );
nand NAND2_6473 ( R2358_U400 , R2358_U371 , R2358_U51 );
nand NAND2_6474 ( R2358_U401 , R2358_U310 , R2358_U53 );
nand NAND2_6475 ( R2358_U402 , R2358_U63 , R2358_U277 );
nand NAND2_6476 ( R2358_U403 , R2358_U77 , R2358_U242 );
nand NAND2_6477 ( R2358_U404 , U2644 , R2358_U242 );
nand NAND2_6478 ( R2358_U405 , U2640 , R2358_U518 );
nand NAND2_6479 ( R2358_U406 , R2358_U8 , R2358_U62 );
nand NAND2_6480 ( R2358_U407 , R2358_U297 , R2358_U9 );
nand NAND2_6481 ( R2358_U408 , R2358_U298 , R2358_U9 );
nand NAND2_6482 ( R2358_U409 , R2358_U159 , R2358_U67 );
nand NAND3_6483 ( R2358_U410 , R2358_U223 , R2358_U224 , R2358_U299 );
nand NAND4_6484 ( R2358_U411 , R2358_U309 , R2358_U311 , R2358_U224 , R2358_U299 );
not NOT1_6485 ( R2358_U412 , R2358_U69 );
nand NAND2_6486 ( R2358_U413 , R2358_U10 , R2358_U176 );
nand NAND2_6487 ( R2358_U414 , R2358_U254 , R2358_U304 );
nand NAND2_6488 ( R2358_U415 , R2358_U13 , R2358_U71 );
nand NAND2_6489 ( R2358_U416 , R2358_U426 , R2358_U67 );
nand NAND2_6490 ( R2358_U417 , R2358_U69 , R2358_U317 );
not NOT1_6491 ( R2358_U418 , R2358_U66 );
nand NAND2_6492 ( R2358_U419 , R2358_U13 , R2358_U71 );
nand NAND3_6493 ( R2358_U420 , R2358_U427 , R2358_U419 , R2358_U428 );
nand NAND2_6494 ( R2358_U421 , R2358_U67 , R2358_U148 );
nand NAND2_6495 ( R2358_U422 , R2358_U66 , R2358_U7 );
not NOT1_6496 ( R2358_U423 , R2358_U73 );
nand NAND2_6497 ( R2358_U424 , R2358_U405 , R2358_U302 );
nand NAND2_6498 ( R2358_U425 , R2358_U424 , R2358_U303 );
not NOT1_6499 ( R2358_U426 , R2358_U55 );
nand NAND2_6500 ( R2358_U427 , R2358_U227 , R2358_U71 );
nand NAND2_6501 ( R2358_U428 , R2358_U534 , R2358_U227 );
nand NAND2_6502 ( R2358_U429 , R2358_U143 , R2358_U435 );
nand NAND2_6503 ( R2358_U430 , R2358_U12 , R2358_U66 );
nand NAND2_6504 ( R2358_U431 , R2358_U136 , R2358_U176 );
nand NAND2_6505 ( R2358_U432 , R2358_U11 , R2358_U73 );
nand NAND2_6506 ( R2358_U433 , R2358_U312 , R2358_U418 );
nand NAND2_6507 ( R2358_U434 , R2358_U418 , R2358_U55 );
nand NAND3_6508 ( R2358_U435 , R2358_U410 , R2358_U219 , R2358_U140 );
nand NAND2_6509 ( R2358_U436 , R2358_U133 , R2358_U327 );
nand NAND2_6510 ( R2358_U437 , R2358_U436 , R2358_U324 );
nand NAND2_6511 ( R2358_U438 , R2358_U134 , R2358_U328 );
not NOT1_6512 ( R2358_U439 , R2358_U62 );
nand NAND2_6513 ( R2358_U440 , U2352 , R2358_U164 );
nand NAND2_6514 ( R2358_U441 , U2612 , R2358_U22 );
not NOT1_6515 ( R2358_U442 , R2358_U76 );
nand NAND2_6516 ( R2358_U443 , R2358_U442 , U2641 );
nand NAND2_6517 ( R2358_U444 , R2358_U76 , R2358_U33 );
nand NAND2_6518 ( R2358_U445 , R2358_U442 , U2641 );
nand NAND2_6519 ( R2358_U446 , R2358_U76 , R2358_U33 );
nand NAND2_6520 ( R2358_U447 , R2358_U446 , R2358_U445 );
nand NAND2_6521 ( R2358_U448 , U2352 , R2358_U166 );
nand NAND2_6522 ( R2358_U449 , U2610 , R2358_U22 );
nand NAND2_6523 ( R2358_U450 , R2358_U449 , R2358_U448 );
nand NAND2_6524 ( R2358_U451 , U2352 , R2358_U166 );
nand NAND2_6525 ( R2358_U452 , U2610 , R2358_U22 );
nand NAND2_6526 ( R2358_U453 , U2352 , R2358_U167 );
nand NAND2_6527 ( R2358_U454 , U2609 , R2358_U22 );
not NOT1_6528 ( R2358_U455 , R2358_U77 );
nand NAND2_6529 ( R2358_U456 , U2352 , R2358_U168 );
nand NAND2_6530 ( R2358_U457 , U2667 , R2358_U22 );
nand NAND2_6531 ( R2358_U458 , R2358_U457 , R2358_U456 );
nand NAND2_6532 ( R2358_U459 , U2352 , R2358_U169 );
nand NAND2_6533 ( R2358_U460 , U2668 , R2358_U22 );
nand NAND2_6534 ( R2358_U461 , R2358_U460 , R2358_U459 );
nand NAND2_6535 ( R2358_U462 , U2352 , R2358_U168 );
nand NAND2_6536 ( R2358_U463 , U2667 , R2358_U22 );
nand NAND2_6537 ( R2358_U464 , U2352 , R2358_U169 );
nand NAND2_6538 ( R2358_U465 , U2668 , R2358_U22 );
nand NAND2_6539 ( R2358_U466 , U2352 , R2358_U170 );
nand NAND2_6540 ( R2358_U467 , U2670 , R2358_U22 );
nand NAND2_6541 ( R2358_U468 , R2358_U467 , R2358_U466 );
nand NAND2_6542 ( R2358_U469 , U2352 , R2358_U171 );
nand NAND2_6543 ( R2358_U470 , U2671 , R2358_U22 );
nand NAND2_6544 ( R2358_U471 , R2358_U470 , R2358_U469 );
nand NAND2_6545 ( R2358_U472 , U2352 , R2358_U172 );
nand NAND2_6546 ( R2358_U473 , U2672 , R2358_U22 );
nand NAND2_6547 ( R2358_U474 , R2358_U473 , R2358_U472 );
nand NAND2_6548 ( R2358_U475 , U2352 , R2358_U171 );
nand NAND2_6549 ( R2358_U476 , U2671 , R2358_U22 );
nand NAND2_6550 ( R2358_U477 , U2352 , R2358_U172 );
nand NAND2_6551 ( R2358_U478 , U2672 , R2358_U22 );
nand NAND2_6552 ( R2358_U479 , U2352 , R2358_U170 );
nand NAND2_6553 ( R2358_U480 , U2670 , R2358_U22 );
nand NAND2_6554 ( R2358_U481 , U2352 , R2358_U173 );
nand NAND2_6555 ( R2358_U482 , U2669 , R2358_U22 );
nand NAND2_6556 ( R2358_U483 , U2352 , R2358_U173 );
nand NAND2_6557 ( R2358_U484 , U2669 , R2358_U22 );
nand NAND2_6558 ( R2358_U485 , R2358_U484 , R2358_U483 );
nand NAND2_6559 ( R2358_U486 , U2352 , R2358_U174 );
nand NAND2_6560 ( R2358_U487 , U2611 , R2358_U22 );
nand NAND2_6561 ( R2358_U488 , U2352 , R2358_U174 );
nand NAND2_6562 ( R2358_U489 , U2611 , R2358_U22 );
nand NAND2_6563 ( R2358_U490 , R2358_U489 , R2358_U488 );
nand NAND2_6564 ( R2358_U491 , R2358_U165 , R2358_U175 );
nand NAND2_6565 ( R2358_U492 , R2358_U256 , R2358_U447 );
nand NAND2_6566 ( R2358_U493 , R2358_U381 , R2358_U176 );
nand NAND2_6567 ( R2358_U494 , R2358_U84 , R2358_U252 );
nand NAND2_6568 ( R2358_U495 , R2358_U455 , U2644 );
nand NAND2_6569 ( R2358_U496 , R2358_U77 , R2358_U24 );
nand NAND2_6570 ( R2358_U497 , R2358_U496 , R2358_U495 );
nand NAND2_6571 ( R2358_U498 , R2358_U382 , R2358_U34 );
nand NAND2_6572 ( R2358_U499 , R2358_U497 , R2358_U260 );
nand NAND2_6573 ( R2358_U500 , R2358_U383 , R2358_U177 );
nand NAND2_6574 ( R2358_U501 , R2358_U87 , R2358_U258 );
nand NAND2_6575 ( R2358_U502 , R2358_U384 , R2358_U178 );
nand NAND2_6576 ( R2358_U503 , R2358_U89 , R2358_U241 );
nand NAND2_6577 ( R2358_U504 , U2352 , R2358_U179 );
nand NAND2_6578 ( R2358_U505 , U2651 , R2358_U22 );
nand NAND2_6579 ( R2358_U506 , U2352 , R2358_U179 );
nand NAND2_6580 ( R2358_U507 , U2651 , R2358_U22 );
nand NAND2_6581 ( R2358_U508 , R2358_U507 , R2358_U506 );
nand NAND2_6582 ( R2358_U509 , U2352 , R2358_U181 );
nand NAND2_6583 ( R2358_U510 , U2613 , R2358_U22 );
nand NAND2_6584 ( R2358_U511 , U2352 , R2358_U182 );
nand NAND2_6585 ( R2358_U512 , U2614 , R2358_U22 );
nand NAND2_6586 ( R2358_U513 , U2352 , R2358_U182 );
nand NAND2_6587 ( R2358_U514 , U2614 , R2358_U22 );
nand NAND2_6588 ( R2358_U515 , R2358_U514 , R2358_U513 );
nand NAND2_6589 ( R2358_U516 , U2352 , R2358_U181 );
nand NAND2_6590 ( R2358_U517 , U2613 , R2358_U22 );
nand NAND2_6591 ( R2358_U518 , R2358_U517 , R2358_U516 );
nand NAND2_6592 ( R2358_U519 , U2352 , R2358_U183 );
nand NAND2_6593 ( R2358_U520 , U2617 , R2358_U22 );
not NOT1_6594 ( R2358_U521 , R2358_U79 );
nand NAND2_6595 ( R2358_U522 , U2352 , R2358_U184 );
nand NAND2_6596 ( R2358_U523 , U2615 , R2358_U22 );
nand NAND2_6597 ( R2358_U524 , U2352 , R2358_U185 );
nand NAND2_6598 ( R2358_U525 , U2616 , R2358_U22 );
not NOT1_6599 ( R2358_U526 , R2358_U80 );
nand NAND2_6600 ( R2358_U527 , U2352 , R2358_U186 );
nand NAND2_6601 ( R2358_U528 , U2618 , R2358_U22 );
nand NAND2_6602 ( R2358_U529 , U2352 , R2358_U184 );
nand NAND2_6603 ( R2358_U530 , U2615 , R2358_U22 );
nand NAND2_6604 ( R2358_U531 , R2358_U530 , R2358_U529 );
nand NAND2_6605 ( R2358_U532 , U2352 , R2358_U186 );
nand NAND2_6606 ( R2358_U533 , U2618 , R2358_U22 );
not NOT1_6607 ( R2358_U534 , R2358_U81 );
nand NAND2_6608 ( R2358_U535 , U2352 , R2358_U187 );
nand NAND2_6609 ( R2358_U536 , U2664 , R2358_U22 );
nand NAND2_6610 ( R2358_U537 , U2352 , R2358_U188 );
nand NAND2_6611 ( R2358_U538 , U2665 , R2358_U22 );
nand NAND2_6612 ( R2358_U539 , U2352 , R2358_U189 );
nand NAND2_6613 ( R2358_U540 , U2666 , R2358_U22 );
nand NAND2_6614 ( R2358_U541 , U2352 , R2358_U190 );
nand NAND2_6615 ( R2358_U542 , U2663 , R2358_U22 );
nand NAND2_6616 ( R2358_U543 , U2352 , R2358_U191 );
nand NAND2_6617 ( R2358_U544 , U2658 , R2358_U22 );
nand NAND2_6618 ( R2358_U545 , U2352 , R2358_U192 );
nand NAND2_6619 ( R2358_U546 , U2659 , R2358_U22 );
nand NAND2_6620 ( R2358_U547 , U2352 , R2358_U193 );
nand NAND2_6621 ( R2358_U548 , U2660 , R2358_U22 );
nand NAND2_6622 ( R2358_U549 , U2352 , R2358_U194 );
nand NAND2_6623 ( R2358_U550 , U2661 , R2358_U22 );
nand NAND2_6624 ( R2358_U551 , U2352 , R2358_U195 );
nand NAND2_6625 ( R2358_U552 , U2662 , R2358_U22 );
not NOT1_6626 ( R2358_U553 , R2358_U78 );
nand NAND2_6627 ( R2358_U554 , U2352 , R2358_U196 );
nand NAND2_6628 ( R2358_U555 , U2654 , R2358_U22 );
nand NAND2_6629 ( R2358_U556 , U2352 , R2358_U197 );
nand NAND2_6630 ( R2358_U557 , U2655 , R2358_U22 );
nand NAND2_6631 ( R2358_U558 , U2352 , R2358_U198 );
nand NAND2_6632 ( R2358_U559 , U2656 , R2358_U22 );
nand NAND2_6633 ( R2358_U560 , U2352 , R2358_U199 );
nand NAND2_6634 ( R2358_U561 , U2657 , R2358_U22 );
nand NAND2_6635 ( R2358_U562 , U2352 , R2358_U200 );
nand NAND2_6636 ( R2358_U563 , U2652 , R2358_U22 );
nand NAND2_6637 ( R2358_U564 , U2352 , R2358_U201 );
nand NAND2_6638 ( R2358_U565 , U2653 , R2358_U22 );
nand NAND2_6639 ( R2358_U566 , U2352 , R2358_U191 );
nand NAND2_6640 ( R2358_U567 , U2658 , R2358_U22 );
nand NAND2_6641 ( R2358_U568 , R2358_U567 , R2358_U566 );
nand NAND2_6642 ( R2358_U569 , U2352 , R2358_U192 );
nand NAND2_6643 ( R2358_U570 , U2659 , R2358_U22 );
nand NAND2_6644 ( R2358_U571 , R2358_U570 , R2358_U569 );
nand NAND2_6645 ( R2358_U572 , U2352 , R2358_U193 );
nand NAND2_6646 ( R2358_U573 , U2660 , R2358_U22 );
nand NAND2_6647 ( R2358_U574 , R2358_U573 , R2358_U572 );
nand NAND2_6648 ( R2358_U575 , U2352 , R2358_U194 );
nand NAND2_6649 ( R2358_U576 , U2661 , R2358_U22 );
nand NAND2_6650 ( R2358_U577 , R2358_U576 , R2358_U575 );
nand NAND2_6651 ( R2358_U578 , U2352 , R2358_U200 );
nand NAND2_6652 ( R2358_U579 , U2652 , R2358_U22 );
nand NAND2_6653 ( R2358_U580 , R2358_U579 , R2358_U578 );
nand NAND2_6654 ( R2358_U581 , U2352 , R2358_U199 );
nand NAND2_6655 ( R2358_U582 , U2657 , R2358_U22 );
nand NAND2_6656 ( R2358_U583 , R2358_U582 , R2358_U581 );
nand NAND2_6657 ( R2358_U584 , U2352 , R2358_U198 );
nand NAND2_6658 ( R2358_U585 , U2656 , R2358_U22 );
nand NAND2_6659 ( R2358_U586 , R2358_U585 , R2358_U584 );
nand NAND2_6660 ( R2358_U587 , U2352 , R2358_U197 );
nand NAND2_6661 ( R2358_U588 , U2655 , R2358_U22 );
nand NAND2_6662 ( R2358_U589 , R2358_U588 , R2358_U587 );
nand NAND2_6663 ( R2358_U590 , U2352 , R2358_U196 );
nand NAND2_6664 ( R2358_U591 , U2654 , R2358_U22 );
nand NAND2_6665 ( R2358_U592 , R2358_U591 , R2358_U590 );
nand NAND2_6666 ( R2358_U593 , U2352 , R2358_U201 );
nand NAND2_6667 ( R2358_U594 , U2653 , R2358_U22 );
nand NAND2_6668 ( R2358_U595 , R2358_U594 , R2358_U593 );
nand NAND2_6669 ( R2358_U596 , U2352 , R2358_U190 );
nand NAND2_6670 ( R2358_U597 , U2663 , R2358_U22 );
nand NAND2_6671 ( R2358_U598 , R2358_U597 , R2358_U596 );
nand NAND2_6672 ( R2358_U599 , U2352 , R2358_U189 );
nand NAND2_6673 ( R2358_U600 , U2666 , R2358_U22 );
nand NAND2_6674 ( R2358_U601 , R2358_U600 , R2358_U599 );
nand NAND2_6675 ( R2358_U602 , U2352 , R2358_U187 );
nand NAND2_6676 ( R2358_U603 , U2664 , R2358_U22 );
nand NAND2_6677 ( R2358_U604 , R2358_U603 , R2358_U602 );
nand NAND2_6678 ( R2358_U605 , U2352 , R2358_U188 );
nand NAND2_6679 ( R2358_U606 , U2665 , R2358_U22 );
nand NAND2_6680 ( R2358_U607 , R2358_U606 , R2358_U605 );
nand NAND2_6681 ( R2358_U608 , R2358_U180 , R2358_U202 );
nand NAND2_6682 ( R2358_U609 , R2358_U330 , R2358_U508 );
nand NAND2_6683 ( R2358_U610 , R2358_U385 , R2358_U203 );
nand NAND2_6684 ( R2358_U611 , R2358_U92 , R2358_U333 );
nand NAND2_6685 ( R2358_U612 , R2358_U386 , R2358_U204 );
nand NAND2_6686 ( R2358_U613 , R2358_U94 , R2358_U339 );
nand NAND2_6687 ( R2358_U614 , R2358_U387 , R2358_U205 );
nand NAND2_6688 ( R2358_U615 , R2358_U96 , R2358_U341 );
nand NAND2_6689 ( R2358_U616 , R2358_U221 , R2358_U388 );
nand NAND2_6690 ( R2358_U617 , R2358_U98 , R2358_U206 );
nand NAND2_6691 ( R2358_U618 , R2358_U389 , R2358_U207 );
nand NAND2_6692 ( R2358_U619 , R2358_U100 , R2358_U343 );
nand NAND2_6693 ( R2358_U620 , R2358_U390 , R2358_U208 );
nand NAND2_6694 ( R2358_U621 , R2358_U102 , R2358_U331 );
nand NAND2_6695 ( R2358_U622 , R2358_U391 , R2358_U209 );
nand NAND2_6696 ( R2358_U623 , R2358_U104 , R2358_U348 );
nand NAND2_6697 ( R2358_U624 , R2358_U392 , R2358_U210 );
nand NAND2_6698 ( R2358_U625 , R2358_U106 , R2358_U346 );
nand NAND2_6699 ( R2358_U626 , R2358_U220 , R2358_U393 );
nand NAND2_6700 ( R2358_U627 , R2358_U108 , R2358_U211 );
nand NAND2_6701 ( R2358_U628 , R2358_U553 , U2630 );
nand NAND2_6702 ( R2358_U629 , R2358_U78 , R2358_U45 );
nand NAND2_6703 ( R2358_U630 , R2358_U629 , R2358_U628 );
nand NAND2_6704 ( R2358_U631 , R2358_U394 , R2358_U68 );
nand NAND2_6705 ( R2358_U632 , R2358_U630 , R2358_U318 );
nand NAND2_6706 ( R2358_U633 , R2358_U395 , R2358_U212 );
nand NAND2_6707 ( R2358_U634 , R2358_U111 , R2358_U269 );
nand NAND2_6708 ( R2358_U635 , R2358_U396 , R2358_U213 );
nand NAND2_6709 ( R2358_U636 , R2358_U113 , R2358_U315 );
nand NAND2_6710 ( R2358_U637 , R2358_U397 , R2358_U214 );
nand NAND2_6711 ( R2358_U638 , R2358_U115 , R2358_U357 );
nand NAND2_6712 ( R2358_U639 , R2358_U398 , R2358_U215 );
nand NAND2_6713 ( R2358_U640 , R2358_U117 , R2358_U355 );
nand NAND2_6714 ( R2358_U641 , R2358_U521 , U2636 );
nand NAND2_6715 ( R2358_U642 , R2358_U79 , R2358_U54 );
nand NAND2_6716 ( R2358_U643 , R2358_U642 , R2358_U641 );
nand NAND2_6717 ( R2358_U644 , R2358_U399 , R2358_U72 );
nand NAND2_6718 ( R2358_U645 , R2358_U643 , R2358_U365 );
nand NAND2_6719 ( R2358_U646 , R2358_U526 , U2637 );
nand NAND2_6720 ( R2358_U647 , R2358_U80 , R2358_U50 );
nand NAND2_6721 ( R2358_U648 , R2358_U647 , R2358_U646 );
nand NAND2_6722 ( R2358_U649 , R2358_U400 , R2358_U216 );
nand NAND2_6723 ( R2358_U650 , R2358_U362 , R2358_U648 );
nand NAND2_6724 ( R2358_U651 , R2358_U401 , R2358_U217 );
nand NAND2_6725 ( R2358_U652 , R2358_U121 , R2358_U308 );
nand NAND2_6726 ( R2358_U653 , U2352 , R2358_U218 );
nand NAND2_6727 ( R2358_U654 , R2358_U380 , R2358_U22 );
not NOT1_6728 ( R2337_U5 , PHYADDRPOINTER_REG_1_ );
not NOT1_6729 ( R2337_U6 , PHYADDRPOINTER_REG_5_ );
not NOT1_6730 ( R2337_U7 , PHYADDRPOINTER_REG_4_ );
not NOT1_6731 ( R2337_U8 , PHYADDRPOINTER_REG_3_ );
not NOT1_6732 ( R2337_U9 , PHYADDRPOINTER_REG_2_ );
nand NAND5_6733 ( R2337_U10 , PHYADDRPOINTER_REG_5_ , PHYADDRPOINTER_REG_1_ , PHYADDRPOINTER_REG_4_ , PHYADDRPOINTER_REG_2_ , PHYADDRPOINTER_REG_3_ );
not NOT1_6734 ( R2337_U11 , PHYADDRPOINTER_REG_7_ );
not NOT1_6735 ( R2337_U12 , PHYADDRPOINTER_REG_6_ );
nand NAND2_6736 ( R2337_U13 , R2337_U81 , R2337_U108 );
not NOT1_6737 ( R2337_U14 , PHYADDRPOINTER_REG_8_ );
not NOT1_6738 ( R2337_U15 , PHYADDRPOINTER_REG_9_ );
nand NAND3_6739 ( R2337_U16 , PHYADDRPOINTER_REG_3_ , PHYADDRPOINTER_REG_1_ , PHYADDRPOINTER_REG_2_ );
nand NAND2_6740 ( R2337_U17 , R2337_U82 , R2337_U110 );
not NOT1_6741 ( R2337_U18 , PHYADDRPOINTER_REG_11_ );
not NOT1_6742 ( R2337_U19 , PHYADDRPOINTER_REG_10_ );
nand NAND2_6743 ( R2337_U20 , R2337_U83 , R2337_U112 );
not NOT1_6744 ( R2337_U21 , PHYADDRPOINTER_REG_13_ );
not NOT1_6745 ( R2337_U22 , PHYADDRPOINTER_REG_12_ );
nand NAND2_6746 ( R2337_U23 , R2337_U84 , R2337_U114 );
not NOT1_6747 ( R2337_U24 , PHYADDRPOINTER_REG_15_ );
not NOT1_6748 ( R2337_U25 , PHYADDRPOINTER_REG_14_ );
nand NAND2_6749 ( R2337_U26 , R2337_U85 , R2337_U116 );
not NOT1_6750 ( R2337_U27 , PHYADDRPOINTER_REG_17_ );
not NOT1_6751 ( R2337_U28 , PHYADDRPOINTER_REG_16_ );
nand NAND2_6752 ( R2337_U29 , R2337_U86 , R2337_U118 );
not NOT1_6753 ( R2337_U30 , PHYADDRPOINTER_REG_19_ );
not NOT1_6754 ( R2337_U31 , PHYADDRPOINTER_REG_18_ );
nand NAND2_6755 ( R2337_U32 , R2337_U87 , R2337_U120 );
not NOT1_6756 ( R2337_U33 , PHYADDRPOINTER_REG_21_ );
not NOT1_6757 ( R2337_U34 , PHYADDRPOINTER_REG_20_ );
nand NAND2_6758 ( R2337_U35 , R2337_U88 , R2337_U122 );
not NOT1_6759 ( R2337_U36 , PHYADDRPOINTER_REG_23_ );
not NOT1_6760 ( R2337_U37 , PHYADDRPOINTER_REG_22_ );
nand NAND2_6761 ( R2337_U38 , R2337_U89 , R2337_U124 );
not NOT1_6762 ( R2337_U39 , PHYADDRPOINTER_REG_25_ );
not NOT1_6763 ( R2337_U40 , PHYADDRPOINTER_REG_24_ );
nand NAND2_6764 ( R2337_U41 , R2337_U90 , R2337_U126 );
not NOT1_6765 ( R2337_U42 , PHYADDRPOINTER_REG_26_ );
nand NAND2_6766 ( R2337_U43 , PHYADDRPOINTER_REG_26_ , R2337_U128 );
not NOT1_6767 ( R2337_U44 , PHYADDRPOINTER_REG_27_ );
nand NAND2_6768 ( R2337_U45 , PHYADDRPOINTER_REG_27_ , R2337_U129 );
not NOT1_6769 ( R2337_U46 , PHYADDRPOINTER_REG_28_ );
nand NAND2_6770 ( R2337_U47 , PHYADDRPOINTER_REG_28_ , R2337_U130 );
not NOT1_6771 ( R2337_U48 , PHYADDRPOINTER_REG_29_ );
nand NAND2_6772 ( R2337_U49 , PHYADDRPOINTER_REG_29_ , R2337_U131 );
not NOT1_6773 ( R2337_U50 , PHYADDRPOINTER_REG_30_ );
nand NAND2_6774 ( R2337_U51 , R2337_U135 , R2337_U134 );
nand NAND2_6775 ( R2337_U52 , R2337_U137 , R2337_U136 );
nand NAND2_6776 ( R2337_U53 , R2337_U139 , R2337_U138 );
nand NAND2_6777 ( R2337_U54 , R2337_U141 , R2337_U140 );
nand NAND2_6778 ( R2337_U55 , R2337_U143 , R2337_U142 );
nand NAND2_6779 ( R2337_U56 , R2337_U145 , R2337_U144 );
nand NAND2_6780 ( R2337_U57 , R2337_U147 , R2337_U146 );
nand NAND2_6781 ( R2337_U58 , R2337_U149 , R2337_U148 );
nand NAND2_6782 ( R2337_U59 , R2337_U151 , R2337_U150 );
nand NAND2_6783 ( R2337_U60 , R2337_U153 , R2337_U152 );
nand NAND2_6784 ( R2337_U61 , R2337_U155 , R2337_U154 );
nand NAND2_6785 ( R2337_U62 , R2337_U157 , R2337_U156 );
nand NAND2_6786 ( R2337_U63 , R2337_U159 , R2337_U158 );
nand NAND2_6787 ( R2337_U64 , R2337_U161 , R2337_U160 );
nand NAND2_6788 ( R2337_U65 , R2337_U163 , R2337_U162 );
nand NAND2_6789 ( R2337_U66 , R2337_U165 , R2337_U164 );
nand NAND2_6790 ( R2337_U67 , R2337_U167 , R2337_U166 );
nand NAND2_6791 ( R2337_U68 , R2337_U169 , R2337_U168 );
nand NAND2_6792 ( R2337_U69 , R2337_U171 , R2337_U170 );
nand NAND2_6793 ( R2337_U70 , R2337_U173 , R2337_U172 );
nand NAND2_6794 ( R2337_U71 , R2337_U175 , R2337_U174 );
nand NAND2_6795 ( R2337_U72 , R2337_U177 , R2337_U176 );
nand NAND2_6796 ( R2337_U73 , R2337_U179 , R2337_U178 );
nand NAND2_6797 ( R2337_U74 , R2337_U181 , R2337_U180 );
nand NAND2_6798 ( R2337_U75 , R2337_U183 , R2337_U182 );
nand NAND2_6799 ( R2337_U76 , R2337_U185 , R2337_U184 );
nand NAND2_6800 ( R2337_U77 , R2337_U187 , R2337_U186 );
nand NAND2_6801 ( R2337_U78 , R2337_U189 , R2337_U188 );
nand NAND2_6802 ( R2337_U79 , R2337_U191 , R2337_U190 );
nand NAND2_6803 ( R2337_U80 , R2337_U193 , R2337_U192 );
and AND2_6804 ( R2337_U81 , PHYADDRPOINTER_REG_7_ , PHYADDRPOINTER_REG_6_ );
and AND2_6805 ( R2337_U82 , PHYADDRPOINTER_REG_8_ , PHYADDRPOINTER_REG_9_ );
and AND2_6806 ( R2337_U83 , PHYADDRPOINTER_REG_11_ , PHYADDRPOINTER_REG_10_ );
and AND2_6807 ( R2337_U84 , PHYADDRPOINTER_REG_13_ , PHYADDRPOINTER_REG_12_ );
and AND2_6808 ( R2337_U85 , PHYADDRPOINTER_REG_15_ , PHYADDRPOINTER_REG_14_ );
and AND2_6809 ( R2337_U86 , PHYADDRPOINTER_REG_17_ , PHYADDRPOINTER_REG_16_ );
and AND2_6810 ( R2337_U87 , PHYADDRPOINTER_REG_19_ , PHYADDRPOINTER_REG_18_ );
and AND2_6811 ( R2337_U88 , PHYADDRPOINTER_REG_21_ , PHYADDRPOINTER_REG_20_ );
and AND2_6812 ( R2337_U89 , PHYADDRPOINTER_REG_23_ , PHYADDRPOINTER_REG_22_ );
and AND2_6813 ( R2337_U90 , PHYADDRPOINTER_REG_25_ , PHYADDRPOINTER_REG_24_ );
nand NAND2_6814 ( R2337_U91 , PHYADDRPOINTER_REG_8_ , R2337_U110 );
nand NAND2_6815 ( R2337_U92 , PHYADDRPOINTER_REG_6_ , R2337_U108 );
nand NAND2_6816 ( R2337_U93 , R2337_U106 , PHYADDRPOINTER_REG_4_ );
nand NAND2_6817 ( R2337_U94 , PHYADDRPOINTER_REG_2_ , PHYADDRPOINTER_REG_1_ );
not NOT1_6818 ( R2337_U95 , PHYADDRPOINTER_REG_31_ );
nand NAND2_6819 ( R2337_U96 , PHYADDRPOINTER_REG_30_ , R2337_U132 );
nand NAND2_6820 ( R2337_U97 , PHYADDRPOINTER_REG_24_ , R2337_U126 );
nand NAND2_6821 ( R2337_U98 , PHYADDRPOINTER_REG_22_ , R2337_U124 );
nand NAND2_6822 ( R2337_U99 , PHYADDRPOINTER_REG_20_ , R2337_U122 );
nand NAND2_6823 ( R2337_U100 , PHYADDRPOINTER_REG_18_ , R2337_U120 );
nand NAND2_6824 ( R2337_U101 , PHYADDRPOINTER_REG_16_ , R2337_U118 );
nand NAND2_6825 ( R2337_U102 , PHYADDRPOINTER_REG_14_ , R2337_U116 );
nand NAND2_6826 ( R2337_U103 , PHYADDRPOINTER_REG_12_ , R2337_U114 );
nand NAND2_6827 ( R2337_U104 , PHYADDRPOINTER_REG_10_ , R2337_U112 );
not NOT1_6828 ( R2337_U105 , R2337_U94 );
not NOT1_6829 ( R2337_U106 , R2337_U16 );
not NOT1_6830 ( R2337_U107 , R2337_U93 );
not NOT1_6831 ( R2337_U108 , R2337_U10 );
not NOT1_6832 ( R2337_U109 , R2337_U92 );
not NOT1_6833 ( R2337_U110 , R2337_U13 );
not NOT1_6834 ( R2337_U111 , R2337_U91 );
not NOT1_6835 ( R2337_U112 , R2337_U17 );
not NOT1_6836 ( R2337_U113 , R2337_U104 );
not NOT1_6837 ( R2337_U114 , R2337_U20 );
not NOT1_6838 ( R2337_U115 , R2337_U103 );
not NOT1_6839 ( R2337_U116 , R2337_U23 );
not NOT1_6840 ( R2337_U117 , R2337_U102 );
not NOT1_6841 ( R2337_U118 , R2337_U26 );
not NOT1_6842 ( R2337_U119 , R2337_U101 );
not NOT1_6843 ( R2337_U120 , R2337_U29 );
not NOT1_6844 ( R2337_U121 , R2337_U100 );
not NOT1_6845 ( R2337_U122 , R2337_U32 );
not NOT1_6846 ( R2337_U123 , R2337_U99 );
not NOT1_6847 ( R2337_U124 , R2337_U35 );
not NOT1_6848 ( R2337_U125 , R2337_U98 );
not NOT1_6849 ( R2337_U126 , R2337_U38 );
not NOT1_6850 ( R2337_U127 , R2337_U97 );
not NOT1_6851 ( R2337_U128 , R2337_U41 );
not NOT1_6852 ( R2337_U129 , R2337_U43 );
not NOT1_6853 ( R2337_U130 , R2337_U45 );
not NOT1_6854 ( R2337_U131 , R2337_U47 );
not NOT1_6855 ( R2337_U132 , R2337_U49 );
not NOT1_6856 ( R2337_U133 , R2337_U96 );
nand NAND2_6857 ( R2337_U134 , PHYADDRPOINTER_REG_9_ , R2337_U91 );
nand NAND2_6858 ( R2337_U135 , R2337_U111 , R2337_U15 );
nand NAND2_6859 ( R2337_U136 , PHYADDRPOINTER_REG_8_ , R2337_U13 );
nand NAND2_6860 ( R2337_U137 , R2337_U110 , R2337_U14 );
nand NAND2_6861 ( R2337_U138 , PHYADDRPOINTER_REG_7_ , R2337_U92 );
nand NAND2_6862 ( R2337_U139 , R2337_U109 , R2337_U11 );
nand NAND2_6863 ( R2337_U140 , PHYADDRPOINTER_REG_6_ , R2337_U10 );
nand NAND2_6864 ( R2337_U141 , R2337_U108 , R2337_U12 );
nand NAND2_6865 ( R2337_U142 , PHYADDRPOINTER_REG_5_ , R2337_U93 );
nand NAND2_6866 ( R2337_U143 , R2337_U107 , R2337_U6 );
nand NAND2_6867 ( R2337_U144 , PHYADDRPOINTER_REG_4_ , R2337_U16 );
nand NAND2_6868 ( R2337_U145 , R2337_U106 , R2337_U7 );
nand NAND2_6869 ( R2337_U146 , PHYADDRPOINTER_REG_3_ , R2337_U94 );
nand NAND2_6870 ( R2337_U147 , R2337_U105 , R2337_U8 );
nand NAND2_6871 ( R2337_U148 , PHYADDRPOINTER_REG_31_ , R2337_U96 );
nand NAND2_6872 ( R2337_U149 , R2337_U133 , R2337_U95 );
nand NAND2_6873 ( R2337_U150 , PHYADDRPOINTER_REG_30_ , R2337_U49 );
nand NAND2_6874 ( R2337_U151 , R2337_U132 , R2337_U50 );
nand NAND2_6875 ( R2337_U152 , PHYADDRPOINTER_REG_1_ , R2337_U9 );
nand NAND2_6876 ( R2337_U153 , PHYADDRPOINTER_REG_2_ , R2337_U5 );
nand NAND2_6877 ( R2337_U154 , PHYADDRPOINTER_REG_29_ , R2337_U47 );
nand NAND2_6878 ( R2337_U155 , R2337_U131 , R2337_U48 );
nand NAND2_6879 ( R2337_U156 , PHYADDRPOINTER_REG_28_ , R2337_U45 );
nand NAND2_6880 ( R2337_U157 , R2337_U130 , R2337_U46 );
nand NAND2_6881 ( R2337_U158 , PHYADDRPOINTER_REG_27_ , R2337_U43 );
nand NAND2_6882 ( R2337_U159 , R2337_U129 , R2337_U44 );
nand NAND2_6883 ( R2337_U160 , PHYADDRPOINTER_REG_26_ , R2337_U41 );
nand NAND2_6884 ( R2337_U161 , R2337_U128 , R2337_U42 );
nand NAND2_6885 ( R2337_U162 , PHYADDRPOINTER_REG_25_ , R2337_U97 );
nand NAND2_6886 ( R2337_U163 , R2337_U127 , R2337_U39 );
nand NAND2_6887 ( R2337_U164 , PHYADDRPOINTER_REG_24_ , R2337_U38 );
nand NAND2_6888 ( R2337_U165 , R2337_U126 , R2337_U40 );
nand NAND2_6889 ( R2337_U166 , PHYADDRPOINTER_REG_23_ , R2337_U98 );
nand NAND2_6890 ( R2337_U167 , R2337_U125 , R2337_U36 );
nand NAND2_6891 ( R2337_U168 , PHYADDRPOINTER_REG_22_ , R2337_U35 );
nand NAND2_6892 ( R2337_U169 , R2337_U124 , R2337_U37 );
nand NAND2_6893 ( R2337_U170 , PHYADDRPOINTER_REG_21_ , R2337_U99 );
nand NAND2_6894 ( R2337_U171 , R2337_U123 , R2337_U33 );
nand NAND2_6895 ( R2337_U172 , PHYADDRPOINTER_REG_20_ , R2337_U32 );
nand NAND2_6896 ( R2337_U173 , R2337_U122 , R2337_U34 );
nand NAND2_6897 ( R2337_U174 , PHYADDRPOINTER_REG_19_ , R2337_U100 );
nand NAND2_6898 ( R2337_U175 , R2337_U121 , R2337_U30 );
nand NAND2_6899 ( R2337_U176 , PHYADDRPOINTER_REG_18_ , R2337_U29 );
nand NAND2_6900 ( R2337_U177 , R2337_U120 , R2337_U31 );
nand NAND2_6901 ( R2337_U178 , PHYADDRPOINTER_REG_17_ , R2337_U101 );
nand NAND2_6902 ( R2337_U179 , R2337_U119 , R2337_U27 );
nand NAND2_6903 ( R2337_U180 , PHYADDRPOINTER_REG_16_ , R2337_U26 );
nand NAND2_6904 ( R2337_U181 , R2337_U118 , R2337_U28 );
nand NAND2_6905 ( R2337_U182 , PHYADDRPOINTER_REG_15_ , R2337_U102 );
nand NAND2_6906 ( R2337_U183 , R2337_U117 , R2337_U24 );
nand NAND2_6907 ( R2337_U184 , PHYADDRPOINTER_REG_14_ , R2337_U23 );
nand NAND2_6908 ( R2337_U185 , R2337_U116 , R2337_U25 );
nand NAND2_6909 ( R2337_U186 , PHYADDRPOINTER_REG_13_ , R2337_U103 );
nand NAND2_6910 ( R2337_U187 , R2337_U115 , R2337_U21 );
nand NAND2_6911 ( R2337_U188 , PHYADDRPOINTER_REG_12_ , R2337_U20 );
nand NAND2_6912 ( R2337_U189 , R2337_U114 , R2337_U22 );
nand NAND2_6913 ( R2337_U190 , PHYADDRPOINTER_REG_11_ , R2337_U104 );
nand NAND2_6914 ( R2337_U191 , R2337_U113 , R2337_U18 );
nand NAND2_6915 ( R2337_U192 , PHYADDRPOINTER_REG_10_ , R2337_U17 );
nand NAND2_6916 ( R2337_U193 , R2337_U112 , R2337_U19 );
and AND2_6917 ( R2182_U5 , R2182_U47 , U2740 );
and AND2_6918 ( R2182_U6 , R2182_U60 , R2182_U16 );
not NOT1_6919 ( R2182_U7 , U2744 );
not NOT1_6920 ( R2182_U8 , U3233 );
nand NAND2_6921 ( R2182_U9 , U3233 , U2744 );
not NOT1_6922 ( R2182_U10 , U2742 );
not NOT1_6923 ( R2182_U11 , U2741 );
not NOT1_6924 ( R2182_U12 , U2740 );
nand NAND2_6925 ( R2182_U13 , R2182_U35 , R2182_U41 );
not NOT1_6926 ( R2182_U14 , U2737 );
not NOT1_6927 ( R2182_U15 , U2738 );
nand NAND2_6928 ( R2182_U16 , U2723 , U2739 );
not NOT1_6929 ( R2182_U17 , U2736 );
not NOT1_6930 ( R2182_U18 , U2735 );
nand NAND2_6931 ( R2182_U19 , R2182_U36 , R2182_U49 );
not NOT1_6932 ( R2182_U20 , U2734 );
nand NAND2_6933 ( R2182_U21 , R2182_U37 , R2182_U46 );
nand NAND2_6934 ( R2182_U22 , R2182_U48 , U2734 );
not NOT1_6935 ( R2182_U23 , U2733 );
nand NAND2_6936 ( R2182_U24 , R2182_U64 , R2182_U63 );
nand NAND2_6937 ( R2182_U25 , R2182_U66 , R2182_U65 );
nand NAND2_6938 ( R2182_U26 , R2182_U68 , R2182_U67 );
nand NAND2_6939 ( R2182_U27 , R2182_U72 , R2182_U71 );
nand NAND2_6940 ( R2182_U28 , R2182_U74 , R2182_U73 );
nand NAND2_6941 ( R2182_U29 , R2182_U76 , R2182_U75 );
nand NAND2_6942 ( R2182_U30 , R2182_U78 , R2182_U77 );
nand NAND2_6943 ( R2182_U31 , R2182_U80 , R2182_U79 );
nand NAND2_6944 ( R2182_U32 , R2182_U82 , R2182_U81 );
nand NAND2_6945 ( R2182_U33 , R2182_U84 , R2182_U83 );
nand NAND2_6946 ( R2182_U34 , R2182_U86 , R2182_U85 );
and AND2_6947 ( R2182_U35 , U2742 , U2741 );
and AND2_6948 ( R2182_U36 , U2738 , U2737 );
and AND2_6949 ( R2182_U37 , U2735 , U2736 );
nand NAND2_6950 ( R2182_U38 , U2742 , R2182_U41 );
not NOT1_6951 ( R2182_U39 , U2732 );
nand NAND2_6952 ( R2182_U40 , U2733 , R2182_U56 );
nand NAND2_6953 ( R2182_U41 , R2182_U52 , R2182_U53 );
and AND2_6954 ( R2182_U42 , R2182_U70 , R2182_U69 );
nand NAND2_6955 ( R2182_U43 , R2182_U46 , U2736 );
nand NAND2_6956 ( R2182_U44 , R2182_U49 , U2738 );
nand NAND2_6957 ( R2182_U45 , R2182_U51 , R2182_U62 );
not NOT1_6958 ( R2182_U46 , R2182_U19 );
not NOT1_6959 ( R2182_U47 , R2182_U13 );
not NOT1_6960 ( R2182_U48 , R2182_U21 );
not NOT1_6961 ( R2182_U49 , R2182_U16 );
not NOT1_6962 ( R2182_U50 , R2182_U9 );
or OR2_6963 ( R2182_U51 , U2743 , U2731 );
nand NAND2_6964 ( R2182_U52 , U2731 , U2743 );
nand NAND2_6965 ( R2182_U53 , R2182_U50 , R2182_U51 );
not NOT1_6966 ( R2182_U54 , R2182_U41 );
not NOT1_6967 ( R2182_U55 , R2182_U38 );
not NOT1_6968 ( R2182_U56 , R2182_U22 );
not NOT1_6969 ( R2182_U57 , R2182_U40 );
not NOT1_6970 ( R2182_U58 , R2182_U43 );
not NOT1_6971 ( R2182_U59 , R2182_U44 );
or OR2_6972 ( R2182_U60 , U2739 , U2723 );
not NOT1_6973 ( R2182_U61 , R2182_U45 );
nand NAND2_6974 ( R2182_U62 , U2731 , U2743 );
nand NAND2_6975 ( R2182_U63 , R2182_U47 , R2182_U12 );
nand NAND2_6976 ( R2182_U64 , U2740 , R2182_U13 );
nand NAND2_6977 ( R2182_U65 , U2741 , R2182_U38 );
nand NAND2_6978 ( R2182_U66 , R2182_U55 , R2182_U11 );
nand NAND2_6979 ( R2182_U67 , U2732 , R2182_U40 );
nand NAND2_6980 ( R2182_U68 , R2182_U57 , R2182_U39 );
nand NAND2_6981 ( R2182_U69 , U2742 , R2182_U41 );
nand NAND2_6982 ( R2182_U70 , R2182_U54 , R2182_U10 );
nand NAND2_6983 ( R2182_U71 , U2733 , R2182_U22 );
nand NAND2_6984 ( R2182_U72 , R2182_U56 , R2182_U23 );
nand NAND2_6985 ( R2182_U73 , R2182_U48 , R2182_U20 );
nand NAND2_6986 ( R2182_U74 , U2734 , R2182_U21 );
nand NAND2_6987 ( R2182_U75 , U2735 , R2182_U43 );
nand NAND2_6988 ( R2182_U76 , R2182_U58 , R2182_U18 );
nand NAND2_6989 ( R2182_U77 , R2182_U46 , R2182_U17 );
nand NAND2_6990 ( R2182_U78 , U2736 , R2182_U19 );
nand NAND2_6991 ( R2182_U79 , U2737 , R2182_U44 );
nand NAND2_6992 ( R2182_U80 , R2182_U59 , R2182_U14 );
nand NAND2_6993 ( R2182_U81 , R2182_U49 , R2182_U15 );
nand NAND2_6994 ( R2182_U82 , U2738 , R2182_U16 );
nand NAND2_6995 ( R2182_U83 , R2182_U50 , R2182_U45 );
nand NAND2_6996 ( R2182_U84 , R2182_U61 , R2182_U9 );
nand NAND2_6997 ( R2182_U85 , U3233 , R2182_U7 );
nand NAND2_6998 ( R2182_U86 , U2744 , R2182_U8 );
and AND2_6999 ( R2144_U5 , R2144_U104 , R2144_U103 );
and AND4_7000 ( R2144_U6 , R2144_U36 , R2144_U35 , R2144_U27 , R2144_U29 );
and AND2_7001 ( R2144_U7 , R2144_U104 , R2144_U81 );
and AND2_7002 ( R2144_U8 , R2144_U138 , R2144_U136 );
and AND2_7003 ( R2144_U9 , R2144_U128 , R2144_U127 );
and AND3_7004 ( R2144_U10 , R2144_U213 , R2144_U212 , R2144_U82 );
nand NAND2_7005 ( R2144_U11 , R2144_U144 , R2144_U146 );
not NOT1_7006 ( R2144_U12 , U2355 );
not NOT1_7007 ( R2144_U13 , U2750 );
not NOT1_7008 ( R2144_U14 , U2751 );
not NOT1_7009 ( R2144_U15 , U2752 );
not NOT1_7010 ( R2144_U16 , U2749 );
not NOT1_7011 ( R2144_U17 , U2745 );
not NOT1_7012 ( R2144_U18 , U2748 );
nand NAND2_7013 ( R2144_U19 , U2748 , R2144_U178 );
not NOT1_7014 ( R2144_U20 , U2747 );
nand NAND2_7015 ( R2144_U21 , U2747 , R2144_U170 );
not NOT1_7016 ( R2144_U22 , U2746 );
nand NAND2_7017 ( R2144_U23 , U2746 , R2144_U173 );
nand NAND2_7018 ( R2144_U24 , R2144_U79 , R2144_U63 );
nand NAND2_7019 ( R2144_U25 , R2144_U6 , R2144_U79 );
nand NAND2_7020 ( R2144_U26 , R2144_U65 , R2144_U141 );
nand NAND2_7021 ( R2144_U27 , R2144_U206 , R2144_U205 );
nand NAND2_7022 ( R2144_U28 , R2144_U186 , R2144_U185 );
nand NAND2_7023 ( R2144_U29 , R2144_U203 , R2144_U202 );
nand NAND2_7024 ( R2144_U30 , R2144_U209 , R2144_U208 );
nand NAND2_7025 ( R2144_U31 , R2144_U224 , R2144_U223 );
nand NAND2_7026 ( R2144_U32 , R2144_U221 , R2144_U220 );
nand NAND2_7027 ( R2144_U33 , R2144_U227 , R2144_U226 );
nand NAND2_7028 ( R2144_U34 , R2144_U230 , R2144_U229 );
nand NAND2_7029 ( R2144_U35 , R2144_U233 , R2144_U232 );
nand NAND2_7030 ( R2144_U36 , R2144_U236 , R2144_U235 );
nand NAND2_7031 ( R2144_U37 , R2144_U248 , R2144_U247 );
nand NAND2_7032 ( R2144_U38 , R2144_U250 , R2144_U249 );
nand NAND2_7033 ( R2144_U39 , R2144_U252 , R2144_U251 );
nand NAND2_7034 ( R2144_U40 , R2144_U254 , R2144_U253 );
nand NAND2_7035 ( R2144_U41 , R2144_U256 , R2144_U255 );
nand NAND2_7036 ( R2144_U42 , R2144_U258 , R2144_U257 );
nand NAND2_7037 ( R2144_U43 , R2144_U260 , R2144_U259 );
and AND2_7038 ( R2144_U44 , R2144_U21 , R2144_U105 );
nand NAND2_7039 ( R2144_U45 , R2144_U217 , R2144_U216 );
and AND2_7040 ( R2144_U46 , R2144_U19 , R2144_U106 );
nand NAND2_7041 ( R2144_U47 , R2144_U219 , R2144_U218 );
and AND2_7042 ( R2144_U48 , R2144_U162 , R2144_U109 );
nand NAND2_7043 ( R2144_U49 , R2144_U239 , R2144_U238 );
nand NAND2_7044 ( R2144_U50 , R2144_U246 , R2144_U245 );
and AND2_7045 ( R2144_U51 , R2144_U110 , R2144_U109 );
and AND2_7046 ( R2144_U52 , R2144_U106 , R2144_U105 );
and AND2_7047 ( R2144_U53 , R2144_U7 , R2144_U52 );
and AND4_7048 ( R2144_U54 , R2144_U103 , R2144_U151 , R2144_U153 , R2144_U152 );
and AND2_7049 ( R2144_U55 , R2144_U109 , R2144_U106 );
and AND2_7050 ( R2144_U56 , R2144_U159 , R2144_U19 );
and AND2_7051 ( R2144_U57 , R2144_U156 , R2144_U21 );
and AND3_7052 ( R2144_U58 , R2144_U19 , R2144_U21 , R2144_U159 );
and AND2_7053 ( R2144_U59 , R2144_U5 , R2144_U105 );
and AND2_7054 ( R2144_U60 , R2144_U126 , R2144_U21 );
and AND2_7055 ( R2144_U61 , R2144_U23 , R2144_U81 );
and AND2_7056 ( R2144_U62 , R2144_U111 , R2144_U110 );
and AND2_7057 ( R2144_U63 , R2144_U6 , R2144_U64 );
and AND4_7058 ( R2144_U64 , R2144_U34 , R2144_U33 , R2144_U31 , R2144_U32 );
and AND2_7059 ( R2144_U65 , R2144_U34 , R2144_U33 );
and AND3_7060 ( R2144_U66 , R2144_U36 , R2144_U27 , R2144_U29 );
and AND2_7061 ( R2144_U67 , R2144_U29 , R2144_U27 );
not NOT1_7062 ( R2144_U68 , U2762 );
not NOT1_7063 ( R2144_U69 , U2761 );
not NOT1_7064 ( R2144_U70 , U2763 );
not NOT1_7065 ( R2144_U71 , U2764 );
not NOT1_7066 ( R2144_U72 , U2766 );
not NOT1_7067 ( R2144_U73 , U2767 );
not NOT1_7068 ( R2144_U74 , U2768 );
not NOT1_7069 ( R2144_U75 , U2765 );
not NOT1_7070 ( R2144_U76 , U2760 );
not NOT1_7071 ( R2144_U77 , U2759 );
nand NAND2_7072 ( R2144_U78 , R2144_U29 , R2144_U79 );
nand NAND2_7073 ( R2144_U79 , R2144_U99 , R2144_U54 );
and AND2_7074 ( R2144_U80 , R2144_U211 , R2144_U210 );
nand NAND3_7075 ( R2144_U81 , R2144_U165 , R2144_U164 , R2144_U22 );
and AND2_7076 ( R2144_U82 , R2144_U215 , R2144_U214 );
nand NAND2_7077 ( R2144_U83 , R2144_U56 , R2144_U158 );
nand NAND2_7078 ( R2144_U84 , R2144_U111 , R2144_U118 );
not NOT1_7079 ( R2144_U85 , U2754 );
not NOT1_7080 ( R2144_U86 , U2753 );
not NOT1_7081 ( R2144_U87 , U2755 );
not NOT1_7082 ( R2144_U88 , U2756 );
not NOT1_7083 ( R2144_U89 , U2757 );
not NOT1_7084 ( R2144_U90 , U2758 );
nand NAND2_7085 ( R2144_U91 , R2144_U100 , R2144_U132 );
and AND2_7086 ( R2144_U92 , R2144_U241 , R2144_U240 );
nand NAND2_7087 ( R2144_U93 , R2144_U129 , R2144_U113 );
nand NAND2_7088 ( R2144_U94 , R2144_U143 , R2144_U32 );
nand NAND2_7089 ( R2144_U95 , R2144_U141 , R2144_U34 );
nand NAND2_7090 ( R2144_U96 , R2144_U79 , R2144_U66 );
nand NAND2_7091 ( R2144_U97 , R2144_U67 , R2144_U79 );
nand NAND2_7092 ( R2144_U98 , R2144_U113 , R2144_U112 );
nand NAND2_7093 ( R2144_U99 , R2144_U53 , R2144_U84 );
nand NAND2_7094 ( R2144_U100 , U2751 , R2144_U28 );
not NOT1_7095 ( R2144_U101 , R2144_U24 );
not NOT1_7096 ( R2144_U102 , R2144_U81 );
nand NAND2_7097 ( R2144_U103 , U2745 , R2144_U181 );
nand NAND3_7098 ( R2144_U104 , R2144_U167 , R2144_U166 , R2144_U17 );
nand NAND3_7099 ( R2144_U105 , R2144_U175 , R2144_U174 , R2144_U20 );
nand NAND3_7100 ( R2144_U106 , R2144_U201 , R2144_U200 , R2144_U18 );
not NOT1_7101 ( R2144_U107 , R2144_U21 );
not NOT1_7102 ( R2144_U108 , R2144_U23 );
nand NAND3_7103 ( R2144_U109 , R2144_U194 , R2144_U193 , R2144_U13 );
nand NAND3_7104 ( R2144_U110 , R2144_U196 , R2144_U195 , R2144_U16 );
nand NAND2_7105 ( R2144_U111 , U2749 , R2144_U199 );
nand NAND3_7106 ( R2144_U112 , R2144_U189 , R2144_U188 , R2144_U15 );
nand NAND2_7107 ( R2144_U113 , U2752 , R2144_U192 );
nand NAND2_7108 ( R2144_U114 , R2144_U187 , R2144_U14 );
nand NAND2_7109 ( R2144_U115 , U2355 , R2144_U112 );
nand NAND2_7110 ( R2144_U116 , U2750 , R2144_U184 );
nand NAND2_7111 ( R2144_U117 , R2144_U155 , R2144_U157 );
nand NAND2_7112 ( R2144_U118 , R2144_U51 , R2144_U117 );
not NOT1_7113 ( R2144_U119 , R2144_U84 );
not NOT1_7114 ( R2144_U120 , R2144_U19 );
not NOT1_7115 ( R2144_U121 , R2144_U79 );
not NOT1_7116 ( R2144_U122 , R2144_U78 );
not NOT1_7117 ( R2144_U123 , R2144_U83 );
nand NAND2_7118 ( R2144_U124 , R2144_U83 , R2144_U105 );
nand NAND2_7119 ( R2144_U125 , R2144_U21 , R2144_U124 );
nand NAND2_7120 ( R2144_U126 , R2144_U23 , R2144_U81 );
nand NAND2_7121 ( R2144_U127 , R2144_U60 , R2144_U124 );
nand NAND2_7122 ( R2144_U128 , R2144_U61 , R2144_U125 );
nand NAND2_7123 ( R2144_U129 , U2355 , R2144_U112 );
not NOT1_7124 ( R2144_U130 , R2144_U93 );
nand NAND2_7125 ( R2144_U131 , R2144_U187 , R2144_U14 );
nand NAND2_7126 ( R2144_U132 , R2144_U131 , R2144_U93 );
not NOT1_7127 ( R2144_U133 , R2144_U91 );
nand NAND2_7128 ( R2144_U134 , R2144_U91 , R2144_U109 );
nand NAND2_7129 ( R2144_U135 , R2144_U134 , R2144_U116 );
nand NAND2_7130 ( R2144_U136 , R2144_U62 , R2144_U135 );
nand NAND2_7131 ( R2144_U137 , R2144_U161 , R2144_U110 );
nand NAND3_7132 ( R2144_U138 , R2144_U134 , R2144_U116 , R2144_U137 );
not NOT1_7133 ( R2144_U139 , R2144_U97 );
not NOT1_7134 ( R2144_U140 , R2144_U96 );
not NOT1_7135 ( R2144_U141 , R2144_U25 );
not NOT1_7136 ( R2144_U142 , R2144_U95 );
not NOT1_7137 ( R2144_U143 , R2144_U26 );
nand NAND2_7138 ( R2144_U144 , U2355 , R2144_U24 );
not NOT1_7139 ( R2144_U145 , R2144_U144 );
nand NAND2_7140 ( R2144_U146 , R2144_U101 , R2144_U12 );
not NOT1_7141 ( R2144_U147 , R2144_U94 );
not NOT1_7142 ( R2144_U148 , R2144_U98 );
nand NAND2_7143 ( R2144_U149 , R2144_U21 , R2144_U105 );
nand NAND2_7144 ( R2144_U150 , R2144_U19 , R2144_U106 );
nand NAND3_7145 ( R2144_U151 , R2144_U120 , R2144_U105 , R2144_U7 );
nand NAND2_7146 ( R2144_U152 , R2144_U107 , R2144_U7 );
nand NAND2_7147 ( R2144_U153 , R2144_U108 , R2144_U7 );
nand NAND3_7148 ( R2144_U154 , R2144_U113 , R2144_U115 , R2144_U100 );
nand NAND2_7149 ( R2144_U155 , R2144_U154 , R2144_U114 );
nand NAND2_7150 ( R2144_U156 , R2144_U104 , R2144_U103 );
nand NAND2_7151 ( R2144_U157 , U2750 , R2144_U184 );
nand NAND3_7152 ( R2144_U158 , R2144_U117 , R2144_U110 , R2144_U55 );
nand NAND3_7153 ( R2144_U159 , U2749 , R2144_U106 , R2144_U199 );
nand NAND2_7154 ( R2144_U160 , R2144_U58 , R2144_U158 );
nand NAND2_7155 ( R2144_U161 , U2749 , R2144_U199 );
nand NAND2_7156 ( R2144_U162 , U2750 , R2144_U184 );
nand NAND2_7157 ( R2144_U163 , R2144_U116 , R2144_U109 );
nand NAND2_7158 ( R2144_U164 , U2355 , R2144_U68 );
nand NAND2_7159 ( R2144_U165 , U2762 , R2144_U12 );
nand NAND2_7160 ( R2144_U166 , U2355 , R2144_U69 );
nand NAND2_7161 ( R2144_U167 , U2761 , R2144_U12 );
nand NAND2_7162 ( R2144_U168 , U2355 , R2144_U70 );
nand NAND2_7163 ( R2144_U169 , U2763 , R2144_U12 );
nand NAND2_7164 ( R2144_U170 , R2144_U169 , R2144_U168 );
nand NAND2_7165 ( R2144_U171 , U2355 , R2144_U68 );
nand NAND2_7166 ( R2144_U172 , U2762 , R2144_U12 );
nand NAND2_7167 ( R2144_U173 , R2144_U172 , R2144_U171 );
nand NAND2_7168 ( R2144_U174 , U2355 , R2144_U70 );
nand NAND2_7169 ( R2144_U175 , U2763 , R2144_U12 );
nand NAND2_7170 ( R2144_U176 , U2355 , R2144_U71 );
nand NAND2_7171 ( R2144_U177 , U2764 , R2144_U12 );
nand NAND2_7172 ( R2144_U178 , R2144_U177 , R2144_U176 );
nand NAND2_7173 ( R2144_U179 , U2355 , R2144_U69 );
nand NAND2_7174 ( R2144_U180 , U2761 , R2144_U12 );
nand NAND2_7175 ( R2144_U181 , R2144_U180 , R2144_U179 );
nand NAND2_7176 ( R2144_U182 , U2355 , R2144_U72 );
nand NAND2_7177 ( R2144_U183 , U2766 , R2144_U12 );
nand NAND2_7178 ( R2144_U184 , R2144_U183 , R2144_U182 );
nand NAND2_7179 ( R2144_U185 , U2355 , R2144_U73 );
nand NAND2_7180 ( R2144_U186 , U2767 , R2144_U12 );
not NOT1_7181 ( R2144_U187 , R2144_U28 );
nand NAND2_7182 ( R2144_U188 , U2355 , R2144_U74 );
nand NAND2_7183 ( R2144_U189 , U2768 , R2144_U12 );
nand NAND2_7184 ( R2144_U190 , U2355 , R2144_U74 );
nand NAND2_7185 ( R2144_U191 , U2768 , R2144_U12 );
nand NAND2_7186 ( R2144_U192 , R2144_U191 , R2144_U190 );
nand NAND2_7187 ( R2144_U193 , U2355 , R2144_U72 );
nand NAND2_7188 ( R2144_U194 , U2766 , R2144_U12 );
nand NAND2_7189 ( R2144_U195 , U2355 , R2144_U75 );
nand NAND2_7190 ( R2144_U196 , U2765 , R2144_U12 );
nand NAND2_7191 ( R2144_U197 , U2355 , R2144_U75 );
nand NAND2_7192 ( R2144_U198 , U2765 , R2144_U12 );
nand NAND2_7193 ( R2144_U199 , R2144_U198 , R2144_U197 );
nand NAND2_7194 ( R2144_U200 , U2355 , R2144_U71 );
nand NAND2_7195 ( R2144_U201 , U2764 , R2144_U12 );
nand NAND2_7196 ( R2144_U202 , U2355 , R2144_U76 );
nand NAND2_7197 ( R2144_U203 , U2760 , R2144_U12 );
not NOT1_7198 ( R2144_U204 , R2144_U29 );
nand NAND2_7199 ( R2144_U205 , U2355 , R2144_U77 );
nand NAND2_7200 ( R2144_U206 , U2759 , R2144_U12 );
not NOT1_7201 ( R2144_U207 , R2144_U27 );
nand NAND2_7202 ( R2144_U208 , R2144_U122 , R2144_U207 );
nand NAND2_7203 ( R2144_U209 , R2144_U27 , R2144_U78 );
nand NAND2_7204 ( R2144_U210 , R2144_U121 , R2144_U204 );
nand NAND2_7205 ( R2144_U211 , R2144_U29 , R2144_U79 );
nand NAND3_7206 ( R2144_U212 , R2144_U57 , R2144_U124 , R2144_U23 );
nand NAND2_7207 ( R2144_U213 , R2144_U5 , R2144_U108 );
nand NAND2_7208 ( R2144_U214 , R2144_U102 , R2144_U156 );
nand NAND3_7209 ( R2144_U215 , R2144_U59 , R2144_U160 , R2144_U81 );
nand NAND2_7210 ( R2144_U216 , R2144_U149 , R2144_U83 );
nand NAND2_7211 ( R2144_U217 , R2144_U44 , R2144_U123 );
nand NAND2_7212 ( R2144_U218 , R2144_U150 , R2144_U84 );
nand NAND2_7213 ( R2144_U219 , R2144_U46 , R2144_U119 );
nand NAND2_7214 ( R2144_U220 , U2355 , R2144_U85 );
nand NAND2_7215 ( R2144_U221 , U2754 , R2144_U12 );
not NOT1_7216 ( R2144_U222 , R2144_U32 );
nand NAND2_7217 ( R2144_U223 , U2355 , R2144_U86 );
nand NAND2_7218 ( R2144_U224 , U2753 , R2144_U12 );
not NOT1_7219 ( R2144_U225 , R2144_U31 );
nand NAND2_7220 ( R2144_U226 , U2355 , R2144_U87 );
nand NAND2_7221 ( R2144_U227 , U2755 , R2144_U12 );
not NOT1_7222 ( R2144_U228 , R2144_U33 );
nand NAND2_7223 ( R2144_U229 , U2355 , R2144_U88 );
nand NAND2_7224 ( R2144_U230 , U2756 , R2144_U12 );
not NOT1_7225 ( R2144_U231 , R2144_U34 );
nand NAND2_7226 ( R2144_U232 , U2355 , R2144_U89 );
nand NAND2_7227 ( R2144_U233 , U2757 , R2144_U12 );
not NOT1_7228 ( R2144_U234 , R2144_U35 );
nand NAND2_7229 ( R2144_U235 , U2355 , R2144_U90 );
nand NAND2_7230 ( R2144_U236 , U2758 , R2144_U12 );
not NOT1_7231 ( R2144_U237 , R2144_U36 );
nand NAND2_7232 ( R2144_U238 , R2144_U163 , R2144_U91 );
nand NAND2_7233 ( R2144_U239 , R2144_U48 , R2144_U133 );
nand NAND2_7234 ( R2144_U240 , R2144_U187 , U2751 );
nand NAND2_7235 ( R2144_U241 , R2144_U28 , R2144_U14 );
nand NAND2_7236 ( R2144_U242 , R2144_U187 , U2751 );
nand NAND2_7237 ( R2144_U243 , R2144_U28 , R2144_U14 );
nand NAND2_7238 ( R2144_U244 , R2144_U243 , R2144_U242 );
nand NAND2_7239 ( R2144_U245 , R2144_U92 , R2144_U93 );
nand NAND2_7240 ( R2144_U246 , R2144_U130 , R2144_U244 );
nand NAND2_7241 ( R2144_U247 , R2144_U147 , R2144_U225 );
nand NAND2_7242 ( R2144_U248 , R2144_U31 , R2144_U94 );
nand NAND2_7243 ( R2144_U249 , R2144_U222 , R2144_U143 );
nand NAND2_7244 ( R2144_U250 , R2144_U32 , R2144_U26 );
nand NAND2_7245 ( R2144_U251 , R2144_U142 , R2144_U228 );
nand NAND2_7246 ( R2144_U252 , R2144_U33 , R2144_U95 );
nand NAND2_7247 ( R2144_U253 , R2144_U231 , R2144_U141 );
nand NAND2_7248 ( R2144_U254 , R2144_U34 , R2144_U25 );
nand NAND2_7249 ( R2144_U255 , R2144_U140 , R2144_U234 );
nand NAND2_7250 ( R2144_U256 , R2144_U35 , R2144_U96 );
nand NAND2_7251 ( R2144_U257 , R2144_U139 , R2144_U237 );
nand NAND2_7252 ( R2144_U258 , R2144_U36 , R2144_U97 );
nand NAND2_7253 ( R2144_U259 , U2355 , R2144_U98 );
nand NAND2_7254 ( R2144_U260 , R2144_U148 , R2144_U12 );
or OR2_7255 ( LT_589_U6 , LT_589_U8 , U2673 );
and AND2_7256 ( LT_589_U7 , R584_U7 , R584_U6 );
nor nor_7257 ( LT_589_U8 , LT_589_U7 , R584_U9 , R584_U8 );
not NOT1_7258 ( R584_U6 , U2676 );
not NOT1_7259 ( R584_U7 , U2677 );
not NOT1_7260 ( R584_U8 , U2674 );
not NOT1_7261 ( R584_U9 , U2675 );
not NOT1_7262 ( R2099_U4 , U4178 );
not NOT1_7263 ( R2099_U5 , U4177 );
not NOT1_7264 ( R2099_U6 , U2678 );
nand NAND2_7265 ( R2099_U7 , R2099_U88 , R2099_U137 );
nand NAND2_7266 ( R2099_U8 , R2099_U89 , R2099_U155 );
nand NAND2_7267 ( R2099_U9 , R2099_U90 , R2099_U157 );
nand NAND2_7268 ( R2099_U10 , R2099_U91 , R2099_U159 );
nand NAND2_7269 ( R2099_U11 , R2099_U92 , R2099_U161 );
nand NAND2_7270 ( R2099_U12 , R2099_U93 , R2099_U163 );
nand NAND2_7271 ( R2099_U13 , R2099_U94 , R2099_U165 );
nand NAND2_7272 ( R2099_U14 , R2099_U95 , R2099_U167 );
nand NAND2_7273 ( R2099_U15 , R2099_U169 , R2099_U55 );
nand NAND2_7274 ( R2099_U16 , R2099_U170 , R2099_U54 );
nand NAND2_7275 ( R2099_U17 , R2099_U171 , R2099_U53 );
nand NAND2_7276 ( R2099_U18 , R2099_U172 , R2099_U52 );
nand NAND2_7277 ( R2099_U19 , R2099_U173 , R2099_U51 );
nand NAND2_7278 ( R2099_U20 , R2099_U174 , R2099_U50 );
nand NAND2_7279 ( R2099_U21 , R2099_U175 , R2099_U49 );
nand NAND2_7280 ( R2099_U22 , R2099_U176 , R2099_U48 );
nand NAND2_7281 ( R2099_U23 , R2099_U177 , R2099_U47 );
nand NAND2_7282 ( R2099_U24 , R2099_U178 , R2099_U46 );
nand NAND2_7283 ( R2099_U25 , R2099_U179 , R2099_U45 );
nand NAND2_7284 ( R2099_U26 , R2099_U210 , R2099_U209 );
nand NAND2_7285 ( R2099_U27 , R2099_U183 , R2099_U182 );
nand NAND2_7286 ( R2099_U28 , R2099_U204 , R2099_U203 );
nand NAND2_7287 ( R2099_U29 , R2099_U207 , R2099_U206 );
nand NAND2_7288 ( R2099_U30 , R2099_U198 , R2099_U197 );
nand NAND2_7289 ( R2099_U31 , R2099_U201 , R2099_U200 );
nand NAND2_7290 ( R2099_U32 , R2099_U186 , R2099_U185 );
nand NAND2_7291 ( R2099_U33 , R2099_U189 , R2099_U188 );
nand NAND2_7292 ( R2099_U34 , R2099_U195 , R2099_U194 );
nand NAND2_7293 ( R2099_U35 , R2099_U192 , R2099_U191 );
nand NAND2_7294 ( R2099_U36 , R2099_U213 , R2099_U212 );
nand NAND2_7295 ( R2099_U37 , R2099_U215 , R2099_U214 );
nand NAND2_7296 ( R2099_U38 , R2099_U217 , R2099_U216 );
nand NAND2_7297 ( R2099_U39 , R2099_U219 , R2099_U218 );
nand NAND2_7298 ( R2099_U40 , R2099_U221 , R2099_U220 );
nand NAND2_7299 ( R2099_U41 , R2099_U223 , R2099_U222 );
nand NAND2_7300 ( R2099_U42 , R2099_U225 , R2099_U224 );
nand NAND2_7301 ( R2099_U43 , R2099_U284 , R2099_U283 );
nand NAND2_7302 ( R2099_U44 , R2099_U287 , R2099_U286 );
nand NAND2_7303 ( R2099_U45 , R2099_U227 , R2099_U226 );
nand NAND2_7304 ( R2099_U46 , R2099_U230 , R2099_U229 );
nand NAND2_7305 ( R2099_U47 , R2099_U233 , R2099_U232 );
nand NAND2_7306 ( R2099_U48 , R2099_U236 , R2099_U235 );
nand NAND2_7307 ( R2099_U49 , R2099_U239 , R2099_U238 );
nand NAND2_7308 ( R2099_U50 , R2099_U242 , R2099_U241 );
nand NAND2_7309 ( R2099_U51 , R2099_U245 , R2099_U244 );
nand NAND2_7310 ( R2099_U52 , R2099_U248 , R2099_U247 );
nand NAND2_7311 ( R2099_U53 , R2099_U251 , R2099_U250 );
nand NAND2_7312 ( R2099_U54 , R2099_U254 , R2099_U253 );
nand NAND2_7313 ( R2099_U55 , R2099_U257 , R2099_U256 );
nand NAND2_7314 ( R2099_U56 , R2099_U278 , R2099_U277 );
nand NAND2_7315 ( R2099_U57 , R2099_U281 , R2099_U280 );
nand NAND2_7316 ( R2099_U58 , R2099_U272 , R2099_U271 );
nand NAND2_7317 ( R2099_U59 , R2099_U275 , R2099_U274 );
nand NAND2_7318 ( R2099_U60 , R2099_U266 , R2099_U265 );
nand NAND2_7319 ( R2099_U61 , R2099_U269 , R2099_U268 );
nand NAND2_7320 ( R2099_U62 , R2099_U260 , R2099_U259 );
nand NAND2_7321 ( R2099_U63 , R2099_U263 , R2099_U262 );
nand NAND2_7322 ( R2099_U64 , R2099_U293 , R2099_U292 );
nand NAND2_7323 ( R2099_U65 , R2099_U295 , R2099_U294 );
nand NAND2_7324 ( R2099_U66 , R2099_U299 , R2099_U298 );
nand NAND2_7325 ( R2099_U67 , R2099_U301 , R2099_U300 );
nand NAND2_7326 ( R2099_U68 , R2099_U303 , R2099_U302 );
nand NAND2_7327 ( R2099_U69 , R2099_U305 , R2099_U304 );
nand NAND2_7328 ( R2099_U70 , R2099_U307 , R2099_U306 );
nand NAND2_7329 ( R2099_U71 , R2099_U309 , R2099_U308 );
nand NAND2_7330 ( R2099_U72 , R2099_U311 , R2099_U310 );
nand NAND2_7331 ( R2099_U73 , R2099_U313 , R2099_U312 );
nand NAND2_7332 ( R2099_U74 , R2099_U315 , R2099_U314 );
nand NAND2_7333 ( R2099_U75 , R2099_U317 , R2099_U316 );
nand NAND2_7334 ( R2099_U76 , R2099_U326 , R2099_U325 );
nand NAND2_7335 ( R2099_U77 , R2099_U328 , R2099_U327 );
nand NAND2_7336 ( R2099_U78 , R2099_U330 , R2099_U329 );
nand NAND2_7337 ( R2099_U79 , R2099_U332 , R2099_U331 );
nand NAND2_7338 ( R2099_U80 , R2099_U334 , R2099_U333 );
nand NAND2_7339 ( R2099_U81 , R2099_U336 , R2099_U335 );
nand NAND2_7340 ( R2099_U82 , R2099_U338 , R2099_U337 );
nand NAND2_7341 ( R2099_U83 , R2099_U340 , R2099_U339 );
nand NAND2_7342 ( R2099_U84 , R2099_U342 , R2099_U341 );
nand NAND2_7343 ( R2099_U85 , R2099_U344 , R2099_U343 );
nand NAND2_7344 ( R2099_U86 , R2099_U349 , R2099_U348 );
nand NAND2_7345 ( R2099_U87 , R2099_U324 , R2099_U323 );
and AND2_7346 ( R2099_U88 , R2099_U34 , R2099_U35 );
and AND2_7347 ( R2099_U89 , R2099_U31 , R2099_U30 );
and AND2_7348 ( R2099_U90 , R2099_U29 , R2099_U28 );
and AND2_7349 ( R2099_U91 , R2099_U26 , R2099_U27 );
and AND2_7350 ( R2099_U92 , R2099_U63 , R2099_U62 );
and AND2_7351 ( R2099_U93 , R2099_U61 , R2099_U60 );
and AND2_7352 ( R2099_U94 , R2099_U59 , R2099_U58 );
and AND2_7353 ( R2099_U95 , R2099_U57 , R2099_U56 );
and AND2_7354 ( R2099_U96 , R2099_U44 , R2099_U43 );
nand NAND2_7355 ( R2099_U97 , R2099_U290 , R2099_U289 );
nand NAND2_7356 ( R2099_U98 , R2099_U346 , R2099_U345 );
not NOT1_7357 ( R2099_U99 , U2702 );
not NOT1_7358 ( R2099_U100 , U2710 );
not NOT1_7359 ( R2099_U101 , U2709 );
not NOT1_7360 ( R2099_U102 , U2708 );
not NOT1_7361 ( R2099_U103 , U2707 );
not NOT1_7362 ( R2099_U104 , U2706 );
not NOT1_7363 ( R2099_U105 , U2705 );
not NOT1_7364 ( R2099_U106 , U2704 );
not NOT1_7365 ( R2099_U107 , U2703 );
not NOT1_7366 ( R2099_U108 , U2701 );
nand NAND2_7367 ( R2099_U109 , R2099_U159 , R2099_U27 );
nand NAND2_7368 ( R2099_U110 , R2099_U157 , R2099_U28 );
nand NAND2_7369 ( R2099_U111 , R2099_U155 , R2099_U30 );
nand NAND2_7370 ( R2099_U112 , R2099_U35 , R2099_U137 );
not NOT1_7371 ( R2099_U113 , U2682 );
not NOT1_7372 ( R2099_U114 , U2683 );
not NOT1_7373 ( R2099_U115 , U2684 );
not NOT1_7374 ( R2099_U116 , U2685 );
not NOT1_7375 ( R2099_U117 , U2686 );
not NOT1_7376 ( R2099_U118 , U2687 );
not NOT1_7377 ( R2099_U119 , U2688 );
not NOT1_7378 ( R2099_U120 , U2689 );
not NOT1_7379 ( R2099_U121 , U2690 );
not NOT1_7380 ( R2099_U122 , U2691 );
not NOT1_7381 ( R2099_U123 , U2692 );
not NOT1_7382 ( R2099_U124 , U2700 );
not NOT1_7383 ( R2099_U125 , U2699 );
not NOT1_7384 ( R2099_U126 , U2698 );
not NOT1_7385 ( R2099_U127 , U2697 );
not NOT1_7386 ( R2099_U128 , U2696 );
not NOT1_7387 ( R2099_U129 , U2695 );
not NOT1_7388 ( R2099_U130 , U2694 );
not NOT1_7389 ( R2099_U131 , U2693 );
not NOT1_7390 ( R2099_U132 , U2680 );
not NOT1_7391 ( R2099_U133 , U2681 );
not NOT1_7392 ( R2099_U134 , U2679 );
nand NAND2_7393 ( R2099_U135 , R2099_U96 , R2099_U180 );
nand NAND2_7394 ( R2099_U136 , R2099_U180 , R2099_U44 );
nand NAND2_7395 ( R2099_U137 , R2099_U152 , R2099_U151 );
and AND2_7396 ( R2099_U138 , R2099_U297 , R2099_U296 );
and AND2_7397 ( R2099_U139 , R2099_U319 , R2099_U318 );
nand NAND2_7398 ( R2099_U140 , R2099_U148 , R2099_U147 );
nand NAND2_7399 ( R2099_U141 , R2099_U167 , R2099_U56 );
nand NAND2_7400 ( R2099_U142 , R2099_U165 , R2099_U58 );
nand NAND2_7401 ( R2099_U143 , R2099_U163 , R2099_U60 );
nand NAND2_7402 ( R2099_U144 , R2099_U161 , R2099_U62 );
not NOT1_7403 ( R2099_U145 , R2099_U135 );
or OR2_7404 ( R2099_U146 , U4178 , U4177 );
nand NAND2_7405 ( R2099_U147 , R2099_U32 , R2099_U146 );
nand NAND2_7406 ( R2099_U148 , U4177 , U4178 );
not NOT1_7407 ( R2099_U149 , R2099_U140 );
nand NAND2_7408 ( R2099_U150 , R2099_U190 , R2099_U6 );
nand NAND2_7409 ( R2099_U151 , R2099_U150 , R2099_U140 );
nand NAND2_7410 ( R2099_U152 , U2678 , R2099_U33 );
not NOT1_7411 ( R2099_U153 , R2099_U137 );
not NOT1_7412 ( R2099_U154 , R2099_U112 );
not NOT1_7413 ( R2099_U155 , R2099_U7 );
not NOT1_7414 ( R2099_U156 , R2099_U111 );
not NOT1_7415 ( R2099_U157 , R2099_U8 );
not NOT1_7416 ( R2099_U158 , R2099_U110 );
not NOT1_7417 ( R2099_U159 , R2099_U9 );
not NOT1_7418 ( R2099_U160 , R2099_U109 );
not NOT1_7419 ( R2099_U161 , R2099_U10 );
not NOT1_7420 ( R2099_U162 , R2099_U144 );
not NOT1_7421 ( R2099_U163 , R2099_U11 );
not NOT1_7422 ( R2099_U164 , R2099_U143 );
not NOT1_7423 ( R2099_U165 , R2099_U12 );
not NOT1_7424 ( R2099_U166 , R2099_U142 );
not NOT1_7425 ( R2099_U167 , R2099_U13 );
not NOT1_7426 ( R2099_U168 , R2099_U141 );
not NOT1_7427 ( R2099_U169 , R2099_U14 );
not NOT1_7428 ( R2099_U170 , R2099_U15 );
not NOT1_7429 ( R2099_U171 , R2099_U16 );
not NOT1_7430 ( R2099_U172 , R2099_U17 );
not NOT1_7431 ( R2099_U173 , R2099_U18 );
not NOT1_7432 ( R2099_U174 , R2099_U19 );
not NOT1_7433 ( R2099_U175 , R2099_U20 );
not NOT1_7434 ( R2099_U176 , R2099_U21 );
not NOT1_7435 ( R2099_U177 , R2099_U22 );
not NOT1_7436 ( R2099_U178 , R2099_U23 );
not NOT1_7437 ( R2099_U179 , R2099_U24 );
not NOT1_7438 ( R2099_U180 , R2099_U25 );
not NOT1_7439 ( R2099_U181 , R2099_U136 );
nand NAND2_7440 ( R2099_U182 , U4178 , R2099_U99 );
nand NAND2_7441 ( R2099_U183 , U2702 , R2099_U4 );
not NOT1_7442 ( R2099_U184 , R2099_U27 );
nand NAND2_7443 ( R2099_U185 , U4178 , R2099_U100 );
nand NAND2_7444 ( R2099_U186 , U2710 , R2099_U4 );
not NOT1_7445 ( R2099_U187 , R2099_U32 );
nand NAND2_7446 ( R2099_U188 , U4178 , R2099_U101 );
nand NAND2_7447 ( R2099_U189 , U2709 , R2099_U4 );
not NOT1_7448 ( R2099_U190 , R2099_U33 );
nand NAND2_7449 ( R2099_U191 , U4178 , R2099_U102 );
nand NAND2_7450 ( R2099_U192 , U2708 , R2099_U4 );
not NOT1_7451 ( R2099_U193 , R2099_U35 );
nand NAND2_7452 ( R2099_U194 , U4178 , R2099_U103 );
nand NAND2_7453 ( R2099_U195 , U2707 , R2099_U4 );
not NOT1_7454 ( R2099_U196 , R2099_U34 );
nand NAND2_7455 ( R2099_U197 , U4178 , R2099_U104 );
nand NAND2_7456 ( R2099_U198 , U2706 , R2099_U4 );
not NOT1_7457 ( R2099_U199 , R2099_U30 );
nand NAND2_7458 ( R2099_U200 , U4178 , R2099_U105 );
nand NAND2_7459 ( R2099_U201 , U2705 , R2099_U4 );
not NOT1_7460 ( R2099_U202 , R2099_U31 );
nand NAND2_7461 ( R2099_U203 , U4178 , R2099_U106 );
nand NAND2_7462 ( R2099_U204 , U2704 , R2099_U4 );
not NOT1_7463 ( R2099_U205 , R2099_U28 );
nand NAND2_7464 ( R2099_U206 , U4178 , R2099_U107 );
nand NAND2_7465 ( R2099_U207 , U2703 , R2099_U4 );
not NOT1_7466 ( R2099_U208 , R2099_U29 );
nand NAND2_7467 ( R2099_U209 , U4178 , R2099_U108 );
nand NAND2_7468 ( R2099_U210 , U2701 , R2099_U4 );
not NOT1_7469 ( R2099_U211 , R2099_U26 );
nand NAND2_7470 ( R2099_U212 , R2099_U160 , R2099_U211 );
nand NAND2_7471 ( R2099_U213 , R2099_U26 , R2099_U109 );
nand NAND2_7472 ( R2099_U214 , R2099_U184 , R2099_U159 );
nand NAND2_7473 ( R2099_U215 , R2099_U27 , R2099_U9 );
nand NAND2_7474 ( R2099_U216 , R2099_U158 , R2099_U208 );
nand NAND2_7475 ( R2099_U217 , R2099_U29 , R2099_U110 );
nand NAND2_7476 ( R2099_U218 , R2099_U205 , R2099_U157 );
nand NAND2_7477 ( R2099_U219 , R2099_U28 , R2099_U8 );
nand NAND2_7478 ( R2099_U220 , R2099_U156 , R2099_U202 );
nand NAND2_7479 ( R2099_U221 , R2099_U31 , R2099_U111 );
nand NAND2_7480 ( R2099_U222 , R2099_U199 , R2099_U155 );
nand NAND2_7481 ( R2099_U223 , R2099_U30 , R2099_U7 );
nand NAND2_7482 ( R2099_U224 , R2099_U154 , R2099_U196 );
nand NAND2_7483 ( R2099_U225 , R2099_U34 , R2099_U112 );
nand NAND2_7484 ( R2099_U226 , U4178 , R2099_U113 );
nand NAND2_7485 ( R2099_U227 , U2682 , R2099_U4 );
not NOT1_7486 ( R2099_U228 , R2099_U45 );
nand NAND2_7487 ( R2099_U229 , U4178 , R2099_U114 );
nand NAND2_7488 ( R2099_U230 , U2683 , R2099_U4 );
not NOT1_7489 ( R2099_U231 , R2099_U46 );
nand NAND2_7490 ( R2099_U232 , U4178 , R2099_U115 );
nand NAND2_7491 ( R2099_U233 , U2684 , R2099_U4 );
not NOT1_7492 ( R2099_U234 , R2099_U47 );
nand NAND2_7493 ( R2099_U235 , U4178 , R2099_U116 );
nand NAND2_7494 ( R2099_U236 , U2685 , R2099_U4 );
not NOT1_7495 ( R2099_U237 , R2099_U48 );
nand NAND2_7496 ( R2099_U238 , U4178 , R2099_U117 );
nand NAND2_7497 ( R2099_U239 , U2686 , R2099_U4 );
not NOT1_7498 ( R2099_U240 , R2099_U49 );
nand NAND2_7499 ( R2099_U241 , U4178 , R2099_U118 );
nand NAND2_7500 ( R2099_U242 , U2687 , R2099_U4 );
not NOT1_7501 ( R2099_U243 , R2099_U50 );
nand NAND2_7502 ( R2099_U244 , U4178 , R2099_U119 );
nand NAND2_7503 ( R2099_U245 , U2688 , R2099_U4 );
not NOT1_7504 ( R2099_U246 , R2099_U51 );
nand NAND2_7505 ( R2099_U247 , U4178 , R2099_U120 );
nand NAND2_7506 ( R2099_U248 , U2689 , R2099_U4 );
not NOT1_7507 ( R2099_U249 , R2099_U52 );
nand NAND2_7508 ( R2099_U250 , U4178 , R2099_U121 );
nand NAND2_7509 ( R2099_U251 , U2690 , R2099_U4 );
not NOT1_7510 ( R2099_U252 , R2099_U53 );
nand NAND2_7511 ( R2099_U253 , U4178 , R2099_U122 );
nand NAND2_7512 ( R2099_U254 , U2691 , R2099_U4 );
not NOT1_7513 ( R2099_U255 , R2099_U54 );
nand NAND2_7514 ( R2099_U256 , U4178 , R2099_U123 );
nand NAND2_7515 ( R2099_U257 , U2692 , R2099_U4 );
not NOT1_7516 ( R2099_U258 , R2099_U55 );
nand NAND2_7517 ( R2099_U259 , U4178 , R2099_U124 );
nand NAND2_7518 ( R2099_U260 , U2700 , R2099_U4 );
not NOT1_7519 ( R2099_U261 , R2099_U62 );
nand NAND2_7520 ( R2099_U262 , U4178 , R2099_U125 );
nand NAND2_7521 ( R2099_U263 , U2699 , R2099_U4 );
not NOT1_7522 ( R2099_U264 , R2099_U63 );
nand NAND2_7523 ( R2099_U265 , U4178 , R2099_U126 );
nand NAND2_7524 ( R2099_U266 , U2698 , R2099_U4 );
not NOT1_7525 ( R2099_U267 , R2099_U60 );
nand NAND2_7526 ( R2099_U268 , U4178 , R2099_U127 );
nand NAND2_7527 ( R2099_U269 , U2697 , R2099_U4 );
not NOT1_7528 ( R2099_U270 , R2099_U61 );
nand NAND2_7529 ( R2099_U271 , U4178 , R2099_U128 );
nand NAND2_7530 ( R2099_U272 , U2696 , R2099_U4 );
not NOT1_7531 ( R2099_U273 , R2099_U58 );
nand NAND2_7532 ( R2099_U274 , U4178 , R2099_U129 );
nand NAND2_7533 ( R2099_U275 , U2695 , R2099_U4 );
not NOT1_7534 ( R2099_U276 , R2099_U59 );
nand NAND2_7535 ( R2099_U277 , U4178 , R2099_U130 );
nand NAND2_7536 ( R2099_U278 , U2694 , R2099_U4 );
not NOT1_7537 ( R2099_U279 , R2099_U56 );
nand NAND2_7538 ( R2099_U280 , U4178 , R2099_U131 );
nand NAND2_7539 ( R2099_U281 , U2693 , R2099_U4 );
not NOT1_7540 ( R2099_U282 , R2099_U57 );
nand NAND2_7541 ( R2099_U283 , U4178 , R2099_U132 );
nand NAND2_7542 ( R2099_U284 , U2680 , R2099_U4 );
not NOT1_7543 ( R2099_U285 , R2099_U43 );
nand NAND2_7544 ( R2099_U286 , U4178 , R2099_U133 );
nand NAND2_7545 ( R2099_U287 , U2681 , R2099_U4 );
not NOT1_7546 ( R2099_U288 , R2099_U44 );
nand NAND2_7547 ( R2099_U289 , U4178 , R2099_U134 );
nand NAND2_7548 ( R2099_U290 , U2679 , R2099_U4 );
not NOT1_7549 ( R2099_U291 , R2099_U97 );
nand NAND2_7550 ( R2099_U292 , R2099_U145 , R2099_U291 );
nand NAND2_7551 ( R2099_U293 , R2099_U97 , R2099_U135 );
nand NAND2_7552 ( R2099_U294 , R2099_U181 , R2099_U285 );
nand NAND2_7553 ( R2099_U295 , R2099_U43 , R2099_U136 );
nand NAND2_7554 ( R2099_U296 , R2099_U153 , R2099_U193 );
nand NAND2_7555 ( R2099_U297 , R2099_U35 , R2099_U137 );
nand NAND2_7556 ( R2099_U298 , R2099_U288 , R2099_U180 );
nand NAND2_7557 ( R2099_U299 , R2099_U44 , R2099_U25 );
nand NAND2_7558 ( R2099_U300 , R2099_U228 , R2099_U179 );
nand NAND2_7559 ( R2099_U301 , R2099_U45 , R2099_U24 );
nand NAND2_7560 ( R2099_U302 , R2099_U231 , R2099_U178 );
nand NAND2_7561 ( R2099_U303 , R2099_U46 , R2099_U23 );
nand NAND2_7562 ( R2099_U304 , R2099_U234 , R2099_U177 );
nand NAND2_7563 ( R2099_U305 , R2099_U47 , R2099_U22 );
nand NAND2_7564 ( R2099_U306 , R2099_U237 , R2099_U176 );
nand NAND2_7565 ( R2099_U307 , R2099_U48 , R2099_U21 );
nand NAND2_7566 ( R2099_U308 , R2099_U240 , R2099_U175 );
nand NAND2_7567 ( R2099_U309 , R2099_U49 , R2099_U20 );
nand NAND2_7568 ( R2099_U310 , R2099_U243 , R2099_U174 );
nand NAND2_7569 ( R2099_U311 , R2099_U50 , R2099_U19 );
nand NAND2_7570 ( R2099_U312 , R2099_U246 , R2099_U173 );
nand NAND2_7571 ( R2099_U313 , R2099_U51 , R2099_U18 );
nand NAND2_7572 ( R2099_U314 , R2099_U249 , R2099_U172 );
nand NAND2_7573 ( R2099_U315 , R2099_U52 , R2099_U17 );
nand NAND2_7574 ( R2099_U316 , R2099_U252 , R2099_U171 );
nand NAND2_7575 ( R2099_U317 , R2099_U53 , R2099_U16 );
nand NAND2_7576 ( R2099_U318 , R2099_U190 , U2678 );
nand NAND2_7577 ( R2099_U319 , R2099_U33 , R2099_U6 );
nand NAND2_7578 ( R2099_U320 , R2099_U190 , U2678 );
nand NAND2_7579 ( R2099_U321 , R2099_U33 , R2099_U6 );
nand NAND2_7580 ( R2099_U322 , R2099_U321 , R2099_U320 );
nand NAND2_7581 ( R2099_U323 , R2099_U139 , R2099_U140 );
nand NAND2_7582 ( R2099_U324 , R2099_U149 , R2099_U322 );
nand NAND2_7583 ( R2099_U325 , R2099_U255 , R2099_U170 );
nand NAND2_7584 ( R2099_U326 , R2099_U54 , R2099_U15 );
nand NAND2_7585 ( R2099_U327 , R2099_U258 , R2099_U169 );
nand NAND2_7586 ( R2099_U328 , R2099_U55 , R2099_U14 );
nand NAND2_7587 ( R2099_U329 , R2099_U168 , R2099_U282 );
nand NAND2_7588 ( R2099_U330 , R2099_U57 , R2099_U141 );
nand NAND2_7589 ( R2099_U331 , R2099_U279 , R2099_U167 );
nand NAND2_7590 ( R2099_U332 , R2099_U56 , R2099_U13 );
nand NAND2_7591 ( R2099_U333 , R2099_U166 , R2099_U276 );
nand NAND2_7592 ( R2099_U334 , R2099_U59 , R2099_U142 );
nand NAND2_7593 ( R2099_U335 , R2099_U273 , R2099_U165 );
nand NAND2_7594 ( R2099_U336 , R2099_U58 , R2099_U12 );
nand NAND2_7595 ( R2099_U337 , R2099_U164 , R2099_U270 );
nand NAND2_7596 ( R2099_U338 , R2099_U61 , R2099_U143 );
nand NAND2_7597 ( R2099_U339 , R2099_U267 , R2099_U163 );
nand NAND2_7598 ( R2099_U340 , R2099_U60 , R2099_U11 );
nand NAND2_7599 ( R2099_U341 , R2099_U162 , R2099_U264 );
nand NAND2_7600 ( R2099_U342 , R2099_U63 , R2099_U144 );
nand NAND2_7601 ( R2099_U343 , R2099_U261 , R2099_U161 );
nand NAND2_7602 ( R2099_U344 , R2099_U62 , R2099_U10 );
nand NAND2_7603 ( R2099_U345 , U4177 , R2099_U4 );
nand NAND2_7604 ( R2099_U346 , U4178 , R2099_U5 );
not NOT1_7605 ( R2099_U347 , R2099_U98 );
nand NAND2_7606 ( R2099_U348 , R2099_U32 , R2099_U347 );
nand NAND2_7607 ( R2099_U349 , R2099_U98 , R2099_U187 );
not NOT1_7608 ( R2167_U6 , U2716 );
not NOT1_7609 ( R2167_U7 , U2714 );
not NOT1_7610 ( R2167_U8 , U2720 );
not NOT1_7611 ( R2167_U9 , U2719 );
not NOT1_7612 ( R2167_U10 , U2713 );
not NOT1_7613 ( R2167_U11 , U2712 );
not NOT1_7614 ( R2167_U12 , U2718 );
not NOT1_7615 ( R2167_U13 , U2717 );
not NOT1_7616 ( R2167_U14 , U2711 );
not NOT1_7617 ( R2167_U15 , U2356 );
not NOT1_7618 ( R2167_U16 , STATE2_REG_0_ );
nand NAND2_7619 ( R2167_U17 , R2167_U50 , R2167_U49 );
and AND2_7620 ( R2167_U18 , R2167_U29 , R2167_U30 );
and AND2_7621 ( R2167_U19 , R2167_U32 , R2167_U33 );
and AND2_7622 ( R2167_U20 , R2167_U35 , R2167_U36 );
and AND2_7623 ( R2167_U21 , R2167_U38 , R2167_U39 );
not NOT1_7624 ( R2167_U22 , U2721 );
not NOT1_7625 ( R2167_U23 , U2722 );
nand NAND2_7626 ( R2167_U24 , U2715 , R2167_U23 );
nand NAND2_7627 ( R2167_U25 , U2715 , R2167_U22 );
or OR2_7628 ( R2167_U26 , U2721 , U2722 );
nand NAND2_7629 ( R2167_U27 , U2714 , R2167_U8 );
nand NAND4_7630 ( R2167_U28 , R2167_U27 , R2167_U26 , R2167_U25 , R2167_U24 );
nand NAND2_7631 ( R2167_U29 , U2720 , R2167_U7 );
nand NAND2_7632 ( R2167_U30 , U2719 , R2167_U10 );
nand NAND2_7633 ( R2167_U31 , R2167_U18 , R2167_U28 );
nand NAND2_7634 ( R2167_U32 , U2713 , R2167_U9 );
nand NAND2_7635 ( R2167_U33 , U2712 , R2167_U12 );
nand NAND2_7636 ( R2167_U34 , R2167_U19 , R2167_U31 );
nand NAND2_7637 ( R2167_U35 , U2718 , R2167_U11 );
nand NAND2_7638 ( R2167_U36 , U2717 , R2167_U14 );
nand NAND2_7639 ( R2167_U37 , R2167_U20 , R2167_U34 );
nand NAND2_7640 ( R2167_U38 , U2711 , R2167_U13 );
nand NAND2_7641 ( R2167_U39 , U2356 , R2167_U6 );
nand NAND2_7642 ( R2167_U40 , R2167_U21 , R2167_U37 );
nand NAND2_7643 ( R2167_U41 , U2716 , R2167_U15 );
nand NAND2_7644 ( R2167_U42 , R2167_U40 , R2167_U41 );
nand NAND2_7645 ( R2167_U43 , U2716 , R2167_U16 );
nand NAND2_7646 ( R2167_U44 , R2167_U42 , R2167_U6 );
nand NAND2_7647 ( R2167_U45 , R2167_U44 , R2167_U43 );
nand NAND2_7648 ( R2167_U46 , STATE2_REG_0_ , R2167_U6 );
nand NAND2_7649 ( R2167_U47 , U2716 , R2167_U42 );
nand NAND2_7650 ( R2167_U48 , R2167_U47 , R2167_U46 );
nand NAND2_7651 ( R2167_U49 , R2167_U45 , R2167_U15 );
nand NAND2_7652 ( R2167_U50 , U2356 , R2167_U48 );
not NOT1_7653 ( SUB_357_U6 , U3220 );
not NOT1_7654 ( SUB_357_U7 , U3215 );
not NOT1_7655 ( SUB_357_U8 , U3221 );
not NOT1_7656 ( SUB_357_U9 , U3219 );
not NOT1_7657 ( SUB_357_U10 , U3214 );
not NOT1_7658 ( SUB_357_U11 , U3217 );
not NOT1_7659 ( SUB_357_U12 , U3216 );
not NOT1_7660 ( SUB_357_U13 , U3218 );
and AND2_7661 ( LT_563_1260_U6 , LT_563_1260_U9 , LT_563_1260_U8 );
not NOT1_7662 ( LT_563_1260_U7 , U2673 );
nand NAND2_7663 ( LT_563_1260_U8 , R584_U8 , LT_563_1260_U7 );
nand NAND2_7664 ( LT_563_1260_U9 , R584_U9 , LT_563_1260_U7 );
nand NAND2_7665 ( SUB_580_U6 , SUB_580_U10 , SUB_580_U9 );
not NOT1_7666 ( SUB_580_U7 , INSTADDRPOINTER_REG_1_ );
not NOT1_7667 ( SUB_580_U8 , INSTADDRPOINTER_REG_0_ );
nand NAND2_7668 ( SUB_580_U9 , INSTADDRPOINTER_REG_1_ , SUB_580_U8 );
nand NAND2_7669 ( SUB_580_U10 , INSTADDRPOINTER_REG_0_ , SUB_580_U7 );
not NOT1_7670 ( R2096_U4 , REIP_REG_1_ );
not NOT1_7671 ( R2096_U5 , REIP_REG_2_ );
nand NAND2_7672 ( R2096_U6 , REIP_REG_2_ , REIP_REG_1_ );
not NOT1_7673 ( R2096_U7 , REIP_REG_3_ );
nand NAND2_7674 ( R2096_U8 , REIP_REG_3_ , R2096_U94 );
not NOT1_7675 ( R2096_U9 , REIP_REG_4_ );
nand NAND2_7676 ( R2096_U10 , REIP_REG_4_ , R2096_U95 );
not NOT1_7677 ( R2096_U11 , REIP_REG_5_ );
nand NAND2_7678 ( R2096_U12 , REIP_REG_5_ , R2096_U96 );
not NOT1_7679 ( R2096_U13 , REIP_REG_6_ );
nand NAND2_7680 ( R2096_U14 , REIP_REG_6_ , R2096_U97 );
not NOT1_7681 ( R2096_U15 , REIP_REG_7_ );
nand NAND2_7682 ( R2096_U16 , REIP_REG_7_ , R2096_U98 );
not NOT1_7683 ( R2096_U17 , REIP_REG_8_ );
not NOT1_7684 ( R2096_U18 , REIP_REG_9_ );
nand NAND2_7685 ( R2096_U19 , REIP_REG_8_ , R2096_U99 );
nand NAND2_7686 ( R2096_U20 , R2096_U100 , REIP_REG_9_ );
not NOT1_7687 ( R2096_U21 , REIP_REG_10_ );
nand NAND2_7688 ( R2096_U22 , REIP_REG_10_ , R2096_U101 );
not NOT1_7689 ( R2096_U23 , REIP_REG_11_ );
nand NAND2_7690 ( R2096_U24 , REIP_REG_11_ , R2096_U102 );
not NOT1_7691 ( R2096_U25 , REIP_REG_12_ );
nand NAND2_7692 ( R2096_U26 , REIP_REG_12_ , R2096_U103 );
not NOT1_7693 ( R2096_U27 , REIP_REG_13_ );
nand NAND2_7694 ( R2096_U28 , REIP_REG_13_ , R2096_U104 );
not NOT1_7695 ( R2096_U29 , REIP_REG_14_ );
nand NAND2_7696 ( R2096_U30 , REIP_REG_14_ , R2096_U105 );
not NOT1_7697 ( R2096_U31 , REIP_REG_15_ );
nand NAND2_7698 ( R2096_U32 , REIP_REG_15_ , R2096_U106 );
not NOT1_7699 ( R2096_U33 , REIP_REG_16_ );
nand NAND2_7700 ( R2096_U34 , REIP_REG_16_ , R2096_U107 );
not NOT1_7701 ( R2096_U35 , REIP_REG_17_ );
nand NAND2_7702 ( R2096_U36 , REIP_REG_17_ , R2096_U108 );
not NOT1_7703 ( R2096_U37 , REIP_REG_18_ );
nand NAND2_7704 ( R2096_U38 , REIP_REG_18_ , R2096_U109 );
not NOT1_7705 ( R2096_U39 , REIP_REG_19_ );
nand NAND2_7706 ( R2096_U40 , REIP_REG_19_ , R2096_U110 );
not NOT1_7707 ( R2096_U41 , REIP_REG_20_ );
nand NAND2_7708 ( R2096_U42 , REIP_REG_20_ , R2096_U111 );
not NOT1_7709 ( R2096_U43 , REIP_REG_21_ );
nand NAND2_7710 ( R2096_U44 , REIP_REG_21_ , R2096_U112 );
not NOT1_7711 ( R2096_U45 , REIP_REG_22_ );
nand NAND2_7712 ( R2096_U46 , REIP_REG_22_ , R2096_U113 );
not NOT1_7713 ( R2096_U47 , REIP_REG_23_ );
nand NAND2_7714 ( R2096_U48 , REIP_REG_23_ , R2096_U114 );
not NOT1_7715 ( R2096_U49 , REIP_REG_24_ );
nand NAND2_7716 ( R2096_U50 , REIP_REG_24_ , R2096_U115 );
not NOT1_7717 ( R2096_U51 , REIP_REG_25_ );
nand NAND2_7718 ( R2096_U52 , REIP_REG_25_ , R2096_U116 );
not NOT1_7719 ( R2096_U53 , REIP_REG_26_ );
nand NAND2_7720 ( R2096_U54 , REIP_REG_26_ , R2096_U117 );
not NOT1_7721 ( R2096_U55 , REIP_REG_27_ );
nand NAND2_7722 ( R2096_U56 , REIP_REG_27_ , R2096_U118 );
not NOT1_7723 ( R2096_U57 , REIP_REG_28_ );
nand NAND2_7724 ( R2096_U58 , REIP_REG_28_ , R2096_U119 );
not NOT1_7725 ( R2096_U59 , REIP_REG_29_ );
nand NAND2_7726 ( R2096_U60 , REIP_REG_29_ , R2096_U120 );
not NOT1_7727 ( R2096_U61 , REIP_REG_30_ );
nand NAND2_7728 ( R2096_U62 , R2096_U124 , R2096_U123 );
nand NAND2_7729 ( R2096_U63 , R2096_U126 , R2096_U125 );
nand NAND2_7730 ( R2096_U64 , R2096_U128 , R2096_U127 );
nand NAND2_7731 ( R2096_U65 , R2096_U130 , R2096_U129 );
nand NAND2_7732 ( R2096_U66 , R2096_U132 , R2096_U131 );
nand NAND2_7733 ( R2096_U67 , R2096_U134 , R2096_U133 );
nand NAND2_7734 ( R2096_U68 , R2096_U136 , R2096_U135 );
nand NAND2_7735 ( R2096_U69 , R2096_U138 , R2096_U137 );
nand NAND2_7736 ( R2096_U70 , R2096_U140 , R2096_U139 );
nand NAND2_7737 ( R2096_U71 , R2096_U142 , R2096_U141 );
nand NAND2_7738 ( R2096_U72 , R2096_U144 , R2096_U143 );
nand NAND2_7739 ( R2096_U73 , R2096_U146 , R2096_U145 );
nand NAND2_7740 ( R2096_U74 , R2096_U148 , R2096_U147 );
nand NAND2_7741 ( R2096_U75 , R2096_U150 , R2096_U149 );
nand NAND2_7742 ( R2096_U76 , R2096_U152 , R2096_U151 );
nand NAND2_7743 ( R2096_U77 , R2096_U154 , R2096_U153 );
nand NAND2_7744 ( R2096_U78 , R2096_U156 , R2096_U155 );
nand NAND2_7745 ( R2096_U79 , R2096_U158 , R2096_U157 );
nand NAND2_7746 ( R2096_U80 , R2096_U160 , R2096_U159 );
nand NAND2_7747 ( R2096_U81 , R2096_U162 , R2096_U161 );
nand NAND2_7748 ( R2096_U82 , R2096_U164 , R2096_U163 );
nand NAND2_7749 ( R2096_U83 , R2096_U166 , R2096_U165 );
nand NAND2_7750 ( R2096_U84 , R2096_U168 , R2096_U167 );
nand NAND2_7751 ( R2096_U85 , R2096_U170 , R2096_U169 );
nand NAND2_7752 ( R2096_U86 , R2096_U172 , R2096_U171 );
nand NAND2_7753 ( R2096_U87 , R2096_U174 , R2096_U173 );
nand NAND2_7754 ( R2096_U88 , R2096_U176 , R2096_U175 );
nand NAND2_7755 ( R2096_U89 , R2096_U178 , R2096_U177 );
nand NAND2_7756 ( R2096_U90 , R2096_U180 , R2096_U179 );
nand NAND2_7757 ( R2096_U91 , R2096_U182 , R2096_U181 );
not NOT1_7758 ( R2096_U92 , REIP_REG_31_ );
nand NAND2_7759 ( R2096_U93 , REIP_REG_30_ , R2096_U121 );
not NOT1_7760 ( R2096_U94 , R2096_U6 );
not NOT1_7761 ( R2096_U95 , R2096_U8 );
not NOT1_7762 ( R2096_U96 , R2096_U10 );
not NOT1_7763 ( R2096_U97 , R2096_U12 );
not NOT1_7764 ( R2096_U98 , R2096_U14 );
not NOT1_7765 ( R2096_U99 , R2096_U16 );
not NOT1_7766 ( R2096_U100 , R2096_U19 );
not NOT1_7767 ( R2096_U101 , R2096_U20 );
not NOT1_7768 ( R2096_U102 , R2096_U22 );
not NOT1_7769 ( R2096_U103 , R2096_U24 );
not NOT1_7770 ( R2096_U104 , R2096_U26 );
not NOT1_7771 ( R2096_U105 , R2096_U28 );
not NOT1_7772 ( R2096_U106 , R2096_U30 );
not NOT1_7773 ( R2096_U107 , R2096_U32 );
not NOT1_7774 ( R2096_U108 , R2096_U34 );
not NOT1_7775 ( R2096_U109 , R2096_U36 );
not NOT1_7776 ( R2096_U110 , R2096_U38 );
not NOT1_7777 ( R2096_U111 , R2096_U40 );
not NOT1_7778 ( R2096_U112 , R2096_U42 );
not NOT1_7779 ( R2096_U113 , R2096_U44 );
not NOT1_7780 ( R2096_U114 , R2096_U46 );
not NOT1_7781 ( R2096_U115 , R2096_U48 );
not NOT1_7782 ( R2096_U116 , R2096_U50 );
not NOT1_7783 ( R2096_U117 , R2096_U52 );
not NOT1_7784 ( R2096_U118 , R2096_U54 );
not NOT1_7785 ( R2096_U119 , R2096_U56 );
not NOT1_7786 ( R2096_U120 , R2096_U58 );
not NOT1_7787 ( R2096_U121 , R2096_U60 );
not NOT1_7788 ( R2096_U122 , R2096_U93 );
nand NAND2_7789 ( R2096_U123 , REIP_REG_9_ , R2096_U19 );
nand NAND2_7790 ( R2096_U124 , R2096_U100 , R2096_U18 );
nand NAND2_7791 ( R2096_U125 , REIP_REG_8_ , R2096_U16 );
nand NAND2_7792 ( R2096_U126 , R2096_U99 , R2096_U17 );
nand NAND2_7793 ( R2096_U127 , REIP_REG_7_ , R2096_U14 );
nand NAND2_7794 ( R2096_U128 , R2096_U98 , R2096_U15 );
nand NAND2_7795 ( R2096_U129 , REIP_REG_6_ , R2096_U12 );
nand NAND2_7796 ( R2096_U130 , R2096_U97 , R2096_U13 );
nand NAND2_7797 ( R2096_U131 , REIP_REG_5_ , R2096_U10 );
nand NAND2_7798 ( R2096_U132 , R2096_U96 , R2096_U11 );
nand NAND2_7799 ( R2096_U133 , REIP_REG_4_ , R2096_U8 );
nand NAND2_7800 ( R2096_U134 , R2096_U95 , R2096_U9 );
nand NAND2_7801 ( R2096_U135 , REIP_REG_3_ , R2096_U6 );
nand NAND2_7802 ( R2096_U136 , R2096_U94 , R2096_U7 );
nand NAND2_7803 ( R2096_U137 , REIP_REG_31_ , R2096_U93 );
nand NAND2_7804 ( R2096_U138 , R2096_U122 , R2096_U92 );
nand NAND2_7805 ( R2096_U139 , REIP_REG_30_ , R2096_U60 );
nand NAND2_7806 ( R2096_U140 , R2096_U121 , R2096_U61 );
nand NAND2_7807 ( R2096_U141 , REIP_REG_2_ , R2096_U4 );
nand NAND2_7808 ( R2096_U142 , REIP_REG_1_ , R2096_U5 );
nand NAND2_7809 ( R2096_U143 , REIP_REG_29_ , R2096_U58 );
nand NAND2_7810 ( R2096_U144 , R2096_U120 , R2096_U59 );
nand NAND2_7811 ( R2096_U145 , REIP_REG_28_ , R2096_U56 );
nand NAND2_7812 ( R2096_U146 , R2096_U119 , R2096_U57 );
nand NAND2_7813 ( R2096_U147 , REIP_REG_27_ , R2096_U54 );
nand NAND2_7814 ( R2096_U148 , R2096_U118 , R2096_U55 );
nand NAND2_7815 ( R2096_U149 , REIP_REG_26_ , R2096_U52 );
nand NAND2_7816 ( R2096_U150 , R2096_U117 , R2096_U53 );
nand NAND2_7817 ( R2096_U151 , REIP_REG_25_ , R2096_U50 );
nand NAND2_7818 ( R2096_U152 , R2096_U116 , R2096_U51 );
nand NAND2_7819 ( R2096_U153 , REIP_REG_24_ , R2096_U48 );
nand NAND2_7820 ( R2096_U154 , R2096_U115 , R2096_U49 );
nand NAND2_7821 ( R2096_U155 , REIP_REG_23_ , R2096_U46 );
nand NAND2_7822 ( R2096_U156 , R2096_U114 , R2096_U47 );
nand NAND2_7823 ( R2096_U157 , REIP_REG_22_ , R2096_U44 );
nand NAND2_7824 ( R2096_U158 , R2096_U113 , R2096_U45 );
nand NAND2_7825 ( R2096_U159 , REIP_REG_21_ , R2096_U42 );
nand NAND2_7826 ( R2096_U160 , R2096_U112 , R2096_U43 );
nand NAND2_7827 ( R2096_U161 , REIP_REG_20_ , R2096_U40 );
nand NAND2_7828 ( R2096_U162 , R2096_U111 , R2096_U41 );
nand NAND2_7829 ( R2096_U163 , REIP_REG_19_ , R2096_U38 );
nand NAND2_7830 ( R2096_U164 , R2096_U110 , R2096_U39 );
nand NAND2_7831 ( R2096_U165 , REIP_REG_18_ , R2096_U36 );
nand NAND2_7832 ( R2096_U166 , R2096_U109 , R2096_U37 );
nand NAND2_7833 ( R2096_U167 , REIP_REG_17_ , R2096_U34 );
nand NAND2_7834 ( R2096_U168 , R2096_U108 , R2096_U35 );
nand NAND2_7835 ( R2096_U169 , REIP_REG_16_ , R2096_U32 );
nand NAND2_7836 ( R2096_U170 , R2096_U107 , R2096_U33 );
nand NAND2_7837 ( R2096_U171 , REIP_REG_15_ , R2096_U30 );
nand NAND2_7838 ( R2096_U172 , R2096_U106 , R2096_U31 );
nand NAND2_7839 ( R2096_U173 , REIP_REG_14_ , R2096_U28 );
nand NAND2_7840 ( R2096_U174 , R2096_U105 , R2096_U29 );
nand NAND2_7841 ( R2096_U175 , REIP_REG_13_ , R2096_U26 );
nand NAND2_7842 ( R2096_U176 , R2096_U104 , R2096_U27 );
nand NAND2_7843 ( R2096_U177 , REIP_REG_12_ , R2096_U24 );
nand NAND2_7844 ( R2096_U178 , R2096_U103 , R2096_U25 );
nand NAND2_7845 ( R2096_U179 , REIP_REG_11_ , R2096_U22 );
nand NAND2_7846 ( R2096_U180 , R2096_U102 , R2096_U23 );
nand NAND2_7847 ( R2096_U181 , REIP_REG_10_ , R2096_U20 );
nand NAND2_7848 ( R2096_U182 , R2096_U101 , R2096_U21 );
and AND2_7849 ( LT_563_U6 , LT_563_U27 , LT_563_U26 );
not NOT1_7850 ( LT_563_U7 , INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_7851 ( LT_563_U8 , U3478 );
not NOT1_7852 ( LT_563_U9 , U3477 );
not NOT1_7853 ( LT_563_U10 , INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_7854 ( LT_563_U11 , INSTQUEUEWR_ADDR_REG_4_ );
not NOT1_7855 ( LT_563_U12 , U3476 );
and AND2_7856 ( LT_563_U13 , LT_563_U21 , LT_563_U22 );
and AND2_7857 ( LT_563_U14 , LT_563_U24 , LT_563_U25 );
not NOT1_7858 ( LT_563_U15 , U3479 );
not NOT1_7859 ( LT_563_U16 , U3480 );
nand NAND3_7860 ( LT_563_U17 , LT_563_U16 , LT_563_U15 , INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_7861 ( LT_563_U18 , INSTQUEUEWR_ADDR_REG_1_ , LT_563_U15 );
nand NAND2_7862 ( LT_563_U19 , INSTQUEUEWR_ADDR_REG_2_ , LT_563_U8 );
nand NAND4_7863 ( LT_563_U20 , LT_563_U28 , LT_563_U19 , LT_563_U18 , LT_563_U17 );
nand NAND2_7864 ( LT_563_U21 , U3478 , LT_563_U7 );
nand NAND2_7865 ( LT_563_U22 , U3477 , LT_563_U10 );
nand NAND2_7866 ( LT_563_U23 , LT_563_U13 , LT_563_U20 );
nand NAND2_7867 ( LT_563_U24 , INSTQUEUEWR_ADDR_REG_3_ , LT_563_U9 );
nand NAND2_7868 ( LT_563_U25 , INSTQUEUEWR_ADDR_REG_4_ , LT_563_U12 );
nand NAND2_7869 ( LT_563_U26 , LT_563_U14 , LT_563_U23 );
nand NAND2_7870 ( LT_563_U27 , U3476 , LT_563_U11 );
nand NAND3_7871 ( LT_563_U28 , INSTQUEUEWR_ADDR_REG_0_ , INSTQUEUEWR_ADDR_REG_1_ , LT_563_U16 );
nand NAND2_7872 ( R2238_U6 , R2238_U45 , R2238_U44 );
nand NAND2_7873 ( R2238_U7 , R2238_U9 , R2238_U46 );
not NOT1_7874 ( R2238_U8 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_7875 ( R2238_U9 , INSTQUEUERD_ADDR_REG_0_ , R2238_U18 );
not NOT1_7876 ( R2238_U10 , INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_7877 ( R2238_U11 , INSTQUEUERD_ADDR_REG_2_ );
not NOT1_7878 ( R2238_U12 , INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_7879 ( R2238_U13 , INSTQUEUERD_ADDR_REG_3_ );
not NOT1_7880 ( R2238_U14 , INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_7881 ( R2238_U15 , INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_7882 ( R2238_U16 , R2238_U41 , R2238_U40 );
not NOT1_7883 ( R2238_U17 , INSTQUEUERD_ADDR_REG_4_ );
not NOT1_7884 ( R2238_U18 , INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_7885 ( R2238_U19 , R2238_U51 , R2238_U50 );
nand NAND2_7886 ( R2238_U20 , R2238_U56 , R2238_U55 );
nand NAND2_7887 ( R2238_U21 , R2238_U61 , R2238_U60 );
nand NAND2_7888 ( R2238_U22 , R2238_U66 , R2238_U65 );
nand NAND2_7889 ( R2238_U23 , R2238_U48 , R2238_U47 );
nand NAND2_7890 ( R2238_U24 , R2238_U53 , R2238_U52 );
nand NAND2_7891 ( R2238_U25 , R2238_U58 , R2238_U57 );
nand NAND2_7892 ( R2238_U26 , R2238_U63 , R2238_U62 );
nand NAND2_7893 ( R2238_U27 , R2238_U37 , R2238_U36 );
nand NAND2_7894 ( R2238_U28 , R2238_U33 , R2238_U32 );
not NOT1_7895 ( R2238_U29 , INSTQUEUERD_ADDR_REG_1_ );
not NOT1_7896 ( R2238_U30 , R2238_U9 );
nand NAND2_7897 ( R2238_U31 , R2238_U30 , R2238_U10 );
nand NAND2_7898 ( R2238_U32 , R2238_U31 , R2238_U29 );
nand NAND2_7899 ( R2238_U33 , INSTQUEUEWR_ADDR_REG_1_ , R2238_U9 );
not NOT1_7900 ( R2238_U34 , R2238_U28 );
nand NAND2_7901 ( R2238_U35 , INSTQUEUERD_ADDR_REG_2_ , R2238_U12 );
nand NAND2_7902 ( R2238_U36 , R2238_U35 , R2238_U28 );
nand NAND2_7903 ( R2238_U37 , INSTQUEUEWR_ADDR_REG_2_ , R2238_U11 );
not NOT1_7904 ( R2238_U38 , R2238_U27 );
nand NAND2_7905 ( R2238_U39 , INSTQUEUERD_ADDR_REG_3_ , R2238_U14 );
nand NAND2_7906 ( R2238_U40 , R2238_U39 , R2238_U27 );
nand NAND2_7907 ( R2238_U41 , INSTQUEUEWR_ADDR_REG_3_ , R2238_U13 );
not NOT1_7908 ( R2238_U42 , R2238_U16 );
nand NAND2_7909 ( R2238_U43 , INSTQUEUEWR_ADDR_REG_4_ , R2238_U17 );
nand NAND2_7910 ( R2238_U44 , R2238_U42 , R2238_U43 );
nand NAND2_7911 ( R2238_U45 , INSTQUEUERD_ADDR_REG_4_ , R2238_U15 );
nand NAND2_7912 ( R2238_U46 , INSTQUEUEWR_ADDR_REG_0_ , R2238_U8 );
nand NAND2_7913 ( R2238_U47 , INSTQUEUERD_ADDR_REG_4_ , R2238_U15 );
nand NAND2_7914 ( R2238_U48 , INSTQUEUEWR_ADDR_REG_4_ , R2238_U17 );
not NOT1_7915 ( R2238_U49 , R2238_U23 );
nand NAND2_7916 ( R2238_U50 , R2238_U49 , R2238_U42 );
nand NAND2_7917 ( R2238_U51 , R2238_U23 , R2238_U16 );
nand NAND2_7918 ( R2238_U52 , INSTQUEUERD_ADDR_REG_3_ , R2238_U14 );
nand NAND2_7919 ( R2238_U53 , INSTQUEUEWR_ADDR_REG_3_ , R2238_U13 );
not NOT1_7920 ( R2238_U54 , R2238_U24 );
nand NAND2_7921 ( R2238_U55 , R2238_U38 , R2238_U54 );
nand NAND2_7922 ( R2238_U56 , R2238_U24 , R2238_U27 );
nand NAND2_7923 ( R2238_U57 , INSTQUEUERD_ADDR_REG_2_ , R2238_U12 );
nand NAND2_7924 ( R2238_U58 , INSTQUEUEWR_ADDR_REG_2_ , R2238_U11 );
not NOT1_7925 ( R2238_U59 , R2238_U25 );
nand NAND2_7926 ( R2238_U60 , R2238_U34 , R2238_U59 );
nand NAND2_7927 ( R2238_U61 , R2238_U25 , R2238_U28 );
nand NAND2_7928 ( R2238_U62 , INSTQUEUERD_ADDR_REG_1_ , R2238_U10 );
nand NAND2_7929 ( R2238_U63 , INSTQUEUEWR_ADDR_REG_1_ , R2238_U29 );
not NOT1_7930 ( R2238_U64 , R2238_U26 );
nand NAND2_7931 ( R2238_U65 , R2238_U64 , R2238_U30 );
nand NAND2_7932 ( R2238_U66 , R2238_U26 , R2238_U9 );
nand NAND2_7933 ( SUB_450_U6 , SUB_450_U45 , SUB_450_U44 );
nand NAND2_7934 ( SUB_450_U7 , SUB_450_U9 , SUB_450_U46 );
not NOT1_7935 ( SUB_450_U8 , INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_7936 ( SUB_450_U9 , INSTQUEUERD_ADDR_REG_0_ , SUB_450_U18 );
not NOT1_7937 ( SUB_450_U10 , INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_7938 ( SUB_450_U11 , INSTQUEUERD_ADDR_REG_2_ );
not NOT1_7939 ( SUB_450_U12 , INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_7940 ( SUB_450_U13 , INSTQUEUERD_ADDR_REG_3_ );
not NOT1_7941 ( SUB_450_U14 , INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_7942 ( SUB_450_U15 , INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_7943 ( SUB_450_U16 , SUB_450_U41 , SUB_450_U40 );
not NOT1_7944 ( SUB_450_U17 , INSTQUEUERD_ADDR_REG_4_ );
not NOT1_7945 ( SUB_450_U18 , INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_7946 ( SUB_450_U19 , SUB_450_U51 , SUB_450_U50 );
nand NAND2_7947 ( SUB_450_U20 , SUB_450_U56 , SUB_450_U55 );
nand NAND2_7948 ( SUB_450_U21 , SUB_450_U61 , SUB_450_U60 );
nand NAND2_7949 ( SUB_450_U22 , SUB_450_U66 , SUB_450_U65 );
nand NAND2_7950 ( SUB_450_U23 , SUB_450_U48 , SUB_450_U47 );
nand NAND2_7951 ( SUB_450_U24 , SUB_450_U53 , SUB_450_U52 );
nand NAND2_7952 ( SUB_450_U25 , SUB_450_U58 , SUB_450_U57 );
nand NAND2_7953 ( SUB_450_U26 , SUB_450_U63 , SUB_450_U62 );
nand NAND2_7954 ( SUB_450_U27 , SUB_450_U37 , SUB_450_U36 );
nand NAND2_7955 ( SUB_450_U28 , SUB_450_U33 , SUB_450_U32 );
not NOT1_7956 ( SUB_450_U29 , INSTQUEUERD_ADDR_REG_1_ );
not NOT1_7957 ( SUB_450_U30 , SUB_450_U9 );
nand NAND2_7958 ( SUB_450_U31 , SUB_450_U30 , SUB_450_U10 );
nand NAND2_7959 ( SUB_450_U32 , SUB_450_U31 , SUB_450_U29 );
nand NAND2_7960 ( SUB_450_U33 , INSTQUEUEWR_ADDR_REG_1_ , SUB_450_U9 );
not NOT1_7961 ( SUB_450_U34 , SUB_450_U28 );
nand NAND2_7962 ( SUB_450_U35 , INSTQUEUERD_ADDR_REG_2_ , SUB_450_U12 );
nand NAND2_7963 ( SUB_450_U36 , SUB_450_U35 , SUB_450_U28 );
nand NAND2_7964 ( SUB_450_U37 , INSTQUEUEWR_ADDR_REG_2_ , SUB_450_U11 );
not NOT1_7965 ( SUB_450_U38 , SUB_450_U27 );
nand NAND2_7966 ( SUB_450_U39 , INSTQUEUERD_ADDR_REG_3_ , SUB_450_U14 );
nand NAND2_7967 ( SUB_450_U40 , SUB_450_U39 , SUB_450_U27 );
nand NAND2_7968 ( SUB_450_U41 , INSTQUEUEWR_ADDR_REG_3_ , SUB_450_U13 );
not NOT1_7969 ( SUB_450_U42 , SUB_450_U16 );
nand NAND2_7970 ( SUB_450_U43 , INSTQUEUEWR_ADDR_REG_4_ , SUB_450_U17 );
nand NAND2_7971 ( SUB_450_U44 , SUB_450_U42 , SUB_450_U43 );
nand NAND2_7972 ( SUB_450_U45 , INSTQUEUERD_ADDR_REG_4_ , SUB_450_U15 );
nand NAND2_7973 ( SUB_450_U46 , INSTQUEUEWR_ADDR_REG_0_ , SUB_450_U8 );
nand NAND2_7974 ( SUB_450_U47 , INSTQUEUERD_ADDR_REG_4_ , SUB_450_U15 );
nand NAND2_7975 ( SUB_450_U48 , INSTQUEUEWR_ADDR_REG_4_ , SUB_450_U17 );
not NOT1_7976 ( SUB_450_U49 , SUB_450_U23 );
nand NAND2_7977 ( SUB_450_U50 , SUB_450_U49 , SUB_450_U42 );
nand NAND2_7978 ( SUB_450_U51 , SUB_450_U23 , SUB_450_U16 );
nand NAND2_7979 ( SUB_450_U52 , INSTQUEUERD_ADDR_REG_3_ , SUB_450_U14 );
nand NAND2_7980 ( SUB_450_U53 , INSTQUEUEWR_ADDR_REG_3_ , SUB_450_U13 );
not NOT1_7981 ( SUB_450_U54 , SUB_450_U24 );
nand NAND2_7982 ( SUB_450_U55 , SUB_450_U38 , SUB_450_U54 );
nand NAND2_7983 ( SUB_450_U56 , SUB_450_U24 , SUB_450_U27 );
nand NAND2_7984 ( SUB_450_U57 , INSTQUEUERD_ADDR_REG_2_ , SUB_450_U12 );
nand NAND2_7985 ( SUB_450_U58 , INSTQUEUEWR_ADDR_REG_2_ , SUB_450_U11 );
not NOT1_7986 ( SUB_450_U59 , SUB_450_U25 );
nand NAND2_7987 ( SUB_450_U60 , SUB_450_U34 , SUB_450_U59 );
nand NAND2_7988 ( SUB_450_U61 , SUB_450_U25 , SUB_450_U28 );
nand NAND2_7989 ( SUB_450_U62 , INSTQUEUERD_ADDR_REG_1_ , SUB_450_U10 );
nand NAND2_7990 ( SUB_450_U63 , INSTQUEUEWR_ADDR_REG_1_ , SUB_450_U29 );
not NOT1_7991 ( SUB_450_U64 , SUB_450_U26 );
nand NAND2_7992 ( SUB_450_U65 , SUB_450_U64 , SUB_450_U30 );
nand NAND2_7993 ( SUB_450_U66 , SUB_450_U26 , SUB_450_U9 );
not NOT1_7994 ( ADD_371_U4 , U3214 );
nand NAND2_7995 ( ADD_371_U5 , ADD_371_U24 , ADD_371_U32 );
and AND2_7996 ( ADD_371_U6 , ADD_371_U22 , ADD_371_U30 );
not NOT1_7997 ( ADD_371_U7 , U3215 );
not NOT1_7998 ( ADD_371_U8 , U3217 );
nand NAND2_7999 ( ADD_371_U9 , U3217 , ADD_371_U24 );
not NOT1_8000 ( ADD_371_U10 , U3218 );
nand NAND2_8001 ( ADD_371_U11 , U3218 , ADD_371_U28 );
not NOT1_8002 ( ADD_371_U12 , U3219 );
nand NAND2_8003 ( ADD_371_U13 , U3219 , ADD_371_U29 );
not NOT1_8004 ( ADD_371_U14 , U3221 );
not NOT1_8005 ( ADD_371_U15 , U3220 );
not NOT1_8006 ( ADD_371_U16 , U3216 );
nand NAND2_8007 ( ADD_371_U17 , ADD_371_U34 , ADD_371_U33 );
nand NAND2_8008 ( ADD_371_U18 , ADD_371_U36 , ADD_371_U35 );
nand NAND2_8009 ( ADD_371_U19 , ADD_371_U38 , ADD_371_U37 );
nand NAND2_8010 ( ADD_371_U20 , ADD_371_U40 , ADD_371_U39 );
nand NAND2_8011 ( ADD_371_U21 , ADD_371_U44 , ADD_371_U43 );
and AND2_8012 ( ADD_371_U22 , U3221 , U3220 );
nand NAND2_8013 ( ADD_371_U23 , U3220 , ADD_371_U30 );
nand NAND2_8014 ( ADD_371_U24 , ADD_371_U16 , ADD_371_U26 );
and AND2_8015 ( ADD_371_U25 , ADD_371_U42 , ADD_371_U41 );
nand NAND2_8016 ( ADD_371_U26 , U3215 , U3214 );
not NOT1_8017 ( ADD_371_U27 , ADD_371_U24 );
not NOT1_8018 ( ADD_371_U28 , ADD_371_U9 );
not NOT1_8019 ( ADD_371_U29 , ADD_371_U11 );
not NOT1_8020 ( ADD_371_U30 , ADD_371_U13 );
not NOT1_8021 ( ADD_371_U31 , ADD_371_U23 );
nand NAND3_8022 ( ADD_371_U32 , U3215 , U3214 , U3216 );
nand NAND2_8023 ( ADD_371_U33 , U3221 , ADD_371_U23 );
nand NAND2_8024 ( ADD_371_U34 , ADD_371_U31 , ADD_371_U14 );
nand NAND2_8025 ( ADD_371_U35 , U3220 , ADD_371_U13 );
nand NAND2_8026 ( ADD_371_U36 , ADD_371_U30 , ADD_371_U15 );
nand NAND2_8027 ( ADD_371_U37 , U3219 , ADD_371_U11 );
nand NAND2_8028 ( ADD_371_U38 , ADD_371_U29 , ADD_371_U12 );
nand NAND2_8029 ( ADD_371_U39 , U3218 , ADD_371_U9 );
nand NAND2_8030 ( ADD_371_U40 , ADD_371_U28 , ADD_371_U10 );
nand NAND2_8031 ( ADD_371_U41 , U3217 , ADD_371_U24 );
nand NAND2_8032 ( ADD_371_U42 , ADD_371_U27 , ADD_371_U8 );
nand NAND2_8033 ( ADD_371_U43 , U3215 , ADD_371_U4 );
nand NAND2_8034 ( ADD_371_U44 , U3214 , ADD_371_U7 );
not NOT1_8035 ( ADD_405_U4 , INSTADDRPOINTER_REG_0_ );
nand NAND2_8036 ( ADD_405_U5 , ADD_405_U92 , ADD_405_U126 );
not NOT1_8037 ( ADD_405_U6 , INSTADDRPOINTER_REG_1_ );
not NOT1_8038 ( ADD_405_U7 , INSTADDRPOINTER_REG_3_ );
nand NAND2_8039 ( ADD_405_U8 , INSTADDRPOINTER_REG_3_ , ADD_405_U92 );
not NOT1_8040 ( ADD_405_U9 , INSTADDRPOINTER_REG_4_ );
nand NAND2_8041 ( ADD_405_U10 , INSTADDRPOINTER_REG_4_ , ADD_405_U98 );
not NOT1_8042 ( ADD_405_U11 , INSTADDRPOINTER_REG_5_ );
nand NAND2_8043 ( ADD_405_U12 , INSTADDRPOINTER_REG_5_ , ADD_405_U99 );
not NOT1_8044 ( ADD_405_U13 , INSTADDRPOINTER_REG_6_ );
nand NAND2_8045 ( ADD_405_U14 , INSTADDRPOINTER_REG_6_ , ADD_405_U100 );
not NOT1_8046 ( ADD_405_U15 , INSTADDRPOINTER_REG_7_ );
nand NAND2_8047 ( ADD_405_U16 , INSTADDRPOINTER_REG_7_ , ADD_405_U101 );
not NOT1_8048 ( ADD_405_U17 , INSTADDRPOINTER_REG_8_ );
not NOT1_8049 ( ADD_405_U18 , INSTADDRPOINTER_REG_9_ );
nand NAND2_8050 ( ADD_405_U19 , INSTADDRPOINTER_REG_8_ , ADD_405_U102 );
nand NAND2_8051 ( ADD_405_U20 , ADD_405_U103 , INSTADDRPOINTER_REG_9_ );
not NOT1_8052 ( ADD_405_U21 , INSTADDRPOINTER_REG_10_ );
nand NAND2_8053 ( ADD_405_U22 , INSTADDRPOINTER_REG_10_ , ADD_405_U104 );
not NOT1_8054 ( ADD_405_U23 , INSTADDRPOINTER_REG_11_ );
nand NAND2_8055 ( ADD_405_U24 , INSTADDRPOINTER_REG_11_ , ADD_405_U105 );
not NOT1_8056 ( ADD_405_U25 , INSTADDRPOINTER_REG_12_ );
nand NAND2_8057 ( ADD_405_U26 , INSTADDRPOINTER_REG_12_ , ADD_405_U106 );
not NOT1_8058 ( ADD_405_U27 , INSTADDRPOINTER_REG_13_ );
nand NAND2_8059 ( ADD_405_U28 , INSTADDRPOINTER_REG_13_ , ADD_405_U107 );
not NOT1_8060 ( ADD_405_U29 , INSTADDRPOINTER_REG_14_ );
nand NAND2_8061 ( ADD_405_U30 , INSTADDRPOINTER_REG_14_ , ADD_405_U108 );
not NOT1_8062 ( ADD_405_U31 , INSTADDRPOINTER_REG_15_ );
nand NAND2_8063 ( ADD_405_U32 , INSTADDRPOINTER_REG_15_ , ADD_405_U109 );
not NOT1_8064 ( ADD_405_U33 , INSTADDRPOINTER_REG_16_ );
nand NAND2_8065 ( ADD_405_U34 , INSTADDRPOINTER_REG_16_ , ADD_405_U110 );
not NOT1_8066 ( ADD_405_U35 , INSTADDRPOINTER_REG_17_ );
nand NAND2_8067 ( ADD_405_U36 , INSTADDRPOINTER_REG_17_ , ADD_405_U111 );
not NOT1_8068 ( ADD_405_U37 , INSTADDRPOINTER_REG_18_ );
nand NAND2_8069 ( ADD_405_U38 , INSTADDRPOINTER_REG_18_ , ADD_405_U112 );
not NOT1_8070 ( ADD_405_U39 , INSTADDRPOINTER_REG_19_ );
nand NAND2_8071 ( ADD_405_U40 , INSTADDRPOINTER_REG_19_ , ADD_405_U113 );
not NOT1_8072 ( ADD_405_U41 , INSTADDRPOINTER_REG_20_ );
nand NAND2_8073 ( ADD_405_U42 , INSTADDRPOINTER_REG_20_ , ADD_405_U114 );
not NOT1_8074 ( ADD_405_U43 , INSTADDRPOINTER_REG_21_ );
nand NAND2_8075 ( ADD_405_U44 , INSTADDRPOINTER_REG_21_ , ADD_405_U115 );
not NOT1_8076 ( ADD_405_U45 , INSTADDRPOINTER_REG_22_ );
nand NAND2_8077 ( ADD_405_U46 , INSTADDRPOINTER_REG_22_ , ADD_405_U116 );
not NOT1_8078 ( ADD_405_U47 , INSTADDRPOINTER_REG_23_ );
nand NAND2_8079 ( ADD_405_U48 , INSTADDRPOINTER_REG_23_ , ADD_405_U117 );
not NOT1_8080 ( ADD_405_U49 , INSTADDRPOINTER_REG_24_ );
nand NAND2_8081 ( ADD_405_U50 , INSTADDRPOINTER_REG_24_ , ADD_405_U118 );
not NOT1_8082 ( ADD_405_U51 , INSTADDRPOINTER_REG_25_ );
nand NAND2_8083 ( ADD_405_U52 , INSTADDRPOINTER_REG_25_ , ADD_405_U119 );
not NOT1_8084 ( ADD_405_U53 , INSTADDRPOINTER_REG_26_ );
nand NAND2_8085 ( ADD_405_U54 , INSTADDRPOINTER_REG_26_ , ADD_405_U120 );
not NOT1_8086 ( ADD_405_U55 , INSTADDRPOINTER_REG_27_ );
nand NAND2_8087 ( ADD_405_U56 , INSTADDRPOINTER_REG_27_ , ADD_405_U121 );
not NOT1_8088 ( ADD_405_U57 , INSTADDRPOINTER_REG_28_ );
nand NAND2_8089 ( ADD_405_U58 , INSTADDRPOINTER_REG_28_ , ADD_405_U122 );
not NOT1_8090 ( ADD_405_U59 , INSTADDRPOINTER_REG_29_ );
nand NAND2_8091 ( ADD_405_U60 , INSTADDRPOINTER_REG_29_ , ADD_405_U123 );
not NOT1_8092 ( ADD_405_U61 , INSTADDRPOINTER_REG_30_ );
not NOT1_8093 ( ADD_405_U62 , INSTADDRPOINTER_REG_2_ );
nand NAND2_8094 ( ADD_405_U63 , ADD_405_U128 , ADD_405_U127 );
nand NAND2_8095 ( ADD_405_U64 , ADD_405_U130 , ADD_405_U129 );
nand NAND2_8096 ( ADD_405_U65 , ADD_405_U132 , ADD_405_U131 );
nand NAND2_8097 ( ADD_405_U66 , ADD_405_U134 , ADD_405_U133 );
nand NAND2_8098 ( ADD_405_U67 , ADD_405_U136 , ADD_405_U135 );
nand NAND2_8099 ( ADD_405_U68 , ADD_405_U138 , ADD_405_U137 );
nand NAND2_8100 ( ADD_405_U69 , ADD_405_U142 , ADD_405_U141 );
nand NAND2_8101 ( ADD_405_U70 , ADD_405_U144 , ADD_405_U143 );
nand NAND2_8102 ( ADD_405_U71 , ADD_405_U146 , ADD_405_U145 );
nand NAND2_8103 ( ADD_405_U72 , ADD_405_U148 , ADD_405_U147 );
nand NAND2_8104 ( ADD_405_U73 , ADD_405_U150 , ADD_405_U149 );
nand NAND2_8105 ( ADD_405_U74 , ADD_405_U152 , ADD_405_U151 );
nand NAND2_8106 ( ADD_405_U75 , ADD_405_U154 , ADD_405_U153 );
nand NAND2_8107 ( ADD_405_U76 , ADD_405_U156 , ADD_405_U155 );
nand NAND2_8108 ( ADD_405_U77 , ADD_405_U158 , ADD_405_U157 );
nand NAND2_8109 ( ADD_405_U78 , ADD_405_U160 , ADD_405_U159 );
nand NAND2_8110 ( ADD_405_U79 , ADD_405_U162 , ADD_405_U161 );
nand NAND2_8111 ( ADD_405_U80 , ADD_405_U164 , ADD_405_U163 );
nand NAND2_8112 ( ADD_405_U81 , ADD_405_U166 , ADD_405_U165 );
nand NAND2_8113 ( ADD_405_U82 , ADD_405_U168 , ADD_405_U167 );
nand NAND2_8114 ( ADD_405_U83 , ADD_405_U170 , ADD_405_U169 );
nand NAND2_8115 ( ADD_405_U84 , ADD_405_U172 , ADD_405_U171 );
nand NAND2_8116 ( ADD_405_U85 , ADD_405_U174 , ADD_405_U173 );
nand NAND2_8117 ( ADD_405_U86 , ADD_405_U176 , ADD_405_U175 );
nand NAND2_8118 ( ADD_405_U87 , ADD_405_U178 , ADD_405_U177 );
nand NAND2_8119 ( ADD_405_U88 , ADD_405_U180 , ADD_405_U179 );
nand NAND2_8120 ( ADD_405_U89 , ADD_405_U182 , ADD_405_U181 );
nand NAND2_8121 ( ADD_405_U90 , ADD_405_U184 , ADD_405_U183 );
nand NAND2_8122 ( ADD_405_U91 , ADD_405_U186 , ADD_405_U185 );
nand NAND2_8123 ( ADD_405_U92 , ADD_405_U62 , ADD_405_U96 );
and AND2_8124 ( ADD_405_U93 , ADD_405_U140 , ADD_405_U139 );
not NOT1_8125 ( ADD_405_U94 , INSTADDRPOINTER_REG_31_ );
nand NAND2_8126 ( ADD_405_U95 , INSTADDRPOINTER_REG_30_ , ADD_405_U124 );
nand NAND2_8127 ( ADD_405_U96 , INSTADDRPOINTER_REG_1_ , INSTADDRPOINTER_REG_0_ );
not NOT1_8128 ( ADD_405_U97 , ADD_405_U92 );
not NOT1_8129 ( ADD_405_U98 , ADD_405_U8 );
not NOT1_8130 ( ADD_405_U99 , ADD_405_U10 );
not NOT1_8131 ( ADD_405_U100 , ADD_405_U12 );
not NOT1_8132 ( ADD_405_U101 , ADD_405_U14 );
not NOT1_8133 ( ADD_405_U102 , ADD_405_U16 );
not NOT1_8134 ( ADD_405_U103 , ADD_405_U19 );
not NOT1_8135 ( ADD_405_U104 , ADD_405_U20 );
not NOT1_8136 ( ADD_405_U105 , ADD_405_U22 );
not NOT1_8137 ( ADD_405_U106 , ADD_405_U24 );
not NOT1_8138 ( ADD_405_U107 , ADD_405_U26 );
not NOT1_8139 ( ADD_405_U108 , ADD_405_U28 );
not NOT1_8140 ( ADD_405_U109 , ADD_405_U30 );
not NOT1_8141 ( ADD_405_U110 , ADD_405_U32 );
not NOT1_8142 ( ADD_405_U111 , ADD_405_U34 );
not NOT1_8143 ( ADD_405_U112 , ADD_405_U36 );
not NOT1_8144 ( ADD_405_U113 , ADD_405_U38 );
not NOT1_8145 ( ADD_405_U114 , ADD_405_U40 );
not NOT1_8146 ( ADD_405_U115 , ADD_405_U42 );
not NOT1_8147 ( ADD_405_U116 , ADD_405_U44 );
not NOT1_8148 ( ADD_405_U117 , ADD_405_U46 );
not NOT1_8149 ( ADD_405_U118 , ADD_405_U48 );
not NOT1_8150 ( ADD_405_U119 , ADD_405_U50 );
not NOT1_8151 ( ADD_405_U120 , ADD_405_U52 );
not NOT1_8152 ( ADD_405_U121 , ADD_405_U54 );
not NOT1_8153 ( ADD_405_U122 , ADD_405_U56 );
not NOT1_8154 ( ADD_405_U123 , ADD_405_U58 );
not NOT1_8155 ( ADD_405_U124 , ADD_405_U60 );
not NOT1_8156 ( ADD_405_U125 , ADD_405_U95 );
nand NAND3_8157 ( ADD_405_U126 , INSTADDRPOINTER_REG_1_ , INSTADDRPOINTER_REG_0_ , INSTADDRPOINTER_REG_2_ );
nand NAND2_8158 ( ADD_405_U127 , INSTADDRPOINTER_REG_9_ , ADD_405_U19 );
nand NAND2_8159 ( ADD_405_U128 , ADD_405_U103 , ADD_405_U18 );
nand NAND2_8160 ( ADD_405_U129 , INSTADDRPOINTER_REG_8_ , ADD_405_U16 );
nand NAND2_8161 ( ADD_405_U130 , ADD_405_U102 , ADD_405_U17 );
nand NAND2_8162 ( ADD_405_U131 , INSTADDRPOINTER_REG_7_ , ADD_405_U14 );
nand NAND2_8163 ( ADD_405_U132 , ADD_405_U101 , ADD_405_U15 );
nand NAND2_8164 ( ADD_405_U133 , INSTADDRPOINTER_REG_6_ , ADD_405_U12 );
nand NAND2_8165 ( ADD_405_U134 , ADD_405_U100 , ADD_405_U13 );
nand NAND2_8166 ( ADD_405_U135 , INSTADDRPOINTER_REG_5_ , ADD_405_U10 );
nand NAND2_8167 ( ADD_405_U136 , ADD_405_U99 , ADD_405_U11 );
nand NAND2_8168 ( ADD_405_U137 , INSTADDRPOINTER_REG_4_ , ADD_405_U8 );
nand NAND2_8169 ( ADD_405_U138 , ADD_405_U98 , ADD_405_U9 );
nand NAND2_8170 ( ADD_405_U139 , INSTADDRPOINTER_REG_3_ , ADD_405_U92 );
nand NAND2_8171 ( ADD_405_U140 , ADD_405_U97 , ADD_405_U7 );
nand NAND2_8172 ( ADD_405_U141 , INSTADDRPOINTER_REG_31_ , ADD_405_U95 );
nand NAND2_8173 ( ADD_405_U142 , ADD_405_U125 , ADD_405_U94 );
nand NAND2_8174 ( ADD_405_U143 , INSTADDRPOINTER_REG_30_ , ADD_405_U60 );
nand NAND2_8175 ( ADD_405_U144 , ADD_405_U124 , ADD_405_U61 );
nand NAND2_8176 ( ADD_405_U145 , INSTADDRPOINTER_REG_29_ , ADD_405_U58 );
nand NAND2_8177 ( ADD_405_U146 , ADD_405_U123 , ADD_405_U59 );
nand NAND2_8178 ( ADD_405_U147 , INSTADDRPOINTER_REG_28_ , ADD_405_U56 );
nand NAND2_8179 ( ADD_405_U148 , ADD_405_U122 , ADD_405_U57 );
nand NAND2_8180 ( ADD_405_U149 , INSTADDRPOINTER_REG_27_ , ADD_405_U54 );
nand NAND2_8181 ( ADD_405_U150 , ADD_405_U121 , ADD_405_U55 );
nand NAND2_8182 ( ADD_405_U151 , INSTADDRPOINTER_REG_26_ , ADD_405_U52 );
nand NAND2_8183 ( ADD_405_U152 , ADD_405_U120 , ADD_405_U53 );
nand NAND2_8184 ( ADD_405_U153 , INSTADDRPOINTER_REG_25_ , ADD_405_U50 );
nand NAND2_8185 ( ADD_405_U154 , ADD_405_U119 , ADD_405_U51 );
nand NAND2_8186 ( ADD_405_U155 , INSTADDRPOINTER_REG_24_ , ADD_405_U48 );
nand NAND2_8187 ( ADD_405_U156 , ADD_405_U118 , ADD_405_U49 );
nand NAND2_8188 ( ADD_405_U157 , INSTADDRPOINTER_REG_23_ , ADD_405_U46 );
nand NAND2_8189 ( ADD_405_U158 , ADD_405_U117 , ADD_405_U47 );
nand NAND2_8190 ( ADD_405_U159 , INSTADDRPOINTER_REG_22_ , ADD_405_U44 );
nand NAND2_8191 ( ADD_405_U160 , ADD_405_U116 , ADD_405_U45 );
nand NAND2_8192 ( ADD_405_U161 , INSTADDRPOINTER_REG_21_ , ADD_405_U42 );
nand NAND2_8193 ( ADD_405_U162 , ADD_405_U115 , ADD_405_U43 );
nand NAND2_8194 ( ADD_405_U163 , INSTADDRPOINTER_REG_20_ , ADD_405_U40 );
nand NAND2_8195 ( ADD_405_U164 , ADD_405_U114 , ADD_405_U41 );
nand NAND2_8196 ( ADD_405_U165 , INSTADDRPOINTER_REG_1_ , ADD_405_U4 );
nand NAND2_8197 ( ADD_405_U166 , INSTADDRPOINTER_REG_0_ , ADD_405_U6 );
nand NAND2_8198 ( ADD_405_U167 , INSTADDRPOINTER_REG_19_ , ADD_405_U38 );
nand NAND2_8199 ( ADD_405_U168 , ADD_405_U113 , ADD_405_U39 );
nand NAND2_8200 ( ADD_405_U169 , INSTADDRPOINTER_REG_18_ , ADD_405_U36 );
nand NAND2_8201 ( ADD_405_U170 , ADD_405_U112 , ADD_405_U37 );
nand NAND2_8202 ( ADD_405_U171 , INSTADDRPOINTER_REG_17_ , ADD_405_U34 );
nand NAND2_8203 ( ADD_405_U172 , ADD_405_U111 , ADD_405_U35 );
nand NAND2_8204 ( ADD_405_U173 , INSTADDRPOINTER_REG_16_ , ADD_405_U32 );
nand NAND2_8205 ( ADD_405_U174 , ADD_405_U110 , ADD_405_U33 );
nand NAND2_8206 ( ADD_405_U175 , INSTADDRPOINTER_REG_15_ , ADD_405_U30 );
nand NAND2_8207 ( ADD_405_U176 , ADD_405_U109 , ADD_405_U31 );
nand NAND2_8208 ( ADD_405_U177 , INSTADDRPOINTER_REG_14_ , ADD_405_U28 );
nand NAND2_8209 ( ADD_405_U178 , ADD_405_U108 , ADD_405_U29 );
nand NAND2_8210 ( ADD_405_U179 , INSTADDRPOINTER_REG_13_ , ADD_405_U26 );
nand NAND2_8211 ( ADD_405_U180 , ADD_405_U107 , ADD_405_U27 );
nand NAND2_8212 ( ADD_405_U181 , INSTADDRPOINTER_REG_12_ , ADD_405_U24 );
nand NAND2_8213 ( ADD_405_U182 , ADD_405_U106 , ADD_405_U25 );
nand NAND2_8214 ( ADD_405_U183 , INSTADDRPOINTER_REG_11_ , ADD_405_U22 );
nand NAND2_8215 ( ADD_405_U184 , ADD_405_U105 , ADD_405_U23 );
nand NAND2_8216 ( ADD_405_U185 , INSTADDRPOINTER_REG_10_ , ADD_405_U20 );
nand NAND2_8217 ( ADD_405_U186 , ADD_405_U104 , ADD_405_U21 );
nor nor_8218 ( GTE_485_U6 , R2238_U6 , GTE_485_U7 );
nor nor_8219 ( GTE_485_U7 , R2238_U19 , R2238_U20 , R2238_U22 , R2238_U21 );
not NOT1_8220 ( ADD_515_U4 , INSTADDRPOINTER_REG_1_ );
not NOT1_8221 ( ADD_515_U5 , INSTADDRPOINTER_REG_2_ );
nand NAND2_8222 ( ADD_515_U6 , INSTADDRPOINTER_REG_2_ , INSTADDRPOINTER_REG_1_ );
not NOT1_8223 ( ADD_515_U7 , INSTADDRPOINTER_REG_3_ );
nand NAND2_8224 ( ADD_515_U8 , INSTADDRPOINTER_REG_3_ , ADD_515_U94 );
not NOT1_8225 ( ADD_515_U9 , INSTADDRPOINTER_REG_4_ );
nand NAND2_8226 ( ADD_515_U10 , INSTADDRPOINTER_REG_4_ , ADD_515_U95 );
not NOT1_8227 ( ADD_515_U11 , INSTADDRPOINTER_REG_5_ );
nand NAND2_8228 ( ADD_515_U12 , INSTADDRPOINTER_REG_5_ , ADD_515_U96 );
not NOT1_8229 ( ADD_515_U13 , INSTADDRPOINTER_REG_6_ );
nand NAND2_8230 ( ADD_515_U14 , INSTADDRPOINTER_REG_6_ , ADD_515_U97 );
not NOT1_8231 ( ADD_515_U15 , INSTADDRPOINTER_REG_7_ );
nand NAND2_8232 ( ADD_515_U16 , INSTADDRPOINTER_REG_7_ , ADD_515_U98 );
not NOT1_8233 ( ADD_515_U17 , INSTADDRPOINTER_REG_8_ );
not NOT1_8234 ( ADD_515_U18 , INSTADDRPOINTER_REG_9_ );
nand NAND2_8235 ( ADD_515_U19 , INSTADDRPOINTER_REG_8_ , ADD_515_U99 );
nand NAND2_8236 ( ADD_515_U20 , ADD_515_U100 , INSTADDRPOINTER_REG_9_ );
not NOT1_8237 ( ADD_515_U21 , INSTADDRPOINTER_REG_10_ );
nand NAND2_8238 ( ADD_515_U22 , INSTADDRPOINTER_REG_10_ , ADD_515_U101 );
not NOT1_8239 ( ADD_515_U23 , INSTADDRPOINTER_REG_11_ );
nand NAND2_8240 ( ADD_515_U24 , INSTADDRPOINTER_REG_11_ , ADD_515_U102 );
not NOT1_8241 ( ADD_515_U25 , INSTADDRPOINTER_REG_12_ );
nand NAND2_8242 ( ADD_515_U26 , INSTADDRPOINTER_REG_12_ , ADD_515_U103 );
not NOT1_8243 ( ADD_515_U27 , INSTADDRPOINTER_REG_13_ );
nand NAND2_8244 ( ADD_515_U28 , INSTADDRPOINTER_REG_13_ , ADD_515_U104 );
not NOT1_8245 ( ADD_515_U29 , INSTADDRPOINTER_REG_14_ );
nand NAND2_8246 ( ADD_515_U30 , INSTADDRPOINTER_REG_14_ , ADD_515_U105 );
not NOT1_8247 ( ADD_515_U31 , INSTADDRPOINTER_REG_15_ );
nand NAND2_8248 ( ADD_515_U32 , INSTADDRPOINTER_REG_15_ , ADD_515_U106 );
not NOT1_8249 ( ADD_515_U33 , INSTADDRPOINTER_REG_16_ );
nand NAND2_8250 ( ADD_515_U34 , INSTADDRPOINTER_REG_16_ , ADD_515_U107 );
not NOT1_8251 ( ADD_515_U35 , INSTADDRPOINTER_REG_17_ );
nand NAND2_8252 ( ADD_515_U36 , INSTADDRPOINTER_REG_17_ , ADD_515_U108 );
not NOT1_8253 ( ADD_515_U37 , INSTADDRPOINTER_REG_18_ );
nand NAND2_8254 ( ADD_515_U38 , INSTADDRPOINTER_REG_18_ , ADD_515_U109 );
not NOT1_8255 ( ADD_515_U39 , INSTADDRPOINTER_REG_19_ );
nand NAND2_8256 ( ADD_515_U40 , INSTADDRPOINTER_REG_19_ , ADD_515_U110 );
not NOT1_8257 ( ADD_515_U41 , INSTADDRPOINTER_REG_20_ );
nand NAND2_8258 ( ADD_515_U42 , INSTADDRPOINTER_REG_20_ , ADD_515_U111 );
not NOT1_8259 ( ADD_515_U43 , INSTADDRPOINTER_REG_21_ );
nand NAND2_8260 ( ADD_515_U44 , INSTADDRPOINTER_REG_21_ , ADD_515_U112 );
not NOT1_8261 ( ADD_515_U45 , INSTADDRPOINTER_REG_22_ );
nand NAND2_8262 ( ADD_515_U46 , INSTADDRPOINTER_REG_22_ , ADD_515_U113 );
not NOT1_8263 ( ADD_515_U47 , INSTADDRPOINTER_REG_23_ );
nand NAND2_8264 ( ADD_515_U48 , INSTADDRPOINTER_REG_23_ , ADD_515_U114 );
not NOT1_8265 ( ADD_515_U49 , INSTADDRPOINTER_REG_24_ );
nand NAND2_8266 ( ADD_515_U50 , INSTADDRPOINTER_REG_24_ , ADD_515_U115 );
not NOT1_8267 ( ADD_515_U51 , INSTADDRPOINTER_REG_25_ );
nand NAND2_8268 ( ADD_515_U52 , INSTADDRPOINTER_REG_25_ , ADD_515_U116 );
not NOT1_8269 ( ADD_515_U53 , INSTADDRPOINTER_REG_26_ );
nand NAND2_8270 ( ADD_515_U54 , INSTADDRPOINTER_REG_26_ , ADD_515_U117 );
not NOT1_8271 ( ADD_515_U55 , INSTADDRPOINTER_REG_27_ );
nand NAND2_8272 ( ADD_515_U56 , INSTADDRPOINTER_REG_27_ , ADD_515_U118 );
not NOT1_8273 ( ADD_515_U57 , INSTADDRPOINTER_REG_28_ );
nand NAND2_8274 ( ADD_515_U58 , INSTADDRPOINTER_REG_28_ , ADD_515_U119 );
not NOT1_8275 ( ADD_515_U59 , INSTADDRPOINTER_REG_29_ );
nand NAND2_8276 ( ADD_515_U60 , INSTADDRPOINTER_REG_29_ , ADD_515_U120 );
not NOT1_8277 ( ADD_515_U61 , INSTADDRPOINTER_REG_30_ );
nand NAND2_8278 ( ADD_515_U62 , ADD_515_U124 , ADD_515_U123 );
nand NAND2_8279 ( ADD_515_U63 , ADD_515_U126 , ADD_515_U125 );
nand NAND2_8280 ( ADD_515_U64 , ADD_515_U128 , ADD_515_U127 );
nand NAND2_8281 ( ADD_515_U65 , ADD_515_U130 , ADD_515_U129 );
nand NAND2_8282 ( ADD_515_U66 , ADD_515_U132 , ADD_515_U131 );
nand NAND2_8283 ( ADD_515_U67 , ADD_515_U134 , ADD_515_U133 );
nand NAND2_8284 ( ADD_515_U68 , ADD_515_U136 , ADD_515_U135 );
nand NAND2_8285 ( ADD_515_U69 , ADD_515_U138 , ADD_515_U137 );
nand NAND2_8286 ( ADD_515_U70 , ADD_515_U140 , ADD_515_U139 );
nand NAND2_8287 ( ADD_515_U71 , ADD_515_U142 , ADD_515_U141 );
nand NAND2_8288 ( ADD_515_U72 , ADD_515_U144 , ADD_515_U143 );
nand NAND2_8289 ( ADD_515_U73 , ADD_515_U146 , ADD_515_U145 );
nand NAND2_8290 ( ADD_515_U74 , ADD_515_U148 , ADD_515_U147 );
nand NAND2_8291 ( ADD_515_U75 , ADD_515_U150 , ADD_515_U149 );
nand NAND2_8292 ( ADD_515_U76 , ADD_515_U152 , ADD_515_U151 );
nand NAND2_8293 ( ADD_515_U77 , ADD_515_U154 , ADD_515_U153 );
nand NAND2_8294 ( ADD_515_U78 , ADD_515_U156 , ADD_515_U155 );
nand NAND2_8295 ( ADD_515_U79 , ADD_515_U158 , ADD_515_U157 );
nand NAND2_8296 ( ADD_515_U80 , ADD_515_U160 , ADD_515_U159 );
nand NAND2_8297 ( ADD_515_U81 , ADD_515_U162 , ADD_515_U161 );
nand NAND2_8298 ( ADD_515_U82 , ADD_515_U164 , ADD_515_U163 );
nand NAND2_8299 ( ADD_515_U83 , ADD_515_U166 , ADD_515_U165 );
nand NAND2_8300 ( ADD_515_U84 , ADD_515_U168 , ADD_515_U167 );
nand NAND2_8301 ( ADD_515_U85 , ADD_515_U170 , ADD_515_U169 );
nand NAND2_8302 ( ADD_515_U86 , ADD_515_U172 , ADD_515_U171 );
nand NAND2_8303 ( ADD_515_U87 , ADD_515_U174 , ADD_515_U173 );
nand NAND2_8304 ( ADD_515_U88 , ADD_515_U176 , ADD_515_U175 );
nand NAND2_8305 ( ADD_515_U89 , ADD_515_U178 , ADD_515_U177 );
nand NAND2_8306 ( ADD_515_U90 , ADD_515_U180 , ADD_515_U179 );
nand NAND2_8307 ( ADD_515_U91 , ADD_515_U182 , ADD_515_U181 );
not NOT1_8308 ( ADD_515_U92 , INSTADDRPOINTER_REG_31_ );
nand NAND2_8309 ( ADD_515_U93 , INSTADDRPOINTER_REG_30_ , ADD_515_U121 );
not NOT1_8310 ( ADD_515_U94 , ADD_515_U6 );
not NOT1_8311 ( ADD_515_U95 , ADD_515_U8 );
not NOT1_8312 ( ADD_515_U96 , ADD_515_U10 );
not NOT1_8313 ( ADD_515_U97 , ADD_515_U12 );
not NOT1_8314 ( ADD_515_U98 , ADD_515_U14 );
not NOT1_8315 ( ADD_515_U99 , ADD_515_U16 );
not NOT1_8316 ( ADD_515_U100 , ADD_515_U19 );
not NOT1_8317 ( ADD_515_U101 , ADD_515_U20 );
not NOT1_8318 ( ADD_515_U102 , ADD_515_U22 );
not NOT1_8319 ( ADD_515_U103 , ADD_515_U24 );
not NOT1_8320 ( ADD_515_U104 , ADD_515_U26 );
not NOT1_8321 ( ADD_515_U105 , ADD_515_U28 );
not NOT1_8322 ( ADD_515_U106 , ADD_515_U30 );
not NOT1_8323 ( ADD_515_U107 , ADD_515_U32 );
not NOT1_8324 ( ADD_515_U108 , ADD_515_U34 );
not NOT1_8325 ( ADD_515_U109 , ADD_515_U36 );
not NOT1_8326 ( ADD_515_U110 , ADD_515_U38 );
not NOT1_8327 ( ADD_515_U111 , ADD_515_U40 );
not NOT1_8328 ( ADD_515_U112 , ADD_515_U42 );
not NOT1_8329 ( ADD_515_U113 , ADD_515_U44 );
not NOT1_8330 ( ADD_515_U114 , ADD_515_U46 );
not NOT1_8331 ( ADD_515_U115 , ADD_515_U48 );
not NOT1_8332 ( ADD_515_U116 , ADD_515_U50 );
not NOT1_8333 ( ADD_515_U117 , ADD_515_U52 );
not NOT1_8334 ( ADD_515_U118 , ADD_515_U54 );
not NOT1_8335 ( ADD_515_U119 , ADD_515_U56 );
not NOT1_8336 ( ADD_515_U120 , ADD_515_U58 );
not NOT1_8337 ( ADD_515_U121 , ADD_515_U60 );
not NOT1_8338 ( ADD_515_U122 , ADD_515_U93 );
nand NAND2_8339 ( ADD_515_U123 , INSTADDRPOINTER_REG_9_ , ADD_515_U19 );
nand NAND2_8340 ( ADD_515_U124 , ADD_515_U100 , ADD_515_U18 );
nand NAND2_8341 ( ADD_515_U125 , INSTADDRPOINTER_REG_8_ , ADD_515_U16 );
nand NAND2_8342 ( ADD_515_U126 , ADD_515_U99 , ADD_515_U17 );
nand NAND2_8343 ( ADD_515_U127 , INSTADDRPOINTER_REG_7_ , ADD_515_U14 );
nand NAND2_8344 ( ADD_515_U128 , ADD_515_U98 , ADD_515_U15 );
nand NAND2_8345 ( ADD_515_U129 , INSTADDRPOINTER_REG_6_ , ADD_515_U12 );
nand NAND2_8346 ( ADD_515_U130 , ADD_515_U97 , ADD_515_U13 );
nand NAND2_8347 ( ADD_515_U131 , INSTADDRPOINTER_REG_5_ , ADD_515_U10 );
nand NAND2_8348 ( ADD_515_U132 , ADD_515_U96 , ADD_515_U11 );
nand NAND2_8349 ( ADD_515_U133 , INSTADDRPOINTER_REG_4_ , ADD_515_U8 );
nand NAND2_8350 ( ADD_515_U134 , ADD_515_U95 , ADD_515_U9 );
nand NAND2_8351 ( ADD_515_U135 , INSTADDRPOINTER_REG_3_ , ADD_515_U6 );
nand NAND2_8352 ( ADD_515_U136 , ADD_515_U94 , ADD_515_U7 );
nand NAND2_8353 ( ADD_515_U137 , INSTADDRPOINTER_REG_31_ , ADD_515_U93 );
nand NAND2_8354 ( ADD_515_U138 , ADD_515_U122 , ADD_515_U92 );
nand NAND2_8355 ( ADD_515_U139 , INSTADDRPOINTER_REG_30_ , ADD_515_U60 );
nand NAND2_8356 ( ADD_515_U140 , ADD_515_U121 , ADD_515_U61 );
nand NAND2_8357 ( ADD_515_U141 , INSTADDRPOINTER_REG_2_ , ADD_515_U4 );
nand NAND2_8358 ( ADD_515_U142 , INSTADDRPOINTER_REG_1_ , ADD_515_U5 );
nand NAND2_8359 ( ADD_515_U143 , INSTADDRPOINTER_REG_29_ , ADD_515_U58 );
nand NAND2_8360 ( ADD_515_U144 , ADD_515_U120 , ADD_515_U59 );
nand NAND2_8361 ( ADD_515_U145 , INSTADDRPOINTER_REG_28_ , ADD_515_U56 );
nand NAND2_8362 ( ADD_515_U146 , ADD_515_U119 , ADD_515_U57 );
nand NAND2_8363 ( ADD_515_U147 , INSTADDRPOINTER_REG_27_ , ADD_515_U54 );
nand NAND2_8364 ( ADD_515_U148 , ADD_515_U118 , ADD_515_U55 );
nand NAND2_8365 ( ADD_515_U149 , INSTADDRPOINTER_REG_26_ , ADD_515_U52 );
nand NAND2_8366 ( ADD_515_U150 , ADD_515_U117 , ADD_515_U53 );
nand NAND2_8367 ( ADD_515_U151 , INSTADDRPOINTER_REG_25_ , ADD_515_U50 );

// 70 Additional buffers.
buf add_BUF1_1 ( BE_N_REG_3_ , BE_N_REG_3__EXTRA );
buf add_BUF1_2 ( BE_N_REG_2_ , BE_N_REG_2__EXTRA );
buf add_BUF1_3 ( BE_N_REG_1_ , BE_N_REG_1__EXTRA );
buf add_BUF1_4 ( BE_N_REG_0_ , BE_N_REG_0__EXTRA );
buf add_BUF1_5 ( ADDRESS_REG_29_ , ADDRESS_REG_29__EXTRA );
buf add_BUF1_6 ( ADDRESS_REG_28_ , ADDRESS_REG_28__EXTRA );
buf add_BUF1_7 ( ADDRESS_REG_27_ , ADDRESS_REG_27__EXTRA );
buf add_BUF1_8 ( ADDRESS_REG_26_ , ADDRESS_REG_26__EXTRA );
buf add_BUF1_9 ( ADDRESS_REG_25_ , ADDRESS_REG_25__EXTRA );
buf add_BUF1_10 ( ADDRESS_REG_24_ , ADDRESS_REG_24__EXTRA );
buf add_BUF1_11 ( ADDRESS_REG_23_ , ADDRESS_REG_23__EXTRA );
buf add_BUF1_12 ( ADDRESS_REG_22_ , ADDRESS_REG_22__EXTRA );
buf add_BUF1_13 ( ADDRESS_REG_21_ , ADDRESS_REG_21__EXTRA );
buf add_BUF1_14 ( ADDRESS_REG_20_ , ADDRESS_REG_20__EXTRA );
buf add_BUF1_15 ( ADDRESS_REG_19_ , ADDRESS_REG_19__EXTRA );
buf add_BUF1_16 ( ADDRESS_REG_18_ , ADDRESS_REG_18__EXTRA );
buf add_BUF1_17 ( ADDRESS_REG_17_ , ADDRESS_REG_17__EXTRA );
buf add_BUF1_18 ( ADDRESS_REG_16_ , ADDRESS_REG_16__EXTRA );
buf add_BUF1_19 ( ADDRESS_REG_15_ , ADDRESS_REG_15__EXTRA );
buf add_BUF1_20 ( ADDRESS_REG_14_ , ADDRESS_REG_14__EXTRA );
buf add_BUF1_21 ( ADDRESS_REG_13_ , ADDRESS_REG_13__EXTRA );
buf add_BUF1_22 ( ADDRESS_REG_12_ , ADDRESS_REG_12__EXTRA );
buf add_BUF1_23 ( ADDRESS_REG_11_ , ADDRESS_REG_11__EXTRA );
buf add_BUF1_24 ( ADDRESS_REG_10_ , ADDRESS_REG_10__EXTRA );
buf add_BUF1_25 ( ADDRESS_REG_9_ , ADDRESS_REG_9__EXTRA );
buf add_BUF1_26 ( ADDRESS_REG_8_ , ADDRESS_REG_8__EXTRA );
buf add_BUF1_27 ( ADDRESS_REG_7_ , ADDRESS_REG_7__EXTRA );
buf add_BUF1_28 ( ADDRESS_REG_6_ , ADDRESS_REG_6__EXTRA );
buf add_BUF1_29 ( ADDRESS_REG_5_ , ADDRESS_REG_5__EXTRA );
buf add_BUF1_30 ( ADDRESS_REG_4_ , ADDRESS_REG_4__EXTRA );
buf add_BUF1_31 ( ADDRESS_REG_3_ , ADDRESS_REG_3__EXTRA );
buf add_BUF1_32 ( ADDRESS_REG_2_ , ADDRESS_REG_2__EXTRA );
buf add_BUF1_33 ( ADDRESS_REG_1_ , ADDRESS_REG_1__EXTRA );
buf add_BUF1_34 ( ADDRESS_REG_0_ , ADDRESS_REG_0__EXTRA );
buf add_BUF1_35 ( DATAO_REG_0_ , DATAO_REG_0__EXTRA );
buf add_BUF1_36 ( DATAO_REG_1_ , DATAO_REG_1__EXTRA );
buf add_BUF1_37 ( DATAO_REG_2_ , DATAO_REG_2__EXTRA );
buf add_BUF1_38 ( DATAO_REG_3_ , DATAO_REG_3__EXTRA );
buf add_BUF1_39 ( DATAO_REG_4_ , DATAO_REG_4__EXTRA );
buf add_BUF1_40 ( DATAO_REG_5_ , DATAO_REG_5__EXTRA );
buf add_BUF1_41 ( DATAO_REG_6_ , DATAO_REG_6__EXTRA );
buf add_BUF1_42 ( DATAO_REG_7_ , DATAO_REG_7__EXTRA );
buf add_BUF1_43 ( DATAO_REG_8_ , DATAO_REG_8__EXTRA );
buf add_BUF1_44 ( DATAO_REG_9_ , DATAO_REG_9__EXTRA );
buf add_BUF1_45 ( DATAO_REG_10_ , DATAO_REG_10__EXTRA );
buf add_BUF1_46 ( DATAO_REG_11_ , DATAO_REG_11__EXTRA );
buf add_BUF1_47 ( DATAO_REG_12_ , DATAO_REG_12__EXTRA );
buf add_BUF1_48 ( DATAO_REG_13_ , DATAO_REG_13__EXTRA );
buf add_BUF1_49 ( DATAO_REG_14_ , DATAO_REG_14__EXTRA );
buf add_BUF1_50 ( DATAO_REG_15_ , DATAO_REG_15__EXTRA );
buf add_BUF1_51 ( DATAO_REG_16_ , DATAO_REG_16__EXTRA );
buf add_BUF1_52 ( DATAO_REG_17_ , DATAO_REG_17__EXTRA );
buf add_BUF1_53 ( DATAO_REG_18_ , DATAO_REG_18__EXTRA );
buf add_BUF1_54 ( DATAO_REG_19_ , DATAO_REG_19__EXTRA );
buf add_BUF1_55 ( DATAO_REG_20_ , DATAO_REG_20__EXTRA );
buf add_BUF1_56 ( DATAO_REG_21_ , DATAO_REG_21__EXTRA );
buf add_BUF1_57 ( DATAO_REG_22_ , DATAO_REG_22__EXTRA );
buf add_BUF1_58 ( DATAO_REG_23_ , DATAO_REG_23__EXTRA );
buf add_BUF1_59 ( DATAO_REG_24_ , DATAO_REG_24__EXTRA );
buf add_BUF1_60 ( DATAO_REG_25_ , DATAO_REG_25__EXTRA );
buf add_BUF1_61 ( DATAO_REG_26_ , DATAO_REG_26__EXTRA );
buf add_BUF1_62 ( DATAO_REG_27_ , DATAO_REG_27__EXTRA );
buf add_BUF1_63 ( DATAO_REG_28_ , DATAO_REG_28__EXTRA );
buf add_BUF1_64 ( DATAO_REG_29_ , DATAO_REG_29__EXTRA );
buf add_BUF1_65 ( DATAO_REG_30_ , DATAO_REG_30__EXTRA );
buf add_BUF1_66 ( DATAO_REG_31_ , DATAO_REG_31__EXTRA );
buf add_BUF1_67 ( W_R_N_REG , W_R_N_REG_EXTRA );
buf add_BUF1_68 ( D_C_N_REG , D_C_N_REG_EXTRA );
buf add_BUF1_69 ( M_IO_N_REG , M_IO_N_REG_EXTRA );
buf add_BUF1_70 ( ADS_N_REG , ADS_N_REG_EXTRA );

endmodule
