// b17
// 1452 inputs  (37 PIs + 1415 PPIs)
// 1512 outputs (97 POs + 1415 PPOs)
// 30844 gates (26303 gates + 4474 inverters + 67 buffers )
// ( 4054 AND + 299 OR + 21815 NAND + 135 NOR + 67 BUFF )
// Time: Wed Mar 25 17:47:48 2009
// All copyrigh from NCKU EE TestLAB, Taiwan. [2008.12. WCL]

module b17_ras ( U247 , U246 , U245 , U244 , U243 , U242 ,
             U241 , U240 , U239 , U238 , U237 , U236 ,
             U235 , U234 , U233 , U232 , U231 , U230 ,
             U229 , U228 , U227 , U226 , U225 , U224 ,
             U223 , U222 , U221 , U220 , U219 , U218 ,
             U217 , U216 , U251 , U252 , U253 , U254 ,
             U255 , U256 , U257 , U258 , U259 , U260 ,
             U261 , U262 , U263 , U264 , U265 , U266 ,
             U267 , U268 , U269 , U270 , U271 , U272 ,
             U273 , U274 , U275 , U276 , U277 , U278 ,
             U279 , U280 , U281 , U282 , U212 , U215 ,
             U213 , U214 , P3_U3274 , P3_U3275 , P3_U3276 , P3_U3277 ,
             P3_U3061 , P3_U3060 , P3_U3059 , P3_U3058 , P3_U3057 , P3_U3056 ,
             P3_U3055 , P3_U3054 , P3_U3053 , P3_U3052 , P3_U3051 , P3_U3050 ,
             P3_U3049 , P3_U3048 , P3_U3047 , P3_U3046 , P3_U3045 , P3_U3044 ,
             P3_U3043 , P3_U3042 , P3_U3041 , P3_U3040 , P3_U3039 , P3_U3038 ,
             P3_U3037 , P3_U3036 , P3_U3035 , P3_U3034 , P3_U3033 , P3_U3032 ,
             P3_U3031 , P3_U3030 , P3_U3029 , P3_U3280 , P3_U3281 , P3_U3028 ,
             P3_U3027 , P3_U3026 , P3_U3025 , P3_U3024 , P3_U3023 , P3_U3022 ,
             P3_U3021 , P3_U3020 , P3_U3019 , P3_U3018 , P3_U3017 , P3_U3016 ,
             P3_U3015 , P3_U3014 , P3_U3013 , P3_U3012 , P3_U3011 , P3_U3010 ,
             P3_U3009 , P3_U3008 , P3_U3007 , P3_U3006 , P3_U3005 , P3_U3004 ,
             P3_U3003 , P3_U3002 , P3_U3001 , P3_U3000 , P3_U2999 , P3_U3282 ,
             P3_U2998 , P3_U2997 , P3_U2996 , P3_U2995 , P3_U2994 , P3_U2993 ,
             P3_U2992 , P3_U2991 , P3_U2990 , P3_U2989 , P3_U2988 , P3_U2987 ,
             P3_U2986 , P3_U2985 , P3_U2984 , P3_U2983 , P3_U2982 , P3_U2981 ,
             P3_U2980 , P3_U2979 , P3_U2978 , P3_U2977 , P3_U2976 , P3_U2975 ,
             P3_U2974 , P3_U2973 , P3_U2972 , P3_U2971 , P3_U2970 , P3_U2969 ,
             P3_U2968 , P3_U2967 , P3_U2966 , P3_U2965 , P3_U2964 , P3_U2963 ,
             P3_U2962 , P3_U2961 , P3_U2960 , P3_U2959 , P3_U2958 , P3_U2957 ,
             P3_U2956 , P3_U2955 , P3_U2954 , P3_U2953 , P3_U2952 , P3_U2951 ,
             P3_U2950 , P3_U2949 , P3_U2948 , P3_U2947 , P3_U2946 , P3_U2945 ,
             P3_U2944 , P3_U2943 , P3_U2942 , P3_U2941 , P3_U2940 , P3_U2939 ,
             P3_U2938 , P3_U2937 , P3_U2936 , P3_U2935 , P3_U2934 , P3_U2933 ,
             P3_U2932 , P3_U2931 , P3_U2930 , P3_U2929 , P3_U2928 , P3_U2927 ,
             P3_U2926 , P3_U2925 , P3_U2924 , P3_U2923 , P3_U2922 , P3_U2921 ,
             P3_U2920 , P3_U2919 , P3_U2918 , P3_U2917 , P3_U2916 , P3_U2915 ,
             P3_U2914 , P3_U2913 , P3_U2912 , P3_U2911 , P3_U2910 , P3_U2909 ,
             P3_U2908 , P3_U2907 , P3_U2906 , P3_U2905 , P3_U2904 , P3_U2903 ,
             P3_U2902 , P3_U2901 , P3_U2900 , P3_U2899 , P3_U2898 , P3_U2897 ,
             P3_U2896 , P3_U2895 , P3_U2894 , P3_U2893 , P3_U2892 , P3_U2891 ,
             P3_U2890 , P3_U2889 , P3_U2888 , P3_U2887 , P3_U2886 , P3_U2885 ,
             P3_U2884 , P3_U2883 , P3_U2882 , P3_U2881 , P3_U2880 , P3_U2879 ,
             P3_U2878 , P3_U2877 , P3_U2876 , P3_U2875 , P3_U2874 , P3_U2873 ,
             P3_U2872 , P3_U2871 , P3_U2870 , P3_U2869 , P3_U2868 , P3_U3284 ,
             P3_U3285 , P3_U3288 , P3_U3289 , P3_U3290 , P3_U2867 , P3_U2866 ,
             P3_U2865 , P3_U2864 , P3_U2863 , P3_U2862 , P3_U2861 , P3_U2860 ,
             P3_U2859 , P3_U2858 , P3_U2857 , P3_U2856 , P3_U2855 , P3_U2854 ,
             P3_U2853 , P3_U2852 , P3_U2851 , P3_U2850 , P3_U2849 , P3_U2848 ,
             P3_U2847 , P3_U2846 , P3_U2845 , P3_U2844 , P3_U2843 , P3_U2842 ,
             P3_U2841 , P3_U2840 , P3_U2839 , P3_U2838 , P3_U2837 , P3_U2836 ,
             P3_U2835 , P3_U2834 , P3_U2833 , P3_U2832 , P3_U2831 , P3_U2830 ,
             P3_U2829 , P3_U2828 , P3_U2827 , P3_U2826 , P3_U2825 , P3_U2824 ,
             P3_U2823 , P3_U2822 , P3_U2821 , P3_U2820 , P3_U2819 , P3_U2818 ,
             P3_U2817 , P3_U2816 , P3_U2815 , P3_U2814 , P3_U2813 , P3_U2812 ,
             P3_U2811 , P3_U2810 , P3_U2809 , P3_U2808 , P3_U2807 , P3_U2806 ,
             P3_U2805 , P3_U2804 , P3_U2803 , P3_U2802 , P3_U2801 , P3_U2800 ,
             P3_U2799 , P3_U2798 , P3_U2797 , P3_U2796 , P3_U2795 , P3_U2794 ,
             P3_U2793 , P3_U2792 , P3_U2791 , P3_U2790 , P3_U2789 , P3_U2788 ,
             P3_U2787 , P3_U2786 , P3_U2785 , P3_U2784 , P3_U2783 , P3_U2782 ,
             P3_U2781 , P3_U2780 , P3_U2779 , P3_U2778 , P3_U2777 , P3_U2776 ,
             P3_U2775 , P3_U2774 , P3_U2773 , P3_U2772 , P3_U2771 , P3_U2770 ,
             P3_U2769 , P3_U2768 , P3_U2767 , P3_U2766 , P3_U2765 , P3_U2764 ,
             P3_U2763 , P3_U2762 , P3_U2761 , P3_U2760 , P3_U2759 , P3_U2758 ,
             P3_U2757 , P3_U2756 , P3_U2755 , P3_U2754 , P3_U2753 , P3_U2752 ,
             P3_U2751 , P3_U2750 , P3_U2749 , P3_U2748 , P3_U2747 , P3_U2746 ,
             P3_U2745 , P3_U2744 , P3_U2743 , P3_U2742 , P3_U2741 , P3_U2740 ,
             P3_U2739 , P3_U2738 , P3_U2737 , P3_U2736 , P3_U2735 , P3_U2734 ,
             P3_U2733 , P3_U2732 , P3_U2731 , P3_U2730 , P3_U2729 , P3_U2728 ,
             P3_U2727 , P3_U2726 , P3_U2725 , P3_U2724 , P3_U2723 , P3_U2722 ,
             P3_U2721 , P3_U2720 , P3_U2719 , P3_U2718 , P3_U2717 , P3_U2716 ,
             P3_U2715 , P3_U2714 , P3_U2713 , P3_U2712 , P3_U2711 , P3_U2710 ,
             P3_U2709 , P3_U2708 , P3_U2707 , P3_U2706 , P3_U2705 , P3_U2704 ,
             P3_U2703 , P3_U2702 , P3_U2701 , P3_U2700 , P3_U2699 , P3_U2698 ,
             P3_U2697 , P3_U2696 , P3_U2695 , P3_U2694 , P3_U2693 , P3_U2692 ,
             P3_U2691 , P3_U2690 , P3_U2689 , P3_U2688 , P3_U2687 , P3_U2686 ,
             P3_U2685 , P3_U2684 , P3_U2683 , P3_U2682 , P3_U2681 , P3_U2680 ,
             P3_U2679 , P3_U2678 , P3_U2677 , P3_U2676 , P3_U2675 , P3_U2674 ,
             P3_U2673 , P3_U2672 , P3_U2671 , P3_U2670 , P3_U2669 , P3_U2668 ,
             P3_U2667 , P3_U2666 , P3_U2665 , P3_U2664 , P3_U2663 , P3_U2662 ,
             P3_U2661 , P3_U2660 , P3_U2659 , P3_U2658 , P3_U2657 , P3_U2656 ,
             P3_U2655 , P3_U2654 , P3_U2653 , P3_U2652 , P3_U2651 , P3_U2650 ,
             P3_U2649 , P3_U2648 , P3_U2647 , P3_U2646 , P3_U2645 , P3_U2644 ,
             P3_U2643 , P3_U2642 , P3_U2641 , P3_U2640 , P3_U2639 , P3_U3292 ,
             P3_U2638 , P3_U3293 , P3_U3294 , P3_U2637 , P3_U3295 , P3_U2636 ,
             P3_U3296 , P3_U2635 , P3_U3297 , P3_U2634 , P3_U2633 , P3_U3298 ,
             P3_U3299 , P2_U3585 , P2_U3586 , P2_U3587 , P2_U3588 , P2_U3241 ,
             P2_U3240 , P2_U3239 , P2_U3238 , P2_U3237 , P2_U3236 , P2_U3235 ,
             P2_U3234 , P2_U3233 , P2_U3232 , P2_U3231 , P2_U3230 , P2_U3229 ,
             P2_U3228 , P2_U3227 , P2_U3226 , P2_U3225 , P2_U3224 , P2_U3223 ,
             P2_U3222 , P2_U3221 , P2_U3220 , P2_U3219 , P2_U3218 , P2_U3217 ,
             P2_U3216 , P2_U3215 , P2_U3214 , P2_U3213 , P2_U3212 , P2_U3211 ,
             P2_U3210 , P2_U3209 , P2_U3591 , P2_U3592 , P2_U3208 , P2_U3207 ,
             P2_U3206 , P2_U3205 , P2_U3204 , P2_U3203 , P2_U3202 , P2_U3201 ,
             P2_U3200 , P2_U3199 , P2_U3198 , P2_U3197 , P2_U3196 , P2_U3195 ,
             P2_U3194 , P2_U3193 , P2_U3192 , P2_U3191 , P2_U3190 , P2_U3189 ,
             P2_U3188 , P2_U3187 , P2_U3186 , P2_U3185 , P2_U3184 , P2_U3183 ,
             P2_U3182 , P2_U3181 , P2_U3180 , P2_U3179 , P2_U3593 , P2_U3178 ,
             P2_U3177 , P2_U3176 , P2_U3175 , P2_U3174 , P2_U3173 , P2_U3172 ,
             P2_U3171 , P2_U3170 , P2_U3169 , P2_U3168 , P2_U3167 , P2_U3166 ,
             P2_U3165 , P2_U3164 , P2_U3163 , P2_U3162 , P2_U3161 , P2_U3160 ,
             P2_U3159 , P2_U3158 , P2_U3157 , P2_U3156 , P2_U3155 , P2_U3154 ,
             P2_U3153 , P2_U3152 , P2_U3151 , P2_U3150 , P2_U3149 , P2_U3148 ,
             P2_U3147 , P2_U3146 , P2_U3145 , P2_U3144 , P2_U3143 , P2_U3142 ,
             P2_U3141 , P2_U3140 , P2_U3139 , P2_U3138 , P2_U3137 , P2_U3136 ,
             P2_U3135 , P2_U3134 , P2_U3133 , P2_U3132 , P2_U3131 , P2_U3130 ,
             P2_U3129 , P2_U3128 , P2_U3127 , P2_U3126 , P2_U3125 , P2_U3124 ,
             P2_U3123 , P2_U3122 , P2_U3121 , P2_U3120 , P2_U3119 , P2_U3118 ,
             P2_U3117 , P2_U3116 , P2_U3115 , P2_U3114 , P2_U3113 , P2_U3112 ,
             P2_U3111 , P2_U3110 , P2_U3109 , P2_U3108 , P2_U3107 , P2_U3106 ,
             P2_U3105 , P2_U3104 , P2_U3103 , P2_U3102 , P2_U3101 , P2_U3100 ,
             P2_U3099 , P2_U3098 , P2_U3097 , P2_U3096 , P2_U3095 , P2_U3094 ,
             P2_U3093 , P2_U3092 , P2_U3091 , P2_U3090 , P2_U3089 , P2_U3088 ,
             P2_U3087 , P2_U3086 , P2_U3085 , P2_U3084 , P2_U3083 , P2_U3082 ,
             P2_U3081 , P2_U3080 , P2_U3079 , P2_U3078 , P2_U3077 , P2_U3076 ,
             P2_U3075 , P2_U3074 , P2_U3073 , P2_U3072 , P2_U3071 , P2_U3070 ,
             P2_U3069 , P2_U3068 , P2_U3067 , P2_U3066 , P2_U3065 , P2_U3064 ,
             P2_U3063 , P2_U3062 , P2_U3061 , P2_U3060 , P2_U3059 , P2_U3058 ,
             P2_U3057 , P2_U3056 , P2_U3055 , P2_U3054 , P2_U3053 , P2_U3052 ,
             P2_U3051 , P2_U3050 , P2_U3049 , P2_U3048 , P2_U3595 , P2_U3596 ,
             P2_U3599 , P2_U3600 , P2_U3601 , P2_U3047 , P2_U3602 , P2_U3603 ,
             P2_U3604 , P2_U3605 , P2_U3046 , P2_U3045 , P2_U3044 , P2_U3043 ,
             P2_U3042 , P2_U3041 , P2_U3040 , P2_U3039 , P2_U3038 , P2_U3037 ,
             P2_U3036 , P2_U3035 , P2_U3034 , P2_U3033 , P2_U3032 , P2_U3031 ,
             P2_U3030 , P2_U3029 , P2_U3028 , P2_U3027 , P2_U3026 , P2_U3025 ,
             P2_U3024 , P2_U3023 , P2_U3022 , P2_U3021 , P2_U3020 , P2_U3019 ,
             P2_U3018 , P2_U3017 , P2_U3016 , P2_U3015 , P2_U3014 , P2_U3013 ,
             P2_U3012 , P2_U3011 , P2_U3010 , P2_U3009 , P2_U3008 , P2_U3007 ,
             P2_U3006 , P2_U3005 , P2_U3004 , P2_U3003 , P2_U3002 , P2_U3001 ,
             P2_U3000 , P2_U2999 , P2_U2998 , P2_U2997 , P2_U2996 , P2_U2995 ,
             P2_U2994 , P2_U2993 , P2_U2992 , P2_U2991 , P2_U2990 , P2_U2989 ,
             P2_U2988 , P2_U2987 , P2_U2986 , P2_U2985 , P2_U2984 , P2_U2983 ,
             P2_U2982 , P2_U2981 , P2_U2980 , P2_U2979 , P2_U2978 , P2_U2977 ,
             P2_U2976 , P2_U2975 , P2_U2974 , P2_U2973 , P2_U2972 , P2_U2971 ,
             P2_U2970 , P2_U2969 , P2_U2968 , P2_U2967 , P2_U2966 , P2_U2965 ,
             P2_U2964 , P2_U2963 , P2_U2962 , P2_U2961 , P2_U2960 , P2_U2959 ,
             P2_U2958 , P2_U2957 , P2_U2956 , P2_U2955 , P2_U2954 , P2_U2953 ,
             P2_U2952 , P2_U2951 , P2_U2950 , P2_U2949 , P2_U2948 , P2_U2947 ,
             P2_U2946 , P2_U2945 , P2_U2944 , P2_U2943 , P2_U2942 , P2_U2941 ,
             P2_U2940 , P2_U2939 , P2_U2938 , P2_U2937 , P2_U2936 , P2_U2935 ,
             P2_U2934 , P2_U2933 , P2_U2932 , P2_U2931 , P2_U2930 , P2_U2929 ,
             P2_U2928 , P2_U2927 , P2_U2926 , P2_U2925 , P2_U2924 , P2_U2923 ,
             P2_U2922 , P2_U2921 , P2_U2920 , P2_U2919 , P2_U2918 , P2_U2917 ,
             P2_U2916 , P2_U2915 , P2_U2914 , P2_U2913 , P2_U2912 , P2_U2911 ,
             P2_U2910 , P2_U2909 , P2_U2908 , P2_U2907 , P2_U2906 , P2_U2905 ,
             P2_U2904 , P2_U2903 , P2_U2902 , P2_U2901 , P2_U2900 , P2_U2899 ,
             P2_U2898 , P2_U2897 , P2_U2896 , P2_U2895 , P2_U2894 , P2_U2893 ,
             P2_U2892 , P2_U2891 , P2_U2890 , P2_U2889 , P2_U2888 , P2_U2887 ,
             P2_U2886 , P2_U2885 , P2_U2884 , P2_U2883 , P2_U2882 , P2_U2881 ,
             P2_U2880 , P2_U2879 , P2_U2878 , P2_U2877 , P2_U2876 , P2_U2875 ,
             P2_U2874 , P2_U2873 , P2_U2872 , P2_U2871 , P2_U2870 , P2_U2869 ,
             P2_U2868 , P2_U2867 , P2_U2866 , P2_U2865 , P2_U2864 , P2_U2863 ,
             P2_U2862 , P2_U2861 , P2_U2860 , P2_U2859 , P2_U2858 , P2_U2857 ,
             P2_U2856 , P2_U2855 , P2_U2854 , P2_U2853 , P2_U2852 , P2_U2851 ,
             P2_U2850 , P2_U2849 , P2_U2848 , P2_U2847 , P2_U2846 , P2_U2845 ,
             P2_U2844 , P2_U2843 , P2_U2842 , P2_U2841 , P2_U2840 , P2_U2839 ,
             P2_U2838 , P2_U2837 , P2_U2836 , P2_U2835 , P2_U2834 , P2_U2833 ,
             P2_U2832 , P2_U2831 , P2_U2830 , P2_U2829 , P2_U2828 , P2_U2827 ,
             P2_U2826 , P2_U2825 , P2_U2824 , P2_U2823 , P2_U2822 , P2_U2821 ,
             P2_U2820 , P2_U3608 , P2_U2819 , P2_U3609 , P2_U2818 , P2_U3610 ,
             P2_U2817 , P2_U3611 , P2_U2816 , P2_U2815 , P2_U3612 , P2_U2814 ,
             P1_U3458 , P1_U3459 , P1_U3460 , P1_U3461 , P1_U3226 , P1_U3225 ,
             P1_U3224 , P1_U3223 , P1_U3222 , P1_U3221 , P1_U3220 , P1_U3219 ,
             P1_U3218 , P1_U3217 , P1_U3216 , P1_U3215 , P1_U3214 , P1_U3213 ,
             P1_U3212 , P1_U3211 , P1_U3210 , P1_U3209 , P1_U3208 , P1_U3207 ,
             P1_U3206 , P1_U3205 , P1_U3204 , P1_U3203 , P1_U3202 , P1_U3201 ,
             P1_U3200 , P1_U3199 , P1_U3198 , P1_U3197 , P1_U3196 , P1_U3195 ,
             P1_U3194 , P1_U3464 , P1_U3465 , P1_U3193 , P1_U3192 , P1_U3191 ,
             P1_U3190 , P1_U3189 , P1_U3188 , P1_U3187 , P1_U3186 , P1_U3185 ,
             P1_U3184 , P1_U3183 , P1_U3182 , P1_U3181 , P1_U3180 , P1_U3179 ,
             P1_U3178 , P1_U3177 , P1_U3176 , P1_U3175 , P1_U3174 , P1_U3173 ,
             P1_U3172 , P1_U3171 , P1_U3170 , P1_U3169 , P1_U3168 , P1_U3167 ,
             P1_U3166 , P1_U3165 , P1_U3164 , P1_U3466 , P1_U3163 , P1_U3162 ,
             P1_U3161 , P1_U3160 , P1_U3159 , P1_U3158 , P1_U3157 , P1_U3156 ,
             P1_U3155 , P1_U3154 , P1_U3153 , P1_U3152 , P1_U3151 , P1_U3150 ,
             P1_U3149 , P1_U3148 , P1_U3147 , P1_U3146 , P1_U3145 , P1_U3144 ,
             P1_U3143 , P1_U3142 , P1_U3141 , P1_U3140 , P1_U3139 , P1_U3138 ,
             P1_U3137 , P1_U3136 , P1_U3135 , P1_U3134 , P1_U3133 , P1_U3132 ,
             P1_U3131 , P1_U3130 , P1_U3129 , P1_U3128 , P1_U3127 , P1_U3126 ,
             P1_U3125 , P1_U3124 , P1_U3123 , P1_U3122 , P1_U3121 , P1_U3120 ,
             P1_U3119 , P1_U3118 , P1_U3117 , P1_U3116 , P1_U3115 , P1_U3114 ,
             P1_U3113 , P1_U3112 , P1_U3111 , P1_U3110 , P1_U3109 , P1_U3108 ,
             P1_U3107 , P1_U3106 , P1_U3105 , P1_U3104 , P1_U3103 , P1_U3102 ,
             P1_U3101 , P1_U3100 , P1_U3099 , P1_U3098 , P1_U3097 , P1_U3096 ,
             P1_U3095 , P1_U3094 , P1_U3093 , P1_U3092 , P1_U3091 , P1_U3090 ,
             P1_U3089 , P1_U3088 , P1_U3087 , P1_U3086 , P1_U3085 , P1_U3084 ,
             P1_U3083 , P1_U3082 , P1_U3081 , P1_U3080 , P1_U3079 , P1_U3078 ,
             P1_U3077 , P1_U3076 , P1_U3075 , P1_U3074 , P1_U3073 , P1_U3072 ,
             P1_U3071 , P1_U3070 , P1_U3069 , P1_U3068 , P1_U3067 , P1_U3066 ,
             P1_U3065 , P1_U3064 , P1_U3063 , P1_U3062 , P1_U3061 , P1_U3060 ,
             P1_U3059 , P1_U3058 , P1_U3057 , P1_U3056 , P1_U3055 , P1_U3054 ,
             P1_U3053 , P1_U3052 , P1_U3051 , P1_U3050 , P1_U3049 , P1_U3048 ,
             P1_U3047 , P1_U3046 , P1_U3045 , P1_U3044 , P1_U3043 , P1_U3042 ,
             P1_U3041 , P1_U3040 , P1_U3039 , P1_U3038 , P1_U3037 , P1_U3036 ,
             P1_U3035 , P1_U3034 , P1_U3033 , P1_U3468 , P1_U3469 , P1_U3472 ,
             P1_U3473 , P1_U3474 , P1_U3032 , P1_U3475 , P1_U3476 , P1_U3477 ,
             P1_U3478 , P1_U3031 , P1_U3030 , P1_U3029 , P1_U3028 , P1_U3027 ,
             P1_U3026 , P1_U3025 , P1_U3024 , P1_U3023 , P1_U3022 , P1_U3021 ,
             P1_U3020 , P1_U3019 , P1_U3018 , P1_U3017 , P1_U3016 , P1_U3015 ,
             P1_U3014 , P1_U3013 , P1_U3012 , P1_U3011 , P1_U3010 , P1_U3009 ,
             P1_U3008 , P1_U3007 , P1_U3006 , P1_U3005 , P1_U3004 , P1_U3003 ,
             P1_U3002 , P1_U3001 , P1_U3000 , P1_U2999 , P1_U2998 , P1_U2997 ,
             P1_U2996 , P1_U2995 , P1_U2994 , P1_U2993 , P1_U2992 , P1_U2991 ,
             P1_U2990 , P1_U2989 , P1_U2988 , P1_U2987 , P1_U2986 , P1_U2985 ,
             P1_U2984 , P1_U2983 , P1_U2982 , P1_U2981 , P1_U2980 , P1_U2979 ,
             P1_U2978 , P1_U2977 , P1_U2976 , P1_U2975 , P1_U2974 , P1_U2973 ,
             P1_U2972 , P1_U2971 , P1_U2970 , P1_U2969 , P1_U2968 , P1_U2967 ,
             P1_U2966 , P1_U2965 , P1_U2964 , P1_U2963 , P1_U2962 , P1_U2961 ,
             P1_U2960 , P1_U2959 , P1_U2958 , P1_U2957 , P1_U2956 , P1_U2955 ,
             P1_U2954 , P1_U2953 , P1_U2952 , P1_U2951 , P1_U2950 , P1_U2949 ,
             P1_U2948 , P1_U2947 , P1_U2946 , P1_U2945 , P1_U2944 , P1_U2943 ,
             P1_U2942 , P1_U2941 , P1_U2940 , P1_U2939 , P1_U2938 , P1_U2937 ,
             P1_U2936 , P1_U2935 , P1_U2934 , P1_U2933 , P1_U2932 , P1_U2931 ,
             P1_U2930 , P1_U2929 , P1_U2928 , P1_U2927 , P1_U2926 , P1_U2925 ,
             P1_U2924 , P1_U2923 , P1_U2922 , P1_U2921 , P1_U2920 , P1_U2919 ,
             P1_U2918 , P1_U2917 , P1_U2916 , P1_U2915 , P1_U2914 , P1_U2913 ,
             P1_U2912 , P1_U2911 , P1_U2910 , P1_U2909 , P1_U2908 , P1_U2907 ,
             P1_U2906 , P1_U2905 , P1_U2904 , P1_U2903 , P1_U2902 , P1_U2901 ,
             P1_U2900 , P1_U2899 , P1_U2898 , P1_U2897 , P1_U2896 , P1_U2895 ,
             P1_U2894 , P1_U2893 , P1_U2892 , P1_U2891 , P1_U2890 , P1_U2889 ,
             P1_U2888 , P1_U2887 , P1_U2886 , P1_U2885 , P1_U2884 , P1_U2883 ,
             P1_U2882 , P1_U2881 , P1_U2880 , P1_U2879 , P1_U2878 , P1_U2877 ,
             P1_U2876 , P1_U2875 , P1_U2874 , P1_U2873 , P1_U2872 , P1_U2871 ,
             P1_U2870 , P1_U2869 , P1_U2868 , P1_U2867 , P1_U2866 , P1_U2865 ,
             P1_U2864 , P1_U2863 , P1_U2862 , P1_U2861 , P1_U2860 , P1_U2859 ,
             P1_U2858 , P1_U2857 , P1_U2856 , P1_U2855 , P1_U2854 , P1_U2853 ,
             P1_U2852 , P1_U2851 , P1_U2850 , P1_U2849 , P1_U2848 , P1_U2847 ,
             P1_U2846 , P1_U2845 , P1_U2844 , P1_U2843 , P1_U2842 , P1_U2841 ,
             P1_U2840 , P1_U2839 , P1_U2838 , P1_U2837 , P1_U2836 , P1_U2835 ,
             P1_U2834 , P1_U2833 , P1_U2832 , P1_U2831 , P1_U2830 , P1_U2829 ,
             P1_U2828 , P1_U2827 , P1_U2826 , P1_U2825 , P1_U2824 , P1_U2823 ,
             P1_U2822 , P1_U2821 , P1_U2820 , P1_U2819 , P1_U2818 , P1_U2817 ,
             P1_U2816 , P1_U2815 , P1_U2814 , P1_U2813 , P1_U2812 , P1_U2811 ,
             P1_U2810 , P1_U2809 , P1_U2808 , P1_U3481 , P1_U2807 , P1_U3482 ,
             P1_U3483 , P1_U2806 , P1_U3484 , P1_U2805 , P1_U3485 , P1_U2804 ,
             P1_U3486 , P1_U2803 , P1_U2802 , P1_U3487 , P1_U2801 , P3_DATAO_REG_31_ ,
             P3_DATAO_REG_30_ , P3_DATAO_REG_29_ , P3_DATAO_REG_28_ , P3_DATAO_REG_27_ , P3_DATAO_REG_26_ , P3_DATAO_REG_25_ ,
             P3_DATAO_REG_24_ , P3_DATAO_REG_23_ , P3_DATAO_REG_22_ , P3_DATAO_REG_21_ , P3_DATAO_REG_20_ , P3_DATAO_REG_19_ ,
             P3_DATAO_REG_18_ , P3_DATAO_REG_17_ , P3_DATAO_REG_16_ , P3_DATAO_REG_15_ , P3_DATAO_REG_14_ , P3_DATAO_REG_13_ ,
             P3_DATAO_REG_12_ , P3_DATAO_REG_11_ , P3_DATAO_REG_10_ , P3_DATAO_REG_9_ , P3_DATAO_REG_8_ , P3_DATAO_REG_7_ ,
             P3_DATAO_REG_6_ , P3_DATAO_REG_5_ , P3_DATAO_REG_4_ , P3_DATAO_REG_3_ , P3_DATAO_REG_2_ , P3_DATAO_REG_1_ ,
             P3_DATAO_REG_0_ , P1_ADDRESS_REG_29_ , P1_ADDRESS_REG_28_ , P1_ADDRESS_REG_27_ , P1_ADDRESS_REG_26_ , P1_ADDRESS_REG_25_ ,
             P1_ADDRESS_REG_24_ , P1_ADDRESS_REG_23_ , P1_ADDRESS_REG_22_ , P1_ADDRESS_REG_21_ , P1_ADDRESS_REG_20_ , P1_ADDRESS_REG_19_ ,
             P1_ADDRESS_REG_18_ , P1_ADDRESS_REG_17_ , P1_ADDRESS_REG_16_ , P1_ADDRESS_REG_15_ , P1_ADDRESS_REG_14_ , P1_ADDRESS_REG_13_ ,
             P1_ADDRESS_REG_12_ , P1_ADDRESS_REG_11_ , P1_ADDRESS_REG_10_ , P1_ADDRESS_REG_9_ , P1_ADDRESS_REG_8_ , P1_ADDRESS_REG_7_ ,
             P1_ADDRESS_REG_6_ , P1_ADDRESS_REG_5_ , P1_ADDRESS_REG_4_ , P1_ADDRESS_REG_3_ , P1_ADDRESS_REG_2_ , P1_ADDRESS_REG_1_ ,
             P1_ADDRESS_REG_0_ , U355 , U356 , U357 , U358 , U359 ,
             U360 , U361 , U362 , U363 , U364 , U366 ,
             U367 , U368 , U369 , U370 , U371 , U372 ,
             U373 , U374 , U375 , U347 , U348 , U349 ,
             U350 , U351 , U352 , U353 , U354 , U365 ,
             U376 , P3_W_R_N_REG , P3_D_C_N_REG , P3_M_IO_N_REG , P1_ADS_N_REG , P3_ADS_N_REG ,
            
             BUF1_REG_0_ , BUF1_REG_1_ , BUF1_REG_2_ , BUF1_REG_3_ , BUF1_REG_4_ , BUF1_REG_5_ ,
             BUF1_REG_6_ , BUF1_REG_7_ , BUF1_REG_8_ , BUF1_REG_9_ , BUF1_REG_10_ , BUF1_REG_11_ ,
             BUF1_REG_12_ , BUF1_REG_13_ , BUF1_REG_14_ , BUF1_REG_15_ , BUF1_REG_16_ , BUF1_REG_17_ ,
             BUF1_REG_18_ , BUF1_REG_19_ , BUF1_REG_20_ , BUF1_REG_21_ , BUF1_REG_22_ , BUF1_REG_23_ ,
             BUF1_REG_24_ , BUF1_REG_25_ , BUF1_REG_26_ , BUF1_REG_27_ , BUF1_REG_28_ , BUF1_REG_29_ ,
             BUF1_REG_30_ , BUF1_REG_31_ , BUF2_REG_0_ , BUF2_REG_1_ , BUF2_REG_2_ , BUF2_REG_3_ ,
             BUF2_REG_4_ , BUF2_REG_5_ , BUF2_REG_6_ , BUF2_REG_7_ , BUF2_REG_8_ , BUF2_REG_9_ ,
             BUF2_REG_10_ , BUF2_REG_11_ , BUF2_REG_12_ , BUF2_REG_13_ , BUF2_REG_14_ , BUF2_REG_15_ ,
             BUF2_REG_16_ , BUF2_REG_17_ , BUF2_REG_18_ , BUF2_REG_19_ , BUF2_REG_20_ , BUF2_REG_21_ ,
             BUF2_REG_22_ , BUF2_REG_23_ , BUF2_REG_24_ , BUF2_REG_25_ , BUF2_REG_26_ , BUF2_REG_27_ ,
             BUF2_REG_28_ , BUF2_REG_29_ , BUF2_REG_30_ , BUF2_REG_31_ , READY12_REG , READY21_REG ,
             READY22_REG , READY11_REG , P3_BE_N_REG_3_ , P3_BE_N_REG_2_ , P3_BE_N_REG_1_ , P3_BE_N_REG_0_ ,
             P3_ADDRESS_REG_29_ , P3_ADDRESS_REG_28_ , P3_ADDRESS_REG_27_ , P3_ADDRESS_REG_26_ , P3_ADDRESS_REG_25_ , P3_ADDRESS_REG_24_ ,
             P3_ADDRESS_REG_23_ , P3_ADDRESS_REG_22_ , P3_ADDRESS_REG_21_ , P3_ADDRESS_REG_20_ , P3_ADDRESS_REG_19_ , P3_ADDRESS_REG_18_ ,
             P3_ADDRESS_REG_17_ , P3_ADDRESS_REG_16_ , P3_ADDRESS_REG_15_ , P3_ADDRESS_REG_14_ , P3_ADDRESS_REG_13_ , P3_ADDRESS_REG_12_ ,
             P3_ADDRESS_REG_11_ , P3_ADDRESS_REG_10_ , P3_ADDRESS_REG_9_ , P3_ADDRESS_REG_8_ , P3_ADDRESS_REG_7_ , P3_ADDRESS_REG_6_ ,
             P3_ADDRESS_REG_5_ , P3_ADDRESS_REG_4_ , P3_ADDRESS_REG_3_ , P3_ADDRESS_REG_2_ , P3_ADDRESS_REG_1_ , P3_ADDRESS_REG_0_ ,
             P3_STATE_REG_2_ , P3_STATE_REG_1_ , P3_STATE_REG_0_ , P3_DATAWIDTH_REG_0_ , P3_DATAWIDTH_REG_1_ , P3_DATAWIDTH_REG_2_ ,
             P3_DATAWIDTH_REG_3_ , P3_DATAWIDTH_REG_4_ , P3_DATAWIDTH_REG_5_ , P3_DATAWIDTH_REG_6_ , P3_DATAWIDTH_REG_7_ , P3_DATAWIDTH_REG_8_ ,
             P3_DATAWIDTH_REG_9_ , P3_DATAWIDTH_REG_10_ , P3_DATAWIDTH_REG_11_ , P3_DATAWIDTH_REG_12_ , P3_DATAWIDTH_REG_13_ , P3_DATAWIDTH_REG_14_ ,
             P3_DATAWIDTH_REG_15_ , P3_DATAWIDTH_REG_16_ , P3_DATAWIDTH_REG_17_ , P3_DATAWIDTH_REG_18_ , P3_DATAWIDTH_REG_19_ , P3_DATAWIDTH_REG_20_ ,
             P3_DATAWIDTH_REG_21_ , P3_DATAWIDTH_REG_22_ , P3_DATAWIDTH_REG_23_ , P3_DATAWIDTH_REG_24_ , P3_DATAWIDTH_REG_25_ , P3_DATAWIDTH_REG_26_ ,
             P3_DATAWIDTH_REG_27_ , P3_DATAWIDTH_REG_28_ , P3_DATAWIDTH_REG_29_ , P3_DATAWIDTH_REG_30_ , P3_DATAWIDTH_REG_31_ , P3_STATE2_REG_3_ ,
             P3_STATE2_REG_2_ , P3_STATE2_REG_1_ , P3_STATE2_REG_0_ , P3_INSTQUEUE_REG_15__7_ , P3_INSTQUEUE_REG_15__6_ , P3_INSTQUEUE_REG_15__5_ ,
             P3_INSTQUEUE_REG_15__4_ , P3_INSTQUEUE_REG_15__3_ , P3_INSTQUEUE_REG_15__2_ , P3_INSTQUEUE_REG_15__1_ , P3_INSTQUEUE_REG_15__0_ , P3_INSTQUEUE_REG_14__7_ ,
             P3_INSTQUEUE_REG_14__6_ , P3_INSTQUEUE_REG_14__5_ , P3_INSTQUEUE_REG_14__4_ , P3_INSTQUEUE_REG_14__3_ , P3_INSTQUEUE_REG_14__2_ , P3_INSTQUEUE_REG_14__1_ ,
             P3_INSTQUEUE_REG_14__0_ , P3_INSTQUEUE_REG_13__7_ , P3_INSTQUEUE_REG_13__6_ , P3_INSTQUEUE_REG_13__5_ , P3_INSTQUEUE_REG_13__4_ , P3_INSTQUEUE_REG_13__3_ ,
             P3_INSTQUEUE_REG_13__2_ , P3_INSTQUEUE_REG_13__1_ , P3_INSTQUEUE_REG_13__0_ , P3_INSTQUEUE_REG_12__7_ , P3_INSTQUEUE_REG_12__6_ , P3_INSTQUEUE_REG_12__5_ ,
             P3_INSTQUEUE_REG_12__4_ , P3_INSTQUEUE_REG_12__3_ , P3_INSTQUEUE_REG_12__2_ , P3_INSTQUEUE_REG_12__1_ , P3_INSTQUEUE_REG_12__0_ , P3_INSTQUEUE_REG_11__7_ ,
             P3_INSTQUEUE_REG_11__6_ , P3_INSTQUEUE_REG_11__5_ , P3_INSTQUEUE_REG_11__4_ , P3_INSTQUEUE_REG_11__3_ , P3_INSTQUEUE_REG_11__2_ , P3_INSTQUEUE_REG_11__1_ ,
             P3_INSTQUEUE_REG_11__0_ , P3_INSTQUEUE_REG_10__7_ , P3_INSTQUEUE_REG_10__6_ , P3_INSTQUEUE_REG_10__5_ , P3_INSTQUEUE_REG_10__4_ , P3_INSTQUEUE_REG_10__3_ ,
             P3_INSTQUEUE_REG_10__2_ , P3_INSTQUEUE_REG_10__1_ , P3_INSTQUEUE_REG_10__0_ , P3_INSTQUEUE_REG_9__7_ , P3_INSTQUEUE_REG_9__6_ , P3_INSTQUEUE_REG_9__5_ ,
             P3_INSTQUEUE_REG_9__4_ , P3_INSTQUEUE_REG_9__3_ , P3_INSTQUEUE_REG_9__2_ , P3_INSTQUEUE_REG_9__1_ , P3_INSTQUEUE_REG_9__0_ , P3_INSTQUEUE_REG_8__7_ ,
             P3_INSTQUEUE_REG_8__6_ , P3_INSTQUEUE_REG_8__5_ , P3_INSTQUEUE_REG_8__4_ , P3_INSTQUEUE_REG_8__3_ , P3_INSTQUEUE_REG_8__2_ , P3_INSTQUEUE_REG_8__1_ ,
             P3_INSTQUEUE_REG_8__0_ , P3_INSTQUEUE_REG_7__7_ , P3_INSTQUEUE_REG_7__6_ , P3_INSTQUEUE_REG_7__5_ , P3_INSTQUEUE_REG_7__4_ , P3_INSTQUEUE_REG_7__3_ ,
             P3_INSTQUEUE_REG_7__2_ , P3_INSTQUEUE_REG_7__1_ , P3_INSTQUEUE_REG_7__0_ , P3_INSTQUEUE_REG_6__7_ , P3_INSTQUEUE_REG_6__6_ , P3_INSTQUEUE_REG_6__5_ ,
             P3_INSTQUEUE_REG_6__4_ , P3_INSTQUEUE_REG_6__3_ , P3_INSTQUEUE_REG_6__2_ , P3_INSTQUEUE_REG_6__1_ , P3_INSTQUEUE_REG_6__0_ , P3_INSTQUEUE_REG_5__7_ ,
             P3_INSTQUEUE_REG_5__6_ , P3_INSTQUEUE_REG_5__5_ , P3_INSTQUEUE_REG_5__4_ , P3_INSTQUEUE_REG_5__3_ , P3_INSTQUEUE_REG_5__2_ , P3_INSTQUEUE_REG_5__1_ ,
             P3_INSTQUEUE_REG_5__0_ , P3_INSTQUEUE_REG_4__7_ , P3_INSTQUEUE_REG_4__6_ , P3_INSTQUEUE_REG_4__5_ , P3_INSTQUEUE_REG_4__4_ , P3_INSTQUEUE_REG_4__3_ ,
             P3_INSTQUEUE_REG_4__2_ , P3_INSTQUEUE_REG_4__1_ , P3_INSTQUEUE_REG_4__0_ , P3_INSTQUEUE_REG_3__7_ , P3_INSTQUEUE_REG_3__6_ , P3_INSTQUEUE_REG_3__5_ ,
             P3_INSTQUEUE_REG_3__4_ , P3_INSTQUEUE_REG_3__3_ , P3_INSTQUEUE_REG_3__2_ , P3_INSTQUEUE_REG_3__1_ , P3_INSTQUEUE_REG_3__0_ , P3_INSTQUEUE_REG_2__7_ ,
             P3_INSTQUEUE_REG_2__6_ , P3_INSTQUEUE_REG_2__5_ , P3_INSTQUEUE_REG_2__4_ , P3_INSTQUEUE_REG_2__3_ , P3_INSTQUEUE_REG_2__2_ , P3_INSTQUEUE_REG_2__1_ ,
             P3_INSTQUEUE_REG_2__0_ , P3_INSTQUEUE_REG_1__7_ , P3_INSTQUEUE_REG_1__6_ , P3_INSTQUEUE_REG_1__5_ , P3_INSTQUEUE_REG_1__4_ , P3_INSTQUEUE_REG_1__3_ ,
             P3_INSTQUEUE_REG_1__2_ , P3_INSTQUEUE_REG_1__1_ , P3_INSTQUEUE_REG_1__0_ , P3_INSTQUEUE_REG_0__7_ , P3_INSTQUEUE_REG_0__6_ , P3_INSTQUEUE_REG_0__5_ ,
             P3_INSTQUEUE_REG_0__4_ , P3_INSTQUEUE_REG_0__3_ , P3_INSTQUEUE_REG_0__2_ , P3_INSTQUEUE_REG_0__1_ , P3_INSTQUEUE_REG_0__0_ , P3_INSTQUEUERD_ADDR_REG_4_ ,
             P3_INSTQUEUERD_ADDR_REG_3_ , P3_INSTQUEUERD_ADDR_REG_2_ , P3_INSTQUEUERD_ADDR_REG_1_ , P3_INSTQUEUERD_ADDR_REG_0_ , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_INSTQUEUEWR_ADDR_REG_3_ ,
             P3_INSTQUEUEWR_ADDR_REG_2_ , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_INSTADDRPOINTER_REG_0_ , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_2_ ,
             P3_INSTADDRPOINTER_REG_3_ , P3_INSTADDRPOINTER_REG_4_ , P3_INSTADDRPOINTER_REG_5_ , P3_INSTADDRPOINTER_REG_6_ , P3_INSTADDRPOINTER_REG_7_ , P3_INSTADDRPOINTER_REG_8_ ,
             P3_INSTADDRPOINTER_REG_9_ , P3_INSTADDRPOINTER_REG_10_ , P3_INSTADDRPOINTER_REG_11_ , P3_INSTADDRPOINTER_REG_12_ , P3_INSTADDRPOINTER_REG_13_ , P3_INSTADDRPOINTER_REG_14_ ,
             P3_INSTADDRPOINTER_REG_15_ , P3_INSTADDRPOINTER_REG_16_ , P3_INSTADDRPOINTER_REG_17_ , P3_INSTADDRPOINTER_REG_18_ , P3_INSTADDRPOINTER_REG_19_ , P3_INSTADDRPOINTER_REG_20_ ,
             P3_INSTADDRPOINTER_REG_21_ , P3_INSTADDRPOINTER_REG_22_ , P3_INSTADDRPOINTER_REG_23_ , P3_INSTADDRPOINTER_REG_24_ , P3_INSTADDRPOINTER_REG_25_ , P3_INSTADDRPOINTER_REG_26_ ,
             P3_INSTADDRPOINTER_REG_27_ , P3_INSTADDRPOINTER_REG_28_ , P3_INSTADDRPOINTER_REG_29_ , P3_INSTADDRPOINTER_REG_30_ , P3_INSTADDRPOINTER_REG_31_ , P3_PHYADDRPOINTER_REG_0_ ,
             P3_PHYADDRPOINTER_REG_1_ , P3_PHYADDRPOINTER_REG_2_ , P3_PHYADDRPOINTER_REG_3_ , P3_PHYADDRPOINTER_REG_4_ , P3_PHYADDRPOINTER_REG_5_ , P3_PHYADDRPOINTER_REG_6_ ,
             P3_PHYADDRPOINTER_REG_7_ , P3_PHYADDRPOINTER_REG_8_ , P3_PHYADDRPOINTER_REG_9_ , P3_PHYADDRPOINTER_REG_10_ , P3_PHYADDRPOINTER_REG_11_ , P3_PHYADDRPOINTER_REG_12_ ,
             P3_PHYADDRPOINTER_REG_13_ , P3_PHYADDRPOINTER_REG_14_ , P3_PHYADDRPOINTER_REG_15_ , P3_PHYADDRPOINTER_REG_16_ , P3_PHYADDRPOINTER_REG_17_ , P3_PHYADDRPOINTER_REG_18_ ,
             P3_PHYADDRPOINTER_REG_19_ , P3_PHYADDRPOINTER_REG_20_ , P3_PHYADDRPOINTER_REG_21_ , P3_PHYADDRPOINTER_REG_22_ , P3_PHYADDRPOINTER_REG_23_ , P3_PHYADDRPOINTER_REG_24_ ,
             P3_PHYADDRPOINTER_REG_25_ , P3_PHYADDRPOINTER_REG_26_ , P3_PHYADDRPOINTER_REG_27_ , P3_PHYADDRPOINTER_REG_28_ , P3_PHYADDRPOINTER_REG_29_ , P3_PHYADDRPOINTER_REG_30_ ,
             P3_PHYADDRPOINTER_REG_31_ , P3_LWORD_REG_15_ , P3_LWORD_REG_14_ , P3_LWORD_REG_13_ , P3_LWORD_REG_12_ , P3_LWORD_REG_11_ ,
             P3_LWORD_REG_10_ , P3_LWORD_REG_9_ , P3_LWORD_REG_8_ , P3_LWORD_REG_7_ , P3_LWORD_REG_6_ , P3_LWORD_REG_5_ ,
             P3_LWORD_REG_4_ , P3_LWORD_REG_3_ , P3_LWORD_REG_2_ , P3_LWORD_REG_1_ , P3_LWORD_REG_0_ , P3_UWORD_REG_14_ ,
             P3_UWORD_REG_13_ , P3_UWORD_REG_12_ , P3_UWORD_REG_11_ , P3_UWORD_REG_10_ , P3_UWORD_REG_9_ , P3_UWORD_REG_8_ ,
             P3_UWORD_REG_7_ , P3_UWORD_REG_6_ , P3_UWORD_REG_5_ , P3_UWORD_REG_4_ , P3_UWORD_REG_3_ , P3_UWORD_REG_2_ ,
             P3_UWORD_REG_1_ , P3_UWORD_REG_0_ , P3_DATAO_REG_0__EXTRA , P3_DATAO_REG_1__EXTRA , P3_DATAO_REG_2__EXTRA , P3_DATAO_REG_3__EXTRA ,
             P3_DATAO_REG_4__EXTRA , P3_DATAO_REG_5__EXTRA , P3_DATAO_REG_6__EXTRA , P3_DATAO_REG_7__EXTRA , P3_DATAO_REG_8__EXTRA , P3_DATAO_REG_9__EXTRA ,
             P3_DATAO_REG_10__EXTRA , P3_DATAO_REG_11__EXTRA , P3_DATAO_REG_12__EXTRA , P3_DATAO_REG_13__EXTRA , P3_DATAO_REG_14__EXTRA , P3_DATAO_REG_15__EXTRA ,
             P3_DATAO_REG_16__EXTRA , P3_DATAO_REG_17__EXTRA , P3_DATAO_REG_18__EXTRA , P3_DATAO_REG_19__EXTRA , P3_DATAO_REG_20__EXTRA , P3_DATAO_REG_21__EXTRA ,
             P3_DATAO_REG_22__EXTRA , P3_DATAO_REG_23__EXTRA , P3_DATAO_REG_24__EXTRA , P3_DATAO_REG_25__EXTRA , P3_DATAO_REG_26__EXTRA , P3_DATAO_REG_27__EXTRA ,
             P3_DATAO_REG_28__EXTRA , P3_DATAO_REG_29__EXTRA , P3_DATAO_REG_30__EXTRA , P3_DATAO_REG_31__EXTRA , P3_EAX_REG_0_ , P3_EAX_REG_1_ ,
             P3_EAX_REG_2_ , P3_EAX_REG_3_ , P3_EAX_REG_4_ , P3_EAX_REG_5_ , P3_EAX_REG_6_ , P3_EAX_REG_7_ ,
             P3_EAX_REG_8_ , P3_EAX_REG_9_ , P3_EAX_REG_10_ , P3_EAX_REG_11_ , P3_EAX_REG_12_ , P3_EAX_REG_13_ ,
             P3_EAX_REG_14_ , P3_EAX_REG_15_ , P3_EAX_REG_16_ , P3_EAX_REG_17_ , P3_EAX_REG_18_ , P3_EAX_REG_19_ ,
             P3_EAX_REG_20_ , P3_EAX_REG_21_ , P3_EAX_REG_22_ , P3_EAX_REG_23_ , P3_EAX_REG_24_ , P3_EAX_REG_25_ ,
             P3_EAX_REG_26_ , P3_EAX_REG_27_ , P3_EAX_REG_28_ , P3_EAX_REG_29_ , P3_EAX_REG_30_ , P3_EAX_REG_31_ ,
             P3_EBX_REG_0_ , P3_EBX_REG_1_ , P3_EBX_REG_2_ , P3_EBX_REG_3_ , P3_EBX_REG_4_ , P3_EBX_REG_5_ ,
             P3_EBX_REG_6_ , P3_EBX_REG_7_ , P3_EBX_REG_8_ , P3_EBX_REG_9_ , P3_EBX_REG_10_ , P3_EBX_REG_11_ ,
             P3_EBX_REG_12_ , P3_EBX_REG_13_ , P3_EBX_REG_14_ , P3_EBX_REG_15_ , P3_EBX_REG_16_ , P3_EBX_REG_17_ ,
             P3_EBX_REG_18_ , P3_EBX_REG_19_ , P3_EBX_REG_20_ , P3_EBX_REG_21_ , P3_EBX_REG_22_ , P3_EBX_REG_23_ ,
             P3_EBX_REG_24_ , P3_EBX_REG_25_ , P3_EBX_REG_26_ , P3_EBX_REG_27_ , P3_EBX_REG_28_ , P3_EBX_REG_29_ ,
             P3_EBX_REG_30_ , P3_EBX_REG_31_ , P3_REIP_REG_0_ , P3_REIP_REG_1_ , P3_REIP_REG_2_ , P3_REIP_REG_3_ ,
             P3_REIP_REG_4_ , P3_REIP_REG_5_ , P3_REIP_REG_6_ , P3_REIP_REG_7_ , P3_REIP_REG_8_ , P3_REIP_REG_9_ ,
             P3_REIP_REG_10_ , P3_REIP_REG_11_ , P3_REIP_REG_12_ , P3_REIP_REG_13_ , P3_REIP_REG_14_ , P3_REIP_REG_15_ ,
             P3_REIP_REG_16_ , P3_REIP_REG_17_ , P3_REIP_REG_18_ , P3_REIP_REG_19_ , P3_REIP_REG_20_ , P3_REIP_REG_21_ ,
             P3_REIP_REG_22_ , P3_REIP_REG_23_ , P3_REIP_REG_24_ , P3_REIP_REG_25_ , P3_REIP_REG_26_ , P3_REIP_REG_27_ ,
             P3_REIP_REG_28_ , P3_REIP_REG_29_ , P3_REIP_REG_30_ , P3_REIP_REG_31_ , P3_BYTEENABLE_REG_3_ , P3_BYTEENABLE_REG_2_ ,
             P3_BYTEENABLE_REG_1_ , P3_BYTEENABLE_REG_0_ , P3_W_R_N_REG_EXTRA , P3_FLUSH_REG , P3_MORE_REG , P3_STATEBS16_REG ,
             P3_REQUESTPENDING_REG , P3_D_C_N_REG_EXTRA , P3_M_IO_N_REG_EXTRA , P3_CODEFETCH_REG , P3_ADS_N_REG_EXTRA , P3_READREQUEST_REG ,
             P3_MEMORYFETCH_REG , P2_BE_N_REG_3_ , P2_BE_N_REG_2_ , P2_BE_N_REG_1_ , P2_BE_N_REG_0_ , P2_ADDRESS_REG_29_ ,
             P2_ADDRESS_REG_28_ , P2_ADDRESS_REG_27_ , P2_ADDRESS_REG_26_ , P2_ADDRESS_REG_25_ , P2_ADDRESS_REG_24_ , P2_ADDRESS_REG_23_ ,
             P2_ADDRESS_REG_22_ , P2_ADDRESS_REG_21_ , P2_ADDRESS_REG_20_ , P2_ADDRESS_REG_19_ , P2_ADDRESS_REG_18_ , P2_ADDRESS_REG_17_ ,
             P2_ADDRESS_REG_16_ , P2_ADDRESS_REG_15_ , P2_ADDRESS_REG_14_ , P2_ADDRESS_REG_13_ , P2_ADDRESS_REG_12_ , P2_ADDRESS_REG_11_ ,
             P2_ADDRESS_REG_10_ , P2_ADDRESS_REG_9_ , P2_ADDRESS_REG_8_ , P2_ADDRESS_REG_7_ , P2_ADDRESS_REG_6_ , P2_ADDRESS_REG_5_ ,
             P2_ADDRESS_REG_4_ , P2_ADDRESS_REG_3_ , P2_ADDRESS_REG_2_ , P2_ADDRESS_REG_1_ , P2_ADDRESS_REG_0_ , P2_STATE_REG_2_ ,
             P2_STATE_REG_1_ , P2_STATE_REG_0_ , P2_DATAWIDTH_REG_0_ , P2_DATAWIDTH_REG_1_ , P2_DATAWIDTH_REG_2_ , P2_DATAWIDTH_REG_3_ ,
             P2_DATAWIDTH_REG_4_ , P2_DATAWIDTH_REG_5_ , P2_DATAWIDTH_REG_6_ , P2_DATAWIDTH_REG_7_ , P2_DATAWIDTH_REG_8_ , P2_DATAWIDTH_REG_9_ ,
             P2_DATAWIDTH_REG_10_ , P2_DATAWIDTH_REG_11_ , P2_DATAWIDTH_REG_12_ , P2_DATAWIDTH_REG_13_ , P2_DATAWIDTH_REG_14_ , P2_DATAWIDTH_REG_15_ ,
             P2_DATAWIDTH_REG_16_ , P2_DATAWIDTH_REG_17_ , P2_DATAWIDTH_REG_18_ , P2_DATAWIDTH_REG_19_ , P2_DATAWIDTH_REG_20_ , P2_DATAWIDTH_REG_21_ ,
             P2_DATAWIDTH_REG_22_ , P2_DATAWIDTH_REG_23_ , P2_DATAWIDTH_REG_24_ , P2_DATAWIDTH_REG_25_ , P2_DATAWIDTH_REG_26_ , P2_DATAWIDTH_REG_27_ ,
             P2_DATAWIDTH_REG_28_ , P2_DATAWIDTH_REG_29_ , P2_DATAWIDTH_REG_30_ , P2_DATAWIDTH_REG_31_ , P2_STATE2_REG_3_ , P2_STATE2_REG_2_ ,
             P2_STATE2_REG_1_ , P2_STATE2_REG_0_ , P2_INSTQUEUE_REG_15__7_ , P2_INSTQUEUE_REG_15__6_ , P2_INSTQUEUE_REG_15__5_ , P2_INSTQUEUE_REG_15__4_ ,
             P2_INSTQUEUE_REG_15__3_ , P2_INSTQUEUE_REG_15__2_ , P2_INSTQUEUE_REG_15__1_ , P2_INSTQUEUE_REG_15__0_ , P2_INSTQUEUE_REG_14__7_ , P2_INSTQUEUE_REG_14__6_ ,
             P2_INSTQUEUE_REG_14__5_ , P2_INSTQUEUE_REG_14__4_ , P2_INSTQUEUE_REG_14__3_ , P2_INSTQUEUE_REG_14__2_ , P2_INSTQUEUE_REG_14__1_ , P2_INSTQUEUE_REG_14__0_ ,
             P2_INSTQUEUE_REG_13__7_ , P2_INSTQUEUE_REG_13__6_ , P2_INSTQUEUE_REG_13__5_ , P2_INSTQUEUE_REG_13__4_ , P2_INSTQUEUE_REG_13__3_ , P2_INSTQUEUE_REG_13__2_ ,
             P2_INSTQUEUE_REG_13__1_ , P2_INSTQUEUE_REG_13__0_ , P2_INSTQUEUE_REG_12__7_ , P2_INSTQUEUE_REG_12__6_ , P2_INSTQUEUE_REG_12__5_ , P2_INSTQUEUE_REG_12__4_ ,
             P2_INSTQUEUE_REG_12__3_ , P2_INSTQUEUE_REG_12__2_ , P2_INSTQUEUE_REG_12__1_ , P2_INSTQUEUE_REG_12__0_ , P2_INSTQUEUE_REG_11__7_ , P2_INSTQUEUE_REG_11__6_ ,
             P2_INSTQUEUE_REG_11__5_ , P2_INSTQUEUE_REG_11__4_ , P2_INSTQUEUE_REG_11__3_ , P2_INSTQUEUE_REG_11__2_ , P2_INSTQUEUE_REG_11__1_ , P2_INSTQUEUE_REG_11__0_ ,
             P2_INSTQUEUE_REG_10__7_ , P2_INSTQUEUE_REG_10__6_ , P2_INSTQUEUE_REG_10__5_ , P2_INSTQUEUE_REG_10__4_ , P2_INSTQUEUE_REG_10__3_ , P2_INSTQUEUE_REG_10__2_ ,
             P2_INSTQUEUE_REG_10__1_ , P2_INSTQUEUE_REG_10__0_ , P2_INSTQUEUE_REG_9__7_ , P2_INSTQUEUE_REG_9__6_ , P2_INSTQUEUE_REG_9__5_ , P2_INSTQUEUE_REG_9__4_ ,
             P2_INSTQUEUE_REG_9__3_ , P2_INSTQUEUE_REG_9__2_ , P2_INSTQUEUE_REG_9__1_ , P2_INSTQUEUE_REG_9__0_ , P2_INSTQUEUE_REG_8__7_ , P2_INSTQUEUE_REG_8__6_ ,
             P2_INSTQUEUE_REG_8__5_ , P2_INSTQUEUE_REG_8__4_ , P2_INSTQUEUE_REG_8__3_ , P2_INSTQUEUE_REG_8__2_ , P2_INSTQUEUE_REG_8__1_ , P2_INSTQUEUE_REG_8__0_ ,
             P2_INSTQUEUE_REG_7__7_ , P2_INSTQUEUE_REG_7__6_ , P2_INSTQUEUE_REG_7__5_ , P2_INSTQUEUE_REG_7__4_ , P2_INSTQUEUE_REG_7__3_ , P2_INSTQUEUE_REG_7__2_ ,
             P2_INSTQUEUE_REG_7__1_ , P2_INSTQUEUE_REG_7__0_ , P2_INSTQUEUE_REG_6__7_ , P2_INSTQUEUE_REG_6__6_ , P2_INSTQUEUE_REG_6__5_ , P2_INSTQUEUE_REG_6__4_ ,
             P2_INSTQUEUE_REG_6__3_ , P2_INSTQUEUE_REG_6__2_ , P2_INSTQUEUE_REG_6__1_ , P2_INSTQUEUE_REG_6__0_ , P2_INSTQUEUE_REG_5__7_ , P2_INSTQUEUE_REG_5__6_ ,
             P2_INSTQUEUE_REG_5__5_ , P2_INSTQUEUE_REG_5__4_ , P2_INSTQUEUE_REG_5__3_ , P2_INSTQUEUE_REG_5__2_ , P2_INSTQUEUE_REG_5__1_ , P2_INSTQUEUE_REG_5__0_ ,
             P2_INSTQUEUE_REG_4__7_ , P2_INSTQUEUE_REG_4__6_ , P2_INSTQUEUE_REG_4__5_ , P2_INSTQUEUE_REG_4__4_ , P2_INSTQUEUE_REG_4__3_ , P2_INSTQUEUE_REG_4__2_ ,
             P2_INSTQUEUE_REG_4__1_ , P2_INSTQUEUE_REG_4__0_ , P2_INSTQUEUE_REG_3__7_ , P2_INSTQUEUE_REG_3__6_ , P2_INSTQUEUE_REG_3__5_ , P2_INSTQUEUE_REG_3__4_ ,
             P2_INSTQUEUE_REG_3__3_ , P2_INSTQUEUE_REG_3__2_ , P2_INSTQUEUE_REG_3__1_ , P2_INSTQUEUE_REG_3__0_ , P2_INSTQUEUE_REG_2__7_ , P2_INSTQUEUE_REG_2__6_ ,
             P2_INSTQUEUE_REG_2__5_ , P2_INSTQUEUE_REG_2__4_ , P2_INSTQUEUE_REG_2__3_ , P2_INSTQUEUE_REG_2__2_ , P2_INSTQUEUE_REG_2__1_ , P2_INSTQUEUE_REG_2__0_ ,
             P2_INSTQUEUE_REG_1__7_ , P2_INSTQUEUE_REG_1__6_ , P2_INSTQUEUE_REG_1__5_ , P2_INSTQUEUE_REG_1__4_ , P2_INSTQUEUE_REG_1__3_ , P2_INSTQUEUE_REG_1__2_ ,
             P2_INSTQUEUE_REG_1__1_ , P2_INSTQUEUE_REG_1__0_ , P2_INSTQUEUE_REG_0__7_ , P2_INSTQUEUE_REG_0__6_ , P2_INSTQUEUE_REG_0__5_ , P2_INSTQUEUE_REG_0__4_ ,
             P2_INSTQUEUE_REG_0__3_ , P2_INSTQUEUE_REG_0__2_ , P2_INSTQUEUE_REG_0__1_ , P2_INSTQUEUE_REG_0__0_ , P2_INSTQUEUERD_ADDR_REG_4_ , P2_INSTQUEUERD_ADDR_REG_3_ ,
             P2_INSTQUEUERD_ADDR_REG_2_ , P2_INSTQUEUERD_ADDR_REG_1_ , P2_INSTQUEUERD_ADDR_REG_0_ , P2_INSTQUEUEWR_ADDR_REG_4_ , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_INSTQUEUEWR_ADDR_REG_2_ ,
             P2_INSTQUEUEWR_ADDR_REG_1_ , P2_INSTQUEUEWR_ADDR_REG_0_ , P2_INSTADDRPOINTER_REG_0_ , P2_INSTADDRPOINTER_REG_1_ , P2_INSTADDRPOINTER_REG_2_ , P2_INSTADDRPOINTER_REG_3_ ,
             P2_INSTADDRPOINTER_REG_4_ , P2_INSTADDRPOINTER_REG_5_ , P2_INSTADDRPOINTER_REG_6_ , P2_INSTADDRPOINTER_REG_7_ , P2_INSTADDRPOINTER_REG_8_ , P2_INSTADDRPOINTER_REG_9_ ,
             P2_INSTADDRPOINTER_REG_10_ , P2_INSTADDRPOINTER_REG_11_ , P2_INSTADDRPOINTER_REG_12_ , P2_INSTADDRPOINTER_REG_13_ , P2_INSTADDRPOINTER_REG_14_ , P2_INSTADDRPOINTER_REG_15_ ,
             P2_INSTADDRPOINTER_REG_16_ , P2_INSTADDRPOINTER_REG_17_ , P2_INSTADDRPOINTER_REG_18_ , P2_INSTADDRPOINTER_REG_19_ , P2_INSTADDRPOINTER_REG_20_ , P2_INSTADDRPOINTER_REG_21_ ,
             P2_INSTADDRPOINTER_REG_22_ , P2_INSTADDRPOINTER_REG_23_ , P2_INSTADDRPOINTER_REG_24_ , P2_INSTADDRPOINTER_REG_25_ , P2_INSTADDRPOINTER_REG_26_ , P2_INSTADDRPOINTER_REG_27_ ,
             P2_INSTADDRPOINTER_REG_28_ , P2_INSTADDRPOINTER_REG_29_ , P2_INSTADDRPOINTER_REG_30_ , P2_INSTADDRPOINTER_REG_31_ , P2_PHYADDRPOINTER_REG_0_ , P2_PHYADDRPOINTER_REG_1_ ,
             P2_PHYADDRPOINTER_REG_2_ , P2_PHYADDRPOINTER_REG_3_ , P2_PHYADDRPOINTER_REG_4_ , P2_PHYADDRPOINTER_REG_5_ , P2_PHYADDRPOINTER_REG_6_ , P2_PHYADDRPOINTER_REG_7_ ,
             P2_PHYADDRPOINTER_REG_8_ , P2_PHYADDRPOINTER_REG_9_ , P2_PHYADDRPOINTER_REG_10_ , P2_PHYADDRPOINTER_REG_11_ , P2_PHYADDRPOINTER_REG_12_ , P2_PHYADDRPOINTER_REG_13_ ,
             P2_PHYADDRPOINTER_REG_14_ , P2_PHYADDRPOINTER_REG_15_ , P2_PHYADDRPOINTER_REG_16_ , P2_PHYADDRPOINTER_REG_17_ , P2_PHYADDRPOINTER_REG_18_ , P2_PHYADDRPOINTER_REG_19_ ,
             P2_PHYADDRPOINTER_REG_20_ , P2_PHYADDRPOINTER_REG_21_ , P2_PHYADDRPOINTER_REG_22_ , P2_PHYADDRPOINTER_REG_23_ , P2_PHYADDRPOINTER_REG_24_ , P2_PHYADDRPOINTER_REG_25_ ,
             P2_PHYADDRPOINTER_REG_26_ , P2_PHYADDRPOINTER_REG_27_ , P2_PHYADDRPOINTER_REG_28_ , P2_PHYADDRPOINTER_REG_29_ , P2_PHYADDRPOINTER_REG_30_ , P2_PHYADDRPOINTER_REG_31_ ,
             P2_LWORD_REG_15_ , P2_LWORD_REG_14_ , P2_LWORD_REG_13_ , P2_LWORD_REG_12_ , P2_LWORD_REG_11_ , P2_LWORD_REG_10_ ,
             P2_LWORD_REG_9_ , P2_LWORD_REG_8_ , P2_LWORD_REG_7_ , P2_LWORD_REG_6_ , P2_LWORD_REG_5_ , P2_LWORD_REG_4_ ,
             P2_LWORD_REG_3_ , P2_LWORD_REG_2_ , P2_LWORD_REG_1_ , P2_LWORD_REG_0_ , P2_UWORD_REG_14_ , P2_UWORD_REG_13_ ,
             P2_UWORD_REG_12_ , P2_UWORD_REG_11_ , P2_UWORD_REG_10_ , P2_UWORD_REG_9_ , P2_UWORD_REG_8_ , P2_UWORD_REG_7_ ,
             P2_UWORD_REG_6_ , P2_UWORD_REG_5_ , P2_UWORD_REG_4_ , P2_UWORD_REG_3_ , P2_UWORD_REG_2_ , P2_UWORD_REG_1_ ,
             P2_UWORD_REG_0_ , P2_DATAO_REG_0_ , P2_DATAO_REG_1_ , P2_DATAO_REG_2_ , P2_DATAO_REG_3_ , P2_DATAO_REG_4_ ,
             P2_DATAO_REG_5_ , P2_DATAO_REG_6_ , P2_DATAO_REG_7_ , P2_DATAO_REG_8_ , P2_DATAO_REG_9_ , P2_DATAO_REG_10_ ,
             P2_DATAO_REG_11_ , P2_DATAO_REG_12_ , P2_DATAO_REG_13_ , P2_DATAO_REG_14_ , P2_DATAO_REG_15_ , P2_DATAO_REG_16_ ,
             P2_DATAO_REG_17_ , P2_DATAO_REG_18_ , P2_DATAO_REG_19_ , P2_DATAO_REG_20_ , P2_DATAO_REG_21_ , P2_DATAO_REG_22_ ,
             P2_DATAO_REG_23_ , P2_DATAO_REG_24_ , P2_DATAO_REG_25_ , P2_DATAO_REG_26_ , P2_DATAO_REG_27_ , P2_DATAO_REG_28_ ,
             P2_DATAO_REG_29_ , P2_DATAO_REG_30_ , P2_DATAO_REG_31_ , P2_EAX_REG_0_ , P2_EAX_REG_1_ , P2_EAX_REG_2_ ,
             P2_EAX_REG_3_ , P2_EAX_REG_4_ , P2_EAX_REG_5_ , P2_EAX_REG_6_ , P2_EAX_REG_7_ , P2_EAX_REG_8_ ,
             P2_EAX_REG_9_ , P2_EAX_REG_10_ , P2_EAX_REG_11_ , P2_EAX_REG_12_ , P2_EAX_REG_13_ , P2_EAX_REG_14_ ,
             P2_EAX_REG_15_ , P2_EAX_REG_16_ , P2_EAX_REG_17_ , P2_EAX_REG_18_ , P2_EAX_REG_19_ , P2_EAX_REG_20_ ,
             P2_EAX_REG_21_ , P2_EAX_REG_22_ , P2_EAX_REG_23_ , P2_EAX_REG_24_ , P2_EAX_REG_25_ , P2_EAX_REG_26_ ,
             P2_EAX_REG_27_ , P2_EAX_REG_28_ , P2_EAX_REG_29_ , P2_EAX_REG_30_ , P2_EAX_REG_31_ , P2_EBX_REG_0_ ,
             P2_EBX_REG_1_ , P2_EBX_REG_2_ , P2_EBX_REG_3_ , P2_EBX_REG_4_ , P2_EBX_REG_5_ , P2_EBX_REG_6_ ,
             P2_EBX_REG_7_ , P2_EBX_REG_8_ , P2_EBX_REG_9_ , P2_EBX_REG_10_ , P2_EBX_REG_11_ , P2_EBX_REG_12_ ,
             P2_EBX_REG_13_ , P2_EBX_REG_14_ , P2_EBX_REG_15_ , P2_EBX_REG_16_ , P2_EBX_REG_17_ , P2_EBX_REG_18_ ,
             P2_EBX_REG_19_ , P2_EBX_REG_20_ , P2_EBX_REG_21_ , P2_EBX_REG_22_ , P2_EBX_REG_23_ , P2_EBX_REG_24_ ,
             P2_EBX_REG_25_ , P2_EBX_REG_26_ , P2_EBX_REG_27_ , P2_EBX_REG_28_ , P2_EBX_REG_29_ , P2_EBX_REG_30_ ,
             P2_EBX_REG_31_ , P2_REIP_REG_0_ , P2_REIP_REG_1_ , P2_REIP_REG_2_ , P2_REIP_REG_3_ , P2_REIP_REG_4_ ,
             P2_REIP_REG_5_ , P2_REIP_REG_6_ , P2_REIP_REG_7_ , P2_REIP_REG_8_ , P2_REIP_REG_9_ , P2_REIP_REG_10_ ,
             P2_REIP_REG_11_ , P2_REIP_REG_12_ , P2_REIP_REG_13_ , P2_REIP_REG_14_ , P2_REIP_REG_15_ , P2_REIP_REG_16_ ,
             P2_REIP_REG_17_ , P2_REIP_REG_18_ , P2_REIP_REG_19_ , P2_REIP_REG_20_ , P2_REIP_REG_21_ , P2_REIP_REG_22_ ,
             P2_REIP_REG_23_ , P2_REIP_REG_24_ , P2_REIP_REG_25_ , P2_REIP_REG_26_ , P2_REIP_REG_27_ , P2_REIP_REG_28_ ,
             P2_REIP_REG_29_ , P2_REIP_REG_30_ , P2_REIP_REG_31_ , P2_BYTEENABLE_REG_3_ , P2_BYTEENABLE_REG_2_ , P2_BYTEENABLE_REG_1_ ,
             P2_BYTEENABLE_REG_0_ , P2_W_R_N_REG , P2_FLUSH_REG , P2_MORE_REG , P2_STATEBS16_REG , P2_REQUESTPENDING_REG ,
             P2_D_C_N_REG , P2_M_IO_N_REG , P2_CODEFETCH_REG , P2_ADS_N_REG , P2_READREQUEST_REG , P2_MEMORYFETCH_REG ,
             P1_BE_N_REG_3_ , P1_BE_N_REG_2_ , P1_BE_N_REG_1_ , P1_BE_N_REG_0_ , P1_ADDRESS_REG_29__EXTRA , P1_ADDRESS_REG_28__EXTRA ,
             P1_ADDRESS_REG_27__EXTRA , P1_ADDRESS_REG_26__EXTRA , P1_ADDRESS_REG_25__EXTRA , P1_ADDRESS_REG_24__EXTRA , P1_ADDRESS_REG_23__EXTRA , P1_ADDRESS_REG_22__EXTRA ,
             P1_ADDRESS_REG_21__EXTRA , P1_ADDRESS_REG_20__EXTRA , P1_ADDRESS_REG_19__EXTRA , P1_ADDRESS_REG_18__EXTRA , P1_ADDRESS_REG_17__EXTRA , P1_ADDRESS_REG_16__EXTRA ,
             P1_ADDRESS_REG_15__EXTRA , P1_ADDRESS_REG_14__EXTRA , P1_ADDRESS_REG_13__EXTRA , P1_ADDRESS_REG_12__EXTRA , P1_ADDRESS_REG_11__EXTRA , P1_ADDRESS_REG_10__EXTRA ,
             P1_ADDRESS_REG_9__EXTRA , P1_ADDRESS_REG_8__EXTRA , P1_ADDRESS_REG_7__EXTRA , P1_ADDRESS_REG_6__EXTRA , P1_ADDRESS_REG_5__EXTRA , P1_ADDRESS_REG_4__EXTRA ,
             P1_ADDRESS_REG_3__EXTRA , P1_ADDRESS_REG_2__EXTRA , P1_ADDRESS_REG_1__EXTRA , P1_ADDRESS_REG_0__EXTRA , P1_STATE_REG_2_ , P1_STATE_REG_1_ ,
             P1_STATE_REG_0_ , P1_DATAWIDTH_REG_0_ , P1_DATAWIDTH_REG_1_ , P1_DATAWIDTH_REG_2_ , P1_DATAWIDTH_REG_3_ , P1_DATAWIDTH_REG_4_ ,
             P1_DATAWIDTH_REG_5_ , P1_DATAWIDTH_REG_6_ , P1_DATAWIDTH_REG_7_ , P1_DATAWIDTH_REG_8_ , P1_DATAWIDTH_REG_9_ , P1_DATAWIDTH_REG_10_ ,
             P1_DATAWIDTH_REG_11_ , P1_DATAWIDTH_REG_12_ , P1_DATAWIDTH_REG_13_ , P1_DATAWIDTH_REG_14_ , P1_DATAWIDTH_REG_15_ , P1_DATAWIDTH_REG_16_ ,
             P1_DATAWIDTH_REG_17_ , P1_DATAWIDTH_REG_18_ , P1_DATAWIDTH_REG_19_ , P1_DATAWIDTH_REG_20_ , P1_DATAWIDTH_REG_21_ , P1_DATAWIDTH_REG_22_ ,
             P1_DATAWIDTH_REG_23_ , P1_DATAWIDTH_REG_24_ , P1_DATAWIDTH_REG_25_ , P1_DATAWIDTH_REG_26_ , P1_DATAWIDTH_REG_27_ , P1_DATAWIDTH_REG_28_ ,
             P1_DATAWIDTH_REG_29_ , P1_DATAWIDTH_REG_30_ , P1_DATAWIDTH_REG_31_ , P1_STATE2_REG_3_ , P1_STATE2_REG_2_ , P1_STATE2_REG_1_ ,
             P1_STATE2_REG_0_ , P1_INSTQUEUE_REG_15__7_ , P1_INSTQUEUE_REG_15__6_ , P1_INSTQUEUE_REG_15__5_ , P1_INSTQUEUE_REG_15__4_ , P1_INSTQUEUE_REG_15__3_ ,
             P1_INSTQUEUE_REG_15__2_ , P1_INSTQUEUE_REG_15__1_ , P1_INSTQUEUE_REG_15__0_ , P1_INSTQUEUE_REG_14__7_ , P1_INSTQUEUE_REG_14__6_ , P1_INSTQUEUE_REG_14__5_ ,
             P1_INSTQUEUE_REG_14__4_ , P1_INSTQUEUE_REG_14__3_ , P1_INSTQUEUE_REG_14__2_ , P1_INSTQUEUE_REG_14__1_ , P1_INSTQUEUE_REG_14__0_ , P1_INSTQUEUE_REG_13__7_ ,
             P1_INSTQUEUE_REG_13__6_ , P1_INSTQUEUE_REG_13__5_ , P1_INSTQUEUE_REG_13__4_ , P1_INSTQUEUE_REG_13__3_ , P1_INSTQUEUE_REG_13__2_ , P1_INSTQUEUE_REG_13__1_ ,
             P1_INSTQUEUE_REG_13__0_ , P1_INSTQUEUE_REG_12__7_ , P1_INSTQUEUE_REG_12__6_ , P1_INSTQUEUE_REG_12__5_ , P1_INSTQUEUE_REG_12__4_ , P1_INSTQUEUE_REG_12__3_ ,
             P1_INSTQUEUE_REG_12__2_ , P1_INSTQUEUE_REG_12__1_ , P1_INSTQUEUE_REG_12__0_ , P1_INSTQUEUE_REG_11__7_ , P1_INSTQUEUE_REG_11__6_ , P1_INSTQUEUE_REG_11__5_ ,
             P1_INSTQUEUE_REG_11__4_ , P1_INSTQUEUE_REG_11__3_ , P1_INSTQUEUE_REG_11__2_ , P1_INSTQUEUE_REG_11__1_ , P1_INSTQUEUE_REG_11__0_ , P1_INSTQUEUE_REG_10__7_ ,
             P1_INSTQUEUE_REG_10__6_ , P1_INSTQUEUE_REG_10__5_ , P1_INSTQUEUE_REG_10__4_ , P1_INSTQUEUE_REG_10__3_ , P1_INSTQUEUE_REG_10__2_ , P1_INSTQUEUE_REG_10__1_ ,
             P1_INSTQUEUE_REG_10__0_ , P1_INSTQUEUE_REG_9__7_ , P1_INSTQUEUE_REG_9__6_ , P1_INSTQUEUE_REG_9__5_ , P1_INSTQUEUE_REG_9__4_ , P1_INSTQUEUE_REG_9__3_ ,
             P1_INSTQUEUE_REG_9__2_ , P1_INSTQUEUE_REG_9__1_ , P1_INSTQUEUE_REG_9__0_ , P1_INSTQUEUE_REG_8__7_ , P1_INSTQUEUE_REG_8__6_ , P1_INSTQUEUE_REG_8__5_ ,
             P1_INSTQUEUE_REG_8__4_ , P1_INSTQUEUE_REG_8__3_ , P1_INSTQUEUE_REG_8__2_ , P1_INSTQUEUE_REG_8__1_ , P1_INSTQUEUE_REG_8__0_ , P1_INSTQUEUE_REG_7__7_ ,
             P1_INSTQUEUE_REG_7__6_ , P1_INSTQUEUE_REG_7__5_ , P1_INSTQUEUE_REG_7__4_ , P1_INSTQUEUE_REG_7__3_ , P1_INSTQUEUE_REG_7__2_ , P1_INSTQUEUE_REG_7__1_ ,
             P1_INSTQUEUE_REG_7__0_ , P1_INSTQUEUE_REG_6__7_ , P1_INSTQUEUE_REG_6__6_ , P1_INSTQUEUE_REG_6__5_ , P1_INSTQUEUE_REG_6__4_ , P1_INSTQUEUE_REG_6__3_ ,
             P1_INSTQUEUE_REG_6__2_ , P1_INSTQUEUE_REG_6__1_ , P1_INSTQUEUE_REG_6__0_ , P1_INSTQUEUE_REG_5__7_ , P1_INSTQUEUE_REG_5__6_ , P1_INSTQUEUE_REG_5__5_ ,
             P1_INSTQUEUE_REG_5__4_ , P1_INSTQUEUE_REG_5__3_ , P1_INSTQUEUE_REG_5__2_ , P1_INSTQUEUE_REG_5__1_ , P1_INSTQUEUE_REG_5__0_ , P1_INSTQUEUE_REG_4__7_ ,
             P1_INSTQUEUE_REG_4__6_ , P1_INSTQUEUE_REG_4__5_ , P1_INSTQUEUE_REG_4__4_ , P1_INSTQUEUE_REG_4__3_ , P1_INSTQUEUE_REG_4__2_ , P1_INSTQUEUE_REG_4__1_ ,
             P1_INSTQUEUE_REG_4__0_ , P1_INSTQUEUE_REG_3__7_ , P1_INSTQUEUE_REG_3__6_ , P1_INSTQUEUE_REG_3__5_ , P1_INSTQUEUE_REG_3__4_ , P1_INSTQUEUE_REG_3__3_ ,
             P1_INSTQUEUE_REG_3__2_ , P1_INSTQUEUE_REG_3__1_ , P1_INSTQUEUE_REG_3__0_ , P1_INSTQUEUE_REG_2__7_ , P1_INSTQUEUE_REG_2__6_ , P1_INSTQUEUE_REG_2__5_ ,
             P1_INSTQUEUE_REG_2__4_ , P1_INSTQUEUE_REG_2__3_ , P1_INSTQUEUE_REG_2__2_ , P1_INSTQUEUE_REG_2__1_ , P1_INSTQUEUE_REG_2__0_ , P1_INSTQUEUE_REG_1__7_ ,
             P1_INSTQUEUE_REG_1__6_ , P1_INSTQUEUE_REG_1__5_ , P1_INSTQUEUE_REG_1__4_ , P1_INSTQUEUE_REG_1__3_ , P1_INSTQUEUE_REG_1__2_ , P1_INSTQUEUE_REG_1__1_ ,
             P1_INSTQUEUE_REG_1__0_ , P1_INSTQUEUE_REG_0__7_ , P1_INSTQUEUE_REG_0__6_ , P1_INSTQUEUE_REG_0__5_ , P1_INSTQUEUE_REG_0__4_ , P1_INSTQUEUE_REG_0__3_ ,
             P1_INSTQUEUE_REG_0__2_ , P1_INSTQUEUE_REG_0__1_ , P1_INSTQUEUE_REG_0__0_ , P1_INSTQUEUERD_ADDR_REG_4_ , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_2_ ,
             P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUEWR_ADDR_REG_4_ , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_INSTQUEUEWR_ADDR_REG_1_ ,
             P1_INSTQUEUEWR_ADDR_REG_0_ , P1_INSTADDRPOINTER_REG_0_ , P1_INSTADDRPOINTER_REG_1_ , P1_INSTADDRPOINTER_REG_2_ , P1_INSTADDRPOINTER_REG_3_ , P1_INSTADDRPOINTER_REG_4_ ,
             P1_INSTADDRPOINTER_REG_5_ , P1_INSTADDRPOINTER_REG_6_ , P1_INSTADDRPOINTER_REG_7_ , P1_INSTADDRPOINTER_REG_8_ , P1_INSTADDRPOINTER_REG_9_ , P1_INSTADDRPOINTER_REG_10_ ,
             P1_INSTADDRPOINTER_REG_11_ , P1_INSTADDRPOINTER_REG_12_ , P1_INSTADDRPOINTER_REG_13_ , P1_INSTADDRPOINTER_REG_14_ , P1_INSTADDRPOINTER_REG_15_ , P1_INSTADDRPOINTER_REG_16_ ,
             P1_INSTADDRPOINTER_REG_17_ , P1_INSTADDRPOINTER_REG_18_ , P1_INSTADDRPOINTER_REG_19_ , P1_INSTADDRPOINTER_REG_20_ , P1_INSTADDRPOINTER_REG_21_ , P1_INSTADDRPOINTER_REG_22_ ,
             P1_INSTADDRPOINTER_REG_23_ , P1_INSTADDRPOINTER_REG_24_ , P1_INSTADDRPOINTER_REG_25_ , P1_INSTADDRPOINTER_REG_26_ , P1_INSTADDRPOINTER_REG_27_ , P1_INSTADDRPOINTER_REG_28_ ,
             P1_INSTADDRPOINTER_REG_29_ , P1_INSTADDRPOINTER_REG_30_ , P1_INSTADDRPOINTER_REG_31_ , P1_PHYADDRPOINTER_REG_0_ , P1_PHYADDRPOINTER_REG_1_ , P1_PHYADDRPOINTER_REG_2_ ,
             P1_PHYADDRPOINTER_REG_3_ , P1_PHYADDRPOINTER_REG_4_ , P1_PHYADDRPOINTER_REG_5_ , P1_PHYADDRPOINTER_REG_6_ , P1_PHYADDRPOINTER_REG_7_ , P1_PHYADDRPOINTER_REG_8_ ,
             P1_PHYADDRPOINTER_REG_9_ , P1_PHYADDRPOINTER_REG_10_ , P1_PHYADDRPOINTER_REG_11_ , P1_PHYADDRPOINTER_REG_12_ , P1_PHYADDRPOINTER_REG_13_ , P1_PHYADDRPOINTER_REG_14_ ,
             P1_PHYADDRPOINTER_REG_15_ , P1_PHYADDRPOINTER_REG_16_ , P1_PHYADDRPOINTER_REG_17_ , P1_PHYADDRPOINTER_REG_18_ , P1_PHYADDRPOINTER_REG_19_ , P1_PHYADDRPOINTER_REG_20_ ,
             P1_PHYADDRPOINTER_REG_21_ , P1_PHYADDRPOINTER_REG_22_ , P1_PHYADDRPOINTER_REG_23_ , P1_PHYADDRPOINTER_REG_24_ , P1_PHYADDRPOINTER_REG_25_ , P1_PHYADDRPOINTER_REG_26_ ,
             P1_PHYADDRPOINTER_REG_27_ , P1_PHYADDRPOINTER_REG_28_ , P1_PHYADDRPOINTER_REG_29_ , P1_PHYADDRPOINTER_REG_30_ , P1_PHYADDRPOINTER_REG_31_ , P1_LWORD_REG_15_ ,
             P1_LWORD_REG_14_ , P1_LWORD_REG_13_ , P1_LWORD_REG_12_ , P1_LWORD_REG_11_ , P1_LWORD_REG_10_ , P1_LWORD_REG_9_ ,
             P1_LWORD_REG_8_ , P1_LWORD_REG_7_ , P1_LWORD_REG_6_ , P1_LWORD_REG_5_ , P1_LWORD_REG_4_ , P1_LWORD_REG_3_ ,
             P1_LWORD_REG_2_ , P1_LWORD_REG_1_ , P1_LWORD_REG_0_ , P1_UWORD_REG_14_ , P1_UWORD_REG_13_ , P1_UWORD_REG_12_ ,
             P1_UWORD_REG_11_ , P1_UWORD_REG_10_ , P1_UWORD_REG_9_ , P1_UWORD_REG_8_ , P1_UWORD_REG_7_ , P1_UWORD_REG_6_ ,
             P1_UWORD_REG_5_ , P1_UWORD_REG_4_ , P1_UWORD_REG_3_ , P1_UWORD_REG_2_ , P1_UWORD_REG_1_ , P1_UWORD_REG_0_ ,
             P1_DATAO_REG_0_ , P1_DATAO_REG_1_ , P1_DATAO_REG_2_ , P1_DATAO_REG_3_ , P1_DATAO_REG_4_ , P1_DATAO_REG_5_ ,
             P1_DATAO_REG_6_ , P1_DATAO_REG_7_ , P1_DATAO_REG_8_ , P1_DATAO_REG_9_ , P1_DATAO_REG_10_ , P1_DATAO_REG_11_ ,
             P1_DATAO_REG_12_ , P1_DATAO_REG_13_ , P1_DATAO_REG_14_ , P1_DATAO_REG_15_ , P1_DATAO_REG_16_ , P1_DATAO_REG_17_ ,
             P1_DATAO_REG_18_ , P1_DATAO_REG_19_ , P1_DATAO_REG_20_ , P1_DATAO_REG_21_ , P1_DATAO_REG_22_ , P1_DATAO_REG_23_ ,
             P1_DATAO_REG_24_ , P1_DATAO_REG_25_ , P1_DATAO_REG_26_ , P1_DATAO_REG_27_ , P1_DATAO_REG_28_ , P1_DATAO_REG_29_ ,
             P1_DATAO_REG_30_ , P1_DATAO_REG_31_ , P1_EAX_REG_0_ , P1_EAX_REG_1_ , P1_EAX_REG_2_ , P1_EAX_REG_3_ ,
             P1_EAX_REG_4_ , P1_EAX_REG_5_ , P1_EAX_REG_6_ , P1_EAX_REG_7_ , P1_EAX_REG_8_ , P1_EAX_REG_9_ ,
             P1_EAX_REG_10_ , P1_EAX_REG_11_ , P1_EAX_REG_12_ , P1_EAX_REG_13_ , P1_EAX_REG_14_ , P1_EAX_REG_15_ ,
             P1_EAX_REG_16_ , P1_EAX_REG_17_ , P1_EAX_REG_18_ , P1_EAX_REG_19_ , P1_EAX_REG_20_ , P1_EAX_REG_21_ ,
             P1_EAX_REG_22_ , P1_EAX_REG_23_ , P1_EAX_REG_24_ , P1_EAX_REG_25_ , P1_EAX_REG_26_ , P1_EAX_REG_27_ ,
             P1_EAX_REG_28_ , P1_EAX_REG_29_ , P1_EAX_REG_30_ , P1_EAX_REG_31_ , P1_EBX_REG_0_ , P1_EBX_REG_1_ ,
             P1_EBX_REG_2_ , P1_EBX_REG_3_ , P1_EBX_REG_4_ , P1_EBX_REG_5_ , P1_EBX_REG_6_ , P1_EBX_REG_7_ ,
             P1_EBX_REG_8_ , P1_EBX_REG_9_ , P1_EBX_REG_10_ , P1_EBX_REG_11_ , P1_EBX_REG_12_ , P1_EBX_REG_13_ ,
             P1_EBX_REG_14_ , P1_EBX_REG_15_ , P1_EBX_REG_16_ , P1_EBX_REG_17_ , P1_EBX_REG_18_ , P1_EBX_REG_19_ ,
             P1_EBX_REG_20_ , P1_EBX_REG_21_ , P1_EBX_REG_22_ , P1_EBX_REG_23_ , P1_EBX_REG_24_ , P1_EBX_REG_25_ ,
             P1_EBX_REG_26_ , P1_EBX_REG_27_ , P1_EBX_REG_28_ , P1_EBX_REG_29_ , P1_EBX_REG_30_ , P1_EBX_REG_31_ ,
             P1_REIP_REG_0_ , P1_REIP_REG_1_ , P1_REIP_REG_2_ , P1_REIP_REG_3_ , P1_REIP_REG_4_ , P1_REIP_REG_5_ ,
             P1_REIP_REG_6_ , P1_REIP_REG_7_ , P1_REIP_REG_8_ , P1_REIP_REG_9_ , P1_REIP_REG_10_ , P1_REIP_REG_11_ ,
             P1_REIP_REG_12_ , P1_REIP_REG_13_ , P1_REIP_REG_14_ , P1_REIP_REG_15_ , P1_REIP_REG_16_ , P1_REIP_REG_17_ ,
             P1_REIP_REG_18_ , P1_REIP_REG_19_ , P1_REIP_REG_20_ , P1_REIP_REG_21_ , P1_REIP_REG_22_ , P1_REIP_REG_23_ ,
             P1_REIP_REG_24_ , P1_REIP_REG_25_ , P1_REIP_REG_26_ , P1_REIP_REG_27_ , P1_REIP_REG_28_ , P1_REIP_REG_29_ ,
             P1_REIP_REG_30_ , P1_REIP_REG_31_ , P1_BYTEENABLE_REG_3_ , P1_BYTEENABLE_REG_2_ , P1_BYTEENABLE_REG_1_ , P1_BYTEENABLE_REG_0_ ,
             P1_W_R_N_REG , P1_FLUSH_REG , P1_MORE_REG , P1_STATEBS16_REG , P1_REQUESTPENDING_REG , P1_D_C_N_REG ,
             P1_M_IO_N_REG , P1_CODEFETCH_REG , P1_ADS_N_REG_EXTRA , P1_READREQUEST_REG , P1_MEMORYFETCH_REG , DATAI_31_ ,
             DATAI_30_ , DATAI_29_ , DATAI_28_ , DATAI_27_ , DATAI_26_ , DATAI_25_ ,
             DATAI_24_ , DATAI_23_ , DATAI_22_ , DATAI_21_ , DATAI_20_ , DATAI_19_ ,
             DATAI_18_ , DATAI_17_ , DATAI_16_ , DATAI_15_ , DATAI_14_ , DATAI_13_ ,
             DATAI_12_ , DATAI_11_ , DATAI_10_ , DATAI_9_ , DATAI_8_ , DATAI_7_ ,
             DATAI_6_ , DATAI_5_ , DATAI_4_ , DATAI_3_ , DATAI_2_ , DATAI_1_ ,
             DATAI_0_ , HOLD , NA , BS16 , READY1 , READY2 );

output P3_DATAO_REG_31_ , P3_DATAO_REG_30_ , P3_DATAO_REG_29_ , P3_DATAO_REG_28_ , P3_DATAO_REG_27_ , P3_DATAO_REG_26_;
output P3_DATAO_REG_25_ , P3_DATAO_REG_24_ , P3_DATAO_REG_23_ , P3_DATAO_REG_22_ , P3_DATAO_REG_21_ , P3_DATAO_REG_20_;
output P3_DATAO_REG_19_ , P3_DATAO_REG_18_ , P3_DATAO_REG_17_ , P3_DATAO_REG_16_ , P3_DATAO_REG_15_ , P3_DATAO_REG_14_;
output P3_DATAO_REG_13_ , P3_DATAO_REG_12_ , P3_DATAO_REG_11_ , P3_DATAO_REG_10_ , P3_DATAO_REG_9_ , P3_DATAO_REG_8_;
output P3_DATAO_REG_7_ , P3_DATAO_REG_6_ , P3_DATAO_REG_5_ , P3_DATAO_REG_4_ , P3_DATAO_REG_3_ , P3_DATAO_REG_2_;
output P3_DATAO_REG_1_ , P3_DATAO_REG_0_ , P1_ADDRESS_REG_29_ , P1_ADDRESS_REG_28_ , P1_ADDRESS_REG_27_ , P1_ADDRESS_REG_26_;
output P1_ADDRESS_REG_25_ , P1_ADDRESS_REG_24_ , P1_ADDRESS_REG_23_ , P1_ADDRESS_REG_22_ , P1_ADDRESS_REG_21_ , P1_ADDRESS_REG_20_;
output P1_ADDRESS_REG_19_ , P1_ADDRESS_REG_18_ , P1_ADDRESS_REG_17_ , P1_ADDRESS_REG_16_ , P1_ADDRESS_REG_15_ , P1_ADDRESS_REG_14_;
output P1_ADDRESS_REG_13_ , P1_ADDRESS_REG_12_ , P1_ADDRESS_REG_11_ , P1_ADDRESS_REG_10_ , P1_ADDRESS_REG_9_ , P1_ADDRESS_REG_8_;
output P1_ADDRESS_REG_7_ , P1_ADDRESS_REG_6_ , P1_ADDRESS_REG_5_ , P1_ADDRESS_REG_4_ , P1_ADDRESS_REG_3_ , P1_ADDRESS_REG_2_;
output P1_ADDRESS_REG_1_ , P1_ADDRESS_REG_0_ , U355 , U356 , U357 , U358;
output U359 , U360 , U361 , U362 , U363 , U364;
output U366 , U367 , U368 , U369 , U370 , U371;
output U372 , U373 , U374 , U375 , U347 , U348;
output U349 , U350 , U351 , U352 , U353 , U354;
output U365 , U376 , P3_W_R_N_REG , P3_D_C_N_REG , P3_M_IO_N_REG , P1_ADS_N_REG;
output P3_ADS_N_REG;
output U247 , U246 , U245 , U244 , U243 , U242 , U241;
output U240 , U239 , U238 , U237 , U236 , U235 , U234;
output U233 , U232 , U231 , U230 , U229 , U228 , U227;
output U226 , U225 , U224 , U223 , U222 , U221 , U220;
output U219 , U218 , U217 , U216 , U251 , U252 , U253;
output U254 , U255 , U256 , U257 , U258 , U259 , U260;
output U261 , U262 , U263 , U264 , U265 , U266 , U267;
output U268 , U269 , U270 , U271 , U272 , U273 , U274;
output U275 , U276 , U277 , U278 , U279 , U280 , U281;
output U282 , U212 , U215 , U213 , U214 , P3_U3274 , P3_U3275;
output P3_U3276 , P3_U3277 , P3_U3061 , P3_U3060 , P3_U3059 , P3_U3058 , P3_U3057;
output P3_U3056 , P3_U3055 , P3_U3054 , P3_U3053 , P3_U3052 , P3_U3051 , P3_U3050;
output P3_U3049 , P3_U3048 , P3_U3047 , P3_U3046 , P3_U3045 , P3_U3044 , P3_U3043;
output P3_U3042 , P3_U3041 , P3_U3040 , P3_U3039 , P3_U3038 , P3_U3037 , P3_U3036;
output P3_U3035 , P3_U3034 , P3_U3033 , P3_U3032 , P3_U3031 , P3_U3030 , P3_U3029;
output P3_U3280 , P3_U3281 , P3_U3028 , P3_U3027 , P3_U3026 , P3_U3025 , P3_U3024;
output P3_U3023 , P3_U3022 , P3_U3021 , P3_U3020 , P3_U3019 , P3_U3018 , P3_U3017;
output P3_U3016 , P3_U3015 , P3_U3014 , P3_U3013 , P3_U3012 , P3_U3011 , P3_U3010;
output P3_U3009 , P3_U3008 , P3_U3007 , P3_U3006 , P3_U3005 , P3_U3004 , P3_U3003;
output P3_U3002 , P3_U3001 , P3_U3000 , P3_U2999 , P3_U3282 , P3_U2998 , P3_U2997;
output P3_U2996 , P3_U2995 , P3_U2994 , P3_U2993 , P3_U2992 , P3_U2991 , P3_U2990;
output P3_U2989 , P3_U2988 , P3_U2987 , P3_U2986 , P3_U2985 , P3_U2984 , P3_U2983;
output P3_U2982 , P3_U2981 , P3_U2980 , P3_U2979 , P3_U2978 , P3_U2977 , P3_U2976;
output P3_U2975 , P3_U2974 , P3_U2973 , P3_U2972 , P3_U2971 , P3_U2970 , P3_U2969;
output P3_U2968 , P3_U2967 , P3_U2966 , P3_U2965 , P3_U2964 , P3_U2963 , P3_U2962;
output P3_U2961 , P3_U2960 , P3_U2959 , P3_U2958 , P3_U2957 , P3_U2956 , P3_U2955;
output P3_U2954 , P3_U2953 , P3_U2952 , P3_U2951 , P3_U2950 , P3_U2949 , P3_U2948;
output P3_U2947 , P3_U2946 , P3_U2945 , P3_U2944 , P3_U2943 , P3_U2942 , P3_U2941;
output P3_U2940 , P3_U2939 , P3_U2938 , P3_U2937 , P3_U2936 , P3_U2935 , P3_U2934;
output P3_U2933 , P3_U2932 , P3_U2931 , P3_U2930 , P3_U2929 , P3_U2928 , P3_U2927;
output P3_U2926 , P3_U2925 , P3_U2924 , P3_U2923 , P3_U2922 , P3_U2921 , P3_U2920;
output P3_U2919 , P3_U2918 , P3_U2917 , P3_U2916 , P3_U2915 , P3_U2914 , P3_U2913;
output P3_U2912 , P3_U2911 , P3_U2910 , P3_U2909 , P3_U2908 , P3_U2907 , P3_U2906;
output P3_U2905 , P3_U2904 , P3_U2903 , P3_U2902 , P3_U2901 , P3_U2900 , P3_U2899;
output P3_U2898 , P3_U2897 , P3_U2896 , P3_U2895 , P3_U2894 , P3_U2893 , P3_U2892;
output P3_U2891 , P3_U2890 , P3_U2889 , P3_U2888 , P3_U2887 , P3_U2886 , P3_U2885;
output P3_U2884 , P3_U2883 , P3_U2882 , P3_U2881 , P3_U2880 , P3_U2879 , P3_U2878;
output P3_U2877 , P3_U2876 , P3_U2875 , P3_U2874 , P3_U2873 , P3_U2872 , P3_U2871;
output P3_U2870 , P3_U2869 , P3_U2868 , P3_U3284 , P3_U3285 , P3_U3288 , P3_U3289;
output P3_U3290 , P3_U2867 , P3_U2866 , P3_U2865 , P3_U2864 , P3_U2863 , P3_U2862;
output P3_U2861 , P3_U2860 , P3_U2859 , P3_U2858 , P3_U2857 , P3_U2856 , P3_U2855;
output P3_U2854 , P3_U2853 , P3_U2852 , P3_U2851 , P3_U2850 , P3_U2849 , P3_U2848;
output P3_U2847 , P3_U2846 , P3_U2845 , P3_U2844 , P3_U2843 , P3_U2842 , P3_U2841;
output P3_U2840 , P3_U2839 , P3_U2838 , P3_U2837 , P3_U2836 , P3_U2835 , P3_U2834;
output P3_U2833 , P3_U2832 , P3_U2831 , P3_U2830 , P3_U2829 , P3_U2828 , P3_U2827;
output P3_U2826 , P3_U2825 , P3_U2824 , P3_U2823 , P3_U2822 , P3_U2821 , P3_U2820;
output P3_U2819 , P3_U2818 , P3_U2817 , P3_U2816 , P3_U2815 , P3_U2814 , P3_U2813;
output P3_U2812 , P3_U2811 , P3_U2810 , P3_U2809 , P3_U2808 , P3_U2807 , P3_U2806;
output P3_U2805 , P3_U2804 , P3_U2803 , P3_U2802 , P3_U2801 , P3_U2800 , P3_U2799;
output P3_U2798 , P3_U2797 , P3_U2796 , P3_U2795 , P3_U2794 , P3_U2793 , P3_U2792;
output P3_U2791 , P3_U2790 , P3_U2789 , P3_U2788 , P3_U2787 , P3_U2786 , P3_U2785;
output P3_U2784 , P3_U2783 , P3_U2782 , P3_U2781 , P3_U2780 , P3_U2779 , P3_U2778;
output P3_U2777 , P3_U2776 , P3_U2775 , P3_U2774 , P3_U2773 , P3_U2772 , P3_U2771;
output P3_U2770 , P3_U2769 , P3_U2768 , P3_U2767 , P3_U2766 , P3_U2765 , P3_U2764;
output P3_U2763 , P3_U2762 , P3_U2761 , P3_U2760 , P3_U2759 , P3_U2758 , P3_U2757;
output P3_U2756 , P3_U2755 , P3_U2754 , P3_U2753 , P3_U2752 , P3_U2751 , P3_U2750;
output P3_U2749 , P3_U2748 , P3_U2747 , P3_U2746 , P3_U2745 , P3_U2744 , P3_U2743;
output P3_U2742 , P3_U2741 , P3_U2740 , P3_U2739 , P3_U2738 , P3_U2737 , P3_U2736;
output P3_U2735 , P3_U2734 , P3_U2733 , P3_U2732 , P3_U2731 , P3_U2730 , P3_U2729;
output P3_U2728 , P3_U2727 , P3_U2726 , P3_U2725 , P3_U2724 , P3_U2723 , P3_U2722;
output P3_U2721 , P3_U2720 , P3_U2719 , P3_U2718 , P3_U2717 , P3_U2716 , P3_U2715;
output P3_U2714 , P3_U2713 , P3_U2712 , P3_U2711 , P3_U2710 , P3_U2709 , P3_U2708;
output P3_U2707 , P3_U2706 , P3_U2705 , P3_U2704 , P3_U2703 , P3_U2702 , P3_U2701;
output P3_U2700 , P3_U2699 , P3_U2698 , P3_U2697 , P3_U2696 , P3_U2695 , P3_U2694;
output P3_U2693 , P3_U2692 , P3_U2691 , P3_U2690 , P3_U2689 , P3_U2688 , P3_U2687;
output P3_U2686 , P3_U2685 , P3_U2684 , P3_U2683 , P3_U2682 , P3_U2681 , P3_U2680;
output P3_U2679 , P3_U2678 , P3_U2677 , P3_U2676 , P3_U2675 , P3_U2674 , P3_U2673;
output P3_U2672 , P3_U2671 , P3_U2670 , P3_U2669 , P3_U2668 , P3_U2667 , P3_U2666;
output P3_U2665 , P3_U2664 , P3_U2663 , P3_U2662 , P3_U2661 , P3_U2660 , P3_U2659;
output P3_U2658 , P3_U2657 , P3_U2656 , P3_U2655 , P3_U2654 , P3_U2653 , P3_U2652;
output P3_U2651 , P3_U2650 , P3_U2649 , P3_U2648 , P3_U2647 , P3_U2646 , P3_U2645;
output P3_U2644 , P3_U2643 , P3_U2642 , P3_U2641 , P3_U2640 , P3_U2639 , P3_U3292;
output P3_U2638 , P3_U3293 , P3_U3294 , P3_U2637 , P3_U3295 , P3_U2636 , P3_U3296;
output P3_U2635 , P3_U3297 , P3_U2634 , P3_U2633 , P3_U3298 , P3_U3299 , P2_U3585;
output P2_U3586 , P2_U3587 , P2_U3588 , P2_U3241 , P2_U3240 , P2_U3239 , P2_U3238;
output P2_U3237 , P2_U3236 , P2_U3235 , P2_U3234 , P2_U3233 , P2_U3232 , P2_U3231;
output P2_U3230 , P2_U3229 , P2_U3228 , P2_U3227 , P2_U3226 , P2_U3225 , P2_U3224;
output P2_U3223 , P2_U3222 , P2_U3221 , P2_U3220 , P2_U3219 , P2_U3218 , P2_U3217;
output P2_U3216 , P2_U3215 , P2_U3214 , P2_U3213 , P2_U3212 , P2_U3211 , P2_U3210;
output P2_U3209 , P2_U3591 , P2_U3592 , P2_U3208 , P2_U3207 , P2_U3206 , P2_U3205;
output P2_U3204 , P2_U3203 , P2_U3202 , P2_U3201 , P2_U3200 , P2_U3199 , P2_U3198;
output P2_U3197 , P2_U3196 , P2_U3195 , P2_U3194 , P2_U3193 , P2_U3192 , P2_U3191;
output P2_U3190 , P2_U3189 , P2_U3188 , P2_U3187 , P2_U3186 , P2_U3185 , P2_U3184;
output P2_U3183 , P2_U3182 , P2_U3181 , P2_U3180 , P2_U3179 , P2_U3593 , P2_U3178;
output P2_U3177 , P2_U3176 , P2_U3175 , P2_U3174 , P2_U3173 , P2_U3172 , P2_U3171;
output P2_U3170 , P2_U3169 , P2_U3168 , P2_U3167 , P2_U3166 , P2_U3165 , P2_U3164;
output P2_U3163 , P2_U3162 , P2_U3161 , P2_U3160 , P2_U3159 , P2_U3158 , P2_U3157;
output P2_U3156 , P2_U3155 , P2_U3154 , P2_U3153 , P2_U3152 , P2_U3151 , P2_U3150;
output P2_U3149 , P2_U3148 , P2_U3147 , P2_U3146 , P2_U3145 , P2_U3144 , P2_U3143;
output P2_U3142 , P2_U3141 , P2_U3140 , P2_U3139 , P2_U3138 , P2_U3137 , P2_U3136;
output P2_U3135 , P2_U3134 , P2_U3133 , P2_U3132 , P2_U3131 , P2_U3130 , P2_U3129;
output P2_U3128 , P2_U3127 , P2_U3126 , P2_U3125 , P2_U3124 , P2_U3123 , P2_U3122;
output P2_U3121 , P2_U3120 , P2_U3119 , P2_U3118 , P2_U3117 , P2_U3116 , P2_U3115;
output P2_U3114 , P2_U3113 , P2_U3112 , P2_U3111 , P2_U3110 , P2_U3109 , P2_U3108;
output P2_U3107 , P2_U3106 , P2_U3105 , P2_U3104 , P2_U3103 , P2_U3102 , P2_U3101;
output P2_U3100 , P2_U3099 , P2_U3098 , P2_U3097 , P2_U3096 , P2_U3095 , P2_U3094;
output P2_U3093 , P2_U3092 , P2_U3091 , P2_U3090 , P2_U3089 , P2_U3088 , P2_U3087;
output P2_U3086 , P2_U3085 , P2_U3084 , P2_U3083 , P2_U3082 , P2_U3081 , P2_U3080;
output P2_U3079 , P2_U3078 , P2_U3077 , P2_U3076 , P2_U3075 , P2_U3074 , P2_U3073;
output P2_U3072 , P2_U3071 , P2_U3070 , P2_U3069 , P2_U3068 , P2_U3067 , P2_U3066;
output P2_U3065 , P2_U3064 , P2_U3063 , P2_U3062 , P2_U3061 , P2_U3060 , P2_U3059;
output P2_U3058 , P2_U3057 , P2_U3056 , P2_U3055 , P2_U3054 , P2_U3053 , P2_U3052;
output P2_U3051 , P2_U3050 , P2_U3049 , P2_U3048 , P2_U3595 , P2_U3596 , P2_U3599;
output P2_U3600 , P2_U3601 , P2_U3047 , P2_U3602 , P2_U3603 , P2_U3604 , P2_U3605;
output P2_U3046 , P2_U3045 , P2_U3044 , P2_U3043 , P2_U3042 , P2_U3041 , P2_U3040;
output P2_U3039 , P2_U3038 , P2_U3037 , P2_U3036 , P2_U3035 , P2_U3034 , P2_U3033;
output P2_U3032 , P2_U3031 , P2_U3030 , P2_U3029 , P2_U3028 , P2_U3027 , P2_U3026;
output P2_U3025 , P2_U3024 , P2_U3023 , P2_U3022 , P2_U3021 , P2_U3020 , P2_U3019;
output P2_U3018 , P2_U3017 , P2_U3016 , P2_U3015 , P2_U3014 , P2_U3013 , P2_U3012;
output P2_U3011 , P2_U3010 , P2_U3009 , P2_U3008 , P2_U3007 , P2_U3006 , P2_U3005;
output P2_U3004 , P2_U3003 , P2_U3002 , P2_U3001 , P2_U3000 , P2_U2999 , P2_U2998;
output P2_U2997 , P2_U2996 , P2_U2995 , P2_U2994 , P2_U2993 , P2_U2992 , P2_U2991;
output P2_U2990 , P2_U2989 , P2_U2988 , P2_U2987 , P2_U2986 , P2_U2985 , P2_U2984;
output P2_U2983 , P2_U2982 , P2_U2981 , P2_U2980 , P2_U2979 , P2_U2978 , P2_U2977;
output P2_U2976 , P2_U2975 , P2_U2974 , P2_U2973 , P2_U2972 , P2_U2971 , P2_U2970;
output P2_U2969 , P2_U2968 , P2_U2967 , P2_U2966 , P2_U2965 , P2_U2964 , P2_U2963;
output P2_U2962 , P2_U2961 , P2_U2960 , P2_U2959 , P2_U2958 , P2_U2957 , P2_U2956;
output P2_U2955 , P2_U2954 , P2_U2953 , P2_U2952 , P2_U2951 , P2_U2950 , P2_U2949;
output P2_U2948 , P2_U2947 , P2_U2946 , P2_U2945 , P2_U2944 , P2_U2943 , P2_U2942;
output P2_U2941 , P2_U2940 , P2_U2939 , P2_U2938 , P2_U2937 , P2_U2936 , P2_U2935;
output P2_U2934 , P2_U2933 , P2_U2932 , P2_U2931 , P2_U2930 , P2_U2929 , P2_U2928;
output P2_U2927 , P2_U2926 , P2_U2925 , P2_U2924 , P2_U2923 , P2_U2922 , P2_U2921;
output P2_U2920 , P2_U2919 , P2_U2918 , P2_U2917 , P2_U2916 , P2_U2915 , P2_U2914;
output P2_U2913 , P2_U2912 , P2_U2911 , P2_U2910 , P2_U2909 , P2_U2908 , P2_U2907;
output P2_U2906 , P2_U2905 , P2_U2904 , P2_U2903 , P2_U2902 , P2_U2901 , P2_U2900;
output P2_U2899 , P2_U2898 , P2_U2897 , P2_U2896 , P2_U2895 , P2_U2894 , P2_U2893;
output P2_U2892 , P2_U2891 , P2_U2890 , P2_U2889 , P2_U2888 , P2_U2887 , P2_U2886;
output P2_U2885 , P2_U2884 , P2_U2883 , P2_U2882 , P2_U2881 , P2_U2880 , P2_U2879;
output P2_U2878 , P2_U2877 , P2_U2876 , P2_U2875 , P2_U2874 , P2_U2873 , P2_U2872;
output P2_U2871 , P2_U2870 , P2_U2869 , P2_U2868 , P2_U2867 , P2_U2866 , P2_U2865;
output P2_U2864 , P2_U2863 , P2_U2862 , P2_U2861 , P2_U2860 , P2_U2859 , P2_U2858;
output P2_U2857 , P2_U2856 , P2_U2855 , P2_U2854 , P2_U2853 , P2_U2852 , P2_U2851;
output P2_U2850 , P2_U2849 , P2_U2848 , P2_U2847 , P2_U2846 , P2_U2845 , P2_U2844;
output P2_U2843 , P2_U2842 , P2_U2841 , P2_U2840 , P2_U2839 , P2_U2838 , P2_U2837;
output P2_U2836 , P2_U2835 , P2_U2834 , P2_U2833 , P2_U2832 , P2_U2831 , P2_U2830;
output P2_U2829 , P2_U2828 , P2_U2827 , P2_U2826 , P2_U2825 , P2_U2824 , P2_U2823;
output P2_U2822 , P2_U2821 , P2_U2820 , P2_U3608 , P2_U2819 , P2_U3609 , P2_U2818;
output P2_U3610 , P2_U2817 , P2_U3611 , P2_U2816 , P2_U2815 , P2_U3612 , P2_U2814;
output P1_U3458 , P1_U3459 , P1_U3460 , P1_U3461 , P1_U3226 , P1_U3225 , P1_U3224;
output P1_U3223 , P1_U3222 , P1_U3221 , P1_U3220 , P1_U3219 , P1_U3218 , P1_U3217;
output P1_U3216 , P1_U3215 , P1_U3214 , P1_U3213 , P1_U3212 , P1_U3211 , P1_U3210;
output P1_U3209 , P1_U3208 , P1_U3207 , P1_U3206 , P1_U3205 , P1_U3204 , P1_U3203;
output P1_U3202 , P1_U3201 , P1_U3200 , P1_U3199 , P1_U3198 , P1_U3197 , P1_U3196;
output P1_U3195 , P1_U3194 , P1_U3464 , P1_U3465 , P1_U3193 , P1_U3192 , P1_U3191;
output P1_U3190 , P1_U3189 , P1_U3188 , P1_U3187 , P1_U3186 , P1_U3185 , P1_U3184;
output P1_U3183 , P1_U3182 , P1_U3181 , P1_U3180 , P1_U3179 , P1_U3178 , P1_U3177;
output P1_U3176 , P1_U3175 , P1_U3174 , P1_U3173 , P1_U3172 , P1_U3171 , P1_U3170;
output P1_U3169 , P1_U3168 , P1_U3167 , P1_U3166 , P1_U3165 , P1_U3164 , P1_U3466;
output P1_U3163 , P1_U3162 , P1_U3161 , P1_U3160 , P1_U3159 , P1_U3158 , P1_U3157;
output P1_U3156 , P1_U3155 , P1_U3154 , P1_U3153 , P1_U3152 , P1_U3151 , P1_U3150;
output P1_U3149 , P1_U3148 , P1_U3147 , P1_U3146 , P1_U3145 , P1_U3144 , P1_U3143;
output P1_U3142 , P1_U3141 , P1_U3140 , P1_U3139 , P1_U3138 , P1_U3137 , P1_U3136;
output P1_U3135 , P1_U3134 , P1_U3133 , P1_U3132 , P1_U3131 , P1_U3130 , P1_U3129;
output P1_U3128 , P1_U3127 , P1_U3126 , P1_U3125 , P1_U3124 , P1_U3123 , P1_U3122;
output P1_U3121 , P1_U3120 , P1_U3119 , P1_U3118 , P1_U3117 , P1_U3116 , P1_U3115;
output P1_U3114 , P1_U3113 , P1_U3112 , P1_U3111 , P1_U3110 , P1_U3109 , P1_U3108;
output P1_U3107 , P1_U3106 , P1_U3105 , P1_U3104 , P1_U3103 , P1_U3102 , P1_U3101;
output P1_U3100 , P1_U3099 , P1_U3098 , P1_U3097 , P1_U3096 , P1_U3095 , P1_U3094;
output P1_U3093 , P1_U3092 , P1_U3091 , P1_U3090 , P1_U3089 , P1_U3088 , P1_U3087;
output P1_U3086 , P1_U3085 , P1_U3084 , P1_U3083 , P1_U3082 , P1_U3081 , P1_U3080;
output P1_U3079 , P1_U3078 , P1_U3077 , P1_U3076 , P1_U3075 , P1_U3074 , P1_U3073;
output P1_U3072 , P1_U3071 , P1_U3070 , P1_U3069 , P1_U3068 , P1_U3067 , P1_U3066;
output P1_U3065 , P1_U3064 , P1_U3063 , P1_U3062 , P1_U3061 , P1_U3060 , P1_U3059;
output P1_U3058 , P1_U3057 , P1_U3056 , P1_U3055 , P1_U3054 , P1_U3053 , P1_U3052;
output P1_U3051 , P1_U3050 , P1_U3049 , P1_U3048 , P1_U3047 , P1_U3046 , P1_U3045;
output P1_U3044 , P1_U3043 , P1_U3042 , P1_U3041 , P1_U3040 , P1_U3039 , P1_U3038;
output P1_U3037 , P1_U3036 , P1_U3035 , P1_U3034 , P1_U3033 , P1_U3468 , P1_U3469;
output P1_U3472 , P1_U3473 , P1_U3474 , P1_U3032 , P1_U3475 , P1_U3476 , P1_U3477;
output P1_U3478 , P1_U3031 , P1_U3030 , P1_U3029 , P1_U3028 , P1_U3027 , P1_U3026;
output P1_U3025 , P1_U3024 , P1_U3023 , P1_U3022 , P1_U3021 , P1_U3020 , P1_U3019;
output P1_U3018 , P1_U3017 , P1_U3016 , P1_U3015 , P1_U3014 , P1_U3013 , P1_U3012;
output P1_U3011 , P1_U3010 , P1_U3009 , P1_U3008 , P1_U3007 , P1_U3006 , P1_U3005;
output P1_U3004 , P1_U3003 , P1_U3002 , P1_U3001 , P1_U3000 , P1_U2999 , P1_U2998;
output P1_U2997 , P1_U2996 , P1_U2995 , P1_U2994 , P1_U2993 , P1_U2992 , P1_U2991;
output P1_U2990 , P1_U2989 , P1_U2988 , P1_U2987 , P1_U2986 , P1_U2985 , P1_U2984;
output P1_U2983 , P1_U2982 , P1_U2981 , P1_U2980 , P1_U2979 , P1_U2978 , P1_U2977;
output P1_U2976 , P1_U2975 , P1_U2974 , P1_U2973 , P1_U2972 , P1_U2971 , P1_U2970;
output P1_U2969 , P1_U2968 , P1_U2967 , P1_U2966 , P1_U2965 , P1_U2964 , P1_U2963;
output P1_U2962 , P1_U2961 , P1_U2960 , P1_U2959 , P1_U2958 , P1_U2957 , P1_U2956;
output P1_U2955 , P1_U2954 , P1_U2953 , P1_U2952 , P1_U2951 , P1_U2950 , P1_U2949;
output P1_U2948 , P1_U2947 , P1_U2946 , P1_U2945 , P1_U2944 , P1_U2943 , P1_U2942;
output P1_U2941 , P1_U2940 , P1_U2939 , P1_U2938 , P1_U2937 , P1_U2936 , P1_U2935;
output P1_U2934 , P1_U2933 , P1_U2932 , P1_U2931 , P1_U2930 , P1_U2929 , P1_U2928;
output P1_U2927 , P1_U2926 , P1_U2925 , P1_U2924 , P1_U2923 , P1_U2922 , P1_U2921;
output P1_U2920 , P1_U2919 , P1_U2918 , P1_U2917 , P1_U2916 , P1_U2915 , P1_U2914;
output P1_U2913 , P1_U2912 , P1_U2911 , P1_U2910 , P1_U2909 , P1_U2908 , P1_U2907;
output P1_U2906 , P1_U2905 , P1_U2904 , P1_U2903 , P1_U2902 , P1_U2901 , P1_U2900;
output P1_U2899 , P1_U2898 , P1_U2897 , P1_U2896 , P1_U2895 , P1_U2894 , P1_U2893;
output P1_U2892 , P1_U2891 , P1_U2890 , P1_U2889 , P1_U2888 , P1_U2887 , P1_U2886;
output P1_U2885 , P1_U2884 , P1_U2883 , P1_U2882 , P1_U2881 , P1_U2880 , P1_U2879;
output P1_U2878 , P1_U2877 , P1_U2876 , P1_U2875 , P1_U2874 , P1_U2873 , P1_U2872;
output P1_U2871 , P1_U2870 , P1_U2869 , P1_U2868 , P1_U2867 , P1_U2866 , P1_U2865;
output P1_U2864 , P1_U2863 , P1_U2862 , P1_U2861 , P1_U2860 , P1_U2859 , P1_U2858;
output P1_U2857 , P1_U2856 , P1_U2855 , P1_U2854 , P1_U2853 , P1_U2852 , P1_U2851;
output P1_U2850 , P1_U2849 , P1_U2848 , P1_U2847 , P1_U2846 , P1_U2845 , P1_U2844;
output P1_U2843 , P1_U2842 , P1_U2841 , P1_U2840 , P1_U2839 , P1_U2838 , P1_U2837;
output P1_U2836 , P1_U2835 , P1_U2834 , P1_U2833 , P1_U2832 , P1_U2831 , P1_U2830;
output P1_U2829 , P1_U2828 , P1_U2827 , P1_U2826 , P1_U2825 , P1_U2824 , P1_U2823;
output P1_U2822 , P1_U2821 , P1_U2820 , P1_U2819 , P1_U2818 , P1_U2817 , P1_U2816;
output P1_U2815 , P1_U2814 , P1_U2813 , P1_U2812 , P1_U2811 , P1_U2810 , P1_U2809;
output P1_U2808 , P1_U3481 , P1_U2807 , P1_U3482 , P1_U3483 , P1_U2806 , P1_U3484;
output P1_U2805 , P1_U3485 , P1_U2804 , P1_U3486 , P1_U2803 , P1_U2802 , P1_U3487;
output P1_U2801;

input DATAI_31_ , DATAI_30_ , DATAI_29_ , DATAI_28_ , DATAI_27_ , DATAI_26_;
input DATAI_25_ , DATAI_24_ , DATAI_23_ , DATAI_22_ , DATAI_21_ , DATAI_20_;
input DATAI_19_ , DATAI_18_ , DATAI_17_ , DATAI_16_ , DATAI_15_ , DATAI_14_;
input DATAI_13_ , DATAI_12_ , DATAI_11_ , DATAI_10_ , DATAI_9_ , DATAI_8_;
input DATAI_7_ , DATAI_6_ , DATAI_5_ , DATAI_4_ , DATAI_3_ , DATAI_2_;
input DATAI_1_ , DATAI_0_ , HOLD , NA , BS16 , READY1;
input READY2;
input BUF1_REG_0_ , BUF1_REG_1_ , BUF1_REG_2_ , BUF1_REG_3_ , BUF1_REG_4_ , BUF1_REG_5_;
input BUF1_REG_6_ , BUF1_REG_7_ , BUF1_REG_8_ , BUF1_REG_9_ , BUF1_REG_10_ , BUF1_REG_11_;
input BUF1_REG_12_ , BUF1_REG_13_ , BUF1_REG_14_ , BUF1_REG_15_ , BUF1_REG_16_ , BUF1_REG_17_;
input BUF1_REG_18_ , BUF1_REG_19_ , BUF1_REG_20_ , BUF1_REG_21_ , BUF1_REG_22_ , BUF1_REG_23_;
input BUF1_REG_24_ , BUF1_REG_25_ , BUF1_REG_26_ , BUF1_REG_27_ , BUF1_REG_28_ , BUF1_REG_29_;
input BUF1_REG_30_ , BUF1_REG_31_ , BUF2_REG_0_ , BUF2_REG_1_ , BUF2_REG_2_ , BUF2_REG_3_;
input BUF2_REG_4_ , BUF2_REG_5_ , BUF2_REG_6_ , BUF2_REG_7_ , BUF2_REG_8_ , BUF2_REG_9_;
input BUF2_REG_10_ , BUF2_REG_11_ , BUF2_REG_12_ , BUF2_REG_13_ , BUF2_REG_14_ , BUF2_REG_15_;
input BUF2_REG_16_ , BUF2_REG_17_ , BUF2_REG_18_ , BUF2_REG_19_ , BUF2_REG_20_ , BUF2_REG_21_;
input BUF2_REG_22_ , BUF2_REG_23_ , BUF2_REG_24_ , BUF2_REG_25_ , BUF2_REG_26_ , BUF2_REG_27_;
input BUF2_REG_28_ , BUF2_REG_29_ , BUF2_REG_30_ , BUF2_REG_31_ , READY12_REG , READY21_REG;
input READY22_REG , READY11_REG , P3_BE_N_REG_3_ , P3_BE_N_REG_2_ , P3_BE_N_REG_1_ , P3_BE_N_REG_0_;
input P3_ADDRESS_REG_29_ , P3_ADDRESS_REG_28_ , P3_ADDRESS_REG_27_ , P3_ADDRESS_REG_26_ , P3_ADDRESS_REG_25_ , P3_ADDRESS_REG_24_;
input P3_ADDRESS_REG_23_ , P3_ADDRESS_REG_22_ , P3_ADDRESS_REG_21_ , P3_ADDRESS_REG_20_ , P3_ADDRESS_REG_19_ , P3_ADDRESS_REG_18_;
input P3_ADDRESS_REG_17_ , P3_ADDRESS_REG_16_ , P3_ADDRESS_REG_15_ , P3_ADDRESS_REG_14_ , P3_ADDRESS_REG_13_ , P3_ADDRESS_REG_12_;
input P3_ADDRESS_REG_11_ , P3_ADDRESS_REG_10_ , P3_ADDRESS_REG_9_ , P3_ADDRESS_REG_8_ , P3_ADDRESS_REG_7_ , P3_ADDRESS_REG_6_;
input P3_ADDRESS_REG_5_ , P3_ADDRESS_REG_4_ , P3_ADDRESS_REG_3_ , P3_ADDRESS_REG_2_ , P3_ADDRESS_REG_1_ , P3_ADDRESS_REG_0_;
input P3_STATE_REG_2_ , P3_STATE_REG_1_ , P3_STATE_REG_0_ , P3_DATAWIDTH_REG_0_ , P3_DATAWIDTH_REG_1_ , P3_DATAWIDTH_REG_2_;
input P3_DATAWIDTH_REG_3_ , P3_DATAWIDTH_REG_4_ , P3_DATAWIDTH_REG_5_ , P3_DATAWIDTH_REG_6_ , P3_DATAWIDTH_REG_7_ , P3_DATAWIDTH_REG_8_;
input P3_DATAWIDTH_REG_9_ , P3_DATAWIDTH_REG_10_ , P3_DATAWIDTH_REG_11_ , P3_DATAWIDTH_REG_12_ , P3_DATAWIDTH_REG_13_ , P3_DATAWIDTH_REG_14_;
input P3_DATAWIDTH_REG_15_ , P3_DATAWIDTH_REG_16_ , P3_DATAWIDTH_REG_17_ , P3_DATAWIDTH_REG_18_ , P3_DATAWIDTH_REG_19_ , P3_DATAWIDTH_REG_20_;
input P3_DATAWIDTH_REG_21_ , P3_DATAWIDTH_REG_22_ , P3_DATAWIDTH_REG_23_ , P3_DATAWIDTH_REG_24_ , P3_DATAWIDTH_REG_25_ , P3_DATAWIDTH_REG_26_;
input P3_DATAWIDTH_REG_27_ , P3_DATAWIDTH_REG_28_ , P3_DATAWIDTH_REG_29_ , P3_DATAWIDTH_REG_30_ , P3_DATAWIDTH_REG_31_ , P3_STATE2_REG_3_;
input P3_STATE2_REG_2_ , P3_STATE2_REG_1_ , P3_STATE2_REG_0_ , P3_INSTQUEUE_REG_15__7_ , P3_INSTQUEUE_REG_15__6_ , P3_INSTQUEUE_REG_15__5_;
input P3_INSTQUEUE_REG_15__4_ , P3_INSTQUEUE_REG_15__3_ , P3_INSTQUEUE_REG_15__2_ , P3_INSTQUEUE_REG_15__1_ , P3_INSTQUEUE_REG_15__0_ , P3_INSTQUEUE_REG_14__7_;
input P3_INSTQUEUE_REG_14__6_ , P3_INSTQUEUE_REG_14__5_ , P3_INSTQUEUE_REG_14__4_ , P3_INSTQUEUE_REG_14__3_ , P3_INSTQUEUE_REG_14__2_ , P3_INSTQUEUE_REG_14__1_;
input P3_INSTQUEUE_REG_14__0_ , P3_INSTQUEUE_REG_13__7_ , P3_INSTQUEUE_REG_13__6_ , P3_INSTQUEUE_REG_13__5_ , P3_INSTQUEUE_REG_13__4_ , P3_INSTQUEUE_REG_13__3_;
input P3_INSTQUEUE_REG_13__2_ , P3_INSTQUEUE_REG_13__1_ , P3_INSTQUEUE_REG_13__0_ , P3_INSTQUEUE_REG_12__7_ , P3_INSTQUEUE_REG_12__6_ , P3_INSTQUEUE_REG_12__5_;
input P3_INSTQUEUE_REG_12__4_ , P3_INSTQUEUE_REG_12__3_ , P3_INSTQUEUE_REG_12__2_ , P3_INSTQUEUE_REG_12__1_ , P3_INSTQUEUE_REG_12__0_ , P3_INSTQUEUE_REG_11__7_;
input P3_INSTQUEUE_REG_11__6_ , P3_INSTQUEUE_REG_11__5_ , P3_INSTQUEUE_REG_11__4_ , P3_INSTQUEUE_REG_11__3_ , P3_INSTQUEUE_REG_11__2_ , P3_INSTQUEUE_REG_11__1_;
input P3_INSTQUEUE_REG_11__0_ , P3_INSTQUEUE_REG_10__7_ , P3_INSTQUEUE_REG_10__6_ , P3_INSTQUEUE_REG_10__5_ , P3_INSTQUEUE_REG_10__4_ , P3_INSTQUEUE_REG_10__3_;
input P3_INSTQUEUE_REG_10__2_ , P3_INSTQUEUE_REG_10__1_ , P3_INSTQUEUE_REG_10__0_ , P3_INSTQUEUE_REG_9__7_ , P3_INSTQUEUE_REG_9__6_ , P3_INSTQUEUE_REG_9__5_;
input P3_INSTQUEUE_REG_9__4_ , P3_INSTQUEUE_REG_9__3_ , P3_INSTQUEUE_REG_9__2_ , P3_INSTQUEUE_REG_9__1_ , P3_INSTQUEUE_REG_9__0_ , P3_INSTQUEUE_REG_8__7_;
input P3_INSTQUEUE_REG_8__6_ , P3_INSTQUEUE_REG_8__5_ , P3_INSTQUEUE_REG_8__4_ , P3_INSTQUEUE_REG_8__3_ , P3_INSTQUEUE_REG_8__2_ , P3_INSTQUEUE_REG_8__1_;
input P3_INSTQUEUE_REG_8__0_ , P3_INSTQUEUE_REG_7__7_ , P3_INSTQUEUE_REG_7__6_ , P3_INSTQUEUE_REG_7__5_ , P3_INSTQUEUE_REG_7__4_ , P3_INSTQUEUE_REG_7__3_;
input P3_INSTQUEUE_REG_7__2_ , P3_INSTQUEUE_REG_7__1_ , P3_INSTQUEUE_REG_7__0_ , P3_INSTQUEUE_REG_6__7_ , P3_INSTQUEUE_REG_6__6_ , P3_INSTQUEUE_REG_6__5_;
input P3_INSTQUEUE_REG_6__4_ , P3_INSTQUEUE_REG_6__3_ , P3_INSTQUEUE_REG_6__2_ , P3_INSTQUEUE_REG_6__1_ , P3_INSTQUEUE_REG_6__0_ , P3_INSTQUEUE_REG_5__7_;
input P3_INSTQUEUE_REG_5__6_ , P3_INSTQUEUE_REG_5__5_ , P3_INSTQUEUE_REG_5__4_ , P3_INSTQUEUE_REG_5__3_ , P3_INSTQUEUE_REG_5__2_ , P3_INSTQUEUE_REG_5__1_;
input P3_INSTQUEUE_REG_5__0_ , P3_INSTQUEUE_REG_4__7_ , P3_INSTQUEUE_REG_4__6_ , P3_INSTQUEUE_REG_4__5_ , P3_INSTQUEUE_REG_4__4_ , P3_INSTQUEUE_REG_4__3_;
input P3_INSTQUEUE_REG_4__2_ , P3_INSTQUEUE_REG_4__1_ , P3_INSTQUEUE_REG_4__0_ , P3_INSTQUEUE_REG_3__7_ , P3_INSTQUEUE_REG_3__6_ , P3_INSTQUEUE_REG_3__5_;
input P3_INSTQUEUE_REG_3__4_ , P3_INSTQUEUE_REG_3__3_ , P3_INSTQUEUE_REG_3__2_ , P3_INSTQUEUE_REG_3__1_ , P3_INSTQUEUE_REG_3__0_ , P3_INSTQUEUE_REG_2__7_;
input P3_INSTQUEUE_REG_2__6_ , P3_INSTQUEUE_REG_2__5_ , P3_INSTQUEUE_REG_2__4_ , P3_INSTQUEUE_REG_2__3_ , P3_INSTQUEUE_REG_2__2_ , P3_INSTQUEUE_REG_2__1_;
input P3_INSTQUEUE_REG_2__0_ , P3_INSTQUEUE_REG_1__7_ , P3_INSTQUEUE_REG_1__6_ , P3_INSTQUEUE_REG_1__5_ , P3_INSTQUEUE_REG_1__4_ , P3_INSTQUEUE_REG_1__3_;
input P3_INSTQUEUE_REG_1__2_ , P3_INSTQUEUE_REG_1__1_ , P3_INSTQUEUE_REG_1__0_ , P3_INSTQUEUE_REG_0__7_ , P3_INSTQUEUE_REG_0__6_ , P3_INSTQUEUE_REG_0__5_;
input P3_INSTQUEUE_REG_0__4_ , P3_INSTQUEUE_REG_0__3_ , P3_INSTQUEUE_REG_0__2_ , P3_INSTQUEUE_REG_0__1_ , P3_INSTQUEUE_REG_0__0_ , P3_INSTQUEUERD_ADDR_REG_4_;
input P3_INSTQUEUERD_ADDR_REG_3_ , P3_INSTQUEUERD_ADDR_REG_2_ , P3_INSTQUEUERD_ADDR_REG_1_ , P3_INSTQUEUERD_ADDR_REG_0_ , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_INSTQUEUEWR_ADDR_REG_3_;
input P3_INSTQUEUEWR_ADDR_REG_2_ , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_INSTADDRPOINTER_REG_0_ , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_2_;
input P3_INSTADDRPOINTER_REG_3_ , P3_INSTADDRPOINTER_REG_4_ , P3_INSTADDRPOINTER_REG_5_ , P3_INSTADDRPOINTER_REG_6_ , P3_INSTADDRPOINTER_REG_7_ , P3_INSTADDRPOINTER_REG_8_;
input P3_INSTADDRPOINTER_REG_9_ , P3_INSTADDRPOINTER_REG_10_ , P3_INSTADDRPOINTER_REG_11_ , P3_INSTADDRPOINTER_REG_12_ , P3_INSTADDRPOINTER_REG_13_ , P3_INSTADDRPOINTER_REG_14_;
input P3_INSTADDRPOINTER_REG_15_ , P3_INSTADDRPOINTER_REG_16_ , P3_INSTADDRPOINTER_REG_17_ , P3_INSTADDRPOINTER_REG_18_ , P3_INSTADDRPOINTER_REG_19_ , P3_INSTADDRPOINTER_REG_20_;
input P3_INSTADDRPOINTER_REG_21_ , P3_INSTADDRPOINTER_REG_22_ , P3_INSTADDRPOINTER_REG_23_ , P3_INSTADDRPOINTER_REG_24_ , P3_INSTADDRPOINTER_REG_25_ , P3_INSTADDRPOINTER_REG_26_;
input P3_INSTADDRPOINTER_REG_27_ , P3_INSTADDRPOINTER_REG_28_ , P3_INSTADDRPOINTER_REG_29_ , P3_INSTADDRPOINTER_REG_30_ , P3_INSTADDRPOINTER_REG_31_ , P3_PHYADDRPOINTER_REG_0_;
input P3_PHYADDRPOINTER_REG_1_ , P3_PHYADDRPOINTER_REG_2_ , P3_PHYADDRPOINTER_REG_3_ , P3_PHYADDRPOINTER_REG_4_ , P3_PHYADDRPOINTER_REG_5_ , P3_PHYADDRPOINTER_REG_6_;
input P3_PHYADDRPOINTER_REG_7_ , P3_PHYADDRPOINTER_REG_8_ , P3_PHYADDRPOINTER_REG_9_ , P3_PHYADDRPOINTER_REG_10_ , P3_PHYADDRPOINTER_REG_11_ , P3_PHYADDRPOINTER_REG_12_;
input P3_PHYADDRPOINTER_REG_13_ , P3_PHYADDRPOINTER_REG_14_ , P3_PHYADDRPOINTER_REG_15_ , P3_PHYADDRPOINTER_REG_16_ , P3_PHYADDRPOINTER_REG_17_ , P3_PHYADDRPOINTER_REG_18_;
input P3_PHYADDRPOINTER_REG_19_ , P3_PHYADDRPOINTER_REG_20_ , P3_PHYADDRPOINTER_REG_21_ , P3_PHYADDRPOINTER_REG_22_ , P3_PHYADDRPOINTER_REG_23_ , P3_PHYADDRPOINTER_REG_24_;
input P3_PHYADDRPOINTER_REG_25_ , P3_PHYADDRPOINTER_REG_26_ , P3_PHYADDRPOINTER_REG_27_ , P3_PHYADDRPOINTER_REG_28_ , P3_PHYADDRPOINTER_REG_29_ , P3_PHYADDRPOINTER_REG_30_;
input P3_PHYADDRPOINTER_REG_31_ , P3_LWORD_REG_15_ , P3_LWORD_REG_14_ , P3_LWORD_REG_13_ , P3_LWORD_REG_12_ , P3_LWORD_REG_11_;
input P3_LWORD_REG_10_ , P3_LWORD_REG_9_ , P3_LWORD_REG_8_ , P3_LWORD_REG_7_ , P3_LWORD_REG_6_ , P3_LWORD_REG_5_;
input P3_LWORD_REG_4_ , P3_LWORD_REG_3_ , P3_LWORD_REG_2_ , P3_LWORD_REG_1_ , P3_LWORD_REG_0_ , P3_UWORD_REG_14_;
input P3_UWORD_REG_13_ , P3_UWORD_REG_12_ , P3_UWORD_REG_11_ , P3_UWORD_REG_10_ , P3_UWORD_REG_9_ , P3_UWORD_REG_8_;
input P3_UWORD_REG_7_ , P3_UWORD_REG_6_ , P3_UWORD_REG_5_ , P3_UWORD_REG_4_ , P3_UWORD_REG_3_ , P3_UWORD_REG_2_;
input P3_UWORD_REG_1_ , P3_UWORD_REG_0_ , P3_DATAO_REG_0__EXTRA , P3_DATAO_REG_1__EXTRA , P3_DATAO_REG_2__EXTRA , P3_DATAO_REG_3__EXTRA;
input P3_DATAO_REG_4__EXTRA , P3_DATAO_REG_5__EXTRA , P3_DATAO_REG_6__EXTRA , P3_DATAO_REG_7__EXTRA , P3_DATAO_REG_8__EXTRA , P3_DATAO_REG_9__EXTRA;
input P3_DATAO_REG_10__EXTRA , P3_DATAO_REG_11__EXTRA , P3_DATAO_REG_12__EXTRA , P3_DATAO_REG_13__EXTRA , P3_DATAO_REG_14__EXTRA , P3_DATAO_REG_15__EXTRA;
input P3_DATAO_REG_16__EXTRA , P3_DATAO_REG_17__EXTRA , P3_DATAO_REG_18__EXTRA , P3_DATAO_REG_19__EXTRA , P3_DATAO_REG_20__EXTRA , P3_DATAO_REG_21__EXTRA;
input P3_DATAO_REG_22__EXTRA , P3_DATAO_REG_23__EXTRA , P3_DATAO_REG_24__EXTRA , P3_DATAO_REG_25__EXTRA , P3_DATAO_REG_26__EXTRA , P3_DATAO_REG_27__EXTRA;
input P3_DATAO_REG_28__EXTRA , P3_DATAO_REG_29__EXTRA , P3_DATAO_REG_30__EXTRA , P3_DATAO_REG_31__EXTRA , P3_EAX_REG_0_ , P3_EAX_REG_1_;
input P3_EAX_REG_2_ , P3_EAX_REG_3_ , P3_EAX_REG_4_ , P3_EAX_REG_5_ , P3_EAX_REG_6_ , P3_EAX_REG_7_;
input P3_EAX_REG_8_ , P3_EAX_REG_9_ , P3_EAX_REG_10_ , P3_EAX_REG_11_ , P3_EAX_REG_12_ , P3_EAX_REG_13_;
input P3_EAX_REG_14_ , P3_EAX_REG_15_ , P3_EAX_REG_16_ , P3_EAX_REG_17_ , P3_EAX_REG_18_ , P3_EAX_REG_19_;
input P3_EAX_REG_20_ , P3_EAX_REG_21_ , P3_EAX_REG_22_ , P3_EAX_REG_23_ , P3_EAX_REG_24_ , P3_EAX_REG_25_;
input P3_EAX_REG_26_ , P3_EAX_REG_27_ , P3_EAX_REG_28_ , P3_EAX_REG_29_ , P3_EAX_REG_30_ , P3_EAX_REG_31_;
input P3_EBX_REG_0_ , P3_EBX_REG_1_ , P3_EBX_REG_2_ , P3_EBX_REG_3_ , P3_EBX_REG_4_ , P3_EBX_REG_5_;
input P3_EBX_REG_6_ , P3_EBX_REG_7_ , P3_EBX_REG_8_ , P3_EBX_REG_9_ , P3_EBX_REG_10_ , P3_EBX_REG_11_;
input P3_EBX_REG_12_ , P3_EBX_REG_13_ , P3_EBX_REG_14_ , P3_EBX_REG_15_ , P3_EBX_REG_16_ , P3_EBX_REG_17_;
input P3_EBX_REG_18_ , P3_EBX_REG_19_ , P3_EBX_REG_20_ , P3_EBX_REG_21_ , P3_EBX_REG_22_ , P3_EBX_REG_23_;
input P3_EBX_REG_24_ , P3_EBX_REG_25_ , P3_EBX_REG_26_ , P3_EBX_REG_27_ , P3_EBX_REG_28_ , P3_EBX_REG_29_;
input P3_EBX_REG_30_ , P3_EBX_REG_31_ , P3_REIP_REG_0_ , P3_REIP_REG_1_ , P3_REIP_REG_2_ , P3_REIP_REG_3_;
input P3_REIP_REG_4_ , P3_REIP_REG_5_ , P3_REIP_REG_6_ , P3_REIP_REG_7_ , P3_REIP_REG_8_ , P3_REIP_REG_9_;
input P3_REIP_REG_10_ , P3_REIP_REG_11_ , P3_REIP_REG_12_ , P3_REIP_REG_13_ , P3_REIP_REG_14_ , P3_REIP_REG_15_;
input P3_REIP_REG_16_ , P3_REIP_REG_17_ , P3_REIP_REG_18_ , P3_REIP_REG_19_ , P3_REIP_REG_20_ , P3_REIP_REG_21_;
input P3_REIP_REG_22_ , P3_REIP_REG_23_ , P3_REIP_REG_24_ , P3_REIP_REG_25_ , P3_REIP_REG_26_ , P3_REIP_REG_27_;
input P3_REIP_REG_28_ , P3_REIP_REG_29_ , P3_REIP_REG_30_ , P3_REIP_REG_31_ , P3_BYTEENABLE_REG_3_ , P3_BYTEENABLE_REG_2_;
input P3_BYTEENABLE_REG_1_ , P3_BYTEENABLE_REG_0_ , P3_W_R_N_REG_EXTRA , P3_FLUSH_REG , P3_MORE_REG , P3_STATEBS16_REG;
input P3_REQUESTPENDING_REG , P3_D_C_N_REG_EXTRA , P3_M_IO_N_REG_EXTRA , P3_CODEFETCH_REG , P3_ADS_N_REG_EXTRA , P3_READREQUEST_REG;
input P3_MEMORYFETCH_REG , P2_BE_N_REG_3_ , P2_BE_N_REG_2_ , P2_BE_N_REG_1_ , P2_BE_N_REG_0_ , P2_ADDRESS_REG_29_;
input P2_ADDRESS_REG_28_ , P2_ADDRESS_REG_27_ , P2_ADDRESS_REG_26_ , P2_ADDRESS_REG_25_ , P2_ADDRESS_REG_24_ , P2_ADDRESS_REG_23_;
input P2_ADDRESS_REG_22_ , P2_ADDRESS_REG_21_ , P2_ADDRESS_REG_20_ , P2_ADDRESS_REG_19_ , P2_ADDRESS_REG_18_ , P2_ADDRESS_REG_17_;
input P2_ADDRESS_REG_16_ , P2_ADDRESS_REG_15_ , P2_ADDRESS_REG_14_ , P2_ADDRESS_REG_13_ , P2_ADDRESS_REG_12_ , P2_ADDRESS_REG_11_;
input P2_ADDRESS_REG_10_ , P2_ADDRESS_REG_9_ , P2_ADDRESS_REG_8_ , P2_ADDRESS_REG_7_ , P2_ADDRESS_REG_6_ , P2_ADDRESS_REG_5_;
input P2_ADDRESS_REG_4_ , P2_ADDRESS_REG_3_ , P2_ADDRESS_REG_2_ , P2_ADDRESS_REG_1_ , P2_ADDRESS_REG_0_ , P2_STATE_REG_2_;
input P2_STATE_REG_1_ , P2_STATE_REG_0_ , P2_DATAWIDTH_REG_0_ , P2_DATAWIDTH_REG_1_ , P2_DATAWIDTH_REG_2_ , P2_DATAWIDTH_REG_3_;
input P2_DATAWIDTH_REG_4_ , P2_DATAWIDTH_REG_5_ , P2_DATAWIDTH_REG_6_ , P2_DATAWIDTH_REG_7_ , P2_DATAWIDTH_REG_8_ , P2_DATAWIDTH_REG_9_;
input P2_DATAWIDTH_REG_10_ , P2_DATAWIDTH_REG_11_ , P2_DATAWIDTH_REG_12_ , P2_DATAWIDTH_REG_13_ , P2_DATAWIDTH_REG_14_ , P2_DATAWIDTH_REG_15_;
input P2_DATAWIDTH_REG_16_ , P2_DATAWIDTH_REG_17_ , P2_DATAWIDTH_REG_18_ , P2_DATAWIDTH_REG_19_ , P2_DATAWIDTH_REG_20_ , P2_DATAWIDTH_REG_21_;
input P2_DATAWIDTH_REG_22_ , P2_DATAWIDTH_REG_23_ , P2_DATAWIDTH_REG_24_ , P2_DATAWIDTH_REG_25_ , P2_DATAWIDTH_REG_26_ , P2_DATAWIDTH_REG_27_;
input P2_DATAWIDTH_REG_28_ , P2_DATAWIDTH_REG_29_ , P2_DATAWIDTH_REG_30_ , P2_DATAWIDTH_REG_31_ , P2_STATE2_REG_3_ , P2_STATE2_REG_2_;
input P2_STATE2_REG_1_ , P2_STATE2_REG_0_ , P2_INSTQUEUE_REG_15__7_ , P2_INSTQUEUE_REG_15__6_ , P2_INSTQUEUE_REG_15__5_ , P2_INSTQUEUE_REG_15__4_;
input P2_INSTQUEUE_REG_15__3_ , P2_INSTQUEUE_REG_15__2_ , P2_INSTQUEUE_REG_15__1_ , P2_INSTQUEUE_REG_15__0_ , P2_INSTQUEUE_REG_14__7_ , P2_INSTQUEUE_REG_14__6_;
input P2_INSTQUEUE_REG_14__5_ , P2_INSTQUEUE_REG_14__4_ , P2_INSTQUEUE_REG_14__3_ , P2_INSTQUEUE_REG_14__2_ , P2_INSTQUEUE_REG_14__1_ , P2_INSTQUEUE_REG_14__0_;
input P2_INSTQUEUE_REG_13__7_ , P2_INSTQUEUE_REG_13__6_ , P2_INSTQUEUE_REG_13__5_ , P2_INSTQUEUE_REG_13__4_ , P2_INSTQUEUE_REG_13__3_ , P2_INSTQUEUE_REG_13__2_;
input P2_INSTQUEUE_REG_13__1_ , P2_INSTQUEUE_REG_13__0_ , P2_INSTQUEUE_REG_12__7_ , P2_INSTQUEUE_REG_12__6_ , P2_INSTQUEUE_REG_12__5_ , P2_INSTQUEUE_REG_12__4_;
input P2_INSTQUEUE_REG_12__3_ , P2_INSTQUEUE_REG_12__2_ , P2_INSTQUEUE_REG_12__1_ , P2_INSTQUEUE_REG_12__0_ , P2_INSTQUEUE_REG_11__7_ , P2_INSTQUEUE_REG_11__6_;
input P2_INSTQUEUE_REG_11__5_ , P2_INSTQUEUE_REG_11__4_ , P2_INSTQUEUE_REG_11__3_ , P2_INSTQUEUE_REG_11__2_ , P2_INSTQUEUE_REG_11__1_ , P2_INSTQUEUE_REG_11__0_;
input P2_INSTQUEUE_REG_10__7_ , P2_INSTQUEUE_REG_10__6_ , P2_INSTQUEUE_REG_10__5_ , P2_INSTQUEUE_REG_10__4_ , P2_INSTQUEUE_REG_10__3_ , P2_INSTQUEUE_REG_10__2_;
input P2_INSTQUEUE_REG_10__1_ , P2_INSTQUEUE_REG_10__0_ , P2_INSTQUEUE_REG_9__7_ , P2_INSTQUEUE_REG_9__6_ , P2_INSTQUEUE_REG_9__5_ , P2_INSTQUEUE_REG_9__4_;
input P2_INSTQUEUE_REG_9__3_ , P2_INSTQUEUE_REG_9__2_ , P2_INSTQUEUE_REG_9__1_ , P2_INSTQUEUE_REG_9__0_ , P2_INSTQUEUE_REG_8__7_ , P2_INSTQUEUE_REG_8__6_;
input P2_INSTQUEUE_REG_8__5_ , P2_INSTQUEUE_REG_8__4_ , P2_INSTQUEUE_REG_8__3_ , P2_INSTQUEUE_REG_8__2_ , P2_INSTQUEUE_REG_8__1_ , P2_INSTQUEUE_REG_8__0_;
input P2_INSTQUEUE_REG_7__7_ , P2_INSTQUEUE_REG_7__6_ , P2_INSTQUEUE_REG_7__5_ , P2_INSTQUEUE_REG_7__4_ , P2_INSTQUEUE_REG_7__3_ , P2_INSTQUEUE_REG_7__2_;
input P2_INSTQUEUE_REG_7__1_ , P2_INSTQUEUE_REG_7__0_ , P2_INSTQUEUE_REG_6__7_ , P2_INSTQUEUE_REG_6__6_ , P2_INSTQUEUE_REG_6__5_ , P2_INSTQUEUE_REG_6__4_;
input P2_INSTQUEUE_REG_6__3_ , P2_INSTQUEUE_REG_6__2_ , P2_INSTQUEUE_REG_6__1_ , P2_INSTQUEUE_REG_6__0_ , P2_INSTQUEUE_REG_5__7_ , P2_INSTQUEUE_REG_5__6_;
input P2_INSTQUEUE_REG_5__5_ , P2_INSTQUEUE_REG_5__4_ , P2_INSTQUEUE_REG_5__3_ , P2_INSTQUEUE_REG_5__2_ , P2_INSTQUEUE_REG_5__1_ , P2_INSTQUEUE_REG_5__0_;
input P2_INSTQUEUE_REG_4__7_ , P2_INSTQUEUE_REG_4__6_ , P2_INSTQUEUE_REG_4__5_ , P2_INSTQUEUE_REG_4__4_ , P2_INSTQUEUE_REG_4__3_ , P2_INSTQUEUE_REG_4__2_;
input P2_INSTQUEUE_REG_4__1_ , P2_INSTQUEUE_REG_4__0_ , P2_INSTQUEUE_REG_3__7_ , P2_INSTQUEUE_REG_3__6_ , P2_INSTQUEUE_REG_3__5_ , P2_INSTQUEUE_REG_3__4_;
input P2_INSTQUEUE_REG_3__3_ , P2_INSTQUEUE_REG_3__2_ , P2_INSTQUEUE_REG_3__1_ , P2_INSTQUEUE_REG_3__0_ , P2_INSTQUEUE_REG_2__7_ , P2_INSTQUEUE_REG_2__6_;
input P2_INSTQUEUE_REG_2__5_ , P2_INSTQUEUE_REG_2__4_ , P2_INSTQUEUE_REG_2__3_ , P2_INSTQUEUE_REG_2__2_ , P2_INSTQUEUE_REG_2__1_ , P2_INSTQUEUE_REG_2__0_;
input P2_INSTQUEUE_REG_1__7_ , P2_INSTQUEUE_REG_1__6_ , P2_INSTQUEUE_REG_1__5_ , P2_INSTQUEUE_REG_1__4_ , P2_INSTQUEUE_REG_1__3_ , P2_INSTQUEUE_REG_1__2_;
input P2_INSTQUEUE_REG_1__1_ , P2_INSTQUEUE_REG_1__0_ , P2_INSTQUEUE_REG_0__7_ , P2_INSTQUEUE_REG_0__6_ , P2_INSTQUEUE_REG_0__5_ , P2_INSTQUEUE_REG_0__4_;
input P2_INSTQUEUE_REG_0__3_ , P2_INSTQUEUE_REG_0__2_ , P2_INSTQUEUE_REG_0__1_ , P2_INSTQUEUE_REG_0__0_ , P2_INSTQUEUERD_ADDR_REG_4_ , P2_INSTQUEUERD_ADDR_REG_3_;
input P2_INSTQUEUERD_ADDR_REG_2_ , P2_INSTQUEUERD_ADDR_REG_1_ , P2_INSTQUEUERD_ADDR_REG_0_ , P2_INSTQUEUEWR_ADDR_REG_4_ , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_INSTQUEUEWR_ADDR_REG_2_;
input P2_INSTQUEUEWR_ADDR_REG_1_ , P2_INSTQUEUEWR_ADDR_REG_0_ , P2_INSTADDRPOINTER_REG_0_ , P2_INSTADDRPOINTER_REG_1_ , P2_INSTADDRPOINTER_REG_2_ , P2_INSTADDRPOINTER_REG_3_;
input P2_INSTADDRPOINTER_REG_4_ , P2_INSTADDRPOINTER_REG_5_ , P2_INSTADDRPOINTER_REG_6_ , P2_INSTADDRPOINTER_REG_7_ , P2_INSTADDRPOINTER_REG_8_ , P2_INSTADDRPOINTER_REG_9_;
input P2_INSTADDRPOINTER_REG_10_ , P2_INSTADDRPOINTER_REG_11_ , P2_INSTADDRPOINTER_REG_12_ , P2_INSTADDRPOINTER_REG_13_ , P2_INSTADDRPOINTER_REG_14_ , P2_INSTADDRPOINTER_REG_15_;
input P2_INSTADDRPOINTER_REG_16_ , P2_INSTADDRPOINTER_REG_17_ , P2_INSTADDRPOINTER_REG_18_ , P2_INSTADDRPOINTER_REG_19_ , P2_INSTADDRPOINTER_REG_20_ , P2_INSTADDRPOINTER_REG_21_;
input P2_INSTADDRPOINTER_REG_22_ , P2_INSTADDRPOINTER_REG_23_ , P2_INSTADDRPOINTER_REG_24_ , P2_INSTADDRPOINTER_REG_25_ , P2_INSTADDRPOINTER_REG_26_ , P2_INSTADDRPOINTER_REG_27_;
input P2_INSTADDRPOINTER_REG_28_ , P2_INSTADDRPOINTER_REG_29_ , P2_INSTADDRPOINTER_REG_30_ , P2_INSTADDRPOINTER_REG_31_ , P2_PHYADDRPOINTER_REG_0_ , P2_PHYADDRPOINTER_REG_1_;
input P2_PHYADDRPOINTER_REG_2_ , P2_PHYADDRPOINTER_REG_3_ , P2_PHYADDRPOINTER_REG_4_ , P2_PHYADDRPOINTER_REG_5_ , P2_PHYADDRPOINTER_REG_6_ , P2_PHYADDRPOINTER_REG_7_;
input P2_PHYADDRPOINTER_REG_8_ , P2_PHYADDRPOINTER_REG_9_ , P2_PHYADDRPOINTER_REG_10_ , P2_PHYADDRPOINTER_REG_11_ , P2_PHYADDRPOINTER_REG_12_ , P2_PHYADDRPOINTER_REG_13_;
input P2_PHYADDRPOINTER_REG_14_ , P2_PHYADDRPOINTER_REG_15_ , P2_PHYADDRPOINTER_REG_16_ , P2_PHYADDRPOINTER_REG_17_ , P2_PHYADDRPOINTER_REG_18_ , P2_PHYADDRPOINTER_REG_19_;
input P2_PHYADDRPOINTER_REG_20_ , P2_PHYADDRPOINTER_REG_21_ , P2_PHYADDRPOINTER_REG_22_ , P2_PHYADDRPOINTER_REG_23_ , P2_PHYADDRPOINTER_REG_24_ , P2_PHYADDRPOINTER_REG_25_;
input P2_PHYADDRPOINTER_REG_26_ , P2_PHYADDRPOINTER_REG_27_ , P2_PHYADDRPOINTER_REG_28_ , P2_PHYADDRPOINTER_REG_29_ , P2_PHYADDRPOINTER_REG_30_ , P2_PHYADDRPOINTER_REG_31_;
input P2_LWORD_REG_15_ , P2_LWORD_REG_14_ , P2_LWORD_REG_13_ , P2_LWORD_REG_12_ , P2_LWORD_REG_11_ , P2_LWORD_REG_10_;
input P2_LWORD_REG_9_ , P2_LWORD_REG_8_ , P2_LWORD_REG_7_ , P2_LWORD_REG_6_ , P2_LWORD_REG_5_ , P2_LWORD_REG_4_;
input P2_LWORD_REG_3_ , P2_LWORD_REG_2_ , P2_LWORD_REG_1_ , P2_LWORD_REG_0_ , P2_UWORD_REG_14_ , P2_UWORD_REG_13_;
input P2_UWORD_REG_12_ , P2_UWORD_REG_11_ , P2_UWORD_REG_10_ , P2_UWORD_REG_9_ , P2_UWORD_REG_8_ , P2_UWORD_REG_7_;
input P2_UWORD_REG_6_ , P2_UWORD_REG_5_ , P2_UWORD_REG_4_ , P2_UWORD_REG_3_ , P2_UWORD_REG_2_ , P2_UWORD_REG_1_;
input P2_UWORD_REG_0_ , P2_DATAO_REG_0_ , P2_DATAO_REG_1_ , P2_DATAO_REG_2_ , P2_DATAO_REG_3_ , P2_DATAO_REG_4_;
input P2_DATAO_REG_5_ , P2_DATAO_REG_6_ , P2_DATAO_REG_7_ , P2_DATAO_REG_8_ , P2_DATAO_REG_9_ , P2_DATAO_REG_10_;
input P2_DATAO_REG_11_ , P2_DATAO_REG_12_ , P2_DATAO_REG_13_ , P2_DATAO_REG_14_ , P2_DATAO_REG_15_ , P2_DATAO_REG_16_;
input P2_DATAO_REG_17_ , P2_DATAO_REG_18_ , P2_DATAO_REG_19_ , P2_DATAO_REG_20_ , P2_DATAO_REG_21_ , P2_DATAO_REG_22_;
input P2_DATAO_REG_23_ , P2_DATAO_REG_24_ , P2_DATAO_REG_25_ , P2_DATAO_REG_26_ , P2_DATAO_REG_27_ , P2_DATAO_REG_28_;
input P2_DATAO_REG_29_ , P2_DATAO_REG_30_ , P2_DATAO_REG_31_ , P2_EAX_REG_0_ , P2_EAX_REG_1_ , P2_EAX_REG_2_;
input P2_EAX_REG_3_ , P2_EAX_REG_4_ , P2_EAX_REG_5_ , P2_EAX_REG_6_ , P2_EAX_REG_7_ , P2_EAX_REG_8_;
input P2_EAX_REG_9_ , P2_EAX_REG_10_ , P2_EAX_REG_11_ , P2_EAX_REG_12_ , P2_EAX_REG_13_ , P2_EAX_REG_14_;
input P2_EAX_REG_15_ , P2_EAX_REG_16_ , P2_EAX_REG_17_ , P2_EAX_REG_18_ , P2_EAX_REG_19_ , P2_EAX_REG_20_;
input P2_EAX_REG_21_ , P2_EAX_REG_22_ , P2_EAX_REG_23_ , P2_EAX_REG_24_ , P2_EAX_REG_25_ , P2_EAX_REG_26_;
input P2_EAX_REG_27_ , P2_EAX_REG_28_ , P2_EAX_REG_29_ , P2_EAX_REG_30_ , P2_EAX_REG_31_ , P2_EBX_REG_0_;
input P2_EBX_REG_1_ , P2_EBX_REG_2_ , P2_EBX_REG_3_ , P2_EBX_REG_4_ , P2_EBX_REG_5_ , P2_EBX_REG_6_;
input P2_EBX_REG_7_ , P2_EBX_REG_8_ , P2_EBX_REG_9_ , P2_EBX_REG_10_ , P2_EBX_REG_11_ , P2_EBX_REG_12_;
input P2_EBX_REG_13_ , P2_EBX_REG_14_ , P2_EBX_REG_15_ , P2_EBX_REG_16_ , P2_EBX_REG_17_ , P2_EBX_REG_18_;
input P2_EBX_REG_19_ , P2_EBX_REG_20_ , P2_EBX_REG_21_ , P2_EBX_REG_22_ , P2_EBX_REG_23_ , P2_EBX_REG_24_;
input P2_EBX_REG_25_ , P2_EBX_REG_26_ , P2_EBX_REG_27_ , P2_EBX_REG_28_ , P2_EBX_REG_29_ , P2_EBX_REG_30_;
input P2_EBX_REG_31_ , P2_REIP_REG_0_ , P2_REIP_REG_1_ , P2_REIP_REG_2_ , P2_REIP_REG_3_ , P2_REIP_REG_4_;
input P2_REIP_REG_5_ , P2_REIP_REG_6_ , P2_REIP_REG_7_ , P2_REIP_REG_8_ , P2_REIP_REG_9_ , P2_REIP_REG_10_;
input P2_REIP_REG_11_ , P2_REIP_REG_12_ , P2_REIP_REG_13_ , P2_REIP_REG_14_ , P2_REIP_REG_15_ , P2_REIP_REG_16_;
input P2_REIP_REG_17_ , P2_REIP_REG_18_ , P2_REIP_REG_19_ , P2_REIP_REG_20_ , P2_REIP_REG_21_ , P2_REIP_REG_22_;
input P2_REIP_REG_23_ , P2_REIP_REG_24_ , P2_REIP_REG_25_ , P2_REIP_REG_26_ , P2_REIP_REG_27_ , P2_REIP_REG_28_;
input P2_REIP_REG_29_ , P2_REIP_REG_30_ , P2_REIP_REG_31_ , P2_BYTEENABLE_REG_3_ , P2_BYTEENABLE_REG_2_ , P2_BYTEENABLE_REG_1_;
input P2_BYTEENABLE_REG_0_ , P2_W_R_N_REG , P2_FLUSH_REG , P2_MORE_REG , P2_STATEBS16_REG , P2_REQUESTPENDING_REG;
input P2_D_C_N_REG , P2_M_IO_N_REG , P2_CODEFETCH_REG , P2_ADS_N_REG , P2_READREQUEST_REG , P2_MEMORYFETCH_REG;
input P1_BE_N_REG_3_ , P1_BE_N_REG_2_ , P1_BE_N_REG_1_ , P1_BE_N_REG_0_ , P1_ADDRESS_REG_29__EXTRA , P1_ADDRESS_REG_28__EXTRA;
input P1_ADDRESS_REG_27__EXTRA , P1_ADDRESS_REG_26__EXTRA , P1_ADDRESS_REG_25__EXTRA , P1_ADDRESS_REG_24__EXTRA , P1_ADDRESS_REG_23__EXTRA , P1_ADDRESS_REG_22__EXTRA;
input P1_ADDRESS_REG_21__EXTRA , P1_ADDRESS_REG_20__EXTRA , P1_ADDRESS_REG_19__EXTRA , P1_ADDRESS_REG_18__EXTRA , P1_ADDRESS_REG_17__EXTRA , P1_ADDRESS_REG_16__EXTRA;
input P1_ADDRESS_REG_15__EXTRA , P1_ADDRESS_REG_14__EXTRA , P1_ADDRESS_REG_13__EXTRA , P1_ADDRESS_REG_12__EXTRA , P1_ADDRESS_REG_11__EXTRA , P1_ADDRESS_REG_10__EXTRA;
input P1_ADDRESS_REG_9__EXTRA , P1_ADDRESS_REG_8__EXTRA , P1_ADDRESS_REG_7__EXTRA , P1_ADDRESS_REG_6__EXTRA , P1_ADDRESS_REG_5__EXTRA , P1_ADDRESS_REG_4__EXTRA;
input P1_ADDRESS_REG_3__EXTRA , P1_ADDRESS_REG_2__EXTRA , P1_ADDRESS_REG_1__EXTRA , P1_ADDRESS_REG_0__EXTRA , P1_STATE_REG_2_ , P1_STATE_REG_1_;
input P1_STATE_REG_0_ , P1_DATAWIDTH_REG_0_ , P1_DATAWIDTH_REG_1_ , P1_DATAWIDTH_REG_2_ , P1_DATAWIDTH_REG_3_ , P1_DATAWIDTH_REG_4_;
input P1_DATAWIDTH_REG_5_ , P1_DATAWIDTH_REG_6_ , P1_DATAWIDTH_REG_7_ , P1_DATAWIDTH_REG_8_ , P1_DATAWIDTH_REG_9_ , P1_DATAWIDTH_REG_10_;
input P1_DATAWIDTH_REG_11_ , P1_DATAWIDTH_REG_12_ , P1_DATAWIDTH_REG_13_ , P1_DATAWIDTH_REG_14_ , P1_DATAWIDTH_REG_15_ , P1_DATAWIDTH_REG_16_;
input P1_DATAWIDTH_REG_17_ , P1_DATAWIDTH_REG_18_ , P1_DATAWIDTH_REG_19_ , P1_DATAWIDTH_REG_20_ , P1_DATAWIDTH_REG_21_ , P1_DATAWIDTH_REG_22_;
input P1_DATAWIDTH_REG_23_ , P1_DATAWIDTH_REG_24_ , P1_DATAWIDTH_REG_25_ , P1_DATAWIDTH_REG_26_ , P1_DATAWIDTH_REG_27_ , P1_DATAWIDTH_REG_28_;
input P1_DATAWIDTH_REG_29_ , P1_DATAWIDTH_REG_30_ , P1_DATAWIDTH_REG_31_ , P1_STATE2_REG_3_ , P1_STATE2_REG_2_ , P1_STATE2_REG_1_;
input P1_STATE2_REG_0_ , P1_INSTQUEUE_REG_15__7_ , P1_INSTQUEUE_REG_15__6_ , P1_INSTQUEUE_REG_15__5_ , P1_INSTQUEUE_REG_15__4_ , P1_INSTQUEUE_REG_15__3_;
input P1_INSTQUEUE_REG_15__2_ , P1_INSTQUEUE_REG_15__1_ , P1_INSTQUEUE_REG_15__0_ , P1_INSTQUEUE_REG_14__7_ , P1_INSTQUEUE_REG_14__6_ , P1_INSTQUEUE_REG_14__5_;
input P1_INSTQUEUE_REG_14__4_ , P1_INSTQUEUE_REG_14__3_ , P1_INSTQUEUE_REG_14__2_ , P1_INSTQUEUE_REG_14__1_ , P1_INSTQUEUE_REG_14__0_ , P1_INSTQUEUE_REG_13__7_;
input P1_INSTQUEUE_REG_13__6_ , P1_INSTQUEUE_REG_13__5_ , P1_INSTQUEUE_REG_13__4_ , P1_INSTQUEUE_REG_13__3_ , P1_INSTQUEUE_REG_13__2_ , P1_INSTQUEUE_REG_13__1_;
input P1_INSTQUEUE_REG_13__0_ , P1_INSTQUEUE_REG_12__7_ , P1_INSTQUEUE_REG_12__6_ , P1_INSTQUEUE_REG_12__5_ , P1_INSTQUEUE_REG_12__4_ , P1_INSTQUEUE_REG_12__3_;
input P1_INSTQUEUE_REG_12__2_ , P1_INSTQUEUE_REG_12__1_ , P1_INSTQUEUE_REG_12__0_ , P1_INSTQUEUE_REG_11__7_ , P1_INSTQUEUE_REG_11__6_ , P1_INSTQUEUE_REG_11__5_;
input P1_INSTQUEUE_REG_11__4_ , P1_INSTQUEUE_REG_11__3_ , P1_INSTQUEUE_REG_11__2_ , P1_INSTQUEUE_REG_11__1_ , P1_INSTQUEUE_REG_11__0_ , P1_INSTQUEUE_REG_10__7_;
input P1_INSTQUEUE_REG_10__6_ , P1_INSTQUEUE_REG_10__5_ , P1_INSTQUEUE_REG_10__4_ , P1_INSTQUEUE_REG_10__3_ , P1_INSTQUEUE_REG_10__2_ , P1_INSTQUEUE_REG_10__1_;
input P1_INSTQUEUE_REG_10__0_ , P1_INSTQUEUE_REG_9__7_ , P1_INSTQUEUE_REG_9__6_ , P1_INSTQUEUE_REG_9__5_ , P1_INSTQUEUE_REG_9__4_ , P1_INSTQUEUE_REG_9__3_;
input P1_INSTQUEUE_REG_9__2_ , P1_INSTQUEUE_REG_9__1_ , P1_INSTQUEUE_REG_9__0_ , P1_INSTQUEUE_REG_8__7_ , P1_INSTQUEUE_REG_8__6_ , P1_INSTQUEUE_REG_8__5_;
input P1_INSTQUEUE_REG_8__4_ , P1_INSTQUEUE_REG_8__3_ , P1_INSTQUEUE_REG_8__2_ , P1_INSTQUEUE_REG_8__1_ , P1_INSTQUEUE_REG_8__0_ , P1_INSTQUEUE_REG_7__7_;
input P1_INSTQUEUE_REG_7__6_ , P1_INSTQUEUE_REG_7__5_ , P1_INSTQUEUE_REG_7__4_ , P1_INSTQUEUE_REG_7__3_ , P1_INSTQUEUE_REG_7__2_ , P1_INSTQUEUE_REG_7__1_;
input P1_INSTQUEUE_REG_7__0_ , P1_INSTQUEUE_REG_6__7_ , P1_INSTQUEUE_REG_6__6_ , P1_INSTQUEUE_REG_6__5_ , P1_INSTQUEUE_REG_6__4_ , P1_INSTQUEUE_REG_6__3_;
input P1_INSTQUEUE_REG_6__2_ , P1_INSTQUEUE_REG_6__1_ , P1_INSTQUEUE_REG_6__0_ , P1_INSTQUEUE_REG_5__7_ , P1_INSTQUEUE_REG_5__6_ , P1_INSTQUEUE_REG_5__5_;
input P1_INSTQUEUE_REG_5__4_ , P1_INSTQUEUE_REG_5__3_ , P1_INSTQUEUE_REG_5__2_ , P1_INSTQUEUE_REG_5__1_ , P1_INSTQUEUE_REG_5__0_ , P1_INSTQUEUE_REG_4__7_;
input P1_INSTQUEUE_REG_4__6_ , P1_INSTQUEUE_REG_4__5_ , P1_INSTQUEUE_REG_4__4_ , P1_INSTQUEUE_REG_4__3_ , P1_INSTQUEUE_REG_4__2_ , P1_INSTQUEUE_REG_4__1_;
input P1_INSTQUEUE_REG_4__0_ , P1_INSTQUEUE_REG_3__7_ , P1_INSTQUEUE_REG_3__6_ , P1_INSTQUEUE_REG_3__5_ , P1_INSTQUEUE_REG_3__4_ , P1_INSTQUEUE_REG_3__3_;
input P1_INSTQUEUE_REG_3__2_ , P1_INSTQUEUE_REG_3__1_ , P1_INSTQUEUE_REG_3__0_ , P1_INSTQUEUE_REG_2__7_ , P1_INSTQUEUE_REG_2__6_ , P1_INSTQUEUE_REG_2__5_;
input P1_INSTQUEUE_REG_2__4_ , P1_INSTQUEUE_REG_2__3_ , P1_INSTQUEUE_REG_2__2_ , P1_INSTQUEUE_REG_2__1_ , P1_INSTQUEUE_REG_2__0_ , P1_INSTQUEUE_REG_1__7_;
input P1_INSTQUEUE_REG_1__6_ , P1_INSTQUEUE_REG_1__5_ , P1_INSTQUEUE_REG_1__4_ , P1_INSTQUEUE_REG_1__3_ , P1_INSTQUEUE_REG_1__2_ , P1_INSTQUEUE_REG_1__1_;
input P1_INSTQUEUE_REG_1__0_ , P1_INSTQUEUE_REG_0__7_ , P1_INSTQUEUE_REG_0__6_ , P1_INSTQUEUE_REG_0__5_ , P1_INSTQUEUE_REG_0__4_ , P1_INSTQUEUE_REG_0__3_;
input P1_INSTQUEUE_REG_0__2_ , P1_INSTQUEUE_REG_0__1_ , P1_INSTQUEUE_REG_0__0_ , P1_INSTQUEUERD_ADDR_REG_4_ , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_2_;
input P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUEWR_ADDR_REG_4_ , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_INSTQUEUEWR_ADDR_REG_1_;
input P1_INSTQUEUEWR_ADDR_REG_0_ , P1_INSTADDRPOINTER_REG_0_ , P1_INSTADDRPOINTER_REG_1_ , P1_INSTADDRPOINTER_REG_2_ , P1_INSTADDRPOINTER_REG_3_ , P1_INSTADDRPOINTER_REG_4_;
input P1_INSTADDRPOINTER_REG_5_ , P1_INSTADDRPOINTER_REG_6_ , P1_INSTADDRPOINTER_REG_7_ , P1_INSTADDRPOINTER_REG_8_ , P1_INSTADDRPOINTER_REG_9_ , P1_INSTADDRPOINTER_REG_10_;
input P1_INSTADDRPOINTER_REG_11_ , P1_INSTADDRPOINTER_REG_12_ , P1_INSTADDRPOINTER_REG_13_ , P1_INSTADDRPOINTER_REG_14_ , P1_INSTADDRPOINTER_REG_15_ , P1_INSTADDRPOINTER_REG_16_;
input P1_INSTADDRPOINTER_REG_17_ , P1_INSTADDRPOINTER_REG_18_ , P1_INSTADDRPOINTER_REG_19_ , P1_INSTADDRPOINTER_REG_20_ , P1_INSTADDRPOINTER_REG_21_ , P1_INSTADDRPOINTER_REG_22_;
input P1_INSTADDRPOINTER_REG_23_ , P1_INSTADDRPOINTER_REG_24_ , P1_INSTADDRPOINTER_REG_25_ , P1_INSTADDRPOINTER_REG_26_ , P1_INSTADDRPOINTER_REG_27_ , P1_INSTADDRPOINTER_REG_28_;
input P1_INSTADDRPOINTER_REG_29_ , P1_INSTADDRPOINTER_REG_30_ , P1_INSTADDRPOINTER_REG_31_ , P1_PHYADDRPOINTER_REG_0_ , P1_PHYADDRPOINTER_REG_1_ , P1_PHYADDRPOINTER_REG_2_;
input P1_PHYADDRPOINTER_REG_3_ , P1_PHYADDRPOINTER_REG_4_ , P1_PHYADDRPOINTER_REG_5_ , P1_PHYADDRPOINTER_REG_6_ , P1_PHYADDRPOINTER_REG_7_ , P1_PHYADDRPOINTER_REG_8_;
input P1_PHYADDRPOINTER_REG_9_ , P1_PHYADDRPOINTER_REG_10_ , P1_PHYADDRPOINTER_REG_11_ , P1_PHYADDRPOINTER_REG_12_ , P1_PHYADDRPOINTER_REG_13_ , P1_PHYADDRPOINTER_REG_14_;
input P1_PHYADDRPOINTER_REG_15_ , P1_PHYADDRPOINTER_REG_16_ , P1_PHYADDRPOINTER_REG_17_ , P1_PHYADDRPOINTER_REG_18_ , P1_PHYADDRPOINTER_REG_19_ , P1_PHYADDRPOINTER_REG_20_;
input P1_PHYADDRPOINTER_REG_21_ , P1_PHYADDRPOINTER_REG_22_ , P1_PHYADDRPOINTER_REG_23_ , P1_PHYADDRPOINTER_REG_24_ , P1_PHYADDRPOINTER_REG_25_ , P1_PHYADDRPOINTER_REG_26_;
input P1_PHYADDRPOINTER_REG_27_ , P1_PHYADDRPOINTER_REG_28_ , P1_PHYADDRPOINTER_REG_29_ , P1_PHYADDRPOINTER_REG_30_ , P1_PHYADDRPOINTER_REG_31_ , P1_LWORD_REG_15_;
input P1_LWORD_REG_14_ , P1_LWORD_REG_13_ , P1_LWORD_REG_12_ , P1_LWORD_REG_11_ , P1_LWORD_REG_10_ , P1_LWORD_REG_9_;
input P1_LWORD_REG_8_ , P1_LWORD_REG_7_ , P1_LWORD_REG_6_ , P1_LWORD_REG_5_ , P1_LWORD_REG_4_ , P1_LWORD_REG_3_;
input P1_LWORD_REG_2_ , P1_LWORD_REG_1_ , P1_LWORD_REG_0_ , P1_UWORD_REG_14_ , P1_UWORD_REG_13_ , P1_UWORD_REG_12_;
input P1_UWORD_REG_11_ , P1_UWORD_REG_10_ , P1_UWORD_REG_9_ , P1_UWORD_REG_8_ , P1_UWORD_REG_7_ , P1_UWORD_REG_6_;
input P1_UWORD_REG_5_ , P1_UWORD_REG_4_ , P1_UWORD_REG_3_ , P1_UWORD_REG_2_ , P1_UWORD_REG_1_ , P1_UWORD_REG_0_;
input P1_DATAO_REG_0_ , P1_DATAO_REG_1_ , P1_DATAO_REG_2_ , P1_DATAO_REG_3_ , P1_DATAO_REG_4_ , P1_DATAO_REG_5_;
input P1_DATAO_REG_6_ , P1_DATAO_REG_7_ , P1_DATAO_REG_8_ , P1_DATAO_REG_9_ , P1_DATAO_REG_10_ , P1_DATAO_REG_11_;
input P1_DATAO_REG_12_ , P1_DATAO_REG_13_ , P1_DATAO_REG_14_ , P1_DATAO_REG_15_ , P1_DATAO_REG_16_ , P1_DATAO_REG_17_;
input P1_DATAO_REG_18_ , P1_DATAO_REG_19_ , P1_DATAO_REG_20_ , P1_DATAO_REG_21_ , P1_DATAO_REG_22_ , P1_DATAO_REG_23_;
input P1_DATAO_REG_24_ , P1_DATAO_REG_25_ , P1_DATAO_REG_26_ , P1_DATAO_REG_27_ , P1_DATAO_REG_28_ , P1_DATAO_REG_29_;
input P1_DATAO_REG_30_ , P1_DATAO_REG_31_ , P1_EAX_REG_0_ , P1_EAX_REG_1_ , P1_EAX_REG_2_ , P1_EAX_REG_3_;
input P1_EAX_REG_4_ , P1_EAX_REG_5_ , P1_EAX_REG_6_ , P1_EAX_REG_7_ , P1_EAX_REG_8_ , P1_EAX_REG_9_;
input P1_EAX_REG_10_ , P1_EAX_REG_11_ , P1_EAX_REG_12_ , P1_EAX_REG_13_ , P1_EAX_REG_14_ , P1_EAX_REG_15_;
input P1_EAX_REG_16_ , P1_EAX_REG_17_ , P1_EAX_REG_18_ , P1_EAX_REG_19_ , P1_EAX_REG_20_ , P1_EAX_REG_21_;
input P1_EAX_REG_22_ , P1_EAX_REG_23_ , P1_EAX_REG_24_ , P1_EAX_REG_25_ , P1_EAX_REG_26_ , P1_EAX_REG_27_;
input P1_EAX_REG_28_ , P1_EAX_REG_29_ , P1_EAX_REG_30_ , P1_EAX_REG_31_ , P1_EBX_REG_0_ , P1_EBX_REG_1_;
input P1_EBX_REG_2_ , P1_EBX_REG_3_ , P1_EBX_REG_4_ , P1_EBX_REG_5_ , P1_EBX_REG_6_ , P1_EBX_REG_7_;
input P1_EBX_REG_8_ , P1_EBX_REG_9_ , P1_EBX_REG_10_ , P1_EBX_REG_11_ , P1_EBX_REG_12_ , P1_EBX_REG_13_;
input P1_EBX_REG_14_ , P1_EBX_REG_15_ , P1_EBX_REG_16_ , P1_EBX_REG_17_ , P1_EBX_REG_18_ , P1_EBX_REG_19_;
input P1_EBX_REG_20_ , P1_EBX_REG_21_ , P1_EBX_REG_22_ , P1_EBX_REG_23_ , P1_EBX_REG_24_ , P1_EBX_REG_25_;
input P1_EBX_REG_26_ , P1_EBX_REG_27_ , P1_EBX_REG_28_ , P1_EBX_REG_29_ , P1_EBX_REG_30_ , P1_EBX_REG_31_;
input P1_REIP_REG_0_ , P1_REIP_REG_1_ , P1_REIP_REG_2_ , P1_REIP_REG_3_ , P1_REIP_REG_4_ , P1_REIP_REG_5_;
input P1_REIP_REG_6_ , P1_REIP_REG_7_ , P1_REIP_REG_8_ , P1_REIP_REG_9_ , P1_REIP_REG_10_ , P1_REIP_REG_11_;
input P1_REIP_REG_12_ , P1_REIP_REG_13_ , P1_REIP_REG_14_ , P1_REIP_REG_15_ , P1_REIP_REG_16_ , P1_REIP_REG_17_;
input P1_REIP_REG_18_ , P1_REIP_REG_19_ , P1_REIP_REG_20_ , P1_REIP_REG_21_ , P1_REIP_REG_22_ , P1_REIP_REG_23_;
input P1_REIP_REG_24_ , P1_REIP_REG_25_ , P1_REIP_REG_26_ , P1_REIP_REG_27_ , P1_REIP_REG_28_ , P1_REIP_REG_29_;
input P1_REIP_REG_30_ , P1_REIP_REG_31_ , P1_BYTEENABLE_REG_3_ , P1_BYTEENABLE_REG_2_ , P1_BYTEENABLE_REG_1_ , P1_BYTEENABLE_REG_0_;
input P1_W_R_N_REG , P1_FLUSH_REG , P1_MORE_REG , P1_STATEBS16_REG , P1_REQUESTPENDING_REG , P1_D_C_N_REG;
input P1_M_IO_N_REG , P1_CODEFETCH_REG , P1_ADS_N_REG_EXTRA , P1_READREQUEST_REG , P1_MEMORYFETCH_REG;

wire P1_ADD_515_U182 , P1_ADD_515_U181 , P1_ADD_515_U180 , U207 , U208 , U209 , U210 , U211 , U248 , U249;
wire U250 , U283 , U284 , U285 , U286 , U287 , U288 , U289 , U290 , U291;
wire U292 , U293 , U294 , U295 , U296 , U297 , U298 , U299 , U300 , U301;
wire U302 , U303 , U304 , U305 , U306 , U307 , U308 , U309 , U310 , U311;
wire U312 , U313 , U314 , U315 , U316 , U317 , U318 , U319 , U320 , U321;
wire U322 , U323 , U324 , U325 , U326 , U327 , U328 , U329 , U330 , U331;
wire U332 , U333 , U334 , U335 , U336 , U337 , U338 , U339 , U340 , U341;
wire U342 , U343 , U344 , U345 , U346 , U377 , U378 , U379 , U380 , U381;
wire U382 , U383 , U384 , U385 , U386 , U387 , U388 , U389 , U390 , U391;
wire U392 , U393 , U394 , U395 , U396 , U397 , U398 , U399 , U400 , U401;
wire U402 , U403 , U404 , U405 , U406 , U407 , U408 , U409 , U410 , U411;
wire U412 , U413 , U414 , U415 , U416 , U417 , U418 , U419 , U420 , U421;
wire U422 , U423 , U424 , U425 , U426 , U427 , U428 , U429 , U430 , U431;
wire U432 , U433 , U434 , U435 , U436 , U437 , U438 , U439 , U440 , U441;
wire U442 , U443 , U444 , U445 , U446 , U447 , U448 , U449 , U450 , U451;
wire U452 , U453 , U454 , U455 , U456 , U457 , U458 , U459 , U460 , U461;
wire U462 , U463 , U464 , U465 , U466 , U467 , U468 , U469 , U470 , U471;
wire U472 , U473 , U474 , U475 , U476 , U477 , U478 , U479 , U480 , U481;
wire U482 , U483 , U484 , U485 , U486 , U487 , U488 , U489 , U490 , U491;
wire U492 , U493 , U494 , U495 , U496 , U497 , U498 , U499 , U500 , U501;
wire U502 , U503 , U504 , U505 , U506 , U507 , U508 , U509 , U510 , U511;
wire U512 , U513 , U514 , U515 , U516 , U517 , U518 , U519 , U520 , U521;
wire U522 , U523 , U524 , U525 , U526 , U527 , U528 , U529 , U530 , U531;
wire U532 , U533 , U534 , U535 , U536 , U537 , U538 , U539 , U540 , U541;
wire U542 , U543 , U544 , U545 , U546 , U547 , U548 , U549 , U550 , U551;
wire U552 , U553 , U554 , U555 , U556 , U557 , U558 , U559 , U560 , U561;
wire U562 , U563 , U564 , U565 , U566 , U567 , U568 , U569 , U570 , U571;
wire U572 , U573 , U574 , U575 , U576 , U577 , U578 , U579 , U580 , U581;
wire U582 , U583 , U584 , U585 , U586 , U587 , U588 , U589 , U590 , U591;
wire U592 , U593 , U594 , U595 , U596 , U597 , U598 , U599 , U600 , U601;
wire U602 , U603 , U604 , U605 , U606 , U607 , U608 , U609 , U610 , U611;
wire U612 , U613 , U614 , U615 , U616 , U617 , U618 , U619 , U620 , U621;
wire U622 , U623 , U624 , U625 , U626 , U627 , U628 , U629 , U630 , U631;
wire U632 , U633 , U634 , U635 , U636 , U637 , U638 , U639 , U640 , U641;
wire U642 , U643 , U644 , U645 , U646 , U647 , U648 , U649 , U650 , U651;
wire U652 , U653 , U654 , U655 , U656 , U657 , U658 , U659 , U660 , U661;
wire U662 , U663 , U664 , U665 , U666 , U667 , U668 , U669 , U670 , U671;
wire U672 , U673 , U674 , U675 , U676 , U677 , U678 , U679 , U680 , U681;
wire U682 , U683 , U684 , U685 , U686 , U687 , U688 , U689 , U690 , U691;
wire U692 , U693 , U694 , U695 , U696 , U697 , U698 , U699 , U700 , U701;
wire U702 , U703 , U704 , U705 , U706 , U707 , U708 , U709 , U710 , U711;
wire U712 , U713 , U714 , U715 , U716 , U717 , U718 , U719 , U720 , U721;
wire U722 , U723 , U724 , U725 , U726 , U727 , U728 , U729 , U730 , U731;
wire U732 , U733 , U734 , U735 , U736 , P1_ADD_515_U179 , P1_ADD_515_U178 , P1_ADD_515_U177 , P1_ADD_515_U176 , P1_ADD_515_U175;
wire P1_ADD_515_U174 , P1_ADD_515_U173 , P1_ADD_515_U172 , P1_ADD_515_U171 , P3_U2352 , P3_U2353 , P3_U2354 , P3_U2355 , P3_U2356 , P3_U2357;
wire P3_U2358 , P3_U2359 , P3_U2360 , P3_U2361 , P3_U2362 , P3_U2363 , P3_U2364 , P3_U2365 , P3_U2366 , P3_U2367;
wire P3_U2368 , P3_U2369 , P3_U2370 , P3_U2371 , P3_U2372 , P3_U2373 , P3_U2374 , P3_U2375 , P3_U2376 , P3_U2377;
wire P3_U2378 , P3_U2379 , P3_U2380 , P3_U2381 , P3_U2382 , P3_U2383 , P3_U2384 , P3_U2385 , P3_U2386 , P3_U2387;
wire P3_U2388 , P3_U2389 , P3_U2390 , P3_U2391 , P3_U2392 , P3_U2393 , P3_U2394 , P3_U2395 , P3_U2396 , P3_U2397;
wire P3_U2398 , P3_U2399 , P3_U2400 , P3_U2401 , P3_U2402 , P3_U2403 , P3_U2404 , P3_U2405 , P3_U2406 , P3_U2407;
wire P3_U2408 , P3_U2409 , P3_U2410 , P3_U2411 , P3_U2412 , P3_U2413 , P3_U2414 , P3_U2415 , P3_U2416 , P3_U2417;
wire P3_U2418 , P3_U2419 , P3_U2420 , P3_U2421 , P3_U2422 , P3_U2423 , P3_U2424 , P3_U2425 , P3_U2426 , P3_U2427;
wire P3_U2428 , P3_U2429 , P3_U2430 , P3_U2431 , P3_U2432 , P3_U2433 , P3_U2434 , P3_U2435 , P3_U2436 , P3_U2437;
wire P3_U2438 , P3_U2439 , P3_U2440 , P3_U2441 , P3_U2442 , P3_U2443 , P3_U2444 , P3_U2445 , P3_U2446 , P3_U2447;
wire P3_U2448 , P3_U2449 , P3_U2450 , P3_U2451 , P3_U2452 , P3_U2453 , P3_U2454 , P3_U2455 , P3_U2456 , P3_U2457;
wire P3_U2458 , P3_U2459 , P3_U2460 , P3_U2461 , P3_U2462 , P3_U2463 , P3_U2464 , P3_U2465 , P3_U2466 , P3_U2467;
wire P3_U2468 , P3_U2469 , P3_U2470 , P3_U2471 , P3_U2472 , P3_U2473 , P3_U2474 , P3_U2475 , P3_U2476 , P3_U2477;
wire P3_U2478 , P3_U2479 , P3_U2480 , P3_U2481 , P3_U2482 , P3_U2483 , P3_U2484 , P3_U2485 , P3_U2486 , P3_U2487;
wire P3_U2488 , P3_U2489 , P3_U2490 , P3_U2491 , P3_U2492 , P3_U2493 , P3_U2494 , P3_U2495 , P3_U2496 , P3_U2497;
wire P3_U2498 , P3_U2499 , P3_U2500 , P3_U2501 , P3_U2502 , P3_U2503 , P3_U2504 , P3_U2505 , P3_U2506 , P3_U2507;
wire P3_U2508 , P3_U2509 , P3_U2510 , P3_U2511 , P3_U2512 , P3_U2513 , P3_U2514 , P3_U2515 , P3_U2516 , P3_U2517;
wire P3_U2518 , P3_U2519 , P3_U2520 , P3_U2521 , P3_U2522 , P3_U2523 , P3_U2524 , P3_U2525 , P3_U2526 , P3_U2527;
wire P3_U2528 , P3_U2529 , P3_U2530 , P3_U2531 , P3_U2532 , P3_U2533 , P3_U2534 , P3_U2535 , P3_U2536 , P3_U2537;
wire P3_U2538 , P3_U2539 , P3_U2540 , P3_U2541 , P3_U2542 , P3_U2543 , P3_U2544 , P3_U2545 , P3_U2546 , P3_U2547;
wire P3_U2548 , P3_U2549 , P3_U2550 , P3_U2551 , P3_U2552 , P3_U2553 , P3_U2554 , P3_U2555 , P3_U2556 , P3_U2557;
wire P3_U2558 , P3_U2559 , P3_U2560 , P3_U2561 , P3_U2562 , P3_U2563 , P3_U2564 , P3_U2565 , P3_U2566 , P3_U2567;
wire P3_U2568 , P3_U2569 , P3_U2570 , P3_U2571 , P3_U2572 , P3_U2573 , P3_U2574 , P3_U2575 , P3_U2576 , P3_U2577;
wire P3_U2578 , P3_U2579 , P3_U2580 , P3_U2581 , P3_U2582 , P3_U2583 , P3_U2584 , P3_U2585 , P3_U2586 , P3_U2587;
wire P3_U2588 , P3_U2589 , P3_U2590 , P3_U2591 , P3_U2592 , P3_U2593 , P3_U2594 , P3_U2595 , P3_U2596 , P3_U2597;
wire P3_U2598 , P3_U2599 , P3_U2600 , P3_U2601 , P3_U2602 , P3_U2603 , P3_U2604 , P3_U2605 , P3_U2606 , P3_U2607;
wire P3_U2608 , P3_U2609 , P3_U2610 , P3_U2611 , P3_U2612 , P3_U2613 , P3_U2614 , P3_U2615 , P3_U2616 , P3_U2617;
wire P3_U2618 , P3_U2619 , P3_U2620 , P3_U2621 , P3_U2622 , P3_U2623 , P3_U2624 , P3_U2625 , P3_U2626 , P3_U2627;
wire P3_U2628 , P3_U2629 , P3_U2630 , P3_U2631 , P3_U2632 , P3_U3062 , P3_U3063 , P3_U3064 , P3_U3065 , P3_U3066;
wire P3_U3067 , P3_U3068 , P3_U3069 , P3_U3070 , P3_U3071 , P3_U3072 , P3_U3073 , P3_U3074 , P3_U3075 , P3_U3076;
wire P3_U3077 , P3_U3078 , P3_U3079 , P3_U3080 , P3_U3081 , P3_U3082 , P3_U3083 , P3_U3084 , P3_U3085 , P3_U3086;
wire P3_U3087 , P3_U3088 , P3_U3089 , P3_U3090 , P3_U3091 , P3_U3092 , P3_U3093 , P3_U3094 , P3_U3095 , P3_U3096;
wire P3_U3097 , P3_U3098 , P3_U3099 , P3_U3100 , P3_U3101 , P3_U3102 , P3_U3103 , P3_U3104 , P3_U3105 , P3_U3106;
wire P3_U3107 , P3_U3108 , P3_U3109 , P3_U3110 , P3_U3111 , P3_U3112 , P3_U3113 , P3_U3114 , P3_U3115 , P3_U3116;
wire P3_U3117 , P3_U3118 , P3_U3119 , P3_U3120 , P3_U3121 , P3_U3122 , P3_U3123 , P3_U3124 , P3_U3125 , P3_U3126;
wire P3_U3127 , P3_U3128 , P3_U3129 , P3_U3130 , P3_U3131 , P3_U3132 , P3_U3133 , P3_U3134 , P3_U3135 , P3_U3136;
wire P3_U3137 , P3_U3138 , P3_U3139 , P3_U3140 , P3_U3141 , P3_U3142 , P3_U3143 , P3_U3144 , P3_U3145 , P3_U3146;
wire P3_U3147 , P3_U3148 , P3_U3149 , P3_U3150 , P3_U3151 , P3_U3152 , P3_U3153 , P3_U3154 , P3_U3155 , P3_U3156;
wire P3_U3157 , P3_U3158 , P3_U3159 , P3_U3160 , P3_U3161 , P3_U3162 , P3_U3163 , P3_U3164 , P3_U3165 , P3_U3166;
wire P3_U3167 , P3_U3168 , P3_U3169 , P3_U3170 , P3_U3171 , P3_U3172 , P3_U3173 , P3_U3174 , P3_U3175 , P3_U3176;
wire P3_U3177 , P3_U3178 , P3_U3179 , P3_U3180 , P3_U3181 , P3_U3182 , P3_U3183 , P3_U3184 , P3_U3185 , P3_U3186;
wire P3_U3187 , P3_U3188 , P3_U3189 , P3_U3190 , P3_U3191 , P3_U3192 , P3_U3193 , P3_U3194 , P3_U3195 , P3_U3196;
wire P3_U3197 , P3_U3198 , P3_U3199 , P3_U3200 , P3_U3201 , P3_U3202 , P3_U3203 , P3_U3204 , P3_U3205 , P3_U3206;
wire P3_U3207 , P3_U3208 , P3_U3209 , P3_U3210 , P3_U3211 , P3_U3212 , P3_U3213 , P3_U3214 , P3_U3215 , P3_U3216;
wire P3_U3217 , P3_U3218 , P3_U3219 , P3_U3220 , P3_U3221 , P3_U3222 , P3_U3223 , P3_U3224 , P3_U3225 , P3_U3226;
wire P3_U3227 , P3_U3228 , P3_U3229 , P3_U3230 , P3_U3231 , P3_U3232 , P3_U3233 , P3_U3234 , P3_U3235 , P3_U3236;
wire P3_U3237 , P3_U3238 , P3_U3239 , P3_U3240 , P3_U3241 , P3_U3242 , P3_U3243 , P3_U3244 , P3_U3245 , P3_U3246;
wire P3_U3247 , P3_U3248 , P3_U3249 , P3_U3250 , P3_U3251 , P3_U3252 , P3_U3253 , P3_U3254 , P3_U3255 , P3_U3256;
wire P3_U3257 , P3_U3258 , P3_U3259 , P3_U3260 , P3_U3261 , P3_U3262 , P3_U3263 , P3_U3264 , P3_U3265 , P3_U3266;
wire P3_U3267 , P3_U3268 , P3_U3269 , P3_U3270 , P3_U3271 , P3_U3272 , P3_U3273 , P3_U3278 , P3_U3279 , P3_U3283;
wire P3_U3286 , P3_U3287 , P3_U3291 , P3_U3300 , P3_U3301 , P3_U3302 , P3_U3303 , P3_U3304 , P3_U3305 , P3_U3306;
wire P3_U3307 , P3_U3308 , P3_U3309 , P3_U3310 , P3_U3311 , P3_U3312 , P3_U3313 , P3_U3314 , P3_U3315 , P3_U3316;
wire P3_U3317 , P3_U3318 , P3_U3319 , P3_U3320 , P3_U3321 , P3_U3322 , P3_U3323 , P3_U3324 , P3_U3325 , P3_U3326;
wire P3_U3327 , P3_U3328 , P3_U3329 , P3_U3330 , P3_U3331 , P3_U3332 , P3_U3333 , P3_U3334 , P3_U3335 , P3_U3336;
wire P3_U3337 , P3_U3338 , P3_U3339 , P3_U3340 , P3_U3341 , P3_U3342 , P3_U3343 , P3_U3344 , P3_U3345 , P3_U3346;
wire P3_U3347 , P3_U3348 , P3_U3349 , P3_U3350 , P3_U3351 , P3_U3352 , P3_U3353 , P3_U3354 , P3_U3355 , P3_U3356;
wire P3_U3357 , P3_U3358 , P3_U3359 , P3_U3360 , P3_U3361 , P3_U3362 , P3_U3363 , P3_U3364 , P3_U3365 , P3_U3366;
wire P3_U3367 , P3_U3368 , P3_U3369 , P3_U3370 , P3_U3371 , P3_U3372 , P3_U3373 , P3_U3374 , P3_U3375 , P3_U3376;
wire P3_U3377 , P3_U3378 , P3_U3379 , P3_U3380 , P3_U3381 , P3_U3382 , P3_U3383 , P3_U3384 , P3_U3385 , P3_U3386;
wire P3_U3387 , P3_U3388 , P3_U3389 , P3_U3390 , P3_U3391 , P3_U3392 , P3_U3393 , P3_U3394 , P3_U3395 , P3_U3396;
wire P3_U3397 , P3_U3398 , P3_U3399 , P3_U3400 , P3_U3401 , P3_U3402 , P3_U3403 , P3_U3404 , P3_U3405 , P3_U3406;
wire P3_U3407 , P3_U3408 , P3_U3409 , P3_U3410 , P3_U3411 , P3_U3412 , P3_U3413 , P3_U3414 , P3_U3415 , P3_U3416;
wire P3_U3417 , P3_U3418 , P3_U3419 , P3_U3420 , P3_U3421 , P3_U3422 , P3_U3423 , P3_U3424 , P3_U3425 , P3_U3426;
wire P3_U3427 , P3_U3428 , P3_U3429 , P3_U3430 , P3_U3431 , P3_U3432 , P3_U3433 , P3_U3434 , P3_U3435 , P3_U3436;
wire P3_U3437 , P3_U3438 , P3_U3439 , P3_U3440 , P3_U3441 , P3_U3442 , P3_U3443 , P3_U3444 , P3_U3445 , P3_U3446;
wire P3_U3447 , P3_U3448 , P3_U3449 , P3_U3450 , P3_U3451 , P3_U3452 , P3_U3453 , P3_U3454 , P3_U3455 , P3_U3456;
wire P3_U3457 , P3_U3458 , P3_U3459 , P3_U3460 , P3_U3461 , P3_U3462 , P3_U3463 , P3_U3464 , P3_U3465 , P3_U3466;
wire P3_U3467 , P3_U3468 , P3_U3469 , P3_U3470 , P3_U3471 , P3_U3472 , P3_U3473 , P3_U3474 , P3_U3475 , P3_U3476;
wire P3_U3477 , P3_U3478 , P3_U3479 , P3_U3480 , P3_U3481 , P3_U3482 , P3_U3483 , P3_U3484 , P3_U3485 , P3_U3486;
wire P3_U3487 , P3_U3488 , P3_U3489 , P3_U3490 , P3_U3491 , P3_U3492 , P3_U3493 , P3_U3494 , P3_U3495 , P3_U3496;
wire P3_U3497 , P3_U3498 , P3_U3499 , P3_U3500 , P3_U3501 , P3_U3502 , P3_U3503 , P3_U3504 , P3_U3505 , P3_U3506;
wire P3_U3507 , P3_U3508 , P3_U3509 , P3_U3510 , P3_U3511 , P3_U3512 , P3_U3513 , P3_U3514 , P3_U3515 , P3_U3516;
wire P3_U3517 , P3_U3518 , P3_U3519 , P3_U3520 , P3_U3521 , P3_U3522 , P3_U3523 , P3_U3524 , P3_U3525 , P3_U3526;
wire P3_U3527 , P3_U3528 , P3_U3529 , P3_U3530 , P3_U3531 , P3_U3532 , P3_U3533 , P3_U3534 , P3_U3535 , P3_U3536;
wire P3_U3537 , P3_U3538 , P3_U3539 , P3_U3540 , P3_U3541 , P3_U3542 , P3_U3543 , P3_U3544 , P3_U3545 , P3_U3546;
wire P3_U3547 , P3_U3548 , P3_U3549 , P3_U3550 , P3_U3551 , P3_U3552 , P3_U3553 , P3_U3554 , P3_U3555 , P3_U3556;
wire P3_U3557 , P3_U3558 , P3_U3559 , P3_U3560 , P3_U3561 , P3_U3562 , P3_U3563 , P3_U3564 , P3_U3565 , P3_U3566;
wire P3_U3567 , P3_U3568 , P3_U3569 , P3_U3570 , P3_U3571 , P3_U3572 , P3_U3573 , P3_U3574 , P3_U3575 , P3_U3576;
wire P3_U3577 , P3_U3578 , P3_U3579 , P3_U3580 , P3_U3581 , P3_U3582 , P3_U3583 , P3_U3584 , P3_U3585 , P3_U3586;
wire P3_U3587 , P3_U3588 , P3_U3589 , P3_U3590 , P3_U3591 , P3_U3592 , P3_U3593 , P3_U3594 , P3_U3595 , P3_U3596;
wire P3_U3597 , P3_U3598 , P3_U3599 , P3_U3600 , P3_U3601 , P3_U3602 , P3_U3603 , P3_U3604 , P3_U3605 , P3_U3606;
wire P3_U3607 , P3_U3608 , P3_U3609 , P3_U3610 , P3_U3611 , P3_U3612 , P3_U3613 , P3_U3614 , P3_U3615 , P3_U3616;
wire P3_U3617 , P3_U3618 , P3_U3619 , P3_U3620 , P3_U3621 , P3_U3622 , P3_U3623 , P3_U3624 , P3_U3625 , P3_U3626;
wire P3_U3627 , P3_U3628 , P3_U3629 , P3_U3630 , P3_U3631 , P3_U3632 , P3_U3633 , P3_U3634 , P3_U3635 , P3_U3636;
wire P3_U3637 , P3_U3638 , P3_U3639 , P3_U3640 , P3_U3641 , P3_U3642 , P3_U3643 , P3_U3644 , P3_U3645 , P3_U3646;
wire P3_U3647 , P3_U3648 , P3_U3649 , P3_U3650 , P3_U3651 , P3_U3652 , P3_U3653 , P3_U3654 , P3_U3655 , P3_U3656;
wire P3_U3657 , P3_U3658 , P3_U3659 , P3_U3660 , P3_U3661 , P3_U3662 , P3_U3663 , P3_U3664 , P3_U3665 , P3_U3666;
wire P3_U3667 , P3_U3668 , P3_U3669 , P3_U3670 , P3_U3671 , P3_U3672 , P3_U3673 , P3_U3674 , P3_U3675 , P3_U3676;
wire P3_U3677 , P3_U3678 , P3_U3679 , P3_U3680 , P3_U3681 , P3_U3682 , P3_U3683 , P3_U3684 , P3_U3685 , P3_U3686;
wire P3_U3687 , P3_U3688 , P3_U3689 , P3_U3690 , P3_U3691 , P3_U3692 , P3_U3693 , P3_U3694 , P3_U3695 , P3_U3696;
wire P3_U3697 , P3_U3698 , P3_U3699 , P3_U3700 , P3_U3701 , P3_U3702 , P3_U3703 , P3_U3704 , P3_U3705 , P3_U3706;
wire P3_U3707 , P3_U3708 , P3_U3709 , P3_U3710 , P3_U3711 , P3_U3712 , P3_U3713 , P3_U3714 , P3_U3715 , P3_U3716;
wire P3_U3717 , P3_U3718 , P3_U3719 , P3_U3720 , P3_U3721 , P3_U3722 , P3_U3723 , P3_U3724 , P3_U3725 , P3_U3726;
wire P3_U3727 , P3_U3728 , P3_U3729 , P3_U3730 , P3_U3731 , P3_U3732 , P3_U3733 , P3_U3734 , P3_U3735 , P3_U3736;
wire P3_U3737 , P3_U3738 , P3_U3739 , P3_U3740 , P3_U3741 , P3_U3742 , P3_U3743 , P3_U3744 , P3_U3745 , P3_U3746;
wire P3_U3747 , P3_U3748 , P3_U3749 , P3_U3750 , P3_U3751 , P3_U3752 , P3_U3753 , P3_U3754 , P3_U3755 , P3_U3756;
wire P3_U3757 , P3_U3758 , P3_U3759 , P3_U3760 , P3_U3761 , P3_U3762 , P3_U3763 , P3_U3764 , P3_U3765 , P3_U3766;
wire P3_U3767 , P3_U3768 , P3_U3769 , P3_U3770 , P3_U3771 , P3_U3772 , P3_U3773 , P3_U3774 , P3_U3775 , P3_U3776;
wire P3_U3777 , P3_U3778 , P3_U3779 , P3_U3780 , P3_U3781 , P3_U3782 , P3_U3783 , P3_U3784 , P3_U3785 , P3_U3786;
wire P3_U3787 , P3_U3788 , P3_U3789 , P3_U3790 , P3_U3791 , P3_U3792 , P3_U3793 , P3_U3794 , P3_U3795 , P3_U3796;
wire P3_U3797 , P3_U3798 , P3_U3799 , P3_U3800 , P3_U3801 , P3_U3802 , P3_U3803 , P3_U3804 , P3_U3805 , P3_U3806;
wire P3_U3807 , P3_U3808 , P3_U3809 , P3_U3810 , P3_U3811 , P3_U3812 , P3_U3813 , P3_U3814 , P3_U3815 , P3_U3816;
wire P3_U3817 , P3_U3818 , P3_U3819 , P3_U3820 , P3_U3821 , P3_U3822 , P3_U3823 , P3_U3824 , P3_U3825 , P3_U3826;
wire P3_U3827 , P3_U3828 , P3_U3829 , P3_U3830 , P3_U3831 , P3_U3832 , P3_U3833 , P3_U3834 , P3_U3835 , P3_U3836;
wire P3_U3837 , P3_U3838 , P3_U3839 , P3_U3840 , P3_U3841 , P3_U3842 , P3_U3843 , P3_U3844 , P3_U3845 , P3_U3846;
wire P3_U3847 , P3_U3848 , P3_U3849 , P3_U3850 , P3_U3851 , P3_U3852 , P3_U3853 , P3_U3854 , P3_U3855 , P3_U3856;
wire P3_U3857 , P3_U3858 , P3_U3859 , P3_U3860 , P3_U3861 , P3_U3862 , P3_U3863 , P3_U3864 , P3_U3865 , P3_U3866;
wire P3_U3867 , P3_U3868 , P3_U3869 , P3_U3870 , P3_U3871 , P3_U3872 , P3_U3873 , P3_U3874 , P3_U3875 , P3_U3876;
wire P3_U3877 , P3_U3878 , P3_U3879 , P3_U3880 , P3_U3881 , P3_U3882 , P3_U3883 , P3_U3884 , P3_U3885 , P3_U3886;
wire P3_U3887 , P3_U3888 , P3_U3889 , P3_U3890 , P3_U3891 , P3_U3892 , P3_U3893 , P3_U3894 , P3_U3895 , P3_U3896;
wire P3_U3897 , P3_U3898 , P3_U3899 , P3_U3900 , P3_U3901 , P3_U3902 , P3_U3903 , P3_U3904 , P3_U3905 , P3_U3906;
wire P3_U3907 , P3_U3908 , P3_U3909 , P3_U3910 , P3_U3911 , P3_U3912 , P3_U3913 , P3_U3914 , P3_U3915 , P3_U3916;
wire P3_U3917 , P3_U3918 , P3_U3919 , P3_U3920 , P3_U3921 , P3_U3922 , P3_U3923 , P3_U3924 , P3_U3925 , P3_U3926;
wire P3_U3927 , P3_U3928 , P3_U3929 , P3_U3930 , P3_U3931 , P3_U3932 , P3_U3933 , P3_U3934 , P3_U3935 , P3_U3936;
wire P3_U3937 , P3_U3938 , P3_U3939 , P3_U3940 , P3_U3941 , P3_U3942 , P3_U3943 , P3_U3944 , P3_U3945 , P3_U3946;
wire P3_U3947 , P3_U3948 , P3_U3949 , P3_U3950 , P3_U3951 , P3_U3952 , P3_U3953 , P3_U3954 , P3_U3955 , P3_U3956;
wire P3_U3957 , P3_U3958 , P3_U3959 , P3_U3960 , P3_U3961 , P3_U3962 , P3_U3963 , P3_U3964 , P3_U3965 , P3_U3966;
wire P3_U3967 , P3_U3968 , P3_U3969 , P3_U3970 , P3_U3971 , P3_U3972 , P3_U3973 , P3_U3974 , P3_U3975 , P3_U3976;
wire P3_U3977 , P3_U3978 , P3_U3979 , P3_U3980 , P3_U3981 , P3_U3982 , P3_U3983 , P3_U3984 , P3_U3985 , P3_U3986;
wire P3_U3987 , P3_U3988 , P3_U3989 , P3_U3990 , P3_U3991 , P3_U3992 , P3_U3993 , P3_U3994 , P3_U3995 , P3_U3996;
wire P3_U3997 , P3_U3998 , P3_U3999 , P3_U4000 , P3_U4001 , P3_U4002 , P3_U4003 , P3_U4004 , P3_U4005 , P3_U4006;
wire P3_U4007 , P3_U4008 , P3_U4009 , P3_U4010 , P3_U4011 , P3_U4012 , P3_U4013 , P3_U4014 , P3_U4015 , P3_U4016;
wire P3_U4017 , P3_U4018 , P3_U4019 , P3_U4020 , P3_U4021 , P3_U4022 , P3_U4023 , P3_U4024 , P3_U4025 , P3_U4026;
wire P3_U4027 , P3_U4028 , P3_U4029 , P3_U4030 , P3_U4031 , P3_U4032 , P3_U4033 , P3_U4034 , P3_U4035 , P3_U4036;
wire P3_U4037 , P3_U4038 , P3_U4039 , P3_U4040 , P3_U4041 , P3_U4042 , P3_U4043 , P3_U4044 , P3_U4045 , P3_U4046;
wire P3_U4047 , P3_U4048 , P3_U4049 , P3_U4050 , P3_U4051 , P3_U4052 , P3_U4053 , P3_U4054 , P3_U4055 , P3_U4056;
wire P3_U4057 , P3_U4058 , P3_U4059 , P3_U4060 , P3_U4061 , P3_U4062 , P3_U4063 , P3_U4064 , P3_U4065 , P3_U4066;
wire P3_U4067 , P3_U4068 , P3_U4069 , P3_U4070 , P3_U4071 , P3_U4072 , P3_U4073 , P3_U4074 , P3_U4075 , P3_U4076;
wire P3_U4077 , P3_U4078 , P3_U4079 , P3_U4080 , P3_U4081 , P3_U4082 , P3_U4083 , P3_U4084 , P3_U4085 , P3_U4086;
wire P3_U4087 , P3_U4088 , P3_U4089 , P3_U4090 , P3_U4091 , P3_U4092 , P3_U4093 , P3_U4094 , P3_U4095 , P3_U4096;
wire P3_U4097 , P3_U4098 , P3_U4099 , P3_U4100 , P3_U4101 , P3_U4102 , P3_U4103 , P3_U4104 , P3_U4105 , P3_U4106;
wire P3_U4107 , P3_U4108 , P3_U4109 , P3_U4110 , P3_U4111 , P3_U4112 , P3_U4113 , P3_U4114 , P3_U4115 , P3_U4116;
wire P3_U4117 , P3_U4118 , P3_U4119 , P3_U4120 , P3_U4121 , P3_U4122 , P3_U4123 , P3_U4124 , P3_U4125 , P3_U4126;
wire P3_U4127 , P3_U4128 , P3_U4129 , P3_U4130 , P3_U4131 , P3_U4132 , P3_U4133 , P3_U4134 , P3_U4135 , P3_U4136;
wire P3_U4137 , P3_U4138 , P3_U4139 , P3_U4140 , P3_U4141 , P3_U4142 , P3_U4143 , P3_U4144 , P3_U4145 , P3_U4146;
wire P3_U4147 , P3_U4148 , P3_U4149 , P3_U4150 , P3_U4151 , P3_U4152 , P3_U4153 , P3_U4154 , P3_U4155 , P3_U4156;
wire P3_U4157 , P3_U4158 , P3_U4159 , P3_U4160 , P3_U4161 , P3_U4162 , P3_U4163 , P3_U4164 , P3_U4165 , P3_U4166;
wire P3_U4167 , P3_U4168 , P3_U4169 , P3_U4170 , P3_U4171 , P3_U4172 , P3_U4173 , P3_U4174 , P3_U4175 , P3_U4176;
wire P3_U4177 , P3_U4178 , P3_U4179 , P3_U4180 , P3_U4181 , P3_U4182 , P3_U4183 , P3_U4184 , P3_U4185 , P3_U4186;
wire P3_U4187 , P3_U4188 , P3_U4189 , P3_U4190 , P3_U4191 , P3_U4192 , P3_U4193 , P3_U4194 , P3_U4195 , P3_U4196;
wire P3_U4197 , P3_U4198 , P3_U4199 , P3_U4200 , P3_U4201 , P3_U4202 , P3_U4203 , P3_U4204 , P3_U4205 , P3_U4206;
wire P3_U4207 , P3_U4208 , P3_U4209 , P3_U4210 , P3_U4211 , P3_U4212 , P3_U4213 , P3_U4214 , P3_U4215 , P3_U4216;
wire P3_U4217 , P3_U4218 , P3_U4219 , P3_U4220 , P3_U4221 , P3_U4222 , P3_U4223 , P3_U4224 , P3_U4225 , P3_U4226;
wire P3_U4227 , P3_U4228 , P3_U4229 , P3_U4230 , P3_U4231 , P3_U4232 , P3_U4233 , P3_U4234 , P3_U4235 , P3_U4236;
wire P3_U4237 , P3_U4238 , P3_U4239 , P3_U4240 , P3_U4241 , P3_U4242 , P3_U4243 , P3_U4244 , P3_U4245 , P3_U4246;
wire P3_U4247 , P3_U4248 , P3_U4249 , P3_U4250 , P3_U4251 , P3_U4252 , P3_U4253 , P3_U4254 , P3_U4255 , P3_U4256;
wire P3_U4257 , P3_U4258 , P3_U4259 , P3_U4260 , P3_U4261 , P3_U4262 , P3_U4263 , P3_U4264 , P3_U4265 , P3_U4266;
wire P3_U4267 , P3_U4268 , P3_U4269 , P3_U4270 , P3_U4271 , P3_U4272 , P3_U4273 , P3_U4274 , P3_U4275 , P3_U4276;
wire P3_U4277 , P3_U4278 , P3_U4279 , P3_U4280 , P3_U4281 , P3_U4282 , P3_U4283 , P3_U4284 , P3_U4285 , P3_U4286;
wire P3_U4287 , P3_U4288 , P3_U4289 , P3_U4290 , P3_U4291 , P3_U4292 , P3_U4293 , P3_U4294 , P3_U4295 , P3_U4296;
wire P3_U4297 , P3_U4298 , P3_U4299 , P3_U4300 , P3_U4301 , P3_U4302 , P3_U4303 , P3_U4304 , P3_U4305 , P3_U4306;
wire P3_U4307 , P3_U4308 , P3_U4309 , P3_U4310 , P3_U4311 , P3_U4312 , P3_U4313 , P3_U4314 , P3_U4315 , P3_U4316;
wire P3_U4317 , P3_U4318 , P3_U4319 , P3_U4320 , P3_U4321 , P3_U4322 , P3_U4323 , P3_U4324 , P3_U4325 , P3_U4326;
wire P3_U4327 , P3_U4328 , P3_U4329 , P3_U4330 , P3_U4331 , P3_U4332 , P3_U4333 , P3_U4334 , P3_U4335 , P3_U4336;
wire P3_U4337 , P3_U4338 , P3_U4339 , P3_U4340 , P3_U4341 , P3_U4342 , P3_U4343 , P3_U4344 , P3_U4345 , P3_U4346;
wire P3_U4347 , P3_U4348 , P3_U4349 , P3_U4350 , P3_U4351 , P3_U4352 , P3_U4353 , P3_U4354 , P3_U4355 , P3_U4356;
wire P3_U4357 , P3_U4358 , P3_U4359 , P3_U4360 , P3_U4361 , P3_U4362 , P3_U4363 , P3_U4364 , P3_U4365 , P3_U4366;
wire P3_U4367 , P3_U4368 , P3_U4369 , P3_U4370 , P3_U4371 , P3_U4372 , P3_U4373 , P3_U4374 , P3_U4375 , P3_U4376;
wire P3_U4377 , P3_U4378 , P3_U4379 , P3_U4380 , P3_U4381 , P3_U4382 , P3_U4383 , P3_U4384 , P3_U4385 , P3_U4386;
wire P3_U4387 , P3_U4388 , P3_U4389 , P3_U4390 , P3_U4391 , P3_U4392 , P3_U4393 , P3_U4394 , P3_U4395 , P3_U4396;
wire P3_U4397 , P3_U4398 , P3_U4399 , P3_U4400 , P3_U4401 , P3_U4402 , P3_U4403 , P3_U4404 , P3_U4405 , P3_U4406;
wire P3_U4407 , P3_U4408 , P3_U4409 , P3_U4410 , P3_U4411 , P3_U4412 , P3_U4413 , P3_U4414 , P3_U4415 , P3_U4416;
wire P3_U4417 , P3_U4418 , P3_U4419 , P3_U4420 , P3_U4421 , P3_U4422 , P3_U4423 , P3_U4424 , P3_U4425 , P3_U4426;
wire P3_U4427 , P3_U4428 , P3_U4429 , P3_U4430 , P3_U4431 , P3_U4432 , P3_U4433 , P3_U4434 , P3_U4435 , P3_U4436;
wire P3_U4437 , P3_U4438 , P3_U4439 , P3_U4440 , P3_U4441 , P3_U4442 , P3_U4443 , P3_U4444 , P3_U4445 , P3_U4446;
wire P3_U4447 , P3_U4448 , P3_U4449 , P3_U4450 , P3_U4451 , P3_U4452 , P3_U4453 , P3_U4454 , P3_U4455 , P3_U4456;
wire P3_U4457 , P3_U4458 , P3_U4459 , P3_U4460 , P3_U4461 , P3_U4462 , P3_U4463 , P3_U4464 , P3_U4465 , P3_U4466;
wire P3_U4467 , P3_U4468 , P3_U4469 , P3_U4470 , P3_U4471 , P3_U4472 , P3_U4473 , P3_U4474 , P3_U4475 , P3_U4476;
wire P3_U4477 , P3_U4478 , P3_U4479 , P3_U4480 , P3_U4481 , P3_U4482 , P3_U4483 , P3_U4484 , P3_U4485 , P3_U4486;
wire P3_U4487 , P3_U4488 , P3_U4489 , P3_U4490 , P3_U4491 , P3_U4492 , P3_U4493 , P3_U4494 , P3_U4495 , P3_U4496;
wire P3_U4497 , P3_U4498 , P3_U4499 , P3_U4500 , P3_U4501 , P3_U4502 , P3_U4503 , P3_U4504 , P3_U4505 , P3_U4506;
wire P3_U4507 , P3_U4508 , P3_U4509 , P3_U4510 , P3_U4511 , P3_U4512 , P3_U4513 , P3_U4514 , P3_U4515 , P3_U4516;
wire P3_U4517 , P3_U4518 , P3_U4519 , P3_U4520 , P3_U4521 , P3_U4522 , P3_U4523 , P3_U4524 , P3_U4525 , P3_U4526;
wire P3_U4527 , P3_U4528 , P3_U4529 , P3_U4530 , P3_U4531 , P3_U4532 , P3_U4533 , P3_U4534 , P3_U4535 , P3_U4536;
wire P3_U4537 , P3_U4538 , P3_U4539 , P3_U4540 , P3_U4541 , P3_U4542 , P3_U4543 , P3_U4544 , P3_U4545 , P3_U4546;
wire P3_U4547 , P3_U4548 , P3_U4549 , P3_U4550 , P3_U4551 , P3_U4552 , P3_U4553 , P3_U4554 , P3_U4555 , P3_U4556;
wire P3_U4557 , P3_U4558 , P3_U4559 , P3_U4560 , P3_U4561 , P3_U4562 , P3_U4563 , P3_U4564 , P3_U4565 , P3_U4566;
wire P3_U4567 , P3_U4568 , P3_U4569 , P3_U4570 , P3_U4571 , P3_U4572 , P3_U4573 , P3_U4574 , P3_U4575 , P3_U4576;
wire P3_U4577 , P3_U4578 , P3_U4579 , P3_U4580 , P3_U4581 , P3_U4582 , P3_U4583 , P3_U4584 , P3_U4585 , P3_U4586;
wire P3_U4587 , P3_U4588 , P3_U4589 , P3_U4590 , P3_U4591 , P3_U4592 , P3_U4593 , P3_U4594 , P3_U4595 , P3_U4596;
wire P3_U4597 , P3_U4598 , P3_U4599 , P3_U4600 , P3_U4601 , P3_U4602 , P3_U4603 , P3_U4604 , P3_U4605 , P3_U4606;
wire P3_U4607 , P3_U4608 , P3_U4609 , P3_U4610 , P3_U4611 , P3_U4612 , P3_U4613 , P3_U4614 , P3_U4615 , P3_U4616;
wire P3_U4617 , P3_U4618 , P3_U4619 , P3_U4620 , P3_U4621 , P3_U4622 , P3_U4623 , P3_U4624 , P3_U4625 , P3_U4626;
wire P3_U4627 , P3_U4628 , P3_U4629 , P3_U4630 , P3_U4631 , P3_U4632 , P3_U4633 , P3_U4634 , P3_U4635 , P3_U4636;
wire P3_U4637 , P3_U4638 , P3_U4639 , P3_U4640 , P3_U4641 , P3_U4642 , P3_U4643 , P3_U4644 , P3_U4645 , P3_U4646;
wire P3_U4647 , P3_U4648 , P3_U4649 , P3_U4650 , P3_U4651 , P3_U4652 , P3_U4653 , P3_U4654 , P3_U4655 , P3_U4656;
wire P3_U4657 , P3_U4658 , P3_U4659 , P3_U4660 , P3_U4661 , P3_U4662 , P3_U4663 , P3_U4664 , P3_U4665 , P3_U4666;
wire P3_U4667 , P3_U4668 , P3_U4669 , P3_U4670 , P3_U4671 , P3_U4672 , P3_U4673 , P3_U4674 , P3_U4675 , P3_U4676;
wire P3_U4677 , P3_U4678 , P3_U4679 , P3_U4680 , P3_U4681 , P3_U4682 , P3_U4683 , P3_U4684 , P3_U4685 , P3_U4686;
wire P3_U4687 , P3_U4688 , P3_U4689 , P3_U4690 , P3_U4691 , P3_U4692 , P3_U4693 , P3_U4694 , P3_U4695 , P3_U4696;
wire P3_U4697 , P3_U4698 , P3_U4699 , P3_U4700 , P3_U4701 , P3_U4702 , P3_U4703 , P3_U4704 , P3_U4705 , P3_U4706;
wire P3_U4707 , P3_U4708 , P3_U4709 , P3_U4710 , P3_U4711 , P3_U4712 , P3_U4713 , P3_U4714 , P3_U4715 , P3_U4716;
wire P3_U4717 , P3_U4718 , P3_U4719 , P3_U4720 , P3_U4721 , P3_U4722 , P3_U4723 , P3_U4724 , P3_U4725 , P3_U4726;
wire P3_U4727 , P3_U4728 , P3_U4729 , P3_U4730 , P3_U4731 , P3_U4732 , P3_U4733 , P3_U4734 , P3_U4735 , P3_U4736;
wire P3_U4737 , P3_U4738 , P3_U4739 , P3_U4740 , P3_U4741 , P3_U4742 , P3_U4743 , P3_U4744 , P3_U4745 , P3_U4746;
wire P3_U4747 , P3_U4748 , P3_U4749 , P3_U4750 , P3_U4751 , P3_U4752 , P3_U4753 , P3_U4754 , P3_U4755 , P3_U4756;
wire P3_U4757 , P3_U4758 , P3_U4759 , P3_U4760 , P3_U4761 , P3_U4762 , P3_U4763 , P3_U4764 , P3_U4765 , P3_U4766;
wire P3_U4767 , P3_U4768 , P3_U4769 , P3_U4770 , P3_U4771 , P3_U4772 , P3_U4773 , P3_U4774 , P3_U4775 , P3_U4776;
wire P3_U4777 , P3_U4778 , P3_U4779 , P3_U4780 , P3_U4781 , P3_U4782 , P3_U4783 , P3_U4784 , P3_U4785 , P3_U4786;
wire P3_U4787 , P3_U4788 , P3_U4789 , P3_U4790 , P3_U4791 , P3_U4792 , P3_U4793 , P3_U4794 , P3_U4795 , P3_U4796;
wire P3_U4797 , P3_U4798 , P3_U4799 , P3_U4800 , P3_U4801 , P3_U4802 , P3_U4803 , P3_U4804 , P3_U4805 , P3_U4806;
wire P3_U4807 , P3_U4808 , P3_U4809 , P3_U4810 , P3_U4811 , P3_U4812 , P3_U4813 , P3_U4814 , P3_U4815 , P3_U4816;
wire P3_U4817 , P3_U4818 , P3_U4819 , P3_U4820 , P3_U4821 , P3_U4822 , P3_U4823 , P3_U4824 , P3_U4825 , P3_U4826;
wire P3_U4827 , P3_U4828 , P3_U4829 , P3_U4830 , P3_U4831 , P3_U4832 , P3_U4833 , P3_U4834 , P3_U4835 , P3_U4836;
wire P3_U4837 , P3_U4838 , P3_U4839 , P3_U4840 , P3_U4841 , P3_U4842 , P3_U4843 , P3_U4844 , P3_U4845 , P3_U4846;
wire P3_U4847 , P3_U4848 , P3_U4849 , P3_U4850 , P3_U4851 , P3_U4852 , P3_U4853 , P3_U4854 , P3_U4855 , P3_U4856;
wire P3_U4857 , P3_U4858 , P3_U4859 , P3_U4860 , P3_U4861 , P3_U4862 , P3_U4863 , P3_U4864 , P3_U4865 , P3_U4866;
wire P3_U4867 , P3_U4868 , P3_U4869 , P3_U4870 , P3_U4871 , P3_U4872 , P3_U4873 , P3_U4874 , P3_U4875 , P3_U4876;
wire P3_U4877 , P3_U4878 , P3_U4879 , P3_U4880 , P3_U4881 , P3_U4882 , P3_U4883 , P3_U4884 , P3_U4885 , P3_U4886;
wire P3_U4887 , P3_U4888 , P3_U4889 , P3_U4890 , P3_U4891 , P3_U4892 , P3_U4893 , P3_U4894 , P3_U4895 , P3_U4896;
wire P3_U4897 , P3_U4898 , P3_U4899 , P3_U4900 , P3_U4901 , P3_U4902 , P3_U4903 , P3_U4904 , P3_U4905 , P3_U4906;
wire P3_U4907 , P3_U4908 , P3_U4909 , P3_U4910 , P3_U4911 , P3_U4912 , P3_U4913 , P3_U4914 , P3_U4915 , P3_U4916;
wire P3_U4917 , P3_U4918 , P3_U4919 , P3_U4920 , P3_U4921 , P3_U4922 , P3_U4923 , P3_U4924 , P3_U4925 , P3_U4926;
wire P3_U4927 , P3_U4928 , P3_U4929 , P3_U4930 , P3_U4931 , P3_U4932 , P3_U4933 , P3_U4934 , P3_U4935 , P3_U4936;
wire P3_U4937 , P3_U4938 , P3_U4939 , P3_U4940 , P3_U4941 , P3_U4942 , P3_U4943 , P3_U4944 , P3_U4945 , P3_U4946;
wire P3_U4947 , P3_U4948 , P3_U4949 , P3_U4950 , P3_U4951 , P3_U4952 , P3_U4953 , P3_U4954 , P3_U4955 , P3_U4956;
wire P3_U4957 , P3_U4958 , P3_U4959 , P3_U4960 , P3_U4961 , P3_U4962 , P3_U4963 , P3_U4964 , P3_U4965 , P3_U4966;
wire P3_U4967 , P3_U4968 , P3_U4969 , P3_U4970 , P3_U4971 , P3_U4972 , P3_U4973 , P3_U4974 , P3_U4975 , P3_U4976;
wire P3_U4977 , P3_U4978 , P3_U4979 , P3_U4980 , P3_U4981 , P3_U4982 , P3_U4983 , P3_U4984 , P3_U4985 , P3_U4986;
wire P3_U4987 , P3_U4988 , P3_U4989 , P3_U4990 , P3_U4991 , P3_U4992 , P3_U4993 , P3_U4994 , P3_U4995 , P3_U4996;
wire P3_U4997 , P3_U4998 , P3_U4999 , P3_U5000 , P3_U5001 , P3_U5002 , P3_U5003 , P3_U5004 , P3_U5005 , P3_U5006;
wire P3_U5007 , P3_U5008 , P3_U5009 , P3_U5010 , P3_U5011 , P3_U5012 , P3_U5013 , P3_U5014 , P3_U5015 , P3_U5016;
wire P3_U5017 , P3_U5018 , P3_U5019 , P3_U5020 , P3_U5021 , P3_U5022 , P3_U5023 , P3_U5024 , P3_U5025 , P3_U5026;
wire P3_U5027 , P3_U5028 , P3_U5029 , P3_U5030 , P3_U5031 , P3_U5032 , P3_U5033 , P3_U5034 , P3_U5035 , P3_U5036;
wire P3_U5037 , P3_U5038 , P3_U5039 , P3_U5040 , P3_U5041 , P3_U5042 , P3_U5043 , P3_U5044 , P3_U5045 , P3_U5046;
wire P3_U5047 , P3_U5048 , P3_U5049 , P3_U5050 , P3_U5051 , P3_U5052 , P3_U5053 , P3_U5054 , P3_U5055 , P3_U5056;
wire P3_U5057 , P3_U5058 , P3_U5059 , P3_U5060 , P3_U5061 , P3_U5062 , P3_U5063 , P3_U5064 , P3_U5065 , P3_U5066;
wire P3_U5067 , P3_U5068 , P3_U5069 , P3_U5070 , P3_U5071 , P3_U5072 , P3_U5073 , P3_U5074 , P3_U5075 , P3_U5076;
wire P3_U5077 , P3_U5078 , P3_U5079 , P3_U5080 , P3_U5081 , P3_U5082 , P3_U5083 , P3_U5084 , P3_U5085 , P3_U5086;
wire P3_U5087 , P3_U5088 , P3_U5089 , P3_U5090 , P3_U5091 , P3_U5092 , P3_U5093 , P3_U5094 , P3_U5095 , P3_U5096;
wire P3_U5097 , P3_U5098 , P3_U5099 , P3_U5100 , P3_U5101 , P3_U5102 , P3_U5103 , P3_U5104 , P3_U5105 , P3_U5106;
wire P3_U5107 , P3_U5108 , P3_U5109 , P3_U5110 , P3_U5111 , P3_U5112 , P3_U5113 , P3_U5114 , P3_U5115 , P3_U5116;
wire P3_U5117 , P3_U5118 , P3_U5119 , P3_U5120 , P3_U5121 , P3_U5122 , P3_U5123 , P3_U5124 , P3_U5125 , P3_U5126;
wire P3_U5127 , P3_U5128 , P3_U5129 , P3_U5130 , P3_U5131 , P3_U5132 , P3_U5133 , P3_U5134 , P3_U5135 , P3_U5136;
wire P3_U5137 , P3_U5138 , P3_U5139 , P3_U5140 , P3_U5141 , P3_U5142 , P3_U5143 , P3_U5144 , P3_U5145 , P3_U5146;
wire P3_U5147 , P3_U5148 , P3_U5149 , P3_U5150 , P3_U5151 , P3_U5152 , P3_U5153 , P3_U5154 , P3_U5155 , P3_U5156;
wire P3_U5157 , P3_U5158 , P3_U5159 , P3_U5160 , P3_U5161 , P3_U5162 , P3_U5163 , P3_U5164 , P3_U5165 , P3_U5166;
wire P3_U5167 , P3_U5168 , P3_U5169 , P3_U5170 , P3_U5171 , P3_U5172 , P3_U5173 , P3_U5174 , P3_U5175 , P3_U5176;
wire P3_U5177 , P3_U5178 , P3_U5179 , P3_U5180 , P3_U5181 , P3_U5182 , P3_U5183 , P3_U5184 , P3_U5185 , P3_U5186;
wire P3_U5187 , P3_U5188 , P3_U5189 , P3_U5190 , P3_U5191 , P3_U5192 , P3_U5193 , P3_U5194 , P3_U5195 , P3_U5196;
wire P3_U5197 , P3_U5198 , P3_U5199 , P3_U5200 , P3_U5201 , P3_U5202 , P3_U5203 , P3_U5204 , P3_U5205 , P3_U5206;
wire P3_U5207 , P3_U5208 , P3_U5209 , P3_U5210 , P3_U5211 , P3_U5212 , P3_U5213 , P3_U5214 , P3_U5215 , P3_U5216;
wire P3_U5217 , P3_U5218 , P3_U5219 , P3_U5220 , P3_U5221 , P3_U5222 , P3_U5223 , P3_U5224 , P3_U5225 , P3_U5226;
wire P3_U5227 , P3_U5228 , P3_U5229 , P3_U5230 , P3_U5231 , P3_U5232 , P3_U5233 , P3_U5234 , P3_U5235 , P3_U5236;
wire P3_U5237 , P3_U5238 , P3_U5239 , P3_U5240 , P3_U5241 , P3_U5242 , P3_U5243 , P3_U5244 , P3_U5245 , P3_U5246;
wire P3_U5247 , P3_U5248 , P3_U5249 , P3_U5250 , P3_U5251 , P3_U5252 , P3_U5253 , P3_U5254 , P3_U5255 , P3_U5256;
wire P3_U5257 , P3_U5258 , P3_U5259 , P3_U5260 , P3_U5261 , P3_U5262 , P3_U5263 , P3_U5264 , P3_U5265 , P3_U5266;
wire P3_U5267 , P3_U5268 , P3_U5269 , P3_U5270 , P3_U5271 , P3_U5272 , P3_U5273 , P3_U5274 , P3_U5275 , P3_U5276;
wire P3_U5277 , P3_U5278 , P3_U5279 , P3_U5280 , P3_U5281 , P3_U5282 , P3_U5283 , P3_U5284 , P3_U5285 , P3_U5286;
wire P3_U5287 , P3_U5288 , P3_U5289 , P3_U5290 , P3_U5291 , P3_U5292 , P3_U5293 , P3_U5294 , P3_U5295 , P3_U5296;
wire P3_U5297 , P3_U5298 , P3_U5299 , P3_U5300 , P3_U5301 , P3_U5302 , P3_U5303 , P3_U5304 , P3_U5305 , P3_U5306;
wire P3_U5307 , P3_U5308 , P3_U5309 , P3_U5310 , P3_U5311 , P3_U5312 , P3_U5313 , P3_U5314 , P3_U5315 , P3_U5316;
wire P3_U5317 , P3_U5318 , P3_U5319 , P3_U5320 , P3_U5321 , P3_U5322 , P3_U5323 , P3_U5324 , P3_U5325 , P3_U5326;
wire P3_U5327 , P3_U5328 , P3_U5329 , P3_U5330 , P3_U5331 , P3_U5332 , P3_U5333 , P3_U5334 , P3_U5335 , P3_U5336;
wire P3_U5337 , P3_U5338 , P3_U5339 , P3_U5340 , P3_U5341 , P3_U5342 , P3_U5343 , P3_U5344 , P3_U5345 , P3_U5346;
wire P3_U5347 , P3_U5348 , P3_U5349 , P3_U5350 , P3_U5351 , P3_U5352 , P3_U5353 , P3_U5354 , P3_U5355 , P3_U5356;
wire P3_U5357 , P3_U5358 , P3_U5359 , P3_U5360 , P3_U5361 , P3_U5362 , P3_U5363 , P3_U5364 , P3_U5365 , P3_U5366;
wire P3_U5367 , P3_U5368 , P3_U5369 , P3_U5370 , P3_U5371 , P3_U5372 , P3_U5373 , P3_U5374 , P3_U5375 , P3_U5376;
wire P3_U5377 , P3_U5378 , P3_U5379 , P3_U5380 , P3_U5381 , P3_U5382 , P3_U5383 , P3_U5384 , P3_U5385 , P3_U5386;
wire P3_U5387 , P3_U5388 , P3_U5389 , P3_U5390 , P3_U5391 , P3_U5392 , P3_U5393 , P3_U5394 , P3_U5395 , P3_U5396;
wire P3_U5397 , P3_U5398 , P3_U5399 , P3_U5400 , P3_U5401 , P3_U5402 , P3_U5403 , P3_U5404 , P3_U5405 , P3_U5406;
wire P3_U5407 , P3_U5408 , P3_U5409 , P3_U5410 , P3_U5411 , P3_U5412 , P3_U5413 , P3_U5414 , P3_U5415 , P3_U5416;
wire P3_U5417 , P3_U5418 , P3_U5419 , P3_U5420 , P3_U5421 , P3_U5422 , P3_U5423 , P3_U5424 , P3_U5425 , P3_U5426;
wire P3_U5427 , P3_U5428 , P3_U5429 , P3_U5430 , P3_U5431 , P3_U5432 , P3_U5433 , P3_U5434 , P3_U5435 , P3_U5436;
wire P3_U5437 , P3_U5438 , P3_U5439 , P3_U5440 , P3_U5441 , P3_U5442 , P3_U5443 , P3_U5444 , P3_U5445 , P3_U5446;
wire P3_U5447 , P3_U5448 , P3_U5449 , P3_U5450 , P3_U5451 , P3_U5452 , P3_U5453 , P3_U5454 , P3_U5455 , P3_U5456;
wire P3_U5457 , P3_U5458 , P3_U5459 , P3_U5460 , P3_U5461 , P3_U5462 , P3_U5463 , P3_U5464 , P3_U5465 , P3_U5466;
wire P3_U5467 , P3_U5468 , P3_U5469 , P3_U5470 , P3_U5471 , P3_U5472 , P3_U5473 , P3_U5474 , P3_U5475 , P3_U5476;
wire P3_U5477 , P3_U5478 , P3_U5479 , P3_U5480 , P3_U5481 , P3_U5482 , P3_U5483 , P3_U5484 , P3_U5485 , P3_U5486;
wire P3_U5487 , P3_U5488 , P3_U5489 , P3_U5490 , P3_U5491 , P3_U5492 , P3_U5493 , P3_U5494 , P3_U5495 , P3_U5496;
wire P3_U5497 , P3_U5498 , P3_U5499 , P3_U5500 , P3_U5501 , P3_U5502 , P3_U5503 , P3_U5504 , P3_U5505 , P3_U5506;
wire P3_U5507 , P3_U5508 , P3_U5509 , P3_U5510 , P3_U5511 , P3_U5512 , P3_U5513 , P3_U5514 , P3_U5515 , P3_U5516;
wire P3_U5517 , P3_U5518 , P3_U5519 , P3_U5520 , P3_U5521 , P3_U5522 , P3_U5523 , P3_U5524 , P3_U5525 , P3_U5526;
wire P3_U5527 , P3_U5528 , P3_U5529 , P3_U5530 , P3_U5531 , P3_U5532 , P3_U5533 , P3_U5534 , P3_U5535 , P3_U5536;
wire P3_U5537 , P3_U5538 , P3_U5539 , P3_U5540 , P3_U5541 , P3_U5542 , P3_U5543 , P3_U5544 , P3_U5545 , P3_U5546;
wire P3_U5547 , P3_U5548 , P3_U5549 , P3_U5550 , P3_U5551 , P3_U5552 , P3_U5553 , P3_U5554 , P3_U5555 , P3_U5556;
wire P3_U5557 , P3_U5558 , P3_U5559 , P3_U5560 , P3_U5561 , P3_U5562 , P3_U5563 , P3_U5564 , P3_U5565 , P3_U5566;
wire P3_U5567 , P3_U5568 , P3_U5569 , P3_U5570 , P3_U5571 , P3_U5572 , P3_U5573 , P3_U5574 , P3_U5575 , P3_U5576;
wire P3_U5577 , P3_U5578 , P3_U5579 , P3_U5580 , P3_U5581 , P3_U5582 , P3_U5583 , P3_U5584 , P3_U5585 , P3_U5586;
wire P3_U5587 , P3_U5588 , P3_U5589 , P3_U5590 , P3_U5591 , P3_U5592 , P3_U5593 , P3_U5594 , P3_U5595 , P3_U5596;
wire P3_U5597 , P3_U5598 , P3_U5599 , P3_U5600 , P3_U5601 , P3_U5602 , P3_U5603 , P3_U5604 , P3_U5605 , P3_U5606;
wire P3_U5607 , P3_U5608 , P3_U5609 , P3_U5610 , P3_U5611 , P3_U5612 , P3_U5613 , P3_U5614 , P3_U5615 , P3_U5616;
wire P3_U5617 , P3_U5618 , P3_U5619 , P3_U5620 , P3_U5621 , P3_U5622 , P3_U5623 , P3_U5624 , P3_U5625 , P3_U5626;
wire P3_U5627 , P3_U5628 , P3_U5629 , P3_U5630 , P3_U5631 , P3_U5632 , P3_U5633 , P3_U5634 , P3_U5635 , P3_U5636;
wire P3_U5637 , P3_U5638 , P3_U5639 , P3_U5640 , P3_U5641 , P3_U5642 , P3_U5643 , P3_U5644 , P3_U5645 , P3_U5646;
wire P3_U5647 , P3_U5648 , P3_U5649 , P3_U5650 , P3_U5651 , P3_U5652 , P3_U5653 , P3_U5654 , P3_U5655 , P3_U5656;
wire P3_U5657 , P3_U5658 , P3_U5659 , P3_U5660 , P3_U5661 , P3_U5662 , P3_U5663 , P3_U5664 , P3_U5665 , P3_U5666;
wire P3_U5667 , P3_U5668 , P3_U5669 , P3_U5670 , P3_U5671 , P3_U5672 , P3_U5673 , P3_U5674 , P3_U5675 , P3_U5676;
wire P3_U5677 , P3_U5678 , P3_U5679 , P3_U5680 , P3_U5681 , P3_U5682 , P3_U5683 , P3_U5684 , P3_U5685 , P3_U5686;
wire P3_U5687 , P3_U5688 , P3_U5689 , P3_U5690 , P3_U5691 , P3_U5692 , P3_U5693 , P3_U5694 , P3_U5695 , P3_U5696;
wire P3_U5697 , P3_U5698 , P3_U5699 , P3_U5700 , P3_U5701 , P3_U5702 , P3_U5703 , P3_U5704 , P3_U5705 , P3_U5706;
wire P3_U5707 , P3_U5708 , P3_U5709 , P3_U5710 , P3_U5711 , P3_U5712 , P3_U5713 , P3_U5714 , P3_U5715 , P3_U5716;
wire P3_U5717 , P3_U5718 , P3_U5719 , P3_U5720 , P3_U5721 , P3_U5722 , P3_U5723 , P3_U5724 , P3_U5725 , P3_U5726;
wire P3_U5727 , P3_U5728 , P3_U5729 , P3_U5730 , P3_U5731 , P3_U5732 , P3_U5733 , P3_U5734 , P3_U5735 , P3_U5736;
wire P3_U5737 , P3_U5738 , P3_U5739 , P3_U5740 , P3_U5741 , P3_U5742 , P3_U5743 , P3_U5744 , P3_U5745 , P3_U5746;
wire P3_U5747 , P3_U5748 , P3_U5749 , P3_U5750 , P3_U5751 , P3_U5752 , P3_U5753 , P3_U5754 , P3_U5755 , P3_U5756;
wire P3_U5757 , P3_U5758 , P3_U5759 , P3_U5760 , P3_U5761 , P3_U5762 , P3_U5763 , P3_U5764 , P3_U5765 , P3_U5766;
wire P3_U5767 , P3_U5768 , P3_U5769 , P3_U5770 , P3_U5771 , P3_U5772 , P3_U5773 , P3_U5774 , P3_U5775 , P3_U5776;
wire P3_U5777 , P3_U5778 , P3_U5779 , P3_U5780 , P3_U5781 , P3_U5782 , P3_U5783 , P3_U5784 , P3_U5785 , P3_U5786;
wire P3_U5787 , P3_U5788 , P3_U5789 , P3_U5790 , P3_U5791 , P3_U5792 , P3_U5793 , P3_U5794 , P3_U5795 , P3_U5796;
wire P3_U5797 , P3_U5798 , P3_U5799 , P3_U5800 , P3_U5801 , P3_U5802 , P3_U5803 , P3_U5804 , P3_U5805 , P3_U5806;
wire P3_U5807 , P3_U5808 , P3_U5809 , P3_U5810 , P3_U5811 , P3_U5812 , P3_U5813 , P3_U5814 , P3_U5815 , P3_U5816;
wire P3_U5817 , P3_U5818 , P3_U5819 , P3_U5820 , P3_U5821 , P3_U5822 , P3_U5823 , P3_U5824 , P3_U5825 , P3_U5826;
wire P3_U5827 , P3_U5828 , P3_U5829 , P3_U5830 , P3_U5831 , P3_U5832 , P3_U5833 , P3_U5834 , P3_U5835 , P3_U5836;
wire P3_U5837 , P3_U5838 , P3_U5839 , P3_U5840 , P3_U5841 , P3_U5842 , P3_U5843 , P3_U5844 , P3_U5845 , P3_U5846;
wire P3_U5847 , P3_U5848 , P3_U5849 , P3_U5850 , P3_U5851 , P3_U5852 , P3_U5853 , P3_U5854 , P3_U5855 , P3_U5856;
wire P3_U5857 , P3_U5858 , P3_U5859 , P3_U5860 , P3_U5861 , P3_U5862 , P3_U5863 , P3_U5864 , P3_U5865 , P3_U5866;
wire P3_U5867 , P3_U5868 , P3_U5869 , P3_U5870 , P3_U5871 , P3_U5872 , P3_U5873 , P3_U5874 , P3_U5875 , P3_U5876;
wire P3_U5877 , P3_U5878 , P3_U5879 , P3_U5880 , P3_U5881 , P3_U5882 , P3_U5883 , P3_U5884 , P3_U5885 , P3_U5886;
wire P3_U5887 , P3_U5888 , P3_U5889 , P3_U5890 , P3_U5891 , P3_U5892 , P3_U5893 , P3_U5894 , P3_U5895 , P3_U5896;
wire P3_U5897 , P3_U5898 , P3_U5899 , P3_U5900 , P3_U5901 , P3_U5902 , P3_U5903 , P3_U5904 , P3_U5905 , P3_U5906;
wire P3_U5907 , P3_U5908 , P3_U5909 , P3_U5910 , P3_U5911 , P3_U5912 , P3_U5913 , P3_U5914 , P3_U5915 , P3_U5916;
wire P3_U5917 , P3_U5918 , P3_U5919 , P3_U5920 , P3_U5921 , P3_U5922 , P3_U5923 , P3_U5924 , P3_U5925 , P3_U5926;
wire P3_U5927 , P3_U5928 , P3_U5929 , P3_U5930 , P3_U5931 , P3_U5932 , P3_U5933 , P3_U5934 , P3_U5935 , P3_U5936;
wire P3_U5937 , P3_U5938 , P3_U5939 , P3_U5940 , P3_U5941 , P3_U5942 , P3_U5943 , P3_U5944 , P3_U5945 , P3_U5946;
wire P3_U5947 , P3_U5948 , P3_U5949 , P3_U5950 , P3_U5951 , P3_U5952 , P3_U5953 , P3_U5954 , P3_U5955 , P3_U5956;
wire P3_U5957 , P3_U5958 , P3_U5959 , P3_U5960 , P3_U5961 , P3_U5962 , P3_U5963 , P3_U5964 , P3_U5965 , P3_U5966;
wire P3_U5967 , P3_U5968 , P3_U5969 , P3_U5970 , P3_U5971 , P3_U5972 , P3_U5973 , P3_U5974 , P3_U5975 , P3_U5976;
wire P3_U5977 , P3_U5978 , P3_U5979 , P3_U5980 , P3_U5981 , P3_U5982 , P3_U5983 , P3_U5984 , P3_U5985 , P3_U5986;
wire P3_U5987 , P3_U5988 , P3_U5989 , P3_U5990 , P3_U5991 , P3_U5992 , P3_U5993 , P3_U5994 , P3_U5995 , P3_U5996;
wire P3_U5997 , P3_U5998 , P3_U5999 , P3_U6000 , P3_U6001 , P3_U6002 , P3_U6003 , P3_U6004 , P3_U6005 , P3_U6006;
wire P3_U6007 , P3_U6008 , P3_U6009 , P3_U6010 , P3_U6011 , P3_U6012 , P3_U6013 , P3_U6014 , P3_U6015 , P3_U6016;
wire P3_U6017 , P3_U6018 , P3_U6019 , P3_U6020 , P3_U6021 , P3_U6022 , P3_U6023 , P3_U6024 , P3_U6025 , P3_U6026;
wire P3_U6027 , P3_U6028 , P3_U6029 , P3_U6030 , P3_U6031 , P3_U6032 , P3_U6033 , P3_U6034 , P3_U6035 , P3_U6036;
wire P3_U6037 , P3_U6038 , P3_U6039 , P3_U6040 , P3_U6041 , P3_U6042 , P3_U6043 , P3_U6044 , P3_U6045 , P3_U6046;
wire P3_U6047 , P3_U6048 , P3_U6049 , P3_U6050 , P3_U6051 , P3_U6052 , P3_U6053 , P3_U6054 , P3_U6055 , P3_U6056;
wire P3_U6057 , P3_U6058 , P3_U6059 , P3_U6060 , P3_U6061 , P3_U6062 , P3_U6063 , P3_U6064 , P3_U6065 , P3_U6066;
wire P3_U6067 , P3_U6068 , P3_U6069 , P3_U6070 , P3_U6071 , P3_U6072 , P3_U6073 , P3_U6074 , P3_U6075 , P3_U6076;
wire P3_U6077 , P3_U6078 , P3_U6079 , P3_U6080 , P3_U6081 , P3_U6082 , P3_U6083 , P3_U6084 , P3_U6085 , P3_U6086;
wire P3_U6087 , P3_U6088 , P3_U6089 , P3_U6090 , P3_U6091 , P3_U6092 , P3_U6093 , P3_U6094 , P3_U6095 , P3_U6096;
wire P3_U6097 , P3_U6098 , P3_U6099 , P3_U6100 , P3_U6101 , P3_U6102 , P3_U6103 , P3_U6104 , P3_U6105 , P3_U6106;
wire P3_U6107 , P3_U6108 , P3_U6109 , P3_U6110 , P3_U6111 , P3_U6112 , P3_U6113 , P3_U6114 , P3_U6115 , P3_U6116;
wire P3_U6117 , P3_U6118 , P3_U6119 , P3_U6120 , P3_U6121 , P3_U6122 , P3_U6123 , P3_U6124 , P3_U6125 , P3_U6126;
wire P3_U6127 , P3_U6128 , P3_U6129 , P3_U6130 , P3_U6131 , P3_U6132 , P3_U6133 , P3_U6134 , P3_U6135 , P3_U6136;
wire P3_U6137 , P3_U6138 , P3_U6139 , P3_U6140 , P3_U6141 , P3_U6142 , P3_U6143 , P3_U6144 , P3_U6145 , P3_U6146;
wire P3_U6147 , P3_U6148 , P3_U6149 , P3_U6150 , P3_U6151 , P3_U6152 , P3_U6153 , P3_U6154 , P3_U6155 , P3_U6156;
wire P3_U6157 , P3_U6158 , P3_U6159 , P3_U6160 , P3_U6161 , P3_U6162 , P3_U6163 , P3_U6164 , P3_U6165 , P3_U6166;
wire P3_U6167 , P3_U6168 , P3_U6169 , P3_U6170 , P3_U6171 , P3_U6172 , P3_U6173 , P3_U6174 , P3_U6175 , P3_U6176;
wire P3_U6177 , P3_U6178 , P3_U6179 , P3_U6180 , P3_U6181 , P3_U6182 , P3_U6183 , P3_U6184 , P3_U6185 , P3_U6186;
wire P3_U6187 , P3_U6188 , P3_U6189 , P3_U6190 , P3_U6191 , P3_U6192 , P3_U6193 , P3_U6194 , P3_U6195 , P3_U6196;
wire P3_U6197 , P3_U6198 , P3_U6199 , P3_U6200 , P3_U6201 , P3_U6202 , P3_U6203 , P3_U6204 , P3_U6205 , P3_U6206;
wire P3_U6207 , P3_U6208 , P3_U6209 , P3_U6210 , P3_U6211 , P3_U6212 , P3_U6213 , P3_U6214 , P3_U6215 , P3_U6216;
wire P3_U6217 , P3_U6218 , P3_U6219 , P3_U6220 , P3_U6221 , P3_U6222 , P3_U6223 , P3_U6224 , P3_U6225 , P3_U6226;
wire P3_U6227 , P3_U6228 , P3_U6229 , P3_U6230 , P3_U6231 , P3_U6232 , P3_U6233 , P3_U6234 , P3_U6235 , P3_U6236;
wire P3_U6237 , P3_U6238 , P3_U6239 , P3_U6240 , P3_U6241 , P3_U6242 , P3_U6243 , P3_U6244 , P3_U6245 , P3_U6246;
wire P3_U6247 , P3_U6248 , P3_U6249 , P3_U6250 , P3_U6251 , P3_U6252 , P3_U6253 , P3_U6254 , P3_U6255 , P3_U6256;
wire P3_U6257 , P3_U6258 , P3_U6259 , P3_U6260 , P3_U6261 , P3_U6262 , P3_U6263 , P3_U6264 , P3_U6265 , P3_U6266;
wire P3_U6267 , P3_U6268 , P3_U6269 , P3_U6270 , P3_U6271 , P3_U6272 , P3_U6273 , P3_U6274 , P3_U6275 , P3_U6276;
wire P3_U6277 , P3_U6278 , P3_U6279 , P3_U6280 , P3_U6281 , P3_U6282 , P3_U6283 , P3_U6284 , P3_U6285 , P3_U6286;
wire P3_U6287 , P3_U6288 , P3_U6289 , P3_U6290 , P3_U6291 , P3_U6292 , P3_U6293 , P3_U6294 , P3_U6295 , P3_U6296;
wire P3_U6297 , P3_U6298 , P3_U6299 , P3_U6300 , P3_U6301 , P3_U6302 , P3_U6303 , P3_U6304 , P3_U6305 , P3_U6306;
wire P3_U6307 , P3_U6308 , P3_U6309 , P3_U6310 , P3_U6311 , P3_U6312 , P3_U6313 , P3_U6314 , P3_U6315 , P3_U6316;
wire P3_U6317 , P3_U6318 , P3_U6319 , P3_U6320 , P3_U6321 , P3_U6322 , P3_U6323 , P3_U6324 , P3_U6325 , P3_U6326;
wire P3_U6327 , P3_U6328 , P3_U6329 , P3_U6330 , P3_U6331 , P3_U6332 , P3_U6333 , P3_U6334 , P3_U6335 , P3_U6336;
wire P3_U6337 , P3_U6338 , P3_U6339 , P3_U6340 , P3_U6341 , P3_U6342 , P3_U6343 , P3_U6344 , P3_U6345 , P3_U6346;
wire P3_U6347 , P3_U6348 , P3_U6349 , P3_U6350 , P3_U6351 , P3_U6352 , P3_U6353 , P3_U6354 , P3_U6355 , P3_U6356;
wire P3_U6357 , P3_U6358 , P3_U6359 , P3_U6360 , P3_U6361 , P3_U6362 , P3_U6363 , P3_U6364 , P3_U6365 , P3_U6366;
wire P3_U6367 , P3_U6368 , P3_U6369 , P3_U6370 , P3_U6371 , P3_U6372 , P3_U6373 , P3_U6374 , P3_U6375 , P3_U6376;
wire P3_U6377 , P3_U6378 , P3_U6379 , P3_U6380 , P3_U6381 , P3_U6382 , P3_U6383 , P3_U6384 , P3_U6385 , P3_U6386;
wire P3_U6387 , P3_U6388 , P3_U6389 , P3_U6390 , P3_U6391 , P3_U6392 , P3_U6393 , P3_U6394 , P3_U6395 , P3_U6396;
wire P3_U6397 , P3_U6398 , P3_U6399 , P3_U6400 , P3_U6401 , P3_U6402 , P3_U6403 , P3_U6404 , P3_U6405 , P3_U6406;
wire P3_U6407 , P3_U6408 , P3_U6409 , P3_U6410 , P3_U6411 , P3_U6412 , P3_U6413 , P3_U6414 , P3_U6415 , P3_U6416;
wire P3_U6417 , P3_U6418 , P3_U6419 , P3_U6420 , P3_U6421 , P3_U6422 , P3_U6423 , P3_U6424 , P3_U6425 , P3_U6426;
wire P3_U6427 , P3_U6428 , P3_U6429 , P3_U6430 , P3_U6431 , P3_U6432 , P3_U6433 , P3_U6434 , P3_U6435 , P3_U6436;
wire P3_U6437 , P3_U6438 , P3_U6439 , P3_U6440 , P3_U6441 , P3_U6442 , P3_U6443 , P3_U6444 , P3_U6445 , P3_U6446;
wire P3_U6447 , P3_U6448 , P3_U6449 , P3_U6450 , P3_U6451 , P3_U6452 , P3_U6453 , P3_U6454 , P3_U6455 , P3_U6456;
wire P3_U6457 , P3_U6458 , P3_U6459 , P3_U6460 , P3_U6461 , P3_U6462 , P3_U6463 , P3_U6464 , P3_U6465 , P3_U6466;
wire P3_U6467 , P3_U6468 , P3_U6469 , P3_U6470 , P3_U6471 , P3_U6472 , P3_U6473 , P3_U6474 , P3_U6475 , P3_U6476;
wire P3_U6477 , P3_U6478 , P3_U6479 , P3_U6480 , P3_U6481 , P3_U6482 , P3_U6483 , P3_U6484 , P3_U6485 , P3_U6486;
wire P3_U6487 , P3_U6488 , P3_U6489 , P3_U6490 , P3_U6491 , P3_U6492 , P3_U6493 , P3_U6494 , P3_U6495 , P3_U6496;
wire P3_U6497 , P3_U6498 , P3_U6499 , P3_U6500 , P3_U6501 , P3_U6502 , P3_U6503 , P3_U6504 , P3_U6505 , P3_U6506;
wire P3_U6507 , P3_U6508 , P3_U6509 , P3_U6510 , P3_U6511 , P3_U6512 , P3_U6513 , P3_U6514 , P3_U6515 , P3_U6516;
wire P3_U6517 , P3_U6518 , P3_U6519 , P3_U6520 , P3_U6521 , P3_U6522 , P3_U6523 , P3_U6524 , P3_U6525 , P3_U6526;
wire P3_U6527 , P3_U6528 , P3_U6529 , P3_U6530 , P3_U6531 , P3_U6532 , P3_U6533 , P3_U6534 , P3_U6535 , P3_U6536;
wire P3_U6537 , P3_U6538 , P3_U6539 , P3_U6540 , P3_U6541 , P3_U6542 , P3_U6543 , P3_U6544 , P3_U6545 , P3_U6546;
wire P3_U6547 , P3_U6548 , P3_U6549 , P3_U6550 , P3_U6551 , P3_U6552 , P3_U6553 , P3_U6554 , P3_U6555 , P3_U6556;
wire P3_U6557 , P3_U6558 , P3_U6559 , P3_U6560 , P3_U6561 , P3_U6562 , P3_U6563 , P3_U6564 , P3_U6565 , P3_U6566;
wire P3_U6567 , P3_U6568 , P3_U6569 , P3_U6570 , P3_U6571 , P3_U6572 , P3_U6573 , P3_U6574 , P3_U6575 , P3_U6576;
wire P3_U6577 , P3_U6578 , P3_U6579 , P3_U6580 , P3_U6581 , P3_U6582 , P3_U6583 , P3_U6584 , P3_U6585 , P3_U6586;
wire P3_U6587 , P3_U6588 , P3_U6589 , P3_U6590 , P3_U6591 , P3_U6592 , P3_U6593 , P3_U6594 , P3_U6595 , P3_U6596;
wire P3_U6597 , P3_U6598 , P3_U6599 , P3_U6600 , P3_U6601 , P3_U6602 , P3_U6603 , P3_U6604 , P3_U6605 , P3_U6606;
wire P3_U6607 , P3_U6608 , P3_U6609 , P3_U6610 , P3_U6611 , P3_U6612 , P3_U6613 , P3_U6614 , P3_U6615 , P3_U6616;
wire P3_U6617 , P3_U6618 , P3_U6619 , P3_U6620 , P3_U6621 , P3_U6622 , P3_U6623 , P3_U6624 , P3_U6625 , P3_U6626;
wire P3_U6627 , P3_U6628 , P3_U6629 , P3_U6630 , P3_U6631 , P3_U6632 , P3_U6633 , P3_U6634 , P3_U6635 , P3_U6636;
wire P3_U6637 , P3_U6638 , P3_U6639 , P3_U6640 , P3_U6641 , P3_U6642 , P3_U6643 , P3_U6644 , P3_U6645 , P3_U6646;
wire P3_U6647 , P3_U6648 , P3_U6649 , P3_U6650 , P3_U6651 , P3_U6652 , P3_U6653 , P3_U6654 , P3_U6655 , P3_U6656;
wire P3_U6657 , P3_U6658 , P3_U6659 , P3_U6660 , P3_U6661 , P3_U6662 , P3_U6663 , P3_U6664 , P3_U6665 , P3_U6666;
wire P3_U6667 , P3_U6668 , P3_U6669 , P3_U6670 , P3_U6671 , P3_U6672 , P3_U6673 , P3_U6674 , P3_U6675 , P3_U6676;
wire P3_U6677 , P3_U6678 , P3_U6679 , P3_U6680 , P3_U6681 , P3_U6682 , P3_U6683 , P3_U6684 , P3_U6685 , P3_U6686;
wire P3_U6687 , P3_U6688 , P3_U6689 , P3_U6690 , P3_U6691 , P3_U6692 , P3_U6693 , P3_U6694 , P3_U6695 , P3_U6696;
wire P3_U6697 , P3_U6698 , P3_U6699 , P3_U6700 , P3_U6701 , P3_U6702 , P3_U6703 , P3_U6704 , P3_U6705 , P3_U6706;
wire P3_U6707 , P3_U6708 , P3_U6709 , P3_U6710 , P3_U6711 , P3_U6712 , P3_U6713 , P3_U6714 , P3_U6715 , P3_U6716;
wire P3_U6717 , P3_U6718 , P3_U6719 , P3_U6720 , P3_U6721 , P3_U6722 , P3_U6723 , P3_U6724 , P3_U6725 , P3_U6726;
wire P3_U6727 , P3_U6728 , P3_U6729 , P3_U6730 , P3_U6731 , P3_U6732 , P3_U6733 , P3_U6734 , P3_U6735 , P3_U6736;
wire P3_U6737 , P3_U6738 , P3_U6739 , P3_U6740 , P3_U6741 , P3_U6742 , P3_U6743 , P3_U6744 , P3_U6745 , P3_U6746;
wire P3_U6747 , P3_U6748 , P3_U6749 , P3_U6750 , P3_U6751 , P3_U6752 , P3_U6753 , P3_U6754 , P3_U6755 , P3_U6756;
wire P3_U6757 , P3_U6758 , P3_U6759 , P3_U6760 , P3_U6761 , P3_U6762 , P3_U6763 , P3_U6764 , P3_U6765 , P3_U6766;
wire P3_U6767 , P3_U6768 , P3_U6769 , P3_U6770 , P3_U6771 , P3_U6772 , P3_U6773 , P3_U6774 , P3_U6775 , P3_U6776;
wire P3_U6777 , P3_U6778 , P3_U6779 , P3_U6780 , P3_U6781 , P3_U6782 , P3_U6783 , P3_U6784 , P3_U6785 , P3_U6786;
wire P3_U6787 , P3_U6788 , P3_U6789 , P3_U6790 , P3_U6791 , P3_U6792 , P3_U6793 , P3_U6794 , P3_U6795 , P3_U6796;
wire P3_U6797 , P3_U6798 , P3_U6799 , P3_U6800 , P3_U6801 , P3_U6802 , P3_U6803 , P3_U6804 , P3_U6805 , P3_U6806;
wire P3_U6807 , P3_U6808 , P3_U6809 , P3_U6810 , P3_U6811 , P3_U6812 , P3_U6813 , P3_U6814 , P3_U6815 , P3_U6816;
wire P3_U6817 , P3_U6818 , P3_U6819 , P3_U6820 , P3_U6821 , P3_U6822 , P3_U6823 , P3_U6824 , P3_U6825 , P3_U6826;
wire P3_U6827 , P3_U6828 , P3_U6829 , P3_U6830 , P3_U6831 , P3_U6832 , P3_U6833 , P3_U6834 , P3_U6835 , P3_U6836;
wire P3_U6837 , P3_U6838 , P3_U6839 , P3_U6840 , P3_U6841 , P3_U6842 , P3_U6843 , P3_U6844 , P3_U6845 , P3_U6846;
wire P3_U6847 , P3_U6848 , P3_U6849 , P3_U6850 , P3_U6851 , P3_U6852 , P3_U6853 , P3_U6854 , P3_U6855 , P3_U6856;
wire P3_U6857 , P3_U6858 , P3_U6859 , P3_U6860 , P3_U6861 , P3_U6862 , P3_U6863 , P3_U6864 , P3_U6865 , P3_U6866;
wire P3_U6867 , P3_U6868 , P3_U6869 , P3_U6870 , P3_U6871 , P3_U6872 , P3_U6873 , P3_U6874 , P3_U6875 , P3_U6876;
wire P3_U6877 , P3_U6878 , P3_U6879 , P3_U6880 , P3_U6881 , P3_U6882 , P3_U6883 , P3_U6884 , P3_U6885 , P3_U6886;
wire P3_U6887 , P3_U6888 , P3_U6889 , P3_U6890 , P3_U6891 , P3_U6892 , P3_U6893 , P3_U6894 , P3_U6895 , P3_U6896;
wire P3_U6897 , P3_U6898 , P3_U6899 , P3_U6900 , P3_U6901 , P3_U6902 , P3_U6903 , P3_U6904 , P3_U6905 , P3_U6906;
wire P3_U6907 , P3_U6908 , P3_U6909 , P3_U6910 , P3_U6911 , P3_U6912 , P3_U6913 , P3_U6914 , P3_U6915 , P3_U6916;
wire P3_U6917 , P3_U6918 , P3_U6919 , P3_U6920 , P3_U6921 , P3_U6922 , P3_U6923 , P3_U6924 , P3_U6925 , P3_U6926;
wire P3_U6927 , P3_U6928 , P3_U6929 , P3_U6930 , P3_U6931 , P3_U6932 , P3_U6933 , P3_U6934 , P3_U6935 , P3_U6936;
wire P3_U6937 , P3_U6938 , P3_U6939 , P3_U6940 , P3_U6941 , P3_U6942 , P3_U6943 , P3_U6944 , P3_U6945 , P3_U6946;
wire P3_U6947 , P3_U6948 , P3_U6949 , P3_U6950 , P3_U6951 , P3_U6952 , P3_U6953 , P3_U6954 , P3_U6955 , P3_U6956;
wire P3_U6957 , P3_U6958 , P3_U6959 , P3_U6960 , P3_U6961 , P3_U6962 , P3_U6963 , P3_U6964 , P3_U6965 , P3_U6966;
wire P3_U6967 , P3_U6968 , P3_U6969 , P3_U6970 , P3_U6971 , P3_U6972 , P3_U6973 , P3_U6974 , P3_U6975 , P3_U6976;
wire P3_U6977 , P3_U6978 , P3_U6979 , P3_U6980 , P3_U6981 , P3_U6982 , P3_U6983 , P3_U6984 , P3_U6985 , P3_U6986;
wire P3_U6987 , P3_U6988 , P3_U6989 , P3_U6990 , P3_U6991 , P3_U6992 , P3_U6993 , P3_U6994 , P3_U6995 , P3_U6996;
wire P3_U6997 , P3_U6998 , P3_U6999 , P3_U7000 , P3_U7001 , P3_U7002 , P3_U7003 , P3_U7004 , P3_U7005 , P3_U7006;
wire P3_U7007 , P3_U7008 , P3_U7009 , P3_U7010 , P3_U7011 , P3_U7012 , P3_U7013 , P3_U7014 , P3_U7015 , P3_U7016;
wire P3_U7017 , P3_U7018 , P3_U7019 , P3_U7020 , P3_U7021 , P3_U7022 , P3_U7023 , P3_U7024 , P3_U7025 , P3_U7026;
wire P3_U7027 , P3_U7028 , P3_U7029 , P3_U7030 , P3_U7031 , P3_U7032 , P3_U7033 , P3_U7034 , P3_U7035 , P3_U7036;
wire P3_U7037 , P3_U7038 , P3_U7039 , P3_U7040 , P3_U7041 , P3_U7042 , P3_U7043 , P3_U7044 , P3_U7045 , P3_U7046;
wire P3_U7047 , P3_U7048 , P3_U7049 , P3_U7050 , P3_U7051 , P3_U7052 , P3_U7053 , P3_U7054 , P3_U7055 , P3_U7056;
wire P3_U7057 , P3_U7058 , P3_U7059 , P3_U7060 , P3_U7061 , P3_U7062 , P3_U7063 , P3_U7064 , P3_U7065 , P3_U7066;
wire P3_U7067 , P3_U7068 , P3_U7069 , P3_U7070 , P3_U7071 , P3_U7072 , P3_U7073 , P3_U7074 , P3_U7075 , P3_U7076;
wire P3_U7077 , P3_U7078 , P3_U7079 , P3_U7080 , P3_U7081 , P3_U7082 , P3_U7083 , P3_U7084 , P3_U7085 , P3_U7086;
wire P3_U7087 , P3_U7088 , P3_U7089 , P3_U7090 , P3_U7091 , P3_U7092 , P3_U7093 , P3_U7094 , P3_U7095 , P3_U7096;
wire P3_U7097 , P3_U7098 , P3_U7099 , P3_U7100 , P3_U7101 , P3_U7102 , P3_U7103 , P3_U7104 , P3_U7105 , P3_U7106;
wire P3_U7107 , P3_U7108 , P3_U7109 , P3_U7110 , P3_U7111 , P3_U7112 , P3_U7113 , P3_U7114 , P3_U7115 , P3_U7116;
wire P3_U7117 , P3_U7118 , P3_U7119 , P3_U7120 , P3_U7121 , P3_U7122 , P3_U7123 , P3_U7124 , P3_U7125 , P3_U7126;
wire P3_U7127 , P3_U7128 , P3_U7129 , P3_U7130 , P3_U7131 , P3_U7132 , P3_U7133 , P3_U7134 , P3_U7135 , P3_U7136;
wire P3_U7137 , P3_U7138 , P3_U7139 , P3_U7140 , P3_U7141 , P3_U7142 , P3_U7143 , P3_U7144 , P3_U7145 , P3_U7146;
wire P3_U7147 , P3_U7148 , P3_U7149 , P3_U7150 , P3_U7151 , P3_U7152 , P3_U7153 , P3_U7154 , P3_U7155 , P3_U7156;
wire P3_U7157 , P3_U7158 , P3_U7159 , P3_U7160 , P3_U7161 , P3_U7162 , P3_U7163 , P3_U7164 , P3_U7165 , P3_U7166;
wire P3_U7167 , P3_U7168 , P3_U7169 , P3_U7170 , P3_U7171 , P3_U7172 , P3_U7173 , P3_U7174 , P3_U7175 , P3_U7176;
wire P3_U7177 , P3_U7178 , P3_U7179 , P3_U7180 , P3_U7181 , P3_U7182 , P3_U7183 , P3_U7184 , P3_U7185 , P3_U7186;
wire P3_U7187 , P3_U7188 , P3_U7189 , P3_U7190 , P3_U7191 , P3_U7192 , P3_U7193 , P3_U7194 , P3_U7195 , P3_U7196;
wire P3_U7197 , P3_U7198 , P3_U7199 , P3_U7200 , P3_U7201 , P3_U7202 , P3_U7203 , P3_U7204 , P3_U7205 , P3_U7206;
wire P3_U7207 , P3_U7208 , P3_U7209 , P3_U7210 , P3_U7211 , P3_U7212 , P3_U7213 , P3_U7214 , P3_U7215 , P3_U7216;
wire P3_U7217 , P3_U7218 , P3_U7219 , P3_U7220 , P3_U7221 , P3_U7222 , P3_U7223 , P3_U7224 , P3_U7225 , P3_U7226;
wire P3_U7227 , P3_U7228 , P3_U7229 , P3_U7230 , P3_U7231 , P3_U7232 , P3_U7233 , P3_U7234 , P3_U7235 , P3_U7236;
wire P3_U7237 , P3_U7238 , P3_U7239 , P3_U7240 , P3_U7241 , P3_U7242 , P3_U7243 , P3_U7244 , P3_U7245 , P3_U7246;
wire P3_U7247 , P3_U7248 , P3_U7249 , P3_U7250 , P3_U7251 , P3_U7252 , P3_U7253 , P3_U7254 , P3_U7255 , P3_U7256;
wire P3_U7257 , P3_U7258 , P3_U7259 , P3_U7260 , P3_U7261 , P3_U7262 , P3_U7263 , P3_U7264 , P3_U7265 , P3_U7266;
wire P3_U7267 , P3_U7268 , P3_U7269 , P3_U7270 , P3_U7271 , P3_U7272 , P3_U7273 , P3_U7274 , P3_U7275 , P3_U7276;
wire P3_U7277 , P3_U7278 , P3_U7279 , P3_U7280 , P3_U7281 , P3_U7282 , P3_U7283 , P3_U7284 , P3_U7285 , P3_U7286;
wire P3_U7287 , P3_U7288 , P3_U7289 , P3_U7290 , P3_U7291 , P3_U7292 , P3_U7293 , P3_U7294 , P3_U7295 , P3_U7296;
wire P3_U7297 , P3_U7298 , P3_U7299 , P3_U7300 , P3_U7301 , P3_U7302 , P3_U7303 , P3_U7304 , P3_U7305 , P3_U7306;
wire P3_U7307 , P3_U7308 , P3_U7309 , P3_U7310 , P3_U7311 , P3_U7312 , P3_U7313 , P3_U7314 , P3_U7315 , P3_U7316;
wire P3_U7317 , P3_U7318 , P3_U7319 , P3_U7320 , P3_U7321 , P3_U7322 , P3_U7323 , P3_U7324 , P3_U7325 , P3_U7326;
wire P3_U7327 , P3_U7328 , P3_U7329 , P3_U7330 , P3_U7331 , P3_U7332 , P3_U7333 , P3_U7334 , P3_U7335 , P3_U7336;
wire P3_U7337 , P3_U7338 , P3_U7339 , P3_U7340 , P3_U7341 , P3_U7342 , P3_U7343 , P3_U7344 , P3_U7345 , P3_U7346;
wire P3_U7347 , P3_U7348 , P3_U7349 , P3_U7350 , P3_U7351 , P3_U7352 , P3_U7353 , P3_U7354 , P3_U7355 , P3_U7356;
wire P3_U7357 , P3_U7358 , P3_U7359 , P3_U7360 , P3_U7361 , P3_U7362 , P3_U7363 , P3_U7364 , P3_U7365 , P3_U7366;
wire P3_U7367 , P3_U7368 , P3_U7369 , P3_U7370 , P3_U7371 , P3_U7372 , P3_U7373 , P3_U7374 , P3_U7375 , P3_U7376;
wire P3_U7377 , P3_U7378 , P3_U7379 , P3_U7380 , P3_U7381 , P3_U7382 , P3_U7383 , P3_U7384 , P3_U7385 , P3_U7386;
wire P3_U7387 , P3_U7388 , P3_U7389 , P3_U7390 , P3_U7391 , P3_U7392 , P3_U7393 , P3_U7394 , P3_U7395 , P3_U7396;
wire P3_U7397 , P3_U7398 , P3_U7399 , P3_U7400 , P3_U7401 , P3_U7402 , P3_U7403 , P3_U7404 , P3_U7405 , P3_U7406;
wire P3_U7407 , P3_U7408 , P3_U7409 , P3_U7410 , P3_U7411 , P3_U7412 , P3_U7413 , P3_U7414 , P3_U7415 , P3_U7416;
wire P3_U7417 , P3_U7418 , P3_U7419 , P3_U7420 , P3_U7421 , P3_U7422 , P3_U7423 , P3_U7424 , P3_U7425 , P3_U7426;
wire P3_U7427 , P3_U7428 , P3_U7429 , P3_U7430 , P3_U7431 , P3_U7432 , P3_U7433 , P3_U7434 , P3_U7435 , P3_U7436;
wire P3_U7437 , P3_U7438 , P3_U7439 , P3_U7440 , P3_U7441 , P3_U7442 , P3_U7443 , P3_U7444 , P3_U7445 , P3_U7446;
wire P3_U7447 , P3_U7448 , P3_U7449 , P3_U7450 , P3_U7451 , P3_U7452 , P3_U7453 , P3_U7454 , P3_U7455 , P3_U7456;
wire P3_U7457 , P3_U7458 , P3_U7459 , P3_U7460 , P3_U7461 , P3_U7462 , P3_U7463 , P3_U7464 , P3_U7465 , P3_U7466;
wire P3_U7467 , P3_U7468 , P3_U7469 , P3_U7470 , P3_U7471 , P3_U7472 , P3_U7473 , P3_U7474 , P3_U7475 , P3_U7476;
wire P3_U7477 , P3_U7478 , P3_U7479 , P3_U7480 , P3_U7481 , P3_U7482 , P3_U7483 , P3_U7484 , P3_U7485 , P3_U7486;
wire P3_U7487 , P3_U7488 , P3_U7489 , P3_U7490 , P3_U7491 , P3_U7492 , P3_U7493 , P3_U7494 , P3_U7495 , P3_U7496;
wire P3_U7497 , P3_U7498 , P3_U7499 , P3_U7500 , P3_U7501 , P3_U7502 , P3_U7503 , P3_U7504 , P3_U7505 , P3_U7506;
wire P3_U7507 , P3_U7508 , P3_U7509 , P3_U7510 , P3_U7511 , P3_U7512 , P3_U7513 , P3_U7514 , P3_U7515 , P3_U7516;
wire P3_U7517 , P3_U7518 , P3_U7519 , P3_U7520 , P3_U7521 , P3_U7522 , P3_U7523 , P3_U7524 , P3_U7525 , P3_U7526;
wire P3_U7527 , P3_U7528 , P3_U7529 , P3_U7530 , P3_U7531 , P3_U7532 , P3_U7533 , P3_U7534 , P3_U7535 , P3_U7536;
wire P3_U7537 , P3_U7538 , P3_U7539 , P3_U7540 , P3_U7541 , P3_U7542 , P3_U7543 , P3_U7544 , P3_U7545 , P3_U7546;
wire P3_U7547 , P3_U7548 , P3_U7549 , P3_U7550 , P3_U7551 , P3_U7552 , P3_U7553 , P3_U7554 , P3_U7555 , P3_U7556;
wire P3_U7557 , P3_U7558 , P3_U7559 , P3_U7560 , P3_U7561 , P3_U7562 , P3_U7563 , P3_U7564 , P3_U7565 , P3_U7566;
wire P3_U7567 , P3_U7568 , P3_U7569 , P3_U7570 , P3_U7571 , P3_U7572 , P3_U7573 , P3_U7574 , P3_U7575 , P3_U7576;
wire P3_U7577 , P3_U7578 , P3_U7579 , P3_U7580 , P3_U7581 , P3_U7582 , P3_U7583 , P3_U7584 , P3_U7585 , P3_U7586;
wire P3_U7587 , P3_U7588 , P3_U7589 , P3_U7590 , P3_U7591 , P3_U7592 , P3_U7593 , P3_U7594 , P3_U7595 , P3_U7596;
wire P3_U7597 , P3_U7598 , P3_U7599 , P3_U7600 , P3_U7601 , P3_U7602 , P3_U7603 , P3_U7604 , P3_U7605 , P3_U7606;
wire P3_U7607 , P3_U7608 , P3_U7609 , P3_U7610 , P3_U7611 , P3_U7612 , P3_U7613 , P3_U7614 , P3_U7615 , P3_U7616;
wire P3_U7617 , P3_U7618 , P3_U7619 , P3_U7620 , P3_U7621 , P3_U7622 , P3_U7623 , P3_U7624 , P3_U7625 , P3_U7626;
wire P3_U7627 , P3_U7628 , P3_U7629 , P3_U7630 , P3_U7631 , P3_U7632 , P3_U7633 , P3_U7634 , P3_U7635 , P3_U7636;
wire P3_U7637 , P3_U7638 , P3_U7639 , P3_U7640 , P3_U7641 , P3_U7642 , P3_U7643 , P3_U7644 , P3_U7645 , P3_U7646;
wire P3_U7647 , P3_U7648 , P3_U7649 , P3_U7650 , P3_U7651 , P3_U7652 , P3_U7653 , P3_U7654 , P3_U7655 , P3_U7656;
wire P3_U7657 , P3_U7658 , P3_U7659 , P3_U7660 , P3_U7661 , P3_U7662 , P3_U7663 , P3_U7664 , P3_U7665 , P3_U7666;
wire P3_U7667 , P3_U7668 , P3_U7669 , P3_U7670 , P3_U7671 , P3_U7672 , P3_U7673 , P3_U7674 , P3_U7675 , P3_U7676;
wire P3_U7677 , P3_U7678 , P3_U7679 , P3_U7680 , P3_U7681 , P3_U7682 , P3_U7683 , P3_U7684 , P3_U7685 , P3_U7686;
wire P3_U7687 , P3_U7688 , P3_U7689 , P3_U7690 , P3_U7691 , P3_U7692 , P3_U7693 , P3_U7694 , P3_U7695 , P3_U7696;
wire P3_U7697 , P3_U7698 , P3_U7699 , P3_U7700 , P3_U7701 , P3_U7702 , P3_U7703 , P3_U7704 , P3_U7705 , P3_U7706;
wire P3_U7707 , P3_U7708 , P3_U7709 , P3_U7710 , P3_U7711 , P3_U7712 , P3_U7713 , P3_U7714 , P3_U7715 , P3_U7716;
wire P3_U7717 , P3_U7718 , P3_U7719 , P3_U7720 , P3_U7721 , P3_U7722 , P3_U7723 , P3_U7724 , P3_U7725 , P3_U7726;
wire P3_U7727 , P3_U7728 , P3_U7729 , P3_U7730 , P3_U7731 , P3_U7732 , P3_U7733 , P3_U7734 , P3_U7735 , P3_U7736;
wire P3_U7737 , P3_U7738 , P3_U7739 , P3_U7740 , P3_U7741 , P3_U7742 , P3_U7743 , P3_U7744 , P3_U7745 , P3_U7746;
wire P3_U7747 , P3_U7748 , P3_U7749 , P3_U7750 , P3_U7751 , P3_U7752 , P3_U7753 , P3_U7754 , P3_U7755 , P3_U7756;
wire P3_U7757 , P3_U7758 , P3_U7759 , P3_U7760 , P3_U7761 , P3_U7762 , P3_U7763 , P3_U7764 , P3_U7765 , P3_U7766;
wire P3_U7767 , P3_U7768 , P3_U7769 , P3_U7770 , P3_U7771 , P3_U7772 , P3_U7773 , P3_U7774 , P3_U7775 , P3_U7776;
wire P3_U7777 , P3_U7778 , P3_U7779 , P3_U7780 , P3_U7781 , P3_U7782 , P3_U7783 , P3_U7784 , P3_U7785 , P3_U7786;
wire P3_U7787 , P3_U7788 , P3_U7789 , P3_U7790 , P3_U7791 , P3_U7792 , P3_U7793 , P3_U7794 , P3_U7795 , P3_U7796;
wire P3_U7797 , P3_U7798 , P3_U7799 , P3_U7800 , P3_U7801 , P3_U7802 , P3_U7803 , P3_U7804 , P3_U7805 , P3_U7806;
wire P3_U7807 , P3_U7808 , P3_U7809 , P3_U7810 , P3_U7811 , P3_U7812 , P3_U7813 , P3_U7814 , P3_U7815 , P3_U7816;
wire P3_U7817 , P3_U7818 , P3_U7819 , P3_U7820 , P3_U7821 , P3_U7822 , P3_U7823 , P3_U7824 , P3_U7825 , P3_U7826;
wire P3_U7827 , P3_U7828 , P3_U7829 , P3_U7830 , P3_U7831 , P3_U7832 , P3_U7833 , P3_U7834 , P3_U7835 , P3_U7836;
wire P3_U7837 , P3_U7838 , P3_U7839 , P3_U7840 , P3_U7841 , P3_U7842 , P3_U7843 , P3_U7844 , P3_U7845 , P3_U7846;
wire P3_U7847 , P3_U7848 , P3_U7849 , P3_U7850 , P3_U7851 , P3_U7852 , P3_U7853 , P3_U7854 , P3_U7855 , P3_U7856;
wire P3_U7857 , P3_U7858 , P3_U7859 , P3_U7860 , P3_U7861 , P3_U7862 , P3_U7863 , P3_U7864 , P3_U7865 , P3_U7866;
wire P3_U7867 , P3_U7868 , P3_U7869 , P3_U7870 , P3_U7871 , P3_U7872 , P3_U7873 , P3_U7874 , P3_U7875 , P3_U7876;
wire P3_U7877 , P3_U7878 , P3_U7879 , P3_U7880 , P3_U7881 , P3_U7882 , P3_U7883 , P3_U7884 , P3_U7885 , P3_U7886;
wire P3_U7887 , P3_U7888 , P3_U7889 , P3_U7890 , P3_U7891 , P3_U7892 , P3_U7893 , P3_U7894 , P3_U7895 , P3_U7896;
wire P3_U7897 , P3_U7898 , P3_U7899 , P3_U7900 , P3_U7901 , P3_U7902 , P3_U7903 , P3_U7904 , P3_U7905 , P3_U7906;
wire P3_U7907 , P3_U7908 , P3_U7909 , P3_U7910 , P3_U7911 , P3_U7912 , P3_U7913 , P3_U7914 , P3_U7915 , P3_U7916;
wire P3_U7917 , P3_U7918 , P3_U7919 , P3_U7920 , P3_U7921 , P3_U7922 , P3_U7923 , P3_U7924 , P3_U7925 , P3_U7926;
wire P3_U7927 , P3_U7928 , P3_U7929 , P3_U7930 , P3_U7931 , P3_U7932 , P3_U7933 , P3_U7934 , P3_U7935 , P3_U7936;
wire P3_U7937 , P3_U7938 , P3_U7939 , P3_U7940 , P3_U7941 , P3_U7942 , P3_U7943 , P3_U7944 , P3_U7945 , P3_U7946;
wire P3_U7947 , P3_U7948 , P3_U7949 , P3_U7950 , P3_U7951 , P3_U7952 , P3_U7953 , P3_U7954 , P3_U7955 , P3_U7956;
wire P3_U7957 , P3_U7958 , P3_U7959 , P3_U7960 , P3_U7961 , P3_U7962 , P3_U7963 , P3_U7964 , P3_U7965 , P3_U7966;
wire P3_U7967 , P3_U7968 , P3_U7969 , P3_U7970 , P3_U7971 , P3_U7972 , P3_U7973 , P3_U7974 , P3_U7975 , P3_U7976;
wire P3_U7977 , P3_U7978 , P3_U7979 , P3_U7980 , P3_U7981 , P3_U7982 , P3_U7983 , P3_U7984 , P3_U7985 , P3_U7986;
wire P3_U7987 , P3_U7988 , P3_U7989 , P3_U7990 , P3_U7991 , P3_U7992 , P3_U7993 , P3_U7994 , P3_U7995 , P3_U7996;
wire P3_U7997 , P3_U7998 , P3_U7999 , P3_U8000 , P3_U8001 , P3_U8002 , P3_U8003 , P3_U8004 , P3_U8005 , P3_U8006;
wire P3_U8007 , P3_U8008 , P3_U8009 , P3_U8010 , P3_U8011 , P3_U8012 , P3_U8013 , P3_U8014 , P3_U8015 , P3_U8016;
wire P3_U8017 , P3_U8018 , P3_U8019 , P3_U8020 , P3_U8021 , P3_U8022 , P3_U8023 , P3_U8024 , P3_U8025 , P3_U8026;
wire P3_U8027 , P3_U8028 , P3_U8029 , P3_U8030 , P3_U8031 , P3_U8032 , P3_U8033 , P3_U8034 , P3_U8035 , P3_U8036;
wire P3_U8037 , P3_U8038 , P3_U8039 , P3_U8040 , P3_U8041 , P3_U8042 , P3_U8043 , P3_U8044 , P3_U8045 , P3_U8046;
wire P3_U8047 , P3_U8048 , P3_U8049 , P3_U8050 , P3_U8051 , P3_U8052 , P3_U8053 , P1_ADD_515_U170 , P1_ADD_515_U169 , P1_ADD_515_U168;
wire P1_ADD_515_U167 , P1_ADD_515_U166 , P1_ADD_515_U165 , P1_ADD_515_U164 , P1_ADD_515_U163 , P1_ADD_515_U162 , P1_ADD_515_U161 , P1_ADD_515_U160 , P1_ADD_515_U159 , P1_ADD_515_U158;
wire P1_ADD_515_U157 , P1_ADD_515_U156 , P1_ADD_515_U155 , P1_ADD_515_U154 , P1_ADD_515_U153 , P1_ADD_515_U152 , P1_ADD_515_U151 , P1_ADD_515_U150 , P1_ADD_515_U149 , P1_ADD_515_U148;
wire P1_ADD_515_U147 , P1_ADD_515_U146 , P1_ADD_515_U145 , P1_ADD_515_U144 , P1_ADD_515_U143 , P1_ADD_515_U142 , P1_ADD_515_U141 , P1_ADD_515_U140 , P1_ADD_515_U139 , P1_ADD_515_U138;
wire P1_ADD_515_U137 , P1_ADD_515_U136 , P1_ADD_515_U135 , P1_ADD_515_U134 , P1_ADD_515_U133 , P1_ADD_515_U132 , P1_ADD_515_U131 , P1_ADD_515_U130 , P1_ADD_515_U129 , P1_ADD_515_U128;
wire P1_ADD_515_U127 , P1_ADD_515_U126 , P1_ADD_515_U125 , P1_ADD_515_U124 , P1_ADD_515_U123 , P1_ADD_515_U122 , P1_ADD_515_U121 , P1_ADD_515_U120 , P1_ADD_515_U119 , P1_ADD_515_U118;
wire P1_ADD_515_U117 , P1_ADD_515_U116 , P1_ADD_515_U115 , P1_ADD_515_U114 , P1_ADD_515_U113 , P1_ADD_515_U112 , P1_ADD_515_U111 , P1_ADD_515_U110 , P1_ADD_515_U109 , P1_ADD_515_U108;
wire P1_ADD_515_U107 , P1_ADD_515_U106 , P1_ADD_515_U105 , P1_ADD_515_U104 , P1_ADD_515_U103 , P1_ADD_515_U102 , P1_ADD_515_U101 , P1_ADD_515_U100 , P1_ADD_515_U99 , P1_ADD_515_U98;
wire P1_ADD_515_U97 , P1_ADD_515_U96 , P1_ADD_515_U95 , P1_ADD_515_U94 , P1_ADD_515_U93 , P1_ADD_515_U92 , P1_ADD_515_U91 , P1_ADD_515_U90 , P1_ADD_515_U89 , P1_ADD_515_U88;
wire P1_ADD_515_U87 , P1_ADD_515_U86 , P1_ADD_515_U85 , P1_ADD_515_U84 , P1_ADD_515_U83 , P1_ADD_515_U82 , P1_ADD_515_U81 , P1_ADD_515_U80 , P1_ADD_515_U79 , P1_ADD_515_U78;
wire P1_ADD_515_U77 , P1_ADD_515_U76 , P1_ADD_515_U75 , P1_ADD_515_U74 , P1_ADD_515_U73 , P1_ADD_515_U72 , P1_ADD_515_U71 , P1_ADD_515_U70 , P1_ADD_515_U69 , P1_ADD_515_U68;
wire P1_ADD_515_U67 , P1_ADD_515_U66 , P1_ADD_515_U65 , P1_ADD_515_U64 , P1_ADD_515_U63 , P1_ADD_515_U62 , P1_ADD_515_U61 , P1_ADD_515_U60 , P1_ADD_515_U59 , P1_ADD_515_U58;
wire P1_ADD_515_U57 , P1_ADD_515_U56 , P1_ADD_515_U55 , P1_ADD_515_U54 , P1_ADD_515_U53 , P1_ADD_515_U52 , P1_ADD_515_U51 , P1_ADD_515_U50 , P1_ADD_515_U49 , P1_ADD_515_U48;
wire P1_ADD_515_U47 , P1_ADD_515_U46 , P1_ADD_515_U45 , P1_ADD_515_U44 , P1_ADD_515_U43 , P1_ADD_515_U42 , P1_ADD_515_U41 , P1_ADD_515_U40 , P1_ADD_515_U39 , P1_ADD_515_U38;
wire P1_ADD_515_U37 , P1_ADD_515_U36 , P1_ADD_515_U35 , P1_ADD_515_U34 , P1_ADD_515_U33 , P1_ADD_515_U32 , P1_ADD_515_U31 , P1_ADD_515_U30 , P1_ADD_515_U29 , P1_ADD_515_U28;
wire P1_ADD_515_U27 , P1_ADD_515_U26 , P1_ADD_515_U25 , P1_ADD_515_U24 , P1_ADD_515_U23 , P1_ADD_515_U22 , P1_ADD_515_U21 , P1_ADD_515_U20 , P1_ADD_515_U19 , P1_ADD_515_U18;
wire P1_ADD_515_U17 , P1_ADD_515_U16 , P1_ADD_515_U15 , P1_ADD_515_U14 , P1_ADD_515_U13 , P1_ADD_515_U12 , P1_ADD_515_U11 , P1_ADD_515_U10 , P1_ADD_515_U9 , P1_ADD_515_U8;
wire P1_ADD_515_U7 , P1_ADD_515_U6 , P1_ADD_515_U5 , P1_ADD_515_U4 , P1_GTE_485_U7 , P1_GTE_485_U6 , P1_ADD_405_U186 , P1_ADD_405_U185 , P1_ADD_405_U184 , P1_ADD_405_U183;
wire P1_ADD_405_U182 , P1_ADD_405_U181 , P1_ADD_405_U180 , P1_ADD_405_U179 , P1_ADD_405_U178 , P1_ADD_405_U177 , P1_ADD_405_U176 , P1_ADD_405_U175 , P1_ADD_405_U174 , P1_ADD_405_U173;
wire P2_U2352 , P2_U2353 , P2_U2354 , P2_U2355 , P2_U2356 , P2_U2357 , P2_U2358 , P2_U2359 , P2_U2360 , P2_U2361;
wire P2_U2362 , P2_U2363 , P2_U2364 , P2_U2365 , P2_U2366 , P2_U2367 , P2_U2368 , P2_U2369 , P2_U2370 , P2_U2371;
wire P2_U2372 , P2_U2373 , P2_U2374 , P2_U2375 , P2_U2376 , P2_U2377 , P2_U2378 , P2_U2379 , P2_U2380 , P2_U2381;
wire P2_U2382 , P2_U2383 , P2_U2384 , P2_U2385 , P2_U2386 , P2_U2387 , P2_U2388 , P2_U2389 , P2_U2390 , P2_U2391;
wire P2_U2392 , P2_U2393 , P2_U2394 , P2_U2395 , P2_U2396 , P2_U2397 , P2_U2398 , P2_U2399 , P2_U2400 , P2_U2401;
wire P2_U2402 , P2_U2403 , P2_U2404 , P2_U2405 , P2_U2406 , P2_U2407 , P2_U2408 , P2_U2409 , P2_U2410 , P2_U2411;
wire P2_U2412 , P2_U2413 , P2_U2414 , P2_U2415 , P2_U2416 , P2_U2417 , P2_U2418 , P2_U2419 , P2_U2420 , P2_U2421;
wire P2_U2422 , P2_U2423 , P2_U2424 , P2_U2425 , P2_U2426 , P2_U2427 , P2_U2428 , P2_U2429 , P2_U2430 , P2_U2431;
wire P2_U2432 , P2_U2433 , P2_U2434 , P2_U2435 , P2_U2436 , P2_U2437 , P2_U2438 , P2_U2439 , P2_U2440 , P2_U2441;
wire P2_U2442 , P2_U2443 , P2_U2444 , P2_U2445 , P2_U2446 , P2_U2447 , P2_U2448 , P2_U2449 , P2_U2450 , P2_U2451;
wire P2_U2452 , P2_U2453 , P2_U2454 , P2_U2455 , P2_U2456 , P2_U2457 , P2_U2458 , P2_U2459 , P2_U2460 , P2_U2461;
wire P2_U2462 , P2_U2463 , P2_U2464 , P2_U2465 , P2_U2466 , P2_U2467 , P2_U2468 , P2_U2469 , P2_U2470 , P2_U2471;
wire P2_U2472 , P2_U2473 , P2_U2474 , P2_U2475 , P2_U2476 , P2_U2477 , P2_U2478 , P2_U2479 , P2_U2480 , P2_U2481;
wire P2_U2482 , P2_U2483 , P2_U2484 , P2_U2485 , P2_U2486 , P2_U2487 , P2_U2488 , P2_U2489 , P2_U2490 , P2_U2491;
wire P2_U2492 , P2_U2493 , P2_U2494 , P2_U2495 , P2_U2496 , P2_U2497 , P2_U2498 , P2_U2499 , P2_U2500 , P2_U2501;
wire P2_U2502 , P2_U2503 , P2_U2504 , P2_U2505 , P2_U2506 , P2_U2507 , P2_U2508 , P2_U2509 , P2_U2510 , P2_U2511;
wire P2_U2512 , P2_U2513 , P2_U2514 , P2_U2515 , P2_U2516 , P2_U2517 , P2_U2518 , P2_U2519 , P2_U2520 , P2_U2521;
wire P2_U2522 , P2_U2523 , P2_U2524 , P2_U2525 , P2_U2526 , P2_U2527 , P2_U2528 , P2_U2529 , P2_U2530 , P2_U2531;
wire P2_U2532 , P2_U2533 , P2_U2534 , P2_U2535 , P2_U2536 , P2_U2537 , P2_U2538 , P2_U2539 , P2_U2540 , P2_U2541;
wire P2_U2542 , P2_U2543 , P2_U2544 , P2_U2545 , P2_U2546 , P2_U2547 , P2_U2548 , P2_U2549 , P2_U2550 , P2_U2551;
wire P2_U2552 , P2_U2553 , P2_U2554 , P2_U2555 , P2_U2556 , P2_U2557 , P2_U2558 , P2_U2559 , P2_U2560 , P2_U2561;
wire P2_U2562 , P2_U2563 , P2_U2564 , P2_U2565 , P2_U2566 , P2_U2567 , P2_U2568 , P2_U2569 , P2_U2570 , P2_U2571;
wire P2_U2572 , P2_U2573 , P2_U2574 , P2_U2575 , P2_U2576 , P2_U2577 , P2_U2578 , P2_U2579 , P2_U2580 , P2_U2581;
wire P2_U2582 , P2_U2583 , P2_U2584 , P2_U2585 , P2_U2586 , P2_U2587 , P2_U2588 , P2_U2589 , P2_U2590 , P2_U2591;
wire P2_U2592 , P2_U2593 , P2_U2594 , P2_U2595 , P2_U2596 , P2_U2597 , P2_U2598 , P2_U2599 , P2_U2600 , P2_U2601;
wire P2_U2602 , P2_U2603 , P2_U2604 , P2_U2605 , P2_U2606 , P2_U2607 , P2_U2608 , P2_U2609 , P2_U2610 , P2_U2611;
wire P2_U2612 , P2_U2613 , P2_U2614 , P2_U2615 , P2_U2616 , P2_U2617 , P2_U2618 , P2_U2619 , P2_U2620 , P2_U2621;
wire P2_U2622 , P2_U2623 , P2_U2624 , P2_U2625 , P2_U2626 , P2_U2627 , P2_U2628 , P2_U2629 , P2_U2630 , P2_U2631;
wire P2_U2632 , P2_U2633 , P2_U2634 , P2_U2635 , P2_U2636 , P2_U2637 , P2_U2638 , P2_U2639 , P2_U2640 , P2_U2641;
wire P2_U2642 , P2_U2643 , P2_U2644 , P2_U2645 , P2_U2646 , P2_U2647 , P2_U2648 , P2_U2649 , P2_U2650 , P2_U2651;
wire P2_U2652 , P2_U2653 , P2_U2654 , P2_U2655 , P2_U2656 , P2_U2657 , P2_U2658 , P2_U2659 , P2_U2660 , P2_U2661;
wire P2_U2662 , P2_U2663 , P2_U2664 , P2_U2665 , P2_U2666 , P2_U2667 , P2_U2668 , P2_U2669 , P2_U2670 , P2_U2671;
wire P2_U2672 , P2_U2673 , P2_U2674 , P2_U2675 , P2_U2676 , P2_U2677 , P2_U2678 , P2_U2679 , P2_U2680 , P2_U2681;
wire P2_U2682 , P2_U2683 , P2_U2684 , P2_U2685 , P2_U2686 , P2_U2687 , P2_U2688 , P2_U2689 , P2_U2690 , P2_U2691;
wire P2_U2692 , P2_U2693 , P2_U2694 , P2_U2695 , P2_U2696 , P1_ADD_405_U172 , P2_U2698 , P2_U2699 , P2_U2700 , P2_U2701;
wire P2_U2702 , P2_U2703 , P2_U2704 , P2_U2705 , P2_U2706 , P2_U2707 , P2_U2708 , P2_U2709 , P2_U2710 , P2_U2711;
wire P2_U2712 , P2_U2713 , P2_U2714 , P2_U2715 , P2_U2716 , P2_U2717 , P2_U2718 , P2_U2719 , P2_U2720 , P2_U2721;
wire P2_U2722 , P2_U2723 , P2_U2724 , P2_U2725 , P2_U2726 , P2_U2727 , P2_U2728 , P2_U2729 , P2_U2730 , P2_U2731;
wire P2_U2732 , P2_U2733 , P2_U2734 , P2_U2735 , P2_U2736 , P2_U2737 , P2_U2738 , P2_U2739 , P2_U2740 , P2_U2741;
wire P2_U2742 , P2_U2743 , P2_U2744 , P2_U2745 , P2_U2746 , P2_U2747 , P2_U2748 , P2_U2749 , P2_U2750 , P2_U2751;
wire P2_U2752 , P2_U2753 , P2_U2754 , P2_U2755 , P2_U2756 , P2_U2757 , P2_U2758 , P2_U2759 , P2_U2760 , P2_U2761;
wire P2_U2762 , P2_U2763 , P2_U2764 , P2_U2765 , P2_U2766 , P2_U2767 , P2_U2768 , P2_U2769 , P2_U2770 , P2_U2771;
wire P2_U2772 , P2_U2773 , P2_U2774 , P2_U2775 , P2_U2776 , P2_U2777 , P2_U2778 , P2_U2779 , P2_U2780 , P2_U2781;
wire P2_U2782 , P2_U2783 , P2_U2784 , P2_U2785 , P2_U2786 , P2_U2787 , P2_U2788 , P2_U2789 , P2_U2790 , P2_U2791;
wire P2_U2792 , P2_U2793 , P2_U2794 , P2_U2795 , P2_U2796 , P2_U2797 , P2_U2798 , P2_U2799 , P2_U2800 , P2_U2801;
wire P2_U2802 , P2_U2803 , P2_U2804 , P2_U2805 , P2_U2806 , P2_U2807 , P2_U2808 , P2_U2809 , P2_U2810 , P2_U2811;
wire P2_U2812 , P2_U2813 , P2_U3242 , P2_U3243 , P2_U3244 , P2_U3245 , P2_U3246 , P2_U3247 , P2_U3248 , P2_U3249;
wire P2_U3250 , P2_U3251 , P2_U3252 , P2_U3253 , P2_U3254 , P2_U3255 , P2_U3256 , P2_U3257 , P2_U3258 , P2_U3259;
wire P2_U3260 , P2_U3261 , P2_U3262 , P2_U3263 , P2_U3264 , P2_U3265 , P2_U3266 , P2_U3267 , P2_U3268 , P2_U3269;
wire P2_U3270 , P2_U3271 , P2_U3272 , P2_U3273 , P2_U3274 , P2_U3275 , P2_U3276 , P2_U3277 , P2_U3278 , P2_U3279;
wire P2_U3280 , P2_U3281 , P2_U3282 , P2_U3283 , P2_U3284 , P2_U3285 , P2_U3286 , P2_U3287 , P2_U3288 , P2_U3289;
wire P2_U3290 , P2_U3291 , P2_U3292 , P2_U3293 , P2_U3294 , P2_U3295 , P2_U3296 , P2_U3297 , P2_U3298 , P2_U3299;
wire P2_U3300 , P2_U3301 , P2_U3302 , P2_U3303 , P2_U3304 , P2_U3305 , P2_U3306 , P2_U3307 , P2_U3308 , P2_U3309;
wire P2_U3310 , P2_U3311 , P2_U3312 , P2_U3313 , P2_U3314 , P2_U3315 , P2_U3316 , P2_U3317 , P2_U3318 , P2_U3319;
wire P2_U3320 , P2_U3321 , P2_U3322 , P2_U3323 , P2_U3324 , P2_U3325 , P2_U3326 , P2_U3327 , P2_U3328 , P2_U3329;
wire P2_U3330 , P2_U3331 , P2_U3332 , P2_U3333 , P2_U3334 , P2_U3335 , P2_U3336 , P2_U3337 , P2_U3338 , P2_U3339;
wire P2_U3340 , P2_U3341 , P2_U3342 , P2_U3343 , P2_U3344 , P2_U3345 , P2_U3346 , P2_U3347 , P2_U3348 , P2_U3349;
wire P2_U3350 , P2_U3351 , P2_U3352 , P2_U3353 , P2_U3354 , P2_U3355 , P2_U3356 , P2_U3357 , P2_U3358 , P2_U3359;
wire P2_U3360 , P2_U3361 , P2_U3362 , P2_U3363 , P2_U3364 , P2_U3365 , P2_U3366 , P2_U3367 , P2_U3368 , P2_U3369;
wire P2_U3370 , P2_U3371 , P2_U3372 , P2_U3373 , P2_U3374 , P2_U3375 , P2_U3376 , P2_U3377 , P2_U3378 , P2_U3379;
wire P2_U3380 , P2_U3381 , P2_U3382 , P2_U3383 , P2_U3384 , P2_U3385 , P2_U3386 , P2_U3387 , P2_U3388 , P2_U3389;
wire P2_U3390 , P2_U3391 , P2_U3392 , P2_U3393 , P2_U3394 , P2_U3395 , P2_U3396 , P2_U3397 , P2_U3398 , P2_U3399;
wire P2_U3400 , P2_U3401 , P2_U3402 , P2_U3403 , P2_U3404 , P2_U3405 , P2_U3406 , P2_U3407 , P2_U3408 , P2_U3409;
wire P2_U3410 , P2_U3411 , P2_U3412 , P2_U3413 , P2_U3414 , P2_U3415 , P2_U3416 , P2_U3417 , P2_U3418 , P2_U3419;
wire P2_U3420 , P2_U3421 , P2_U3422 , P2_U3423 , P2_U3424 , P2_U3425 , P2_U3426 , P2_U3427 , P2_U3428 , P2_U3429;
wire P2_U3430 , P2_U3431 , P2_U3432 , P2_U3433 , P2_U3434 , P2_U3435 , P2_U3436 , P2_U3437 , P2_U3438 , P2_U3439;
wire P2_U3440 , P2_U3441 , P2_U3442 , P2_U3443 , P2_U3444 , P2_U3445 , P2_U3446 , P2_U3447 , P2_U3448 , P2_U3449;
wire P2_U3450 , P2_U3451 , P2_U3452 , P2_U3453 , P2_U3454 , P2_U3455 , P2_U3456 , P2_U3457 , P2_U3458 , P2_U3459;
wire P2_U3460 , P2_U3461 , P2_U3462 , P2_U3463 , P2_U3464 , P2_U3465 , P2_U3466 , P2_U3467 , P2_U3468 , P2_U3469;
wire P2_U3470 , P2_U3471 , P2_U3472 , P2_U3473 , P2_U3474 , P2_U3475 , P2_U3476 , P2_U3477 , P2_U3478 , P2_U3479;
wire P2_U3480 , P2_U3481 , P2_U3482 , P2_U3483 , P2_U3484 , P2_U3485 , P2_U3486 , P2_U3487 , P2_U3488 , P2_U3489;
wire P2_U3490 , P2_U3491 , P2_U3492 , P2_U3493 , P2_U3494 , P2_U3495 , P2_U3496 , P2_U3497 , P2_U3498 , P2_U3499;
wire P2_U3500 , P2_U3501 , P2_U3502 , P2_U3503 , P2_U3504 , P2_U3505 , P2_U3506 , P2_U3507 , P2_U3508 , P2_U3509;
wire P2_U3510 , P2_U3511 , P2_U3512 , P2_U3513 , P2_U3514 , P2_U3515 , P2_U3516 , P2_U3517 , P2_U3518 , P2_U3519;
wire P2_U3520 , P2_U3521 , P2_U3522 , P2_U3523 , P2_U3524 , P2_U3525 , P2_U3526 , P2_U3527 , P2_U3528 , P2_U3529;
wire P2_U3530 , P2_U3531 , P2_U3532 , P2_U3533 , P2_U3534 , P2_U3535 , P2_U3536 , P2_U3537 , P2_U3538 , P2_U3539;
wire P2_U3540 , P2_U3541 , P2_U3542 , P2_U3543 , P2_U3544 , P2_U3545 , P2_U3546 , P2_U3547 , P2_U3548 , P2_U3549;
wire P2_U3550 , P2_U3551 , P2_U3552 , P2_U3553 , P2_U3554 , P2_U3555 , P2_U3556 , P2_U3557 , P2_U3558 , P2_U3559;
wire P2_U3560 , P2_U3561 , P2_U3562 , P2_U3563 , P2_U3564 , P2_U3565 , P2_U3566 , P2_U3567 , P2_U3568 , P2_U3569;
wire P2_U3570 , P2_U3571 , P2_U3572 , P2_U3573 , P2_U3574 , P2_U3575 , P2_U3576 , P2_U3577 , P2_U3578 , P2_U3579;
wire P2_U3580 , P2_U3581 , P2_U3582 , P2_U3583 , P2_U3584 , P2_U3589 , P2_U3590 , P2_U3594 , P2_U3597 , P2_U3598;
wire P2_U3606 , P2_U3607 , P2_U3613 , P2_U3614 , P2_U3615 , P2_U3616 , P2_U3617 , P2_U3618 , P2_U3619 , P2_U3620;
wire P2_U3621 , P2_U3622 , P2_U3623 , P2_U3624 , P2_U3625 , P2_U3626 , P2_U3627 , P2_U3628 , P2_U3629 , P2_U3630;
wire P2_U3631 , P2_U3632 , P2_U3633 , P2_U3634 , P2_U3635 , P2_U3636 , P2_U3637 , P2_U3638 , P2_U3639 , P2_U3640;
wire P2_U3641 , P2_U3642 , P2_U3643 , P2_U3644 , P2_U3645 , P2_U3646 , P2_U3647 , P2_U3648 , P2_U3649 , P2_U3650;
wire P2_U3651 , P2_U3652 , P2_U3653 , P2_U3654 , P2_U3655 , P2_U3656 , P2_U3657 , P2_U3658 , P2_U3659 , P2_U3660;
wire P2_U3661 , P2_U3662 , P2_U3663 , P2_U3664 , P2_U3665 , P2_U3666 , P2_U3667 , P2_U3668 , P2_U3669 , P2_U3670;
wire P2_U3671 , P2_U3672 , P2_U3673 , P2_U3674 , P2_U3675 , P2_U3676 , P2_U3677 , P2_U3678 , P2_U3679 , P2_U3680;
wire P2_U3681 , P2_U3682 , P2_U3683 , P2_U3684 , P2_U3685 , P2_U3686 , P2_U3687 , P2_U3688 , P2_U3689 , P2_U3690;
wire P2_U3691 , P2_U3692 , P2_U3693 , P2_U3694 , P2_U3695 , P2_U3696 , P2_U3697 , P2_U3698 , P2_U3699 , P2_U3700;
wire P2_U3701 , P2_U3702 , P2_U3703 , P2_U3704 , P2_U3705 , P2_U3706 , P2_U3707 , P2_U3708 , P2_U3709 , P2_U3710;
wire P2_U3711 , P2_U3712 , P2_U3713 , P2_U3714 , P2_U3715 , P2_U3716 , P2_U3717 , P2_U3718 , P2_U3719 , P2_U3720;
wire P2_U3721 , P2_U3722 , P2_U3723 , P2_U3724 , P2_U3725 , P2_U3726 , P2_U3727 , P2_U3728 , P2_U3729 , P2_U3730;
wire P2_U3731 , P2_U3732 , P2_U3733 , P2_U3734 , P2_U3735 , P2_U3736 , P2_U3737 , P2_U3738 , P2_U3739 , P2_U3740;
wire P2_U3741 , P2_U3742 , P2_U3743 , P2_U3744 , P2_U3745 , P2_U3746 , P2_U3747 , P2_U3748 , P2_U3749 , P2_U3750;
wire P2_U3751 , P2_U3752 , P2_U3753 , P2_U3754 , P2_U3755 , P2_U3756 , P2_U3757 , P2_U3758 , P2_U3759 , P2_U3760;
wire P2_U3761 , P2_U3762 , P2_U3763 , P2_U3764 , P2_U3765 , P2_U3766 , P2_U3767 , P2_U3768 , P2_U3769 , P2_U3770;
wire P2_U3771 , P2_U3772 , P2_U3773 , P2_U3774 , P2_U3775 , P2_U3776 , P2_U3777 , P2_U3778 , P2_U3779 , P2_U3780;
wire P2_U3781 , P2_U3782 , P2_U3783 , P2_U3784 , P2_U3785 , P2_U3786 , P2_U3787 , P2_U3788 , P2_U3789 , P2_U3790;
wire P2_U3791 , P2_U3792 , P2_U3793 , P2_U3794 , P2_U3795 , P2_U3796 , P2_U3797 , P2_U3798 , P2_U3799 , P2_U3800;
wire P2_U3801 , P2_U3802 , P2_U3803 , P2_U3804 , P2_U3805 , P2_U3806 , P2_U3807 , P2_U3808 , P2_U3809 , P2_U3810;
wire P2_U3811 , P2_U3812 , P2_U3813 , P2_U3814 , P2_U3815 , P2_U3816 , P2_U3817 , P2_U3818 , P2_U3819 , P2_U3820;
wire P2_U3821 , P2_U3822 , P2_U3823 , P2_U3824 , P2_U3825 , P2_U3826 , P2_U3827 , P2_U3828 , P2_U3829 , P2_U3830;
wire P2_U3831 , P2_U3832 , P2_U3833 , P2_U3834 , P2_U3835 , P2_U3836 , P2_U3837 , P2_U3838 , P2_U3839 , P2_U3840;
wire P2_U3841 , P2_U3842 , P2_U3843 , P2_U3844 , P2_U3845 , P2_U3846 , P2_U3847 , P2_U3848 , P2_U3849 , P2_U3850;
wire P2_U3851 , P2_U3852 , P2_U3853 , P2_U3854 , P2_U3855 , P2_U3856 , P2_U3857 , P2_U3858 , P2_U3859 , P2_U3860;
wire P2_U3861 , P2_U3862 , P2_U3863 , P2_U3864 , P2_U3865 , P2_U3866 , P2_U3867 , P2_U3868 , P2_U3869 , P2_U3870;
wire P2_U3871 , P2_U3872 , P2_U3873 , P2_U3874 , P2_U3875 , P2_U3876 , P2_U3877 , P2_U3878 , P2_U3879 , P2_U3880;
wire P2_U3881 , P2_U3882 , P2_U3883 , P2_U3884 , P2_U3885 , P2_U3886 , P2_U3887 , P2_U3888 , P2_U3889 , P2_U3890;
wire P2_U3891 , P2_U3892 , P2_U3893 , P2_U3894 , P2_U3895 , P2_U3896 , P2_U3897 , P2_U3898 , P2_U3899 , P2_U3900;
wire P2_U3901 , P2_U3902 , P2_U3903 , P2_U3904 , P2_U3905 , P2_U3906 , P2_U3907 , P2_U3908 , P2_U3909 , P2_U3910;
wire P2_U3911 , P2_U3912 , P2_U3913 , P2_U3914 , P2_U3915 , P2_U3916 , P2_U3917 , P2_U3918 , P2_U3919 , P2_U3920;
wire P2_U3921 , P2_U3922 , P2_U3923 , P2_U3924 , P2_U3925 , P2_U3926 , P2_U3927 , P2_U3928 , P2_U3929 , P2_U3930;
wire P2_U3931 , P2_U3932 , P2_U3933 , P2_U3934 , P2_U3935 , P2_U3936 , P2_U3937 , P2_U3938 , P2_U3939 , P2_U3940;
wire P2_U3941 , P2_U3942 , P2_U3943 , P2_U3944 , P2_U3945 , P2_U3946 , P2_U3947 , P2_U3948 , P2_U3949 , P2_U3950;
wire P2_U3951 , P2_U3952 , P2_U3953 , P2_U3954 , P2_U3955 , P2_U3956 , P2_U3957 , P2_U3958 , P2_U3959 , P2_U3960;
wire P2_U3961 , P2_U3962 , P2_U3963 , P2_U3964 , P2_U3965 , P2_U3966 , P2_U3967 , P2_U3968 , P2_U3969 , P2_U3970;
wire P2_U3971 , P2_U3972 , P2_U3973 , P2_U3974 , P2_U3975 , P2_U3976 , P2_U3977 , P2_U3978 , P2_U3979 , P2_U3980;
wire P2_U3981 , P2_U3982 , P2_U3983 , P2_U3984 , P2_U3985 , P2_U3986 , P2_U3987 , P2_U3988 , P2_U3989 , P2_U3990;
wire P2_U3991 , P2_U3992 , P2_U3993 , P2_U3994 , P2_U3995 , P2_U3996 , P2_U3997 , P2_U3998 , P2_U3999 , P2_U4000;
wire P2_U4001 , P2_U4002 , P2_U4003 , P2_U4004 , P2_U4005 , P2_U4006 , P2_U4007 , P2_U4008 , P2_U4009 , P2_U4010;
wire P2_U4011 , P2_U4012 , P2_U4013 , P2_U4014 , P2_U4015 , P2_U4016 , P2_U4017 , P2_U4018 , P2_U4019 , P2_U4020;
wire P2_U4021 , P2_U4022 , P2_U4023 , P2_U4024 , P2_U4025 , P2_U4026 , P2_U4027 , P2_U4028 , P2_U4029 , P2_U4030;
wire P2_U4031 , P2_U4032 , P2_U4033 , P2_U4034 , P2_U4035 , P2_U4036 , P2_U4037 , P2_U4038 , P2_U4039 , P2_U4040;
wire P2_U4041 , P2_U4042 , P2_U4043 , P2_U4044 , P2_U4045 , P2_U4046 , P2_U4047 , P2_U4048 , P2_U4049 , P2_U4050;
wire P2_U4051 , P2_U4052 , P2_U4053 , P2_U4054 , P2_U4055 , P2_U4056 , P2_U4057 , P2_U4058 , P2_U4059 , P2_U4060;
wire P2_U4061 , P2_U4062 , P2_U4063 , P2_U4064 , P2_U4065 , P2_U4066 , P2_U4067 , P2_U4068 , P2_U4069 , P2_U4070;
wire P2_U4071 , P2_U4072 , P2_U4073 , P2_U4074 , P2_U4075 , P2_U4076 , P2_U4077 , P2_U4078 , P2_U4079 , P2_U4080;
wire P2_U4081 , P2_U4082 , P2_U4083 , P2_U4084 , P2_U4085 , P2_U4086 , P2_U4087 , P2_U4088 , P2_U4089 , P2_U4090;
wire P2_U4091 , P2_U4092 , P2_U4093 , P2_U4094 , P2_U4095 , P2_U4096 , P2_U4097 , P2_U4098 , P2_U4099 , P2_U4100;
wire P2_U4101 , P2_U4102 , P2_U4103 , P2_U4104 , P2_U4105 , P2_U4106 , P2_U4107 , P2_U4108 , P2_U4109 , P2_U4110;
wire P2_U4111 , P2_U4112 , P2_U4113 , P2_U4114 , P2_U4115 , P2_U4116 , P2_U4117 , P2_U4118 , P2_U4119 , P2_U4120;
wire P2_U4121 , P2_U4122 , P2_U4123 , P2_U4124 , P2_U4125 , P2_U4126 , P2_U4127 , P2_U4128 , P2_U4129 , P2_U4130;
wire P2_U4131 , P2_U4132 , P2_U4133 , P2_U4134 , P2_U4135 , P2_U4136 , P2_U4137 , P2_U4138 , P2_U4139 , P2_U4140;
wire P2_U4141 , P2_U4142 , P2_U4143 , P2_U4144 , P2_U4145 , P2_U4146 , P2_U4147 , P2_U4148 , P2_U4149 , P2_U4150;
wire P2_U4151 , P2_U4152 , P2_U4153 , P2_U4154 , P2_U4155 , P2_U4156 , P2_U4157 , P2_U4158 , P2_U4159 , P2_U4160;
wire P2_U4161 , P2_U4162 , P2_U4163 , P2_U4164 , P2_U4165 , P2_U4166 , P2_U4167 , P2_U4168 , P2_U4169 , P2_U4170;
wire P2_U4171 , P2_U4172 , P2_U4173 , P2_U4174 , P2_U4175 , P2_U4176 , P2_U4177 , P2_U4178 , P2_U4179 , P2_U4180;
wire P2_U4181 , P2_U4182 , P2_U4183 , P2_U4184 , P2_U4185 , P2_U4186 , P2_U4187 , P2_U4188 , P2_U4189 , P2_U4190;
wire P2_U4191 , P2_U4192 , P2_U4193 , P2_U4194 , P2_U4195 , P2_U4196 , P2_U4197 , P2_U4198 , P2_U4199 , P2_U4200;
wire P2_U4201 , P2_U4202 , P2_U4203 , P2_U4204 , P2_U4205 , P2_U4206 , P2_U4207 , P2_U4208 , P2_U4209 , P2_U4210;
wire P2_U4211 , P2_U4212 , P2_U4213 , P2_U4214 , P2_U4215 , P2_U4216 , P2_U4217 , P2_U4218 , P2_U4219 , P2_U4220;
wire P2_U4221 , P2_U4222 , P2_U4223 , P2_U4224 , P2_U4225 , P2_U4226 , P2_U4227 , P2_U4228 , P2_U4229 , P2_U4230;
wire P2_U4231 , P2_U4232 , P2_U4233 , P2_U4234 , P2_U4235 , P2_U4236 , P2_U4237 , P2_U4238 , P2_U4239 , P2_U4240;
wire P2_U4241 , P2_U4242 , P2_U4243 , P2_U4244 , P2_U4245 , P2_U4246 , P2_U4247 , P2_U4248 , P2_U4249 , P2_U4250;
wire P2_U4251 , P2_U4252 , P2_U4253 , P2_U4254 , P2_U4255 , P2_U4256 , P2_U4257 , P2_U4258 , P2_U4259 , P2_U4260;
wire P2_U4261 , P2_U4262 , P2_U4263 , P2_U4264 , P2_U4265 , P2_U4266 , P2_U4267 , P2_U4268 , P2_U4269 , P2_U4270;
wire P2_U4271 , P2_U4272 , P2_U4273 , P2_U4274 , P2_U4275 , P2_U4276 , P2_U4277 , P2_U4278 , P2_U4279 , P2_U4280;
wire P2_U4281 , P2_U4282 , P2_U4283 , P2_U4284 , P2_U4285 , P2_U4286 , P2_U4287 , P2_U4288 , P2_U4289 , P2_U4290;
wire P2_U4291 , P2_U4292 , P2_U4293 , P2_U4294 , P2_U4295 , P2_U4296 , P2_U4297 , P2_U4298 , P2_U4299 , P2_U4300;
wire P2_U4301 , P2_U4302 , P2_U4303 , P2_U4304 , P2_U4305 , P2_U4306 , P2_U4307 , P2_U4308 , P2_U4309 , P2_U4310;
wire P2_U4311 , P2_U4312 , P2_U4313 , P2_U4314 , P2_U4315 , P2_U4316 , P2_U4317 , P2_U4318 , P2_U4319 , P2_U4320;
wire P2_U4321 , P2_U4322 , P2_U4323 , P2_U4324 , P2_U4325 , P2_U4326 , P2_U4327 , P2_U4328 , P2_U4329 , P2_U4330;
wire P2_U4331 , P2_U4332 , P2_U4333 , P2_U4334 , P2_U4335 , P2_U4336 , P2_U4337 , P2_U4338 , P2_U4339 , P2_U4340;
wire P2_U4341 , P2_U4342 , P2_U4343 , P2_U4344 , P2_U4345 , P2_U4346 , P2_U4347 , P2_U4348 , P2_U4349 , P2_U4350;
wire P2_U4351 , P2_U4352 , P2_U4353 , P2_U4354 , P2_U4355 , P2_U4356 , P2_U4357 , P2_U4358 , P2_U4359 , P2_U4360;
wire P2_U4361 , P2_U4362 , P2_U4363 , P2_U4364 , P2_U4365 , P2_U4366 , P2_U4367 , P2_U4368 , P2_U4369 , P2_U4370;
wire P2_U4371 , P2_U4372 , P2_U4373 , P2_U4374 , P2_U4375 , P2_U4376 , P2_U4377 , P2_U4378 , P2_U4379 , P2_U4380;
wire P2_U4381 , P2_U4382 , P2_U4383 , P2_U4384 , P2_U4385 , P2_U4386 , P2_U4387 , P2_U4388 , P2_U4389 , P2_U4390;
wire P2_U4391 , P2_U4392 , P2_U4393 , P2_U4394 , P2_U4395 , P2_U4396 , P2_U4397 , P2_U4398 , P2_U4399 , P2_U4400;
wire P2_U4401 , P2_U4402 , P2_U4403 , P2_U4404 , P2_U4405 , P2_U4406 , P2_U4407 , P2_U4408 , P2_U4409 , P2_U4410;
wire P2_U4411 , P2_U4412 , P2_U4413 , P2_U4414 , P2_U4415 , P2_U4416 , P2_U4417 , P2_U4418 , P2_U4419 , P2_U4420;
wire P2_U4421 , P2_U4422 , P2_U4423 , P2_U4424 , P2_U4425 , P2_U4426 , P2_U4427 , P2_U4428 , P2_U4429 , P2_U4430;
wire P2_U4431 , P2_U4432 , P2_U4433 , P2_U4434 , P2_U4435 , P2_U4436 , P2_U4437 , P2_U4438 , P2_U4439 , P2_U4440;
wire P2_U4441 , P2_U4442 , P2_U4443 , P2_U4444 , P2_U4445 , P2_U4446 , P2_U4447 , P2_U4448 , P2_U4449 , P2_U4450;
wire P2_U4451 , P2_U4452 , P2_U4453 , P2_U4454 , P2_U4455 , P2_U4456 , P2_U4457 , P2_U4458 , P2_U4459 , P2_U4460;
wire P2_U4461 , P2_U4462 , P2_U4463 , P2_U4464 , P2_U4465 , P2_U4466 , P2_U4467 , P2_U4468 , P2_U4469 , P2_U4470;
wire P2_U4471 , P2_U4472 , P2_U4473 , P2_U4474 , P2_U4475 , P2_U4476 , P2_U4477 , P2_U4478 , P2_U4479 , P2_U4480;
wire P2_U4481 , P2_U4482 , P2_U4483 , P2_U4484 , P2_U4485 , P2_U4486 , P2_U4487 , P2_U4488 , P2_U4489 , P2_U4490;
wire P2_U4491 , P2_U4492 , P2_U4493 , P2_U4494 , P2_U4495 , P2_U4496 , P2_U4497 , P2_U4498 , P2_U4499 , P2_U4500;
wire P2_U4501 , P2_U4502 , P2_U4503 , P2_U4504 , P2_U4505 , P2_U4506 , P2_U4507 , P2_U4508 , P2_U4509 , P2_U4510;
wire P2_U4511 , P2_U4512 , P2_U4513 , P2_U4514 , P2_U4515 , P2_U4516 , P2_U4517 , P2_U4518 , P2_U4519 , P2_U4520;
wire P2_U4521 , P2_U4522 , P2_U4523 , P2_U4524 , P2_U4525 , P2_U4526 , P2_U4527 , P2_U4528 , P2_U4529 , P2_U4530;
wire P2_U4531 , P2_U4532 , P2_U4533 , P2_U4534 , P2_U4535 , P2_U4536 , P2_U4537 , P2_U4538 , P2_U4539 , P2_U4540;
wire P2_U4541 , P2_U4542 , P2_U4543 , P2_U4544 , P2_U4545 , P2_U4546 , P2_U4547 , P2_U4548 , P2_U4549 , P2_U4550;
wire P2_U4551 , P2_U4552 , P2_U4553 , P2_U4554 , P2_U4555 , P2_U4556 , P2_U4557 , P2_U4558 , P2_U4559 , P2_U4560;
wire P2_U4561 , P2_U4562 , P2_U4563 , P2_U4564 , P2_U4565 , P2_U4566 , P2_U4567 , P2_U4568 , P2_U4569 , P2_U4570;
wire P2_U4571 , P2_U4572 , P2_U4573 , P2_U4574 , P2_U4575 , P2_U4576 , P2_U4577 , P2_U4578 , P2_U4579 , P2_U4580;
wire P2_U4581 , P2_U4582 , P2_U4583 , P2_U4584 , P2_U4585 , P2_U4586 , P2_U4587 , P2_U4588 , P2_U4589 , P2_U4590;
wire P2_U4591 , P2_U4592 , P2_U4593 , P2_U4594 , P2_U4595 , P2_U4596 , P2_U4597 , P2_U4598 , P2_U4599 , P2_U4600;
wire P2_U4601 , P2_U4602 , P2_U4603 , P2_U4604 , P2_U4605 , P2_U4606 , P2_U4607 , P2_U4608 , P2_U4609 , P2_U4610;
wire P2_U4611 , P2_U4612 , P2_U4613 , P2_U4614 , P2_U4615 , P2_U4616 , P2_U4617 , P2_U4618 , P2_U4619 , P2_U4620;
wire P2_U4621 , P2_U4622 , P2_U4623 , P2_U4624 , P2_U4625 , P2_U4626 , P2_U4627 , P2_U4628 , P2_U4629 , P2_U4630;
wire P2_U4631 , P2_U4632 , P2_U4633 , P2_U4634 , P2_U4635 , P2_U4636 , P2_U4637 , P2_U4638 , P2_U4639 , P2_U4640;
wire P2_U4641 , P2_U4642 , P2_U4643 , P2_U4644 , P2_U4645 , P2_U4646 , P2_U4647 , P2_U4648 , P2_U4649 , P2_U4650;
wire P2_U4651 , P2_U4652 , P2_U4653 , P2_U4654 , P2_U4655 , P2_U4656 , P2_U4657 , P2_U4658 , P2_U4659 , P2_U4660;
wire P2_U4661 , P2_U4662 , P2_U4663 , P2_U4664 , P2_U4665 , P2_U4666 , P2_U4667 , P2_U4668 , P2_U4669 , P2_U4670;
wire P2_U4671 , P2_U4672 , P2_U4673 , P2_U4674 , P2_U4675 , P2_U4676 , P2_U4677 , P2_U4678 , P2_U4679 , P2_U4680;
wire P2_U4681 , P2_U4682 , P2_U4683 , P2_U4684 , P2_U4685 , P2_U4686 , P2_U4687 , P2_U4688 , P2_U4689 , P2_U4690;
wire P2_U4691 , P2_U4692 , P2_U4693 , P2_U4694 , P2_U4695 , P2_U4696 , P2_U4697 , P2_U4698 , P2_U4699 , P2_U4700;
wire P2_U4701 , P2_U4702 , P2_U4703 , P2_U4704 , P2_U4705 , P2_U4706 , P2_U4707 , P2_U4708 , P2_U4709 , P2_U4710;
wire P2_U4711 , P2_U4712 , P2_U4713 , P2_U4714 , P2_U4715 , P2_U4716 , P2_U4717 , P2_U4718 , P2_U4719 , P2_U4720;
wire P2_U4721 , P2_U4722 , P2_U4723 , P2_U4724 , P2_U4725 , P2_U4726 , P2_U4727 , P2_U4728 , P2_U4729 , P2_U4730;
wire P2_U4731 , P2_U4732 , P2_U4733 , P2_U4734 , P2_U4735 , P2_U4736 , P2_U4737 , P2_U4738 , P2_U4739 , P2_U4740;
wire P2_U4741 , P2_U4742 , P2_U4743 , P2_U4744 , P2_U4745 , P2_U4746 , P2_U4747 , P2_U4748 , P2_U4749 , P2_U4750;
wire P2_U4751 , P2_U4752 , P2_U4753 , P2_U4754 , P2_U4755 , P2_U4756 , P2_U4757 , P2_U4758 , P2_U4759 , P2_U4760;
wire P2_U4761 , P2_U4762 , P2_U4763 , P2_U4764 , P2_U4765 , P2_U4766 , P2_U4767 , P2_U4768 , P2_U4769 , P2_U4770;
wire P2_U4771 , P2_U4772 , P2_U4773 , P2_U4774 , P2_U4775 , P2_U4776 , P2_U4777 , P2_U4778 , P2_U4779 , P2_U4780;
wire P2_U4781 , P2_U4782 , P2_U4783 , P2_U4784 , P2_U4785 , P2_U4786 , P2_U4787 , P2_U4788 , P2_U4789 , P2_U4790;
wire P2_U4791 , P2_U4792 , P2_U4793 , P2_U4794 , P2_U4795 , P2_U4796 , P2_U4797 , P2_U4798 , P2_U4799 , P2_U4800;
wire P2_U4801 , P2_U4802 , P2_U4803 , P2_U4804 , P2_U4805 , P2_U4806 , P2_U4807 , P2_U4808 , P2_U4809 , P2_U4810;
wire P2_U4811 , P2_U4812 , P2_U4813 , P2_U4814 , P2_U4815 , P2_U4816 , P2_U4817 , P2_U4818 , P2_U4819 , P2_U4820;
wire P2_U4821 , P2_U4822 , P2_U4823 , P2_U4824 , P2_U4825 , P2_U4826 , P2_U4827 , P2_U4828 , P2_U4829 , P2_U4830;
wire P2_U4831 , P2_U4832 , P2_U4833 , P2_U4834 , P2_U4835 , P2_U4836 , P2_U4837 , P2_U4838 , P2_U4839 , P2_U4840;
wire P2_U4841 , P2_U4842 , P2_U4843 , P2_U4844 , P2_U4845 , P2_U4846 , P2_U4847 , P2_U4848 , P2_U4849 , P2_U4850;
wire P2_U4851 , P2_U4852 , P2_U4853 , P2_U4854 , P2_U4855 , P2_U4856 , P2_U4857 , P2_U4858 , P2_U4859 , P2_U4860;
wire P2_U4861 , P2_U4862 , P2_U4863 , P2_U4864 , P2_U4865 , P2_U4866 , P2_U4867 , P2_U4868 , P2_U4869 , P2_U4870;
wire P2_U4871 , P2_U4872 , P2_U4873 , P2_U4874 , P2_U4875 , P2_U4876 , P2_U4877 , P2_U4878 , P2_U4879 , P2_U4880;
wire P2_U4881 , P2_U4882 , P2_U4883 , P2_U4884 , P2_U4885 , P2_U4886 , P2_U4887 , P2_U4888 , P2_U4889 , P2_U4890;
wire P2_U4891 , P2_U4892 , P2_U4893 , P2_U4894 , P2_U4895 , P2_U4896 , P2_U4897 , P2_U4898 , P2_U4899 , P2_U4900;
wire P2_U4901 , P2_U4902 , P2_U4903 , P2_U4904 , P2_U4905 , P2_U4906 , P2_U4907 , P2_U4908 , P2_U4909 , P2_U4910;
wire P2_U4911 , P2_U4912 , P2_U4913 , P2_U4914 , P2_U4915 , P2_U4916 , P2_U4917 , P2_U4918 , P2_U4919 , P2_U4920;
wire P2_U4921 , P2_U4922 , P2_U4923 , P2_U4924 , P2_U4925 , P2_U4926 , P2_U4927 , P2_U4928 , P2_U4929 , P2_U4930;
wire P2_U4931 , P2_U4932 , P2_U4933 , P2_U4934 , P2_U4935 , P2_U4936 , P2_U4937 , P2_U4938 , P2_U4939 , P2_U4940;
wire P2_U4941 , P2_U4942 , P2_U4943 , P2_U4944 , P2_U4945 , P2_U4946 , P2_U4947 , P2_U4948 , P2_U4949 , P2_U4950;
wire P2_U4951 , P2_U4952 , P2_U4953 , P2_U4954 , P2_U4955 , P2_U4956 , P2_U4957 , P2_U4958 , P2_U4959 , P2_U4960;
wire P2_U4961 , P2_U4962 , P2_U4963 , P2_U4964 , P2_U4965 , P2_U4966 , P2_U4967 , P2_U4968 , P2_U4969 , P2_U4970;
wire P2_U4971 , P2_U4972 , P2_U4973 , P2_U4974 , P2_U4975 , P2_U4976 , P2_U4977 , P2_U4978 , P2_U4979 , P2_U4980;
wire P2_U4981 , P2_U4982 , P2_U4983 , P2_U4984 , P2_U4985 , P2_U4986 , P2_U4987 , P2_U4988 , P2_U4989 , P2_U4990;
wire P2_U4991 , P2_U4992 , P2_U4993 , P2_U4994 , P2_U4995 , P2_U4996 , P2_U4997 , P2_U4998 , P2_U4999 , P2_U5000;
wire P2_U5001 , P2_U5002 , P2_U5003 , P2_U5004 , P2_U5005 , P2_U5006 , P2_U5007 , P2_U5008 , P2_U5009 , P2_U5010;
wire P2_U5011 , P2_U5012 , P2_U5013 , P2_U5014 , P2_U5015 , P2_U5016 , P2_U5017 , P2_U5018 , P2_U5019 , P2_U5020;
wire P2_U5021 , P2_U5022 , P2_U5023 , P2_U5024 , P2_U5025 , P2_U5026 , P2_U5027 , P2_U5028 , P2_U5029 , P2_U5030;
wire P2_U5031 , P2_U5032 , P2_U5033 , P2_U5034 , P2_U5035 , P2_U5036 , P2_U5037 , P2_U5038 , P2_U5039 , P2_U5040;
wire P2_U5041 , P2_U5042 , P2_U5043 , P2_U5044 , P2_U5045 , P2_U5046 , P2_U5047 , P2_U5048 , P2_U5049 , P2_U5050;
wire P2_U5051 , P2_U5052 , P2_U5053 , P2_U5054 , P2_U5055 , P2_U5056 , P2_U5057 , P2_U5058 , P2_U5059 , P2_U5060;
wire P2_U5061 , P2_U5062 , P2_U5063 , P2_U5064 , P2_U5065 , P2_U5066 , P2_U5067 , P2_U5068 , P2_U5069 , P2_U5070;
wire P2_U5071 , P2_U5072 , P2_U5073 , P2_U5074 , P2_U5075 , P2_U5076 , P2_U5077 , P2_U5078 , P2_U5079 , P2_U5080;
wire P2_U5081 , P2_U5082 , P2_U5083 , P2_U5084 , P2_U5085 , P2_U5086 , P2_U5087 , P2_U5088 , P2_U5089 , P2_U5090;
wire P2_U5091 , P2_U5092 , P2_U5093 , P2_U5094 , P2_U5095 , P2_U5096 , P2_U5097 , P2_U5098 , P2_U5099 , P2_U5100;
wire P2_U5101 , P2_U5102 , P2_U5103 , P2_U5104 , P2_U5105 , P2_U5106 , P2_U5107 , P2_U5108 , P2_U5109 , P2_U5110;
wire P2_U5111 , P2_U5112 , P2_U5113 , P2_U5114 , P2_U5115 , P2_U5116 , P2_U5117 , P2_U5118 , P2_U5119 , P2_U5120;
wire P2_U5121 , P2_U5122 , P2_U5123 , P2_U5124 , P2_U5125 , P2_U5126 , P2_U5127 , P2_U5128 , P2_U5129 , P2_U5130;
wire P2_U5131 , P2_U5132 , P2_U5133 , P2_U5134 , P2_U5135 , P2_U5136 , P2_U5137 , P2_U5138 , P2_U5139 , P2_U5140;
wire P2_U5141 , P2_U5142 , P2_U5143 , P2_U5144 , P2_U5145 , P2_U5146 , P2_U5147 , P2_U5148 , P2_U5149 , P2_U5150;
wire P2_U5151 , P2_U5152 , P2_U5153 , P2_U5154 , P2_U5155 , P2_U5156 , P2_U5157 , P2_U5158 , P2_U5159 , P2_U5160;
wire P2_U5161 , P2_U5162 , P2_U5163 , P2_U5164 , P2_U5165 , P2_U5166 , P2_U5167 , P2_U5168 , P2_U5169 , P2_U5170;
wire P2_U5171 , P2_U5172 , P2_U5173 , P2_U5174 , P2_U5175 , P2_U5176 , P2_U5177 , P2_U5178 , P2_U5179 , P2_U5180;
wire P2_U5181 , P2_U5182 , P2_U5183 , P2_U5184 , P2_U5185 , P2_U5186 , P2_U5187 , P2_U5188 , P2_U5189 , P2_U5190;
wire P2_U5191 , P2_U5192 , P2_U5193 , P2_U5194 , P2_U5195 , P2_U5196 , P2_U5197 , P2_U5198 , P2_U5199 , P2_U5200;
wire P2_U5201 , P2_U5202 , P2_U5203 , P2_U5204 , P2_U5205 , P2_U5206 , P2_U5207 , P2_U5208 , P2_U5209 , P2_U5210;
wire P2_U5211 , P2_U5212 , P2_U5213 , P2_U5214 , P2_U5215 , P2_U5216 , P2_U5217 , P2_U5218 , P2_U5219 , P2_U5220;
wire P2_U5221 , P2_U5222 , P2_U5223 , P2_U5224 , P2_U5225 , P2_U5226 , P2_U5227 , P2_U5228 , P2_U5229 , P2_U5230;
wire P2_U5231 , P2_U5232 , P2_U5233 , P2_U5234 , P2_U5235 , P2_U5236 , P2_U5237 , P2_U5238 , P2_U5239 , P2_U5240;
wire P2_U5241 , P2_U5242 , P2_U5243 , P2_U5244 , P2_U5245 , P2_U5246 , P2_U5247 , P2_U5248 , P2_U5249 , P2_U5250;
wire P2_U5251 , P2_U5252 , P2_U5253 , P2_U5254 , P2_U5255 , P2_U5256 , P2_U5257 , P2_U5258 , P2_U5259 , P2_U5260;
wire P2_U5261 , P2_U5262 , P2_U5263 , P2_U5264 , P2_U5265 , P2_U5266 , P2_U5267 , P2_U5268 , P2_U5269 , P2_U5270;
wire P2_U5271 , P2_U5272 , P2_U5273 , P2_U5274 , P2_U5275 , P2_U5276 , P2_U5277 , P2_U5278 , P2_U5279 , P2_U5280;
wire P2_U5281 , P2_U5282 , P2_U5283 , P2_U5284 , P2_U5285 , P2_U5286 , P2_U5287 , P2_U5288 , P2_U5289 , P2_U5290;
wire P2_U5291 , P2_U5292 , P2_U5293 , P2_U5294 , P2_U5295 , P2_U5296 , P2_U5297 , P2_U5298 , P2_U5299 , P2_U5300;
wire P2_U5301 , P2_U5302 , P2_U5303 , P2_U5304 , P2_U5305 , P2_U5306 , P2_U5307 , P2_U5308 , P2_U5309 , P2_U5310;
wire P2_U5311 , P2_U5312 , P2_U5313 , P2_U5314 , P2_U5315 , P2_U5316 , P2_U5317 , P2_U5318 , P2_U5319 , P2_U5320;
wire P2_U5321 , P2_U5322 , P2_U5323 , P2_U5324 , P2_U5325 , P2_U5326 , P2_U5327 , P2_U5328 , P2_U5329 , P2_U5330;
wire P2_U5331 , P2_U5332 , P2_U5333 , P2_U5334 , P2_U5335 , P2_U5336 , P2_U5337 , P2_U5338 , P2_U5339 , P2_U5340;
wire P2_U5341 , P2_U5342 , P2_U5343 , P2_U5344 , P2_U5345 , P2_U5346 , P2_U5347 , P2_U5348 , P2_U5349 , P2_U5350;
wire P2_U5351 , P2_U5352 , P2_U5353 , P2_U5354 , P2_U5355 , P2_U5356 , P2_U5357 , P2_U5358 , P2_U5359 , P2_U5360;
wire P2_U5361 , P2_U5362 , P2_U5363 , P2_U5364 , P2_U5365 , P2_U5366 , P2_U5367 , P2_U5368 , P2_U5369 , P2_U5370;
wire P2_U5371 , P2_U5372 , P2_U5373 , P2_U5374 , P2_U5375 , P2_U5376 , P2_U5377 , P2_U5378 , P2_U5379 , P2_U5380;
wire P2_U5381 , P2_U5382 , P2_U5383 , P2_U5384 , P2_U5385 , P2_U5386 , P2_U5387 , P2_U5388 , P2_U5389 , P2_U5390;
wire P2_U5391 , P2_U5392 , P2_U5393 , P2_U5394 , P2_U5395 , P2_U5396 , P2_U5397 , P2_U5398 , P2_U5399 , P2_U5400;
wire P2_U5401 , P2_U5402 , P2_U5403 , P2_U5404 , P2_U5405 , P2_U5406 , P2_U5407 , P2_U5408 , P2_U5409 , P2_U5410;
wire P2_U5411 , P2_U5412 , P2_U5413 , P2_U5414 , P2_U5415 , P2_U5416 , P2_U5417 , P2_U5418 , P2_U5419 , P2_U5420;
wire P2_U5421 , P2_U5422 , P2_U5423 , P2_U5424 , P2_U5425 , P2_U5426 , P2_U5427 , P2_U5428 , P2_U5429 , P2_U5430;
wire P2_U5431 , P2_U5432 , P2_U5433 , P2_U5434 , P2_U5435 , P2_U5436 , P2_U5437 , P2_U5438 , P2_U5439 , P2_U5440;
wire P2_U5441 , P2_U5442 , P2_U5443 , P2_U5444 , P2_U5445 , P2_U5446 , P2_U5447 , P2_U5448 , P2_U5449 , P2_U5450;
wire P2_U5451 , P2_U5452 , P2_U5453 , P2_U5454 , P2_U5455 , P2_U5456 , P2_U5457 , P2_U5458 , P2_U5459 , P2_U5460;
wire P2_U5461 , P2_U5462 , P2_U5463 , P2_U5464 , P2_U5465 , P2_U5466 , P2_U5467 , P2_U5468 , P2_U5469 , P2_U5470;
wire P2_U5471 , P2_U5472 , P2_U5473 , P2_U5474 , P2_U5475 , P2_U5476 , P2_U5477 , P2_U5478 , P2_U5479 , P2_U5480;
wire P2_U5481 , P2_U5482 , P2_U5483 , P2_U5484 , P2_U5485 , P2_U5486 , P2_U5487 , P2_U5488 , P2_U5489 , P2_U5490;
wire P2_U5491 , P2_U5492 , P2_U5493 , P2_U5494 , P2_U5495 , P2_U5496 , P2_U5497 , P2_U5498 , P2_U5499 , P2_U5500;
wire P2_U5501 , P2_U5502 , P2_U5503 , P2_U5504 , P2_U5505 , P2_U5506 , P2_U5507 , P2_U5508 , P2_U5509 , P2_U5510;
wire P2_U5511 , P2_U5512 , P2_U5513 , P2_U5514 , P2_U5515 , P2_U5516 , P2_U5517 , P2_U5518 , P2_U5519 , P2_U5520;
wire P2_U5521 , P2_U5522 , P2_U5523 , P2_U5524 , P2_U5525 , P2_U5526 , P2_U5527 , P2_U5528 , P2_U5529 , P2_U5530;
wire P2_U5531 , P2_U5532 , P2_U5533 , P2_U5534 , P2_U5535 , P2_U5536 , P2_U5537 , P2_U5538 , P2_U5539 , P2_U5540;
wire P2_U5541 , P2_U5542 , P2_U5543 , P2_U5544 , P2_U5545 , P2_U5546 , P2_U5547 , P2_U5548 , P2_U5549 , P2_U5550;
wire P2_U5551 , P2_U5552 , P2_U5553 , P2_U5554 , P2_U5555 , P2_U5556 , P2_U5557 , P2_U5558 , P2_U5559 , P2_U5560;
wire P2_U5561 , P2_U5562 , P2_U5563 , P2_U5564 , P2_U5565 , P2_U5566 , P2_U5567 , P2_U5568 , P2_U5569 , P2_U5570;
wire P2_U5571 , P2_U5572 , P2_U5573 , P2_U5574 , P2_U5575 , P2_U5576 , P2_U5577 , P2_U5578 , P2_U5579 , P2_U5580;
wire P2_U5581 , P2_U5582 , P2_U5583 , P2_U5584 , P2_U5585 , P2_U5586 , P2_U5587 , P2_U5588 , P2_U5589 , P2_U5590;
wire P2_U5591 , P2_U5592 , P2_U5593 , P2_U5594 , P2_U5595 , P2_U5596 , P2_U5597 , P2_U5598 , P2_U5599 , P2_U5600;
wire P2_U5601 , P2_U5602 , P2_U5603 , P2_U5604 , P2_U5605 , P2_U5606 , P2_U5607 , P2_U5608 , P2_U5609 , P2_U5610;
wire P2_U5611 , P2_U5612 , P2_U5613 , P2_U5614 , P2_U5615 , P2_U5616 , P2_U5617 , P2_U5618 , P2_U5619 , P2_U5620;
wire P2_U5621 , P2_U5622 , P2_U5623 , P2_U5624 , P2_U5625 , P2_U5626 , P2_U5627 , P2_U5628 , P2_U5629 , P2_U5630;
wire P2_U5631 , P2_U5632 , P2_U5633 , P2_U5634 , P2_U5635 , P2_U5636 , P2_U5637 , P2_U5638 , P2_U5639 , P2_U5640;
wire P2_U5641 , P2_U5642 , P2_U5643 , P2_U5644 , P2_U5645 , P2_U5646 , P2_U5647 , P2_U5648 , P2_U5649 , P2_U5650;
wire P2_U5651 , P2_U5652 , P2_U5653 , P2_U5654 , P2_U5655 , P2_U5656 , P2_U5657 , P2_U5658 , P2_U5659 , P2_U5660;
wire P2_U5661 , P2_U5662 , P2_U5663 , P2_U5664 , P2_U5665 , P2_U5666 , P2_U5667 , P2_U5668 , P2_U5669 , P2_U5670;
wire P2_U5671 , P2_U5672 , P2_U5673 , P2_U5674 , P2_U5675 , P2_U5676 , P2_U5677 , P2_U5678 , P2_U5679 , P2_U5680;
wire P2_U5681 , P2_U5682 , P2_U5683 , P2_U5684 , P2_U5685 , P2_U5686 , P2_U5687 , P2_U5688 , P2_U5689 , P2_U5690;
wire P2_U5691 , P2_U5692 , P2_U5693 , P2_U5694 , P2_U5695 , P2_U5696 , P2_U5697 , P2_U5698 , P2_U5699 , P2_U5700;
wire P2_U5701 , P2_U5702 , P2_U5703 , P2_U5704 , P2_U5705 , P2_U5706 , P2_U5707 , P2_U5708 , P2_U5709 , P2_U5710;
wire P2_U5711 , P2_U5712 , P2_U5713 , P2_U5714 , P2_U5715 , P2_U5716 , P2_U5717 , P2_U5718 , P2_U5719 , P2_U5720;
wire P2_U5721 , P2_U5722 , P2_U5723 , P2_U5724 , P2_U5725 , P2_U5726 , P2_U5727 , P2_U5728 , P2_U5729 , P2_U5730;
wire P2_U5731 , P2_U5732 , P2_U5733 , P2_U5734 , P2_U5735 , P2_U5736 , P2_U5737 , P2_U5738 , P2_U5739 , P2_U5740;
wire P2_U5741 , P2_U5742 , P2_U5743 , P2_U5744 , P2_U5745 , P2_U5746 , P2_U5747 , P2_U5748 , P2_U5749 , P2_U5750;
wire P2_U5751 , P2_U5752 , P2_U5753 , P2_U5754 , P2_U5755 , P2_U5756 , P2_U5757 , P2_U5758 , P2_U5759 , P2_U5760;
wire P2_U5761 , P2_U5762 , P2_U5763 , P2_U5764 , P2_U5765 , P2_U5766 , P2_U5767 , P2_U5768 , P2_U5769 , P2_U5770;
wire P2_U5771 , P2_U5772 , P2_U5773 , P2_U5774 , P2_U5775 , P2_U5776 , P2_U5777 , P2_U5778 , P2_U5779 , P2_U5780;
wire P2_U5781 , P2_U5782 , P2_U5783 , P2_U5784 , P2_U5785 , P2_U5786 , P2_U5787 , P2_U5788 , P2_U5789 , P2_U5790;
wire P2_U5791 , P2_U5792 , P2_U5793 , P2_U5794 , P2_U5795 , P2_U5796 , P2_U5797 , P2_U5798 , P2_U5799 , P2_U5800;
wire P2_U5801 , P2_U5802 , P2_U5803 , P2_U5804 , P2_U5805 , P2_U5806 , P2_U5807 , P2_U5808 , P2_U5809 , P2_U5810;
wire P2_U5811 , P2_U5812 , P2_U5813 , P2_U5814 , P2_U5815 , P2_U5816 , P2_U5817 , P2_U5818 , P2_U5819 , P2_U5820;
wire P2_U5821 , P2_U5822 , P2_U5823 , P2_U5824 , P2_U5825 , P2_U5826 , P2_U5827 , P2_U5828 , P2_U5829 , P2_U5830;
wire P2_U5831 , P2_U5832 , P2_U5833 , P2_U5834 , P2_U5835 , P2_U5836 , P2_U5837 , P2_U5838 , P2_U5839 , P2_U5840;
wire P2_U5841 , P2_U5842 , P2_U5843 , P2_U5844 , P2_U5845 , P2_U5846 , P2_U5847 , P2_U5848 , P2_U5849 , P2_U5850;
wire P2_U5851 , P2_U5852 , P2_U5853 , P2_U5854 , P2_U5855 , P2_U5856 , P2_U5857 , P2_U5858 , P2_U5859 , P2_U5860;
wire P2_U5861 , P2_U5862 , P2_U5863 , P2_U5864 , P2_U5865 , P2_U5866 , P2_U5867 , P2_U5868 , P2_U5869 , P2_U5870;
wire P2_U5871 , P2_U5872 , P2_U5873 , P2_U5874 , P2_U5875 , P2_U5876 , P2_U5877 , P2_U5878 , P2_U5879 , P2_U5880;
wire P2_U5881 , P2_U5882 , P2_U5883 , P2_U5884 , P2_U5885 , P2_U5886 , P2_U5887 , P2_U5888 , P2_U5889 , P2_U5890;
wire P2_U5891 , P2_U5892 , P2_U5893 , P2_U5894 , P2_U5895 , P2_U5896 , P2_U5897 , P2_U5898 , P2_U5899 , P2_U5900;
wire P2_U5901 , P2_U5902 , P2_U5903 , P2_U5904 , P2_U5905 , P2_U5906 , P2_U5907 , P2_U5908 , P2_U5909 , P2_U5910;
wire P2_U5911 , P2_U5912 , P2_U5913 , P2_U5914 , P2_U5915 , P2_U5916 , P2_U5917 , P2_U5918 , P2_U5919 , P2_U5920;
wire P2_U5921 , P2_U5922 , P2_U5923 , P2_U5924 , P2_U5925 , P2_U5926 , P2_U5927 , P2_U5928 , P2_U5929 , P2_U5930;
wire P2_U5931 , P2_U5932 , P2_U5933 , P2_U5934 , P2_U5935 , P2_U5936 , P2_U5937 , P2_U5938 , P2_U5939 , P2_U5940;
wire P2_U5941 , P2_U5942 , P2_U5943 , P2_U5944 , P2_U5945 , P2_U5946 , P2_U5947 , P2_U5948 , P2_U5949 , P2_U5950;
wire P2_U5951 , P2_U5952 , P2_U5953 , P2_U5954 , P2_U5955 , P2_U5956 , P2_U5957 , P2_U5958 , P2_U5959 , P2_U5960;
wire P2_U5961 , P2_U5962 , P2_U5963 , P2_U5964 , P2_U5965 , P2_U5966 , P2_U5967 , P2_U5968 , P2_U5969 , P2_U5970;
wire P2_U5971 , P2_U5972 , P2_U5973 , P2_U5974 , P2_U5975 , P2_U5976 , P2_U5977 , P2_U5978 , P2_U5979 , P2_U5980;
wire P2_U5981 , P2_U5982 , P2_U5983 , P2_U5984 , P2_U5985 , P2_U5986 , P2_U5987 , P2_U5988 , P2_U5989 , P2_U5990;
wire P2_U5991 , P2_U5992 , P2_U5993 , P2_U5994 , P2_U5995 , P2_U5996 , P2_U5997 , P2_U5998 , P2_U5999 , P2_U6000;
wire P2_U6001 , P2_U6002 , P2_U6003 , P2_U6004 , P2_U6005 , P2_U6006 , P2_U6007 , P2_U6008 , P2_U6009 , P2_U6010;
wire P2_U6011 , P2_U6012 , P2_U6013 , P2_U6014 , P2_U6015 , P2_U6016 , P2_U6017 , P2_U6018 , P2_U6019 , P2_U6020;
wire P2_U6021 , P2_U6022 , P2_U6023 , P2_U6024 , P2_U6025 , P2_U6026 , P2_U6027 , P2_U6028 , P2_U6029 , P2_U6030;
wire P2_U6031 , P2_U6032 , P2_U6033 , P2_U6034 , P2_U6035 , P2_U6036 , P2_U6037 , P2_U6038 , P2_U6039 , P2_U6040;
wire P2_U6041 , P2_U6042 , P2_U6043 , P2_U6044 , P2_U6045 , P2_U6046 , P2_U6047 , P2_U6048 , P2_U6049 , P2_U6050;
wire P2_U6051 , P2_U6052 , P2_U6053 , P2_U6054 , P2_U6055 , P2_U6056 , P2_U6057 , P2_U6058 , P2_U6059 , P2_U6060;
wire P2_U6061 , P2_U6062 , P2_U6063 , P2_U6064 , P2_U6065 , P2_U6066 , P2_U6067 , P2_U6068 , P2_U6069 , P2_U6070;
wire P2_U6071 , P2_U6072 , P2_U6073 , P2_U6074 , P2_U6075 , P2_U6076 , P2_U6077 , P2_U6078 , P2_U6079 , P2_U6080;
wire P2_U6081 , P2_U6082 , P2_U6083 , P2_U6084 , P2_U6085 , P2_U6086 , P2_U6087 , P2_U6088 , P2_U6089 , P2_U6090;
wire P2_U6091 , P2_U6092 , P2_U6093 , P2_U6094 , P2_U6095 , P2_U6096 , P2_U6097 , P2_U6098 , P2_U6099 , P2_U6100;
wire P2_U6101 , P2_U6102 , P2_U6103 , P2_U6104 , P2_U6105 , P2_U6106 , P2_U6107 , P2_U6108 , P2_U6109 , P2_U6110;
wire P2_U6111 , P2_U6112 , P2_U6113 , P2_U6114 , P2_U6115 , P2_U6116 , P2_U6117 , P2_U6118 , P2_U6119 , P2_U6120;
wire P2_U6121 , P2_U6122 , P2_U6123 , P2_U6124 , P2_U6125 , P2_U6126 , P2_U6127 , P2_U6128 , P2_U6129 , P2_U6130;
wire P2_U6131 , P2_U6132 , P2_U6133 , P2_U6134 , P2_U6135 , P2_U6136 , P2_U6137 , P2_U6138 , P2_U6139 , P2_U6140;
wire P2_U6141 , P2_U6142 , P2_U6143 , P2_U6144 , P2_U6145 , P2_U6146 , P2_U6147 , P2_U6148 , P2_U6149 , P2_U6150;
wire P2_U6151 , P2_U6152 , P2_U6153 , P2_U6154 , P2_U6155 , P2_U6156 , P2_U6157 , P2_U6158 , P2_U6159 , P2_U6160;
wire P2_U6161 , P2_U6162 , P2_U6163 , P2_U6164 , P2_U6165 , P2_U6166 , P2_U6167 , P2_U6168 , P2_U6169 , P2_U6170;
wire P2_U6171 , P2_U6172 , P2_U6173 , P2_U6174 , P2_U6175 , P2_U6176 , P2_U6177 , P2_U6178 , P2_U6179 , P2_U6180;
wire P2_U6181 , P2_U6182 , P2_U6183 , P2_U6184 , P2_U6185 , P2_U6186 , P2_U6187 , P2_U6188 , P2_U6189 , P2_U6190;
wire P2_U6191 , P2_U6192 , P2_U6193 , P2_U6194 , P2_U6195 , P2_U6196 , P2_U6197 , P2_U6198 , P2_U6199 , P2_U6200;
wire P2_U6201 , P2_U6202 , P2_U6203 , P2_U6204 , P2_U6205 , P2_U6206 , P2_U6207 , P2_U6208 , P2_U6209 , P2_U6210;
wire P2_U6211 , P2_U6212 , P2_U6213 , P2_U6214 , P2_U6215 , P2_U6216 , P2_U6217 , P2_U6218 , P2_U6219 , P2_U6220;
wire P2_U6221 , P2_U6222 , P2_U6223 , P2_U6224 , P2_U6225 , P2_U6226 , P2_U6227 , P2_U6228 , P2_U6229 , P2_U6230;
wire P2_U6231 , P2_U6232 , P2_U6233 , P2_U6234 , P2_U6235 , P2_U6236 , P2_U6237 , P2_U6238 , P2_U6239 , P2_U6240;
wire P2_U6241 , P2_U6242 , P2_U6243 , P2_U6244 , P2_U6245 , P2_U6246 , P2_U6247 , P2_U6248 , P2_U6249 , P2_U6250;
wire P2_U6251 , P2_U6252 , P2_U6253 , P2_U6254 , P2_U6255 , P2_U6256 , P2_U6257 , P2_U6258 , P2_U6259 , P2_U6260;
wire P2_U6261 , P2_U6262 , P2_U6263 , P2_U6264 , P2_U6265 , P2_U6266 , P2_U6267 , P2_U6268 , P2_U6269 , P2_U6270;
wire P2_U6271 , P2_U6272 , P2_U6273 , P2_U6274 , P2_U6275 , P2_U6276 , P2_U6277 , P2_U6278 , P2_U6279 , P2_U6280;
wire P2_U6281 , P2_U6282 , P2_U6283 , P2_U6284 , P2_U6285 , P2_U6286 , P2_U6287 , P2_U6288 , P2_U6289 , P2_U6290;
wire P2_U6291 , P2_U6292 , P2_U6293 , P2_U6294 , P2_U6295 , P2_U6296 , P2_U6297 , P2_U6298 , P2_U6299 , P2_U6300;
wire P2_U6301 , P2_U6302 , P2_U6303 , P2_U6304 , P2_U6305 , P2_U6306 , P2_U6307 , P2_U6308 , P2_U6309 , P2_U6310;
wire P2_U6311 , P2_U6312 , P2_U6313 , P2_U6314 , P2_U6315 , P2_U6316 , P2_U6317 , P2_U6318 , P2_U6319 , P2_U6320;
wire P2_U6321 , P2_U6322 , P2_U6323 , P2_U6324 , P2_U6325 , P2_U6326 , P2_U6327 , P2_U6328 , P2_U6329 , P2_U6330;
wire P2_U6331 , P2_U6332 , P2_U6333 , P2_U6334 , P2_U6335 , P2_U6336 , P2_U6337 , P2_U6338 , P2_U6339 , P2_U6340;
wire P2_U6341 , P2_U6342 , P2_U6343 , P2_U6344 , P2_U6345 , P2_U6346 , P2_U6347 , P2_U6348 , P2_U6349 , P2_U6350;
wire P2_U6351 , P2_U6352 , P2_U6353 , P2_U6354 , P2_U6355 , P2_U6356 , P2_U6357 , P2_U6358 , P2_U6359 , P2_U6360;
wire P2_U6361 , P2_U6362 , P2_U6363 , P2_U6364 , P2_U6365 , P2_U6366 , P2_U6367 , P2_U6368 , P2_U6369 , P2_U6370;
wire P2_U6371 , P2_U6372 , P2_U6373 , P2_U6374 , P2_U6375 , P2_U6376 , P2_U6377 , P2_U6378 , P2_U6379 , P2_U6380;
wire P2_U6381 , P2_U6382 , P2_U6383 , P2_U6384 , P2_U6385 , P2_U6386 , P2_U6387 , P2_U6388 , P2_U6389 , P2_U6390;
wire P2_U6391 , P2_U6392 , P2_U6393 , P2_U6394 , P2_U6395 , P2_U6396 , P2_U6397 , P2_U6398 , P2_U6399 , P2_U6400;
wire P2_U6401 , P2_U6402 , P2_U6403 , P2_U6404 , P2_U6405 , P2_U6406 , P2_U6407 , P2_U6408 , P2_U6409 , P2_U6410;
wire P2_U6411 , P2_U6412 , P2_U6413 , P2_U6414 , P2_U6415 , P2_U6416 , P2_U6417 , P2_U6418 , P2_U6419 , P2_U6420;
wire P2_U6421 , P2_U6422 , P2_U6423 , P2_U6424 , P2_U6425 , P2_U6426 , P2_U6427 , P2_U6428 , P2_U6429 , P2_U6430;
wire P2_U6431 , P2_U6432 , P2_U6433 , P2_U6434 , P2_U6435 , P2_U6436 , P2_U6437 , P2_U6438 , P2_U6439 , P2_U6440;
wire P2_U6441 , P2_U6442 , P2_U6443 , P2_U6444 , P2_U6445 , P2_U6446 , P2_U6447 , P2_U6448 , P2_U6449 , P2_U6450;
wire P2_U6451 , P2_U6452 , P2_U6453 , P2_U6454 , P2_U6455 , P2_U6456 , P2_U6457 , P2_U6458 , P2_U6459 , P2_U6460;
wire P2_U6461 , P2_U6462 , P2_U6463 , P2_U6464 , P2_U6465 , P2_U6466 , P2_U6467 , P2_U6468 , P2_U6469 , P2_U6470;
wire P2_U6471 , P2_U6472 , P2_U6473 , P2_U6474 , P2_U6475 , P2_U6476 , P2_U6477 , P2_U6478 , P2_U6479 , P2_U6480;
wire P2_U6481 , P2_U6482 , P2_U6483 , P2_U6484 , P2_U6485 , P2_U6486 , P2_U6487 , P2_U6488 , P2_U6489 , P2_U6490;
wire P2_U6491 , P2_U6492 , P2_U6493 , P2_U6494 , P2_U6495 , P2_U6496 , P2_U6497 , P2_U6498 , P2_U6499 , P2_U6500;
wire P2_U6501 , P2_U6502 , P2_U6503 , P2_U6504 , P2_U6505 , P2_U6506 , P2_U6507 , P2_U6508 , P2_U6509 , P2_U6510;
wire P2_U6511 , P2_U6512 , P2_U6513 , P2_U6514 , P2_U6515 , P2_U6516 , P2_U6517 , P2_U6518 , P2_U6519 , P2_U6520;
wire P2_U6521 , P2_U6522 , P2_U6523 , P2_U6524 , P2_U6525 , P2_U6526 , P2_U6527 , P2_U6528 , P2_U6529 , P2_U6530;
wire P2_U6531 , P2_U6532 , P2_U6533 , P2_U6534 , P2_U6535 , P2_U6536 , P2_U6537 , P2_U6538 , P2_U6539 , P2_U6540;
wire P2_U6541 , P2_U6542 , P2_U6543 , P2_U6544 , P2_U6545 , P2_U6546 , P2_U6547 , P2_U6548 , P2_U6549 , P2_U6550;
wire P2_U6551 , P2_U6552 , P2_U6553 , P2_U6554 , P2_U6555 , P2_U6556 , P2_U6557 , P2_U6558 , P2_U6559 , P2_U6560;
wire P2_U6561 , P2_U6562 , P2_U6563 , P2_U6564 , P2_U6565 , P2_U6566 , P2_U6567 , P2_U6568 , P2_U6569 , P2_U6570;
wire P2_U6571 , P2_U6572 , P2_U6573 , P2_U6574 , P2_U6575 , P2_U6576 , P2_U6577 , P2_U6578 , P2_U6579 , P2_U6580;
wire P2_U6581 , P2_U6582 , P2_U6583 , P2_U6584 , P2_U6585 , P2_U6586 , P2_U6587 , P2_U6588 , P2_U6589 , P2_U6590;
wire P2_U6591 , P2_U6592 , P2_U6593 , P2_U6594 , P2_U6595 , P2_U6596 , P2_U6597 , P2_U6598 , P2_U6599 , P2_U6600;
wire P2_U6601 , P2_U6602 , P2_U6603 , P2_U6604 , P2_U6605 , P2_U6606 , P2_U6607 , P2_U6608 , P2_U6609 , P2_U6610;
wire P2_U6611 , P2_U6612 , P2_U6613 , P2_U6614 , P2_U6615 , P2_U6616 , P2_U6617 , P2_U6618 , P2_U6619 , P2_U6620;
wire P2_U6621 , P2_U6622 , P2_U6623 , P2_U6624 , P2_U6625 , P2_U6626 , P2_U6627 , P2_U6628 , P2_U6629 , P2_U6630;
wire P2_U6631 , P2_U6632 , P2_U6633 , P2_U6634 , P2_U6635 , P2_U6636 , P2_U6637 , P2_U6638 , P2_U6639 , P2_U6640;
wire P2_U6641 , P2_U6642 , P2_U6643 , P2_U6644 , P2_U6645 , P2_U6646 , P2_U6647 , P2_U6648 , P2_U6649 , P2_U6650;
wire P2_U6651 , P2_U6652 , P2_U6653 , P2_U6654 , P2_U6655 , P2_U6656 , P2_U6657 , P2_U6658 , P2_U6659 , P2_U6660;
wire P2_U6661 , P2_U6662 , P2_U6663 , P2_U6664 , P2_U6665 , P2_U6666 , P2_U6667 , P2_U6668 , P2_U6669 , P2_U6670;
wire P2_U6671 , P2_U6672 , P2_U6673 , P2_U6674 , P2_U6675 , P2_U6676 , P2_U6677 , P2_U6678 , P2_U6679 , P2_U6680;
wire P2_U6681 , P2_U6682 , P2_U6683 , P2_U6684 , P2_U6685 , P2_U6686 , P2_U6687 , P2_U6688 , P2_U6689 , P2_U6690;
wire P2_U6691 , P2_U6692 , P2_U6693 , P2_U6694 , P2_U6695 , P2_U6696 , P2_U6697 , P2_U6698 , P2_U6699 , P2_U6700;
wire P2_U6701 , P2_U6702 , P2_U6703 , P2_U6704 , P2_U6705 , P2_U6706 , P2_U6707 , P2_U6708 , P2_U6709 , P2_U6710;
wire P2_U6711 , P2_U6712 , P2_U6713 , P2_U6714 , P2_U6715 , P2_U6716 , P2_U6717 , P2_U6718 , P2_U6719 , P2_U6720;
wire P2_U6721 , P2_U6722 , P2_U6723 , P2_U6724 , P2_U6725 , P2_U6726 , P2_U6727 , P2_U6728 , P2_U6729 , P2_U6730;
wire P2_U6731 , P2_U6732 , P2_U6733 , P2_U6734 , P2_U6735 , P2_U6736 , P2_U6737 , P2_U6738 , P2_U6739 , P2_U6740;
wire P2_U6741 , P2_U6742 , P2_U6743 , P2_U6744 , P2_U6745 , P2_U6746 , P2_U6747 , P2_U6748 , P2_U6749 , P2_U6750;
wire P2_U6751 , P2_U6752 , P2_U6753 , P2_U6754 , P2_U6755 , P2_U6756 , P2_U6757 , P2_U6758 , P2_U6759 , P2_U6760;
wire P2_U6761 , P2_U6762 , P2_U6763 , P2_U6764 , P2_U6765 , P2_U6766 , P2_U6767 , P2_U6768 , P2_U6769 , P2_U6770;
wire P2_U6771 , P2_U6772 , P2_U6773 , P2_U6774 , P2_U6775 , P2_U6776 , P2_U6777 , P2_U6778 , P2_U6779 , P2_U6780;
wire P2_U6781 , P2_U6782 , P2_U6783 , P2_U6784 , P2_U6785 , P2_U6786 , P2_U6787 , P2_U6788 , P2_U6789 , P2_U6790;
wire P2_U6791 , P2_U6792 , P2_U6793 , P2_U6794 , P2_U6795 , P2_U6796 , P2_U6797 , P2_U6798 , P2_U6799 , P2_U6800;
wire P2_U6801 , P2_U6802 , P2_U6803 , P2_U6804 , P2_U6805 , P2_U6806 , P2_U6807 , P2_U6808 , P2_U6809 , P2_U6810;
wire P2_U6811 , P2_U6812 , P2_U6813 , P2_U6814 , P2_U6815 , P2_U6816 , P2_U6817 , P2_U6818 , P2_U6819 , P2_U6820;
wire P2_U6821 , P2_U6822 , P2_U6823 , P2_U6824 , P2_U6825 , P2_U6826 , P2_U6827 , P2_U6828 , P2_U6829 , P2_U6830;
wire P2_U6831 , P2_U6832 , P2_U6833 , P2_U6834 , P2_U6835 , P2_U6836 , P2_U6837 , P2_U6838 , P2_U6839 , P2_U6840;
wire P2_U6841 , P2_U6842 , P2_U6843 , P2_U6844 , P2_U6845 , P2_U6846 , P2_U6847 , P2_U6848 , P2_U6849 , P2_U6850;
wire P2_U6851 , P2_U6852 , P2_U6853 , P2_U6854 , P2_U6855 , P2_U6856 , P2_U6857 , P2_U6858 , P2_U6859 , P2_U6860;
wire P2_U6861 , P2_U6862 , P2_U6863 , P2_U6864 , P2_U6865 , P2_U6866 , P2_U6867 , P2_U6868 , P2_U6869 , P2_U6870;
wire P2_U6871 , P2_U6872 , P2_U6873 , P2_U6874 , P2_U6875 , P2_U6876 , P2_U6877 , P2_U6878 , P2_U6879 , P2_U6880;
wire P2_U6881 , P2_U6882 , P2_U6883 , P2_U6884 , P2_U6885 , P2_U6886 , P2_U6887 , P2_U6888 , P2_U6889 , P2_U6890;
wire P2_U6891 , P2_U6892 , P2_U6893 , P2_U6894 , P2_U6895 , P2_U6896 , P2_U6897 , P2_U6898 , P2_U6899 , P2_U6900;
wire P2_U6901 , P2_U6902 , P2_U6903 , P2_U6904 , P2_U6905 , P2_U6906 , P2_U6907 , P2_U6908 , P2_U6909 , P2_U6910;
wire P2_U6911 , P2_U6912 , P2_U6913 , P2_U6914 , P2_U6915 , P2_U6916 , P2_U6917 , P2_U6918 , P2_U6919 , P2_U6920;
wire P2_U6921 , P2_U6922 , P2_U6923 , P2_U6924 , P2_U6925 , P2_U6926 , P2_U6927 , P2_U6928 , P2_U6929 , P2_U6930;
wire P2_U6931 , P2_U6932 , P2_U6933 , P2_U6934 , P2_U6935 , P2_U6936 , P2_U6937 , P2_U6938 , P2_U6939 , P2_U6940;
wire P2_U6941 , P2_U6942 , P2_U6943 , P2_U6944 , P2_U6945 , P2_U6946 , P2_U6947 , P2_U6948 , P2_U6949 , P2_U6950;
wire P2_U6951 , P2_U6952 , P2_U6953 , P2_U6954 , P2_U6955 , P2_U6956 , P2_U6957 , P2_U6958 , P2_U6959 , P2_U6960;
wire P2_U6961 , P2_U6962 , P2_U6963 , P2_U6964 , P2_U6965 , P2_U6966 , P2_U6967 , P2_U6968 , P2_U6969 , P2_U6970;
wire P2_U6971 , P2_U6972 , P2_U6973 , P2_U6974 , P2_U6975 , P2_U6976 , P2_U6977 , P2_U6978 , P2_U6979 , P2_U6980;
wire P2_U6981 , P2_U6982 , P2_U6983 , P2_U6984 , P2_U6985 , P2_U6986 , P2_U6987 , P2_U6988 , P2_U6989 , P2_U6990;
wire P2_U6991 , P2_U6992 , P2_U6993 , P2_U6994 , P2_U6995 , P2_U6996 , P2_U6997 , P2_U6998 , P2_U6999 , P2_U7000;
wire P2_U7001 , P2_U7002 , P2_U7003 , P2_U7004 , P2_U7005 , P2_U7006 , P2_U7007 , P2_U7008 , P2_U7009 , P2_U7010;
wire P2_U7011 , P2_U7012 , P2_U7013 , P2_U7014 , P2_U7015 , P2_U7016 , P2_U7017 , P2_U7018 , P2_U7019 , P2_U7020;
wire P2_U7021 , P2_U7022 , P2_U7023 , P2_U7024 , P2_U7025 , P2_U7026 , P2_U7027 , P2_U7028 , P2_U7029 , P2_U7030;
wire P2_U7031 , P2_U7032 , P2_U7033 , P2_U7034 , P2_U7035 , P2_U7036 , P2_U7037 , P2_U7038 , P2_U7039 , P2_U7040;
wire P2_U7041 , P2_U7042 , P2_U7043 , P2_U7044 , P2_U7045 , P2_U7046 , P2_U7047 , P2_U7048 , P2_U7049 , P2_U7050;
wire P2_U7051 , P2_U7052 , P2_U7053 , P2_U7054 , P2_U7055 , P2_U7056 , P2_U7057 , P2_U7058 , P2_U7059 , P2_U7060;
wire P2_U7061 , P2_U7062 , P2_U7063 , P2_U7064 , P2_U7065 , P2_U7066 , P2_U7067 , P2_U7068 , P2_U7069 , P2_U7070;
wire P2_U7071 , P2_U7072 , P2_U7073 , P2_U7074 , P2_U7075 , P2_U7076 , P2_U7077 , P2_U7078 , P2_U7079 , P2_U7080;
wire P2_U7081 , P2_U7082 , P2_U7083 , P2_U7084 , P2_U7085 , P2_U7086 , P2_U7087 , P2_U7088 , P2_U7089 , P2_U7090;
wire P2_U7091 , P2_U7092 , P2_U7093 , P2_U7094 , P2_U7095 , P2_U7096 , P2_U7097 , P2_U7098 , P2_U7099 , P2_U7100;
wire P2_U7101 , P2_U7102 , P2_U7103 , P2_U7104 , P2_U7105 , P2_U7106 , P2_U7107 , P2_U7108 , P2_U7109 , P2_U7110;
wire P2_U7111 , P2_U7112 , P2_U7113 , P2_U7114 , P2_U7115 , P2_U7116 , P2_U7117 , P2_U7118 , P2_U7119 , P2_U7120;
wire P2_U7121 , P2_U7122 , P2_U7123 , P2_U7124 , P2_U7125 , P2_U7126 , P2_U7127 , P2_U7128 , P2_U7129 , P2_U7130;
wire P2_U7131 , P2_U7132 , P2_U7133 , P2_U7134 , P2_U7135 , P2_U7136 , P2_U7137 , P2_U7138 , P2_U7139 , P2_U7140;
wire P2_U7141 , P2_U7142 , P2_U7143 , P2_U7144 , P2_U7145 , P2_U7146 , P2_U7147 , P2_U7148 , P2_U7149 , P2_U7150;
wire P2_U7151 , P2_U7152 , P2_U7153 , P2_U7154 , P2_U7155 , P2_U7156 , P2_U7157 , P2_U7158 , P2_U7159 , P2_U7160;
wire P2_U7161 , P2_U7162 , P2_U7163 , P2_U7164 , P2_U7165 , P2_U7166 , P2_U7167 , P2_U7168 , P2_U7169 , P2_U7170;
wire P2_U7171 , P2_U7172 , P2_U7173 , P2_U7174 , P2_U7175 , P2_U7176 , P2_U7177 , P2_U7178 , P2_U7179 , P2_U7180;
wire P2_U7181 , P2_U7182 , P2_U7183 , P2_U7184 , P2_U7185 , P2_U7186 , P2_U7187 , P2_U7188 , P2_U7189 , P2_U7190;
wire P2_U7191 , P2_U7192 , P2_U7193 , P2_U7194 , P2_U7195 , P2_U7196 , P2_U7197 , P2_U7198 , P2_U7199 , P2_U7200;
wire P2_U7201 , P2_U7202 , P2_U7203 , P2_U7204 , P2_U7205 , P2_U7206 , P2_U7207 , P2_U7208 , P2_U7209 , P2_U7210;
wire P2_U7211 , P2_U7212 , P2_U7213 , P2_U7214 , P2_U7215 , P2_U7216 , P2_U7217 , P2_U7218 , P2_U7219 , P2_U7220;
wire P2_U7221 , P2_U7222 , P2_U7223 , P2_U7224 , P2_U7225 , P2_U7226 , P2_U7227 , P2_U7228 , P2_U7229 , P2_U7230;
wire P2_U7231 , P2_U7232 , P2_U7233 , P2_U7234 , P2_U7235 , P2_U7236 , P2_U7237 , P2_U7238 , P2_U7239 , P2_U7240;
wire P2_U7241 , P2_U7242 , P2_U7243 , P2_U7244 , P2_U7245 , P2_U7246 , P2_U7247 , P2_U7248 , P2_U7249 , P2_U7250;
wire P2_U7251 , P2_U7252 , P2_U7253 , P2_U7254 , P2_U7255 , P2_U7256 , P2_U7257 , P2_U7258 , P2_U7259 , P2_U7260;
wire P2_U7261 , P2_U7262 , P2_U7263 , P2_U7264 , P2_U7265 , P2_U7266 , P2_U7267 , P2_U7268 , P2_U7269 , P2_U7270;
wire P2_U7271 , P2_U7272 , P2_U7273 , P2_U7274 , P2_U7275 , P2_U7276 , P2_U7277 , P2_U7278 , P2_U7279 , P2_U7280;
wire P2_U7281 , P2_U7282 , P2_U7283 , P2_U7284 , P2_U7285 , P2_U7286 , P2_U7287 , P2_U7288 , P2_U7289 , P2_U7290;
wire P2_U7291 , P2_U7292 , P2_U7293 , P2_U7294 , P2_U7295 , P2_U7296 , P2_U7297 , P2_U7298 , P2_U7299 , P2_U7300;
wire P2_U7301 , P2_U7302 , P2_U7303 , P2_U7304 , P2_U7305 , P2_U7306 , P2_U7307 , P2_U7308 , P2_U7309 , P2_U7310;
wire P2_U7311 , P2_U7312 , P2_U7313 , P2_U7314 , P2_U7315 , P2_U7316 , P2_U7317 , P2_U7318 , P2_U7319 , P2_U7320;
wire P2_U7321 , P2_U7322 , P2_U7323 , P2_U7324 , P2_U7325 , P2_U7326 , P2_U7327 , P2_U7328 , P2_U7329 , P2_U7330;
wire P2_U7331 , P2_U7332 , P2_U7333 , P2_U7334 , P2_U7335 , P2_U7336 , P2_U7337 , P2_U7338 , P2_U7339 , P2_U7340;
wire P2_U7341 , P2_U7342 , P2_U7343 , P2_U7344 , P2_U7345 , P2_U7346 , P2_U7347 , P2_U7348 , P2_U7349 , P2_U7350;
wire P2_U7351 , P2_U7352 , P2_U7353 , P2_U7354 , P2_U7355 , P2_U7356 , P2_U7357 , P2_U7358 , P2_U7359 , P2_U7360;
wire P2_U7361 , P2_U7362 , P2_U7363 , P2_U7364 , P2_U7365 , P2_U7366 , P2_U7367 , P2_U7368 , P2_U7369 , P2_U7370;
wire P2_U7371 , P2_U7372 , P2_U7373 , P2_U7374 , P2_U7375 , P2_U7376 , P2_U7377 , P2_U7378 , P2_U7379 , P2_U7380;
wire P2_U7381 , P2_U7382 , P2_U7383 , P2_U7384 , P2_U7385 , P2_U7386 , P2_U7387 , P2_U7388 , P2_U7389 , P2_U7390;
wire P2_U7391 , P2_U7392 , P2_U7393 , P2_U7394 , P2_U7395 , P2_U7396 , P2_U7397 , P2_U7398 , P2_U7399 , P2_U7400;
wire P2_U7401 , P2_U7402 , P2_U7403 , P2_U7404 , P2_U7405 , P2_U7406 , P2_U7407 , P2_U7408 , P2_U7409 , P2_U7410;
wire P2_U7411 , P2_U7412 , P2_U7413 , P2_U7414 , P2_U7415 , P2_U7416 , P2_U7417 , P2_U7418 , P2_U7419 , P2_U7420;
wire P2_U7421 , P2_U7422 , P2_U7423 , P2_U7424 , P2_U7425 , P2_U7426 , P2_U7427 , P2_U7428 , P2_U7429 , P2_U7430;
wire P2_U7431 , P2_U7432 , P2_U7433 , P2_U7434 , P2_U7435 , P2_U7436 , P2_U7437 , P2_U7438 , P2_U7439 , P2_U7440;
wire P2_U7441 , P2_U7442 , P2_U7443 , P2_U7444 , P2_U7445 , P2_U7446 , P2_U7447 , P2_U7448 , P2_U7449 , P2_U7450;
wire P2_U7451 , P2_U7452 , P2_U7453 , P2_U7454 , P2_U7455 , P2_U7456 , P2_U7457 , P2_U7458 , P2_U7459 , P2_U7460;
wire P2_U7461 , P2_U7462 , P2_U7463 , P2_U7464 , P2_U7465 , P2_U7466 , P2_U7467 , P2_U7468 , P2_U7469 , P2_U7470;
wire P2_U7471 , P2_U7472 , P2_U7473 , P2_U7474 , P2_U7475 , P2_U7476 , P2_U7477 , P2_U7478 , P2_U7479 , P2_U7480;
wire P2_U7481 , P2_U7482 , P2_U7483 , P2_U7484 , P2_U7485 , P2_U7486 , P2_U7487 , P2_U7488 , P2_U7489 , P2_U7490;
wire P2_U7491 , P2_U7492 , P2_U7493 , P2_U7494 , P2_U7495 , P2_U7496 , P2_U7497 , P2_U7498 , P2_U7499 , P2_U7500;
wire P2_U7501 , P2_U7502 , P2_U7503 , P2_U7504 , P2_U7505 , P2_U7506 , P2_U7507 , P2_U7508 , P2_U7509 , P2_U7510;
wire P2_U7511 , P2_U7512 , P2_U7513 , P2_U7514 , P2_U7515 , P2_U7516 , P2_U7517 , P2_U7518 , P2_U7519 , P2_U7520;
wire P2_U7521 , P2_U7522 , P2_U7523 , P2_U7524 , P2_U7525 , P2_U7526 , P2_U7527 , P2_U7528 , P2_U7529 , P2_U7530;
wire P2_U7531 , P2_U7532 , P2_U7533 , P2_U7534 , P2_U7535 , P2_U7536 , P2_U7537 , P2_U7538 , P2_U7539 , P2_U7540;
wire P2_U7541 , P2_U7542 , P2_U7543 , P2_U7544 , P2_U7545 , P2_U7546 , P2_U7547 , P2_U7548 , P2_U7549 , P2_U7550;
wire P2_U7551 , P2_U7552 , P2_U7553 , P2_U7554 , P2_U7555 , P2_U7556 , P2_U7557 , P2_U7558 , P2_U7559 , P2_U7560;
wire P2_U7561 , P2_U7562 , P2_U7563 , P2_U7564 , P2_U7565 , P2_U7566 , P2_U7567 , P2_U7568 , P2_U7569 , P2_U7570;
wire P2_U7571 , P2_U7572 , P2_U7573 , P2_U7574 , P2_U7575 , P2_U7576 , P2_U7577 , P2_U7578 , P2_U7579 , P2_U7580;
wire P2_U7581 , P2_U7582 , P2_U7583 , P2_U7584 , P2_U7585 , P2_U7586 , P2_U7587 , P2_U7588 , P2_U7589 , P2_U7590;
wire P2_U7591 , P2_U7592 , P2_U7593 , P2_U7594 , P2_U7595 , P2_U7596 , P2_U7597 , P2_U7598 , P2_U7599 , P2_U7600;
wire P2_U7601 , P2_U7602 , P2_U7603 , P2_U7604 , P2_U7605 , P2_U7606 , P2_U7607 , P2_U7608 , P2_U7609 , P2_U7610;
wire P2_U7611 , P2_U7612 , P2_U7613 , P2_U7614 , P2_U7615 , P2_U7616 , P2_U7617 , P2_U7618 , P2_U7619 , P2_U7620;
wire P2_U7621 , P2_U7622 , P2_U7623 , P2_U7624 , P2_U7625 , P2_U7626 , P2_U7627 , P2_U7628 , P2_U7629 , P2_U7630;
wire P2_U7631 , P2_U7632 , P2_U7633 , P2_U7634 , P2_U7635 , P2_U7636 , P2_U7637 , P2_U7638 , P2_U7639 , P2_U7640;
wire P2_U7641 , P2_U7642 , P2_U7643 , P2_U7644 , P2_U7645 , P2_U7646 , P2_U7647 , P2_U7648 , P2_U7649 , P2_U7650;
wire P2_U7651 , P2_U7652 , P2_U7653 , P2_U7654 , P2_U7655 , P2_U7656 , P2_U7657 , P2_U7658 , P2_U7659 , P2_U7660;
wire P2_U7661 , P2_U7662 , P2_U7663 , P2_U7664 , P2_U7665 , P2_U7666 , P2_U7667 , P2_U7668 , P2_U7669 , P2_U7670;
wire P2_U7671 , P2_U7672 , P2_U7673 , P2_U7674 , P2_U7675 , P2_U7676 , P2_U7677 , P2_U7678 , P2_U7679 , P2_U7680;
wire P2_U7681 , P2_U7682 , P2_U7683 , P2_U7684 , P2_U7685 , P2_U7686 , P2_U7687 , P2_U7688 , P2_U7689 , P2_U7690;
wire P2_U7691 , P2_U7692 , P2_U7693 , P2_U7694 , P2_U7695 , P2_U7696 , P2_U7697 , P2_U7698 , P2_U7699 , P2_U7700;
wire P2_U7701 , P2_U7702 , P2_U7703 , P2_U7704 , P2_U7705 , P2_U7706 , P2_U7707 , P2_U7708 , P2_U7709 , P2_U7710;
wire P2_U7711 , P2_U7712 , P2_U7713 , P2_U7714 , P2_U7715 , P2_U7716 , P2_U7717 , P2_U7718 , P2_U7719 , P2_U7720;
wire P2_U7721 , P2_U7722 , P2_U7723 , P2_U7724 , P2_U7725 , P2_U7726 , P2_U7727 , P2_U7728 , P2_U7729 , P2_U7730;
wire P2_U7731 , P2_U7732 , P2_U7733 , P2_U7734 , P2_U7735 , P2_U7736 , P2_U7737 , P2_U7738 , P2_U7739 , P2_U7740;
wire P2_U7741 , P2_U7742 , P2_U7743 , P2_U7744 , P2_U7745 , P2_U7746 , P2_U7747 , P2_U7748 , P2_U7749 , P2_U7750;
wire P2_U7751 , P2_U7752 , P2_U7753 , P2_U7754 , P2_U7755 , P2_U7756 , P2_U7757 , P2_U7758 , P2_U7759 , P2_U7760;
wire P2_U7761 , P2_U7762 , P2_U7763 , P2_U7764 , P2_U7765 , P2_U7766 , P2_U7767 , P2_U7768 , P2_U7769 , P2_U7770;
wire P2_U7771 , P2_U7772 , P2_U7773 , P2_U7774 , P2_U7775 , P2_U7776 , P2_U7777 , P2_U7778 , P2_U7779 , P2_U7780;
wire P2_U7781 , P2_U7782 , P2_U7783 , P2_U7784 , P2_U7785 , P2_U7786 , P2_U7787 , P2_U7788 , P2_U7789 , P2_U7790;
wire P2_U7791 , P2_U7792 , P2_U7793 , P2_U7794 , P2_U7795 , P2_U7796 , P2_U7797 , P2_U7798 , P2_U7799 , P2_U7800;
wire P2_U7801 , P2_U7802 , P2_U7803 , P2_U7804 , P2_U7805 , P2_U7806 , P2_U7807 , P2_U7808 , P2_U7809 , P2_U7810;
wire P2_U7811 , P2_U7812 , P2_U7813 , P2_U7814 , P2_U7815 , P2_U7816 , P2_U7817 , P2_U7818 , P2_U7819 , P2_U7820;
wire P2_U7821 , P2_U7822 , P2_U7823 , P2_U7824 , P2_U7825 , P2_U7826 , P2_U7827 , P2_U7828 , P2_U7829 , P2_U7830;
wire P2_U7831 , P2_U7832 , P2_U7833 , P2_U7834 , P2_U7835 , P2_U7836 , P2_U7837 , P2_U7838 , P2_U7839 , P2_U7840;
wire P2_U7841 , P2_U7842 , P2_U7843 , P2_U7844 , P2_U7845 , P2_U7846 , P2_U7847 , P2_U7848 , P2_U7849 , P2_U7850;
wire P2_U7851 , P2_U7852 , P2_U7853 , P2_U7854 , P2_U7855 , P2_U7856 , P2_U7857 , P2_U7858 , P2_U7859 , P2_U7860;
wire P2_U7861 , P2_U7862 , P2_U7863 , P2_U7864 , P2_U7865 , P2_U7866 , P2_U7867 , P2_U7868 , P2_U7869 , P2_U7870;
wire P2_U7871 , P2_U7872 , P2_U7873 , P2_U7874 , P2_U7875 , P2_U7876 , P2_U7877 , P2_U7878 , P2_U7879 , P2_U7880;
wire P2_U7881 , P2_U7882 , P2_U7883 , P2_U7884 , P2_U7885 , P2_U7886 , P2_U7887 , P2_U7888 , P2_U7889 , P2_U7890;
wire P2_U7891 , P2_U7892 , P2_U7893 , P2_U7894 , P2_U7895 , P2_U7896 , P2_U7897 , P2_U7898 , P2_U7899 , P2_U7900;
wire P2_U7901 , P2_U7902 , P2_U7903 , P2_U7904 , P2_U7905 , P2_U7906 , P2_U7907 , P2_U7908 , P2_U7909 , P2_U7910;
wire P2_U7911 , P2_U7912 , P2_U7913 , P2_U7914 , P2_U7915 , P2_U7916 , P2_U7917 , P2_U7918 , P2_U7919 , P2_U7920;
wire P2_U7921 , P2_U7922 , P2_U7923 , P2_U7924 , P2_U7925 , P2_U7926 , P2_U7927 , P2_U7928 , P2_U7929 , P2_U7930;
wire P2_U7931 , P2_U7932 , P2_U7933 , P2_U7934 , P2_U7935 , P2_U7936 , P2_U7937 , P2_U7938 , P2_U7939 , P2_U7940;
wire P2_U7941 , P2_U7942 , P2_U7943 , P2_U7944 , P2_U7945 , P2_U7946 , P2_U7947 , P2_U7948 , P2_U7949 , P2_U7950;
wire P2_U7951 , P2_U7952 , P2_U7953 , P2_U7954 , P2_U7955 , P2_U7956 , P2_U7957 , P2_U7958 , P2_U7959 , P2_U7960;
wire P2_U7961 , P2_U7962 , P2_U7963 , P2_U7964 , P2_U7965 , P2_U7966 , P2_U7967 , P2_U7968 , P2_U7969 , P2_U7970;
wire P2_U7971 , P2_U7972 , P2_U7973 , P2_U7974 , P2_U7975 , P2_U7976 , P2_U7977 , P2_U7978 , P2_U7979 , P2_U7980;
wire P2_U7981 , P2_U7982 , P2_U7983 , P2_U7984 , P2_U7985 , P2_U7986 , P2_U7987 , P2_U7988 , P2_U7989 , P2_U7990;
wire P2_U7991 , P2_U7992 , P2_U7993 , P2_U7994 , P2_U7995 , P2_U7996 , P2_U7997 , P2_U7998 , P2_U7999 , P2_U8000;
wire P2_U8001 , P2_U8002 , P2_U8003 , P2_U8004 , P2_U8005 , P2_U8006 , P2_U8007 , P2_U8008 , P2_U8009 , P2_U8010;
wire P2_U8011 , P2_U8012 , P2_U8013 , P2_U8014 , P2_U8015 , P2_U8016 , P2_U8017 , P2_U8018 , P2_U8019 , P2_U8020;
wire P2_U8021 , P2_U8022 , P2_U8023 , P2_U8024 , P2_U8025 , P2_U8026 , P2_U8027 , P2_U8028 , P2_U8029 , P2_U8030;
wire P2_U8031 , P2_U8032 , P2_U8033 , P2_U8034 , P2_U8035 , P2_U8036 , P2_U8037 , P2_U8038 , P2_U8039 , P2_U8040;
wire P2_U8041 , P2_U8042 , P2_U8043 , P2_U8044 , P2_U8045 , P2_U8046 , P2_U8047 , P2_U8048 , P2_U8049 , P2_U8050;
wire P2_U8051 , P2_U8052 , P2_U8053 , P2_U8054 , P2_U8055 , P2_U8056 , P2_U8057 , P2_U8058 , P2_U8059 , P2_U8060;
wire P2_U8061 , P2_U8062 , P2_U8063 , P2_U8064 , P2_U8065 , P2_U8066 , P2_U8067 , P2_U8068 , P2_U8069 , P2_U8070;
wire P2_U8071 , P2_U8072 , P2_U8073 , P2_U8074 , P2_U8075 , P2_U8076 , P2_U8077 , P2_U8078 , P2_U8079 , P2_U8080;
wire P2_U8081 , P2_U8082 , P2_U8083 , P2_U8084 , P2_U8085 , P2_U8086 , P2_U8087 , P2_U8088 , P2_U8089 , P2_U8090;
wire P2_U8091 , P2_U8092 , P2_U8093 , P2_U8094 , P2_U8095 , P2_U8096 , P2_U8097 , P2_U8098 , P2_U8099 , P2_U8100;
wire P2_U8101 , P2_U8102 , P2_U8103 , P2_U8104 , P2_U8105 , P2_U8106 , P2_U8107 , P2_U8108 , P2_U8109 , P2_U8110;
wire P2_U8111 , P2_U8112 , P2_U8113 , P2_U8114 , P2_U8115 , P2_U8116 , P2_U8117 , P2_U8118 , P2_U8119 , P2_U8120;
wire P2_U8121 , P2_U8122 , P2_U8123 , P2_U8124 , P2_U8125 , P2_U8126 , P2_U8127 , P2_U8128 , P2_U8129 , P2_U8130;
wire P2_U8131 , P2_U8132 , P2_U8133 , P2_U8134 , P2_U8135 , P2_U8136 , P2_U8137 , P2_U8138 , P2_U8139 , P2_U8140;
wire P2_U8141 , P2_U8142 , P2_U8143 , P2_U8144 , P2_U8145 , P2_U8146 , P2_U8147 , P2_U8148 , P2_U8149 , P2_U8150;
wire P2_U8151 , P2_U8152 , P2_U8153 , P2_U8154 , P2_U8155 , P2_U8156 , P2_U8157 , P2_U8158 , P2_U8159 , P2_U8160;
wire P2_U8161 , P2_U8162 , P2_U8163 , P2_U8164 , P2_U8165 , P2_U8166 , P2_U8167 , P2_U8168 , P2_U8169 , P2_U8170;
wire P2_U8171 , P2_U8172 , P2_U8173 , P2_U8174 , P2_U8175 , P2_U8176 , P2_U8177 , P2_U8178 , P2_U8179 , P2_U8180;
wire P2_U8181 , P2_U8182 , P2_U8183 , P2_U8184 , P2_U8185 , P2_U8186 , P2_U8187 , P2_U8188 , P2_U8189 , P2_U8190;
wire P2_U8191 , P2_U8192 , P2_U8193 , P2_U8194 , P2_U8195 , P2_U8196 , P2_U8197 , P2_U8198 , P2_U8199 , P2_U8200;
wire P2_U8201 , P2_U8202 , P2_U8203 , P2_U8204 , P2_U8205 , P2_U8206 , P2_U8207 , P2_U8208 , P2_U8209 , P2_U8210;
wire P2_U8211 , P2_U8212 , P2_U8213 , P2_U8214 , P2_U8215 , P2_U8216 , P2_U8217 , P2_U8218 , P2_U8219 , P2_U8220;
wire P2_U8221 , P2_U8222 , P2_U8223 , P2_U8224 , P2_U8225 , P2_U8226 , P2_U8227 , P2_U8228 , P2_U8229 , P2_U8230;
wire P2_U8231 , P2_U8232 , P2_U8233 , P2_U8234 , P2_U8235 , P2_U8236 , P2_U8237 , P2_U8238 , P2_U8239 , P2_U8240;
wire P2_U8241 , P2_U8242 , P2_U8243 , P2_U8244 , P2_U8245 , P2_U8246 , P2_U8247 , P2_U8248 , P2_U8249 , P2_U8250;
wire P2_U8251 , P2_U8252 , P2_U8253 , P2_U8254 , P2_U8255 , P2_U8256 , P2_U8257 , P2_U8258 , P2_U8259 , P2_U8260;
wire P2_U8261 , P2_U8262 , P2_U8263 , P2_U8264 , P2_U8265 , P2_U8266 , P2_U8267 , P2_U8268 , P2_U8269 , P2_U8270;
wire P2_U8271 , P2_U8272 , P2_U8273 , P2_U8274 , P2_U8275 , P2_U8276 , P2_U8277 , P2_U8278 , P2_U8279 , P2_U8280;
wire P2_U8281 , P2_U8282 , P2_U8283 , P2_U8284 , P2_U8285 , P2_U8286 , P2_U8287 , P2_U8288 , P2_U8289 , P2_U8290;
wire P2_U8291 , P2_U8292 , P2_U8293 , P2_U8294 , P2_U8295 , P2_U8296 , P2_U8297 , P2_U8298 , P2_U8299 , P2_U8300;
wire P2_U8301 , P2_U8302 , P2_U8303 , P2_U8304 , P2_U8305 , P2_U8306 , P2_U8307 , P2_U8308 , P2_U8309 , P2_U8310;
wire P2_U8311 , P2_U8312 , P2_U8313 , P2_U8314 , P2_U8315 , P2_U8316 , P2_U8317 , P2_U8318 , P2_U8319 , P2_U8320;
wire P2_U8321 , P2_U8322 , P2_U8323 , P2_U8324 , P2_U8325 , P2_U8326 , P2_U8327 , P2_U8328 , P2_U8329 , P2_U8330;
wire P2_U8331 , P2_U8332 , P2_U8333 , P2_U8334 , P2_U8335 , P2_U8336 , P2_U8337 , P2_U8338 , P2_U8339 , P2_U8340;
wire P2_U8341 , P2_U8342 , P2_U8343 , P2_U8344 , P2_U8345 , P2_U8346 , P2_U8347 , P2_U8348 , P2_U8349 , P2_U8350;
wire P2_U8351 , P2_U8352 , P2_U8353 , P2_U8354 , P2_U8355 , P2_U8356 , P2_U8357 , P2_U8358 , P2_U8359 , P2_U8360;
wire P2_U8361 , P2_U8362 , P2_U8363 , P2_U8364 , P2_U8365 , P2_U8366 , P2_U8367 , P2_U8368 , P2_U8369 , P2_U8370;
wire P2_U8371 , P2_U8372 , P2_U8373 , P2_U8374 , P2_U8375 , P2_U8376 , P2_U8377 , P2_U8378 , P2_U8379 , P2_U8380;
wire P2_U8381 , P2_U8382 , P2_U8383 , P2_U8384 , P2_U8385 , P2_U8386 , P2_U8387 , P2_U8388 , P2_U8389 , P2_U8390;
wire P2_U8391 , P2_U8392 , P2_U8393 , P2_U8394 , P2_U8395 , P2_U8396 , P2_U8397 , P2_U8398 , P2_U8399 , P2_U8400;
wire P2_U8401 , P2_U8402 , P2_U8403 , P2_U8404 , P2_U8405 , P2_U8406 , P2_U8407 , P2_U8408 , P2_U8409 , P2_U8410;
wire P2_U8411 , P2_U8412 , P2_U8413 , P2_U8414 , P2_U8415 , P2_U8416 , P2_U8417 , P2_U8418 , P2_U8419 , P2_U8420;
wire P2_U8421 , P2_U8422 , P2_U8423 , P2_U8424 , P2_U8425 , P2_U8426 , P2_U8427 , P2_U8428 , P2_U8429 , P2_U8430;
wire P2_U8431 , P2_U8432 , P2_U8433 , P2_U8434 , P1_ADD_405_U171 , P1_ADD_405_U170 , P1_ADD_405_U169 , P1_ADD_405_U168 , P1_ADD_405_U167 , P1_ADD_405_U166;
wire P1_ADD_405_U165 , P1_ADD_405_U164 , P1_ADD_405_U163 , P1_ADD_405_U162 , P1_ADD_405_U161 , P1_ADD_405_U160 , P1_ADD_405_U159 , P1_ADD_405_U158 , P1_ADD_405_U157 , P1_ADD_405_U156;
wire P1_ADD_405_U155 , P1_ADD_405_U154 , P1_ADD_405_U153 , P1_ADD_405_U152 , P1_ADD_405_U151 , P1_ADD_405_U150 , P1_ADD_405_U149 , P1_ADD_405_U148 , P1_ADD_405_U147 , P1_ADD_405_U146;
wire P1_ADD_405_U145 , P1_ADD_405_U144 , P1_ADD_405_U143 , P1_ADD_405_U142 , P1_ADD_405_U141 , P1_ADD_405_U140 , P1_ADD_405_U139 , P1_ADD_405_U138 , P1_ADD_405_U137 , P1_ADD_405_U136;
wire P1_ADD_405_U135 , P1_ADD_405_U134 , P1_ADD_405_U133 , P1_ADD_405_U132 , P1_ADD_405_U131 , P1_ADD_405_U130 , P1_ADD_405_U129 , P1_ADD_405_U128 , P1_ADD_405_U127 , P1_ADD_405_U126;
wire P1_ADD_405_U125 , P1_ADD_405_U124 , P1_ADD_405_U123 , P1_ADD_405_U122 , P1_ADD_405_U121 , P1_ADD_405_U120 , P1_ADD_405_U119 , P1_ADD_405_U118 , P1_ADD_405_U117 , P1_ADD_405_U116;
wire P1_ADD_405_U115 , P1_U2352 , P1_U2353 , P1_U2354 , P1_U2355 , P1_U2356 , P1_U2357 , P1_U2358 , P1_U2359 , P1_U2360;
wire P1_U2361 , P1_U2362 , P1_U2363 , P1_U2364 , P1_U2365 , P1_U2366 , P1_U2367 , P1_U2368 , P1_U2369 , P1_U2370;
wire P1_U2371 , P1_U2372 , P1_U2373 , P1_U2374 , P1_U2375 , P1_U2376 , P1_U2377 , P1_U2378 , P1_U2379 , P1_U2380;
wire P1_U2381 , P1_U2382 , P1_U2383 , P1_U2384 , P1_U2385 , P1_U2386 , P1_U2387 , P1_U2388 , P1_U2389 , P1_U2390;
wire P1_U2391 , P1_U2392 , P1_U2393 , P1_U2394 , P1_U2395 , P1_U2396 , P1_U2397 , P1_U2398 , P1_U2399 , P1_U2400;
wire P1_U2401 , P1_U2402 , P1_U2403 , P1_U2404 , P1_U2405 , P1_U2406 , P1_U2407 , P1_U2408 , P1_U2409 , P1_U2410;
wire P1_U2411 , P1_U2412 , P1_U2413 , P1_U2414 , P1_U2415 , P1_U2416 , P1_U2417 , P1_U2418 , P1_U2419 , P1_U2420;
wire P1_U2421 , P1_U2422 , P1_U2423 , P1_U2424 , P1_U2425 , P1_U2426 , P1_U2427 , P1_U2428 , P1_U2429 , P1_U2430;
wire P1_U2431 , P1_U2432 , P1_U2433 , P1_U2434 , P1_U2435 , P1_U2436 , P1_U2437 , P1_U2438 , P1_U2439 , P1_U2440;
wire P1_U2441 , P1_U2442 , P1_U2443 , P1_U2444 , P1_U2445 , P1_U2446 , P1_U2447 , P1_U2448 , P1_U2449 , P1_U2450;
wire P1_U2451 , P1_U2452 , P1_U2453 , P1_U2454 , P1_U2455 , P1_U2456 , P1_U2457 , P1_U2458 , P1_U2459 , P1_U2460;
wire P1_U2461 , P1_U2462 , P1_U2463 , P1_U2464 , P1_U2465 , P1_U2466 , P1_U2467 , P1_U2468 , P1_U2469 , P1_U2470;
wire P1_U2471 , P1_U2472 , P1_U2473 , P1_U2474 , P1_U2475 , P1_U2476 , P1_U2477 , P1_U2478 , P1_U2479 , P1_U2480;
wire P1_U2481 , P1_U2482 , P1_U2483 , P1_U2484 , P1_U2485 , P1_U2486 , P1_U2487 , P1_U2488 , P1_U2489 , P1_U2490;
wire P1_U2491 , P1_U2492 , P1_U2493 , P1_U2494 , P1_U2495 , P1_U2496 , P1_U2497 , P1_U2498 , P1_U2499 , P1_U2500;
wire P1_U2501 , P1_U2502 , P1_U2503 , P1_U2504 , P1_U2505 , P1_U2506 , P1_U2507 , P1_U2508 , P1_U2509 , P1_U2510;
wire P1_U2511 , P1_U2512 , P1_U2513 , P1_U2514 , P1_U2515 , P1_U2516 , P1_U2517 , P1_U2518 , P1_U2519 , P1_U2520;
wire P1_U2521 , P1_U2522 , P1_U2523 , P1_U2524 , P1_U2525 , P1_U2526 , P1_U2527 , P1_U2528 , P1_U2529 , P1_U2530;
wire P1_U2531 , P1_U2532 , P1_U2533 , P1_U2534 , P1_U2535 , P1_U2536 , P1_U2537 , P1_U2538 , P1_U2539 , P1_U2540;
wire P1_U2541 , P1_U2542 , P1_U2543 , P1_U2544 , P1_U2545 , P1_U2546 , P1_U2547 , P1_U2548 , P1_U2549 , P1_U2550;
wire P1_U2551 , P1_U2552 , P1_U2553 , P1_U2554 , P1_U2555 , P1_U2556 , P1_U2557 , P1_U2558 , P1_U2559 , P1_U2560;
wire P1_U2561 , P1_U2562 , P1_U2563 , P1_U2564 , P1_U2565 , P1_U2566 , P1_U2567 , P1_U2568 , P1_U2569 , P1_U2570;
wire P1_U2571 , P1_U2572 , P1_U2573 , P1_U2574 , P1_U2575 , P1_U2576 , P1_U2577 , P1_U2578 , P1_U2579 , P1_U2580;
wire P1_U2581 , P1_U2582 , P1_U2583 , P1_U2584 , P1_U2585 , P1_U2586 , P1_U2587 , P1_U2588 , P1_U2589 , P1_U2590;
wire P1_U2591 , P1_U2592 , P1_U2593 , P1_U2594 , P1_U2595 , P1_U2596 , P1_U2597 , P1_U2598 , P1_U2599 , P1_U2600;
wire P1_U2601 , P1_U2602 , P1_U2603 , P1_U2604 , P1_U2605 , P1_U2606 , P1_U2607 , P1_U2608 , P1_U2609 , P1_U2610;
wire P1_U2611 , P1_U2612 , P1_U2613 , P1_U2614 , P1_U2615 , P1_U2616 , P1_U2617 , P1_U2618 , P1_ADD_405_U114 , P1_U2620;
wire P1_U2621 , P1_U2622 , P1_U2623 , P1_U2624 , P1_U2625 , P1_U2626 , P1_U2627 , P1_U2628 , P1_U2629 , P1_U2630;
wire P1_U2631 , P1_U2632 , P1_U2633 , P1_U2634 , P1_U2635 , P1_U2636 , P1_U2637 , P1_U2638 , P1_U2639 , P1_U2640;
wire P1_U2641 , P1_U2642 , P1_U2643 , P1_U2644 , P1_U2645 , P1_U2646 , P1_U2647 , P1_U2648 , P1_U2649 , P1_U2650;
wire P1_U2651 , P1_U2652 , P1_U2653 , P1_U2654 , P1_U2655 , P1_U2656 , P1_U2657 , P1_U2658 , P1_U2659 , P1_U2660;
wire P1_U2661 , P1_U2662 , P1_U2663 , P1_U2664 , P1_U2665 , P1_U2666 , P1_U2667 , P1_U2668 , P1_U2669 , P1_U2670;
wire P1_U2671 , P1_U2672 , P1_U2673 , P1_U2674 , P1_U2675 , P1_U2676 , P1_U2677 , P1_U2678 , P1_U2679 , P1_U2680;
wire P1_U2681 , P1_U2682 , P1_U2683 , P1_U2684 , P1_U2685 , P1_U2686 , P1_U2687 , P1_U2688 , P1_U2689 , P1_U2690;
wire P1_U2691 , P1_U2692 , P1_U2693 , P1_U2694 , P1_U2695 , P1_U2696 , P1_U2697 , P1_U2698 , P1_U2699 , P1_U2700;
wire P1_U2701 , P1_U2702 , P1_U2703 , P1_U2704 , P1_U2705 , P1_U2706 , P1_U2707 , P1_U2708 , P1_U2709 , P1_U2710;
wire P1_U2711 , P1_U2712 , P1_U2713 , P1_U2714 , P1_U2715 , P1_U2716 , P1_U2717 , P1_U2718 , P1_U2719 , P1_U2720;
wire P1_U2721 , P1_U2722 , P1_U2723 , P1_U2724 , P1_U2725 , P1_U2726 , P1_U2727 , P1_U2728 , P1_U2729 , P1_U2730;
wire P1_U2731 , P1_U2732 , P1_U2733 , P1_U2734 , P1_U2735 , P1_U2736 , P1_U2737 , P1_U2738 , P1_U2739 , P1_U2740;
wire P1_U2741 , P1_U2742 , P1_U2743 , P1_U2744 , P1_U2745 , P1_U2746 , P1_U2747 , P1_U2748 , P1_U2749 , P1_U2750;
wire P1_U2751 , P1_U2752 , P1_U2753 , P1_U2754 , P1_U2755 , P1_U2756 , P1_U2757 , P1_U2758 , P1_U2759 , P1_U2760;
wire P1_U2761 , P1_U2762 , P1_U2763 , P1_U2764 , P1_U2765 , P1_U2766 , P1_U2767 , P1_U2768 , P1_U2769 , P1_U2770;
wire P1_U2771 , P1_U2772 , P1_U2773 , P1_U2774 , P1_U2775 , P1_U2776 , P1_U2777 , P1_U2778 , P1_U2779 , P1_U2780;
wire P1_U2781 , P1_U2782 , P1_U2783 , P1_U2784 , P1_U2785 , P1_U2786 , P1_U2787 , P1_U2788 , P1_U2789 , P1_U2790;
wire P1_U2791 , P1_U2792 , P1_U2793 , P1_U2794 , P1_U2795 , P1_U2796 , P1_U2797 , P1_U2798 , P1_U2799 , P1_U2800;
wire P1_U3227 , P1_U3228 , P1_U3229 , P1_U3230 , P1_U3231 , P1_U3232 , P1_U3233 , P1_U3234 , P1_U3235 , P1_U3236;
wire P1_U3237 , P1_U3238 , P1_U3239 , P1_U3240 , P1_U3241 , P1_U3242 , P1_U3243 , P1_U3244 , P1_U3245 , P1_U3246;
wire P1_U3247 , P1_U3248 , P1_U3249 , P1_U3250 , P1_U3251 , P1_U3252 , P1_U3253 , P1_U3254 , P1_U3255 , P1_U3256;
wire P1_U3257 , P1_U3258 , P1_U3259 , P1_U3260 , P1_U3261 , P1_U3262 , P1_U3263 , P1_U3264 , P1_U3265 , P1_U3266;
wire P1_U3267 , P1_U3268 , P1_U3269 , P1_U3270 , P1_U3271 , P1_U3272 , P1_U3273 , P1_U3274 , P1_U3275 , P1_U3276;
wire P1_U3277 , P1_U3278 , P1_U3279 , P1_U3280 , P1_U3281 , P1_U3282 , P1_U3283 , P1_U3284 , P1_U3285 , P1_U3286;
wire P1_U3287 , P1_U3288 , P1_U3289 , P1_U3290 , P1_U3291 , P1_U3292 , P1_U3293 , P1_U3294 , P1_U3295 , P1_U3296;
wire P1_U3297 , P1_U3298 , P1_U3299 , P1_U3300 , P1_U3301 , P1_U3302 , P1_U3303 , P1_U3304 , P1_U3305 , P1_U3306;
wire P1_U3307 , P1_U3308 , P1_U3309 , P1_U3310 , P1_U3311 , P1_U3312 , P1_U3313 , P1_U3314 , P1_U3315 , P1_U3316;
wire P1_U3317 , P1_U3318 , P1_U3319 , P1_U3320 , P1_U3321 , P1_U3322 , P1_U3323 , P1_U3324 , P1_U3325 , P1_U3326;
wire P1_U3327 , P1_U3328 , P1_U3329 , P1_U3330 , P1_U3331 , P1_U3332 , P1_U3333 , P1_U3334 , P1_U3335 , P1_U3336;
wire P1_U3337 , P1_U3338 , P1_U3339 , P1_U3340 , P1_U3341 , P1_U3342 , P1_U3343 , P1_U3344 , P1_U3345 , P1_U3346;
wire P1_U3347 , P1_U3348 , P1_U3349 , P1_U3350 , P1_U3351 , P1_U3352 , P1_U3353 , P1_U3354 , P1_U3355 , P1_U3356;
wire P1_U3357 , P1_U3358 , P1_U3359 , P1_U3360 , P1_U3361 , P1_U3362 , P1_U3363 , P1_U3364 , P1_U3365 , P1_U3366;
wire P1_U3367 , P1_U3368 , P1_U3369 , P1_U3370 , P1_U3371 , P1_U3372 , P1_U3373 , P1_U3374 , P1_U3375 , P1_U3376;
wire P1_U3377 , P1_U3378 , P1_U3379 , P1_U3380 , P1_U3381 , P1_U3382 , P1_U3383 , P1_U3384 , P1_U3385 , P1_U3386;
wire P1_U3387 , P1_U3388 , P1_U3389 , P1_U3390 , P1_U3391 , P1_U3392 , P1_U3393 , P1_U3394 , P1_U3395 , P1_U3396;
wire P1_U3397 , P1_U3398 , P1_U3399 , P1_U3400 , P1_U3401 , P1_U3402 , P1_U3403 , P1_U3404 , P1_U3405 , P1_U3406;
wire P1_U3407 , P1_U3408 , P1_U3409 , P1_U3410 , P1_U3411 , P1_U3412 , P1_U3413 , P1_U3414 , P1_U3415 , P1_U3416;
wire P1_U3417 , P1_U3418 , P1_U3419 , P1_U3420 , P1_U3421 , P1_U3422 , P1_U3423 , P1_U3424 , P1_U3425 , P1_U3426;
wire P1_U3427 , P1_U3428 , P1_U3429 , P1_U3430 , P1_U3431 , P1_U3432 , P1_U3433 , P1_U3434 , P1_U3435 , P1_U3436;
wire P1_U3437 , P1_U3438 , P1_U3439 , P1_U3440 , P1_U3441 , P1_U3442 , P1_U3443 , P1_U3444 , P1_U3445 , P1_U3446;
wire P1_U3447 , P1_U3448 , P1_U3449 , P1_U3450 , P1_U3451 , P1_U3452 , P1_U3453 , P1_U3454 , P1_U3455 , P1_U3456;
wire P1_U3457 , P1_U3462 , P1_U3463 , P1_U3467 , P1_U3470 , P1_U3471 , P1_U3479 , P1_U3480 , P1_U3488 , P1_U3489;
wire P1_U3490 , P1_U3491 , P1_U3492 , P1_U3493 , P1_U3494 , P1_U3495 , P1_U3496 , P1_U3497 , P1_U3498 , P1_U3499;
wire P1_U3500 , P1_U3501 , P1_U3502 , P1_U3503 , P1_U3504 , P1_U3505 , P1_U3506 , P1_U3507 , P1_U3508 , P1_U3509;
wire P1_U3510 , P1_U3511 , P1_U3512 , P1_U3513 , P1_U3514 , P1_U3515 , P1_U3516 , P1_U3517 , P1_U3518 , P1_U3519;
wire P1_U3520 , P1_U3521 , P1_U3522 , P1_U3523 , P1_U3524 , P1_U3525 , P1_U3526 , P1_U3527 , P1_U3528 , P1_U3529;
wire P1_U3530 , P1_U3531 , P1_U3532 , P1_U3533 , P1_U3534 , P1_U3535 , P1_U3536 , P1_U3537 , P1_U3538 , P1_U3539;
wire P1_U3540 , P1_U3541 , P1_U3542 , P1_U3543 , P1_U3544 , P1_U3545 , P1_U3546 , P1_U3547 , P1_U3548 , P1_U3549;
wire P1_U3550 , P1_U3551 , P1_U3552 , P1_U3553 , P1_U3554 , P1_U3555 , P1_U3556 , P1_U3557 , P1_U3558 , P1_U3559;
wire P1_U3560 , P1_U3561 , P1_U3562 , P1_U3563 , P1_U3564 , P1_U3565 , P1_U3566 , P1_U3567 , P1_U3568 , P1_U3569;
wire P1_U3570 , P1_U3571 , P1_U3572 , P1_U3573 , P1_U3574 , P1_U3575 , P1_U3576 , P1_U3577 , P1_U3578 , P1_U3579;
wire P1_U3580 , P1_U3581 , P1_U3582 , P1_U3583 , P1_U3584 , P1_U3585 , P1_U3586 , P1_U3587 , P1_U3588 , P1_U3589;
wire P1_U3590 , P1_U3591 , P1_U3592 , P1_U3593 , P1_U3594 , P1_U3595 , P1_U3596 , P1_U3597 , P1_U3598 , P1_U3599;
wire P1_U3600 , P1_U3601 , P1_U3602 , P1_U3603 , P1_U3604 , P1_U3605 , P1_U3606 , P1_U3607 , P1_U3608 , P1_U3609;
wire P1_U3610 , P1_U3611 , P1_U3612 , P1_U3613 , P1_U3614 , P1_U3615 , P1_U3616 , P1_U3617 , P1_U3618 , P1_U3619;
wire P1_U3620 , P1_U3621 , P1_U3622 , P1_U3623 , P1_U3624 , P1_U3625 , P1_U3626 , P1_U3627 , P1_U3628 , P1_U3629;
wire P1_U3630 , P1_U3631 , P1_U3632 , P1_U3633 , P1_U3634 , P1_U3635 , P1_U3636 , P1_U3637 , P1_U3638 , P1_U3639;
wire P1_U3640 , P1_U3641 , P1_U3642 , P1_U3643 , P1_U3644 , P1_U3645 , P1_U3646 , P1_U3647 , P1_U3648 , P1_U3649;
wire P1_U3650 , P1_U3651 , P1_U3652 , P1_U3653 , P1_U3654 , P1_U3655 , P1_U3656 , P1_U3657 , P1_U3658 , P1_U3659;
wire P1_U3660 , P1_U3661 , P1_U3662 , P1_U3663 , P1_U3664 , P1_U3665 , P1_U3666 , P1_U3667 , P1_U3668 , P1_U3669;
wire P1_U3670 , P1_U3671 , P1_U3672 , P1_U3673 , P1_U3674 , P1_U3675 , P1_U3676 , P1_U3677 , P1_U3678 , P1_U3679;
wire P1_U3680 , P1_U3681 , P1_U3682 , P1_U3683 , P1_U3684 , P1_U3685 , P1_U3686 , P1_U3687 , P1_U3688 , P1_U3689;
wire P1_U3690 , P1_U3691 , P1_U3692 , P1_U3693 , P1_U3694 , P1_U3695 , P1_U3696 , P1_U3697 , P1_U3698 , P1_U3699;
wire P1_U3700 , P1_U3701 , P1_U3702 , P1_U3703 , P1_U3704 , P1_U3705 , P1_U3706 , P1_U3707 , P1_U3708 , P1_U3709;
wire P1_U3710 , P1_U3711 , P1_U3712 , P1_U3713 , P1_U3714 , P1_U3715 , P1_U3716 , P1_U3717 , P1_U3718 , P1_U3719;
wire P1_U3720 , P1_U3721 , P1_U3722 , P1_U3723 , P1_U3724 , P1_U3725 , P1_U3726 , P1_U3727 , P1_U3728 , P1_U3729;
wire P1_U3730 , P1_U3731 , P1_U3732 , P1_U3733 , P1_U3734 , P1_U3735 , P1_U3736 , P1_U3737 , P1_U3738 , P1_U3739;
wire P1_U3740 , P1_U3741 , P1_U3742 , P1_U3743 , P1_U3744 , P1_U3745 , P1_U3746 , P1_U3747 , P1_U3748 , P1_U3749;
wire P1_U3750 , P1_U3751 , P1_U3752 , P1_U3753 , P1_U3754 , P1_U3755 , P1_U3756 , P1_U3757 , P1_U3758 , P1_U3759;
wire P1_U3760 , P1_U3761 , P1_U3762 , P1_U3763 , P1_U3764 , P1_U3765 , P1_U3766 , P1_U3767 , P1_U3768 , P1_U3769;
wire P1_U3770 , P1_U3771 , P1_U3772 , P1_U3773 , P1_U3774 , P1_U3775 , P1_U3776 , P1_U3777 , P1_U3778 , P1_U3779;
wire P1_U3780 , P1_U3781 , P1_U3782 , P1_U3783 , P1_U3784 , P1_U3785 , P1_U3786 , P1_U3787 , P1_U3788 , P1_U3789;
wire P1_U3790 , P1_U3791 , P1_U3792 , P1_U3793 , P1_U3794 , P1_U3795 , P1_U3796 , P1_U3797 , P1_U3798 , P1_U3799;
wire P1_U3800 , P1_U3801 , P1_U3802 , P1_U3803 , P1_U3804 , P1_U3805 , P1_U3806 , P1_U3807 , P1_U3808 , P1_U3809;
wire P1_U3810 , P1_U3811 , P1_U3812 , P1_U3813 , P1_U3814 , P1_U3815 , P1_U3816 , P1_U3817 , P1_U3818 , P1_U3819;
wire P1_U3820 , P1_U3821 , P1_U3822 , P1_U3823 , P1_U3824 , P1_U3825 , P1_U3826 , P1_U3827 , P1_U3828 , P1_U3829;
wire P1_U3830 , P1_U3831 , P1_U3832 , P1_U3833 , P1_U3834 , P1_U3835 , P1_U3836 , P1_U3837 , P1_U3838 , P1_U3839;
wire P1_U3840 , P1_U3841 , P1_U3842 , P1_U3843 , P1_U3844 , P1_U3845 , P1_U3846 , P1_U3847 , P1_U3848 , P1_U3849;
wire P1_U3850 , P1_U3851 , P1_U3852 , P1_U3853 , P1_U3854 , P1_U3855 , P1_U3856 , P1_U3857 , P1_U3858 , P1_U3859;
wire P1_U3860 , P1_U3861 , P1_U3862 , P1_U3863 , P1_U3864 , P1_U3865 , P1_U3866 , P1_U3867 , P1_U3868 , P1_U3869;
wire P1_U3870 , P1_U3871 , P1_U3872 , P1_U3873 , P1_U3874 , P1_U3875 , P1_U3876 , P1_U3877 , P1_U3878 , P1_U3879;
wire P1_U3880 , P1_U3881 , P1_U3882 , P1_U3883 , P1_U3884 , P1_U3885 , P1_U3886 , P1_U3887 , P1_U3888 , P1_U3889;
wire P1_U3890 , P1_U3891 , P1_U3892 , P1_U3893 , P1_U3894 , P1_U3895 , P1_U3896 , P1_U3897 , P1_U3898 , P1_U3899;
wire P1_U3900 , P1_U3901 , P1_U3902 , P1_U3903 , P1_U3904 , P1_U3905 , P1_U3906 , P1_U3907 , P1_U3908 , P1_U3909;
wire P1_U3910 , P1_U3911 , P1_U3912 , P1_U3913 , P1_U3914 , P1_U3915 , P1_U3916 , P1_U3917 , P1_U3918 , P1_U3919;
wire P1_U3920 , P1_U3921 , P1_U3922 , P1_U3923 , P1_U3924 , P1_U3925 , P1_U3926 , P1_U3927 , P1_U3928 , P1_U3929;
wire P1_U3930 , P1_U3931 , P1_U3932 , P1_U3933 , P1_U3934 , P1_U3935 , P1_U3936 , P1_U3937 , P1_U3938 , P1_U3939;
wire P1_U3940 , P1_U3941 , P1_U3942 , P1_U3943 , P1_U3944 , P1_U3945 , P1_U3946 , P1_U3947 , P1_U3948 , P1_U3949;
wire P1_U3950 , P1_U3951 , P1_U3952 , P1_U3953 , P1_U3954 , P1_U3955 , P1_U3956 , P1_U3957 , P1_U3958 , P1_U3959;
wire P1_U3960 , P1_U3961 , P1_U3962 , P1_U3963 , P1_U3964 , P1_U3965 , P1_U3966 , P1_U3967 , P1_U3968 , P1_U3969;
wire P1_U3970 , P1_U3971 , P1_U3972 , P1_U3973 , P1_U3974 , P1_U3975 , P1_U3976 , P1_U3977 , P1_U3978 , P1_U3979;
wire P1_U3980 , P1_U3981 , P1_U3982 , P1_U3983 , P1_U3984 , P1_U3985 , P1_U3986 , P1_U3987 , P1_U3988 , P1_U3989;
wire P1_U3990 , P1_U3991 , P1_U3992 , P1_U3993 , P1_U3994 , P1_U3995 , P1_U3996 , P1_U3997 , P1_U3998 , P1_U3999;
wire P1_U4000 , P1_U4001 , P1_U4002 , P1_U4003 , P1_U4004 , P1_U4005 , P1_U4006 , P1_U4007 , P1_U4008 , P1_U4009;
wire P1_U4010 , P1_U4011 , P1_U4012 , P1_U4013 , P1_U4014 , P1_U4015 , P1_U4016 , P1_U4017 , P1_U4018 , P1_U4019;
wire P1_U4020 , P1_U4021 , P1_U4022 , P1_U4023 , P1_U4024 , P1_U4025 , P1_U4026 , P1_U4027 , P1_U4028 , P1_U4029;
wire P1_U4030 , P1_U4031 , P1_U4032 , P1_U4033 , P1_U4034 , P1_U4035 , P1_U4036 , P1_U4037 , P1_U4038 , P1_U4039;
wire P1_U4040 , P1_U4041 , P1_U4042 , P1_U4043 , P1_U4044 , P1_U4045 , P1_U4046 , P1_U4047 , P1_U4048 , P1_U4049;
wire P1_U4050 , P1_U4051 , P1_U4052 , P1_U4053 , P1_U4054 , P1_U4055 , P1_U4056 , P1_U4057 , P1_U4058 , P1_U4059;
wire P1_U4060 , P1_U4061 , P1_U4062 , P1_U4063 , P1_U4064 , P1_U4065 , P1_U4066 , P1_U4067 , P1_U4068 , P1_U4069;
wire P1_U4070 , P1_U4071 , P1_U4072 , P1_U4073 , P1_U4074 , P1_U4075 , P1_U4076 , P1_U4077 , P1_U4078 , P1_U4079;
wire P1_U4080 , P1_U4081 , P1_U4082 , P1_U4083 , P1_U4084 , P1_U4085 , P1_U4086 , P1_U4087 , P1_U4088 , P1_U4089;
wire P1_U4090 , P1_U4091 , P1_U4092 , P1_U4093 , P1_U4094 , P1_U4095 , P1_U4096 , P1_U4097 , P1_U4098 , P1_U4099;
wire P1_U4100 , P1_U4101 , P1_U4102 , P1_U4103 , P1_U4104 , P1_U4105 , P1_U4106 , P1_U4107 , P1_U4108 , P1_U4109;
wire P1_U4110 , P1_U4111 , P1_U4112 , P1_U4113 , P1_U4114 , P1_U4115 , P1_U4116 , P1_U4117 , P1_U4118 , P1_U4119;
wire P1_U4120 , P1_U4121 , P1_U4122 , P1_U4123 , P1_U4124 , P1_U4125 , P1_U4126 , P1_U4127 , P1_U4128 , P1_U4129;
wire P1_U4130 , P1_U4131 , P1_U4132 , P1_U4133 , P1_U4134 , P1_U4135 , P1_U4136 , P1_U4137 , P1_U4138 , P1_U4139;
wire P1_U4140 , P1_U4141 , P1_U4142 , P1_U4143 , P1_U4144 , P1_U4145 , P1_U4146 , P1_U4147 , P1_U4148 , P1_U4149;
wire P1_U4150 , P1_U4151 , P1_U4152 , P1_U4153 , P1_U4154 , P1_U4155 , P1_U4156 , P1_U4157 , P1_U4158 , P1_U4159;
wire P1_U4160 , P1_U4161 , P1_U4162 , P1_U4163 , P1_U4164 , P1_U4165 , P1_U4166 , P1_U4167 , P1_U4168 , P1_U4169;
wire P1_U4170 , P1_U4171 , P1_U4172 , P1_U4173 , P1_U4174 , P1_U4175 , P1_U4176 , P1_U4177 , P1_U4178 , P1_U4179;
wire P1_U4180 , P1_U4181 , P1_U4182 , P1_U4183 , P1_U4184 , P1_U4185 , P1_U4186 , P1_U4187 , P1_U4188 , P1_U4189;
wire P1_U4190 , P1_U4191 , P1_U4192 , P1_U4193 , P1_U4194 , P1_U4195 , P1_U4196 , P1_U4197 , P1_U4198 , P1_U4199;
wire P1_U4200 , P1_U4201 , P1_U4202 , P1_U4203 , P1_U4204 , P1_U4205 , P1_U4206 , P1_U4207 , P1_U4208 , P1_U4209;
wire P1_U4210 , P1_U4211 , P1_U4212 , P1_U4213 , P1_U4214 , P1_U4215 , P1_U4216 , P1_U4217 , P1_U4218 , P1_U4219;
wire P1_U4220 , P1_U4221 , P1_U4222 , P1_U4223 , P1_U4224 , P1_U4225 , P1_U4226 , P1_U4227 , P1_U4228 , P1_U4229;
wire P1_U4230 , P1_U4231 , P1_U4232 , P1_U4233 , P1_U4234 , P1_U4235 , P1_U4236 , P1_U4237 , P1_U4238 , P1_U4239;
wire P1_U4240 , P1_U4241 , P1_U4242 , P1_U4243 , P1_U4244 , P1_U4245 , P1_U4246 , P1_U4247 , P1_U4248 , P1_U4249;
wire P1_U4250 , P1_U4251 , P1_U4252 , P1_U4253 , P1_U4254 , P1_U4255 , P1_U4256 , P1_U4257 , P1_U4258 , P1_U4259;
wire P1_U4260 , P1_U4261 , P1_U4262 , P1_U4263 , P1_U4264 , P1_U4265 , P1_U4266 , P1_U4267 , P1_U4268 , P1_U4269;
wire P1_U4270 , P1_U4271 , P1_U4272 , P1_U4273 , P1_U4274 , P1_U4275 , P1_U4276 , P1_U4277 , P1_U4278 , P1_U4279;
wire P1_U4280 , P1_U4281 , P1_U4282 , P1_U4283 , P1_U4284 , P1_U4285 , P1_U4286 , P1_U4287 , P1_U4288 , P1_U4289;
wire P1_U4290 , P1_U4291 , P1_U4292 , P1_U4293 , P1_U4294 , P1_U4295 , P1_U4296 , P1_U4297 , P1_U4298 , P1_U4299;
wire P1_U4300 , P1_U4301 , P1_U4302 , P1_U4303 , P1_U4304 , P1_U4305 , P1_U4306 , P1_U4307 , P1_U4308 , P1_U4309;
wire P1_U4310 , P1_U4311 , P1_U4312 , P1_U4313 , P1_U4314 , P1_U4315 , P1_U4316 , P1_U4317 , P1_U4318 , P1_U4319;
wire P1_U4320 , P1_U4321 , P1_U4322 , P1_U4323 , P1_U4324 , P1_U4325 , P1_U4326 , P1_U4327 , P1_U4328 , P1_U4329;
wire P1_U4330 , P1_U4331 , P1_U4332 , P1_U4333 , P1_U4334 , P1_U4335 , P1_U4336 , P1_U4337 , P1_U4338 , P1_U4339;
wire P1_U4340 , P1_U4341 , P1_U4342 , P1_U4343 , P1_U4344 , P1_U4345 , P1_U4346 , P1_U4347 , P1_U4348 , P1_U4349;
wire P1_U4350 , P1_U4351 , P1_U4352 , P1_U4353 , P1_U4354 , P1_U4355 , P1_U4356 , P1_U4357 , P1_U4358 , P1_U4359;
wire P1_U4360 , P1_U4361 , P1_U4362 , P1_U4363 , P1_U4364 , P1_U4365 , P1_U4366 , P1_U4367 , P1_U4368 , P1_U4369;
wire P1_U4370 , P1_U4371 , P1_U4372 , P1_U4373 , P1_U4374 , P1_U4375 , P1_U4376 , P1_U4377 , P1_U4378 , P1_U4379;
wire P1_U4380 , P1_U4381 , P1_U4382 , P1_U4383 , P1_U4384 , P1_U4385 , P1_U4386 , P1_U4387 , P1_U4388 , P1_U4389;
wire P1_U4390 , P1_U4391 , P1_U4392 , P1_U4393 , P1_U4394 , P1_U4395 , P1_U4396 , P1_U4397 , P1_U4398 , P1_U4399;
wire P1_U4400 , P1_U4401 , P1_U4402 , P1_U4403 , P1_U4404 , P1_U4405 , P1_U4406 , P1_U4407 , P1_U4408 , P1_U4409;
wire P1_U4410 , P1_U4411 , P1_U4412 , P1_U4413 , P1_U4414 , P1_U4415 , P1_U4416 , P1_U4417 , P1_U4418 , P1_U4419;
wire P1_U4420 , P1_U4421 , P1_U4422 , P1_U4423 , P1_U4424 , P1_U4425 , P1_U4426 , P1_U4427 , P1_U4428 , P1_U4429;
wire P1_U4430 , P1_U4431 , P1_U4432 , P1_U4433 , P1_U4434 , P1_U4435 , P1_U4436 , P1_U4437 , P1_U4438 , P1_U4439;
wire P1_U4440 , P1_U4441 , P1_U4442 , P1_U4443 , P1_U4444 , P1_U4445 , P1_U4446 , P1_U4447 , P1_U4448 , P1_U4449;
wire P1_U4450 , P1_U4451 , P1_U4452 , P1_U4453 , P1_U4454 , P1_U4455 , P1_U4456 , P1_U4457 , P1_U4458 , P1_U4459;
wire P1_U4460 , P1_U4461 , P1_U4462 , P1_U4463 , P1_U4464 , P1_U4465 , P1_U4466 , P1_U4467 , P1_U4468 , P1_U4469;
wire P1_U4470 , P1_U4471 , P1_U4472 , P1_U4473 , P1_U4474 , P1_U4475 , P1_U4476 , P1_U4477 , P1_U4478 , P1_U4479;
wire P1_U4480 , P1_U4481 , P1_U4482 , P1_U4483 , P1_U4484 , P1_U4485 , P1_U4486 , P1_U4487 , P1_U4488 , P1_U4489;
wire P1_U4490 , P1_U4491 , P1_U4492 , P1_U4493 , P1_U4494 , P1_U4495 , P1_U4496 , P1_U4497 , P1_U4498 , P1_U4499;
wire P1_U4500 , P1_U4501 , P1_U4502 , P1_U4503 , P1_U4504 , P1_U4505 , P1_U4506 , P1_U4507 , P1_U4508 , P1_U4509;
wire P1_U4510 , P1_U4511 , P1_U4512 , P1_U4513 , P1_U4514 , P1_U4515 , P1_U4516 , P1_U4517 , P1_U4518 , P1_U4519;
wire P1_U4520 , P1_U4521 , P1_U4522 , P1_U4523 , P1_U4524 , P1_U4525 , P1_U4526 , P1_U4527 , P1_U4528 , P1_U4529;
wire P1_U4530 , P1_U4531 , P1_U4532 , P1_U4533 , P1_U4534 , P1_U4535 , P1_U4536 , P1_U4537 , P1_U4538 , P1_U4539;
wire P1_U4540 , P1_U4541 , P1_U4542 , P1_U4543 , P1_U4544 , P1_U4545 , P1_U4546 , P1_U4547 , P1_U4548 , P1_U4549;
wire P1_U4550 , P1_U4551 , P1_U4552 , P1_U4553 , P1_U4554 , P1_U4555 , P1_U4556 , P1_U4557 , P1_U4558 , P1_U4559;
wire P1_U4560 , P1_U4561 , P1_U4562 , P1_U4563 , P1_U4564 , P1_U4565 , P1_U4566 , P1_U4567 , P1_U4568 , P1_U4569;
wire P1_U4570 , P1_U4571 , P1_U4572 , P1_U4573 , P1_U4574 , P1_U4575 , P1_U4576 , P1_U4577 , P1_U4578 , P1_U4579;
wire P1_U4580 , P1_U4581 , P1_U4582 , P1_U4583 , P1_U4584 , P1_U4585 , P1_U4586 , P1_U4587 , P1_U4588 , P1_U4589;
wire P1_U4590 , P1_U4591 , P1_U4592 , P1_U4593 , P1_U4594 , P1_U4595 , P1_U4596 , P1_U4597 , P1_U4598 , P1_U4599;
wire P1_U4600 , P1_U4601 , P1_U4602 , P1_U4603 , P1_U4604 , P1_U4605 , P1_U4606 , P1_U4607 , P1_U4608 , P1_U4609;
wire P1_U4610 , P1_U4611 , P1_U4612 , P1_U4613 , P1_U4614 , P1_U4615 , P1_U4616 , P1_U4617 , P1_U4618 , P1_U4619;
wire P1_U4620 , P1_U4621 , P1_U4622 , P1_U4623 , P1_U4624 , P1_U4625 , P1_U4626 , P1_U4627 , P1_U4628 , P1_U4629;
wire P1_U4630 , P1_U4631 , P1_U4632 , P1_U4633 , P1_U4634 , P1_U4635 , P1_U4636 , P1_U4637 , P1_U4638 , P1_U4639;
wire P1_U4640 , P1_U4641 , P1_U4642 , P1_U4643 , P1_U4644 , P1_U4645 , P1_U4646 , P1_U4647 , P1_U4648 , P1_U4649;
wire P1_U4650 , P1_U4651 , P1_U4652 , P1_U4653 , P1_U4654 , P1_U4655 , P1_U4656 , P1_U4657 , P1_U4658 , P1_U4659;
wire P1_U4660 , P1_U4661 , P1_U4662 , P1_U4663 , P1_U4664 , P1_U4665 , P1_U4666 , P1_U4667 , P1_U4668 , P1_U4669;
wire P1_U4670 , P1_U4671 , P1_U4672 , P1_U4673 , P1_U4674 , P1_U4675 , P1_U4676 , P1_U4677 , P1_U4678 , P1_U4679;
wire P1_U4680 , P1_U4681 , P1_U4682 , P1_U4683 , P1_U4684 , P1_U4685 , P1_U4686 , P1_U4687 , P1_U4688 , P1_U4689;
wire P1_U4690 , P1_U4691 , P1_U4692 , P1_U4693 , P1_U4694 , P1_U4695 , P1_U4696 , P1_U4697 , P1_U4698 , P1_U4699;
wire P1_U4700 , P1_U4701 , P1_U4702 , P1_U4703 , P1_U4704 , P1_U4705 , P1_U4706 , P1_U4707 , P1_U4708 , P1_U4709;
wire P1_U4710 , P1_U4711 , P1_U4712 , P1_U4713 , P1_U4714 , P1_U4715 , P1_U4716 , P1_U4717 , P1_U4718 , P1_U4719;
wire P1_U4720 , P1_U4721 , P1_U4722 , P1_U4723 , P1_U4724 , P1_U4725 , P1_U4726 , P1_U4727 , P1_U4728 , P1_U4729;
wire P1_U4730 , P1_U4731 , P1_U4732 , P1_U4733 , P1_U4734 , P1_U4735 , P1_U4736 , P1_U4737 , P1_U4738 , P1_U4739;
wire P1_U4740 , P1_U4741 , P1_U4742 , P1_U4743 , P1_U4744 , P1_U4745 , P1_U4746 , P1_U4747 , P1_U4748 , P1_U4749;
wire P1_U4750 , P1_U4751 , P1_U4752 , P1_U4753 , P1_U4754 , P1_U4755 , P1_U4756 , P1_U4757 , P1_U4758 , P1_U4759;
wire P1_U4760 , P1_U4761 , P1_U4762 , P1_U4763 , P1_U4764 , P1_U4765 , P1_U4766 , P1_U4767 , P1_U4768 , P1_U4769;
wire P1_U4770 , P1_U4771 , P1_U4772 , P1_U4773 , P1_U4774 , P1_U4775 , P1_U4776 , P1_U4777 , P1_U4778 , P1_U4779;
wire P1_U4780 , P1_U4781 , P1_U4782 , P1_U4783 , P1_U4784 , P1_U4785 , P1_U4786 , P1_U4787 , P1_U4788 , P1_U4789;
wire P1_U4790 , P1_U4791 , P1_U4792 , P1_U4793 , P1_U4794 , P1_U4795 , P1_U4796 , P1_U4797 , P1_U4798 , P1_U4799;
wire P1_U4800 , P1_U4801 , P1_U4802 , P1_U4803 , P1_U4804 , P1_U4805 , P1_U4806 , P1_U4807 , P1_U4808 , P1_U4809;
wire P1_U4810 , P1_U4811 , P1_U4812 , P1_U4813 , P1_U4814 , P1_U4815 , P1_U4816 , P1_U4817 , P1_U4818 , P1_U4819;
wire P1_U4820 , P1_U4821 , P1_U4822 , P1_U4823 , P1_U4824 , P1_U4825 , P1_U4826 , P1_U4827 , P1_U4828 , P1_U4829;
wire P1_U4830 , P1_U4831 , P1_U4832 , P1_U4833 , P1_U4834 , P1_U4835 , P1_U4836 , P1_U4837 , P1_U4838 , P1_U4839;
wire P1_U4840 , P1_U4841 , P1_U4842 , P1_U4843 , P1_U4844 , P1_U4845 , P1_U4846 , P1_U4847 , P1_U4848 , P1_U4849;
wire P1_U4850 , P1_U4851 , P1_U4852 , P1_U4853 , P1_U4854 , P1_U4855 , P1_U4856 , P1_U4857 , P1_U4858 , P1_U4859;
wire P1_U4860 , P1_U4861 , P1_U4862 , P1_U4863 , P1_U4864 , P1_U4865 , P1_U4866 , P1_U4867 , P1_U4868 , P1_U4869;
wire P1_U4870 , P1_U4871 , P1_U4872 , P1_U4873 , P1_U4874 , P1_U4875 , P1_U4876 , P1_U4877 , P1_U4878 , P1_U4879;
wire P1_U4880 , P1_U4881 , P1_U4882 , P1_U4883 , P1_U4884 , P1_U4885 , P1_U4886 , P1_U4887 , P1_U4888 , P1_U4889;
wire P1_U4890 , P1_U4891 , P1_U4892 , P1_U4893 , P1_U4894 , P1_U4895 , P1_U4896 , P1_U4897 , P1_U4898 , P1_U4899;
wire P1_U4900 , P1_U4901 , P1_U4902 , P1_U4903 , P1_U4904 , P1_U4905 , P1_U4906 , P1_U4907 , P1_U4908 , P1_U4909;
wire P1_U4910 , P1_U4911 , P1_U4912 , P1_U4913 , P1_U4914 , P1_U4915 , P1_U4916 , P1_U4917 , P1_U4918 , P1_U4919;
wire P1_U4920 , P1_U4921 , P1_U4922 , P1_U4923 , P1_U4924 , P1_U4925 , P1_U4926 , P1_U4927 , P1_U4928 , P1_U4929;
wire P1_U4930 , P1_U4931 , P1_U4932 , P1_U4933 , P1_U4934 , P1_U4935 , P1_U4936 , P1_U4937 , P1_U4938 , P1_U4939;
wire P1_U4940 , P1_U4941 , P1_U4942 , P1_U4943 , P1_U4944 , P1_U4945 , P1_U4946 , P1_U4947 , P1_U4948 , P1_U4949;
wire P1_U4950 , P1_U4951 , P1_U4952 , P1_U4953 , P1_U4954 , P1_U4955 , P1_U4956 , P1_U4957 , P1_U4958 , P1_U4959;
wire P1_U4960 , P1_U4961 , P1_U4962 , P1_U4963 , P1_U4964 , P1_U4965 , P1_U4966 , P1_U4967 , P1_U4968 , P1_U4969;
wire P1_U4970 , P1_U4971 , P1_U4972 , P1_U4973 , P1_U4974 , P1_U4975 , P1_U4976 , P1_U4977 , P1_U4978 , P1_U4979;
wire P1_U4980 , P1_U4981 , P1_U4982 , P1_U4983 , P1_U4984 , P1_U4985 , P1_U4986 , P1_U4987 , P1_U4988 , P1_U4989;
wire P1_U4990 , P1_U4991 , P1_U4992 , P1_U4993 , P1_U4994 , P1_U4995 , P1_U4996 , P1_U4997 , P1_U4998 , P1_U4999;
wire P1_U5000 , P1_U5001 , P1_U5002 , P1_U5003 , P1_U5004 , P1_U5005 , P1_U5006 , P1_U5007 , P1_U5008 , P1_U5009;
wire P1_U5010 , P1_U5011 , P1_U5012 , P1_U5013 , P1_U5014 , P1_U5015 , P1_U5016 , P1_U5017 , P1_U5018 , P1_U5019;
wire P1_U5020 , P1_U5021 , P1_U5022 , P1_U5023 , P1_U5024 , P1_U5025 , P1_U5026 , P1_U5027 , P1_U5028 , P1_U5029;
wire P1_U5030 , P1_U5031 , P1_U5032 , P1_U5033 , P1_U5034 , P1_U5035 , P1_U5036 , P1_U5037 , P1_U5038 , P1_U5039;
wire P1_U5040 , P1_U5041 , P1_U5042 , P1_U5043 , P1_U5044 , P1_U5045 , P1_U5046 , P1_U5047 , P1_U5048 , P1_U5049;
wire P1_U5050 , P1_U5051 , P1_U5052 , P1_U5053 , P1_U5054 , P1_U5055 , P1_U5056 , P1_U5057 , P1_U5058 , P1_U5059;
wire P1_U5060 , P1_U5061 , P1_U5062 , P1_U5063 , P1_U5064 , P1_U5065 , P1_U5066 , P1_U5067 , P1_U5068 , P1_U5069;
wire P1_U5070 , P1_U5071 , P1_U5072 , P1_U5073 , P1_U5074 , P1_U5075 , P1_U5076 , P1_U5077 , P1_U5078 , P1_U5079;
wire P1_U5080 , P1_U5081 , P1_U5082 , P1_U5083 , P1_U5084 , P1_U5085 , P1_U5086 , P1_U5087 , P1_U5088 , P1_U5089;
wire P1_U5090 , P1_U5091 , P1_U5092 , P1_U5093 , P1_U5094 , P1_U5095 , P1_U5096 , P1_U5097 , P1_U5098 , P1_U5099;
wire P1_U5100 , P1_U5101 , P1_U5102 , P1_U5103 , P1_U5104 , P1_U5105 , P1_U5106 , P1_U5107 , P1_U5108 , P1_U5109;
wire P1_U5110 , P1_U5111 , P1_U5112 , P1_U5113 , P1_U5114 , P1_U5115 , P1_U5116 , P1_U5117 , P1_U5118 , P1_U5119;
wire P1_U5120 , P1_U5121 , P1_U5122 , P1_U5123 , P1_U5124 , P1_U5125 , P1_U5126 , P1_U5127 , P1_U5128 , P1_U5129;
wire P1_U5130 , P1_U5131 , P1_U5132 , P1_U5133 , P1_U5134 , P1_U5135 , P1_U5136 , P1_U5137 , P1_U5138 , P1_U5139;
wire P1_U5140 , P1_U5141 , P1_U5142 , P1_U5143 , P1_U5144 , P1_U5145 , P1_U5146 , P1_U5147 , P1_U5148 , P1_U5149;
wire P1_U5150 , P1_U5151 , P1_U5152 , P1_U5153 , P1_U5154 , P1_U5155 , P1_U5156 , P1_U5157 , P1_U5158 , P1_U5159;
wire P1_U5160 , P1_U5161 , P1_U5162 , P1_U5163 , P1_U5164 , P1_U5165 , P1_U5166 , P1_U5167 , P1_U5168 , P1_U5169;
wire P1_U5170 , P1_U5171 , P1_U5172 , P1_U5173 , P1_U5174 , P1_U5175 , P1_U5176 , P1_U5177 , P1_U5178 , P1_U5179;
wire P1_U5180 , P1_U5181 , P1_U5182 , P1_U5183 , P1_U5184 , P1_U5185 , P1_U5186 , P1_U5187 , P1_U5188 , P1_U5189;
wire P1_U5190 , P1_U5191 , P1_U5192 , P1_U5193 , P1_U5194 , P1_U5195 , P1_U5196 , P1_U5197 , P1_U5198 , P1_U5199;
wire P1_U5200 , P1_U5201 , P1_U5202 , P1_U5203 , P1_U5204 , P1_U5205 , P1_U5206 , P1_U5207 , P1_U5208 , P1_U5209;
wire P1_U5210 , P1_U5211 , P1_U5212 , P1_U5213 , P1_U5214 , P1_U5215 , P1_U5216 , P1_U5217 , P1_U5218 , P1_U5219;
wire P1_U5220 , P1_U5221 , P1_U5222 , P1_U5223 , P1_U5224 , P1_U5225 , P1_U5226 , P1_U5227 , P1_U5228 , P1_U5229;
wire P1_U5230 , P1_U5231 , P1_U5232 , P1_U5233 , P1_U5234 , P1_U5235 , P1_U5236 , P1_U5237 , P1_U5238 , P1_U5239;
wire P1_U5240 , P1_U5241 , P1_U5242 , P1_U5243 , P1_U5244 , P1_U5245 , P1_U5246 , P1_U5247 , P1_U5248 , P1_U5249;
wire P1_U5250 , P1_U5251 , P1_U5252 , P1_U5253 , P1_U5254 , P1_U5255 , P1_U5256 , P1_U5257 , P1_U5258 , P1_U5259;
wire P1_U5260 , P1_U5261 , P1_U5262 , P1_U5263 , P1_U5264 , P1_U5265 , P1_U5266 , P1_U5267 , P1_U5268 , P1_U5269;
wire P1_U5270 , P1_U5271 , P1_U5272 , P1_U5273 , P1_U5274 , P1_U5275 , P1_U5276 , P1_U5277 , P1_U5278 , P1_U5279;
wire P1_U5280 , P1_U5281 , P1_U5282 , P1_U5283 , P1_U5284 , P1_U5285 , P1_U5286 , P1_U5287 , P1_U5288 , P1_U5289;
wire P1_U5290 , P1_U5291 , P1_U5292 , P1_U5293 , P1_U5294 , P1_U5295 , P1_U5296 , P1_U5297 , P1_U5298 , P1_U5299;
wire P1_U5300 , P1_U5301 , P1_U5302 , P1_U5303 , P1_U5304 , P1_U5305 , P1_U5306 , P1_U5307 , P1_U5308 , P1_U5309;
wire P1_U5310 , P1_U5311 , P1_U5312 , P1_U5313 , P1_U5314 , P1_U5315 , P1_U5316 , P1_U5317 , P1_U5318 , P1_U5319;
wire P1_U5320 , P1_U5321 , P1_U5322 , P1_U5323 , P1_U5324 , P1_U5325 , P1_U5326 , P1_U5327 , P1_U5328 , P1_U5329;
wire P1_U5330 , P1_U5331 , P1_U5332 , P1_U5333 , P1_U5334 , P1_U5335 , P1_U5336 , P1_U5337 , P1_U5338 , P1_U5339;
wire P1_U5340 , P1_U5341 , P1_U5342 , P1_U5343 , P1_U5344 , P1_U5345 , P1_U5346 , P1_U5347 , P1_U5348 , P1_U5349;
wire P1_U5350 , P1_U5351 , P1_U5352 , P1_U5353 , P1_U5354 , P1_U5355 , P1_U5356 , P1_U5357 , P1_U5358 , P1_U5359;
wire P1_U5360 , P1_U5361 , P1_U5362 , P1_U5363 , P1_U5364 , P1_U5365 , P1_U5366 , P1_U5367 , P1_U5368 , P1_U5369;
wire P1_U5370 , P1_U5371 , P1_U5372 , P1_U5373 , P1_U5374 , P1_U5375 , P1_U5376 , P1_U5377 , P1_U5378 , P1_U5379;
wire P1_U5380 , P1_U5381 , P1_U5382 , P1_U5383 , P1_U5384 , P1_U5385 , P1_U5386 , P1_U5387 , P1_U5388 , P1_U5389;
wire P1_U5390 , P1_U5391 , P1_U5392 , P1_U5393 , P1_U5394 , P1_U5395 , P1_U5396 , P1_U5397 , P1_U5398 , P1_U5399;
wire P1_U5400 , P1_U5401 , P1_U5402 , P1_U5403 , P1_U5404 , P1_U5405 , P1_U5406 , P1_U5407 , P1_U5408 , P1_U5409;
wire P1_U5410 , P1_U5411 , P1_U5412 , P1_U5413 , P1_U5414 , P1_U5415 , P1_U5416 , P1_U5417 , P1_U5418 , P1_U5419;
wire P1_U5420 , P1_U5421 , P1_U5422 , P1_U5423 , P1_U5424 , P1_U5425 , P1_U5426 , P1_U5427 , P1_U5428 , P1_U5429;
wire P1_U5430 , P1_U5431 , P1_U5432 , P1_U5433 , P1_U5434 , P1_U5435 , P1_U5436 , P1_U5437 , P1_U5438 , P1_U5439;
wire P1_U5440 , P1_U5441 , P1_U5442 , P1_U5443 , P1_U5444 , P1_U5445 , P1_U5446 , P1_U5447 , P1_U5448 , P1_U5449;
wire P1_U5450 , P1_U5451 , P1_U5452 , P1_U5453 , P1_U5454 , P1_U5455 , P1_U5456 , P1_U5457 , P1_U5458 , P1_U5459;
wire P1_U5460 , P1_U5461 , P1_U5462 , P1_U5463 , P1_U5464 , P1_U5465 , P1_U5466 , P1_U5467 , P1_U5468 , P1_U5469;
wire P1_U5470 , P1_U5471 , P1_U5472 , P1_U5473 , P1_U5474 , P1_U5475 , P1_U5476 , P1_U5477 , P1_U5478 , P1_U5479;
wire P1_U5480 , P1_U5481 , P1_U5482 , P1_U5483 , P1_U5484 , P1_U5485 , P1_U5486 , P1_U5487 , P1_U5488 , P1_U5489;
wire P1_U5490 , P1_U5491 , P1_U5492 , P1_U5493 , P1_U5494 , P1_U5495 , P1_U5496 , P1_U5497 , P1_U5498 , P1_U5499;
wire P1_U5500 , P1_U5501 , P1_U5502 , P1_U5503 , P1_U5504 , P1_U5505 , P1_U5506 , P1_U5507 , P1_U5508 , P1_U5509;
wire P1_U5510 , P1_U5511 , P1_U5512 , P1_U5513 , P1_U5514 , P1_U5515 , P1_U5516 , P1_U5517 , P1_U5518 , P1_U5519;
wire P1_U5520 , P1_U5521 , P1_U5522 , P1_U5523 , P1_U5524 , P1_U5525 , P1_U5526 , P1_U5527 , P1_U5528 , P1_U5529;
wire P1_U5530 , P1_U5531 , P1_U5532 , P1_U5533 , P1_U5534 , P1_U5535 , P1_U5536 , P1_U5537 , P1_U5538 , P1_U5539;
wire P1_U5540 , P1_U5541 , P1_U5542 , P1_U5543 , P1_U5544 , P1_U5545 , P1_U5546 , P1_U5547 , P1_U5548 , P1_U5549;
wire P1_U5550 , P1_U5551 , P1_U5552 , P1_U5553 , P1_U5554 , P1_U5555 , P1_U5556 , P1_U5557 , P1_U5558 , P1_U5559;
wire P1_U5560 , P1_U5561 , P1_U5562 , P1_U5563 , P1_U5564 , P1_U5565 , P1_U5566 , P1_U5567 , P1_U5568 , P1_U5569;
wire P1_U5570 , P1_U5571 , P1_U5572 , P1_U5573 , P1_U5574 , P1_U5575 , P1_U5576 , P1_U5577 , P1_U5578 , P1_U5579;
wire P1_U5580 , P1_U5581 , P1_U5582 , P1_U5583 , P1_U5584 , P1_U5585 , P1_U5586 , P1_U5587 , P1_U5588 , P1_U5589;
wire P1_U5590 , P1_U5591 , P1_U5592 , P1_U5593 , P1_U5594 , P1_U5595 , P1_U5596 , P1_U5597 , P1_U5598 , P1_U5599;
wire P1_U5600 , P1_U5601 , P1_U5602 , P1_U5603 , P1_U5604 , P1_U5605 , P1_U5606 , P1_U5607 , P1_U5608 , P1_U5609;
wire P1_U5610 , P1_U5611 , P1_U5612 , P1_U5613 , P1_U5614 , P1_U5615 , P1_U5616 , P1_U5617 , P1_U5618 , P1_U5619;
wire P1_U5620 , P1_U5621 , P1_U5622 , P1_U5623 , P1_U5624 , P1_U5625 , P1_U5626 , P1_U5627 , P1_U5628 , P1_U5629;
wire P1_U5630 , P1_U5631 , P1_U5632 , P1_U5633 , P1_U5634 , P1_U5635 , P1_U5636 , P1_U5637 , P1_U5638 , P1_U5639;
wire P1_U5640 , P1_U5641 , P1_U5642 , P1_U5643 , P1_U5644 , P1_U5645 , P1_U5646 , P1_U5647 , P1_U5648 , P1_U5649;
wire P1_U5650 , P1_U5651 , P1_U5652 , P1_U5653 , P1_U5654 , P1_U5655 , P1_U5656 , P1_U5657 , P1_U5658 , P1_U5659;
wire P1_U5660 , P1_U5661 , P1_U5662 , P1_U5663 , P1_U5664 , P1_U5665 , P1_U5666 , P1_U5667 , P1_U5668 , P1_U5669;
wire P1_U5670 , P1_U5671 , P1_U5672 , P1_U5673 , P1_U5674 , P1_U5675 , P1_U5676 , P1_U5677 , P1_U5678 , P1_U5679;
wire P1_U5680 , P1_U5681 , P1_U5682 , P1_U5683 , P1_U5684 , P1_U5685 , P1_U5686 , P1_U5687 , P1_U5688 , P1_U5689;
wire P1_U5690 , P1_U5691 , P1_U5692 , P1_U5693 , P1_U5694 , P1_U5695 , P1_U5696 , P1_U5697 , P1_U5698 , P1_U5699;
wire P1_U5700 , P1_U5701 , P1_U5702 , P1_U5703 , P1_U5704 , P1_U5705 , P1_U5706 , P1_U5707 , P1_U5708 , P1_U5709;
wire P1_U5710 , P1_U5711 , P1_U5712 , P1_U5713 , P1_U5714 , P1_U5715 , P1_U5716 , P1_U5717 , P1_U5718 , P1_U5719;
wire P1_U5720 , P1_U5721 , P1_U5722 , P1_U5723 , P1_U5724 , P1_U5725 , P1_U5726 , P1_U5727 , P1_U5728 , P1_U5729;
wire P1_U5730 , P1_U5731 , P1_U5732 , P1_U5733 , P1_U5734 , P1_U5735 , P1_U5736 , P1_U5737 , P1_U5738 , P1_U5739;
wire P1_U5740 , P1_U5741 , P1_U5742 , P1_U5743 , P1_U5744 , P1_U5745 , P1_U5746 , P1_U5747 , P1_U5748 , P1_U5749;
wire P1_U5750 , P1_U5751 , P1_U5752 , P1_U5753 , P1_U5754 , P1_U5755 , P1_U5756 , P1_U5757 , P1_U5758 , P1_U5759;
wire P1_U5760 , P1_U5761 , P1_U5762 , P1_U5763 , P1_U5764 , P1_U5765 , P1_U5766 , P1_U5767 , P1_U5768 , P1_U5769;
wire P1_U5770 , P1_U5771 , P1_U5772 , P1_U5773 , P1_U5774 , P1_U5775 , P1_U5776 , P1_U5777 , P1_U5778 , P1_U5779;
wire P1_U5780 , P1_U5781 , P1_U5782 , P1_U5783 , P1_U5784 , P1_U5785 , P1_U5786 , P1_U5787 , P1_U5788 , P1_U5789;
wire P1_U5790 , P1_U5791 , P1_U5792 , P1_U5793 , P1_U5794 , P1_U5795 , P1_U5796 , P1_U5797 , P1_U5798 , P1_U5799;
wire P1_U5800 , P1_U5801 , P1_U5802 , P1_U5803 , P1_U5804 , P1_U5805 , P1_U5806 , P1_U5807 , P1_U5808 , P1_U5809;
wire P1_U5810 , P1_U5811 , P1_U5812 , P1_U5813 , P1_U5814 , P1_U5815 , P1_U5816 , P1_U5817 , P1_U5818 , P1_U5819;
wire P1_U5820 , P1_U5821 , P1_U5822 , P1_U5823 , P1_U5824 , P1_U5825 , P1_U5826 , P1_U5827 , P1_U5828 , P1_U5829;
wire P1_U5830 , P1_U5831 , P1_U5832 , P1_U5833 , P1_U5834 , P1_U5835 , P1_U5836 , P1_U5837 , P1_U5838 , P1_U5839;
wire P1_U5840 , P1_U5841 , P1_U5842 , P1_U5843 , P1_U5844 , P1_U5845 , P1_U5846 , P1_U5847 , P1_U5848 , P1_U5849;
wire P1_U5850 , P1_U5851 , P1_U5852 , P1_U5853 , P1_U5854 , P1_U5855 , P1_U5856 , P1_U5857 , P1_U5858 , P1_U5859;
wire P1_U5860 , P1_U5861 , P1_U5862 , P1_U5863 , P1_U5864 , P1_U5865 , P1_U5866 , P1_U5867 , P1_U5868 , P1_U5869;
wire P1_U5870 , P1_U5871 , P1_U5872 , P1_U5873 , P1_U5874 , P1_U5875 , P1_U5876 , P1_U5877 , P1_U5878 , P1_U5879;
wire P1_U5880 , P1_U5881 , P1_U5882 , P1_U5883 , P1_U5884 , P1_U5885 , P1_U5886 , P1_U5887 , P1_U5888 , P1_U5889;
wire P1_U5890 , P1_U5891 , P1_U5892 , P1_U5893 , P1_U5894 , P1_U5895 , P1_U5896 , P1_U5897 , P1_U5898 , P1_U5899;
wire P1_U5900 , P1_U5901 , P1_U5902 , P1_U5903 , P1_U5904 , P1_U5905 , P1_U5906 , P1_U5907 , P1_U5908 , P1_U5909;
wire P1_U5910 , P1_U5911 , P1_U5912 , P1_U5913 , P1_U5914 , P1_U5915 , P1_U5916 , P1_U5917 , P1_U5918 , P1_U5919;
wire P1_U5920 , P1_U5921 , P1_U5922 , P1_U5923 , P1_U5924 , P1_U5925 , P1_U5926 , P1_U5927 , P1_U5928 , P1_U5929;
wire P1_U5930 , P1_U5931 , P1_U5932 , P1_U5933 , P1_U5934 , P1_U5935 , P1_U5936 , P1_U5937 , P1_U5938 , P1_U5939;
wire P1_U5940 , P1_U5941 , P1_U5942 , P1_U5943 , P1_U5944 , P1_U5945 , P1_U5946 , P1_U5947 , P1_U5948 , P1_U5949;
wire P1_U5950 , P1_U5951 , P1_U5952 , P1_U5953 , P1_U5954 , P1_U5955 , P1_U5956 , P1_U5957 , P1_U5958 , P1_U5959;
wire P1_U5960 , P1_U5961 , P1_U5962 , P1_U5963 , P1_U5964 , P1_U5965 , P1_U5966 , P1_U5967 , P1_U5968 , P1_U5969;
wire P1_U5970 , P1_U5971 , P1_U5972 , P1_U5973 , P1_U5974 , P1_U5975 , P1_U5976 , P1_U5977 , P1_U5978 , P1_U5979;
wire P1_U5980 , P1_U5981 , P1_U5982 , P1_U5983 , P1_U5984 , P1_U5985 , P1_U5986 , P1_U5987 , P1_U5988 , P1_U5989;
wire P1_U5990 , P1_U5991 , P1_U5992 , P1_U5993 , P1_U5994 , P1_U5995 , P1_U5996 , P1_U5997 , P1_U5998 , P1_U5999;
wire P1_U6000 , P1_U6001 , P1_U6002 , P1_U6003 , P1_U6004 , P1_U6005 , P1_U6006 , P1_U6007 , P1_U6008 , P1_U6009;
wire P1_U6010 , P1_U6011 , P1_U6012 , P1_U6013 , P1_U6014 , P1_U6015 , P1_U6016 , P1_U6017 , P1_U6018 , P1_U6019;
wire P1_U6020 , P1_U6021 , P1_U6022 , P1_U6023 , P1_U6024 , P1_U6025 , P1_U6026 , P1_U6027 , P1_U6028 , P1_U6029;
wire P1_U6030 , P1_U6031 , P1_U6032 , P1_U6033 , P1_U6034 , P1_U6035 , P1_U6036 , P1_U6037 , P1_U6038 , P1_U6039;
wire P1_U6040 , P1_U6041 , P1_U6042 , P1_U6043 , P1_U6044 , P1_U6045 , P1_U6046 , P1_U6047 , P1_U6048 , P1_U6049;
wire P1_U6050 , P1_U6051 , P1_U6052 , P1_U6053 , P1_U6054 , P1_U6055 , P1_U6056 , P1_U6057 , P1_U6058 , P1_U6059;
wire P1_U6060 , P1_U6061 , P1_U6062 , P1_U6063 , P1_U6064 , P1_U6065 , P1_U6066 , P1_U6067 , P1_U6068 , P1_U6069;
wire P1_U6070 , P1_U6071 , P1_U6072 , P1_U6073 , P1_U6074 , P1_U6075 , P1_U6076 , P1_U6077 , P1_U6078 , P1_U6079;
wire P1_U6080 , P1_U6081 , P1_U6082 , P1_U6083 , P1_U6084 , P1_U6085 , P1_U6086 , P1_U6087 , P1_U6088 , P1_U6089;
wire P1_U6090 , P1_U6091 , P1_U6092 , P1_U6093 , P1_U6094 , P1_U6095 , P1_U6096 , P1_U6097 , P1_U6098 , P1_U6099;
wire P1_U6100 , P1_U6101 , P1_U6102 , P1_U6103 , P1_U6104 , P1_U6105 , P1_U6106 , P1_U6107 , P1_U6108 , P1_U6109;
wire P1_U6110 , P1_U6111 , P1_U6112 , P1_U6113 , P1_U6114 , P1_U6115 , P1_U6116 , P1_U6117 , P1_U6118 , P1_U6119;
wire P1_U6120 , P1_U6121 , P1_U6122 , P1_U6123 , P1_U6124 , P1_U6125 , P1_U6126 , P1_U6127 , P1_U6128 , P1_U6129;
wire P1_U6130 , P1_U6131 , P1_U6132 , P1_U6133 , P1_U6134 , P1_U6135 , P1_U6136 , P1_U6137 , P1_U6138 , P1_U6139;
wire P1_U6140 , P1_U6141 , P1_U6142 , P1_U6143 , P1_U6144 , P1_U6145 , P1_U6146 , P1_U6147 , P1_U6148 , P1_U6149;
wire P1_U6150 , P1_U6151 , P1_U6152 , P1_U6153 , P1_U6154 , P1_U6155 , P1_U6156 , P1_U6157 , P1_U6158 , P1_U6159;
wire P1_U6160 , P1_U6161 , P1_U6162 , P1_U6163 , P1_U6164 , P1_U6165 , P1_U6166 , P1_U6167 , P1_U6168 , P1_U6169;
wire P1_U6170 , P1_U6171 , P1_U6172 , P1_U6173 , P1_U6174 , P1_U6175 , P1_U6176 , P1_U6177 , P1_U6178 , P1_U6179;
wire P1_U6180 , P1_U6181 , P1_U6182 , P1_U6183 , P1_U6184 , P1_U6185 , P1_U6186 , P1_U6187 , P1_U6188 , P1_U6189;
wire P1_U6190 , P1_U6191 , P1_U6192 , P1_U6193 , P1_U6194 , P1_U6195 , P1_U6196 , P1_U6197 , P1_U6198 , P1_U6199;
wire P1_U6200 , P1_U6201 , P1_U6202 , P1_U6203 , P1_U6204 , P1_U6205 , P1_U6206 , P1_U6207 , P1_U6208 , P1_U6209;
wire P1_U6210 , P1_U6211 , P1_U6212 , P1_U6213 , P1_U6214 , P1_U6215 , P1_U6216 , P1_U6217 , P1_U6218 , P1_U6219;
wire P1_U6220 , P1_U6221 , P1_U6222 , P1_U6223 , P1_U6224 , P1_U6225 , P1_U6226 , P1_U6227 , P1_U6228 , P1_U6229;
wire P1_U6230 , P1_U6231 , P1_U6232 , P1_U6233 , P1_U6234 , P1_U6235 , P1_U6236 , P1_U6237 , P1_U6238 , P1_U6239;
wire P1_U6240 , P1_U6241 , P1_U6242 , P1_U6243 , P1_U6244 , P1_U6245 , P1_U6246 , P1_U6247 , P1_U6248 , P1_U6249;
wire P1_U6250 , P1_U6251 , P1_U6252 , P1_U6253 , P1_U6254 , P1_U6255 , P1_U6256 , P1_U6257 , P1_U6258 , P1_U6259;
wire P1_U6260 , P1_U6261 , P1_U6262 , P1_U6263 , P1_U6264 , P1_U6265 , P1_U6266 , P1_U6267 , P1_U6268 , P1_U6269;
wire P1_U6270 , P1_U6271 , P1_U6272 , P1_U6273 , P1_U6274 , P1_U6275 , P1_U6276 , P1_U6277 , P1_U6278 , P1_U6279;
wire P1_U6280 , P1_U6281 , P1_U6282 , P1_U6283 , P1_U6284 , P1_U6285 , P1_U6286 , P1_U6287 , P1_U6288 , P1_U6289;
wire P1_U6290 , P1_U6291 , P1_U6292 , P1_U6293 , P1_U6294 , P1_U6295 , P1_U6296 , P1_U6297 , P1_U6298 , P1_U6299;
wire P1_U6300 , P1_U6301 , P1_U6302 , P1_U6303 , P1_U6304 , P1_U6305 , P1_U6306 , P1_U6307 , P1_U6308 , P1_U6309;
wire P1_U6310 , P1_U6311 , P1_U6312 , P1_U6313 , P1_U6314 , P1_U6315 , P1_U6316 , P1_U6317 , P1_U6318 , P1_U6319;
wire P1_U6320 , P1_U6321 , P1_U6322 , P1_U6323 , P1_U6324 , P1_U6325 , P1_U6326 , P1_U6327 , P1_U6328 , P1_U6329;
wire P1_U6330 , P1_U6331 , P1_U6332 , P1_U6333 , P1_U6334 , P1_U6335 , P1_U6336 , P1_U6337 , P1_U6338 , P1_U6339;
wire P1_U6340 , P1_U6341 , P1_U6342 , P1_U6343 , P1_U6344 , P1_U6345 , P1_U6346 , P1_U6347 , P1_U6348 , P1_U6349;
wire P1_U6350 , P1_U6351 , P1_U6352 , P1_U6353 , P1_U6354 , P1_U6355 , P1_U6356 , P1_U6357 , P1_U6358 , P1_U6359;
wire P1_U6360 , P1_U6361 , P1_U6362 , P1_U6363 , P1_U6364 , P1_U6365 , P1_U6366 , P1_U6367 , P1_U6368 , P1_U6369;
wire P1_U6370 , P1_U6371 , P1_U6372 , P1_U6373 , P1_U6374 , P1_U6375 , P1_U6376 , P1_U6377 , P1_U6378 , P1_U6379;
wire P1_U6380 , P1_U6381 , P1_U6382 , P1_U6383 , P1_U6384 , P1_U6385 , P1_U6386 , P1_U6387 , P1_U6388 , P1_U6389;
wire P1_U6390 , P1_U6391 , P1_U6392 , P1_U6393 , P1_U6394 , P1_U6395 , P1_U6396 , P1_U6397 , P1_U6398 , P1_U6399;
wire P1_U6400 , P1_U6401 , P1_U6402 , P1_U6403 , P1_U6404 , P1_U6405 , P1_U6406 , P1_U6407 , P1_U6408 , P1_U6409;
wire P1_U6410 , P1_U6411 , P1_U6412 , P1_U6413 , P1_U6414 , P1_U6415 , P1_U6416 , P1_U6417 , P1_U6418 , P1_U6419;
wire P1_U6420 , P1_U6421 , P1_U6422 , P1_U6423 , P1_U6424 , P1_U6425 , P1_U6426 , P1_U6427 , P1_U6428 , P1_U6429;
wire P1_U6430 , P1_U6431 , P1_U6432 , P1_U6433 , P1_U6434 , P1_U6435 , P1_U6436 , P1_U6437 , P1_U6438 , P1_U6439;
wire P1_U6440 , P1_U6441 , P1_U6442 , P1_U6443 , P1_U6444 , P1_U6445 , P1_U6446 , P1_U6447 , P1_U6448 , P1_U6449;
wire P1_U6450 , P1_U6451 , P1_U6452 , P1_U6453 , P1_U6454 , P1_U6455 , P1_U6456 , P1_U6457 , P1_U6458 , P1_U6459;
wire P1_U6460 , P1_U6461 , P1_U6462 , P1_U6463 , P1_U6464 , P1_U6465 , P1_U6466 , P1_U6467 , P1_U6468 , P1_U6469;
wire P1_U6470 , P1_U6471 , P1_U6472 , P1_U6473 , P1_U6474 , P1_U6475 , P1_U6476 , P1_U6477 , P1_U6478 , P1_U6479;
wire P1_U6480 , P1_U6481 , P1_U6482 , P1_U6483 , P1_U6484 , P1_U6485 , P1_U6486 , P1_U6487 , P1_U6488 , P1_U6489;
wire P1_U6490 , P1_U6491 , P1_U6492 , P1_U6493 , P1_U6494 , P1_U6495 , P1_U6496 , P1_U6497 , P1_U6498 , P1_U6499;
wire P1_U6500 , P1_U6501 , P1_U6502 , P1_U6503 , P1_U6504 , P1_U6505 , P1_U6506 , P1_U6507 , P1_U6508 , P1_U6509;
wire P1_U6510 , P1_U6511 , P1_U6512 , P1_U6513 , P1_U6514 , P1_U6515 , P1_U6516 , P1_U6517 , P1_U6518 , P1_U6519;
wire P1_U6520 , P1_U6521 , P1_U6522 , P1_U6523 , P1_U6524 , P1_U6525 , P1_U6526 , P1_U6527 , P1_U6528 , P1_U6529;
wire P1_U6530 , P1_U6531 , P1_U6532 , P1_U6533 , P1_U6534 , P1_U6535 , P1_U6536 , P1_U6537 , P1_U6538 , P1_U6539;
wire P1_U6540 , P1_U6541 , P1_U6542 , P1_U6543 , P1_U6544 , P1_U6545 , P1_U6546 , P1_U6547 , P1_U6548 , P1_U6549;
wire P1_U6550 , P1_U6551 , P1_U6552 , P1_U6553 , P1_U6554 , P1_U6555 , P1_U6556 , P1_U6557 , P1_U6558 , P1_U6559;
wire P1_U6560 , P1_U6561 , P1_U6562 , P1_U6563 , P1_U6564 , P1_U6565 , P1_U6566 , P1_U6567 , P1_U6568 , P1_U6569;
wire P1_U6570 , P1_U6571 , P1_U6572 , P1_U6573 , P1_U6574 , P1_U6575 , P1_U6576 , P1_U6577 , P1_U6578 , P1_U6579;
wire P1_U6580 , P1_U6581 , P1_U6582 , P1_U6583 , P1_U6584 , P1_U6585 , P1_U6586 , P1_U6587 , P1_U6588 , P1_U6589;
wire P1_U6590 , P1_U6591 , P1_U6592 , P1_U6593 , P1_U6594 , P1_U6595 , P1_U6596 , P1_U6597 , P1_U6598 , P1_U6599;
wire P1_U6600 , P1_U6601 , P1_U6602 , P1_U6603 , P1_U6604 , P1_U6605 , P1_U6606 , P1_U6607 , P1_U6608 , P1_U6609;
wire P1_U6610 , P1_U6611 , P1_U6612 , P1_U6613 , P1_U6614 , P1_U6615 , P1_U6616 , P1_U6617 , P1_U6618 , P1_U6619;
wire P1_U6620 , P1_U6621 , P1_U6622 , P1_U6623 , P1_U6624 , P1_U6625 , P1_U6626 , P1_U6627 , P1_U6628 , P1_U6629;
wire P1_U6630 , P1_U6631 , P1_U6632 , P1_U6633 , P1_U6634 , P1_U6635 , P1_U6636 , P1_U6637 , P1_U6638 , P1_U6639;
wire P1_U6640 , P1_U6641 , P1_U6642 , P1_U6643 , P1_U6644 , P1_U6645 , P1_U6646 , P1_U6647 , P1_U6648 , P1_U6649;
wire P1_U6650 , P1_U6651 , P1_U6652 , P1_U6653 , P1_U6654 , P1_U6655 , P1_U6656 , P1_U6657 , P1_U6658 , P1_U6659;
wire P1_U6660 , P1_U6661 , P1_U6662 , P1_U6663 , P1_U6664 , P1_U6665 , P1_U6666 , P1_U6667 , P1_U6668 , P1_U6669;
wire P1_U6670 , P1_U6671 , P1_U6672 , P1_U6673 , P1_U6674 , P1_U6675 , P1_U6676 , P1_U6677 , P1_U6678 , P1_U6679;
wire P1_U6680 , P1_U6681 , P1_U6682 , P1_U6683 , P1_U6684 , P1_U6685 , P1_U6686 , P1_U6687 , P1_U6688 , P1_U6689;
wire P1_U6690 , P1_U6691 , P1_U6692 , P1_U6693 , P1_U6694 , P1_U6695 , P1_U6696 , P1_U6697 , P1_U6698 , P1_U6699;
wire P1_U6700 , P1_U6701 , P1_U6702 , P1_U6703 , P1_U6704 , P1_U6705 , P1_U6706 , P1_U6707 , P1_U6708 , P1_U6709;
wire P1_U6710 , P1_U6711 , P1_U6712 , P1_U6713 , P1_U6714 , P1_U6715 , P1_U6716 , P1_U6717 , P1_U6718 , P1_U6719;
wire P1_U6720 , P1_U6721 , P1_U6722 , P1_U6723 , P1_U6724 , P1_U6725 , P1_U6726 , P1_U6727 , P1_U6728 , P1_U6729;
wire P1_U6730 , P1_U6731 , P1_U6732 , P1_U6733 , P1_U6734 , P1_U6735 , P1_U6736 , P1_U6737 , P1_U6738 , P1_U6739;
wire P1_U6740 , P1_U6741 , P1_U6742 , P1_U6743 , P1_U6744 , P1_U6745 , P1_U6746 , P1_U6747 , P1_U6748 , P1_U6749;
wire P1_U6750 , P1_U6751 , P1_U6752 , P1_U6753 , P1_U6754 , P1_U6755 , P1_U6756 , P1_U6757 , P1_U6758 , P1_U6759;
wire P1_U6760 , P1_U6761 , P1_U6762 , P1_U6763 , P1_U6764 , P1_U6765 , P1_U6766 , P1_U6767 , P1_U6768 , P1_U6769;
wire P1_U6770 , P1_U6771 , P1_U6772 , P1_U6773 , P1_U6774 , P1_U6775 , P1_U6776 , P1_U6777 , P1_U6778 , P1_U6779;
wire P1_U6780 , P1_U6781 , P1_U6782 , P1_U6783 , P1_U6784 , P1_U6785 , P1_U6786 , P1_U6787 , P1_U6788 , P1_U6789;
wire P1_U6790 , P1_U6791 , P1_U6792 , P1_U6793 , P1_U6794 , P1_U6795 , P1_U6796 , P1_U6797 , P1_U6798 , P1_U6799;
wire P1_U6800 , P1_U6801 , P1_U6802 , P1_U6803 , P1_U6804 , P1_U6805 , P1_U6806 , P1_U6807 , P1_U6808 , P1_U6809;
wire P1_U6810 , P1_U6811 , P1_U6812 , P1_U6813 , P1_U6814 , P1_U6815 , P1_U6816 , P1_U6817 , P1_U6818 , P1_U6819;
wire P1_U6820 , P1_U6821 , P1_U6822 , P1_U6823 , P1_U6824 , P1_U6825 , P1_U6826 , P1_U6827 , P1_U6828 , P1_U6829;
wire P1_U6830 , P1_U6831 , P1_U6832 , P1_U6833 , P1_U6834 , P1_U6835 , P1_U6836 , P1_U6837 , P1_U6838 , P1_U6839;
wire P1_U6840 , P1_U6841 , P1_U6842 , P1_U6843 , P1_U6844 , P1_U6845 , P1_U6846 , P1_U6847 , P1_U6848 , P1_U6849;
wire P1_U6850 , P1_U6851 , P1_U6852 , P1_U6853 , P1_U6854 , P1_U6855 , P1_U6856 , P1_U6857 , P1_U6858 , P1_U6859;
wire P1_U6860 , P1_U6861 , P1_U6862 , P1_U6863 , P1_U6864 , P1_U6865 , P1_U6866 , P1_U6867 , P1_U6868 , P1_U6869;
wire P1_U6870 , P1_U6871 , P1_U6872 , P1_U6873 , P1_U6874 , P1_U6875 , P1_U6876 , P1_U6877 , P1_U6878 , P1_U6879;
wire P1_U6880 , P1_U6881 , P1_U6882 , P1_U6883 , P1_U6884 , P1_U6885 , P1_U6886 , P1_U6887 , P1_U6888 , P1_U6889;
wire P1_U6890 , P1_U6891 , P1_U6892 , P1_U6893 , P1_U6894 , P1_U6895 , P1_U6896 , P1_U6897 , P1_U6898 , P1_U6899;
wire P1_U6900 , P1_U6901 , P1_U6902 , P1_U6903 , P1_U6904 , P1_U6905 , P1_U6906 , P1_U6907 , P1_U6908 , P1_U6909;
wire P1_U6910 , P1_U6911 , P1_U6912 , P1_U6913 , P1_U6914 , P1_U6915 , P1_U6916 , P1_U6917 , P1_U6918 , P1_U6919;
wire P1_U6920 , P1_U6921 , P1_U6922 , P1_U6923 , P1_U6924 , P1_U6925 , P1_U6926 , P1_U6927 , P1_U6928 , P1_U6929;
wire P1_U6930 , P1_U6931 , P1_U6932 , P1_U6933 , P1_U6934 , P1_U6935 , P1_U6936 , P1_U6937 , P1_U6938 , P1_U6939;
wire P1_U6940 , P1_U6941 , P1_U6942 , P1_U6943 , P1_U6944 , P1_U6945 , P1_U6946 , P1_U6947 , P1_U6948 , P1_U6949;
wire P1_U6950 , P1_U6951 , P1_U6952 , P1_U6953 , P1_U6954 , P1_U6955 , P1_U6956 , P1_U6957 , P1_U6958 , P1_U6959;
wire P1_U6960 , P1_U6961 , P1_U6962 , P1_U6963 , P1_U6964 , P1_U6965 , P1_U6966 , P1_U6967 , P1_U6968 , P1_U6969;
wire P1_U6970 , P1_U6971 , P1_U6972 , P1_U6973 , P1_U6974 , P1_U6975 , P1_U6976 , P1_U6977 , P1_U6978 , P1_U6979;
wire P1_U6980 , P1_U6981 , P1_U6982 , P1_U6983 , P1_U6984 , P1_U6985 , P1_U6986 , P1_U6987 , P1_U6988 , P1_U6989;
wire P1_U6990 , P1_U6991 , P1_U6992 , P1_U6993 , P1_U6994 , P1_U6995 , P1_U6996 , P1_U6997 , P1_U6998 , P1_U6999;
wire P1_U7000 , P1_U7001 , P1_U7002 , P1_U7003 , P1_U7004 , P1_U7005 , P1_U7006 , P1_U7007 , P1_U7008 , P1_U7009;
wire P1_U7010 , P1_U7011 , P1_U7012 , P1_U7013 , P1_U7014 , P1_U7015 , P1_U7016 , P1_U7017 , P1_U7018 , P1_U7019;
wire P1_U7020 , P1_U7021 , P1_U7022 , P1_U7023 , P1_U7024 , P1_U7025 , P1_U7026 , P1_U7027 , P1_U7028 , P1_U7029;
wire P1_U7030 , P1_U7031 , P1_U7032 , P1_U7033 , P1_U7034 , P1_U7035 , P1_U7036 , P1_U7037 , P1_U7038 , P1_U7039;
wire P1_U7040 , P1_U7041 , P1_U7042 , P1_U7043 , P1_U7044 , P1_U7045 , P1_U7046 , P1_U7047 , P1_U7048 , P1_U7049;
wire P1_U7050 , P1_U7051 , P1_U7052 , P1_U7053 , P1_U7054 , P1_U7055 , P1_U7056 , P1_U7057 , P1_U7058 , P1_U7059;
wire P1_U7060 , P1_U7061 , P1_U7062 , P1_U7063 , P1_U7064 , P1_U7065 , P1_U7066 , P1_U7067 , P1_U7068 , P1_U7069;
wire P1_U7070 , P1_U7071 , P1_U7072 , P1_U7073 , P1_U7074 , P1_U7075 , P1_U7076 , P1_U7077 , P1_U7078 , P1_U7079;
wire P1_U7080 , P1_U7081 , P1_U7082 , P1_U7083 , P1_U7084 , P1_U7085 , P1_U7086 , P1_U7087 , P1_U7088 , P1_U7089;
wire P1_U7090 , P1_U7091 , P1_U7092 , P1_U7093 , P1_U7094 , P1_U7095 , P1_U7096 , P1_U7097 , P1_U7098 , P1_U7099;
wire P1_U7100 , P1_U7101 , P1_U7102 , P1_U7103 , P1_U7104 , P1_U7105 , P1_U7106 , P1_U7107 , P1_U7108 , P1_U7109;
wire P1_U7110 , P1_U7111 , P1_U7112 , P1_U7113 , P1_U7114 , P1_U7115 , P1_U7116 , P1_U7117 , P1_U7118 , P1_U7119;
wire P1_U7120 , P1_U7121 , P1_U7122 , P1_U7123 , P1_U7124 , P1_U7125 , P1_U7126 , P1_U7127 , P1_U7128 , P1_U7129;
wire P1_U7130 , P1_U7131 , P1_U7132 , P1_U7133 , P1_U7134 , P1_U7135 , P1_U7136 , P1_U7137 , P1_U7138 , P1_U7139;
wire P1_U7140 , P1_U7141 , P1_U7142 , P1_U7143 , P1_U7144 , P1_U7145 , P1_U7146 , P1_U7147 , P1_U7148 , P1_U7149;
wire P1_U7150 , P1_U7151 , P1_U7152 , P1_U7153 , P1_U7154 , P1_U7155 , P1_U7156 , P1_U7157 , P1_U7158 , P1_U7159;
wire P1_U7160 , P1_U7161 , P1_U7162 , P1_U7163 , P1_U7164 , P1_U7165 , P1_U7166 , P1_U7167 , P1_U7168 , P1_U7169;
wire P1_U7170 , P1_U7171 , P1_U7172 , P1_U7173 , P1_U7174 , P1_U7175 , P1_U7176 , P1_U7177 , P1_U7178 , P1_U7179;
wire P1_U7180 , P1_U7181 , P1_U7182 , P1_U7183 , P1_U7184 , P1_U7185 , P1_U7186 , P1_U7187 , P1_U7188 , P1_U7189;
wire P1_U7190 , P1_U7191 , P1_U7192 , P1_U7193 , P1_U7194 , P1_U7195 , P1_U7196 , P1_U7197 , P1_U7198 , P1_U7199;
wire P1_U7200 , P1_U7201 , P1_U7202 , P1_U7203 , P1_U7204 , P1_U7205 , P1_U7206 , P1_U7207 , P1_U7208 , P1_U7209;
wire P1_U7210 , P1_U7211 , P1_U7212 , P1_U7213 , P1_U7214 , P1_U7215 , P1_U7216 , P1_U7217 , P1_U7218 , P1_U7219;
wire P1_U7220 , P1_U7221 , P1_U7222 , P1_U7223 , P1_U7224 , P1_U7225 , P1_U7226 , P1_U7227 , P1_U7228 , P1_U7229;
wire P1_U7230 , P1_U7231 , P1_U7232 , P1_U7233 , P1_U7234 , P1_U7235 , P1_U7236 , P1_U7237 , P1_U7238 , P1_U7239;
wire P1_U7240 , P1_U7241 , P1_U7242 , P1_U7243 , P1_U7244 , P1_U7245 , P1_U7246 , P1_U7247 , P1_U7248 , P1_U7249;
wire P1_U7250 , P1_U7251 , P1_U7252 , P1_U7253 , P1_U7254 , P1_U7255 , P1_U7256 , P1_U7257 , P1_U7258 , P1_U7259;
wire P1_U7260 , P1_U7261 , P1_U7262 , P1_U7263 , P1_U7264 , P1_U7265 , P1_U7266 , P1_U7267 , P1_U7268 , P1_U7269;
wire P1_U7270 , P1_U7271 , P1_U7272 , P1_U7273 , P1_U7274 , P1_U7275 , P1_U7276 , P1_U7277 , P1_U7278 , P1_U7279;
wire P1_U7280 , P1_U7281 , P1_U7282 , P1_U7283 , P1_U7284 , P1_U7285 , P1_U7286 , P1_U7287 , P1_U7288 , P1_U7289;
wire P1_U7290 , P1_U7291 , P1_U7292 , P1_U7293 , P1_U7294 , P1_U7295 , P1_U7296 , P1_U7297 , P1_U7298 , P1_U7299;
wire P1_U7300 , P1_U7301 , P1_U7302 , P1_U7303 , P1_U7304 , P1_U7305 , P1_U7306 , P1_U7307 , P1_U7308 , P1_U7309;
wire P1_U7310 , P1_U7311 , P1_U7312 , P1_U7313 , P1_U7314 , P1_U7315 , P1_U7316 , P1_U7317 , P1_U7318 , P1_U7319;
wire P1_U7320 , P1_U7321 , P1_U7322 , P1_U7323 , P1_U7324 , P1_U7325 , P1_U7326 , P1_U7327 , P1_U7328 , P1_U7329;
wire P1_U7330 , P1_U7331 , P1_U7332 , P1_U7333 , P1_U7334 , P1_U7335 , P1_U7336 , P1_U7337 , P1_U7338 , P1_U7339;
wire P1_U7340 , P1_U7341 , P1_U7342 , P1_U7343 , P1_U7344 , P1_U7345 , P1_U7346 , P1_U7347 , P1_U7348 , P1_U7349;
wire P1_U7350 , P1_U7351 , P1_U7352 , P1_U7353 , P1_U7354 , P1_U7355 , P1_U7356 , P1_U7357 , P1_U7358 , P1_U7359;
wire P1_U7360 , P1_U7361 , P1_U7362 , P1_U7363 , P1_U7364 , P1_U7365 , P1_U7366 , P1_U7367 , P1_U7368 , P1_U7369;
wire P1_U7370 , P1_U7371 , P1_U7372 , P1_U7373 , P1_U7374 , P1_U7375 , P1_U7376 , P1_U7377 , P1_U7378 , P1_U7379;
wire P1_U7380 , P1_U7381 , P1_U7382 , P1_U7383 , P1_U7384 , P1_U7385 , P1_U7386 , P1_U7387 , P1_U7388 , P1_U7389;
wire P1_U7390 , P1_U7391 , P1_U7392 , P1_U7393 , P1_U7394 , P1_U7395 , P1_U7396 , P1_U7397 , P1_U7398 , P1_U7399;
wire P1_U7400 , P1_U7401 , P1_U7402 , P1_U7403 , P1_U7404 , P1_U7405 , P1_U7406 , P1_U7407 , P1_U7408 , P1_U7409;
wire P1_U7410 , P1_U7411 , P1_U7412 , P1_U7413 , P1_U7414 , P1_U7415 , P1_U7416 , P1_U7417 , P1_U7418 , P1_U7419;
wire P1_U7420 , P1_U7421 , P1_U7422 , P1_U7423 , P1_U7424 , P1_U7425 , P1_U7426 , P1_U7427 , P1_U7428 , P1_U7429;
wire P1_U7430 , P1_U7431 , P1_U7432 , P1_U7433 , P1_U7434 , P1_U7435 , P1_U7436 , P1_U7437 , P1_U7438 , P1_U7439;
wire P1_U7440 , P1_U7441 , P1_U7442 , P1_U7443 , P1_U7444 , P1_U7445 , P1_U7446 , P1_U7447 , P1_U7448 , P1_U7449;
wire P1_U7450 , P1_U7451 , P1_U7452 , P1_U7453 , P1_U7454 , P1_U7455 , P1_U7456 , P1_U7457 , P1_U7458 , P1_U7459;
wire P1_U7460 , P1_U7461 , P1_U7462 , P1_U7463 , P1_U7464 , P1_U7465 , P1_U7466 , P1_U7467 , P1_U7468 , P1_U7469;
wire P1_U7470 , P1_U7471 , P1_U7472 , P1_U7473 , P1_U7474 , P1_U7475 , P1_U7476 , P1_U7477 , P1_U7478 , P1_U7479;
wire P1_U7480 , P1_U7481 , P1_U7482 , P1_U7483 , P1_U7484 , P1_U7485 , P1_U7486 , P1_U7487 , P1_U7488 , P1_U7489;
wire P1_U7490 , P1_U7491 , P1_U7492 , P1_U7493 , P1_U7494 , P1_U7495 , P1_U7496 , P1_U7497 , P1_U7498 , P1_U7499;
wire P1_U7500 , P1_U7501 , P1_U7502 , P1_U7503 , P1_U7504 , P1_U7505 , P1_U7506 , P1_U7507 , P1_U7508 , P1_U7509;
wire P1_U7510 , P1_U7511 , P1_U7512 , P1_U7513 , P1_U7514 , P1_U7515 , P1_U7516 , P1_U7517 , P1_U7518 , P1_U7519;
wire P1_U7520 , P1_U7521 , P1_U7522 , P1_U7523 , P1_U7524 , P1_U7525 , P1_U7526 , P1_U7527 , P1_U7528 , P1_U7529;
wire P1_U7530 , P1_U7531 , P1_U7532 , P1_U7533 , P1_U7534 , P1_U7535 , P1_U7536 , P1_U7537 , P1_U7538 , P1_U7539;
wire P1_U7540 , P1_U7541 , P1_U7542 , P1_U7543 , P1_U7544 , P1_U7545 , P1_U7546 , P1_U7547 , P1_U7548 , P1_U7549;
wire P1_U7550 , P1_U7551 , P1_U7552 , P1_U7553 , P1_U7554 , P1_U7555 , P1_U7556 , P1_U7557 , P1_U7558 , P1_U7559;
wire P1_U7560 , P1_U7561 , P1_U7562 , P1_U7563 , P1_U7564 , P1_U7565 , P1_U7566 , P1_U7567 , P1_U7568 , P1_U7569;
wire P1_U7570 , P1_U7571 , P1_U7572 , P1_U7573 , P1_U7574 , P1_U7575 , P1_U7576 , P1_U7577 , P1_U7578 , P1_U7579;
wire P1_U7580 , P1_U7581 , P1_U7582 , P1_U7583 , P1_U7584 , P1_U7585 , P1_U7586 , P1_U7587 , P1_U7588 , P1_U7589;
wire P1_U7590 , P1_U7591 , P1_U7592 , P1_U7593 , P1_U7594 , P1_U7595 , P1_U7596 , P1_U7597 , P1_U7598 , P1_U7599;
wire P1_U7600 , P1_U7601 , P1_U7602 , P1_U7603 , P1_U7604 , P1_U7605 , P1_U7606 , P1_U7607 , P1_U7608 , P1_U7609;
wire P1_U7610 , P1_U7611 , P1_U7612 , P1_U7613 , P1_U7614 , P1_U7615 , P1_U7616 , P1_U7617 , P1_U7618 , P1_U7619;
wire P1_U7620 , P1_U7621 , P1_U7622 , P1_U7623 , P1_U7624 , P1_U7625 , P1_U7626 , P1_U7627 , P1_U7628 , P1_U7629;
wire P1_U7630 , P1_U7631 , P1_U7632 , P1_U7633 , P1_U7634 , P1_U7635 , P1_U7636 , P1_U7637 , P1_U7638 , P1_U7639;
wire P1_U7640 , P1_U7641 , P1_U7642 , P1_U7643 , P1_U7644 , P1_U7645 , P1_U7646 , P1_U7647 , P1_U7648 , P1_U7649;
wire P1_U7650 , P1_U7651 , P1_U7652 , P1_U7653 , P1_U7654 , P1_U7655 , P1_U7656 , P1_U7657 , P1_U7658 , P1_U7659;
wire P1_U7660 , P1_U7661 , P1_U7662 , P1_U7663 , P1_U7664 , P1_U7665 , P1_U7666 , P1_U7667 , P1_U7668 , P1_U7669;
wire P1_U7670 , P1_U7671 , P1_U7672 , P1_U7673 , P1_U7674 , P1_U7675 , P1_U7676 , P1_U7677 , P1_U7678 , P1_U7679;
wire P1_U7680 , P1_U7681 , P1_U7682 , P1_U7683 , P1_U7684 , P1_U7685 , P1_U7686 , P1_U7687 , P1_U7688 , P1_U7689;
wire P1_U7690 , P1_U7691 , P1_U7692 , P1_U7693 , P1_U7694 , P1_U7695 , P1_U7696 , P1_U7697 , P1_U7698 , P1_U7699;
wire P1_U7700 , P1_U7701 , P1_U7702 , P1_U7703 , P1_U7704 , P1_U7705 , P1_U7706 , P1_U7707 , P1_U7708 , P1_U7709;
wire P1_U7710 , P1_U7711 , P1_U7712 , P1_U7713 , P1_U7714 , P1_U7715 , P1_U7716 , P1_U7717 , P1_U7718 , P1_U7719;
wire P1_U7720 , P1_U7721 , P1_U7722 , P1_U7723 , P1_U7724 , P1_U7725 , P1_U7726 , P1_U7727 , P1_U7728 , P1_U7729;
wire P1_U7730 , P1_U7731 , P1_U7732 , P1_U7733 , P1_U7734 , P1_U7735 , P1_U7736 , P1_U7737 , P1_U7738 , P1_U7739;
wire P1_U7740 , P1_U7741 , P1_U7742 , P1_U7743 , P1_U7744 , P1_U7745 , P1_U7746 , P1_U7747 , P1_U7748 , P1_U7749;
wire P1_U7750 , P1_U7751 , P1_U7752 , P1_U7753 , P1_U7754 , P1_U7755 , P1_U7756 , P1_U7757 , P1_U7758 , P1_U7759;
wire P1_U7760 , P1_U7761 , P1_U7762 , P1_U7763 , P1_U7764 , P1_U7765 , P1_U7766 , P1_U7767 , P1_U7768 , P1_U7769;
wire P1_U7770 , P1_U7771 , P1_U7772 , P1_U7773 , P1_U7774 , P1_U7775 , P1_U7776 , P1_U7777 , P1_U7778 , P1_U7779;
wire P1_U7780 , P1_U7781 , P1_U7782 , P1_U7783 , P1_U7784 , P1_U7785 , P1_U7786 , P1_U7787 , P1_U7788 , P1_U7789;
wire P1_U7790 , P1_U7791 , P1_U7792 , P1_U7793 , P1_U7794 , P1_ADD_405_U113 , P1_ADD_405_U112 , P1_ADD_405_U111 , P1_ADD_405_U110 , P1_ADD_405_U109;
wire P1_ADD_405_U108 , P1_ADD_405_U107 , P1_ADD_405_U106 , P1_ADD_405_U105 , P1_ADD_405_U104 , P1_ADD_405_U103 , P1_ADD_405_U102 , P1_ADD_405_U101 , P1_ADD_405_U100 , P1_ADD_405_U99;
wire P1_ADD_405_U98 , P1_ADD_405_U97 , P1_ADD_405_U96 , P1_ADD_405_U95 , P1_ADD_405_U94 , P1_ADD_405_U93 , P1_ADD_405_U92 , P1_ADD_405_U91 , P1_ADD_405_U90 , P1_ADD_405_U89;
wire P1_ADD_405_U88 , P1_ADD_405_U87 , LT_782_120_U6 , LT_782_120_U7 , LT_782_U6 , LT_782_U7 , LT_748_U6 , R170_U6 , R170_U7 , R170_U8;
wire R170_U9 , R170_U10 , R170_U11 , R170_U12 , R170_U13 , R170_U14 , R170_U15 , R165_U6 , R165_U7 , R165_U8;
wire R165_U9 , R165_U10 , R165_U11 , R165_U12 , R165_U13 , R165_U14 , R165_U15 , LT_782_119_U6 , LT_782_119_U7 , P3_ADD_526_U5;
wire P3_ADD_526_U6 , P3_ADD_526_U7 , P3_ADD_526_U8 , P3_ADD_526_U9 , P3_ADD_526_U10 , P3_ADD_526_U11 , P3_ADD_526_U12 , P3_ADD_526_U13 , P3_ADD_526_U14 , P3_ADD_526_U15;
wire P3_ADD_526_U16 , P3_ADD_526_U17 , P3_ADD_526_U18 , P3_ADD_526_U19 , P3_ADD_526_U20 , P3_ADD_526_U21 , P3_ADD_526_U22 , P3_ADD_526_U23 , P3_ADD_526_U24 , P3_ADD_526_U25;
wire P3_ADD_526_U26 , P3_ADD_526_U27 , P3_ADD_526_U28 , P3_ADD_526_U29 , P3_ADD_526_U30 , P3_ADD_526_U31 , P3_ADD_526_U32 , P3_ADD_526_U33 , P3_ADD_526_U34 , P3_ADD_526_U35;
wire P3_ADD_526_U36 , P3_ADD_526_U37 , P3_ADD_526_U38 , P3_ADD_526_U39 , P3_ADD_526_U40 , P3_ADD_526_U41 , P3_ADD_526_U42 , P3_ADD_526_U43 , P3_ADD_526_U44 , P3_ADD_526_U45;
wire P3_ADD_526_U46 , P3_ADD_526_U47 , P3_ADD_526_U48 , P3_ADD_526_U49 , P3_ADD_526_U50 , P3_ADD_526_U51 , P3_ADD_526_U52 , P3_ADD_526_U53 , P3_ADD_526_U54 , P3_ADD_526_U55;
wire P3_ADD_526_U56 , P3_ADD_526_U57 , P3_ADD_526_U58 , P3_ADD_526_U59 , P3_ADD_526_U60 , P3_ADD_526_U61 , P3_ADD_526_U62 , P3_ADD_526_U63 , P3_ADD_526_U64 , P3_ADD_526_U65;
wire P3_ADD_526_U66 , P3_ADD_526_U67 , P3_ADD_526_U68 , P3_ADD_526_U69 , P3_ADD_526_U70 , P3_ADD_526_U71 , P3_ADD_526_U72 , P3_ADD_526_U73 , P3_ADD_526_U74 , P3_ADD_526_U75;
wire P3_ADD_526_U76 , P3_ADD_526_U77 , P3_ADD_526_U78 , P3_ADD_526_U79 , P3_ADD_526_U80 , P3_ADD_526_U81 , P3_ADD_526_U82 , P3_ADD_526_U83 , P3_ADD_526_U84 , P3_ADD_526_U85;
wire P3_ADD_526_U86 , P3_ADD_526_U87 , P3_ADD_526_U88 , P3_ADD_526_U89 , P3_ADD_526_U90 , P3_ADD_526_U91 , P3_ADD_526_U92 , P3_ADD_526_U93 , P3_ADD_526_U94 , P3_ADD_526_U95;
wire P3_ADD_526_U96 , P3_ADD_526_U97 , P3_ADD_526_U98 , P3_ADD_526_U99 , P3_ADD_526_U100 , P3_ADD_526_U101 , P3_ADD_526_U102 , P3_ADD_526_U103 , P3_ADD_526_U104 , P3_ADD_526_U105;
wire P3_ADD_526_U106 , P3_ADD_526_U107 , P3_ADD_526_U108 , P3_ADD_526_U109 , P3_ADD_526_U110 , P3_ADD_526_U111 , P3_ADD_526_U112 , P3_ADD_526_U113 , P3_ADD_526_U114 , P3_ADD_526_U115;
wire P3_ADD_526_U116 , P3_ADD_526_U117 , P3_ADD_526_U118 , P3_ADD_526_U119 , P3_ADD_526_U120 , P3_ADD_526_U121 , P3_ADD_526_U122 , P3_ADD_526_U123 , P3_ADD_526_U124 , P3_ADD_526_U125;
wire P3_ADD_526_U126 , P3_ADD_526_U127 , P3_ADD_526_U128 , P3_ADD_526_U129 , P3_ADD_526_U130 , P3_ADD_526_U131 , P3_ADD_526_U132 , P3_ADD_526_U133 , P3_ADD_526_U134 , P3_ADD_526_U135;
wire P3_ADD_526_U136 , P3_ADD_526_U137 , P3_ADD_526_U138 , P3_ADD_526_U139 , P3_ADD_526_U140 , P3_ADD_526_U141 , P3_ADD_526_U142 , P3_ADD_526_U143 , P3_ADD_526_U144 , P3_ADD_526_U145;
wire P3_ADD_526_U146 , P3_ADD_526_U147 , P3_ADD_526_U148 , P3_ADD_526_U149 , P3_ADD_526_U150 , P3_ADD_526_U151 , P3_ADD_526_U152 , P3_ADD_526_U153 , P3_ADD_526_U154 , P3_ADD_526_U155;
wire P3_ADD_526_U156 , P3_ADD_526_U157 , P3_ADD_526_U158 , P3_ADD_526_U159 , P3_ADD_526_U160 , P3_ADD_526_U161 , P3_ADD_526_U162 , P3_ADD_526_U163 , P3_ADD_526_U164 , P3_ADD_526_U165;
wire P3_ADD_526_U166 , P3_ADD_526_U167 , P3_ADD_526_U168 , P3_ADD_526_U169 , P3_ADD_526_U170 , P3_ADD_526_U171 , P3_ADD_526_U172 , P3_ADD_526_U173 , P3_ADD_526_U174 , P3_ADD_526_U175;
wire P3_ADD_526_U176 , P3_ADD_526_U177 , P3_ADD_526_U178 , P3_ADD_526_U179 , P3_ADD_526_U180 , P3_ADD_526_U181 , P3_ADD_526_U182 , P3_ADD_526_U183 , P3_ADD_526_U184 , P3_ADD_526_U185;
wire P3_ADD_526_U186 , P3_ADD_526_U187 , P3_ADD_526_U188 , P3_ADD_526_U189 , P3_ADD_526_U190 , P3_ADD_526_U191 , P3_ADD_526_U192 , P3_ADD_526_U193 , P3_ADD_526_U194 , P3_ADD_526_U195;
wire P3_ADD_526_U196 , P3_ADD_526_U197 , P3_ADD_526_U198 , P3_ADD_526_U199 , P3_ADD_526_U200 , P3_ADD_526_U201 , P3_ADD_526_U202 , P3_ADD_552_U5 , P3_ADD_552_U6 , P3_ADD_552_U7;
wire P3_ADD_552_U8 , P3_ADD_552_U9 , P3_ADD_552_U10 , P3_ADD_552_U11 , P3_ADD_552_U12 , P3_ADD_552_U13 , P3_ADD_552_U14 , P3_ADD_552_U15 , P3_ADD_552_U16 , P3_ADD_552_U17;
wire P3_ADD_552_U18 , P3_ADD_552_U19 , P3_ADD_552_U20 , P3_ADD_552_U21 , P3_ADD_552_U22 , P3_ADD_552_U23 , P3_ADD_552_U24 , P3_ADD_552_U25 , P3_ADD_552_U26 , P3_ADD_552_U27;
wire P3_ADD_552_U28 , P3_ADD_552_U29 , P3_ADD_552_U30 , P3_ADD_552_U31 , P3_ADD_552_U32 , P3_ADD_552_U33 , P3_ADD_552_U34 , P3_ADD_552_U35 , P3_ADD_552_U36 , P3_ADD_552_U37;
wire P3_ADD_552_U38 , P3_ADD_552_U39 , P3_ADD_552_U40 , P3_ADD_552_U41 , P3_ADD_552_U42 , P3_ADD_552_U43 , P3_ADD_552_U44 , P3_ADD_552_U45 , P3_ADD_552_U46 , P3_ADD_552_U47;
wire P3_ADD_552_U48 , P3_ADD_552_U49 , P3_ADD_552_U50 , P3_ADD_552_U51 , P3_ADD_552_U52 , P3_ADD_552_U53 , P3_ADD_552_U54 , P3_ADD_552_U55 , P3_ADD_552_U56 , P3_ADD_552_U57;
wire P3_ADD_552_U58 , P3_ADD_552_U59 , P3_ADD_552_U60 , P3_ADD_552_U61 , P3_ADD_552_U62 , P3_ADD_552_U63 , P3_ADD_552_U64 , P3_ADD_552_U65 , P3_ADD_552_U66 , P3_ADD_552_U67;
wire P3_ADD_552_U68 , P3_ADD_552_U69 , P3_ADD_552_U70 , P3_ADD_552_U71 , P3_ADD_552_U72 , P3_ADD_552_U73 , P3_ADD_552_U74 , P3_ADD_552_U75 , P3_ADD_552_U76 , P3_ADD_552_U77;
wire P3_ADD_552_U78 , P3_ADD_552_U79 , P3_ADD_552_U80 , P3_ADD_552_U81 , P3_ADD_552_U82 , P3_ADD_552_U83 , P3_ADD_552_U84 , P3_ADD_552_U85 , P3_ADD_552_U86 , P3_ADD_552_U87;
wire P3_ADD_552_U88 , P3_ADD_552_U89 , P3_ADD_552_U90 , P3_ADD_552_U91 , P3_ADD_552_U92 , P3_ADD_552_U93 , P3_ADD_552_U94 , P3_ADD_552_U95 , P3_ADD_552_U96 , P3_ADD_552_U97;
wire P3_ADD_552_U98 , P3_ADD_552_U99 , P3_ADD_552_U100 , P3_ADD_552_U101 , P3_ADD_552_U102 , P3_ADD_552_U103 , P3_ADD_552_U104 , P3_ADD_552_U105 , P3_ADD_552_U106 , P3_ADD_552_U107;
wire P3_ADD_552_U108 , P3_ADD_552_U109 , P3_ADD_552_U110 , P3_ADD_552_U111 , P3_ADD_552_U112 , P3_ADD_552_U113 , P3_ADD_552_U114 , P3_ADD_552_U115 , P3_ADD_552_U116 , P3_ADD_552_U117;
wire P3_ADD_552_U118 , P3_ADD_552_U119 , P3_ADD_552_U120 , P3_ADD_552_U121 , P3_ADD_552_U122 , P3_ADD_552_U123 , P3_ADD_552_U124 , P3_ADD_552_U125 , P3_ADD_552_U126 , P3_ADD_552_U127;
wire P3_ADD_552_U128 , P3_ADD_552_U129 , P3_ADD_552_U130 , P3_ADD_552_U131 , P3_ADD_552_U132 , P3_ADD_552_U133 , P3_ADD_552_U134 , P3_ADD_552_U135 , P3_ADD_552_U136 , P3_ADD_552_U137;
wire P3_ADD_552_U138 , P3_ADD_552_U139 , P3_ADD_552_U140 , P3_ADD_552_U141 , P3_ADD_552_U142 , P3_ADD_552_U143 , P3_ADD_552_U144 , P3_ADD_552_U145 , P3_ADD_552_U146 , P3_ADD_552_U147;
wire P3_ADD_552_U148 , P3_ADD_552_U149 , P3_ADD_552_U150 , P3_ADD_552_U151 , P3_ADD_552_U152 , P3_ADD_552_U153 , P3_ADD_552_U154 , P3_ADD_552_U155 , P3_ADD_552_U156 , P3_ADD_552_U157;
wire P3_ADD_552_U158 , P3_ADD_552_U159 , P3_ADD_552_U160 , P3_ADD_552_U161 , P3_ADD_552_U162 , P3_ADD_552_U163 , P3_ADD_552_U164 , P3_ADD_552_U165 , P3_ADD_552_U166 , P3_ADD_552_U167;
wire P3_ADD_552_U168 , P3_ADD_552_U169 , P3_ADD_552_U170 , P3_ADD_552_U171 , P3_ADD_552_U172 , P3_ADD_552_U173 , P3_ADD_552_U174 , P3_ADD_552_U175 , P3_ADD_552_U176 , P3_ADD_552_U177;
wire P3_ADD_552_U178 , P3_ADD_552_U179 , P3_ADD_552_U180 , P3_ADD_552_U181 , P3_ADD_552_U182 , P3_ADD_552_U183 , P3_ADD_552_U184 , P3_ADD_552_U185 , P3_ADD_552_U186 , P3_ADD_552_U187;
wire P3_ADD_552_U188 , P3_ADD_552_U189 , P3_ADD_552_U190 , P3_ADD_552_U191 , P3_ADD_552_U192 , P3_ADD_552_U193 , P3_ADD_552_U194 , P3_ADD_552_U195 , P3_ADD_552_U196 , P3_ADD_552_U197;
wire P3_ADD_552_U198 , P3_ADD_552_U199 , P3_ADD_552_U200 , P3_ADD_552_U201 , P3_ADD_552_U202 , P3_ADD_546_U5 , P3_ADD_546_U6 , P3_ADD_546_U7 , P3_ADD_546_U8 , P3_ADD_546_U9;
wire P3_ADD_546_U10 , P3_ADD_546_U11 , P3_ADD_546_U12 , P3_ADD_546_U13 , P3_ADD_546_U14 , P3_ADD_546_U15 , P3_ADD_546_U16 , P3_ADD_546_U17 , P3_ADD_546_U18 , P3_ADD_546_U19;
wire P3_ADD_546_U20 , P3_ADD_546_U21 , P3_ADD_546_U22 , P3_ADD_546_U23 , P3_ADD_546_U24 , P3_ADD_546_U25 , P3_ADD_546_U26 , P3_ADD_546_U27 , P3_ADD_546_U28 , P3_ADD_546_U29;
wire P3_ADD_546_U30 , P3_ADD_546_U31 , P3_ADD_546_U32 , P3_ADD_546_U33 , P3_ADD_546_U34 , P3_ADD_546_U35 , P3_ADD_546_U36 , P3_ADD_546_U37 , P3_ADD_546_U38 , P3_ADD_546_U39;
wire P3_ADD_546_U40 , P3_ADD_546_U41 , P3_ADD_546_U42 , P3_ADD_546_U43 , P3_ADD_546_U44 , P3_ADD_546_U45 , P3_ADD_546_U46 , P3_ADD_546_U47 , P3_ADD_546_U48 , P3_ADD_546_U49;
wire P3_ADD_546_U50 , P3_ADD_546_U51 , P3_ADD_546_U52 , P3_ADD_546_U53 , P3_ADD_546_U54 , P3_ADD_546_U55 , P3_ADD_546_U56 , P3_ADD_546_U57 , P3_ADD_546_U58 , P3_ADD_546_U59;
wire P3_ADD_546_U60 , P3_ADD_546_U61 , P3_ADD_546_U62 , P3_ADD_546_U63 , P3_ADD_546_U64 , P3_ADD_546_U65 , P3_ADD_546_U66 , P3_ADD_546_U67 , P3_ADD_546_U68 , P3_ADD_546_U69;
wire P3_ADD_546_U70 , P3_ADD_546_U71 , P3_ADD_546_U72 , P3_ADD_546_U73 , P3_ADD_546_U74 , P3_ADD_546_U75 , P3_ADD_546_U76 , P3_ADD_546_U77 , P3_ADD_546_U78 , P3_ADD_546_U79;
wire P3_ADD_546_U80 , P3_ADD_546_U81 , P3_ADD_546_U82 , P3_ADD_546_U83 , P3_ADD_546_U84 , P3_ADD_546_U85 , P3_ADD_546_U86 , P3_ADD_546_U87 , P3_ADD_546_U88 , P3_ADD_546_U89;
wire P3_ADD_546_U90 , P3_ADD_546_U91 , P3_ADD_546_U92 , P3_ADD_546_U93 , P3_ADD_546_U94 , P3_ADD_546_U95 , P3_ADD_546_U96 , P3_ADD_546_U97 , P3_ADD_546_U98 , P3_ADD_546_U99;
wire P3_ADD_546_U100 , P3_ADD_546_U101 , P3_ADD_546_U102 , P3_ADD_546_U103 , P3_ADD_546_U104 , P3_ADD_546_U105 , P3_ADD_546_U106 , P3_ADD_546_U107 , P3_ADD_546_U108 , P3_ADD_546_U109;
wire P3_ADD_546_U110 , P3_ADD_546_U111 , P3_ADD_546_U112 , P3_ADD_546_U113 , P3_ADD_546_U114 , P3_ADD_546_U115 , P3_ADD_546_U116 , P3_ADD_546_U117 , P3_ADD_546_U118 , P3_ADD_546_U119;
wire P3_ADD_546_U120 , P3_ADD_546_U121 , P3_ADD_546_U122 , P3_ADD_546_U123 , P3_ADD_546_U124 , P3_ADD_546_U125 , P3_ADD_546_U126 , P3_ADD_546_U127 , P3_ADD_546_U128 , P3_ADD_546_U129;
wire P3_ADD_546_U130 , P3_ADD_546_U131 , P3_ADD_546_U132 , P3_ADD_546_U133 , P3_ADD_546_U134 , P3_ADD_546_U135 , P3_ADD_546_U136 , P3_ADD_546_U137 , P3_ADD_546_U138 , P3_ADD_546_U139;
wire P3_ADD_546_U140 , P3_ADD_546_U141 , P3_ADD_546_U142 , P3_ADD_546_U143 , P3_ADD_546_U144 , P3_ADD_546_U145 , P3_ADD_546_U146 , P3_ADD_546_U147 , P3_ADD_546_U148 , P3_ADD_546_U149;
wire P3_ADD_546_U150 , P3_ADD_546_U151 , P3_ADD_546_U152 , P3_ADD_546_U153 , P3_ADD_546_U154 , P3_ADD_546_U155 , P3_ADD_546_U156 , P3_ADD_546_U157 , P3_ADD_546_U158 , P3_ADD_546_U159;
wire P3_ADD_546_U160 , P3_ADD_546_U161 , P3_ADD_546_U162 , P3_ADD_546_U163 , P3_ADD_546_U164 , P3_ADD_546_U165 , P3_ADD_546_U166 , P3_ADD_546_U167 , P3_ADD_546_U168 , P3_ADD_546_U169;
wire P3_ADD_546_U170 , P3_ADD_546_U171 , P3_ADD_546_U172 , P3_ADD_546_U173 , P3_ADD_546_U174 , P3_ADD_546_U175 , P3_ADD_546_U176 , P3_ADD_546_U177 , P3_ADD_546_U178 , P3_ADD_546_U179;
wire P3_ADD_546_U180 , P3_ADD_546_U181 , P3_ADD_546_U182 , P3_ADD_546_U183 , P3_ADD_546_U184 , P3_ADD_546_U185 , P3_ADD_546_U186 , P3_ADD_546_U187 , P3_ADD_546_U188 , P3_ADD_546_U189;
wire P3_ADD_546_U190 , P3_ADD_546_U191 , P3_ADD_546_U192 , P3_ADD_546_U193 , P3_ADD_546_U194 , P3_ADD_546_U195 , P3_ADD_546_U196 , P3_ADD_546_U197 , P3_ADD_546_U198 , P3_ADD_546_U199;
wire P3_ADD_546_U200 , P3_ADD_546_U201 , P3_ADD_546_U202 , P3_GTE_401_U6 , P3_GTE_401_U7 , P3_GTE_401_U8 , P3_GTE_401_U9 , P3_ADD_391_1180_U4 , P3_ADD_391_1180_U5 , P3_ADD_391_1180_U6;
wire P3_ADD_391_1180_U7 , P3_ADD_391_1180_U8 , P3_ADD_391_1180_U9 , P3_ADD_391_1180_U10 , P3_ADD_391_1180_U11 , P3_ADD_391_1180_U12 , P3_ADD_391_1180_U13 , P3_ADD_391_1180_U14 , P3_ADD_391_1180_U15 , P3_ADD_391_1180_U16;
wire P3_ADD_391_1180_U17 , P3_ADD_391_1180_U18 , P3_ADD_391_1180_U19 , P3_ADD_391_1180_U20 , P3_ADD_391_1180_U21 , P3_ADD_391_1180_U22 , P3_ADD_391_1180_U23 , P3_ADD_391_1180_U24 , P3_ADD_391_1180_U25 , P3_ADD_391_1180_U26;
wire P3_ADD_391_1180_U27 , P3_ADD_391_1180_U28 , P3_ADD_391_1180_U29 , P3_ADD_391_1180_U30 , P3_ADD_391_1180_U31 , P3_ADD_391_1180_U32 , P3_ADD_391_1180_U33 , P3_ADD_391_1180_U34 , P3_ADD_391_1180_U35 , P3_ADD_391_1180_U36;
wire P3_ADD_391_1180_U37 , P3_ADD_391_1180_U38 , P3_ADD_391_1180_U39 , P3_ADD_391_1180_U40 , P3_ADD_391_1180_U41 , P3_ADD_391_1180_U42 , P3_ADD_391_1180_U43 , P3_ADD_391_1180_U44 , P3_ADD_391_1180_U45 , P3_ADD_391_1180_U46;
wire P3_ADD_391_1180_U47 , P3_ADD_391_1180_U48 , P3_ADD_391_1180_U49 , P3_ADD_391_1180_U50 , P3_ADD_476_U4 , P3_ADD_476_U5 , P3_ADD_476_U6 , P3_ADD_476_U7 , P3_ADD_476_U8 , P3_ADD_476_U9;
wire P3_ADD_476_U10 , P3_ADD_476_U11 , P3_ADD_476_U12 , P3_ADD_476_U13 , P3_ADD_476_U14 , P3_ADD_476_U15 , P3_ADD_476_U16 , P3_ADD_476_U17 , P3_ADD_476_U18 , P3_ADD_476_U19;
wire P3_ADD_476_U20 , P3_ADD_476_U21 , P3_ADD_476_U22 , P3_ADD_476_U23 , P3_ADD_476_U24 , P3_ADD_476_U25 , P3_ADD_476_U26 , P3_ADD_476_U27 , P3_ADD_476_U28 , P3_ADD_476_U29;
wire P3_ADD_476_U30 , P3_ADD_476_U31 , P3_ADD_476_U32 , P3_ADD_476_U33 , P3_ADD_476_U34 , P3_ADD_476_U35 , P3_ADD_476_U36 , P3_ADD_476_U37 , P3_ADD_476_U38 , P3_ADD_476_U39;
wire P3_ADD_476_U40 , P3_ADD_476_U41 , P3_ADD_476_U42 , P3_ADD_476_U43 , P3_ADD_476_U44 , P3_ADD_476_U45 , P3_ADD_476_U46 , P3_ADD_476_U47 , P3_ADD_476_U48 , P3_ADD_476_U49;
wire P3_ADD_476_U50 , P3_ADD_476_U51 , P3_ADD_476_U52 , P3_ADD_476_U53 , P3_ADD_476_U54 , P3_ADD_476_U55 , P3_ADD_476_U56 , P3_ADD_476_U57 , P3_ADD_476_U58 , P3_ADD_476_U59;
wire P3_ADD_476_U60 , P3_ADD_476_U61 , P3_ADD_476_U62 , P3_ADD_476_U63 , P3_ADD_476_U64 , P3_ADD_476_U65 , P3_ADD_476_U66 , P3_ADD_476_U67 , P3_ADD_476_U68 , P3_ADD_476_U69;
wire P3_ADD_476_U70 , P3_ADD_476_U71 , P3_ADD_476_U72 , P3_ADD_476_U73 , P3_ADD_476_U74 , P3_ADD_476_U75 , P3_ADD_476_U76 , P3_ADD_476_U77 , P3_ADD_476_U78 , P3_ADD_476_U79;
wire P3_ADD_476_U80 , P3_ADD_476_U81 , P3_ADD_476_U82 , P3_ADD_476_U83 , P3_ADD_476_U84 , P3_ADD_476_U85 , P3_ADD_476_U86 , P3_ADD_476_U87 , P3_ADD_476_U88 , P3_ADD_476_U89;
wire P3_ADD_476_U90 , P3_ADD_476_U91 , P3_ADD_476_U92 , P3_ADD_476_U93 , P3_ADD_476_U94 , P3_ADD_476_U95 , P3_ADD_476_U96 , P3_ADD_476_U97 , P3_ADD_476_U98 , P3_ADD_476_U99;
wire P3_ADD_476_U100 , P3_ADD_476_U101 , P3_ADD_476_U102 , P3_ADD_476_U103 , P3_ADD_476_U104 , P3_ADD_476_U105 , P3_ADD_476_U106 , P3_ADD_476_U107 , P3_ADD_476_U108 , P3_ADD_476_U109;
wire P3_ADD_476_U110 , P3_ADD_476_U111 , P3_ADD_476_U112 , P3_ADD_476_U113 , P3_ADD_476_U114 , P3_ADD_476_U115 , P3_ADD_476_U116 , P3_ADD_476_U117 , P3_ADD_476_U118 , P3_ADD_476_U119;
wire P3_ADD_476_U120 , P3_ADD_476_U121 , P3_ADD_476_U122 , P3_ADD_476_U123 , P3_ADD_476_U124 , P3_ADD_476_U125 , P3_ADD_476_U126 , P3_ADD_476_U127 , P3_ADD_476_U128 , P3_ADD_476_U129;
wire P3_ADD_476_U130 , P3_ADD_476_U131 , P3_ADD_476_U132 , P3_ADD_476_U133 , P3_ADD_476_U134 , P3_ADD_476_U135 , P3_ADD_476_U136 , P3_ADD_476_U137 , P3_ADD_476_U138 , P3_ADD_476_U139;
wire P3_ADD_476_U140 , P3_ADD_476_U141 , P3_ADD_476_U142 , P3_ADD_476_U143 , P3_ADD_476_U144 , P3_ADD_476_U145 , P3_ADD_476_U146 , P3_ADD_476_U147 , P3_ADD_476_U148 , P3_ADD_476_U149;
wire P3_ADD_476_U150 , P3_ADD_476_U151 , P3_ADD_476_U152 , P3_ADD_476_U153 , P3_ADD_476_U154 , P3_ADD_476_U155 , P3_ADD_476_U156 , P3_ADD_476_U157 , P3_ADD_476_U158 , P3_ADD_476_U159;
wire P3_ADD_476_U160 , P3_ADD_476_U161 , P3_ADD_476_U162 , P3_ADD_476_U163 , P3_ADD_476_U164 , P3_ADD_476_U165 , P3_ADD_476_U166 , P3_ADD_476_U167 , P3_ADD_476_U168 , P3_ADD_476_U169;
wire P3_ADD_476_U170 , P3_ADD_476_U171 , P3_ADD_476_U172 , P3_ADD_476_U173 , P3_ADD_476_U174 , P3_ADD_476_U175 , P3_ADD_476_U176 , P3_ADD_476_U177 , P3_ADD_476_U178 , P3_ADD_476_U179;
wire P3_ADD_476_U180 , P3_ADD_476_U181 , P3_ADD_476_U182 , P3_GTE_390_U6 , P3_GTE_390_U7 , P3_GTE_390_U8 , P3_GTE_390_U9 , P3_ADD_531_U5 , P3_ADD_531_U6 , P3_ADD_531_U7;
wire P3_ADD_531_U8 , P3_ADD_531_U9 , P3_ADD_531_U10 , P3_ADD_531_U11 , P3_ADD_531_U12 , P3_ADD_531_U13 , P3_ADD_531_U14 , P3_ADD_531_U15 , P3_ADD_531_U16 , P3_ADD_531_U17;
wire P3_ADD_531_U18 , P3_ADD_531_U19 , P3_ADD_531_U20 , P3_ADD_531_U21 , P3_ADD_531_U22 , P3_ADD_531_U23 , P3_ADD_531_U24 , P3_ADD_531_U25 , P3_ADD_531_U26 , P3_ADD_531_U27;
wire P3_ADD_531_U28 , P3_ADD_531_U29 , P3_ADD_531_U30 , P3_ADD_531_U31 , P3_ADD_531_U32 , P3_ADD_531_U33 , P3_ADD_531_U34 , P3_ADD_531_U35 , P3_ADD_531_U36 , P3_ADD_531_U37;
wire P3_ADD_531_U38 , P3_ADD_531_U39 , P3_ADD_531_U40 , P3_ADD_531_U41 , P3_ADD_531_U42 , P3_ADD_531_U43 , P3_ADD_531_U44 , P3_ADD_531_U45 , P3_ADD_531_U46 , P3_ADD_531_U47;
wire P3_ADD_531_U48 , P3_ADD_531_U49 , P3_ADD_531_U50 , P3_ADD_531_U51 , P3_ADD_531_U52 , P3_ADD_531_U53 , P3_ADD_531_U54 , P3_ADD_531_U55 , P3_ADD_531_U56 , P3_ADD_531_U57;
wire P3_ADD_531_U58 , P3_ADD_531_U59 , P3_ADD_531_U60 , P3_ADD_531_U61 , P3_ADD_531_U62 , P3_ADD_531_U63 , P3_ADD_531_U64 , P3_ADD_531_U65 , P3_ADD_531_U66 , P3_ADD_531_U67;
wire P3_ADD_531_U68 , P3_ADD_531_U69 , P3_ADD_531_U70 , P3_ADD_531_U71 , P3_ADD_531_U72 , P3_ADD_531_U73 , P3_ADD_531_U74 , P3_ADD_531_U75 , P3_ADD_531_U76 , P3_ADD_531_U77;
wire P3_ADD_531_U78 , P3_ADD_531_U79 , P3_ADD_531_U80 , P3_ADD_531_U81 , P3_ADD_531_U82 , P3_ADD_531_U83 , P3_ADD_531_U84 , P3_ADD_531_U85 , P3_ADD_531_U86 , P3_ADD_531_U87;
wire P3_ADD_531_U88 , P3_ADD_531_U89 , P3_ADD_531_U90 , P3_ADD_531_U91 , P3_ADD_531_U92 , P3_ADD_531_U93 , P3_ADD_531_U94 , P3_ADD_531_U95 , P3_ADD_531_U96 , P3_ADD_531_U97;
wire P3_ADD_531_U98 , P3_ADD_531_U99 , P3_ADD_531_U100 , P3_ADD_531_U101 , P3_ADD_531_U102 , P3_ADD_531_U103 , P3_ADD_531_U104 , P3_ADD_531_U105 , P3_ADD_531_U106 , P3_ADD_531_U107;
wire P3_ADD_531_U108 , P3_ADD_531_U109 , P3_ADD_531_U110 , P3_ADD_531_U111 , P3_ADD_531_U112 , P3_ADD_531_U113 , P3_ADD_531_U114 , P3_ADD_531_U115 , P3_ADD_531_U116 , P3_ADD_531_U117;
wire P3_ADD_531_U118 , P3_ADD_531_U119 , P3_ADD_531_U120 , P3_ADD_531_U121 , P3_ADD_531_U122 , P3_ADD_531_U123 , P3_ADD_531_U124 , P3_ADD_531_U125 , P3_ADD_531_U126 , P3_ADD_531_U127;
wire P3_ADD_531_U128 , P3_ADD_531_U129 , P3_ADD_531_U130 , P3_ADD_531_U131 , P3_ADD_531_U132 , P3_ADD_531_U133 , P3_ADD_531_U134 , P3_ADD_531_U135 , P3_ADD_531_U136 , P3_ADD_531_U137;
wire P3_ADD_531_U138 , P3_ADD_531_U139 , P3_ADD_531_U140 , P3_ADD_531_U141 , P3_ADD_531_U142 , P3_ADD_531_U143 , P3_ADD_531_U144 , P3_ADD_531_U145 , P3_ADD_531_U146 , P3_ADD_531_U147;
wire P3_ADD_531_U148 , P3_ADD_531_U149 , P3_ADD_531_U150 , P3_ADD_531_U151 , P3_ADD_531_U152 , P3_ADD_531_U153 , P3_ADD_531_U154 , P3_ADD_531_U155 , P3_ADD_531_U156 , P3_ADD_531_U157;
wire P3_ADD_531_U158 , P3_ADD_531_U159 , P3_ADD_531_U160 , P3_ADD_531_U161 , P3_ADD_531_U162 , P3_ADD_531_U163 , P3_ADD_531_U164 , P3_ADD_531_U165 , P3_ADD_531_U166 , P3_ADD_531_U167;
wire P3_ADD_531_U168 , P3_ADD_531_U169 , P3_ADD_531_U170 , P3_ADD_531_U171 , P3_ADD_531_U172 , P3_ADD_531_U173 , P3_ADD_531_U174 , P3_ADD_531_U175 , P3_ADD_531_U176 , P3_ADD_531_U177;
wire P3_ADD_531_U178 , P3_ADD_531_U179 , P3_ADD_531_U180 , P3_ADD_531_U181 , P3_ADD_531_U182 , P3_ADD_531_U183 , P3_ADD_531_U184 , P3_ADD_531_U185 , P3_ADD_531_U186 , P3_ADD_531_U187;
wire P3_ADD_531_U188 , P3_ADD_531_U189 , P3_SUB_320_U6 , P3_SUB_320_U7 , P3_SUB_320_U8 , P3_SUB_320_U9 , P3_SUB_320_U10 , P3_SUB_320_U11 , P3_SUB_320_U12 , P3_SUB_320_U13;
wire P3_SUB_320_U14 , P3_SUB_320_U15 , P3_SUB_320_U16 , P3_SUB_320_U17 , P3_SUB_320_U18 , P3_SUB_320_U19 , P3_SUB_320_U20 , P3_SUB_320_U21 , P3_SUB_320_U22 , P3_SUB_320_U23;
wire P3_SUB_320_U24 , P3_SUB_320_U25 , P3_SUB_320_U26 , P3_SUB_320_U27 , P3_SUB_320_U28 , P3_SUB_320_U29 , P3_SUB_320_U30 , P3_SUB_320_U31 , P3_SUB_320_U32 , P3_SUB_320_U33;
wire P3_SUB_320_U34 , P3_SUB_320_U35 , P3_SUB_320_U36 , P3_SUB_320_U37 , P3_SUB_320_U38 , P3_SUB_320_U39 , P3_SUB_320_U40 , P3_SUB_320_U41 , P3_SUB_320_U42 , P3_SUB_320_U43;
wire P3_SUB_320_U44 , P3_SUB_320_U45 , P3_SUB_320_U46 , P3_SUB_320_U47 , P3_SUB_320_U48 , P3_SUB_320_U49 , P3_SUB_320_U50 , P3_SUB_320_U51 , P3_SUB_320_U52 , P3_SUB_320_U53;
wire P3_SUB_320_U54 , P3_SUB_320_U55 , P3_SUB_320_U56 , P3_SUB_320_U57 , P3_SUB_320_U58 , P3_SUB_320_U59 , P3_SUB_320_U60 , P3_SUB_320_U61 , P3_SUB_320_U62 , P3_SUB_320_U63;
wire P3_SUB_320_U64 , P3_SUB_320_U65 , P3_SUB_320_U66 , P3_SUB_320_U67 , P3_SUB_320_U68 , P3_SUB_320_U69 , P3_SUB_320_U70 , P3_SUB_320_U71 , P3_SUB_320_U72 , P3_SUB_320_U73;
wire P3_SUB_320_U74 , P3_SUB_320_U75 , P3_SUB_320_U76 , P3_SUB_320_U77 , P3_SUB_320_U78 , P3_SUB_320_U79 , P3_SUB_320_U80 , P3_SUB_320_U81 , P3_SUB_320_U82 , P3_SUB_320_U83;
wire P3_SUB_320_U84 , P3_SUB_320_U85 , P3_SUB_320_U86 , P3_SUB_320_U87 , P3_SUB_320_U88 , P3_SUB_320_U89 , P3_SUB_320_U90 , P3_SUB_320_U91 , P3_SUB_320_U92 , P3_SUB_320_U93;
wire P3_SUB_320_U94 , P3_SUB_320_U95 , P3_SUB_320_U96 , P3_SUB_320_U97 , P3_SUB_320_U98 , P3_SUB_320_U99 , P3_SUB_320_U100 , P3_SUB_320_U101 , P3_SUB_320_U102 , P3_SUB_320_U103;
wire P3_SUB_320_U104 , P3_SUB_320_U105 , P3_SUB_320_U106 , P3_SUB_320_U107 , P3_SUB_320_U108 , P3_SUB_320_U109 , P3_SUB_320_U110 , P3_SUB_320_U111 , P3_SUB_320_U112 , P3_SUB_320_U113;
wire P3_SUB_320_U114 , P3_SUB_320_U115 , P3_SUB_320_U116 , P3_SUB_320_U117 , P3_SUB_320_U118 , P3_SUB_320_U119 , P3_SUB_320_U120 , P3_SUB_320_U121 , P3_SUB_320_U122 , P3_SUB_320_U123;
wire P3_SUB_320_U124 , P3_SUB_320_U125 , P3_SUB_320_U126 , P3_SUB_320_U127 , P3_SUB_320_U128 , P3_SUB_320_U129 , P3_SUB_320_U130 , P3_SUB_320_U131 , P3_SUB_320_U132 , P3_SUB_320_U133;
wire P3_SUB_320_U134 , P3_SUB_320_U135 , P3_SUB_320_U136 , P3_SUB_320_U137 , P3_SUB_320_U138 , P3_SUB_320_U139 , P3_SUB_320_U140 , P3_SUB_320_U141 , P3_SUB_320_U142 , P3_SUB_320_U143;
wire P3_SUB_320_U144 , P3_SUB_320_U145 , P3_SUB_320_U146 , P3_SUB_320_U147 , P3_SUB_320_U148 , P3_SUB_320_U149 , P3_SUB_320_U150 , P3_SUB_320_U151 , P3_SUB_320_U152 , P3_SUB_320_U153;
wire P3_SUB_320_U154 , P3_SUB_320_U155 , P3_SUB_320_U156 , P3_SUB_320_U157 , P3_SUB_320_U158 , P3_SUB_320_U159 , P3_ADD_505_U5 , P3_ADD_505_U6 , P3_ADD_505_U7 , P3_ADD_505_U8;
wire P3_ADD_505_U9 , P3_ADD_505_U10 , P3_ADD_505_U11 , P3_ADD_505_U12 , P3_ADD_505_U13 , P3_ADD_505_U14 , P3_ADD_505_U15 , P3_ADD_505_U16 , P3_ADD_505_U17 , P3_ADD_505_U18;
wire P3_ADD_505_U19 , P3_ADD_505_U20 , P3_ADD_505_U21 , P3_ADD_505_U22 , P3_ADD_505_U23 , P3_ADD_505_U24 , P3_ADD_505_U25 , P3_ADD_505_U26 , P3_ADD_505_U27 , P3_ADD_505_U28;
wire P3_GTE_485_U6 , P3_GTE_485_U7 , P3_ADD_318_U4 , P3_ADD_318_U5 , P3_ADD_318_U6 , P3_ADD_318_U7 , P3_ADD_318_U8 , P3_ADD_318_U9 , P3_ADD_318_U10 , P3_ADD_318_U11;
wire P3_ADD_318_U12 , P3_ADD_318_U13 , P3_ADD_318_U14 , P3_ADD_318_U15 , P3_ADD_318_U16 , P3_ADD_318_U17 , P3_ADD_318_U18 , P3_ADD_318_U19 , P3_ADD_318_U20 , P3_ADD_318_U21;
wire P3_ADD_318_U22 , P3_ADD_318_U23 , P3_ADD_318_U24 , P3_ADD_318_U25 , P3_ADD_318_U26 , P3_ADD_318_U27 , P3_ADD_318_U28 , P3_ADD_318_U29 , P3_ADD_318_U30 , P3_ADD_318_U31;
wire P3_ADD_318_U32 , P3_ADD_318_U33 , P3_ADD_318_U34 , P3_ADD_318_U35 , P3_ADD_318_U36 , P3_ADD_318_U37 , P3_ADD_318_U38 , P3_ADD_318_U39 , P3_ADD_318_U40 , P3_ADD_318_U41;
wire P3_ADD_318_U42 , P3_ADD_318_U43 , P3_ADD_318_U44 , P3_ADD_318_U45 , P3_ADD_318_U46 , P3_ADD_318_U47 , P3_ADD_318_U48 , P3_ADD_318_U49 , P3_ADD_318_U50 , P3_ADD_318_U51;
wire P3_ADD_318_U52 , P3_ADD_318_U53 , P3_ADD_318_U54 , P3_ADD_318_U55 , P3_ADD_318_U56 , P3_ADD_318_U57 , P3_ADD_318_U58 , P3_ADD_318_U59 , P3_ADD_318_U60 , P3_ADD_318_U61;
wire P3_ADD_318_U62 , P3_ADD_318_U63 , P3_ADD_318_U64 , P3_ADD_318_U65 , P3_ADD_318_U66 , P3_ADD_318_U67 , P3_ADD_318_U68 , P3_ADD_318_U69 , P3_ADD_318_U70 , P3_ADD_318_U71;
wire P3_ADD_318_U72 , P3_ADD_318_U73 , P3_ADD_318_U74 , P3_ADD_318_U75 , P3_ADD_318_U76 , P3_ADD_318_U77 , P3_ADD_318_U78 , P3_ADD_318_U79 , P3_ADD_318_U80 , P3_ADD_318_U81;
wire P3_ADD_318_U82 , P3_ADD_318_U83 , P3_ADD_318_U84 , P3_ADD_318_U85 , P3_ADD_318_U86 , P3_ADD_318_U87 , P3_ADD_318_U88 , P3_ADD_318_U89 , P3_ADD_318_U90 , P3_ADD_318_U91;
wire P3_ADD_318_U92 , P3_ADD_318_U93 , P3_ADD_318_U94 , P3_ADD_318_U95 , P3_ADD_318_U96 , P3_ADD_318_U97 , P3_ADD_318_U98 , P3_ADD_318_U99 , P3_ADD_318_U100 , P3_ADD_318_U101;
wire P3_ADD_318_U102 , P3_ADD_318_U103 , P3_ADD_318_U104 , P3_ADD_318_U105 , P3_ADD_318_U106 , P3_ADD_318_U107 , P3_ADD_318_U108 , P3_ADD_318_U109 , P3_ADD_318_U110 , P3_ADD_318_U111;
wire P3_ADD_318_U112 , P3_ADD_318_U113 , P3_ADD_318_U114 , P3_ADD_318_U115 , P3_ADD_318_U116 , P3_ADD_318_U117 , P3_ADD_318_U118 , P3_ADD_318_U119 , P3_ADD_318_U120 , P3_ADD_318_U121;
wire P3_ADD_318_U122 , P3_ADD_318_U123 , P3_ADD_318_U124 , P3_ADD_318_U125 , P3_ADD_318_U126 , P3_ADD_318_U127 , P3_ADD_318_U128 , P3_ADD_318_U129 , P3_ADD_318_U130 , P3_ADD_318_U131;
wire P3_ADD_318_U132 , P3_ADD_318_U133 , P3_ADD_318_U134 , P3_ADD_318_U135 , P3_ADD_318_U136 , P3_ADD_318_U137 , P3_ADD_318_U138 , P3_ADD_318_U139 , P3_ADD_318_U140 , P3_ADD_318_U141;
wire P3_ADD_318_U142 , P3_ADD_318_U143 , P3_ADD_318_U144 , P3_ADD_318_U145 , P3_ADD_318_U146 , P3_ADD_318_U147 , P3_ADD_318_U148 , P3_ADD_318_U149 , P3_ADD_318_U150 , P3_ADD_318_U151;
wire P3_ADD_318_U152 , P3_ADD_318_U153 , P3_ADD_318_U154 , P3_ADD_318_U155 , P3_ADD_318_U156 , P3_ADD_318_U157 , P3_ADD_318_U158 , P3_ADD_318_U159 , P3_ADD_318_U160 , P3_ADD_318_U161;
wire P3_ADD_318_U162 , P3_ADD_318_U163 , P3_ADD_318_U164 , P3_ADD_318_U165 , P3_ADD_318_U166 , P3_ADD_318_U167 , P3_ADD_318_U168 , P3_ADD_318_U169 , P3_ADD_318_U170 , P3_ADD_318_U171;
wire P3_ADD_318_U172 , P3_ADD_318_U173 , P3_ADD_318_U174 , P3_ADD_318_U175 , P3_ADD_318_U176 , P3_ADD_318_U177 , P3_ADD_318_U178 , P3_ADD_318_U179 , P3_ADD_318_U180 , P3_ADD_318_U181;
wire P3_ADD_318_U182 , P3_SUB_370_U6 , P3_SUB_370_U7 , P3_SUB_370_U8 , P3_SUB_370_U9 , P3_SUB_370_U10 , P3_SUB_370_U11 , P3_SUB_370_U12 , P3_SUB_370_U13 , P3_SUB_370_U14;
wire P3_SUB_370_U15 , P3_SUB_370_U16 , P3_SUB_370_U17 , P3_SUB_370_U18 , P3_SUB_370_U19 , P3_SUB_370_U20 , P3_SUB_370_U21 , P3_SUB_370_U22 , P3_SUB_370_U23 , P3_SUB_370_U24;
wire P3_SUB_370_U25 , P3_SUB_370_U26 , P3_SUB_370_U27 , P3_SUB_370_U28 , P3_SUB_370_U29 , P3_SUB_370_U30 , P3_SUB_370_U31 , P3_SUB_370_U32 , P3_SUB_370_U33 , P3_SUB_370_U34;
wire P3_SUB_370_U35 , P3_SUB_370_U36 , P3_SUB_370_U37 , P3_SUB_370_U38 , P3_SUB_370_U39 , P3_SUB_370_U40 , P3_SUB_370_U41 , P3_SUB_370_U42 , P3_SUB_370_U43 , P3_SUB_370_U44;
wire P3_SUB_370_U45 , P3_SUB_370_U46 , P3_SUB_370_U47 , P3_SUB_370_U48 , P3_SUB_370_U49 , P3_SUB_370_U50 , P3_SUB_370_U51 , P3_SUB_370_U52 , P3_SUB_370_U53 , P3_SUB_370_U54;
wire P3_SUB_370_U55 , P3_SUB_370_U56 , P3_SUB_370_U57 , P3_SUB_370_U58 , P3_SUB_370_U59 , P3_SUB_370_U60 , P3_SUB_370_U61 , P3_SUB_370_U62 , P3_SUB_370_U63 , P3_SUB_370_U64;
wire P3_SUB_370_U65 , P3_SUB_370_U66 , P3_ADD_315_U4 , P3_ADD_315_U5 , P3_ADD_315_U6 , P3_ADD_315_U7 , P3_ADD_315_U8 , P3_ADD_315_U9 , P3_ADD_315_U10 , P3_ADD_315_U11;
wire P3_ADD_315_U12 , P3_ADD_315_U13 , P3_ADD_315_U14 , P3_ADD_315_U15 , P3_ADD_315_U16 , P3_ADD_315_U17 , P3_ADD_315_U18 , P3_ADD_315_U19 , P3_ADD_315_U20 , P3_ADD_315_U21;
wire P3_ADD_315_U22 , P3_ADD_315_U23 , P3_ADD_315_U24 , P3_ADD_315_U25 , P3_ADD_315_U26 , P3_ADD_315_U27 , P3_ADD_315_U28 , P3_ADD_315_U29 , P3_ADD_315_U30 , P3_ADD_315_U31;
wire P3_ADD_315_U32 , P3_ADD_315_U33 , P3_ADD_315_U34 , P3_ADD_315_U35 , P3_ADD_315_U36 , P3_ADD_315_U37 , P3_ADD_315_U38 , P3_ADD_315_U39 , P3_ADD_315_U40 , P3_ADD_315_U41;
wire P3_ADD_315_U42 , P3_ADD_315_U43 , P3_ADD_315_U44 , P3_ADD_315_U45 , P3_ADD_315_U46 , P3_ADD_315_U47 , P3_ADD_315_U48 , P3_ADD_315_U49 , P3_ADD_315_U50 , P3_ADD_315_U51;
wire P3_ADD_315_U52 , P3_ADD_315_U53 , P3_ADD_315_U54 , P3_ADD_315_U55 , P3_ADD_315_U56 , P3_ADD_315_U57 , P3_ADD_315_U58 , P3_ADD_315_U59 , P3_ADD_315_U60 , P3_ADD_315_U61;
wire P3_ADD_315_U62 , P3_ADD_315_U63 , P3_ADD_315_U64 , P3_ADD_315_U65 , P3_ADD_315_U66 , P3_ADD_315_U67 , P3_ADD_315_U68 , P3_ADD_315_U69 , P3_ADD_315_U70 , P3_ADD_315_U71;
wire P3_ADD_315_U72 , P3_ADD_315_U73 , P3_ADD_315_U74 , P3_ADD_315_U75 , P3_ADD_315_U76 , P3_ADD_315_U77 , P3_ADD_315_U78 , P3_ADD_315_U79 , P3_ADD_315_U80 , P3_ADD_315_U81;
wire P3_ADD_315_U82 , P3_ADD_315_U83 , P3_ADD_315_U84 , P3_ADD_315_U85 , P3_ADD_315_U86 , P3_ADD_315_U87 , P3_ADD_315_U88 , P3_ADD_315_U89 , P3_ADD_315_U90 , P3_ADD_315_U91;
wire P3_ADD_315_U92 , P3_ADD_315_U93 , P3_ADD_315_U94 , P3_ADD_315_U95 , P3_ADD_315_U96 , P3_ADD_315_U97 , P3_ADD_315_U98 , P3_ADD_315_U99 , P3_ADD_315_U100 , P3_ADD_315_U101;
wire P3_ADD_315_U102 , P3_ADD_315_U103 , P3_ADD_315_U104 , P3_ADD_315_U105 , P3_ADD_315_U106 , P3_ADD_315_U107 , P3_ADD_315_U108 , P3_ADD_315_U109 , P3_ADD_315_U110 , P3_ADD_315_U111;
wire P3_ADD_315_U112 , P3_ADD_315_U113 , P3_ADD_315_U114 , P3_ADD_315_U115 , P3_ADD_315_U116 , P3_ADD_315_U117 , P3_ADD_315_U118 , P3_ADD_315_U119 , P3_ADD_315_U120 , P3_ADD_315_U121;
wire P3_ADD_315_U122 , P3_ADD_315_U123 , P3_ADD_315_U124 , P3_ADD_315_U125 , P3_ADD_315_U126 , P3_ADD_315_U127 , P3_ADD_315_U128 , P3_ADD_315_U129 , P3_ADD_315_U130 , P3_ADD_315_U131;
wire P3_ADD_315_U132 , P3_ADD_315_U133 , P3_ADD_315_U134 , P3_ADD_315_U135 , P3_ADD_315_U136 , P3_ADD_315_U137 , P3_ADD_315_U138 , P3_ADD_315_U139 , P3_ADD_315_U140 , P3_ADD_315_U141;
wire P3_ADD_315_U142 , P3_ADD_315_U143 , P3_ADD_315_U144 , P3_ADD_315_U145 , P3_ADD_315_U146 , P3_ADD_315_U147 , P3_ADD_315_U148 , P3_ADD_315_U149 , P3_ADD_315_U150 , P3_ADD_315_U151;
wire P3_ADD_315_U152 , P3_ADD_315_U153 , P3_ADD_315_U154 , P3_ADD_315_U155 , P3_ADD_315_U156 , P3_ADD_315_U157 , P3_ADD_315_U158 , P3_ADD_315_U159 , P3_ADD_315_U160 , P3_ADD_315_U161;
wire P3_ADD_315_U162 , P3_ADD_315_U163 , P3_ADD_315_U164 , P3_ADD_315_U165 , P3_ADD_315_U166 , P3_ADD_315_U167 , P3_ADD_315_U168 , P3_ADD_315_U169 , P3_ADD_315_U170 , P3_ADD_315_U171;
wire P3_ADD_315_U172 , P3_ADD_315_U173 , P3_ADD_315_U174 , P3_ADD_315_U175 , P3_ADD_315_U176 , P3_GTE_355_U6 , P3_GTE_355_U7 , P3_GTE_355_U8 , P3_ADD_360_1242_U4 , P3_ADD_360_1242_U5;
wire P3_ADD_360_1242_U6 , P3_ADD_360_1242_U7 , P3_ADD_360_1242_U8 , P3_ADD_360_1242_U9 , P3_ADD_360_1242_U10 , P3_ADD_360_1242_U11 , P3_ADD_360_1242_U12 , P3_ADD_360_1242_U13 , P3_ADD_360_1242_U14 , P3_ADD_360_1242_U15;
wire P3_ADD_360_1242_U16 , P3_ADD_360_1242_U17 , P3_ADD_360_1242_U18 , P3_ADD_360_1242_U19 , P3_ADD_360_1242_U20 , P3_ADD_360_1242_U21 , P3_ADD_360_1242_U22 , P3_ADD_360_1242_U23 , P3_ADD_360_1242_U24 , P3_ADD_360_1242_U25;
wire P3_ADD_360_1242_U26 , P3_ADD_360_1242_U27 , P3_ADD_360_1242_U28 , P3_ADD_360_1242_U29 , P3_ADD_360_1242_U30 , P3_ADD_360_1242_U31 , P3_ADD_360_1242_U32 , P3_ADD_360_1242_U33 , P3_ADD_360_1242_U34 , P3_ADD_360_1242_U35;
wire P3_ADD_360_1242_U36 , P3_ADD_360_1242_U37 , P3_ADD_360_1242_U38 , P3_ADD_360_1242_U39 , P3_ADD_360_1242_U40 , P3_ADD_360_1242_U41 , P3_ADD_360_1242_U42 , P3_ADD_360_1242_U43 , P3_ADD_360_1242_U44 , P3_ADD_360_1242_U45;
wire P3_ADD_360_1242_U46 , P3_ADD_360_1242_U47 , P3_ADD_360_1242_U48 , P3_ADD_360_1242_U49 , P3_ADD_360_1242_U50 , P3_ADD_360_1242_U51 , P3_ADD_360_1242_U52 , P3_ADD_360_1242_U53 , P3_ADD_360_1242_U54 , P3_ADD_360_1242_U55;
wire P3_ADD_360_1242_U56 , P3_ADD_360_1242_U57 , P3_ADD_360_1242_U58 , P3_ADD_360_1242_U59 , P3_ADD_360_1242_U60 , P3_ADD_360_1242_U61 , P3_ADD_360_1242_U62 , P3_ADD_360_1242_U63 , P3_ADD_360_1242_U64 , P3_ADD_360_1242_U65;
wire P3_ADD_360_1242_U66 , P3_ADD_360_1242_U67 , P3_ADD_360_1242_U68 , P3_ADD_360_1242_U69 , P3_ADD_360_1242_U70 , P3_ADD_360_1242_U71 , P3_ADD_360_1242_U72 , P3_ADD_360_1242_U73 , P3_ADD_360_1242_U74 , P3_ADD_360_1242_U75;
wire P3_ADD_360_1242_U76 , P3_ADD_360_1242_U77 , P3_ADD_360_1242_U78 , P3_ADD_360_1242_U79 , P3_ADD_360_1242_U80 , P3_ADD_360_1242_U81 , P3_ADD_360_1242_U82 , P3_ADD_360_1242_U83 , P3_ADD_360_1242_U84 , P3_ADD_360_1242_U85;
wire P3_ADD_360_1242_U86 , P3_ADD_360_1242_U87 , P3_ADD_360_1242_U88 , P3_ADD_360_1242_U89 , P3_ADD_360_1242_U90 , P3_ADD_360_1242_U91 , P3_ADD_360_1242_U92 , P3_ADD_360_1242_U93 , P3_ADD_360_1242_U94 , P3_ADD_360_1242_U95;
wire P3_ADD_360_1242_U96 , P3_ADD_360_1242_U97 , P3_ADD_360_1242_U98 , P3_ADD_360_1242_U99 , P3_ADD_360_1242_U100 , P3_ADD_360_1242_U101 , P3_ADD_360_1242_U102 , P3_ADD_360_1242_U103 , P3_ADD_360_1242_U104 , P3_ADD_360_1242_U105;
wire P3_ADD_360_1242_U106 , P3_ADD_360_1242_U107 , P3_ADD_360_1242_U108 , P3_ADD_360_1242_U109 , P3_ADD_360_1242_U110 , P3_ADD_360_1242_U111 , P3_ADD_360_1242_U112 , P3_ADD_360_1242_U113 , P3_ADD_360_1242_U114 , P3_ADD_360_1242_U115;
wire P3_ADD_360_1242_U116 , P3_ADD_360_1242_U117 , P3_ADD_360_1242_U118 , P3_ADD_360_1242_U119 , P3_ADD_360_1242_U120 , P3_ADD_360_1242_U121 , P3_ADD_360_1242_U122 , P3_ADD_360_1242_U123 , P3_ADD_360_1242_U124 , P3_ADD_360_1242_U125;
wire P3_ADD_360_1242_U126 , P3_ADD_360_1242_U127 , P3_ADD_360_1242_U128 , P3_ADD_360_1242_U129 , P3_ADD_360_1242_U130 , P3_ADD_360_1242_U131 , P3_ADD_360_1242_U132 , P3_ADD_360_1242_U133 , P3_ADD_360_1242_U134 , P3_ADD_360_1242_U135;
wire P3_ADD_360_1242_U136 , P3_ADD_360_1242_U137 , P3_ADD_360_1242_U138 , P3_ADD_360_1242_U139 , P3_ADD_360_1242_U140 , P3_ADD_360_1242_U141 , P3_ADD_360_1242_U142 , P3_ADD_360_1242_U143 , P3_ADD_360_1242_U144 , P3_ADD_360_1242_U145;
wire P3_ADD_360_1242_U146 , P3_ADD_360_1242_U147 , P3_ADD_360_1242_U148 , P3_ADD_360_1242_U149 , P3_ADD_360_1242_U150 , P3_ADD_360_1242_U151 , P3_ADD_360_1242_U152 , P3_ADD_360_1242_U153 , P3_ADD_360_1242_U154 , P3_ADD_360_1242_U155;
wire P3_ADD_360_1242_U156 , P3_ADD_360_1242_U157 , P3_ADD_360_1242_U158 , P3_ADD_360_1242_U159 , P3_ADD_360_1242_U160 , P3_ADD_360_1242_U161 , P3_ADD_360_1242_U162 , P3_ADD_360_1242_U163 , P3_ADD_360_1242_U164 , P3_ADD_360_1242_U165;
wire P3_ADD_360_1242_U166 , P3_ADD_360_1242_U167 , P3_ADD_360_1242_U168 , P3_ADD_360_1242_U169 , P3_ADD_360_1242_U170 , P3_ADD_360_1242_U171 , P3_ADD_360_1242_U172 , P3_ADD_360_1242_U173 , P3_ADD_360_1242_U174 , P3_ADD_360_1242_U175;
wire P3_ADD_360_1242_U176 , P3_ADD_360_1242_U177 , P3_ADD_360_1242_U178 , P3_ADD_360_1242_U179 , P3_ADD_360_1242_U180 , P3_ADD_360_1242_U181 , P3_ADD_360_1242_U182 , P3_ADD_360_1242_U183 , P3_ADD_360_1242_U184 , P3_ADD_360_1242_U185;
wire P3_ADD_360_1242_U186 , P3_ADD_360_1242_U187 , P3_ADD_360_1242_U188 , P3_ADD_360_1242_U189 , P3_ADD_360_1242_U190 , P3_ADD_360_1242_U191 , P3_ADD_360_1242_U192 , P3_ADD_360_1242_U193 , P3_ADD_360_1242_U194 , P3_ADD_360_1242_U195;
wire P3_ADD_360_1242_U196 , P3_ADD_360_1242_U197 , P3_ADD_360_1242_U198 , P3_ADD_360_1242_U199 , P3_ADD_360_1242_U200 , P3_ADD_360_1242_U201 , P3_ADD_360_1242_U202 , P3_ADD_360_1242_U203 , P3_ADD_360_1242_U204 , P3_ADD_360_1242_U205;
wire P3_ADD_360_1242_U206 , P3_ADD_360_1242_U207 , P3_ADD_360_1242_U208 , P3_ADD_360_1242_U209 , P3_ADD_360_1242_U210 , P3_ADD_360_1242_U211 , P3_ADD_360_1242_U212 , P3_ADD_360_1242_U213 , P3_ADD_360_1242_U214 , P3_ADD_360_1242_U215;
wire P3_ADD_360_1242_U216 , P3_ADD_360_1242_U217 , P3_ADD_360_1242_U218 , P3_ADD_360_1242_U219 , P3_ADD_360_1242_U220 , P3_ADD_360_1242_U221 , P3_ADD_360_1242_U222 , P3_ADD_360_1242_U223 , P3_ADD_360_1242_U224 , P3_ADD_360_1242_U225;
wire P3_ADD_360_1242_U226 , P3_ADD_360_1242_U227 , P3_ADD_360_1242_U228 , P3_ADD_360_1242_U229 , P3_ADD_360_1242_U230 , P3_ADD_360_1242_U231 , P3_ADD_360_1242_U232 , P3_ADD_360_1242_U233 , P3_ADD_360_1242_U234 , P3_ADD_360_1242_U235;
wire P3_ADD_360_1242_U236 , P3_ADD_360_1242_U237 , P3_ADD_360_1242_U238 , P3_ADD_360_1242_U239 , P3_ADD_360_1242_U240 , P3_ADD_360_1242_U241 , P3_ADD_360_1242_U242 , P3_ADD_360_1242_U243 , P3_ADD_360_1242_U244 , P3_ADD_360_1242_U245;
wire P3_ADD_360_1242_U246 , P3_ADD_360_1242_U247 , P3_ADD_360_1242_U248 , P3_ADD_360_1242_U249 , P3_ADD_360_1242_U250 , P3_ADD_360_1242_U251 , P3_ADD_360_1242_U252 , P3_ADD_360_1242_U253 , P3_ADD_360_1242_U254 , P3_ADD_360_1242_U255;
wire P3_ADD_360_1242_U256 , P3_ADD_360_1242_U257 , P3_ADD_360_1242_U258 , P3_LT_563_1260_U6 , P3_LT_563_1260_U7 , P3_SUB_589_U6 , P3_SUB_589_U7 , P3_SUB_589_U8 , P3_SUB_589_U9 , P3_ADD_467_U4;
wire P3_ADD_467_U5 , P3_ADD_467_U6 , P3_ADD_467_U7 , P3_ADD_467_U8 , P3_ADD_467_U9 , P3_ADD_467_U10 , P3_ADD_467_U11 , P3_ADD_467_U12 , P3_ADD_467_U13 , P3_ADD_467_U14;
wire P3_ADD_467_U15 , P3_ADD_467_U16 , P3_ADD_467_U17 , P3_ADD_467_U18 , P3_ADD_467_U19 , P3_ADD_467_U20 , P3_ADD_467_U21 , P3_ADD_467_U22 , P3_ADD_467_U23 , P3_ADD_467_U24;
wire P3_ADD_467_U25 , P3_ADD_467_U26 , P3_ADD_467_U27 , P3_ADD_467_U28 , P3_ADD_467_U29 , P3_ADD_467_U30 , P3_ADD_467_U31 , P3_ADD_467_U32 , P3_ADD_467_U33 , P3_ADD_467_U34;
wire P3_ADD_467_U35 , P3_ADD_467_U36 , P3_ADD_467_U37 , P3_ADD_467_U38 , P3_ADD_467_U39 , P3_ADD_467_U40 , P3_ADD_467_U41 , P3_ADD_467_U42 , P3_ADD_467_U43 , P3_ADD_467_U44;
wire P3_ADD_467_U45 , P3_ADD_467_U46 , P3_ADD_467_U47 , P3_ADD_467_U48 , P3_ADD_467_U49 , P3_ADD_467_U50 , P3_ADD_467_U51 , P3_ADD_467_U52 , P3_ADD_467_U53 , P3_ADD_467_U54;
wire P3_ADD_467_U55 , P3_ADD_467_U56 , P3_ADD_467_U57 , P3_ADD_467_U58 , P3_ADD_467_U59 , P3_ADD_467_U60 , P3_ADD_467_U61 , P3_ADD_467_U62 , P3_ADD_467_U63 , P3_ADD_467_U64;
wire P3_ADD_467_U65 , P3_ADD_467_U66 , P3_ADD_467_U67 , P3_ADD_467_U68 , P3_ADD_467_U69 , P3_ADD_467_U70 , P3_ADD_467_U71 , P3_ADD_467_U72 , P3_ADD_467_U73 , P3_ADD_467_U74;
wire P3_ADD_467_U75 , P3_ADD_467_U76 , P3_ADD_467_U77 , P3_ADD_467_U78 , P3_ADD_467_U79 , P3_ADD_467_U80 , P3_ADD_467_U81 , P3_ADD_467_U82 , P3_ADD_467_U83 , P3_ADD_467_U84;
wire P3_ADD_467_U85 , P3_ADD_467_U86 , P3_ADD_467_U87 , P3_ADD_467_U88 , P3_ADD_467_U89 , P3_ADD_467_U90 , P3_ADD_467_U91 , P3_ADD_467_U92 , P3_ADD_467_U93 , P3_ADD_467_U94;
wire P3_ADD_467_U95 , P3_ADD_467_U96 , P3_ADD_467_U97 , P3_ADD_467_U98 , P3_ADD_467_U99 , P3_ADD_467_U100 , P3_ADD_467_U101 , P3_ADD_467_U102 , P3_ADD_467_U103 , P3_ADD_467_U104;
wire P3_ADD_467_U105 , P3_ADD_467_U106 , P3_ADD_467_U107 , P3_ADD_467_U108 , P3_ADD_467_U109 , P3_ADD_467_U110 , P3_ADD_467_U111 , P3_ADD_467_U112 , P3_ADD_467_U113 , P3_ADD_467_U114;
wire P3_ADD_467_U115 , P3_ADD_467_U116 , P3_ADD_467_U117 , P3_ADD_467_U118 , P3_ADD_467_U119 , P3_ADD_467_U120 , P3_ADD_467_U121 , P3_ADD_467_U122 , P3_ADD_467_U123 , P3_ADD_467_U124;
wire P3_ADD_467_U125 , P3_ADD_467_U126 , P3_ADD_467_U127 , P3_ADD_467_U128 , P3_ADD_467_U129 , P3_ADD_467_U130 , P3_ADD_467_U131 , P3_ADD_467_U132 , P3_ADD_467_U133 , P3_ADD_467_U134;
wire P3_ADD_467_U135 , P3_ADD_467_U136 , P3_ADD_467_U137 , P3_ADD_467_U138 , P3_ADD_467_U139 , P3_ADD_467_U140 , P3_ADD_467_U141 , P3_ADD_467_U142 , P3_ADD_467_U143 , P3_ADD_467_U144;
wire P3_ADD_467_U145 , P3_ADD_467_U146 , P3_ADD_467_U147 , P3_ADD_467_U148 , P3_ADD_467_U149 , P3_ADD_467_U150 , P3_ADD_467_U151 , P3_ADD_467_U152 , P3_ADD_467_U153 , P3_ADD_467_U154;
wire P3_ADD_467_U155 , P3_ADD_467_U156 , P3_ADD_467_U157 , P3_ADD_467_U158 , P3_ADD_467_U159 , P3_ADD_467_U160 , P3_ADD_467_U161 , P3_ADD_467_U162 , P3_ADD_467_U163 , P3_ADD_467_U164;
wire P3_ADD_467_U165 , P3_ADD_467_U166 , P3_ADD_467_U167 , P3_ADD_467_U168 , P3_ADD_467_U169 , P3_ADD_467_U170 , P3_ADD_467_U171 , P3_ADD_467_U172 , P3_ADD_467_U173 , P3_ADD_467_U174;
wire P3_ADD_467_U175 , P3_ADD_467_U176 , P3_ADD_467_U177 , P3_ADD_467_U178 , P3_ADD_467_U179 , P3_ADD_467_U180 , P3_ADD_467_U181 , P3_ADD_467_U182 , P3_ADD_430_U4 , P3_ADD_430_U5;
wire P3_ADD_430_U6 , P3_ADD_430_U7 , P3_ADD_430_U8 , P3_ADD_430_U9 , P3_ADD_430_U10 , P3_ADD_430_U11 , P3_ADD_430_U12 , P3_ADD_430_U13 , P3_ADD_430_U14 , P3_ADD_430_U15;
wire P3_ADD_430_U16 , P3_ADD_430_U17 , P3_ADD_430_U18 , P3_ADD_430_U19 , P3_ADD_430_U20 , P3_ADD_430_U21 , P3_ADD_430_U22 , P3_ADD_430_U23 , P3_ADD_430_U24 , P3_ADD_430_U25;
wire P3_ADD_430_U26 , P3_ADD_430_U27 , P3_ADD_430_U28 , P3_ADD_430_U29 , P3_ADD_430_U30 , P3_ADD_430_U31 , P3_ADD_430_U32 , P3_ADD_430_U33 , P3_ADD_430_U34 , P3_ADD_430_U35;
wire P3_ADD_430_U36 , P3_ADD_430_U37 , P3_ADD_430_U38 , P3_ADD_430_U39 , P3_ADD_430_U40 , P3_ADD_430_U41 , P3_ADD_430_U42 , P3_ADD_430_U43 , P3_ADD_430_U44 , P3_ADD_430_U45;
wire P3_ADD_430_U46 , P3_ADD_430_U47 , P3_ADD_430_U48 , P3_ADD_430_U49 , P3_ADD_430_U50 , P3_ADD_430_U51 , P3_ADD_430_U52 , P3_ADD_430_U53 , P3_ADD_430_U54 , P3_ADD_430_U55;
wire P3_ADD_430_U56 , P3_ADD_430_U57 , P3_ADD_430_U58 , P3_ADD_430_U59 , P3_ADD_430_U60 , P3_ADD_430_U61 , P3_ADD_430_U62 , P3_ADD_430_U63 , P3_ADD_430_U64 , P3_ADD_430_U65;
wire P3_ADD_430_U66 , P3_ADD_430_U67 , P3_ADD_430_U68 , P3_ADD_430_U69 , P3_ADD_430_U70 , P3_ADD_430_U71 , P3_ADD_430_U72 , P3_ADD_430_U73 , P3_ADD_430_U74 , P3_ADD_430_U75;
wire P3_ADD_430_U76 , P3_ADD_430_U77 , P3_ADD_430_U78 , P3_ADD_430_U79 , P3_ADD_430_U80 , P3_ADD_430_U81 , P3_ADD_430_U82 , P3_ADD_430_U83 , P3_ADD_430_U84 , P3_ADD_430_U85;
wire P3_ADD_430_U86 , P3_ADD_430_U87 , P3_ADD_430_U88 , P3_ADD_430_U89 , P3_ADD_430_U90 , P3_ADD_430_U91 , P3_ADD_430_U92 , P3_ADD_430_U93 , P3_ADD_430_U94 , P3_ADD_430_U95;
wire P3_ADD_430_U96 , P3_ADD_430_U97 , P3_ADD_430_U98 , P3_ADD_430_U99 , P3_ADD_430_U100 , P3_ADD_430_U101 , P3_ADD_430_U102 , P3_ADD_430_U103 , P3_ADD_430_U104 , P3_ADD_430_U105;
wire P3_ADD_430_U106 , P3_ADD_430_U107 , P3_ADD_430_U108 , P3_ADD_430_U109 , P3_ADD_430_U110 , P3_ADD_430_U111 , P3_ADD_430_U112 , P3_ADD_430_U113 , P3_ADD_430_U114 , P3_ADD_430_U115;
wire P3_ADD_430_U116 , P3_ADD_430_U117 , P3_ADD_430_U118 , P3_ADD_430_U119 , P3_ADD_430_U120 , P3_ADD_430_U121 , P3_ADD_430_U122 , P3_ADD_430_U123 , P3_ADD_430_U124 , P3_ADD_430_U125;
wire P3_ADD_430_U126 , P3_ADD_430_U127 , P3_ADD_430_U128 , P3_ADD_430_U129 , P3_ADD_430_U130 , P3_ADD_430_U131 , P3_ADD_430_U132 , P3_ADD_430_U133 , P3_ADD_430_U134 , P3_ADD_430_U135;
wire P3_ADD_430_U136 , P3_ADD_430_U137 , P3_ADD_430_U138 , P3_ADD_430_U139 , P3_ADD_430_U140 , P3_ADD_430_U141 , P3_ADD_430_U142 , P3_ADD_430_U143 , P3_ADD_430_U144 , P3_ADD_430_U145;
wire P3_ADD_430_U146 , P3_ADD_430_U147 , P3_ADD_430_U148 , P3_ADD_430_U149 , P3_ADD_430_U150 , P3_ADD_430_U151 , P3_ADD_430_U152 , P3_ADD_430_U153 , P3_ADD_430_U154 , P3_ADD_430_U155;
wire P3_ADD_430_U156 , P3_ADD_430_U157 , P3_ADD_430_U158 , P3_ADD_430_U159 , P3_ADD_430_U160 , P3_ADD_430_U161 , P3_ADD_430_U162 , P3_ADD_430_U163 , P3_ADD_430_U164 , P3_ADD_430_U165;
wire P3_ADD_430_U166 , P3_ADD_430_U167 , P3_ADD_430_U168 , P3_ADD_430_U169 , P3_ADD_430_U170 , P3_ADD_430_U171 , P3_ADD_430_U172 , P3_ADD_430_U173 , P3_ADD_430_U174 , P3_ADD_430_U175;
wire P3_ADD_430_U176 , P3_ADD_430_U177 , P3_ADD_430_U178 , P3_ADD_430_U179 , P3_ADD_430_U180 , P3_ADD_430_U181 , P3_ADD_430_U182 , P3_ADD_380_U5 , P3_ADD_380_U6 , P3_ADD_380_U7;
wire P3_ADD_380_U8 , P3_ADD_380_U9 , P3_ADD_380_U10 , P3_ADD_380_U11 , P3_ADD_380_U12 , P3_ADD_380_U13 , P3_ADD_380_U14 , P3_ADD_380_U15 , P3_ADD_380_U16 , P3_ADD_380_U17;
wire P3_ADD_380_U18 , P3_ADD_380_U19 , P3_ADD_380_U20 , P3_ADD_380_U21 , P3_ADD_380_U22 , P3_ADD_380_U23 , P3_ADD_380_U24 , P3_ADD_380_U25 , P3_ADD_380_U26 , P3_ADD_380_U27;
wire P3_ADD_380_U28 , P3_ADD_380_U29 , P3_ADD_380_U30 , P3_ADD_380_U31 , P3_ADD_380_U32 , P3_ADD_380_U33 , P3_ADD_380_U34 , P3_ADD_380_U35 , P3_ADD_380_U36 , P3_ADD_380_U37;
wire P3_ADD_380_U38 , P3_ADD_380_U39 , P3_ADD_380_U40 , P3_ADD_380_U41 , P3_ADD_380_U42 , P3_ADD_380_U43 , P3_ADD_380_U44 , P3_ADD_380_U45 , P3_ADD_380_U46 , P3_ADD_380_U47;
wire P3_ADD_380_U48 , P3_ADD_380_U49 , P3_ADD_380_U50 , P3_ADD_380_U51 , P3_ADD_380_U52 , P3_ADD_380_U53 , P3_ADD_380_U54 , P3_ADD_380_U55 , P3_ADD_380_U56 , P3_ADD_380_U57;
wire P3_ADD_380_U58 , P3_ADD_380_U59 , P3_ADD_380_U60 , P3_ADD_380_U61 , P3_ADD_380_U62 , P3_ADD_380_U63 , P3_ADD_380_U64 , P3_ADD_380_U65 , P3_ADD_380_U66 , P3_ADD_380_U67;
wire P3_ADD_380_U68 , P3_ADD_380_U69 , P3_ADD_380_U70 , P3_ADD_380_U71 , P3_ADD_380_U72 , P3_ADD_380_U73 , P3_ADD_380_U74 , P3_ADD_380_U75 , P3_ADD_380_U76 , P3_ADD_380_U77;
wire P3_ADD_380_U78 , P3_ADD_380_U79 , P3_ADD_380_U80 , P3_ADD_380_U81 , P3_ADD_380_U82 , P3_ADD_380_U83 , P3_ADD_380_U84 , P3_ADD_380_U85 , P3_ADD_380_U86 , P3_ADD_380_U87;
wire P3_ADD_380_U88 , P3_ADD_380_U89 , P3_ADD_380_U90 , P3_ADD_380_U91 , P3_ADD_380_U92 , P3_ADD_380_U93 , P3_ADD_380_U94 , P3_ADD_380_U95 , P3_ADD_380_U96 , P3_ADD_380_U97;
wire P3_ADD_380_U98 , P3_ADD_380_U99 , P3_ADD_380_U100 , P3_ADD_380_U101 , P3_ADD_380_U102 , P3_ADD_380_U103 , P3_ADD_380_U104 , P3_ADD_380_U105 , P3_ADD_380_U106 , P3_ADD_380_U107;
wire P3_ADD_380_U108 , P3_ADD_380_U109 , P3_ADD_380_U110 , P3_ADD_380_U111 , P3_ADD_380_U112 , P3_ADD_380_U113 , P3_ADD_380_U114 , P3_ADD_380_U115 , P3_ADD_380_U116 , P3_ADD_380_U117;
wire P3_ADD_380_U118 , P3_ADD_380_U119 , P3_ADD_380_U120 , P3_ADD_380_U121 , P3_ADD_380_U122 , P3_ADD_380_U123 , P3_ADD_380_U124 , P3_ADD_380_U125 , P3_ADD_380_U126 , P3_ADD_380_U127;
wire P3_ADD_380_U128 , P3_ADD_380_U129 , P3_ADD_380_U130 , P3_ADD_380_U131 , P3_ADD_380_U132 , P3_ADD_380_U133 , P3_ADD_380_U134 , P3_ADD_380_U135 , P3_ADD_380_U136 , P3_ADD_380_U137;
wire P3_ADD_380_U138 , P3_ADD_380_U139 , P3_ADD_380_U140 , P3_ADD_380_U141 , P3_ADD_380_U142 , P3_ADD_380_U143 , P3_ADD_380_U144 , P3_ADD_380_U145 , P3_ADD_380_U146 , P3_ADD_380_U147;
wire P3_ADD_380_U148 , P3_ADD_380_U149 , P3_ADD_380_U150 , P3_ADD_380_U151 , P3_ADD_380_U152 , P3_ADD_380_U153 , P3_ADD_380_U154 , P3_ADD_380_U155 , P3_ADD_380_U156 , P3_ADD_380_U157;
wire P3_ADD_380_U158 , P3_ADD_380_U159 , P3_ADD_380_U160 , P3_ADD_380_U161 , P3_ADD_380_U162 , P3_ADD_380_U163 , P3_ADD_380_U164 , P3_ADD_380_U165 , P3_ADD_380_U166 , P3_ADD_380_U167;
wire P3_ADD_380_U168 , P3_ADD_380_U169 , P3_ADD_380_U170 , P3_ADD_380_U171 , P3_ADD_380_U172 , P3_ADD_380_U173 , P3_ADD_380_U174 , P3_ADD_380_U175 , P3_ADD_380_U176 , P3_ADD_380_U177;
wire P3_ADD_380_U178 , P3_ADD_380_U179 , P3_ADD_380_U180 , P3_ADD_380_U181 , P3_ADD_380_U182 , P3_ADD_380_U183 , P3_ADD_380_U184 , P3_ADD_380_U185 , P3_ADD_380_U186 , P3_ADD_380_U187;
wire P3_ADD_380_U188 , P3_ADD_380_U189 , P3_GTE_370_U6 , P3_GTE_370_U7 , P3_GTE_370_U8 , P3_GTE_370_U9 , P3_ADD_344_U5 , P3_ADD_344_U6 , P3_ADD_344_U7 , P3_ADD_344_U8;
wire P3_ADD_344_U9 , P3_ADD_344_U10 , P3_ADD_344_U11 , P3_ADD_344_U12 , P3_ADD_344_U13 , P3_ADD_344_U14 , P3_ADD_344_U15 , P3_ADD_344_U16 , P3_ADD_344_U17 , P3_ADD_344_U18;
wire P3_ADD_344_U19 , P3_ADD_344_U20 , P3_ADD_344_U21 , P3_ADD_344_U22 , P3_ADD_344_U23 , P3_ADD_344_U24 , P3_ADD_344_U25 , P3_ADD_344_U26 , P3_ADD_344_U27 , P3_ADD_344_U28;
wire P3_ADD_344_U29 , P3_ADD_344_U30 , P3_ADD_344_U31 , P3_ADD_344_U32 , P3_ADD_344_U33 , P3_ADD_344_U34 , P3_ADD_344_U35 , P3_ADD_344_U36 , P3_ADD_344_U37 , P3_ADD_344_U38;
wire P3_ADD_344_U39 , P3_ADD_344_U40 , P3_ADD_344_U41 , P3_ADD_344_U42 , P3_ADD_344_U43 , P3_ADD_344_U44 , P3_ADD_344_U45 , P3_ADD_344_U46 , P3_ADD_344_U47 , P3_ADD_344_U48;
wire P3_ADD_344_U49 , P3_ADD_344_U50 , P3_ADD_344_U51 , P3_ADD_344_U52 , P3_ADD_344_U53 , P3_ADD_344_U54 , P3_ADD_344_U55 , P3_ADD_344_U56 , P3_ADD_344_U57 , P3_ADD_344_U58;
wire P3_ADD_344_U59 , P3_ADD_344_U60 , P3_ADD_344_U61 , P3_ADD_344_U62 , P3_ADD_344_U63 , P3_ADD_344_U64 , P3_ADD_344_U65 , P3_ADD_344_U66 , P3_ADD_344_U67 , P3_ADD_344_U68;
wire P3_ADD_344_U69 , P3_ADD_344_U70 , P3_ADD_344_U71 , P3_ADD_344_U72 , P3_ADD_344_U73 , P3_ADD_344_U74 , P3_ADD_344_U75 , P3_ADD_344_U76 , P3_ADD_344_U77 , P3_ADD_344_U78;
wire P3_ADD_344_U79 , P3_ADD_344_U80 , P3_ADD_344_U81 , P3_ADD_344_U82 , P3_ADD_344_U83 , P3_ADD_344_U84 , P3_ADD_344_U85 , P3_ADD_344_U86 , P3_ADD_344_U87 , P3_ADD_344_U88;
wire P3_ADD_344_U89 , P3_ADD_344_U90 , P3_ADD_344_U91 , P3_ADD_344_U92 , P3_ADD_344_U93 , P3_ADD_344_U94 , P3_ADD_344_U95 , P3_ADD_344_U96 , P3_ADD_344_U97 , P3_ADD_344_U98;
wire P3_ADD_344_U99 , P3_ADD_344_U100 , P3_ADD_344_U101 , P3_ADD_344_U102 , P3_ADD_344_U103 , P3_ADD_344_U104 , P3_ADD_344_U105 , P3_ADD_344_U106 , P3_ADD_344_U107 , P3_ADD_344_U108;
wire P3_ADD_344_U109 , P3_ADD_344_U110 , P3_ADD_344_U111 , P3_ADD_344_U112 , P3_ADD_344_U113 , P3_ADD_344_U114 , P3_ADD_344_U115 , P3_ADD_344_U116 , P3_ADD_344_U117 , P3_ADD_344_U118;
wire P3_ADD_344_U119 , P3_ADD_344_U120 , P3_ADD_344_U121 , P3_ADD_344_U122 , P3_ADD_344_U123 , P3_ADD_344_U124 , P3_ADD_344_U125 , P3_ADD_344_U126 , P3_ADD_344_U127 , P3_ADD_344_U128;
wire P3_ADD_344_U129 , P3_ADD_344_U130 , P3_ADD_344_U131 , P3_ADD_344_U132 , P3_ADD_344_U133 , P3_ADD_344_U134 , P3_ADD_344_U135 , P3_ADD_344_U136 , P3_ADD_344_U137 , P3_ADD_344_U138;
wire P3_ADD_344_U139 , P3_ADD_344_U140 , P3_ADD_344_U141 , P3_ADD_344_U142 , P3_ADD_344_U143 , P3_ADD_344_U144 , P3_ADD_344_U145 , P3_ADD_344_U146 , P3_ADD_344_U147 , P3_ADD_344_U148;
wire P3_ADD_344_U149 , P3_ADD_344_U150 , P3_ADD_344_U151 , P3_ADD_344_U152 , P3_ADD_344_U153 , P3_ADD_344_U154 , P3_ADD_344_U155 , P3_ADD_344_U156 , P3_ADD_344_U157 , P3_ADD_344_U158;
wire P3_ADD_344_U159 , P3_ADD_344_U160 , P3_ADD_344_U161 , P3_ADD_344_U162 , P3_ADD_344_U163 , P3_ADD_344_U164 , P3_ADD_344_U165 , P3_ADD_344_U166 , P3_ADD_344_U167 , P3_ADD_344_U168;
wire P3_ADD_344_U169 , P3_ADD_344_U170 , P3_ADD_344_U171 , P3_ADD_344_U172 , P3_ADD_344_U173 , P3_ADD_344_U174 , P3_ADD_344_U175 , P3_ADD_344_U176 , P3_ADD_344_U177 , P3_ADD_344_U178;
wire P3_ADD_344_U179 , P3_ADD_344_U180 , P3_ADD_344_U181 , P3_ADD_344_U182 , P3_ADD_344_U183 , P3_ADD_344_U184 , P3_ADD_344_U185 , P3_ADD_344_U186 , P3_ADD_344_U187 , P3_ADD_344_U188;
wire P3_ADD_344_U189 , P3_LT_563_U6 , P3_LT_563_U7 , P3_LT_563_U8 , P3_LT_563_U9 , P3_LT_563_U10 , P3_LT_563_U11 , P3_LT_563_U12 , P3_LT_563_U13 , P3_LT_563_U14;
wire P3_LT_563_U15 , P3_LT_563_U16 , P3_LT_563_U17 , P3_LT_563_U18 , P3_LT_563_U19 , P3_LT_563_U20 , P3_LT_563_U21 , P3_LT_563_U22 , P3_LT_563_U23 , P3_LT_563_U24;
wire P3_LT_563_U25 , P3_LT_563_U26 , P3_LT_563_U27 , P3_LT_563_U28 , P3_ADD_339_U4 , P3_ADD_339_U5 , P3_ADD_339_U6 , P3_ADD_339_U7 , P3_ADD_339_U8 , P3_ADD_339_U9;
wire P3_ADD_339_U10 , P3_ADD_339_U11 , P3_ADD_339_U12 , P3_ADD_339_U13 , P3_ADD_339_U14 , P3_ADD_339_U15 , P3_ADD_339_U16 , P3_ADD_339_U17 , P3_ADD_339_U18 , P3_ADD_339_U19;
wire P3_ADD_339_U20 , P3_ADD_339_U21 , P3_ADD_339_U22 , P3_ADD_339_U23 , P3_ADD_339_U24 , P3_ADD_339_U25 , P3_ADD_339_U26 , P3_ADD_339_U27 , P3_ADD_339_U28 , P3_ADD_339_U29;
wire P3_ADD_339_U30 , P3_ADD_339_U31 , P3_ADD_339_U32 , P3_ADD_339_U33 , P3_ADD_339_U34 , P3_ADD_339_U35 , P3_ADD_339_U36 , P3_ADD_339_U37 , P3_ADD_339_U38 , P3_ADD_339_U39;
wire P3_ADD_339_U40 , P3_ADD_339_U41 , P3_ADD_339_U42 , P3_ADD_339_U43 , P3_ADD_339_U44 , P3_ADD_339_U45 , P3_ADD_339_U46 , P3_ADD_339_U47 , P3_ADD_339_U48 , P3_ADD_339_U49;
wire P3_ADD_339_U50 , P3_ADD_339_U51 , P3_ADD_339_U52 , P3_ADD_339_U53 , P3_ADD_339_U54 , P3_ADD_339_U55 , P3_ADD_339_U56 , P3_ADD_339_U57 , P3_ADD_339_U58 , P3_ADD_339_U59;
wire P3_ADD_339_U60 , P3_ADD_339_U61 , P3_ADD_339_U62 , P3_ADD_339_U63 , P3_ADD_339_U64 , P3_ADD_339_U65 , P3_ADD_339_U66 , P3_ADD_339_U67 , P3_ADD_339_U68 , P3_ADD_339_U69;
wire P3_ADD_339_U70 , P3_ADD_339_U71 , P3_ADD_339_U72 , P3_ADD_339_U73 , P3_ADD_339_U74 , P3_ADD_339_U75 , P3_ADD_339_U76 , P3_ADD_339_U77 , P3_ADD_339_U78 , P3_ADD_339_U79;
wire P3_ADD_339_U80 , P3_ADD_339_U81 , P3_ADD_339_U82 , P3_ADD_339_U83 , P3_ADD_339_U84 , P3_ADD_339_U85 , P3_ADD_339_U86 , P3_ADD_339_U87 , P3_ADD_339_U88 , P3_ADD_339_U89;
wire P3_ADD_339_U90 , P3_ADD_339_U91 , P3_ADD_339_U92 , P3_ADD_339_U93 , P3_ADD_339_U94 , P3_ADD_339_U95 , P3_ADD_339_U96 , P3_ADD_339_U97 , P3_ADD_339_U98 , P3_ADD_339_U99;
wire P3_ADD_339_U100 , P3_ADD_339_U101 , P3_ADD_339_U102 , P3_ADD_339_U103 , P3_ADD_339_U104 , P3_ADD_339_U105 , P3_ADD_339_U106 , P3_ADD_339_U107 , P3_ADD_339_U108 , P3_ADD_339_U109;
wire P3_ADD_339_U110 , P3_ADD_339_U111 , P3_ADD_339_U112 , P3_ADD_339_U113 , P3_ADD_339_U114 , P3_ADD_339_U115 , P3_ADD_339_U116 , P3_ADD_339_U117 , P3_ADD_339_U118 , P3_ADD_339_U119;
wire P3_ADD_339_U120 , P3_ADD_339_U121 , P3_ADD_339_U122 , P3_ADD_339_U123 , P3_ADD_339_U124 , P3_ADD_339_U125 , P3_ADD_339_U126 , P3_ADD_339_U127 , P3_ADD_339_U128 , P3_ADD_339_U129;
wire P3_ADD_339_U130 , P3_ADD_339_U131 , P3_ADD_339_U132 , P3_ADD_339_U133 , P3_ADD_339_U134 , P3_ADD_339_U135 , P3_ADD_339_U136 , P3_ADD_339_U137 , P3_ADD_339_U138 , P3_ADD_339_U139;
wire P3_ADD_339_U140 , P3_ADD_339_U141 , P3_ADD_339_U142 , P3_ADD_339_U143 , P3_ADD_339_U144 , P3_ADD_339_U145 , P3_ADD_339_U146 , P3_ADD_339_U147 , P3_ADD_339_U148 , P3_ADD_339_U149;
wire P3_ADD_339_U150 , P3_ADD_339_U151 , P3_ADD_339_U152 , P3_ADD_339_U153 , P3_ADD_339_U154 , P3_ADD_339_U155 , P3_ADD_339_U156 , P3_ADD_339_U157 , P3_ADD_339_U158 , P3_ADD_339_U159;
wire P3_ADD_339_U160 , P3_ADD_339_U161 , P3_ADD_339_U162 , P3_ADD_339_U163 , P3_ADD_339_U164 , P3_ADD_339_U165 , P3_ADD_339_U166 , P3_ADD_339_U167 , P3_ADD_339_U168 , P3_ADD_339_U169;
wire P3_ADD_339_U170 , P3_ADD_339_U171 , P3_ADD_339_U172 , P3_ADD_339_U173 , P3_ADD_339_U174 , P3_ADD_339_U175 , P3_ADD_339_U176 , P3_ADD_339_U177 , P3_ADD_339_U178 , P3_ADD_339_U179;
wire P3_ADD_339_U180 , P3_ADD_339_U181 , P3_ADD_339_U182 , P3_ADD_360_U4 , P3_ADD_360_U5 , P3_ADD_360_U6 , P3_ADD_360_U7 , P3_ADD_360_U8 , P3_ADD_360_U9 , P3_ADD_360_U10;
wire P3_ADD_360_U11 , P3_ADD_360_U12 , P3_ADD_360_U13 , P3_ADD_360_U14 , P3_ADD_360_U15 , P3_ADD_360_U16 , P3_ADD_360_U17 , P3_ADD_360_U18 , P3_ADD_360_U19 , P3_ADD_360_U20;
wire P3_ADD_360_U21 , P3_ADD_360_U22 , P3_ADD_360_U23 , P3_ADD_360_U24 , P3_ADD_360_U25 , P3_ADD_360_U26 , P3_ADD_360_U27 , P3_ADD_360_U28 , P3_ADD_360_U29 , P3_ADD_360_U30;
wire P3_ADD_360_U31 , P3_ADD_360_U32 , P3_ADD_360_U33 , P3_ADD_360_U34 , P3_ADD_360_U35 , P3_ADD_360_U36 , P3_ADD_360_U37 , P3_ADD_360_U38 , P3_ADD_360_U39 , P3_ADD_360_U40;
wire P3_LTE_597_U6 , P3_SUB_580_U6 , P3_SUB_580_U7 , P3_SUB_580_U8 , P3_SUB_580_U9 , P3_SUB_580_U10 , P3_LT_589_U6 , P3_LT_589_U7 , P3_LT_589_U8 , P3_ADD_541_U4;
wire P3_ADD_541_U5 , P3_ADD_541_U6 , P3_ADD_541_U7 , P3_ADD_541_U8 , P3_ADD_541_U9 , P3_ADD_541_U10 , P3_ADD_541_U11 , P3_ADD_541_U12 , P3_ADD_541_U13 , P3_ADD_541_U14;
wire P3_ADD_541_U15 , P3_ADD_541_U16 , P3_ADD_541_U17 , P3_ADD_541_U18 , P3_ADD_541_U19 , P3_ADD_541_U20 , P3_ADD_541_U21 , P3_ADD_541_U22 , P3_ADD_541_U23 , P3_ADD_541_U24;
wire P3_ADD_541_U25 , P3_ADD_541_U26 , P3_ADD_541_U27 , P3_ADD_541_U28 , P3_ADD_541_U29 , P3_ADD_541_U30 , P3_ADD_541_U31 , P3_ADD_541_U32 , P3_ADD_541_U33 , P3_ADD_541_U34;
wire P3_ADD_541_U35 , P3_ADD_541_U36 , P3_ADD_541_U37 , P3_ADD_541_U38 , P3_ADD_541_U39 , P3_ADD_541_U40 , P3_ADD_541_U41 , P3_ADD_541_U42 , P3_ADD_541_U43 , P3_ADD_541_U44;
wire P3_ADD_541_U45 , P3_ADD_541_U46 , P3_ADD_541_U47 , P3_ADD_541_U48 , P3_ADD_541_U49 , P3_ADD_541_U50 , P3_ADD_541_U51 , P3_ADD_541_U52 , P3_ADD_541_U53 , P3_ADD_541_U54;
wire P3_ADD_541_U55 , P3_ADD_541_U56 , P3_ADD_541_U57 , P3_ADD_541_U58 , P3_ADD_541_U59 , P3_ADD_541_U60 , P3_ADD_541_U61 , P3_ADD_541_U62 , P3_ADD_541_U63 , P3_ADD_541_U64;
wire P3_ADD_541_U65 , P3_ADD_541_U66 , P3_ADD_541_U67 , P3_ADD_541_U68 , P3_ADD_541_U69 , P3_ADD_541_U70 , P3_ADD_541_U71 , P3_ADD_541_U72 , P3_ADD_541_U73 , P3_ADD_541_U74;
wire P3_ADD_541_U75 , P3_ADD_541_U76 , P3_ADD_541_U77 , P3_ADD_541_U78 , P3_ADD_541_U79 , P3_ADD_541_U80 , P3_ADD_541_U81 , P3_ADD_541_U82 , P3_ADD_541_U83 , P3_ADD_541_U84;
wire P3_ADD_541_U85 , P3_ADD_541_U86 , P3_ADD_541_U87 , P3_ADD_541_U88 , P3_ADD_541_U89 , P3_ADD_541_U90 , P3_ADD_541_U91 , P3_ADD_541_U92 , P3_ADD_541_U93 , P3_ADD_541_U94;
wire P3_ADD_541_U95 , P3_ADD_541_U96 , P3_ADD_541_U97 , P3_ADD_541_U98 , P3_ADD_541_U99 , P3_ADD_541_U100 , P3_ADD_541_U101 , P3_ADD_541_U102 , P3_ADD_541_U103 , P3_ADD_541_U104;
wire P3_ADD_541_U105 , P3_ADD_541_U106 , P3_ADD_541_U107 , P3_ADD_541_U108 , P3_ADD_541_U109 , P3_ADD_541_U110 , P3_ADD_541_U111 , P3_ADD_541_U112 , P3_ADD_541_U113 , P3_ADD_541_U114;
wire P3_ADD_541_U115 , P3_ADD_541_U116 , P3_ADD_541_U117 , P3_ADD_541_U118 , P3_ADD_541_U119 , P3_ADD_541_U120 , P3_ADD_541_U121 , P3_ADD_541_U122 , P3_ADD_541_U123 , P3_ADD_541_U124;
wire P3_ADD_541_U125 , P3_ADD_541_U126 , P3_ADD_541_U127 , P3_ADD_541_U128 , P3_ADD_541_U129 , P3_ADD_541_U130 , P3_ADD_541_U131 , P3_ADD_541_U132 , P3_ADD_541_U133 , P3_ADD_541_U134;
wire P3_ADD_541_U135 , P3_ADD_541_U136 , P3_ADD_541_U137 , P3_ADD_541_U138 , P3_ADD_541_U139 , P3_ADD_541_U140 , P3_ADD_541_U141 , P3_ADD_541_U142 , P3_ADD_541_U143 , P3_ADD_541_U144;
wire P3_ADD_541_U145 , P3_ADD_541_U146 , P3_ADD_541_U147 , P3_ADD_541_U148 , P3_ADD_541_U149 , P3_ADD_541_U150 , P3_ADD_541_U151 , P3_ADD_541_U152 , P3_ADD_541_U153 , P3_ADD_541_U154;
wire P3_ADD_541_U155 , P3_ADD_541_U156 , P3_ADD_541_U157 , P3_ADD_541_U158 , P3_ADD_541_U159 , P3_ADD_541_U160 , P3_ADD_541_U161 , P3_ADD_541_U162 , P3_ADD_541_U163 , P3_ADD_541_U164;
wire P3_ADD_541_U165 , P3_ADD_541_U166 , P3_ADD_541_U167 , P3_ADD_541_U168 , P3_ADD_541_U169 , P3_ADD_541_U170 , P3_ADD_541_U171 , P3_ADD_541_U172 , P3_ADD_541_U173 , P3_ADD_541_U174;
wire P3_ADD_541_U175 , P3_ADD_541_U176 , P3_ADD_541_U177 , P3_ADD_541_U178 , P3_ADD_541_U179 , P3_ADD_541_U180 , P3_ADD_541_U181 , P3_ADD_541_U182 , P3_SUB_355_U6 , P3_SUB_355_U7;
wire P3_SUB_355_U8 , P3_SUB_355_U9 , P3_SUB_355_U10 , P3_SUB_355_U11 , P3_SUB_355_U12 , P3_SUB_355_U13 , P3_SUB_355_U14 , P3_SUB_355_U15 , P3_SUB_355_U16 , P3_SUB_355_U17;
wire P3_SUB_355_U18 , P3_SUB_355_U19 , P3_SUB_355_U20 , P3_SUB_355_U21 , P3_SUB_355_U22 , P3_SUB_355_U23 , P3_SUB_355_U24 , P3_SUB_355_U25 , P3_SUB_355_U26 , P3_SUB_355_U27;
wire P3_SUB_355_U28 , P3_SUB_355_U29 , P3_SUB_355_U30 , P3_SUB_355_U31 , P3_SUB_355_U32 , P3_SUB_355_U33 , P3_SUB_355_U34 , P3_SUB_355_U35 , P3_SUB_355_U36 , P3_SUB_355_U37;
wire P3_SUB_355_U38 , P3_SUB_355_U39 , P3_SUB_355_U40 , P3_SUB_355_U41 , P3_SUB_355_U42 , P3_SUB_355_U43 , P3_SUB_355_U44 , P3_SUB_355_U45 , P3_SUB_355_U46 , P3_SUB_355_U47;
wire P3_SUB_355_U48 , P3_SUB_355_U49 , P3_SUB_355_U50 , P3_SUB_355_U51 , P3_SUB_355_U52 , P3_SUB_355_U53 , P3_SUB_355_U54 , P3_SUB_355_U55 , P3_SUB_355_U56 , P3_SUB_355_U57;
wire P3_SUB_355_U58 , P3_SUB_355_U59 , P3_SUB_355_U60 , P3_SUB_355_U61 , P3_SUB_355_U62 , P3_SUB_355_U63 , P3_SUB_355_U64 , P3_SUB_355_U65 , P3_SUB_355_U66 , P3_SUB_450_U6;
wire P3_SUB_450_U7 , P3_SUB_450_U8 , P3_SUB_450_U9 , P3_SUB_450_U10 , P3_SUB_450_U11 , P3_SUB_450_U12 , P3_SUB_450_U13 , P3_SUB_450_U14 , P3_SUB_450_U15 , P3_SUB_450_U16;
wire P3_SUB_450_U17 , P3_SUB_450_U18 , P3_SUB_450_U19 , P3_SUB_450_U20 , P3_SUB_450_U21 , P3_SUB_450_U22 , P3_SUB_450_U23 , P3_SUB_450_U24 , P3_SUB_450_U25 , P3_SUB_450_U26;
wire P3_SUB_450_U27 , P3_SUB_450_U28 , P3_SUB_450_U29 , P3_SUB_450_U30 , P3_SUB_450_U31 , P3_SUB_450_U32 , P3_SUB_450_U33 , P3_SUB_450_U34 , P3_SUB_450_U35 , P3_SUB_450_U36;
wire P3_SUB_450_U37 , P3_SUB_450_U38 , P3_SUB_450_U39 , P3_SUB_450_U40 , P3_SUB_450_U41 , P3_SUB_450_U42 , P3_SUB_450_U43 , P3_SUB_450_U44 , P3_SUB_450_U45 , P3_SUB_450_U46;
wire P3_SUB_450_U47 , P3_SUB_450_U48 , P3_SUB_450_U49 , P3_SUB_450_U50 , P3_SUB_450_U51 , P3_SUB_450_U52 , P3_SUB_450_U53 , P3_SUB_450_U54 , P3_SUB_450_U55 , P3_SUB_450_U56;
wire P3_SUB_450_U57 , P3_SUB_450_U58 , P3_SUB_450_U59 , P3_SUB_450_U60 , P3_SUB_450_U61 , P3_SUB_450_U62 , P3_SUB_450_U63 , P3_SUB_357_1258_U4 , P3_SUB_357_1258_U5 , P3_SUB_357_1258_U6;
wire P3_SUB_357_1258_U7 , P3_SUB_357_1258_U8 , P3_SUB_357_1258_U9 , P3_SUB_357_1258_U10 , P3_SUB_357_1258_U11 , P3_SUB_357_1258_U12 , P3_SUB_357_1258_U13 , P3_SUB_357_1258_U14 , P3_SUB_357_1258_U15 , P3_SUB_357_1258_U16;
wire P3_SUB_357_1258_U17 , P3_SUB_357_1258_U18 , P3_SUB_357_1258_U19 , P3_SUB_357_1258_U20 , P3_SUB_357_1258_U21 , P3_SUB_357_1258_U22 , P3_SUB_357_1258_U23 , P3_SUB_357_1258_U24 , P3_SUB_357_1258_U25 , P3_SUB_357_1258_U26;
wire P3_SUB_357_1258_U27 , P3_SUB_357_1258_U28 , P3_SUB_357_1258_U29 , P3_SUB_357_1258_U30 , P3_SUB_357_1258_U31 , P3_SUB_357_1258_U32 , P3_SUB_357_1258_U33 , P3_SUB_357_1258_U34 , P3_SUB_357_1258_U35 , P3_SUB_357_1258_U36;
wire P3_SUB_357_1258_U37 , P3_SUB_357_1258_U38 , P3_SUB_357_1258_U39 , P3_SUB_357_1258_U40 , P3_SUB_357_1258_U41 , P3_SUB_357_1258_U42 , P3_SUB_357_1258_U43 , P3_SUB_357_1258_U44 , P3_SUB_357_1258_U45 , P3_SUB_357_1258_U46;
wire P3_SUB_357_1258_U47 , P3_SUB_357_1258_U48 , P3_SUB_357_1258_U49 , P3_SUB_357_1258_U50 , P3_SUB_357_1258_U51 , P3_SUB_357_1258_U52 , P3_SUB_357_1258_U53 , P3_SUB_357_1258_U54 , P3_SUB_357_1258_U55 , P3_SUB_357_1258_U56;
wire P3_SUB_357_1258_U57 , P3_SUB_357_1258_U58 , P3_SUB_357_1258_U59 , P3_SUB_357_1258_U60 , P3_SUB_357_1258_U61 , P3_SUB_357_1258_U62 , P3_SUB_357_1258_U63 , P3_SUB_357_1258_U64 , P3_SUB_357_1258_U65 , P3_SUB_357_1258_U66;
wire P3_SUB_357_1258_U67 , P3_SUB_357_1258_U68 , P3_SUB_357_1258_U69 , P3_SUB_357_1258_U70 , P3_SUB_357_1258_U71 , P3_SUB_357_1258_U72 , P3_SUB_357_1258_U73 , P3_SUB_357_1258_U74 , P3_SUB_357_1258_U75 , P3_SUB_357_1258_U76;
wire P3_SUB_357_1258_U77 , P3_SUB_357_1258_U78 , P3_SUB_357_1258_U79 , P3_SUB_357_1258_U80 , P3_SUB_357_1258_U81 , P3_SUB_357_1258_U82 , P3_SUB_357_1258_U83 , P3_SUB_357_1258_U84 , P3_SUB_357_1258_U85 , P3_SUB_357_1258_U86;
wire P3_SUB_357_1258_U87 , P3_SUB_357_1258_U88 , P3_SUB_357_1258_U89 , P3_SUB_357_1258_U90 , P3_SUB_357_1258_U91 , P3_SUB_357_1258_U92 , P3_SUB_357_1258_U93 , P3_SUB_357_1258_U94 , P3_SUB_357_1258_U95 , P3_SUB_357_1258_U96;
wire P3_SUB_357_1258_U97 , P3_SUB_357_1258_U98 , P3_SUB_357_1258_U99 , P3_SUB_357_1258_U100 , P3_SUB_357_1258_U101 , P3_SUB_357_1258_U102 , P3_SUB_357_1258_U103 , P3_SUB_357_1258_U104 , P3_SUB_357_1258_U105 , P3_SUB_357_1258_U106;
wire P3_SUB_357_1258_U107 , P3_SUB_357_1258_U108 , P3_SUB_357_1258_U109 , P3_SUB_357_1258_U110 , P3_SUB_357_1258_U111 , P3_SUB_357_1258_U112 , P3_SUB_357_1258_U113 , P3_SUB_357_1258_U114 , P3_SUB_357_1258_U115 , P3_SUB_357_1258_U116;
wire P3_SUB_357_1258_U117 , P3_SUB_357_1258_U118 , P3_SUB_357_1258_U119 , P3_SUB_357_1258_U120 , P3_SUB_357_1258_U121 , P3_SUB_357_1258_U122 , P3_SUB_357_1258_U123 , P3_SUB_357_1258_U124 , P3_SUB_357_1258_U125 , P3_SUB_357_1258_U126;
wire P3_SUB_357_1258_U127 , P3_SUB_357_1258_U128 , P3_SUB_357_1258_U129 , P3_SUB_357_1258_U130 , P3_SUB_357_1258_U131 , P3_SUB_357_1258_U132 , P3_SUB_357_1258_U133 , P3_SUB_357_1258_U134 , P3_SUB_357_1258_U135 , P3_SUB_357_1258_U136;
wire P3_SUB_357_1258_U137 , P3_SUB_357_1258_U138 , P3_SUB_357_1258_U139 , P3_SUB_357_1258_U140 , P3_SUB_357_1258_U141 , P3_SUB_357_1258_U142 , P3_SUB_357_1258_U143 , P3_SUB_357_1258_U144 , P3_SUB_357_1258_U145 , P3_SUB_357_1258_U146;
wire P3_SUB_357_1258_U147 , P3_SUB_357_1258_U148 , P3_SUB_357_1258_U149 , P3_SUB_357_1258_U150 , P3_SUB_357_1258_U151 , P3_SUB_357_1258_U152 , P3_SUB_357_1258_U153 , P3_SUB_357_1258_U154 , P3_SUB_357_1258_U155 , P3_SUB_357_1258_U156;
wire P3_SUB_357_1258_U157 , P3_SUB_357_1258_U158 , P3_SUB_357_1258_U159 , P3_SUB_357_1258_U160 , P3_SUB_357_1258_U161 , P3_SUB_357_1258_U162 , P3_SUB_357_1258_U163 , P3_SUB_357_1258_U164 , P3_SUB_357_1258_U165 , P3_SUB_357_1258_U166;
wire P3_SUB_357_1258_U167 , P3_SUB_357_1258_U168 , P3_SUB_357_1258_U169 , P3_SUB_357_1258_U170 , P3_SUB_357_1258_U171 , P3_SUB_357_1258_U172 , P3_SUB_357_1258_U173 , P3_SUB_357_1258_U174 , P3_SUB_357_1258_U175 , P3_SUB_357_1258_U176;
wire P3_SUB_357_1258_U177 , P3_SUB_357_1258_U178 , P3_SUB_357_1258_U179 , P3_SUB_357_1258_U180 , P3_SUB_357_1258_U181 , P3_SUB_357_1258_U182 , P3_SUB_357_1258_U183 , P3_SUB_357_1258_U184 , P3_SUB_357_1258_U185 , P3_SUB_357_1258_U186;
wire P3_SUB_357_1258_U187 , P3_SUB_357_1258_U188 , P3_SUB_357_1258_U189 , P3_SUB_357_1258_U190 , P3_SUB_357_1258_U191 , P3_SUB_357_1258_U192 , P3_SUB_357_1258_U193 , P3_SUB_357_1258_U194 , P3_SUB_357_1258_U195 , P3_SUB_357_1258_U196;
wire P3_SUB_357_1258_U197 , P3_SUB_357_1258_U198 , P3_SUB_357_1258_U199 , P3_SUB_357_1258_U200 , P3_SUB_357_1258_U201 , P3_SUB_357_1258_U202 , P3_SUB_357_1258_U203 , P3_SUB_357_1258_U204 , P3_SUB_357_1258_U205 , P3_SUB_357_1258_U206;
wire P3_SUB_357_1258_U207 , P3_SUB_357_1258_U208 , P3_SUB_357_1258_U209 , P3_SUB_357_1258_U210 , P3_SUB_357_1258_U211 , P3_SUB_357_1258_U212 , P3_SUB_357_1258_U213 , P3_SUB_357_1258_U214 , P3_SUB_357_1258_U215 , P3_SUB_357_1258_U216;
wire P3_SUB_357_1258_U217 , P3_SUB_357_1258_U218 , P3_SUB_357_1258_U219 , P3_SUB_357_1258_U220 , P3_SUB_357_1258_U221 , P3_SUB_357_1258_U222 , P3_SUB_357_1258_U223 , P3_SUB_357_1258_U224 , P3_SUB_357_1258_U225 , P3_SUB_357_1258_U226;
wire P3_SUB_357_1258_U227 , P3_SUB_357_1258_U228 , P3_SUB_357_1258_U229 , P3_SUB_357_1258_U230 , P3_SUB_357_1258_U231 , P3_SUB_357_1258_U232 , P3_SUB_357_1258_U233 , P3_SUB_357_1258_U234 , P3_SUB_357_1258_U235 , P3_SUB_357_1258_U236;
wire P3_SUB_357_1258_U237 , P3_SUB_357_1258_U238 , P3_SUB_357_1258_U239 , P3_SUB_357_1258_U240 , P3_SUB_357_1258_U241 , P3_SUB_357_1258_U242 , P3_SUB_357_1258_U243 , P3_SUB_357_1258_U244 , P3_SUB_357_1258_U245 , P3_SUB_357_1258_U246;
wire P3_SUB_357_1258_U247 , P3_SUB_357_1258_U248 , P3_SUB_357_1258_U249 , P3_SUB_357_1258_U250 , P3_SUB_357_1258_U251 , P3_SUB_357_1258_U252 , P3_SUB_357_1258_U253 , P3_SUB_357_1258_U254 , P3_SUB_357_1258_U255 , P3_SUB_357_1258_U256;
wire P3_SUB_357_1258_U257 , P3_SUB_357_1258_U258 , P3_SUB_357_1258_U259 , P3_SUB_357_1258_U260 , P3_SUB_357_1258_U261 , P3_SUB_357_1258_U262 , P3_SUB_357_1258_U263 , P3_SUB_357_1258_U264 , P3_SUB_357_1258_U265 , P3_SUB_357_1258_U266;
wire P3_SUB_357_1258_U267 , P3_SUB_357_1258_U268 , P3_SUB_357_1258_U269 , P3_SUB_357_1258_U270 , P3_SUB_357_1258_U271 , P3_SUB_357_1258_U272 , P3_SUB_357_1258_U273 , P3_SUB_357_1258_U274 , P3_SUB_357_1258_U275 , P3_SUB_357_1258_U276;
wire P3_SUB_357_1258_U277 , P3_SUB_357_1258_U278 , P3_SUB_357_1258_U279 , P3_SUB_357_1258_U280 , P3_SUB_357_1258_U281 , P3_SUB_357_1258_U282 , P3_SUB_357_1258_U283 , P3_SUB_357_1258_U284 , P3_SUB_357_1258_U285 , P3_SUB_357_1258_U286;
wire P3_SUB_357_1258_U287 , P3_SUB_357_1258_U288 , P3_SUB_357_1258_U289 , P3_SUB_357_1258_U290 , P3_SUB_357_1258_U291 , P3_SUB_357_1258_U292 , P3_SUB_357_1258_U293 , P3_SUB_357_1258_U294 , P3_SUB_357_1258_U295 , P3_SUB_357_1258_U296;
wire P3_SUB_357_1258_U297 , P3_SUB_357_1258_U298 , P3_SUB_357_1258_U299 , P3_SUB_357_1258_U300 , P3_SUB_357_1258_U301 , P3_SUB_357_1258_U302 , P3_SUB_357_1258_U303 , P3_SUB_357_1258_U304 , P3_SUB_357_1258_U305 , P3_SUB_357_1258_U306;
wire P3_SUB_357_1258_U307 , P3_SUB_357_1258_U308 , P3_SUB_357_1258_U309 , P3_SUB_357_1258_U310 , P3_SUB_357_1258_U311 , P3_SUB_357_1258_U312 , P3_SUB_357_1258_U313 , P3_SUB_357_1258_U314 , P3_SUB_357_1258_U315 , P3_SUB_357_1258_U316;
wire P3_SUB_357_1258_U317 , P3_SUB_357_1258_U318 , P3_SUB_357_1258_U319 , P3_SUB_357_1258_U320 , P3_SUB_357_1258_U321 , P3_SUB_357_1258_U322 , P3_SUB_357_1258_U323 , P3_SUB_357_1258_U324 , P3_SUB_357_1258_U325 , P3_SUB_357_1258_U326;
wire P3_SUB_357_1258_U327 , P3_SUB_357_1258_U328 , P3_SUB_357_1258_U329 , P3_SUB_357_1258_U330 , P3_SUB_357_1258_U331 , P3_SUB_357_1258_U332 , P3_SUB_357_1258_U333 , P3_SUB_357_1258_U334 , P3_SUB_357_1258_U335 , P3_SUB_357_1258_U336;
wire P3_SUB_357_1258_U337 , P3_SUB_357_1258_U338 , P3_SUB_357_1258_U339 , P3_SUB_357_1258_U340 , P3_SUB_357_1258_U341 , P3_SUB_357_1258_U342 , P3_SUB_357_1258_U343 , P3_SUB_357_1258_U344 , P3_SUB_357_1258_U345 , P3_SUB_357_1258_U346;
wire P3_SUB_357_1258_U347 , P3_SUB_357_1258_U348 , P3_SUB_357_1258_U349 , P3_SUB_357_1258_U350 , P3_SUB_357_1258_U351 , P3_SUB_357_1258_U352 , P3_SUB_357_1258_U353 , P3_SUB_357_1258_U354 , P3_SUB_357_1258_U355 , P3_SUB_357_1258_U356;
wire P3_SUB_357_1258_U357 , P3_SUB_357_1258_U358 , P3_SUB_357_1258_U359 , P3_SUB_357_1258_U360 , P3_SUB_357_1258_U361 , P3_SUB_357_1258_U362 , P3_SUB_357_1258_U363 , P3_SUB_357_1258_U364 , P3_SUB_357_1258_U365 , P3_SUB_357_1258_U366;
wire P3_SUB_357_1258_U367 , P3_SUB_357_1258_U368 , P3_SUB_357_1258_U369 , P3_SUB_357_1258_U370 , P3_SUB_357_1258_U371 , P3_SUB_357_1258_U372 , P3_SUB_357_1258_U373 , P3_SUB_357_1258_U374 , P3_SUB_357_1258_U375 , P3_SUB_357_1258_U376;
wire P3_SUB_357_1258_U377 , P3_SUB_357_1258_U378 , P3_SUB_357_1258_U379 , P3_SUB_357_1258_U380 , P3_SUB_357_1258_U381 , P3_SUB_357_1258_U382 , P3_SUB_357_1258_U383 , P3_SUB_357_1258_U384 , P3_SUB_357_1258_U385 , P3_SUB_357_1258_U386;
wire P3_SUB_357_1258_U387 , P3_SUB_357_1258_U388 , P3_SUB_357_1258_U389 , P3_SUB_357_1258_U390 , P3_SUB_357_1258_U391 , P3_SUB_357_1258_U392 , P3_SUB_357_1258_U393 , P3_SUB_357_1258_U394 , P3_SUB_357_1258_U395 , P3_SUB_357_1258_U396;
wire P3_SUB_357_1258_U397 , P3_SUB_357_1258_U398 , P3_SUB_357_1258_U399 , P3_SUB_357_1258_U400 , P3_SUB_357_1258_U401 , P3_SUB_357_1258_U402 , P3_SUB_357_1258_U403 , P3_SUB_357_1258_U404 , P3_SUB_357_1258_U405 , P3_SUB_357_1258_U406;
wire P3_SUB_357_1258_U407 , P3_SUB_357_1258_U408 , P3_SUB_357_1258_U409 , P3_SUB_357_1258_U410 , P3_SUB_357_1258_U411 , P3_SUB_357_1258_U412 , P3_SUB_357_1258_U413 , P3_SUB_357_1258_U414 , P3_SUB_357_1258_U415 , P3_SUB_357_1258_U416;
wire P3_SUB_357_1258_U417 , P3_SUB_357_1258_U418 , P3_SUB_357_1258_U419 , P3_SUB_357_1258_U420 , P3_SUB_357_1258_U421 , P3_SUB_357_1258_U422 , P3_SUB_357_1258_U423 , P3_SUB_357_1258_U424 , P3_SUB_357_1258_U425 , P3_SUB_357_1258_U426;
wire P3_SUB_357_1258_U427 , P3_SUB_357_1258_U428 , P3_SUB_357_1258_U429 , P3_SUB_357_1258_U430 , P3_SUB_357_1258_U431 , P3_SUB_357_1258_U432 , P3_SUB_357_1258_U433 , P3_SUB_357_1258_U434 , P3_SUB_357_1258_U435 , P3_SUB_357_1258_U436;
wire P3_SUB_357_1258_U437 , P3_SUB_357_1258_U438 , P3_SUB_357_1258_U439 , P3_SUB_357_1258_U440 , P3_SUB_357_1258_U441 , P3_SUB_357_1258_U442 , P3_SUB_357_1258_U443 , P3_SUB_357_1258_U444 , P3_SUB_357_1258_U445 , P3_SUB_357_1258_U446;
wire P3_SUB_357_1258_U447 , P3_SUB_357_1258_U448 , P3_SUB_357_1258_U449 , P3_SUB_357_1258_U450 , P3_SUB_357_1258_U451 , P3_SUB_357_1258_U452 , P3_SUB_357_1258_U453 , P3_SUB_357_1258_U454 , P3_SUB_357_1258_U455 , P3_SUB_357_1258_U456;
wire P3_SUB_357_1258_U457 , P3_SUB_357_1258_U458 , P3_SUB_357_1258_U459 , P3_SUB_357_1258_U460 , P3_SUB_357_1258_U461 , P3_SUB_357_1258_U462 , P3_SUB_357_1258_U463 , P3_SUB_357_1258_U464 , P3_SUB_357_1258_U465 , P3_SUB_357_1258_U466;
wire P3_SUB_357_1258_U467 , P3_SUB_357_1258_U468 , P3_SUB_357_1258_U469 , P3_SUB_357_1258_U470 , P3_SUB_357_1258_U471 , P3_SUB_357_1258_U472 , P3_SUB_357_1258_U473 , P3_SUB_357_1258_U474 , P3_SUB_357_1258_U475 , P3_SUB_357_1258_U476;
wire P3_SUB_357_1258_U477 , P3_SUB_357_1258_U478 , P3_SUB_357_1258_U479 , P3_SUB_357_1258_U480 , P3_SUB_357_1258_U481 , P3_SUB_357_1258_U482 , P3_SUB_357_1258_U483 , P3_SUB_357_1258_U484 , P3_ADD_486_U5 , P3_ADD_486_U6;
wire P3_ADD_486_U7 , P3_ADD_486_U8 , P3_ADD_486_U9 , P3_ADD_486_U10 , P3_ADD_486_U11 , P3_ADD_486_U12 , P3_ADD_486_U13 , P3_ADD_486_U14 , P3_ADD_486_U15 , P3_ADD_486_U16;
wire P3_ADD_486_U17 , P3_ADD_486_U18 , P3_ADD_486_U19 , P3_ADD_486_U20 , P3_ADD_486_U21 , P3_ADD_486_U22 , P3_ADD_486_U23 , P3_ADD_486_U24 , P3_ADD_486_U25 , P3_ADD_486_U26;
wire P3_ADD_486_U27 , P3_ADD_486_U28 , P3_SUB_485_U6 , P3_SUB_485_U7 , P3_SUB_485_U8 , P3_SUB_485_U9 , P3_SUB_485_U10 , P3_SUB_485_U11 , P3_SUB_485_U12 , P3_SUB_485_U13;
wire P3_SUB_485_U14 , P3_SUB_485_U15 , P3_SUB_485_U16 , P3_SUB_485_U17 , P3_SUB_485_U18 , P3_SUB_485_U19 , P3_SUB_485_U20 , P3_SUB_485_U21 , P3_SUB_485_U22 , P3_SUB_485_U23;
wire P3_SUB_485_U24 , P3_SUB_485_U25 , P3_SUB_485_U26 , P3_SUB_485_U27 , P3_SUB_485_U28 , P3_SUB_485_U29 , P3_SUB_485_U30 , P3_SUB_485_U31 , P3_SUB_485_U32 , P3_SUB_485_U33;
wire P3_SUB_485_U34 , P3_SUB_485_U35 , P3_SUB_485_U36 , P3_SUB_485_U37 , P3_SUB_485_U38 , P3_SUB_485_U39 , P3_SUB_485_U40 , P3_SUB_485_U41 , P3_SUB_485_U42 , P3_SUB_485_U43;
wire P3_SUB_485_U44 , P3_SUB_485_U45 , P3_SUB_485_U46 , P3_SUB_485_U47 , P3_SUB_485_U48 , P3_SUB_485_U49 , P3_SUB_485_U50 , P3_SUB_485_U51 , P3_SUB_485_U52 , P3_SUB_485_U53;
wire P3_SUB_485_U54 , P3_SUB_485_U55 , P3_SUB_485_U56 , P3_SUB_485_U57 , P3_SUB_485_U58 , P3_SUB_485_U59 , P3_SUB_485_U60 , P3_SUB_485_U61 , P3_SUB_485_U62 , P3_SUB_485_U63;
wire P3_SUB_563_U6 , P3_SUB_563_U7 , P3_ADD_515_U4 , P3_ADD_515_U5 , P3_ADD_515_U6 , P3_ADD_515_U7 , P3_ADD_515_U8 , P3_ADD_515_U9 , P3_ADD_515_U10 , P3_ADD_515_U11;
wire P3_ADD_515_U12 , P3_ADD_515_U13 , P3_ADD_515_U14 , P3_ADD_515_U15 , P3_ADD_515_U16 , P3_ADD_515_U17 , P3_ADD_515_U18 , P3_ADD_515_U19 , P3_ADD_515_U20 , P3_ADD_515_U21;
wire P3_ADD_515_U22 , P3_ADD_515_U23 , P3_ADD_515_U24 , P3_ADD_515_U25 , P3_ADD_515_U26 , P3_ADD_515_U27 , P3_ADD_515_U28 , P3_ADD_515_U29 , P3_ADD_515_U30 , P3_ADD_515_U31;
wire P3_ADD_515_U32 , P3_ADD_515_U33 , P3_ADD_515_U34 , P3_ADD_515_U35 , P3_ADD_515_U36 , P3_ADD_515_U37 , P3_ADD_515_U38 , P3_ADD_515_U39 , P3_ADD_515_U40 , P3_ADD_515_U41;
wire P3_ADD_515_U42 , P3_ADD_515_U43 , P3_ADD_515_U44 , P3_ADD_515_U45 , P3_ADD_515_U46 , P3_ADD_515_U47 , P3_ADD_515_U48 , P3_ADD_515_U49 , P3_ADD_515_U50 , P3_ADD_515_U51;
wire P3_ADD_515_U52 , P3_ADD_515_U53 , P3_ADD_515_U54 , P3_ADD_515_U55 , P3_ADD_515_U56 , P3_ADD_515_U57 , P3_ADD_515_U58 , P3_ADD_515_U59 , P3_ADD_515_U60 , P3_ADD_515_U61;
wire P3_ADD_515_U62 , P3_ADD_515_U63 , P3_ADD_515_U64 , P3_ADD_515_U65 , P3_ADD_515_U66 , P3_ADD_515_U67 , P3_ADD_515_U68 , P3_ADD_515_U69 , P3_ADD_515_U70 , P3_ADD_515_U71;
wire P3_ADD_515_U72 , P3_ADD_515_U73 , P3_ADD_515_U74 , P3_ADD_515_U75 , P3_ADD_515_U76 , P3_ADD_515_U77 , P3_ADD_515_U78 , P3_ADD_515_U79 , P3_ADD_515_U80 , P3_ADD_515_U81;
wire P3_ADD_515_U82 , P3_ADD_515_U83 , P3_ADD_515_U84 , P3_ADD_515_U85 , P3_ADD_515_U86 , P3_ADD_515_U87 , P3_ADD_515_U88 , P3_ADD_515_U89 , P3_ADD_515_U90 , P3_ADD_515_U91;
wire P3_ADD_515_U92 , P3_ADD_515_U93 , P3_ADD_515_U94 , P3_ADD_515_U95 , P3_ADD_515_U96 , P3_ADD_515_U97 , P3_ADD_515_U98 , P3_ADD_515_U99 , P3_ADD_515_U100 , P3_ADD_515_U101;
wire P3_ADD_515_U102 , P3_ADD_515_U103 , P3_ADD_515_U104 , P3_ADD_515_U105 , P3_ADD_515_U106 , P3_ADD_515_U107 , P3_ADD_515_U108 , P3_ADD_515_U109 , P3_ADD_515_U110 , P3_ADD_515_U111;
wire P3_ADD_515_U112 , P3_ADD_515_U113 , P3_ADD_515_U114 , P3_ADD_515_U115 , P3_ADD_515_U116 , P3_ADD_515_U117 , P3_ADD_515_U118 , P3_ADD_515_U119 , P3_ADD_515_U120 , P3_ADD_515_U121;
wire P3_ADD_515_U122 , P3_ADD_515_U123 , P3_ADD_515_U124 , P3_ADD_515_U125 , P3_ADD_515_U126 , P3_ADD_515_U127 , P3_ADD_515_U128 , P3_ADD_515_U129 , P3_ADD_515_U130 , P3_ADD_515_U131;
wire P3_ADD_515_U132 , P3_ADD_515_U133 , P3_ADD_515_U134 , P3_ADD_515_U135 , P3_ADD_515_U136 , P3_ADD_515_U137 , P3_ADD_515_U138 , P3_ADD_515_U139 , P3_ADD_515_U140 , P3_ADD_515_U141;
wire P3_ADD_515_U142 , P3_ADD_515_U143 , P3_ADD_515_U144 , P3_ADD_515_U145 , P3_ADD_515_U146 , P3_ADD_515_U147 , P3_ADD_515_U148 , P3_ADD_515_U149 , P3_ADD_515_U150 , P3_ADD_515_U151;
wire P3_ADD_515_U152 , P3_ADD_515_U153 , P3_ADD_515_U154 , P3_ADD_515_U155 , P3_ADD_515_U156 , P3_ADD_515_U157 , P3_ADD_515_U158 , P3_ADD_515_U159 , P3_ADD_515_U160 , P3_ADD_515_U161;
wire P3_ADD_515_U162 , P3_ADD_515_U163 , P3_ADD_515_U164 , P3_ADD_515_U165 , P3_ADD_515_U166 , P3_ADD_515_U167 , P3_ADD_515_U168 , P3_ADD_515_U169 , P3_ADD_515_U170 , P3_ADD_515_U171;
wire P3_ADD_515_U172 , P3_ADD_515_U173 , P3_ADD_515_U174 , P3_ADD_515_U175 , P3_ADD_515_U176 , P3_ADD_515_U177 , P3_ADD_515_U178 , P3_ADD_515_U179 , P3_ADD_515_U180 , P3_ADD_515_U181;
wire P3_ADD_515_U182 , P3_ADD_394_U4 , P3_ADD_394_U5 , P3_ADD_394_U6 , P3_ADD_394_U7 , P3_ADD_394_U8 , P3_ADD_394_U9 , P3_ADD_394_U10 , P3_ADD_394_U11 , P3_ADD_394_U12;
wire P3_ADD_394_U13 , P3_ADD_394_U14 , P3_ADD_394_U15 , P3_ADD_394_U16 , P3_ADD_394_U17 , P3_ADD_394_U18 , P3_ADD_394_U19 , P3_ADD_394_U20 , P3_ADD_394_U21 , P3_ADD_394_U22;
wire P3_ADD_394_U23 , P3_ADD_394_U24 , P3_ADD_394_U25 , P3_ADD_394_U26 , P3_ADD_394_U27 , P3_ADD_394_U28 , P3_ADD_394_U29 , P3_ADD_394_U30 , P3_ADD_394_U31 , P3_ADD_394_U32;
wire P3_ADD_394_U33 , P3_ADD_394_U34 , P3_ADD_394_U35 , P3_ADD_394_U36 , P3_ADD_394_U37 , P3_ADD_394_U38 , P3_ADD_394_U39 , P3_ADD_394_U40 , P3_ADD_394_U41 , P3_ADD_394_U42;
wire P3_ADD_394_U43 , P3_ADD_394_U44 , P3_ADD_394_U45 , P3_ADD_394_U46 , P3_ADD_394_U47 , P3_ADD_394_U48 , P3_ADD_394_U49 , P3_ADD_394_U50 , P3_ADD_394_U51 , P3_ADD_394_U52;
wire P3_ADD_394_U53 , P3_ADD_394_U54 , P3_ADD_394_U55 , P3_ADD_394_U56 , P3_ADD_394_U57 , P3_ADD_394_U58 , P3_ADD_394_U59 , P3_ADD_394_U60 , P3_ADD_394_U61 , P3_ADD_394_U62;
wire P3_ADD_394_U63 , P3_ADD_394_U64 , P3_ADD_394_U65 , P3_ADD_394_U66 , P3_ADD_394_U67 , P3_ADD_394_U68 , P3_ADD_394_U69 , P3_ADD_394_U70 , P3_ADD_394_U71 , P3_ADD_394_U72;
wire P3_ADD_394_U73 , P3_ADD_394_U74 , P3_ADD_394_U75 , P3_ADD_394_U76 , P3_ADD_394_U77 , P3_ADD_394_U78 , P3_ADD_394_U79 , P3_ADD_394_U80 , P3_ADD_394_U81 , P3_ADD_394_U82;
wire P3_ADD_394_U83 , P3_ADD_394_U84 , P3_ADD_394_U85 , P3_ADD_394_U86 , P3_ADD_394_U87 , P3_ADD_394_U88 , P3_ADD_394_U89 , P3_ADD_394_U90 , P3_ADD_394_U91 , P3_ADD_394_U92;
wire P3_ADD_394_U93 , P3_ADD_394_U94 , P3_ADD_394_U95 , P3_ADD_394_U96 , P3_ADD_394_U97 , P3_ADD_394_U98 , P3_ADD_394_U99 , P3_ADD_394_U100 , P3_ADD_394_U101 , P3_ADD_394_U102;
wire P3_ADD_394_U103 , P3_ADD_394_U104 , P3_ADD_394_U105 , P3_ADD_394_U106 , P3_ADD_394_U107 , P3_ADD_394_U108 , P3_ADD_394_U109 , P3_ADD_394_U110 , P3_ADD_394_U111 , P3_ADD_394_U112;
wire P3_ADD_394_U113 , P3_ADD_394_U114 , P3_ADD_394_U115 , P3_ADD_394_U116 , P3_ADD_394_U117 , P3_ADD_394_U118 , P3_ADD_394_U119 , P3_ADD_394_U120 , P3_ADD_394_U121 , P3_ADD_394_U122;
wire P3_ADD_394_U123 , P3_ADD_394_U124 , P3_ADD_394_U125 , P3_ADD_394_U126 , P3_ADD_394_U127 , P3_ADD_394_U128 , P3_ADD_394_U129 , P3_ADD_394_U130 , P3_ADD_394_U131 , P3_ADD_394_U132;
wire P3_ADD_394_U133 , P3_ADD_394_U134 , P3_ADD_394_U135 , P3_ADD_394_U136 , P3_ADD_394_U137 , P3_ADD_394_U138 , P3_ADD_394_U139 , P3_ADD_394_U140 , P3_ADD_394_U141 , P3_ADD_394_U142;
wire P3_ADD_394_U143 , P3_ADD_394_U144 , P3_ADD_394_U145 , P3_ADD_394_U146 , P3_ADD_394_U147 , P3_ADD_394_U148 , P3_ADD_394_U149 , P3_ADD_394_U150 , P3_ADD_394_U151 , P3_ADD_394_U152;
wire P3_ADD_394_U153 , P3_ADD_394_U154 , P3_ADD_394_U155 , P3_ADD_394_U156 , P3_ADD_394_U157 , P3_ADD_394_U158 , P3_ADD_394_U159 , P3_ADD_394_U160 , P3_ADD_394_U161 , P3_ADD_394_U162;
wire P3_ADD_394_U163 , P3_ADD_394_U164 , P3_ADD_394_U165 , P3_ADD_394_U166 , P3_ADD_394_U167 , P3_ADD_394_U168 , P3_ADD_394_U169 , P3_ADD_394_U170 , P3_ADD_394_U171 , P3_ADD_394_U172;
wire P3_ADD_394_U173 , P3_ADD_394_U174 , P3_ADD_394_U175 , P3_ADD_394_U176 , P3_ADD_394_U177 , P3_ADD_394_U178 , P3_ADD_394_U179 , P3_ADD_394_U180 , P3_ADD_394_U181 , P3_ADD_394_U182;
wire P3_ADD_394_U183 , P3_ADD_394_U184 , P3_ADD_394_U185 , P3_ADD_394_U186 , P3_GTE_450_U6 , P3_GTE_450_U7 , P3_SUB_414_U6 , P3_SUB_414_U7 , P3_SUB_414_U8 , P3_SUB_414_U9;
wire P3_SUB_414_U10 , P3_SUB_414_U11 , P3_SUB_414_U12 , P3_SUB_414_U13 , P3_SUB_414_U14 , P3_SUB_414_U15 , P3_SUB_414_U16 , P3_SUB_414_U17 , P3_SUB_414_U18 , P3_SUB_414_U19;
wire P3_SUB_414_U20 , P3_SUB_414_U21 , P3_SUB_414_U22 , P3_SUB_414_U23 , P3_SUB_414_U24 , P3_SUB_414_U25 , P3_SUB_414_U26 , P3_SUB_414_U27 , P3_SUB_414_U28 , P3_SUB_414_U29;
wire P3_SUB_414_U30 , P3_SUB_414_U31 , P3_SUB_414_U32 , P3_SUB_414_U33 , P3_SUB_414_U34 , P3_SUB_414_U35 , P3_SUB_414_U36 , P3_SUB_414_U37 , P3_SUB_414_U38 , P3_SUB_414_U39;
wire P3_SUB_414_U40 , P3_SUB_414_U41 , P3_SUB_414_U42 , P3_SUB_414_U43 , P3_SUB_414_U44 , P3_SUB_414_U45 , P3_SUB_414_U46 , P3_SUB_414_U47 , P3_SUB_414_U48 , P3_SUB_414_U49;
wire P3_SUB_414_U50 , P3_SUB_414_U51 , P3_SUB_414_U52 , P3_SUB_414_U53 , P3_SUB_414_U54 , P3_SUB_414_U55 , P3_SUB_414_U56 , P3_SUB_414_U57 , P3_SUB_414_U58 , P3_SUB_414_U59;
wire P3_SUB_414_U60 , P3_SUB_414_U61 , P3_SUB_414_U62 , P3_SUB_414_U63 , P3_SUB_414_U64 , P3_SUB_414_U65 , P3_SUB_414_U66 , P3_SUB_414_U67 , P3_SUB_414_U68 , P3_SUB_414_U69;
wire P3_SUB_414_U70 , P3_SUB_414_U71 , P3_SUB_414_U72 , P3_SUB_414_U73 , P3_SUB_414_U74 , P3_SUB_414_U75 , P3_SUB_414_U76 , P3_SUB_414_U77 , P3_SUB_414_U78 , P3_SUB_414_U79;
wire P3_SUB_414_U80 , P3_SUB_414_U81 , P3_SUB_414_U82 , P3_SUB_414_U83 , P3_SUB_414_U84 , P3_SUB_414_U85 , P3_SUB_414_U86 , P3_SUB_414_U87 , P3_SUB_414_U88 , P3_SUB_414_U89;
wire P3_SUB_414_U90 , P3_SUB_414_U91 , P3_SUB_414_U92 , P3_SUB_414_U93 , P3_SUB_414_U94 , P3_SUB_414_U95 , P3_SUB_414_U96 , P3_SUB_414_U97 , P3_SUB_414_U98 , P3_SUB_414_U99;
wire P3_SUB_414_U100 , P3_SUB_414_U101 , P3_SUB_414_U102 , P3_SUB_414_U103 , P3_SUB_414_U104 , P3_SUB_414_U105 , P3_SUB_414_U106 , P3_SUB_414_U107 , P3_SUB_414_U108 , P3_SUB_414_U109;
wire P3_SUB_414_U110 , P3_SUB_414_U111 , P3_SUB_414_U112 , P3_SUB_414_U113 , P3_SUB_414_U114 , P3_SUB_414_U115 , P3_SUB_414_U116 , P3_SUB_414_U117 , P3_SUB_414_U118 , P3_SUB_414_U119;
wire P3_SUB_414_U120 , P3_SUB_414_U121 , P3_SUB_414_U122 , P3_SUB_414_U123 , P3_SUB_414_U124 , P3_SUB_414_U125 , P3_SUB_414_U126 , P3_SUB_414_U127 , P3_SUB_414_U128 , P3_SUB_414_U129;
wire P3_SUB_414_U130 , P3_SUB_414_U131 , P3_SUB_414_U132 , P3_SUB_414_U133 , P3_SUB_414_U134 , P3_SUB_414_U135 , P3_SUB_414_U136 , P3_SUB_414_U137 , P3_SUB_414_U138 , P3_SUB_414_U139;
wire P3_SUB_414_U140 , P3_SUB_414_U141 , P3_SUB_414_U142 , P3_SUB_414_U143 , P3_SUB_414_U144 , P3_SUB_414_U145 , P3_SUB_414_U146 , P3_SUB_414_U147 , P3_SUB_414_U148 , P3_SUB_414_U149;
wire P3_SUB_414_U150 , P3_SUB_414_U151 , P3_SUB_414_U152 , P3_SUB_414_U153 , P3_SUB_414_U154 , P3_SUB_414_U155 , P3_SUB_414_U156 , P3_SUB_414_U157 , P3_SUB_414_U158 , P3_SUB_414_U159;
wire P3_ADD_441_U4 , P3_ADD_441_U5 , P3_ADD_441_U6 , P3_ADD_441_U7 , P3_ADD_441_U8 , P3_ADD_441_U9 , P3_ADD_441_U10 , P3_ADD_441_U11 , P3_ADD_441_U12 , P3_ADD_441_U13;
wire P3_ADD_441_U14 , P3_ADD_441_U15 , P3_ADD_441_U16 , P3_ADD_441_U17 , P3_ADD_441_U18 , P3_ADD_441_U19 , P3_ADD_441_U20 , P3_ADD_441_U21 , P3_ADD_441_U22 , P3_ADD_441_U23;
wire P3_ADD_441_U24 , P3_ADD_441_U25 , P3_ADD_441_U26 , P3_ADD_441_U27 , P3_ADD_441_U28 , P3_ADD_441_U29 , P3_ADD_441_U30 , P3_ADD_441_U31 , P3_ADD_441_U32 , P3_ADD_441_U33;
wire P3_ADD_441_U34 , P3_ADD_441_U35 , P3_ADD_441_U36 , P3_ADD_441_U37 , P3_ADD_441_U38 , P3_ADD_441_U39 , P3_ADD_441_U40 , P3_ADD_441_U41 , P3_ADD_441_U42 , P3_ADD_441_U43;
wire P3_ADD_441_U44 , P3_ADD_441_U45 , P3_ADD_441_U46 , P3_ADD_441_U47 , P3_ADD_441_U48 , P3_ADD_441_U49 , P3_ADD_441_U50 , P3_ADD_441_U51 , P3_ADD_441_U52 , P3_ADD_441_U53;
wire P3_ADD_441_U54 , P3_ADD_441_U55 , P3_ADD_441_U56 , P3_ADD_441_U57 , P3_ADD_441_U58 , P3_ADD_441_U59 , P3_ADD_441_U60 , P3_ADD_441_U61 , P3_ADD_441_U62 , P3_ADD_441_U63;
wire P3_ADD_441_U64 , P3_ADD_441_U65 , P3_ADD_441_U66 , P3_ADD_441_U67 , P3_ADD_441_U68 , P3_ADD_441_U69 , P3_ADD_441_U70 , P3_ADD_441_U71 , P3_ADD_441_U72 , P3_ADD_441_U73;
wire P3_ADD_441_U74 , P3_ADD_441_U75 , P3_ADD_441_U76 , P3_ADD_441_U77 , P3_ADD_441_U78 , P3_ADD_441_U79 , P3_ADD_441_U80 , P3_ADD_441_U81 , P3_ADD_441_U82 , P3_ADD_441_U83;
wire P3_ADD_441_U84 , P3_ADD_441_U85 , P3_ADD_441_U86 , P3_ADD_441_U87 , P3_ADD_441_U88 , P3_ADD_441_U89 , P3_ADD_441_U90 , P3_ADD_441_U91 , P3_ADD_441_U92 , P3_ADD_441_U93;
wire P3_ADD_441_U94 , P3_ADD_441_U95 , P3_ADD_441_U96 , P3_ADD_441_U97 , P3_ADD_441_U98 , P3_ADD_441_U99 , P3_ADD_441_U100 , P3_ADD_441_U101 , P3_ADD_441_U102 , P3_ADD_441_U103;
wire P3_ADD_441_U104 , P3_ADD_441_U105 , P3_ADD_441_U106 , P3_ADD_441_U107 , P3_ADD_441_U108 , P3_ADD_441_U109 , P3_ADD_441_U110 , P3_ADD_441_U111 , P3_ADD_441_U112 , P3_ADD_441_U113;
wire P3_ADD_441_U114 , P3_ADD_441_U115 , P3_ADD_441_U116 , P3_ADD_441_U117 , P3_ADD_441_U118 , P3_ADD_441_U119 , P3_ADD_441_U120 , P3_ADD_441_U121 , P3_ADD_441_U122 , P3_ADD_441_U123;
wire P3_ADD_441_U124 , P3_ADD_441_U125 , P3_ADD_441_U126 , P3_ADD_441_U127 , P3_ADD_441_U128 , P3_ADD_441_U129 , P3_ADD_441_U130 , P3_ADD_441_U131 , P3_ADD_441_U132 , P3_ADD_441_U133;
wire P3_ADD_441_U134 , P3_ADD_441_U135 , P3_ADD_441_U136 , P3_ADD_441_U137 , P3_ADD_441_U138 , P3_ADD_441_U139 , P3_ADD_441_U140 , P3_ADD_441_U141 , P3_ADD_441_U142 , P3_ADD_441_U143;
wire P3_ADD_441_U144 , P3_ADD_441_U145 , P3_ADD_441_U146 , P3_ADD_441_U147 , P3_ADD_441_U148 , P3_ADD_441_U149 , P3_ADD_441_U150 , P3_ADD_441_U151 , P3_ADD_441_U152 , P3_ADD_441_U153;
wire P3_ADD_441_U154 , P3_ADD_441_U155 , P3_ADD_441_U156 , P3_ADD_441_U157 , P3_ADD_441_U158 , P3_ADD_441_U159 , P3_ADD_441_U160 , P3_ADD_441_U161 , P3_ADD_441_U162 , P3_ADD_441_U163;
wire P3_ADD_441_U164 , P3_ADD_441_U165 , P3_ADD_441_U166 , P3_ADD_441_U167 , P3_ADD_441_U168 , P3_ADD_441_U169 , P3_ADD_441_U170 , P3_ADD_441_U171 , P3_ADD_441_U172 , P3_ADD_441_U173;
wire P3_ADD_441_U174 , P3_ADD_441_U175 , P3_ADD_441_U176 , P3_ADD_441_U177 , P3_ADD_441_U178 , P3_ADD_441_U179 , P3_ADD_441_U180 , P3_ADD_441_U181 , P3_ADD_441_U182 , P3_ADD_349_U5;
wire P3_ADD_349_U6 , P3_ADD_349_U7 , P3_ADD_349_U8 , P3_ADD_349_U9 , P3_ADD_349_U10 , P3_ADD_349_U11 , P3_ADD_349_U12 , P3_ADD_349_U13 , P3_ADD_349_U14 , P3_ADD_349_U15;
wire P3_ADD_349_U16 , P3_ADD_349_U17 , P3_ADD_349_U18 , P3_ADD_349_U19 , P3_ADD_349_U20 , P3_ADD_349_U21 , P3_ADD_349_U22 , P3_ADD_349_U23 , P3_ADD_349_U24 , P3_ADD_349_U25;
wire P3_ADD_349_U26 , P3_ADD_349_U27 , P3_ADD_349_U28 , P3_ADD_349_U29 , P3_ADD_349_U30 , P3_ADD_349_U31 , P3_ADD_349_U32 , P3_ADD_349_U33 , P3_ADD_349_U34 , P3_ADD_349_U35;
wire P3_ADD_349_U36 , P3_ADD_349_U37 , P3_ADD_349_U38 , P3_ADD_349_U39 , P3_ADD_349_U40 , P3_ADD_349_U41 , P3_ADD_349_U42 , P3_ADD_349_U43 , P3_ADD_349_U44 , P3_ADD_349_U45;
wire P3_ADD_349_U46 , P3_ADD_349_U47 , P3_ADD_349_U48 , P3_ADD_349_U49 , P3_ADD_349_U50 , P3_ADD_349_U51 , P3_ADD_349_U52 , P3_ADD_349_U53 , P3_ADD_349_U54 , P3_ADD_349_U55;
wire P3_ADD_349_U56 , P3_ADD_349_U57 , P3_ADD_349_U58 , P3_ADD_349_U59 , P3_ADD_349_U60 , P3_ADD_349_U61 , P3_ADD_349_U62 , P3_ADD_349_U63 , P3_ADD_349_U64 , P3_ADD_349_U65;
wire P3_ADD_349_U66 , P3_ADD_349_U67 , P3_ADD_349_U68 , P3_ADD_349_U69 , P3_ADD_349_U70 , P3_ADD_349_U71 , P3_ADD_349_U72 , P3_ADD_349_U73 , P3_ADD_349_U74 , P3_ADD_349_U75;
wire P3_ADD_349_U76 , P3_ADD_349_U77 , P3_ADD_349_U78 , P3_ADD_349_U79 , P3_ADD_349_U80 , P3_ADD_349_U81 , P3_ADD_349_U82 , P3_ADD_349_U83 , P3_ADD_349_U84 , P3_ADD_349_U85;
wire P3_ADD_349_U86 , P3_ADD_349_U87 , P3_ADD_349_U88 , P3_ADD_349_U89 , P3_ADD_349_U90 , P3_ADD_349_U91 , P3_ADD_349_U92 , P3_ADD_349_U93 , P3_ADD_349_U94 , P3_ADD_349_U95;
wire P3_ADD_349_U96 , P3_ADD_349_U97 , P3_ADD_349_U98 , P3_ADD_349_U99 , P3_ADD_349_U100 , P3_ADD_349_U101 , P3_ADD_349_U102 , P3_ADD_349_U103 , P3_ADD_349_U104 , P3_ADD_349_U105;
wire P3_ADD_349_U106 , P3_ADD_349_U107 , P3_ADD_349_U108 , P3_ADD_349_U109 , P3_ADD_349_U110 , P3_ADD_349_U111 , P3_ADD_349_U112 , P3_ADD_349_U113 , P3_ADD_349_U114 , P3_ADD_349_U115;
wire P3_ADD_349_U116 , P3_ADD_349_U117 , P3_ADD_349_U118 , P3_ADD_349_U119 , P3_ADD_349_U120 , P3_ADD_349_U121 , P3_ADD_349_U122 , P3_ADD_349_U123 , P3_ADD_349_U124 , P3_ADD_349_U125;
wire P3_ADD_349_U126 , P3_ADD_349_U127 , P3_ADD_349_U128 , P3_ADD_349_U129 , P3_ADD_349_U130 , P3_ADD_349_U131 , P3_ADD_349_U132 , P3_ADD_349_U133 , P3_ADD_349_U134 , P3_ADD_349_U135;
wire P3_ADD_349_U136 , P3_ADD_349_U137 , P3_ADD_349_U138 , P3_ADD_349_U139 , P3_ADD_349_U140 , P3_ADD_349_U141 , P3_ADD_349_U142 , P3_ADD_349_U143 , P3_ADD_349_U144 , P3_ADD_349_U145;
wire P3_ADD_349_U146 , P3_ADD_349_U147 , P3_ADD_349_U148 , P3_ADD_349_U149 , P3_ADD_349_U150 , P3_ADD_349_U151 , P3_ADD_349_U152 , P3_ADD_349_U153 , P3_ADD_349_U154 , P3_ADD_349_U155;
wire P3_ADD_349_U156 , P3_ADD_349_U157 , P3_ADD_349_U158 , P3_ADD_349_U159 , P3_ADD_349_U160 , P3_ADD_349_U161 , P3_ADD_349_U162 , P3_ADD_349_U163 , P3_ADD_349_U164 , P3_ADD_349_U165;
wire P3_ADD_349_U166 , P3_ADD_349_U167 , P3_ADD_349_U168 , P3_ADD_349_U169 , P3_ADD_349_U170 , P3_ADD_349_U171 , P3_ADD_349_U172 , P3_ADD_349_U173 , P3_ADD_349_U174 , P3_ADD_349_U175;
wire P3_ADD_349_U176 , P3_ADD_349_U177 , P3_ADD_349_U178 , P3_ADD_349_U179 , P3_ADD_349_U180 , P3_ADD_349_U181 , P3_ADD_349_U182 , P3_ADD_349_U183 , P3_ADD_349_U184 , P3_ADD_349_U185;
wire P3_ADD_349_U186 , P3_ADD_349_U187 , P3_ADD_349_U188 , P3_ADD_349_U189 , P3_ADD_405_U4 , P3_ADD_405_U5 , P3_ADD_405_U6 , P3_ADD_405_U7 , P3_ADD_405_U8 , P3_ADD_405_U9;
wire P3_ADD_405_U10 , P3_ADD_405_U11 , P3_ADD_405_U12 , P3_ADD_405_U13 , P3_ADD_405_U14 , P3_ADD_405_U15 , P3_ADD_405_U16 , P3_ADD_405_U17 , P3_ADD_405_U18 , P3_ADD_405_U19;
wire P3_ADD_405_U20 , P3_ADD_405_U21 , P3_ADD_405_U22 , P3_ADD_405_U23 , P3_ADD_405_U24 , P3_ADD_405_U25 , P3_ADD_405_U26 , P3_ADD_405_U27 , P3_ADD_405_U28 , P3_ADD_405_U29;
wire P3_ADD_405_U30 , P3_ADD_405_U31 , P3_ADD_405_U32 , P3_ADD_405_U33 , P3_ADD_405_U34 , P3_ADD_405_U35 , P3_ADD_405_U36 , P3_ADD_405_U37 , P3_ADD_405_U38 , P3_ADD_405_U39;
wire P3_ADD_405_U40 , P3_ADD_405_U41 , P3_ADD_405_U42 , P3_ADD_405_U43 , P3_ADD_405_U44 , P3_ADD_405_U45 , P3_ADD_405_U46 , P3_ADD_405_U47 , P3_ADD_405_U48 , P3_ADD_405_U49;
wire P3_ADD_405_U50 , P3_ADD_405_U51 , P3_ADD_405_U52 , P3_ADD_405_U53 , P3_ADD_405_U54 , P3_ADD_405_U55 , P3_ADD_405_U56 , P3_ADD_405_U57 , P3_ADD_405_U58 , P3_ADD_405_U59;
wire P3_ADD_405_U60 , P3_ADD_405_U61 , P3_ADD_405_U62 , P3_ADD_405_U63 , P3_ADD_405_U64 , P3_ADD_405_U65 , P3_ADD_405_U66 , P3_ADD_405_U67 , P3_ADD_405_U68 , P3_ADD_405_U69;
wire P3_ADD_405_U70 , P3_ADD_405_U71 , P3_ADD_405_U72 , P3_ADD_405_U73 , P3_ADD_405_U74 , P3_ADD_405_U75 , P3_ADD_405_U76 , P3_ADD_405_U77 , P3_ADD_405_U78 , P3_ADD_405_U79;
wire P3_ADD_405_U80 , P3_ADD_405_U81 , P3_ADD_405_U82 , P3_ADD_405_U83 , P3_ADD_405_U84 , P3_ADD_405_U85 , P3_ADD_405_U86 , P3_ADD_405_U87 , P3_ADD_405_U88 , P3_ADD_405_U89;
wire P3_ADD_405_U90 , P3_ADD_405_U91 , P3_ADD_405_U92 , P3_ADD_405_U93 , P3_ADD_405_U94 , P3_ADD_405_U95 , P3_ADD_405_U96 , P3_ADD_405_U97 , P3_ADD_405_U98 , P3_ADD_405_U99;
wire P3_ADD_405_U100 , P3_ADD_405_U101 , P3_ADD_405_U102 , P3_ADD_405_U103 , P3_ADD_405_U104 , P3_ADD_405_U105 , P3_ADD_405_U106 , P3_ADD_405_U107 , P3_ADD_405_U108 , P3_ADD_405_U109;
wire P3_ADD_405_U110 , P3_ADD_405_U111 , P3_ADD_405_U112 , P3_ADD_405_U113 , P3_ADD_405_U114 , P3_ADD_405_U115 , P3_ADD_405_U116 , P3_ADD_405_U117 , P3_ADD_405_U118 , P3_ADD_405_U119;
wire P3_ADD_405_U120 , P3_ADD_405_U121 , P3_ADD_405_U122 , P3_ADD_405_U123 , P3_ADD_405_U124 , P3_ADD_405_U125 , P3_ADD_405_U126 , P3_ADD_405_U127 , P3_ADD_405_U128 , P3_ADD_405_U129;
wire P3_ADD_405_U130 , P3_ADD_405_U131 , P3_ADD_405_U132 , P3_ADD_405_U133 , P3_ADD_405_U134 , P3_ADD_405_U135 , P3_ADD_405_U136 , P3_ADD_405_U137 , P3_ADD_405_U138 , P3_ADD_405_U139;
wire P3_ADD_405_U140 , P3_ADD_405_U141 , P3_ADD_405_U142 , P3_ADD_405_U143 , P3_ADD_405_U144 , P3_ADD_405_U145 , P3_ADD_405_U146 , P3_ADD_405_U147 , P3_ADD_405_U148 , P3_ADD_405_U149;
wire P3_ADD_405_U150 , P3_ADD_405_U151 , P3_ADD_405_U152 , P3_ADD_405_U153 , P3_ADD_405_U154 , P3_ADD_405_U155 , P3_ADD_405_U156 , P3_ADD_405_U157 , P3_ADD_405_U158 , P3_ADD_405_U159;
wire P3_ADD_405_U160 , P3_ADD_405_U161 , P3_ADD_405_U162 , P3_ADD_405_U163 , P3_ADD_405_U164 , P3_ADD_405_U165 , P3_ADD_405_U166 , P3_ADD_405_U167 , P3_ADD_405_U168 , P3_ADD_405_U169;
wire P3_ADD_405_U170 , P3_ADD_405_U171 , P3_ADD_405_U172 , P3_ADD_405_U173 , P3_ADD_405_U174 , P3_ADD_405_U175 , P3_ADD_405_U176 , P3_ADD_405_U177 , P3_ADD_405_U178 , P3_ADD_405_U179;
wire P3_ADD_405_U180 , P3_ADD_405_U181 , P3_ADD_405_U182 , P3_ADD_405_U183 , P3_ADD_405_U184 , P3_ADD_405_U185 , P3_ADD_405_U186 , P3_ADD_553_U5 , P3_ADD_553_U6 , P3_ADD_553_U7;
wire P3_ADD_553_U8 , P3_ADD_553_U9 , P3_ADD_553_U10 , P3_ADD_553_U11 , P3_ADD_553_U12 , P3_ADD_553_U13 , P3_ADD_553_U14 , P3_ADD_553_U15 , P3_ADD_553_U16 , P3_ADD_553_U17;
wire P3_ADD_553_U18 , P3_ADD_553_U19 , P3_ADD_553_U20 , P3_ADD_553_U21 , P3_ADD_553_U22 , P3_ADD_553_U23 , P3_ADD_553_U24 , P3_ADD_553_U25 , P3_ADD_553_U26 , P3_ADD_553_U27;
wire P3_ADD_553_U28 , P3_ADD_553_U29 , P3_ADD_553_U30 , P3_ADD_553_U31 , P3_ADD_553_U32 , P3_ADD_553_U33 , P3_ADD_553_U34 , P3_ADD_553_U35 , P3_ADD_553_U36 , P3_ADD_553_U37;
wire P3_ADD_553_U38 , P3_ADD_553_U39 , P3_ADD_553_U40 , P3_ADD_553_U41 , P3_ADD_553_U42 , P3_ADD_553_U43 , P3_ADD_553_U44 , P3_ADD_553_U45 , P3_ADD_553_U46 , P3_ADD_553_U47;
wire P3_ADD_553_U48 , P3_ADD_553_U49 , P3_ADD_553_U50 , P3_ADD_553_U51 , P3_ADD_553_U52 , P3_ADD_553_U53 , P3_ADD_553_U54 , P3_ADD_553_U55 , P3_ADD_553_U56 , P3_ADD_553_U57;
wire P3_ADD_553_U58 , P3_ADD_553_U59 , P3_ADD_553_U60 , P3_ADD_553_U61 , P3_ADD_553_U62 , P3_ADD_553_U63 , P3_ADD_553_U64 , P3_ADD_553_U65 , P3_ADD_553_U66 , P3_ADD_553_U67;
wire P3_ADD_553_U68 , P3_ADD_553_U69 , P3_ADD_553_U70 , P3_ADD_553_U71 , P3_ADD_553_U72 , P3_ADD_553_U73 , P3_ADD_553_U74 , P3_ADD_553_U75 , P3_ADD_553_U76 , P3_ADD_553_U77;
wire P3_ADD_553_U78 , P3_ADD_553_U79 , P3_ADD_553_U80 , P3_ADD_553_U81 , P3_ADD_553_U82 , P3_ADD_553_U83 , P3_ADD_553_U84 , P3_ADD_553_U85 , P3_ADD_553_U86 , P3_ADD_553_U87;
wire P3_ADD_553_U88 , P3_ADD_553_U89 , P3_ADD_553_U90 , P3_ADD_553_U91 , P3_ADD_553_U92 , P3_ADD_553_U93 , P3_ADD_553_U94 , P3_ADD_553_U95 , P3_ADD_553_U96 , P3_ADD_553_U97;
wire P3_ADD_553_U98 , P3_ADD_553_U99 , P3_ADD_553_U100 , P3_ADD_553_U101 , P3_ADD_553_U102 , P3_ADD_553_U103 , P3_ADD_553_U104 , P3_ADD_553_U105 , P3_ADD_553_U106 , P3_ADD_553_U107;
wire P3_ADD_553_U108 , P3_ADD_553_U109 , P3_ADD_553_U110 , P3_ADD_553_U111 , P3_ADD_553_U112 , P3_ADD_553_U113 , P3_ADD_553_U114 , P3_ADD_553_U115 , P3_ADD_553_U116 , P3_ADD_553_U117;
wire P3_ADD_553_U118 , P3_ADD_553_U119 , P3_ADD_553_U120 , P3_ADD_553_U121 , P3_ADD_553_U122 , P3_ADD_553_U123 , P3_ADD_553_U124 , P3_ADD_553_U125 , P3_ADD_553_U126 , P3_ADD_553_U127;
wire P3_ADD_553_U128 , P3_ADD_553_U129 , P3_ADD_553_U130 , P3_ADD_553_U131 , P3_ADD_553_U132 , P3_ADD_553_U133 , P3_ADD_553_U134 , P3_ADD_553_U135 , P3_ADD_553_U136 , P3_ADD_553_U137;
wire P3_ADD_553_U138 , P3_ADD_553_U139 , P3_ADD_553_U140 , P3_ADD_553_U141 , P3_ADD_553_U142 , P3_ADD_553_U143 , P3_ADD_553_U144 , P3_ADD_553_U145 , P3_ADD_553_U146 , P3_ADD_553_U147;
wire P3_ADD_553_U148 , P3_ADD_553_U149 , P3_ADD_553_U150 , P3_ADD_553_U151 , P3_ADD_553_U152 , P3_ADD_553_U153 , P3_ADD_553_U154 , P3_ADD_553_U155 , P3_ADD_553_U156 , P3_ADD_553_U157;
wire P3_ADD_553_U158 , P3_ADD_553_U159 , P3_ADD_553_U160 , P3_ADD_553_U161 , P3_ADD_553_U162 , P3_ADD_553_U163 , P3_ADD_553_U164 , P3_ADD_553_U165 , P3_ADD_553_U166 , P3_ADD_553_U167;
wire P3_ADD_553_U168 , P3_ADD_553_U169 , P3_ADD_553_U170 , P3_ADD_553_U171 , P3_ADD_553_U172 , P3_ADD_553_U173 , P3_ADD_553_U174 , P3_ADD_553_U175 , P3_ADD_553_U176 , P3_ADD_553_U177;
wire P3_ADD_553_U178 , P3_ADD_553_U179 , P3_ADD_553_U180 , P3_ADD_553_U181 , P3_ADD_553_U182 , P3_ADD_553_U183 , P3_ADD_553_U184 , P3_ADD_553_U185 , P3_ADD_553_U186 , P3_ADD_553_U187;
wire P3_ADD_553_U188 , P3_ADD_553_U189 , P3_ADD_558_U5 , P3_ADD_558_U6 , P3_ADD_558_U7 , P3_ADD_558_U8 , P3_ADD_558_U9 , P3_ADD_558_U10 , P3_ADD_558_U11 , P3_ADD_558_U12;
wire P3_ADD_558_U13 , P3_ADD_558_U14 , P3_ADD_558_U15 , P3_ADD_558_U16 , P3_ADD_558_U17 , P3_ADD_558_U18 , P3_ADD_558_U19 , P3_ADD_558_U20 , P3_ADD_558_U21 , P3_ADD_558_U22;
wire P3_ADD_558_U23 , P3_ADD_558_U24 , P3_ADD_558_U25 , P3_ADD_558_U26 , P3_ADD_558_U27 , P3_ADD_558_U28 , P3_ADD_558_U29 , P3_ADD_558_U30 , P3_ADD_558_U31 , P3_ADD_558_U32;
wire P3_ADD_558_U33 , P3_ADD_558_U34 , P3_ADD_558_U35 , P3_ADD_558_U36 , P3_ADD_558_U37 , P3_ADD_558_U38 , P3_ADD_558_U39 , P3_ADD_558_U40 , P3_ADD_558_U41 , P3_ADD_558_U42;
wire P3_ADD_558_U43 , P3_ADD_558_U44 , P3_ADD_558_U45 , P3_ADD_558_U46 , P3_ADD_558_U47 , P3_ADD_558_U48 , P3_ADD_558_U49 , P3_ADD_558_U50 , P3_ADD_558_U51 , P3_ADD_558_U52;
wire P3_ADD_558_U53 , P3_ADD_558_U54 , P3_ADD_558_U55 , P3_ADD_558_U56 , P3_ADD_558_U57 , P3_ADD_558_U58 , P3_ADD_558_U59 , P3_ADD_558_U60 , P3_ADD_558_U61 , P3_ADD_558_U62;
wire P3_ADD_558_U63 , P3_ADD_558_U64 , P3_ADD_558_U65 , P3_ADD_558_U66 , P3_ADD_558_U67 , P3_ADD_558_U68 , P3_ADD_558_U69 , P3_ADD_558_U70 , P3_ADD_558_U71 , P3_ADD_558_U72;
wire P3_ADD_558_U73 , P3_ADD_558_U74 , P3_ADD_558_U75 , P3_ADD_558_U76 , P3_ADD_558_U77 , P3_ADD_558_U78 , P3_ADD_558_U79 , P3_ADD_558_U80 , P3_ADD_558_U81 , P3_ADD_558_U82;
wire P3_ADD_558_U83 , P3_ADD_558_U84 , P3_ADD_558_U85 , P3_ADD_558_U86 , P3_ADD_558_U87 , P3_ADD_558_U88 , P3_ADD_558_U89 , P3_ADD_558_U90 , P3_ADD_558_U91 , P3_ADD_558_U92;
wire P3_ADD_558_U93 , P3_ADD_558_U94 , P3_ADD_558_U95 , P3_ADD_558_U96 , P3_ADD_558_U97 , P3_ADD_558_U98 , P3_ADD_558_U99 , P3_ADD_558_U100 , P3_ADD_558_U101 , P3_ADD_558_U102;
wire P3_ADD_558_U103 , P3_ADD_558_U104 , P3_ADD_558_U105 , P3_ADD_558_U106 , P3_ADD_558_U107 , P3_ADD_558_U108 , P3_ADD_558_U109 , P3_ADD_558_U110 , P3_ADD_558_U111 , P3_ADD_558_U112;
wire P3_ADD_558_U113 , P3_ADD_558_U114 , P3_ADD_558_U115 , P3_ADD_558_U116 , P3_ADD_558_U117 , P3_ADD_558_U118 , P3_ADD_558_U119 , P3_ADD_558_U120 , P3_ADD_558_U121 , P3_ADD_558_U122;
wire P3_ADD_558_U123 , P3_ADD_558_U124 , P3_ADD_558_U125 , P3_ADD_558_U126 , P3_ADD_558_U127 , P3_ADD_558_U128 , P3_ADD_558_U129 , P3_ADD_558_U130 , P3_ADD_558_U131 , P3_ADD_558_U132;
wire P3_ADD_558_U133 , P3_ADD_558_U134 , P3_ADD_558_U135 , P3_ADD_558_U136 , P3_ADD_558_U137 , P3_ADD_558_U138 , P3_ADD_558_U139 , P3_ADD_558_U140 , P3_ADD_558_U141 , P3_ADD_558_U142;
wire P3_ADD_558_U143 , P3_ADD_558_U144 , P3_ADD_558_U145 , P3_ADD_558_U146 , P3_ADD_558_U147 , P3_ADD_558_U148 , P3_ADD_558_U149 , P3_ADD_558_U150 , P3_ADD_558_U151 , P3_ADD_558_U152;
wire P3_ADD_558_U153 , P3_ADD_558_U154 , P3_ADD_558_U155 , P3_ADD_558_U156 , P3_ADD_558_U157 , P3_ADD_558_U158 , P3_ADD_558_U159 , P3_ADD_558_U160 , P3_ADD_558_U161 , P3_ADD_558_U162;
wire P3_ADD_558_U163 , P3_ADD_558_U164 , P3_ADD_558_U165 , P3_ADD_558_U166 , P3_ADD_558_U167 , P3_ADD_558_U168 , P3_ADD_558_U169 , P3_ADD_558_U170 , P3_ADD_558_U171 , P3_ADD_558_U172;
wire P3_ADD_558_U173 , P3_ADD_558_U174 , P3_ADD_558_U175 , P3_ADD_558_U176 , P3_ADD_558_U177 , P3_ADD_558_U178 , P3_ADD_558_U179 , P3_ADD_558_U180 , P3_ADD_558_U181 , P3_ADD_558_U182;
wire P3_ADD_558_U183 , P3_ADD_558_U184 , P3_ADD_558_U185 , P3_ADD_558_U186 , P3_ADD_558_U187 , P3_ADD_558_U188 , P3_ADD_558_U189 , P3_ADD_385_U5 , P3_ADD_385_U6 , P3_ADD_385_U7;
wire P3_ADD_385_U8 , P3_ADD_385_U9 , P3_ADD_385_U10 , P3_ADD_385_U11 , P3_ADD_385_U12 , P3_ADD_385_U13 , P3_ADD_385_U14 , P3_ADD_385_U15 , P3_ADD_385_U16 , P3_ADD_385_U17;
wire P3_ADD_385_U18 , P3_ADD_385_U19 , P3_ADD_385_U20 , P3_ADD_385_U21 , P3_ADD_385_U22 , P3_ADD_385_U23 , P3_ADD_385_U24 , P3_ADD_385_U25 , P3_ADD_385_U26 , P3_ADD_385_U27;
wire P3_ADD_385_U28 , P3_ADD_385_U29 , P3_ADD_385_U30 , P3_ADD_385_U31 , P3_ADD_385_U32 , P3_ADD_385_U33 , P3_ADD_385_U34 , P3_ADD_385_U35 , P3_ADD_385_U36 , P3_ADD_385_U37;
wire P3_ADD_385_U38 , P3_ADD_385_U39 , P3_ADD_385_U40 , P3_ADD_385_U41 , P3_ADD_385_U42 , P3_ADD_385_U43 , P3_ADD_385_U44 , P3_ADD_385_U45 , P3_ADD_385_U46 , P3_ADD_385_U47;
wire P3_ADD_385_U48 , P3_ADD_385_U49 , P3_ADD_385_U50 , P3_ADD_385_U51 , P3_ADD_385_U52 , P3_ADD_385_U53 , P3_ADD_385_U54 , P3_ADD_385_U55 , P3_ADD_385_U56 , P3_ADD_385_U57;
wire P3_ADD_385_U58 , P3_ADD_385_U59 , P3_ADD_385_U60 , P3_ADD_385_U61 , P3_ADD_385_U62 , P3_ADD_385_U63 , P3_ADD_385_U64 , P3_ADD_385_U65 , P3_ADD_385_U66 , P3_ADD_385_U67;
wire P3_ADD_385_U68 , P3_ADD_385_U69 , P3_ADD_385_U70 , P3_ADD_385_U71 , P3_ADD_385_U72 , P3_ADD_385_U73 , P3_ADD_385_U74 , P3_ADD_385_U75 , P3_ADD_385_U76 , P3_ADD_385_U77;
wire P3_ADD_385_U78 , P3_ADD_385_U79 , P3_ADD_385_U80 , P3_ADD_385_U81 , P3_ADD_385_U82 , P3_ADD_385_U83 , P3_ADD_385_U84 , P3_ADD_385_U85 , P3_ADD_385_U86 , P3_ADD_385_U87;
wire P3_ADD_385_U88 , P3_ADD_385_U89 , P3_ADD_385_U90 , P3_ADD_385_U91 , P3_ADD_385_U92 , P3_ADD_385_U93 , P3_ADD_385_U94 , P3_ADD_385_U95 , P3_ADD_385_U96 , P3_ADD_385_U97;
wire P3_ADD_385_U98 , P3_ADD_385_U99 , P3_ADD_385_U100 , P3_ADD_385_U101 , P3_ADD_385_U102 , P3_ADD_385_U103 , P3_ADD_385_U104 , P3_ADD_385_U105 , P3_ADD_385_U106 , P3_ADD_385_U107;
wire P3_ADD_385_U108 , P3_ADD_385_U109 , P3_ADD_385_U110 , P3_ADD_385_U111 , P3_ADD_385_U112 , P3_ADD_385_U113 , P3_ADD_385_U114 , P3_ADD_385_U115 , P3_ADD_385_U116 , P3_ADD_385_U117;
wire P3_ADD_385_U118 , P3_ADD_385_U119 , P3_ADD_385_U120 , P3_ADD_385_U121 , P3_ADD_385_U122 , P3_ADD_385_U123 , P3_ADD_385_U124 , P3_ADD_385_U125 , P3_ADD_385_U126 , P3_ADD_385_U127;
wire P3_ADD_385_U128 , P3_ADD_385_U129 , P3_ADD_385_U130 , P3_ADD_385_U131 , P3_ADD_385_U132 , P3_ADD_385_U133 , P3_ADD_385_U134 , P3_ADD_385_U135 , P3_ADD_385_U136 , P3_ADD_385_U137;
wire P3_ADD_385_U138 , P3_ADD_385_U139 , P3_ADD_385_U140 , P3_ADD_385_U141 , P3_ADD_385_U142 , P3_ADD_385_U143 , P3_ADD_385_U144 , P3_ADD_385_U145 , P3_ADD_385_U146 , P3_ADD_385_U147;
wire P3_ADD_385_U148 , P3_ADD_385_U149 , P3_ADD_385_U150 , P3_ADD_385_U151 , P3_ADD_385_U152 , P3_ADD_385_U153 , P3_ADD_385_U154 , P3_ADD_385_U155 , P3_ADD_385_U156 , P3_ADD_385_U157;
wire P3_ADD_385_U158 , P3_ADD_385_U159 , P3_ADD_385_U160 , P3_ADD_385_U161 , P3_ADD_385_U162 , P3_ADD_385_U163 , P3_ADD_385_U164 , P3_ADD_385_U165 , P3_ADD_385_U166 , P3_ADD_385_U167;
wire P3_ADD_385_U168 , P3_ADD_385_U169 , P3_ADD_385_U170 , P3_ADD_385_U171 , P3_ADD_385_U172 , P3_ADD_385_U173 , P3_ADD_385_U174 , P3_ADD_385_U175 , P3_ADD_385_U176 , P3_ADD_385_U177;
wire P3_ADD_385_U178 , P3_ADD_385_U179 , P3_ADD_385_U180 , P3_ADD_385_U181 , P3_ADD_385_U182 , P3_ADD_385_U183 , P3_ADD_385_U184 , P3_ADD_385_U185 , P3_ADD_385_U186 , P3_ADD_385_U187;
wire P3_ADD_385_U188 , P3_ADD_385_U189 , P3_ADD_357_U6 , P3_ADD_357_U7 , P3_ADD_357_U8 , P3_ADD_357_U9 , P3_ADD_357_U10 , P3_ADD_357_U11 , P3_ADD_357_U12 , P3_ADD_357_U13;
wire P3_ADD_357_U14 , P3_ADD_357_U15 , P3_ADD_357_U16 , P3_ADD_357_U17 , P3_ADD_357_U18 , P3_ADD_357_U19 , P3_ADD_357_U20 , P3_ADD_357_U21 , P3_ADD_357_U22 , P3_ADD_357_U23;
wire P3_ADD_357_U24 , P3_ADD_357_U25 , P3_ADD_357_U26 , P3_ADD_357_U27 , P3_ADD_357_U28 , P3_ADD_357_U29 , P3_ADD_357_U30 , P3_ADD_357_U31 , P3_ADD_357_U32 , P3_ADD_357_U33;
wire P3_ADD_357_U34 , P3_ADD_357_U35 , P3_ADD_547_U5 , P3_ADD_547_U6 , P3_ADD_547_U7 , P3_ADD_547_U8 , P3_ADD_547_U9 , P3_ADD_547_U10 , P3_ADD_547_U11 , P3_ADD_547_U12;
wire P3_ADD_547_U13 , P3_ADD_547_U14 , P3_ADD_547_U15 , P3_ADD_547_U16 , P3_ADD_547_U17 , P3_ADD_547_U18 , P3_ADD_547_U19 , P3_ADD_547_U20 , P3_ADD_547_U21 , P3_ADD_547_U22;
wire P3_ADD_547_U23 , P3_ADD_547_U24 , P3_ADD_547_U25 , P3_ADD_547_U26 , P3_ADD_547_U27 , P3_ADD_547_U28 , P3_ADD_547_U29 , P3_ADD_547_U30 , P3_ADD_547_U31 , P3_ADD_547_U32;
wire P3_ADD_547_U33 , P3_ADD_547_U34 , P3_ADD_547_U35 , P3_ADD_547_U36 , P3_ADD_547_U37 , P3_ADD_547_U38 , P3_ADD_547_U39 , P3_ADD_547_U40 , P3_ADD_547_U41 , P3_ADD_547_U42;
wire P3_ADD_547_U43 , P3_ADD_547_U44 , P3_ADD_547_U45 , P3_ADD_547_U46 , P3_ADD_547_U47 , P3_ADD_547_U48 , P3_ADD_547_U49 , P3_ADD_547_U50 , P3_ADD_547_U51 , P3_ADD_547_U52;
wire P3_ADD_547_U53 , P3_ADD_547_U54 , P3_ADD_547_U55 , P3_ADD_547_U56 , P3_ADD_547_U57 , P3_ADD_547_U58 , P3_ADD_547_U59 , P3_ADD_547_U60 , P3_ADD_547_U61 , P3_ADD_547_U62;
wire P3_ADD_547_U63 , P3_ADD_547_U64 , P3_ADD_547_U65 , P3_ADD_547_U66 , P3_ADD_547_U67 , P3_ADD_547_U68 , P3_ADD_547_U69 , P3_ADD_547_U70 , P3_ADD_547_U71 , P3_ADD_547_U72;
wire P3_ADD_547_U73 , P3_ADD_547_U74 , P3_ADD_547_U75 , P3_ADD_547_U76 , P3_ADD_547_U77 , P3_ADD_547_U78 , P3_ADD_547_U79 , P3_ADD_547_U80 , P3_ADD_547_U81 , P3_ADD_547_U82;
wire P3_ADD_547_U83 , P3_ADD_547_U84 , P3_ADD_547_U85 , P3_ADD_547_U86 , P3_ADD_547_U87 , P3_ADD_547_U88 , P3_ADD_547_U89 , P3_ADD_547_U90 , P3_ADD_547_U91 , P3_ADD_547_U92;
wire P3_ADD_547_U93 , P3_ADD_547_U94 , P3_ADD_547_U95 , P3_ADD_547_U96 , P3_ADD_547_U97 , P3_ADD_547_U98 , P3_ADD_547_U99 , P3_ADD_547_U100 , P3_ADD_547_U101 , P3_ADD_547_U102;
wire P3_ADD_547_U103 , P3_ADD_547_U104 , P3_ADD_547_U105 , P3_ADD_547_U106 , P3_ADD_547_U107 , P3_ADD_547_U108 , P3_ADD_547_U109 , P3_ADD_547_U110 , P3_ADD_547_U111 , P3_ADD_547_U112;
wire P3_ADD_547_U113 , P3_ADD_547_U114 , P3_ADD_547_U115 , P3_ADD_547_U116 , P3_ADD_547_U117 , P3_ADD_547_U118 , P3_ADD_547_U119 , P3_ADD_547_U120 , P3_ADD_547_U121 , P3_ADD_547_U122;
wire P3_ADD_547_U123 , P3_ADD_547_U124 , P3_ADD_547_U125 , P3_ADD_547_U126 , P3_ADD_547_U127 , P3_ADD_547_U128 , P3_ADD_547_U129 , P3_ADD_547_U130 , P3_ADD_547_U131 , P3_ADD_547_U132;
wire P3_ADD_547_U133 , P3_ADD_547_U134 , P3_ADD_547_U135 , P3_ADD_547_U136 , P3_ADD_547_U137 , P3_ADD_547_U138 , P3_ADD_547_U139 , P3_ADD_547_U140 , P3_ADD_547_U141 , P3_ADD_547_U142;
wire P3_ADD_547_U143 , P3_ADD_547_U144 , P3_ADD_547_U145 , P3_ADD_547_U146 , P3_ADD_547_U147 , P3_ADD_547_U148 , P3_ADD_547_U149 , P3_ADD_547_U150 , P3_ADD_547_U151 , P3_ADD_547_U152;
wire P3_ADD_547_U153 , P3_ADD_547_U154 , P3_ADD_547_U155 , P3_ADD_547_U156 , P3_ADD_547_U157 , P3_ADD_547_U158 , P3_ADD_547_U159 , P3_ADD_547_U160 , P3_ADD_547_U161 , P3_ADD_547_U162;
wire P3_ADD_547_U163 , P3_ADD_547_U164 , P3_ADD_547_U165 , P3_ADD_547_U166 , P3_ADD_547_U167 , P3_ADD_547_U168 , P3_ADD_547_U169 , P3_ADD_547_U170 , P3_ADD_547_U171 , P3_ADD_547_U172;
wire P3_ADD_547_U173 , P3_ADD_547_U174 , P3_ADD_547_U175 , P3_ADD_547_U176 , P3_ADD_547_U177 , P3_ADD_547_U178 , P3_ADD_547_U179 , P3_ADD_547_U180 , P3_ADD_547_U181 , P3_ADD_547_U182;
wire P3_ADD_547_U183 , P3_ADD_547_U184 , P3_ADD_547_U185 , P3_ADD_547_U186 , P3_ADD_547_U187 , P3_ADD_547_U188 , P3_ADD_547_U189 , P3_SUB_412_U6 , P3_SUB_412_U7 , P3_SUB_412_U8;
wire P3_SUB_412_U9 , P3_SUB_412_U10 , P3_SUB_412_U11 , P3_SUB_412_U12 , P3_SUB_412_U13 , P3_SUB_412_U14 , P3_SUB_412_U15 , P3_SUB_412_U16 , P3_SUB_412_U17 , P3_SUB_412_U18;
wire P3_SUB_412_U19 , P3_SUB_412_U20 , P3_SUB_412_U21 , P3_SUB_412_U22 , P3_SUB_412_U23 , P3_SUB_412_U24 , P3_SUB_412_U25 , P3_SUB_412_U26 , P3_SUB_412_U27 , P3_SUB_412_U28;
wire P3_SUB_412_U29 , P3_SUB_412_U30 , P3_SUB_412_U31 , P3_SUB_412_U32 , P3_SUB_412_U33 , P3_SUB_412_U34 , P3_SUB_412_U35 , P3_SUB_412_U36 , P3_SUB_412_U37 , P3_SUB_412_U38;
wire P3_SUB_412_U39 , P3_SUB_412_U40 , P3_SUB_412_U41 , P3_SUB_412_U42 , P3_SUB_412_U43 , P3_SUB_412_U44 , P3_SUB_412_U45 , P3_SUB_412_U46 , P3_SUB_412_U47 , P3_SUB_412_U48;
wire P3_SUB_412_U49 , P3_SUB_412_U50 , P3_SUB_412_U51 , P3_SUB_412_U52 , P3_SUB_412_U53 , P3_SUB_412_U54 , P3_SUB_412_U55 , P3_SUB_412_U56 , P3_SUB_412_U57 , P3_SUB_412_U58;
wire P3_SUB_412_U59 , P3_SUB_412_U60 , P3_SUB_412_U61 , P3_SUB_412_U62 , P3_SUB_412_U63 , P3_ADD_371_1212_U4 , P3_ADD_371_1212_U5 , P3_ADD_371_1212_U6 , P3_ADD_371_1212_U7 , P3_ADD_371_1212_U8;
wire P3_ADD_371_1212_U9 , P3_ADD_371_1212_U10 , P3_ADD_371_1212_U11 , P3_ADD_371_1212_U12 , P3_ADD_371_1212_U13 , P3_ADD_371_1212_U14 , P3_ADD_371_1212_U15 , P3_ADD_371_1212_U16 , P3_ADD_371_1212_U17 , P3_ADD_371_1212_U18;
wire P3_ADD_371_1212_U19 , P3_ADD_371_1212_U20 , P3_ADD_371_1212_U21 , P3_ADD_371_1212_U22 , P3_ADD_371_1212_U23 , P3_ADD_371_1212_U24 , P3_ADD_371_1212_U25 , P3_ADD_371_1212_U26 , P3_ADD_371_1212_U27 , P3_ADD_371_1212_U28;
wire P3_ADD_371_1212_U29 , P3_ADD_371_1212_U30 , P3_ADD_371_1212_U31 , P3_ADD_371_1212_U32 , P3_ADD_371_1212_U33 , P3_ADD_371_1212_U34 , P3_ADD_371_1212_U35 , P3_ADD_371_1212_U36 , P3_ADD_371_1212_U37 , P3_ADD_371_1212_U38;
wire P3_ADD_371_1212_U39 , P3_ADD_371_1212_U40 , P3_ADD_371_1212_U41 , P3_ADD_371_1212_U42 , P3_ADD_371_1212_U43 , P3_ADD_371_1212_U44 , P3_ADD_371_1212_U45 , P3_ADD_371_1212_U46 , P3_ADD_371_1212_U47 , P3_ADD_371_1212_U48;
wire P3_ADD_371_1212_U49 , P3_ADD_371_1212_U50 , P3_ADD_371_1212_U51 , P3_ADD_371_1212_U52 , P3_ADD_371_1212_U53 , P3_ADD_371_1212_U54 , P3_ADD_371_1212_U55 , P3_ADD_371_1212_U56 , P3_ADD_371_1212_U57 , P3_ADD_371_1212_U58;
wire P3_ADD_371_1212_U59 , P3_ADD_371_1212_U60 , P3_ADD_371_1212_U61 , P3_ADD_371_1212_U62 , P3_ADD_371_1212_U63 , P3_ADD_371_1212_U64 , P3_ADD_371_1212_U65 , P3_ADD_371_1212_U66 , P3_ADD_371_1212_U67 , P3_ADD_371_1212_U68;
wire P3_ADD_371_1212_U69 , P3_ADD_371_1212_U70 , P3_ADD_371_1212_U71 , P3_ADD_371_1212_U72 , P3_ADD_371_1212_U73 , P3_ADD_371_1212_U74 , P3_ADD_371_1212_U75 , P3_ADD_371_1212_U76 , P3_ADD_371_1212_U77 , P3_ADD_371_1212_U78;
wire P3_ADD_371_1212_U79 , P3_ADD_371_1212_U80 , P3_ADD_371_1212_U81 , P3_ADD_371_1212_U82 , P3_ADD_371_1212_U83 , P3_ADD_371_1212_U84 , P3_ADD_371_1212_U85 , P3_ADD_371_1212_U86 , P3_ADD_371_1212_U87 , P3_ADD_371_1212_U88;
wire P3_ADD_371_1212_U89 , P3_ADD_371_1212_U90 , P3_ADD_371_1212_U91 , P3_ADD_371_1212_U92 , P3_ADD_371_1212_U93 , P3_ADD_371_1212_U94 , P3_ADD_371_1212_U95 , P3_ADD_371_1212_U96 , P3_ADD_371_1212_U97 , P3_ADD_371_1212_U98;
wire P3_ADD_371_1212_U99 , P3_ADD_371_1212_U100 , P3_ADD_371_1212_U101 , P3_ADD_371_1212_U102 , P3_ADD_371_1212_U103 , P3_ADD_371_1212_U104 , P3_ADD_371_1212_U105 , P3_ADD_371_1212_U106 , P3_ADD_371_1212_U107 , P3_ADD_371_1212_U108;
wire P3_ADD_371_1212_U109 , P3_ADD_371_1212_U110 , P3_ADD_371_1212_U111 , P3_ADD_371_1212_U112 , P3_ADD_371_1212_U113 , P3_ADD_371_1212_U114 , P3_ADD_371_1212_U115 , P3_ADD_371_1212_U116 , P3_ADD_371_1212_U117 , P3_ADD_371_1212_U118;
wire P3_ADD_371_1212_U119 , P3_ADD_371_1212_U120 , P3_ADD_371_1212_U121 , P3_ADD_371_1212_U122 , P3_ADD_371_1212_U123 , P3_ADD_371_1212_U124 , P3_ADD_371_1212_U125 , P3_ADD_371_1212_U126 , P3_ADD_371_1212_U127 , P3_ADD_371_1212_U128;
wire P3_ADD_371_1212_U129 , P3_ADD_371_1212_U130 , P3_ADD_371_1212_U131 , P3_ADD_371_1212_U132 , P3_ADD_371_1212_U133 , P3_ADD_371_1212_U134 , P3_ADD_371_1212_U135 , P3_ADD_371_1212_U136 , P3_ADD_371_1212_U137 , P3_ADD_371_1212_U138;
wire P3_ADD_371_1212_U139 , P3_ADD_371_1212_U140 , P3_ADD_371_1212_U141 , P3_ADD_371_1212_U142 , P3_ADD_371_1212_U143 , P3_ADD_371_1212_U144 , P3_ADD_371_1212_U145 , P3_ADD_371_1212_U146 , P3_ADD_371_1212_U147 , P3_ADD_371_1212_U148;
wire P3_ADD_371_1212_U149 , P3_ADD_371_1212_U150 , P3_ADD_371_1212_U151 , P3_ADD_371_1212_U152 , P3_ADD_371_1212_U153 , P3_ADD_371_1212_U154 , P3_ADD_371_1212_U155 , P3_ADD_371_1212_U156 , P3_ADD_371_1212_U157 , P3_ADD_371_1212_U158;
wire P3_ADD_371_1212_U159 , P3_ADD_371_1212_U160 , P3_ADD_371_1212_U161 , P3_ADD_371_1212_U162 , P3_ADD_371_1212_U163 , P3_ADD_371_1212_U164 , P3_ADD_371_1212_U165 , P3_ADD_371_1212_U166 , P3_ADD_371_1212_U167 , P3_ADD_371_1212_U168;
wire P3_ADD_371_1212_U169 , P3_ADD_371_1212_U170 , P3_ADD_371_1212_U171 , P3_ADD_371_1212_U172 , P3_ADD_371_1212_U173 , P3_ADD_371_1212_U174 , P3_ADD_371_1212_U175 , P3_ADD_371_1212_U176 , P3_ADD_371_1212_U177 , P3_ADD_371_1212_U178;
wire P3_ADD_371_1212_U179 , P3_ADD_371_1212_U180 , P3_ADD_371_1212_U181 , P3_ADD_371_1212_U182 , P3_ADD_371_1212_U183 , P3_ADD_371_1212_U184 , P3_ADD_371_1212_U185 , P3_ADD_371_1212_U186 , P3_ADD_371_1212_U187 , P3_ADD_371_1212_U188;
wire P3_ADD_371_1212_U189 , P3_ADD_371_1212_U190 , P3_ADD_371_1212_U191 , P3_ADD_371_1212_U192 , P3_ADD_371_1212_U193 , P3_ADD_371_1212_U194 , P3_ADD_371_1212_U195 , P3_ADD_371_1212_U196 , P3_ADD_371_1212_U197 , P3_ADD_371_1212_U198;
wire P3_ADD_371_1212_U199 , P3_ADD_371_1212_U200 , P3_ADD_371_1212_U201 , P3_ADD_371_1212_U202 , P3_ADD_371_1212_U203 , P3_ADD_371_1212_U204 , P3_ADD_371_1212_U205 , P3_ADD_371_1212_U206 , P3_ADD_371_1212_U207 , P3_ADD_371_1212_U208;
wire P3_ADD_371_1212_U209 , P3_ADD_371_1212_U210 , P3_ADD_371_1212_U211 , P3_ADD_371_1212_U212 , P3_ADD_371_1212_U213 , P3_ADD_371_1212_U214 , P3_ADD_371_1212_U215 , P3_ADD_371_1212_U216 , P3_ADD_371_1212_U217 , P3_ADD_371_1212_U218;
wire P3_ADD_371_1212_U219 , P3_ADD_371_1212_U220 , P3_ADD_371_1212_U221 , P3_ADD_371_1212_U222 , P3_ADD_371_1212_U223 , P3_ADD_371_1212_U224 , P3_ADD_371_1212_U225 , P3_ADD_371_1212_U226 , P3_ADD_371_1212_U227 , P3_ADD_371_1212_U228;
wire P3_ADD_371_1212_U229 , P3_ADD_371_1212_U230 , P3_ADD_371_1212_U231 , P3_ADD_371_1212_U232 , P3_ADD_371_1212_U233 , P3_ADD_371_1212_U234 , P3_ADD_371_1212_U235 , P3_ADD_371_1212_U236 , P3_ADD_371_1212_U237 , P3_ADD_371_1212_U238;
wire P3_ADD_371_1212_U239 , P3_ADD_371_1212_U240 , P3_ADD_371_1212_U241 , P3_ADD_371_1212_U242 , P3_ADD_371_1212_U243 , P3_ADD_371_1212_U244 , P3_ADD_371_1212_U245 , P3_ADD_371_1212_U246 , P3_ADD_371_1212_U247 , P3_ADD_371_1212_U248;
wire P3_ADD_371_1212_U249 , P3_ADD_371_1212_U250 , P3_ADD_371_1212_U251 , P3_ADD_371_1212_U252 , P3_ADD_371_1212_U253 , P3_ADD_371_1212_U254 , P3_ADD_371_1212_U255 , P3_ADD_371_1212_U256 , P3_ADD_371_1212_U257 , P3_ADD_371_1212_U258;
wire P3_ADD_371_1212_U259 , P3_ADD_371_1212_U260 , P3_ADD_371_1212_U261 , P3_ADD_371_1212_U262 , P3_ADD_371_1212_U263 , P3_ADD_371_1212_U264 , P3_ADD_371_1212_U265 , P3_SUB_504_U6 , P3_SUB_504_U7 , P3_SUB_504_U8;
wire P3_SUB_504_U9 , P3_SUB_504_U10 , P3_SUB_504_U11 , P3_SUB_504_U12 , P3_SUB_504_U13 , P3_SUB_504_U14 , P3_SUB_504_U15 , P3_SUB_504_U16 , P3_SUB_504_U17 , P3_SUB_504_U18;
wire P3_SUB_504_U19 , P3_SUB_504_U20 , P3_SUB_504_U21 , P3_SUB_504_U22 , P3_SUB_504_U23 , P3_SUB_504_U24 , P3_SUB_504_U25 , P3_SUB_504_U26 , P3_SUB_504_U27 , P3_SUB_504_U28;
wire P3_SUB_504_U29 , P3_SUB_504_U30 , P3_SUB_504_U31 , P3_SUB_504_U32 , P3_SUB_504_U33 , P3_SUB_504_U34 , P3_SUB_504_U35 , P3_SUB_504_U36 , P3_SUB_504_U37 , P3_SUB_504_U38;
wire P3_SUB_504_U39 , P3_SUB_504_U40 , P3_SUB_504_U41 , P3_SUB_504_U42 , P3_SUB_504_U43 , P3_SUB_504_U44 , P3_SUB_504_U45 , P3_SUB_504_U46 , P3_SUB_504_U47 , P3_SUB_504_U48;
wire P3_SUB_504_U49 , P3_SUB_504_U50 , P3_SUB_504_U51 , P3_SUB_504_U52 , P3_SUB_504_U53 , P3_SUB_504_U54 , P3_SUB_504_U55 , P3_SUB_504_U56 , P3_SUB_504_U57 , P3_SUB_504_U58;
wire P3_SUB_504_U59 , P3_SUB_504_U60 , P3_SUB_504_U61 , P3_SUB_504_U62 , P3_SUB_504_U63 , P3_SUB_401_U6 , P3_SUB_401_U7 , P3_SUB_401_U8 , P3_SUB_401_U9 , P3_SUB_401_U10;
wire P3_SUB_401_U11 , P3_SUB_401_U12 , P3_SUB_401_U13 , P3_SUB_401_U14 , P3_SUB_401_U15 , P3_SUB_401_U16 , P3_SUB_401_U17 , P3_SUB_401_U18 , P3_SUB_401_U19 , P3_SUB_401_U20;
wire P3_SUB_401_U21 , P3_SUB_401_U22 , P3_SUB_401_U23 , P3_SUB_401_U24 , P3_SUB_401_U25 , P3_SUB_401_U26 , P3_SUB_401_U27 , P3_SUB_401_U28 , P3_SUB_401_U29 , P3_SUB_401_U30;
wire P3_SUB_401_U31 , P3_SUB_401_U32 , P3_SUB_401_U33 , P3_SUB_401_U34 , P3_SUB_401_U35 , P3_SUB_401_U36 , P3_SUB_401_U37 , P3_SUB_401_U38 , P3_SUB_401_U39 , P3_SUB_401_U40;
wire P3_SUB_401_U41 , P3_SUB_401_U42 , P3_SUB_401_U43 , P3_SUB_401_U44 , P3_SUB_401_U45 , P3_SUB_401_U46 , P3_SUB_401_U47 , P3_SUB_401_U48 , P3_SUB_401_U49 , P3_SUB_401_U50;
wire P3_SUB_401_U51 , P3_SUB_401_U52 , P3_SUB_401_U53 , P3_SUB_401_U54 , P3_SUB_401_U55 , P3_SUB_401_U56 , P3_SUB_401_U57 , P3_SUB_401_U58 , P3_SUB_401_U59 , P3_SUB_401_U60;
wire P3_SUB_401_U61 , P3_SUB_401_U62 , P3_SUB_401_U63 , P3_SUB_401_U64 , P3_SUB_401_U65 , P3_SUB_401_U66 , P3_ADD_371_U4 , P3_ADD_371_U5 , P3_ADD_371_U6 , P3_ADD_371_U7;
wire P3_ADD_371_U8 , P3_ADD_371_U9 , P3_ADD_371_U10 , P3_ADD_371_U11 , P3_ADD_371_U12 , P3_ADD_371_U13 , P3_ADD_371_U14 , P3_ADD_371_U15 , P3_ADD_371_U16 , P3_ADD_371_U17;
wire P3_ADD_371_U18 , P3_ADD_371_U19 , P3_ADD_371_U20 , P3_ADD_371_U21 , P3_ADD_371_U22 , P3_ADD_371_U23 , P3_ADD_371_U24 , P3_ADD_371_U25 , P3_ADD_371_U26 , P3_ADD_371_U27;
wire P3_ADD_371_U28 , P3_ADD_371_U29 , P3_ADD_371_U30 , P3_ADD_371_U31 , P3_ADD_371_U32 , P3_ADD_371_U33 , P3_ADD_371_U34 , P3_ADD_371_U35 , P3_ADD_371_U36 , P3_ADD_371_U37;
wire P3_ADD_371_U38 , P3_ADD_371_U39 , P3_ADD_371_U40 , P3_ADD_371_U41 , P3_ADD_371_U42 , P3_ADD_371_U43 , P3_ADD_371_U44 , P3_SUB_390_U6 , P3_SUB_390_U7 , P3_SUB_390_U8;
wire P3_SUB_390_U9 , P3_SUB_390_U10 , P3_SUB_390_U11 , P3_SUB_390_U12 , P3_SUB_390_U13 , P3_SUB_390_U14 , P3_SUB_390_U15 , P3_SUB_390_U16 , P3_SUB_390_U17 , P3_SUB_390_U18;
wire P3_SUB_390_U19 , P3_SUB_390_U20 , P3_SUB_390_U21 , P3_SUB_390_U22 , P3_SUB_390_U23 , P3_SUB_390_U24 , P3_SUB_390_U25 , P3_SUB_390_U26 , P3_SUB_390_U27 , P3_SUB_390_U28;
wire P3_SUB_390_U29 , P3_SUB_390_U30 , P3_SUB_390_U31 , P3_SUB_390_U32 , P3_SUB_390_U33 , P3_SUB_390_U34 , P3_SUB_390_U35 , P3_SUB_390_U36 , P3_SUB_390_U37 , P3_SUB_390_U38;
wire P3_SUB_390_U39 , P3_SUB_390_U40 , P3_SUB_390_U41 , P3_SUB_390_U42 , P3_SUB_390_U43 , P3_SUB_390_U44 , P3_SUB_390_U45 , P3_SUB_390_U46 , P3_SUB_390_U47 , P3_SUB_390_U48;
wire P3_SUB_390_U49 , P3_SUB_390_U50 , P3_SUB_390_U51 , P3_SUB_390_U52 , P3_SUB_390_U53 , P3_SUB_390_U54 , P3_SUB_390_U55 , P3_SUB_390_U56 , P3_SUB_390_U57 , P3_SUB_390_U58;
wire P3_SUB_390_U59 , P3_SUB_390_U60 , P3_SUB_390_U61 , P3_SUB_390_U62 , P3_SUB_390_U63 , P3_SUB_390_U64 , P3_SUB_390_U65 , P3_SUB_390_U66 , P3_SUB_357_U6 , P3_SUB_357_U7;
wire P3_SUB_357_U8 , P3_SUB_357_U9 , P3_SUB_357_U10 , P3_SUB_357_U11 , P3_SUB_357_U12 , P3_SUB_357_U13 , P3_ADD_495_U4 , P3_ADD_495_U5 , P3_ADD_495_U6 , P3_ADD_495_U7;
wire P3_ADD_495_U8 , P3_ADD_495_U9 , P3_ADD_495_U10 , P3_ADD_495_U11 , P3_ADD_495_U12 , P3_ADD_495_U13 , P3_ADD_495_U14 , P3_ADD_495_U15 , P3_ADD_495_U16 , P3_ADD_495_U17;
wire P3_ADD_495_U18 , P3_ADD_495_U19 , P3_ADD_495_U20 , P3_GTE_412_U6 , P3_GTE_412_U7 , P3_GTE_504_U6 , P3_GTE_504_U7 , P3_ADD_494_U4 , P3_ADD_494_U5 , P3_ADD_494_U6;
wire P3_ADD_494_U7 , P3_ADD_494_U8 , P3_ADD_494_U9 , P3_ADD_494_U10 , P3_ADD_494_U11 , P3_ADD_494_U12 , P3_ADD_494_U13 , P3_ADD_494_U14 , P3_ADD_494_U15 , P3_ADD_494_U16;
wire P3_ADD_494_U17 , P3_ADD_494_U18 , P3_ADD_494_U19 , P3_ADD_494_U20 , P3_ADD_494_U21 , P3_ADD_494_U22 , P3_ADD_494_U23 , P3_ADD_494_U24 , P3_ADD_494_U25 , P3_ADD_494_U26;
wire P3_ADD_494_U27 , P3_ADD_494_U28 , P3_ADD_494_U29 , P3_ADD_494_U30 , P3_ADD_494_U31 , P3_ADD_494_U32 , P3_ADD_494_U33 , P3_ADD_494_U34 , P3_ADD_494_U35 , P3_ADD_494_U36;
wire P3_ADD_494_U37 , P3_ADD_494_U38 , P3_ADD_494_U39 , P3_ADD_494_U40 , P3_ADD_494_U41 , P3_ADD_494_U42 , P3_ADD_494_U43 , P3_ADD_494_U44 , P3_ADD_494_U45 , P3_ADD_494_U46;
wire P3_ADD_494_U47 , P3_ADD_494_U48 , P3_ADD_494_U49 , P3_ADD_494_U50 , P3_ADD_494_U51 , P3_ADD_494_U52 , P3_ADD_494_U53 , P3_ADD_494_U54 , P3_ADD_494_U55 , P3_ADD_494_U56;
wire P3_ADD_494_U57 , P3_ADD_494_U58 , P3_ADD_494_U59 , P3_ADD_494_U60 , P3_ADD_494_U61 , P3_ADD_494_U62 , P3_ADD_494_U63 , P3_ADD_494_U64 , P3_ADD_494_U65 , P3_ADD_494_U66;
wire P3_ADD_494_U67 , P3_ADD_494_U68 , P3_ADD_494_U69 , P3_ADD_494_U70 , P3_ADD_494_U71 , P3_ADD_494_U72 , P3_ADD_494_U73 , P3_ADD_494_U74 , P3_ADD_494_U75 , P3_ADD_494_U76;
wire P3_ADD_494_U77 , P3_ADD_494_U78 , P3_ADD_494_U79 , P3_ADD_494_U80 , P3_ADD_494_U81 , P3_ADD_494_U82 , P3_ADD_494_U83 , P3_ADD_494_U84 , P3_ADD_494_U85 , P3_ADD_494_U86;
wire P3_ADD_494_U87 , P3_ADD_494_U88 , P3_ADD_494_U89 , P3_ADD_494_U90 , P3_ADD_494_U91 , P3_ADD_494_U92 , P3_ADD_494_U93 , P3_ADD_494_U94 , P3_ADD_494_U95 , P3_ADD_494_U96;
wire P3_ADD_494_U97 , P3_ADD_494_U98 , P3_ADD_494_U99 , P3_ADD_494_U100 , P3_ADD_494_U101 , P3_ADD_494_U102 , P3_ADD_494_U103 , P3_ADD_494_U104 , P3_ADD_494_U105 , P3_ADD_494_U106;
wire P3_ADD_494_U107 , P3_ADD_494_U108 , P3_ADD_494_U109 , P3_ADD_494_U110 , P3_ADD_494_U111 , P3_ADD_494_U112 , P3_ADD_494_U113 , P3_ADD_494_U114 , P3_ADD_494_U115 , P3_ADD_494_U116;
wire P3_ADD_494_U117 , P3_ADD_494_U118 , P3_ADD_494_U119 , P3_ADD_494_U120 , P3_ADD_494_U121 , P3_ADD_494_U122 , P3_ADD_494_U123 , P3_ADD_494_U124 , P3_ADD_494_U125 , P3_ADD_494_U126;
wire P3_ADD_494_U127 , P3_ADD_494_U128 , P3_ADD_494_U129 , P3_ADD_494_U130 , P3_ADD_494_U131 , P3_ADD_494_U132 , P3_ADD_494_U133 , P3_ADD_494_U134 , P3_ADD_494_U135 , P3_ADD_494_U136;
wire P3_ADD_494_U137 , P3_ADD_494_U138 , P3_ADD_494_U139 , P3_ADD_494_U140 , P3_ADD_494_U141 , P3_ADD_494_U142 , P3_ADD_494_U143 , P3_ADD_494_U144 , P3_ADD_494_U145 , P3_ADD_494_U146;
wire P3_ADD_494_U147 , P3_ADD_494_U148 , P3_ADD_494_U149 , P3_ADD_494_U150 , P3_ADD_494_U151 , P3_ADD_494_U152 , P3_ADD_494_U153 , P3_ADD_494_U154 , P3_ADD_494_U155 , P3_ADD_494_U156;
wire P3_ADD_494_U157 , P3_ADD_494_U158 , P3_ADD_494_U159 , P3_ADD_494_U160 , P3_ADD_494_U161 , P3_ADD_494_U162 , P3_ADD_494_U163 , P3_ADD_494_U164 , P3_ADD_494_U165 , P3_ADD_494_U166;
wire P3_ADD_494_U167 , P3_ADD_494_U168 , P3_ADD_494_U169 , P3_ADD_494_U170 , P3_ADD_494_U171 , P3_ADD_494_U172 , P3_ADD_494_U173 , P3_ADD_494_U174 , P3_ADD_494_U175 , P3_ADD_494_U176;
wire P3_ADD_494_U177 , P3_ADD_494_U178 , P3_ADD_494_U179 , P3_ADD_494_U180 , P3_ADD_494_U181 , P3_ADD_494_U182 , P3_ADD_536_U4 , P3_ADD_536_U5 , P3_ADD_536_U6 , P3_ADD_536_U7;
wire P3_ADD_536_U8 , P3_ADD_536_U9 , P3_ADD_536_U10 , P3_ADD_536_U11 , P3_ADD_536_U12 , P3_ADD_536_U13 , P3_ADD_536_U14 , P3_ADD_536_U15 , P3_ADD_536_U16 , P3_ADD_536_U17;
wire P3_ADD_536_U18 , P3_ADD_536_U19 , P3_ADD_536_U20 , P3_ADD_536_U21 , P3_ADD_536_U22 , P3_ADD_536_U23 , P3_ADD_536_U24 , P3_ADD_536_U25 , P3_ADD_536_U26 , P3_ADD_536_U27;
wire P3_ADD_536_U28 , P3_ADD_536_U29 , P3_ADD_536_U30 , P3_ADD_536_U31 , P3_ADD_536_U32 , P3_ADD_536_U33 , P3_ADD_536_U34 , P3_ADD_536_U35 , P3_ADD_536_U36 , P3_ADD_536_U37;
wire P3_ADD_536_U38 , P3_ADD_536_U39 , P3_ADD_536_U40 , P3_ADD_536_U41 , P3_ADD_536_U42 , P3_ADD_536_U43 , P3_ADD_536_U44 , P3_ADD_536_U45 , P3_ADD_536_U46 , P3_ADD_536_U47;
wire P3_ADD_536_U48 , P3_ADD_536_U49 , P3_ADD_536_U50 , P3_ADD_536_U51 , P3_ADD_536_U52 , P3_ADD_536_U53 , P3_ADD_536_U54 , P3_ADD_536_U55 , P3_ADD_536_U56 , P3_ADD_536_U57;
wire P3_ADD_536_U58 , P3_ADD_536_U59 , P3_ADD_536_U60 , P3_ADD_536_U61 , P3_ADD_536_U62 , P3_ADD_536_U63 , P3_ADD_536_U64 , P3_ADD_536_U65 , P3_ADD_536_U66 , P3_ADD_536_U67;
wire P3_ADD_536_U68 , P3_ADD_536_U69 , P3_ADD_536_U70 , P3_ADD_536_U71 , P3_ADD_536_U72 , P3_ADD_536_U73 , P3_ADD_536_U74 , P3_ADD_536_U75 , P3_ADD_536_U76 , P3_ADD_536_U77;
wire P3_ADD_536_U78 , P3_ADD_536_U79 , P3_ADD_536_U80 , P3_ADD_536_U81 , P3_ADD_536_U82 , P3_ADD_536_U83 , P3_ADD_536_U84 , P3_ADD_536_U85 , P3_ADD_536_U86 , P3_ADD_536_U87;
wire P3_ADD_536_U88 , P3_ADD_536_U89 , P3_ADD_536_U90 , P3_ADD_536_U91 , P3_ADD_536_U92 , P3_ADD_536_U93 , P3_ADD_536_U94 , P3_ADD_536_U95 , P3_ADD_536_U96 , P3_ADD_536_U97;
wire P3_ADD_536_U98 , P3_ADD_536_U99 , P3_ADD_536_U100 , P3_ADD_536_U101 , P3_ADD_536_U102 , P3_ADD_536_U103 , P3_ADD_536_U104 , P3_ADD_536_U105 , P3_ADD_536_U106 , P3_ADD_536_U107;
wire P3_ADD_536_U108 , P3_ADD_536_U109 , P3_ADD_536_U110 , P3_ADD_536_U111 , P3_ADD_536_U112 , P3_ADD_536_U113 , P3_ADD_536_U114 , P3_ADD_536_U115 , P3_ADD_536_U116 , P3_ADD_536_U117;
wire P3_ADD_536_U118 , P3_ADD_536_U119 , P3_ADD_536_U120 , P3_ADD_536_U121 , P3_ADD_536_U122 , P3_ADD_536_U123 , P3_ADD_536_U124 , P3_ADD_536_U125 , P3_ADD_536_U126 , P3_ADD_536_U127;
wire P3_ADD_536_U128 , P3_ADD_536_U129 , P3_ADD_536_U130 , P3_ADD_536_U131 , P3_ADD_536_U132 , P3_ADD_536_U133 , P3_ADD_536_U134 , P3_ADD_536_U135 , P3_ADD_536_U136 , P3_ADD_536_U137;
wire P3_ADD_536_U138 , P3_ADD_536_U139 , P3_ADD_536_U140 , P3_ADD_536_U141 , P3_ADD_536_U142 , P3_ADD_536_U143 , P3_ADD_536_U144 , P3_ADD_536_U145 , P3_ADD_536_U146 , P3_ADD_536_U147;
wire P3_ADD_536_U148 , P3_ADD_536_U149 , P3_ADD_536_U150 , P3_ADD_536_U151 , P3_ADD_536_U152 , P3_ADD_536_U153 , P3_ADD_536_U154 , P3_ADD_536_U155 , P3_ADD_536_U156 , P3_ADD_536_U157;
wire P3_ADD_536_U158 , P3_ADD_536_U159 , P3_ADD_536_U160 , P3_ADD_536_U161 , P3_ADD_536_U162 , P3_ADD_536_U163 , P3_ADD_536_U164 , P3_ADD_536_U165 , P3_ADD_536_U166 , P3_ADD_536_U167;
wire P3_ADD_536_U168 , P3_ADD_536_U169 , P3_ADD_536_U170 , P3_ADD_536_U171 , P3_ADD_536_U172 , P3_ADD_536_U173 , P3_ADD_536_U174 , P3_ADD_536_U175 , P3_ADD_536_U176 , P3_ADD_536_U177;
wire P3_ADD_536_U178 , P3_ADD_536_U179 , P3_ADD_536_U180 , P3_ADD_536_U181 , P3_ADD_536_U182 , P3_ADD_402_1132_U4 , P3_ADD_402_1132_U5 , P3_ADD_402_1132_U6 , P3_ADD_402_1132_U7 , P3_ADD_402_1132_U8;
wire P3_ADD_402_1132_U9 , P3_ADD_402_1132_U10 , P3_ADD_402_1132_U11 , P3_ADD_402_1132_U12 , P3_ADD_402_1132_U13 , P3_ADD_402_1132_U14 , P3_ADD_402_1132_U15 , P3_ADD_402_1132_U16 , P3_ADD_402_1132_U17 , P3_ADD_402_1132_U18;
wire P3_ADD_402_1132_U19 , P3_ADD_402_1132_U20 , P3_ADD_402_1132_U21 , P3_ADD_402_1132_U22 , P3_ADD_402_1132_U23 , P3_ADD_402_1132_U24 , P3_ADD_402_1132_U25 , P3_ADD_402_1132_U26 , P3_ADD_402_1132_U27 , P3_ADD_402_1132_U28;
wire P3_ADD_402_1132_U29 , P3_ADD_402_1132_U30 , P3_ADD_402_1132_U31 , P3_ADD_402_1132_U32 , P3_ADD_402_1132_U33 , P3_ADD_402_1132_U34 , P3_ADD_402_1132_U35 , P3_ADD_402_1132_U36 , P3_ADD_402_1132_U37 , P3_ADD_402_1132_U38;
wire P3_ADD_402_1132_U39 , P3_ADD_402_1132_U40 , P3_ADD_402_1132_U41 , P3_ADD_402_1132_U42 , P3_ADD_402_1132_U43 , P3_ADD_402_1132_U44 , P3_ADD_402_1132_U45 , P3_ADD_402_1132_U46 , P3_ADD_402_1132_U47 , P3_ADD_402_1132_U48;
wire P3_ADD_402_1132_U49 , P3_ADD_402_1132_U50 , P2_R2099_U5 , P2_R2099_U6 , P2_R2099_U7 , P2_R2099_U8 , P2_R2099_U9 , P2_R2099_U10 , P2_R2099_U11 , P2_R2099_U12;
wire P2_R2099_U13 , P2_R2099_U14 , P2_R2099_U15 , P2_R2099_U16 , P2_R2099_U17 , P2_R2099_U18 , P2_R2099_U19 , P2_R2099_U20 , P2_R2099_U21 , P2_R2099_U22;
wire P2_R2099_U23 , P2_R2099_U24 , P2_R2099_U25 , P2_R2099_U26 , P2_R2099_U27 , P2_R2099_U28 , P2_R2099_U29 , P2_R2099_U30 , P2_R2099_U31 , P2_R2099_U32;
wire P2_R2099_U33 , P2_R2099_U34 , P2_R2099_U35 , P2_R2099_U36 , P2_R2099_U37 , P2_R2099_U38 , P2_R2099_U39 , P2_R2099_U40 , P2_R2099_U41 , P2_R2099_U42;
wire P2_R2099_U43 , P2_R2099_U44 , P2_R2099_U45 , P2_R2099_U46 , P2_R2099_U47 , P2_R2099_U48 , P2_R2099_U49 , P2_R2099_U50 , P2_R2099_U51 , P2_R2099_U52;
wire P2_R2099_U53 , P2_R2099_U54 , P2_R2099_U55 , P2_R2099_U56 , P2_R2099_U57 , P2_R2099_U58 , P2_R2099_U59 , P2_R2099_U60 , P2_R2099_U61 , P2_R2099_U62;
wire P2_R2099_U63 , P2_R2099_U64 , P2_R2099_U65 , P2_R2099_U66 , P2_R2099_U67 , P2_R2099_U68 , P2_R2099_U69 , P2_R2099_U70 , P2_R2099_U71 , P2_R2099_U72;
wire P2_R2099_U73 , P2_R2099_U74 , P2_R2099_U75 , P2_R2099_U76 , P2_R2099_U77 , P2_R2099_U78 , P2_R2099_U79 , P2_R2099_U80 , P2_R2099_U81 , P2_R2099_U82;
wire P2_R2099_U83 , P2_R2099_U84 , P2_R2099_U85 , P2_R2099_U86 , P2_R2099_U87 , P2_R2099_U88 , P2_R2099_U89 , P2_R2099_U90 , P2_R2099_U91 , P2_R2099_U92;
wire P2_R2099_U93 , P2_R2099_U94 , P2_R2099_U95 , P2_R2099_U96 , P2_R2099_U97 , P2_R2099_U98 , P2_R2099_U99 , P2_R2099_U100 , P2_R2099_U101 , P2_R2099_U102;
wire P2_R2099_U103 , P2_R2099_U104 , P2_R2099_U105 , P2_R2099_U106 , P2_R2099_U107 , P2_R2099_U108 , P2_R2099_U109 , P2_R2099_U110 , P2_R2099_U111 , P2_R2099_U112;
wire P2_R2099_U113 , P2_R2099_U114 , P2_R2099_U115 , P2_R2099_U116 , P2_R2099_U117 , P2_R2099_U118 , P2_R2099_U119 , P2_R2099_U120 , P2_R2099_U121 , P2_R2099_U122;
wire P2_R2099_U123 , P2_R2099_U124 , P2_R2099_U125 , P2_R2099_U126 , P2_R2099_U127 , P2_R2099_U128 , P2_R2099_U129 , P2_R2099_U130 , P2_R2099_U131 , P2_R2099_U132;
wire P2_R2099_U133 , P2_R2099_U134 , P2_R2099_U135 , P2_R2099_U136 , P2_R2099_U137 , P2_R2099_U138 , P2_R2099_U139 , P2_R2099_U140 , P2_R2099_U141 , P2_R2099_U142;
wire P2_R2099_U143 , P2_R2099_U144 , P2_R2099_U145 , P2_R2099_U146 , P2_R2099_U147 , P2_R2099_U148 , P2_R2099_U149 , P2_R2099_U150 , P2_R2099_U151 , P2_R2099_U152;
wire P2_R2099_U153 , P2_R2099_U154 , P2_R2099_U155 , P2_R2099_U156 , P2_R2099_U157 , P2_R2099_U158 , P2_R2099_U159 , P2_R2099_U160 , P2_R2099_U161 , P2_R2099_U162;
wire P2_R2099_U163 , P2_R2099_U164 , P2_R2099_U165 , P2_R2099_U166 , P2_R2099_U167 , P2_R2099_U168 , P2_R2099_U169 , P2_R2099_U170 , P2_R2099_U171 , P2_R2099_U172;
wire P2_R2099_U173 , P2_R2099_U174 , P2_R2099_U175 , P2_R2099_U176 , P2_R2099_U177 , P2_R2099_U178 , P2_R2099_U179 , P2_R2099_U180 , P2_R2099_U181 , P2_R2099_U182;
wire P2_R2099_U183 , P2_R2099_U184 , P2_R2099_U185 , P2_R2099_U186 , P2_R2099_U187 , P2_R2099_U188 , P2_R2099_U189 , P2_R2099_U190 , P2_R2099_U191 , P2_R2099_U192;
wire P2_R2099_U193 , P2_R2099_U194 , P2_R2099_U195 , P2_R2099_U196 , P2_R2099_U197 , P2_R2099_U198 , P2_R2099_U199 , P2_R2099_U200 , P2_R2099_U201 , P2_R2099_U202;
wire P2_R2099_U203 , P2_R2099_U204 , P2_R2099_U205 , P2_R2099_U206 , P2_R2099_U207 , P2_R2099_U208 , P2_R2099_U209 , P2_R2099_U210 , P2_R2099_U211 , P2_R2099_U212;
wire P2_R2099_U213 , P2_R2099_U214 , P2_R2099_U215 , P2_R2099_U216 , P2_R2099_U217 , P2_R2099_U218 , P2_R2099_U219 , P2_R2099_U220 , P2_R2099_U221 , P2_R2099_U222;
wire P2_R2099_U223 , P2_R2099_U224 , P2_R2099_U225 , P2_ADD_391_1196_U5 , P2_ADD_391_1196_U6 , P2_ADD_391_1196_U7 , P2_ADD_391_1196_U8 , P2_ADD_391_1196_U9 , P2_ADD_391_1196_U10 , P2_ADD_391_1196_U11;
wire P2_ADD_391_1196_U12 , P2_ADD_391_1196_U13 , P2_ADD_391_1196_U14 , P2_ADD_391_1196_U15 , P2_ADD_391_1196_U16 , P2_ADD_391_1196_U17 , P2_ADD_391_1196_U18 , P2_ADD_391_1196_U19 , P2_ADD_391_1196_U20 , P2_ADD_391_1196_U21;
wire P2_ADD_391_1196_U22 , P2_ADD_391_1196_U23 , P2_ADD_391_1196_U24 , P2_ADD_391_1196_U25 , P2_ADD_391_1196_U26 , P2_ADD_391_1196_U27 , P2_ADD_391_1196_U28 , P2_ADD_391_1196_U29 , P2_ADD_391_1196_U30 , P2_ADD_391_1196_U31;
wire P2_ADD_391_1196_U32 , P2_ADD_391_1196_U33 , P2_ADD_391_1196_U34 , P2_ADD_391_1196_U35 , P2_ADD_391_1196_U36 , P2_ADD_391_1196_U37 , P2_ADD_391_1196_U38 , P2_ADD_391_1196_U39 , P2_ADD_391_1196_U40 , P2_ADD_391_1196_U41;
wire P2_ADD_391_1196_U42 , P2_ADD_391_1196_U43 , P2_ADD_391_1196_U44 , P2_ADD_391_1196_U45 , P2_ADD_391_1196_U46 , P2_ADD_391_1196_U47 , P2_ADD_391_1196_U48 , P2_ADD_391_1196_U49 , P2_ADD_391_1196_U50 , P2_ADD_391_1196_U51;
wire P2_ADD_391_1196_U52 , P2_ADD_391_1196_U53 , P2_ADD_391_1196_U54 , P2_ADD_391_1196_U55 , P2_ADD_391_1196_U56 , P2_ADD_391_1196_U57 , P2_ADD_391_1196_U58 , P2_ADD_391_1196_U59 , P2_ADD_391_1196_U60 , P2_ADD_391_1196_U61;
wire P2_ADD_391_1196_U62 , P2_ADD_391_1196_U63 , P2_ADD_391_1196_U64 , P2_ADD_391_1196_U65 , P2_ADD_391_1196_U66 , P2_ADD_391_1196_U67 , P2_ADD_391_1196_U68 , P2_ADD_391_1196_U69 , P2_ADD_391_1196_U70 , P2_ADD_391_1196_U71;
wire P2_ADD_391_1196_U72 , P2_ADD_391_1196_U73 , P2_ADD_391_1196_U74 , P2_ADD_391_1196_U75 , P2_ADD_391_1196_U76 , P2_ADD_391_1196_U77 , P2_ADD_391_1196_U78 , P2_ADD_391_1196_U79 , P2_ADD_391_1196_U80 , P2_ADD_391_1196_U81;
wire P2_ADD_391_1196_U82 , P2_ADD_391_1196_U83 , P2_ADD_391_1196_U84 , P2_ADD_391_1196_U85 , P2_ADD_391_1196_U86 , P2_ADD_391_1196_U87 , P2_ADD_391_1196_U88 , P2_ADD_391_1196_U89 , P2_ADD_391_1196_U90 , P2_ADD_391_1196_U91;
wire P2_ADD_391_1196_U92 , P2_ADD_391_1196_U93 , P2_ADD_391_1196_U94 , P2_ADD_391_1196_U95 , P2_ADD_391_1196_U96 , P2_ADD_391_1196_U97 , P2_ADD_391_1196_U98 , P2_ADD_391_1196_U99 , P2_ADD_391_1196_U100 , P2_ADD_391_1196_U101;
wire P2_ADD_391_1196_U102 , P2_ADD_391_1196_U103 , P2_ADD_391_1196_U104 , P2_ADD_391_1196_U105 , P2_ADD_391_1196_U106 , P2_ADD_391_1196_U107 , P2_ADD_391_1196_U108 , P2_ADD_391_1196_U109 , P2_ADD_391_1196_U110 , P2_ADD_391_1196_U111;
wire P2_ADD_391_1196_U112 , P2_ADD_391_1196_U113 , P2_ADD_391_1196_U114 , P2_ADD_391_1196_U115 , P2_ADD_391_1196_U116 , P2_ADD_391_1196_U117 , P2_ADD_391_1196_U118 , P2_ADD_391_1196_U119 , P2_ADD_391_1196_U120 , P2_ADD_391_1196_U121;
wire P2_ADD_391_1196_U122 , P2_ADD_391_1196_U123 , P2_ADD_391_1196_U124 , P2_ADD_391_1196_U125 , P2_ADD_391_1196_U126 , P2_ADD_391_1196_U127 , P2_ADD_391_1196_U128 , P2_ADD_391_1196_U129 , P2_ADD_391_1196_U130 , P2_ADD_391_1196_U131;
wire P2_ADD_391_1196_U132 , P2_ADD_391_1196_U133 , P2_ADD_391_1196_U134 , P2_ADD_391_1196_U135 , P2_ADD_391_1196_U136 , P2_ADD_391_1196_U137 , P2_ADD_391_1196_U138 , P2_ADD_391_1196_U139 , P2_ADD_391_1196_U140 , P2_ADD_391_1196_U141;
wire P2_ADD_391_1196_U142 , P2_ADD_391_1196_U143 , P2_ADD_391_1196_U144 , P2_ADD_391_1196_U145 , P2_ADD_391_1196_U146 , P2_ADD_391_1196_U147 , P2_ADD_391_1196_U148 , P2_ADD_391_1196_U149 , P2_ADD_391_1196_U150 , P2_ADD_391_1196_U151;
wire P2_ADD_391_1196_U152 , P2_ADD_391_1196_U153 , P2_ADD_391_1196_U154 , P2_ADD_391_1196_U155 , P2_ADD_391_1196_U156 , P2_ADD_391_1196_U157 , P2_ADD_391_1196_U158 , P2_ADD_391_1196_U159 , P2_ADD_391_1196_U160 , P2_ADD_391_1196_U161;
wire P2_ADD_391_1196_U162 , P2_ADD_391_1196_U163 , P2_ADD_391_1196_U164 , P2_ADD_391_1196_U165 , P2_ADD_391_1196_U166 , P2_ADD_391_1196_U167 , P2_ADD_391_1196_U168 , P2_ADD_391_1196_U169 , P2_ADD_391_1196_U170 , P2_ADD_391_1196_U171;
wire P2_ADD_391_1196_U172 , P2_ADD_391_1196_U173 , P2_ADD_391_1196_U174 , P2_ADD_391_1196_U175 , P2_ADD_391_1196_U176 , P2_ADD_391_1196_U177 , P2_ADD_391_1196_U178 , P2_ADD_391_1196_U179 , P2_ADD_391_1196_U180 , P2_ADD_391_1196_U181;
wire P2_ADD_391_1196_U182 , P2_ADD_391_1196_U183 , P2_ADD_391_1196_U184 , P2_ADD_391_1196_U185 , P2_ADD_391_1196_U186 , P2_ADD_391_1196_U187 , P2_ADD_391_1196_U188 , P2_ADD_391_1196_U189 , P2_ADD_391_1196_U190 , P2_ADD_391_1196_U191;
wire P2_ADD_391_1196_U192 , P2_ADD_391_1196_U193 , P2_ADD_391_1196_U194 , P2_ADD_391_1196_U195 , P2_ADD_391_1196_U196 , P2_ADD_391_1196_U197 , P2_ADD_391_1196_U198 , P2_ADD_391_1196_U199 , P2_ADD_391_1196_U200 , P2_ADD_391_1196_U201;
wire P2_ADD_391_1196_U202 , P2_ADD_391_1196_U203 , P2_ADD_391_1196_U204 , P2_ADD_391_1196_U205 , P2_ADD_391_1196_U206 , P2_ADD_391_1196_U207 , P2_ADD_391_1196_U208 , P2_ADD_391_1196_U209 , P2_ADD_391_1196_U210 , P2_ADD_391_1196_U211;
wire P2_ADD_391_1196_U212 , P2_ADD_391_1196_U213 , P2_ADD_391_1196_U214 , P2_ADD_391_1196_U215 , P2_ADD_391_1196_U216 , P2_ADD_391_1196_U217 , P2_ADD_391_1196_U218 , P2_ADD_391_1196_U219 , P2_ADD_391_1196_U220 , P2_ADD_391_1196_U221;
wire P2_ADD_391_1196_U222 , P2_ADD_391_1196_U223 , P2_ADD_391_1196_U224 , P2_ADD_391_1196_U225 , P2_ADD_391_1196_U226 , P2_ADD_391_1196_U227 , P2_ADD_391_1196_U228 , P2_ADD_391_1196_U229 , P2_ADD_391_1196_U230 , P2_ADD_391_1196_U231;
wire P2_ADD_391_1196_U232 , P2_ADD_391_1196_U233 , P2_ADD_391_1196_U234 , P2_ADD_391_1196_U235 , P2_ADD_391_1196_U236 , P2_ADD_391_1196_U237 , P2_ADD_391_1196_U238 , P2_ADD_391_1196_U239 , P2_ADD_391_1196_U240 , P2_ADD_391_1196_U241;
wire P2_ADD_391_1196_U242 , P2_ADD_391_1196_U243 , P2_ADD_391_1196_U244 , P2_ADD_391_1196_U245 , P2_ADD_391_1196_U246 , P2_ADD_391_1196_U247 , P2_ADD_391_1196_U248 , P2_ADD_391_1196_U249 , P2_ADD_391_1196_U250 , P2_ADD_391_1196_U251;
wire P2_ADD_391_1196_U252 , P2_ADD_391_1196_U253 , P2_ADD_391_1196_U254 , P2_ADD_391_1196_U255 , P2_ADD_391_1196_U256 , P2_ADD_391_1196_U257 , P2_ADD_391_1196_U258 , P2_ADD_391_1196_U259 , P2_ADD_391_1196_U260 , P2_ADD_391_1196_U261;
wire P2_ADD_391_1196_U262 , P2_ADD_391_1196_U263 , P2_ADD_391_1196_U264 , P2_ADD_391_1196_U265 , P2_ADD_391_1196_U266 , P2_ADD_391_1196_U267 , P2_ADD_391_1196_U268 , P2_ADD_391_1196_U269 , P2_ADD_391_1196_U270 , P2_ADD_391_1196_U271;
wire P2_ADD_391_1196_U272 , P2_ADD_391_1196_U273 , P2_ADD_391_1196_U274 , P2_ADD_391_1196_U275 , P2_ADD_391_1196_U276 , P2_ADD_391_1196_U277 , P2_ADD_391_1196_U278 , P2_ADD_391_1196_U279 , P2_ADD_391_1196_U280 , P2_ADD_391_1196_U281;
wire P2_ADD_391_1196_U282 , P2_ADD_391_1196_U283 , P2_ADD_391_1196_U284 , P2_ADD_391_1196_U285 , P2_ADD_391_1196_U286 , P2_ADD_391_1196_U287 , P2_ADD_391_1196_U288 , P2_ADD_391_1196_U289 , P2_ADD_391_1196_U290 , P2_ADD_391_1196_U291;
wire P2_ADD_391_1196_U292 , P2_ADD_391_1196_U293 , P2_ADD_391_1196_U294 , P2_ADD_391_1196_U295 , P2_ADD_391_1196_U296 , P2_ADD_391_1196_U297 , P2_ADD_391_1196_U298 , P2_ADD_391_1196_U299 , P2_ADD_391_1196_U300 , P2_ADD_391_1196_U301;
wire P2_ADD_391_1196_U302 , P2_ADD_391_1196_U303 , P2_ADD_391_1196_U304 , P2_ADD_391_1196_U305 , P2_ADD_391_1196_U306 , P2_ADD_391_1196_U307 , P2_ADD_391_1196_U308 , P2_ADD_391_1196_U309 , P2_ADD_391_1196_U310 , P2_ADD_391_1196_U311;
wire P2_ADD_391_1196_U312 , P2_ADD_391_1196_U313 , P2_ADD_391_1196_U314 , P2_ADD_391_1196_U315 , P2_ADD_391_1196_U316 , P2_ADD_391_1196_U317 , P2_ADD_391_1196_U318 , P2_ADD_391_1196_U319 , P2_ADD_391_1196_U320 , P2_ADD_391_1196_U321;
wire P2_ADD_391_1196_U322 , P2_ADD_391_1196_U323 , P2_ADD_391_1196_U324 , P2_ADD_391_1196_U325 , P2_ADD_391_1196_U326 , P2_ADD_391_1196_U327 , P2_ADD_391_1196_U328 , P2_ADD_391_1196_U329 , P2_ADD_391_1196_U330 , P2_ADD_391_1196_U331;
wire P2_ADD_391_1196_U332 , P2_ADD_391_1196_U333 , P2_ADD_391_1196_U334 , P2_ADD_391_1196_U335 , P2_ADD_391_1196_U336 , P2_ADD_391_1196_U337 , P2_ADD_391_1196_U338 , P2_ADD_391_1196_U339 , P2_ADD_391_1196_U340 , P2_ADD_391_1196_U341;
wire P2_ADD_391_1196_U342 , P2_ADD_391_1196_U343 , P2_ADD_391_1196_U344 , P2_ADD_391_1196_U345 , P2_ADD_391_1196_U346 , P2_ADD_391_1196_U347 , P2_ADD_391_1196_U348 , P2_ADD_391_1196_U349 , P2_ADD_391_1196_U350 , P2_ADD_391_1196_U351;
wire P2_ADD_391_1196_U352 , P2_ADD_391_1196_U353 , P2_ADD_391_1196_U354 , P2_ADD_391_1196_U355 , P2_ADD_391_1196_U356 , P2_ADD_391_1196_U357 , P2_ADD_391_1196_U358 , P2_ADD_391_1196_U359 , P2_ADD_391_1196_U360 , P2_ADD_391_1196_U361;
wire P2_ADD_391_1196_U362 , P2_ADD_391_1196_U363 , P2_ADD_391_1196_U364 , P2_ADD_391_1196_U365 , P2_ADD_391_1196_U366 , P2_ADD_391_1196_U367 , P2_ADD_391_1196_U368 , P2_ADD_391_1196_U369 , P2_ADD_391_1196_U370 , P2_ADD_391_1196_U371;
wire P2_ADD_391_1196_U372 , P2_ADD_391_1196_U373 , P2_ADD_391_1196_U374 , P2_ADD_391_1196_U375 , P2_ADD_391_1196_U376 , P2_ADD_391_1196_U377 , P2_ADD_391_1196_U378 , P2_ADD_391_1196_U379 , P2_ADD_391_1196_U380 , P2_ADD_391_1196_U381;
wire P2_ADD_391_1196_U382 , P2_ADD_391_1196_U383 , P2_ADD_391_1196_U384 , P2_ADD_391_1196_U385 , P2_ADD_391_1196_U386 , P2_ADD_391_1196_U387 , P2_ADD_391_1196_U388 , P2_ADD_391_1196_U389 , P2_ADD_391_1196_U390 , P2_ADD_391_1196_U391;
wire P2_ADD_391_1196_U392 , P2_ADD_391_1196_U393 , P2_ADD_391_1196_U394 , P2_ADD_391_1196_U395 , P2_ADD_391_1196_U396 , P2_ADD_391_1196_U397 , P2_ADD_391_1196_U398 , P2_ADD_391_1196_U399 , P2_ADD_391_1196_U400 , P2_ADD_391_1196_U401;
wire P2_ADD_391_1196_U402 , P2_ADD_391_1196_U403 , P2_ADD_391_1196_U404 , P2_ADD_391_1196_U405 , P2_ADD_391_1196_U406 , P2_ADD_391_1196_U407 , P2_ADD_391_1196_U408 , P2_ADD_391_1196_U409 , P2_ADD_391_1196_U410 , P2_ADD_391_1196_U411;
wire P2_ADD_391_1196_U412 , P2_ADD_391_1196_U413 , P2_ADD_391_1196_U414 , P2_ADD_391_1196_U415 , P2_ADD_391_1196_U416 , P2_ADD_391_1196_U417 , P2_ADD_391_1196_U418 , P2_ADD_391_1196_U419 , P2_ADD_391_1196_U420 , P2_ADD_391_1196_U421;
wire P2_ADD_391_1196_U422 , P2_ADD_391_1196_U423 , P2_ADD_391_1196_U424 , P2_ADD_391_1196_U425 , P2_ADD_391_1196_U426 , P2_ADD_391_1196_U427 , P2_ADD_391_1196_U428 , P2_ADD_391_1196_U429 , P2_ADD_391_1196_U430 , P2_ADD_391_1196_U431;
wire P2_ADD_391_1196_U432 , P2_ADD_391_1196_U433 , P2_ADD_391_1196_U434 , P2_ADD_391_1196_U435 , P2_ADD_391_1196_U436 , P2_ADD_391_1196_U437 , P2_ADD_391_1196_U438 , P2_ADD_391_1196_U439 , P2_ADD_391_1196_U440 , P2_ADD_391_1196_U441;
wire P2_ADD_391_1196_U442 , P2_ADD_391_1196_U443 , P2_ADD_391_1196_U444 , P2_ADD_391_1196_U445 , P2_ADD_391_1196_U446 , P2_ADD_391_1196_U447 , P2_ADD_391_1196_U448 , P2_ADD_391_1196_U449 , P2_ADD_391_1196_U450 , P2_ADD_391_1196_U451;
wire P2_ADD_391_1196_U452 , P2_ADD_391_1196_U453 , P2_ADD_391_1196_U454 , P2_ADD_391_1196_U455 , P2_ADD_391_1196_U456 , P2_ADD_391_1196_U457 , P2_ADD_391_1196_U458 , P2_ADD_391_1196_U459 , P2_ADD_391_1196_U460 , P2_ADD_391_1196_U461;
wire P2_ADD_391_1196_U462 , P2_ADD_391_1196_U463 , P2_ADD_391_1196_U464 , P2_ADD_391_1196_U465 , P2_ADD_391_1196_U466 , P2_ADD_391_1196_U467 , P2_ADD_391_1196_U468 , P2_ADD_391_1196_U469 , P2_ADD_391_1196_U470 , P2_ADD_391_1196_U471;
wire P2_ADD_391_1196_U472 , P2_ADD_391_1196_U473 , P2_ADD_391_1196_U474 , P2_ADD_391_1196_U475 , P2_ADD_391_1196_U476 , P2_ADD_391_1196_U477 , P2_ADD_391_1196_U478 , P2_ADD_402_1132_U4 , P2_ADD_402_1132_U5 , P2_ADD_402_1132_U6;
wire P2_ADD_402_1132_U7 , P2_ADD_402_1132_U8 , P2_ADD_402_1132_U9 , P2_ADD_402_1132_U10 , P2_ADD_402_1132_U11 , P2_ADD_402_1132_U12 , P2_ADD_402_1132_U13 , P2_ADD_402_1132_U14 , P2_ADD_402_1132_U15 , P2_ADD_402_1132_U16;
wire P2_ADD_402_1132_U17 , P2_ADD_402_1132_U18 , P2_ADD_402_1132_U19 , P2_ADD_402_1132_U20 , P2_ADD_402_1132_U21 , P2_ADD_402_1132_U22 , P2_ADD_402_1132_U23 , P2_ADD_402_1132_U24 , P2_ADD_402_1132_U25 , P2_ADD_402_1132_U26;
wire P2_ADD_402_1132_U27 , P2_ADD_402_1132_U28 , P2_ADD_402_1132_U29 , P2_ADD_402_1132_U30 , P2_ADD_402_1132_U31 , P2_ADD_402_1132_U32 , P2_ADD_402_1132_U33 , P2_ADD_402_1132_U34 , P2_ADD_402_1132_U35 , P2_ADD_402_1132_U36;
wire P2_ADD_402_1132_U37 , P2_ADD_402_1132_U38 , P2_ADD_402_1132_U39 , P2_ADD_402_1132_U40 , P2_ADD_402_1132_U41 , P2_ADD_402_1132_U42 , P2_ADD_402_1132_U43 , P2_ADD_402_1132_U44 , P2_ADD_402_1132_U45 , P2_ADD_402_1132_U46;
wire P2_ADD_402_1132_U47 , P2_ADD_402_1132_U48 , P2_ADD_402_1132_U49 , P2_ADD_402_1132_U50 , P2_SUB_563_U6 , P2_SUB_563_U7 , P2_R2182_U4 , P2_R2182_U5 , P2_R2182_U6 , P2_R2182_U7;
wire P2_R2182_U8 , P2_R2182_U9 , P2_R2182_U10 , P2_R2182_U11 , P2_R2182_U12 , P2_R2182_U13 , P2_R2182_U14 , P2_R2182_U15 , P2_R2182_U16 , P2_R2182_U17;
wire P2_R2182_U18 , P2_R2182_U19 , P2_R2182_U20 , P2_R2182_U21 , P2_R2182_U22 , P2_R2182_U23 , P2_R2182_U24 , P2_R2182_U25 , P2_R2182_U26 , P2_R2182_U27;
wire P2_R2182_U28 , P2_R2182_U29 , P2_R2182_U30 , P2_R2182_U31 , P2_R2182_U32 , P2_R2182_U33 , P2_R2182_U34 , P2_R2182_U35 , P2_R2182_U36 , P2_R2182_U37;
wire P2_R2182_U38 , P2_R2182_U39 , P2_R2182_U40 , P2_R2182_U41 , P2_R2182_U42 , P2_R2182_U43 , P2_R2182_U44 , P2_R2182_U45 , P2_R2182_U46 , P2_R2182_U47;
wire P2_R2182_U48 , P2_R2182_U49 , P2_R2182_U50 , P2_R2182_U51 , P2_R2182_U52 , P2_R2182_U53 , P2_R2182_U54 , P2_R2182_U55 , P2_R2182_U56 , P2_R2182_U57;
wire P2_R2182_U58 , P2_R2182_U59 , P2_R2182_U60 , P2_R2182_U61 , P2_R2182_U62 , P2_R2182_U63 , P2_R2182_U64 , P2_R2182_U65 , P2_R2182_U66 , P2_R2182_U67;
wire P2_R2182_U68 , P2_R2182_U69 , P2_R2182_U70 , P2_R2182_U71 , P2_R2182_U72 , P2_R2182_U73 , P2_R2182_U74 , P2_R2182_U75 , P2_R2182_U76 , P2_R2182_U77;
wire P2_R2182_U78 , P2_R2182_U79 , P2_R2182_U80 , P2_R2182_U81 , P2_R2182_U82 , P2_R2182_U83 , P2_R2182_U84 , P2_R2182_U85 , P2_R2182_U86 , P2_R2182_U87;
wire P2_R2182_U88 , P2_R2182_U89 , P2_R2182_U90 , P2_R2182_U91 , P2_R2182_U92 , P2_R2182_U93 , P2_R2182_U94 , P2_R2182_U95 , P2_R2182_U96 , P2_R2182_U97;
wire P2_R2182_U98 , P2_R2182_U99 , P2_R2182_U100 , P2_R2182_U101 , P2_R2182_U102 , P2_R2182_U103 , P2_R2182_U104 , P2_R2182_U105 , P2_R2182_U106 , P2_R2182_U107;
wire P2_R2182_U108 , P2_R2182_U109 , P2_R2182_U110 , P2_R2182_U111 , P2_R2182_U112 , P2_R2182_U113 , P2_R2182_U114 , P2_R2182_U115 , P2_R2182_U116 , P2_R2182_U117;
wire P2_R2182_U118 , P2_R2182_U119 , P2_R2182_U120 , P2_R2182_U121 , P2_R2182_U122 , P2_R2182_U123 , P2_R2182_U124 , P2_R2182_U125 , P2_R2182_U126 , P2_R2182_U127;
wire P2_R2182_U128 , P2_R2182_U129 , P2_R2182_U130 , P2_R2182_U131 , P2_R2182_U132 , P2_R2182_U133 , P2_R2182_U134 , P2_R2182_U135 , P2_R2182_U136 , P2_R2182_U137;
wire P2_R2182_U138 , P2_R2182_U139 , P2_R2182_U140 , P2_R2182_U141 , P2_R2182_U142 , P2_R2182_U143 , P2_R2182_U144 , P2_R2182_U145 , P2_R2182_U146 , P2_R2182_U147;
wire P2_R2182_U148 , P2_R2182_U149 , P2_R2182_U150 , P2_R2182_U151 , P2_R2182_U152 , P2_R2182_U153 , P2_R2182_U154 , P2_R2182_U155 , P2_R2182_U156 , P2_R2182_U157;
wire P2_R2182_U158 , P2_R2182_U159 , P2_R2182_U160 , P2_R2182_U161 , P2_R2182_U162 , P2_R2182_U163 , P2_R2182_U164 , P2_R2182_U165 , P2_R2182_U166 , P2_R2182_U167;
wire P2_R2182_U168 , P2_R2182_U169 , P2_R2182_U170 , P2_R2182_U171 , P2_R2182_U172 , P2_R2182_U173 , P2_R2182_U174 , P2_R2182_U175 , P2_R2182_U176 , P2_R2182_U177;
wire P2_R2182_U178 , P2_R2182_U179 , P2_R2182_U180 , P2_R2182_U181 , P2_R2182_U182 , P2_R2182_U183 , P2_R2182_U184 , P2_R2182_U185 , P2_R2182_U186 , P2_R2182_U187;
wire P2_R2182_U188 , P2_R2182_U189 , P2_R2182_U190 , P2_R2182_U191 , P2_R2182_U192 , P2_R2182_U193 , P2_R2182_U194 , P2_R2182_U195 , P2_R2182_U196 , P2_R2182_U197;
wire P2_R2182_U198 , P2_R2182_U199 , P2_R2182_U200 , P2_R2182_U201 , P2_R2182_U202 , P2_R2182_U203 , P2_R2182_U204 , P2_R2182_U205 , P2_R2182_U206 , P2_R2182_U207;
wire P2_R2182_U208 , P2_R2182_U209 , P2_R2182_U210 , P2_R2182_U211 , P2_R2182_U212 , P2_R2182_U213 , P2_R2182_U214 , P2_R2182_U215 , P2_R2182_U216 , P2_R2182_U217;
wire P2_R2182_U218 , P2_R2182_U219 , P2_R2182_U220 , P2_R2182_U221 , P2_R2182_U222 , P2_R2182_U223 , P2_R2182_U224 , P2_R2182_U225 , P2_R2182_U226 , P2_R2182_U227;
wire P2_R2182_U228 , P2_R2182_U229 , P2_R2182_U230 , P2_R2182_U231 , P2_R2182_U232 , P2_R2182_U233 , P2_R2182_U234 , P2_R2182_U235 , P2_R2182_U236 , P2_R2182_U237;
wire P2_R2182_U238 , P2_R2182_U239 , P2_R2182_U240 , P2_R2182_U241 , P2_R2182_U242 , P2_R2182_U243 , P2_R2182_U244 , P2_R2182_U245 , P2_R2182_U246 , P2_R2182_U247;
wire P2_R2182_U248 , P2_R2182_U249 , P2_R2182_U250 , P2_R2182_U251 , P2_R2182_U252 , P2_R2182_U253 , P2_R2182_U254 , P2_R2182_U255 , P2_R2182_U256 , P2_R2182_U257;
wire P2_R2182_U258 , P2_R2182_U259 , P2_R2182_U260 , P2_R2182_U261 , P2_R2182_U262 , P2_R2182_U263 , P2_R2182_U264 , P2_R2182_U265 , P2_R2182_U266 , P2_R2182_U267;
wire P2_R2182_U268 , P2_R2182_U269 , P2_R2182_U270 , P2_R2182_U271 , P2_R2182_U272 , P2_R2182_U273 , P2_R2182_U274 , P2_R2182_U275 , P2_R2182_U276 , P2_R2182_U277;
wire P2_R2182_U278 , P2_R2182_U279 , P2_R2182_U280 , P2_R2182_U281 , P2_R2182_U282 , P2_R2182_U283 , P2_R2182_U284 , P2_R2182_U285 , P2_R2182_U286 , P2_R2182_U287;
wire P2_R2182_U288 , P2_R2182_U289 , P2_R2182_U290 , P2_R2182_U291 , P2_R2182_U292 , P2_R2182_U293 , P2_R2182_U294 , P2_R2182_U295 , P2_R2182_U296 , P2_R2182_U297;
wire P2_R2182_U298 , P2_R2182_U299 , P2_R2182_U300 , P2_R2182_U301 , P2_R2182_U302 , P2_R2182_U303 , P2_R2182_U304 , P2_R2182_U305 , P2_R2167_U6 , P2_R2167_U7;
wire P2_R2167_U8 , P2_R2167_U9 , P2_R2167_U10 , P2_R2167_U11 , P2_R2167_U12 , P2_R2167_U13 , P2_R2167_U14 , P2_R2167_U15 , P2_R2167_U16 , P2_R2167_U17;
wire P2_R2167_U18 , P2_R2167_U19 , P2_R2167_U20 , P2_R2167_U21 , P2_R2167_U22 , P2_R2167_U23 , P2_R2167_U24 , P2_R2167_U25 , P2_R2167_U26 , P2_R2167_U27;
wire P2_R2167_U28 , P2_R2167_U29 , P2_R2167_U30 , P2_R2167_U31 , P2_R2167_U32 , P2_R2167_U33 , P2_R2167_U34 , P2_R2167_U35 , P2_R2167_U36 , P2_R2167_U37;
wire P2_R2167_U38 , P2_R2167_U39 , P2_R2167_U40 , P2_R2167_U41 , P2_R2167_U42 , P2_R2027_U5 , P2_R2027_U6 , P2_R2027_U7 , P2_R2027_U8 , P2_R2027_U9;
wire P2_R2027_U10 , P2_R2027_U11 , P2_R2027_U12 , P2_R2027_U13 , P2_R2027_U14 , P2_R2027_U15 , P2_R2027_U16 , P2_R2027_U17 , P2_R2027_U18 , P2_R2027_U19;
wire P2_R2027_U20 , P2_R2027_U21 , P2_R2027_U22 , P2_R2027_U23 , P2_R2027_U24 , P2_R2027_U25 , P2_R2027_U26 , P2_R2027_U27 , P2_R2027_U28 , P2_R2027_U29;
wire P2_R2027_U30 , P2_R2027_U31 , P2_R2027_U32 , P2_R2027_U33 , P2_R2027_U34 , P2_R2027_U35 , P2_R2027_U36 , P2_R2027_U37 , P2_R2027_U38 , P2_R2027_U39;
wire P2_R2027_U40 , P2_R2027_U41 , P2_R2027_U42 , P2_R2027_U43 , P2_R2027_U44 , P2_R2027_U45 , P2_R2027_U46 , P2_R2027_U47 , P2_R2027_U48 , P2_R2027_U49;
wire P2_R2027_U50 , P2_R2027_U51 , P2_R2027_U52 , P2_R2027_U53 , P2_R2027_U54 , P2_R2027_U55 , P2_R2027_U56 , P2_R2027_U57 , P2_R2027_U58 , P2_R2027_U59;
wire P2_R2027_U60 , P2_R2027_U61 , P2_R2027_U62 , P2_R2027_U63 , P2_R2027_U64 , P2_R2027_U65 , P2_R2027_U66 , P2_R2027_U67 , P2_R2027_U68 , P2_R2027_U69;
wire P2_R2027_U70 , P2_R2027_U71 , P2_R2027_U72 , P2_R2027_U73 , P2_R2027_U74 , P2_R2027_U75 , P2_R2027_U76 , P2_R2027_U77 , P2_R2027_U78 , P2_R2027_U79;
wire P2_R2027_U80 , P2_R2027_U81 , P2_R2027_U82 , P2_R2027_U83 , P2_R2027_U84 , P2_R2027_U85 , P2_R2027_U86 , P2_R2027_U87 , P2_R2027_U88 , P2_R2027_U89;
wire P2_R2027_U90 , P2_R2027_U91 , P2_R2027_U92 , P2_R2027_U93 , P2_R2027_U94 , P2_R2027_U95 , P2_R2027_U96 , P2_R2027_U97 , P2_R2027_U98 , P2_R2027_U99;
wire P2_R2027_U100 , P2_R2027_U101 , P2_R2027_U102 , P2_R2027_U103 , P2_R2027_U104 , P2_R2027_U105 , P2_R2027_U106 , P2_R2027_U107 , P2_R2027_U108 , P2_R2027_U109;
wire P2_R2027_U110 , P2_R2027_U111 , P2_R2027_U112 , P2_R2027_U113 , P2_R2027_U114 , P2_R2027_U115 , P2_R2027_U116 , P2_R2027_U117 , P2_R2027_U118 , P2_R2027_U119;
wire P2_R2027_U120 , P2_R2027_U121 , P2_R2027_U122 , P2_R2027_U123 , P2_R2027_U124 , P2_R2027_U125 , P2_R2027_U126 , P2_R2027_U127 , P2_R2027_U128 , P2_R2027_U129;
wire P2_R2027_U130 , P2_R2027_U131 , P2_R2027_U132 , P2_R2027_U133 , P2_R2027_U134 , P2_R2027_U135 , P2_R2027_U136 , P2_R2027_U137 , P2_R2027_U138 , P2_R2027_U139;
wire P2_R2027_U140 , P2_R2027_U141 , P2_R2027_U142 , P2_R2027_U143 , P2_R2027_U144 , P2_R2027_U145 , P2_R2027_U146 , P2_R2027_U147 , P2_R2027_U148 , P2_R2027_U149;
wire P2_R2027_U150 , P2_R2027_U151 , P2_R2027_U152 , P2_R2027_U153 , P2_R2027_U154 , P2_R2027_U155 , P2_R2027_U156 , P2_R2027_U157 , P2_R2027_U158 , P2_R2027_U159;
wire P2_R2027_U160 , P2_R2027_U161 , P2_R2027_U162 , P2_R2027_U163 , P2_R2027_U164 , P2_R2027_U165 , P2_R2027_U166 , P2_R2027_U167 , P2_R2027_U168 , P2_R2027_U169;
wire P2_R2027_U170 , P2_R2027_U171 , P2_R2027_U172 , P2_R2027_U173 , P2_R2027_U174 , P2_R2027_U175 , P2_R2027_U176 , P2_R2027_U177 , P2_R2027_U178 , P2_R2027_U179;
wire P2_R2027_U180 , P2_R2027_U181 , P2_R2027_U182 , P2_R2027_U183 , P2_R2027_U184 , P2_R2027_U185 , P2_R2027_U186 , P2_R2027_U187 , P2_R2027_U188 , P2_R2027_U189;
wire P2_LT_563_1260_U6 , P2_LT_563_1260_U7 , P2_R2337_U4 , P2_R2337_U5 , P2_R2337_U6 , P2_R2337_U7 , P2_R2337_U8 , P2_R2337_U9 , P2_R2337_U10 , P2_R2337_U11;
wire P2_R2337_U12 , P2_R2337_U13 , P2_R2337_U14 , P2_R2337_U15 , P2_R2337_U16 , P2_R2337_U17 , P2_R2337_U18 , P2_R2337_U19 , P2_R2337_U20 , P2_R2337_U21;
wire P2_R2337_U22 , P2_R2337_U23 , P2_R2337_U24 , P2_R2337_U25 , P2_R2337_U26 , P2_R2337_U27 , P2_R2337_U28 , P2_R2337_U29 , P2_R2337_U30 , P2_R2337_U31;
wire P2_R2337_U32 , P2_R2337_U33 , P2_R2337_U34 , P2_R2337_U35 , P2_R2337_U36 , P2_R2337_U37 , P2_R2337_U38 , P2_R2337_U39 , P2_R2337_U40 , P2_R2337_U41;
wire P2_R2337_U42 , P2_R2337_U43 , P2_R2337_U44 , P2_R2337_U45 , P2_R2337_U46 , P2_R2337_U47 , P2_R2337_U48 , P2_R2337_U49 , P2_R2337_U50 , P2_R2337_U51;
wire P2_R2337_U52 , P2_R2337_U53 , P2_R2337_U54 , P2_R2337_U55 , P2_R2337_U56 , P2_R2337_U57 , P2_R2337_U58 , P2_R2337_U59 , P2_R2337_U60 , P2_R2337_U61;
wire P2_R2337_U62 , P2_R2337_U63 , P2_R2337_U64 , P2_R2337_U65 , P2_R2337_U66 , P2_R2337_U67 , P2_R2337_U68 , P2_R2337_U69 , P2_R2337_U70 , P2_R2337_U71;
wire P2_R2337_U72 , P2_R2337_U73 , P2_R2337_U74 , P2_R2337_U75 , P2_R2337_U76 , P2_R2337_U77 , P2_R2337_U78 , P2_R2337_U79 , P2_R2337_U80 , P2_R2337_U81;
wire P2_R2337_U82 , P2_R2337_U83 , P2_R2337_U84 , P2_R2337_U85 , P2_R2337_U86 , P2_R2337_U87 , P2_R2337_U88 , P2_R2337_U89 , P2_R2337_U90 , P2_R2337_U91;
wire P2_R2337_U92 , P2_R2337_U93 , P2_R2337_U94 , P2_R2337_U95 , P2_R2337_U96 , P2_R2337_U97 , P2_R2337_U98 , P2_R2337_U99 , P2_R2337_U100 , P2_R2337_U101;
wire P2_R2337_U102 , P2_R2337_U103 , P2_R2337_U104 , P2_R2337_U105 , P2_R2337_U106 , P2_R2337_U107 , P2_R2337_U108 , P2_R2337_U109 , P2_R2337_U110 , P2_R2337_U111;
wire P2_R2337_U112 , P2_R2337_U113 , P2_R2337_U114 , P2_R2337_U115 , P2_R2337_U116 , P2_R2337_U117 , P2_R2337_U118 , P2_R2337_U119 , P2_R2337_U120 , P2_R2337_U121;
wire P2_R2337_U122 , P2_R2337_U123 , P2_R2337_U124 , P2_R2337_U125 , P2_R2337_U126 , P2_R2337_U127 , P2_R2337_U128 , P2_R2337_U129 , P2_R2337_U130 , P2_R2337_U131;
wire P2_R2337_U132 , P2_R2337_U133 , P2_R2337_U134 , P2_R2337_U135 , P2_R2337_U136 , P2_R2337_U137 , P2_R2337_U138 , P2_R2337_U139 , P2_R2337_U140 , P2_R2337_U141;
wire P2_R2337_U142 , P2_R2337_U143 , P2_R2337_U144 , P2_R2337_U145 , P2_R2337_U146 , P2_R2337_U147 , P2_R2337_U148 , P2_R2337_U149 , P2_R2337_U150 , P2_R2337_U151;
wire P2_R2337_U152 , P2_R2337_U153 , P2_R2337_U154 , P2_R2337_U155 , P2_R2337_U156 , P2_R2337_U157 , P2_R2337_U158 , P2_R2337_U159 , P2_R2337_U160 , P2_R2337_U161;
wire P2_R2337_U162 , P2_R2337_U163 , P2_R2337_U164 , P2_R2337_U165 , P2_R2337_U166 , P2_R2337_U167 , P2_R2337_U168 , P2_R2337_U169 , P2_R2337_U170 , P2_R2337_U171;
wire P2_R2337_U172 , P2_R2337_U173 , P2_R2337_U174 , P2_R2337_U175 , P2_R2337_U176 , P2_R2337_U177 , P2_R2337_U178 , P2_R2337_U179 , P2_R2337_U180 , P2_R2337_U181;
wire P2_R2337_U182 , P2_R2147_U4 , P2_R2147_U5 , P2_R2147_U6 , P2_R2147_U7 , P2_R2147_U8 , P2_R2147_U9 , P2_R2147_U10 , P2_R2147_U11 , P2_R2147_U12;
wire P2_R2147_U13 , P2_R2147_U14 , P2_R2147_U15 , P2_R2147_U16 , P2_R2147_U17 , P2_R2147_U18 , P2_R2147_U19 , P2_R2147_U20 , P2_R2219_U6 , P2_R2219_U7;
wire P2_R2219_U8 , P2_R2219_U9 , P2_R2219_U10 , P2_R2219_U11 , P2_R2219_U12 , P2_R2219_U13 , P2_R2219_U14 , P2_R2219_U15 , P2_R2219_U16 , P2_R2219_U17;
wire P2_R2219_U18 , P2_R2219_U19 , P2_R2219_U20 , P2_R2219_U21 , P2_R2219_U22 , P2_R2219_U23 , P2_R2219_U24 , P2_R2219_U25 , P2_R2219_U26 , P2_R2219_U27;
wire P2_R2219_U28 , P2_R2219_U29 , P2_R2219_U30 , P2_R2219_U31 , P2_R2219_U32 , P2_R2219_U33 , P2_R2219_U34 , P2_R2219_U35 , P2_R2219_U36 , P2_R2219_U37;
wire P2_R2219_U38 , P2_R2219_U39 , P2_R2219_U40 , P2_R2219_U41 , P2_R2219_U42 , P2_R2219_U43 , P2_R2219_U44 , P2_R2219_U45 , P2_R2219_U46 , P2_R2219_U47;
wire P2_R2219_U48 , P2_R2219_U49 , P2_R2219_U50 , P2_R2219_U51 , P2_R2219_U52 , P2_R2219_U53 , P2_R2219_U54 , P2_R2219_U55 , P2_R2219_U56 , P2_R2219_U57;
wire P2_R2219_U58 , P2_R2219_U59 , P2_R2219_U60 , P2_R2219_U61 , P2_R2219_U62 , P2_R2219_U63 , P2_R2219_U64 , P2_R2219_U65 , P2_R2219_U66 , P2_R2219_U67;
wire P2_R2219_U68 , P2_R2219_U69 , P2_R2219_U70 , P2_R2219_U71 , P2_R2219_U72 , P2_R2219_U73 , P2_R2219_U74 , P2_R2219_U75 , P2_R2219_U76 , P2_R2219_U77;
wire P2_R2219_U78 , P2_R2219_U79 , P2_R2219_U80 , P2_R2219_U81 , P2_R2219_U82 , P2_R2219_U83 , P2_R2219_U84 , P2_R2219_U85 , P2_R2219_U86 , P2_R2219_U87;
wire P2_R2219_U88 , P2_R2219_U89 , P2_R2219_U90 , P2_R2219_U91 , P2_R2219_U92 , P2_R2219_U93 , P2_R2219_U94 , P2_R2219_U95 , P2_R2219_U96 , P2_R2219_U97;
wire P2_R2219_U98 , P2_R2219_U99 , P2_R2219_U100 , P2_R2219_U101 , P2_R2219_U102 , P2_R2219_U103 , P2_R2219_U104 , P2_R2219_U105 , P2_R2219_U106 , P2_R2219_U107;
wire P2_R2219_U108 , P2_R2219_U109 , P2_R2219_U110 , P2_R2219_U111 , P2_R2219_U112 , P2_R2219_U113 , P2_R2219_U114 , P2_R2219_U115 , P2_R2219_U116 , P2_R2243_U6;
wire P2_R2243_U7 , P2_R2243_U8 , P2_R2243_U9 , P2_R2243_U10 , P2_R2243_U11 , P2_SUB_589_U6 , P2_SUB_589_U7 , P2_SUB_589_U8 , P2_SUB_589_U9 , P2_R2096_U4;
wire P2_R2096_U5 , P2_R2096_U6 , P2_R2096_U7 , P2_R2096_U8 , P2_R2096_U9 , P2_R2096_U10 , P2_R2096_U11 , P2_R2096_U12 , P2_R2096_U13 , P2_R2096_U14;
wire P2_R2096_U15 , P2_R2096_U16 , P2_R2096_U17 , P2_R2096_U18 , P2_R2096_U19 , P2_R2096_U20 , P2_R2096_U21 , P2_R2096_U22 , P2_R2096_U23 , P2_R2096_U24;
wire P2_R2096_U25 , P2_R2096_U26 , P2_R2096_U27 , P2_R2096_U28 , P2_R2096_U29 , P2_R2096_U30 , P2_R2096_U31 , P2_R2096_U32 , P2_R2096_U33 , P2_R2096_U34;
wire P2_R2096_U35 , P2_R2096_U36 , P2_R2096_U37 , P2_R2096_U38 , P2_R2096_U39 , P2_R2096_U40 , P2_R2096_U41 , P2_R2096_U42 , P2_R2096_U43 , P2_R2096_U44;
wire P2_R2096_U45 , P2_R2096_U46 , P2_R2096_U47 , P2_R2096_U48 , P2_R2096_U49 , P2_R2096_U50 , P2_R2096_U51 , P2_R2096_U52 , P2_R2096_U53 , P2_R2096_U54;
wire P2_R2096_U55 , P2_R2096_U56 , P2_R2096_U57 , P2_R2096_U58 , P2_R2096_U59 , P2_R2096_U60 , P2_R2096_U61 , P2_R2096_U62 , P2_R2096_U63 , P2_R2096_U64;
wire P2_R2096_U65 , P2_R2096_U66 , P2_R2096_U67 , P2_R2096_U68 , P2_R2096_U69 , P2_R2096_U70 , P2_R2096_U71 , P2_R2096_U72 , P2_R2096_U73 , P2_R2096_U74;
wire P2_R2096_U75 , P2_R2096_U76 , P2_R2096_U77 , P2_R2096_U78 , P2_R2096_U79 , P2_R2096_U80 , P2_R2096_U81 , P2_R2096_U82 , P2_R2096_U83 , P2_R2096_U84;
wire P2_R2096_U85 , P2_R2096_U86 , P2_R2096_U87 , P2_R2096_U88 , P2_R2096_U89 , P2_R2096_U90 , P2_R2096_U91 , P2_R2096_U92 , P2_R2096_U93 , P2_R2096_U94;
wire P2_R2096_U95 , P2_R2096_U96 , P2_R2096_U97 , P2_R2096_U98 , P2_R2096_U99 , P2_R2096_U100 , P2_R2096_U101 , P2_R2096_U102 , P2_R2096_U103 , P2_R2096_U104;
wire P2_R2096_U105 , P2_R2096_U106 , P2_R2096_U107 , P2_R2096_U108 , P2_R2096_U109 , P2_R2096_U110 , P2_R2096_U111 , P2_R2096_U112 , P2_R2096_U113 , P2_R2096_U114;
wire P2_R2096_U115 , P2_R2096_U116 , P2_R2096_U117 , P2_R2096_U118 , P2_R2096_U119 , P2_R2096_U120 , P2_R2096_U121 , P2_R2096_U122 , P2_R2096_U123 , P2_R2096_U124;
wire P2_R2096_U125 , P2_R2096_U126 , P2_R2096_U127 , P2_R2096_U128 , P2_R2096_U129 , P2_R2096_U130 , P2_R2096_U131 , P2_R2096_U132 , P2_R2096_U133 , P2_R2096_U134;
wire P2_R2096_U135 , P2_R2096_U136 , P2_R2096_U137 , P2_R2096_U138 , P2_R2096_U139 , P2_R2096_U140 , P2_R2096_U141 , P2_R2096_U142 , P2_R2096_U143 , P2_R2096_U144;
wire P2_R2096_U145 , P2_R2096_U146 , P2_R2096_U147 , P2_R2096_U148 , P2_R2096_U149 , P2_R2096_U150 , P2_R2096_U151 , P2_R2096_U152 , P2_R2096_U153 , P2_R2096_U154;
wire P2_R2096_U155 , P2_R2096_U156 , P2_R2096_U157 , P2_R2096_U158 , P2_R2096_U159 , P2_R2096_U160 , P2_R2096_U161 , P2_R2096_U162 , P2_R2096_U163 , P2_R2096_U164;
wire P2_R2096_U165 , P2_R2096_U166 , P2_R2096_U167 , P2_R2096_U168 , P2_R2096_U169 , P2_R2096_U170 , P2_R2096_U171 , P2_R2096_U172 , P2_R2096_U173 , P2_R2096_U174;
wire P2_R2096_U175 , P2_R2096_U176 , P2_R2096_U177 , P2_R2096_U178 , P2_R2096_U179 , P2_R2096_U180 , P2_R2096_U181 , P2_R2096_U182 , P2_R2096_U183 , P2_R2096_U184;
wire P2_R2096_U185 , P2_R2096_U186 , P2_R2096_U187 , P2_R2096_U188 , P2_R2096_U189 , P2_R2096_U190 , P2_R2096_U191 , P2_R2096_U192 , P2_R2096_U193 , P2_R2096_U194;
wire P2_R2096_U195 , P2_R2096_U196 , P2_R2096_U197 , P2_R2096_U198 , P2_R2096_U199 , P2_R2096_U200 , P2_R2096_U201 , P2_R2096_U202 , P2_R2096_U203 , P2_R2096_U204;
wire P2_R2096_U205 , P2_R2096_U206 , P2_R2096_U207 , P2_R2096_U208 , P2_R2096_U209 , P2_R2096_U210 , P2_R2096_U211 , P2_R2096_U212 , P2_R2096_U213 , P2_R2096_U214;
wire P2_R2096_U215 , P2_R2096_U216 , P2_R2096_U217 , P2_R2096_U218 , P2_R2096_U219 , P2_R2096_U220 , P2_R2096_U221 , P2_R2096_U222 , P2_R2096_U223 , P2_R2096_U224;
wire P2_R2096_U225 , P2_R2096_U226 , P2_R2096_U227 , P2_R2096_U228 , P2_R2096_U229 , P2_R2096_U230 , P2_R2096_U231 , P2_R2096_U232 , P2_R2096_U233 , P2_R2096_U234;
wire P2_R2096_U235 , P2_R2096_U236 , P2_R2096_U237 , P2_R2096_U238 , P2_R2096_U239 , P2_R2096_U240 , P2_R2096_U241 , P2_R2096_U242 , P2_R2096_U243 , P2_R2096_U244;
wire P2_R2096_U245 , P2_R2096_U246 , P2_R2096_U247 , P2_R2096_U248 , P2_R2096_U249 , P2_R2096_U250 , P2_R2096_U251 , P2_R2096_U252 , P2_R2096_U253 , P2_R2096_U254;
wire P2_R2096_U255 , P2_R2096_U256 , P2_R2096_U257 , P2_R2096_U258 , P2_R2096_U259 , P2_R2096_U260 , P2_R2096_U261 , P2_R2096_U262 , P2_R2096_U263 , P2_R2096_U264;
wire P2_R2096_U265 , P2_GTE_370_U6 , P2_GTE_370_U7 , P2_GTE_370_U8 , P2_GTE_370_U9 , P2_LT_563_U6 , P2_LT_563_U7 , P2_LT_563_U8 , P2_LT_563_U9 , P2_LT_563_U10;
wire P2_LT_563_U11 , P2_LT_563_U12 , P2_LT_563_U13 , P2_LT_563_U14 , P2_LT_563_U15 , P2_LT_563_U16 , P2_LT_563_U17 , P2_LT_563_U18 , P2_LT_563_U19 , P2_LT_563_U20;
wire P2_LT_563_U21 , P2_LT_563_U22 , P2_LT_563_U23 , P2_LT_563_U24 , P2_LT_563_U25 , P2_LT_563_U26 , P2_LT_563_U27 , P2_R2256_U4 , P2_R2256_U5 , P2_R2256_U6;
wire P2_R2256_U7 , P2_R2256_U8 , P2_R2256_U9 , P2_R2256_U10 , P2_R2256_U11 , P2_R2256_U12 , P2_R2256_U13 , P2_R2256_U14 , P2_R2256_U15 , P2_R2256_U16;
wire P2_R2256_U17 , P2_R2256_U18 , P2_R2256_U19 , P2_R2256_U20 , P2_R2256_U21 , P2_R2256_U22 , P2_R2256_U23 , P2_R2256_U24 , P2_R2256_U25 , P2_R2256_U26;
wire P2_R2256_U27 , P2_R2256_U28 , P2_R2256_U29 , P2_R2256_U30 , P2_R2256_U31 , P2_R2256_U32 , P2_R2256_U33 , P2_R2256_U34 , P2_R2256_U35 , P2_R2256_U36;
wire P2_R2256_U37 , P2_R2256_U38 , P2_R2256_U39 , P2_R2256_U40 , P2_R2256_U41 , P2_R2256_U42 , P2_R2256_U43 , P2_R2256_U44 , P2_R2256_U45 , P2_R2256_U46;
wire P2_R2256_U47 , P2_R2256_U48 , P2_R2256_U49 , P2_R2256_U50 , P2_R2256_U51 , P2_R2256_U52 , P2_R2256_U53 , P2_R2256_U54 , P2_R2256_U55 , P2_R2256_U56;
wire P2_R2256_U57 , P2_R2256_U58 , P2_R2256_U59 , P2_R2256_U60 , P2_R2256_U61 , P2_R2256_U62 , P2_R2256_U63 , P2_R2256_U64 , P2_R2256_U65 , P2_R2256_U66;
wire P2_R2256_U67 , P2_R2256_U68 , P2_R2256_U69 , P2_R2256_U70 , P2_R2238_U6 , P2_R2238_U7 , P2_R2238_U8 , P2_R2238_U9 , P2_R2238_U10 , P2_R2238_U11;
wire P2_R2238_U12 , P2_R2238_U13 , P2_R2238_U14 , P2_R2238_U15 , P2_R2238_U16 , P2_R2238_U17 , P2_R2238_U18 , P2_R2238_U19 , P2_R2238_U20 , P2_R2238_U21;
wire P2_R2238_U22 , P2_R2238_U23 , P2_R2238_U24 , P2_R2238_U25 , P2_R2238_U26 , P2_R2238_U27 , P2_R2238_U28 , P2_R2238_U29 , P2_R2238_U30 , P2_R2238_U31;
wire P2_R2238_U32 , P2_R2238_U33 , P2_R2238_U34 , P2_R2238_U35 , P2_R2238_U36 , P2_R2238_U37 , P2_R2238_U38 , P2_R2238_U39 , P2_R2238_U40 , P2_R2238_U41;
wire P2_R2238_U42 , P2_R2238_U43 , P2_R2238_U44 , P2_R2238_U45 , P2_R2238_U46 , P2_R2238_U47 , P2_R2238_U48 , P2_R2238_U49 , P2_R2238_U50 , P2_R2238_U51;
wire P2_R2238_U52 , P2_R2238_U53 , P2_R2238_U54 , P2_R2238_U55 , P2_R2238_U56 , P2_R2238_U57 , P2_R2238_U58 , P2_R2238_U59 , P2_R2238_U60 , P2_R2238_U61;
wire P2_R2238_U62 , P2_R2238_U63 , P2_R2238_U64 , P2_R2238_U65 , P2_R2238_U66 , P2_R1957_U6 , P2_R1957_U7 , P2_R1957_U8 , P2_R1957_U9 , P2_R1957_U10;
wire P2_R1957_U11 , P2_R1957_U12 , P2_R1957_U13 , P2_R1957_U14 , P2_R1957_U15 , P2_R1957_U16 , P2_R1957_U17 , P2_R1957_U18 , P2_R1957_U19 , P2_R1957_U20;
wire P2_R1957_U21 , P2_R1957_U22 , P2_R1957_U23 , P2_R1957_U24 , P2_R1957_U25 , P2_R1957_U26 , P2_R1957_U27 , P2_R1957_U28 , P2_R1957_U29 , P2_R1957_U30;
wire P2_R1957_U31 , P2_R1957_U32 , P2_R1957_U33 , P2_R1957_U34 , P2_R1957_U35 , P2_R1957_U36 , P2_R1957_U37 , P2_R1957_U38 , P2_R1957_U39 , P2_R1957_U40;
wire P2_R1957_U41 , P2_R1957_U42 , P2_R1957_U43 , P2_R1957_U44 , P2_R1957_U45 , P2_R1957_U46 , P2_R1957_U47 , P2_R1957_U48 , P2_R1957_U49 , P2_R1957_U50;
wire P2_R1957_U51 , P2_R1957_U52 , P2_R1957_U53 , P2_R1957_U54 , P2_R1957_U55 , P2_R1957_U56 , P2_R1957_U57 , P2_R1957_U58 , P2_R1957_U59 , P2_R1957_U60;
wire P2_R1957_U61 , P2_R1957_U62 , P2_R1957_U63 , P2_R1957_U64 , P2_R1957_U65 , P2_R1957_U66 , P2_R1957_U67 , P2_R1957_U68 , P2_R1957_U69 , P2_R1957_U70;
wire P2_R1957_U71 , P2_R1957_U72 , P2_R1957_U73 , P2_R1957_U74 , P2_R1957_U75 , P2_R1957_U76 , P2_R1957_U77 , P2_R1957_U78 , P2_R1957_U79 , P2_R1957_U80;
wire P2_R1957_U81 , P2_R1957_U82 , P2_R1957_U83 , P2_R1957_U84 , P2_R1957_U85 , P2_R1957_U86 , P2_R1957_U87 , P2_R1957_U88 , P2_R1957_U89 , P2_R1957_U90;
wire P2_R1957_U91 , P2_R1957_U92 , P2_R1957_U93 , P2_R1957_U94 , P2_R1957_U95 , P2_R1957_U96 , P2_R1957_U97 , P2_R1957_U98 , P2_R1957_U99 , P2_R1957_U100;
wire P2_R1957_U101 , P2_R1957_U102 , P2_R1957_U103 , P2_R1957_U104 , P2_R1957_U105 , P2_R1957_U106 , P2_R1957_U107 , P2_R1957_U108 , P2_R1957_U109 , P2_R1957_U110;
wire P2_R1957_U111 , P2_R1957_U112 , P2_R1957_U113 , P2_R1957_U114 , P2_R1957_U115 , P2_R1957_U116 , P2_R1957_U117 , P2_R1957_U118 , P2_R1957_U119 , P2_R1957_U120;
wire P2_R1957_U121 , P2_R1957_U122 , P2_R1957_U123 , P2_R1957_U124 , P2_R1957_U125 , P2_R1957_U126 , P2_R1957_U127 , P2_R1957_U128 , P2_R1957_U129 , P2_R1957_U130;
wire P2_R1957_U131 , P2_R1957_U132 , P2_R1957_U133 , P2_R1957_U134 , P2_R1957_U135 , P2_R1957_U136 , P2_R1957_U137 , P2_R1957_U138 , P2_R1957_U139 , P2_R1957_U140;
wire P2_R1957_U141 , P2_R1957_U142 , P2_R1957_U143 , P2_R1957_U144 , P2_R1957_U145 , P2_R1957_U146 , P2_R1957_U147 , P2_R1957_U148 , P2_R1957_U149 , P2_R1957_U150;
wire P2_R1957_U151 , P2_R1957_U152 , P2_R1957_U153 , P2_R1957_U154 , P2_R1957_U155 , P2_R1957_U156 , P2_R1957_U157 , P2_R1957_U158 , P2_R1957_U159 , P2_R2278_U4;
wire P2_R2278_U5 , P2_R2278_U6 , P2_R2278_U7 , P2_R2278_U8 , P2_R2278_U9 , P2_R2278_U10 , P2_R2278_U11 , P2_R2278_U12 , P2_R2278_U13 , P2_R2278_U14;
wire P2_R2278_U15 , P2_R2278_U16 , P2_R2278_U17 , P2_R2278_U18 , P2_R2278_U19 , P2_R2278_U20 , P2_R2278_U21 , P2_R2278_U22 , P2_R2278_U23 , P2_R2278_U24;
wire P2_R2278_U25 , P2_R2278_U26 , P2_R2278_U27 , P2_R2278_U28 , P2_R2278_U29 , P2_R2278_U30 , P2_R2278_U31 , P2_R2278_U32 , P2_R2278_U33 , P2_R2278_U34;
wire P2_R2278_U35 , P2_R2278_U36 , P2_R2278_U37 , P2_R2278_U38 , P2_R2278_U39 , P2_R2278_U40 , P2_R2278_U41 , P2_R2278_U42 , P2_R2278_U43 , P2_R2278_U44;
wire P2_R2278_U45 , P2_R2278_U46 , P2_R2278_U47 , P2_R2278_U48 , P2_R2278_U49 , P2_R2278_U50 , P2_R2278_U51 , P2_R2278_U52 , P2_R2278_U53 , P2_R2278_U54;
wire P2_R2278_U55 , P2_R2278_U56 , P2_R2278_U57 , P2_R2278_U58 , P2_R2278_U59 , P2_R2278_U60 , P2_R2278_U61 , P2_R2278_U62 , P2_R2278_U63 , P2_R2278_U64;
wire P2_R2278_U65 , P2_R2278_U66 , P2_R2278_U67 , P2_R2278_U68 , P2_R2278_U69 , P2_R2278_U70 , P2_R2278_U71 , P2_R2278_U72 , P2_R2278_U73 , P2_R2278_U74;
wire P2_R2278_U75 , P2_R2278_U76 , P2_R2278_U77 , P2_R2278_U78 , P2_R2278_U79 , P2_R2278_U80 , P2_R2278_U81 , P2_R2278_U82 , P2_R2278_U83 , P2_R2278_U84;
wire P2_R2278_U85 , P2_R2278_U86 , P2_R2278_U87 , P2_R2278_U88 , P2_R2278_U89 , P2_R2278_U90 , P2_R2278_U91 , P2_R2278_U92 , P2_R2278_U93 , P2_R2278_U94;
wire P2_R2278_U95 , P2_R2278_U96 , P2_R2278_U97 , P2_R2278_U98 , P2_R2278_U99 , P2_R2278_U100 , P2_R2278_U101 , P2_R2278_U102 , P2_R2278_U103 , P2_R2278_U104;
wire P2_R2278_U105 , P2_R2278_U106 , P2_R2278_U107 , P2_R2278_U108 , P2_R2278_U109 , P2_R2278_U110 , P2_R2278_U111 , P2_R2278_U112 , P2_R2278_U113 , P2_R2278_U114;
wire P2_R2278_U115 , P2_R2278_U116 , P2_R2278_U117 , P2_R2278_U118 , P2_R2278_U119 , P2_R2278_U120 , P2_R2278_U121 , P2_R2278_U122 , P2_R2278_U123 , P2_R2278_U124;
wire P2_R2278_U125 , P2_R2278_U126 , P2_R2278_U127 , P2_R2278_U128 , P2_R2278_U129 , P2_R2278_U130 , P2_R2278_U131 , P2_R2278_U132 , P2_R2278_U133 , P2_R2278_U134;
wire P2_R2278_U135 , P2_R2278_U136 , P2_R2278_U137 , P2_R2278_U138 , P2_R2278_U139 , P2_R2278_U140 , P2_R2278_U141 , P2_R2278_U142 , P2_R2278_U143 , P2_R2278_U144;
wire P2_R2278_U145 , P2_R2278_U146 , P2_R2278_U147 , P2_R2278_U148 , P2_R2278_U149 , P2_R2278_U150 , P2_R2278_U151 , P2_R2278_U152 , P2_R2278_U153 , P2_R2278_U154;
wire P2_R2278_U155 , P2_R2278_U156 , P2_R2278_U157 , P2_R2278_U158 , P2_R2278_U159 , P2_R2278_U160 , P2_R2278_U161 , P2_R2278_U162 , P2_R2278_U163 , P2_R2278_U164;
wire P2_R2278_U165 , P2_R2278_U166 , P2_R2278_U167 , P2_R2278_U168 , P2_R2278_U169 , P2_R2278_U170 , P2_R2278_U171 , P2_R2278_U172 , P2_R2278_U173 , P2_R2278_U174;
wire P2_R2278_U175 , P2_R2278_U176 , P2_R2278_U177 , P2_R2278_U178 , P2_R2278_U179 , P2_R2278_U180 , P2_R2278_U181 , P2_R2278_U182 , P2_R2278_U183 , P2_R2278_U184;
wire P2_R2278_U185 , P2_R2278_U186 , P2_R2278_U187 , P2_R2278_U188 , P2_R2278_U189 , P2_R2278_U190 , P2_R2278_U191 , P2_R2278_U192 , P2_R2278_U193 , P2_R2278_U194;
wire P2_R2278_U195 , P2_R2278_U196 , P2_R2278_U197 , P2_R2278_U198 , P2_R2278_U199 , P2_R2278_U200 , P2_R2278_U201 , P2_R2278_U202 , P2_R2278_U203 , P2_R2278_U204;
wire P2_R2278_U205 , P2_R2278_U206 , P2_R2278_U207 , P2_R2278_U208 , P2_R2278_U209 , P2_R2278_U210 , P2_R2278_U211 , P2_R2278_U212 , P2_R2278_U213 , P2_R2278_U214;
wire P2_R2278_U215 , P2_R2278_U216 , P2_R2278_U217 , P2_R2278_U218 , P2_R2278_U219 , P2_R2278_U220 , P2_R2278_U221 , P2_R2278_U222 , P2_R2278_U223 , P2_R2278_U224;
wire P2_R2278_U225 , P2_R2278_U226 , P2_R2278_U227 , P2_R2278_U228 , P2_R2278_U229 , P2_R2278_U230 , P2_R2278_U231 , P2_R2278_U232 , P2_R2278_U233 , P2_R2278_U234;
wire P2_R2278_U235 , P2_R2278_U236 , P2_R2278_U237 , P2_R2278_U238 , P2_R2278_U239 , P2_R2278_U240 , P2_R2278_U241 , P2_R2278_U242 , P2_R2278_U243 , P2_R2278_U244;
wire P2_R2278_U245 , P2_R2278_U246 , P2_R2278_U247 , P2_R2278_U248 , P2_R2278_U249 , P2_R2278_U250 , P2_R2278_U251 , P2_R2278_U252 , P2_R2278_U253 , P2_R2278_U254;
wire P2_R2278_U255 , P2_R2278_U256 , P2_R2278_U257 , P2_R2278_U258 , P2_R2278_U259 , P2_R2278_U260 , P2_R2278_U261 , P2_R2278_U262 , P2_R2278_U263 , P2_R2278_U264;
wire P2_R2278_U265 , P2_R2278_U266 , P2_R2278_U267 , P2_R2278_U268 , P2_R2278_U269 , P2_R2278_U270 , P2_R2278_U271 , P2_R2278_U272 , P2_R2278_U273 , P2_R2278_U274;
wire P2_R2278_U275 , P2_R2278_U276 , P2_R2278_U277 , P2_R2278_U278 , P2_R2278_U279 , P2_R2278_U280 , P2_R2278_U281 , P2_R2278_U282 , P2_R2278_U283 , P2_R2278_U284;
wire P2_R2278_U285 , P2_R2278_U286 , P2_R2278_U287 , P2_R2278_U288 , P2_R2278_U289 , P2_R2278_U290 , P2_R2278_U291 , P2_R2278_U292 , P2_R2278_U293 , P2_R2278_U294;
wire P2_R2278_U295 , P2_R2278_U296 , P2_R2278_U297 , P2_R2278_U298 , P2_R2278_U299 , P2_R2278_U300 , P2_R2278_U301 , P2_R2278_U302 , P2_R2278_U303 , P2_R2278_U304;
wire P2_R2278_U305 , P2_R2278_U306 , P2_R2278_U307 , P2_R2278_U308 , P2_R2278_U309 , P2_R2278_U310 , P2_R2278_U311 , P2_R2278_U312 , P2_R2278_U313 , P2_R2278_U314;
wire P2_R2278_U315 , P2_R2278_U316 , P2_R2278_U317 , P2_R2278_U318 , P2_R2278_U319 , P2_R2278_U320 , P2_R2278_U321 , P2_R2278_U322 , P2_R2278_U323 , P2_R2278_U324;
wire P2_R2278_U325 , P2_R2278_U326 , P2_R2278_U327 , P2_R2278_U328 , P2_R2278_U329 , P2_R2278_U330 , P2_R2278_U331 , P2_R2278_U332 , P2_R2278_U333 , P2_R2278_U334;
wire P2_R2278_U335 , P2_R2278_U336 , P2_R2278_U337 , P2_R2278_U338 , P2_R2278_U339 , P2_R2278_U340 , P2_R2278_U341 , P2_R2278_U342 , P2_R2278_U343 , P2_R2278_U344;
wire P2_R2278_U345 , P2_R2278_U346 , P2_R2278_U347 , P2_R2278_U348 , P2_R2278_U349 , P2_R2278_U350 , P2_R2278_U351 , P2_R2278_U352 , P2_R2278_U353 , P2_R2278_U354;
wire P2_R2278_U355 , P2_R2278_U356 , P2_R2278_U357 , P2_R2278_U358 , P2_R2278_U359 , P2_R2278_U360 , P2_R2278_U361 , P2_R2278_U362 , P2_R2278_U363 , P2_R2278_U364;
wire P2_R2278_U365 , P2_R2278_U366 , P2_R2278_U367 , P2_R2278_U368 , P2_R2278_U369 , P2_R2278_U370 , P2_R2278_U371 , P2_R2278_U372 , P2_R2278_U373 , P2_R2278_U374;
wire P2_R2278_U375 , P2_R2278_U376 , P2_R2278_U377 , P2_R2278_U378 , P2_R2278_U379 , P2_R2278_U380 , P2_R2278_U381 , P2_R2278_U382 , P2_R2278_U383 , P2_R2278_U384;
wire P2_R2278_U385 , P2_R2278_U386 , P2_R2278_U387 , P2_R2278_U388 , P2_R2278_U389 , P2_R2278_U390 , P2_R2278_U391 , P2_R2278_U392 , P2_R2278_U393 , P2_R2278_U394;
wire P2_R2278_U395 , P2_R2278_U396 , P2_R2278_U397 , P2_R2278_U398 , P2_R2278_U399 , P2_R2278_U400 , P2_R2278_U401 , P2_R2278_U402 , P2_R2278_U403 , P2_R2278_U404;
wire P2_R2278_U405 , P2_R2278_U406 , P2_R2278_U407 , P2_R2278_U408 , P2_R2278_U409 , P2_R2278_U410 , P2_R2278_U411 , P2_R2278_U412 , P2_R2278_U413 , P2_R2278_U414;
wire P2_R2278_U415 , P2_R2278_U416 , P2_R2278_U417 , P2_R2278_U418 , P2_R2278_U419 , P2_R2278_U420 , P2_R2278_U421 , P2_R2278_U422 , P2_R2278_U423 , P2_R2278_U424;
wire P2_R2278_U425 , P2_R2278_U426 , P2_R2278_U427 , P2_R2278_U428 , P2_R2278_U429 , P2_R2278_U430 , P2_R2278_U431 , P2_R2278_U432 , P2_R2278_U433 , P2_R2278_U434;
wire P2_R2278_U435 , P2_R2278_U436 , P2_R2278_U437 , P2_R2278_U438 , P2_R2278_U439 , P2_R2278_U440 , P2_R2278_U441 , P2_R2278_U442 , P2_R2278_U443 , P2_R2278_U444;
wire P2_R2278_U445 , P2_R2278_U446 , P2_R2278_U447 , P2_R2278_U448 , P2_R2278_U449 , P2_R2278_U450 , P2_R2278_U451 , P2_R2278_U452 , P2_R2278_U453 , P2_R2278_U454;
wire P2_R2278_U455 , P2_R2278_U456 , P2_R2278_U457 , P2_R2278_U458 , P2_R2278_U459 , P2_R2278_U460 , P2_R2278_U461 , P2_R2278_U462 , P2_R2278_U463 , P2_R2278_U464;
wire P2_R2278_U465 , P2_R2278_U466 , P2_R2278_U467 , P2_R2278_U468 , P2_R2278_U469 , P2_R2278_U470 , P2_R2278_U471 , P2_R2278_U472 , P2_R2278_U473 , P2_R2278_U474;
wire P2_R2278_U475 , P2_R2278_U476 , P2_R2278_U477 , P2_R2278_U478 , P2_R2278_U479 , P2_R2278_U480 , P2_R2278_U481 , P2_R2278_U482 , P2_R2278_U483 , P2_R2278_U484;
wire P2_R2278_U485 , P2_R2278_U486 , P2_R2278_U487 , P2_R2278_U488 , P2_R2278_U489 , P2_R2278_U490 , P2_R2278_U491 , P2_R2278_U492 , P2_R2278_U493 , P2_R2278_U494;
wire P2_R2278_U495 , P2_R2278_U496 , P2_R2278_U497 , P2_R2278_U498 , P2_R2278_U499 , P2_R2278_U500 , P2_R2278_U501 , P2_R2278_U502 , P2_R2278_U503 , P2_R2278_U504;
wire P2_R2278_U505 , P2_R2278_U506 , P2_R2278_U507 , P2_R2278_U508 , P2_R2278_U509 , P2_R2278_U510 , P2_R2278_U511 , P2_R2278_U512 , P2_R2278_U513 , P2_R2278_U514;
wire P2_R2278_U515 , P2_R2278_U516 , P2_R2278_U517 , P2_R2278_U518 , P2_R2278_U519 , P2_R2278_U520 , P2_R2278_U521 , P2_R2278_U522 , P2_R2278_U523 , P2_R2278_U524;
wire P2_R2278_U525 , P2_R2278_U526 , P2_R2278_U527 , P2_R2278_U528 , P2_R2278_U529 , P2_R2278_U530 , P2_R2278_U531 , P2_R2278_U532 , P2_R2278_U533 , P2_R2278_U534;
wire P2_R2278_U535 , P2_R2278_U536 , P2_R2278_U537 , P2_R2278_U538 , P2_R2278_U539 , P2_R2278_U540 , P2_R2278_U541 , P2_R2278_U542 , P2_R2278_U543 , P2_R2278_U544;
wire P2_R2278_U545 , P2_R2278_U546 , P2_R2278_U547 , P2_R2278_U548 , P2_R2278_U549 , P2_R2278_U550 , P2_R2278_U551 , P2_R2278_U552 , P2_R2278_U553 , P2_R2278_U554;
wire P2_R2278_U555 , P2_R2278_U556 , P2_R2278_U557 , P2_R2278_U558 , P2_R2278_U559 , P2_R2278_U560 , P2_R2278_U561 , P2_R2278_U562 , P2_SUB_450_U6 , P2_SUB_450_U7;
wire P2_SUB_450_U8 , P2_SUB_450_U9 , P2_SUB_450_U10 , P2_SUB_450_U11 , P2_SUB_450_U12 , P2_SUB_450_U13 , P2_SUB_450_U14 , P2_SUB_450_U15 , P2_SUB_450_U16 , P2_SUB_450_U17;
wire P2_SUB_450_U18 , P2_SUB_450_U19 , P2_SUB_450_U20 , P2_SUB_450_U21 , P2_SUB_450_U22 , P2_SUB_450_U23 , P2_SUB_450_U24 , P2_SUB_450_U25 , P2_SUB_450_U26 , P2_SUB_450_U27;
wire P2_SUB_450_U28 , P2_SUB_450_U29 , P2_SUB_450_U30 , P2_SUB_450_U31 , P2_SUB_450_U32 , P2_SUB_450_U33 , P2_SUB_450_U34 , P2_SUB_450_U35 , P2_SUB_450_U36 , P2_SUB_450_U37;
wire P2_SUB_450_U38 , P2_SUB_450_U39 , P2_SUB_450_U40 , P2_SUB_450_U41 , P2_SUB_450_U42 , P2_SUB_450_U43 , P2_SUB_450_U44 , P2_SUB_450_U45 , P2_SUB_450_U46 , P2_SUB_450_U47;
wire P2_SUB_450_U48 , P2_SUB_450_U49 , P2_SUB_450_U50 , P2_SUB_450_U51 , P2_SUB_450_U52 , P2_SUB_450_U53 , P2_SUB_450_U54 , P2_SUB_450_U55 , P2_SUB_450_U56 , P2_SUB_450_U57;
wire P2_SUB_450_U58 , P2_SUB_450_U59 , P2_SUB_450_U60 , P2_SUB_450_U61 , P2_SUB_450_U62 , P2_SUB_450_U63 , P2_R2088_U6 , P2_R2088_U7 , P2_ADD_394_U4 , P2_ADD_394_U5;
wire P2_ADD_394_U6 , P2_ADD_394_U7 , P2_ADD_394_U8 , P2_ADD_394_U9 , P2_ADD_394_U10 , P2_ADD_394_U11 , P2_ADD_394_U12 , P2_ADD_394_U13 , P2_ADD_394_U14 , P2_ADD_394_U15;
wire P2_ADD_394_U16 , P2_ADD_394_U17 , P2_ADD_394_U18 , P2_ADD_394_U19 , P2_ADD_394_U20 , P2_ADD_394_U21 , P2_ADD_394_U22 , P2_ADD_394_U23 , P2_ADD_394_U24 , P2_ADD_394_U25;
wire P2_ADD_394_U26 , P2_ADD_394_U27 , P2_ADD_394_U28 , P2_ADD_394_U29 , P2_ADD_394_U30 , P2_ADD_394_U31 , P2_ADD_394_U32 , P2_ADD_394_U33 , P2_ADD_394_U34 , P2_ADD_394_U35;
wire P2_ADD_394_U36 , P2_ADD_394_U37 , P2_ADD_394_U38 , P2_ADD_394_U39 , P2_ADD_394_U40 , P2_ADD_394_U41 , P2_ADD_394_U42 , P2_ADD_394_U43 , P2_ADD_394_U44 , P2_ADD_394_U45;
wire P2_ADD_394_U46 , P2_ADD_394_U47 , P2_ADD_394_U48 , P2_ADD_394_U49 , P2_ADD_394_U50 , P2_ADD_394_U51 , P2_ADD_394_U52 , P2_ADD_394_U53 , P2_ADD_394_U54 , P2_ADD_394_U55;
wire P2_ADD_394_U56 , P2_ADD_394_U57 , P2_ADD_394_U58 , P2_ADD_394_U59 , P2_ADD_394_U60 , P2_ADD_394_U61 , P2_ADD_394_U62 , P2_ADD_394_U63 , P2_ADD_394_U64 , P2_ADD_394_U65;
wire P2_ADD_394_U66 , P2_ADD_394_U67 , P2_ADD_394_U68 , P2_ADD_394_U69 , P2_ADD_394_U70 , P2_ADD_394_U71 , P2_ADD_394_U72 , P2_ADD_394_U73 , P2_ADD_394_U74 , P2_ADD_394_U75;
wire P2_ADD_394_U76 , P2_ADD_394_U77 , P2_ADD_394_U78 , P2_ADD_394_U79 , P2_ADD_394_U80 , P2_ADD_394_U81 , P2_ADD_394_U82 , P2_ADD_394_U83 , P2_ADD_394_U84 , P2_ADD_394_U85;
wire P2_ADD_394_U86 , P2_ADD_394_U87 , P2_ADD_394_U88 , P2_ADD_394_U89 , P2_ADD_394_U90 , P2_ADD_394_U91 , P2_ADD_394_U92 , P2_ADD_394_U93 , P2_ADD_394_U94 , P2_ADD_394_U95;
wire P2_ADD_394_U96 , P2_ADD_394_U97 , P2_ADD_394_U98 , P2_ADD_394_U99 , P2_ADD_394_U100 , P2_ADD_394_U101 , P2_ADD_394_U102 , P2_ADD_394_U103 , P2_ADD_394_U104 , P2_ADD_394_U105;
wire P2_ADD_394_U106 , P2_ADD_394_U107 , P2_ADD_394_U108 , P2_ADD_394_U109 , P2_ADD_394_U110 , P2_ADD_394_U111 , P2_ADD_394_U112 , P2_ADD_394_U113 , P2_ADD_394_U114 , P2_ADD_394_U115;
wire P2_ADD_394_U116 , P2_ADD_394_U117 , P2_ADD_394_U118 , P2_ADD_394_U119 , P2_ADD_394_U120 , P2_ADD_394_U121 , P2_ADD_394_U122 , P2_ADD_394_U123 , P2_ADD_394_U124 , P2_ADD_394_U125;
wire P2_ADD_394_U126 , P2_ADD_394_U127 , P2_ADD_394_U128 , P2_ADD_394_U129 , P2_ADD_394_U130 , P2_ADD_394_U131 , P2_ADD_394_U132 , P2_ADD_394_U133 , P2_ADD_394_U134 , P2_ADD_394_U135;
wire P2_ADD_394_U136 , P2_ADD_394_U137 , P2_ADD_394_U138 , P2_ADD_394_U139 , P2_ADD_394_U140 , P2_ADD_394_U141 , P2_ADD_394_U142 , P2_ADD_394_U143 , P2_ADD_394_U144 , P2_ADD_394_U145;
wire P2_ADD_394_U146 , P2_ADD_394_U147 , P2_ADD_394_U148 , P2_ADD_394_U149 , P2_ADD_394_U150 , P2_ADD_394_U151 , P2_ADD_394_U152 , P2_ADD_394_U153 , P2_ADD_394_U154 , P2_ADD_394_U155;
wire P2_ADD_394_U156 , P2_ADD_394_U157 , P2_ADD_394_U158 , P2_ADD_394_U159 , P2_ADD_394_U160 , P2_ADD_394_U161 , P2_ADD_394_U162 , P2_ADD_394_U163 , P2_ADD_394_U164 , P2_ADD_394_U165;
wire P2_ADD_394_U166 , P2_ADD_394_U167 , P2_ADD_394_U168 , P2_ADD_394_U169 , P2_ADD_394_U170 , P2_ADD_394_U171 , P2_ADD_394_U172 , P2_ADD_394_U173 , P2_ADD_394_U174 , P2_ADD_394_U175;
wire P2_ADD_394_U176 , P2_ADD_394_U177 , P2_ADD_394_U178 , P2_ADD_394_U179 , P2_ADD_394_U180 , P2_ADD_394_U181 , P2_ADD_394_U182 , P2_ADD_394_U183 , P2_ADD_394_U184 , P2_ADD_394_U185;
wire P2_ADD_394_U186 , P2_R2267_U6 , P2_R2267_U7 , P2_R2267_U8 , P2_R2267_U9 , P2_R2267_U10 , P2_R2267_U11 , P2_R2267_U12 , P2_R2267_U13 , P2_R2267_U14;
wire P2_R2267_U15 , P2_R2267_U16 , P2_R2267_U17 , P2_R2267_U18 , P2_R2267_U19 , P2_R2267_U20 , P2_R2267_U21 , P2_R2267_U22 , P2_R2267_U23 , P2_R2267_U24;
wire P2_R2267_U25 , P2_R2267_U26 , P2_R2267_U27 , P2_R2267_U28 , P2_R2267_U29 , P2_R2267_U30 , P2_R2267_U31 , P2_R2267_U32 , P2_R2267_U33 , P2_R2267_U34;
wire P2_R2267_U35 , P2_R2267_U36 , P2_R2267_U37 , P2_R2267_U38 , P2_R2267_U39 , P2_R2267_U40 , P2_R2267_U41 , P2_R2267_U42 , P2_R2267_U43 , P2_R2267_U44;
wire P2_R2267_U45 , P2_R2267_U46 , P2_R2267_U47 , P2_R2267_U48 , P2_R2267_U49 , P2_R2267_U50 , P2_R2267_U51 , P2_R2267_U52 , P2_R2267_U53 , P2_R2267_U54;
wire P2_R2267_U55 , P2_R2267_U56 , P2_R2267_U57 , P2_R2267_U58 , P2_R2267_U59 , P2_R2267_U60 , P2_R2267_U61 , P2_R2267_U62 , P2_R2267_U63 , P2_R2267_U64;
wire P2_R2267_U65 , P2_R2267_U66 , P2_R2267_U67 , P2_R2267_U68 , P2_R2267_U69 , P2_R2267_U70 , P2_R2267_U71 , P2_R2267_U72 , P2_R2267_U73 , P2_R2267_U74;
wire P2_R2267_U75 , P2_R2267_U76 , P2_R2267_U77 , P2_R2267_U78 , P2_R2267_U79 , P2_R2267_U80 , P2_R2267_U81 , P2_R2267_U82 , P2_R2267_U83 , P2_R2267_U84;
wire P2_R2267_U85 , P2_R2267_U86 , P2_R2267_U87 , P2_R2267_U88 , P2_R2267_U89 , P2_R2267_U90 , P2_R2267_U91 , P2_R2267_U92 , P2_R2267_U93 , P2_R2267_U94;
wire P2_R2267_U95 , P2_R2267_U96 , P2_R2267_U97 , P2_R2267_U98 , P2_R2267_U99 , P2_R2267_U100 , P2_R2267_U101 , P2_R2267_U102 , P2_R2267_U103 , P2_R2267_U104;
wire P2_R2267_U105 , P2_R2267_U106 , P2_R2267_U107 , P2_R2267_U108 , P2_R2267_U109 , P2_R2267_U110 , P2_R2267_U111 , P2_R2267_U112 , P2_R2267_U113 , P2_R2267_U114;
wire P2_R2267_U115 , P2_R2267_U116 , P2_R2267_U117 , P2_R2267_U118 , P2_R2267_U119 , P2_R2267_U120 , P2_R2267_U121 , P2_R2267_U122 , P2_R2267_U123 , P2_R2267_U124;
wire P2_R2267_U125 , P2_R2267_U126 , P2_R2267_U127 , P2_R2267_U128 , P2_R2267_U129 , P2_R2267_U130 , P2_R2267_U131 , P2_R2267_U132 , P2_R2267_U133 , P2_R2267_U134;
wire P2_R2267_U135 , P2_R2267_U136 , P2_R2267_U137 , P2_R2267_U138 , P2_R2267_U139 , P2_R2267_U140 , P2_R2267_U141 , P2_R2267_U142 , P2_R2267_U143 , P2_R2267_U144;
wire P2_R2267_U145 , P2_R2267_U146 , P2_R2267_U147 , P2_R2267_U148 , P2_R2267_U149 , P2_R2267_U150 , P2_R2267_U151 , P2_R2267_U152 , P2_R2267_U153 , P2_R2267_U154;
wire P2_R2267_U155 , P2_R2267_U156 , P2_R2267_U157 , P2_R2267_U158 , P2_R2267_U159 , P2_R2267_U160 , P2_R2267_U161 , P2_R2267_U162 , P2_R2267_U163 , P2_R2267_U164;
wire P2_R2267_U165 , P2_R2267_U166 , P2_ADD_371_1212_U4 , P2_ADD_371_1212_U5 , P2_ADD_371_1212_U6 , P2_ADD_371_1212_U7 , P2_ADD_371_1212_U8 , P2_ADD_371_1212_U9 , P2_ADD_371_1212_U10 , P2_ADD_371_1212_U11;
wire P2_ADD_371_1212_U12 , P2_ADD_371_1212_U13 , P2_ADD_371_1212_U14 , P2_ADD_371_1212_U15 , P2_ADD_371_1212_U16 , P2_ADD_371_1212_U17 , P2_ADD_371_1212_U18 , P2_ADD_371_1212_U19 , P2_ADD_371_1212_U20 , P2_ADD_371_1212_U21;
wire P2_ADD_371_1212_U22 , P2_ADD_371_1212_U23 , P2_ADD_371_1212_U24 , P2_ADD_371_1212_U25 , P2_ADD_371_1212_U26 , P2_ADD_371_1212_U27 , P2_ADD_371_1212_U28 , P2_ADD_371_1212_U29 , P2_ADD_371_1212_U30 , P2_ADD_371_1212_U31;
wire P2_ADD_371_1212_U32 , P2_ADD_371_1212_U33 , P2_ADD_371_1212_U34 , P2_ADD_371_1212_U35 , P2_ADD_371_1212_U36 , P2_ADD_371_1212_U37 , P2_ADD_371_1212_U38 , P2_ADD_371_1212_U39 , P2_ADD_371_1212_U40 , P2_ADD_371_1212_U41;
wire P2_ADD_371_1212_U42 , P2_ADD_371_1212_U43 , P2_ADD_371_1212_U44 , P2_ADD_371_1212_U45 , P2_ADD_371_1212_U46 , P2_ADD_371_1212_U47 , P2_ADD_371_1212_U48 , P2_ADD_371_1212_U49 , P2_ADD_371_1212_U50 , P2_ADD_371_1212_U51;
wire P2_ADD_371_1212_U52 , P2_ADD_371_1212_U53 , P2_ADD_371_1212_U54 , P2_ADD_371_1212_U55 , P2_ADD_371_1212_U56 , P2_ADD_371_1212_U57 , P2_ADD_371_1212_U58 , P2_ADD_371_1212_U59 , P2_ADD_371_1212_U60 , P2_ADD_371_1212_U61;
wire P2_ADD_371_1212_U62 , P2_ADD_371_1212_U63 , P2_ADD_371_1212_U64 , P2_ADD_371_1212_U65 , P2_ADD_371_1212_U66 , P2_ADD_371_1212_U67 , P2_ADD_371_1212_U68 , P2_ADD_371_1212_U69 , P2_ADD_371_1212_U70 , P2_ADD_371_1212_U71;
wire P2_ADD_371_1212_U72 , P2_ADD_371_1212_U73 , P2_ADD_371_1212_U74 , P2_ADD_371_1212_U75 , P2_ADD_371_1212_U76 , P2_ADD_371_1212_U77 , P2_ADD_371_1212_U78 , P2_ADD_371_1212_U79 , P2_ADD_371_1212_U80 , P2_ADD_371_1212_U81;
wire P2_ADD_371_1212_U82 , P2_ADD_371_1212_U83 , P2_ADD_371_1212_U84 , P2_ADD_371_1212_U85 , P2_ADD_371_1212_U86 , P2_ADD_371_1212_U87 , P2_ADD_371_1212_U88 , P2_ADD_371_1212_U89 , P2_ADD_371_1212_U90 , P2_ADD_371_1212_U91;
wire P2_ADD_371_1212_U92 , P2_ADD_371_1212_U93 , P2_ADD_371_1212_U94 , P2_ADD_371_1212_U95 , P2_ADD_371_1212_U96 , P2_ADD_371_1212_U97 , P2_ADD_371_1212_U98 , P2_ADD_371_1212_U99 , P2_ADD_371_1212_U100 , P2_ADD_371_1212_U101;
wire P2_ADD_371_1212_U102 , P2_ADD_371_1212_U103 , P2_ADD_371_1212_U104 , P2_ADD_371_1212_U105 , P2_ADD_371_1212_U106 , P2_ADD_371_1212_U107 , P2_ADD_371_1212_U108 , P2_ADD_371_1212_U109 , P2_ADD_371_1212_U110 , P2_ADD_371_1212_U111;
wire P2_ADD_371_1212_U112 , P2_ADD_371_1212_U113 , P2_ADD_371_1212_U114 , P2_ADD_371_1212_U115 , P2_ADD_371_1212_U116 , P2_ADD_371_1212_U117 , P2_ADD_371_1212_U118 , P2_ADD_371_1212_U119 , P2_ADD_371_1212_U120 , P2_ADD_371_1212_U121;
wire P2_ADD_371_1212_U122 , P2_ADD_371_1212_U123 , P2_ADD_371_1212_U124 , P2_ADD_371_1212_U125 , P2_ADD_371_1212_U126 , P2_ADD_371_1212_U127 , P2_ADD_371_1212_U128 , P2_ADD_371_1212_U129 , P2_ADD_371_1212_U130 , P2_ADD_371_1212_U131;
wire P2_ADD_371_1212_U132 , P2_ADD_371_1212_U133 , P2_ADD_371_1212_U134 , P2_ADD_371_1212_U135 , P2_ADD_371_1212_U136 , P2_ADD_371_1212_U137 , P2_ADD_371_1212_U138 , P2_ADD_371_1212_U139 , P2_ADD_371_1212_U140 , P2_ADD_371_1212_U141;
wire P2_ADD_371_1212_U142 , P2_ADD_371_1212_U143 , P2_ADD_371_1212_U144 , P2_ADD_371_1212_U145 , P2_ADD_371_1212_U146 , P2_ADD_371_1212_U147 , P2_ADD_371_1212_U148 , P2_ADD_371_1212_U149 , P2_ADD_371_1212_U150 , P2_ADD_371_1212_U151;
wire P2_ADD_371_1212_U152 , P2_ADD_371_1212_U153 , P2_ADD_371_1212_U154 , P2_ADD_371_1212_U155 , P2_ADD_371_1212_U156 , P2_ADD_371_1212_U157 , P2_ADD_371_1212_U158 , P2_ADD_371_1212_U159 , P2_ADD_371_1212_U160 , P2_ADD_371_1212_U161;
wire P2_ADD_371_1212_U162 , P2_ADD_371_1212_U163 , P2_ADD_371_1212_U164 , P2_ADD_371_1212_U165 , P2_ADD_371_1212_U166 , P2_ADD_371_1212_U167 , P2_ADD_371_1212_U168 , P2_ADD_371_1212_U169 , P2_ADD_371_1212_U170 , P2_ADD_371_1212_U171;
wire P2_ADD_371_1212_U172 , P2_ADD_371_1212_U173 , P2_ADD_371_1212_U174 , P2_ADD_371_1212_U175 , P2_ADD_371_1212_U176 , P2_ADD_371_1212_U177 , P2_ADD_371_1212_U178 , P2_ADD_371_1212_U179 , P2_ADD_371_1212_U180 , P2_ADD_371_1212_U181;
wire P2_ADD_371_1212_U182 , P2_ADD_371_1212_U183 , P2_ADD_371_1212_U184 , P2_ADD_371_1212_U185 , P2_ADD_371_1212_U186 , P2_ADD_371_1212_U187 , P2_ADD_371_1212_U188 , P2_ADD_371_1212_U189 , P2_ADD_371_1212_U190 , P2_ADD_371_1212_U191;
wire P2_ADD_371_1212_U192 , P2_ADD_371_1212_U193 , P2_ADD_371_1212_U194 , P2_ADD_371_1212_U195 , P2_ADD_371_1212_U196 , P2_ADD_371_1212_U197 , P2_ADD_371_1212_U198 , P2_ADD_371_1212_U199 , P2_ADD_371_1212_U200 , P2_ADD_371_1212_U201;
wire P2_ADD_371_1212_U202 , P2_ADD_371_1212_U203 , P2_ADD_371_1212_U204 , P2_ADD_371_1212_U205 , P2_ADD_371_1212_U206 , P2_ADD_371_1212_U207 , P2_ADD_371_1212_U208 , P2_ADD_371_1212_U209 , P2_ADD_371_1212_U210 , P2_ADD_371_1212_U211;
wire P2_ADD_371_1212_U212 , P2_ADD_371_1212_U213 , P2_ADD_371_1212_U214 , P2_ADD_371_1212_U215 , P2_ADD_371_1212_U216 , P2_ADD_371_1212_U217 , P2_ADD_371_1212_U218 , P2_ADD_371_1212_U219 , P2_ADD_371_1212_U220 , P2_ADD_371_1212_U221;
wire P2_ADD_371_1212_U222 , P2_ADD_371_1212_U223 , P2_ADD_371_1212_U224 , P2_ADD_371_1212_U225 , P2_ADD_371_1212_U226 , P2_ADD_371_1212_U227 , P2_ADD_371_1212_U228 , P2_ADD_371_1212_U229 , P2_ADD_371_1212_U230 , P2_ADD_371_1212_U231;
wire P2_ADD_371_1212_U232 , P2_ADD_371_1212_U233 , P2_ADD_371_1212_U234 , P2_ADD_371_1212_U235 , P2_ADD_371_1212_U236 , P2_ADD_371_1212_U237 , P2_ADD_371_1212_U238 , P2_ADD_371_1212_U239 , P2_ADD_371_1212_U240 , P2_ADD_371_1212_U241;
wire P2_ADD_371_1212_U242 , P2_ADD_371_1212_U243 , P2_ADD_371_1212_U244 , P2_ADD_371_1212_U245 , P2_ADD_371_1212_U246 , P2_ADD_371_1212_U247 , P2_ADD_371_1212_U248 , P2_ADD_371_1212_U249 , P2_ADD_371_1212_U250 , P2_ADD_371_1212_U251;
wire P2_ADD_371_1212_U252 , P2_ADD_371_1212_U253 , P2_ADD_371_1212_U254 , P2_ADD_371_1212_U255 , P2_ADD_371_1212_U256 , P2_ADD_371_1212_U257 , P2_ADD_371_1212_U258 , P2_ADD_371_1212_U259 , P2_ADD_371_1212_U260 , P2_ADD_371_1212_U261;
wire P2_ADD_371_1212_U262 , P2_ADD_371_1212_U263 , P2_ADD_371_1212_U264 , P2_ADD_371_1212_U265 , P2_ADD_371_1212_U266 , P2_ADD_371_1212_U267 , P2_ADD_371_1212_U268 , P2_ADD_371_1212_U269 , P2_ADD_371_1212_U270 , P2_ADD_371_1212_U271;
wire P2_ADD_371_1212_U272 , P2_ADD_371_1212_U273 , P2_ADD_371_1212_U274 , P2_ADD_371_1212_U275 , P2_ADD_371_1212_U276 , P2_ADD_371_1212_U277 , P2_ADD_371_1212_U278 , P2_ADD_371_1212_U279 , P2_ADD_371_1212_U280 , P2_ADD_371_1212_U281;
wire P2_ADD_371_1212_U282 , P1_R2027_U5 , P1_R2027_U6 , P1_R2027_U7 , P1_R2027_U8 , P1_R2027_U9 , P1_R2027_U10 , P1_R2027_U11 , P1_R2027_U12 , P1_R2027_U13;
wire P1_R2027_U14 , P1_R2027_U15 , P1_R2027_U16 , P1_R2027_U17 , P1_R2027_U18 , P1_R2027_U19 , P1_R2027_U20 , P1_R2027_U21 , P1_R2027_U22 , P1_R2027_U23;
wire P1_R2027_U24 , P1_R2027_U25 , P1_R2027_U26 , P1_R2027_U27 , P1_R2027_U28 , P1_R2027_U29 , P1_R2027_U30 , P1_R2027_U31 , P1_R2027_U32 , P1_R2027_U33;
wire P1_R2027_U34 , P1_R2027_U35 , P1_R2027_U36 , P1_R2027_U37 , P1_R2027_U38 , P1_R2027_U39 , P1_R2027_U40 , P1_R2027_U41 , P1_R2027_U42 , P1_R2027_U43;
wire P1_R2027_U44 , P1_R2027_U45 , P1_R2027_U46 , P1_R2027_U47 , P1_R2027_U48 , P1_R2027_U49 , P1_R2027_U50 , P1_R2027_U51 , P1_R2027_U52 , P1_R2027_U53;
wire P1_R2027_U54 , P1_R2027_U55 , P1_R2027_U56 , P1_R2027_U57 , P1_R2027_U58 , P1_R2027_U59 , P1_R2027_U60 , P1_R2027_U61 , P1_R2027_U62 , P1_R2027_U63;
wire P1_R2027_U64 , P1_R2027_U65 , P1_R2027_U66 , P1_R2027_U67 , P1_R2027_U68 , P1_R2027_U69 , P1_R2027_U70 , P1_R2027_U71 , P1_R2027_U72 , P1_R2027_U73;
wire P1_R2027_U74 , P1_R2027_U75 , P1_R2027_U76 , P1_R2027_U77 , P1_R2027_U78 , P1_R2027_U79 , P1_R2027_U80 , P1_R2027_U81 , P1_R2027_U82 , P1_R2027_U83;
wire P1_R2027_U84 , P1_R2027_U85 , P1_R2027_U86 , P1_R2027_U87 , P1_R2027_U88 , P1_R2027_U89 , P1_R2027_U90 , P1_R2027_U91 , P1_R2027_U92 , P1_R2027_U93;
wire P1_R2027_U94 , P1_R2027_U95 , P1_R2027_U96 , P1_R2027_U97 , P1_R2027_U98 , P1_R2027_U99 , P1_R2027_U100 , P1_R2027_U101 , P1_R2027_U102 , P1_R2027_U103;
wire P1_R2027_U104 , P1_R2027_U105 , P1_R2027_U106 , P1_R2027_U107 , P1_R2027_U108 , P1_R2027_U109 , P1_R2027_U110 , P1_R2027_U111 , P1_R2027_U112 , P1_R2027_U113;
wire P1_R2027_U114 , P1_R2027_U115 , P1_R2027_U116 , P1_R2027_U117 , P1_R2027_U118 , P1_R2027_U119 , P1_R2027_U120 , P1_R2027_U121 , P1_R2027_U122 , P1_R2027_U123;
wire P1_R2027_U124 , P1_R2027_U125 , P1_R2027_U126 , P1_R2027_U127 , P1_R2027_U128 , P1_R2027_U129 , P1_R2027_U130 , P1_R2027_U131 , P1_R2027_U132 , P1_R2027_U133;
wire P1_R2027_U134 , P1_R2027_U135 , P1_R2027_U136 , P1_R2027_U137 , P1_R2027_U138 , P1_R2027_U139 , P1_R2027_U140 , P1_R2027_U141 , P1_R2027_U142 , P1_R2027_U143;
wire P1_R2027_U144 , P1_R2027_U145 , P1_R2027_U146 , P1_R2027_U147 , P1_R2027_U148 , P1_R2027_U149 , P1_R2027_U150 , P1_R2027_U151 , P1_R2027_U152 , P1_R2027_U153;
wire P1_R2027_U154 , P1_R2027_U155 , P1_R2027_U156 , P1_R2027_U157 , P1_R2027_U158 , P1_R2027_U159 , P1_R2027_U160 , P1_R2027_U161 , P1_R2027_U162 , P1_R2027_U163;
wire P1_R2027_U164 , P1_R2027_U165 , P1_R2027_U166 , P1_R2027_U167 , P1_R2027_U168 , P1_R2027_U169 , P1_R2027_U170 , P1_R2027_U171 , P1_R2027_U172 , P1_R2027_U173;
wire P1_R2027_U174 , P1_R2027_U175 , P1_R2027_U176 , P1_R2027_U177 , P1_R2027_U178 , P1_R2027_U179 , P1_R2027_U180 , P1_R2027_U181 , P1_R2027_U182 , P1_R2027_U183;
wire P1_R2027_U184 , P1_R2027_U185 , P1_R2027_U186 , P1_R2027_U187 , P1_R2027_U188 , P1_R2027_U189 , P1_R2027_U190 , P1_R2027_U191 , P1_R2027_U192 , P1_R2027_U193;
wire P1_R2027_U194 , P1_R2027_U195 , P1_R2027_U196 , P1_R2027_U197 , P1_R2027_U198 , P1_R2027_U199 , P1_R2027_U200 , P1_R2027_U201 , P1_R2027_U202 , P1_R2182_U5;
wire P1_R2182_U6 , P1_R2182_U7 , P1_R2182_U8 , P1_R2182_U9 , P1_R2182_U10 , P1_R2182_U11 , P1_R2182_U12 , P1_R2182_U13 , P1_R2182_U14 , P1_R2182_U15;
wire P1_R2182_U16 , P1_R2182_U17 , P1_R2182_U18 , P1_R2182_U19 , P1_R2182_U20 , P1_R2182_U21 , P1_R2182_U22 , P1_R2182_U23 , P1_R2182_U24 , P1_R2182_U25;
wire P1_R2182_U26 , P1_R2182_U27 , P1_R2182_U28 , P1_R2182_U29 , P1_R2182_U30 , P1_R2182_U31 , P1_R2182_U32 , P1_R2182_U33 , P1_R2182_U34 , P1_R2182_U35;
wire P1_R2182_U36 , P1_R2182_U37 , P1_R2182_U38 , P1_R2182_U39 , P1_R2182_U40 , P1_R2182_U41 , P1_R2182_U42 , P1_R2182_U43 , P1_R2182_U44 , P1_R2182_U45;
wire P1_R2182_U46 , P1_R2182_U47 , P1_R2182_U48 , P1_R2182_U49 , P1_R2182_U50 , P1_R2182_U51 , P1_R2182_U52 , P1_R2182_U53 , P1_R2182_U54 , P1_R2182_U55;
wire P1_R2182_U56 , P1_R2182_U57 , P1_R2182_U58 , P1_R2182_U59 , P1_R2182_U60 , P1_R2182_U61 , P1_R2182_U62 , P1_R2182_U63 , P1_R2182_U64 , P1_R2182_U65;
wire P1_R2182_U66 , P1_R2182_U67 , P1_R2182_U68 , P1_R2182_U69 , P1_R2182_U70 , P1_R2182_U71 , P1_R2182_U72 , P1_R2182_U73 , P1_R2182_U74 , P1_R2182_U75;
wire P1_R2182_U76 , P1_R2182_U77 , P1_R2182_U78 , P1_R2182_U79 , P1_R2182_U80 , P1_R2182_U81 , P1_R2182_U82 , P1_R2182_U83 , P1_R2182_U84 , P1_R2182_U85;
wire P1_R2182_U86 , P1_R2144_U5 , P1_R2144_U6 , P1_R2144_U7 , P1_R2144_U8 , P1_R2144_U9 , P1_R2144_U10 , P1_R2144_U11 , P1_R2144_U12 , P1_R2144_U13;
wire P1_R2144_U14 , P1_R2144_U15 , P1_R2144_U16 , P1_R2144_U17 , P1_R2144_U18 , P1_R2144_U19 , P1_R2144_U20 , P1_R2144_U21 , P1_R2144_U22 , P1_R2144_U23;
wire P1_R2144_U24 , P1_R2144_U25 , P1_R2144_U26 , P1_R2144_U27 , P1_R2144_U28 , P1_R2144_U29 , P1_R2144_U30 , P1_R2144_U31 , P1_R2144_U32 , P1_R2144_U33;
wire P1_R2144_U34 , P1_R2144_U35 , P1_R2144_U36 , P1_R2144_U37 , P1_R2144_U38 , P1_R2144_U39 , P1_R2144_U40 , P1_R2144_U41 , P1_R2144_U42 , P1_R2144_U43;
wire P1_R2144_U44 , P1_R2144_U45 , P1_R2144_U46 , P1_R2144_U47 , P1_R2144_U48 , P1_R2144_U49 , P1_R2144_U50 , P1_R2144_U51 , P1_R2144_U52 , P1_R2144_U53;
wire P1_R2144_U54 , P1_R2144_U55 , P1_R2144_U56 , P1_R2144_U57 , P1_R2144_U58 , P1_R2144_U59 , P1_R2144_U60 , P1_R2144_U61 , P1_R2144_U62 , P1_R2144_U63;
wire P1_R2144_U64 , P1_R2144_U65 , P1_R2144_U66 , P1_R2144_U67 , P1_R2144_U68 , P1_R2144_U69 , P1_R2144_U70 , P1_R2144_U71 , P1_R2144_U72 , P1_R2144_U73;
wire P1_R2144_U74 , P1_R2144_U75 , P1_R2144_U76 , P1_R2144_U77 , P1_R2144_U78 , P1_R2144_U79 , P1_R2144_U80 , P1_R2144_U81 , P1_R2144_U82 , P1_R2144_U83;
wire P1_R2144_U84 , P1_R2144_U85 , P1_R2144_U86 , P1_R2144_U87 , P1_R2144_U88 , P1_R2144_U89 , P1_R2144_U90 , P1_R2144_U91 , P1_R2144_U92 , P1_R2144_U93;
wire P1_R2144_U94 , P1_R2144_U95 , P1_R2144_U96 , P1_R2144_U97 , P1_R2144_U98 , P1_R2144_U99 , P1_R2144_U100 , P1_R2144_U101 , P1_R2144_U102 , P1_R2144_U103;
wire P1_R2144_U104 , P1_R2144_U105 , P1_R2144_U106 , P1_R2144_U107 , P1_R2144_U108 , P1_R2144_U109 , P1_R2144_U110 , P1_R2144_U111 , P1_R2144_U112 , P1_R2144_U113;
wire P1_R2144_U114 , P1_R2144_U115 , P1_R2144_U116 , P1_R2144_U117 , P1_R2144_U118 , P1_R2144_U119 , P1_R2144_U120 , P1_R2144_U121 , P1_R2144_U122 , P1_R2144_U123;
wire P1_R2144_U124 , P1_R2144_U125 , P1_R2144_U126 , P1_R2144_U127 , P1_R2144_U128 , P1_R2144_U129 , P1_R2144_U130 , P1_R2144_U131 , P1_R2144_U132 , P1_R2144_U133;
wire P1_R2144_U134 , P1_R2144_U135 , P1_R2144_U136 , P1_R2144_U137 , P1_R2144_U138 , P1_R2144_U139 , P1_R2144_U140 , P1_R2144_U141 , P1_R2144_U142 , P1_R2144_U143;
wire P1_R2144_U144 , P1_R2144_U145 , P1_R2144_U146 , P1_R2144_U147 , P1_R2144_U148 , P1_R2144_U149 , P1_R2144_U150 , P1_R2144_U151 , P1_R2144_U152 , P1_R2144_U153;
wire P1_R2144_U154 , P1_R2144_U155 , P1_R2144_U156 , P1_R2144_U157 , P1_R2144_U158 , P1_R2144_U159 , P1_R2144_U160 , P1_R2144_U161 , P1_R2144_U162 , P1_R2144_U163;
wire P1_R2144_U164 , P1_R2144_U165 , P1_R2144_U166 , P1_R2144_U167 , P1_R2144_U168 , P1_R2144_U169 , P1_R2144_U170 , P1_R2144_U171 , P1_R2144_U172 , P1_R2144_U173;
wire P1_R2144_U174 , P1_R2144_U175 , P1_R2144_U176 , P1_R2144_U177 , P1_R2144_U178 , P1_R2144_U179 , P1_R2144_U180 , P1_R2144_U181 , P1_R2144_U182 , P1_R2144_U183;
wire P1_R2144_U184 , P1_R2144_U185 , P1_R2144_U186 , P1_R2144_U187 , P1_R2144_U188 , P1_R2144_U189 , P1_R2144_U190 , P1_R2144_U191 , P1_R2144_U192 , P1_R2144_U193;
wire P1_R2144_U194 , P1_R2144_U195 , P1_R2144_U196 , P1_R2144_U197 , P1_R2144_U198 , P1_R2144_U199 , P1_R2144_U200 , P1_R2144_U201 , P1_R2144_U202 , P1_R2144_U203;
wire P1_R2144_U204 , P1_R2144_U205 , P1_R2144_U206 , P1_R2144_U207 , P1_R2144_U208 , P1_R2144_U209 , P1_R2144_U210 , P1_R2144_U211 , P1_R2144_U212 , P1_R2144_U213;
wire P1_R2144_U214 , P1_R2144_U215 , P1_R2144_U216 , P1_R2144_U217 , P1_R2144_U218 , P1_R2144_U219 , P1_R2144_U220 , P1_R2144_U221 , P1_R2144_U222 , P1_R2144_U223;
wire P1_R2144_U224 , P1_R2144_U225 , P1_R2144_U226 , P1_R2144_U227 , P1_R2144_U228 , P1_R2144_U229 , P1_R2144_U230 , P1_R2144_U231 , P1_R2144_U232 , P1_R2144_U233;
wire P1_R2144_U234 , P1_R2144_U235 , P1_R2144_U236 , P1_R2144_U237 , P1_R2144_U238 , P1_R2144_U239 , P1_R2144_U240 , P1_R2144_U241 , P1_R2144_U242 , P1_R2144_U243;
wire P1_R2144_U244 , P1_R2144_U245 , P1_R2144_U246 , P1_R2144_U247 , P1_R2144_U248 , P1_R2144_U249 , P1_R2144_U250 , P1_R2144_U251 , P1_R2144_U252 , P1_R2144_U253;
wire P1_R2144_U254 , P1_R2144_U255 , P1_R2144_U256 , P1_R2144_U257 , P1_R2144_U258 , P1_R2144_U259 , P1_R2144_U260 , P1_R2278_U5 , P1_R2278_U6 , P1_R2278_U7;
wire P1_R2278_U8 , P1_R2278_U9 , P1_R2278_U10 , P1_R2278_U11 , P1_R2278_U12 , P1_R2278_U13 , P1_R2278_U14 , P1_R2278_U15 , P1_R2278_U16 , P1_R2278_U17;
wire P1_R2278_U18 , P1_R2278_U19 , P1_R2278_U20 , P1_R2278_U21 , P1_R2278_U22 , P1_R2278_U23 , P1_R2278_U24 , P1_R2278_U25 , P1_R2278_U26 , P1_R2278_U27;
wire P1_R2278_U28 , P1_R2278_U29 , P1_R2278_U30 , P1_R2278_U31 , P1_R2278_U32 , P1_R2278_U33 , P1_R2278_U34 , P1_R2278_U35 , P1_R2278_U36 , P1_R2278_U37;
wire P1_R2278_U38 , P1_R2278_U39 , P1_R2278_U40 , P1_R2278_U41 , P1_R2278_U42 , P1_R2278_U43 , P1_R2278_U44 , P1_R2278_U45 , P1_R2278_U46 , P1_R2278_U47;
wire P1_R2278_U48 , P1_R2278_U49 , P1_R2278_U50 , P1_R2278_U51 , P1_R2278_U52 , P1_R2278_U53 , P1_R2278_U54 , P1_R2278_U55 , P1_R2278_U56 , P1_R2278_U57;
wire P1_R2278_U58 , P1_R2278_U59 , P1_R2278_U60 , P1_R2278_U61 , P1_R2278_U62 , P1_R2278_U63 , P1_R2278_U64 , P1_R2278_U65 , P1_R2278_U66 , P1_R2278_U67;
wire P1_R2278_U68 , P1_R2278_U69 , P1_R2278_U70 , P1_R2278_U71 , P1_R2278_U72 , P1_R2278_U73 , P1_R2278_U74 , P1_R2278_U75 , P1_R2278_U76 , P1_R2278_U77;
wire P1_R2278_U78 , P1_R2278_U79 , P1_R2278_U80 , P1_R2278_U81 , P1_R2278_U82 , P1_R2278_U83 , P1_R2278_U84 , P1_R2278_U85 , P1_R2278_U86 , P1_R2278_U87;
wire P1_R2278_U88 , P1_R2278_U89 , P1_R2278_U90 , P1_R2278_U91 , P1_R2278_U92 , P1_R2278_U93 , P1_R2278_U94 , P1_R2278_U95 , P1_R2278_U96 , P1_R2278_U97;
wire P1_R2278_U98 , P1_R2278_U99 , P1_R2278_U100 , P1_R2278_U101 , P1_R2278_U102 , P1_R2278_U103 , P1_R2278_U104 , P1_R2278_U105 , P1_R2278_U106 , P1_R2278_U107;
wire P1_R2278_U108 , P1_R2278_U109 , P1_R2278_U110 , P1_R2278_U111 , P1_R2278_U112 , P1_R2278_U113 , P1_R2278_U114 , P1_R2278_U115 , P1_R2278_U116 , P1_R2278_U117;
wire P1_R2278_U118 , P1_R2278_U119 , P1_R2278_U120 , P1_R2278_U121 , P1_R2278_U122 , P1_R2278_U123 , P1_R2278_U124 , P1_R2278_U125 , P1_R2278_U126 , P1_R2278_U127;
wire P1_R2278_U128 , P1_R2278_U129 , P1_R2278_U130 , P1_R2278_U131 , P1_R2278_U132 , P1_R2278_U133 , P1_R2278_U134 , P1_R2278_U135 , P1_R2278_U136 , P1_R2278_U137;
wire P1_R2278_U138 , P1_R2278_U139 , P1_R2278_U140 , P1_R2278_U141 , P1_R2278_U142 , P1_R2278_U143 , P1_R2278_U144 , P1_R2278_U145 , P1_R2278_U146 , P1_R2278_U147;
wire P1_R2278_U148 , P1_R2278_U149 , P1_R2278_U150 , P1_R2278_U151 , P1_R2278_U152 , P1_R2278_U153 , P1_R2278_U154 , P1_R2278_U155 , P1_R2278_U156 , P1_R2278_U157;
wire P1_R2278_U158 , P1_R2278_U159 , P1_R2278_U160 , P1_R2278_U161 , P1_R2278_U162 , P1_R2278_U163 , P1_R2278_U164 , P1_R2278_U165 , P1_R2278_U166 , P1_R2278_U167;
wire P1_R2278_U168 , P1_R2278_U169 , P1_R2278_U170 , P1_R2278_U171 , P1_R2278_U172 , P1_R2278_U173 , P1_R2278_U174 , P1_R2278_U175 , P1_R2278_U176 , P1_R2278_U177;
wire P1_R2278_U178 , P1_R2278_U179 , P1_R2278_U180 , P1_R2278_U181 , P1_R2278_U182 , P1_R2278_U183 , P1_R2278_U184 , P1_R2278_U185 , P1_R2278_U186 , P1_R2278_U187;
wire P1_R2278_U188 , P1_R2278_U189 , P1_R2278_U190 , P1_R2278_U191 , P1_R2278_U192 , P1_R2278_U193 , P1_R2278_U194 , P1_R2278_U195 , P1_R2278_U196 , P1_R2278_U197;
wire P1_R2278_U198 , P1_R2278_U199 , P1_R2278_U200 , P1_R2278_U201 , P1_R2278_U202 , P1_R2278_U203 , P1_R2278_U204 , P1_R2278_U205 , P1_R2278_U206 , P1_R2278_U207;
wire P1_R2278_U208 , P1_R2278_U209 , P1_R2278_U210 , P1_R2278_U211 , P1_R2278_U212 , P1_R2278_U213 , P1_R2278_U214 , P1_R2278_U215 , P1_R2278_U216 , P1_R2278_U217;
wire P1_R2278_U218 , P1_R2278_U219 , P1_R2278_U220 , P1_R2278_U221 , P1_R2278_U222 , P1_R2278_U223 , P1_R2278_U224 , P1_R2278_U225 , P1_R2278_U226 , P1_R2278_U227;
wire P1_R2278_U228 , P1_R2278_U229 , P1_R2278_U230 , P1_R2278_U231 , P1_R2278_U232 , P1_R2278_U233 , P1_R2278_U234 , P1_R2278_U235 , P1_R2278_U236 , P1_R2278_U237;
wire P1_R2278_U238 , P1_R2278_U239 , P1_R2278_U240 , P1_R2278_U241 , P1_R2278_U242 , P1_R2278_U243 , P1_R2278_U244 , P1_R2278_U245 , P1_R2278_U246 , P1_R2278_U247;
wire P1_R2278_U248 , P1_R2278_U249 , P1_R2278_U250 , P1_R2278_U251 , P1_R2278_U252 , P1_R2278_U253 , P1_R2278_U254 , P1_R2278_U255 , P1_R2278_U256 , P1_R2278_U257;
wire P1_R2278_U258 , P1_R2278_U259 , P1_R2278_U260 , P1_R2278_U261 , P1_R2278_U262 , P1_R2278_U263 , P1_R2278_U264 , P1_R2278_U265 , P1_R2278_U266 , P1_R2278_U267;
wire P1_R2278_U268 , P1_R2278_U269 , P1_R2278_U270 , P1_R2278_U271 , P1_R2278_U272 , P1_R2278_U273 , P1_R2278_U274 , P1_R2278_U275 , P1_R2278_U276 , P1_R2278_U277;
wire P1_R2278_U278 , P1_R2278_U279 , P1_R2278_U280 , P1_R2278_U281 , P1_R2278_U282 , P1_R2278_U283 , P1_R2278_U284 , P1_R2278_U285 , P1_R2278_U286 , P1_R2278_U287;
wire P1_R2278_U288 , P1_R2278_U289 , P1_R2278_U290 , P1_R2278_U291 , P1_R2278_U292 , P1_R2278_U293 , P1_R2278_U294 , P1_R2278_U295 , P1_R2278_U296 , P1_R2278_U297;
wire P1_R2278_U298 , P1_R2278_U299 , P1_R2278_U300 , P1_R2278_U301 , P1_R2278_U302 , P1_R2278_U303 , P1_R2278_U304 , P1_R2278_U305 , P1_R2278_U306 , P1_R2278_U307;
wire P1_R2278_U308 , P1_R2278_U309 , P1_R2278_U310 , P1_R2278_U311 , P1_R2278_U312 , P1_R2278_U313 , P1_R2278_U314 , P1_R2278_U315 , P1_R2278_U316 , P1_R2278_U317;
wire P1_R2278_U318 , P1_R2278_U319 , P1_R2278_U320 , P1_R2278_U321 , P1_R2278_U322 , P1_R2278_U323 , P1_R2278_U324 , P1_R2278_U325 , P1_R2278_U326 , P1_R2278_U327;
wire P1_R2278_U328 , P1_R2278_U329 , P1_R2278_U330 , P1_R2278_U331 , P1_R2278_U332 , P1_R2278_U333 , P1_R2278_U334 , P1_R2278_U335 , P1_R2278_U336 , P1_R2278_U337;
wire P1_R2278_U338 , P1_R2278_U339 , P1_R2278_U340 , P1_R2278_U341 , P1_R2278_U342 , P1_R2278_U343 , P1_R2278_U344 , P1_R2278_U345 , P1_R2278_U346 , P1_R2278_U347;
wire P1_R2278_U348 , P1_R2278_U349 , P1_R2278_U350 , P1_R2278_U351 , P1_R2278_U352 , P1_R2278_U353 , P1_R2278_U354 , P1_R2278_U355 , P1_R2278_U356 , P1_R2278_U357;
wire P1_R2278_U358 , P1_R2278_U359 , P1_R2278_U360 , P1_R2278_U361 , P1_R2278_U362 , P1_R2278_U363 , P1_R2278_U364 , P1_R2278_U365 , P1_R2278_U366 , P1_R2278_U367;
wire P1_R2278_U368 , P1_R2278_U369 , P1_R2278_U370 , P1_R2278_U371 , P1_R2278_U372 , P1_R2278_U373 , P1_R2278_U374 , P1_R2278_U375 , P1_R2278_U376 , P1_R2278_U377;
wire P1_R2278_U378 , P1_R2278_U379 , P1_R2278_U380 , P1_R2278_U381 , P1_R2278_U382 , P1_R2278_U383 , P1_R2278_U384 , P1_R2278_U385 , P1_R2278_U386 , P1_R2278_U387;
wire P1_R2278_U388 , P1_R2278_U389 , P1_R2278_U390 , P1_R2278_U391 , P1_R2278_U392 , P1_R2278_U393 , P1_R2278_U394 , P1_R2278_U395 , P1_R2278_U396 , P1_R2278_U397;
wire P1_R2278_U398 , P1_R2278_U399 , P1_R2278_U400 , P1_R2278_U401 , P1_R2278_U402 , P1_R2278_U403 , P1_R2278_U404 , P1_R2278_U405 , P1_R2278_U406 , P1_R2278_U407;
wire P1_R2278_U408 , P1_R2278_U409 , P1_R2278_U410 , P1_R2278_U411 , P1_R2278_U412 , P1_R2278_U413 , P1_R2278_U414 , P1_R2278_U415 , P1_R2278_U416 , P1_R2278_U417;
wire P1_R2278_U418 , P1_R2278_U419 , P1_R2278_U420 , P1_R2278_U421 , P1_R2278_U422 , P1_R2278_U423 , P1_R2278_U424 , P1_R2278_U425 , P1_R2278_U426 , P1_R2278_U427;
wire P1_R2278_U428 , P1_R2278_U429 , P1_R2278_U430 , P1_R2278_U431 , P1_R2278_U432 , P1_R2278_U433 , P1_R2278_U434 , P1_R2278_U435 , P1_R2278_U436 , P1_R2278_U437;
wire P1_R2278_U438 , P1_R2278_U439 , P1_R2278_U440 , P1_R2278_U441 , P1_R2278_U442 , P1_R2278_U443 , P1_R2278_U444 , P1_R2278_U445 , P1_R2278_U446 , P1_R2278_U447;
wire P1_R2278_U448 , P1_R2278_U449 , P1_R2278_U450 , P1_R2278_U451 , P1_R2278_U452 , P1_R2278_U453 , P1_R2278_U454 , P1_R2278_U455 , P1_R2278_U456 , P1_R2278_U457;
wire P1_R2278_U458 , P1_R2278_U459 , P1_R2278_U460 , P1_R2278_U461 , P1_R2278_U462 , P1_R2278_U463 , P1_R2278_U464 , P1_R2278_U465 , P1_R2278_U466 , P1_R2278_U467;
wire P1_R2278_U468 , P1_R2278_U469 , P1_R2278_U470 , P1_R2278_U471 , P1_R2278_U472 , P1_R2278_U473 , P1_R2278_U474 , P1_R2278_U475 , P1_R2278_U476 , P1_R2278_U477;
wire P1_R2278_U478 , P1_R2278_U479 , P1_R2278_U480 , P1_R2278_U481 , P1_R2278_U482 , P1_R2278_U483 , P1_R2278_U484 , P1_R2278_U485 , P1_R2278_U486 , P1_R2278_U487;
wire P1_R2278_U488 , P1_R2278_U489 , P1_R2278_U490 , P1_R2278_U491 , P1_R2278_U492 , P1_R2278_U493 , P1_R2278_U494 , P1_R2278_U495 , P1_R2278_U496 , P1_R2278_U497;
wire P1_R2278_U498 , P1_R2278_U499 , P1_R2278_U500 , P1_R2278_U501 , P1_R2278_U502 , P1_R2278_U503 , P1_R2278_U504 , P1_R2278_U505 , P1_R2278_U506 , P1_R2278_U507;
wire P1_R2278_U508 , P1_R2278_U509 , P1_R2278_U510 , P1_R2278_U511 , P1_R2278_U512 , P1_R2278_U513 , P1_R2278_U514 , P1_R2278_U515 , P1_R2278_U516 , P1_R2278_U517;
wire P1_R2278_U518 , P1_R2278_U519 , P1_R2278_U520 , P1_R2278_U521 , P1_R2278_U522 , P1_R2278_U523 , P1_R2278_U524 , P1_R2278_U525 , P1_R2278_U526 , P1_R2278_U527;
wire P1_R2278_U528 , P1_R2278_U529 , P1_R2278_U530 , P1_R2278_U531 , P1_R2278_U532 , P1_R2278_U533 , P1_R2278_U534 , P1_R2278_U535 , P1_R2278_U536 , P1_R2278_U537;
wire P1_R2278_U538 , P1_R2278_U539 , P1_R2278_U540 , P1_R2278_U541 , P1_R2278_U542 , P1_R2278_U543 , P1_R2278_U544 , P1_R2278_U545 , P1_R2278_U546 , P1_R2278_U547;
wire P1_R2278_U548 , P1_R2278_U549 , P1_R2278_U550 , P1_R2278_U551 , P1_R2278_U552 , P1_R2278_U553 , P1_R2278_U554 , P1_R2278_U555 , P1_R2278_U556 , P1_R2278_U557;
wire P1_R2278_U558 , P1_R2278_U559 , P1_R2278_U560 , P1_R2278_U561 , P1_R2278_U562 , P1_R2278_U563 , P1_R2278_U564 , P1_R2278_U565 , P1_R2278_U566 , P1_R2278_U567;
wire P1_R2278_U568 , P1_R2278_U569 , P1_R2278_U570 , P1_R2278_U571 , P1_R2278_U572 , P1_R2278_U573 , P1_R2278_U574 , P1_R2278_U575 , P1_R2278_U576 , P1_R2278_U577;
wire P1_R2278_U578 , P1_R2278_U579 , P1_R2278_U580 , P1_R2278_U581 , P1_R2278_U582 , P1_R2278_U583 , P1_R2278_U584 , P1_R2278_U585 , P1_R2278_U586 , P1_R2278_U587;
wire P1_R2278_U588 , P1_R2278_U589 , P1_R2278_U590 , P1_R2278_U591 , P1_R2278_U592 , P1_R2278_U593 , P1_R2278_U594 , P1_R2278_U595 , P1_R2278_U596 , P1_R2278_U597;
wire P1_R2278_U598 , P1_R2278_U599 , P1_R2278_U600 , P1_R2278_U601 , P1_R2278_U602 , P1_R2278_U603 , P1_R2278_U604 , P1_R2278_U605 , P1_R2278_U606 , P1_R2278_U607;
wire P1_R2278_U608 , P1_R2278_U609 , P1_R2278_U610 , P1_R2358_U5 , P1_R2358_U6 , P1_R2358_U7 , P1_R2358_U8 , P1_R2358_U9 , P1_R2358_U10 , P1_R2358_U11;
wire P1_R2358_U12 , P1_R2358_U13 , P1_R2358_U14 , P1_R2358_U15 , P1_R2358_U16 , P1_R2358_U17 , P1_R2358_U18 , P1_R2358_U19 , P1_R2358_U20 , P1_R2358_U21;
wire P1_R2358_U22 , P1_R2358_U23 , P1_R2358_U24 , P1_R2358_U25 , P1_R2358_U26 , P1_R2358_U27 , P1_R2358_U28 , P1_R2358_U29 , P1_R2358_U30 , P1_R2358_U31;
wire P1_R2358_U32 , P1_R2358_U33 , P1_R2358_U34 , P1_R2358_U35 , P1_R2358_U36 , P1_R2358_U37 , P1_R2358_U38 , P1_R2358_U39 , P1_R2358_U40 , P1_R2358_U41;
wire P1_R2358_U42 , P1_R2358_U43 , P1_R2358_U44 , P1_R2358_U45 , P1_R2358_U46 , P1_R2358_U47 , P1_R2358_U48 , P1_R2358_U49 , P1_R2358_U50 , P1_R2358_U51;
wire P1_R2358_U52 , P1_R2358_U53 , P1_R2358_U54 , P1_R2358_U55 , P1_R2358_U56 , P1_R2358_U57 , P1_R2358_U58 , P1_R2358_U59 , P1_R2358_U60 , P1_R2358_U61;
wire P1_R2358_U62 , P1_R2358_U63 , P1_R2358_U64 , P1_R2358_U65 , P1_R2358_U66 , P1_R2358_U67 , P1_R2358_U68 , P1_R2358_U69 , P1_R2358_U70 , P1_R2358_U71;
wire P1_R2358_U72 , P1_R2358_U73 , P1_R2358_U74 , P1_R2358_U75 , P1_R2358_U76 , P1_R2358_U77 , P1_R2358_U78 , P1_R2358_U79 , P1_R2358_U80 , P1_R2358_U81;
wire P1_R2358_U82 , P1_R2358_U83 , P1_R2358_U84 , P1_R2358_U85 , P1_R2358_U86 , P1_R2358_U87 , P1_R2358_U88 , P1_R2358_U89 , P1_R2358_U90 , P1_R2358_U91;
wire P1_R2358_U92 , P1_R2358_U93 , P1_R2358_U94 , P1_R2358_U95 , P1_R2358_U96 , P1_R2358_U97 , P1_R2358_U98 , P1_R2358_U99 , P1_R2358_U100 , P1_R2358_U101;
wire P1_R2358_U102 , P1_R2358_U103 , P1_R2358_U104 , P1_R2358_U105 , P1_R2358_U106 , P1_R2358_U107 , P1_R2358_U108 , P1_R2358_U109 , P1_R2358_U110 , P1_R2358_U111;
wire P1_R2358_U112 , P1_R2358_U113 , P1_R2358_U114 , P1_R2358_U115 , P1_R2358_U116 , P1_R2358_U117 , P1_R2358_U118 , P1_R2358_U119 , P1_R2358_U120 , P1_R2358_U121;
wire P1_R2358_U122 , P1_R2358_U123 , P1_R2358_U124 , P1_R2358_U125 , P1_R2358_U126 , P1_R2358_U127 , P1_R2358_U128 , P1_R2358_U129 , P1_R2358_U130 , P1_R2358_U131;
wire P1_R2358_U132 , P1_R2358_U133 , P1_R2358_U134 , P1_R2358_U135 , P1_R2358_U136 , P1_R2358_U137 , P1_R2358_U138 , P1_R2358_U139 , P1_R2358_U140 , P1_R2358_U141;
wire P1_R2358_U142 , P1_R2358_U143 , P1_R2358_U144 , P1_R2358_U145 , P1_R2358_U146 , P1_R2358_U147 , P1_R2358_U148 , P1_R2358_U149 , P1_R2358_U150 , P1_R2358_U151;
wire P1_R2358_U152 , P1_R2358_U153 , P1_R2358_U154 , P1_R2358_U155 , P1_R2358_U156 , P1_R2358_U157 , P1_R2358_U158 , P1_R2358_U159 , P1_R2358_U160 , P1_R2358_U161;
wire P1_R2358_U162 , P1_R2358_U163 , P1_R2358_U164 , P1_R2358_U165 , P1_R2358_U166 , P1_R2358_U167 , P1_R2358_U168 , P1_R2358_U169 , P1_R2358_U170 , P1_R2358_U171;
wire P1_R2358_U172 , P1_R2358_U173 , P1_R2358_U174 , P1_R2358_U175 , P1_R2358_U176 , P1_R2358_U177 , P1_R2358_U178 , P1_R2358_U179 , P1_R2358_U180 , P1_R2358_U181;
wire P1_R2358_U182 , P1_R2358_U183 , P1_R2358_U184 , P1_R2358_U185 , P1_R2358_U186 , P1_R2358_U187 , P1_R2358_U188 , P1_R2358_U189 , P1_R2358_U190 , P1_R2358_U191;
wire P1_R2358_U192 , P1_R2358_U193 , P1_R2358_U194 , P1_R2358_U195 , P1_R2358_U196 , P1_R2358_U197 , P1_R2358_U198 , P1_R2358_U199 , P1_R2358_U200 , P1_R2358_U201;
wire P1_R2358_U202 , P1_R2358_U203 , P1_R2358_U204 , P1_R2358_U205 , P1_R2358_U206 , P1_R2358_U207 , P1_R2358_U208 , P1_R2358_U209 , P1_R2358_U210 , P1_R2358_U211;
wire P1_R2358_U212 , P1_R2358_U213 , P1_R2358_U214 , P1_R2358_U215 , P1_R2358_U216 , P1_R2358_U217 , P1_R2358_U218 , P1_R2358_U219 , P1_R2358_U220 , P1_R2358_U221;
wire P1_R2358_U222 , P1_R2358_U223 , P1_R2358_U224 , P1_R2358_U225 , P1_R2358_U226 , P1_R2358_U227 , P1_R2358_U228 , P1_R2358_U229 , P1_R2358_U230 , P1_R2358_U231;
wire P1_R2358_U232 , P1_R2358_U233 , P1_R2358_U234 , P1_R2358_U235 , P1_R2358_U236 , P1_R2358_U237 , P1_R2358_U238 , P1_R2358_U239 , P1_R2358_U240 , P1_R2358_U241;
wire P1_R2358_U242 , P1_R2358_U243 , P1_R2358_U244 , P1_R2358_U245 , P1_R2358_U246 , P1_R2358_U247 , P1_R2358_U248 , P1_R2358_U249 , P1_R2358_U250 , P1_R2358_U251;
wire P1_R2358_U252 , P1_R2358_U253 , P1_R2358_U254 , P1_R2358_U255 , P1_R2358_U256 , P1_R2358_U257 , P1_R2358_U258 , P1_R2358_U259 , P1_R2358_U260 , P1_R2358_U261;
wire P1_R2358_U262 , P1_R2358_U263 , P1_R2358_U264 , P1_R2358_U265 , P1_R2358_U266 , P1_R2358_U267 , P1_R2358_U268 , P1_R2358_U269 , P1_R2358_U270 , P1_R2358_U271;
wire P1_R2358_U272 , P1_R2358_U273 , P1_R2358_U274 , P1_R2358_U275 , P1_R2358_U276 , P1_R2358_U277 , P1_R2358_U278 , P1_R2358_U279 , P1_R2358_U280 , P1_R2358_U281;
wire P1_R2358_U282 , P1_R2358_U283 , P1_R2358_U284 , P1_R2358_U285 , P1_R2358_U286 , P1_R2358_U287 , P1_R2358_U288 , P1_R2358_U289 , P1_R2358_U290 , P1_R2358_U291;
wire P1_R2358_U292 , P1_R2358_U293 , P1_R2358_U294 , P1_R2358_U295 , P1_R2358_U296 , P1_R2358_U297 , P1_R2358_U298 , P1_R2358_U299 , P1_R2358_U300 , P1_R2358_U301;
wire P1_R2358_U302 , P1_R2358_U303 , P1_R2358_U304 , P1_R2358_U305 , P1_R2358_U306 , P1_R2358_U307 , P1_R2358_U308 , P1_R2358_U309 , P1_R2358_U310 , P1_R2358_U311;
wire P1_R2358_U312 , P1_R2358_U313 , P1_R2358_U314 , P1_R2358_U315 , P1_R2358_U316 , P1_R2358_U317 , P1_R2358_U318 , P1_R2358_U319 , P1_R2358_U320 , P1_R2358_U321;
wire P1_R2358_U322 , P1_R2358_U323 , P1_R2358_U324 , P1_R2358_U325 , P1_R2358_U326 , P1_R2358_U327 , P1_R2358_U328 , P1_R2358_U329 , P1_R2358_U330 , P1_R2358_U331;
wire P1_R2358_U332 , P1_R2358_U333 , P1_R2358_U334 , P1_R2358_U335 , P1_R2358_U336 , P1_R2358_U337 , P1_R2358_U338 , P1_R2358_U339 , P1_R2358_U340 , P1_R2358_U341;
wire P1_R2358_U342 , P1_R2358_U343 , P1_R2358_U344 , P1_R2358_U345 , P1_R2358_U346 , P1_R2358_U347 , P1_R2358_U348 , P1_R2358_U349 , P1_R2358_U350 , P1_R2358_U351;
wire P1_R2358_U352 , P1_R2358_U353 , P1_R2358_U354 , P1_R2358_U355 , P1_R2358_U356 , P1_R2358_U357 , P1_R2358_U358 , P1_R2358_U359 , P1_R2358_U360 , P1_R2358_U361;
wire P1_R2358_U362 , P1_R2358_U363 , P1_R2358_U364 , P1_R2358_U365 , P1_R2358_U366 , P1_R2358_U367 , P1_R2358_U368 , P1_R2358_U369 , P1_R2358_U370 , P1_R2358_U371;
wire P1_R2358_U372 , P1_R2358_U373 , P1_R2358_U374 , P1_R2358_U375 , P1_R2358_U376 , P1_R2358_U377 , P1_R2358_U378 , P1_R2358_U379 , P1_R2358_U380 , P1_R2358_U381;
wire P1_R2358_U382 , P1_R2358_U383 , P1_R2358_U384 , P1_R2358_U385 , P1_R2358_U386 , P1_R2358_U387 , P1_R2358_U388 , P1_R2358_U389 , P1_R2358_U390 , P1_R2358_U391;
wire P1_R2358_U392 , P1_R2358_U393 , P1_R2358_U394 , P1_R2358_U395 , P1_R2358_U396 , P1_R2358_U397 , P1_R2358_U398 , P1_R2358_U399 , P1_R2358_U400 , P1_R2358_U401;
wire P1_R2358_U402 , P1_R2358_U403 , P1_R2358_U404 , P1_R2358_U405 , P1_R2358_U406 , P1_R2358_U407 , P1_R2358_U408 , P1_R2358_U409 , P1_R2358_U410 , P1_R2358_U411;
wire P1_R2358_U412 , P1_R2358_U413 , P1_R2358_U414 , P1_R2358_U415 , P1_R2358_U416 , P1_R2358_U417 , P1_R2358_U418 , P1_R2358_U419 , P1_R2358_U420 , P1_R2358_U421;
wire P1_R2358_U422 , P1_R2358_U423 , P1_R2358_U424 , P1_R2358_U425 , P1_R2358_U426 , P1_R2358_U427 , P1_R2358_U428 , P1_R2358_U429 , P1_R2358_U430 , P1_R2358_U431;
wire P1_R2358_U432 , P1_R2358_U433 , P1_R2358_U434 , P1_R2358_U435 , P1_R2358_U436 , P1_R2358_U437 , P1_R2358_U438 , P1_R2358_U439 , P1_R2358_U440 , P1_R2358_U441;
wire P1_R2358_U442 , P1_R2358_U443 , P1_R2358_U444 , P1_R2358_U445 , P1_R2358_U446 , P1_R2358_U447 , P1_R2358_U448 , P1_R2358_U449 , P1_R2358_U450 , P1_R2358_U451;
wire P1_R2358_U452 , P1_R2358_U453 , P1_R2358_U454 , P1_R2358_U455 , P1_R2358_U456 , P1_R2358_U457 , P1_R2358_U458 , P1_R2358_U459 , P1_R2358_U460 , P1_R2358_U461;
wire P1_R2358_U462 , P1_R2358_U463 , P1_R2358_U464 , P1_R2358_U465 , P1_R2358_U466 , P1_R2358_U467 , P1_R2358_U468 , P1_R2358_U469 , P1_R2358_U470 , P1_R2358_U471;
wire P1_R2358_U472 , P1_R2358_U473 , P1_R2358_U474 , P1_R2358_U475 , P1_R2358_U476 , P1_R2358_U477 , P1_R2358_U478 , P1_R2358_U479 , P1_R2358_U480 , P1_R2358_U481;
wire P1_R2358_U482 , P1_R2358_U483 , P1_R2358_U484 , P1_R2358_U485 , P1_R2358_U486 , P1_R2358_U487 , P1_R2358_U488 , P1_R2358_U489 , P1_R2358_U490 , P1_R2358_U491;
wire P1_R2358_U492 , P1_R2358_U493 , P1_R2358_U494 , P1_R2358_U495 , P1_R2358_U496 , P1_R2358_U497 , P1_R2358_U498 , P1_R2358_U499 , P1_R2358_U500 , P1_R2358_U501;
wire P1_R2358_U502 , P1_R2358_U503 , P1_R2358_U504 , P1_R2358_U505 , P1_R2358_U506 , P1_R2358_U507 , P1_R2358_U508 , P1_R2358_U509 , P1_R2358_U510 , P1_R2358_U511;
wire P1_R2358_U512 , P1_R2358_U513 , P1_R2358_U514 , P1_R2358_U515 , P1_R2358_U516 , P1_R2358_U517 , P1_R2358_U518 , P1_R2358_U519 , P1_R2358_U520 , P1_R2358_U521;
wire P1_R2358_U522 , P1_R2358_U523 , P1_R2358_U524 , P1_R2358_U525 , P1_R2358_U526 , P1_R2358_U527 , P1_R2358_U528 , P1_R2358_U529 , P1_R2358_U530 , P1_R2358_U531;
wire P1_R2358_U532 , P1_R2358_U533 , P1_R2358_U534 , P1_R2358_U535 , P1_R2358_U536 , P1_R2358_U537 , P1_R2358_U538 , P1_R2358_U539 , P1_R2358_U540 , P1_R2358_U541;
wire P1_R2358_U542 , P1_R2358_U543 , P1_R2358_U544 , P1_R2358_U545 , P1_R2358_U546 , P1_R2358_U547 , P1_R2358_U548 , P1_R2358_U549 , P1_R2358_U550 , P1_R2358_U551;
wire P1_R2358_U552 , P1_R2358_U553 , P1_R2358_U554 , P1_R2358_U555 , P1_R2358_U556 , P1_R2358_U557 , P1_R2358_U558 , P1_R2358_U559 , P1_R2358_U560 , P1_R2358_U561;
wire P1_R2358_U562 , P1_R2358_U563 , P1_R2358_U564 , P1_R2358_U565 , P1_R2358_U566 , P1_R2358_U567 , P1_R2358_U568 , P1_R2358_U569 , P1_R2358_U570 , P1_R2358_U571;
wire P1_R2358_U572 , P1_R2358_U573 , P1_R2358_U574 , P1_R2358_U575 , P1_R2358_U576 , P1_R2358_U577 , P1_R2358_U578 , P1_R2358_U579 , P1_R2358_U580 , P1_R2358_U581;
wire P1_R2358_U582 , P1_R2358_U583 , P1_R2358_U584 , P1_R2358_U585 , P1_R2358_U586 , P1_R2358_U587 , P1_R2358_U588 , P1_R2358_U589 , P1_R2358_U590 , P1_R2358_U591;
wire P1_R2358_U592 , P1_R2358_U593 , P1_R2358_U594 , P1_R2358_U595 , P1_R2358_U596 , P1_R2358_U597 , P1_R2358_U598 , P1_R2358_U599 , P1_R2358_U600 , P1_R2358_U601;
wire P1_R2358_U602 , P1_R2358_U603 , P1_R2358_U604 , P1_R2358_U605 , P1_R2358_U606 , P1_R2358_U607 , P1_R2358_U608 , P1_R2358_U609 , P1_R2358_U610 , P1_R2358_U611;
wire P1_LT_589_U6 , P1_LT_589_U7 , P1_LT_589_U8 , P1_R584_U6 , P1_R584_U7 , P1_R584_U8 , P1_R584_U9 , P1_R2099_U4 , P1_R2099_U5 , P1_R2099_U6;
wire P1_R2099_U7 , P1_R2099_U8 , P1_R2099_U9 , P1_R2099_U10 , P1_R2099_U11 , P1_R2099_U12 , P1_R2099_U13 , P1_R2099_U14 , P1_R2099_U15 , P1_R2099_U16;
wire P1_R2099_U17 , P1_R2099_U18 , P1_R2099_U19 , P1_R2099_U20 , P1_R2099_U21 , P1_R2099_U22 , P1_R2099_U23 , P1_R2099_U24 , P1_R2099_U25 , P1_R2099_U26;
wire P1_R2099_U27 , P1_R2099_U28 , P1_R2099_U29 , P1_R2099_U30 , P1_R2099_U31 , P1_R2099_U32 , P1_R2099_U33 , P1_R2099_U34 , P1_R2099_U35 , P1_R2099_U36;
wire P1_R2099_U37 , P1_R2099_U38 , P1_R2099_U39 , P1_R2099_U40 , P1_R2099_U41 , P1_R2099_U42 , P1_R2099_U43 , P1_R2099_U44 , P1_R2099_U45 , P1_R2099_U46;
wire P1_R2099_U47 , P1_R2099_U48 , P1_R2099_U49 , P1_R2099_U50 , P1_R2099_U51 , P1_R2099_U52 , P1_R2099_U53 , P1_R2099_U54 , P1_R2099_U55 , P1_R2099_U56;
wire P1_R2099_U57 , P1_R2099_U58 , P1_R2099_U59 , P1_R2099_U60 , P1_R2099_U61 , P1_R2099_U62 , P1_R2099_U63 , P1_R2099_U64 , P1_R2099_U65 , P1_R2099_U66;
wire P1_R2099_U67 , P1_R2099_U68 , P1_R2099_U69 , P1_R2099_U70 , P1_R2099_U71 , P1_R2099_U72 , P1_R2099_U73 , P1_R2099_U74 , P1_R2099_U75 , P1_R2099_U76;
wire P1_R2099_U77 , P1_R2099_U78 , P1_R2099_U79 , P1_R2099_U80 , P1_R2099_U81 , P1_R2099_U82 , P1_R2099_U83 , P1_R2099_U84 , P1_R2099_U85 , P1_R2099_U86;
wire P1_R2099_U87 , P1_R2099_U88 , P1_R2099_U89 , P1_R2099_U90 , P1_R2099_U91 , P1_R2099_U92 , P1_R2099_U93 , P1_R2099_U94 , P1_R2099_U95 , P1_R2099_U96;
wire P1_R2099_U97 , P1_R2099_U98 , P1_R2099_U99 , P1_R2099_U100 , P1_R2099_U101 , P1_R2099_U102 , P1_R2099_U103 , P1_R2099_U104 , P1_R2099_U105 , P1_R2099_U106;
wire P1_R2099_U107 , P1_R2099_U108 , P1_R2099_U109 , P1_R2099_U110 , P1_R2099_U111 , P1_R2099_U112 , P1_R2099_U113 , P1_R2099_U114 , P1_R2099_U115 , P1_R2099_U116;
wire P1_R2099_U117 , P1_R2099_U118 , P1_R2099_U119 , P1_R2099_U120 , P1_R2099_U121 , P1_R2099_U122 , P1_R2099_U123 , P1_R2099_U124 , P1_R2099_U125 , P1_R2099_U126;
wire P1_R2099_U127 , P1_R2099_U128 , P1_R2099_U129 , P1_R2099_U130 , P1_R2099_U131 , P1_R2099_U132 , P1_R2099_U133 , P1_R2099_U134 , P1_R2099_U135 , P1_R2099_U136;
wire P1_R2099_U137 , P1_R2099_U138 , P1_R2099_U139 , P1_R2099_U140 , P1_R2099_U141 , P1_R2099_U142 , P1_R2099_U143 , P1_R2099_U144 , P1_R2099_U145 , P1_R2099_U146;
wire P1_R2099_U147 , P1_R2099_U148 , P1_R2099_U149 , P1_R2099_U150 , P1_R2099_U151 , P1_R2099_U152 , P1_R2099_U153 , P1_R2099_U154 , P1_R2099_U155 , P1_R2099_U156;
wire P1_R2099_U157 , P1_R2099_U158 , P1_R2099_U159 , P1_R2099_U160 , P1_R2099_U161 , P1_R2099_U162 , P1_R2099_U163 , P1_R2099_U164 , P1_R2099_U165 , P1_R2099_U166;
wire P1_R2099_U167 , P1_R2099_U168 , P1_R2099_U169 , P1_R2099_U170 , P1_R2099_U171 , P1_R2099_U172 , P1_R2099_U173 , P1_R2099_U174 , P1_R2099_U175 , P1_R2099_U176;
wire P1_R2099_U177 , P1_R2099_U178 , P1_R2099_U179 , P1_R2099_U180 , P1_R2099_U181 , P1_R2099_U182 , P1_R2099_U183 , P1_R2099_U184 , P1_R2099_U185 , P1_R2099_U186;
wire P1_R2099_U187 , P1_R2099_U188 , P1_R2099_U189 , P1_R2099_U190 , P1_R2099_U191 , P1_R2099_U192 , P1_R2099_U193 , P1_R2099_U194 , P1_R2099_U195 , P1_R2099_U196;
wire P1_R2099_U197 , P1_R2099_U198 , P1_R2099_U199 , P1_R2099_U200 , P1_R2099_U201 , P1_R2099_U202 , P1_R2099_U203 , P1_R2099_U204 , P1_R2099_U205 , P1_R2099_U206;
wire P1_R2099_U207 , P1_R2099_U208 , P1_R2099_U209 , P1_R2099_U210 , P1_R2099_U211 , P1_R2099_U212 , P1_R2099_U213 , P1_R2099_U214 , P1_R2099_U215 , P1_R2099_U216;
wire P1_R2099_U217 , P1_R2099_U218 , P1_R2099_U219 , P1_R2099_U220 , P1_R2099_U221 , P1_R2099_U222 , P1_R2099_U223 , P1_R2099_U224 , P1_R2099_U225 , P1_R2099_U226;
wire P1_R2099_U227 , P1_R2099_U228 , P1_R2099_U229 , P1_R2099_U230 , P1_R2099_U231 , P1_R2099_U232 , P1_R2099_U233 , P1_R2099_U234 , P1_R2099_U235 , P1_R2099_U236;
wire P1_R2099_U237 , P1_R2099_U238 , P1_R2099_U239 , P1_R2099_U240 , P1_R2099_U241 , P1_R2099_U242 , P1_R2099_U243 , P1_R2099_U244 , P1_R2099_U245 , P1_R2099_U246;
wire P1_R2099_U247 , P1_R2099_U248 , P1_R2099_U249 , P1_R2099_U250 , P1_R2099_U251 , P1_R2099_U252 , P1_R2099_U253 , P1_R2099_U254 , P1_R2099_U255 , P1_R2099_U256;
wire P1_R2099_U257 , P1_R2099_U258 , P1_R2099_U259 , P1_R2099_U260 , P1_R2099_U261 , P1_R2099_U262 , P1_R2099_U263 , P1_R2099_U264 , P1_R2099_U265 , P1_R2099_U266;
wire P1_R2099_U267 , P1_R2099_U268 , P1_R2099_U269 , P1_R2099_U270 , P1_R2099_U271 , P1_R2099_U272 , P1_R2099_U273 , P1_R2099_U274 , P1_R2099_U275 , P1_R2099_U276;
wire P1_R2099_U277 , P1_R2099_U278 , P1_R2099_U279 , P1_R2099_U280 , P1_R2099_U281 , P1_R2099_U282 , P1_R2099_U283 , P1_R2099_U284 , P1_R2099_U285 , P1_R2099_U286;
wire P1_R2099_U287 , P1_R2099_U288 , P1_R2099_U289 , P1_R2099_U290 , P1_R2099_U291 , P1_R2099_U292 , P1_R2099_U293 , P1_R2099_U294 , P1_R2099_U295 , P1_R2099_U296;
wire P1_R2099_U297 , P1_R2099_U298 , P1_R2099_U299 , P1_R2099_U300 , P1_R2099_U301 , P1_R2099_U302 , P1_R2099_U303 , P1_R2099_U304 , P1_R2099_U305 , P1_R2099_U306;
wire P1_R2099_U307 , P1_R2099_U308 , P1_R2099_U309 , P1_R2099_U310 , P1_R2099_U311 , P1_R2099_U312 , P1_R2099_U313 , P1_R2099_U314 , P1_R2099_U315 , P1_R2099_U316;
wire P1_R2099_U317 , P1_R2099_U318 , P1_R2099_U319 , P1_R2099_U320 , P1_R2099_U321 , P1_R2099_U322 , P1_R2099_U323 , P1_R2099_U324 , P1_R2099_U325 , P1_R2099_U326;
wire P1_R2099_U327 , P1_R2099_U328 , P1_R2099_U329 , P1_R2099_U330 , P1_R2099_U331 , P1_R2099_U332 , P1_R2099_U333 , P1_R2099_U334 , P1_R2099_U335 , P1_R2099_U336;
wire P1_R2099_U337 , P1_R2099_U338 , P1_R2099_U339 , P1_R2099_U340 , P1_R2099_U341 , P1_R2099_U342 , P1_R2099_U343 , P1_R2099_U344 , P1_R2099_U345 , P1_R2099_U346;
wire P1_R2099_U347 , P1_R2099_U348 , P1_R2099_U349 , P1_R2167_U6 , P1_R2167_U7 , P1_R2167_U8 , P1_R2167_U9 , P1_R2167_U10 , P1_R2167_U11 , P1_R2167_U12;
wire P1_R2167_U13 , P1_R2167_U14 , P1_R2167_U15 , P1_R2167_U16 , P1_R2167_U17 , P1_R2167_U18 , P1_R2167_U19 , P1_R2167_U20 , P1_R2167_U21 , P1_R2167_U22;
wire P1_R2167_U23 , P1_R2167_U24 , P1_R2167_U25 , P1_R2167_U26 , P1_R2167_U27 , P1_R2167_U28 , P1_R2167_U29 , P1_R2167_U30 , P1_R2167_U31 , P1_R2167_U32;
wire P1_R2167_U33 , P1_R2167_U34 , P1_R2167_U35 , P1_R2167_U36 , P1_R2167_U37 , P1_R2167_U38 , P1_R2167_U39 , P1_R2167_U40 , P1_R2167_U41 , P1_R2167_U42;
wire P1_R2167_U43 , P1_R2167_U44 , P1_R2167_U45 , P1_R2167_U46 , P1_R2167_U47 , P1_R2167_U48 , P1_R2167_U49 , P1_R2167_U50 , P1_R2337_U4 , P1_R2337_U5;
wire P1_R2337_U6 , P1_R2337_U7 , P1_R2337_U8 , P1_R2337_U9 , P1_R2337_U10 , P1_R2337_U11 , P1_R2337_U12 , P1_R2337_U13 , P1_R2337_U14 , P1_R2337_U15;
wire P1_R2337_U16 , P1_R2337_U17 , P1_R2337_U18 , P1_R2337_U19 , P1_R2337_U20 , P1_R2337_U21 , P1_R2337_U22 , P1_R2337_U23 , P1_R2337_U24 , P1_R2337_U25;
wire P1_R2337_U26 , P1_R2337_U27 , P1_R2337_U28 , P1_R2337_U29 , P1_R2337_U30 , P1_R2337_U31 , P1_R2337_U32 , P1_R2337_U33 , P1_R2337_U34 , P1_R2337_U35;
wire P1_R2337_U36 , P1_R2337_U37 , P1_R2337_U38 , P1_R2337_U39 , P1_R2337_U40 , P1_R2337_U41 , P1_R2337_U42 , P1_R2337_U43 , P1_R2337_U44 , P1_R2337_U45;
wire P1_R2337_U46 , P1_R2337_U47 , P1_R2337_U48 , P1_R2337_U49 , P1_R2337_U50 , P1_R2337_U51 , P1_R2337_U52 , P1_R2337_U53 , P1_R2337_U54 , P1_R2337_U55;
wire P1_R2337_U56 , P1_R2337_U57 , P1_R2337_U58 , P1_R2337_U59 , P1_R2337_U60 , P1_R2337_U61 , P1_R2337_U62 , P1_R2337_U63 , P1_R2337_U64 , P1_R2337_U65;
wire P1_R2337_U66 , P1_R2337_U67 , P1_R2337_U68 , P1_R2337_U69 , P1_R2337_U70 , P1_R2337_U71 , P1_R2337_U72 , P1_R2337_U73 , P1_R2337_U74 , P1_R2337_U75;
wire P1_R2337_U76 , P1_R2337_U77 , P1_R2337_U78 , P1_R2337_U79 , P1_R2337_U80 , P1_R2337_U81 , P1_R2337_U82 , P1_R2337_U83 , P1_R2337_U84 , P1_R2337_U85;
wire P1_R2337_U86 , P1_R2337_U87 , P1_R2337_U88 , P1_R2337_U89 , P1_R2337_U90 , P1_R2337_U91 , P1_R2337_U92 , P1_R2337_U93 , P1_R2337_U94 , P1_R2337_U95;
wire P1_R2337_U96 , P1_R2337_U97 , P1_R2337_U98 , P1_R2337_U99 , P1_R2337_U100 , P1_R2337_U101 , P1_R2337_U102 , P1_R2337_U103 , P1_R2337_U104 , P1_R2337_U105;
wire P1_R2337_U106 , P1_R2337_U107 , P1_R2337_U108 , P1_R2337_U109 , P1_R2337_U110 , P1_R2337_U111 , P1_R2337_U112 , P1_R2337_U113 , P1_R2337_U114 , P1_R2337_U115;
wire P1_R2337_U116 , P1_R2337_U117 , P1_R2337_U118 , P1_R2337_U119 , P1_R2337_U120 , P1_R2337_U121 , P1_R2337_U122 , P1_R2337_U123 , P1_R2337_U124 , P1_R2337_U125;
wire P1_R2337_U126 , P1_R2337_U127 , P1_R2337_U128 , P1_R2337_U129 , P1_R2337_U130 , P1_R2337_U131 , P1_R2337_U132 , P1_R2337_U133 , P1_R2337_U134 , P1_R2337_U135;
wire P1_R2337_U136 , P1_R2337_U137 , P1_R2337_U138 , P1_R2337_U139 , P1_R2337_U140 , P1_R2337_U141 , P1_R2337_U142 , P1_R2337_U143 , P1_R2337_U144 , P1_R2337_U145;
wire P1_R2337_U146 , P1_R2337_U147 , P1_R2337_U148 , P1_R2337_U149 , P1_R2337_U150 , P1_R2337_U151 , P1_R2337_U152 , P1_R2337_U153 , P1_R2337_U154 , P1_R2337_U155;
wire P1_R2337_U156 , P1_R2337_U157 , P1_R2337_U158 , P1_R2337_U159 , P1_R2337_U160 , P1_R2337_U161 , P1_R2337_U162 , P1_R2337_U163 , P1_R2337_U164 , P1_R2337_U165;
wire P1_R2337_U166 , P1_R2337_U167 , P1_R2337_U168 , P1_R2337_U169 , P1_R2337_U170 , P1_R2337_U171 , P1_R2337_U172 , P1_R2337_U173 , P1_R2337_U174 , P1_R2337_U175;
wire P1_R2337_U176 , P1_R2337_U177 , P1_R2337_U178 , P1_R2337_U179 , P1_R2337_U180 , P1_R2337_U181 , P1_R2337_U182 , P1_SUB_357_U6 , P1_SUB_357_U7 , P1_SUB_357_U8;
wire P1_SUB_357_U9 , P1_SUB_357_U10 , P1_SUB_357_U11 , P1_SUB_357_U12 , P1_SUB_357_U13 , P1_LT_563_1260_U6 , P1_LT_563_1260_U7 , P1_LT_563_1260_U8 , P1_LT_563_1260_U9 , P1_SUB_580_U6;
wire P1_SUB_580_U7 , P1_SUB_580_U8 , P1_SUB_580_U9 , P1_SUB_580_U10 , P1_R2096_U4 , P1_R2096_U5 , P1_R2096_U6 , P1_R2096_U7 , P1_R2096_U8 , P1_R2096_U9;
wire P1_R2096_U10 , P1_R2096_U11 , P1_R2096_U12 , P1_R2096_U13 , P1_R2096_U14 , P1_R2096_U15 , P1_R2096_U16 , P1_R2096_U17 , P1_R2096_U18 , P1_R2096_U19;
wire P1_R2096_U20 , P1_R2096_U21 , P1_R2096_U22 , P1_R2096_U23 , P1_R2096_U24 , P1_R2096_U25 , P1_R2096_U26 , P1_R2096_U27 , P1_R2096_U28 , P1_R2096_U29;
wire P1_R2096_U30 , P1_R2096_U31 , P1_R2096_U32 , P1_R2096_U33 , P1_R2096_U34 , P1_R2096_U35 , P1_R2096_U36 , P1_R2096_U37 , P1_R2096_U38 , P1_R2096_U39;
wire P1_R2096_U40 , P1_R2096_U41 , P1_R2096_U42 , P1_R2096_U43 , P1_R2096_U44 , P1_R2096_U45 , P1_R2096_U46 , P1_R2096_U47 , P1_R2096_U48 , P1_R2096_U49;
wire P1_R2096_U50 , P1_R2096_U51 , P1_R2096_U52 , P1_R2096_U53 , P1_R2096_U54 , P1_R2096_U55 , P1_R2096_U56 , P1_R2096_U57 , P1_R2096_U58 , P1_R2096_U59;
wire P1_R2096_U60 , P1_R2096_U61 , P1_R2096_U62 , P1_R2096_U63 , P1_R2096_U64 , P1_R2096_U65 , P1_R2096_U66 , P1_R2096_U67 , P1_R2096_U68 , P1_R2096_U69;
wire P1_R2096_U70 , P1_R2096_U71 , P1_R2096_U72 , P1_R2096_U73 , P1_R2096_U74 , P1_R2096_U75 , P1_R2096_U76 , P1_R2096_U77 , P1_R2096_U78 , P1_R2096_U79;
wire P1_R2096_U80 , P1_R2096_U81 , P1_R2096_U82 , P1_R2096_U83 , P1_R2096_U84 , P1_R2096_U85 , P1_R2096_U86 , P1_R2096_U87 , P1_R2096_U88 , P1_R2096_U89;
wire P1_R2096_U90 , P1_R2096_U91 , P1_R2096_U92 , P1_R2096_U93 , P1_R2096_U94 , P1_R2096_U95 , P1_R2096_U96 , P1_R2096_U97 , P1_R2096_U98 , P1_R2096_U99;
wire P1_R2096_U100 , P1_R2096_U101 , P1_R2096_U102 , P1_R2096_U103 , P1_R2096_U104 , P1_R2096_U105 , P1_R2096_U106 , P1_R2096_U107 , P1_R2096_U108 , P1_R2096_U109;
wire P1_R2096_U110 , P1_R2096_U111 , P1_R2096_U112 , P1_R2096_U113 , P1_R2096_U114 , P1_R2096_U115 , P1_R2096_U116 , P1_R2096_U117 , P1_R2096_U118 , P1_R2096_U119;
wire P1_R2096_U120 , P1_R2096_U121 , P1_R2096_U122 , P1_R2096_U123 , P1_R2096_U124 , P1_R2096_U125 , P1_R2096_U126 , P1_R2096_U127 , P1_R2096_U128 , P1_R2096_U129;
wire P1_R2096_U130 , P1_R2096_U131 , P1_R2096_U132 , P1_R2096_U133 , P1_R2096_U134 , P1_R2096_U135 , P1_R2096_U136 , P1_R2096_U137 , P1_R2096_U138 , P1_R2096_U139;
wire P1_R2096_U140 , P1_R2096_U141 , P1_R2096_U142 , P1_R2096_U143 , P1_R2096_U144 , P1_R2096_U145 , P1_R2096_U146 , P1_R2096_U147 , P1_R2096_U148 , P1_R2096_U149;
wire P1_R2096_U150 , P1_R2096_U151 , P1_R2096_U152 , P1_R2096_U153 , P1_R2096_U154 , P1_R2096_U155 , P1_R2096_U156 , P1_R2096_U157 , P1_R2096_U158 , P1_R2096_U159;
wire P1_R2096_U160 , P1_R2096_U161 , P1_R2096_U162 , P1_R2096_U163 , P1_R2096_U164 , P1_R2096_U165 , P1_R2096_U166 , P1_R2096_U167 , P1_R2096_U168 , P1_R2096_U169;
wire P1_R2096_U170 , P1_R2096_U171 , P1_R2096_U172 , P1_R2096_U173 , P1_R2096_U174 , P1_R2096_U175 , P1_R2096_U176 , P1_R2096_U177 , P1_R2096_U178 , P1_R2096_U179;
wire P1_R2096_U180 , P1_R2096_U181 , P1_R2096_U182 , P1_LT_563_U6 , P1_LT_563_U7 , P1_LT_563_U8 , P1_LT_563_U9 , P1_LT_563_U10 , P1_LT_563_U11 , P1_LT_563_U12;
wire P1_LT_563_U13 , P1_LT_563_U14 , P1_LT_563_U15 , P1_LT_563_U16 , P1_LT_563_U17 , P1_LT_563_U18 , P1_LT_563_U19 , P1_LT_563_U20 , P1_LT_563_U21 , P1_LT_563_U22;
wire P1_LT_563_U23 , P1_LT_563_U24 , P1_LT_563_U25 , P1_LT_563_U26 , P1_LT_563_U27 , P1_LT_563_U28 , P1_R2238_U6 , P1_R2238_U7 , P1_R2238_U8 , P1_R2238_U9;
wire P1_R2238_U10 , P1_R2238_U11 , P1_R2238_U12 , P1_R2238_U13 , P1_R2238_U14 , P1_R2238_U15 , P1_R2238_U16 , P1_R2238_U17 , P1_R2238_U18 , P1_R2238_U19;
wire P1_R2238_U20 , P1_R2238_U21 , P1_R2238_U22 , P1_R2238_U23 , P1_R2238_U24 , P1_R2238_U25 , P1_R2238_U26 , P1_R2238_U27 , P1_R2238_U28 , P1_R2238_U29;
wire P1_R2238_U30 , P1_R2238_U31 , P1_R2238_U32 , P1_R2238_U33 , P1_R2238_U34 , P1_R2238_U35 , P1_R2238_U36 , P1_R2238_U37 , P1_R2238_U38 , P1_R2238_U39;
wire P1_R2238_U40 , P1_R2238_U41 , P1_R2238_U42 , P1_R2238_U43 , P1_R2238_U44 , P1_R2238_U45 , P1_R2238_U46 , P1_R2238_U47 , P1_R2238_U48 , P1_R2238_U49;
wire P1_R2238_U50 , P1_R2238_U51 , P1_R2238_U52 , P1_R2238_U53 , P1_R2238_U54 , P1_R2238_U55 , P1_R2238_U56 , P1_R2238_U57 , P1_R2238_U58 , P1_R2238_U59;
wire P1_R2238_U60 , P1_R2238_U61 , P1_R2238_U62 , P1_R2238_U63 , P1_R2238_U64 , P1_R2238_U65 , P1_R2238_U66 , P1_SUB_450_U6 , P1_SUB_450_U7 , P1_SUB_450_U8;
wire P1_SUB_450_U9 , P1_SUB_450_U10 , P1_SUB_450_U11 , P1_SUB_450_U12 , P1_SUB_450_U13 , P1_SUB_450_U14 , P1_SUB_450_U15 , P1_SUB_450_U16 , P1_SUB_450_U17 , P1_SUB_450_U18;
wire P1_SUB_450_U19 , P1_SUB_450_U20 , P1_SUB_450_U21 , P1_SUB_450_U22 , P1_SUB_450_U23 , P1_SUB_450_U24 , P1_SUB_450_U25 , P1_SUB_450_U26 , P1_SUB_450_U27 , P1_SUB_450_U28;
wire P1_SUB_450_U29 , P1_SUB_450_U30 , P1_SUB_450_U31 , P1_SUB_450_U32 , P1_SUB_450_U33 , P1_SUB_450_U34 , P1_SUB_450_U35 , P1_SUB_450_U36 , P1_SUB_450_U37 , P1_SUB_450_U38;
wire P1_SUB_450_U39 , P1_SUB_450_U40 , P1_SUB_450_U41 , P1_SUB_450_U42 , P1_SUB_450_U43 , P1_SUB_450_U44 , P1_SUB_450_U45 , P1_SUB_450_U46 , P1_SUB_450_U47 , P1_SUB_450_U48;
wire P1_SUB_450_U49 , P1_SUB_450_U50 , P1_SUB_450_U51 , P1_SUB_450_U52 , P1_SUB_450_U53 , P1_SUB_450_U54 , P1_SUB_450_U55 , P1_SUB_450_U56 , P1_SUB_450_U57 , P1_SUB_450_U58;
wire P1_SUB_450_U59 , P1_SUB_450_U60 , P1_SUB_450_U61 , P1_SUB_450_U62 , P1_SUB_450_U63 , P1_SUB_450_U64 , P1_SUB_450_U65 , P1_SUB_450_U66 , P1_ADD_371_U4 , P1_ADD_371_U5;
wire P1_ADD_371_U6 , P1_ADD_371_U7 , P1_ADD_371_U8 , P1_ADD_371_U9 , P1_ADD_371_U10 , P1_ADD_371_U11 , P1_ADD_371_U12 , P1_ADD_371_U13 , P1_ADD_371_U14 , P1_ADD_371_U15;
wire P1_ADD_371_U16 , P1_ADD_371_U17 , P1_ADD_371_U18 , P1_ADD_371_U19 , P1_ADD_371_U20 , P1_ADD_371_U21 , P1_ADD_371_U22 , P1_ADD_371_U23 , P1_ADD_371_U24 , P1_ADD_371_U25;
wire P1_ADD_371_U26 , P1_ADD_371_U27 , P1_ADD_371_U28 , P1_ADD_371_U29 , P1_ADD_371_U30 , P1_ADD_371_U31 , P1_ADD_371_U32 , P1_ADD_371_U33 , P1_ADD_371_U34 , P1_ADD_371_U35;
wire P1_ADD_371_U36 , P1_ADD_371_U37 , P1_ADD_371_U38 , P1_ADD_371_U39 , P1_ADD_371_U40 , P1_ADD_371_U41 , P1_ADD_371_U42 , P1_ADD_371_U43 , P1_ADD_371_U44 , P1_ADD_405_U4;
wire P1_ADD_405_U5 , P1_ADD_405_U6 , P1_ADD_405_U7 , P1_ADD_405_U8 , P1_ADD_405_U9 , P1_ADD_405_U10 , P1_ADD_405_U11 , P1_ADD_405_U12 , P1_ADD_405_U13 , P1_ADD_405_U14;
wire P1_ADD_405_U15 , P1_ADD_405_U16 , P1_ADD_405_U17 , P1_ADD_405_U18 , P1_ADD_405_U19 , P1_ADD_405_U20 , P1_ADD_405_U21 , P1_ADD_405_U22 , P1_ADD_405_U23 , P1_ADD_405_U24;
wire P1_ADD_405_U25 , P1_ADD_405_U26 , P1_ADD_405_U27 , P1_ADD_405_U28 , P1_ADD_405_U29 , P1_ADD_405_U30 , P1_ADD_405_U31 , P1_ADD_405_U32 , P1_ADD_405_U33 , P1_ADD_405_U34;
wire P1_ADD_405_U35 , P1_ADD_405_U36 , P1_ADD_405_U37 , P1_ADD_405_U38 , P1_ADD_405_U39 , P1_ADD_405_U40 , P1_ADD_405_U41 , P1_ADD_405_U42 , P1_ADD_405_U43 , P1_ADD_405_U44;
wire P1_ADD_405_U45 , P1_ADD_405_U46 , P1_ADD_405_U47 , P1_ADD_405_U48 , P1_ADD_405_U49 , P1_ADD_405_U50 , P1_ADD_405_U51 , P1_ADD_405_U52 , P1_ADD_405_U53 , P1_ADD_405_U54;
wire P1_ADD_405_U55 , P1_ADD_405_U56 , P1_ADD_405_U57 , P1_ADD_405_U58 , P1_ADD_405_U59 , P1_ADD_405_U60 , P1_ADD_405_U61 , P1_ADD_405_U62 , P1_ADD_405_U63 , P1_ADD_405_U64;
wire P1_ADD_405_U65 , P1_ADD_405_U66 , P1_ADD_405_U67 , P1_ADD_405_U68 , P1_ADD_405_U69 , P1_ADD_405_U70 , P1_ADD_405_U71 , P1_ADD_405_U72 , P1_ADD_405_U73 , P1_ADD_405_U74;
wire P1_ADD_405_U75 , P1_ADD_405_U76 , P1_ADD_405_U77 , P1_ADD_405_U78 , P1_ADD_405_U79 , P1_ADD_405_U80 , P1_ADD_405_U81 , P1_ADD_405_U82 , P1_ADD_405_U83 , P1_ADD_405_U84;
wire P1_ADD_405_U85 , P1_ADD_405_U86;


nand NAND2_1 ( P1_ADD_515_U182 , P1_ADD_515_U107 , P1_ADD_515_U33 );
nand NAND2_2 ( P1_ADD_515_U181 , P1_INSTADDRPOINTER_REG_16_ , P1_ADD_515_U32 );
nand NAND2_3 ( P1_ADD_515_U180 , P1_ADD_515_U116 , P1_ADD_515_U51 );
and AND2_4 ( U207 , U250 , U214 );
and AND4_5 ( U208 , P2_W_R_N_REG , P2_M_IO_N_REG , U378 , U377 );
and AND2_6 ( U209 , READY22_REG , READY2 );
and AND2_7 ( U210 , READY11_REG , READY1 );
and AND2_8 ( U211 , READY12_REG , READY21_REG );
nand NAND3_9 ( U212 , U208 , R170_U6 , U214 );
nand NAND4_10 ( U213 , P3_M_IO_N_REG , U380 , U379 , U215 );
nand NAND5_11 ( U214 , P1_M_IO_N_REG , U383 , P1_W_R_N_REG , U381 , R165_U6 );
nand NAND2_12 ( U215 , LT_748_U6 , U208 );
nand NAND3_13 ( U216 , U483 , U484 , U482 );
nand NAND3_14 ( U217 , U480 , U481 , U479 );
nand NAND3_15 ( U218 , U477 , U478 , U476 );
nand NAND3_16 ( U219 , U474 , U475 , U473 );
nand NAND3_17 ( U220 , U471 , U472 , U470 );
nand NAND3_18 ( U221 , U468 , U469 , U467 );
nand NAND3_19 ( U222 , U465 , U466 , U464 );
nand NAND3_20 ( U223 , U462 , U463 , U461 );
nand NAND3_21 ( U224 , U459 , U460 , U458 );
nand NAND3_22 ( U225 , U456 , U457 , U455 );
nand NAND3_23 ( U226 , U453 , U454 , U452 );
nand NAND3_24 ( U227 , U450 , U451 , U449 );
nand NAND3_25 ( U228 , U447 , U448 , U446 );
nand NAND3_26 ( U229 , U444 , U445 , U443 );
nand NAND3_27 ( U230 , U441 , U442 , U440 );
nand NAND3_28 ( U231 , U438 , U439 , U437 );
nand NAND3_29 ( U232 , U435 , U436 , U434 );
nand NAND3_30 ( U233 , U432 , U433 , U431 );
nand NAND3_31 ( U234 , U429 , U430 , U428 );
nand NAND3_32 ( U235 , U426 , U427 , U425 );
nand NAND3_33 ( U236 , U423 , U424 , U422 );
nand NAND3_34 ( U237 , U420 , U421 , U419 );
nand NAND3_35 ( U238 , U417 , U418 , U416 );
nand NAND3_36 ( U239 , U414 , U415 , U413 );
nand NAND3_37 ( U240 , U411 , U412 , U410 );
nand NAND3_38 ( U241 , U408 , U409 , U407 );
nand NAND3_39 ( U242 , U405 , U406 , U404 );
nand NAND3_40 ( U243 , U402 , U403 , U401 );
nand NAND3_41 ( U244 , U399 , U400 , U398 );
nand NAND3_42 ( U245 , U396 , U397 , U395 );
nand NAND3_43 ( U246 , U393 , U394 , U392 );
nand NAND3_44 ( U247 , U390 , U391 , U389 );
not NOT1_45 ( U248 , R165_U6 );
not NOT1_46 ( U249 , R170_U6 );
nand NAND2_47 ( U250 , U214 , U387 );
nand NAND2_48 ( U251 , U486 , U485 );
nand NAND2_49 ( U252 , U488 , U487 );
nand NAND2_50 ( U253 , U490 , U489 );
nand NAND2_51 ( U254 , U492 , U491 );
nand NAND2_52 ( U255 , U494 , U493 );
nand NAND2_53 ( U256 , U496 , U495 );
nand NAND2_54 ( U257 , U498 , U497 );
nand NAND2_55 ( U258 , U500 , U499 );
nand NAND2_56 ( U259 , U502 , U501 );
nand NAND2_57 ( U260 , U504 , U503 );
nand NAND2_58 ( U261 , U506 , U505 );
nand NAND2_59 ( U262 , U508 , U507 );
nand NAND2_60 ( U263 , U510 , U509 );
nand NAND2_61 ( U264 , U512 , U511 );
nand NAND2_62 ( U265 , U514 , U513 );
nand NAND2_63 ( U266 , U516 , U515 );
nand NAND2_64 ( U267 , U518 , U517 );
nand NAND2_65 ( U268 , U520 , U519 );
nand NAND2_66 ( U269 , U522 , U521 );
nand NAND2_67 ( U270 , U524 , U523 );
nand NAND2_68 ( U271 , U526 , U525 );
nand NAND2_69 ( U272 , U528 , U527 );
nand NAND2_70 ( U273 , U530 , U529 );
nand NAND2_71 ( U274 , U532 , U531 );
nand NAND2_72 ( U275 , U534 , U533 );
nand NAND2_73 ( U276 , U536 , U535 );
nand NAND2_74 ( U277 , U538 , U537 );
nand NAND2_75 ( U278 , U540 , U539 );
nand NAND2_76 ( U279 , U542 , U541 );
nand NAND2_77 ( U280 , U544 , U543 );
nand NAND2_78 ( U281 , U546 , U545 );
nand NAND2_79 ( U282 , U548 , U547 );
nand NAND2_80 ( U283 , U550 , U549 );
nand NAND2_81 ( U284 , U552 , U551 );
nand NAND2_82 ( U285 , U554 , U553 );
nand NAND2_83 ( U286 , U556 , U555 );
nand NAND2_84 ( U287 , U558 , U557 );
nand NAND2_85 ( U288 , U560 , U559 );
nand NAND2_86 ( U289 , U562 , U561 );
nand NAND2_87 ( U290 , U564 , U563 );
nand NAND2_88 ( U291 , U566 , U565 );
nand NAND2_89 ( U292 , U568 , U567 );
nand NAND2_90 ( U293 , U570 , U569 );
nand NAND2_91 ( U294 , U572 , U571 );
nand NAND2_92 ( U295 , U574 , U573 );
nand NAND2_93 ( U296 , U576 , U575 );
nand NAND2_94 ( U297 , U578 , U577 );
nand NAND2_95 ( U298 , U580 , U579 );
nand NAND2_96 ( U299 , U582 , U581 );
nand NAND2_97 ( U300 , U584 , U583 );
nand NAND2_98 ( U301 , U586 , U585 );
nand NAND2_99 ( U302 , U588 , U587 );
nand NAND2_100 ( U303 , U590 , U589 );
nand NAND2_101 ( U304 , U592 , U591 );
nand NAND2_102 ( U305 , U594 , U593 );
nand NAND2_103 ( U306 , U596 , U595 );
nand NAND2_104 ( U307 , U598 , U597 );
nand NAND2_105 ( U308 , U600 , U599 );
nand NAND2_106 ( U309 , U602 , U601 );
nand NAND2_107 ( U310 , U604 , U603 );
nand NAND2_108 ( U311 , U606 , U605 );
nand NAND2_109 ( U312 , U608 , U607 );
nand NAND2_110 ( U313 , U610 , U609 );
nand NAND2_111 ( U314 , U612 , U611 );
nand NAND2_112 ( U315 , U614 , U613 );
nand NAND2_113 ( U316 , U616 , U615 );
nand NAND2_114 ( U317 , U618 , U617 );
nand NAND2_115 ( U318 , U620 , U619 );
nand NAND2_116 ( U319 , U622 , U621 );
nand NAND2_117 ( U320 , U624 , U623 );
nand NAND2_118 ( U321 , U626 , U625 );
nand NAND2_119 ( U322 , U628 , U627 );
nand NAND2_120 ( U323 , U630 , U629 );
nand NAND2_121 ( U324 , U632 , U631 );
nand NAND2_122 ( U325 , U634 , U633 );
nand NAND2_123 ( U326 , U636 , U635 );
nand NAND2_124 ( U327 , U638 , U637 );
nand NAND2_125 ( U328 , U640 , U639 );
nand NAND2_126 ( U329 , U642 , U641 );
nand NAND2_127 ( U330 , U644 , U643 );
nand NAND2_128 ( U331 , U646 , U645 );
nand NAND2_129 ( U332 , U648 , U647 );
nand NAND2_130 ( U333 , U650 , U649 );
nand NAND2_131 ( U334 , U652 , U651 );
nand NAND2_132 ( U335 , U654 , U653 );
nand NAND2_133 ( U336 , U656 , U655 );
nand NAND2_134 ( U337 , U658 , U657 );
nand NAND2_135 ( U338 , U660 , U659 );
nand NAND2_136 ( U339 , U662 , U661 );
nand NAND2_137 ( U340 , U664 , U663 );
nand NAND2_138 ( U341 , U666 , U665 );
nand NAND2_139 ( U342 , U668 , U667 );
nand NAND2_140 ( U343 , U670 , U669 );
nand NAND2_141 ( U344 , U672 , U671 );
nand NAND2_142 ( U345 , U674 , U673 );
nand NAND2_143 ( U346 , U676 , U675 );
nand NAND2_144 ( U347 , U678 , U677 );
nand NAND2_145 ( U348 , U680 , U679 );
nand NAND2_146 ( U349 , U682 , U681 );
nand NAND2_147 ( U350 , U684 , U683 );
nand NAND2_148 ( U351 , U686 , U685 );
nand NAND2_149 ( U352 , U688 , U687 );
nand NAND2_150 ( U353 , U690 , U689 );
nand NAND2_151 ( U354 , U692 , U691 );
nand NAND2_152 ( U355 , U694 , U693 );
nand NAND2_153 ( U356 , U696 , U695 );
nand NAND2_154 ( U357 , U698 , U697 );
nand NAND2_155 ( U358 , U700 , U699 );
nand NAND2_156 ( U359 , U702 , U701 );
nand NAND2_157 ( U360 , U704 , U703 );
nand NAND2_158 ( U361 , U706 , U705 );
nand NAND2_159 ( U362 , U708 , U707 );
nand NAND2_160 ( U363 , U710 , U709 );
nand NAND2_161 ( U364 , U712 , U711 );
nand NAND2_162 ( U365 , U714 , U713 );
nand NAND2_163 ( U366 , U716 , U715 );
nand NAND2_164 ( U367 , U718 , U717 );
nand NAND2_165 ( U368 , U720 , U719 );
nand NAND2_166 ( U369 , U722 , U721 );
nand NAND2_167 ( U370 , U724 , U723 );
nand NAND2_168 ( U371 , U726 , U725 );
nand NAND2_169 ( U372 , U728 , U727 );
nand NAND2_170 ( U373 , U730 , U729 );
nand NAND2_171 ( U374 , U732 , U731 );
nand NAND2_172 ( U375 , U734 , U733 );
nand NAND2_173 ( U376 , U736 , U735 );
nor nor_174 ( U377 , P2_BE_N_REG_0_ , P2_ADS_N_REG , P2_BE_N_REG_2_ , P2_BE_N_REG_1_ );
nor nor_175 ( U378 , P2_D_C_N_REG , P2_BE_N_REG_3_ );
nor nor_176 ( U379 , P3_BE_N_REG_1_ , P3_BE_N_REG_0_ , P3_ADS_N_REG , P3_D_C_N_REG , P3_W_R_N_REG );
nor nor_177 ( U380 , P3_BE_N_REG_3_ , P3_BE_N_REG_2_ );
nor nor_178 ( U381 , P1_BE_N_REG_1_ , P1_BE_N_REG_3_ , P1_D_C_N_REG , P1_ADS_N_REG , P1_BE_N_REG_0_ );
nand NAND3_179 ( U382 , LT_782_120_U6 , LT_782_U6 , LT_782_119_U6 );
not NOT1_180 ( U383 , P1_BE_N_REG_2_ );
not NOT1_181 ( U384 , U382 );
not NOT1_182 ( U385 , U214 );
not NOT1_183 ( U386 , U215 );
nand NAND2_184 ( U387 , R170_U6 , U208 );
not NOT1_185 ( U388 , U250 );
nand NAND2_186 ( U389 , P2_DATAO_REG_0_ , U207 );
nand NAND2_187 ( U390 , P1_DATAO_REG_0_ , U385 );
nand NAND2_188 ( U391 , BUF1_REG_0_ , U388 );
nand NAND2_189 ( U392 , P2_DATAO_REG_1_ , U207 );
nand NAND2_190 ( U393 , P1_DATAO_REG_1_ , U385 );
nand NAND2_191 ( U394 , BUF1_REG_1_ , U388 );
nand NAND2_192 ( U395 , P2_DATAO_REG_2_ , U207 );
nand NAND2_193 ( U396 , P1_DATAO_REG_2_ , U385 );
nand NAND2_194 ( U397 , BUF1_REG_2_ , U388 );
nand NAND2_195 ( U398 , P2_DATAO_REG_3_ , U207 );
nand NAND2_196 ( U399 , P1_DATAO_REG_3_ , U385 );
nand NAND2_197 ( U400 , BUF1_REG_3_ , U388 );
nand NAND2_198 ( U401 , P2_DATAO_REG_4_ , U207 );
nand NAND2_199 ( U402 , P1_DATAO_REG_4_ , U385 );
nand NAND2_200 ( U403 , BUF1_REG_4_ , U388 );
nand NAND2_201 ( U404 , P2_DATAO_REG_5_ , U207 );
nand NAND2_202 ( U405 , P1_DATAO_REG_5_ , U385 );
nand NAND2_203 ( U406 , BUF1_REG_5_ , U388 );
nand NAND2_204 ( U407 , P2_DATAO_REG_6_ , U207 );
nand NAND2_205 ( U408 , P1_DATAO_REG_6_ , U385 );
nand NAND2_206 ( U409 , BUF1_REG_6_ , U388 );
nand NAND2_207 ( U410 , P2_DATAO_REG_7_ , U207 );
nand NAND2_208 ( U411 , P1_DATAO_REG_7_ , U385 );
nand NAND2_209 ( U412 , BUF1_REG_7_ , U388 );
nand NAND2_210 ( U413 , P2_DATAO_REG_8_ , U207 );
nand NAND2_211 ( U414 , P1_DATAO_REG_8_ , U385 );
nand NAND2_212 ( U415 , BUF1_REG_8_ , U388 );
nand NAND2_213 ( U416 , P2_DATAO_REG_9_ , U207 );
nand NAND2_214 ( U417 , P1_DATAO_REG_9_ , U385 );
nand NAND2_215 ( U418 , BUF1_REG_9_ , U388 );
nand NAND2_216 ( U419 , P2_DATAO_REG_10_ , U207 );
nand NAND2_217 ( U420 , P1_DATAO_REG_10_ , U385 );
nand NAND2_218 ( U421 , BUF1_REG_10_ , U388 );
nand NAND2_219 ( U422 , P2_DATAO_REG_11_ , U207 );
nand NAND2_220 ( U423 , P1_DATAO_REG_11_ , U385 );
nand NAND2_221 ( U424 , BUF1_REG_11_ , U388 );
nand NAND2_222 ( U425 , P2_DATAO_REG_12_ , U207 );
nand NAND2_223 ( U426 , P1_DATAO_REG_12_ , U385 );
nand NAND2_224 ( U427 , BUF1_REG_12_ , U388 );
nand NAND2_225 ( U428 , P2_DATAO_REG_13_ , U207 );
nand NAND2_226 ( U429 , P1_DATAO_REG_13_ , U385 );
nand NAND2_227 ( U430 , BUF1_REG_13_ , U388 );
nand NAND2_228 ( U431 , P2_DATAO_REG_14_ , U207 );
nand NAND2_229 ( U432 , P1_DATAO_REG_14_ , U385 );
nand NAND2_230 ( U433 , BUF1_REG_14_ , U388 );
nand NAND2_231 ( U434 , P2_DATAO_REG_15_ , U207 );
nand NAND2_232 ( U435 , P1_DATAO_REG_15_ , U385 );
nand NAND2_233 ( U436 , BUF1_REG_15_ , U388 );
nand NAND2_234 ( U437 , P2_DATAO_REG_16_ , U207 );
nand NAND2_235 ( U438 , P1_DATAO_REG_16_ , U385 );
nand NAND2_236 ( U439 , BUF1_REG_16_ , U388 );
nand NAND2_237 ( U440 , P2_DATAO_REG_17_ , U207 );
nand NAND2_238 ( U441 , P1_DATAO_REG_17_ , U385 );
nand NAND2_239 ( U442 , BUF1_REG_17_ , U388 );
nand NAND2_240 ( U443 , P2_DATAO_REG_18_ , U207 );
nand NAND2_241 ( U444 , P1_DATAO_REG_18_ , U385 );
nand NAND2_242 ( U445 , BUF1_REG_18_ , U388 );
nand NAND2_243 ( U446 , P2_DATAO_REG_19_ , U207 );
nand NAND2_244 ( U447 , P1_DATAO_REG_19_ , U385 );
nand NAND2_245 ( U448 , BUF1_REG_19_ , U388 );
nand NAND2_246 ( U449 , P2_DATAO_REG_20_ , U207 );
nand NAND2_247 ( U450 , P1_DATAO_REG_20_ , U385 );
nand NAND2_248 ( U451 , BUF1_REG_20_ , U388 );
nand NAND2_249 ( U452 , P2_DATAO_REG_21_ , U207 );
nand NAND2_250 ( U453 , P1_DATAO_REG_21_ , U385 );
nand NAND2_251 ( U454 , BUF1_REG_21_ , U388 );
nand NAND2_252 ( U455 , P2_DATAO_REG_22_ , U207 );
nand NAND2_253 ( U456 , P1_DATAO_REG_22_ , U385 );
nand NAND2_254 ( U457 , BUF1_REG_22_ , U388 );
nand NAND2_255 ( U458 , P2_DATAO_REG_23_ , U207 );
nand NAND2_256 ( U459 , P1_DATAO_REG_23_ , U385 );
nand NAND2_257 ( U460 , BUF1_REG_23_ , U388 );
nand NAND2_258 ( U461 , P2_DATAO_REG_24_ , U207 );
nand NAND2_259 ( U462 , P1_DATAO_REG_24_ , U385 );
nand NAND2_260 ( U463 , BUF1_REG_24_ , U388 );
nand NAND2_261 ( U464 , P2_DATAO_REG_25_ , U207 );
nand NAND2_262 ( U465 , P1_DATAO_REG_25_ , U385 );
nand NAND2_263 ( U466 , BUF1_REG_25_ , U388 );
nand NAND2_264 ( U467 , P2_DATAO_REG_26_ , U207 );
nand NAND2_265 ( U468 , P1_DATAO_REG_26_ , U385 );
nand NAND2_266 ( U469 , BUF1_REG_26_ , U388 );
nand NAND2_267 ( U470 , P2_DATAO_REG_27_ , U207 );
nand NAND2_268 ( U471 , P1_DATAO_REG_27_ , U385 );
nand NAND2_269 ( U472 , BUF1_REG_27_ , U388 );
nand NAND2_270 ( U473 , P2_DATAO_REG_28_ , U207 );
nand NAND2_271 ( U474 , P1_DATAO_REG_28_ , U385 );
nand NAND2_272 ( U475 , BUF1_REG_28_ , U388 );
nand NAND2_273 ( U476 , P2_DATAO_REG_29_ , U207 );
nand NAND2_274 ( U477 , P1_DATAO_REG_29_ , U385 );
nand NAND2_275 ( U478 , BUF1_REG_29_ , U388 );
nand NAND2_276 ( U479 , P2_DATAO_REG_30_ , U207 );
nand NAND2_277 ( U480 , P1_DATAO_REG_30_ , U385 );
nand NAND2_278 ( U481 , BUF1_REG_30_ , U388 );
nand NAND2_279 ( U482 , P2_DATAO_REG_31_ , U207 );
nand NAND2_280 ( U483 , P1_DATAO_REG_31_ , U385 );
nand NAND2_281 ( U484 , BUF1_REG_31_ , U388 );
nand NAND2_282 ( U485 , BUF2_REG_0_ , U215 );
nand NAND2_283 ( U486 , P2_DATAO_REG_0_ , U386 );
nand NAND2_284 ( U487 , BUF2_REG_1_ , U215 );
nand NAND2_285 ( U488 , P2_DATAO_REG_1_ , U386 );
nand NAND2_286 ( U489 , BUF2_REG_2_ , U215 );
nand NAND2_287 ( U490 , P2_DATAO_REG_2_ , U386 );
nand NAND2_288 ( U491 , BUF2_REG_3_ , U215 );
nand NAND2_289 ( U492 , P2_DATAO_REG_3_ , U386 );
nand NAND2_290 ( U493 , BUF2_REG_4_ , U215 );
nand NAND2_291 ( U494 , P2_DATAO_REG_4_ , U386 );
nand NAND2_292 ( U495 , BUF2_REG_5_ , U215 );
nand NAND2_293 ( U496 , P2_DATAO_REG_5_ , U386 );
nand NAND2_294 ( U497 , BUF2_REG_6_ , U215 );
nand NAND2_295 ( U498 , P2_DATAO_REG_6_ , U386 );
nand NAND2_296 ( U499 , BUF2_REG_7_ , U215 );
nand NAND2_297 ( U500 , P2_DATAO_REG_7_ , U386 );
nand NAND2_298 ( U501 , BUF2_REG_8_ , U215 );
nand NAND2_299 ( U502 , P2_DATAO_REG_8_ , U386 );
nand NAND2_300 ( U503 , BUF2_REG_9_ , U215 );
nand NAND2_301 ( U504 , P2_DATAO_REG_9_ , U386 );
nand NAND2_302 ( U505 , BUF2_REG_10_ , U215 );
nand NAND2_303 ( U506 , P2_DATAO_REG_10_ , U386 );
nand NAND2_304 ( U507 , BUF2_REG_11_ , U215 );
nand NAND2_305 ( U508 , P2_DATAO_REG_11_ , U386 );
nand NAND2_306 ( U509 , BUF2_REG_12_ , U215 );
nand NAND2_307 ( U510 , P2_DATAO_REG_12_ , U386 );
nand NAND2_308 ( U511 , BUF2_REG_13_ , U215 );
nand NAND2_309 ( U512 , P2_DATAO_REG_13_ , U386 );
nand NAND2_310 ( U513 , BUF2_REG_14_ , U215 );
nand NAND2_311 ( U514 , P2_DATAO_REG_14_ , U386 );
nand NAND2_312 ( U515 , BUF2_REG_15_ , U215 );
nand NAND2_313 ( U516 , P2_DATAO_REG_15_ , U386 );
nand NAND2_314 ( U517 , BUF2_REG_16_ , U215 );
nand NAND2_315 ( U518 , P2_DATAO_REG_16_ , U386 );
nand NAND2_316 ( U519 , BUF2_REG_17_ , U215 );
nand NAND2_317 ( U520 , P2_DATAO_REG_17_ , U386 );
nand NAND2_318 ( U521 , BUF2_REG_18_ , U215 );
nand NAND2_319 ( U522 , P2_DATAO_REG_18_ , U386 );
nand NAND2_320 ( U523 , BUF2_REG_19_ , U215 );
nand NAND2_321 ( U524 , P2_DATAO_REG_19_ , U386 );
nand NAND2_322 ( U525 , BUF2_REG_20_ , U215 );
nand NAND2_323 ( U526 , P2_DATAO_REG_20_ , U386 );
nand NAND2_324 ( U527 , BUF2_REG_21_ , U215 );
nand NAND2_325 ( U528 , P2_DATAO_REG_21_ , U386 );
nand NAND2_326 ( U529 , BUF2_REG_22_ , U215 );
nand NAND2_327 ( U530 , P2_DATAO_REG_22_ , U386 );
nand NAND2_328 ( U531 , BUF2_REG_23_ , U215 );
nand NAND2_329 ( U532 , P2_DATAO_REG_23_ , U386 );
nand NAND2_330 ( U533 , BUF2_REG_24_ , U215 );
nand NAND2_331 ( U534 , P2_DATAO_REG_24_ , U386 );
nand NAND2_332 ( U535 , BUF2_REG_25_ , U215 );
nand NAND2_333 ( U536 , P2_DATAO_REG_25_ , U386 );
nand NAND2_334 ( U537 , BUF2_REG_26_ , U215 );
nand NAND2_335 ( U538 , P2_DATAO_REG_26_ , U386 );
nand NAND2_336 ( U539 , BUF2_REG_27_ , U215 );
nand NAND2_337 ( U540 , P2_DATAO_REG_27_ , U386 );
nand NAND2_338 ( U541 , BUF2_REG_28_ , U215 );
nand NAND2_339 ( U542 , P2_DATAO_REG_28_ , U386 );
nand NAND2_340 ( U543 , BUF2_REG_29_ , U215 );
nand NAND2_341 ( U544 , P2_DATAO_REG_29_ , U386 );
nand NAND2_342 ( U545 , BUF2_REG_30_ , U215 );
nand NAND2_343 ( U546 , P2_DATAO_REG_30_ , U386 );
nand NAND2_344 ( U547 , BUF2_REG_31_ , U215 );
nand NAND2_345 ( U548 , P2_DATAO_REG_31_ , U386 );
nand NAND2_346 ( U549 , BUF2_REG_9_ , U249 );
nand NAND2_347 ( U550 , BUF1_REG_9_ , R170_U6 );
nand NAND2_348 ( U551 , BUF2_REG_8_ , U249 );
nand NAND2_349 ( U552 , BUF1_REG_8_ , R170_U6 );
nand NAND2_350 ( U553 , BUF2_REG_7_ , U249 );
nand NAND2_351 ( U554 , BUF1_REG_7_ , R170_U6 );
nand NAND2_352 ( U555 , BUF2_REG_6_ , U249 );
nand NAND2_353 ( U556 , BUF1_REG_6_ , R170_U6 );
nand NAND2_354 ( U557 , BUF2_REG_5_ , U249 );
nand NAND2_355 ( U558 , BUF1_REG_5_ , R170_U6 );
nand NAND2_356 ( U559 , BUF2_REG_4_ , U249 );
nand NAND2_357 ( U560 , BUF1_REG_4_ , R170_U6 );
nand NAND2_358 ( U561 , BUF2_REG_3_ , U249 );
nand NAND2_359 ( U562 , BUF1_REG_3_ , R170_U6 );
nand NAND2_360 ( U563 , BUF2_REG_31_ , U249 );
nand NAND2_361 ( U564 , BUF1_REG_31_ , R170_U6 );
nand NAND2_362 ( U565 , BUF2_REG_30_ , U249 );
nand NAND2_363 ( U566 , BUF1_REG_30_ , R170_U6 );
nand NAND2_364 ( U567 , BUF2_REG_2_ , U249 );
nand NAND2_365 ( U568 , BUF1_REG_2_ , R170_U6 );
nand NAND2_366 ( U569 , BUF2_REG_29_ , U249 );
nand NAND2_367 ( U570 , BUF1_REG_29_ , R170_U6 );
nand NAND2_368 ( U571 , BUF2_REG_28_ , U249 );
nand NAND2_369 ( U572 , BUF1_REG_28_ , R170_U6 );
nand NAND2_370 ( U573 , BUF2_REG_27_ , U249 );
nand NAND2_371 ( U574 , BUF1_REG_27_ , R170_U6 );
nand NAND2_372 ( U575 , BUF2_REG_26_ , U249 );
nand NAND2_373 ( U576 , BUF1_REG_26_ , R170_U6 );
nand NAND2_374 ( U577 , BUF2_REG_25_ , U249 );
nand NAND2_375 ( U578 , BUF1_REG_25_ , R170_U6 );
nand NAND2_376 ( U579 , BUF2_REG_24_ , U249 );
nand NAND2_377 ( U580 , BUF1_REG_24_ , R170_U6 );
nand NAND2_378 ( U581 , BUF2_REG_23_ , U249 );
nand NAND2_379 ( U582 , BUF1_REG_23_ , R170_U6 );
nand NAND2_380 ( U583 , BUF2_REG_22_ , U249 );
nand NAND2_381 ( U584 , BUF1_REG_22_ , R170_U6 );
nand NAND2_382 ( U585 , BUF2_REG_21_ , U249 );
nand NAND2_383 ( U586 , BUF1_REG_21_ , R170_U6 );
nand NAND2_384 ( U587 , BUF2_REG_20_ , U249 );
nand NAND2_385 ( U588 , BUF1_REG_20_ , R170_U6 );
nand NAND2_386 ( U589 , BUF2_REG_1_ , U249 );
nand NAND2_387 ( U590 , BUF1_REG_1_ , R170_U6 );
nand NAND2_388 ( U591 , BUF2_REG_19_ , U249 );
nand NAND2_389 ( U592 , BUF1_REG_19_ , R170_U6 );
nand NAND2_390 ( U593 , BUF2_REG_18_ , U249 );
nand NAND2_391 ( U594 , BUF1_REG_18_ , R170_U6 );
nand NAND2_392 ( U595 , BUF2_REG_17_ , U249 );
nand NAND2_393 ( U596 , BUF1_REG_17_ , R170_U6 );
nand NAND2_394 ( U597 , BUF2_REG_16_ , U249 );
nand NAND2_395 ( U598 , BUF1_REG_16_ , R170_U6 );
nand NAND2_396 ( U599 , BUF2_REG_15_ , U249 );
nand NAND2_397 ( U600 , BUF1_REG_15_ , R170_U6 );
nand NAND2_398 ( U601 , BUF2_REG_14_ , U249 );
nand NAND2_399 ( U602 , BUF1_REG_14_ , R170_U6 );
nand NAND2_400 ( U603 , BUF2_REG_13_ , U249 );
nand NAND2_401 ( U604 , BUF1_REG_13_ , R170_U6 );
nand NAND2_402 ( U605 , BUF2_REG_12_ , U249 );
nand NAND2_403 ( U606 , BUF1_REG_12_ , R170_U6 );
nand NAND2_404 ( U607 , BUF2_REG_11_ , U249 );
nand NAND2_405 ( U608 , BUF1_REG_11_ , R170_U6 );
nand NAND2_406 ( U609 , BUF2_REG_10_ , U249 );
nand NAND2_407 ( U610 , BUF1_REG_10_ , R170_U6 );
nand NAND2_408 ( U611 , BUF2_REG_0_ , U249 );
nand NAND2_409 ( U612 , BUF1_REG_0_ , R170_U6 );
nand NAND2_410 ( U613 , DATAI_9_ , U248 );
nand NAND2_411 ( U614 , BUF1_REG_9_ , R165_U6 );
nand NAND2_412 ( U615 , DATAI_8_ , U248 );
nand NAND2_413 ( U616 , BUF1_REG_8_ , R165_U6 );
nand NAND2_414 ( U617 , DATAI_7_ , U248 );
nand NAND2_415 ( U618 , BUF1_REG_7_ , R165_U6 );
nand NAND2_416 ( U619 , DATAI_6_ , U248 );
nand NAND2_417 ( U620 , BUF1_REG_6_ , R165_U6 );
nand NAND2_418 ( U621 , DATAI_5_ , U248 );
nand NAND2_419 ( U622 , BUF1_REG_5_ , R165_U6 );
nand NAND2_420 ( U623 , DATAI_4_ , U248 );
nand NAND2_421 ( U624 , BUF1_REG_4_ , R165_U6 );
nand NAND2_422 ( U625 , DATAI_3_ , U248 );
nand NAND2_423 ( U626 , BUF1_REG_3_ , R165_U6 );
nand NAND2_424 ( U627 , DATAI_31_ , U248 );
nand NAND2_425 ( U628 , BUF1_REG_31_ , R165_U6 );
nand NAND2_426 ( U629 , DATAI_30_ , U248 );
nand NAND2_427 ( U630 , BUF1_REG_30_ , R165_U6 );
nand NAND2_428 ( U631 , DATAI_2_ , U248 );
nand NAND2_429 ( U632 , BUF1_REG_2_ , R165_U6 );
nand NAND2_430 ( U633 , DATAI_29_ , U248 );
nand NAND2_431 ( U634 , BUF1_REG_29_ , R165_U6 );
nand NAND2_432 ( U635 , DATAI_28_ , U248 );
nand NAND2_433 ( U636 , BUF1_REG_28_ , R165_U6 );
nand NAND2_434 ( U637 , DATAI_27_ , U248 );
nand NAND2_435 ( U638 , BUF1_REG_27_ , R165_U6 );
nand NAND2_436 ( U639 , DATAI_26_ , U248 );
nand NAND2_437 ( U640 , BUF1_REG_26_ , R165_U6 );
nand NAND2_438 ( U641 , DATAI_25_ , U248 );
nand NAND2_439 ( U642 , BUF1_REG_25_ , R165_U6 );
nand NAND2_440 ( U643 , DATAI_24_ , U248 );
nand NAND2_441 ( U644 , BUF1_REG_24_ , R165_U6 );
nand NAND2_442 ( U645 , DATAI_23_ , U248 );
nand NAND2_443 ( U646 , BUF1_REG_23_ , R165_U6 );
nand NAND2_444 ( U647 , DATAI_22_ , U248 );
nand NAND2_445 ( U648 , BUF1_REG_22_ , R165_U6 );
nand NAND2_446 ( U649 , DATAI_21_ , U248 );
nand NAND2_447 ( U650 , BUF1_REG_21_ , R165_U6 );
nand NAND2_448 ( U651 , DATAI_20_ , U248 );
nand NAND2_449 ( U652 , BUF1_REG_20_ , R165_U6 );
nand NAND2_450 ( U653 , DATAI_1_ , U248 );
nand NAND2_451 ( U654 , BUF1_REG_1_ , R165_U6 );
nand NAND2_452 ( U655 , DATAI_19_ , U248 );
nand NAND2_453 ( U656 , BUF1_REG_19_ , R165_U6 );
nand NAND2_454 ( U657 , DATAI_18_ , U248 );
nand NAND2_455 ( U658 , BUF1_REG_18_ , R165_U6 );
nand NAND2_456 ( U659 , DATAI_17_ , U248 );
nand NAND2_457 ( U660 , BUF1_REG_17_ , R165_U6 );
nand NAND2_458 ( U661 , DATAI_16_ , U248 );
nand NAND2_459 ( U662 , BUF1_REG_16_ , R165_U6 );
nand NAND2_460 ( U663 , DATAI_15_ , U248 );
nand NAND2_461 ( U664 , BUF1_REG_15_ , R165_U6 );
nand NAND2_462 ( U665 , DATAI_14_ , U248 );
nand NAND2_463 ( U666 , BUF1_REG_14_ , R165_U6 );
nand NAND2_464 ( U667 , DATAI_13_ , U248 );
nand NAND2_465 ( U668 , BUF1_REG_13_ , R165_U6 );
nand NAND2_466 ( U669 , DATAI_12_ , U248 );
nand NAND2_467 ( U670 , BUF1_REG_12_ , R165_U6 );
nand NAND2_468 ( U671 , DATAI_11_ , U248 );
nand NAND2_469 ( U672 , BUF1_REG_11_ , R165_U6 );
nand NAND2_470 ( U673 , DATAI_10_ , U248 );
nand NAND2_471 ( U674 , BUF1_REG_10_ , R165_U6 );
nand NAND2_472 ( U675 , DATAI_0_ , U248 );
nand NAND2_473 ( U676 , BUF1_REG_0_ , R165_U6 );
nand NAND2_474 ( U677 , P2_ADDRESS_REG_9_ , U382 );
nand NAND2_475 ( U678 , P3_ADDRESS_REG_9_ , U384 );
nand NAND2_476 ( U679 , P2_ADDRESS_REG_8_ , U382 );
nand NAND2_477 ( U680 , P3_ADDRESS_REG_8_ , U384 );
nand NAND2_478 ( U681 , P2_ADDRESS_REG_7_ , U382 );
nand NAND2_479 ( U682 , P3_ADDRESS_REG_7_ , U384 );
nand NAND2_480 ( U683 , P2_ADDRESS_REG_6_ , U382 );
nand NAND2_481 ( U684 , P3_ADDRESS_REG_6_ , U384 );
nand NAND2_482 ( U685 , P2_ADDRESS_REG_5_ , U382 );
nand NAND2_483 ( U686 , P3_ADDRESS_REG_5_ , U384 );
nand NAND2_484 ( U687 , P2_ADDRESS_REG_4_ , U382 );
nand NAND2_485 ( U688 , P3_ADDRESS_REG_4_ , U384 );
nand NAND2_486 ( U689 , P2_ADDRESS_REG_3_ , U382 );
nand NAND2_487 ( U690 , P3_ADDRESS_REG_3_ , U384 );
nand NAND2_488 ( U691 , P2_ADDRESS_REG_2_ , U382 );
nand NAND2_489 ( U692 , P3_ADDRESS_REG_2_ , U384 );
nand NAND2_490 ( U693 , P2_ADDRESS_REG_29_ , U382 );
nand NAND2_491 ( U694 , P3_ADDRESS_REG_29_ , U384 );
nand NAND2_492 ( U695 , P2_ADDRESS_REG_28_ , U382 );
nand NAND2_493 ( U696 , P3_ADDRESS_REG_28_ , U384 );
nand NAND2_494 ( U697 , P2_ADDRESS_REG_27_ , U382 );
nand NAND2_495 ( U698 , P3_ADDRESS_REG_27_ , U384 );
nand NAND2_496 ( U699 , P2_ADDRESS_REG_26_ , U382 );
nand NAND2_497 ( U700 , P3_ADDRESS_REG_26_ , U384 );
nand NAND2_498 ( U701 , P2_ADDRESS_REG_25_ , U382 );
nand NAND2_499 ( U702 , P3_ADDRESS_REG_25_ , U384 );
nand NAND2_500 ( U703 , P2_ADDRESS_REG_24_ , U382 );
nand NAND2_501 ( U704 , P3_ADDRESS_REG_24_ , U384 );
nand NAND2_502 ( U705 , P2_ADDRESS_REG_23_ , U382 );
nand NAND2_503 ( U706 , P3_ADDRESS_REG_23_ , U384 );
nand NAND2_504 ( U707 , P2_ADDRESS_REG_22_ , U382 );
nand NAND2_505 ( U708 , P3_ADDRESS_REG_22_ , U384 );
nand NAND2_506 ( U709 , P2_ADDRESS_REG_21_ , U382 );
nand NAND2_507 ( U710 , P3_ADDRESS_REG_21_ , U384 );
nand NAND2_508 ( U711 , P2_ADDRESS_REG_20_ , U382 );
nand NAND2_509 ( U712 , P3_ADDRESS_REG_20_ , U384 );
nand NAND2_510 ( U713 , P2_ADDRESS_REG_1_ , U382 );
nand NAND2_511 ( U714 , P3_ADDRESS_REG_1_ , U384 );
nand NAND2_512 ( U715 , P2_ADDRESS_REG_19_ , U382 );
nand NAND2_513 ( U716 , P3_ADDRESS_REG_19_ , U384 );
nand NAND2_514 ( U717 , P2_ADDRESS_REG_18_ , U382 );
nand NAND2_515 ( U718 , P3_ADDRESS_REG_18_ , U384 );
nand NAND2_516 ( U719 , P2_ADDRESS_REG_17_ , U382 );
nand NAND2_517 ( U720 , P3_ADDRESS_REG_17_ , U384 );
nand NAND2_518 ( U721 , P2_ADDRESS_REG_16_ , U382 );
nand NAND2_519 ( U722 , P3_ADDRESS_REG_16_ , U384 );
nand NAND2_520 ( U723 , P2_ADDRESS_REG_15_ , U382 );
nand NAND2_521 ( U724 , P3_ADDRESS_REG_15_ , U384 );
nand NAND2_522 ( U725 , P2_ADDRESS_REG_14_ , U382 );
nand NAND2_523 ( U726 , P3_ADDRESS_REG_14_ , U384 );
nand NAND2_524 ( U727 , P2_ADDRESS_REG_13_ , U382 );
nand NAND2_525 ( U728 , P3_ADDRESS_REG_13_ , U384 );
nand NAND2_526 ( U729 , P2_ADDRESS_REG_12_ , U382 );
nand NAND2_527 ( U730 , P3_ADDRESS_REG_12_ , U384 );
nand NAND2_528 ( U731 , P2_ADDRESS_REG_11_ , U382 );
nand NAND2_529 ( U732 , P3_ADDRESS_REG_11_ , U384 );
nand NAND2_530 ( U733 , P2_ADDRESS_REG_10_ , U382 );
nand NAND2_531 ( U734 , P3_ADDRESS_REG_10_ , U384 );
nand NAND2_532 ( U735 , P2_ADDRESS_REG_0_ , U382 );
nand NAND2_533 ( U736 , P3_ADDRESS_REG_0_ , U384 );
nand NAND2_534 ( P1_ADD_515_U179 , P1_INSTADDRPOINTER_REG_25_ , P1_ADD_515_U50 );
nand NAND2_535 ( P1_ADD_515_U178 , P1_ADD_515_U98 , P1_ADD_515_U15 );
nand NAND2_536 ( P1_ADD_515_U177 , P1_INSTADDRPOINTER_REG_7_ , P1_ADD_515_U14 );
nand NAND2_537 ( P1_ADD_515_U176 , P1_ADD_515_U103 , P1_ADD_515_U25 );
nand NAND2_538 ( P1_ADD_515_U175 , P1_INSTADDRPOINTER_REG_12_ , P1_ADD_515_U24 );
nand NAND2_539 ( P1_ADD_515_U174 , P1_ADD_515_U112 , P1_ADD_515_U43 );
nand NAND2_540 ( P1_ADD_515_U173 , P1_INSTADDRPOINTER_REG_21_ , P1_ADD_515_U42 );
nand NAND2_541 ( P1_ADD_515_U172 , P1_ADD_515_U119 , P1_ADD_515_U57 );
nand NAND2_542 ( P1_ADD_515_U171 , P1_INSTADDRPOINTER_REG_28_ , P1_ADD_515_U56 );
nor nor_543 ( P3_U2352 , U209 , P3_STATEBS16_REG );
and AND2_544 ( P3_U2353 , P3_U3354 , P3_U2449 );
and AND2_545 ( P3_U2354 , P3_U3688 , P3_U4325 );
and AND2_546 ( P3_U2355 , P3_U3689 , P3_U4325 );
and AND2_547 ( P3_U2356 , P3_U3355 , P3_U2353 );
and AND2_548 ( P3_U2357 , P3_U4323 , P3_U2451 );
and AND2_549 ( P3_U2358 , P3_U3690 , P3_U4341 );
and AND2_550 ( P3_U2359 , P3_U4324 , P3_U2462 );
and AND2_551 ( P3_U2360 , P3_U4296 , P3_U2462 );
and AND2_552 ( P3_U2361 , P3_U4297 , P3_U2462 );
and AND2_553 ( P3_U2362 , P3_U3691 , P3_U4341 );
and AND2_554 ( P3_U2363 , P3_U5442 , P3_U5435 );
and AND2_555 ( P3_U2364 , P3_U5392 , P3_U3204 );
and AND2_556 ( P3_U2365 , P3_U5341 , P3_U3201 );
and AND2_557 ( P3_U2366 , P3_U5290 , P3_U3198 );
and AND2_558 ( P3_U2367 , P3_U5239 , P3_U5232 );
and AND2_559 ( P3_U2368 , P3_U5189 , P3_U3193 );
and AND2_560 ( P3_U2369 , P3_U5137 , P3_U3189 );
and AND2_561 ( P3_U2370 , P3_U5085 , P3_U3185 );
and AND2_562 ( P3_U2371 , P3_U5036 , P3_U5028 );
and AND2_563 ( P3_U2372 , P3_U4985 , P3_U3176 );
and AND2_564 ( P3_U2373 , P3_U4933 , P3_U3172 );
and AND2_565 ( P3_U2374 , P3_U4881 , P3_U3168 );
and AND2_566 ( P3_U2375 , P3_U4829 , P3_U4821 );
and AND2_567 ( P3_U2376 , P3_U4778 , P3_U3160 );
and AND2_568 ( P3_U2377 , P3_U4726 , P3_U3152 );
and AND2_569 ( P3_U2378 , P3_U4674 , P3_U3146 );
and AND2_570 ( P3_U2379 , P3_U4322 , P3_U4312 );
and AND2_571 ( P3_U2380 , P3_STATE2_REG_2_ , P3_U3260 );
and AND2_572 ( P3_U2381 , P3_U4312 , P3_STATE2_REG_3_ );
and AND2_573 ( P3_U2382 , P3_U3951 , P3_U3249 );
and AND2_574 ( P3_U2383 , P3_U2380 , P3_U4296 );
and AND2_575 ( P3_U2384 , P3_U2380 , P3_U4297 );
and AND2_576 ( P3_U2385 , P3_STATE2_REG_1_ , P3_U3260 );
and AND2_577 ( P3_U2386 , P3_STATE2_REG_1_ , P3_U3249 );
and AND2_578 ( P3_U2387 , P3_U3953 , P3_U3249 );
and AND2_579 ( P3_U2388 , P3_U3952 , P3_U3249 );
and AND2_580 ( P3_U2389 , P3_U4354 , P3_U3249 );
and AND2_581 ( P3_U2390 , P3_U4353 , P3_STATE2_REG_0_ );
and AND2_582 ( P3_U2391 , P3_U4310 , P3_U3218 );
and AND2_583 ( P3_U2392 , P3_U2383 , P3_U4293 );
and AND2_584 ( P3_U2393 , P3_U2628 , P3_U2361 );
and AND2_585 ( P3_U2394 , P3_U2382 , P3_U2628 );
and AND2_586 ( P3_U2395 , P3_U2361 , P3_U3241 );
and AND2_587 ( P3_U2396 , P3_U2382 , P3_U3241 );
and AND2_588 ( P3_U2397 , P3_U2386 , P3_STATEBS16_REG );
and AND2_589 ( P3_U2398 , P3_U2386 , P3_U2631 );
and AND2_590 ( P3_U2399 , P3_U4309 , P3_U4573 );
and AND2_591 ( P3_U2400 , P3_U4310 , P3_U4573 );
and AND2_592 ( P3_U2401 , P3_STATE2_REG_3_ , P3_U3260 );
and AND2_593 ( P3_U2402 , P3_U3248 , P3_U3090 );
and AND2_594 ( P3_U2403 , P3_U2385 , P3_U3258 );
and AND2_595 ( P3_U2404 , P3_U2384 , P3_U3257 );
and AND2_596 ( P3_U2405 , P3_U7095 , P3_U2384 );
and AND2_597 ( P3_U2406 , P3_U4311 , P3_U3104 );
and AND2_598 ( P3_U2407 , P3_U4311 , P3_U4505 );
and AND2_599 ( P3_U2408 , P3_U4309 , P3_U3218 );
and AND2_600 ( P3_U2409 , P3_STATE2_REG_0_ , P3_U3251 );
and AND2_601 ( P3_U2410 , P3_U3251 , P3_U3121 );
and AND2_602 ( P3_U2411 , P3_U4310 , P3_U4608 );
and AND3_603 ( P3_U2412 , P3_U3218 , P3_U3107 , P3_U4539 );
and AND2_604 ( P3_U2413 , BUF2_REG_0_ , P3_U4312 );
and AND2_605 ( P3_U2414 , BUF2_REG_1_ , P3_U4312 );
and AND2_606 ( P3_U2415 , BUF2_REG_2_ , P3_U4312 );
and AND2_607 ( P3_U2416 , BUF2_REG_3_ , P3_U4312 );
and AND2_608 ( P3_U2417 , BUF2_REG_4_ , P3_U4312 );
and AND2_609 ( P3_U2418 , BUF2_REG_5_ , P3_U4312 );
and AND2_610 ( P3_U2419 , BUF2_REG_6_ , P3_U4312 );
and AND2_611 ( P3_U2420 , BUF2_REG_7_ , P3_U4312 );
and AND2_612 ( P3_U2421 , BUF2_REG_24_ , P3_U2379 );
and AND2_613 ( P3_U2422 , BUF2_REG_16_ , P3_U2379 );
and AND2_614 ( P3_U2423 , BUF2_REG_25_ , P3_U2379 );
and AND2_615 ( P3_U2424 , BUF2_REG_17_ , P3_U2379 );
and AND2_616 ( P3_U2425 , BUF2_REG_26_ , P3_U2379 );
and AND2_617 ( P3_U2426 , BUF2_REG_18_ , P3_U2379 );
and AND2_618 ( P3_U2427 , BUF2_REG_27_ , P3_U2379 );
and AND2_619 ( P3_U2428 , BUF2_REG_19_ , P3_U2379 );
and AND2_620 ( P3_U2429 , BUF2_REG_28_ , P3_U2379 );
and AND2_621 ( P3_U2430 , BUF2_REG_20_ , P3_U2379 );
and AND2_622 ( P3_U2431 , BUF2_REG_29_ , P3_U2379 );
and AND2_623 ( P3_U2432 , BUF2_REG_21_ , P3_U2379 );
and AND2_624 ( P3_U2433 , BUF2_REG_30_ , P3_U2379 );
and AND2_625 ( P3_U2434 , BUF2_REG_22_ , P3_U2379 );
and AND2_626 ( P3_U2435 , BUF2_REG_31_ , P3_U2379 );
and AND2_627 ( P3_U2436 , BUF2_REG_23_ , P3_U2379 );
and AND2_628 ( P3_U2437 , P3_U2381 , P3_U3108 );
and AND2_629 ( P3_U2438 , P3_U2381 , P3_U3104 );
and AND2_630 ( P3_U2439 , P3_U2381 , P3_U3101 );
and AND2_631 ( P3_U2440 , P3_U2381 , P3_U3107 );
and AND2_632 ( P3_U2441 , P3_U2381 , P3_U3102 );
and AND2_633 ( P3_U2442 , P3_U2381 , P3_U3110 );
and AND2_634 ( P3_U2443 , P3_U2381 , P3_U3074 );
and AND2_635 ( P3_U2444 , P3_U2391 , P3_U3074 );
and AND2_636 ( P3_U2445 , P3_U2381 , P3_U3218 );
and AND2_637 ( P3_U2446 , P3_U2391 , P3_U3113 );
and AND2_638 ( P3_U2447 , P3_U2409 , P3_U3108 );
and AND2_639 ( P3_U2448 , P3_U2391 , P3_U4590 );
and AND2_640 ( P3_U2449 , P3_U4344 , P3_U4522 );
and AND2_641 ( P3_U2450 , P3_U3660 , P3_U4351 );
and AND3_642 ( P3_U2451 , P3_U4608 , P3_U3102 , P3_U2412 );
and AND3_643 ( P3_U2452 , P3_U2463 , P3_U4522 , P3_U2412 );
and AND2_644 ( P3_U2453 , P3_STATE2_REG_2_ , P3_STATE2_REG_1_ );
and AND2_645 ( P3_U2454 , P3_U2380 , P3_U4323 );
and AND2_646 ( P3_U2455 , P3_U2380 , P3_U4324 );
and AND2_647 ( P3_U2456 , P3_U4556 , P3_U4607 );
and AND2_648 ( P3_U2457 , P3_U3269 , P3_U3139 );
and AND2_649 ( P3_U2458 , P3_U4652 , P3_U3269 );
and AND2_650 ( P3_U2459 , P3_U7962 , P3_U3139 );
and AND2_651 ( P3_U2460 , P3_U7962 , P3_U4652 );
and AND2_652 ( P3_U2461 , P3_U4573 , P3_U4522 );
and AND2_653 ( P3_U2462 , P3_U2412 , P3_U2449 );
and AND2_654 ( P3_U2463 , P3_U4590 , P3_U4607 );
and AND2_655 ( P3_U2464 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_INSTQUEUERD_ADDR_REG_2_ );
and AND2_656 ( P3_U2465 , P3_U2464 , P3_U4332 );
and AND2_657 ( P3_U2466 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_U3093 );
and AND2_658 ( P3_U2467 , P3_U2464 , P3_U2466 );
and AND2_659 ( P3_U2468 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_U3094 );
and AND2_660 ( P3_U2469 , P3_U2464 , P3_U2468 );
and AND2_661 ( P3_U2470 , P3_U2464 , P3_U4467 );
and AND2_662 ( P3_U2471 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_U4468 );
and AND2_663 ( P3_U2472 , P3_U2466 , P3_U3097 );
and AND2_664 ( P3_U2473 , P3_U2472 , P3_INSTQUEUERD_ADDR_REG_3_ );
and AND2_665 ( P3_U2474 , P3_U2468 , P3_U3097 );
and AND2_666 ( P3_U2475 , P3_U2474 , P3_INSTQUEUERD_ADDR_REG_3_ );
and AND2_667 ( P3_U2476 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_U4469 );
and AND2_668 ( P3_U2477 , P3_U4470 , P3_U2466 );
and AND2_669 ( P3_U2478 , P3_U4470 , P3_U2468 );
and AND2_670 ( P3_U2479 , P3_U4470 , P3_U4467 );
and AND2_671 ( P3_U2480 , P3_U4468 , P3_U3100 );
nor nor_672 ( P3_U2481 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_INSTQUEUERD_ADDR_REG_2_ );
and AND2_673 ( P3_U2482 , P3_U2466 , P3_U2481 );
and AND2_674 ( P3_U2483 , P3_U2468 , P3_U2481 );
and AND2_675 ( P3_U2484 , P3_U4469 , P3_U3100 );
and AND2_676 ( P3_U2485 , P3_U4656 , P3_U3270 );
and AND2_677 ( P3_U2486 , P3_U3271 , P3_U3182 );
and AND2_678 ( P3_U2487 , P3_U3270 , P3_U3142 );
and AND2_679 ( P3_U2488 , P3_U4657 , P3_U2487 );
and AND2_680 ( P3_U2489 , P3_U3090 , P3_U4315 );
and AND2_681 ( P3_U2490 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_U3156 );
and AND2_682 ( P3_U2491 , P3_U4644 , P3_U2487 );
and AND2_683 ( P3_U2492 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_U3128 );
and AND2_684 ( P3_U2493 , P3_U4646 , P3_U3128 );
and AND2_685 ( P3_U2494 , P3_U4645 , P3_U2487 );
and AND2_686 ( P3_U2495 , P3_U4646 , P3_INSTQUEUEWR_ADDR_REG_0_ );
and AND2_687 ( P3_U2496 , P3_U4643 , P3_U3128 );
and AND2_688 ( P3_U2497 , P3_U2496 , P3_U2487 );
and AND2_689 ( P3_U2498 , P3_U7968 , P3_U3182 );
and AND2_690 ( P3_U2499 , P3_U4658 , P3_U4657 );
and AND2_691 ( P3_U2500 , P3_U4658 , P3_U4644 );
nor nor_692 ( P3_U2501 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_INSTQUEUEWR_ADDR_REG_2_ );
and AND2_693 ( P3_U2502 , P3_U4658 , P3_U4645 );
and AND2_694 ( P3_U2503 , P3_U4658 , P3_U2496 );
and AND2_695 ( P3_U2504 , P3_U4660 , P3_U3271 );
and AND2_696 ( P3_U2505 , P3_U4644 , P3_U2485 );
and AND2_697 ( P3_U2506 , P3_U4645 , P3_U2485 );
and AND2_698 ( P3_U2507 , P3_U2496 , P3_U2485 );
and AND2_699 ( P3_U2508 , P3_U4660 , P3_U7968 );
and AND2_700 ( P3_U2509 , P3_U7965 , P3_U4656 );
and AND2_701 ( P3_U2510 , P3_U2509 , P3_U4657 );
and AND2_702 ( P3_U2511 , P3_U2509 , P3_U4644 );
and AND2_703 ( P3_U2512 , P3_U2509 , P3_U4645 );
and AND2_704 ( P3_U2513 , P3_U2509 , P3_U2496 );
and AND2_705 ( P3_U2514 , P3_U3218 , P3_U3216 );
and AND3_706 ( P3_U2515 , P3_U7970 , P3_U7969 , P3_U5485 );
and AND2_707 ( P3_U2516 , P3_U5493 , P3_U5492 );
and AND2_708 ( P3_U2517 , P3_U3246 , P3_U5526 );
and AND2_709 ( P3_U2518 , P3_U3668 , P3_U5522 );
and AND2_710 ( P3_U2519 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_U3228 );
and AND2_711 ( P3_U2520 , P3_U5543 , P3_U5548 );
and AND2_712 ( P3_U2521 , P3_U2520 , P3_U2519 );
and AND2_713 ( P3_U2522 , P3_U3093 , P3_U3228 );
and AND2_714 ( P3_U2523 , P3_U2520 , P3_U2522 );
and AND2_715 ( P3_U2524 , P3_U5558 , P3_INSTQUEUERD_ADDR_REG_0_ );
and AND2_716 ( P3_U2525 , P3_U2520 , P3_U2524 );
and AND2_717 ( P3_U2526 , P3_U5558 , P3_U3093 );
and AND2_718 ( P3_U2527 , P3_U2520 , P3_U2526 );
and AND2_719 ( P3_U2528 , P3_U5543 , P3_U3225 );
and AND2_720 ( P3_U2529 , P3_U2528 , P3_U2519 );
and AND2_721 ( P3_U2530 , P3_U2528 , P3_U2522 );
and AND2_722 ( P3_U2531 , P3_U2528 , P3_U2524 );
and AND2_723 ( P3_U2532 , P3_U2528 , P3_U2526 );
and AND2_724 ( P3_U2533 , P3_U5548 , P3_U3265 );
and AND2_725 ( P3_U2534 , P3_U2533 , P3_U2519 );
and AND2_726 ( P3_U2535 , P3_U2533 , P3_U2522 );
and AND2_727 ( P3_U2536 , P3_U2533 , P3_U2524 );
and AND2_728 ( P3_U2537 , P3_U2533 , P3_U2526 );
and AND2_729 ( P3_U2538 , P3_U3265 , P3_U3225 );
and AND2_730 ( P3_U2539 , P3_U2519 , P3_U2538 );
and AND2_731 ( P3_U2540 , P3_U2522 , P3_U2538 );
and AND2_732 ( P3_U2541 , P3_U2524 , P3_U2538 );
and AND2_733 ( P3_U2542 , P3_U2526 , P3_U2538 );
and AND2_734 ( P3_U2543 , P3_U3272 , P3_U3266 );
and AND2_735 ( P3_U2544 , P3_U2543 , P3_U2468 );
and AND2_736 ( P3_U2545 , P3_U2543 , P3_U4467 );
and AND2_737 ( P3_U2546 , P3_U2543 , P3_U4332 );
and AND2_738 ( P3_U2547 , P3_U2543 , P3_U2466 );
and AND2_739 ( P3_U2548 , P3_U8034 , P3_U3266 );
and AND2_740 ( P3_U2549 , P3_U2548 , P3_U2468 );
and AND2_741 ( P3_U2550 , P3_U2548 , P3_U4467 );
and AND2_742 ( P3_U2551 , P3_U2548 , P3_U4332 );
and AND2_743 ( P3_U2552 , P3_U2548 , P3_U2466 );
and AND2_744 ( P3_U2553 , P3_U7516 , P3_U3272 );
and AND2_745 ( P3_U2554 , P3_U2553 , P3_U2468 );
and AND2_746 ( P3_U2555 , P3_U2553 , P3_U4467 );
and AND2_747 ( P3_U2556 , P3_U2553 , P3_U4332 );
and AND2_748 ( P3_U2557 , P3_U2553 , P3_U2466 );
and AND2_749 ( P3_U2558 , P3_U7516 , P3_U8034 );
and AND2_750 ( P3_U2559 , P3_U2558 , P3_U2468 );
and AND2_751 ( P3_U2560 , P3_U2558 , P3_U4467 );
and AND2_752 ( P3_U2561 , P3_U2558 , P3_U4332 );
and AND2_753 ( P3_U2562 , P3_U2558 , P3_U2466 );
and AND2_754 ( P3_U2563 , P3_U8037 , P3_U4291 );
and AND2_755 ( P3_U2564 , P3_U2563 , P3_U2522 );
and AND2_756 ( P3_U2565 , P3_U2563 , P3_U2519 );
and AND2_757 ( P3_U2566 , P3_U2563 , P3_U2526 );
and AND2_758 ( P3_U2567 , P3_U2563 , P3_U2524 );
and AND2_759 ( P3_U2568 , P3_U8037 , P3_U3267 );
and AND2_760 ( P3_U2569 , P3_U2568 , P3_U2522 );
and AND2_761 ( P3_U2570 , P3_U2568 , P3_U2519 );
and AND2_762 ( P3_U2571 , P3_U2568 , P3_U2526 );
and AND2_763 ( P3_U2572 , P3_U2568 , P3_U2524 );
and AND2_764 ( P3_U2573 , P3_U4291 , P3_U3273 );
and AND2_765 ( P3_U2574 , P3_U2573 , P3_U2522 );
and AND2_766 ( P3_U2575 , P3_U2573 , P3_U2519 );
and AND2_767 ( P3_U2576 , P3_U2573 , P3_U2526 );
and AND2_768 ( P3_U2577 , P3_U2573 , P3_U2524 );
and AND2_769 ( P3_U2578 , P3_U3273 , P3_U3267 );
and AND2_770 ( P3_U2579 , P3_U2578 , P3_U2522 );
and AND2_771 ( P3_U2580 , P3_U2578 , P3_U2519 );
and AND2_772 ( P3_U2581 , P3_U2578 , P3_U2526 );
and AND2_773 ( P3_U2582 , P3_U2578 , P3_U2524 );
and AND2_774 ( P3_U2583 , P3_U7775 , P3_U4468 );
and AND2_775 ( P3_U2584 , P3_U7775 , P3_U2472 );
and AND2_776 ( P3_U2585 , P3_U7775 , P3_U2474 );
and AND2_777 ( P3_U2586 , P3_U7775 , P3_U4469 );
and AND2_778 ( P3_U2587 , P3_U7775 , P3_INSTQUEUERD_ADDR_REG_2_ );
and AND2_779 ( P3_U2588 , P3_U2587 , P3_U4332 );
and AND2_780 ( P3_U2589 , P3_U2587 , P3_U2466 );
and AND2_781 ( P3_U2590 , P3_U2587 , P3_U2468 );
and AND2_782 ( P3_U2591 , P3_U2587 , P3_U4467 );
and AND2_783 ( P3_U2592 , P3_U4468 , P3_U3268 );
and AND2_784 ( P3_U2593 , P3_U2472 , P3_U3268 );
and AND2_785 ( P3_U2594 , P3_U2474 , P3_U3268 );
and AND2_786 ( P3_U2595 , P3_U4469 , P3_U3268 );
and AND2_787 ( P3_U2596 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_U3268 );
and AND2_788 ( P3_U2597 , P3_U2596 , P3_U4332 );
and AND2_789 ( P3_U2598 , P3_U2596 , P3_U2466 );
and AND2_790 ( P3_U2599 , P3_U2596 , P3_U2468 );
and AND2_791 ( P3_U2600 , P3_U2596 , P3_U4467 );
and AND2_792 ( P3_U2601 , P3_U2392 , P3_U2352 );
and AND2_793 ( P3_U2602 , P3_EBX_REG_31_ , P3_U2404 );
and AND4_794 ( P3_U2603 , P3_U7360 , P3_U7358 , P3_U7359 , P3_U4133 );
and AND2_795 ( P3_U2604 , P3_U7947 , P3_U7946 );
nand NAND4_796 ( P3_U2605 , P3_U4215 , P3_U4214 , P3_U4213 , P3_U4212 );
nand NAND4_797 ( P3_U2606 , P3_U4211 , P3_U4210 , P3_U4209 , P3_U4208 );
nand NAND4_798 ( P3_U2607 , P3_U4207 , P3_U4206 , P3_U4205 , P3_U4204 );
nand NAND4_799 ( P3_U2608 , P3_U4203 , P3_U4202 , P3_U4201 , P3_U4200 );
nand NAND4_800 ( P3_U2609 , P3_U4199 , P3_U4198 , P3_U4197 , P3_U4196 );
nand NAND4_801 ( P3_U2610 , P3_U4195 , P3_U4194 , P3_U4193 , P3_U4192 );
nand NAND4_802 ( P3_U2611 , P3_U4191 , P3_U4190 , P3_U4189 , P3_U4188 );
nand NAND4_803 ( P3_U2612 , P3_U4187 , P3_U4186 , P3_U4185 , P3_U4184 );
nand NAND4_804 ( P3_U2613 , P3_U4279 , P3_U4278 , P3_U4277 , P3_U4276 );
nand NAND4_805 ( P3_U2614 , P3_U4275 , P3_U4274 , P3_U4273 , P3_U4272 );
nand NAND4_806 ( P3_U2615 , P3_U4271 , P3_U4270 , P3_U4269 , P3_U4268 );
nand NAND4_807 ( P3_U2616 , P3_U4267 , P3_U4266 , P3_U4265 , P3_U4264 );
nand NAND4_808 ( P3_U2617 , P3_U4263 , P3_U4262 , P3_U4261 , P3_U4260 );
nand NAND4_809 ( P3_U2618 , P3_U4259 , P3_U4258 , P3_U4257 , P3_U4256 );
nand NAND4_810 ( P3_U2619 , P3_U4255 , P3_U4254 , P3_U4253 , P3_U4252 );
nand NAND4_811 ( P3_U2620 , P3_U4251 , P3_U4250 , P3_U4249 , P3_U4248 );
nand NAND4_812 ( P3_U2621 , P3_U4183 , P3_U4182 , P3_U4181 , P3_U4180 );
nand NAND4_813 ( P3_U2622 , P3_U4179 , P3_U4178 , P3_U4177 , P3_U4176 );
nand NAND4_814 ( P3_U2623 , P3_U4175 , P3_U4174 , P3_U4173 , P3_U4172 );
nand NAND4_815 ( P3_U2624 , P3_U4171 , P3_U4170 , P3_U4169 , P3_U4168 );
nand NAND4_816 ( P3_U2625 , P3_U4167 , P3_U4166 , P3_U4165 , P3_U4164 );
nand NAND4_817 ( P3_U2626 , P3_U4163 , P3_U4162 , P3_U4161 , P3_U4160 );
nand NAND4_818 ( P3_U2627 , P3_U4159 , P3_U4158 , P3_U4157 , P3_U4156 );
nand NAND4_819 ( P3_U2628 , P3_U4155 , P3_U4154 , P3_U4153 , P3_U4152 );
and AND2_820 ( P3_U2629 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_U3207 );
not NOT1_821 ( P3_U2630 , U209 );
not NOT1_822 ( P3_U2631 , P3_STATEBS16_REG );
and AND2_823 ( P3_U2632 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_U3207 );
nand NAND2_824 ( P3_U2633 , P3_U7937 , P3_U7383 );
nand NAND2_825 ( P3_U2634 , P3_U7382 , P3_U7381 );
nand NAND3_826 ( P3_U2635 , P3_U8025 , P3_U8024 , P3_U4335 );
nand NAND3_827 ( P3_U2636 , P3_U8021 , P3_U8020 , P3_U4335 );
nand NAND2_828 ( P3_U2637 , P3_U7370 , P3_U7369 );
nand NAND3_829 ( P3_U2638 , P3_U8013 , P3_U8012 , P3_U4327 );
nand NAND3_830 ( P3_U2639 , P3_U8003 , P3_U8002 , P3_U4327 );
and AND2_831 ( P3_U2640 , P3_U7357 , P3_U7907 );
nand NAND5_832 ( P3_U2641 , P3_U7352 , P3_U7351 , P3_U4129 , P3_U7354 , P3_U4130 );
nand NAND5_833 ( P3_U2642 , P3_U7344 , P3_U7343 , P3_U4126 , P3_U7346 , P3_U4127 );
nand NAND5_834 ( P3_U2643 , P3_U7336 , P3_U7335 , P3_U4123 , P3_U7338 , P3_U4124 );
nand NAND5_835 ( P3_U2644 , P3_U7328 , P3_U7327 , P3_U4120 , P3_U7330 , P3_U4121 );
nand NAND5_836 ( P3_U2645 , P3_U7320 , P3_U7319 , P3_U4117 , P3_U7322 , P3_U4118 );
nand NAND5_837 ( P3_U2646 , P3_U7312 , P3_U7311 , P3_U4114 , P3_U7314 , P3_U4115 );
nand NAND5_838 ( P3_U2647 , P3_U7304 , P3_U7303 , P3_U4111 , P3_U7306 , P3_U4112 );
nand NAND5_839 ( P3_U2648 , P3_U7296 , P3_U7295 , P3_U4108 , P3_U7298 , P3_U4109 );
nand NAND5_840 ( P3_U2649 , P3_U7288 , P3_U7287 , P3_U4105 , P3_U7290 , P3_U4106 );
nand NAND5_841 ( P3_U2650 , P3_U7280 , P3_U7279 , P3_U4102 , P3_U7282 , P3_U4103 );
nand NAND5_842 ( P3_U2651 , P3_U7272 , P3_U7271 , P3_U4099 , P3_U7274 , P3_U4100 );
nand NAND5_843 ( P3_U2652 , P3_U7264 , P3_U7263 , P3_U4096 , P3_U7266 , P3_U4097 );
nand NAND5_844 ( P3_U2653 , P3_U7256 , P3_U7255 , P3_U4093 , P3_U7258 , P3_U4094 );
nand NAND5_845 ( P3_U2654 , P3_U7248 , P3_U7247 , P3_U4090 , P3_U7250 , P3_U4091 );
nand NAND5_846 ( P3_U2655 , P3_U7240 , P3_U7239 , P3_U4087 , P3_U7242 , P3_U4088 );
nand NAND5_847 ( P3_U2656 , P3_U7232 , P3_U7231 , P3_U4084 , P3_U7234 , P3_U4085 );
nand NAND5_848 ( P3_U2657 , P3_U7224 , P3_U7223 , P3_U4081 , P3_U7226 , P3_U4082 );
nand NAND5_849 ( P3_U2658 , P3_U7216 , P3_U7215 , P3_U4078 , P3_U7218 , P3_U4079 );
nand NAND5_850 ( P3_U2659 , P3_U7208 , P3_U7207 , P3_U4075 , P3_U7210 , P3_U4076 );
nand NAND5_851 ( P3_U2660 , P3_U7200 , P3_U7199 , P3_U4072 , P3_U7202 , P3_U4073 );
nand NAND5_852 ( P3_U2661 , P3_U7192 , P3_U7191 , P3_U4069 , P3_U7194 , P3_U4070 );
nand NAND5_853 ( P3_U2662 , P3_U7184 , P3_U7183 , P3_U4066 , P3_U7186 , P3_U4067 );
nand NAND5_854 ( P3_U2663 , P3_U7176 , P3_U7175 , P3_U4063 , P3_U7178 , P3_U4064 );
nand NAND5_855 ( P3_U2664 , P3_U7168 , P3_U7167 , P3_U4060 , P3_U7170 , P3_U4061 );
nand NAND5_856 ( P3_U2665 , P3_U7160 , P3_U7159 , P3_U4057 , P3_U7162 , P3_U4058 );
nand NAND2_857 ( P3_U2666 , P3_U4056 , P3_U4054 );
nand NAND2_858 ( P3_U2667 , P3_U4051 , P3_U4049 );
nand NAND5_859 ( P3_U2668 , P3_U7129 , P3_U4043 , P3_U7132 , P3_U7133 , P3_U4045 );
nand NAND5_860 ( P3_U2669 , P3_U7119 , P3_U4039 , P3_U7122 , P3_U7123 , P3_U4041 );
nand NAND5_861 ( P3_U2670 , P3_U7109 , P3_U4035 , P3_U7112 , P3_U7113 , P3_U4037 );
nand NAND5_862 ( P3_U2671 , P3_U7099 , P3_U4031 , P3_U7102 , P3_U7103 , P3_U4033 );
nand NAND2_863 ( P3_U2672 , P3_U7092 , P3_U7091 );
nand NAND3_864 ( P3_U2673 , P3_U7090 , P3_U7088 , P3_U7089 );
nand NAND3_865 ( P3_U2674 , P3_U7087 , P3_U7085 , P3_U7086 );
nand NAND3_866 ( P3_U2675 , P3_U7084 , P3_U7082 , P3_U7083 );
nand NAND3_867 ( P3_U2676 , P3_U7081 , P3_U7079 , P3_U7080 );
nand NAND3_868 ( P3_U2677 , P3_U7078 , P3_U7076 , P3_U7077 );
nand NAND3_869 ( P3_U2678 , P3_U7075 , P3_U7073 , P3_U7074 );
nand NAND3_870 ( P3_U2679 , P3_U7072 , P3_U7070 , P3_U7071 );
nand NAND3_871 ( P3_U2680 , P3_U7069 , P3_U7067 , P3_U7068 );
nand NAND3_872 ( P3_U2681 , P3_U7066 , P3_U7064 , P3_U7065 );
nand NAND3_873 ( P3_U2682 , P3_U7063 , P3_U7061 , P3_U7062 );
nand NAND3_874 ( P3_U2683 , P3_U7060 , P3_U7058 , P3_U7059 );
nand NAND3_875 ( P3_U2684 , P3_U7057 , P3_U7055 , P3_U7056 );
nand NAND3_876 ( P3_U2685 , P3_U7054 , P3_U7052 , P3_U7053 );
nand NAND3_877 ( P3_U2686 , P3_U7051 , P3_U7049 , P3_U7050 );
nand NAND3_878 ( P3_U2687 , P3_U7048 , P3_U7046 , P3_U7047 );
nand NAND3_879 ( P3_U2688 , P3_U7045 , P3_U7043 , P3_U7044 );
nand NAND3_880 ( P3_U2689 , P3_U7042 , P3_U7040 , P3_U7041 );
nand NAND3_881 ( P3_U2690 , P3_U7039 , P3_U7037 , P3_U7038 );
nand NAND3_882 ( P3_U2691 , P3_U7036 , P3_U7034 , P3_U7035 );
nand NAND3_883 ( P3_U2692 , P3_U7033 , P3_U7031 , P3_U7032 );
nand NAND3_884 ( P3_U2693 , P3_U7030 , P3_U7028 , P3_U7029 );
nand NAND3_885 ( P3_U2694 , P3_U7026 , P3_U7025 , P3_U7027 );
nand NAND3_886 ( P3_U2695 , P3_U7023 , P3_U7022 , P3_U7024 );
nand NAND3_887 ( P3_U2696 , P3_U7020 , P3_U7019 , P3_U7021 );
nand NAND3_888 ( P3_U2697 , P3_U7017 , P3_U7016 , P3_U7018 );
nand NAND3_889 ( P3_U2698 , P3_U7014 , P3_U7013 , P3_U7015 );
nand NAND3_890 ( P3_U2699 , P3_U7011 , P3_U7010 , P3_U7012 );
nand NAND3_891 ( P3_U2700 , P3_U7008 , P3_U7007 , P3_U7009 );
nand NAND3_892 ( P3_U2701 , P3_U7005 , P3_U7004 , P3_U7006 );
nand NAND3_893 ( P3_U2702 , P3_U7002 , P3_U7001 , P3_U7003 );
nand NAND3_894 ( P3_U2703 , P3_U6999 , P3_U6998 , P3_U7000 );
nand NAND3_895 ( P3_U2704 , P3_U6995 , P3_U6993 , P3_U6994 );
nand NAND5_896 ( P3_U2705 , P3_U6989 , P3_U6988 , P3_U6992 , P3_U6990 , P3_U6991 );
nand NAND5_897 ( P3_U2706 , P3_U6984 , P3_U6983 , P3_U6987 , P3_U6985 , P3_U6986 );
nand NAND5_898 ( P3_U2707 , P3_U6979 , P3_U6978 , P3_U6982 , P3_U6980 , P3_U6981 );
nand NAND4_899 ( P3_U2708 , P3_U6974 , P3_U6973 , P3_U4029 , P3_U6976 );
nand NAND4_900 ( P3_U2709 , P3_U6969 , P3_U6968 , P3_U4028 , P3_U6971 );
nand NAND4_901 ( P3_U2710 , P3_U6964 , P3_U6963 , P3_U4027 , P3_U6966 );
nand NAND4_902 ( P3_U2711 , P3_U6959 , P3_U6958 , P3_U4026 , P3_U6961 );
nand NAND4_903 ( P3_U2712 , P3_U6954 , P3_U6953 , P3_U4025 , P3_U6956 );
nand NAND4_904 ( P3_U2713 , P3_U6949 , P3_U6948 , P3_U4024 , P3_U6951 );
nand NAND4_905 ( P3_U2714 , P3_U6944 , P3_U6943 , P3_U4023 , P3_U6946 );
nand NAND4_906 ( P3_U2715 , P3_U6939 , P3_U6938 , P3_U4022 , P3_U6941 );
nand NAND4_907 ( P3_U2716 , P3_U6934 , P3_U6933 , P3_U4021 , P3_U6936 );
nand NAND4_908 ( P3_U2717 , P3_U6929 , P3_U6928 , P3_U4020 , P3_U6931 );
nand NAND4_909 ( P3_U2718 , P3_U6924 , P3_U6923 , P3_U4019 , P3_U6926 );
nand NAND4_910 ( P3_U2719 , P3_U6919 , P3_U6918 , P3_U4018 , P3_U6921 );
nand NAND3_911 ( P3_U2720 , P3_U6914 , P3_U4017 , P3_U6916 );
nand NAND3_912 ( P3_U2721 , P3_U6910 , P3_U4016 , P3_U6912 );
nand NAND3_913 ( P3_U2722 , P3_U6906 , P3_U4015 , P3_U6908 );
nand NAND3_914 ( P3_U2723 , P3_U6903 , P3_U6902 , P3_U4014 );
nand NAND3_915 ( P3_U2724 , P3_U6899 , P3_U6898 , P3_U4013 );
nand NAND3_916 ( P3_U2725 , P3_U6895 , P3_U6894 , P3_U4012 );
nand NAND3_917 ( P3_U2726 , P3_U6891 , P3_U6890 , P3_U4011 );
nand NAND3_918 ( P3_U2727 , P3_U6887 , P3_U6886 , P3_U4010 );
nand NAND3_919 ( P3_U2728 , P3_U6883 , P3_U6882 , P3_U4009 );
nand NAND3_920 ( P3_U2729 , P3_U6879 , P3_U6878 , P3_U4008 );
nand NAND3_921 ( P3_U2730 , P3_U6875 , P3_U6874 , P3_U4007 );
nand NAND3_922 ( P3_U2731 , P3_U6871 , P3_U6870 , P3_U4006 );
nand NAND3_923 ( P3_U2732 , P3_U6867 , P3_U6866 , P3_U4005 );
nand NAND3_924 ( P3_U2733 , P3_U6863 , P3_U6862 , P3_U4004 );
nand NAND3_925 ( P3_U2734 , P3_U6859 , P3_U6858 , P3_U4003 );
nand NAND3_926 ( P3_U2735 , P3_U6855 , P3_U6854 , P3_U4002 );
and AND2_927 ( P3_U2736 , P3_DATAO_REG_31_ , P3_U6759 );
nand NAND2_928 ( P3_U2737 , P3_U4001 , P3_U6850 );
nand NAND2_929 ( P3_U2738 , P3_U4000 , P3_U6847 );
nand NAND2_930 ( P3_U2739 , P3_U3999 , P3_U6844 );
nand NAND2_931 ( P3_U2740 , P3_U3998 , P3_U6841 );
nand NAND2_932 ( P3_U2741 , P3_U3997 , P3_U6838 );
nand NAND2_933 ( P3_U2742 , P3_U3996 , P3_U6835 );
nand NAND2_934 ( P3_U2743 , P3_U3995 , P3_U6832 );
nand NAND2_935 ( P3_U2744 , P3_U3994 , P3_U6829 );
nand NAND2_936 ( P3_U2745 , P3_U3993 , P3_U6826 );
nand NAND2_937 ( P3_U2746 , P3_U3992 , P3_U6823 );
nand NAND2_938 ( P3_U2747 , P3_U3991 , P3_U6820 );
nand NAND2_939 ( P3_U2748 , P3_U3990 , P3_U6817 );
nand NAND2_940 ( P3_U2749 , P3_U3989 , P3_U6814 );
nand NAND2_941 ( P3_U2750 , P3_U3988 , P3_U6811 );
nand NAND2_942 ( P3_U2751 , P3_U3987 , P3_U6808 );
nand NAND3_943 ( P3_U2752 , P3_U6806 , P3_U6805 , P3_U6807 );
nand NAND3_944 ( P3_U2753 , P3_U6803 , P3_U6802 , P3_U6804 );
nand NAND3_945 ( P3_U2754 , P3_U6800 , P3_U6799 , P3_U6801 );
nand NAND3_946 ( P3_U2755 , P3_U6797 , P3_U6796 , P3_U6798 );
nand NAND3_947 ( P3_U2756 , P3_U6794 , P3_U6793 , P3_U6795 );
nand NAND3_948 ( P3_U2757 , P3_U6791 , P3_U6790 , P3_U6792 );
nand NAND3_949 ( P3_U2758 , P3_U6788 , P3_U6787 , P3_U6789 );
nand NAND3_950 ( P3_U2759 , P3_U6785 , P3_U6784 , P3_U6786 );
nand NAND3_951 ( P3_U2760 , P3_U6782 , P3_U6781 , P3_U6783 );
nand NAND3_952 ( P3_U2761 , P3_U6779 , P3_U6778 , P3_U6780 );
nand NAND3_953 ( P3_U2762 , P3_U6776 , P3_U6775 , P3_U6777 );
nand NAND3_954 ( P3_U2763 , P3_U6773 , P3_U6772 , P3_U6774 );
nand NAND3_955 ( P3_U2764 , P3_U6770 , P3_U6769 , P3_U6771 );
nand NAND3_956 ( P3_U2765 , P3_U6767 , P3_U6766 , P3_U6768 );
nand NAND3_957 ( P3_U2766 , P3_U6764 , P3_U6763 , P3_U6765 );
nand NAND3_958 ( P3_U2767 , P3_U6761 , P3_U6760 , P3_U6762 );
nand NAND3_959 ( P3_U2768 , P3_U6755 , P3_U6754 , P3_U6756 );
nand NAND3_960 ( P3_U2769 , P3_U6752 , P3_U6751 , P3_U6753 );
nand NAND3_961 ( P3_U2770 , P3_U6749 , P3_U6748 , P3_U6750 );
nand NAND3_962 ( P3_U2771 , P3_U6746 , P3_U6745 , P3_U6747 );
nand NAND3_963 ( P3_U2772 , P3_U6743 , P3_U6742 , P3_U6744 );
nand NAND3_964 ( P3_U2773 , P3_U6740 , P3_U6739 , P3_U6741 );
nand NAND3_965 ( P3_U2774 , P3_U6737 , P3_U6736 , P3_U6738 );
nand NAND3_966 ( P3_U2775 , P3_U6734 , P3_U6733 , P3_U6735 );
nand NAND3_967 ( P3_U2776 , P3_U6731 , P3_U6730 , P3_U6732 );
nand NAND3_968 ( P3_U2777 , P3_U6728 , P3_U6727 , P3_U6729 );
nand NAND3_969 ( P3_U2778 , P3_U6725 , P3_U6724 , P3_U6726 );
nand NAND3_970 ( P3_U2779 , P3_U6722 , P3_U6721 , P3_U6723 );
nand NAND3_971 ( P3_U2780 , P3_U6719 , P3_U6718 , P3_U6720 );
nand NAND3_972 ( P3_U2781 , P3_U6716 , P3_U6715 , P3_U6717 );
nand NAND3_973 ( P3_U2782 , P3_U6713 , P3_U6712 , P3_U6714 );
nand NAND3_974 ( P3_U2783 , P3_U6710 , P3_U6709 , P3_U6711 );
nand NAND3_975 ( P3_U2784 , P3_U6707 , P3_U6706 , P3_U6708 );
nand NAND3_976 ( P3_U2785 , P3_U6704 , P3_U6703 , P3_U6705 );
nand NAND3_977 ( P3_U2786 , P3_U6701 , P3_U6700 , P3_U6702 );
nand NAND3_978 ( P3_U2787 , P3_U6698 , P3_U6697 , P3_U6699 );
nand NAND3_979 ( P3_U2788 , P3_U6695 , P3_U6694 , P3_U6696 );
nand NAND3_980 ( P3_U2789 , P3_U6692 , P3_U6691 , P3_U6693 );
nand NAND3_981 ( P3_U2790 , P3_U6689 , P3_U6688 , P3_U6690 );
nand NAND3_982 ( P3_U2791 , P3_U6686 , P3_U6685 , P3_U6687 );
nand NAND3_983 ( P3_U2792 , P3_U6683 , P3_U6682 , P3_U6684 );
nand NAND3_984 ( P3_U2793 , P3_U6680 , P3_U6679 , P3_U6681 );
nand NAND3_985 ( P3_U2794 , P3_U6677 , P3_U6676 , P3_U6678 );
nand NAND3_986 ( P3_U2795 , P3_U6674 , P3_U6673 , P3_U6675 );
nand NAND3_987 ( P3_U2796 , P3_U6671 , P3_U6670 , P3_U6672 );
nand NAND3_988 ( P3_U2797 , P3_U6668 , P3_U6667 , P3_U6669 );
nand NAND3_989 ( P3_U2798 , P3_U6665 , P3_U6664 , P3_U6666 );
nand NAND5_990 ( P3_U2799 , P3_U6656 , P3_U6654 , P3_U6655 , P3_U6653 , P3_U3985 );
nand NAND5_991 ( P3_U2800 , P3_U6648 , P3_U6647 , P3_U6646 , P3_U6645 , P3_U3984 );
nand NAND5_992 ( P3_U2801 , P3_U6640 , P3_U6639 , P3_U6638 , P3_U6637 , P3_U3983 );
nand NAND5_993 ( P3_U2802 , P3_U6632 , P3_U6631 , P3_U6630 , P3_U6629 , P3_U3982 );
nand NAND5_994 ( P3_U2803 , P3_U6622 , P3_U6624 , P3_U6621 , P3_U6623 , P3_U3981 );
nand NAND5_995 ( P3_U2804 , P3_U6614 , P3_U6616 , P3_U6613 , P3_U6615 , P3_U3980 );
nand NAND5_996 ( P3_U2805 , P3_U6606 , P3_U6608 , P3_U6605 , P3_U6607 , P3_U3979 );
nand NAND5_997 ( P3_U2806 , P3_U6598 , P3_U6600 , P3_U6597 , P3_U6599 , P3_U3978 );
nand NAND5_998 ( P3_U2807 , P3_U6590 , P3_U6589 , P3_U6592 , P3_U6591 , P3_U3977 );
nand NAND5_999 ( P3_U2808 , P3_U6582 , P3_U6581 , P3_U6584 , P3_U6583 , P3_U3976 );
nand NAND5_1000 ( P3_U2809 , P3_U6574 , P3_U6573 , P3_U6575 , P3_U3975 , P3_U6576 );
nand NAND5_1001 ( P3_U2810 , P3_U6566 , P3_U6565 , P3_U6567 , P3_U3974 , P3_U6568 );
nand NAND5_1002 ( P3_U2811 , P3_U6558 , P3_U6557 , P3_U6559 , P3_U6560 , P3_U3973 );
nand NAND5_1003 ( P3_U2812 , P3_U6550 , P3_U6549 , P3_U6551 , P3_U6552 , P3_U3972 );
nand NAND5_1004 ( P3_U2813 , P3_U6542 , P3_U6541 , P3_U6543 , P3_U6544 , P3_U3971 );
nand NAND5_1005 ( P3_U2814 , P3_U6534 , P3_U6533 , P3_U6535 , P3_U6536 , P3_U3970 );
nand NAND5_1006 ( P3_U2815 , P3_U6526 , P3_U6525 , P3_U6528 , P3_U6527 , P3_U3969 );
nand NAND5_1007 ( P3_U2816 , P3_U6518 , P3_U6517 , P3_U6520 , P3_U6519 , P3_U3968 );
nand NAND5_1008 ( P3_U2817 , P3_U6510 , P3_U6509 , P3_U6512 , P3_U6511 , P3_U3967 );
nand NAND5_1009 ( P3_U2818 , P3_U6502 , P3_U6501 , P3_U6504 , P3_U6503 , P3_U3966 );
nand NAND5_1010 ( P3_U2819 , P3_U6494 , P3_U6493 , P3_U6495 , P3_U6496 , P3_U3965 );
nand NAND5_1011 ( P3_U2820 , P3_U6486 , P3_U6485 , P3_U6487 , P3_U6488 , P3_U3964 );
nand NAND5_1012 ( P3_U2821 , P3_U6478 , P3_U6477 , P3_U6480 , P3_U6479 , P3_U3963 );
nand NAND5_1013 ( P3_U2822 , P3_U6470 , P3_U6469 , P3_U6472 , P3_U6471 , P3_U3962 );
nand NAND5_1014 ( P3_U2823 , P3_U6462 , P3_U6461 , P3_U6464 , P3_U6463 , P3_U3961 );
nand NAND5_1015 ( P3_U2824 , P3_U6454 , P3_U6453 , P3_U6456 , P3_U6455 , P3_U3960 );
nand NAND5_1016 ( P3_U2825 , P3_U6446 , P3_U6445 , P3_U6448 , P3_U6447 , P3_U3959 );
nand NAND5_1017 ( P3_U2826 , P3_U6438 , P3_U6437 , P3_U6439 , P3_U6440 , P3_U3958 );
nand NAND5_1018 ( P3_U2827 , P3_U6432 , P3_U6431 , P3_U6430 , P3_U6429 , P3_U3957 );
nand NAND5_1019 ( P3_U2828 , P3_U6424 , P3_U6423 , P3_U6422 , P3_U6421 , P3_U3956 );
nand NAND5_1020 ( P3_U2829 , P3_U6416 , P3_U6415 , P3_U6414 , P3_U6413 , P3_U3955 );
nand NAND5_1021 ( P3_U2830 , P3_U6408 , P3_U6407 , P3_U6406 , P3_U6405 , P3_U3954 );
and AND2_1022 ( P3_U2831 , P3_U6396 , P3_U7906 );
nand NAND3_1023 ( P3_U2832 , P3_U6375 , P3_U6373 , P3_U6374 );
nand NAND3_1024 ( P3_U2833 , P3_U6351 , P3_U6349 , P3_U6350 );
nand NAND3_1025 ( P3_U2834 , P3_U6327 , P3_U6325 , P3_U6326 );
nand NAND3_1026 ( P3_U2835 , P3_U6303 , P3_U6301 , P3_U6302 );
nand NAND3_1027 ( P3_U2836 , P3_U6279 , P3_U6277 , P3_U6278 );
nand NAND2_1028 ( P3_U2837 , P3_U3893 , P3_U6254 );
nand NAND2_1029 ( P3_U2838 , P3_U3883 , P3_U6230 );
nand NAND2_1030 ( P3_U2839 , P3_U3873 , P3_U6206 );
nand NAND2_1031 ( P3_U2840 , P3_U3863 , P3_U6182 );
nand NAND2_1032 ( P3_U2841 , P3_U3853 , P3_U6158 );
nand NAND2_1033 ( P3_U2842 , P3_U3845 , P3_U6134 );
nand NAND3_1034 ( P3_U2843 , P3_U6111 , P3_U6109 , P3_U6110 );
nand NAND3_1035 ( P3_U2844 , P3_U6087 , P3_U6085 , P3_U6086 );
nand NAND3_1036 ( P3_U2845 , P3_U6063 , P3_U6061 , P3_U6062 );
nand NAND3_1037 ( P3_U2846 , P3_U6039 , P3_U6037 , P3_U6038 );
nand NAND2_1038 ( P3_U2847 , P3_U3811 , P3_U6014 );
nand NAND2_1039 ( P3_U2848 , P3_U3803 , P3_U5990 );
nand NAND3_1040 ( P3_U2849 , P3_U5967 , P3_U5965 , P3_U5966 );
nand NAND3_1041 ( P3_U2850 , P3_U5943 , P3_U5941 , P3_U5942 );
nand NAND3_1042 ( P3_U2851 , P3_U5919 , P3_U5917 , P3_U5918 );
nand NAND3_1043 ( P3_U2852 , P3_U5895 , P3_U5893 , P3_U5894 );
nand NAND3_1044 ( P3_U2853 , P3_U5871 , P3_U5869 , P3_U5870 );
nand NAND3_1045 ( P3_U2854 , P3_U5847 , P3_U5845 , P3_U5846 );
nand NAND3_1046 ( P3_U2855 , P3_U5823 , P3_U5821 , P3_U5822 );
nand NAND3_1047 ( P3_U2856 , P3_U5799 , P3_U5797 , P3_U5798 );
nand NAND3_1048 ( P3_U2857 , P3_U5775 , P3_U5773 , P3_U5774 );
nand NAND3_1049 ( P3_U2858 , P3_U5751 , P3_U5749 , P3_U5750 );
nand NAND3_1050 ( P3_U2859 , P3_U5727 , P3_U5725 , P3_U5726 );
nand NAND3_1051 ( P3_U2860 , P3_U5703 , P3_U5701 , P3_U5702 );
nand NAND3_1052 ( P3_U2861 , P3_U5679 , P3_U5677 , P3_U5678 );
nand NAND3_1053 ( P3_U2862 , P3_U5654 , P3_U5653 , P3_U5655 );
nand NAND2_1054 ( P3_U2863 , P3_U5616 , P3_U5615 );
nand NAND2_1055 ( P3_U2864 , P3_U5610 , P3_U5609 );
nand NAND2_1056 ( P3_U2865 , P3_U5599 , P3_U5598 );
nand NAND2_1057 ( P3_U2866 , P3_U5591 , P3_U5590 );
and AND2_1058 ( P3_U2867 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_U5579 );
nand NAND2_1059 ( P3_U2868 , P3_U3651 , P3_U5482 );
nand NAND2_1060 ( P3_U2869 , P3_U3649 , P3_U5477 );
nand NAND2_1061 ( P3_U2870 , P3_U3647 , P3_U5472 );
nand NAND2_1062 ( P3_U2871 , P3_U3645 , P3_U5467 );
nand NAND2_1063 ( P3_U2872 , P3_U3643 , P3_U5462 );
nand NAND2_1064 ( P3_U2873 , P3_U3641 , P3_U5457 );
nand NAND2_1065 ( P3_U2874 , P3_U3639 , P3_U5452 );
nand NAND2_1066 ( P3_U2875 , P3_U3637 , P3_U5447 );
nand NAND2_1067 ( P3_U2876 , P3_U3633 , P3_U5432 );
nand NAND2_1068 ( P3_U2877 , P3_U3631 , P3_U5427 );
nand NAND2_1069 ( P3_U2878 , P3_U3629 , P3_U5422 );
nand NAND2_1070 ( P3_U2879 , P3_U3627 , P3_U5417 );
nand NAND2_1071 ( P3_U2880 , P3_U3625 , P3_U5412 );
nand NAND2_1072 ( P3_U2881 , P3_U3623 , P3_U5407 );
nand NAND2_1073 ( P3_U2882 , P3_U3621 , P3_U5402 );
nand NAND2_1074 ( P3_U2883 , P3_U3619 , P3_U5397 );
nand NAND2_1075 ( P3_U2884 , P3_U3615 , P3_U5381 );
nand NAND2_1076 ( P3_U2885 , P3_U3613 , P3_U5376 );
nand NAND2_1077 ( P3_U2886 , P3_U3611 , P3_U5371 );
nand NAND2_1078 ( P3_U2887 , P3_U3609 , P3_U5366 );
nand NAND2_1079 ( P3_U2888 , P3_U3607 , P3_U5361 );
nand NAND2_1080 ( P3_U2889 , P3_U3605 , P3_U5356 );
nand NAND2_1081 ( P3_U2890 , P3_U3603 , P3_U5351 );
nand NAND2_1082 ( P3_U2891 , P3_U3601 , P3_U5346 );
nand NAND2_1083 ( P3_U2892 , P3_U3598 , P3_U5330 );
nand NAND2_1084 ( P3_U2893 , P3_U3596 , P3_U5325 );
nand NAND2_1085 ( P3_U2894 , P3_U3594 , P3_U5320 );
nand NAND2_1086 ( P3_U2895 , P3_U3592 , P3_U5315 );
nand NAND2_1087 ( P3_U2896 , P3_U3590 , P3_U5310 );
nand NAND2_1088 ( P3_U2897 , P3_U3588 , P3_U5305 );
nand NAND2_1089 ( P3_U2898 , P3_U3586 , P3_U5300 );
nand NAND2_1090 ( P3_U2899 , P3_U3584 , P3_U5295 );
nand NAND2_1091 ( P3_U2900 , P3_U3580 , P3_U5279 );
nand NAND2_1092 ( P3_U2901 , P3_U3578 , P3_U5274 );
nand NAND2_1093 ( P3_U2902 , P3_U3576 , P3_U5269 );
nand NAND2_1094 ( P3_U2903 , P3_U3574 , P3_U5264 );
nand NAND2_1095 ( P3_U2904 , P3_U3572 , P3_U5259 );
nand NAND2_1096 ( P3_U2905 , P3_U3570 , P3_U5254 );
nand NAND2_1097 ( P3_U2906 , P3_U3568 , P3_U5249 );
nand NAND2_1098 ( P3_U2907 , P3_U3566 , P3_U5244 );
nand NAND3_1099 ( P3_U2908 , P3_U5229 , P3_U3562 , P3_U5228 );
nand NAND3_1100 ( P3_U2909 , P3_U5224 , P3_U3560 , P3_U5223 );
nand NAND3_1101 ( P3_U2910 , P3_U5219 , P3_U3558 , P3_U5218 );
nand NAND3_1102 ( P3_U2911 , P3_U5214 , P3_U3556 , P3_U5213 );
nand NAND3_1103 ( P3_U2912 , P3_U5209 , P3_U3554 , P3_U5208 );
nand NAND3_1104 ( P3_U2913 , P3_U5204 , P3_U3552 , P3_U5203 );
nand NAND3_1105 ( P3_U2914 , P3_U5199 , P3_U3550 , P3_U5198 );
nand NAND3_1106 ( P3_U2915 , P3_U5194 , P3_U3548 , P3_U5193 );
nand NAND3_1107 ( P3_U2916 , P3_U5177 , P3_U3544 , P3_U5176 );
nand NAND3_1108 ( P3_U2917 , P3_U5172 , P3_U3542 , P3_U5171 );
nand NAND3_1109 ( P3_U2918 , P3_U5167 , P3_U3540 , P3_U5166 );
nand NAND3_1110 ( P3_U2919 , P3_U5162 , P3_U3538 , P3_U5161 );
nand NAND3_1111 ( P3_U2920 , P3_U5157 , P3_U3536 , P3_U5156 );
nand NAND3_1112 ( P3_U2921 , P3_U5152 , P3_U3534 , P3_U5151 );
nand NAND3_1113 ( P3_U2922 , P3_U5147 , P3_U3532 , P3_U5146 );
nand NAND3_1114 ( P3_U2923 , P3_U5142 , P3_U3530 , P3_U5141 );
nand NAND3_1115 ( P3_U2924 , P3_U5125 , P3_U3526 , P3_U5124 );
nand NAND3_1116 ( P3_U2925 , P3_U5120 , P3_U3524 , P3_U5119 );
nand NAND3_1117 ( P3_U2926 , P3_U5115 , P3_U3522 , P3_U5114 );
nand NAND3_1118 ( P3_U2927 , P3_U5110 , P3_U3520 , P3_U5109 );
nand NAND3_1119 ( P3_U2928 , P3_U5105 , P3_U3518 , P3_U5104 );
nand NAND3_1120 ( P3_U2929 , P3_U5100 , P3_U3516 , P3_U5099 );
nand NAND3_1121 ( P3_U2930 , P3_U5095 , P3_U3514 , P3_U5094 );
nand NAND3_1122 ( P3_U2931 , P3_U5090 , P3_U3512 , P3_U5089 );
nand NAND3_1123 ( P3_U2932 , P3_U5076 , P3_U3509 , P3_U5075 );
nand NAND3_1124 ( P3_U2933 , P3_U5071 , P3_U3507 , P3_U5070 );
nand NAND3_1125 ( P3_U2934 , P3_U5066 , P3_U3505 , P3_U5065 );
nand NAND3_1126 ( P3_U2935 , P3_U5061 , P3_U3503 , P3_U5060 );
nand NAND3_1127 ( P3_U2936 , P3_U5056 , P3_U3501 , P3_U5055 );
nand NAND3_1128 ( P3_U2937 , P3_U5051 , P3_U3499 , P3_U5050 );
nand NAND3_1129 ( P3_U2938 , P3_U5046 , P3_U3497 , P3_U5045 );
nand NAND3_1130 ( P3_U2939 , P3_U5041 , P3_U3495 , P3_U5040 );
nand NAND3_1131 ( P3_U2940 , P3_U5025 , P3_U3492 , P3_U5024 );
nand NAND3_1132 ( P3_U2941 , P3_U5020 , P3_U3490 , P3_U5019 );
nand NAND3_1133 ( P3_U2942 , P3_U5015 , P3_U3488 , P3_U5014 );
nand NAND3_1134 ( P3_U2943 , P3_U5010 , P3_U3486 , P3_U5009 );
nand NAND3_1135 ( P3_U2944 , P3_U5005 , P3_U3484 , P3_U5004 );
nand NAND3_1136 ( P3_U2945 , P3_U5000 , P3_U3482 , P3_U4999 );
nand NAND3_1137 ( P3_U2946 , P3_U4995 , P3_U3480 , P3_U4994 );
nand NAND3_1138 ( P3_U2947 , P3_U4990 , P3_U3478 , P3_U4989 );
nand NAND3_1139 ( P3_U2948 , P3_U4973 , P3_U3474 , P3_U4972 );
nand NAND3_1140 ( P3_U2949 , P3_U4968 , P3_U3472 , P3_U4967 );
nand NAND3_1141 ( P3_U2950 , P3_U4963 , P3_U3470 , P3_U4962 );
nand NAND3_1142 ( P3_U2951 , P3_U4958 , P3_U3468 , P3_U4957 );
nand NAND3_1143 ( P3_U2952 , P3_U4953 , P3_U3466 , P3_U4952 );
nand NAND3_1144 ( P3_U2953 , P3_U4948 , P3_U3464 , P3_U4947 );
nand NAND3_1145 ( P3_U2954 , P3_U4943 , P3_U3462 , P3_U4942 );
nand NAND3_1146 ( P3_U2955 , P3_U4938 , P3_U3460 , P3_U4937 );
nand NAND3_1147 ( P3_U2956 , P3_U4921 , P3_U3456 , P3_U4920 );
nand NAND3_1148 ( P3_U2957 , P3_U4916 , P3_U3454 , P3_U4915 );
nand NAND3_1149 ( P3_U2958 , P3_U4911 , P3_U3452 , P3_U4910 );
nand NAND3_1150 ( P3_U2959 , P3_U4906 , P3_U3450 , P3_U4905 );
nand NAND3_1151 ( P3_U2960 , P3_U4901 , P3_U3448 , P3_U4900 );
nand NAND3_1152 ( P3_U2961 , P3_U4896 , P3_U3446 , P3_U4895 );
nand NAND3_1153 ( P3_U2962 , P3_U4891 , P3_U3444 , P3_U4890 );
nand NAND3_1154 ( P3_U2963 , P3_U4886 , P3_U3442 , P3_U4885 );
nand NAND3_1155 ( P3_U2964 , P3_U4869 , P3_U3439 , P3_U4868 );
nand NAND3_1156 ( P3_U2965 , P3_U4864 , P3_U3437 , P3_U4863 );
nand NAND3_1157 ( P3_U2966 , P3_U4859 , P3_U3435 , P3_U4858 );
nand NAND3_1158 ( P3_U2967 , P3_U4854 , P3_U3433 , P3_U4853 );
nand NAND3_1159 ( P3_U2968 , P3_U4849 , P3_U3431 , P3_U4848 );
nand NAND3_1160 ( P3_U2969 , P3_U4844 , P3_U3429 , P3_U4843 );
nand NAND3_1161 ( P3_U2970 , P3_U4839 , P3_U3427 , P3_U4838 );
nand NAND3_1162 ( P3_U2971 , P3_U4834 , P3_U3425 , P3_U4833 );
nand NAND3_1163 ( P3_U2972 , P3_U4818 , P3_U3421 , P3_U4817 );
nand NAND3_1164 ( P3_U2973 , P3_U4813 , P3_U3419 , P3_U4812 );
nand NAND3_1165 ( P3_U2974 , P3_U4808 , P3_U3417 , P3_U4807 );
nand NAND3_1166 ( P3_U2975 , P3_U4803 , P3_U3415 , P3_U4802 );
nand NAND3_1167 ( P3_U2976 , P3_U4798 , P3_U3413 , P3_U4797 );
nand NAND3_1168 ( P3_U2977 , P3_U4793 , P3_U3411 , P3_U4792 );
nand NAND3_1169 ( P3_U2978 , P3_U4788 , P3_U3409 , P3_U4787 );
nand NAND3_1170 ( P3_U2979 , P3_U4783 , P3_U3407 , P3_U4782 );
nand NAND3_1171 ( P3_U2980 , P3_U4766 , P3_U3403 , P3_U4765 );
nand NAND3_1172 ( P3_U2981 , P3_U4761 , P3_U3401 , P3_U4760 );
nand NAND3_1173 ( P3_U2982 , P3_U4756 , P3_U3399 , P3_U4755 );
nand NAND3_1174 ( P3_U2983 , P3_U4751 , P3_U3397 , P3_U4750 );
nand NAND3_1175 ( P3_U2984 , P3_U4746 , P3_U3395 , P3_U4745 );
nand NAND3_1176 ( P3_U2985 , P3_U4741 , P3_U3393 , P3_U4740 );
nand NAND3_1177 ( P3_U2986 , P3_U4736 , P3_U3391 , P3_U4735 );
nand NAND3_1178 ( P3_U2987 , P3_U4731 , P3_U3389 , P3_U4730 );
nand NAND3_1179 ( P3_U2988 , P3_U4714 , P3_U3385 , P3_U4713 );
nand NAND3_1180 ( P3_U2989 , P3_U4709 , P3_U3383 , P3_U4708 );
nand NAND3_1181 ( P3_U2990 , P3_U4704 , P3_U3381 , P3_U4703 );
nand NAND3_1182 ( P3_U2991 , P3_U4699 , P3_U3379 , P3_U4698 );
nand NAND3_1183 ( P3_U2992 , P3_U4694 , P3_U3377 , P3_U4693 );
nand NAND3_1184 ( P3_U2993 , P3_U4689 , P3_U3375 , P3_U4688 );
nand NAND3_1185 ( P3_U2994 , P3_U4684 , P3_U3373 , P3_U4683 );
nand NAND3_1186 ( P3_U2995 , P3_U4679 , P3_U3371 , P3_U4678 );
nand NAND3_1187 ( P3_U2996 , P3_U7959 , P3_U7958 , P3_U3367 );
nand NAND4_1188 ( P3_U2997 , P3_U4636 , P3_U4635 , P3_U4634 , P3_U4329 );
nand NAND2_1189 ( P3_U2998 , P3_U3363 , P3_U4632 );
and AND2_1190 ( P3_U2999 , P3_DATAWIDTH_REG_31_ , P3_U7937 );
and AND2_1191 ( P3_U3000 , P3_DATAWIDTH_REG_30_ , P3_U7937 );
and AND2_1192 ( P3_U3001 , P3_DATAWIDTH_REG_29_ , P3_U7937 );
and AND2_1193 ( P3_U3002 , P3_DATAWIDTH_REG_28_ , P3_U7937 );
and AND2_1194 ( P3_U3003 , P3_DATAWIDTH_REG_27_ , P3_U7937 );
and AND2_1195 ( P3_U3004 , P3_DATAWIDTH_REG_26_ , P3_U7937 );
and AND2_1196 ( P3_U3005 , P3_DATAWIDTH_REG_25_ , P3_U7937 );
and AND2_1197 ( P3_U3006 , P3_DATAWIDTH_REG_24_ , P3_U7937 );
and AND2_1198 ( P3_U3007 , P3_DATAWIDTH_REG_23_ , P3_U7937 );
and AND2_1199 ( P3_U3008 , P3_DATAWIDTH_REG_22_ , P3_U7937 );
and AND2_1200 ( P3_U3009 , P3_DATAWIDTH_REG_21_ , P3_U7937 );
and AND2_1201 ( P3_U3010 , P3_DATAWIDTH_REG_20_ , P3_U7937 );
and AND2_1202 ( P3_U3011 , P3_DATAWIDTH_REG_19_ , P3_U7937 );
and AND2_1203 ( P3_U3012 , P3_DATAWIDTH_REG_18_ , P3_U7937 );
and AND2_1204 ( P3_U3013 , P3_DATAWIDTH_REG_17_ , P3_U7937 );
and AND2_1205 ( P3_U3014 , P3_DATAWIDTH_REG_16_ , P3_U7937 );
and AND2_1206 ( P3_U3015 , P3_DATAWIDTH_REG_15_ , P3_U7937 );
and AND2_1207 ( P3_U3016 , P3_DATAWIDTH_REG_14_ , P3_U7937 );
and AND2_1208 ( P3_U3017 , P3_DATAWIDTH_REG_13_ , P3_U7937 );
and AND2_1209 ( P3_U3018 , P3_DATAWIDTH_REG_12_ , P3_U7937 );
and AND2_1210 ( P3_U3019 , P3_DATAWIDTH_REG_11_ , P3_U7937 );
and AND2_1211 ( P3_U3020 , P3_DATAWIDTH_REG_10_ , P3_U7937 );
and AND2_1212 ( P3_U3021 , P3_DATAWIDTH_REG_9_ , P3_U7937 );
and AND2_1213 ( P3_U3022 , P3_DATAWIDTH_REG_8_ , P3_U7937 );
and AND2_1214 ( P3_U3023 , P3_DATAWIDTH_REG_7_ , P3_U7937 );
and AND2_1215 ( P3_U3024 , P3_DATAWIDTH_REG_6_ , P3_U7937 );
and AND2_1216 ( P3_U3025 , P3_DATAWIDTH_REG_5_ , P3_U7937 );
and AND2_1217 ( P3_U3026 , P3_DATAWIDTH_REG_4_ , P3_U7937 );
and AND2_1218 ( P3_U3027 , P3_DATAWIDTH_REG_3_ , P3_U7937 );
and AND2_1219 ( P3_U3028 , P3_DATAWIDTH_REG_2_ , P3_U7937 );
nand NAND3_1220 ( P3_U3029 , P3_U7934 , P3_U7933 , P3_U4463 );
nand NAND3_1221 ( P3_U3030 , P3_U7932 , P3_U7931 , P3_U3311 );
nand NAND2_1222 ( P3_U3031 , P3_U3310 , P3_U4457 );
nand NAND3_1223 ( P3_U3032 , P3_U4443 , P3_U4442 , P3_U4444 );
nand NAND3_1224 ( P3_U3033 , P3_U4440 , P3_U4439 , P3_U4441 );
nand NAND3_1225 ( P3_U3034 , P3_U4437 , P3_U4436 , P3_U4438 );
nand NAND3_1226 ( P3_U3035 , P3_U4434 , P3_U4433 , P3_U4435 );
nand NAND3_1227 ( P3_U3036 , P3_U4431 , P3_U4430 , P3_U4432 );
nand NAND3_1228 ( P3_U3037 , P3_U4428 , P3_U4427 , P3_U4429 );
nand NAND3_1229 ( P3_U3038 , P3_U4425 , P3_U4424 , P3_U4426 );
nand NAND3_1230 ( P3_U3039 , P3_U4422 , P3_U4421 , P3_U4423 );
nand NAND3_1231 ( P3_U3040 , P3_U4419 , P3_U4418 , P3_U4420 );
nand NAND3_1232 ( P3_U3041 , P3_U4416 , P3_U4415 , P3_U4417 );
nand NAND3_1233 ( P3_U3042 , P3_U4413 , P3_U4412 , P3_U4414 );
nand NAND3_1234 ( P3_U3043 , P3_U4410 , P3_U4409 , P3_U4411 );
nand NAND3_1235 ( P3_U3044 , P3_U4407 , P3_U4406 , P3_U4408 );
nand NAND3_1236 ( P3_U3045 , P3_U4404 , P3_U4403 , P3_U4405 );
nand NAND3_1237 ( P3_U3046 , P3_U4401 , P3_U4400 , P3_U4402 );
nand NAND3_1238 ( P3_U3047 , P3_U4398 , P3_U4397 , P3_U4399 );
nand NAND3_1239 ( P3_U3048 , P3_U4395 , P3_U4394 , P3_U4396 );
nand NAND3_1240 ( P3_U3049 , P3_U4392 , P3_U4391 , P3_U4393 );
nand NAND3_1241 ( P3_U3050 , P3_U4389 , P3_U4388 , P3_U4390 );
nand NAND3_1242 ( P3_U3051 , P3_U4386 , P3_U4385 , P3_U4387 );
nand NAND3_1243 ( P3_U3052 , P3_U4383 , P3_U4382 , P3_U4384 );
nand NAND3_1244 ( P3_U3053 , P3_U4380 , P3_U4379 , P3_U4381 );
nand NAND3_1245 ( P3_U3054 , P3_U4377 , P3_U4376 , P3_U4378 );
nand NAND3_1246 ( P3_U3055 , P3_U4374 , P3_U4373 , P3_U4375 );
nand NAND3_1247 ( P3_U3056 , P3_U4371 , P3_U4370 , P3_U4372 );
nand NAND3_1248 ( P3_U3057 , P3_U4368 , P3_U4367 , P3_U4369 );
nand NAND3_1249 ( P3_U3058 , P3_U4365 , P3_U4364 , P3_U4366 );
nand NAND3_1250 ( P3_U3059 , P3_U4362 , P3_U4361 , P3_U4363 );
nand NAND3_1251 ( P3_U3060 , P3_U4359 , P3_U4358 , P3_U4360 );
nand NAND3_1252 ( P3_U3061 , P3_U4356 , P3_U4355 , P3_U4357 );
nand NAND4_1253 ( P3_U3062 , P3_U4247 , P3_U4246 , P3_U4245 , P3_U4244 );
nand NAND4_1254 ( P3_U3063 , P3_U4243 , P3_U4242 , P3_U4241 , P3_U4240 );
nand NAND4_1255 ( P3_U3064 , P3_U4239 , P3_U4238 , P3_U4237 , P3_U4236 );
nand NAND4_1256 ( P3_U3065 , P3_U4235 , P3_U4234 , P3_U4233 , P3_U4232 );
nand NAND4_1257 ( P3_U3066 , P3_U4231 , P3_U4230 , P3_U4229 , P3_U4228 );
nand NAND4_1258 ( P3_U3067 , P3_U4227 , P3_U4226 , P3_U4225 , P3_U4224 );
nand NAND4_1259 ( P3_U3068 , P3_U4223 , P3_U4222 , P3_U4221 , P3_U4220 );
nand NAND4_1260 ( P3_U3069 , P3_U4219 , P3_U4218 , P3_U4217 , P3_U4216 );
nand NAND2_1261 ( P3_U3070 , P3_U2457 , P3_U4642 );
nand NAND2_1262 ( P3_U3071 , P3_U2459 , P3_U4642 );
nand NAND2_1263 ( P3_U3072 , P3_U2458 , P3_U4642 );
nand NAND2_1264 ( P3_U3073 , P3_U2460 , P3_U4642 );
nand NAND5_1265 ( P3_U3074 , P3_U3346 , P3_U3345 , P3_U3347 , P3_U3344 , P3_U3343 );
not NOT1_1266 ( P3_U3075 , P3_REQUESTPENDING_REG );
not NOT1_1267 ( P3_U3076 , P3_STATE_REG_1_ );
nand NAND2_1268 ( P3_U3077 , P3_STATE_REG_1_ , P3_U3085 );
nand NAND2_1269 ( P3_U3078 , P3_U4308 , P3_U3079 );
not NOT1_1270 ( P3_U3079 , P3_STATE_REG_2_ );
nand NAND2_1271 ( P3_U3080 , P3_STATE_REG_2_ , P3_U4308 );
not NOT1_1272 ( P3_U3081 , P3_REIP_REG_1_ );
nand NAND2_1273 ( P3_U3082 , P3_STATE_REG_1_ , P3_U3079 );
or OR2_1274 ( P3_U3083 , P3_STATE_REG_1_ , P3_STATE_REG_2_ );
not NOT1_1275 ( P3_U3084 , HOLD );
not NOT1_1276 ( P3_U3085 , P3_STATE_REG_0_ );
nand NAND2_1277 ( P3_U3086 , P3_STATE_REG_0_ , P3_U3087 );
nand NAND2_1278 ( P3_U3087 , P3_REQUESTPENDING_REG , P3_U3084 );
or OR2_1279 ( P3_U3088 , HOLD , P3_REQUESTPENDING_REG );
not NOT1_1280 ( P3_U3089 , P3_STATE2_REG_1_ );
not NOT1_1281 ( P3_U3090 , P3_STATE2_REG_2_ );
or OR2_1282 ( P3_U3091 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_1283 ( P3_U3092 , P3_U4467 , P3_U3097 );
not NOT1_1284 ( P3_U3093 , P3_INSTQUEUERD_ADDR_REG_0_ );
not NOT1_1285 ( P3_U3094 , P3_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_1286 ( P3_U3095 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_1287 ( P3_U3096 , P3_U4332 , P3_U3097 );
not NOT1_1288 ( P3_U3097 , P3_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_1289 ( P3_U3098 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_U3100 );
nand NAND2_1290 ( P3_U3099 , P3_U4470 , P3_U4332 );
not NOT1_1291 ( P3_U3100 , P3_INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_1292 ( P3_U3101 , P3_U3341 , P3_U3340 , P3_U3342 , P3_U3339 , P3_U3338 );
nand NAND5_1293 ( P3_U3102 , P3_U3326 , P3_U3325 , P3_U3327 , P3_U3324 , P3_U3323 );
nand NAND2_1294 ( P3_U3103 , P3_U3074 , P3_U3110 );
nand NAND5_1295 ( P3_U3104 , P3_U3321 , P3_U3320 , P3_U3322 , P3_U3319 , P3_U3318 );
nand NAND2_1296 ( P3_U3105 , P3_U4466 , P3_U3085 );
nand NAND2_1297 ( P3_U3106 , P3_U4293 , P3_U2630 );
nand NAND5_1298 ( P3_U3107 , P3_U3331 , P3_U3330 , P3_U3332 , P3_U3329 , P3_U3328 );
nand NAND5_1299 ( P3_U3108 , P3_U3316 , P3_U3315 , P3_U3317 , P3_U3314 , P3_U3313 );
nand NAND2_1300 ( P3_U3109 , P3_U2353 , P3_U4488 );
nand NAND5_1301 ( P3_U3110 , P3_U3351 , P3_U3350 , P3_U3352 , P3_U3349 , P3_U3348 );
nand NAND2_1302 ( P3_U3111 , P3_U3104 , P3_U3108 );
nand NAND2_1303 ( P3_U3112 , P3_U4505 , P3_U3108 );
nand NAND2_1304 ( P3_U3113 , P3_U4607 , P3_U3110 );
nand NAND2_1305 ( P3_U3114 , P3_U4488 , P3_U4505 );
nand NAND2_1306 ( P3_U3115 , P3_U2451 , P3_U4297 );
nand NAND2_1307 ( P3_U3116 , P3_U2452 , P3_U4297 );
nand NAND2_1308 ( P3_U3117 , P3_U2452 , P3_U4296 );
nand NAND2_1309 ( P3_U3118 , P3_U4488 , P3_U3104 );
nand NAND2_1310 ( P3_U3119 , P3_U3356 , P3_U2353 );
nand NAND5_1311 ( P3_U3120 , P3_U7949 , P3_U7948 , P3_U3262 , P3_U4313 , P3_LT_563_U6 );
not NOT1_1312 ( P3_U3121 , P3_STATE2_REG_0_ );
nand NAND2_1313 ( P3_U3122 , P3_STATE2_REG_0_ , P3_U4629 );
or OR2_1314 ( P3_U3123 , P3_STATE2_REG_3_ , P3_STATE2_REG_1_ );
nand NAND2_1315 ( P3_U3124 , P3_STATE2_REG_2_ , P3_U3089 );
or OR2_1316 ( P3_U3125 , P3_STATE2_REG_2_ , P3_STATE2_REG_1_ );
nand NAND2_1317 ( P3_U3126 , P3_LTE_597_U6 , P3_STATE2_REG_3_ );
nand NAND2_1318 ( P3_U3127 , P3_U4666 , P3_U3121 );
not NOT1_1319 ( P3_U3128 , P3_INSTQUEUEWR_ADDR_REG_0_ );
not NOT1_1320 ( P3_U3129 , P3_INSTQUEUEWR_ADDR_REG_1_ );
nand NAND2_1321 ( P3_U3130 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_INSTQUEUEWR_ADDR_REG_0_ );
not NOT1_1322 ( P3_U3131 , P3_INSTQUEUEWR_ADDR_REG_2_ );
nand NAND2_1323 ( P3_U3132 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_U4648 );
not NOT1_1324 ( P3_U3133 , P3_INSTQUEUEWR_ADDR_REG_3_ );
nand NAND2_1325 ( P3_U3134 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_U4649 );
or OR2_1326 ( P3_U3135 , P3_STATE2_REG_3_ , P3_STATE2_REG_2_ );
nand NAND2_1327 ( P3_U3136 , P3_U4295 , P3_STATEBS16_REG );
nand NAND2_1328 ( P3_U3137 , P3_U3153 , P3_U4641 );
nand NAND2_1329 ( P3_U3138 , P3_U3137 , P3_U3128 );
nand NAND2_1330 ( P3_U3139 , P3_U3180 , P3_U4651 );
nand NAND2_1331 ( P3_U3140 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_U3141 );
nand NAND2_1332 ( P3_U3141 , P3_U3150 , P3_U3158 );
nand NAND2_1333 ( P3_U3142 , P3_U4331 , P3_U4655 );
nand NAND2_1334 ( P3_U3143 , P3_U3156 , P3_U3128 );
nand NAND2_1335 ( P3_U3144 , P3_U4647 , P3_U2486 );
nand NAND2_1336 ( P3_U3145 , P3_U3144 , P3_U4667 );
nand NAND2_1337 ( P3_U3146 , P3_U3134 , P3_U4663 );
nand NAND2_1338 ( P3_U3147 , P3_U3386 , P3_U2492 );
nand NAND2_1339 ( P3_U3148 , P3_U3141 , P3_U3128 );
nand NAND2_1340 ( P3_U3149 , P3_U2490 , P3_U2486 );
nand NAND2_1341 ( P3_U3150 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_U3137 );
nand NAND2_1342 ( P3_U3151 , P3_U3149 , P3_U4719 );
nand NAND2_1343 ( P3_U3152 , P3_U3147 , P3_U4717 );
nand NAND2_1344 ( P3_U3153 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_U3129 );
nand NAND2_1345 ( P3_U3154 , P3_U3404 , P3_U4640 );
nand NAND2_1346 ( P3_U3155 , P3_U4643 , P3_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_1347 ( P3_U3156 , P3_U3148 , P3_U3155 );
nand NAND2_1348 ( P3_U3157 , P3_U2493 , P3_U2486 );
nand NAND2_1349 ( P3_U3158 , P3_U4642 , P3_U3128 );
nand NAND2_1350 ( P3_U3159 , P3_U3157 , P3_U4771 );
nand NAND2_1351 ( P3_U3160 , P3_U3154 , P3_U4769 );
nand NAND2_1352 ( P3_U3161 , P3_U3422 , P3_U2492 );
nand NAND2_1353 ( P3_U3162 , P3_U2495 , P3_U2486 );
nand NAND2_1354 ( P3_U3163 , P3_U3162 , P3_U4822 );
nand NAND3_1355 ( P3_U3164 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_U3131 , P3_U4648 );
nand NAND2_1356 ( P3_U3165 , P3_U7965 , P3_U3142 );
nand NAND2_1357 ( P3_U3166 , P3_U2498 , P3_U4647 );
nand NAND2_1358 ( P3_U3167 , P3_U3166 , P3_U4874 );
nand NAND2_1359 ( P3_U3168 , P3_U3164 , P3_U4872 );
nand NAND2_1360 ( P3_U3169 , P3_U3457 , P3_U2501 );
nand NAND2_1361 ( P3_U3170 , P3_U2498 , P3_U2490 );
nand NAND2_1362 ( P3_U3171 , P3_U3170 , P3_U4926 );
nand NAND2_1363 ( P3_U3172 , P3_U3169 , P3_U4924 );
nand NAND2_1364 ( P3_U3173 , P3_U3475 , P3_U4640 );
nand NAND2_1365 ( P3_U3174 , P3_U2498 , P3_U2493 );
nand NAND2_1366 ( P3_U3175 , P3_U3174 , P3_U4978 );
nand NAND2_1367 ( P3_U3176 , P3_U3173 , P3_U4976 );
nand NAND3_1368 ( P3_U3177 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_U3129 , P3_U2501 );
nand NAND2_1369 ( P3_U3178 , P3_U2498 , P3_U2495 );
nand NAND2_1370 ( P3_U3179 , P3_U3178 , P3_U5029 );
nand NAND2_1371 ( P3_U3180 , P3_U4649 , P3_U3133 );
nand NAND2_1372 ( P3_U3181 , P3_U2485 , P3_U4657 );
nand NAND2_1373 ( P3_U3182 , P3_U3368 , P3_U3181 );
nand NAND2_1374 ( P3_U3183 , P3_U2504 , P3_U4647 );
nand NAND2_1375 ( P3_U3184 , P3_U3183 , P3_U3181 );
nand NAND2_1376 ( P3_U3185 , P3_U3180 , P3_U4331 );
nand NAND2_1377 ( P3_U3186 , P3_U3527 , P3_U2492 );
nand NAND2_1378 ( P3_U3187 , P3_U2504 , P3_U2490 );
nand NAND2_1379 ( P3_U3188 , P3_U3187 , P3_U5130 );
nand NAND2_1380 ( P3_U3189 , P3_U3186 , P3_U5128 );
nand NAND2_1381 ( P3_U3190 , P3_U3545 , P3_U4640 );
nand NAND2_1382 ( P3_U3191 , P3_U2504 , P3_U2493 );
nand NAND2_1383 ( P3_U3192 , P3_U3191 , P3_U5182 );
nand NAND2_1384 ( P3_U3193 , P3_U3190 , P3_U5180 );
nand NAND2_1385 ( P3_U3194 , P3_U3563 , P3_U2492 );
nand NAND2_1386 ( P3_U3195 , P3_U2504 , P3_U2495 );
nand NAND2_1387 ( P3_U3196 , P3_U3581 , P3_U4648 );
nand NAND2_1388 ( P3_U3197 , P3_U2508 , P3_U4647 );
nand NAND2_1389 ( P3_U3198 , P3_U3196 , P3_U5282 );
nand NAND3_1390 ( P3_U3199 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_U3133 , P3_U2501 );
nand NAND2_1391 ( P3_U3200 , P3_U2508 , P3_U2490 );
nand NAND2_1392 ( P3_U3201 , P3_U3199 , P3_U5333 );
nand NAND2_1393 ( P3_U3202 , P3_U3616 , P3_U4640 );
nand NAND2_1394 ( P3_U3203 , P3_U2508 , P3_U2493 );
nand NAND2_1395 ( P3_U3204 , P3_U3202 , P3_U5384 );
nand NAND2_1396 ( P3_U3205 , P3_U3634 , P3_U2501 );
nand NAND2_1397 ( P3_U3206 , P3_U2508 , P3_U2495 );
not NOT1_1398 ( P3_U3207 , P3_FLUSH_REG );
nand NAND2_1399 ( P3_U3208 , P3_U4539 , P3_U3102 );
nand NAND2_1400 ( P3_U3209 , P3_U2514 , P3_U3113 );
not NOT1_1401 ( P3_U3210 , P3_GTE_412_U6 );
not NOT1_1402 ( P3_U3211 , P3_GTE_485_U6 );
not NOT1_1403 ( P3_U3212 , P3_GTE_390_U6 );
not NOT1_1404 ( P3_U3213 , P3_GTE_450_U6 );
not NOT1_1405 ( P3_U3214 , P3_GTE_504_U6 );
not NOT1_1406 ( P3_U3215 , P3_GTE_401_U6 );
nand NAND2_1407 ( P3_U3216 , P3_U4590 , P3_U3074 );
nand NAND2_1408 ( P3_U3217 , P3_U2450 , P3_U4323 );
nand NAND5_1409 ( P3_U3218 , P3_U3336 , P3_U3335 , P3_U3337 , P3_U3334 , P3_U3333 );
nand NAND2_1410 ( P3_U3219 , P3_U3662 , P3_U2461 );
nand NAND3_1411 ( P3_U3220 , P3_U7976 , P3_U7975 , P3_U3667 );
nand NAND3_1412 ( P3_U3221 , P3_U3222 , P3_U3119 , P3_U5524 );
nand NAND2_1413 ( P3_U3222 , P3_U4314 , P3_U3218 );
nand NAND2_1414 ( P3_U3223 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_U5503 );
nand NAND2_1415 ( P3_U3224 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_U5505 );
nand NAND2_1416 ( P3_U3225 , P3_U3096 , P3_U3227 );
nand NAND2_1417 ( P3_U3226 , P3_U3674 , P3_U2517 );
nand NAND2_1418 ( P3_U3227 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_U3095 );
nand NAND2_1419 ( P3_U3228 , P3_U3091 , P3_U3095 );
nand NAND3_1420 ( P3_U3229 , P3_U4323 , P3_U3218 , P3_U4350 );
nand NAND2_1421 ( P3_U3230 , P3_U2518 , P3_U3243 );
nand NAND2_1422 ( P3_U3231 , P3_U3115 , P3_U5559 );
not NOT1_1423 ( P3_U3232 , P3_LT_589_U6 );
nand NAND3_1424 ( P3_U3233 , P3_U4330 , P3_U3127 , P3_U5578 );
nand NAND2_1425 ( P3_U3234 , P3_U3135 , P3_U3123 );
nand NAND3_1426 ( P3_U3235 , P3_U3101 , P3_U3104 , P3_U4294 );
nand NAND3_1427 ( P3_U3236 , P3_U3101 , P3_U2630 , P3_U4505 );
not NOT1_1428 ( P3_U3237 , P3_GTE_370_U6 );
not NOT1_1429 ( P3_U3238 , P3_GTE_355_U6 );
nand NAND2_1430 ( P3_U3239 , P3_U4295 , P3_U3089 );
not NOT1_1431 ( P3_U3240 , P3_REIP_REG_0_ );
not NOT1_1432 ( P3_U3241 , P3_U2628 );
nand NAND2_1433 ( P3_U3242 , P3_U3661 , P3_U2450 );
nand NAND2_1434 ( P3_U3243 , P3_U2461 , P3_U4314 );
nand NAND2_1435 ( P3_U3244 , P3_U4352 , P3_U4522 );
nand NAND2_1436 ( P3_U3245 , P3_U4352 , P3_U3102 );
nand NAND3_1437 ( P3_U3246 , P3_U3663 , P3_U2449 , P3_U3664 );
nand NAND2_1438 ( P3_U3247 , P3_STATE2_REG_2_ , P3_U3248 );
nand NAND2_1439 ( P3_U3248 , P3_U4336 , P3_U5630 );
nand NAND2_1440 ( P3_U3249 , P3_U6403 , P3_U6402 );
nand NAND2_1441 ( P3_U3250 , P3_U2390 , P3_U6663 );
nand NAND2_1442 ( P3_U3251 , P3_U6758 , P3_U6757 );
nand NAND2_1443 ( P3_U3252 , P3_U2390 , P3_U6853 );
nand NAND2_1444 ( P3_U3253 , P3_U2390 , P3_U6997 );
nand NAND2_1445 ( P3_U3254 , P3_U5490 , P3_U5489 );
nand NAND2_1446 ( P3_U3255 , P3_U5487 , P3_U5486 );
not NOT1_1447 ( P3_U3256 , P3_EBX_REG_31_ );
or OR2_1448 ( P3_U3257 , P3_STATEBS16_REG , U209 );
not NOT1_1449 ( P3_U3258 , P3_ADD_318_U69 );
nand NAND2_1450 ( P3_U3259 , P3_ADD_318_U69 , P3_U2385 );
nand NAND2_1451 ( P3_U3260 , P3_U4030 , P3_U4334 );
nand NAND4_1452 ( P3_U3261 , P3_U4148 , P3_U4144 , P3_U4141 , P3_U4138 );
nand NAND3_1453 ( P3_U3262 , P3_U2462 , P3_U3108 , P3_U4282 );
not NOT1_1454 ( P3_U3263 , P3_CODEFETCH_REG );
not NOT1_1455 ( P3_U3264 , P3_READREQUEST_REG );
nand NAND2_1456 ( P3_U3265 , P3_U3099 , P3_U3224 );
nand NAND2_1457 ( P3_U3266 , P3_U3223 , P3_U7515 );
nand NAND2_1458 ( P3_U3267 , P3_U4289 , P3_U3092 );
nand NAND2_1459 ( P3_U3268 , P3_U3098 , P3_U7774 );
nand NAND2_1460 ( P3_U3269 , P3_U7961 , P3_U7960 );
nand NAND2_1461 ( P3_U3270 , P3_U7964 , P3_U7963 );
nand NAND2_1462 ( P3_U3271 , P3_U7967 , P3_U7966 );
nand NAND2_1463 ( P3_U3272 , P3_U8033 , P3_U8032 );
nand NAND2_1464 ( P3_U3273 , P3_U8036 , P3_U8035 );
nand NAND2_1465 ( P3_U3274 , P3_U7921 , P3_U7920 );
nand NAND2_1466 ( P3_U3275 , P3_U7923 , P3_U7922 );
nand NAND2_1467 ( P3_U3276 , P3_U7925 , P3_U7924 );
nand NAND2_1468 ( P3_U3277 , P3_U7927 , P3_U7926 );
nand NAND2_1469 ( P3_U3278 , P3_U7936 , P3_U7935 );
and AND2_1470 ( P3_U3279 , P3_U3083 , P3_U4286 );
nand NAND2_1471 ( P3_U3280 , P3_U7939 , P3_U7938 );
nand NAND2_1472 ( P3_U3281 , P3_U7941 , P3_U7940 );
nand NAND2_1473 ( P3_U3282 , P3_U7955 , P3_U7954 );
and AND2_1474 ( P3_U3283 , P3_U3652 , P3_U2356 );
nand NAND2_1475 ( P3_U3284 , P3_U7972 , P3_U7971 );
nand NAND2_1476 ( P3_U3285 , P3_U7980 , P3_U7979 );
nand NAND2_1477 ( P3_U3286 , P3_U7987 , P3_U7986 );
nand NAND2_1478 ( P3_U3287 , P3_U7984 , P3_U7983 );
nand NAND2_1479 ( P3_U3288 , P3_U7990 , P3_U7989 );
nand NAND2_1480 ( P3_U3289 , P3_U7992 , P3_U7991 );
nand NAND2_1481 ( P3_U3290 , P3_U7996 , P3_U7995 );
nor nor_1482 ( P3_U3291 , P3_DATAWIDTH_REG_1_ , P3_REIP_REG_1_ );
nand NAND2_1483 ( P3_U3292 , P3_U8011 , P3_U8010 );
nand NAND2_1484 ( P3_U3293 , P3_U8015 , P3_U8014 );
nand NAND2_1485 ( P3_U3294 , P3_U8017 , P3_U8016 );
nand NAND2_1486 ( P3_U3295 , P3_U8019 , P3_U8018 );
nand NAND2_1487 ( P3_U3296 , P3_U8023 , P3_U8022 );
nand NAND2_1488 ( P3_U3297 , P3_U8027 , P3_U8026 );
nand NAND2_1489 ( P3_U3298 , P3_U8029 , P3_U8028 );
nand NAND2_1490 ( P3_U3299 , P3_U8031 , P3_U8030 );
nand NAND2_1491 ( P3_U3300 , P3_U8039 , P3_U8038 );
nand NAND2_1492 ( P3_U3301 , P3_U8041 , P3_U8040 );
nand NAND2_1493 ( P3_U3302 , P3_U8043 , P3_U8042 );
and AND2_1494 ( P3_U3303 , P3_ADD_495_U8 , P3_U2356 );
nand NAND2_1495 ( P3_U3304 , P3_U8045 , P3_U8044 );
nand NAND2_1496 ( P3_U3305 , P3_U8047 , P3_U8046 );
nand NAND2_1497 ( P3_U3306 , P3_U8049 , P3_U8048 );
nand NAND2_1498 ( P3_U3307 , P3_U8051 , P3_U8050 );
nand NAND2_1499 ( P3_U3308 , P3_U8053 , P3_U8052 );
and AND2_1500 ( P3_U3309 , P3_STATE_REG_0_ , P3_U4447 );
and AND2_1501 ( P3_U3310 , P3_U4456 , P3_U3080 );
and AND2_1502 ( P3_U3311 , P3_U4458 , P3_U3078 );
and AND2_1503 ( P3_U3312 , P3_REQUESTPENDING_REG , P3_STATE_REG_0_ );
and AND4_1504 ( P3_U3313 , P3_U4475 , P3_U4474 , P3_U4473 , P3_U4472 );
and AND4_1505 ( P3_U3314 , P3_U4479 , P3_U4478 , P3_U4477 , P3_U4476 );
and AND2_1506 ( P3_U3315 , P3_U4481 , P3_U4480 );
and AND2_1507 ( P3_U3316 , P3_U4483 , P3_U4482 );
and AND4_1508 ( P3_U3317 , P3_U4487 , P3_U4486 , P3_U4485 , P3_U4484 );
and AND4_1509 ( P3_U3318 , P3_U4492 , P3_U4491 , P3_U4490 , P3_U4489 );
and AND4_1510 ( P3_U3319 , P3_U4496 , P3_U4495 , P3_U4494 , P3_U4493 );
and AND2_1511 ( P3_U3320 , P3_U4498 , P3_U4497 );
and AND2_1512 ( P3_U3321 , P3_U4500 , P3_U4499 );
and AND4_1513 ( P3_U3322 , P3_U4504 , P3_U4503 , P3_U4502 , P3_U4501 );
and AND4_1514 ( P3_U3323 , P3_U4509 , P3_U4508 , P3_U4507 , P3_U4506 );
and AND4_1515 ( P3_U3324 , P3_U4513 , P3_U4512 , P3_U4511 , P3_U4510 );
and AND2_1516 ( P3_U3325 , P3_U4515 , P3_U4514 );
and AND2_1517 ( P3_U3326 , P3_U4517 , P3_U4516 );
and AND4_1518 ( P3_U3327 , P3_U4521 , P3_U4520 , P3_U4519 , P3_U4518 );
and AND4_1519 ( P3_U3328 , P3_U4543 , P3_U4542 , P3_U4541 , P3_U4540 );
and AND4_1520 ( P3_U3329 , P3_U4547 , P3_U4546 , P3_U4545 , P3_U4544 );
and AND2_1521 ( P3_U3330 , P3_U4549 , P3_U4548 );
and AND2_1522 ( P3_U3331 , P3_U4551 , P3_U4550 );
and AND4_1523 ( P3_U3332 , P3_U4555 , P3_U4554 , P3_U4553 , P3_U4552 );
and AND4_1524 ( P3_U3333 , P3_U4560 , P3_U4559 , P3_U4558 , P3_U4557 );
and AND4_1525 ( P3_U3334 , P3_U4564 , P3_U4563 , P3_U4562 , P3_U4561 );
and AND2_1526 ( P3_U3335 , P3_U4566 , P3_U4565 );
and AND2_1527 ( P3_U3336 , P3_U4568 , P3_U4567 );
and AND4_1528 ( P3_U3337 , P3_U4572 , P3_U4571 , P3_U4570 , P3_U4569 );
and AND4_1529 ( P3_U3338 , P3_U4526 , P3_U4525 , P3_U4524 , P3_U4523 );
and AND4_1530 ( P3_U3339 , P3_U4530 , P3_U4529 , P3_U4528 , P3_U4527 );
and AND2_1531 ( P3_U3340 , P3_U4532 , P3_U4531 );
and AND2_1532 ( P3_U3341 , P3_U4534 , P3_U4533 );
and AND4_1533 ( P3_U3342 , P3_U4538 , P3_U4537 , P3_U4536 , P3_U4535 );
and AND4_1534 ( P3_U3343 , P3_U4594 , P3_U4593 , P3_U4592 , P3_U4591 );
and AND4_1535 ( P3_U3344 , P3_U4598 , P3_U4597 , P3_U4596 , P3_U4595 );
and AND2_1536 ( P3_U3345 , P3_U4600 , P3_U4599 );
and AND2_1537 ( P3_U3346 , P3_U4602 , P3_U4601 );
and AND4_1538 ( P3_U3347 , P3_U4606 , P3_U4605 , P3_U4604 , P3_U4603 );
and AND4_1539 ( P3_U3348 , P3_U4577 , P3_U4576 , P3_U4575 , P3_U4574 );
and AND4_1540 ( P3_U3349 , P3_U4581 , P3_U4580 , P3_U4579 , P3_U4578 );
and AND2_1541 ( P3_U3350 , P3_U4583 , P3_U4582 );
and AND2_1542 ( P3_U3351 , P3_U4585 , P3_U4584 );
and AND4_1543 ( P3_U3352 , P3_U4589 , P3_U4588 , P3_U4587 , P3_U4586 );
and AND2_1544 ( P3_U3353 , P3_U2352 , P3_U4293 );
and AND2_1545 ( P3_U3354 , P3_U4556 , P3_U3218 );
and AND2_1546 ( P3_U3355 , P3_U4323 , P3_U3101 );
and AND2_1547 ( P3_U3356 , P3_U4324 , P3_U3101 );
and AND4_1548 ( P3_U3357 , P3_U4612 , P3_U4611 , P3_U4610 , P3_U4609 );
and AND4_1549 ( P3_U3358 , P3_U4616 , P3_U4615 , P3_U4614 , P3_U4613 );
and AND2_1550 ( P3_U3359 , P3_U4539 , P3_U2630 );
and AND3_1551 ( P3_U3360 , P3_U3107 , P3_U3108 , P3_U3218 );
and AND3_1552 ( P3_U3361 , P3_U3235 , P3_U3236 , P3_U4621 );
and AND2_1553 ( P3_U3362 , P3_U4626 , P3_U3089 );
and AND2_1554 ( P3_U3363 , P3_U4631 , P3_U3124 );
and AND2_1555 ( P3_U3364 , P3_U4340 , P3_U2630 );
and AND2_1556 ( P3_U3365 , P3_STATE2_REG_3_ , P3_STATE2_REG_0_ );
and AND2_1557 ( P3_U3366 , P3_U4338 , P3_U4328 );
and AND2_1558 ( P3_U3367 , P3_U3366 , P3_U4639 );
and AND2_1559 ( P3_U3368 , P3_U3165 , P3_U4659 );
and AND2_1560 ( P3_U3369 , P3_U4671 , P3_U4312 );
and AND2_1561 ( P3_U3370 , P3_U4676 , P3_U4675 );
and AND2_1562 ( P3_U3371 , P3_U3370 , P3_U4677 );
and AND2_1563 ( P3_U3372 , P3_U4681 , P3_U4680 );
and AND2_1564 ( P3_U3373 , P3_U3372 , P3_U4682 );
and AND2_1565 ( P3_U3374 , P3_U4686 , P3_U4685 );
and AND2_1566 ( P3_U3375 , P3_U3374 , P3_U4687 );
and AND2_1567 ( P3_U3376 , P3_U4691 , P3_U4690 );
and AND2_1568 ( P3_U3377 , P3_U3376 , P3_U4692 );
and AND2_1569 ( P3_U3378 , P3_U4696 , P3_U4695 );
and AND2_1570 ( P3_U3379 , P3_U3378 , P3_U4697 );
and AND2_1571 ( P3_U3380 , P3_U4701 , P3_U4700 );
and AND2_1572 ( P3_U3381 , P3_U3380 , P3_U4702 );
and AND2_1573 ( P3_U3382 , P3_U4706 , P3_U4705 );
and AND2_1574 ( P3_U3383 , P3_U3382 , P3_U4707 );
and AND2_1575 ( P3_U3384 , P3_U4711 , P3_U4710 );
and AND2_1576 ( P3_U3385 , P3_U3384 , P3_U4712 );
and AND2_1577 ( P3_U3386 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_INSTQUEUEWR_ADDR_REG_1_ );
and AND2_1578 ( P3_U3387 , P3_U4723 , P3_U4312 );
and AND2_1579 ( P3_U3388 , P3_U4728 , P3_U4727 );
and AND2_1580 ( P3_U3389 , P3_U3388 , P3_U4729 );
and AND2_1581 ( P3_U3390 , P3_U4733 , P3_U4732 );
and AND2_1582 ( P3_U3391 , P3_U3390 , P3_U4734 );
and AND2_1583 ( P3_U3392 , P3_U4738 , P3_U4737 );
and AND2_1584 ( P3_U3393 , P3_U3392 , P3_U4739 );
and AND2_1585 ( P3_U3394 , P3_U4743 , P3_U4742 );
and AND2_1586 ( P3_U3395 , P3_U3394 , P3_U4744 );
and AND2_1587 ( P3_U3396 , P3_U4748 , P3_U4747 );
and AND2_1588 ( P3_U3397 , P3_U3396 , P3_U4749 );
and AND2_1589 ( P3_U3398 , P3_U4753 , P3_U4752 );
and AND2_1590 ( P3_U3399 , P3_U3398 , P3_U4754 );
and AND2_1591 ( P3_U3400 , P3_U4758 , P3_U4757 );
and AND2_1592 ( P3_U3401 , P3_U3400 , P3_U4759 );
and AND2_1593 ( P3_U3402 , P3_U4763 , P3_U4762 );
and AND2_1594 ( P3_U3403 , P3_U3402 , P3_U4764 );
and AND2_1595 ( P3_U3404 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_INSTQUEUEWR_ADDR_REG_2_ );
and AND2_1596 ( P3_U3405 , P3_U4775 , P3_U4312 );
and AND2_1597 ( P3_U3406 , P3_U4780 , P3_U4779 );
and AND2_1598 ( P3_U3407 , P3_U3406 , P3_U4781 );
and AND2_1599 ( P3_U3408 , P3_U4785 , P3_U4784 );
and AND2_1600 ( P3_U3409 , P3_U3408 , P3_U4786 );
and AND2_1601 ( P3_U3410 , P3_U4790 , P3_U4789 );
and AND2_1602 ( P3_U3411 , P3_U3410 , P3_U4791 );
and AND2_1603 ( P3_U3412 , P3_U4795 , P3_U4794 );
and AND2_1604 ( P3_U3413 , P3_U3412 , P3_U4796 );
and AND2_1605 ( P3_U3414 , P3_U4800 , P3_U4799 );
and AND2_1606 ( P3_U3415 , P3_U3414 , P3_U4801 );
and AND2_1607 ( P3_U3416 , P3_U4805 , P3_U4804 );
and AND2_1608 ( P3_U3417 , P3_U3416 , P3_U4806 );
and AND2_1609 ( P3_U3418 , P3_U4810 , P3_U4809 );
and AND2_1610 ( P3_U3419 , P3_U3418 , P3_U4811 );
and AND2_1611 ( P3_U3420 , P3_U4815 , P3_U4814 );
and AND2_1612 ( P3_U3421 , P3_U3420 , P3_U4816 );
and AND2_1613 ( P3_U3422 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_U3129 );
and AND2_1614 ( P3_U3423 , P3_U4826 , P3_U4312 );
and AND2_1615 ( P3_U3424 , P3_U4831 , P3_U4830 );
and AND2_1616 ( P3_U3425 , P3_U3424 , P3_U4832 );
and AND2_1617 ( P3_U3426 , P3_U4836 , P3_U4835 );
and AND2_1618 ( P3_U3427 , P3_U3426 , P3_U4837 );
and AND2_1619 ( P3_U3428 , P3_U4841 , P3_U4840 );
and AND2_1620 ( P3_U3429 , P3_U3428 , P3_U4842 );
and AND2_1621 ( P3_U3430 , P3_U4846 , P3_U4845 );
and AND2_1622 ( P3_U3431 , P3_U3430 , P3_U4847 );
and AND2_1623 ( P3_U3432 , P3_U4851 , P3_U4850 );
and AND2_1624 ( P3_U3433 , P3_U3432 , P3_U4852 );
and AND2_1625 ( P3_U3434 , P3_U4856 , P3_U4855 );
and AND2_1626 ( P3_U3435 , P3_U3434 , P3_U4857 );
and AND2_1627 ( P3_U3436 , P3_U4861 , P3_U4860 );
and AND2_1628 ( P3_U3437 , P3_U3436 , P3_U4862 );
and AND2_1629 ( P3_U3438 , P3_U4866 , P3_U4865 );
and AND2_1630 ( P3_U3439 , P3_U3438 , P3_U4867 );
and AND2_1631 ( P3_U3440 , P3_U4878 , P3_U4312 );
and AND2_1632 ( P3_U3441 , P3_U4883 , P3_U4882 );
and AND2_1633 ( P3_U3442 , P3_U3441 , P3_U4884 );
and AND2_1634 ( P3_U3443 , P3_U4888 , P3_U4887 );
and AND2_1635 ( P3_U3444 , P3_U3443 , P3_U4889 );
and AND2_1636 ( P3_U3445 , P3_U4893 , P3_U4892 );
and AND2_1637 ( P3_U3446 , P3_U3445 , P3_U4894 );
and AND2_1638 ( P3_U3447 , P3_U4898 , P3_U4897 );
and AND2_1639 ( P3_U3448 , P3_U3447 , P3_U4899 );
and AND2_1640 ( P3_U3449 , P3_U4903 , P3_U4902 );
and AND2_1641 ( P3_U3450 , P3_U3449 , P3_U4904 );
and AND2_1642 ( P3_U3451 , P3_U4908 , P3_U4907 );
and AND2_1643 ( P3_U3452 , P3_U3451 , P3_U4909 );
and AND2_1644 ( P3_U3453 , P3_U4913 , P3_U4912 );
and AND2_1645 ( P3_U3454 , P3_U3453 , P3_U4914 );
and AND2_1646 ( P3_U3455 , P3_U4918 , P3_U4917 );
and AND2_1647 ( P3_U3456 , P3_U3455 , P3_U4919 );
and AND2_1648 ( P3_U3457 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_INSTQUEUEWR_ADDR_REG_1_ );
and AND2_1649 ( P3_U3458 , P3_U4930 , P3_U4312 );
and AND2_1650 ( P3_U3459 , P3_U4935 , P3_U4934 );
and AND2_1651 ( P3_U3460 , P3_U3459 , P3_U4936 );
and AND2_1652 ( P3_U3461 , P3_U4940 , P3_U4939 );
and AND2_1653 ( P3_U3462 , P3_U3461 , P3_U4941 );
and AND2_1654 ( P3_U3463 , P3_U4945 , P3_U4944 );
and AND2_1655 ( P3_U3464 , P3_U3463 , P3_U4946 );
and AND2_1656 ( P3_U3465 , P3_U4950 , P3_U4949 );
and AND2_1657 ( P3_U3466 , P3_U3465 , P3_U4951 );
and AND2_1658 ( P3_U3467 , P3_U4955 , P3_U4954 );
and AND2_1659 ( P3_U3468 , P3_U3467 , P3_U4956 );
and AND2_1660 ( P3_U3469 , P3_U4960 , P3_U4959 );
and AND2_1661 ( P3_U3470 , P3_U3469 , P3_U4961 );
and AND2_1662 ( P3_U3471 , P3_U4965 , P3_U4964 );
and AND2_1663 ( P3_U3472 , P3_U3471 , P3_U4966 );
and AND2_1664 ( P3_U3473 , P3_U4970 , P3_U4969 );
and AND2_1665 ( P3_U3474 , P3_U3473 , P3_U4971 );
and AND2_1666 ( P3_U3475 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_U3131 );
and AND2_1667 ( P3_U3476 , P3_U4982 , P3_U4312 );
and AND2_1668 ( P3_U3477 , P3_U4987 , P3_U4986 );
and AND2_1669 ( P3_U3478 , P3_U3477 , P3_U4988 );
and AND2_1670 ( P3_U3479 , P3_U4992 , P3_U4991 );
and AND2_1671 ( P3_U3480 , P3_U3479 , P3_U4993 );
and AND2_1672 ( P3_U3481 , P3_U4997 , P3_U4996 );
and AND2_1673 ( P3_U3482 , P3_U3481 , P3_U4998 );
and AND2_1674 ( P3_U3483 , P3_U5002 , P3_U5001 );
and AND2_1675 ( P3_U3484 , P3_U3483 , P3_U5003 );
and AND2_1676 ( P3_U3485 , P3_U5007 , P3_U5006 );
and AND2_1677 ( P3_U3486 , P3_U3485 , P3_U5008 );
and AND2_1678 ( P3_U3487 , P3_U5012 , P3_U5011 );
and AND2_1679 ( P3_U3488 , P3_U3487 , P3_U5013 );
and AND2_1680 ( P3_U3489 , P3_U5017 , P3_U5016 );
and AND2_1681 ( P3_U3490 , P3_U3489 , P3_U5018 );
and AND2_1682 ( P3_U3491 , P3_U5022 , P3_U5021 );
and AND2_1683 ( P3_U3492 , P3_U3491 , P3_U5023 );
and AND2_1684 ( P3_U3493 , P3_U5033 , P3_U4312 );
and AND2_1685 ( P3_U3494 , P3_U5038 , P3_U5037 );
and AND2_1686 ( P3_U3495 , P3_U3494 , P3_U5039 );
and AND2_1687 ( P3_U3496 , P3_U5043 , P3_U5042 );
and AND2_1688 ( P3_U3497 , P3_U3496 , P3_U5044 );
and AND2_1689 ( P3_U3498 , P3_U5048 , P3_U5047 );
and AND2_1690 ( P3_U3499 , P3_U3498 , P3_U5049 );
and AND2_1691 ( P3_U3500 , P3_U5053 , P3_U5052 );
and AND2_1692 ( P3_U3501 , P3_U3500 , P3_U5054 );
and AND2_1693 ( P3_U3502 , P3_U5058 , P3_U5057 );
and AND2_1694 ( P3_U3503 , P3_U3502 , P3_U5059 );
and AND2_1695 ( P3_U3504 , P3_U5063 , P3_U5062 );
and AND2_1696 ( P3_U3505 , P3_U3504 , P3_U5064 );
and AND2_1697 ( P3_U3506 , P3_U5068 , P3_U5067 );
and AND2_1698 ( P3_U3507 , P3_U3506 , P3_U5069 );
and AND2_1699 ( P3_U3508 , P3_U5073 , P3_U5072 );
and AND2_1700 ( P3_U3509 , P3_U3508 , P3_U5074 );
and AND2_1701 ( P3_U3510 , P3_U5082 , P3_U4312 );
and AND2_1702 ( P3_U3511 , P3_U5087 , P3_U5086 );
and AND2_1703 ( P3_U3512 , P3_U3511 , P3_U5088 );
and AND2_1704 ( P3_U3513 , P3_U5092 , P3_U5091 );
and AND2_1705 ( P3_U3514 , P3_U3513 , P3_U5093 );
and AND2_1706 ( P3_U3515 , P3_U5097 , P3_U5096 );
and AND2_1707 ( P3_U3516 , P3_U3515 , P3_U5098 );
and AND2_1708 ( P3_U3517 , P3_U5102 , P3_U5101 );
and AND2_1709 ( P3_U3518 , P3_U3517 , P3_U5103 );
and AND2_1710 ( P3_U3519 , P3_U5107 , P3_U5106 );
and AND2_1711 ( P3_U3520 , P3_U3519 , P3_U5108 );
and AND2_1712 ( P3_U3521 , P3_U5112 , P3_U5111 );
and AND2_1713 ( P3_U3522 , P3_U3521 , P3_U5113 );
and AND2_1714 ( P3_U3523 , P3_U5117 , P3_U5116 );
and AND2_1715 ( P3_U3524 , P3_U3523 , P3_U5118 );
and AND2_1716 ( P3_U3525 , P3_U5122 , P3_U5121 );
and AND2_1717 ( P3_U3526 , P3_U3525 , P3_U5123 );
and AND2_1718 ( P3_U3527 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_U3133 );
and AND2_1719 ( P3_U3528 , P3_U5134 , P3_U4312 );
and AND2_1720 ( P3_U3529 , P3_U5139 , P3_U5138 );
and AND2_1721 ( P3_U3530 , P3_U3529 , P3_U5140 );
and AND2_1722 ( P3_U3531 , P3_U5144 , P3_U5143 );
and AND2_1723 ( P3_U3532 , P3_U3531 , P3_U5145 );
and AND2_1724 ( P3_U3533 , P3_U5149 , P3_U5148 );
and AND2_1725 ( P3_U3534 , P3_U3533 , P3_U5150 );
and AND2_1726 ( P3_U3535 , P3_U5154 , P3_U5153 );
and AND2_1727 ( P3_U3536 , P3_U3535 , P3_U5155 );
and AND2_1728 ( P3_U3537 , P3_U5159 , P3_U5158 );
and AND2_1729 ( P3_U3538 , P3_U3537 , P3_U5160 );
and AND2_1730 ( P3_U3539 , P3_U5164 , P3_U5163 );
and AND2_1731 ( P3_U3540 , P3_U3539 , P3_U5165 );
and AND2_1732 ( P3_U3541 , P3_U5169 , P3_U5168 );
and AND2_1733 ( P3_U3542 , P3_U3541 , P3_U5170 );
and AND2_1734 ( P3_U3543 , P3_U5174 , P3_U5173 );
and AND2_1735 ( P3_U3544 , P3_U3543 , P3_U5175 );
and AND2_1736 ( P3_U3545 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_U3133 );
and AND2_1737 ( P3_U3546 , P3_U5186 , P3_U4312 );
and AND2_1738 ( P3_U3547 , P3_U5191 , P3_U5190 );
and AND2_1739 ( P3_U3548 , P3_U3547 , P3_U5192 );
and AND2_1740 ( P3_U3549 , P3_U5196 , P3_U5195 );
and AND2_1741 ( P3_U3550 , P3_U3549 , P3_U5197 );
and AND2_1742 ( P3_U3551 , P3_U5201 , P3_U5200 );
and AND2_1743 ( P3_U3552 , P3_U3551 , P3_U5202 );
and AND2_1744 ( P3_U3553 , P3_U5206 , P3_U5205 );
and AND2_1745 ( P3_U3554 , P3_U3553 , P3_U5207 );
and AND2_1746 ( P3_U3555 , P3_U5211 , P3_U5210 );
and AND2_1747 ( P3_U3556 , P3_U3555 , P3_U5212 );
and AND2_1748 ( P3_U3557 , P3_U5216 , P3_U5215 );
and AND2_1749 ( P3_U3558 , P3_U3557 , P3_U5217 );
and AND2_1750 ( P3_U3559 , P3_U5221 , P3_U5220 );
and AND2_1751 ( P3_U3560 , P3_U3559 , P3_U5222 );
and AND2_1752 ( P3_U3561 , P3_U5226 , P3_U5225 );
and AND2_1753 ( P3_U3562 , P3_U3561 , P3_U5227 );
nor nor_1754 ( P3_U3563 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_INSTQUEUEWR_ADDR_REG_1_ );
and AND2_1755 ( P3_U3564 , P3_U5237 , P3_U4312 );
and AND3_1756 ( P3_U3565 , P3_U5241 , P3_U5240 , P3_U5243 );
and AND2_1757 ( P3_U3566 , P3_U3565 , P3_U5242 );
and AND3_1758 ( P3_U3567 , P3_U5246 , P3_U5245 , P3_U5248 );
and AND2_1759 ( P3_U3568 , P3_U3567 , P3_U5247 );
and AND3_1760 ( P3_U3569 , P3_U5251 , P3_U5250 , P3_U5253 );
and AND2_1761 ( P3_U3570 , P3_U3569 , P3_U5252 );
and AND3_1762 ( P3_U3571 , P3_U5256 , P3_U5255 , P3_U5258 );
and AND2_1763 ( P3_U3572 , P3_U3571 , P3_U5257 );
and AND3_1764 ( P3_U3573 , P3_U5261 , P3_U5260 , P3_U5263 );
and AND2_1765 ( P3_U3574 , P3_U3573 , P3_U5262 );
and AND3_1766 ( P3_U3575 , P3_U5266 , P3_U5265 , P3_U5268 );
and AND2_1767 ( P3_U3576 , P3_U3575 , P3_U5267 );
and AND3_1768 ( P3_U3577 , P3_U5271 , P3_U5270 , P3_U5273 );
and AND2_1769 ( P3_U3578 , P3_U3577 , P3_U5272 );
and AND3_1770 ( P3_U3579 , P3_U5276 , P3_U5275 , P3_U5278 );
and AND2_1771 ( P3_U3580 , P3_U3579 , P3_U5277 );
nor nor_1772 ( P3_U3581 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_INSTQUEUEWR_ADDR_REG_3_ );
and AND2_1773 ( P3_U3582 , P3_U5288 , P3_U4312 );
and AND3_1774 ( P3_U3583 , P3_U5292 , P3_U5291 , P3_U5294 );
and AND2_1775 ( P3_U3584 , P3_U3583 , P3_U5293 );
and AND3_1776 ( P3_U3585 , P3_U5297 , P3_U5296 , P3_U5299 );
and AND2_1777 ( P3_U3586 , P3_U3585 , P3_U5298 );
and AND3_1778 ( P3_U3587 , P3_U5302 , P3_U5301 , P3_U5304 );
and AND2_1779 ( P3_U3588 , P3_U3587 , P3_U5303 );
and AND3_1780 ( P3_U3589 , P3_U5307 , P3_U5306 , P3_U5309 );
and AND2_1781 ( P3_U3590 , P3_U3589 , P3_U5308 );
and AND3_1782 ( P3_U3591 , P3_U5312 , P3_U5311 , P3_U5314 );
and AND2_1783 ( P3_U3592 , P3_U3591 , P3_U5313 );
and AND3_1784 ( P3_U3593 , P3_U5317 , P3_U5316 , P3_U5319 );
and AND2_1785 ( P3_U3594 , P3_U3593 , P3_U5318 );
and AND3_1786 ( P3_U3595 , P3_U5322 , P3_U5321 , P3_U5324 );
and AND2_1787 ( P3_U3596 , P3_U3595 , P3_U5323 );
and AND3_1788 ( P3_U3597 , P3_U5327 , P3_U5326 , P3_U5329 );
and AND2_1789 ( P3_U3598 , P3_U3597 , P3_U5328 );
and AND2_1790 ( P3_U3599 , P3_U5339 , P3_U4312 );
and AND3_1791 ( P3_U3600 , P3_U5343 , P3_U5342 , P3_U5345 );
and AND2_1792 ( P3_U3601 , P3_U3600 , P3_U5344 );
and AND3_1793 ( P3_U3602 , P3_U5348 , P3_U5347 , P3_U5350 );
and AND2_1794 ( P3_U3603 , P3_U3602 , P3_U5349 );
and AND3_1795 ( P3_U3604 , P3_U5353 , P3_U5352 , P3_U5355 );
and AND2_1796 ( P3_U3605 , P3_U3604 , P3_U5354 );
and AND3_1797 ( P3_U3606 , P3_U5358 , P3_U5357 , P3_U5360 );
and AND2_1798 ( P3_U3607 , P3_U3606 , P3_U5359 );
and AND3_1799 ( P3_U3608 , P3_U5363 , P3_U5362 , P3_U5365 );
and AND2_1800 ( P3_U3609 , P3_U3608 , P3_U5364 );
and AND3_1801 ( P3_U3610 , P3_U5368 , P3_U5367 , P3_U5370 );
and AND2_1802 ( P3_U3611 , P3_U3610 , P3_U5369 );
and AND3_1803 ( P3_U3612 , P3_U5373 , P3_U5372 , P3_U5375 );
and AND2_1804 ( P3_U3613 , P3_U3612 , P3_U5374 );
and AND3_1805 ( P3_U3614 , P3_U5378 , P3_U5377 , P3_U5380 );
and AND2_1806 ( P3_U3615 , P3_U3614 , P3_U5379 );
nor nor_1807 ( P3_U3616 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_INSTQUEUEWR_ADDR_REG_3_ );
and AND2_1808 ( P3_U3617 , P3_U5390 , P3_U4312 );
and AND3_1809 ( P3_U3618 , P3_U5394 , P3_U5393 , P3_U5396 );
and AND2_1810 ( P3_U3619 , P3_U3618 , P3_U5395 );
and AND3_1811 ( P3_U3620 , P3_U5399 , P3_U5398 , P3_U5401 );
and AND2_1812 ( P3_U3621 , P3_U3620 , P3_U5400 );
and AND3_1813 ( P3_U3622 , P3_U5404 , P3_U5403 , P3_U5406 );
and AND2_1814 ( P3_U3623 , P3_U3622 , P3_U5405 );
and AND3_1815 ( P3_U3624 , P3_U5409 , P3_U5408 , P3_U5411 );
and AND2_1816 ( P3_U3625 , P3_U3624 , P3_U5410 );
and AND3_1817 ( P3_U3626 , P3_U5414 , P3_U5413 , P3_U5416 );
and AND2_1818 ( P3_U3627 , P3_U3626 , P3_U5415 );
and AND3_1819 ( P3_U3628 , P3_U5419 , P3_U5418 , P3_U5421 );
and AND2_1820 ( P3_U3629 , P3_U3628 , P3_U5420 );
and AND3_1821 ( P3_U3630 , P3_U5424 , P3_U5423 , P3_U5426 );
and AND2_1822 ( P3_U3631 , P3_U3630 , P3_U5425 );
and AND3_1823 ( P3_U3632 , P3_U5429 , P3_U5428 , P3_U5431 );
and AND2_1824 ( P3_U3633 , P3_U3632 , P3_U5430 );
nor nor_1825 ( P3_U3634 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_INSTQUEUEWR_ADDR_REG_1_ );
and AND2_1826 ( P3_U3635 , P3_U5440 , P3_U4312 );
and AND3_1827 ( P3_U3636 , P3_U5444 , P3_U5443 , P3_U5446 );
and AND2_1828 ( P3_U3637 , P3_U3636 , P3_U5445 );
and AND3_1829 ( P3_U3638 , P3_U5449 , P3_U5448 , P3_U5451 );
and AND2_1830 ( P3_U3639 , P3_U3638 , P3_U5450 );
and AND3_1831 ( P3_U3640 , P3_U5454 , P3_U5453 , P3_U5456 );
and AND2_1832 ( P3_U3641 , P3_U3640 , P3_U5455 );
and AND3_1833 ( P3_U3642 , P3_U5459 , P3_U5458 , P3_U5461 );
and AND2_1834 ( P3_U3643 , P3_U3642 , P3_U5460 );
and AND3_1835 ( P3_U3644 , P3_U5464 , P3_U5463 , P3_U5466 );
and AND2_1836 ( P3_U3645 , P3_U3644 , P3_U5465 );
and AND3_1837 ( P3_U3646 , P3_U5469 , P3_U5468 , P3_U5471 );
and AND2_1838 ( P3_U3647 , P3_U3646 , P3_U5470 );
and AND3_1839 ( P3_U3648 , P3_U5474 , P3_U5473 , P3_U5476 );
and AND2_1840 ( P3_U3649 , P3_U3648 , P3_U5475 );
and AND3_1841 ( P3_U3650 , P3_U5479 , P3_U5478 , P3_U5481 );
and AND2_1842 ( P3_U3651 , P3_U3650 , P3_U5480 );
and AND2_1843 ( P3_U3652 , P3_U4340 , P3_ADD_495_U8 );
and AND2_1844 ( P3_U3653 , P3_FLUSH_REG , P3_STATE2_REG_0_ );
and AND2_1845 ( P3_U3654 , P3_U4522 , P3_U3104 );
and AND2_1846 ( P3_U3655 , P3_U3107 , P3_U3118 );
and AND2_1847 ( P3_U3656 , P3_U5495 , P3_U4333 );
and AND2_1848 ( P3_U3657 , P3_U3656 , P3_U5494 );
and AND2_1849 ( P3_U3658 , P3_U5498 , P3_U4330 );
and AND2_1850 ( P3_U3659 , P3_U5502 , P3_U5501 );
and AND2_1851 ( P3_U3660 , P3_U4556 , P3_U4539 );
and AND2_1852 ( P3_U3661 , P3_U2461 , P3_U4297 );
and AND2_1853 ( P3_U3662 , P3_U4590 , P3_U3101 );
and AND2_1854 ( P3_U3663 , P3_U4556 , P3_U3101 );
and AND2_1855 ( P3_U3664 , P3_U4573 , P3_U4324 );
and AND3_1856 ( P3_U3665 , P3_U5511 , P3_U5510 , P3_U5508 );
and AND3_1857 ( P3_U3666 , P3_U5519 , P3_U4339 , P3_U5520 );
and AND4_1858 ( P3_U3667 , P3_U7978 , P3_U7977 , P3_U5521 , P3_U3666 );
and AND3_1859 ( P3_U3668 , P3_U5528 , P3_U3242 , P3_U2517 );
and AND2_1860 ( P3_U3669 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_U4470 );
and AND2_1861 ( P3_U3670 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_U3093 );
and AND3_1862 ( P3_U3671 , P3_U3116 , P3_U3117 , P3_U3119 );
and AND3_1863 ( P3_U3672 , P3_U3245 , P3_U3244 , P3_U3671 );
and AND2_1864 ( P3_U3673 , P3_U4505 , P3_U2456 );
and AND2_1865 ( P3_U3674 , P3_U5533 , P3_U5532 );
and AND2_1866 ( P3_U3675 , P3_U5538 , P3_U5536 );
and AND3_1867 ( P3_U3676 , P3_U3677 , P3_U5539 , P3_U3675 );
and AND2_1868 ( P3_U3677 , P3_U5540 , P3_U5541 );
and AND2_1869 ( P3_U3678 , P3_U5552 , P3_U5550 );
and AND2_1870 ( P3_U3679 , P3_U3678 , P3_U5551 );
and AND2_1871 ( P3_U3680 , P3_U5555 , P3_U5554 );
and AND2_1872 ( P3_U3681 , P3_U3682 , P3_U5562 );
and AND2_1873 ( P3_U3682 , P3_U5565 , P3_U5564 );
and AND2_1874 ( P3_U3683 , P3_U5568 , P3_U5567 );
and AND2_1875 ( P3_U3684 , P3_U5576 , P3_U5574 );
and AND2_1876 ( P3_U3685 , P3_U5587 , P3_U5588 );
and AND2_1877 ( P3_U3686 , P3_U5594 , P3_U5592 );
and AND3_1878 ( P3_U3687 , P3_U5625 , P3_U4333 , P3_U5626 );
and AND2_1879 ( P3_U3688 , P3_U2456 , P3_U4296 );
and AND2_1880 ( P3_U3689 , P3_U2456 , P3_U4323 );
and AND2_1881 ( P3_U3690 , P3_U4608 , P3_U4556 );
and AND2_1882 ( P3_U3691 , P3_U2456 , P3_U4590 );
and AND2_1883 ( P3_U3692 , P3_U5636 , P3_U5635 );
and AND5_1884 ( P3_U3693 , P3_U5638 , P3_U5637 , P3_U3694 , P3_U5633 , P3_U5632 );
and AND2_1885 ( P3_U3694 , P3_U3695 , P3_U5641 );
and AND2_1886 ( P3_U3695 , P3_U5639 , P3_U5640 );
and AND5_1887 ( P3_U3696 , P3_U5643 , P3_U5642 , P3_U5644 , P3_U5646 , P3_U5645 );
and AND5_1888 ( P3_U3697 , P3_U5648 , P3_U5649 , P3_U5647 , P3_U5651 , P3_U5650 );
and AND2_1889 ( P3_U3698 , P3_U3697 , P3_U3696 );
and AND2_1890 ( P3_U3699 , P3_U5660 , P3_U5659 );
and AND4_1891 ( P3_U3700 , P3_U5662 , P3_U5661 , P3_U3701 , P3_U5657 );
and AND2_1892 ( P3_U3701 , P3_U3702 , P3_U5665 );
and AND2_1893 ( P3_U3702 , P3_U5663 , P3_U5664 );
and AND5_1894 ( P3_U3703 , P3_U5667 , P3_U5666 , P3_U5668 , P3_U5670 , P3_U5669 );
and AND4_1895 ( P3_U3704 , P3_U5674 , P3_U5671 , P3_U5672 , P3_U5673 );
and AND3_1896 ( P3_U3705 , P3_U3704 , P3_U3703 , P3_U5675 );
and AND2_1897 ( P3_U3706 , P3_U3707 , P3_U5681 );
and AND2_1898 ( P3_U3707 , P3_U5684 , P3_U5683 );
and AND2_1899 ( P3_U3708 , P3_U3709 , P3_U5689 );
and AND2_1900 ( P3_U3709 , P3_U5687 , P3_U5688 );
and AND3_1901 ( P3_U3710 , P3_U5686 , P3_U5685 , P3_U3708 );
and AND5_1902 ( P3_U3711 , P3_U5691 , P3_U5690 , P3_U5692 , P3_U5694 , P3_U5693 );
and AND4_1903 ( P3_U3712 , P3_U5698 , P3_U5695 , P3_U5696 , P3_U5697 );
and AND3_1904 ( P3_U3713 , P3_U3712 , P3_U3711 , P3_U5699 );
and AND2_1905 ( P3_U3714 , P3_U5705 , P3_U5704 );
and AND2_1906 ( P3_U3715 , P3_U5708 , P3_U5707 );
and AND2_1907 ( P3_U3716 , P3_U3717 , P3_U5713 );
and AND2_1908 ( P3_U3717 , P3_U5711 , P3_U5712 );
and AND3_1909 ( P3_U3718 , P3_U5710 , P3_U5709 , P3_U3716 );
and AND5_1910 ( P3_U3719 , P3_U5715 , P3_U5714 , P3_U5716 , P3_U5718 , P3_U5717 );
and AND4_1911 ( P3_U3720 , P3_U5722 , P3_U5719 , P3_U5720 , P3_U5721 );
and AND3_1912 ( P3_U3721 , P3_U3720 , P3_U3719 , P3_U5723 );
and AND2_1913 ( P3_U3722 , P3_U3723 , P3_U5729 );
and AND2_1914 ( P3_U3723 , P3_U5732 , P3_U5731 );
and AND2_1915 ( P3_U3724 , P3_U3725 , P3_U5737 );
and AND2_1916 ( P3_U3725 , P3_U5735 , P3_U5736 );
and AND3_1917 ( P3_U3726 , P3_U5734 , P3_U5733 , P3_U3724 );
and AND5_1918 ( P3_U3727 , P3_U5739 , P3_U5738 , P3_U5740 , P3_U5742 , P3_U5741 );
and AND4_1919 ( P3_U3728 , P3_U5746 , P3_U5743 , P3_U5744 , P3_U5745 );
and AND3_1920 ( P3_U3729 , P3_U3728 , P3_U3727 , P3_U5747 );
and AND2_1921 ( P3_U3730 , P3_U3731 , P3_U5752 );
and AND2_1922 ( P3_U3731 , P3_U5756 , P3_U5755 );
and AND2_1923 ( P3_U3732 , P3_U3733 , P3_U5761 );
and AND2_1924 ( P3_U3733 , P3_U5759 , P3_U5760 );
and AND3_1925 ( P3_U3734 , P3_U5758 , P3_U5757 , P3_U3732 );
and AND5_1926 ( P3_U3735 , P3_U5763 , P3_U5762 , P3_U5764 , P3_U5766 , P3_U5765 );
and AND4_1927 ( P3_U3736 , P3_U5770 , P3_U5767 , P3_U5768 , P3_U5769 );
and AND3_1928 ( P3_U3737 , P3_U3736 , P3_U3735 , P3_U5771 );
and AND2_1929 ( P3_U3738 , P3_U3739 , P3_U5776 );
and AND2_1930 ( P3_U3739 , P3_U5780 , P3_U5779 );
and AND2_1931 ( P3_U3740 , P3_U3741 , P3_U5785 );
and AND2_1932 ( P3_U3741 , P3_U5783 , P3_U5784 );
and AND3_1933 ( P3_U3742 , P3_U5782 , P3_U5781 , P3_U3740 );
and AND5_1934 ( P3_U3743 , P3_U5787 , P3_U5786 , P3_U5788 , P3_U5790 , P3_U5789 );
and AND4_1935 ( P3_U3744 , P3_U5794 , P3_U5791 , P3_U5792 , P3_U5793 );
and AND3_1936 ( P3_U3745 , P3_U3744 , P3_U3743 , P3_U5795 );
and AND2_1937 ( P3_U3746 , P3_U3747 , P3_U5800 );
and AND2_1938 ( P3_U3747 , P3_U5804 , P3_U5803 );
and AND2_1939 ( P3_U3748 , P3_U3749 , P3_U5809 );
and AND2_1940 ( P3_U3749 , P3_U5807 , P3_U5808 );
and AND3_1941 ( P3_U3750 , P3_U5806 , P3_U5805 , P3_U3748 );
and AND5_1942 ( P3_U3751 , P3_U5811 , P3_U5810 , P3_U5812 , P3_U5814 , P3_U5813 );
and AND4_1943 ( P3_U3752 , P3_U5818 , P3_U5815 , P3_U5816 , P3_U5817 );
and AND3_1944 ( P3_U3753 , P3_U3752 , P3_U3751 , P3_U5819 );
and AND2_1945 ( P3_U3754 , P3_U3755 , P3_U5824 );
and AND2_1946 ( P3_U3755 , P3_U5828 , P3_U5827 );
and AND3_1947 ( P3_U3756 , P3_U5833 , P3_U5832 , P3_U5831 );
and AND3_1948 ( P3_U3757 , P3_U5830 , P3_U5829 , P3_U3756 );
and AND5_1949 ( P3_U3758 , P3_U5835 , P3_U5834 , P3_U5836 , P3_U5838 , P3_U5837 );
and AND4_1950 ( P3_U3759 , P3_U5842 , P3_U5841 , P3_U5840 , P3_U5839 );
and AND3_1951 ( P3_U3760 , P3_U3759 , P3_U3758 , P3_U5843 );
and AND2_1952 ( P3_U3761 , P3_U3762 , P3_U5848 );
and AND2_1953 ( P3_U3762 , P3_U5852 , P3_U5851 );
and AND2_1954 ( P3_U3763 , P3_U5857 , P3_U5856 );
and AND4_1955 ( P3_U3764 , P3_U5854 , P3_U5853 , P3_U5855 , P3_U3763 );
and AND5_1956 ( P3_U3765 , P3_U5859 , P3_U5858 , P3_U5860 , P3_U5862 , P3_U5861 );
and AND4_1957 ( P3_U3766 , P3_U5866 , P3_U5865 , P3_U5864 , P3_U5863 );
and AND3_1958 ( P3_U3767 , P3_U3766 , P3_U3765 , P3_U5867 );
and AND2_1959 ( P3_U3768 , P3_U3769 , P3_U5873 );
and AND2_1960 ( P3_U3769 , P3_U5876 , P3_U5875 );
and AND2_1961 ( P3_U3770 , P3_U5881 , P3_U5880 );
and AND4_1962 ( P3_U3771 , P3_U5878 , P3_U5877 , P3_U5879 , P3_U3770 );
and AND5_1963 ( P3_U3772 , P3_U5883 , P3_U5882 , P3_U5884 , P3_U5886 , P3_U5885 );
and AND4_1964 ( P3_U3773 , P3_U5890 , P3_U5889 , P3_U5888 , P3_U5887 );
and AND3_1965 ( P3_U3774 , P3_U3773 , P3_U3772 , P3_U5891 );
and AND2_1966 ( P3_U3775 , P3_U3776 , P3_U5897 );
and AND2_1967 ( P3_U3776 , P3_U5900 , P3_U5899 );
and AND2_1968 ( P3_U3777 , P3_U5905 , P3_U5904 );
and AND4_1969 ( P3_U3778 , P3_U5902 , P3_U5901 , P3_U5903 , P3_U3777 );
and AND5_1970 ( P3_U3779 , P3_U5907 , P3_U5906 , P3_U5908 , P3_U5910 , P3_U5909 );
and AND4_1971 ( P3_U3780 , P3_U5914 , P3_U5913 , P3_U5912 , P3_U5911 );
and AND3_1972 ( P3_U3781 , P3_U3780 , P3_U3779 , P3_U5915 );
and AND2_1973 ( P3_U3782 , P3_U3783 , P3_U5920 );
and AND2_1974 ( P3_U3783 , P3_U5924 , P3_U5923 );
and AND2_1975 ( P3_U3784 , P3_U5929 , P3_U5928 );
and AND4_1976 ( P3_U3785 , P3_U5926 , P3_U5925 , P3_U5927 , P3_U3784 );
and AND5_1977 ( P3_U3786 , P3_U5931 , P3_U5930 , P3_U5932 , P3_U5934 , P3_U5933 );
and AND4_1978 ( P3_U3787 , P3_U5938 , P3_U5937 , P3_U5936 , P3_U5935 );
and AND3_1979 ( P3_U3788 , P3_U3787 , P3_U3786 , P3_U5939 );
and AND2_1980 ( P3_U3789 , P3_U3790 , P3_U5944 );
and AND2_1981 ( P3_U3790 , P3_U5948 , P3_U5947 );
and AND2_1982 ( P3_U3791 , P3_U5953 , P3_U5952 );
and AND4_1983 ( P3_U3792 , P3_U5950 , P3_U5949 , P3_U5951 , P3_U3791 );
and AND5_1984 ( P3_U3793 , P3_U5955 , P3_U5954 , P3_U5956 , P3_U5958 , P3_U5957 );
and AND4_1985 ( P3_U3794 , P3_U5962 , P3_U5961 , P3_U5960 , P3_U5959 );
and AND3_1986 ( P3_U3795 , P3_U3794 , P3_U3793 , P3_U5963 );
and AND2_1987 ( P3_U3796 , P3_U5972 , P3_U5971 );
and AND2_1988 ( P3_U3797 , P3_U5977 , P3_U5976 );
and AND4_1989 ( P3_U3798 , P3_U5974 , P3_U5973 , P3_U5975 , P3_U3797 );
and AND5_1990 ( P3_U3799 , P3_U3796 , P3_U5970 , P3_U3798 , P3_U5969 , P3_U5968 );
and AND5_1991 ( P3_U3800 , P3_U5979 , P3_U5978 , P3_U5980 , P3_U5982 , P3_U5981 );
and AND4_1992 ( P3_U3801 , P3_U5986 , P3_U5985 , P3_U5984 , P3_U5983 );
and AND3_1993 ( P3_U3802 , P3_U3801 , P3_U3800 , P3_U5987 );
and AND2_1994 ( P3_U3803 , P3_U5991 , P3_U5989 );
and AND2_1995 ( P3_U3804 , P3_U5996 , P3_U5995 );
and AND2_1996 ( P3_U3805 , P3_U6001 , P3_U6000 );
and AND4_1997 ( P3_U3806 , P3_U5998 , P3_U5997 , P3_U5999 , P3_U3805 );
and AND5_1998 ( P3_U3807 , P3_U3804 , P3_U5994 , P3_U3806 , P3_U5993 , P3_U5992 );
and AND5_1999 ( P3_U3808 , P3_U6003 , P3_U6002 , P3_U6004 , P3_U6006 , P3_U6005 );
and AND4_2000 ( P3_U3809 , P3_U6010 , P3_U6009 , P3_U6008 , P3_U6007 );
and AND3_2001 ( P3_U3810 , P3_U3809 , P3_U3808 , P3_U6011 );
and AND2_2002 ( P3_U3811 , P3_U6015 , P3_U6013 );
and AND2_2003 ( P3_U3812 , P3_U3813 , P3_U6017 );
and AND2_2004 ( P3_U3813 , P3_U6020 , P3_U6019 );
and AND2_2005 ( P3_U3814 , P3_U6025 , P3_U6024 );
and AND4_2006 ( P3_U3815 , P3_U6022 , P3_U6021 , P3_U6023 , P3_U3814 );
and AND5_2007 ( P3_U3816 , P3_U6027 , P3_U6026 , P3_U6028 , P3_U6030 , P3_U6029 );
and AND4_2008 ( P3_U3817 , P3_U6034 , P3_U6033 , P3_U6032 , P3_U6031 );
and AND3_2009 ( P3_U3818 , P3_U3817 , P3_U3816 , P3_U6035 );
and AND2_2010 ( P3_U3819 , P3_U6044 , P3_U6043 );
and AND5_2011 ( P3_U3820 , P3_U6046 , P3_U6045 , P3_U6047 , P3_U3821 , P3_U6041 );
and AND2_2012 ( P3_U3821 , P3_U6049 , P3_U6048 );
and AND5_2013 ( P3_U3822 , P3_U6051 , P3_U6050 , P3_U6052 , P3_U6054 , P3_U6053 );
and AND4_2014 ( P3_U3823 , P3_U6058 , P3_U6057 , P3_U6056 , P3_U6055 );
and AND3_2015 ( P3_U3824 , P3_U3823 , P3_U3822 , P3_U6059 );
and AND2_2016 ( P3_U3825 , P3_U3826 , P3_U6065 );
and AND2_2017 ( P3_U3826 , P3_U6068 , P3_U6067 );
and AND2_2018 ( P3_U3827 , P3_U6073 , P3_U6072 );
and AND4_2019 ( P3_U3828 , P3_U6070 , P3_U6069 , P3_U6071 , P3_U3827 );
and AND5_2020 ( P3_U3829 , P3_U6075 , P3_U6074 , P3_U6076 , P3_U6078 , P3_U6077 );
and AND4_2021 ( P3_U3830 , P3_U6082 , P3_U6081 , P3_U6080 , P3_U6079 );
and AND3_2022 ( P3_U3831 , P3_U3830 , P3_U3829 , P3_U6083 );
and AND2_2023 ( P3_U3832 , P3_U6092 , P3_U6091 );
and AND5_2024 ( P3_U3833 , P3_U6094 , P3_U6093 , P3_U6095 , P3_U3834 , P3_U6089 );
and AND2_2025 ( P3_U3834 , P3_U6097 , P3_U6096 );
and AND5_2026 ( P3_U3835 , P3_U6099 , P3_U6098 , P3_U6100 , P3_U6102 , P3_U6101 );
and AND4_2027 ( P3_U3836 , P3_U6106 , P3_U6105 , P3_U6104 , P3_U6103 );
and AND3_2028 ( P3_U3837 , P3_U3836 , P3_U3835 , P3_U6107 );
and AND2_2029 ( P3_U3838 , P3_U6116 , P3_U6115 );
and AND2_2030 ( P3_U3839 , P3_U6121 , P3_U6120 );
and AND4_2031 ( P3_U3840 , P3_U6118 , P3_U6117 , P3_U6119 , P3_U3839 );
and AND5_2032 ( P3_U3841 , P3_U6114 , P3_U3838 , P3_U3840 , P3_U6112 , P3_U3844 );
and AND5_2033 ( P3_U3842 , P3_U6123 , P3_U6122 , P3_U6124 , P3_U6126 , P3_U6125 );
and AND4_2034 ( P3_U3843 , P3_U6130 , P3_U6129 , P3_U6128 , P3_U6127 );
and AND3_2035 ( P3_U3844 , P3_U3843 , P3_U3842 , P3_U6131 );
and AND2_2036 ( P3_U3845 , P3_U6135 , P3_U6133 );
and AND2_2037 ( P3_U3846 , P3_U6140 , P3_U6139 );
and AND2_2038 ( P3_U3847 , P3_U6145 , P3_U6144 );
and AND4_2039 ( P3_U3848 , P3_U6142 , P3_U6141 , P3_U6143 , P3_U3847 );
and AND5_2040 ( P3_U3849 , P3_U6138 , P3_U3846 , P3_U3848 , P3_U6136 , P3_U3852 );
and AND5_2041 ( P3_U3850 , P3_U6147 , P3_U6146 , P3_U6148 , P3_U6150 , P3_U6149 );
and AND4_2042 ( P3_U3851 , P3_U6154 , P3_U6153 , P3_U6152 , P3_U6151 );
and AND3_2043 ( P3_U3852 , P3_U3850 , P3_U3851 , P3_U6155 );
and AND2_2044 ( P3_U3853 , P3_U6159 , P3_U6157 );
and AND2_2045 ( P3_U3854 , P3_U6164 , P3_U6163 );
and AND2_2046 ( P3_U3855 , P3_U6169 , P3_U6168 );
and AND4_2047 ( P3_U3856 , P3_U6166 , P3_U6165 , P3_U6167 , P3_U3855 );
and AND5_2048 ( P3_U3857 , P3_U6161 , P3_U6162 , P3_U3854 , P3_U3856 , P3_U6160 );
and AND3_2049 ( P3_U3858 , P3_U6171 , P3_U6170 , P3_U6172 );
and AND2_2050 ( P3_U3859 , P3_U6174 , P3_U6173 );
and AND3_2051 ( P3_U3860 , P3_U6176 , P3_U6175 , P3_U6177 );
and AND2_2052 ( P3_U3861 , P3_U6179 , P3_U6178 );
and AND4_2053 ( P3_U3862 , P3_U3859 , P3_U3858 , P3_U3860 , P3_U3861 );
and AND2_2054 ( P3_U3863 , P3_U6183 , P3_U6181 );
and AND2_2055 ( P3_U3864 , P3_U6188 , P3_U6187 );
and AND2_2056 ( P3_U3865 , P3_U6193 , P3_U6192 );
and AND4_2057 ( P3_U3866 , P3_U6190 , P3_U6189 , P3_U6191 , P3_U3865 );
and AND5_2058 ( P3_U3867 , P3_U6185 , P3_U6186 , P3_U3864 , P3_U3866 , P3_U6184 );
and AND3_2059 ( P3_U3868 , P3_U6195 , P3_U6194 , P3_U6196 );
and AND2_2060 ( P3_U3869 , P3_U6198 , P3_U6197 );
and AND3_2061 ( P3_U3870 , P3_U6200 , P3_U6199 , P3_U6201 );
and AND2_2062 ( P3_U3871 , P3_U6203 , P3_U6202 );
and AND4_2063 ( P3_U3872 , P3_U3869 , P3_U3868 , P3_U3870 , P3_U3871 );
and AND2_2064 ( P3_U3873 , P3_U6207 , P3_U6205 );
and AND2_2065 ( P3_U3874 , P3_U6212 , P3_U6211 );
and AND2_2066 ( P3_U3875 , P3_U6217 , P3_U6216 );
and AND4_2067 ( P3_U3876 , P3_U6214 , P3_U6213 , P3_U6215 , P3_U3875 );
and AND5_2068 ( P3_U3877 , P3_U6209 , P3_U6210 , P3_U3874 , P3_U6208 , P3_U3876 );
and AND3_2069 ( P3_U3878 , P3_U6219 , P3_U6218 , P3_U6220 );
and AND2_2070 ( P3_U3879 , P3_U6222 , P3_U6221 );
and AND3_2071 ( P3_U3880 , P3_U6224 , P3_U6223 , P3_U6225 );
and AND2_2072 ( P3_U3881 , P3_U6227 , P3_U6226 );
and AND4_2073 ( P3_U3882 , P3_U3879 , P3_U3878 , P3_U3881 , P3_U3880 );
and AND2_2074 ( P3_U3883 , P3_U6231 , P3_U6229 );
and AND2_2075 ( P3_U3884 , P3_U6236 , P3_U6235 );
and AND2_2076 ( P3_U3885 , P3_U6241 , P3_U6240 );
and AND4_2077 ( P3_U3886 , P3_U6238 , P3_U6237 , P3_U6239 , P3_U3885 );
and AND5_2078 ( P3_U3887 , P3_U6233 , P3_U6234 , P3_U6232 , P3_U3884 , P3_U3886 );
and AND3_2079 ( P3_U3888 , P3_U6243 , P3_U6242 , P3_U6244 );
and AND2_2080 ( P3_U3889 , P3_U6246 , P3_U6245 );
and AND3_2081 ( P3_U3890 , P3_U6248 , P3_U6247 , P3_U6249 );
and AND2_2082 ( P3_U3891 , P3_U6251 , P3_U6250 );
and AND4_2083 ( P3_U3892 , P3_U3889 , P3_U3888 , P3_U3891 , P3_U3890 );
and AND2_2084 ( P3_U3893 , P3_U6255 , P3_U6253 );
and AND2_2085 ( P3_U3894 , P3_U6257 , P3_U6256 );
and AND2_2086 ( P3_U3895 , P3_U6260 , P3_U6259 );
and AND2_2087 ( P3_U3896 , P3_U6265 , P3_U6264 );
and AND4_2088 ( P3_U3897 , P3_U6262 , P3_U6261 , P3_U6263 , P3_U3896 );
and AND3_2089 ( P3_U3898 , P3_U6267 , P3_U6266 , P3_U6268 );
and AND2_2090 ( P3_U3899 , P3_U6270 , P3_U6269 );
and AND3_2091 ( P3_U3900 , P3_U6272 , P3_U6271 , P3_U6273 );
and AND2_2092 ( P3_U3901 , P3_U6275 , P3_U6274 );
and AND4_2093 ( P3_U3902 , P3_U3899 , P3_U3898 , P3_U3901 , P3_U3900 );
and AND2_2094 ( P3_U3903 , P3_U6281 , P3_U6280 );
and AND2_2095 ( P3_U3904 , P3_U6284 , P3_U6283 );
and AND2_2096 ( P3_U3905 , P3_U6289 , P3_U6288 );
and AND4_2097 ( P3_U3906 , P3_U6286 , P3_U6285 , P3_U6287 , P3_U3905 );
and AND3_2098 ( P3_U3907 , P3_U6291 , P3_U6290 , P3_U6292 );
and AND2_2099 ( P3_U3908 , P3_U6294 , P3_U6293 );
and AND3_2100 ( P3_U3909 , P3_U6296 , P3_U6295 , P3_U6297 );
and AND2_2101 ( P3_U3910 , P3_U6299 , P3_U6298 );
and AND4_2102 ( P3_U3911 , P3_U3908 , P3_U3907 , P3_U3910 , P3_U3909 );
and AND2_2103 ( P3_U3912 , P3_U6305 , P3_U6304 );
and AND2_2104 ( P3_U3913 , P3_U6308 , P3_U6307 );
and AND2_2105 ( P3_U3914 , P3_U6313 , P3_U6312 );
and AND4_2106 ( P3_U3915 , P3_U6310 , P3_U6309 , P3_U6311 , P3_U3914 );
and AND3_2107 ( P3_U3916 , P3_U6315 , P3_U6314 , P3_U6316 );
and AND2_2108 ( P3_U3917 , P3_U6318 , P3_U6317 );
and AND3_2109 ( P3_U3918 , P3_U6320 , P3_U6319 , P3_U6321 );
and AND2_2110 ( P3_U3919 , P3_U6323 , P3_U6322 );
and AND4_2111 ( P3_U3920 , P3_U3917 , P3_U3916 , P3_U3919 , P3_U3918 );
and AND2_2112 ( P3_U3921 , P3_U6329 , P3_U6328 );
and AND2_2113 ( P3_U3922 , P3_U6332 , P3_U6331 );
and AND2_2114 ( P3_U3923 , P3_U6337 , P3_U6336 );
and AND4_2115 ( P3_U3924 , P3_U6334 , P3_U6333 , P3_U6335 , P3_U3923 );
and AND3_2116 ( P3_U3925 , P3_U6339 , P3_U6338 , P3_U6340 );
and AND2_2117 ( P3_U3926 , P3_U6342 , P3_U6341 );
and AND3_2118 ( P3_U3927 , P3_U6344 , P3_U6343 , P3_U6345 );
and AND2_2119 ( P3_U3928 , P3_U6347 , P3_U6346 );
and AND4_2120 ( P3_U3929 , P3_U3926 , P3_U3925 , P3_U3928 , P3_U3927 );
and AND2_2121 ( P3_U3930 , P3_U6353 , P3_U6352 );
and AND2_2122 ( P3_U3931 , P3_U6356 , P3_U6355 );
and AND2_2123 ( P3_U3932 , P3_U6361 , P3_U6360 );
and AND4_2124 ( P3_U3933 , P3_U6358 , P3_U6357 , P3_U6359 , P3_U3932 );
and AND3_2125 ( P3_U3934 , P3_U6363 , P3_U6362 , P3_U6364 );
and AND2_2126 ( P3_U3935 , P3_U6366 , P3_U6365 );
and AND3_2127 ( P3_U3936 , P3_U6368 , P3_U6367 , P3_U6369 );
and AND2_2128 ( P3_U3937 , P3_U6371 , P3_U6370 );
and AND4_2129 ( P3_U3938 , P3_U3935 , P3_U3934 , P3_U3937 , P3_U3936 );
and AND2_2130 ( P3_U3939 , P3_U6398 , P3_U3247 );
and AND2_2131 ( P3_U3940 , P3_U6377 , P3_U6376 );
and AND2_2132 ( P3_U3941 , P3_U6380 , P3_U6379 );
and AND2_2133 ( P3_U3942 , P3_U3941 , P3_U6381 );
and AND3_2134 ( P3_U3943 , P3_U6386 , P3_U6385 , P3_U6384 );
and AND3_2135 ( P3_U3944 , P3_U6383 , P3_U6382 , P3_U3943 );
and AND4_2136 ( P3_U3945 , P3_U3940 , P3_U6378 , P3_U3942 , P3_U3944 );
and AND3_2137 ( P3_U3946 , P3_U6388 , P3_U6387 , P3_U6389 );
and AND2_2138 ( P3_U3947 , P3_U6391 , P3_U6390 );
and AND3_2139 ( P3_U3948 , P3_U3946 , P3_U6392 , P3_U3947 );
and AND2_2140 ( P3_U3949 , P3_U6394 , P3_U6393 );
and AND5_2141 ( P3_U3950 , P3_U6398 , P3_U6397 , P3_U6395 , P3_U3949 , P3_U3948 );
and AND2_2142 ( P3_U3951 , P3_STATE2_REG_0_ , P3_U3104 );
and AND2_2143 ( P3_U3952 , P3_STATE2_REG_2_ , P3_U3121 );
and AND2_2144 ( P3_U3953 , P3_U4505 , P3_STATE2_REG_0_ );
and AND4_2145 ( P3_U3954 , P3_U6412 , P3_U6411 , P3_U6410 , P3_U6409 );
and AND4_2146 ( P3_U3955 , P3_U6420 , P3_U6419 , P3_U6418 , P3_U6417 );
and AND4_2147 ( P3_U3956 , P3_U6426 , P3_U6425 , P3_U6428 , P3_U6427 );
and AND4_2148 ( P3_U3957 , P3_U6434 , P3_U6433 , P3_U6436 , P3_U6435 );
and AND4_2149 ( P3_U3958 , P3_U6442 , P3_U6441 , P3_U6444 , P3_U6443 );
and AND4_2150 ( P3_U3959 , P3_U6450 , P3_U6449 , P3_U6452 , P3_U6451 );
and AND4_2151 ( P3_U3960 , P3_U6458 , P3_U6457 , P3_U6460 , P3_U6459 );
and AND4_2152 ( P3_U3961 , P3_U6466 , P3_U6465 , P3_U6468 , P3_U6467 );
and AND4_2153 ( P3_U3962 , P3_U6474 , P3_U6473 , P3_U6476 , P3_U6475 );
and AND4_2154 ( P3_U3963 , P3_U6482 , P3_U6481 , P3_U6484 , P3_U6483 );
and AND4_2155 ( P3_U3964 , P3_U6490 , P3_U6489 , P3_U6492 , P3_U6491 );
and AND4_2156 ( P3_U3965 , P3_U6498 , P3_U6497 , P3_U6500 , P3_U6499 );
and AND4_2157 ( P3_U3966 , P3_U6508 , P3_U6505 , P3_U6506 , P3_U6507 );
and AND4_2158 ( P3_U3967 , P3_U6516 , P3_U6513 , P3_U6514 , P3_U6515 );
and AND4_2159 ( P3_U3968 , P3_U6524 , P3_U6521 , P3_U6522 , P3_U6523 );
and AND4_2160 ( P3_U3969 , P3_U6532 , P3_U6529 , P3_U6530 , P3_U6531 );
and AND4_2161 ( P3_U3970 , P3_U6540 , P3_U6537 , P3_U6538 , P3_U6539 );
and AND4_2162 ( P3_U3971 , P3_U6548 , P3_U6545 , P3_U6546 , P3_U6547 );
and AND4_2163 ( P3_U3972 , P3_U6556 , P3_U6553 , P3_U6554 , P3_U6555 );
and AND4_2164 ( P3_U3973 , P3_U6564 , P3_U6561 , P3_U6562 , P3_U6563 );
and AND4_2165 ( P3_U3974 , P3_U6572 , P3_U6569 , P3_U6570 , P3_U6571 );
and AND4_2166 ( P3_U3975 , P3_U6580 , P3_U6577 , P3_U6578 , P3_U6579 );
and AND4_2167 ( P3_U3976 , P3_U6588 , P3_U6585 , P3_U6586 , P3_U6587 );
and AND4_2168 ( P3_U3977 , P3_U6596 , P3_U6593 , P3_U6594 , P3_U6595 );
and AND4_2169 ( P3_U3978 , P3_U6604 , P3_U6601 , P3_U6602 , P3_U6603 );
and AND4_2170 ( P3_U3979 , P3_U6612 , P3_U6609 , P3_U6610 , P3_U6611 );
and AND4_2171 ( P3_U3980 , P3_U6620 , P3_U6619 , P3_U6618 , P3_U6617 );
and AND4_2172 ( P3_U3981 , P3_U6628 , P3_U6627 , P3_U6626 , P3_U6625 );
and AND4_2173 ( P3_U3982 , P3_U6636 , P3_U6635 , P3_U6634 , P3_U6633 );
and AND4_2174 ( P3_U3983 , P3_U6644 , P3_U6641 , P3_U6643 , P3_U6642 );
and AND4_2175 ( P3_U3984 , P3_U6652 , P3_U6649 , P3_U6651 , P3_U6650 );
and AND4_2176 ( P3_U3985 , P3_U6660 , P3_U6657 , P3_U6659 , P3_U6658 );
and AND2_2177 ( P3_U3986 , P3_U4293 , P3_U2390 );
and AND2_2178 ( P3_U3987 , P3_U6809 , P3_U6810 );
and AND2_2179 ( P3_U3988 , P3_U6812 , P3_U6813 );
and AND2_2180 ( P3_U3989 , P3_U6815 , P3_U6816 );
and AND2_2181 ( P3_U3990 , P3_U6818 , P3_U6819 );
and AND2_2182 ( P3_U3991 , P3_U6821 , P3_U6822 );
and AND2_2183 ( P3_U3992 , P3_U6824 , P3_U6825 );
and AND2_2184 ( P3_U3993 , P3_U6827 , P3_U6828 );
and AND2_2185 ( P3_U3994 , P3_U6830 , P3_U6831 );
and AND2_2186 ( P3_U3995 , P3_U6833 , P3_U6834 );
and AND2_2187 ( P3_U3996 , P3_U6836 , P3_U6837 );
and AND2_2188 ( P3_U3997 , P3_U6839 , P3_U6840 );
and AND2_2189 ( P3_U3998 , P3_U6842 , P3_U6843 );
and AND2_2190 ( P3_U3999 , P3_U6845 , P3_U6846 );
and AND2_2191 ( P3_U4000 , P3_U6848 , P3_U6849 );
and AND2_2192 ( P3_U4001 , P3_U6851 , P3_U6852 );
and AND2_2193 ( P3_U4002 , P3_U6857 , P3_U6856 );
and AND2_2194 ( P3_U4003 , P3_U6861 , P3_U6860 );
and AND2_2195 ( P3_U4004 , P3_U6865 , P3_U6864 );
and AND2_2196 ( P3_U4005 , P3_U6869 , P3_U6868 );
and AND2_2197 ( P3_U4006 , P3_U6873 , P3_U6872 );
and AND2_2198 ( P3_U4007 , P3_U6877 , P3_U6876 );
and AND2_2199 ( P3_U4008 , P3_U6881 , P3_U6880 );
and AND2_2200 ( P3_U4009 , P3_U6885 , P3_U6884 );
and AND2_2201 ( P3_U4010 , P3_U6889 , P3_U6888 );
and AND2_2202 ( P3_U4011 , P3_U6893 , P3_U6892 );
and AND2_2203 ( P3_U4012 , P3_U6897 , P3_U6896 );
and AND2_2204 ( P3_U4013 , P3_U6901 , P3_U6900 );
and AND2_2205 ( P3_U4014 , P3_U6905 , P3_U6904 );
and AND2_2206 ( P3_U4015 , P3_U6907 , P3_U6909 );
and AND2_2207 ( P3_U4016 , P3_U6911 , P3_U6913 );
and AND2_2208 ( P3_U4017 , P3_U6915 , P3_U6917 );
and AND2_2209 ( P3_U4018 , P3_U6922 , P3_U6920 );
and AND2_2210 ( P3_U4019 , P3_U6927 , P3_U6925 );
and AND2_2211 ( P3_U4020 , P3_U6932 , P3_U6930 );
and AND2_2212 ( P3_U4021 , P3_U6937 , P3_U6935 );
and AND2_2213 ( P3_U4022 , P3_U6942 , P3_U6940 );
and AND2_2214 ( P3_U4023 , P3_U6947 , P3_U6945 );
and AND2_2215 ( P3_U4024 , P3_U6952 , P3_U6950 );
and AND2_2216 ( P3_U4025 , P3_U6957 , P3_U6955 );
and AND2_2217 ( P3_U4026 , P3_U6962 , P3_U6960 );
and AND2_2218 ( P3_U4027 , P3_U6967 , P3_U6965 );
and AND2_2219 ( P3_U4028 , P3_U6972 , P3_U6970 );
and AND2_2220 ( P3_U4029 , P3_U6977 , P3_U6975 );
and AND3_2221 ( P3_U4030 , P3_U4329 , P3_U4328 , P3_U4336 );
and AND3_2222 ( P3_U4031 , P3_U7098 , P3_U7097 , P3_U4032 );
and AND2_2223 ( P3_U4032 , P3_U7101 , P3_U7100 );
and AND2_2224 ( P3_U4033 , P3_U4034 , P3_U7104 );
and AND2_2225 ( P3_U4034 , P3_U7106 , P3_U7105 );
and AND3_2226 ( P3_U4035 , P3_U7108 , P3_U7107 , P3_U4036 );
and AND2_2227 ( P3_U4036 , P3_U7111 , P3_U7110 );
and AND2_2228 ( P3_U4037 , P3_U4038 , P3_U7114 );
and AND2_2229 ( P3_U4038 , P3_U7116 , P3_U7115 );
and AND3_2230 ( P3_U4039 , P3_U7118 , P3_U7117 , P3_U4040 );
and AND2_2231 ( P3_U4040 , P3_U7121 , P3_U7120 );
and AND2_2232 ( P3_U4041 , P3_U4042 , P3_U7124 );
and AND2_2233 ( P3_U4042 , P3_U7126 , P3_U7125 );
and AND3_2234 ( P3_U4043 , P3_U7128 , P3_U7127 , P3_U4044 );
and AND2_2235 ( P3_U4044 , P3_U7131 , P3_U7130 );
and AND2_2236 ( P3_U4045 , P3_U4046 , P3_U7134 );
and AND2_2237 ( P3_U4046 , P3_U7136 , P3_U7135 );
and AND3_2238 ( P3_U4047 , P3_U7137 , P3_U4316 , P3_U7138 );
and AND2_2239 ( P3_U4048 , P3_U7140 , P3_U7141 );
and AND2_2240 ( P3_U4049 , P3_U4050 , P3_U7144 );
and AND2_2241 ( P3_U4050 , P3_U7146 , P3_U7145 );
and AND5_2242 ( P3_U4051 , P3_U4048 , P3_U7139 , P3_U4047 , P3_U7142 , P3_U7143 );
and AND3_2243 ( P3_U4052 , P3_U7147 , P3_U4316 , P3_U7148 );
and AND2_2244 ( P3_U4053 , P3_U7150 , P3_U7151 );
and AND2_2245 ( P3_U4054 , P3_U4055 , P3_U7154 );
and AND2_2246 ( P3_U4055 , P3_U7156 , P3_U7155 );
and AND5_2247 ( P3_U4056 , P3_U4053 , P3_U7149 , P3_U4052 , P3_U7152 , P3_U7153 );
and AND3_2248 ( P3_U4057 , P3_U7157 , P3_U4316 , P3_U7158 );
and AND2_2249 ( P3_U4058 , P3_U4059 , P3_U7161 );
and AND2_2250 ( P3_U4059 , P3_U7164 , P3_U7163 );
and AND3_2251 ( P3_U4060 , P3_U7165 , P3_U4316 , P3_U7166 );
and AND2_2252 ( P3_U4061 , P3_U4062 , P3_U7169 );
and AND2_2253 ( P3_U4062 , P3_U7172 , P3_U7171 );
and AND3_2254 ( P3_U4063 , P3_U7173 , P3_U4316 , P3_U7174 );
and AND2_2255 ( P3_U4064 , P3_U4065 , P3_U7177 );
and AND2_2256 ( P3_U4065 , P3_U7180 , P3_U7179 );
and AND3_2257 ( P3_U4066 , P3_U7181 , P3_U4316 , P3_U7182 );
and AND2_2258 ( P3_U4067 , P3_U4068 , P3_U7185 );
and AND2_2259 ( P3_U4068 , P3_U7188 , P3_U7187 );
and AND3_2260 ( P3_U4069 , P3_U7189 , P3_U4316 , P3_U7190 );
and AND2_2261 ( P3_U4070 , P3_U4071 , P3_U7193 );
and AND2_2262 ( P3_U4071 , P3_U7196 , P3_U7195 );
and AND3_2263 ( P3_U4072 , P3_U7197 , P3_U4316 , P3_U7198 );
and AND2_2264 ( P3_U4073 , P3_U4074 , P3_U7201 );
and AND2_2265 ( P3_U4074 , P3_U7204 , P3_U7203 );
and AND3_2266 ( P3_U4075 , P3_U7205 , P3_U4316 , P3_U7206 );
and AND2_2267 ( P3_U4076 , P3_U4077 , P3_U7209 );
and AND2_2268 ( P3_U4077 , P3_U7212 , P3_U7211 );
and AND3_2269 ( P3_U4078 , P3_U7213 , P3_U4316 , P3_U7214 );
and AND2_2270 ( P3_U4079 , P3_U4080 , P3_U7217 );
and AND2_2271 ( P3_U4080 , P3_U7220 , P3_U7219 );
and AND3_2272 ( P3_U4081 , P3_U7221 , P3_U4316 , P3_U7222 );
and AND2_2273 ( P3_U4082 , P3_U4083 , P3_U7225 );
and AND2_2274 ( P3_U4083 , P3_U7228 , P3_U7227 );
and AND3_2275 ( P3_U4084 , P3_U7229 , P3_U4316 , P3_U7230 );
and AND2_2276 ( P3_U4085 , P3_U4086 , P3_U7233 );
and AND2_2277 ( P3_U4086 , P3_U7236 , P3_U7235 );
and AND3_2278 ( P3_U4087 , P3_U7237 , P3_U4316 , P3_U7238 );
and AND2_2279 ( P3_U4088 , P3_U4089 , P3_U7241 );
and AND2_2280 ( P3_U4089 , P3_U7244 , P3_U7243 );
and AND3_2281 ( P3_U4090 , P3_U7245 , P3_U4316 , P3_U7246 );
and AND2_2282 ( P3_U4091 , P3_U4092 , P3_U7249 );
and AND2_2283 ( P3_U4092 , P3_U7252 , P3_U7251 );
and AND3_2284 ( P3_U4093 , P3_U7253 , P3_U4316 , P3_U7254 );
and AND2_2285 ( P3_U4094 , P3_U4095 , P3_U7257 );
and AND2_2286 ( P3_U4095 , P3_U7260 , P3_U7259 );
and AND3_2287 ( P3_U4096 , P3_U7261 , P3_U4316 , P3_U7262 );
and AND2_2288 ( P3_U4097 , P3_U4098 , P3_U7265 );
and AND2_2289 ( P3_U4098 , P3_U7268 , P3_U7267 );
and AND2_2290 ( P3_U4099 , P3_U7270 , P3_U7269 );
and AND2_2291 ( P3_U4100 , P3_U4101 , P3_U7273 );
and AND2_2292 ( P3_U4101 , P3_U7276 , P3_U7275 );
and AND2_2293 ( P3_U4102 , P3_U7278 , P3_U7277 );
and AND2_2294 ( P3_U4103 , P3_U4104 , P3_U7281 );
and AND2_2295 ( P3_U4104 , P3_U7284 , P3_U7283 );
and AND2_2296 ( P3_U4105 , P3_U7286 , P3_U7285 );
and AND2_2297 ( P3_U4106 , P3_U4107 , P3_U7289 );
and AND2_2298 ( P3_U4107 , P3_U7292 , P3_U7291 );
and AND2_2299 ( P3_U4108 , P3_U7294 , P3_U7293 );
and AND2_2300 ( P3_U4109 , P3_U4110 , P3_U7297 );
and AND2_2301 ( P3_U4110 , P3_U7300 , P3_U7299 );
and AND2_2302 ( P3_U4111 , P3_U7302 , P3_U7301 );
and AND2_2303 ( P3_U4112 , P3_U4113 , P3_U7305 );
and AND2_2304 ( P3_U4113 , P3_U7308 , P3_U7307 );
and AND2_2305 ( P3_U4114 , P3_U7310 , P3_U7309 );
and AND2_2306 ( P3_U4115 , P3_U4116 , P3_U7313 );
and AND2_2307 ( P3_U4116 , P3_U7316 , P3_U7315 );
and AND2_2308 ( P3_U4117 , P3_U7318 , P3_U7317 );
and AND2_2309 ( P3_U4118 , P3_U4119 , P3_U7321 );
and AND2_2310 ( P3_U4119 , P3_U7324 , P3_U7323 );
and AND2_2311 ( P3_U4120 , P3_U7326 , P3_U7325 );
and AND2_2312 ( P3_U4121 , P3_U4122 , P3_U7329 );
and AND2_2313 ( P3_U4122 , P3_U7332 , P3_U7331 );
and AND2_2314 ( P3_U4123 , P3_U7334 , P3_U7333 );
and AND2_2315 ( P3_U4124 , P3_U4125 , P3_U7337 );
and AND2_2316 ( P3_U4125 , P3_U7340 , P3_U7339 );
and AND2_2317 ( P3_U4126 , P3_U7342 , P3_U7341 );
and AND2_2318 ( P3_U4127 , P3_U4128 , P3_U7345 );
and AND2_2319 ( P3_U4128 , P3_U7348 , P3_U7347 );
and AND2_2320 ( P3_U4129 , P3_U7350 , P3_U7349 );
and AND2_2321 ( P3_U4130 , P3_U4131 , P3_U7353 );
and AND2_2322 ( P3_U4131 , P3_U7356 , P3_U7355 );
and AND2_2323 ( P3_U4132 , P3_U7364 , P3_U7365 );
and AND2_2324 ( P3_U4133 , P3_U4132 , P3_U7361 );
and AND2_2325 ( P3_U4134 , P3_U7362 , P3_U3259 );
nor nor_2326 ( P3_U4135 , P3_SUB_320_U51 , P3_U7363 );
nor nor_2327 ( P3_U4136 , P3_DATAWIDTH_REG_2_ , P3_DATAWIDTH_REG_3_ , P3_DATAWIDTH_REG_4_ , P3_DATAWIDTH_REG_5_ );
nor nor_2328 ( P3_U4137 , P3_DATAWIDTH_REG_6_ , P3_DATAWIDTH_REG_7_ , P3_DATAWIDTH_REG_8_ , P3_DATAWIDTH_REG_9_ );
and AND2_2329 ( P3_U4138 , P3_U4137 , P3_U4136 );
nor nor_2330 ( P3_U4139 , P3_DATAWIDTH_REG_10_ , P3_DATAWIDTH_REG_11_ , P3_DATAWIDTH_REG_12_ , P3_DATAWIDTH_REG_13_ );
nor nor_2331 ( P3_U4140 , P3_DATAWIDTH_REG_14_ , P3_DATAWIDTH_REG_15_ , P3_DATAWIDTH_REG_16_ , P3_DATAWIDTH_REG_17_ );
and AND2_2332 ( P3_U4141 , P3_U4140 , P3_U4139 );
nor nor_2333 ( P3_U4142 , P3_DATAWIDTH_REG_18_ , P3_DATAWIDTH_REG_19_ , P3_DATAWIDTH_REG_20_ , P3_DATAWIDTH_REG_21_ );
nor nor_2334 ( P3_U4143 , P3_DATAWIDTH_REG_22_ , P3_DATAWIDTH_REG_23_ , P3_DATAWIDTH_REG_24_ , P3_DATAWIDTH_REG_25_ );
and AND2_2335 ( P3_U4144 , P3_U4143 , P3_U4142 );
nor nor_2336 ( P3_U4145 , P3_DATAWIDTH_REG_26_ , P3_DATAWIDTH_REG_27_ );
nor nor_2337 ( P3_U4146 , P3_DATAWIDTH_REG_28_ , P3_DATAWIDTH_REG_29_ );
nor nor_2338 ( P3_U4147 , P3_DATAWIDTH_REG_30_ , P3_DATAWIDTH_REG_31_ );
and AND4_2339 ( P3_U4148 , P3_U4147 , P3_U7366 , P3_U4146 , P3_U4145 );
nor nor_2340 ( P3_U4149 , P3_REIP_REG_0_ , P3_DATAWIDTH_REG_0_ , P3_DATAWIDTH_REG_1_ );
and AND2_2341 ( P3_U4150 , P3_U7375 , P3_U2630 );
and AND2_2342 ( P3_U4151 , P3_U7373 , P3_U3135 );
and AND4_2343 ( P3_U4152 , P3_U7390 , P3_U7389 , P3_U7388 , P3_U7387 );
and AND4_2344 ( P3_U4153 , P3_U7394 , P3_U7393 , P3_U7392 , P3_U7391 );
and AND4_2345 ( P3_U4154 , P3_U7398 , P3_U7397 , P3_U7396 , P3_U7395 );
and AND4_2346 ( P3_U4155 , P3_U7402 , P3_U7401 , P3_U7400 , P3_U7399 );
and AND4_2347 ( P3_U4156 , P3_U7406 , P3_U7405 , P3_U7404 , P3_U7403 );
and AND4_2348 ( P3_U4157 , P3_U7410 , P3_U7409 , P3_U7408 , P3_U7407 );
and AND4_2349 ( P3_U4158 , P3_U7414 , P3_U7413 , P3_U7412 , P3_U7411 );
and AND4_2350 ( P3_U4159 , P3_U7418 , P3_U7417 , P3_U7416 , P3_U7415 );
and AND4_2351 ( P3_U4160 , P3_U7422 , P3_U7421 , P3_U7420 , P3_U7419 );
and AND4_2352 ( P3_U4161 , P3_U7426 , P3_U7425 , P3_U7424 , P3_U7423 );
and AND4_2353 ( P3_U4162 , P3_U7430 , P3_U7429 , P3_U7428 , P3_U7427 );
and AND4_2354 ( P3_U4163 , P3_U7434 , P3_U7433 , P3_U7432 , P3_U7431 );
and AND4_2355 ( P3_U4164 , P3_U7438 , P3_U7437 , P3_U7436 , P3_U7435 );
and AND4_2356 ( P3_U4165 , P3_U7442 , P3_U7441 , P3_U7440 , P3_U7439 );
and AND4_2357 ( P3_U4166 , P3_U7446 , P3_U7445 , P3_U7444 , P3_U7443 );
and AND4_2358 ( P3_U4167 , P3_U7450 , P3_U7449 , P3_U7448 , P3_U7447 );
and AND4_2359 ( P3_U4168 , P3_U7454 , P3_U7453 , P3_U7452 , P3_U7451 );
and AND4_2360 ( P3_U4169 , P3_U7458 , P3_U7457 , P3_U7456 , P3_U7455 );
and AND4_2361 ( P3_U4170 , P3_U7462 , P3_U7461 , P3_U7460 , P3_U7459 );
and AND4_2362 ( P3_U4171 , P3_U7466 , P3_U7465 , P3_U7464 , P3_U7463 );
and AND4_2363 ( P3_U4172 , P3_U7470 , P3_U7469 , P3_U7468 , P3_U7467 );
and AND4_2364 ( P3_U4173 , P3_U7474 , P3_U7473 , P3_U7472 , P3_U7471 );
and AND4_2365 ( P3_U4174 , P3_U7478 , P3_U7477 , P3_U7476 , P3_U7475 );
and AND4_2366 ( P3_U4175 , P3_U7482 , P3_U7481 , P3_U7480 , P3_U7479 );
and AND4_2367 ( P3_U4176 , P3_U7486 , P3_U7485 , P3_U7484 , P3_U7483 );
and AND4_2368 ( P3_U4177 , P3_U7490 , P3_U7489 , P3_U7488 , P3_U7487 );
and AND4_2369 ( P3_U4178 , P3_U7494 , P3_U7493 , P3_U7492 , P3_U7491 );
and AND4_2370 ( P3_U4179 , P3_U7498 , P3_U7497 , P3_U7496 , P3_U7495 );
and AND4_2371 ( P3_U4180 , P3_U7502 , P3_U7501 , P3_U7500 , P3_U7499 );
and AND4_2372 ( P3_U4181 , P3_U7506 , P3_U7505 , P3_U7504 , P3_U7503 );
and AND4_2373 ( P3_U4182 , P3_U7510 , P3_U7509 , P3_U7508 , P3_U7507 );
and AND4_2374 ( P3_U4183 , P3_U7514 , P3_U7513 , P3_U7512 , P3_U7511 );
and AND4_2375 ( P3_U4184 , P3_U7520 , P3_U7519 , P3_U7518 , P3_U7517 );
and AND4_2376 ( P3_U4185 , P3_U7524 , P3_U7523 , P3_U7522 , P3_U7521 );
and AND4_2377 ( P3_U4186 , P3_U7528 , P3_U7527 , P3_U7526 , P3_U7525 );
and AND4_2378 ( P3_U4187 , P3_U7532 , P3_U7531 , P3_U7530 , P3_U7529 );
and AND4_2379 ( P3_U4188 , P3_U7536 , P3_U7535 , P3_U7534 , P3_U7533 );
and AND4_2380 ( P3_U4189 , P3_U7540 , P3_U7539 , P3_U7538 , P3_U7537 );
and AND4_2381 ( P3_U4190 , P3_U7544 , P3_U7543 , P3_U7542 , P3_U7541 );
and AND4_2382 ( P3_U4191 , P3_U7548 , P3_U7547 , P3_U7546 , P3_U7545 );
and AND4_2383 ( P3_U4192 , P3_U7552 , P3_U7551 , P3_U7550 , P3_U7549 );
and AND4_2384 ( P3_U4193 , P3_U7556 , P3_U7555 , P3_U7554 , P3_U7553 );
and AND4_2385 ( P3_U4194 , P3_U7560 , P3_U7559 , P3_U7558 , P3_U7557 );
and AND4_2386 ( P3_U4195 , P3_U7564 , P3_U7563 , P3_U7562 , P3_U7561 );
and AND4_2387 ( P3_U4196 , P3_U7568 , P3_U7567 , P3_U7566 , P3_U7565 );
and AND4_2388 ( P3_U4197 , P3_U7572 , P3_U7571 , P3_U7570 , P3_U7569 );
and AND4_2389 ( P3_U4198 , P3_U7576 , P3_U7575 , P3_U7574 , P3_U7573 );
and AND4_2390 ( P3_U4199 , P3_U7580 , P3_U7579 , P3_U7578 , P3_U7577 );
and AND4_2391 ( P3_U4200 , P3_U7584 , P3_U7583 , P3_U7582 , P3_U7581 );
and AND4_2392 ( P3_U4201 , P3_U7588 , P3_U7587 , P3_U7586 , P3_U7585 );
and AND4_2393 ( P3_U4202 , P3_U7592 , P3_U7591 , P3_U7590 , P3_U7589 );
and AND4_2394 ( P3_U4203 , P3_U7596 , P3_U7595 , P3_U7594 , P3_U7593 );
and AND4_2395 ( P3_U4204 , P3_U7600 , P3_U7599 , P3_U7598 , P3_U7597 );
and AND4_2396 ( P3_U4205 , P3_U7604 , P3_U7603 , P3_U7602 , P3_U7601 );
and AND4_2397 ( P3_U4206 , P3_U7608 , P3_U7607 , P3_U7606 , P3_U7605 );
and AND4_2398 ( P3_U4207 , P3_U7612 , P3_U7611 , P3_U7610 , P3_U7609 );
and AND4_2399 ( P3_U4208 , P3_U7616 , P3_U7615 , P3_U7614 , P3_U7613 );
and AND4_2400 ( P3_U4209 , P3_U7620 , P3_U7619 , P3_U7618 , P3_U7617 );
and AND4_2401 ( P3_U4210 , P3_U7624 , P3_U7623 , P3_U7622 , P3_U7621 );
and AND4_2402 ( P3_U4211 , P3_U7628 , P3_U7627 , P3_U7626 , P3_U7625 );
and AND4_2403 ( P3_U4212 , P3_U7632 , P3_U7631 , P3_U7630 , P3_U7629 );
and AND4_2404 ( P3_U4213 , P3_U7636 , P3_U7635 , P3_U7634 , P3_U7633 );
and AND4_2405 ( P3_U4214 , P3_U7640 , P3_U7639 , P3_U7638 , P3_U7637 );
and AND4_2406 ( P3_U4215 , P3_U7644 , P3_U7643 , P3_U7642 , P3_U7641 );
and AND4_2407 ( P3_U4216 , P3_U7649 , P3_U7648 , P3_U7647 , P3_U7646 );
and AND4_2408 ( P3_U4217 , P3_U7653 , P3_U7652 , P3_U7651 , P3_U7650 );
and AND4_2409 ( P3_U4218 , P3_U7657 , P3_U7656 , P3_U7655 , P3_U7654 );
and AND4_2410 ( P3_U4219 , P3_U7661 , P3_U7660 , P3_U7659 , P3_U7658 );
and AND4_2411 ( P3_U4220 , P3_U7665 , P3_U7664 , P3_U7663 , P3_U7662 );
and AND4_2412 ( P3_U4221 , P3_U7669 , P3_U7668 , P3_U7667 , P3_U7666 );
and AND4_2413 ( P3_U4222 , P3_U7673 , P3_U7672 , P3_U7671 , P3_U7670 );
and AND4_2414 ( P3_U4223 , P3_U7677 , P3_U7676 , P3_U7675 , P3_U7674 );
and AND4_2415 ( P3_U4224 , P3_U7681 , P3_U7680 , P3_U7679 , P3_U7678 );
and AND4_2416 ( P3_U4225 , P3_U7685 , P3_U7684 , P3_U7683 , P3_U7682 );
and AND4_2417 ( P3_U4226 , P3_U7689 , P3_U7688 , P3_U7687 , P3_U7686 );
and AND4_2418 ( P3_U4227 , P3_U7693 , P3_U7692 , P3_U7691 , P3_U7690 );
and AND4_2419 ( P3_U4228 , P3_U7697 , P3_U7696 , P3_U7695 , P3_U7694 );
and AND4_2420 ( P3_U4229 , P3_U7701 , P3_U7700 , P3_U7699 , P3_U7698 );
and AND4_2421 ( P3_U4230 , P3_U7705 , P3_U7704 , P3_U7703 , P3_U7702 );
and AND4_2422 ( P3_U4231 , P3_U7709 , P3_U7708 , P3_U7707 , P3_U7706 );
and AND4_2423 ( P3_U4232 , P3_U7713 , P3_U7712 , P3_U7711 , P3_U7710 );
and AND4_2424 ( P3_U4233 , P3_U7717 , P3_U7716 , P3_U7715 , P3_U7714 );
and AND4_2425 ( P3_U4234 , P3_U7721 , P3_U7720 , P3_U7719 , P3_U7718 );
and AND4_2426 ( P3_U4235 , P3_U7725 , P3_U7724 , P3_U7723 , P3_U7722 );
and AND4_2427 ( P3_U4236 , P3_U7729 , P3_U7728 , P3_U7727 , P3_U7726 );
and AND4_2428 ( P3_U4237 , P3_U7733 , P3_U7732 , P3_U7731 , P3_U7730 );
and AND4_2429 ( P3_U4238 , P3_U7737 , P3_U7736 , P3_U7735 , P3_U7734 );
and AND4_2430 ( P3_U4239 , P3_U7741 , P3_U7740 , P3_U7739 , P3_U7738 );
and AND4_2431 ( P3_U4240 , P3_U7745 , P3_U7744 , P3_U7743 , P3_U7742 );
and AND4_2432 ( P3_U4241 , P3_U7749 , P3_U7748 , P3_U7747 , P3_U7746 );
and AND4_2433 ( P3_U4242 , P3_U7753 , P3_U7752 , P3_U7751 , P3_U7750 );
and AND4_2434 ( P3_U4243 , P3_U7757 , P3_U7756 , P3_U7755 , P3_U7754 );
and AND4_2435 ( P3_U4244 , P3_U7761 , P3_U7760 , P3_U7759 , P3_U7758 );
and AND4_2436 ( P3_U4245 , P3_U7765 , P3_U7764 , P3_U7763 , P3_U7762 );
and AND4_2437 ( P3_U4246 , P3_U7769 , P3_U7768 , P3_U7767 , P3_U7766 );
and AND4_2438 ( P3_U4247 , P3_U7773 , P3_U7772 , P3_U7771 , P3_U7770 );
and AND4_2439 ( P3_U4248 , P3_U7779 , P3_U7778 , P3_U7777 , P3_U7776 );
and AND4_2440 ( P3_U4249 , P3_U7783 , P3_U7782 , P3_U7781 , P3_U7780 );
and AND4_2441 ( P3_U4250 , P3_U7787 , P3_U7786 , P3_U7785 , P3_U7784 );
and AND4_2442 ( P3_U4251 , P3_U7791 , P3_U7790 , P3_U7789 , P3_U7788 );
and AND4_2443 ( P3_U4252 , P3_U7795 , P3_U7794 , P3_U7793 , P3_U7792 );
and AND4_2444 ( P3_U4253 , P3_U7799 , P3_U7798 , P3_U7797 , P3_U7796 );
and AND4_2445 ( P3_U4254 , P3_U7803 , P3_U7802 , P3_U7801 , P3_U7800 );
and AND4_2446 ( P3_U4255 , P3_U7807 , P3_U7806 , P3_U7805 , P3_U7804 );
and AND4_2447 ( P3_U4256 , P3_U7811 , P3_U7810 , P3_U7809 , P3_U7808 );
and AND4_2448 ( P3_U4257 , P3_U7815 , P3_U7814 , P3_U7813 , P3_U7812 );
and AND4_2449 ( P3_U4258 , P3_U7819 , P3_U7818 , P3_U7817 , P3_U7816 );
and AND4_2450 ( P3_U4259 , P3_U7823 , P3_U7822 , P3_U7821 , P3_U7820 );
and AND4_2451 ( P3_U4260 , P3_U7827 , P3_U7826 , P3_U7825 , P3_U7824 );
and AND4_2452 ( P3_U4261 , P3_U7831 , P3_U7830 , P3_U7829 , P3_U7828 );
and AND4_2453 ( P3_U4262 , P3_U7835 , P3_U7834 , P3_U7833 , P3_U7832 );
and AND4_2454 ( P3_U4263 , P3_U7839 , P3_U7838 , P3_U7837 , P3_U7836 );
and AND4_2455 ( P3_U4264 , P3_U7843 , P3_U7842 , P3_U7841 , P3_U7840 );
and AND4_2456 ( P3_U4265 , P3_U7847 , P3_U7846 , P3_U7845 , P3_U7844 );
and AND4_2457 ( P3_U4266 , P3_U7851 , P3_U7850 , P3_U7849 , P3_U7848 );
and AND4_2458 ( P3_U4267 , P3_U7855 , P3_U7854 , P3_U7853 , P3_U7852 );
and AND4_2459 ( P3_U4268 , P3_U7859 , P3_U7858 , P3_U7857 , P3_U7856 );
and AND4_2460 ( P3_U4269 , P3_U7863 , P3_U7862 , P3_U7861 , P3_U7860 );
and AND4_2461 ( P3_U4270 , P3_U7867 , P3_U7866 , P3_U7865 , P3_U7864 );
and AND4_2462 ( P3_U4271 , P3_U7871 , P3_U7870 , P3_U7869 , P3_U7868 );
and AND4_2463 ( P3_U4272 , P3_U7875 , P3_U7874 , P3_U7873 , P3_U7872 );
and AND4_2464 ( P3_U4273 , P3_U7879 , P3_U7878 , P3_U7877 , P3_U7876 );
and AND4_2465 ( P3_U4274 , P3_U7883 , P3_U7882 , P3_U7881 , P3_U7880 );
and AND4_2466 ( P3_U4275 , P3_U7887 , P3_U7886 , P3_U7885 , P3_U7884 );
and AND4_2467 ( P3_U4276 , P3_U7891 , P3_U7890 , P3_U7889 , P3_U7888 );
and AND4_2468 ( P3_U4277 , P3_U7895 , P3_U7894 , P3_U7893 , P3_U7892 );
and AND4_2469 ( P3_U4278 , P3_U7899 , P3_U7898 , P3_U7897 , P3_U7896 );
and AND4_2470 ( P3_U4279 , P3_U7903 , P3_U7902 , P3_U7901 , P3_U7900 );
and AND2_2471 ( P3_U4280 , P3_U7943 , P3_U7942 );
nand NAND2_2472 ( P3_U4281 , P3_U3361 , P3_U2604 );
and AND2_2473 ( P3_U4282 , P3_U7951 , P3_U7950 );
nand NAND2_2474 ( P3_U4283 , P3_U3658 , P3_U5497 );
not NOT1_2475 ( P3_U4284 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_2476 ( P3_U4285 , P3_U2390 , P3_U4281 );
not NOT1_2477 ( P3_U4286 , BS16 );
nand NAND2_2478 ( P3_U4287 , P3_U4151 , P3_U4334 );
nand NAND2_2479 ( P3_U4288 , P3_U4334 , P3_U3239 );
nand NAND2_2480 ( P3_U4289 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_U3091 );
nand NAND3_2481 ( P3_U4290 , P3_U2515 , P3_U2516 , P3_U3657 );
not NOT1_2482 ( P3_U4291 , P3_U3267 );
nand NAND2_2483 ( P3_U4292 , HOLD , P3_U2630 );
not NOT1_2484 ( P3_U4293 , P3_U3105 );
not NOT1_2485 ( P3_U4294 , P3_U3106 );
not NOT1_2486 ( P3_U4295 , P3_U3135 );
not NOT1_2487 ( P3_U4296 , P3_U3112 );
not NOT1_2488 ( P3_U4297 , P3_U3111 );
not NOT1_2489 ( P3_U4298 , P3_U3242 );
not NOT1_2490 ( P3_U4299 , P3_U3243 );
not NOT1_2491 ( P3_U4300 , P3_U3244 );
not NOT1_2492 ( P3_U4301 , P3_U3245 );
not NOT1_2493 ( P3_U4302 , P3_U3119 );
not NOT1_2494 ( P3_U4303 , P3_U3117 );
not NOT1_2495 ( P3_U4304 , P3_U3116 );
not NOT1_2496 ( P3_U4305 , P3_U3115 );
not NOT1_2497 ( P3_U4306 , P3_U3246 );
not NOT1_2498 ( P3_U4307 , P3_U3261 );
not NOT1_2499 ( P3_U4308 , P3_U3077 );
not NOT1_2500 ( P3_U4309 , P3_U3253 );
not NOT1_2501 ( P3_U4310 , P3_U3252 );
not NOT1_2502 ( P3_U4311 , P3_U3250 );
not NOT1_2503 ( P3_U4312 , P3_U3127 );
not NOT1_2504 ( P3_U4313 , P3_LT_563_1260_U6 );
not NOT1_2505 ( P3_U4314 , P3_U3217 );
nand NAND2_2506 ( P3_U4315 , P3_U4295 , P3_U2631 );
nand NAND2_2507 ( P3_U4316 , P3_U4347 , P3_U3260 );
nand NAND2_2508 ( P3_U4317 , P3_U2383 , P3_U3105 );
not NOT1_2509 ( P3_U4318 , P3_U3247 );
not NOT1_2510 ( P3_U4319 , P3_U3259 );
not NOT1_2511 ( P3_U4320 , P3_U3080 );
not NOT1_2512 ( P3_U4321 , P3_U3078 );
not NOT1_2513 ( P3_U4322 , P3_U3136 );
not NOT1_2514 ( P3_U4323 , P3_U3114 );
not NOT1_2515 ( P3_U4324 , P3_U3118 );
not NOT1_2516 ( P3_U4325 , P3_U3219 );
not NOT1_2517 ( P3_U4326 , P3_U3181 );
nand NAND2_2518 ( P3_U4327 , P3_U4149 , P3_U4307 );
nand NAND2_2519 ( P3_U4328 , P3_U3365 , P3_U4354 );
nand NAND4_2520 ( P3_U4329 , P3_STATE2_REG_1_ , P3_U3121 , P3_U3090 , P3_U2631 );
nand NAND2_2521 ( P3_U4330 , P3_U3653 , P3_U2453 );
nand NAND2_2522 ( P3_U4331 , P3_U2458 , P3_U4653 );
not NOT1_2523 ( P3_U4332 , P3_U3095 );
nand NAND2_2524 ( P3_U4333 , P3_U4350 , P3_U3113 );
nand NAND2_2525 ( P3_U4334 , P3_U2390 , P3_U7093 );
nand NAND2_2526 ( P3_U4335 , P3_U4452 , P3_U3085 );
nand NAND2_2527 ( P3_U4336 , P3_U4347 , P3_U3121 );
nand NAND2_2528 ( P3_U4337 , P3_U2453 , P3_U3232 );
nand NAND3_2529 ( P3_U4338 , P3_U3090 , P3_STATE2_REG_0_ , U209 );
nand NAND2_2530 ( P3_U4339 , P3_U3654 , P3_U4608 );
not NOT1_2531 ( P3_U4340 , P3_U3123 );
not NOT1_2532 ( P3_U4341 , P3_U3229 );
not NOT1_2533 ( P3_U4342 , P3_U3150 );
not NOT1_2534 ( P3_U4343 , P3_U3158 );
not NOT1_2535 ( P3_U4344 , P3_U3103 );
not NOT1_2536 ( P3_U4345 , P3_U3126 );
not NOT1_2537 ( P3_U4346 , P3_U3082 );
not NOT1_2538 ( P3_U4347 , P3_U3239 );
not NOT1_2539 ( P3_U4348 , P3_U3236 );
not NOT1_2540 ( P3_U4349 , P3_U3235 );
not NOT1_2541 ( P3_U4350 , P3_U3208 );
not NOT1_2542 ( P3_U4351 , P3_U3216 );
not NOT1_2543 ( P3_U4352 , P3_U3222 );
not NOT1_2544 ( P3_U4353 , P3_U3124 );
not NOT1_2545 ( P3_U4354 , P3_U3125 );
nand NAND2_2546 ( P3_U4355 , P3_REIP_REG_31_ , P3_U4321 );
nand NAND2_2547 ( P3_U4356 , P3_REIP_REG_30_ , P3_U4320 );
nand NAND2_2548 ( P3_U4357 , P3_ADDRESS_REG_29_ , P3_U3077 );
nand NAND2_2549 ( P3_U4358 , P3_REIP_REG_30_ , P3_U4321 );
nand NAND2_2550 ( P3_U4359 , P3_REIP_REG_29_ , P3_U4320 );
nand NAND2_2551 ( P3_U4360 , P3_ADDRESS_REG_28_ , P3_U3077 );
nand NAND2_2552 ( P3_U4361 , P3_REIP_REG_29_ , P3_U4321 );
nand NAND2_2553 ( P3_U4362 , P3_REIP_REG_28_ , P3_U4320 );
nand NAND2_2554 ( P3_U4363 , P3_ADDRESS_REG_27_ , P3_U3077 );
nand NAND2_2555 ( P3_U4364 , P3_REIP_REG_28_ , P3_U4321 );
nand NAND2_2556 ( P3_U4365 , P3_REIP_REG_27_ , P3_U4320 );
nand NAND2_2557 ( P3_U4366 , P3_ADDRESS_REG_26_ , P3_U3077 );
nand NAND2_2558 ( P3_U4367 , P3_REIP_REG_27_ , P3_U4321 );
nand NAND2_2559 ( P3_U4368 , P3_REIP_REG_26_ , P3_U4320 );
nand NAND2_2560 ( P3_U4369 , P3_ADDRESS_REG_25_ , P3_U3077 );
nand NAND2_2561 ( P3_U4370 , P3_REIP_REG_26_ , P3_U4321 );
nand NAND2_2562 ( P3_U4371 , P3_REIP_REG_25_ , P3_U4320 );
nand NAND2_2563 ( P3_U4372 , P3_ADDRESS_REG_24_ , P3_U3077 );
nand NAND2_2564 ( P3_U4373 , P3_REIP_REG_25_ , P3_U4321 );
nand NAND2_2565 ( P3_U4374 , P3_REIP_REG_24_ , P3_U4320 );
nand NAND2_2566 ( P3_U4375 , P3_ADDRESS_REG_23_ , P3_U3077 );
nand NAND2_2567 ( P3_U4376 , P3_REIP_REG_24_ , P3_U4321 );
nand NAND2_2568 ( P3_U4377 , P3_REIP_REG_23_ , P3_U4320 );
nand NAND2_2569 ( P3_U4378 , P3_ADDRESS_REG_22_ , P3_U3077 );
nand NAND2_2570 ( P3_U4379 , P3_REIP_REG_23_ , P3_U4321 );
nand NAND2_2571 ( P3_U4380 , P3_REIP_REG_22_ , P3_U4320 );
nand NAND2_2572 ( P3_U4381 , P3_ADDRESS_REG_21_ , P3_U3077 );
nand NAND2_2573 ( P3_U4382 , P3_REIP_REG_22_ , P3_U4321 );
nand NAND2_2574 ( P3_U4383 , P3_REIP_REG_21_ , P3_U4320 );
nand NAND2_2575 ( P3_U4384 , P3_ADDRESS_REG_20_ , P3_U3077 );
nand NAND2_2576 ( P3_U4385 , P3_REIP_REG_21_ , P3_U4321 );
nand NAND2_2577 ( P3_U4386 , P3_REIP_REG_20_ , P3_U4320 );
nand NAND2_2578 ( P3_U4387 , P3_ADDRESS_REG_19_ , P3_U3077 );
nand NAND2_2579 ( P3_U4388 , P3_REIP_REG_20_ , P3_U4321 );
nand NAND2_2580 ( P3_U4389 , P3_REIP_REG_19_ , P3_U4320 );
nand NAND2_2581 ( P3_U4390 , P3_ADDRESS_REG_18_ , P3_U3077 );
nand NAND2_2582 ( P3_U4391 , P3_REIP_REG_19_ , P3_U4321 );
nand NAND2_2583 ( P3_U4392 , P3_REIP_REG_18_ , P3_U4320 );
nand NAND2_2584 ( P3_U4393 , P3_ADDRESS_REG_17_ , P3_U3077 );
nand NAND2_2585 ( P3_U4394 , P3_REIP_REG_18_ , P3_U4321 );
nand NAND2_2586 ( P3_U4395 , P3_REIP_REG_17_ , P3_U4320 );
nand NAND2_2587 ( P3_U4396 , P3_ADDRESS_REG_16_ , P3_U3077 );
nand NAND2_2588 ( P3_U4397 , P3_REIP_REG_17_ , P3_U4321 );
nand NAND2_2589 ( P3_U4398 , P3_REIP_REG_16_ , P3_U4320 );
nand NAND2_2590 ( P3_U4399 , P3_ADDRESS_REG_15_ , P3_U3077 );
nand NAND2_2591 ( P3_U4400 , P3_REIP_REG_16_ , P3_U4321 );
nand NAND2_2592 ( P3_U4401 , P3_REIP_REG_15_ , P3_U4320 );
nand NAND2_2593 ( P3_U4402 , P3_ADDRESS_REG_14_ , P3_U3077 );
nand NAND2_2594 ( P3_U4403 , P3_REIP_REG_15_ , P3_U4321 );
nand NAND2_2595 ( P3_U4404 , P3_REIP_REG_14_ , P3_U4320 );
nand NAND2_2596 ( P3_U4405 , P3_ADDRESS_REG_13_ , P3_U3077 );
nand NAND2_2597 ( P3_U4406 , P3_REIP_REG_14_ , P3_U4321 );
nand NAND2_2598 ( P3_U4407 , P3_REIP_REG_13_ , P3_U4320 );
nand NAND2_2599 ( P3_U4408 , P3_ADDRESS_REG_12_ , P3_U3077 );
nand NAND2_2600 ( P3_U4409 , P3_REIP_REG_13_ , P3_U4321 );
nand NAND2_2601 ( P3_U4410 , P3_REIP_REG_12_ , P3_U4320 );
nand NAND2_2602 ( P3_U4411 , P3_ADDRESS_REG_11_ , P3_U3077 );
nand NAND2_2603 ( P3_U4412 , P3_REIP_REG_12_ , P3_U4321 );
nand NAND2_2604 ( P3_U4413 , P3_REIP_REG_11_ , P3_U4320 );
nand NAND2_2605 ( P3_U4414 , P3_ADDRESS_REG_10_ , P3_U3077 );
nand NAND2_2606 ( P3_U4415 , P3_REIP_REG_11_ , P3_U4321 );
nand NAND2_2607 ( P3_U4416 , P3_REIP_REG_10_ , P3_U4320 );
nand NAND2_2608 ( P3_U4417 , P3_ADDRESS_REG_9_ , P3_U3077 );
nand NAND2_2609 ( P3_U4418 , P3_REIP_REG_10_ , P3_U4321 );
nand NAND2_2610 ( P3_U4419 , P3_REIP_REG_9_ , P3_U4320 );
nand NAND2_2611 ( P3_U4420 , P3_ADDRESS_REG_8_ , P3_U3077 );
nand NAND2_2612 ( P3_U4421 , P3_REIP_REG_9_ , P3_U4321 );
nand NAND2_2613 ( P3_U4422 , P3_REIP_REG_8_ , P3_U4320 );
nand NAND2_2614 ( P3_U4423 , P3_ADDRESS_REG_7_ , P3_U3077 );
nand NAND2_2615 ( P3_U4424 , P3_REIP_REG_8_ , P3_U4321 );
nand NAND2_2616 ( P3_U4425 , P3_REIP_REG_7_ , P3_U4320 );
nand NAND2_2617 ( P3_U4426 , P3_ADDRESS_REG_6_ , P3_U3077 );
nand NAND2_2618 ( P3_U4427 , P3_REIP_REG_7_ , P3_U4321 );
nand NAND2_2619 ( P3_U4428 , P3_REIP_REG_6_ , P3_U4320 );
nand NAND2_2620 ( P3_U4429 , P3_ADDRESS_REG_5_ , P3_U3077 );
nand NAND2_2621 ( P3_U4430 , P3_REIP_REG_6_ , P3_U4321 );
nand NAND2_2622 ( P3_U4431 , P3_REIP_REG_5_ , P3_U4320 );
nand NAND2_2623 ( P3_U4432 , P3_ADDRESS_REG_4_ , P3_U3077 );
nand NAND2_2624 ( P3_U4433 , P3_REIP_REG_5_ , P3_U4321 );
nand NAND2_2625 ( P3_U4434 , P3_REIP_REG_4_ , P3_U4320 );
nand NAND2_2626 ( P3_U4435 , P3_ADDRESS_REG_3_ , P3_U3077 );
nand NAND2_2627 ( P3_U4436 , P3_REIP_REG_4_ , P3_U4321 );
nand NAND2_2628 ( P3_U4437 , P3_REIP_REG_3_ , P3_U4320 );
nand NAND2_2629 ( P3_U4438 , P3_ADDRESS_REG_2_ , P3_U3077 );
nand NAND2_2630 ( P3_U4439 , P3_REIP_REG_3_ , P3_U4321 );
nand NAND2_2631 ( P3_U4440 , P3_REIP_REG_2_ , P3_U4320 );
nand NAND2_2632 ( P3_U4441 , P3_ADDRESS_REG_1_ , P3_U3077 );
nand NAND2_2633 ( P3_U4442 , P3_REIP_REG_2_ , P3_U4321 );
nand NAND2_2634 ( P3_U4443 , P3_REIP_REG_1_ , P3_U4320 );
nand NAND2_2635 ( P3_U4444 , P3_ADDRESS_REG_0_ , P3_U3077 );
not NOT1_2636 ( P3_U4445 , P3_U3087 );
nand NAND2_2637 ( P3_U4446 , P3_U4445 , P3_U2630 );
nand NAND2_2638 ( P3_U4447 , NA , P3_U4346 );
not NOT1_2639 ( P3_U4448 , P3_U3088 );
nand NAND2_2640 ( P3_U4449 , P3_U4448 , P3_U2630 );
or OR2_2641 ( P3_U4450 , P3_STATE_REG_0_ , NA );
nand NAND3_2642 ( P3_U4451 , P3_U7912 , P3_U4450 , P3_U7913 );
not NOT1_2643 ( P3_U4452 , P3_U3083 );
nand NAND3_2644 ( P3_U4453 , P3_U3088 , U209 , P3_U4346 );
nand NAND3_2645 ( P3_U4454 , HOLD , P3_U3075 , P3_U4452 );
nand NAND2_2646 ( P3_U4455 , P3_U4453 , P3_U4454 );
nand NAND2_2647 ( P3_U4456 , P3_U3309 , P3_U4455 );
nand NAND2_2648 ( P3_U4457 , P3_STATE_REG_2_ , P3_U4451 );
nand NAND2_2649 ( P3_U4458 , P3_U4308 , U209 );
nand NAND2_2650 ( P3_U4459 , P3_U3312 , P3_U7915 );
nand NAND2_2651 ( P3_U4460 , P3_STATE_REG_2_ , P3_U3087 );
nand NAND2_2652 ( P3_U4461 , NA , P3_U3085 );
nand NAND2_2653 ( P3_U4462 , P3_U4461 , P3_U4460 );
nand NAND2_2654 ( P3_U4463 , P3_U4462 , P3_U3076 );
nand NAND2_2655 ( P3_U4464 , P3_U4286 , P3_U3083 );
nand NAND2_2656 ( P3_U4465 , P3_STATE_REG_2_ , P3_U3076 );
nand NAND2_2657 ( P3_U4466 , P3_U3082 , P3_U4465 );
not NOT1_2658 ( P3_U4467 , P3_U3091 );
not NOT1_2659 ( P3_U4468 , P3_U3096 );
not NOT1_2660 ( P3_U4469 , P3_U3092 );
not NOT1_2661 ( P3_U4470 , P3_U3098 );
not NOT1_2662 ( P3_U4471 , P3_U3099 );
nand NAND2_2663 ( P3_U4472 , P3_INSTQUEUE_REG_0__0_ , P3_U2484 );
nand NAND2_2664 ( P3_U4473 , P3_INSTQUEUE_REG_1__0_ , P3_U2483 );
nand NAND2_2665 ( P3_U4474 , P3_INSTQUEUE_REG_2__0_ , P3_U2482 );
nand NAND2_2666 ( P3_U4475 , P3_INSTQUEUE_REG_3__0_ , P3_U2480 );
nand NAND2_2667 ( P3_U4476 , P3_INSTQUEUE_REG_4__0_ , P3_U2479 );
nand NAND2_2668 ( P3_U4477 , P3_INSTQUEUE_REG_5__0_ , P3_U2478 );
nand NAND2_2669 ( P3_U4478 , P3_INSTQUEUE_REG_6__0_ , P3_U2477 );
nand NAND2_2670 ( P3_U4479 , P3_INSTQUEUE_REG_7__0_ , P3_U4471 );
nand NAND2_2671 ( P3_U4480 , P3_INSTQUEUE_REG_8__0_ , P3_U2476 );
nand NAND2_2672 ( P3_U4481 , P3_INSTQUEUE_REG_9__0_ , P3_U2475 );
nand NAND2_2673 ( P3_U4482 , P3_INSTQUEUE_REG_10__0_ , P3_U2473 );
nand NAND2_2674 ( P3_U4483 , P3_INSTQUEUE_REG_11__0_ , P3_U2471 );
nand NAND2_2675 ( P3_U4484 , P3_INSTQUEUE_REG_12__0_ , P3_U2470 );
nand NAND2_2676 ( P3_U4485 , P3_INSTQUEUE_REG_13__0_ , P3_U2469 );
nand NAND2_2677 ( P3_U4486 , P3_INSTQUEUE_REG_14__0_ , P3_U2467 );
nand NAND2_2678 ( P3_U4487 , P3_INSTQUEUE_REG_15__0_ , P3_U2465 );
not NOT1_2679 ( P3_U4488 , P3_U3108 );
nand NAND2_2680 ( P3_U4489 , P3_INSTQUEUE_REG_0__1_ , P3_U2484 );
nand NAND2_2681 ( P3_U4490 , P3_INSTQUEUE_REG_1__1_ , P3_U2483 );
nand NAND2_2682 ( P3_U4491 , P3_INSTQUEUE_REG_2__1_ , P3_U2482 );
nand NAND2_2683 ( P3_U4492 , P3_INSTQUEUE_REG_3__1_ , P3_U2480 );
nand NAND2_2684 ( P3_U4493 , P3_INSTQUEUE_REG_4__1_ , P3_U2479 );
nand NAND2_2685 ( P3_U4494 , P3_INSTQUEUE_REG_5__1_ , P3_U2478 );
nand NAND2_2686 ( P3_U4495 , P3_INSTQUEUE_REG_6__1_ , P3_U2477 );
nand NAND2_2687 ( P3_U4496 , P3_INSTQUEUE_REG_7__1_ , P3_U4471 );
nand NAND2_2688 ( P3_U4497 , P3_INSTQUEUE_REG_8__1_ , P3_U2476 );
nand NAND2_2689 ( P3_U4498 , P3_INSTQUEUE_REG_9__1_ , P3_U2475 );
nand NAND2_2690 ( P3_U4499 , P3_INSTQUEUE_REG_10__1_ , P3_U2473 );
nand NAND2_2691 ( P3_U4500 , P3_INSTQUEUE_REG_11__1_ , P3_U2471 );
nand NAND2_2692 ( P3_U4501 , P3_INSTQUEUE_REG_12__1_ , P3_U2470 );
nand NAND2_2693 ( P3_U4502 , P3_INSTQUEUE_REG_13__1_ , P3_U2469 );
nand NAND2_2694 ( P3_U4503 , P3_INSTQUEUE_REG_14__1_ , P3_U2467 );
nand NAND2_2695 ( P3_U4504 , P3_INSTQUEUE_REG_15__1_ , P3_U2465 );
not NOT1_2696 ( P3_U4505 , P3_U3104 );
nand NAND2_2697 ( P3_U4506 , P3_INSTQUEUE_REG_0__4_ , P3_U2484 );
nand NAND2_2698 ( P3_U4507 , P3_INSTQUEUE_REG_1__4_ , P3_U2483 );
nand NAND2_2699 ( P3_U4508 , P3_INSTQUEUE_REG_2__4_ , P3_U2482 );
nand NAND2_2700 ( P3_U4509 , P3_INSTQUEUE_REG_3__4_ , P3_U2480 );
nand NAND2_2701 ( P3_U4510 , P3_INSTQUEUE_REG_4__4_ , P3_U2479 );
nand NAND2_2702 ( P3_U4511 , P3_INSTQUEUE_REG_5__4_ , P3_U2478 );
nand NAND2_2703 ( P3_U4512 , P3_INSTQUEUE_REG_6__4_ , P3_U2477 );
nand NAND2_2704 ( P3_U4513 , P3_INSTQUEUE_REG_7__4_ , P3_U4471 );
nand NAND2_2705 ( P3_U4514 , P3_INSTQUEUE_REG_8__4_ , P3_U2476 );
nand NAND2_2706 ( P3_U4515 , P3_INSTQUEUE_REG_9__4_ , P3_U2475 );
nand NAND2_2707 ( P3_U4516 , P3_INSTQUEUE_REG_10__4_ , P3_U2473 );
nand NAND2_2708 ( P3_U4517 , P3_INSTQUEUE_REG_11__4_ , P3_U2471 );
nand NAND2_2709 ( P3_U4518 , P3_INSTQUEUE_REG_12__4_ , P3_U2470 );
nand NAND2_2710 ( P3_U4519 , P3_INSTQUEUE_REG_13__4_ , P3_U2469 );
nand NAND2_2711 ( P3_U4520 , P3_INSTQUEUE_REG_14__4_ , P3_U2467 );
nand NAND2_2712 ( P3_U4521 , P3_INSTQUEUE_REG_15__4_ , P3_U2465 );
not NOT1_2713 ( P3_U4522 , P3_U3102 );
nand NAND2_2714 ( P3_U4523 , P3_INSTQUEUE_REG_0__2_ , P3_U2484 );
nand NAND2_2715 ( P3_U4524 , P3_INSTQUEUE_REG_1__2_ , P3_U2483 );
nand NAND2_2716 ( P3_U4525 , P3_INSTQUEUE_REG_2__2_ , P3_U2482 );
nand NAND2_2717 ( P3_U4526 , P3_INSTQUEUE_REG_3__2_ , P3_U2480 );
nand NAND2_2718 ( P3_U4527 , P3_INSTQUEUE_REG_4__2_ , P3_U2479 );
nand NAND2_2719 ( P3_U4528 , P3_INSTQUEUE_REG_5__2_ , P3_U2478 );
nand NAND2_2720 ( P3_U4529 , P3_INSTQUEUE_REG_6__2_ , P3_U2477 );
nand NAND2_2721 ( P3_U4530 , P3_INSTQUEUE_REG_7__2_ , P3_U4471 );
nand NAND2_2722 ( P3_U4531 , P3_INSTQUEUE_REG_8__2_ , P3_U2476 );
nand NAND2_2723 ( P3_U4532 , P3_INSTQUEUE_REG_9__2_ , P3_U2475 );
nand NAND2_2724 ( P3_U4533 , P3_INSTQUEUE_REG_10__2_ , P3_U2473 );
nand NAND2_2725 ( P3_U4534 , P3_INSTQUEUE_REG_11__2_ , P3_U2471 );
nand NAND2_2726 ( P3_U4535 , P3_INSTQUEUE_REG_12__2_ , P3_U2470 );
nand NAND2_2727 ( P3_U4536 , P3_INSTQUEUE_REG_13__2_ , P3_U2469 );
nand NAND2_2728 ( P3_U4537 , P3_INSTQUEUE_REG_14__2_ , P3_U2467 );
nand NAND2_2729 ( P3_U4538 , P3_INSTQUEUE_REG_15__2_ , P3_U2465 );
not NOT1_2730 ( P3_U4539 , P3_U3101 );
nand NAND2_2731 ( P3_U4540 , P3_INSTQUEUE_REG_0__3_ , P3_U2484 );
nand NAND2_2732 ( P3_U4541 , P3_INSTQUEUE_REG_1__3_ , P3_U2483 );
nand NAND2_2733 ( P3_U4542 , P3_INSTQUEUE_REG_2__3_ , P3_U2482 );
nand NAND2_2734 ( P3_U4543 , P3_INSTQUEUE_REG_3__3_ , P3_U2480 );
nand NAND2_2735 ( P3_U4544 , P3_INSTQUEUE_REG_4__3_ , P3_U2479 );
nand NAND2_2736 ( P3_U4545 , P3_INSTQUEUE_REG_5__3_ , P3_U2478 );
nand NAND2_2737 ( P3_U4546 , P3_INSTQUEUE_REG_6__3_ , P3_U2477 );
nand NAND2_2738 ( P3_U4547 , P3_INSTQUEUE_REG_7__3_ , P3_U4471 );
nand NAND2_2739 ( P3_U4548 , P3_INSTQUEUE_REG_8__3_ , P3_U2476 );
nand NAND2_2740 ( P3_U4549 , P3_INSTQUEUE_REG_9__3_ , P3_U2475 );
nand NAND2_2741 ( P3_U4550 , P3_INSTQUEUE_REG_10__3_ , P3_U2473 );
nand NAND2_2742 ( P3_U4551 , P3_INSTQUEUE_REG_11__3_ , P3_U2471 );
nand NAND2_2743 ( P3_U4552 , P3_INSTQUEUE_REG_12__3_ , P3_U2470 );
nand NAND2_2744 ( P3_U4553 , P3_INSTQUEUE_REG_13__3_ , P3_U2469 );
nand NAND2_2745 ( P3_U4554 , P3_INSTQUEUE_REG_14__3_ , P3_U2467 );
nand NAND2_2746 ( P3_U4555 , P3_INSTQUEUE_REG_15__3_ , P3_U2465 );
not NOT1_2747 ( P3_U4556 , P3_U3107 );
nand NAND2_2748 ( P3_U4557 , P3_INSTQUEUE_REG_0__7_ , P3_U2484 );
nand NAND2_2749 ( P3_U4558 , P3_INSTQUEUE_REG_1__7_ , P3_U2483 );
nand NAND2_2750 ( P3_U4559 , P3_INSTQUEUE_REG_2__7_ , P3_U2482 );
nand NAND2_2751 ( P3_U4560 , P3_INSTQUEUE_REG_3__7_ , P3_U2480 );
nand NAND2_2752 ( P3_U4561 , P3_INSTQUEUE_REG_4__7_ , P3_U2479 );
nand NAND2_2753 ( P3_U4562 , P3_INSTQUEUE_REG_5__7_ , P3_U2478 );
nand NAND2_2754 ( P3_U4563 , P3_INSTQUEUE_REG_6__7_ , P3_U2477 );
nand NAND2_2755 ( P3_U4564 , P3_INSTQUEUE_REG_7__7_ , P3_U4471 );
nand NAND2_2756 ( P3_U4565 , P3_INSTQUEUE_REG_8__7_ , P3_U2476 );
nand NAND2_2757 ( P3_U4566 , P3_INSTQUEUE_REG_9__7_ , P3_U2475 );
nand NAND2_2758 ( P3_U4567 , P3_INSTQUEUE_REG_10__7_ , P3_U2473 );
nand NAND2_2759 ( P3_U4568 , P3_INSTQUEUE_REG_11__7_ , P3_U2471 );
nand NAND2_2760 ( P3_U4569 , P3_INSTQUEUE_REG_12__7_ , P3_U2470 );
nand NAND2_2761 ( P3_U4570 , P3_INSTQUEUE_REG_13__7_ , P3_U2469 );
nand NAND2_2762 ( P3_U4571 , P3_INSTQUEUE_REG_14__7_ , P3_U2467 );
nand NAND2_2763 ( P3_U4572 , P3_INSTQUEUE_REG_15__7_ , P3_U2465 );
not NOT1_2764 ( P3_U4573 , P3_U3218 );
nand NAND2_2765 ( P3_U4574 , P3_INSTQUEUE_REG_0__5_ , P3_U2484 );
nand NAND2_2766 ( P3_U4575 , P3_INSTQUEUE_REG_1__5_ , P3_U2483 );
nand NAND2_2767 ( P3_U4576 , P3_INSTQUEUE_REG_2__5_ , P3_U2482 );
nand NAND2_2768 ( P3_U4577 , P3_INSTQUEUE_REG_3__5_ , P3_U2480 );
nand NAND2_2769 ( P3_U4578 , P3_INSTQUEUE_REG_4__5_ , P3_U2479 );
nand NAND2_2770 ( P3_U4579 , P3_INSTQUEUE_REG_5__5_ , P3_U2478 );
nand NAND2_2771 ( P3_U4580 , P3_INSTQUEUE_REG_6__5_ , P3_U2477 );
nand NAND2_2772 ( P3_U4581 , P3_INSTQUEUE_REG_7__5_ , P3_U4471 );
nand NAND2_2773 ( P3_U4582 , P3_INSTQUEUE_REG_8__5_ , P3_U2476 );
nand NAND2_2774 ( P3_U4583 , P3_INSTQUEUE_REG_9__5_ , P3_U2475 );
nand NAND2_2775 ( P3_U4584 , P3_INSTQUEUE_REG_10__5_ , P3_U2473 );
nand NAND2_2776 ( P3_U4585 , P3_INSTQUEUE_REG_11__5_ , P3_U2471 );
nand NAND2_2777 ( P3_U4586 , P3_INSTQUEUE_REG_12__5_ , P3_U2470 );
nand NAND2_2778 ( P3_U4587 , P3_INSTQUEUE_REG_13__5_ , P3_U2469 );
nand NAND2_2779 ( P3_U4588 , P3_INSTQUEUE_REG_14__5_ , P3_U2467 );
nand NAND2_2780 ( P3_U4589 , P3_INSTQUEUE_REG_15__5_ , P3_U2465 );
not NOT1_2781 ( P3_U4590 , P3_U3110 );
nand NAND2_2782 ( P3_U4591 , P3_INSTQUEUE_REG_0__6_ , P3_U2484 );
nand NAND2_2783 ( P3_U4592 , P3_INSTQUEUE_REG_1__6_ , P3_U2483 );
nand NAND2_2784 ( P3_U4593 , P3_INSTQUEUE_REG_2__6_ , P3_U2482 );
nand NAND2_2785 ( P3_U4594 , P3_INSTQUEUE_REG_3__6_ , P3_U2480 );
nand NAND2_2786 ( P3_U4595 , P3_INSTQUEUE_REG_4__6_ , P3_U2479 );
nand NAND2_2787 ( P3_U4596 , P3_INSTQUEUE_REG_5__6_ , P3_U2478 );
nand NAND2_2788 ( P3_U4597 , P3_INSTQUEUE_REG_6__6_ , P3_U2477 );
nand NAND2_2789 ( P3_U4598 , P3_INSTQUEUE_REG_7__6_ , P3_U4471 );
nand NAND2_2790 ( P3_U4599 , P3_INSTQUEUE_REG_8__6_ , P3_U2476 );
nand NAND2_2791 ( P3_U4600 , P3_INSTQUEUE_REG_9__6_ , P3_U2475 );
nand NAND2_2792 ( P3_U4601 , P3_INSTQUEUE_REG_10__6_ , P3_U2473 );
nand NAND2_2793 ( P3_U4602 , P3_INSTQUEUE_REG_11__6_ , P3_U2471 );
nand NAND2_2794 ( P3_U4603 , P3_INSTQUEUE_REG_12__6_ , P3_U2470 );
nand NAND2_2795 ( P3_U4604 , P3_INSTQUEUE_REG_13__6_ , P3_U2469 );
nand NAND2_2796 ( P3_U4605 , P3_INSTQUEUE_REG_14__6_ , P3_U2467 );
nand NAND2_2797 ( P3_U4606 , P3_INSTQUEUE_REG_15__6_ , P3_U2465 );
not NOT1_2798 ( P3_U4607 , P3_U3074 );
not NOT1_2799 ( P3_U4608 , P3_U3113 );
nand NAND2_2800 ( P3_U4609 , P3_U2361 , P3_U3238 );
nand NAND2_2801 ( P3_U4610 , P3_U2360 , P3_U3237 );
nand NAND2_2802 ( P3_U4611 , P3_U2357 , P3_U3212 );
nand NAND2_2803 ( P3_U4612 , P3_U4305 , P3_U3215 );
nand NAND2_2804 ( P3_U4613 , P3_U4304 , P3_U3210 );
nand NAND2_2805 ( P3_U4614 , P3_U4303 , P3_U3213 );
nand NAND2_2806 ( P3_U4615 , P3_U2356 , P3_U3211 );
nand NAND2_2807 ( P3_U4616 , P3_U4302 , P3_U3214 );
nand NAND2_2808 ( P3_U4617 , P3_U3358 , P3_U3357 );
nand NAND5_2809 ( P3_U4618 , P3_U2463 , P3_U4522 , P3_U3360 , P3_U7945 , P3_U7944 );
not NOT1_2810 ( P3_U4619 , P3_U3109 );
nand NAND2_2811 ( P3_U4620 , P3_U4280 , P3_U4619 );
nand NAND2_2812 ( P3_U4621 , P3_U3359 , P3_U7916 );
not NOT1_2813 ( P3_U4622 , P3_U4281 );
not NOT1_2814 ( P3_U4623 , P3_U3262 );
or OR2_2815 ( P3_U4624 , P3_MORE_REG , P3_FLUSH_REG );
not NOT1_2816 ( P3_U4625 , P3_U3120 );
nand NAND2_2817 ( P3_U4626 , P3_U3353 , P3_U4303 );
nand NAND2_2818 ( P3_U4627 , P3_U3362 , P3_U4625 );
nand NAND2_2819 ( P3_U4628 , P3_STATE2_REG_1_ , U209 );
nand NAND3_2820 ( P3_U4629 , P3_U7953 , P3_U7952 , P3_STATE2_REG_2_ );
not NOT1_2821 ( P3_U4630 , P3_U3122 );
nand NAND3_2822 ( P3_U4631 , P3_U7957 , P3_U7956 , P3_STATE2_REG_1_ );
nand NAND2_2823 ( P3_U4632 , P3_STATE2_REG_2_ , P3_U3122 );
nand NAND2_2824 ( P3_U4633 , P3_U4629 , P3_U4338 );
nand NAND2_2825 ( P3_U4634 , P3_U3364 , P3_U4630 );
nand NAND2_2826 ( P3_U4635 , P3_STATE2_REG_1_ , P3_U4633 );
nand NAND2_2827 ( P3_U4636 , P3_U2390 , P3_U4629 );
nand NAND2_2828 ( P3_U4637 , P3_U4345 , P3_U4354 );
nand NAND2_2829 ( P3_U4638 , P3_U4629 , P3_U4337 );
nand NAND2_2830 ( P3_U4639 , P3_U2390 , P3_U3120 );
not NOT1_2831 ( P3_U4640 , P3_U3153 );
nand NAND2_2832 ( P3_U4641 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_U3128 );
not NOT1_2833 ( P3_U4642 , P3_U3137 );
not NOT1_2834 ( P3_U4643 , P3_U3141 );
not NOT1_2835 ( P3_U4644 , P3_U3148 );
not NOT1_2836 ( P3_U4645 , P3_U3155 );
not NOT1_2837 ( P3_U4646 , P3_U3156 );
not NOT1_2838 ( P3_U4647 , P3_U3143 );
not NOT1_2839 ( P3_U4648 , P3_U3130 );
not NOT1_2840 ( P3_U4649 , P3_U3132 );
not NOT1_2841 ( P3_U4650 , P3_U3180 );
nand NAND2_2842 ( P3_U4651 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_U3132 );
not NOT1_2843 ( P3_U4652 , P3_U3139 );
not NOT1_2844 ( P3_U4653 , P3_U3138 );
nand NAND2_2845 ( P3_U4654 , P3_U4653 , P3_U3269 );
nand NAND2_2846 ( P3_U4655 , P3_U4654 , P3_U3139 );
not NOT1_2847 ( P3_U4656 , P3_U3142 );
not NOT1_2848 ( P3_U4657 , P3_U3140 );
not NOT1_2849 ( P3_U4658 , P3_U3165 );
nand NAND2_2850 ( P3_U4659 , P3_U3140 , P3_U3142 );
not NOT1_2851 ( P3_U4660 , P3_U3182 );
not NOT1_2852 ( P3_U4661 , P3_U3144 );
not NOT1_2853 ( P3_U4662 , P3_U3134 );
nand NAND2_2854 ( P3_U4663 , P3_U2457 , P3_U4653 );
not NOT1_2855 ( P3_U4664 , P3_U3146 );
nand NAND2_2856 ( P3_U4665 , P3_STATE2_REG_1_ , P3_U3090 );
nand NAND3_2857 ( P3_U4666 , P3_U3124 , P3_U4665 , P3_U3126 );
nand NAND2_2858 ( P3_U4667 , P3_U4657 , P3_U2487 );
not NOT1_2859 ( P3_U4668 , P3_U3145 );
nand NAND2_2860 ( P3_U4669 , P3_U2489 , P3_U3145 );
nand NAND2_2861 ( P3_U4670 , P3_U4664 , P3_U4669 );
nand NAND2_2862 ( P3_U4671 , P3_STATE2_REG_3_ , P3_U3134 );
nand NAND2_2863 ( P3_U4672 , P3_U3369 , P3_U4670 );
nand NAND2_2864 ( P3_U4673 , P3_U4668 , P3_U4322 );
nand NAND2_2865 ( P3_U4674 , P3_U2489 , P3_U4673 );
nand NAND2_2866 ( P3_U4675 , P3_U2445 , P3_U4662 );
nand NAND2_2867 ( P3_U4676 , P3_U2436 , P3_U2488 );
nand NAND2_2868 ( P3_U4677 , P3_U2435 , P3_U4661 );
nand NAND2_2869 ( P3_U4678 , P3_U2378 , P3_U2420 );
nand NAND2_2870 ( P3_U4679 , P3_INSTQUEUE_REG_15__7_ , P3_U4672 );
nand NAND2_2871 ( P3_U4680 , P3_U2443 , P3_U4662 );
nand NAND2_2872 ( P3_U4681 , P3_U2434 , P3_U2488 );
nand NAND2_2873 ( P3_U4682 , P3_U2433 , P3_U4661 );
nand NAND2_2874 ( P3_U4683 , P3_U2419 , P3_U2378 );
nand NAND2_2875 ( P3_U4684 , P3_INSTQUEUE_REG_15__6_ , P3_U4672 );
nand NAND2_2876 ( P3_U4685 , P3_U2442 , P3_U4662 );
nand NAND2_2877 ( P3_U4686 , P3_U2432 , P3_U2488 );
nand NAND2_2878 ( P3_U4687 , P3_U2431 , P3_U4661 );
nand NAND2_2879 ( P3_U4688 , P3_U2418 , P3_U2378 );
nand NAND2_2880 ( P3_U4689 , P3_INSTQUEUE_REG_15__5_ , P3_U4672 );
nand NAND2_2881 ( P3_U4690 , P3_U2441 , P3_U4662 );
nand NAND2_2882 ( P3_U4691 , P3_U2430 , P3_U2488 );
nand NAND2_2883 ( P3_U4692 , P3_U2429 , P3_U4661 );
nand NAND2_2884 ( P3_U4693 , P3_U2417 , P3_U2378 );
nand NAND2_2885 ( P3_U4694 , P3_INSTQUEUE_REG_15__4_ , P3_U4672 );
nand NAND2_2886 ( P3_U4695 , P3_U2440 , P3_U4662 );
nand NAND2_2887 ( P3_U4696 , P3_U2428 , P3_U2488 );
nand NAND2_2888 ( P3_U4697 , P3_U2427 , P3_U4661 );
nand NAND2_2889 ( P3_U4698 , P3_U2416 , P3_U2378 );
nand NAND2_2890 ( P3_U4699 , P3_INSTQUEUE_REG_15__3_ , P3_U4672 );
nand NAND2_2891 ( P3_U4700 , P3_U2439 , P3_U4662 );
nand NAND2_2892 ( P3_U4701 , P3_U2426 , P3_U2488 );
nand NAND2_2893 ( P3_U4702 , P3_U2425 , P3_U4661 );
nand NAND2_2894 ( P3_U4703 , P3_U2415 , P3_U2378 );
nand NAND2_2895 ( P3_U4704 , P3_INSTQUEUE_REG_15__2_ , P3_U4672 );
nand NAND2_2896 ( P3_U4705 , P3_U2438 , P3_U4662 );
nand NAND2_2897 ( P3_U4706 , P3_U2424 , P3_U2488 );
nand NAND2_2898 ( P3_U4707 , P3_U2423 , P3_U4661 );
nand NAND2_2899 ( P3_U4708 , P3_U2414 , P3_U2378 );
nand NAND2_2900 ( P3_U4709 , P3_INSTQUEUE_REG_15__1_ , P3_U4672 );
nand NAND2_2901 ( P3_U4710 , P3_U2437 , P3_U4662 );
nand NAND2_2902 ( P3_U4711 , P3_U2422 , P3_U2488 );
nand NAND2_2903 ( P3_U4712 , P3_U2421 , P3_U4661 );
nand NAND2_2904 ( P3_U4713 , P3_U2413 , P3_U2378 );
nand NAND2_2905 ( P3_U4714 , P3_INSTQUEUE_REG_15__0_ , P3_U4672 );
not NOT1_2906 ( P3_U4715 , P3_U3149 );
not NOT1_2907 ( P3_U4716 , P3_U3147 );
nand NAND2_2908 ( P3_U4717 , P3_U4342 , P3_U2457 );
not NOT1_2909 ( P3_U4718 , P3_U3152 );
nand NAND2_2910 ( P3_U4719 , P3_U4644 , P3_U2487 );
not NOT1_2911 ( P3_U4720 , P3_U3151 );
nand NAND2_2912 ( P3_U4721 , P3_U2489 , P3_U3151 );
nand NAND2_2913 ( P3_U4722 , P3_U4718 , P3_U4721 );
nand NAND2_2914 ( P3_U4723 , P3_STATE2_REG_3_ , P3_U3147 );
nand NAND2_2915 ( P3_U4724 , P3_U3387 , P3_U4722 );
nand NAND2_2916 ( P3_U4725 , P3_U4720 , P3_U4322 );
nand NAND2_2917 ( P3_U4726 , P3_U2489 , P3_U4725 );
nand NAND2_2918 ( P3_U4727 , P3_U4716 , P3_U2445 );
nand NAND2_2919 ( P3_U4728 , P3_U2491 , P3_U2436 );
nand NAND2_2920 ( P3_U4729 , P3_U4715 , P3_U2435 );
nand NAND2_2921 ( P3_U4730 , P3_U2377 , P3_U2420 );
nand NAND2_2922 ( P3_U4731 , P3_INSTQUEUE_REG_14__7_ , P3_U4724 );
nand NAND2_2923 ( P3_U4732 , P3_U4716 , P3_U2443 );
nand NAND2_2924 ( P3_U4733 , P3_U2491 , P3_U2434 );
nand NAND2_2925 ( P3_U4734 , P3_U4715 , P3_U2433 );
nand NAND2_2926 ( P3_U4735 , P3_U2377 , P3_U2419 );
nand NAND2_2927 ( P3_U4736 , P3_INSTQUEUE_REG_14__6_ , P3_U4724 );
nand NAND2_2928 ( P3_U4737 , P3_U4716 , P3_U2442 );
nand NAND2_2929 ( P3_U4738 , P3_U2491 , P3_U2432 );
nand NAND2_2930 ( P3_U4739 , P3_U4715 , P3_U2431 );
nand NAND2_2931 ( P3_U4740 , P3_U2377 , P3_U2418 );
nand NAND2_2932 ( P3_U4741 , P3_INSTQUEUE_REG_14__5_ , P3_U4724 );
nand NAND2_2933 ( P3_U4742 , P3_U4716 , P3_U2441 );
nand NAND2_2934 ( P3_U4743 , P3_U2491 , P3_U2430 );
nand NAND2_2935 ( P3_U4744 , P3_U4715 , P3_U2429 );
nand NAND2_2936 ( P3_U4745 , P3_U2377 , P3_U2417 );
nand NAND2_2937 ( P3_U4746 , P3_INSTQUEUE_REG_14__4_ , P3_U4724 );
nand NAND2_2938 ( P3_U4747 , P3_U4716 , P3_U2440 );
nand NAND2_2939 ( P3_U4748 , P3_U2491 , P3_U2428 );
nand NAND2_2940 ( P3_U4749 , P3_U4715 , P3_U2427 );
nand NAND2_2941 ( P3_U4750 , P3_U2377 , P3_U2416 );
nand NAND2_2942 ( P3_U4751 , P3_INSTQUEUE_REG_14__3_ , P3_U4724 );
nand NAND2_2943 ( P3_U4752 , P3_U4716 , P3_U2439 );
nand NAND2_2944 ( P3_U4753 , P3_U2491 , P3_U2426 );
nand NAND2_2945 ( P3_U4754 , P3_U4715 , P3_U2425 );
nand NAND2_2946 ( P3_U4755 , P3_U2377 , P3_U2415 );
nand NAND2_2947 ( P3_U4756 , P3_INSTQUEUE_REG_14__2_ , P3_U4724 );
nand NAND2_2948 ( P3_U4757 , P3_U4716 , P3_U2438 );
nand NAND2_2949 ( P3_U4758 , P3_U2491 , P3_U2424 );
nand NAND2_2950 ( P3_U4759 , P3_U4715 , P3_U2423 );
nand NAND2_2951 ( P3_U4760 , P3_U2377 , P3_U2414 );
nand NAND2_2952 ( P3_U4761 , P3_INSTQUEUE_REG_14__1_ , P3_U4724 );
nand NAND2_2953 ( P3_U4762 , P3_U4716 , P3_U2437 );
nand NAND2_2954 ( P3_U4763 , P3_U2491 , P3_U2422 );
nand NAND2_2955 ( P3_U4764 , P3_U4715 , P3_U2421 );
nand NAND2_2956 ( P3_U4765 , P3_U2377 , P3_U2413 );
nand NAND2_2957 ( P3_U4766 , P3_INSTQUEUE_REG_14__0_ , P3_U4724 );
not NOT1_2958 ( P3_U4767 , P3_U3157 );
not NOT1_2959 ( P3_U4768 , P3_U3154 );
nand NAND2_2960 ( P3_U4769 , P3_U4343 , P3_U2457 );
not NOT1_2961 ( P3_U4770 , P3_U3160 );
nand NAND2_2962 ( P3_U4771 , P3_U4645 , P3_U2487 );
not NOT1_2963 ( P3_U4772 , P3_U3159 );
nand NAND2_2964 ( P3_U4773 , P3_U2489 , P3_U3159 );
nand NAND2_2965 ( P3_U4774 , P3_U4770 , P3_U4773 );
nand NAND2_2966 ( P3_U4775 , P3_STATE2_REG_3_ , P3_U3154 );
nand NAND2_2967 ( P3_U4776 , P3_U3405 , P3_U4774 );
nand NAND2_2968 ( P3_U4777 , P3_U4772 , P3_U4322 );
nand NAND2_2969 ( P3_U4778 , P3_U2489 , P3_U4777 );
nand NAND2_2970 ( P3_U4779 , P3_U4768 , P3_U2445 );
nand NAND2_2971 ( P3_U4780 , P3_U2494 , P3_U2436 );
nand NAND2_2972 ( P3_U4781 , P3_U4767 , P3_U2435 );
nand NAND2_2973 ( P3_U4782 , P3_U2376 , P3_U2420 );
nand NAND2_2974 ( P3_U4783 , P3_INSTQUEUE_REG_13__7_ , P3_U4776 );
nand NAND2_2975 ( P3_U4784 , P3_U4768 , P3_U2443 );
nand NAND2_2976 ( P3_U4785 , P3_U2494 , P3_U2434 );
nand NAND2_2977 ( P3_U4786 , P3_U4767 , P3_U2433 );
nand NAND2_2978 ( P3_U4787 , P3_U2376 , P3_U2419 );
nand NAND2_2979 ( P3_U4788 , P3_INSTQUEUE_REG_13__6_ , P3_U4776 );
nand NAND2_2980 ( P3_U4789 , P3_U4768 , P3_U2442 );
nand NAND2_2981 ( P3_U4790 , P3_U2494 , P3_U2432 );
nand NAND2_2982 ( P3_U4791 , P3_U4767 , P3_U2431 );
nand NAND2_2983 ( P3_U4792 , P3_U2376 , P3_U2418 );
nand NAND2_2984 ( P3_U4793 , P3_INSTQUEUE_REG_13__5_ , P3_U4776 );
nand NAND2_2985 ( P3_U4794 , P3_U4768 , P3_U2441 );
nand NAND2_2986 ( P3_U4795 , P3_U2494 , P3_U2430 );
nand NAND2_2987 ( P3_U4796 , P3_U4767 , P3_U2429 );
nand NAND2_2988 ( P3_U4797 , P3_U2376 , P3_U2417 );
nand NAND2_2989 ( P3_U4798 , P3_INSTQUEUE_REG_13__4_ , P3_U4776 );
nand NAND2_2990 ( P3_U4799 , P3_U4768 , P3_U2440 );
nand NAND2_2991 ( P3_U4800 , P3_U2494 , P3_U2428 );
nand NAND2_2992 ( P3_U4801 , P3_U4767 , P3_U2427 );
nand NAND2_2993 ( P3_U4802 , P3_U2376 , P3_U2416 );
nand NAND2_2994 ( P3_U4803 , P3_INSTQUEUE_REG_13__3_ , P3_U4776 );
nand NAND2_2995 ( P3_U4804 , P3_U4768 , P3_U2439 );
nand NAND2_2996 ( P3_U4805 , P3_U2494 , P3_U2426 );
nand NAND2_2997 ( P3_U4806 , P3_U4767 , P3_U2425 );
nand NAND2_2998 ( P3_U4807 , P3_U2376 , P3_U2415 );
nand NAND2_2999 ( P3_U4808 , P3_INSTQUEUE_REG_13__2_ , P3_U4776 );
nand NAND2_3000 ( P3_U4809 , P3_U4768 , P3_U2438 );
nand NAND2_3001 ( P3_U4810 , P3_U2494 , P3_U2424 );
nand NAND2_3002 ( P3_U4811 , P3_U4767 , P3_U2423 );
nand NAND2_3003 ( P3_U4812 , P3_U2376 , P3_U2414 );
nand NAND2_3004 ( P3_U4813 , P3_INSTQUEUE_REG_13__1_ , P3_U4776 );
nand NAND2_3005 ( P3_U4814 , P3_U4768 , P3_U2437 );
nand NAND2_3006 ( P3_U4815 , P3_U2494 , P3_U2422 );
nand NAND2_3007 ( P3_U4816 , P3_U4767 , P3_U2421 );
nand NAND2_3008 ( P3_U4817 , P3_U2376 , P3_U2413 );
nand NAND2_3009 ( P3_U4818 , P3_INSTQUEUE_REG_13__0_ , P3_U4776 );
not NOT1_3010 ( P3_U4819 , P3_U3162 );
not NOT1_3011 ( P3_U4820 , P3_U3161 );
not NOT1_3012 ( P3_U4821 , P3_U3070 );
nand NAND2_3013 ( P3_U4822 , P3_U2496 , P3_U2487 );
not NOT1_3014 ( P3_U4823 , P3_U3163 );
nand NAND2_3015 ( P3_U4824 , P3_U2489 , P3_U3163 );
nand NAND2_3016 ( P3_U4825 , P3_U4824 , P3_U3070 );
nand NAND2_3017 ( P3_U4826 , P3_STATE2_REG_3_ , P3_U3161 );
nand NAND2_3018 ( P3_U4827 , P3_U3423 , P3_U4825 );
nand NAND2_3019 ( P3_U4828 , P3_U4823 , P3_U4322 );
nand NAND2_3020 ( P3_U4829 , P3_U2489 , P3_U4828 );
nand NAND2_3021 ( P3_U4830 , P3_U4820 , P3_U2445 );
nand NAND2_3022 ( P3_U4831 , P3_U2497 , P3_U2436 );
nand NAND2_3023 ( P3_U4832 , P3_U4819 , P3_U2435 );
nand NAND2_3024 ( P3_U4833 , P3_U2375 , P3_U2420 );
nand NAND2_3025 ( P3_U4834 , P3_INSTQUEUE_REG_12__7_ , P3_U4827 );
nand NAND2_3026 ( P3_U4835 , P3_U4820 , P3_U2443 );
nand NAND2_3027 ( P3_U4836 , P3_U2497 , P3_U2434 );
nand NAND2_3028 ( P3_U4837 , P3_U4819 , P3_U2433 );
nand NAND2_3029 ( P3_U4838 , P3_U2375 , P3_U2419 );
nand NAND2_3030 ( P3_U4839 , P3_INSTQUEUE_REG_12__6_ , P3_U4827 );
nand NAND2_3031 ( P3_U4840 , P3_U4820 , P3_U2442 );
nand NAND2_3032 ( P3_U4841 , P3_U2497 , P3_U2432 );
nand NAND2_3033 ( P3_U4842 , P3_U4819 , P3_U2431 );
nand NAND2_3034 ( P3_U4843 , P3_U2375 , P3_U2418 );
nand NAND2_3035 ( P3_U4844 , P3_INSTQUEUE_REG_12__5_ , P3_U4827 );
nand NAND2_3036 ( P3_U4845 , P3_U4820 , P3_U2441 );
nand NAND2_3037 ( P3_U4846 , P3_U2497 , P3_U2430 );
nand NAND2_3038 ( P3_U4847 , P3_U4819 , P3_U2429 );
nand NAND2_3039 ( P3_U4848 , P3_U2375 , P3_U2417 );
nand NAND2_3040 ( P3_U4849 , P3_INSTQUEUE_REG_12__4_ , P3_U4827 );
nand NAND2_3041 ( P3_U4850 , P3_U4820 , P3_U2440 );
nand NAND2_3042 ( P3_U4851 , P3_U2497 , P3_U2428 );
nand NAND2_3043 ( P3_U4852 , P3_U4819 , P3_U2427 );
nand NAND2_3044 ( P3_U4853 , P3_U2375 , P3_U2416 );
nand NAND2_3045 ( P3_U4854 , P3_INSTQUEUE_REG_12__3_ , P3_U4827 );
nand NAND2_3046 ( P3_U4855 , P3_U4820 , P3_U2439 );
nand NAND2_3047 ( P3_U4856 , P3_U2497 , P3_U2426 );
nand NAND2_3048 ( P3_U4857 , P3_U4819 , P3_U2425 );
nand NAND2_3049 ( P3_U4858 , P3_U2375 , P3_U2415 );
nand NAND2_3050 ( P3_U4859 , P3_INSTQUEUE_REG_12__2_ , P3_U4827 );
nand NAND2_3051 ( P3_U4860 , P3_U4820 , P3_U2438 );
nand NAND2_3052 ( P3_U4861 , P3_U2497 , P3_U2424 );
nand NAND2_3053 ( P3_U4862 , P3_U4819 , P3_U2423 );
nand NAND2_3054 ( P3_U4863 , P3_U2375 , P3_U2414 );
nand NAND2_3055 ( P3_U4864 , P3_INSTQUEUE_REG_12__1_ , P3_U4827 );
nand NAND2_3056 ( P3_U4865 , P3_U4820 , P3_U2437 );
nand NAND2_3057 ( P3_U4866 , P3_U2497 , P3_U2422 );
nand NAND2_3058 ( P3_U4867 , P3_U4819 , P3_U2421 );
nand NAND2_3059 ( P3_U4868 , P3_U2375 , P3_U2413 );
nand NAND2_3060 ( P3_U4869 , P3_INSTQUEUE_REG_12__0_ , P3_U4827 );
not NOT1_3061 ( P3_U4870 , P3_U3166 );
not NOT1_3062 ( P3_U4871 , P3_U3164 );
nand NAND2_3063 ( P3_U4872 , P3_U2459 , P3_U4653 );
not NOT1_3064 ( P3_U4873 , P3_U3168 );
nand NAND2_3065 ( P3_U4874 , P3_U4658 , P3_U4657 );
not NOT1_3066 ( P3_U4875 , P3_U3167 );
nand NAND2_3067 ( P3_U4876 , P3_U2489 , P3_U3167 );
nand NAND2_3068 ( P3_U4877 , P3_U4873 , P3_U4876 );
nand NAND2_3069 ( P3_U4878 , P3_STATE2_REG_3_ , P3_U3164 );
nand NAND2_3070 ( P3_U4879 , P3_U3440 , P3_U4877 );
nand NAND2_3071 ( P3_U4880 , P3_U4875 , P3_U4322 );
nand NAND2_3072 ( P3_U4881 , P3_U2489 , P3_U4880 );
nand NAND2_3073 ( P3_U4882 , P3_U4871 , P3_U2445 );
nand NAND2_3074 ( P3_U4883 , P3_U2499 , P3_U2436 );
nand NAND2_3075 ( P3_U4884 , P3_U4870 , P3_U2435 );
nand NAND2_3076 ( P3_U4885 , P3_U2374 , P3_U2420 );
nand NAND2_3077 ( P3_U4886 , P3_INSTQUEUE_REG_11__7_ , P3_U4879 );
nand NAND2_3078 ( P3_U4887 , P3_U4871 , P3_U2443 );
nand NAND2_3079 ( P3_U4888 , P3_U2499 , P3_U2434 );
nand NAND2_3080 ( P3_U4889 , P3_U4870 , P3_U2433 );
nand NAND2_3081 ( P3_U4890 , P3_U2374 , P3_U2419 );
nand NAND2_3082 ( P3_U4891 , P3_INSTQUEUE_REG_11__6_ , P3_U4879 );
nand NAND2_3083 ( P3_U4892 , P3_U4871 , P3_U2442 );
nand NAND2_3084 ( P3_U4893 , P3_U2499 , P3_U2432 );
nand NAND2_3085 ( P3_U4894 , P3_U4870 , P3_U2431 );
nand NAND2_3086 ( P3_U4895 , P3_U2374 , P3_U2418 );
nand NAND2_3087 ( P3_U4896 , P3_INSTQUEUE_REG_11__5_ , P3_U4879 );
nand NAND2_3088 ( P3_U4897 , P3_U4871 , P3_U2441 );
nand NAND2_3089 ( P3_U4898 , P3_U2499 , P3_U2430 );
nand NAND2_3090 ( P3_U4899 , P3_U4870 , P3_U2429 );
nand NAND2_3091 ( P3_U4900 , P3_U2374 , P3_U2417 );
nand NAND2_3092 ( P3_U4901 , P3_INSTQUEUE_REG_11__4_ , P3_U4879 );
nand NAND2_3093 ( P3_U4902 , P3_U4871 , P3_U2440 );
nand NAND2_3094 ( P3_U4903 , P3_U2499 , P3_U2428 );
nand NAND2_3095 ( P3_U4904 , P3_U4870 , P3_U2427 );
nand NAND2_3096 ( P3_U4905 , P3_U2374 , P3_U2416 );
nand NAND2_3097 ( P3_U4906 , P3_INSTQUEUE_REG_11__3_ , P3_U4879 );
nand NAND2_3098 ( P3_U4907 , P3_U4871 , P3_U2439 );
nand NAND2_3099 ( P3_U4908 , P3_U2499 , P3_U2426 );
nand NAND2_3100 ( P3_U4909 , P3_U4870 , P3_U2425 );
nand NAND2_3101 ( P3_U4910 , P3_U2374 , P3_U2415 );
nand NAND2_3102 ( P3_U4911 , P3_INSTQUEUE_REG_11__2_ , P3_U4879 );
nand NAND2_3103 ( P3_U4912 , P3_U4871 , P3_U2438 );
nand NAND2_3104 ( P3_U4913 , P3_U2499 , P3_U2424 );
nand NAND2_3105 ( P3_U4914 , P3_U4870 , P3_U2423 );
nand NAND2_3106 ( P3_U4915 , P3_U2374 , P3_U2414 );
nand NAND2_3107 ( P3_U4916 , P3_INSTQUEUE_REG_11__1_ , P3_U4879 );
nand NAND2_3108 ( P3_U4917 , P3_U4871 , P3_U2437 );
nand NAND2_3109 ( P3_U4918 , P3_U2499 , P3_U2422 );
nand NAND2_3110 ( P3_U4919 , P3_U4870 , P3_U2421 );
nand NAND2_3111 ( P3_U4920 , P3_U2374 , P3_U2413 );
nand NAND2_3112 ( P3_U4921 , P3_INSTQUEUE_REG_11__0_ , P3_U4879 );
not NOT1_3113 ( P3_U4922 , P3_U3170 );
not NOT1_3114 ( P3_U4923 , P3_U3169 );
nand NAND2_3115 ( P3_U4924 , P3_U2459 , P3_U4342 );
not NOT1_3116 ( P3_U4925 , P3_U3172 );
nand NAND2_3117 ( P3_U4926 , P3_U4658 , P3_U4644 );
not NOT1_3118 ( P3_U4927 , P3_U3171 );
nand NAND2_3119 ( P3_U4928 , P3_U2489 , P3_U3171 );
nand NAND2_3120 ( P3_U4929 , P3_U4925 , P3_U4928 );
nand NAND2_3121 ( P3_U4930 , P3_STATE2_REG_3_ , P3_U3169 );
nand NAND2_3122 ( P3_U4931 , P3_U3458 , P3_U4929 );
nand NAND2_3123 ( P3_U4932 , P3_U4927 , P3_U4322 );
nand NAND2_3124 ( P3_U4933 , P3_U2489 , P3_U4932 );
nand NAND2_3125 ( P3_U4934 , P3_U4923 , P3_U2445 );
nand NAND2_3126 ( P3_U4935 , P3_U2500 , P3_U2436 );
nand NAND2_3127 ( P3_U4936 , P3_U4922 , P3_U2435 );
nand NAND2_3128 ( P3_U4937 , P3_U2373 , P3_U2420 );
nand NAND2_3129 ( P3_U4938 , P3_INSTQUEUE_REG_10__7_ , P3_U4931 );
nand NAND2_3130 ( P3_U4939 , P3_U4923 , P3_U2443 );
nand NAND2_3131 ( P3_U4940 , P3_U2500 , P3_U2434 );
nand NAND2_3132 ( P3_U4941 , P3_U4922 , P3_U2433 );
nand NAND2_3133 ( P3_U4942 , P3_U2373 , P3_U2419 );
nand NAND2_3134 ( P3_U4943 , P3_INSTQUEUE_REG_10__6_ , P3_U4931 );
nand NAND2_3135 ( P3_U4944 , P3_U4923 , P3_U2442 );
nand NAND2_3136 ( P3_U4945 , P3_U2500 , P3_U2432 );
nand NAND2_3137 ( P3_U4946 , P3_U4922 , P3_U2431 );
nand NAND2_3138 ( P3_U4947 , P3_U2373 , P3_U2418 );
nand NAND2_3139 ( P3_U4948 , P3_INSTQUEUE_REG_10__5_ , P3_U4931 );
nand NAND2_3140 ( P3_U4949 , P3_U4923 , P3_U2441 );
nand NAND2_3141 ( P3_U4950 , P3_U2500 , P3_U2430 );
nand NAND2_3142 ( P3_U4951 , P3_U4922 , P3_U2429 );
nand NAND2_3143 ( P3_U4952 , P3_U2373 , P3_U2417 );
nand NAND2_3144 ( P3_U4953 , P3_INSTQUEUE_REG_10__4_ , P3_U4931 );
nand NAND2_3145 ( P3_U4954 , P3_U4923 , P3_U2440 );
nand NAND2_3146 ( P3_U4955 , P3_U2500 , P3_U2428 );
nand NAND2_3147 ( P3_U4956 , P3_U4922 , P3_U2427 );
nand NAND2_3148 ( P3_U4957 , P3_U2373 , P3_U2416 );
nand NAND2_3149 ( P3_U4958 , P3_INSTQUEUE_REG_10__3_ , P3_U4931 );
nand NAND2_3150 ( P3_U4959 , P3_U4923 , P3_U2439 );
nand NAND2_3151 ( P3_U4960 , P3_U2500 , P3_U2426 );
nand NAND2_3152 ( P3_U4961 , P3_U4922 , P3_U2425 );
nand NAND2_3153 ( P3_U4962 , P3_U2373 , P3_U2415 );
nand NAND2_3154 ( P3_U4963 , P3_INSTQUEUE_REG_10__2_ , P3_U4931 );
nand NAND2_3155 ( P3_U4964 , P3_U4923 , P3_U2438 );
nand NAND2_3156 ( P3_U4965 , P3_U2500 , P3_U2424 );
nand NAND2_3157 ( P3_U4966 , P3_U4922 , P3_U2423 );
nand NAND2_3158 ( P3_U4967 , P3_U2373 , P3_U2414 );
nand NAND2_3159 ( P3_U4968 , P3_INSTQUEUE_REG_10__1_ , P3_U4931 );
nand NAND2_3160 ( P3_U4969 , P3_U4923 , P3_U2437 );
nand NAND2_3161 ( P3_U4970 , P3_U2500 , P3_U2422 );
nand NAND2_3162 ( P3_U4971 , P3_U4922 , P3_U2421 );
nand NAND2_3163 ( P3_U4972 , P3_U2373 , P3_U2413 );
nand NAND2_3164 ( P3_U4973 , P3_INSTQUEUE_REG_10__0_ , P3_U4931 );
not NOT1_3165 ( P3_U4974 , P3_U3174 );
not NOT1_3166 ( P3_U4975 , P3_U3173 );
nand NAND2_3167 ( P3_U4976 , P3_U2459 , P3_U4343 );
not NOT1_3168 ( P3_U4977 , P3_U3176 );
nand NAND2_3169 ( P3_U4978 , P3_U4658 , P3_U4645 );
not NOT1_3170 ( P3_U4979 , P3_U3175 );
nand NAND2_3171 ( P3_U4980 , P3_U2489 , P3_U3175 );
nand NAND2_3172 ( P3_U4981 , P3_U4977 , P3_U4980 );
nand NAND2_3173 ( P3_U4982 , P3_STATE2_REG_3_ , P3_U3173 );
nand NAND2_3174 ( P3_U4983 , P3_U3476 , P3_U4981 );
nand NAND2_3175 ( P3_U4984 , P3_U4979 , P3_U4322 );
nand NAND2_3176 ( P3_U4985 , P3_U2489 , P3_U4984 );
nand NAND2_3177 ( P3_U4986 , P3_U4975 , P3_U2445 );
nand NAND2_3178 ( P3_U4987 , P3_U2502 , P3_U2436 );
nand NAND2_3179 ( P3_U4988 , P3_U4974 , P3_U2435 );
nand NAND2_3180 ( P3_U4989 , P3_U2372 , P3_U2420 );
nand NAND2_3181 ( P3_U4990 , P3_INSTQUEUE_REG_9__7_ , P3_U4983 );
nand NAND2_3182 ( P3_U4991 , P3_U4975 , P3_U2443 );
nand NAND2_3183 ( P3_U4992 , P3_U2502 , P3_U2434 );
nand NAND2_3184 ( P3_U4993 , P3_U4974 , P3_U2433 );
nand NAND2_3185 ( P3_U4994 , P3_U2372 , P3_U2419 );
nand NAND2_3186 ( P3_U4995 , P3_INSTQUEUE_REG_9__6_ , P3_U4983 );
nand NAND2_3187 ( P3_U4996 , P3_U4975 , P3_U2442 );
nand NAND2_3188 ( P3_U4997 , P3_U2502 , P3_U2432 );
nand NAND2_3189 ( P3_U4998 , P3_U4974 , P3_U2431 );
nand NAND2_3190 ( P3_U4999 , P3_U2372 , P3_U2418 );
nand NAND2_3191 ( P3_U5000 , P3_INSTQUEUE_REG_9__5_ , P3_U4983 );
nand NAND2_3192 ( P3_U5001 , P3_U4975 , P3_U2441 );
nand NAND2_3193 ( P3_U5002 , P3_U2502 , P3_U2430 );
nand NAND2_3194 ( P3_U5003 , P3_U4974 , P3_U2429 );
nand NAND2_3195 ( P3_U5004 , P3_U2372 , P3_U2417 );
nand NAND2_3196 ( P3_U5005 , P3_INSTQUEUE_REG_9__4_ , P3_U4983 );
nand NAND2_3197 ( P3_U5006 , P3_U4975 , P3_U2440 );
nand NAND2_3198 ( P3_U5007 , P3_U2502 , P3_U2428 );
nand NAND2_3199 ( P3_U5008 , P3_U4974 , P3_U2427 );
nand NAND2_3200 ( P3_U5009 , P3_U2372 , P3_U2416 );
nand NAND2_3201 ( P3_U5010 , P3_INSTQUEUE_REG_9__3_ , P3_U4983 );
nand NAND2_3202 ( P3_U5011 , P3_U4975 , P3_U2439 );
nand NAND2_3203 ( P3_U5012 , P3_U2502 , P3_U2426 );
nand NAND2_3204 ( P3_U5013 , P3_U4974 , P3_U2425 );
nand NAND2_3205 ( P3_U5014 , P3_U2372 , P3_U2415 );
nand NAND2_3206 ( P3_U5015 , P3_INSTQUEUE_REG_9__2_ , P3_U4983 );
nand NAND2_3207 ( P3_U5016 , P3_U4975 , P3_U2438 );
nand NAND2_3208 ( P3_U5017 , P3_U2502 , P3_U2424 );
nand NAND2_3209 ( P3_U5018 , P3_U4974 , P3_U2423 );
nand NAND2_3210 ( P3_U5019 , P3_U2372 , P3_U2414 );
nand NAND2_3211 ( P3_U5020 , P3_INSTQUEUE_REG_9__1_ , P3_U4983 );
nand NAND2_3212 ( P3_U5021 , P3_U4975 , P3_U2437 );
nand NAND2_3213 ( P3_U5022 , P3_U2502 , P3_U2422 );
nand NAND2_3214 ( P3_U5023 , P3_U4974 , P3_U2421 );
nand NAND2_3215 ( P3_U5024 , P3_U2372 , P3_U2413 );
nand NAND2_3216 ( P3_U5025 , P3_INSTQUEUE_REG_9__0_ , P3_U4983 );
not NOT1_3217 ( P3_U5026 , P3_U3178 );
not NOT1_3218 ( P3_U5027 , P3_U3177 );
not NOT1_3219 ( P3_U5028 , P3_U3071 );
nand NAND2_3220 ( P3_U5029 , P3_U4658 , P3_U2496 );
not NOT1_3221 ( P3_U5030 , P3_U3179 );
nand NAND2_3222 ( P3_U5031 , P3_U2489 , P3_U3179 );
nand NAND2_3223 ( P3_U5032 , P3_U5031 , P3_U3071 );
nand NAND2_3224 ( P3_U5033 , P3_STATE2_REG_3_ , P3_U3177 );
nand NAND2_3225 ( P3_U5034 , P3_U3493 , P3_U5032 );
nand NAND2_3226 ( P3_U5035 , P3_U5030 , P3_U4322 );
nand NAND2_3227 ( P3_U5036 , P3_U2489 , P3_U5035 );
nand NAND2_3228 ( P3_U5037 , P3_U5027 , P3_U2445 );
nand NAND2_3229 ( P3_U5038 , P3_U2503 , P3_U2436 );
nand NAND2_3230 ( P3_U5039 , P3_U5026 , P3_U2435 );
nand NAND2_3231 ( P3_U5040 , P3_U2371 , P3_U2420 );
nand NAND2_3232 ( P3_U5041 , P3_INSTQUEUE_REG_8__7_ , P3_U5034 );
nand NAND2_3233 ( P3_U5042 , P3_U5027 , P3_U2443 );
nand NAND2_3234 ( P3_U5043 , P3_U2503 , P3_U2434 );
nand NAND2_3235 ( P3_U5044 , P3_U5026 , P3_U2433 );
nand NAND2_3236 ( P3_U5045 , P3_U2371 , P3_U2419 );
nand NAND2_3237 ( P3_U5046 , P3_INSTQUEUE_REG_8__6_ , P3_U5034 );
nand NAND2_3238 ( P3_U5047 , P3_U5027 , P3_U2442 );
nand NAND2_3239 ( P3_U5048 , P3_U2503 , P3_U2432 );
nand NAND2_3240 ( P3_U5049 , P3_U5026 , P3_U2431 );
nand NAND2_3241 ( P3_U5050 , P3_U2371 , P3_U2418 );
nand NAND2_3242 ( P3_U5051 , P3_INSTQUEUE_REG_8__5_ , P3_U5034 );
nand NAND2_3243 ( P3_U5052 , P3_U5027 , P3_U2441 );
nand NAND2_3244 ( P3_U5053 , P3_U2503 , P3_U2430 );
nand NAND2_3245 ( P3_U5054 , P3_U5026 , P3_U2429 );
nand NAND2_3246 ( P3_U5055 , P3_U2371 , P3_U2417 );
nand NAND2_3247 ( P3_U5056 , P3_INSTQUEUE_REG_8__4_ , P3_U5034 );
nand NAND2_3248 ( P3_U5057 , P3_U5027 , P3_U2440 );
nand NAND2_3249 ( P3_U5058 , P3_U2503 , P3_U2428 );
nand NAND2_3250 ( P3_U5059 , P3_U5026 , P3_U2427 );
nand NAND2_3251 ( P3_U5060 , P3_U2371 , P3_U2416 );
nand NAND2_3252 ( P3_U5061 , P3_INSTQUEUE_REG_8__3_ , P3_U5034 );
nand NAND2_3253 ( P3_U5062 , P3_U5027 , P3_U2439 );
nand NAND2_3254 ( P3_U5063 , P3_U2503 , P3_U2426 );
nand NAND2_3255 ( P3_U5064 , P3_U5026 , P3_U2425 );
nand NAND2_3256 ( P3_U5065 , P3_U2371 , P3_U2415 );
nand NAND2_3257 ( P3_U5066 , P3_INSTQUEUE_REG_8__2_ , P3_U5034 );
nand NAND2_3258 ( P3_U5067 , P3_U5027 , P3_U2438 );
nand NAND2_3259 ( P3_U5068 , P3_U2503 , P3_U2424 );
nand NAND2_3260 ( P3_U5069 , P3_U5026 , P3_U2423 );
nand NAND2_3261 ( P3_U5070 , P3_U2371 , P3_U2414 );
nand NAND2_3262 ( P3_U5071 , P3_INSTQUEUE_REG_8__1_ , P3_U5034 );
nand NAND2_3263 ( P3_U5072 , P3_U5027 , P3_U2437 );
nand NAND2_3264 ( P3_U5073 , P3_U2503 , P3_U2422 );
nand NAND2_3265 ( P3_U5074 , P3_U5026 , P3_U2421 );
nand NAND2_3266 ( P3_U5075 , P3_U2371 , P3_U2413 );
nand NAND2_3267 ( P3_U5076 , P3_INSTQUEUE_REG_8__0_ , P3_U5034 );
not NOT1_3268 ( P3_U5077 , P3_U3183 );
not NOT1_3269 ( P3_U5078 , P3_U3185 );
not NOT1_3270 ( P3_U5079 , P3_U3184 );
nand NAND2_3271 ( P3_U5080 , P3_U2489 , P3_U3184 );
nand NAND2_3272 ( P3_U5081 , P3_U5078 , P3_U5080 );
nand NAND2_3273 ( P3_U5082 , P3_STATE2_REG_3_ , P3_U3180 );
nand NAND2_3274 ( P3_U5083 , P3_U3510 , P3_U5081 );
nand NAND2_3275 ( P3_U5084 , P3_U5079 , P3_U4322 );
nand NAND2_3276 ( P3_U5085 , P3_U2489 , P3_U5084 );
nand NAND2_3277 ( P3_U5086 , P3_U4650 , P3_U2445 );
nand NAND2_3278 ( P3_U5087 , P3_U4326 , P3_U2436 );
nand NAND2_3279 ( P3_U5088 , P3_U5077 , P3_U2435 );
nand NAND2_3280 ( P3_U5089 , P3_U2370 , P3_U2420 );
nand NAND2_3281 ( P3_U5090 , P3_INSTQUEUE_REG_7__7_ , P3_U5083 );
nand NAND2_3282 ( P3_U5091 , P3_U4650 , P3_U2443 );
nand NAND2_3283 ( P3_U5092 , P3_U4326 , P3_U2434 );
nand NAND2_3284 ( P3_U5093 , P3_U5077 , P3_U2433 );
nand NAND2_3285 ( P3_U5094 , P3_U2370 , P3_U2419 );
nand NAND2_3286 ( P3_U5095 , P3_INSTQUEUE_REG_7__6_ , P3_U5083 );
nand NAND2_3287 ( P3_U5096 , P3_U4650 , P3_U2442 );
nand NAND2_3288 ( P3_U5097 , P3_U4326 , P3_U2432 );
nand NAND2_3289 ( P3_U5098 , P3_U5077 , P3_U2431 );
nand NAND2_3290 ( P3_U5099 , P3_U2370 , P3_U2418 );
nand NAND2_3291 ( P3_U5100 , P3_INSTQUEUE_REG_7__5_ , P3_U5083 );
nand NAND2_3292 ( P3_U5101 , P3_U4650 , P3_U2441 );
nand NAND2_3293 ( P3_U5102 , P3_U4326 , P3_U2430 );
nand NAND2_3294 ( P3_U5103 , P3_U5077 , P3_U2429 );
nand NAND2_3295 ( P3_U5104 , P3_U2370 , P3_U2417 );
nand NAND2_3296 ( P3_U5105 , P3_INSTQUEUE_REG_7__4_ , P3_U5083 );
nand NAND2_3297 ( P3_U5106 , P3_U4650 , P3_U2440 );
nand NAND2_3298 ( P3_U5107 , P3_U4326 , P3_U2428 );
nand NAND2_3299 ( P3_U5108 , P3_U5077 , P3_U2427 );
nand NAND2_3300 ( P3_U5109 , P3_U2370 , P3_U2416 );
nand NAND2_3301 ( P3_U5110 , P3_INSTQUEUE_REG_7__3_ , P3_U5083 );
nand NAND2_3302 ( P3_U5111 , P3_U4650 , P3_U2439 );
nand NAND2_3303 ( P3_U5112 , P3_U4326 , P3_U2426 );
nand NAND2_3304 ( P3_U5113 , P3_U5077 , P3_U2425 );
nand NAND2_3305 ( P3_U5114 , P3_U2370 , P3_U2415 );
nand NAND2_3306 ( P3_U5115 , P3_INSTQUEUE_REG_7__2_ , P3_U5083 );
nand NAND2_3307 ( P3_U5116 , P3_U4650 , P3_U2438 );
nand NAND2_3308 ( P3_U5117 , P3_U4326 , P3_U2424 );
nand NAND2_3309 ( P3_U5118 , P3_U5077 , P3_U2423 );
nand NAND2_3310 ( P3_U5119 , P3_U2370 , P3_U2414 );
nand NAND2_3311 ( P3_U5120 , P3_INSTQUEUE_REG_7__1_ , P3_U5083 );
nand NAND2_3312 ( P3_U5121 , P3_U4650 , P3_U2437 );
nand NAND2_3313 ( P3_U5122 , P3_U4326 , P3_U2422 );
nand NAND2_3314 ( P3_U5123 , P3_U5077 , P3_U2421 );
nand NAND2_3315 ( P3_U5124 , P3_U2370 , P3_U2413 );
nand NAND2_3316 ( P3_U5125 , P3_INSTQUEUE_REG_7__0_ , P3_U5083 );
not NOT1_3317 ( P3_U5126 , P3_U3187 );
not NOT1_3318 ( P3_U5127 , P3_U3186 );
nand NAND2_3319 ( P3_U5128 , P3_U4342 , P3_U2458 );
not NOT1_3320 ( P3_U5129 , P3_U3189 );
nand NAND2_3321 ( P3_U5130 , P3_U4644 , P3_U2485 );
not NOT1_3322 ( P3_U5131 , P3_U3188 );
nand NAND2_3323 ( P3_U5132 , P3_U2489 , P3_U3188 );
nand NAND2_3324 ( P3_U5133 , P3_U5129 , P3_U5132 );
nand NAND2_3325 ( P3_U5134 , P3_STATE2_REG_3_ , P3_U3186 );
nand NAND2_3326 ( P3_U5135 , P3_U3528 , P3_U5133 );
nand NAND2_3327 ( P3_U5136 , P3_U5131 , P3_U4322 );
nand NAND2_3328 ( P3_U5137 , P3_U2489 , P3_U5136 );
nand NAND2_3329 ( P3_U5138 , P3_U5127 , P3_U2445 );
nand NAND2_3330 ( P3_U5139 , P3_U2505 , P3_U2436 );
nand NAND2_3331 ( P3_U5140 , P3_U5126 , P3_U2435 );
nand NAND2_3332 ( P3_U5141 , P3_U2369 , P3_U2420 );
nand NAND2_3333 ( P3_U5142 , P3_INSTQUEUE_REG_6__7_ , P3_U5135 );
nand NAND2_3334 ( P3_U5143 , P3_U5127 , P3_U2443 );
nand NAND2_3335 ( P3_U5144 , P3_U2505 , P3_U2434 );
nand NAND2_3336 ( P3_U5145 , P3_U5126 , P3_U2433 );
nand NAND2_3337 ( P3_U5146 , P3_U2369 , P3_U2419 );
nand NAND2_3338 ( P3_U5147 , P3_INSTQUEUE_REG_6__6_ , P3_U5135 );
nand NAND2_3339 ( P3_U5148 , P3_U5127 , P3_U2442 );
nand NAND2_3340 ( P3_U5149 , P3_U2505 , P3_U2432 );
nand NAND2_3341 ( P3_U5150 , P3_U5126 , P3_U2431 );
nand NAND2_3342 ( P3_U5151 , P3_U2369 , P3_U2418 );
nand NAND2_3343 ( P3_U5152 , P3_INSTQUEUE_REG_6__5_ , P3_U5135 );
nand NAND2_3344 ( P3_U5153 , P3_U5127 , P3_U2441 );
nand NAND2_3345 ( P3_U5154 , P3_U2505 , P3_U2430 );
nand NAND2_3346 ( P3_U5155 , P3_U5126 , P3_U2429 );
nand NAND2_3347 ( P3_U5156 , P3_U2369 , P3_U2417 );
nand NAND2_3348 ( P3_U5157 , P3_INSTQUEUE_REG_6__4_ , P3_U5135 );
nand NAND2_3349 ( P3_U5158 , P3_U5127 , P3_U2440 );
nand NAND2_3350 ( P3_U5159 , P3_U2505 , P3_U2428 );
nand NAND2_3351 ( P3_U5160 , P3_U5126 , P3_U2427 );
nand NAND2_3352 ( P3_U5161 , P3_U2369 , P3_U2416 );
nand NAND2_3353 ( P3_U5162 , P3_INSTQUEUE_REG_6__3_ , P3_U5135 );
nand NAND2_3354 ( P3_U5163 , P3_U5127 , P3_U2439 );
nand NAND2_3355 ( P3_U5164 , P3_U2505 , P3_U2426 );
nand NAND2_3356 ( P3_U5165 , P3_U5126 , P3_U2425 );
nand NAND2_3357 ( P3_U5166 , P3_U2369 , P3_U2415 );
nand NAND2_3358 ( P3_U5167 , P3_INSTQUEUE_REG_6__2_ , P3_U5135 );
nand NAND2_3359 ( P3_U5168 , P3_U5127 , P3_U2438 );
nand NAND2_3360 ( P3_U5169 , P3_U2505 , P3_U2424 );
nand NAND2_3361 ( P3_U5170 , P3_U5126 , P3_U2423 );
nand NAND2_3362 ( P3_U5171 , P3_U2369 , P3_U2414 );
nand NAND2_3363 ( P3_U5172 , P3_INSTQUEUE_REG_6__1_ , P3_U5135 );
nand NAND2_3364 ( P3_U5173 , P3_U5127 , P3_U2437 );
nand NAND2_3365 ( P3_U5174 , P3_U2505 , P3_U2422 );
nand NAND2_3366 ( P3_U5175 , P3_U5126 , P3_U2421 );
nand NAND2_3367 ( P3_U5176 , P3_U2369 , P3_U2413 );
nand NAND2_3368 ( P3_U5177 , P3_INSTQUEUE_REG_6__0_ , P3_U5135 );
not NOT1_3369 ( P3_U5178 , P3_U3191 );
not NOT1_3370 ( P3_U5179 , P3_U3190 );
nand NAND2_3371 ( P3_U5180 , P3_U4343 , P3_U2458 );
not NOT1_3372 ( P3_U5181 , P3_U3193 );
nand NAND2_3373 ( P3_U5182 , P3_U4645 , P3_U2485 );
not NOT1_3374 ( P3_U5183 , P3_U3192 );
nand NAND2_3375 ( P3_U5184 , P3_U2489 , P3_U3192 );
nand NAND2_3376 ( P3_U5185 , P3_U5181 , P3_U5184 );
nand NAND2_3377 ( P3_U5186 , P3_STATE2_REG_3_ , P3_U3190 );
nand NAND2_3378 ( P3_U5187 , P3_U3546 , P3_U5185 );
nand NAND2_3379 ( P3_U5188 , P3_U5183 , P3_U4322 );
nand NAND2_3380 ( P3_U5189 , P3_U2489 , P3_U5188 );
nand NAND2_3381 ( P3_U5190 , P3_U5179 , P3_U2445 );
nand NAND2_3382 ( P3_U5191 , P3_U2506 , P3_U2436 );
nand NAND2_3383 ( P3_U5192 , P3_U5178 , P3_U2435 );
nand NAND2_3384 ( P3_U5193 , P3_U2368 , P3_U2420 );
nand NAND2_3385 ( P3_U5194 , P3_INSTQUEUE_REG_5__7_ , P3_U5187 );
nand NAND2_3386 ( P3_U5195 , P3_U5179 , P3_U2443 );
nand NAND2_3387 ( P3_U5196 , P3_U2506 , P3_U2434 );
nand NAND2_3388 ( P3_U5197 , P3_U5178 , P3_U2433 );
nand NAND2_3389 ( P3_U5198 , P3_U2368 , P3_U2419 );
nand NAND2_3390 ( P3_U5199 , P3_INSTQUEUE_REG_5__6_ , P3_U5187 );
nand NAND2_3391 ( P3_U5200 , P3_U5179 , P3_U2442 );
nand NAND2_3392 ( P3_U5201 , P3_U2506 , P3_U2432 );
nand NAND2_3393 ( P3_U5202 , P3_U5178 , P3_U2431 );
nand NAND2_3394 ( P3_U5203 , P3_U2368 , P3_U2418 );
nand NAND2_3395 ( P3_U5204 , P3_INSTQUEUE_REG_5__5_ , P3_U5187 );
nand NAND2_3396 ( P3_U5205 , P3_U5179 , P3_U2441 );
nand NAND2_3397 ( P3_U5206 , P3_U2506 , P3_U2430 );
nand NAND2_3398 ( P3_U5207 , P3_U5178 , P3_U2429 );
nand NAND2_3399 ( P3_U5208 , P3_U2368 , P3_U2417 );
nand NAND2_3400 ( P3_U5209 , P3_INSTQUEUE_REG_5__4_ , P3_U5187 );
nand NAND2_3401 ( P3_U5210 , P3_U5179 , P3_U2440 );
nand NAND2_3402 ( P3_U5211 , P3_U2506 , P3_U2428 );
nand NAND2_3403 ( P3_U5212 , P3_U5178 , P3_U2427 );
nand NAND2_3404 ( P3_U5213 , P3_U2368 , P3_U2416 );
nand NAND2_3405 ( P3_U5214 , P3_INSTQUEUE_REG_5__3_ , P3_U5187 );
nand NAND2_3406 ( P3_U5215 , P3_U5179 , P3_U2439 );
nand NAND2_3407 ( P3_U5216 , P3_U2506 , P3_U2426 );
nand NAND2_3408 ( P3_U5217 , P3_U5178 , P3_U2425 );
nand NAND2_3409 ( P3_U5218 , P3_U2368 , P3_U2415 );
nand NAND2_3410 ( P3_U5219 , P3_INSTQUEUE_REG_5__2_ , P3_U5187 );
nand NAND2_3411 ( P3_U5220 , P3_U5179 , P3_U2438 );
nand NAND2_3412 ( P3_U5221 , P3_U2506 , P3_U2424 );
nand NAND2_3413 ( P3_U5222 , P3_U5178 , P3_U2423 );
nand NAND2_3414 ( P3_U5223 , P3_U2368 , P3_U2414 );
nand NAND2_3415 ( P3_U5224 , P3_INSTQUEUE_REG_5__1_ , P3_U5187 );
nand NAND2_3416 ( P3_U5225 , P3_U5179 , P3_U2437 );
nand NAND2_3417 ( P3_U5226 , P3_U2506 , P3_U2422 );
nand NAND2_3418 ( P3_U5227 , P3_U5178 , P3_U2421 );
nand NAND2_3419 ( P3_U5228 , P3_U2368 , P3_U2413 );
nand NAND2_3420 ( P3_U5229 , P3_INSTQUEUE_REG_5__0_ , P3_U5187 );
not NOT1_3421 ( P3_U5230 , P3_U3195 );
not NOT1_3422 ( P3_U5231 , P3_U3194 );
not NOT1_3423 ( P3_U5232 , P3_U3072 );
nand NAND2_3424 ( P3_U5233 , P3_U2496 , P3_U2485 );
nand NAND2_3425 ( P3_U5234 , P3_U3195 , P3_U5233 );
nand NAND2_3426 ( P3_U5235 , P3_U2489 , P3_U5234 );
nand NAND2_3427 ( P3_U5236 , P3_U5235 , P3_U3072 );
nand NAND2_3428 ( P3_U5237 , P3_STATE2_REG_3_ , P3_U3194 );
nand NAND2_3429 ( P3_U5238 , P3_U3564 , P3_U5236 );
nand NAND2_3430 ( P3_U5239 , P3_U2489 , P3_U3136 );
nand NAND2_3431 ( P3_U5240 , P3_U5231 , P3_U2445 );
nand NAND2_3432 ( P3_U5241 , P3_U2507 , P3_U2436 );
nand NAND2_3433 ( P3_U5242 , P3_U5230 , P3_U2435 );
nand NAND2_3434 ( P3_U5243 , P3_U2367 , P3_U2420 );
nand NAND2_3435 ( P3_U5244 , P3_INSTQUEUE_REG_4__7_ , P3_U5238 );
nand NAND2_3436 ( P3_U5245 , P3_U5231 , P3_U2443 );
nand NAND2_3437 ( P3_U5246 , P3_U2507 , P3_U2434 );
nand NAND2_3438 ( P3_U5247 , P3_U5230 , P3_U2433 );
nand NAND2_3439 ( P3_U5248 , P3_U2367 , P3_U2419 );
nand NAND2_3440 ( P3_U5249 , P3_INSTQUEUE_REG_4__6_ , P3_U5238 );
nand NAND2_3441 ( P3_U5250 , P3_U5231 , P3_U2442 );
nand NAND2_3442 ( P3_U5251 , P3_U2507 , P3_U2432 );
nand NAND2_3443 ( P3_U5252 , P3_U5230 , P3_U2431 );
nand NAND2_3444 ( P3_U5253 , P3_U2367 , P3_U2418 );
nand NAND2_3445 ( P3_U5254 , P3_INSTQUEUE_REG_4__5_ , P3_U5238 );
nand NAND2_3446 ( P3_U5255 , P3_U5231 , P3_U2441 );
nand NAND2_3447 ( P3_U5256 , P3_U2507 , P3_U2430 );
nand NAND2_3448 ( P3_U5257 , P3_U5230 , P3_U2429 );
nand NAND2_3449 ( P3_U5258 , P3_U2367 , P3_U2417 );
nand NAND2_3450 ( P3_U5259 , P3_INSTQUEUE_REG_4__4_ , P3_U5238 );
nand NAND2_3451 ( P3_U5260 , P3_U5231 , P3_U2440 );
nand NAND2_3452 ( P3_U5261 , P3_U2507 , P3_U2428 );
nand NAND2_3453 ( P3_U5262 , P3_U5230 , P3_U2427 );
nand NAND2_3454 ( P3_U5263 , P3_U2367 , P3_U2416 );
nand NAND2_3455 ( P3_U5264 , P3_INSTQUEUE_REG_4__3_ , P3_U5238 );
nand NAND2_3456 ( P3_U5265 , P3_U5231 , P3_U2439 );
nand NAND2_3457 ( P3_U5266 , P3_U2507 , P3_U2426 );
nand NAND2_3458 ( P3_U5267 , P3_U5230 , P3_U2425 );
nand NAND2_3459 ( P3_U5268 , P3_U2367 , P3_U2415 );
nand NAND2_3460 ( P3_U5269 , P3_INSTQUEUE_REG_4__2_ , P3_U5238 );
nand NAND2_3461 ( P3_U5270 , P3_U5231 , P3_U2438 );
nand NAND2_3462 ( P3_U5271 , P3_U2507 , P3_U2424 );
nand NAND2_3463 ( P3_U5272 , P3_U5230 , P3_U2423 );
nand NAND2_3464 ( P3_U5273 , P3_U2367 , P3_U2414 );
nand NAND2_3465 ( P3_U5274 , P3_INSTQUEUE_REG_4__1_ , P3_U5238 );
nand NAND2_3466 ( P3_U5275 , P3_U5231 , P3_U2437 );
nand NAND2_3467 ( P3_U5276 , P3_U2507 , P3_U2422 );
nand NAND2_3468 ( P3_U5277 , P3_U5230 , P3_U2421 );
nand NAND2_3469 ( P3_U5278 , P3_U2367 , P3_U2413 );
nand NAND2_3470 ( P3_U5279 , P3_INSTQUEUE_REG_4__0_ , P3_U5238 );
not NOT1_3471 ( P3_U5280 , P3_U3197 );
not NOT1_3472 ( P3_U5281 , P3_U3196 );
nand NAND2_3473 ( P3_U5282 , P3_U2460 , P3_U4653 );
not NOT1_3474 ( P3_U5283 , P3_U3198 );
nand NAND2_3475 ( P3_U5284 , P3_U2509 , P3_U4657 );
nand NAND2_3476 ( P3_U5285 , P3_U3197 , P3_U5284 );
nand NAND2_3477 ( P3_U5286 , P3_U2489 , P3_U5285 );
nand NAND2_3478 ( P3_U5287 , P3_U5283 , P3_U5286 );
nand NAND2_3479 ( P3_U5288 , P3_STATE2_REG_3_ , P3_U3196 );
nand NAND2_3480 ( P3_U5289 , P3_U3582 , P3_U5287 );
nand NAND2_3481 ( P3_U5290 , P3_U2489 , P3_U3136 );
nand NAND2_3482 ( P3_U5291 , P3_U5281 , P3_U2445 );
nand NAND2_3483 ( P3_U5292 , P3_U2510 , P3_U2436 );
nand NAND2_3484 ( P3_U5293 , P3_U5280 , P3_U2435 );
nand NAND2_3485 ( P3_U5294 , P3_U2366 , P3_U2420 );
nand NAND2_3486 ( P3_U5295 , P3_INSTQUEUE_REG_3__7_ , P3_U5289 );
nand NAND2_3487 ( P3_U5296 , P3_U5281 , P3_U2443 );
nand NAND2_3488 ( P3_U5297 , P3_U2510 , P3_U2434 );
nand NAND2_3489 ( P3_U5298 , P3_U5280 , P3_U2433 );
nand NAND2_3490 ( P3_U5299 , P3_U2366 , P3_U2419 );
nand NAND2_3491 ( P3_U5300 , P3_INSTQUEUE_REG_3__6_ , P3_U5289 );
nand NAND2_3492 ( P3_U5301 , P3_U5281 , P3_U2442 );
nand NAND2_3493 ( P3_U5302 , P3_U2510 , P3_U2432 );
nand NAND2_3494 ( P3_U5303 , P3_U5280 , P3_U2431 );
nand NAND2_3495 ( P3_U5304 , P3_U2366 , P3_U2418 );
nand NAND2_3496 ( P3_U5305 , P3_INSTQUEUE_REG_3__5_ , P3_U5289 );
nand NAND2_3497 ( P3_U5306 , P3_U5281 , P3_U2441 );
nand NAND2_3498 ( P3_U5307 , P3_U2510 , P3_U2430 );
nand NAND2_3499 ( P3_U5308 , P3_U5280 , P3_U2429 );
nand NAND2_3500 ( P3_U5309 , P3_U2366 , P3_U2417 );
nand NAND2_3501 ( P3_U5310 , P3_INSTQUEUE_REG_3__4_ , P3_U5289 );
nand NAND2_3502 ( P3_U5311 , P3_U5281 , P3_U2440 );
nand NAND2_3503 ( P3_U5312 , P3_U2510 , P3_U2428 );
nand NAND2_3504 ( P3_U5313 , P3_U5280 , P3_U2427 );
nand NAND2_3505 ( P3_U5314 , P3_U2366 , P3_U2416 );
nand NAND2_3506 ( P3_U5315 , P3_INSTQUEUE_REG_3__3_ , P3_U5289 );
nand NAND2_3507 ( P3_U5316 , P3_U5281 , P3_U2439 );
nand NAND2_3508 ( P3_U5317 , P3_U2510 , P3_U2426 );
nand NAND2_3509 ( P3_U5318 , P3_U5280 , P3_U2425 );
nand NAND2_3510 ( P3_U5319 , P3_U2366 , P3_U2415 );
nand NAND2_3511 ( P3_U5320 , P3_INSTQUEUE_REG_3__2_ , P3_U5289 );
nand NAND2_3512 ( P3_U5321 , P3_U5281 , P3_U2438 );
nand NAND2_3513 ( P3_U5322 , P3_U2510 , P3_U2424 );
nand NAND2_3514 ( P3_U5323 , P3_U5280 , P3_U2423 );
nand NAND2_3515 ( P3_U5324 , P3_U2366 , P3_U2414 );
nand NAND2_3516 ( P3_U5325 , P3_INSTQUEUE_REG_3__1_ , P3_U5289 );
nand NAND2_3517 ( P3_U5326 , P3_U5281 , P3_U2437 );
nand NAND2_3518 ( P3_U5327 , P3_U2510 , P3_U2422 );
nand NAND2_3519 ( P3_U5328 , P3_U5280 , P3_U2421 );
nand NAND2_3520 ( P3_U5329 , P3_U2366 , P3_U2413 );
nand NAND2_3521 ( P3_U5330 , P3_INSTQUEUE_REG_3__0_ , P3_U5289 );
not NOT1_3522 ( P3_U5331 , P3_U3200 );
not NOT1_3523 ( P3_U5332 , P3_U3199 );
nand NAND2_3524 ( P3_U5333 , P3_U2460 , P3_U4342 );
not NOT1_3525 ( P3_U5334 , P3_U3201 );
nand NAND2_3526 ( P3_U5335 , P3_U2509 , P3_U4644 );
nand NAND2_3527 ( P3_U5336 , P3_U3200 , P3_U5335 );
nand NAND2_3528 ( P3_U5337 , P3_U2489 , P3_U5336 );
nand NAND2_3529 ( P3_U5338 , P3_U5334 , P3_U5337 );
nand NAND2_3530 ( P3_U5339 , P3_STATE2_REG_3_ , P3_U3199 );
nand NAND2_3531 ( P3_U5340 , P3_U3599 , P3_U5338 );
nand NAND2_3532 ( P3_U5341 , P3_U2489 , P3_U3136 );
nand NAND2_3533 ( P3_U5342 , P3_U5332 , P3_U2445 );
nand NAND2_3534 ( P3_U5343 , P3_U2511 , P3_U2436 );
nand NAND2_3535 ( P3_U5344 , P3_U5331 , P3_U2435 );
nand NAND2_3536 ( P3_U5345 , P3_U2365 , P3_U2420 );
nand NAND2_3537 ( P3_U5346 , P3_INSTQUEUE_REG_2__7_ , P3_U5340 );
nand NAND2_3538 ( P3_U5347 , P3_U5332 , P3_U2443 );
nand NAND2_3539 ( P3_U5348 , P3_U2511 , P3_U2434 );
nand NAND2_3540 ( P3_U5349 , P3_U5331 , P3_U2433 );
nand NAND2_3541 ( P3_U5350 , P3_U2365 , P3_U2419 );
nand NAND2_3542 ( P3_U5351 , P3_INSTQUEUE_REG_2__6_ , P3_U5340 );
nand NAND2_3543 ( P3_U5352 , P3_U5332 , P3_U2442 );
nand NAND2_3544 ( P3_U5353 , P3_U2511 , P3_U2432 );
nand NAND2_3545 ( P3_U5354 , P3_U5331 , P3_U2431 );
nand NAND2_3546 ( P3_U5355 , P3_U2365 , P3_U2418 );
nand NAND2_3547 ( P3_U5356 , P3_INSTQUEUE_REG_2__5_ , P3_U5340 );
nand NAND2_3548 ( P3_U5357 , P3_U5332 , P3_U2441 );
nand NAND2_3549 ( P3_U5358 , P3_U2511 , P3_U2430 );
nand NAND2_3550 ( P3_U5359 , P3_U5331 , P3_U2429 );
nand NAND2_3551 ( P3_U5360 , P3_U2365 , P3_U2417 );
nand NAND2_3552 ( P3_U5361 , P3_INSTQUEUE_REG_2__4_ , P3_U5340 );
nand NAND2_3553 ( P3_U5362 , P3_U5332 , P3_U2440 );
nand NAND2_3554 ( P3_U5363 , P3_U2511 , P3_U2428 );
nand NAND2_3555 ( P3_U5364 , P3_U5331 , P3_U2427 );
nand NAND2_3556 ( P3_U5365 , P3_U2365 , P3_U2416 );
nand NAND2_3557 ( P3_U5366 , P3_INSTQUEUE_REG_2__3_ , P3_U5340 );
nand NAND2_3558 ( P3_U5367 , P3_U5332 , P3_U2439 );
nand NAND2_3559 ( P3_U5368 , P3_U2511 , P3_U2426 );
nand NAND2_3560 ( P3_U5369 , P3_U5331 , P3_U2425 );
nand NAND2_3561 ( P3_U5370 , P3_U2365 , P3_U2415 );
nand NAND2_3562 ( P3_U5371 , P3_INSTQUEUE_REG_2__2_ , P3_U5340 );
nand NAND2_3563 ( P3_U5372 , P3_U5332 , P3_U2438 );
nand NAND2_3564 ( P3_U5373 , P3_U2511 , P3_U2424 );
nand NAND2_3565 ( P3_U5374 , P3_U5331 , P3_U2423 );
nand NAND2_3566 ( P3_U5375 , P3_U2365 , P3_U2414 );
nand NAND2_3567 ( P3_U5376 , P3_INSTQUEUE_REG_2__1_ , P3_U5340 );
nand NAND2_3568 ( P3_U5377 , P3_U5332 , P3_U2437 );
nand NAND2_3569 ( P3_U5378 , P3_U2511 , P3_U2422 );
nand NAND2_3570 ( P3_U5379 , P3_U5331 , P3_U2421 );
nand NAND2_3571 ( P3_U5380 , P3_U2365 , P3_U2413 );
nand NAND2_3572 ( P3_U5381 , P3_INSTQUEUE_REG_2__0_ , P3_U5340 );
not NOT1_3573 ( P3_U5382 , P3_U3203 );
not NOT1_3574 ( P3_U5383 , P3_U3202 );
nand NAND2_3575 ( P3_U5384 , P3_U2460 , P3_U4343 );
not NOT1_3576 ( P3_U5385 , P3_U3204 );
nand NAND2_3577 ( P3_U5386 , P3_U2509 , P3_U4645 );
nand NAND2_3578 ( P3_U5387 , P3_U3203 , P3_U5386 );
nand NAND2_3579 ( P3_U5388 , P3_U2489 , P3_U5387 );
nand NAND2_3580 ( P3_U5389 , P3_U5385 , P3_U5388 );
nand NAND2_3581 ( P3_U5390 , P3_STATE2_REG_3_ , P3_U3202 );
nand NAND2_3582 ( P3_U5391 , P3_U3617 , P3_U5389 );
nand NAND2_3583 ( P3_U5392 , P3_U2489 , P3_U3136 );
nand NAND2_3584 ( P3_U5393 , P3_U5383 , P3_U2445 );
nand NAND2_3585 ( P3_U5394 , P3_U2512 , P3_U2436 );
nand NAND2_3586 ( P3_U5395 , P3_U5382 , P3_U2435 );
nand NAND2_3587 ( P3_U5396 , P3_U2364 , P3_U2420 );
nand NAND2_3588 ( P3_U5397 , P3_INSTQUEUE_REG_1__7_ , P3_U5391 );
nand NAND2_3589 ( P3_U5398 , P3_U5383 , P3_U2443 );
nand NAND2_3590 ( P3_U5399 , P3_U2512 , P3_U2434 );
nand NAND2_3591 ( P3_U5400 , P3_U5382 , P3_U2433 );
nand NAND2_3592 ( P3_U5401 , P3_U2364 , P3_U2419 );
nand NAND2_3593 ( P3_U5402 , P3_INSTQUEUE_REG_1__6_ , P3_U5391 );
nand NAND2_3594 ( P3_U5403 , P3_U5383 , P3_U2442 );
nand NAND2_3595 ( P3_U5404 , P3_U2512 , P3_U2432 );
nand NAND2_3596 ( P3_U5405 , P3_U5382 , P3_U2431 );
nand NAND2_3597 ( P3_U5406 , P3_U2364 , P3_U2418 );
nand NAND2_3598 ( P3_U5407 , P3_INSTQUEUE_REG_1__5_ , P3_U5391 );
nand NAND2_3599 ( P3_U5408 , P3_U5383 , P3_U2441 );
nand NAND2_3600 ( P3_U5409 , P3_U2512 , P3_U2430 );
nand NAND2_3601 ( P3_U5410 , P3_U5382 , P3_U2429 );
nand NAND2_3602 ( P3_U5411 , P3_U2364 , P3_U2417 );
nand NAND2_3603 ( P3_U5412 , P3_INSTQUEUE_REG_1__4_ , P3_U5391 );
nand NAND2_3604 ( P3_U5413 , P3_U5383 , P3_U2440 );
nand NAND2_3605 ( P3_U5414 , P3_U2512 , P3_U2428 );
nand NAND2_3606 ( P3_U5415 , P3_U5382 , P3_U2427 );
nand NAND2_3607 ( P3_U5416 , P3_U2364 , P3_U2416 );
nand NAND2_3608 ( P3_U5417 , P3_INSTQUEUE_REG_1__3_ , P3_U5391 );
nand NAND2_3609 ( P3_U5418 , P3_U5383 , P3_U2439 );
nand NAND2_3610 ( P3_U5419 , P3_U2512 , P3_U2426 );
nand NAND2_3611 ( P3_U5420 , P3_U5382 , P3_U2425 );
nand NAND2_3612 ( P3_U5421 , P3_U2364 , P3_U2415 );
nand NAND2_3613 ( P3_U5422 , P3_INSTQUEUE_REG_1__2_ , P3_U5391 );
nand NAND2_3614 ( P3_U5423 , P3_U5383 , P3_U2438 );
nand NAND2_3615 ( P3_U5424 , P3_U2512 , P3_U2424 );
nand NAND2_3616 ( P3_U5425 , P3_U5382 , P3_U2423 );
nand NAND2_3617 ( P3_U5426 , P3_U2364 , P3_U2414 );
nand NAND2_3618 ( P3_U5427 , P3_INSTQUEUE_REG_1__1_ , P3_U5391 );
nand NAND2_3619 ( P3_U5428 , P3_U5383 , P3_U2437 );
nand NAND2_3620 ( P3_U5429 , P3_U2512 , P3_U2422 );
nand NAND2_3621 ( P3_U5430 , P3_U5382 , P3_U2421 );
nand NAND2_3622 ( P3_U5431 , P3_U2364 , P3_U2413 );
nand NAND2_3623 ( P3_U5432 , P3_INSTQUEUE_REG_1__0_ , P3_U5391 );
not NOT1_3624 ( P3_U5433 , P3_U3206 );
not NOT1_3625 ( P3_U5434 , P3_U3205 );
not NOT1_3626 ( P3_U5435 , P3_U3073 );
nand NAND2_3627 ( P3_U5436 , P3_U2509 , P3_U2496 );
nand NAND2_3628 ( P3_U5437 , P3_U3206 , P3_U5436 );
nand NAND2_3629 ( P3_U5438 , P3_U2489 , P3_U5437 );
nand NAND2_3630 ( P3_U5439 , P3_U5438 , P3_U3073 );
nand NAND2_3631 ( P3_U5440 , P3_STATE2_REG_3_ , P3_U3205 );
nand NAND2_3632 ( P3_U5441 , P3_U3635 , P3_U5439 );
nand NAND2_3633 ( P3_U5442 , P3_U2489 , P3_U3136 );
nand NAND2_3634 ( P3_U5443 , P3_U5434 , P3_U2445 );
nand NAND2_3635 ( P3_U5444 , P3_U2513 , P3_U2436 );
nand NAND2_3636 ( P3_U5445 , P3_U5433 , P3_U2435 );
nand NAND2_3637 ( P3_U5446 , P3_U2363 , P3_U2420 );
nand NAND2_3638 ( P3_U5447 , P3_INSTQUEUE_REG_0__7_ , P3_U5441 );
nand NAND2_3639 ( P3_U5448 , P3_U5434 , P3_U2443 );
nand NAND2_3640 ( P3_U5449 , P3_U2513 , P3_U2434 );
nand NAND2_3641 ( P3_U5450 , P3_U5433 , P3_U2433 );
nand NAND2_3642 ( P3_U5451 , P3_U2363 , P3_U2419 );
nand NAND2_3643 ( P3_U5452 , P3_INSTQUEUE_REG_0__6_ , P3_U5441 );
nand NAND2_3644 ( P3_U5453 , P3_U5434 , P3_U2442 );
nand NAND2_3645 ( P3_U5454 , P3_U2513 , P3_U2432 );
nand NAND2_3646 ( P3_U5455 , P3_U5433 , P3_U2431 );
nand NAND2_3647 ( P3_U5456 , P3_U2363 , P3_U2418 );
nand NAND2_3648 ( P3_U5457 , P3_INSTQUEUE_REG_0__5_ , P3_U5441 );
nand NAND2_3649 ( P3_U5458 , P3_U5434 , P3_U2441 );
nand NAND2_3650 ( P3_U5459 , P3_U2513 , P3_U2430 );
nand NAND2_3651 ( P3_U5460 , P3_U5433 , P3_U2429 );
nand NAND2_3652 ( P3_U5461 , P3_U2363 , P3_U2417 );
nand NAND2_3653 ( P3_U5462 , P3_INSTQUEUE_REG_0__4_ , P3_U5441 );
nand NAND2_3654 ( P3_U5463 , P3_U5434 , P3_U2440 );
nand NAND2_3655 ( P3_U5464 , P3_U2513 , P3_U2428 );
nand NAND2_3656 ( P3_U5465 , P3_U5433 , P3_U2427 );
nand NAND2_3657 ( P3_U5466 , P3_U2363 , P3_U2416 );
nand NAND2_3658 ( P3_U5467 , P3_INSTQUEUE_REG_0__3_ , P3_U5441 );
nand NAND2_3659 ( P3_U5468 , P3_U5434 , P3_U2439 );
nand NAND2_3660 ( P3_U5469 , P3_U2513 , P3_U2426 );
nand NAND2_3661 ( P3_U5470 , P3_U5433 , P3_U2425 );
nand NAND2_3662 ( P3_U5471 , P3_U2363 , P3_U2415 );
nand NAND2_3663 ( P3_U5472 , P3_INSTQUEUE_REG_0__2_ , P3_U5441 );
nand NAND2_3664 ( P3_U5473 , P3_U5434 , P3_U2438 );
nand NAND2_3665 ( P3_U5474 , P3_U2513 , P3_U2424 );
nand NAND2_3666 ( P3_U5475 , P3_U5433 , P3_U2423 );
nand NAND2_3667 ( P3_U5476 , P3_U2363 , P3_U2414 );
nand NAND2_3668 ( P3_U5477 , P3_INSTQUEUE_REG_0__1_ , P3_U5441 );
nand NAND2_3669 ( P3_U5478 , P3_U5434 , P3_U2437 );
nand NAND2_3670 ( P3_U5479 , P3_U2513 , P3_U2422 );
nand NAND2_3671 ( P3_U5480 , P3_U5433 , P3_U2421 );
nand NAND2_3672 ( P3_U5481 , P3_U2363 , P3_U2413 );
nand NAND2_3673 ( P3_U5482 , P3_INSTQUEUE_REG_0__0_ , P3_U5441 );
nand NAND4_3674 ( P3_U5483 , P3_U7917 , P3_U2514 , P3_U3655 , P3_U4339 );
not NOT1_3675 ( P3_U5484 , P3_U3209 );
nand NAND2_3676 ( P3_U5485 , P3_U4296 , P3_U3209 );
nand NAND2_3677 ( P3_U5486 , P3_GTE_450_U6 , P3_U4303 );
nand NAND2_3678 ( P3_U5487 , P3_GTE_504_U6 , P3_U4302 );
not NOT1_3679 ( P3_U5488 , P3_U3255 );
nand NAND2_3680 ( P3_U5489 , P3_GTE_412_U6 , P3_U4304 );
nand NAND2_3681 ( P3_U5490 , P3_GTE_485_U6 , P3_U2356 );
not NOT1_3682 ( P3_U5491 , P3_U3254 );
nand NAND2_3683 ( P3_U5492 , P3_U3254 , P3_U2630 );
nand NAND2_3684 ( P3_U5493 , P3_GTE_390_U6 , P3_U2357 );
nand NAND2_3685 ( P3_U5494 , P3_U4294 , P3_U3255 );
nand NAND2_3686 ( P3_U5495 , P3_GTE_401_U6 , P3_U4305 );
not NOT1_3687 ( P3_U5496 , P3_U4290 );
nand NAND2_3688 ( P3_U5497 , P3_U2390 , P3_U4290 );
nand NAND2_3689 ( P3_U5498 , P3_STATE2_REG_3_ , P3_U3121 );
not NOT1_3690 ( P3_U5499 , P3_U4283 );
nand NAND2_3691 ( P3_U5500 , P3_U3095 , P3_U3097 );
nand NAND2_3692 ( P3_U5501 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_U5500 );
nand NAND2_3693 ( P3_U5502 , P3_U2481 , P3_U3095 );
nand NAND2_3694 ( P3_U5503 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_3695 ( P3_U5504 , P3_U3223 );
nand NAND2_3696 ( P3_U5505 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_U4332 );
not NOT1_3697 ( P3_U5506 , P3_U3224 );
nand NAND2_3698 ( P3_U5507 , P3_U5484 , P3_U3107 );
nand NAND3_3699 ( P3_U5508 , P3_U4522 , P3_U4607 , P3_U4488 );
nand NAND2_3700 ( P3_U5509 , P3_U4296 , P3_U5507 );
nand NAND3_3701 ( P3_U5510 , P3_U7974 , P3_U7973 , P3_U3104 );
nand NAND2_3702 ( P3_U5511 , P3_U4323 , P3_U4344 );
nand NAND2_3703 ( P3_U5512 , P3_U5509 , P3_U3665 );
nand NAND2_3704 ( P3_U5513 , P3_U4522 , P3_U4607 );
nand NAND2_3705 ( P3_U5514 , P3_U4607 , P3_U3218 );
nand NAND3_3706 ( P3_U5515 , P3_U5514 , P3_U3216 , P3_U4556 );
nand NAND2_3707 ( P3_U5516 , P3_U4573 , P3_U4505 );
nand NAND2_3708 ( P3_U5517 , P3_U4488 , P3_U5516 );
nand NAND3_3709 ( P3_U5518 , P3_U3103 , P3_U3218 , P3_U3112 );
nand NAND3_3710 ( P3_U5519 , P3_U4607 , P3_U3104 , P3_U4573 );
nand NAND2_3711 ( P3_U5520 , P3_U4324 , P3_U3103 );
nand NAND2_3712 ( P3_U5521 , P3_U5518 , P3_U3102 );
not NOT1_3713 ( P3_U5522 , P3_U3220 );
nand NAND2_3714 ( P3_U5523 , P3_U3111 , P3_U3114 );
nand NAND2_3715 ( P3_U5524 , P3_U2452 , P3_U3108 );
not NOT1_3716 ( P3_U5525 , P3_U3221 );
nand NAND2_3717 ( P3_U5526 , P3_U2462 , P3_U3104 );
nand NAND2_3718 ( P3_U5527 , P3_U3229 , P3_U3219 );
nand NAND2_3719 ( P3_U5528 , P3_U2456 , P3_U5527 );
nand NAND2_3720 ( P3_U5529 , P3_U2518 , P3_U3217 );
nand NAND2_3721 ( P3_U5530 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_U5529 );
nand NAND2_3722 ( P3_U5531 , P3_U5525 , P3_U5530 );
nand NAND3_3723 ( P3_U5532 , P3_U2461 , P3_U5523 , P3_U2450 );
nand NAND2_3724 ( P3_U5533 , P3_U3673 , P3_U7918 );
not NOT1_3725 ( P3_U5534 , P3_U3226 );
nand NAND2_3726 ( P3_U5535 , P3_U3672 , P3_U5522 );
nand NAND3_3727 ( P3_U5536 , P3_U3659 , P3_U5523 , P3_U2451 );
nand NAND2_3728 ( P3_U5537 , P3_U3669 , P3_U5531 );
nand NAND2_3729 ( P3_U5538 , P3_U3670 , P3_U3220 );
nand NAND2_3730 ( P3_U5539 , P3_U5504 , P3_U5535 );
nand NAND2_3731 ( P3_U5540 , P3_U5506 , P3_U3226 );
nand NAND2_3732 ( P3_U5541 , P3_ADD_495_U9 , P3_U2356 );
nand NAND2_3733 ( P3_U5542 , P3_U5537 , P3_U3676 );
not NOT1_3734 ( P3_U5543 , P3_U3265 );
nand NAND2_3735 ( P3_U5544 , P3_U4345 , P3_U3265 );
nand NAND2_3736 ( P3_U5545 , P3_U4340 , P3_U5542 );
nand NAND2_3737 ( P3_U5546 , P3_U5545 , P3_U5544 );
not NOT1_3738 ( P3_U5547 , P3_U3227 );
not NOT1_3739 ( P3_U5548 , P3_U3225 );
nand NAND2_3740 ( P3_U5549 , P3_U5534 , P3_U5522 );
nand NAND3_3741 ( P3_U5550 , P3_U5548 , P3_U5523 , P3_U2451 );
nand NAND2_3742 ( P3_U5551 , P3_U5547 , P3_U5549 );
nand NAND2_3743 ( P3_U5552 , P3_ADD_495_U10 , P3_U2356 );
nand NAND3_3744 ( P3_U5553 , P3_U7982 , P3_U7981 , P3_U3679 );
nand NAND3_3745 ( P3_U5554 , P3_STATE2_REG_1_ , P3_U3286 , P3_U3287 );
nand NAND2_3746 ( P3_U5555 , P3_U4345 , P3_U3225 );
nand NAND2_3747 ( P3_U5556 , P3_U4340 , P3_U5553 );
nand NAND2_3748 ( P3_U5557 , P3_U3680 , P3_U5556 );
not NOT1_3749 ( P3_U5558 , P3_U3228 );
nand NAND2_3750 ( P3_U5559 , P3_U4341 , P3_U4608 );
not NOT1_3751 ( P3_U5560 , P3_U3231 );
not NOT1_3752 ( P3_U5561 , P3_U3230 );
nand NAND2_3753 ( P3_U5562 , P3_U2466 , P3_U3230 );
nand NAND2_3754 ( P3_U5563 , P3_U5531 , P3_U3094 );
nand NAND2_3755 ( P3_U5564 , P3_U5558 , P3_U3231 );
nand NAND2_3756 ( P3_U5565 , P3_ADD_495_U4 , P3_U2356 );
nand NAND2_3757 ( P3_U5566 , P3_U5563 , P3_U3681 );
nand NAND3_3758 ( P3_U5567 , P3_STATE2_REG_1_ , P3_U3286 , P3_U7985 );
nand NAND2_3759 ( P3_U5568 , P3_U5558 , P3_U4345 );
nand NAND2_3760 ( P3_U5569 , P3_U4340 , P3_U5566 );
nand NAND2_3761 ( P3_U5570 , P3_U3683 , P3_U5569 );
nand NAND2_3762 ( P3_U5571 , P3_U5560 , P3_U5561 );
nand NAND2_3763 ( P3_U5572 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_U2356 );
nand NAND3_3764 ( P3_U5573 , P3_U7994 , P3_U7993 , P3_U5572 );
nand NAND2_3765 ( P3_U5574 , P3_U4345 , P3_U3093 );
nand NAND2_3766 ( P3_U5575 , P3_U4340 , P3_U5573 );
nand NAND2_3767 ( P3_U5576 , P3_U7988 , P3_STATE2_REG_1_ );
nand NAND2_3768 ( P3_U5577 , P3_U3684 , P3_U5575 );
nand NAND3_3769 ( P3_U5578 , P3_U2453 , P3_STATE2_REG_0_ , P3_LT_589_U6 );
not NOT1_3770 ( P3_U5579 , P3_U3233 );
nand NAND2_3771 ( P3_U5580 , P3_STATE2_REG_3_ , P3_U3132 );
nand NAND2_3772 ( P3_U5581 , P3_U3233 , P3_U5580 );
nand NAND2_3773 ( P3_U5582 , P3_U4315 , P3_U3123 );
nand NAND2_3774 ( P3_U5583 , P3_U4647 , P3_U3271 );
nand NAND2_3775 ( P3_U5584 , P3_U3182 , P3_U5583 );
nand NAND2_3776 ( P3_U5585 , P3_U3183 , P3_U5584 );
nand NAND2_3777 ( P3_U5586 , P3_U4322 , P3_U5585 );
nand NAND2_3778 ( P3_U5587 , P3_U5582 , P3_U3142 );
nand NAND2_3779 ( P3_U5588 , P3_U4650 , P3_STATE2_REG_3_ );
nand NAND2_3780 ( P3_U5589 , P3_U3685 , P3_U5586 );
nand NAND2_3781 ( P3_U5590 , P3_U5589 , P3_U3233 );
nand NAND2_3782 ( P3_U5591 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_U5581 );
nand NAND3_3783 ( P3_U5592 , P3_STATE2_REG_3_ , P3_U3131 , P3_U4648 );
nand NAND2_3784 ( P3_U5593 , P3_U4322 , P3_U7999 );
nand NAND2_3785 ( P3_U5594 , P3_U3270 , P3_U5582 );
nand NAND2_3786 ( P3_U5595 , P3_U3686 , P3_U5593 );
nand NAND2_3787 ( P3_U5596 , P3_STATE2_REG_3_ , P3_U3130 );
nand NAND2_3788 ( P3_U5597 , P3_U3233 , P3_U5596 );
nand NAND2_3789 ( P3_U5598 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_U5597 );
nand NAND2_3790 ( P3_U5599 , P3_U5595 , P3_U3233 );
nand NAND2_3791 ( P3_U5600 , P3_U4322 , P3_U3156 );
nand NAND2_3792 ( P3_U5601 , P3_STATE2_REG_3_ , P3_U3129 );
nand NAND2_3793 ( P3_U5602 , P3_U5601 , P3_U5600 );
nand NAND2_3794 ( P3_U5603 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_U5602 );
nand NAND2_3795 ( P3_U5604 , P3_U2493 , P3_U4322 );
nand NAND2_3796 ( P3_U5605 , P3_U5582 , P3_U3141 );
nand NAND3_3797 ( P3_U5606 , P3_U5605 , P3_U5603 , P3_U5604 );
nand NAND2_3798 ( P3_U5607 , P3_STATE2_REG_3_ , P3_U3128 );
nand NAND2_3799 ( P3_U5608 , P3_U3233 , P3_U5607 );
nand NAND2_3800 ( P3_U5609 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_U5608 );
nand NAND2_3801 ( P3_U5610 , P3_U5606 , P3_U3233 );
not NOT1_3802 ( P3_U5611 , P3_U3234 );
nand NAND2_3803 ( P3_U5612 , P3_U5611 , P3_U3233 );
nand NAND2_3804 ( P3_U5613 , P3_STATE2_REG_3_ , P3_U3128 );
nand NAND2_3805 ( P3_U5614 , P3_U4337 , P3_U5613 );
nand NAND2_3806 ( P3_U5615 , P3_U5614 , P3_U3233 );
nand NAND2_3807 ( P3_U5616 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_U5612 );
nand NAND3_3808 ( P3_U5617 , P3_U2463 , P3_U4294 , P3_GTE_450_U6 );
nand NAND2_3809 ( P3_U5618 , P3_GTE_370_U6 , P3_U4344 );
nand NAND2_3810 ( P3_U5619 , P3_U5618 , P3_U5617 );
nand NAND3_3811 ( P3_U5620 , P3_U4590 , P3_U2630 , P3_GTE_412_U6 );
nand NAND2_3812 ( P3_U5621 , P3_GTE_355_U6 , P3_U3074 );
nand NAND2_3813 ( P3_U5622 , P3_U5621 , P3_U5620 );
nand NAND2_3814 ( P3_U5623 , P3_GTE_390_U6 , P3_U4488 );
nand NAND3_3815 ( P3_U5624 , P3_U8001 , P3_U8000 , P3_U5623 );
nand NAND3_3816 ( P3_U5625 , P3_U3102 , P3_U3108 , P3_GTE_401_U6 );
nand NAND2_3817 ( P3_U5626 , P3_U4349 , P3_GTE_504_U6 );
nand NAND2_3818 ( P3_U5627 , P3_U4348 , P3_GTE_485_U6 );
nand NAND2_3819 ( P3_U5628 , P3_U4539 , P3_U5624 );
nand NAND4_3820 ( P3_U5629 , P3_U2515 , P3_U5627 , P3_U3687 , P3_U5628 );
nand NAND2_3821 ( P3_U5630 , P3_U2390 , P3_U5629 );
not NOT1_3822 ( P3_U5631 , P3_U3248 );
nand NAND2_3823 ( P3_U5632 , P3_ADD_360_1242_U85 , P3_U2395 );
nand NAND2_3824 ( P3_U5633 , P3_SUB_357_1258_U69 , P3_U2393 );
nand NAND2_3825 ( P3_U5634 , P3_ADD_558_U5 , P3_U3220 );
nand NAND2_3826 ( P3_U5635 , P3_U4298 , P3_ADD_553_U5 );
nand NAND2_3827 ( P3_U5636 , P3_U4299 , P3_ADD_547_U5 );
nand NAND2_3828 ( P3_U5637 , P3_U4300 , P3_INSTADDRPOINTER_REG_0_ );
nand NAND2_3829 ( P3_U5638 , P3_U4301 , P3_INSTADDRPOINTER_REG_0_ );
nand NAND2_3830 ( P3_U5639 , P3_U2354 , P3_ADD_531_U5 );
nand NAND2_3831 ( P3_U5640 , P3_U2355 , P3_ADD_526_U5 );
nand NAND2_3832 ( P3_U5641 , P3_INSTADDRPOINTER_REG_0_ , P3_U4302 );
nand NAND2_3833 ( P3_U5642 , P3_INSTADDRPOINTER_REG_0_ , P3_U2356 );
nand NAND2_3834 ( P3_U5643 , P3_INSTADDRPOINTER_REG_0_ , P3_U4303 );
nand NAND2_3835 ( P3_U5644 , P3_INSTADDRPOINTER_REG_0_ , P3_U4304 );
nand NAND2_3836 ( P3_U5645 , P3_ADD_405_U4 , P3_U4305 );
nand NAND2_3837 ( P3_U5646 , P3_ADD_394_U4 , P3_U2357 );
nand NAND2_3838 ( P3_U5647 , P3_U2358 , P3_ADD_385_U5 );
nand NAND2_3839 ( P3_U5648 , P3_U2359 , P3_ADD_380_U5 );
nand NAND2_3840 ( P3_U5649 , P3_U4306 , P3_ADD_349_U5 );
nand NAND2_3841 ( P3_U5650 , P3_U2362 , P3_ADD_344_U5 );
nand NAND2_3842 ( P3_U5651 , P3_ADD_371_1212_U87 , P3_U2360 );
nand NAND4_3843 ( P3_U5652 , P3_U3692 , P3_U5634 , P3_U3693 , P3_U3698 );
nand NAND2_3844 ( P3_U5653 , P3_REIP_REG_0_ , P3_U2402 );
nand NAND2_3845 ( P3_U5654 , P3_U4318 , P3_U5652 );
nand NAND2_3846 ( P3_U5655 , P3_U5631 , P3_INSTADDRPOINTER_REG_0_ );
nand NAND2_3847 ( P3_U5656 , P3_ADD_360_1242_U19 , P3_U2395 );
nand NAND2_3848 ( P3_U5657 , P3_SUB_357_1258_U21 , P3_U2393 );
nand NAND2_3849 ( P3_U5658 , P3_ADD_558_U85 , P3_U3220 );
nand NAND2_3850 ( P3_U5659 , P3_ADD_553_U85 , P3_U4298 );
nand NAND2_3851 ( P3_U5660 , P3_ADD_547_U85 , P3_U4299 );
nand NAND2_3852 ( P3_U5661 , P3_ADD_541_U4 , P3_U4300 );
nand NAND2_3853 ( P3_U5662 , P3_ADD_536_U4 , P3_U4301 );
nand NAND2_3854 ( P3_U5663 , P3_ADD_531_U85 , P3_U2354 );
nand NAND2_3855 ( P3_U5664 , P3_ADD_526_U71 , P3_U2355 );
nand NAND2_3856 ( P3_U5665 , P3_ADD_515_U4 , P3_U4302 );
nand NAND2_3857 ( P3_U5666 , P3_ADD_494_U4 , P3_U2356 );
nand NAND2_3858 ( P3_U5667 , P3_ADD_476_U4 , P3_U4303 );
nand NAND2_3859 ( P3_U5668 , P3_ADD_441_U4 , P3_U4304 );
nand NAND2_3860 ( P3_U5669 , P3_ADD_405_U81 , P3_U4305 );
nand NAND2_3861 ( P3_U5670 , P3_ADD_394_U81 , P3_U2357 );
nand NAND2_3862 ( P3_U5671 , P3_ADD_385_U85 , P3_U2358 );
nand NAND2_3863 ( P3_U5672 , P3_ADD_380_U85 , P3_U2359 );
nand NAND2_3864 ( P3_U5673 , P3_ADD_349_U85 , P3_U4306 );
nand NAND2_3865 ( P3_U5674 , P3_ADD_344_U85 , P3_U2362 );
nand NAND2_3866 ( P3_U5675 , P3_ADD_371_1212_U20 , P3_U2360 );
nand NAND5_3867 ( P3_U5676 , P3_U5658 , P3_U3699 , P3_U5656 , P3_U3705 , P3_U3700 );
nand NAND2_3868 ( P3_U5677 , P3_U2402 , P3_REIP_REG_1_ );
nand NAND2_3869 ( P3_U5678 , P3_U4318 , P3_U5676 );
nand NAND2_3870 ( P3_U5679 , P3_U5631 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_3871 ( P3_U5680 , P3_ADD_360_1242_U91 , P3_U2395 );
nand NAND2_3872 ( P3_U5681 , P3_SUB_357_1258_U78 , P3_U2393 );
nand NAND2_3873 ( P3_U5682 , P3_ADD_558_U74 , P3_U3220 );
nand NAND2_3874 ( P3_U5683 , P3_ADD_553_U74 , P3_U4298 );
nand NAND2_3875 ( P3_U5684 , P3_ADD_547_U74 , P3_U4299 );
nand NAND2_3876 ( P3_U5685 , P3_ADD_541_U71 , P3_U4300 );
nand NAND2_3877 ( P3_U5686 , P3_ADD_536_U71 , P3_U4301 );
nand NAND2_3878 ( P3_U5687 , P3_ADD_531_U74 , P3_U2354 );
nand NAND2_3879 ( P3_U5688 , P3_ADD_526_U60 , P3_U2355 );
nand NAND2_3880 ( P3_U5689 , P3_ADD_515_U71 , P3_U4302 );
nand NAND2_3881 ( P3_U5690 , P3_ADD_494_U71 , P3_U2356 );
nand NAND2_3882 ( P3_U5691 , P3_ADD_476_U71 , P3_U4303 );
nand NAND2_3883 ( P3_U5692 , P3_ADD_441_U71 , P3_U4304 );
nand NAND2_3884 ( P3_U5693 , P3_ADD_405_U5 , P3_U4305 );
nand NAND2_3885 ( P3_U5694 , P3_ADD_394_U5 , P3_U2357 );
nand NAND2_3886 ( P3_U5695 , P3_ADD_385_U74 , P3_U2358 );
nand NAND2_3887 ( P3_U5696 , P3_ADD_380_U74 , P3_U2359 );
nand NAND2_3888 ( P3_U5697 , P3_ADD_349_U74 , P3_U4306 );
nand NAND2_3889 ( P3_U5698 , P3_ADD_344_U74 , P3_U2362 );
nand NAND2_3890 ( P3_U5699 , P3_ADD_371_1212_U93 , P3_U2360 );
nand NAND5_3891 ( P3_U5700 , P3_U5682 , P3_U3710 , P3_U5680 , P3_U3706 , P3_U3713 );
nand NAND2_3892 ( P3_U5701 , P3_U2402 , P3_REIP_REG_2_ );
nand NAND2_3893 ( P3_U5702 , P3_U4318 , P3_U5700 );
nand NAND2_3894 ( P3_U5703 , P3_INSTADDRPOINTER_REG_2_ , P3_U5631 );
nand NAND2_3895 ( P3_U5704 , P3_ADD_360_1242_U17 , P3_U2395 );
nand NAND2_3896 ( P3_U5705 , P3_SUB_357_1258_U76 , P3_U2393 );
nand NAND2_3897 ( P3_U5706 , P3_ADD_558_U71 , P3_U3220 );
nand NAND2_3898 ( P3_U5707 , P3_ADD_553_U71 , P3_U4298 );
nand NAND2_3899 ( P3_U5708 , P3_ADD_547_U71 , P3_U4299 );
nand NAND2_3900 ( P3_U5709 , P3_ADD_541_U68 , P3_U4300 );
nand NAND2_3901 ( P3_U5710 , P3_ADD_536_U68 , P3_U4301 );
nand NAND2_3902 ( P3_U5711 , P3_ADD_531_U71 , P3_U2354 );
nand NAND2_3903 ( P3_U5712 , P3_ADD_526_U57 , P3_U2355 );
nand NAND2_3904 ( P3_U5713 , P3_ADD_515_U68 , P3_U4302 );
nand NAND2_3905 ( P3_U5714 , P3_ADD_494_U68 , P3_U2356 );
nand NAND2_3906 ( P3_U5715 , P3_ADD_476_U68 , P3_U4303 );
nand NAND2_3907 ( P3_U5716 , P3_ADD_441_U68 , P3_U4304 );
nand NAND2_3908 ( P3_U5717 , P3_ADD_405_U93 , P3_U4305 );
nand NAND2_3909 ( P3_U5718 , P3_ADD_394_U93 , P3_U2357 );
nand NAND2_3910 ( P3_U5719 , P3_ADD_385_U71 , P3_U2358 );
nand NAND2_3911 ( P3_U5720 , P3_ADD_380_U71 , P3_U2359 );
nand NAND2_3912 ( P3_U5721 , P3_ADD_349_U71 , P3_U4306 );
nand NAND2_3913 ( P3_U5722 , P3_ADD_344_U71 , P3_U2362 );
nand NAND2_3914 ( P3_U5723 , P3_ADD_371_1212_U18 , P3_U2360 );
nand NAND5_3915 ( P3_U5724 , P3_U3715 , P3_U5706 , P3_U3718 , P3_U3714 , P3_U3721 );
nand NAND2_3916 ( P3_U5725 , P3_U2402 , P3_REIP_REG_3_ );
nand NAND2_3917 ( P3_U5726 , P3_U4318 , P3_U5724 );
nand NAND2_3918 ( P3_U5727 , P3_INSTADDRPOINTER_REG_3_ , P3_U5631 );
nand NAND2_3919 ( P3_U5728 , P3_ADD_360_1242_U18 , P3_U2395 );
nand NAND2_3920 ( P3_U5729 , P3_SUB_357_1258_U75 , P3_U2393 );
nand NAND2_3921 ( P3_U5730 , P3_ADD_558_U70 , P3_U3220 );
nand NAND2_3922 ( P3_U5731 , P3_ADD_553_U70 , P3_U4298 );
nand NAND2_3923 ( P3_U5732 , P3_ADD_547_U70 , P3_U4299 );
nand NAND2_3924 ( P3_U5733 , P3_ADD_541_U67 , P3_U4300 );
nand NAND2_3925 ( P3_U5734 , P3_ADD_536_U67 , P3_U4301 );
nand NAND2_3926 ( P3_U5735 , P3_ADD_531_U70 , P3_U2354 );
nand NAND2_3927 ( P3_U5736 , P3_ADD_526_U56 , P3_U2355 );
nand NAND2_3928 ( P3_U5737 , P3_ADD_515_U67 , P3_U4302 );
nand NAND2_3929 ( P3_U5738 , P3_ADD_494_U67 , P3_U2356 );
nand NAND2_3930 ( P3_U5739 , P3_ADD_476_U67 , P3_U4303 );
nand NAND2_3931 ( P3_U5740 , P3_ADD_441_U67 , P3_U4304 );
nand NAND2_3932 ( P3_U5741 , P3_ADD_405_U68 , P3_U4305 );
nand NAND2_3933 ( P3_U5742 , P3_ADD_394_U68 , P3_U2357 );
nand NAND2_3934 ( P3_U5743 , P3_ADD_385_U70 , P3_U2358 );
nand NAND2_3935 ( P3_U5744 , P3_ADD_380_U70 , P3_U2359 );
nand NAND2_3936 ( P3_U5745 , P3_ADD_349_U70 , P3_U4306 );
nand NAND2_3937 ( P3_U5746 , P3_ADD_344_U70 , P3_U2362 );
nand NAND2_3938 ( P3_U5747 , P3_ADD_371_1212_U91 , P3_U2360 );
nand NAND5_3939 ( P3_U5748 , P3_U5730 , P3_U3726 , P3_U5728 , P3_U3722 , P3_U3729 );
nand NAND2_3940 ( P3_U5749 , P3_U2402 , P3_REIP_REG_4_ );
nand NAND2_3941 ( P3_U5750 , P3_U4318 , P3_U5748 );
nand NAND2_3942 ( P3_U5751 , P3_INSTADDRPOINTER_REG_4_ , P3_U5631 );
nand NAND2_3943 ( P3_U5752 , P3_ADD_360_1242_U89 , P3_U2395 );
nand NAND2_3944 ( P3_U5753 , P3_SUB_357_1258_U74 , P3_U2393 );
nand NAND2_3945 ( P3_U5754 , P3_ADD_558_U69 , P3_U3220 );
nand NAND2_3946 ( P3_U5755 , P3_ADD_553_U69 , P3_U4298 );
nand NAND2_3947 ( P3_U5756 , P3_ADD_547_U69 , P3_U4299 );
nand NAND2_3948 ( P3_U5757 , P3_ADD_541_U66 , P3_U4300 );
nand NAND2_3949 ( P3_U5758 , P3_ADD_536_U66 , P3_U4301 );
nand NAND2_3950 ( P3_U5759 , P3_ADD_531_U69 , P3_U2354 );
nand NAND2_3951 ( P3_U5760 , P3_ADD_526_U55 , P3_U2355 );
nand NAND2_3952 ( P3_U5761 , P3_ADD_515_U66 , P3_U4302 );
nand NAND2_3953 ( P3_U5762 , P3_ADD_494_U66 , P3_U2356 );
nand NAND2_3954 ( P3_U5763 , P3_ADD_476_U66 , P3_U4303 );
nand NAND2_3955 ( P3_U5764 , P3_ADD_441_U66 , P3_U4304 );
nand NAND2_3956 ( P3_U5765 , P3_ADD_405_U67 , P3_U4305 );
nand NAND2_3957 ( P3_U5766 , P3_ADD_394_U67 , P3_U2357 );
nand NAND2_3958 ( P3_U5767 , P3_ADD_385_U69 , P3_U2358 );
nand NAND2_3959 ( P3_U5768 , P3_ADD_380_U69 , P3_U2359 );
nand NAND2_3960 ( P3_U5769 , P3_ADD_349_U69 , P3_U4306 );
nand NAND2_3961 ( P3_U5770 , P3_ADD_344_U69 , P3_U2362 );
nand NAND2_3962 ( P3_U5771 , P3_ADD_371_1212_U19 , P3_U2360 );
nand NAND5_3963 ( P3_U5772 , P3_U3734 , P3_U5754 , P3_U5753 , P3_U3730 , P3_U3737 );
nand NAND2_3964 ( P3_U5773 , P3_U2402 , P3_REIP_REG_5_ );
nand NAND2_3965 ( P3_U5774 , P3_U4318 , P3_U5772 );
nand NAND2_3966 ( P3_U5775 , P3_INSTADDRPOINTER_REG_5_ , P3_U5631 );
nand NAND2_3967 ( P3_U5776 , P3_ADD_360_1242_U88 , P3_U2395 );
nand NAND2_3968 ( P3_U5777 , P3_SUB_357_1258_U73 , P3_U2393 );
nand NAND2_3969 ( P3_U5778 , P3_ADD_558_U68 , P3_U3220 );
nand NAND2_3970 ( P3_U5779 , P3_ADD_553_U68 , P3_U4298 );
nand NAND2_3971 ( P3_U5780 , P3_ADD_547_U68 , P3_U4299 );
nand NAND2_3972 ( P3_U5781 , P3_ADD_541_U65 , P3_U4300 );
nand NAND2_3973 ( P3_U5782 , P3_ADD_536_U65 , P3_U4301 );
nand NAND2_3974 ( P3_U5783 , P3_ADD_531_U68 , P3_U2354 );
nand NAND2_3975 ( P3_U5784 , P3_ADD_526_U54 , P3_U2355 );
nand NAND2_3976 ( P3_U5785 , P3_ADD_515_U65 , P3_U4302 );
nand NAND2_3977 ( P3_U5786 , P3_ADD_494_U65 , P3_U2356 );
nand NAND2_3978 ( P3_U5787 , P3_ADD_476_U65 , P3_U4303 );
nand NAND2_3979 ( P3_U5788 , P3_ADD_441_U65 , P3_U4304 );
nand NAND2_3980 ( P3_U5789 , P3_ADD_405_U66 , P3_U4305 );
nand NAND2_3981 ( P3_U5790 , P3_ADD_394_U66 , P3_U2357 );
nand NAND2_3982 ( P3_U5791 , P3_ADD_385_U68 , P3_U2358 );
nand NAND2_3983 ( P3_U5792 , P3_ADD_380_U68 , P3_U2359 );
nand NAND2_3984 ( P3_U5793 , P3_ADD_349_U68 , P3_U4306 );
nand NAND2_3985 ( P3_U5794 , P3_ADD_344_U68 , P3_U2362 );
nand NAND2_3986 ( P3_U5795 , P3_ADD_371_1212_U90 , P3_U2360 );
nand NAND5_3987 ( P3_U5796 , P3_U3742 , P3_U5778 , P3_U5777 , P3_U3738 , P3_U3745 );
nand NAND2_3988 ( P3_U5797 , P3_U2402 , P3_REIP_REG_6_ );
nand NAND2_3989 ( P3_U5798 , P3_U4318 , P3_U5796 );
nand NAND2_3990 ( P3_U5799 , P3_INSTADDRPOINTER_REG_6_ , P3_U5631 );
nand NAND2_3991 ( P3_U5800 , P3_ADD_360_1242_U87 , P3_U2395 );
nand NAND2_3992 ( P3_U5801 , P3_SUB_357_1258_U72 , P3_U2393 );
nand NAND2_3993 ( P3_U5802 , P3_ADD_558_U67 , P3_U3220 );
nand NAND2_3994 ( P3_U5803 , P3_ADD_553_U67 , P3_U4298 );
nand NAND2_3995 ( P3_U5804 , P3_ADD_547_U67 , P3_U4299 );
nand NAND2_3996 ( P3_U5805 , P3_ADD_541_U64 , P3_U4300 );
nand NAND2_3997 ( P3_U5806 , P3_ADD_536_U64 , P3_U4301 );
nand NAND2_3998 ( P3_U5807 , P3_ADD_531_U67 , P3_U2354 );
nand NAND2_3999 ( P3_U5808 , P3_ADD_526_U53 , P3_U2355 );
nand NAND2_4000 ( P3_U5809 , P3_ADD_515_U64 , P3_U4302 );
nand NAND2_4001 ( P3_U5810 , P3_ADD_494_U64 , P3_U2356 );
nand NAND2_4002 ( P3_U5811 , P3_ADD_476_U64 , P3_U4303 );
nand NAND2_4003 ( P3_U5812 , P3_ADD_441_U64 , P3_U4304 );
nand NAND2_4004 ( P3_U5813 , P3_ADD_405_U65 , P3_U4305 );
nand NAND2_4005 ( P3_U5814 , P3_ADD_394_U65 , P3_U2357 );
nand NAND2_4006 ( P3_U5815 , P3_ADD_385_U67 , P3_U2358 );
nand NAND2_4007 ( P3_U5816 , P3_ADD_380_U67 , P3_U2359 );
nand NAND2_4008 ( P3_U5817 , P3_ADD_349_U67 , P3_U4306 );
nand NAND2_4009 ( P3_U5818 , P3_ADD_344_U67 , P3_U2362 );
nand NAND2_4010 ( P3_U5819 , P3_ADD_371_1212_U89 , P3_U2360 );
nand NAND5_4011 ( P3_U5820 , P3_U3750 , P3_U5802 , P3_U5801 , P3_U3746 , P3_U3753 );
nand NAND2_4012 ( P3_U5821 , P3_U2402 , P3_REIP_REG_7_ );
nand NAND2_4013 ( P3_U5822 , P3_U4318 , P3_U5820 );
nand NAND2_4014 ( P3_U5823 , P3_INSTADDRPOINTER_REG_7_ , P3_U5631 );
nand NAND2_4015 ( P3_U5824 , P3_ADD_360_1242_U86 , P3_U2395 );
nand NAND2_4016 ( P3_U5825 , P3_SUB_357_1258_U71 , P3_U2393 );
nand NAND2_4017 ( P3_U5826 , P3_ADD_558_U66 , P3_U3220 );
nand NAND2_4018 ( P3_U5827 , P3_ADD_553_U66 , P3_U4298 );
nand NAND2_4019 ( P3_U5828 , P3_ADD_547_U66 , P3_U4299 );
nand NAND2_4020 ( P3_U5829 , P3_ADD_541_U63 , P3_U4300 );
nand NAND2_4021 ( P3_U5830 , P3_ADD_536_U63 , P3_U4301 );
nand NAND2_4022 ( P3_U5831 , P3_ADD_531_U66 , P3_U2354 );
nand NAND2_4023 ( P3_U5832 , P3_ADD_526_U52 , P3_U2355 );
nand NAND2_4024 ( P3_U5833 , P3_ADD_515_U63 , P3_U4302 );
nand NAND2_4025 ( P3_U5834 , P3_ADD_494_U63 , P3_U2356 );
nand NAND2_4026 ( P3_U5835 , P3_ADD_476_U63 , P3_U4303 );
nand NAND2_4027 ( P3_U5836 , P3_ADD_441_U63 , P3_U4304 );
nand NAND2_4028 ( P3_U5837 , P3_ADD_405_U64 , P3_U4305 );
nand NAND2_4029 ( P3_U5838 , P3_ADD_394_U64 , P3_U2357 );
nand NAND2_4030 ( P3_U5839 , P3_ADD_385_U66 , P3_U2358 );
nand NAND2_4031 ( P3_U5840 , P3_ADD_380_U66 , P3_U2359 );
nand NAND2_4032 ( P3_U5841 , P3_ADD_349_U66 , P3_U4306 );
nand NAND2_4033 ( P3_U5842 , P3_ADD_344_U66 , P3_U2362 );
nand NAND2_4034 ( P3_U5843 , P3_ADD_371_1212_U88 , P3_U2360 );
nand NAND5_4035 ( P3_U5844 , P3_U3757 , P3_U5826 , P3_U5825 , P3_U3754 , P3_U3760 );
nand NAND2_4036 ( P3_U5845 , P3_U2402 , P3_REIP_REG_8_ );
nand NAND2_4037 ( P3_U5846 , P3_U4318 , P3_U5844 );
nand NAND2_4038 ( P3_U5847 , P3_INSTADDRPOINTER_REG_8_ , P3_U5631 );
nand NAND2_4039 ( P3_U5848 , P3_ADD_360_1242_U106 , P3_U2395 );
nand NAND2_4040 ( P3_U5849 , P3_SUB_357_1258_U70 , P3_U2393 );
nand NAND2_4041 ( P3_U5850 , P3_ADD_558_U65 , P3_U3220 );
nand NAND2_4042 ( P3_U5851 , P3_ADD_553_U65 , P3_U4298 );
nand NAND2_4043 ( P3_U5852 , P3_ADD_547_U65 , P3_U4299 );
nand NAND2_4044 ( P3_U5853 , P3_ADD_541_U62 , P3_U4300 );
nand NAND2_4045 ( P3_U5854 , P3_ADD_536_U62 , P3_U4301 );
nand NAND2_4046 ( P3_U5855 , P3_ADD_531_U65 , P3_U2354 );
nand NAND2_4047 ( P3_U5856 , P3_ADD_526_U51 , P3_U2355 );
nand NAND2_4048 ( P3_U5857 , P3_ADD_515_U62 , P3_U4302 );
nand NAND2_4049 ( P3_U5858 , P3_ADD_494_U62 , P3_U2356 );
nand NAND2_4050 ( P3_U5859 , P3_ADD_476_U62 , P3_U4303 );
nand NAND2_4051 ( P3_U5860 , P3_ADD_441_U62 , P3_U4304 );
nand NAND2_4052 ( P3_U5861 , P3_ADD_405_U63 , P3_U4305 );
nand NAND2_4053 ( P3_U5862 , P3_ADD_394_U63 , P3_U2357 );
nand NAND2_4054 ( P3_U5863 , P3_ADD_385_U65 , P3_U2358 );
nand NAND2_4055 ( P3_U5864 , P3_ADD_380_U65 , P3_U2359 );
nand NAND2_4056 ( P3_U5865 , P3_ADD_349_U65 , P3_U4306 );
nand NAND2_4057 ( P3_U5866 , P3_ADD_344_U65 , P3_U2362 );
nand NAND2_4058 ( P3_U5867 , P3_ADD_371_1212_U109 , P3_U2360 );
nand NAND5_4059 ( P3_U5868 , P3_U3764 , P3_U5850 , P3_U5849 , P3_U3761 , P3_U3767 );
nand NAND2_4060 ( P3_U5869 , P3_U2402 , P3_REIP_REG_9_ );
nand NAND2_4061 ( P3_U5870 , P3_U4318 , P3_U5868 );
nand NAND2_4062 ( P3_U5871 , P3_INSTADDRPOINTER_REG_9_ , P3_U5631 );
nand NAND2_4063 ( P3_U5872 , P3_ADD_360_1242_U4 , P3_U2395 );
nand NAND2_4064 ( P3_U5873 , P3_SUB_357_1258_U93 , P3_U2393 );
nand NAND2_4065 ( P3_U5874 , P3_ADD_558_U95 , P3_U3220 );
nand NAND2_4066 ( P3_U5875 , P3_ADD_553_U95 , P3_U4298 );
nand NAND2_4067 ( P3_U5876 , P3_ADD_547_U95 , P3_U4299 );
nand NAND2_4068 ( P3_U5877 , P3_ADD_541_U91 , P3_U4300 );
nand NAND2_4069 ( P3_U5878 , P3_ADD_536_U91 , P3_U4301 );
nand NAND2_4070 ( P3_U5879 , P3_ADD_531_U95 , P3_U2354 );
nand NAND2_4071 ( P3_U5880 , P3_ADD_526_U81 , P3_U2355 );
nand NAND2_4072 ( P3_U5881 , P3_ADD_515_U91 , P3_U4302 );
nand NAND2_4073 ( P3_U5882 , P3_ADD_494_U91 , P3_U2356 );
nand NAND2_4074 ( P3_U5883 , P3_ADD_476_U91 , P3_U4303 );
nand NAND2_4075 ( P3_U5884 , P3_ADD_441_U91 , P3_U4304 );
nand NAND2_4076 ( P3_U5885 , P3_ADD_405_U91 , P3_U4305 );
nand NAND2_4077 ( P3_U5886 , P3_ADD_394_U91 , P3_U2357 );
nand NAND2_4078 ( P3_U5887 , P3_ADD_385_U95 , P3_U2358 );
nand NAND2_4079 ( P3_U5888 , P3_ADD_380_U95 , P3_U2359 );
nand NAND2_4080 ( P3_U5889 , P3_ADD_349_U95 , P3_U4306 );
nand NAND2_4081 ( P3_U5890 , P3_ADD_344_U95 , P3_U2362 );
nand NAND2_4082 ( P3_U5891 , P3_ADD_371_1212_U5 , P3_U2360 );
nand NAND5_4083 ( P3_U5892 , P3_U5874 , P3_U3771 , P3_U5872 , P3_U3774 , P3_U3768 );
nand NAND2_4084 ( P3_U5893 , P3_U2402 , P3_REIP_REG_10_ );
nand NAND2_4085 ( P3_U5894 , P3_U4318 , P3_U5892 );
nand NAND2_4086 ( P3_U5895 , P3_INSTADDRPOINTER_REG_10_ , P3_U5631 );
nand NAND2_4087 ( P3_U5896 , P3_ADD_360_1242_U84 , P3_U2395 );
nand NAND2_4088 ( P3_U5897 , P3_SUB_357_1258_U92 , P3_U2393 );
nand NAND2_4089 ( P3_U5898 , P3_ADD_558_U94 , P3_U3220 );
nand NAND2_4090 ( P3_U5899 , P3_ADD_553_U94 , P3_U4298 );
nand NAND2_4091 ( P3_U5900 , P3_ADD_547_U94 , P3_U4299 );
nand NAND2_4092 ( P3_U5901 , P3_ADD_541_U90 , P3_U4300 );
nand NAND2_4093 ( P3_U5902 , P3_ADD_536_U90 , P3_U4301 );
nand NAND2_4094 ( P3_U5903 , P3_ADD_531_U94 , P3_U2354 );
nand NAND2_4095 ( P3_U5904 , P3_ADD_526_U80 , P3_U2355 );
nand NAND2_4096 ( P3_U5905 , P3_ADD_515_U90 , P3_U4302 );
nand NAND2_4097 ( P3_U5906 , P3_ADD_494_U90 , P3_U2356 );
nand NAND2_4098 ( P3_U5907 , P3_ADD_476_U90 , P3_U4303 );
nand NAND2_4099 ( P3_U5908 , P3_ADD_441_U90 , P3_U4304 );
nand NAND2_4100 ( P3_U5909 , P3_ADD_405_U90 , P3_U4305 );
nand NAND2_4101 ( P3_U5910 , P3_ADD_394_U90 , P3_U2357 );
nand NAND2_4102 ( P3_U5911 , P3_ADD_385_U94 , P3_U2358 );
nand NAND2_4103 ( P3_U5912 , P3_ADD_380_U94 , P3_U2359 );
nand NAND2_4104 ( P3_U5913 , P3_ADD_349_U94 , P3_U4306 );
nand NAND2_4105 ( P3_U5914 , P3_ADD_344_U94 , P3_U2362 );
nand NAND2_4106 ( P3_U5915 , P3_ADD_371_1212_U86 , P3_U2360 );
nand NAND5_4107 ( P3_U5916 , P3_U5898 , P3_U3778 , P3_U5896 , P3_U3775 , P3_U3781 );
nand NAND2_4108 ( P3_U5917 , P3_U2402 , P3_REIP_REG_11_ );
nand NAND2_4109 ( P3_U5918 , P3_U4318 , P3_U5916 );
nand NAND2_4110 ( P3_U5919 , P3_INSTADDRPOINTER_REG_11_ , P3_U5631 );
nand NAND2_4111 ( P3_U5920 , P3_ADD_360_1242_U5 , P3_U2395 );
nand NAND2_4112 ( P3_U5921 , P3_SUB_357_1258_U91 , P3_U2393 );
nand NAND2_4113 ( P3_U5922 , P3_ADD_558_U93 , P3_U3220 );
nand NAND2_4114 ( P3_U5923 , P3_ADD_553_U93 , P3_U4298 );
nand NAND2_4115 ( P3_U5924 , P3_ADD_547_U93 , P3_U4299 );
nand NAND2_4116 ( P3_U5925 , P3_ADD_541_U89 , P3_U4300 );
nand NAND2_4117 ( P3_U5926 , P3_ADD_536_U89 , P3_U4301 );
nand NAND2_4118 ( P3_U5927 , P3_ADD_531_U93 , P3_U2354 );
nand NAND2_4119 ( P3_U5928 , P3_ADD_526_U79 , P3_U2355 );
nand NAND2_4120 ( P3_U5929 , P3_ADD_515_U89 , P3_U4302 );
nand NAND2_4121 ( P3_U5930 , P3_ADD_494_U89 , P3_U2356 );
nand NAND2_4122 ( P3_U5931 , P3_ADD_476_U89 , P3_U4303 );
nand NAND2_4123 ( P3_U5932 , P3_ADD_441_U89 , P3_U4304 );
nand NAND2_4124 ( P3_U5933 , P3_ADD_405_U89 , P3_U4305 );
nand NAND2_4125 ( P3_U5934 , P3_ADD_394_U89 , P3_U2357 );
nand NAND2_4126 ( P3_U5935 , P3_ADD_385_U93 , P3_U2358 );
nand NAND2_4127 ( P3_U5936 , P3_ADD_380_U93 , P3_U2359 );
nand NAND2_4128 ( P3_U5937 , P3_ADD_349_U93 , P3_U4306 );
nand NAND2_4129 ( P3_U5938 , P3_ADD_344_U93 , P3_U2362 );
nand NAND2_4130 ( P3_U5939 , P3_ADD_371_1212_U6 , P3_U2360 );
nand NAND5_4131 ( P3_U5940 , P3_U3785 , P3_U5922 , P3_U5921 , P3_U3782 , P3_U3788 );
nand NAND2_4132 ( P3_U5941 , P3_U2402 , P3_REIP_REG_12_ );
nand NAND2_4133 ( P3_U5942 , P3_U4318 , P3_U5940 );
nand NAND2_4134 ( P3_U5943 , P3_INSTADDRPOINTER_REG_12_ , P3_U5631 );
nand NAND2_4135 ( P3_U5944 , P3_ADD_360_1242_U6 , P3_U2395 );
nand NAND2_4136 ( P3_U5945 , P3_SUB_357_1258_U15 , P3_U2393 );
nand NAND2_4137 ( P3_U5946 , P3_ADD_558_U92 , P3_U3220 );
nand NAND2_4138 ( P3_U5947 , P3_ADD_553_U92 , P3_U4298 );
nand NAND2_4139 ( P3_U5948 , P3_ADD_547_U92 , P3_U4299 );
nand NAND2_4140 ( P3_U5949 , P3_ADD_541_U88 , P3_U4300 );
nand NAND2_4141 ( P3_U5950 , P3_ADD_536_U88 , P3_U4301 );
nand NAND2_4142 ( P3_U5951 , P3_ADD_531_U92 , P3_U2354 );
nand NAND2_4143 ( P3_U5952 , P3_ADD_526_U78 , P3_U2355 );
nand NAND2_4144 ( P3_U5953 , P3_ADD_515_U88 , P3_U4302 );
nand NAND2_4145 ( P3_U5954 , P3_ADD_494_U88 , P3_U2356 );
nand NAND2_4146 ( P3_U5955 , P3_ADD_476_U88 , P3_U4303 );
nand NAND2_4147 ( P3_U5956 , P3_ADD_441_U88 , P3_U4304 );
nand NAND2_4148 ( P3_U5957 , P3_ADD_405_U88 , P3_U4305 );
nand NAND2_4149 ( P3_U5958 , P3_ADD_394_U88 , P3_U2357 );
nand NAND2_4150 ( P3_U5959 , P3_ADD_385_U92 , P3_U2358 );
nand NAND2_4151 ( P3_U5960 , P3_ADD_380_U92 , P3_U2359 );
nand NAND2_4152 ( P3_U5961 , P3_ADD_349_U92 , P3_U4306 );
nand NAND2_4153 ( P3_U5962 , P3_ADD_344_U92 , P3_U2362 );
nand NAND2_4154 ( P3_U5963 , P3_ADD_371_1212_U7 , P3_U2360 );
nand NAND5_4155 ( P3_U5964 , P3_U3792 , P3_U5946 , P3_U5945 , P3_U3789 , P3_U3795 );
nand NAND2_4156 ( P3_U5965 , P3_U2402 , P3_REIP_REG_13_ );
nand NAND2_4157 ( P3_U5966 , P3_U4318 , P3_U5964 );
nand NAND2_4158 ( P3_U5967 , P3_INSTADDRPOINTER_REG_13_ , P3_U5631 );
nand NAND2_4159 ( P3_U5968 , P3_ADD_360_1242_U83 , P3_U2395 );
nand NAND2_4160 ( P3_U5969 , P3_SUB_357_1258_U90 , P3_U2393 );
nand NAND2_4161 ( P3_U5970 , P3_ADD_558_U91 , P3_U3220 );
nand NAND2_4162 ( P3_U5971 , P3_ADD_553_U91 , P3_U4298 );
nand NAND2_4163 ( P3_U5972 , P3_ADD_547_U91 , P3_U4299 );
nand NAND2_4164 ( P3_U5973 , P3_ADD_541_U87 , P3_U4300 );
nand NAND2_4165 ( P3_U5974 , P3_ADD_536_U87 , P3_U4301 );
nand NAND2_4166 ( P3_U5975 , P3_ADD_531_U91 , P3_U2354 );
nand NAND2_4167 ( P3_U5976 , P3_ADD_526_U77 , P3_U2355 );
nand NAND2_4168 ( P3_U5977 , P3_ADD_515_U87 , P3_U4302 );
nand NAND2_4169 ( P3_U5978 , P3_ADD_494_U87 , P3_U2356 );
nand NAND2_4170 ( P3_U5979 , P3_ADD_476_U87 , P3_U4303 );
nand NAND2_4171 ( P3_U5980 , P3_ADD_441_U87 , P3_U4304 );
nand NAND2_4172 ( P3_U5981 , P3_ADD_405_U87 , P3_U4305 );
nand NAND2_4173 ( P3_U5982 , P3_ADD_394_U87 , P3_U2357 );
nand NAND2_4174 ( P3_U5983 , P3_ADD_385_U91 , P3_U2358 );
nand NAND2_4175 ( P3_U5984 , P3_ADD_380_U91 , P3_U2359 );
nand NAND2_4176 ( P3_U5985 , P3_ADD_349_U91 , P3_U4306 );
nand NAND2_4177 ( P3_U5986 , P3_ADD_344_U91 , P3_U2362 );
nand NAND2_4178 ( P3_U5987 , P3_ADD_371_1212_U85 , P3_U2360 );
nand NAND2_4179 ( P3_U5988 , P3_U3802 , P3_U3799 );
nand NAND2_4180 ( P3_U5989 , P3_U2402 , P3_REIP_REG_14_ );
nand NAND2_4181 ( P3_U5990 , P3_U4318 , P3_U5988 );
nand NAND2_4182 ( P3_U5991 , P3_INSTADDRPOINTER_REG_14_ , P3_U5631 );
nand NAND2_4183 ( P3_U5992 , P3_ADD_360_1242_U7 , P3_U2395 );
nand NAND2_4184 ( P3_U5993 , P3_SUB_357_1258_U89 , P3_U2393 );
nand NAND2_4185 ( P3_U5994 , P3_ADD_558_U90 , P3_U3220 );
nand NAND2_4186 ( P3_U5995 , P3_ADD_553_U90 , P3_U4298 );
nand NAND2_4187 ( P3_U5996 , P3_ADD_547_U90 , P3_U4299 );
nand NAND2_4188 ( P3_U5997 , P3_ADD_541_U86 , P3_U4300 );
nand NAND2_4189 ( P3_U5998 , P3_ADD_536_U86 , P3_U4301 );
nand NAND2_4190 ( P3_U5999 , P3_ADD_531_U90 , P3_U2354 );
nand NAND2_4191 ( P3_U6000 , P3_ADD_526_U76 , P3_U2355 );
nand NAND2_4192 ( P3_U6001 , P3_ADD_515_U86 , P3_U4302 );
nand NAND2_4193 ( P3_U6002 , P3_ADD_494_U86 , P3_U2356 );
nand NAND2_4194 ( P3_U6003 , P3_ADD_476_U86 , P3_U4303 );
nand NAND2_4195 ( P3_U6004 , P3_ADD_441_U86 , P3_U4304 );
nand NAND2_4196 ( P3_U6005 , P3_ADD_405_U86 , P3_U4305 );
nand NAND2_4197 ( P3_U6006 , P3_ADD_394_U86 , P3_U2357 );
nand NAND2_4198 ( P3_U6007 , P3_ADD_385_U90 , P3_U2358 );
nand NAND2_4199 ( P3_U6008 , P3_ADD_380_U90 , P3_U2359 );
nand NAND2_4200 ( P3_U6009 , P3_ADD_349_U90 , P3_U4306 );
nand NAND2_4201 ( P3_U6010 , P3_ADD_344_U90 , P3_U2362 );
nand NAND2_4202 ( P3_U6011 , P3_ADD_371_1212_U8 , P3_U2360 );
nand NAND2_4203 ( P3_U6012 , P3_U3810 , P3_U3807 );
nand NAND2_4204 ( P3_U6013 , P3_U2402 , P3_REIP_REG_15_ );
nand NAND2_4205 ( P3_U6014 , P3_U4318 , P3_U6012 );
nand NAND2_4206 ( P3_U6015 , P3_INSTADDRPOINTER_REG_15_ , P3_U5631 );
nand NAND2_4207 ( P3_U6016 , P3_ADD_360_1242_U82 , P3_U2395 );
nand NAND2_4208 ( P3_U6017 , P3_SUB_357_1258_U88 , P3_U2393 );
nand NAND2_4209 ( P3_U6018 , P3_ADD_558_U89 , P3_U3220 );
nand NAND2_4210 ( P3_U6019 , P3_ADD_553_U89 , P3_U4298 );
nand NAND2_4211 ( P3_U6020 , P3_ADD_547_U89 , P3_U4299 );
nand NAND2_4212 ( P3_U6021 , P3_ADD_541_U85 , P3_U4300 );
nand NAND2_4213 ( P3_U6022 , P3_ADD_536_U85 , P3_U4301 );
nand NAND2_4214 ( P3_U6023 , P3_ADD_531_U89 , P3_U2354 );
nand NAND2_4215 ( P3_U6024 , P3_ADD_526_U75 , P3_U2355 );
nand NAND2_4216 ( P3_U6025 , P3_ADD_515_U85 , P3_U4302 );
nand NAND2_4217 ( P3_U6026 , P3_ADD_494_U85 , P3_U2356 );
nand NAND2_4218 ( P3_U6027 , P3_ADD_476_U85 , P3_U4303 );
nand NAND2_4219 ( P3_U6028 , P3_ADD_441_U85 , P3_U4304 );
nand NAND2_4220 ( P3_U6029 , P3_ADD_405_U85 , P3_U4305 );
nand NAND2_4221 ( P3_U6030 , P3_ADD_394_U85 , P3_U2357 );
nand NAND2_4222 ( P3_U6031 , P3_ADD_385_U89 , P3_U2358 );
nand NAND2_4223 ( P3_U6032 , P3_ADD_380_U89 , P3_U2359 );
nand NAND2_4224 ( P3_U6033 , P3_ADD_349_U89 , P3_U4306 );
nand NAND2_4225 ( P3_U6034 , P3_ADD_344_U89 , P3_U2362 );
nand NAND2_4226 ( P3_U6035 , P3_ADD_371_1212_U84 , P3_U2360 );
nand NAND5_4227 ( P3_U6036 , P3_U6018 , P3_U3815 , P3_U6016 , P3_U3812 , P3_U3818 );
nand NAND2_4228 ( P3_U6037 , P3_U2402 , P3_REIP_REG_16_ );
nand NAND2_4229 ( P3_U6038 , P3_U4318 , P3_U6036 );
nand NAND2_4230 ( P3_U6039 , P3_INSTADDRPOINTER_REG_16_ , P3_U5631 );
nand NAND2_4231 ( P3_U6040 , P3_ADD_360_1242_U8 , P3_U2395 );
nand NAND2_4232 ( P3_U6041 , P3_SUB_357_1258_U16 , P3_U2393 );
nand NAND2_4233 ( P3_U6042 , P3_ADD_558_U88 , P3_U3220 );
nand NAND2_4234 ( P3_U6043 , P3_ADD_553_U88 , P3_U4298 );
nand NAND2_4235 ( P3_U6044 , P3_ADD_547_U88 , P3_U4299 );
nand NAND2_4236 ( P3_U6045 , P3_ADD_541_U84 , P3_U4300 );
nand NAND2_4237 ( P3_U6046 , P3_ADD_536_U84 , P3_U4301 );
nand NAND2_4238 ( P3_U6047 , P3_ADD_531_U88 , P3_U2354 );
nand NAND2_4239 ( P3_U6048 , P3_ADD_526_U74 , P3_U2355 );
nand NAND2_4240 ( P3_U6049 , P3_ADD_515_U84 , P3_U4302 );
nand NAND2_4241 ( P3_U6050 , P3_ADD_494_U84 , P3_U2356 );
nand NAND2_4242 ( P3_U6051 , P3_ADD_476_U84 , P3_U4303 );
nand NAND2_4243 ( P3_U6052 , P3_ADD_441_U84 , P3_U4304 );
nand NAND2_4244 ( P3_U6053 , P3_ADD_405_U84 , P3_U4305 );
nand NAND2_4245 ( P3_U6054 , P3_ADD_394_U84 , P3_U2357 );
nand NAND2_4246 ( P3_U6055 , P3_ADD_385_U88 , P3_U2358 );
nand NAND2_4247 ( P3_U6056 , P3_ADD_380_U88 , P3_U2359 );
nand NAND2_4248 ( P3_U6057 , P3_ADD_349_U88 , P3_U4306 );
nand NAND2_4249 ( P3_U6058 , P3_ADD_344_U88 , P3_U2362 );
nand NAND2_4250 ( P3_U6059 , P3_ADD_371_1212_U9 , P3_U2360 );
nand NAND5_4251 ( P3_U6060 , P3_U6042 , P3_U3819 , P3_U6040 , P3_U3824 , P3_U3820 );
nand NAND2_4252 ( P3_U6061 , P3_U2402 , P3_REIP_REG_17_ );
nand NAND2_4253 ( P3_U6062 , P3_U4318 , P3_U6060 );
nand NAND2_4254 ( P3_U6063 , P3_INSTADDRPOINTER_REG_17_ , P3_U5631 );
nand NAND2_4255 ( P3_U6064 , P3_ADD_360_1242_U81 , P3_U2395 );
nand NAND2_4256 ( P3_U6065 , P3_SUB_357_1258_U87 , P3_U2393 );
nand NAND2_4257 ( P3_U6066 , P3_ADD_558_U87 , P3_U3220 );
nand NAND2_4258 ( P3_U6067 , P3_ADD_553_U87 , P3_U4298 );
nand NAND2_4259 ( P3_U6068 , P3_ADD_547_U87 , P3_U4299 );
nand NAND2_4260 ( P3_U6069 , P3_ADD_541_U83 , P3_U4300 );
nand NAND2_4261 ( P3_U6070 , P3_ADD_536_U83 , P3_U4301 );
nand NAND2_4262 ( P3_U6071 , P3_ADD_531_U87 , P3_U2354 );
nand NAND2_4263 ( P3_U6072 , P3_ADD_526_U73 , P3_U2355 );
nand NAND2_4264 ( P3_U6073 , P3_ADD_515_U83 , P3_U4302 );
nand NAND2_4265 ( P3_U6074 , P3_ADD_494_U83 , P3_U2356 );
nand NAND2_4266 ( P3_U6075 , P3_ADD_476_U83 , P3_U4303 );
nand NAND2_4267 ( P3_U6076 , P3_ADD_441_U83 , P3_U4304 );
nand NAND2_4268 ( P3_U6077 , P3_ADD_405_U83 , P3_U4305 );
nand NAND2_4269 ( P3_U6078 , P3_ADD_394_U83 , P3_U2357 );
nand NAND2_4270 ( P3_U6079 , P3_ADD_385_U87 , P3_U2358 );
nand NAND2_4271 ( P3_U6080 , P3_ADD_380_U87 , P3_U2359 );
nand NAND2_4272 ( P3_U6081 , P3_ADD_349_U87 , P3_U4306 );
nand NAND2_4273 ( P3_U6082 , P3_ADD_344_U87 , P3_U2362 );
nand NAND2_4274 ( P3_U6083 , P3_ADD_371_1212_U83 , P3_U2360 );
nand NAND5_4275 ( P3_U6084 , P3_U6066 , P3_U3828 , P3_U6064 , P3_U3825 , P3_U3831 );
nand NAND2_4276 ( P3_U6085 , P3_U2402 , P3_REIP_REG_18_ );
nand NAND2_4277 ( P3_U6086 , P3_U4318 , P3_U6084 );
nand NAND2_4278 ( P3_U6087 , P3_INSTADDRPOINTER_REG_18_ , P3_U5631 );
nand NAND2_4279 ( P3_U6088 , P3_ADD_360_1242_U9 , P3_U2395 );
nand NAND2_4280 ( P3_U6089 , P3_SUB_357_1258_U86 , P3_U2393 );
nand NAND2_4281 ( P3_U6090 , P3_ADD_558_U86 , P3_U3220 );
nand NAND2_4282 ( P3_U6091 , P3_ADD_553_U86 , P3_U4298 );
nand NAND2_4283 ( P3_U6092 , P3_ADD_547_U86 , P3_U4299 );
nand NAND2_4284 ( P3_U6093 , P3_ADD_541_U82 , P3_U4300 );
nand NAND2_4285 ( P3_U6094 , P3_ADD_536_U82 , P3_U4301 );
nand NAND2_4286 ( P3_U6095 , P3_ADD_531_U86 , P3_U2354 );
nand NAND2_4287 ( P3_U6096 , P3_ADD_526_U72 , P3_U2355 );
nand NAND2_4288 ( P3_U6097 , P3_ADD_515_U82 , P3_U4302 );
nand NAND2_4289 ( P3_U6098 , P3_ADD_494_U82 , P3_U2356 );
nand NAND2_4290 ( P3_U6099 , P3_ADD_476_U82 , P3_U4303 );
nand NAND2_4291 ( P3_U6100 , P3_ADD_441_U82 , P3_U4304 );
nand NAND2_4292 ( P3_U6101 , P3_ADD_405_U82 , P3_U4305 );
nand NAND2_4293 ( P3_U6102 , P3_ADD_394_U82 , P3_U2357 );
nand NAND2_4294 ( P3_U6103 , P3_ADD_385_U86 , P3_U2358 );
nand NAND2_4295 ( P3_U6104 , P3_ADD_380_U86 , P3_U2359 );
nand NAND2_4296 ( P3_U6105 , P3_ADD_349_U86 , P3_U4306 );
nand NAND2_4297 ( P3_U6106 , P3_ADD_344_U86 , P3_U2362 );
nand NAND2_4298 ( P3_U6107 , P3_ADD_371_1212_U10 , P3_U2360 );
nand NAND5_4299 ( P3_U6108 , P3_U6090 , P3_U3832 , P3_U6088 , P3_U3837 , P3_U3833 );
nand NAND2_4300 ( P3_U6109 , P3_U2402 , P3_REIP_REG_19_ );
nand NAND2_4301 ( P3_U6110 , P3_U4318 , P3_U6108 );
nand NAND2_4302 ( P3_U6111 , P3_INSTADDRPOINTER_REG_19_ , P3_U5631 );
nand NAND2_4303 ( P3_U6112 , P3_ADD_360_1242_U10 , P3_U2395 );
nand NAND2_4304 ( P3_U6113 , P3_SUB_357_1258_U17 , P3_U2393 );
nand NAND2_4305 ( P3_U6114 , P3_ADD_558_U84 , P3_U3220 );
nand NAND2_4306 ( P3_U6115 , P3_ADD_553_U84 , P3_U4298 );
nand NAND2_4307 ( P3_U6116 , P3_ADD_547_U84 , P3_U4299 );
nand NAND2_4308 ( P3_U6117 , P3_ADD_541_U81 , P3_U4300 );
nand NAND2_4309 ( P3_U6118 , P3_ADD_536_U81 , P3_U4301 );
nand NAND2_4310 ( P3_U6119 , P3_ADD_531_U84 , P3_U2354 );
nand NAND2_4311 ( P3_U6120 , P3_ADD_526_U70 , P3_U2355 );
nand NAND2_4312 ( P3_U6121 , P3_ADD_515_U81 , P3_U4302 );
nand NAND2_4313 ( P3_U6122 , P3_ADD_494_U81 , P3_U2356 );
nand NAND2_4314 ( P3_U6123 , P3_ADD_476_U81 , P3_U4303 );
nand NAND2_4315 ( P3_U6124 , P3_ADD_441_U81 , P3_U4304 );
nand NAND2_4316 ( P3_U6125 , P3_ADD_405_U80 , P3_U4305 );
nand NAND2_4317 ( P3_U6126 , P3_ADD_394_U80 , P3_U2357 );
nand NAND2_4318 ( P3_U6127 , P3_ADD_385_U84 , P3_U2358 );
nand NAND2_4319 ( P3_U6128 , P3_ADD_380_U84 , P3_U2359 );
nand NAND2_4320 ( P3_U6129 , P3_ADD_349_U84 , P3_U4306 );
nand NAND2_4321 ( P3_U6130 , P3_ADD_344_U84 , P3_U2362 );
nand NAND2_4322 ( P3_U6131 , P3_ADD_371_1212_U11 , P3_U2360 );
nand NAND2_4323 ( P3_U6132 , P3_U6113 , P3_U3841 );
nand NAND2_4324 ( P3_U6133 , P3_U2402 , P3_REIP_REG_20_ );
nand NAND2_4325 ( P3_U6134 , P3_U4318 , P3_U6132 );
nand NAND2_4326 ( P3_U6135 , P3_INSTADDRPOINTER_REG_20_ , P3_U5631 );
nand NAND2_4327 ( P3_U6136 , P3_ADD_360_1242_U11 , P3_U2395 );
nand NAND2_4328 ( P3_U6137 , P3_SUB_357_1258_U85 , P3_U2393 );
nand NAND2_4329 ( P3_U6138 , P3_ADD_558_U83 , P3_U3220 );
nand NAND2_4330 ( P3_U6139 , P3_ADD_553_U83 , P3_U4298 );
nand NAND2_4331 ( P3_U6140 , P3_ADD_547_U83 , P3_U4299 );
nand NAND2_4332 ( P3_U6141 , P3_ADD_541_U80 , P3_U4300 );
nand NAND2_4333 ( P3_U6142 , P3_ADD_536_U80 , P3_U4301 );
nand NAND2_4334 ( P3_U6143 , P3_ADD_531_U83 , P3_U2354 );
nand NAND2_4335 ( P3_U6144 , P3_ADD_526_U69 , P3_U2355 );
nand NAND2_4336 ( P3_U6145 , P3_ADD_515_U80 , P3_U4302 );
nand NAND2_4337 ( P3_U6146 , P3_ADD_494_U80 , P3_U2356 );
nand NAND2_4338 ( P3_U6147 , P3_ADD_476_U80 , P3_U4303 );
nand NAND2_4339 ( P3_U6148 , P3_ADD_441_U80 , P3_U4304 );
nand NAND2_4340 ( P3_U6149 , P3_ADD_405_U79 , P3_U4305 );
nand NAND2_4341 ( P3_U6150 , P3_ADD_394_U79 , P3_U2357 );
nand NAND2_4342 ( P3_U6151 , P3_ADD_385_U83 , P3_U2358 );
nand NAND2_4343 ( P3_U6152 , P3_ADD_380_U83 , P3_U2359 );
nand NAND2_4344 ( P3_U6153 , P3_ADD_349_U83 , P3_U4306 );
nand NAND2_4345 ( P3_U6154 , P3_ADD_344_U83 , P3_U2362 );
nand NAND2_4346 ( P3_U6155 , P3_ADD_371_1212_U12 , P3_U2360 );
nand NAND2_4347 ( P3_U6156 , P3_U6137 , P3_U3849 );
nand NAND2_4348 ( P3_U6157 , P3_U2402 , P3_REIP_REG_21_ );
nand NAND2_4349 ( P3_U6158 , P3_U4318 , P3_U6156 );
nand NAND2_4350 ( P3_U6159 , P3_INSTADDRPOINTER_REG_21_ , P3_U5631 );
nand NAND2_4351 ( P3_U6160 , P3_ADD_360_1242_U80 , P3_U2395 );
nand NAND2_4352 ( P3_U6161 , P3_SUB_357_1258_U84 , P3_U2393 );
nand NAND2_4353 ( P3_U6162 , P3_ADD_558_U82 , P3_U3220 );
nand NAND2_4354 ( P3_U6163 , P3_ADD_553_U82 , P3_U4298 );
nand NAND2_4355 ( P3_U6164 , P3_ADD_547_U82 , P3_U4299 );
nand NAND2_4356 ( P3_U6165 , P3_ADD_541_U79 , P3_U4300 );
nand NAND2_4357 ( P3_U6166 , P3_ADD_536_U79 , P3_U4301 );
nand NAND2_4358 ( P3_U6167 , P3_ADD_531_U82 , P3_U2354 );
nand NAND2_4359 ( P3_U6168 , P3_ADD_526_U68 , P3_U2355 );
nand NAND2_4360 ( P3_U6169 , P3_ADD_515_U79 , P3_U4302 );
nand NAND2_4361 ( P3_U6170 , P3_ADD_494_U79 , P3_U2356 );
nand NAND2_4362 ( P3_U6171 , P3_ADD_476_U79 , P3_U4303 );
nand NAND2_4363 ( P3_U6172 , P3_ADD_441_U79 , P3_U4304 );
nand NAND2_4364 ( P3_U6173 , P3_ADD_405_U78 , P3_U4305 );
nand NAND2_4365 ( P3_U6174 , P3_ADD_394_U78 , P3_U2357 );
nand NAND2_4366 ( P3_U6175 , P3_ADD_385_U82 , P3_U2358 );
nand NAND2_4367 ( P3_U6176 , P3_ADD_380_U82 , P3_U2359 );
nand NAND2_4368 ( P3_U6177 , P3_ADD_349_U82 , P3_U4306 );
nand NAND2_4369 ( P3_U6178 , P3_ADD_344_U82 , P3_U2362 );
nand NAND2_4370 ( P3_U6179 , P3_ADD_371_1212_U82 , P3_U2360 );
nand NAND2_4371 ( P3_U6180 , P3_U3862 , P3_U3857 );
nand NAND2_4372 ( P3_U6181 , P3_U2402 , P3_REIP_REG_22_ );
nand NAND2_4373 ( P3_U6182 , P3_U4318 , P3_U6180 );
nand NAND2_4374 ( P3_U6183 , P3_INSTADDRPOINTER_REG_22_ , P3_U5631 );
nand NAND2_4375 ( P3_U6184 , P3_ADD_360_1242_U12 , P3_U2395 );
nand NAND2_4376 ( P3_U6185 , P3_SUB_357_1258_U83 , P3_U2393 );
nand NAND2_4377 ( P3_U6186 , P3_ADD_558_U81 , P3_U3220 );
nand NAND2_4378 ( P3_U6187 , P3_ADD_553_U81 , P3_U4298 );
nand NAND2_4379 ( P3_U6188 , P3_ADD_547_U81 , P3_U4299 );
nand NAND2_4380 ( P3_U6189 , P3_ADD_541_U78 , P3_U4300 );
nand NAND2_4381 ( P3_U6190 , P3_ADD_536_U78 , P3_U4301 );
nand NAND2_4382 ( P3_U6191 , P3_ADD_531_U81 , P3_U2354 );
nand NAND2_4383 ( P3_U6192 , P3_ADD_526_U67 , P3_U2355 );
nand NAND2_4384 ( P3_U6193 , P3_ADD_515_U78 , P3_U4302 );
nand NAND2_4385 ( P3_U6194 , P3_ADD_494_U78 , P3_U2356 );
nand NAND2_4386 ( P3_U6195 , P3_ADD_476_U78 , P3_U4303 );
nand NAND2_4387 ( P3_U6196 , P3_ADD_441_U78 , P3_U4304 );
nand NAND2_4388 ( P3_U6197 , P3_ADD_405_U77 , P3_U4305 );
nand NAND2_4389 ( P3_U6198 , P3_ADD_394_U77 , P3_U2357 );
nand NAND2_4390 ( P3_U6199 , P3_ADD_385_U81 , P3_U2358 );
nand NAND2_4391 ( P3_U6200 , P3_ADD_380_U81 , P3_U2359 );
nand NAND2_4392 ( P3_U6201 , P3_ADD_349_U81 , P3_U4306 );
nand NAND2_4393 ( P3_U6202 , P3_ADD_344_U81 , P3_U2362 );
nand NAND2_4394 ( P3_U6203 , P3_ADD_371_1212_U13 , P3_U2360 );
nand NAND2_4395 ( P3_U6204 , P3_U3872 , P3_U3867 );
nand NAND2_4396 ( P3_U6205 , P3_U2402 , P3_REIP_REG_23_ );
nand NAND2_4397 ( P3_U6206 , P3_U4318 , P3_U6204 );
nand NAND2_4398 ( P3_U6207 , P3_INSTADDRPOINTER_REG_23_ , P3_U5631 );
nand NAND2_4399 ( P3_U6208 , P3_ADD_360_1242_U79 , P3_U2395 );
nand NAND2_4400 ( P3_U6209 , P3_SUB_357_1258_U82 , P3_U2393 );
nand NAND2_4401 ( P3_U6210 , P3_ADD_558_U80 , P3_U3220 );
nand NAND2_4402 ( P3_U6211 , P3_ADD_553_U80 , P3_U4298 );
nand NAND2_4403 ( P3_U6212 , P3_ADD_547_U80 , P3_U4299 );
nand NAND2_4404 ( P3_U6213 , P3_ADD_541_U77 , P3_U4300 );
nand NAND2_4405 ( P3_U6214 , P3_ADD_536_U77 , P3_U4301 );
nand NAND2_4406 ( P3_U6215 , P3_ADD_531_U80 , P3_U2354 );
nand NAND2_4407 ( P3_U6216 , P3_ADD_526_U66 , P3_U2355 );
nand NAND2_4408 ( P3_U6217 , P3_ADD_515_U77 , P3_U4302 );
nand NAND2_4409 ( P3_U6218 , P3_ADD_494_U77 , P3_U2356 );
nand NAND2_4410 ( P3_U6219 , P3_ADD_476_U77 , P3_U4303 );
nand NAND2_4411 ( P3_U6220 , P3_ADD_441_U77 , P3_U4304 );
nand NAND2_4412 ( P3_U6221 , P3_ADD_405_U76 , P3_U4305 );
nand NAND2_4413 ( P3_U6222 , P3_ADD_394_U76 , P3_U2357 );
nand NAND2_4414 ( P3_U6223 , P3_ADD_385_U80 , P3_U2358 );
nand NAND2_4415 ( P3_U6224 , P3_ADD_380_U80 , P3_U2359 );
nand NAND2_4416 ( P3_U6225 , P3_ADD_349_U80 , P3_U4306 );
nand NAND2_4417 ( P3_U6226 , P3_ADD_344_U80 , P3_U2362 );
nand NAND2_4418 ( P3_U6227 , P3_ADD_371_1212_U81 , P3_U2360 );
nand NAND2_4419 ( P3_U6228 , P3_U3882 , P3_U3877 );
nand NAND2_4420 ( P3_U6229 , P3_U2402 , P3_REIP_REG_24_ );
nand NAND2_4421 ( P3_U6230 , P3_U4318 , P3_U6228 );
nand NAND2_4422 ( P3_U6231 , P3_INSTADDRPOINTER_REG_24_ , P3_U5631 );
nand NAND2_4423 ( P3_U6232 , P3_ADD_360_1242_U13 , P3_U2395 );
nand NAND2_4424 ( P3_U6233 , P3_SUB_357_1258_U81 , P3_U2393 );
nand NAND2_4425 ( P3_U6234 , P3_ADD_558_U79 , P3_U3220 );
nand NAND2_4426 ( P3_U6235 , P3_ADD_553_U79 , P3_U4298 );
nand NAND2_4427 ( P3_U6236 , P3_ADD_547_U79 , P3_U4299 );
nand NAND2_4428 ( P3_U6237 , P3_ADD_541_U76 , P3_U4300 );
nand NAND2_4429 ( P3_U6238 , P3_ADD_536_U76 , P3_U4301 );
nand NAND2_4430 ( P3_U6239 , P3_ADD_531_U79 , P3_U2354 );
nand NAND2_4431 ( P3_U6240 , P3_ADD_526_U65 , P3_U2355 );
nand NAND2_4432 ( P3_U6241 , P3_ADD_515_U76 , P3_U4302 );
nand NAND2_4433 ( P3_U6242 , P3_ADD_494_U76 , P3_U2356 );
nand NAND2_4434 ( P3_U6243 , P3_ADD_476_U76 , P3_U4303 );
nand NAND2_4435 ( P3_U6244 , P3_ADD_441_U76 , P3_U4304 );
nand NAND2_4436 ( P3_U6245 , P3_ADD_405_U75 , P3_U4305 );
nand NAND2_4437 ( P3_U6246 , P3_ADD_394_U75 , P3_U2357 );
nand NAND2_4438 ( P3_U6247 , P3_ADD_385_U79 , P3_U2358 );
nand NAND2_4439 ( P3_U6248 , P3_ADD_380_U79 , P3_U2359 );
nand NAND2_4440 ( P3_U6249 , P3_ADD_349_U79 , P3_U4306 );
nand NAND2_4441 ( P3_U6250 , P3_ADD_344_U79 , P3_U2362 );
nand NAND2_4442 ( P3_U6251 , P3_ADD_371_1212_U14 , P3_U2360 );
nand NAND2_4443 ( P3_U6252 , P3_U3892 , P3_U3887 );
nand NAND2_4444 ( P3_U6253 , P3_U2402 , P3_REIP_REG_25_ );
nand NAND2_4445 ( P3_U6254 , P3_U4318 , P3_U6252 );
nand NAND2_4446 ( P3_U6255 , P3_INSTADDRPOINTER_REG_25_ , P3_U5631 );
nand NAND2_4447 ( P3_U6256 , P3_ADD_360_1242_U14 , P3_U2395 );
nand NAND2_4448 ( P3_U6257 , P3_SUB_357_1258_U18 , P3_U2393 );
nand NAND2_4449 ( P3_U6258 , P3_ADD_558_U78 , P3_U3220 );
nand NAND2_4450 ( P3_U6259 , P3_ADD_553_U78 , P3_U4298 );
nand NAND2_4451 ( P3_U6260 , P3_ADD_547_U78 , P3_U4299 );
nand NAND2_4452 ( P3_U6261 , P3_ADD_541_U75 , P3_U4300 );
nand NAND2_4453 ( P3_U6262 , P3_ADD_536_U75 , P3_U4301 );
nand NAND2_4454 ( P3_U6263 , P3_ADD_531_U78 , P3_U2354 );
nand NAND2_4455 ( P3_U6264 , P3_ADD_526_U64 , P3_U2355 );
nand NAND2_4456 ( P3_U6265 , P3_ADD_515_U75 , P3_U4302 );
nand NAND2_4457 ( P3_U6266 , P3_ADD_494_U75 , P3_U2356 );
nand NAND2_4458 ( P3_U6267 , P3_ADD_476_U75 , P3_U4303 );
nand NAND2_4459 ( P3_U6268 , P3_ADD_441_U75 , P3_U4304 );
nand NAND2_4460 ( P3_U6269 , P3_ADD_405_U74 , P3_U4305 );
nand NAND2_4461 ( P3_U6270 , P3_ADD_394_U74 , P3_U2357 );
nand NAND2_4462 ( P3_U6271 , P3_ADD_385_U78 , P3_U2358 );
nand NAND2_4463 ( P3_U6272 , P3_ADD_380_U78 , P3_U2359 );
nand NAND2_4464 ( P3_U6273 , P3_ADD_349_U78 , P3_U4306 );
nand NAND2_4465 ( P3_U6274 , P3_ADD_344_U78 , P3_U2362 );
nand NAND2_4466 ( P3_U6275 , P3_ADD_371_1212_U15 , P3_U2360 );
nand NAND5_4467 ( P3_U6276 , P3_U3894 , P3_U6258 , P3_U3895 , P3_U3897 , P3_U3902 );
nand NAND2_4468 ( P3_U6277 , P3_U2402 , P3_REIP_REG_26_ );
nand NAND2_4469 ( P3_U6278 , P3_U4318 , P3_U6276 );
nand NAND2_4470 ( P3_U6279 , P3_INSTADDRPOINTER_REG_26_ , P3_U5631 );
nand NAND2_4471 ( P3_U6280 , P3_ADD_360_1242_U78 , P3_U2395 );
nand NAND2_4472 ( P3_U6281 , P3_SUB_357_1258_U80 , P3_U2393 );
nand NAND2_4473 ( P3_U6282 , P3_ADD_558_U77 , P3_U3220 );
nand NAND2_4474 ( P3_U6283 , P3_ADD_553_U77 , P3_U4298 );
nand NAND2_4475 ( P3_U6284 , P3_ADD_547_U77 , P3_U4299 );
nand NAND2_4476 ( P3_U6285 , P3_ADD_541_U74 , P3_U4300 );
nand NAND2_4477 ( P3_U6286 , P3_ADD_536_U74 , P3_U4301 );
nand NAND2_4478 ( P3_U6287 , P3_ADD_531_U77 , P3_U2354 );
nand NAND2_4479 ( P3_U6288 , P3_ADD_526_U63 , P3_U2355 );
nand NAND2_4480 ( P3_U6289 , P3_ADD_515_U74 , P3_U4302 );
nand NAND2_4481 ( P3_U6290 , P3_ADD_494_U74 , P3_U2356 );
nand NAND2_4482 ( P3_U6291 , P3_ADD_476_U74 , P3_U4303 );
nand NAND2_4483 ( P3_U6292 , P3_ADD_441_U74 , P3_U4304 );
nand NAND2_4484 ( P3_U6293 , P3_ADD_405_U73 , P3_U4305 );
nand NAND2_4485 ( P3_U6294 , P3_ADD_394_U73 , P3_U2357 );
nand NAND2_4486 ( P3_U6295 , P3_ADD_385_U77 , P3_U2358 );
nand NAND2_4487 ( P3_U6296 , P3_ADD_380_U77 , P3_U2359 );
nand NAND2_4488 ( P3_U6297 , P3_ADD_349_U77 , P3_U4306 );
nand NAND2_4489 ( P3_U6298 , P3_ADD_344_U77 , P3_U2362 );
nand NAND2_4490 ( P3_U6299 , P3_ADD_371_1212_U80 , P3_U2360 );
nand NAND5_4491 ( P3_U6300 , P3_U3903 , P3_U6282 , P3_U3904 , P3_U3906 , P3_U3911 );
nand NAND2_4492 ( P3_U6301 , P3_U2402 , P3_REIP_REG_27_ );
nand NAND2_4493 ( P3_U6302 , P3_U4318 , P3_U6300 );
nand NAND2_4494 ( P3_U6303 , P3_INSTADDRPOINTER_REG_27_ , P3_U5631 );
nand NAND2_4495 ( P3_U6304 , P3_ADD_360_1242_U15 , P3_U2395 );
nand NAND2_4496 ( P3_U6305 , P3_SUB_357_1258_U19 , P3_U2393 );
nand NAND2_4497 ( P3_U6306 , P3_ADD_558_U76 , P3_U3220 );
nand NAND2_4498 ( P3_U6307 , P3_ADD_553_U76 , P3_U4298 );
nand NAND2_4499 ( P3_U6308 , P3_ADD_547_U76 , P3_U4299 );
nand NAND2_4500 ( P3_U6309 , P3_ADD_541_U73 , P3_U4300 );
nand NAND2_4501 ( P3_U6310 , P3_ADD_536_U73 , P3_U4301 );
nand NAND2_4502 ( P3_U6311 , P3_ADD_531_U76 , P3_U2354 );
nand NAND2_4503 ( P3_U6312 , P3_ADD_526_U62 , P3_U2355 );
nand NAND2_4504 ( P3_U6313 , P3_ADD_515_U73 , P3_U4302 );
nand NAND2_4505 ( P3_U6314 , P3_ADD_494_U73 , P3_U2356 );
nand NAND2_4506 ( P3_U6315 , P3_ADD_476_U73 , P3_U4303 );
nand NAND2_4507 ( P3_U6316 , P3_ADD_441_U73 , P3_U4304 );
nand NAND2_4508 ( P3_U6317 , P3_ADD_405_U72 , P3_U4305 );
nand NAND2_4509 ( P3_U6318 , P3_ADD_394_U72 , P3_U2357 );
nand NAND2_4510 ( P3_U6319 , P3_ADD_385_U76 , P3_U2358 );
nand NAND2_4511 ( P3_U6320 , P3_ADD_380_U76 , P3_U2359 );
nand NAND2_4512 ( P3_U6321 , P3_ADD_349_U76 , P3_U4306 );
nand NAND2_4513 ( P3_U6322 , P3_ADD_344_U76 , P3_U2362 );
nand NAND2_4514 ( P3_U6323 , P3_ADD_371_1212_U16 , P3_U2360 );
nand NAND5_4515 ( P3_U6324 , P3_U3912 , P3_U6306 , P3_U3913 , P3_U3915 , P3_U3920 );
nand NAND2_4516 ( P3_U6325 , P3_U2402 , P3_REIP_REG_28_ );
nand NAND2_4517 ( P3_U6326 , P3_U4318 , P3_U6324 );
nand NAND2_4518 ( P3_U6327 , P3_INSTADDRPOINTER_REG_28_ , P3_U5631 );
nand NAND2_4519 ( P3_U6328 , P3_ADD_360_1242_U16 , P3_U2395 );
nand NAND2_4520 ( P3_U6329 , P3_SUB_357_1258_U79 , P3_U2393 );
nand NAND2_4521 ( P3_U6330 , P3_ADD_558_U75 , P3_U3220 );
nand NAND2_4522 ( P3_U6331 , P3_ADD_553_U75 , P3_U4298 );
nand NAND2_4523 ( P3_U6332 , P3_ADD_547_U75 , P3_U4299 );
nand NAND2_4524 ( P3_U6333 , P3_ADD_541_U72 , P3_U4300 );
nand NAND2_4525 ( P3_U6334 , P3_ADD_536_U72 , P3_U4301 );
nand NAND2_4526 ( P3_U6335 , P3_ADD_531_U75 , P3_U2354 );
nand NAND2_4527 ( P3_U6336 , P3_ADD_526_U61 , P3_U2355 );
nand NAND2_4528 ( P3_U6337 , P3_ADD_515_U72 , P3_U4302 );
nand NAND2_4529 ( P3_U6338 , P3_ADD_494_U72 , P3_U2356 );
nand NAND2_4530 ( P3_U6339 , P3_ADD_476_U72 , P3_U4303 );
nand NAND2_4531 ( P3_U6340 , P3_ADD_441_U72 , P3_U4304 );
nand NAND2_4532 ( P3_U6341 , P3_ADD_405_U71 , P3_U4305 );
nand NAND2_4533 ( P3_U6342 , P3_ADD_394_U71 , P3_U2357 );
nand NAND2_4534 ( P3_U6343 , P3_ADD_385_U75 , P3_U2358 );
nand NAND2_4535 ( P3_U6344 , P3_ADD_380_U75 , P3_U2359 );
nand NAND2_4536 ( P3_U6345 , P3_ADD_349_U75 , P3_U4306 );
nand NAND2_4537 ( P3_U6346 , P3_ADD_344_U75 , P3_U2362 );
nand NAND2_4538 ( P3_U6347 , P3_ADD_371_1212_U17 , P3_U2360 );
nand NAND5_4539 ( P3_U6348 , P3_U3921 , P3_U6330 , P3_U3922 , P3_U3924 , P3_U3929 );
nand NAND2_4540 ( P3_U6349 , P3_U2402 , P3_REIP_REG_29_ );
nand NAND2_4541 ( P3_U6350 , P3_U4318 , P3_U6348 );
nand NAND2_4542 ( P3_U6351 , P3_INSTADDRPOINTER_REG_29_ , P3_U5631 );
nand NAND2_4543 ( P3_U6352 , P3_ADD_360_1242_U77 , P3_U2395 );
nand NAND2_4544 ( P3_U6353 , P3_SUB_357_1258_U77 , P3_U2393 );
nand NAND2_4545 ( P3_U6354 , P3_ADD_558_U73 , P3_U3220 );
nand NAND2_4546 ( P3_U6355 , P3_ADD_553_U73 , P3_U4298 );
nand NAND2_4547 ( P3_U6356 , P3_ADD_547_U73 , P3_U4299 );
nand NAND2_4548 ( P3_U6357 , P3_ADD_541_U70 , P3_U4300 );
nand NAND2_4549 ( P3_U6358 , P3_ADD_536_U70 , P3_U4301 );
nand NAND2_4550 ( P3_U6359 , P3_ADD_531_U73 , P3_U2354 );
nand NAND2_4551 ( P3_U6360 , P3_ADD_526_U59 , P3_U2355 );
nand NAND2_4552 ( P3_U6361 , P3_ADD_515_U70 , P3_U4302 );
nand NAND2_4553 ( P3_U6362 , P3_ADD_494_U70 , P3_U2356 );
nand NAND2_4554 ( P3_U6363 , P3_ADD_476_U70 , P3_U4303 );
nand NAND2_4555 ( P3_U6364 , P3_ADD_441_U70 , P3_U4304 );
nand NAND2_4556 ( P3_U6365 , P3_ADD_405_U70 , P3_U4305 );
nand NAND2_4557 ( P3_U6366 , P3_ADD_394_U70 , P3_U2357 );
nand NAND2_4558 ( P3_U6367 , P3_ADD_385_U73 , P3_U2358 );
nand NAND2_4559 ( P3_U6368 , P3_ADD_380_U73 , P3_U2359 );
nand NAND2_4560 ( P3_U6369 , P3_ADD_349_U73 , P3_U4306 );
nand NAND2_4561 ( P3_U6370 , P3_ADD_344_U73 , P3_U2362 );
nand NAND2_4562 ( P3_U6371 , P3_ADD_371_1212_U79 , P3_U2360 );
nand NAND5_4563 ( P3_U6372 , P3_U3930 , P3_U6354 , P3_U3931 , P3_U3933 , P3_U3938 );
nand NAND2_4564 ( P3_U6373 , P3_U2402 , P3_REIP_REG_30_ );
nand NAND2_4565 ( P3_U6374 , P3_U4318 , P3_U6372 );
nand NAND2_4566 ( P3_U6375 , P3_INSTADDRPOINTER_REG_30_ , P3_U5631 );
nand NAND2_4567 ( P3_U6376 , P3_ADD_360_1242_U90 , P3_U2395 );
nand NAND2_4568 ( P3_U6377 , P3_SUB_357_1258_U20 , P3_U2393 );
nand NAND2_4569 ( P3_U6378 , P3_ADD_558_U72 , P3_U3220 );
nand NAND2_4570 ( P3_U6379 , P3_ADD_553_U72 , P3_U4298 );
nand NAND2_4571 ( P3_U6380 , P3_ADD_547_U72 , P3_U4299 );
nand NAND2_4572 ( P3_U6381 , P3_ADD_541_U69 , P3_U4300 );
nand NAND2_4573 ( P3_U6382 , P3_ADD_536_U69 , P3_U4301 );
nand NAND2_4574 ( P3_U6383 , P3_ADD_531_U72 , P3_U2354 );
nand NAND2_4575 ( P3_U6384 , P3_ADD_526_U58 , P3_U2355 );
nand NAND2_4576 ( P3_U6385 , P3_ADD_515_U69 , P3_U4302 );
nand NAND2_4577 ( P3_U6386 , P3_ADD_494_U69 , P3_U2356 );
nand NAND2_4578 ( P3_U6387 , P3_ADD_476_U69 , P3_U4303 );
nand NAND2_4579 ( P3_U6388 , P3_ADD_441_U69 , P3_U4304 );
nand NAND2_4580 ( P3_U6389 , P3_ADD_405_U69 , P3_U4305 );
nand NAND2_4581 ( P3_U6390 , P3_ADD_394_U69 , P3_U2357 );
nand NAND2_4582 ( P3_U6391 , P3_ADD_385_U72 , P3_U2358 );
nand NAND2_4583 ( P3_U6392 , P3_ADD_380_U72 , P3_U2359 );
nand NAND2_4584 ( P3_U6393 , P3_ADD_349_U72 , P3_U4306 );
nand NAND2_4585 ( P3_U6394 , P3_ADD_344_U72 , P3_U2362 );
nand NAND2_4586 ( P3_U6395 , P3_ADD_371_1212_U92 , P3_U2360 );
nand NAND2_4587 ( P3_U6396 , P3_U3950 , P3_U3945 );
nand NAND2_4588 ( P3_U6397 , P3_U2402 , P3_REIP_REG_31_ );
nand NAND2_4589 ( P3_U6398 , P3_INSTADDRPOINTER_REG_31_ , P3_U5631 );
nand NAND2_4590 ( P3_U6399 , P3_GTE_355_U6 , P3_U2361 );
nand NAND2_4591 ( P3_U6400 , P3_GTE_370_U6 , P3_U2360 );
nand NAND2_4592 ( P3_U6401 , P3_U6400 , P3_U6399 );
nand NAND2_4593 ( P3_U6402 , P3_U2390 , P3_U6401 );
nand NAND2_4594 ( P3_U6403 , P3_U3234 , P3_U3121 );
not NOT1_4595 ( P3_U6404 , P3_U3249 );
nand NAND2_4596 ( P3_U6405 , P3_PHYADDRPOINTER_REG_0_ , P3_U2398 );
nand NAND2_4597 ( P3_U6406 , P3_PHYADDRPOINTER_REG_0_ , P3_U2397 );
nand NAND2_4598 ( P3_U6407 , P3_U2396 , P3_ADD_360_1242_U85 );
nand NAND2_4599 ( P3_U6408 , P3_U2394 , P3_SUB_357_1258_U69 );
nand NAND2_4600 ( P3_U6409 , P3_U2389 , P3_REIP_REG_0_ );
nand NAND2_4601 ( P3_U6410 , P3_PHYADDRPOINTER_REG_0_ , P3_U2388 );
nand NAND2_4602 ( P3_U6411 , P3_U2387 , P3_ADD_371_1212_U87 );
nand NAND2_4603 ( P3_U6412 , P3_PHYADDRPOINTER_REG_0_ , P3_U6404 );
nand NAND2_4604 ( P3_U6413 , P3_ADD_318_U4 , P3_U2398 );
nand NAND2_4605 ( P3_U6414 , P3_PHYADDRPOINTER_REG_1_ , P3_U2397 );
nand NAND2_4606 ( P3_U6415 , P3_U2396 , P3_ADD_360_1242_U19 );
nand NAND2_4607 ( P3_U6416 , P3_U2394 , P3_SUB_357_1258_U21 );
nand NAND2_4608 ( P3_U6417 , P3_U2389 , P3_REIP_REG_1_ );
nand NAND2_4609 ( P3_U6418 , P3_ADD_339_U4 , P3_U2388 );
nand NAND2_4610 ( P3_U6419 , P3_U2387 , P3_ADD_371_1212_U20 );
nand NAND2_4611 ( P3_U6420 , P3_PHYADDRPOINTER_REG_1_ , P3_U6404 );
nand NAND2_4612 ( P3_U6421 , P3_ADD_318_U71 , P3_U2398 );
nand NAND2_4613 ( P3_U6422 , P3_ADD_315_U4 , P3_U2397 );
nand NAND2_4614 ( P3_U6423 , P3_U2396 , P3_ADD_360_1242_U91 );
nand NAND2_4615 ( P3_U6424 , P3_U2394 , P3_SUB_357_1258_U78 );
nand NAND2_4616 ( P3_U6425 , P3_U2389 , P3_REIP_REG_2_ );
nand NAND2_4617 ( P3_U6426 , P3_ADD_339_U71 , P3_U2388 );
nand NAND2_4618 ( P3_U6427 , P3_U2387 , P3_ADD_371_1212_U93 );
nand NAND2_4619 ( P3_U6428 , P3_PHYADDRPOINTER_REG_2_ , P3_U6404 );
nand NAND2_4620 ( P3_U6429 , P3_ADD_318_U68 , P3_U2398 );
nand NAND2_4621 ( P3_U6430 , P3_ADD_315_U66 , P3_U2397 );
nand NAND2_4622 ( P3_U6431 , P3_U2396 , P3_ADD_360_1242_U17 );
nand NAND2_4623 ( P3_U6432 , P3_U2394 , P3_SUB_357_1258_U76 );
nand NAND2_4624 ( P3_U6433 , P3_U2389 , P3_REIP_REG_3_ );
nand NAND2_4625 ( P3_U6434 , P3_ADD_339_U68 , P3_U2388 );
nand NAND2_4626 ( P3_U6435 , P3_U2387 , P3_ADD_371_1212_U18 );
nand NAND2_4627 ( P3_U6436 , P3_PHYADDRPOINTER_REG_3_ , P3_U6404 );
nand NAND2_4628 ( P3_U6437 , P3_ADD_318_U67 , P3_U2398 );
nand NAND2_4629 ( P3_U6438 , P3_ADD_315_U65 , P3_U2397 );
nand NAND2_4630 ( P3_U6439 , P3_U2396 , P3_ADD_360_1242_U18 );
nand NAND2_4631 ( P3_U6440 , P3_U2394 , P3_SUB_357_1258_U75 );
nand NAND2_4632 ( P3_U6441 , P3_U2389 , P3_REIP_REG_4_ );
nand NAND2_4633 ( P3_U6442 , P3_ADD_339_U67 , P3_U2388 );
nand NAND2_4634 ( P3_U6443 , P3_U2387 , P3_ADD_371_1212_U91 );
nand NAND2_4635 ( P3_U6444 , P3_PHYADDRPOINTER_REG_4_ , P3_U6404 );
nand NAND2_4636 ( P3_U6445 , P3_ADD_318_U66 , P3_U2398 );
nand NAND2_4637 ( P3_U6446 , P3_ADD_315_U64 , P3_U2397 );
nand NAND2_4638 ( P3_U6447 , P3_U2396 , P3_ADD_360_1242_U89 );
nand NAND2_4639 ( P3_U6448 , P3_U2394 , P3_SUB_357_1258_U74 );
nand NAND2_4640 ( P3_U6449 , P3_U2389 , P3_REIP_REG_5_ );
nand NAND2_4641 ( P3_U6450 , P3_ADD_339_U66 , P3_U2388 );
nand NAND2_4642 ( P3_U6451 , P3_U2387 , P3_ADD_371_1212_U19 );
nand NAND2_4643 ( P3_U6452 , P3_PHYADDRPOINTER_REG_5_ , P3_U6404 );
nand NAND2_4644 ( P3_U6453 , P3_ADD_318_U65 , P3_U2398 );
nand NAND2_4645 ( P3_U6454 , P3_ADD_315_U63 , P3_U2397 );
nand NAND2_4646 ( P3_U6455 , P3_U2396 , P3_ADD_360_1242_U88 );
nand NAND2_4647 ( P3_U6456 , P3_U2394 , P3_SUB_357_1258_U73 );
nand NAND2_4648 ( P3_U6457 , P3_U2389 , P3_REIP_REG_6_ );
nand NAND2_4649 ( P3_U6458 , P3_ADD_339_U65 , P3_U2388 );
nand NAND2_4650 ( P3_U6459 , P3_U2387 , P3_ADD_371_1212_U90 );
nand NAND2_4651 ( P3_U6460 , P3_PHYADDRPOINTER_REG_6_ , P3_U6404 );
nand NAND2_4652 ( P3_U6461 , P3_ADD_318_U64 , P3_U2398 );
nand NAND2_4653 ( P3_U6462 , P3_ADD_315_U62 , P3_U2397 );
nand NAND2_4654 ( P3_U6463 , P3_U2396 , P3_ADD_360_1242_U87 );
nand NAND2_4655 ( P3_U6464 , P3_U2394 , P3_SUB_357_1258_U72 );
nand NAND2_4656 ( P3_U6465 , P3_U2389 , P3_REIP_REG_7_ );
nand NAND2_4657 ( P3_U6466 , P3_ADD_339_U64 , P3_U2388 );
nand NAND2_4658 ( P3_U6467 , P3_U2387 , P3_ADD_371_1212_U89 );
nand NAND2_4659 ( P3_U6468 , P3_PHYADDRPOINTER_REG_7_ , P3_U6404 );
nand NAND2_4660 ( P3_U6469 , P3_ADD_318_U63 , P3_U2398 );
nand NAND2_4661 ( P3_U6470 , P3_ADD_315_U61 , P3_U2397 );
nand NAND2_4662 ( P3_U6471 , P3_U2396 , P3_ADD_360_1242_U86 );
nand NAND2_4663 ( P3_U6472 , P3_U2394 , P3_SUB_357_1258_U71 );
nand NAND2_4664 ( P3_U6473 , P3_U2389 , P3_REIP_REG_8_ );
nand NAND2_4665 ( P3_U6474 , P3_ADD_339_U63 , P3_U2388 );
nand NAND2_4666 ( P3_U6475 , P3_U2387 , P3_ADD_371_1212_U88 );
nand NAND2_4667 ( P3_U6476 , P3_PHYADDRPOINTER_REG_8_ , P3_U6404 );
nand NAND2_4668 ( P3_U6477 , P3_ADD_318_U62 , P3_U2398 );
nand NAND2_4669 ( P3_U6478 , P3_ADD_315_U60 , P3_U2397 );
nand NAND2_4670 ( P3_U6479 , P3_U2396 , P3_ADD_360_1242_U106 );
nand NAND2_4671 ( P3_U6480 , P3_U2394 , P3_SUB_357_1258_U70 );
nand NAND2_4672 ( P3_U6481 , P3_U2389 , P3_REIP_REG_9_ );
nand NAND2_4673 ( P3_U6482 , P3_ADD_339_U62 , P3_U2388 );
nand NAND2_4674 ( P3_U6483 , P3_U2387 , P3_ADD_371_1212_U109 );
nand NAND2_4675 ( P3_U6484 , P3_PHYADDRPOINTER_REG_9_ , P3_U6404 );
nand NAND2_4676 ( P3_U6485 , P3_ADD_318_U91 , P3_U2398 );
nand NAND2_4677 ( P3_U6486 , P3_ADD_315_U88 , P3_U2397 );
nand NAND2_4678 ( P3_U6487 , P3_U2396 , P3_ADD_360_1242_U4 );
nand NAND2_4679 ( P3_U6488 , P3_U2394 , P3_SUB_357_1258_U93 );
nand NAND2_4680 ( P3_U6489 , P3_U2389 , P3_REIP_REG_10_ );
nand NAND2_4681 ( P3_U6490 , P3_ADD_339_U91 , P3_U2388 );
nand NAND2_4682 ( P3_U6491 , P3_U2387 , P3_ADD_371_1212_U5 );
nand NAND2_4683 ( P3_U6492 , P3_PHYADDRPOINTER_REG_10_ , P3_U6404 );
nand NAND2_4684 ( P3_U6493 , P3_ADD_318_U90 , P3_U2398 );
nand NAND2_4685 ( P3_U6494 , P3_ADD_315_U87 , P3_U2397 );
nand NAND2_4686 ( P3_U6495 , P3_U2396 , P3_ADD_360_1242_U84 );
nand NAND2_4687 ( P3_U6496 , P3_U2394 , P3_SUB_357_1258_U92 );
nand NAND2_4688 ( P3_U6497 , P3_U2389 , P3_REIP_REG_11_ );
nand NAND2_4689 ( P3_U6498 , P3_ADD_339_U90 , P3_U2388 );
nand NAND2_4690 ( P3_U6499 , P3_U2387 , P3_ADD_371_1212_U86 );
nand NAND2_4691 ( P3_U6500 , P3_PHYADDRPOINTER_REG_11_ , P3_U6404 );
nand NAND2_4692 ( P3_U6501 , P3_ADD_318_U89 , P3_U2398 );
nand NAND2_4693 ( P3_U6502 , P3_ADD_315_U86 , P3_U2397 );
nand NAND2_4694 ( P3_U6503 , P3_U2396 , P3_ADD_360_1242_U5 );
nand NAND2_4695 ( P3_U6504 , P3_U2394 , P3_SUB_357_1258_U91 );
nand NAND2_4696 ( P3_U6505 , P3_U2389 , P3_REIP_REG_12_ );
nand NAND2_4697 ( P3_U6506 , P3_ADD_339_U89 , P3_U2388 );
nand NAND2_4698 ( P3_U6507 , P3_U2387 , P3_ADD_371_1212_U6 );
nand NAND2_4699 ( P3_U6508 , P3_PHYADDRPOINTER_REG_12_ , P3_U6404 );
nand NAND2_4700 ( P3_U6509 , P3_ADD_318_U88 , P3_U2398 );
nand NAND2_4701 ( P3_U6510 , P3_ADD_315_U85 , P3_U2397 );
nand NAND2_4702 ( P3_U6511 , P3_U2396 , P3_ADD_360_1242_U6 );
nand NAND2_4703 ( P3_U6512 , P3_U2394 , P3_SUB_357_1258_U15 );
nand NAND2_4704 ( P3_U6513 , P3_U2389 , P3_REIP_REG_13_ );
nand NAND2_4705 ( P3_U6514 , P3_ADD_339_U88 , P3_U2388 );
nand NAND2_4706 ( P3_U6515 , P3_U2387 , P3_ADD_371_1212_U7 );
nand NAND2_4707 ( P3_U6516 , P3_PHYADDRPOINTER_REG_13_ , P3_U6404 );
nand NAND2_4708 ( P3_U6517 , P3_ADD_318_U87 , P3_U2398 );
nand NAND2_4709 ( P3_U6518 , P3_ADD_315_U84 , P3_U2397 );
nand NAND2_4710 ( P3_U6519 , P3_U2396 , P3_ADD_360_1242_U83 );
nand NAND2_4711 ( P3_U6520 , P3_U2394 , P3_SUB_357_1258_U90 );
nand NAND2_4712 ( P3_U6521 , P3_U2389 , P3_REIP_REG_14_ );
nand NAND2_4713 ( P3_U6522 , P3_ADD_339_U87 , P3_U2388 );
nand NAND2_4714 ( P3_U6523 , P3_U2387 , P3_ADD_371_1212_U85 );
nand NAND2_4715 ( P3_U6524 , P3_PHYADDRPOINTER_REG_14_ , P3_U6404 );
nand NAND2_4716 ( P3_U6525 , P3_ADD_318_U86 , P3_U2398 );
nand NAND2_4717 ( P3_U6526 , P3_ADD_315_U83 , P3_U2397 );
nand NAND2_4718 ( P3_U6527 , P3_U2396 , P3_ADD_360_1242_U7 );
nand NAND2_4719 ( P3_U6528 , P3_U2394 , P3_SUB_357_1258_U89 );
nand NAND2_4720 ( P3_U6529 , P3_U2389 , P3_REIP_REG_15_ );
nand NAND2_4721 ( P3_U6530 , P3_ADD_339_U86 , P3_U2388 );
nand NAND2_4722 ( P3_U6531 , P3_U2387 , P3_ADD_371_1212_U8 );
nand NAND2_4723 ( P3_U6532 , P3_PHYADDRPOINTER_REG_15_ , P3_U6404 );
nand NAND2_4724 ( P3_U6533 , P3_ADD_318_U85 , P3_U2398 );
nand NAND2_4725 ( P3_U6534 , P3_ADD_315_U82 , P3_U2397 );
nand NAND2_4726 ( P3_U6535 , P3_U2396 , P3_ADD_360_1242_U82 );
nand NAND2_4727 ( P3_U6536 , P3_U2394 , P3_SUB_357_1258_U88 );
nand NAND2_4728 ( P3_U6537 , P3_U2389 , P3_REIP_REG_16_ );
nand NAND2_4729 ( P3_U6538 , P3_ADD_339_U85 , P3_U2388 );
nand NAND2_4730 ( P3_U6539 , P3_U2387 , P3_ADD_371_1212_U84 );
nand NAND2_4731 ( P3_U6540 , P3_PHYADDRPOINTER_REG_16_ , P3_U6404 );
nand NAND2_4732 ( P3_U6541 , P3_ADD_318_U84 , P3_U2398 );
nand NAND2_4733 ( P3_U6542 , P3_ADD_315_U81 , P3_U2397 );
nand NAND2_4734 ( P3_U6543 , P3_U2396 , P3_ADD_360_1242_U8 );
nand NAND2_4735 ( P3_U6544 , P3_U2394 , P3_SUB_357_1258_U16 );
nand NAND2_4736 ( P3_U6545 , P3_U2389 , P3_REIP_REG_17_ );
nand NAND2_4737 ( P3_U6546 , P3_ADD_339_U84 , P3_U2388 );
nand NAND2_4738 ( P3_U6547 , P3_U2387 , P3_ADD_371_1212_U9 );
nand NAND2_4739 ( P3_U6548 , P3_PHYADDRPOINTER_REG_17_ , P3_U6404 );
nand NAND2_4740 ( P3_U6549 , P3_ADD_318_U83 , P3_U2398 );
nand NAND2_4741 ( P3_U6550 , P3_ADD_315_U80 , P3_U2397 );
nand NAND2_4742 ( P3_U6551 , P3_U2396 , P3_ADD_360_1242_U81 );
nand NAND2_4743 ( P3_U6552 , P3_U2394 , P3_SUB_357_1258_U87 );
nand NAND2_4744 ( P3_U6553 , P3_U2389 , P3_REIP_REG_18_ );
nand NAND2_4745 ( P3_U6554 , P3_ADD_339_U83 , P3_U2388 );
nand NAND2_4746 ( P3_U6555 , P3_U2387 , P3_ADD_371_1212_U83 );
nand NAND2_4747 ( P3_U6556 , P3_PHYADDRPOINTER_REG_18_ , P3_U6404 );
nand NAND2_4748 ( P3_U6557 , P3_ADD_318_U82 , P3_U2398 );
nand NAND2_4749 ( P3_U6558 , P3_ADD_315_U79 , P3_U2397 );
nand NAND2_4750 ( P3_U6559 , P3_U2396 , P3_ADD_360_1242_U9 );
nand NAND2_4751 ( P3_U6560 , P3_U2394 , P3_SUB_357_1258_U86 );
nand NAND2_4752 ( P3_U6561 , P3_U2389 , P3_REIP_REG_19_ );
nand NAND2_4753 ( P3_U6562 , P3_ADD_339_U82 , P3_U2388 );
nand NAND2_4754 ( P3_U6563 , P3_U2387 , P3_ADD_371_1212_U10 );
nand NAND2_4755 ( P3_U6564 , P3_PHYADDRPOINTER_REG_19_ , P3_U6404 );
nand NAND2_4756 ( P3_U6565 , P3_ADD_318_U81 , P3_U2398 );
nand NAND2_4757 ( P3_U6566 , P3_ADD_315_U78 , P3_U2397 );
nand NAND2_4758 ( P3_U6567 , P3_U2396 , P3_ADD_360_1242_U10 );
nand NAND2_4759 ( P3_U6568 , P3_U2394 , P3_SUB_357_1258_U17 );
nand NAND2_4760 ( P3_U6569 , P3_U2389 , P3_REIP_REG_20_ );
nand NAND2_4761 ( P3_U6570 , P3_ADD_339_U81 , P3_U2388 );
nand NAND2_4762 ( P3_U6571 , P3_U2387 , P3_ADD_371_1212_U11 );
nand NAND2_4763 ( P3_U6572 , P3_PHYADDRPOINTER_REG_20_ , P3_U6404 );
nand NAND2_4764 ( P3_U6573 , P3_ADD_318_U80 , P3_U2398 );
nand NAND2_4765 ( P3_U6574 , P3_ADD_315_U77 , P3_U2397 );
nand NAND2_4766 ( P3_U6575 , P3_U2396 , P3_ADD_360_1242_U11 );
nand NAND2_4767 ( P3_U6576 , P3_U2394 , P3_SUB_357_1258_U85 );
nand NAND2_4768 ( P3_U6577 , P3_U2389 , P3_REIP_REG_21_ );
nand NAND2_4769 ( P3_U6578 , P3_ADD_339_U80 , P3_U2388 );
nand NAND2_4770 ( P3_U6579 , P3_U2387 , P3_ADD_371_1212_U12 );
nand NAND2_4771 ( P3_U6580 , P3_PHYADDRPOINTER_REG_21_ , P3_U6404 );
nand NAND2_4772 ( P3_U6581 , P3_ADD_318_U79 , P3_U2398 );
nand NAND2_4773 ( P3_U6582 , P3_ADD_315_U76 , P3_U2397 );
nand NAND2_4774 ( P3_U6583 , P3_U2396 , P3_ADD_360_1242_U80 );
nand NAND2_4775 ( P3_U6584 , P3_U2394 , P3_SUB_357_1258_U84 );
nand NAND2_4776 ( P3_U6585 , P3_U2389 , P3_REIP_REG_22_ );
nand NAND2_4777 ( P3_U6586 , P3_ADD_339_U79 , P3_U2388 );
nand NAND2_4778 ( P3_U6587 , P3_U2387 , P3_ADD_371_1212_U82 );
nand NAND2_4779 ( P3_U6588 , P3_PHYADDRPOINTER_REG_22_ , P3_U6404 );
nand NAND2_4780 ( P3_U6589 , P3_ADD_318_U78 , P3_U2398 );
nand NAND2_4781 ( P3_U6590 , P3_ADD_315_U75 , P3_U2397 );
nand NAND2_4782 ( P3_U6591 , P3_U2396 , P3_ADD_360_1242_U12 );
nand NAND2_4783 ( P3_U6592 , P3_U2394 , P3_SUB_357_1258_U83 );
nand NAND2_4784 ( P3_U6593 , P3_U2389 , P3_REIP_REG_23_ );
nand NAND2_4785 ( P3_U6594 , P3_ADD_339_U78 , P3_U2388 );
nand NAND2_4786 ( P3_U6595 , P3_U2387 , P3_ADD_371_1212_U13 );
nand NAND2_4787 ( P3_U6596 , P3_PHYADDRPOINTER_REG_23_ , P3_U6404 );
nand NAND2_4788 ( P3_U6597 , P3_ADD_318_U77 , P3_U2398 );
nand NAND2_4789 ( P3_U6598 , P3_ADD_315_U74 , P3_U2397 );
nand NAND2_4790 ( P3_U6599 , P3_U2396 , P3_ADD_360_1242_U79 );
nand NAND2_4791 ( P3_U6600 , P3_U2394 , P3_SUB_357_1258_U82 );
nand NAND2_4792 ( P3_U6601 , P3_U2389 , P3_REIP_REG_24_ );
nand NAND2_4793 ( P3_U6602 , P3_ADD_339_U77 , P3_U2388 );
nand NAND2_4794 ( P3_U6603 , P3_U2387 , P3_ADD_371_1212_U81 );
nand NAND2_4795 ( P3_U6604 , P3_PHYADDRPOINTER_REG_24_ , P3_U6404 );
nand NAND2_4796 ( P3_U6605 , P3_ADD_318_U76 , P3_U2398 );
nand NAND2_4797 ( P3_U6606 , P3_ADD_315_U73 , P3_U2397 );
nand NAND2_4798 ( P3_U6607 , P3_U2396 , P3_ADD_360_1242_U13 );
nand NAND2_4799 ( P3_U6608 , P3_U2394 , P3_SUB_357_1258_U81 );
nand NAND2_4800 ( P3_U6609 , P3_U2389 , P3_REIP_REG_25_ );
nand NAND2_4801 ( P3_U6610 , P3_ADD_339_U76 , P3_U2388 );
nand NAND2_4802 ( P3_U6611 , P3_U2387 , P3_ADD_371_1212_U14 );
nand NAND2_4803 ( P3_U6612 , P3_PHYADDRPOINTER_REG_25_ , P3_U6404 );
nand NAND2_4804 ( P3_U6613 , P3_ADD_318_U75 , P3_U2398 );
nand NAND2_4805 ( P3_U6614 , P3_ADD_315_U72 , P3_U2397 );
nand NAND2_4806 ( P3_U6615 , P3_U2396 , P3_ADD_360_1242_U14 );
nand NAND2_4807 ( P3_U6616 , P3_U2394 , P3_SUB_357_1258_U18 );
nand NAND2_4808 ( P3_U6617 , P3_U2389 , P3_REIP_REG_26_ );
nand NAND2_4809 ( P3_U6618 , P3_ADD_339_U75 , P3_U2388 );
nand NAND2_4810 ( P3_U6619 , P3_U2387 , P3_ADD_371_1212_U15 );
nand NAND2_4811 ( P3_U6620 , P3_PHYADDRPOINTER_REG_26_ , P3_U6404 );
nand NAND2_4812 ( P3_U6621 , P3_ADD_318_U74 , P3_U2398 );
nand NAND2_4813 ( P3_U6622 , P3_ADD_315_U71 , P3_U2397 );
nand NAND2_4814 ( P3_U6623 , P3_U2396 , P3_ADD_360_1242_U78 );
nand NAND2_4815 ( P3_U6624 , P3_U2394 , P3_SUB_357_1258_U80 );
nand NAND2_4816 ( P3_U6625 , P3_U2389 , P3_REIP_REG_27_ );
nand NAND2_4817 ( P3_U6626 , P3_ADD_339_U74 , P3_U2388 );
nand NAND2_4818 ( P3_U6627 , P3_U2387 , P3_ADD_371_1212_U80 );
nand NAND2_4819 ( P3_U6628 , P3_PHYADDRPOINTER_REG_27_ , P3_U6404 );
nand NAND2_4820 ( P3_U6629 , P3_ADD_318_U73 , P3_U2398 );
nand NAND2_4821 ( P3_U6630 , P3_ADD_315_U70 , P3_U2397 );
nand NAND2_4822 ( P3_U6631 , P3_U2396 , P3_ADD_360_1242_U15 );
nand NAND2_4823 ( P3_U6632 , P3_U2394 , P3_SUB_357_1258_U19 );
nand NAND2_4824 ( P3_U6633 , P3_U2389 , P3_REIP_REG_28_ );
nand NAND2_4825 ( P3_U6634 , P3_ADD_339_U73 , P3_U2388 );
nand NAND2_4826 ( P3_U6635 , P3_U2387 , P3_ADD_371_1212_U16 );
nand NAND2_4827 ( P3_U6636 , P3_PHYADDRPOINTER_REG_28_ , P3_U6404 );
nand NAND2_4828 ( P3_U6637 , P3_ADD_318_U72 , P3_U2398 );
nand NAND2_4829 ( P3_U6638 , P3_ADD_315_U69 , P3_U2397 );
nand NAND2_4830 ( P3_U6639 , P3_U2396 , P3_ADD_360_1242_U16 );
nand NAND2_4831 ( P3_U6640 , P3_U2394 , P3_SUB_357_1258_U79 );
nand NAND2_4832 ( P3_U6641 , P3_U2389 , P3_REIP_REG_29_ );
nand NAND2_4833 ( P3_U6642 , P3_ADD_339_U72 , P3_U2388 );
nand NAND2_4834 ( P3_U6643 , P3_U2387 , P3_ADD_371_1212_U17 );
nand NAND2_4835 ( P3_U6644 , P3_PHYADDRPOINTER_REG_29_ , P3_U6404 );
nand NAND2_4836 ( P3_U6645 , P3_ADD_318_U70 , P3_U2398 );
nand NAND2_4837 ( P3_U6646 , P3_ADD_315_U68 , P3_U2397 );
nand NAND2_4838 ( P3_U6647 , P3_U2396 , P3_ADD_360_1242_U77 );
nand NAND2_4839 ( P3_U6648 , P3_U2394 , P3_SUB_357_1258_U77 );
nand NAND2_4840 ( P3_U6649 , P3_U2389 , P3_REIP_REG_30_ );
nand NAND2_4841 ( P3_U6650 , P3_ADD_339_U70 , P3_U2388 );
nand NAND2_4842 ( P3_U6651 , P3_U2387 , P3_ADD_371_1212_U79 );
nand NAND2_4843 ( P3_U6652 , P3_PHYADDRPOINTER_REG_30_ , P3_U6404 );
nand NAND2_4844 ( P3_U6653 , P3_ADD_318_U69 , P3_U2398 );
nand NAND2_4845 ( P3_U6654 , P3_ADD_315_U67 , P3_U2397 );
nand NAND2_4846 ( P3_U6655 , P3_U2396 , P3_ADD_360_1242_U90 );
nand NAND2_4847 ( P3_U6656 , P3_U2394 , P3_SUB_357_1258_U20 );
nand NAND2_4848 ( P3_U6657 , P3_U2389 , P3_REIP_REG_31_ );
nand NAND2_4849 ( P3_U6658 , P3_ADD_339_U69 , P3_U2388 );
nand NAND2_4850 ( P3_U6659 , P3_U2387 , P3_ADD_371_1212_U92 );
nand NAND2_4851 ( P3_U6660 , P3_PHYADDRPOINTER_REG_31_ , P3_U6404 );
nand NAND3_4852 ( P3_U6661 , P3_U4304 , P3_U2630 , P3_GTE_412_U6 );
nand NAND2_4853 ( P3_U6662 , P3_GTE_450_U6 , P3_U4303 );
nand NAND2_4854 ( P3_U6663 , P3_U6662 , P3_U6661 );
nand NAND2_4855 ( P3_U6664 , P3_EAX_REG_15_ , P3_U2407 );
nand NAND2_4856 ( P3_U6665 , BUF2_REG_15_ , P3_U2406 );
nand NAND2_4857 ( P3_U6666 , P3_LWORD_REG_15_ , P3_U3250 );
nand NAND2_4858 ( P3_U6667 , P3_EAX_REG_14_ , P3_U2407 );
nand NAND2_4859 ( P3_U6668 , BUF2_REG_14_ , P3_U2406 );
nand NAND2_4860 ( P3_U6669 , P3_LWORD_REG_14_ , P3_U3250 );
nand NAND2_4861 ( P3_U6670 , P3_EAX_REG_13_ , P3_U2407 );
nand NAND2_4862 ( P3_U6671 , BUF2_REG_13_ , P3_U2406 );
nand NAND2_4863 ( P3_U6672 , P3_LWORD_REG_13_ , P3_U3250 );
nand NAND2_4864 ( P3_U6673 , P3_EAX_REG_12_ , P3_U2407 );
nand NAND2_4865 ( P3_U6674 , BUF2_REG_12_ , P3_U2406 );
nand NAND2_4866 ( P3_U6675 , P3_LWORD_REG_12_ , P3_U3250 );
nand NAND2_4867 ( P3_U6676 , P3_EAX_REG_11_ , P3_U2407 );
nand NAND2_4868 ( P3_U6677 , BUF2_REG_11_ , P3_U2406 );
nand NAND2_4869 ( P3_U6678 , P3_LWORD_REG_11_ , P3_U3250 );
nand NAND2_4870 ( P3_U6679 , P3_EAX_REG_10_ , P3_U2407 );
nand NAND2_4871 ( P3_U6680 , BUF2_REG_10_ , P3_U2406 );
nand NAND2_4872 ( P3_U6681 , P3_LWORD_REG_10_ , P3_U3250 );
nand NAND2_4873 ( P3_U6682 , P3_EAX_REG_9_ , P3_U2407 );
nand NAND2_4874 ( P3_U6683 , BUF2_REG_9_ , P3_U2406 );
nand NAND2_4875 ( P3_U6684 , P3_LWORD_REG_9_ , P3_U3250 );
nand NAND2_4876 ( P3_U6685 , P3_EAX_REG_8_ , P3_U2407 );
nand NAND2_4877 ( P3_U6686 , BUF2_REG_8_ , P3_U2406 );
nand NAND2_4878 ( P3_U6687 , P3_LWORD_REG_8_ , P3_U3250 );
nand NAND2_4879 ( P3_U6688 , P3_EAX_REG_7_ , P3_U2407 );
nand NAND2_4880 ( P3_U6689 , P3_U2406 , BUF2_REG_7_ );
nand NAND2_4881 ( P3_U6690 , P3_LWORD_REG_7_ , P3_U3250 );
nand NAND2_4882 ( P3_U6691 , P3_EAX_REG_6_ , P3_U2407 );
nand NAND2_4883 ( P3_U6692 , P3_U2406 , BUF2_REG_6_ );
nand NAND2_4884 ( P3_U6693 , P3_LWORD_REG_6_ , P3_U3250 );
nand NAND2_4885 ( P3_U6694 , P3_EAX_REG_5_ , P3_U2407 );
nand NAND2_4886 ( P3_U6695 , P3_U2406 , BUF2_REG_5_ );
nand NAND2_4887 ( P3_U6696 , P3_LWORD_REG_5_ , P3_U3250 );
nand NAND2_4888 ( P3_U6697 , P3_EAX_REG_4_ , P3_U2407 );
nand NAND2_4889 ( P3_U6698 , P3_U2406 , BUF2_REG_4_ );
nand NAND2_4890 ( P3_U6699 , P3_LWORD_REG_4_ , P3_U3250 );
nand NAND2_4891 ( P3_U6700 , P3_EAX_REG_3_ , P3_U2407 );
nand NAND2_4892 ( P3_U6701 , P3_U2406 , BUF2_REG_3_ );
nand NAND2_4893 ( P3_U6702 , P3_LWORD_REG_3_ , P3_U3250 );
nand NAND2_4894 ( P3_U6703 , P3_EAX_REG_2_ , P3_U2407 );
nand NAND2_4895 ( P3_U6704 , P3_U2406 , BUF2_REG_2_ );
nand NAND2_4896 ( P3_U6705 , P3_LWORD_REG_2_ , P3_U3250 );
nand NAND2_4897 ( P3_U6706 , P3_EAX_REG_1_ , P3_U2407 );
nand NAND2_4898 ( P3_U6707 , P3_U2406 , BUF2_REG_1_ );
nand NAND2_4899 ( P3_U6708 , P3_LWORD_REG_1_ , P3_U3250 );
nand NAND2_4900 ( P3_U6709 , P3_EAX_REG_0_ , P3_U2407 );
nand NAND2_4901 ( P3_U6710 , P3_U2406 , BUF2_REG_0_ );
nand NAND2_4902 ( P3_U6711 , P3_LWORD_REG_0_ , P3_U3250 );
nand NAND2_4903 ( P3_U6712 , P3_EAX_REG_30_ , P3_U2407 );
nand NAND2_4904 ( P3_U6713 , BUF2_REG_14_ , P3_U2406 );
nand NAND2_4905 ( P3_U6714 , P3_UWORD_REG_14_ , P3_U3250 );
nand NAND2_4906 ( P3_U6715 , P3_EAX_REG_29_ , P3_U2407 );
nand NAND2_4907 ( P3_U6716 , BUF2_REG_13_ , P3_U2406 );
nand NAND2_4908 ( P3_U6717 , P3_UWORD_REG_13_ , P3_U3250 );
nand NAND2_4909 ( P3_U6718 , P3_EAX_REG_28_ , P3_U2407 );
nand NAND2_4910 ( P3_U6719 , BUF2_REG_12_ , P3_U2406 );
nand NAND2_4911 ( P3_U6720 , P3_UWORD_REG_12_ , P3_U3250 );
nand NAND2_4912 ( P3_U6721 , P3_EAX_REG_27_ , P3_U2407 );
nand NAND2_4913 ( P3_U6722 , BUF2_REG_11_ , P3_U2406 );
nand NAND2_4914 ( P3_U6723 , P3_UWORD_REG_11_ , P3_U3250 );
nand NAND2_4915 ( P3_U6724 , P3_EAX_REG_26_ , P3_U2407 );
nand NAND2_4916 ( P3_U6725 , BUF2_REG_10_ , P3_U2406 );
nand NAND2_4917 ( P3_U6726 , P3_UWORD_REG_10_ , P3_U3250 );
nand NAND2_4918 ( P3_U6727 , P3_EAX_REG_25_ , P3_U2407 );
nand NAND2_4919 ( P3_U6728 , BUF2_REG_9_ , P3_U2406 );
nand NAND2_4920 ( P3_U6729 , P3_UWORD_REG_9_ , P3_U3250 );
nand NAND2_4921 ( P3_U6730 , P3_EAX_REG_24_ , P3_U2407 );
nand NAND2_4922 ( P3_U6731 , BUF2_REG_8_ , P3_U2406 );
nand NAND2_4923 ( P3_U6732 , P3_UWORD_REG_8_ , P3_U3250 );
nand NAND2_4924 ( P3_U6733 , P3_EAX_REG_23_ , P3_U2407 );
nand NAND2_4925 ( P3_U6734 , P3_U2406 , BUF2_REG_7_ );
nand NAND2_4926 ( P3_U6735 , P3_UWORD_REG_7_ , P3_U3250 );
nand NAND2_4927 ( P3_U6736 , P3_EAX_REG_22_ , P3_U2407 );
nand NAND2_4928 ( P3_U6737 , P3_U2406 , BUF2_REG_6_ );
nand NAND2_4929 ( P3_U6738 , P3_UWORD_REG_6_ , P3_U3250 );
nand NAND2_4930 ( P3_U6739 , P3_EAX_REG_21_ , P3_U2407 );
nand NAND2_4931 ( P3_U6740 , P3_U2406 , BUF2_REG_5_ );
nand NAND2_4932 ( P3_U6741 , P3_UWORD_REG_5_ , P3_U3250 );
nand NAND2_4933 ( P3_U6742 , P3_EAX_REG_20_ , P3_U2407 );
nand NAND2_4934 ( P3_U6743 , P3_U2406 , BUF2_REG_4_ );
nand NAND2_4935 ( P3_U6744 , P3_UWORD_REG_4_ , P3_U3250 );
nand NAND2_4936 ( P3_U6745 , P3_EAX_REG_19_ , P3_U2407 );
nand NAND2_4937 ( P3_U6746 , P3_U2406 , BUF2_REG_3_ );
nand NAND2_4938 ( P3_U6747 , P3_UWORD_REG_3_ , P3_U3250 );
nand NAND2_4939 ( P3_U6748 , P3_EAX_REG_18_ , P3_U2407 );
nand NAND2_4940 ( P3_U6749 , P3_U2406 , BUF2_REG_2_ );
nand NAND2_4941 ( P3_U6750 , P3_UWORD_REG_2_ , P3_U3250 );
nand NAND2_4942 ( P3_U6751 , P3_EAX_REG_17_ , P3_U2407 );
nand NAND2_4943 ( P3_U6752 , P3_U2406 , BUF2_REG_1_ );
nand NAND2_4944 ( P3_U6753 , P3_UWORD_REG_1_ , P3_U3250 );
nand NAND2_4945 ( P3_U6754 , P3_EAX_REG_16_ , P3_U2407 );
nand NAND2_4946 ( P3_U6755 , P3_U2406 , BUF2_REG_0_ );
nand NAND2_4947 ( P3_U6756 , P3_UWORD_REG_0_ , P3_U3250 );
nand NAND2_4948 ( P3_U6757 , P3_U3986 , P3_U3255 );
nand NAND2_4949 ( P3_U6758 , P3_U2453 , P3_U3121 );
not NOT1_4950 ( P3_U6759 , P3_U3251 );
nand NAND2_4951 ( P3_U6760 , P3_U2410 , P3_LWORD_REG_0_ );
nand NAND2_4952 ( P3_U6761 , P3_U2409 , P3_EAX_REG_0_ );
nand NAND2_4953 ( P3_U6762 , P3_DATAO_REG_0_ , P3_U6759 );
nand NAND2_4954 ( P3_U6763 , P3_U2410 , P3_LWORD_REG_1_ );
nand NAND2_4955 ( P3_U6764 , P3_U2409 , P3_EAX_REG_1_ );
nand NAND2_4956 ( P3_U6765 , P3_DATAO_REG_1_ , P3_U6759 );
nand NAND2_4957 ( P3_U6766 , P3_U2410 , P3_LWORD_REG_2_ );
nand NAND2_4958 ( P3_U6767 , P3_U2409 , P3_EAX_REG_2_ );
nand NAND2_4959 ( P3_U6768 , P3_DATAO_REG_2_ , P3_U6759 );
nand NAND2_4960 ( P3_U6769 , P3_U2410 , P3_LWORD_REG_3_ );
nand NAND2_4961 ( P3_U6770 , P3_U2409 , P3_EAX_REG_3_ );
nand NAND2_4962 ( P3_U6771 , P3_DATAO_REG_3_ , P3_U6759 );
nand NAND2_4963 ( P3_U6772 , P3_U2410 , P3_LWORD_REG_4_ );
nand NAND2_4964 ( P3_U6773 , P3_U2409 , P3_EAX_REG_4_ );
nand NAND2_4965 ( P3_U6774 , P3_DATAO_REG_4_ , P3_U6759 );
nand NAND2_4966 ( P3_U6775 , P3_U2410 , P3_LWORD_REG_5_ );
nand NAND2_4967 ( P3_U6776 , P3_U2409 , P3_EAX_REG_5_ );
nand NAND2_4968 ( P3_U6777 , P3_DATAO_REG_5_ , P3_U6759 );
nand NAND2_4969 ( P3_U6778 , P3_U2410 , P3_LWORD_REG_6_ );
nand NAND2_4970 ( P3_U6779 , P3_U2409 , P3_EAX_REG_6_ );
nand NAND2_4971 ( P3_U6780 , P3_DATAO_REG_6_ , P3_U6759 );
nand NAND2_4972 ( P3_U6781 , P3_U2410 , P3_LWORD_REG_7_ );
nand NAND2_4973 ( P3_U6782 , P3_U2409 , P3_EAX_REG_7_ );
nand NAND2_4974 ( P3_U6783 , P3_DATAO_REG_7_ , P3_U6759 );
nand NAND2_4975 ( P3_U6784 , P3_U2410 , P3_LWORD_REG_8_ );
nand NAND2_4976 ( P3_U6785 , P3_U2409 , P3_EAX_REG_8_ );
nand NAND2_4977 ( P3_U6786 , P3_DATAO_REG_8_ , P3_U6759 );
nand NAND2_4978 ( P3_U6787 , P3_U2410 , P3_LWORD_REG_9_ );
nand NAND2_4979 ( P3_U6788 , P3_U2409 , P3_EAX_REG_9_ );
nand NAND2_4980 ( P3_U6789 , P3_DATAO_REG_9_ , P3_U6759 );
nand NAND2_4981 ( P3_U6790 , P3_U2410 , P3_LWORD_REG_10_ );
nand NAND2_4982 ( P3_U6791 , P3_U2409 , P3_EAX_REG_10_ );
nand NAND2_4983 ( P3_U6792 , P3_DATAO_REG_10_ , P3_U6759 );
nand NAND2_4984 ( P3_U6793 , P3_U2410 , P3_LWORD_REG_11_ );
nand NAND2_4985 ( P3_U6794 , P3_U2409 , P3_EAX_REG_11_ );
nand NAND2_4986 ( P3_U6795 , P3_DATAO_REG_11_ , P3_U6759 );
nand NAND2_4987 ( P3_U6796 , P3_U2410 , P3_LWORD_REG_12_ );
nand NAND2_4988 ( P3_U6797 , P3_U2409 , P3_EAX_REG_12_ );
nand NAND2_4989 ( P3_U6798 , P3_DATAO_REG_12_ , P3_U6759 );
nand NAND2_4990 ( P3_U6799 , P3_U2410 , P3_LWORD_REG_13_ );
nand NAND2_4991 ( P3_U6800 , P3_U2409 , P3_EAX_REG_13_ );
nand NAND2_4992 ( P3_U6801 , P3_DATAO_REG_13_ , P3_U6759 );
nand NAND2_4993 ( P3_U6802 , P3_U2410 , P3_LWORD_REG_14_ );
nand NAND2_4994 ( P3_U6803 , P3_U2409 , P3_EAX_REG_14_ );
nand NAND2_4995 ( P3_U6804 , P3_DATAO_REG_14_ , P3_U6759 );
nand NAND2_4996 ( P3_U6805 , P3_U2410 , P3_LWORD_REG_15_ );
nand NAND2_4997 ( P3_U6806 , P3_U2409 , P3_EAX_REG_15_ );
nand NAND2_4998 ( P3_U6807 , P3_DATAO_REG_15_ , P3_U6759 );
nand NAND2_4999 ( P3_U6808 , P3_U2447 , P3_EAX_REG_16_ );
nand NAND2_5000 ( P3_U6809 , P3_U2410 , P3_UWORD_REG_0_ );
nand NAND2_5001 ( P3_U6810 , P3_DATAO_REG_16_ , P3_U6759 );
nand NAND2_5002 ( P3_U6811 , P3_U2447 , P3_EAX_REG_17_ );
nand NAND2_5003 ( P3_U6812 , P3_U2410 , P3_UWORD_REG_1_ );
nand NAND2_5004 ( P3_U6813 , P3_DATAO_REG_17_ , P3_U6759 );
nand NAND2_5005 ( P3_U6814 , P3_U2447 , P3_EAX_REG_18_ );
nand NAND2_5006 ( P3_U6815 , P3_U2410 , P3_UWORD_REG_2_ );
nand NAND2_5007 ( P3_U6816 , P3_DATAO_REG_18_ , P3_U6759 );
nand NAND2_5008 ( P3_U6817 , P3_U2447 , P3_EAX_REG_19_ );
nand NAND2_5009 ( P3_U6818 , P3_U2410 , P3_UWORD_REG_3_ );
nand NAND2_5010 ( P3_U6819 , P3_DATAO_REG_19_ , P3_U6759 );
nand NAND2_5011 ( P3_U6820 , P3_U2447 , P3_EAX_REG_20_ );
nand NAND2_5012 ( P3_U6821 , P3_U2410 , P3_UWORD_REG_4_ );
nand NAND2_5013 ( P3_U6822 , P3_DATAO_REG_20_ , P3_U6759 );
nand NAND2_5014 ( P3_U6823 , P3_U2447 , P3_EAX_REG_21_ );
nand NAND2_5015 ( P3_U6824 , P3_U2410 , P3_UWORD_REG_5_ );
nand NAND2_5016 ( P3_U6825 , P3_DATAO_REG_21_ , P3_U6759 );
nand NAND2_5017 ( P3_U6826 , P3_U2447 , P3_EAX_REG_22_ );
nand NAND2_5018 ( P3_U6827 , P3_U2410 , P3_UWORD_REG_6_ );
nand NAND2_5019 ( P3_U6828 , P3_DATAO_REG_22_ , P3_U6759 );
nand NAND2_5020 ( P3_U6829 , P3_U2447 , P3_EAX_REG_23_ );
nand NAND2_5021 ( P3_U6830 , P3_U2410 , P3_UWORD_REG_7_ );
nand NAND2_5022 ( P3_U6831 , P3_DATAO_REG_23_ , P3_U6759 );
nand NAND2_5023 ( P3_U6832 , P3_U2447 , P3_EAX_REG_24_ );
nand NAND2_5024 ( P3_U6833 , P3_U2410 , P3_UWORD_REG_8_ );
nand NAND2_5025 ( P3_U6834 , P3_DATAO_REG_24_ , P3_U6759 );
nand NAND2_5026 ( P3_U6835 , P3_U2447 , P3_EAX_REG_25_ );
nand NAND2_5027 ( P3_U6836 , P3_U2410 , P3_UWORD_REG_9_ );
nand NAND2_5028 ( P3_U6837 , P3_DATAO_REG_25_ , P3_U6759 );
nand NAND2_5029 ( P3_U6838 , P3_U2447 , P3_EAX_REG_26_ );
nand NAND2_5030 ( P3_U6839 , P3_U2410 , P3_UWORD_REG_10_ );
nand NAND2_5031 ( P3_U6840 , P3_DATAO_REG_26_ , P3_U6759 );
nand NAND2_5032 ( P3_U6841 , P3_U2447 , P3_EAX_REG_27_ );
nand NAND2_5033 ( P3_U6842 , P3_U2410 , P3_UWORD_REG_11_ );
nand NAND2_5034 ( P3_U6843 , P3_DATAO_REG_27_ , P3_U6759 );
nand NAND2_5035 ( P3_U6844 , P3_U2447 , P3_EAX_REG_28_ );
nand NAND2_5036 ( P3_U6845 , P3_U2410 , P3_UWORD_REG_12_ );
nand NAND2_5037 ( P3_U6846 , P3_DATAO_REG_28_ , P3_U6759 );
nand NAND2_5038 ( P3_U6847 , P3_U2447 , P3_EAX_REG_29_ );
nand NAND2_5039 ( P3_U6848 , P3_U2410 , P3_UWORD_REG_13_ );
nand NAND2_5040 ( P3_U6849 , P3_DATAO_REG_29_ , P3_U6759 );
nand NAND2_5041 ( P3_U6850 , P3_U2447 , P3_EAX_REG_30_ );
nand NAND2_5042 ( P3_U6851 , P3_U2410 , P3_UWORD_REG_14_ );
nand NAND2_5043 ( P3_U6852 , P3_DATAO_REG_30_ , P3_U6759 );
nand NAND2_5044 ( P3_U6853 , P3_U2516 , P3_U3243 );
nand NAND2_5045 ( P3_U6854 , P3_U2446 , BUF2_REG_0_ );
nand NAND2_5046 ( P3_U6855 , P3_U2621 , P3_U2411 );
nand NAND2_5047 ( P3_U6856 , P3_ADD_546_U5 , P3_U2400 );
nand NAND2_5048 ( P3_U6857 , P3_EAX_REG_0_ , P3_U3252 );
nand NAND2_5049 ( P3_U6858 , P3_U2446 , BUF2_REG_1_ );
nand NAND2_5050 ( P3_U6859 , P3_U2622 , P3_U2411 );
nand NAND2_5051 ( P3_U6860 , P3_ADD_546_U71 , P3_U2400 );
nand NAND2_5052 ( P3_U6861 , P3_EAX_REG_1_ , P3_U3252 );
nand NAND2_5053 ( P3_U6862 , P3_U2446 , BUF2_REG_2_ );
nand NAND2_5054 ( P3_U6863 , P3_U2623 , P3_U2411 );
nand NAND2_5055 ( P3_U6864 , P3_ADD_546_U60 , P3_U2400 );
nand NAND2_5056 ( P3_U6865 , P3_EAX_REG_2_ , P3_U3252 );
nand NAND2_5057 ( P3_U6866 , P3_U2446 , BUF2_REG_3_ );
nand NAND2_5058 ( P3_U6867 , P3_U2624 , P3_U2411 );
nand NAND2_5059 ( P3_U6868 , P3_ADD_546_U57 , P3_U2400 );
nand NAND2_5060 ( P3_U6869 , P3_EAX_REG_3_ , P3_U3252 );
nand NAND2_5061 ( P3_U6870 , P3_U2446 , BUF2_REG_4_ );
nand NAND2_5062 ( P3_U6871 , P3_U2625 , P3_U2411 );
nand NAND2_5063 ( P3_U6872 , P3_ADD_546_U56 , P3_U2400 );
nand NAND2_5064 ( P3_U6873 , P3_EAX_REG_4_ , P3_U3252 );
nand NAND2_5065 ( P3_U6874 , P3_U2446 , BUF2_REG_5_ );
nand NAND2_5066 ( P3_U6875 , P3_U2626 , P3_U2411 );
nand NAND2_5067 ( P3_U6876 , P3_ADD_546_U55 , P3_U2400 );
nand NAND2_5068 ( P3_U6877 , P3_EAX_REG_5_ , P3_U3252 );
nand NAND2_5069 ( P3_U6878 , P3_U2446 , BUF2_REG_6_ );
nand NAND2_5070 ( P3_U6879 , P3_U2627 , P3_U2411 );
nand NAND2_5071 ( P3_U6880 , P3_ADD_546_U54 , P3_U2400 );
nand NAND2_5072 ( P3_U6881 , P3_EAX_REG_6_ , P3_U3252 );
nand NAND2_5073 ( P3_U6882 , P3_U2446 , BUF2_REG_7_ );
nand NAND2_5074 ( P3_U6883 , P3_U2628 , P3_U2411 );
nand NAND2_5075 ( P3_U6884 , P3_ADD_546_U53 , P3_U2400 );
nand NAND2_5076 ( P3_U6885 , P3_EAX_REG_7_ , P3_U3252 );
nand NAND2_5077 ( P3_U6886 , P3_U2446 , BUF2_REG_8_ );
nand NAND2_5078 ( P3_U6887 , P3_U2605 , P3_U2411 );
nand NAND2_5079 ( P3_U6888 , P3_ADD_546_U52 , P3_U2400 );
nand NAND2_5080 ( P3_U6889 , P3_EAX_REG_8_ , P3_U3252 );
nand NAND2_5081 ( P3_U6890 , P3_U2446 , BUF2_REG_9_ );
nand NAND2_5082 ( P3_U6891 , P3_U2606 , P3_U2411 );
nand NAND2_5083 ( P3_U6892 , P3_ADD_546_U51 , P3_U2400 );
nand NAND2_5084 ( P3_U6893 , P3_EAX_REG_9_ , P3_U3252 );
nand NAND2_5085 ( P3_U6894 , P3_U2446 , BUF2_REG_10_ );
nand NAND2_5086 ( P3_U6895 , P3_U2607 , P3_U2411 );
nand NAND2_5087 ( P3_U6896 , P3_ADD_546_U81 , P3_U2400 );
nand NAND2_5088 ( P3_U6897 , P3_EAX_REG_10_ , P3_U3252 );
nand NAND2_5089 ( P3_U6898 , P3_U2446 , BUF2_REG_11_ );
nand NAND2_5090 ( P3_U6899 , P3_U2608 , P3_U2411 );
nand NAND2_5091 ( P3_U6900 , P3_ADD_546_U80 , P3_U2400 );
nand NAND2_5092 ( P3_U6901 , P3_EAX_REG_11_ , P3_U3252 );
nand NAND2_5093 ( P3_U6902 , P3_U2446 , BUF2_REG_12_ );
nand NAND2_5094 ( P3_U6903 , P3_U2609 , P3_U2411 );
nand NAND2_5095 ( P3_U6904 , P3_ADD_546_U79 , P3_U2400 );
nand NAND2_5096 ( P3_U6905 , P3_EAX_REG_12_ , P3_U3252 );
nand NAND2_5097 ( P3_U6906 , P3_U2446 , BUF2_REG_13_ );
nand NAND2_5098 ( P3_U6907 , P3_U2610 , P3_U2411 );
nand NAND2_5099 ( P3_U6908 , P3_ADD_546_U78 , P3_U2400 );
nand NAND2_5100 ( P3_U6909 , P3_EAX_REG_13_ , P3_U3252 );
nand NAND2_5101 ( P3_U6910 , P3_U2446 , BUF2_REG_14_ );
nand NAND2_5102 ( P3_U6911 , P3_U2611 , P3_U2411 );
nand NAND2_5103 ( P3_U6912 , P3_ADD_546_U77 , P3_U2400 );
nand NAND2_5104 ( P3_U6913 , P3_EAX_REG_14_ , P3_U3252 );
nand NAND2_5105 ( P3_U6914 , P3_U2446 , BUF2_REG_15_ );
nand NAND2_5106 ( P3_U6915 , P3_U2612 , P3_U2411 );
nand NAND2_5107 ( P3_U6916 , P3_ADD_546_U76 , P3_U2400 );
nand NAND2_5108 ( P3_U6917 , P3_EAX_REG_15_ , P3_U3252 );
nand NAND2_5109 ( P3_U6918 , P3_U2448 , BUF2_REG_0_ );
nand NAND2_5110 ( P3_U6919 , P3_U2444 , BUF2_REG_16_ );
nand NAND2_5111 ( P3_U6920 , P3_U3062 , P3_U2411 );
nand NAND2_5112 ( P3_U6921 , P3_ADD_546_U75 , P3_U2400 );
nand NAND2_5113 ( P3_U6922 , P3_EAX_REG_16_ , P3_U3252 );
nand NAND2_5114 ( P3_U6923 , P3_U2448 , BUF2_REG_1_ );
nand NAND2_5115 ( P3_U6924 , P3_U2444 , BUF2_REG_17_ );
nand NAND2_5116 ( P3_U6925 , P3_U3063 , P3_U2411 );
nand NAND2_5117 ( P3_U6926 , P3_ADD_546_U74 , P3_U2400 );
nand NAND2_5118 ( P3_U6927 , P3_EAX_REG_17_ , P3_U3252 );
nand NAND2_5119 ( P3_U6928 , P3_U2448 , BUF2_REG_2_ );
nand NAND2_5120 ( P3_U6929 , P3_U2444 , BUF2_REG_18_ );
nand NAND2_5121 ( P3_U6930 , P3_U3064 , P3_U2411 );
nand NAND2_5122 ( P3_U6931 , P3_ADD_546_U73 , P3_U2400 );
nand NAND2_5123 ( P3_U6932 , P3_EAX_REG_18_ , P3_U3252 );
nand NAND2_5124 ( P3_U6933 , P3_U2448 , BUF2_REG_3_ );
nand NAND2_5125 ( P3_U6934 , P3_U2444 , BUF2_REG_19_ );
nand NAND2_5126 ( P3_U6935 , P3_U3065 , P3_U2411 );
nand NAND2_5127 ( P3_U6936 , P3_ADD_546_U72 , P3_U2400 );
nand NAND2_5128 ( P3_U6937 , P3_EAX_REG_19_ , P3_U3252 );
nand NAND2_5129 ( P3_U6938 , P3_U2448 , BUF2_REG_4_ );
nand NAND2_5130 ( P3_U6939 , P3_U2444 , BUF2_REG_20_ );
nand NAND2_5131 ( P3_U6940 , P3_U3066 , P3_U2411 );
nand NAND2_5132 ( P3_U6941 , P3_ADD_546_U70 , P3_U2400 );
nand NAND2_5133 ( P3_U6942 , P3_EAX_REG_20_ , P3_U3252 );
nand NAND2_5134 ( P3_U6943 , P3_U2448 , BUF2_REG_5_ );
nand NAND2_5135 ( P3_U6944 , P3_U2444 , BUF2_REG_21_ );
nand NAND2_5136 ( P3_U6945 , P3_U3067 , P3_U2411 );
nand NAND2_5137 ( P3_U6946 , P3_ADD_546_U69 , P3_U2400 );
nand NAND2_5138 ( P3_U6947 , P3_EAX_REG_21_ , P3_U3252 );
nand NAND2_5139 ( P3_U6948 , P3_U2448 , BUF2_REG_6_ );
nand NAND2_5140 ( P3_U6949 , P3_U2444 , BUF2_REG_22_ );
nand NAND2_5141 ( P3_U6950 , P3_U3068 , P3_U2411 );
nand NAND2_5142 ( P3_U6951 , P3_ADD_546_U68 , P3_U2400 );
nand NAND2_5143 ( P3_U6952 , P3_EAX_REG_22_ , P3_U3252 );
nand NAND2_5144 ( P3_U6953 , P3_U2448 , BUF2_REG_7_ );
nand NAND2_5145 ( P3_U6954 , P3_U2444 , BUF2_REG_23_ );
nand NAND2_5146 ( P3_U6955 , P3_ADD_391_1180_U25 , P3_U2411 );
nand NAND2_5147 ( P3_U6956 , P3_ADD_546_U67 , P3_U2400 );
nand NAND2_5148 ( P3_U6957 , P3_EAX_REG_23_ , P3_U3252 );
nand NAND2_5149 ( P3_U6958 , P3_U2448 , BUF2_REG_8_ );
nand NAND2_5150 ( P3_U6959 , P3_U2444 , BUF2_REG_24_ );
nand NAND2_5151 ( P3_U6960 , P3_ADD_391_1180_U24 , P3_U2411 );
nand NAND2_5152 ( P3_U6961 , P3_ADD_546_U66 , P3_U2400 );
nand NAND2_5153 ( P3_U6962 , P3_EAX_REG_24_ , P3_U3252 );
nand NAND2_5154 ( P3_U6963 , P3_U2448 , BUF2_REG_9_ );
nand NAND2_5155 ( P3_U6964 , P3_U2444 , BUF2_REG_25_ );
nand NAND2_5156 ( P3_U6965 , P3_ADD_391_1180_U23 , P3_U2411 );
nand NAND2_5157 ( P3_U6966 , P3_ADD_546_U65 , P3_U2400 );
nand NAND2_5158 ( P3_U6967 , P3_EAX_REG_25_ , P3_U3252 );
nand NAND2_5159 ( P3_U6968 , P3_U2448 , BUF2_REG_10_ );
nand NAND2_5160 ( P3_U6969 , P3_U2444 , BUF2_REG_26_ );
nand NAND2_5161 ( P3_U6970 , P3_ADD_391_1180_U22 , P3_U2411 );
nand NAND2_5162 ( P3_U6971 , P3_ADD_546_U64 , P3_U2400 );
nand NAND2_5163 ( P3_U6972 , P3_EAX_REG_26_ , P3_U3252 );
nand NAND2_5164 ( P3_U6973 , P3_U2448 , BUF2_REG_11_ );
nand NAND2_5165 ( P3_U6974 , P3_U2444 , BUF2_REG_27_ );
nand NAND2_5166 ( P3_U6975 , P3_ADD_391_1180_U21 , P3_U2411 );
nand NAND2_5167 ( P3_U6976 , P3_ADD_546_U63 , P3_U2400 );
nand NAND2_5168 ( P3_U6977 , P3_EAX_REG_27_ , P3_U3252 );
nand NAND2_5169 ( P3_U6978 , P3_U2448 , BUF2_REG_12_ );
nand NAND2_5170 ( P3_U6979 , P3_U2444 , BUF2_REG_28_ );
nand NAND2_5171 ( P3_U6980 , P3_ADD_391_1180_U20 , P3_U2411 );
nand NAND2_5172 ( P3_U6981 , P3_ADD_546_U62 , P3_U2400 );
nand NAND2_5173 ( P3_U6982 , P3_EAX_REG_28_ , P3_U3252 );
nand NAND2_5174 ( P3_U6983 , P3_U2448 , BUF2_REG_13_ );
nand NAND2_5175 ( P3_U6984 , P3_U2444 , BUF2_REG_29_ );
nand NAND2_5176 ( P3_U6985 , P3_ADD_391_1180_U19 , P3_U2411 );
nand NAND2_5177 ( P3_U6986 , P3_ADD_546_U61 , P3_U2400 );
nand NAND2_5178 ( P3_U6987 , P3_EAX_REG_29_ , P3_U3252 );
nand NAND2_5179 ( P3_U6988 , P3_U2448 , BUF2_REG_14_ );
nand NAND2_5180 ( P3_U6989 , P3_U2444 , BUF2_REG_30_ );
nand NAND2_5181 ( P3_U6990 , P3_ADD_391_1180_U18 , P3_U2411 );
nand NAND2_5182 ( P3_U6991 , P3_ADD_546_U59 , P3_U2400 );
nand NAND2_5183 ( P3_U6992 , P3_EAX_REG_30_ , P3_U3252 );
nand NAND2_5184 ( P3_U6993 , P3_U2444 , BUF2_REG_31_ );
nand NAND2_5185 ( P3_U6994 , P3_ADD_546_U58 , P3_U2400 );
nand NAND2_5186 ( P3_U6995 , P3_EAX_REG_31_ , P3_U3252 );
nand NAND2_5187 ( P3_U6996 , P3_GTE_401_U6 , P3_U4305 );
nand NAND2_5188 ( P3_U6997 , P3_U3242 , P3_U6996 );
nand NAND2_5189 ( P3_U6998 , P3_INSTQUEUE_REG_0__0_ , P3_U2408 );
nand NAND2_5190 ( P3_U6999 , P3_ADD_552_U5 , P3_U2399 );
nand NAND2_5191 ( P3_U7000 , P3_EBX_REG_0_ , P3_U3253 );
nand NAND2_5192 ( P3_U7001 , P3_INSTQUEUE_REG_0__1_ , P3_U2408 );
nand NAND2_5193 ( P3_U7002 , P3_ADD_552_U71 , P3_U2399 );
nand NAND2_5194 ( P3_U7003 , P3_EBX_REG_1_ , P3_U3253 );
nand NAND2_5195 ( P3_U7004 , P3_INSTQUEUE_REG_0__2_ , P3_U2408 );
nand NAND2_5196 ( P3_U7005 , P3_ADD_552_U60 , P3_U2399 );
nand NAND2_5197 ( P3_U7006 , P3_EBX_REG_2_ , P3_U3253 );
nand NAND2_5198 ( P3_U7007 , P3_INSTQUEUE_REG_0__3_ , P3_U2408 );
nand NAND2_5199 ( P3_U7008 , P3_ADD_552_U57 , P3_U2399 );
nand NAND2_5200 ( P3_U7009 , P3_EBX_REG_3_ , P3_U3253 );
nand NAND2_5201 ( P3_U7010 , P3_INSTQUEUE_REG_0__4_ , P3_U2408 );
nand NAND2_5202 ( P3_U7011 , P3_ADD_552_U56 , P3_U2399 );
nand NAND2_5203 ( P3_U7012 , P3_EBX_REG_4_ , P3_U3253 );
nand NAND2_5204 ( P3_U7013 , P3_INSTQUEUE_REG_0__5_ , P3_U2408 );
nand NAND2_5205 ( P3_U7014 , P3_ADD_552_U55 , P3_U2399 );
nand NAND2_5206 ( P3_U7015 , P3_EBX_REG_5_ , P3_U3253 );
nand NAND2_5207 ( P3_U7016 , P3_INSTQUEUE_REG_0__6_ , P3_U2408 );
nand NAND2_5208 ( P3_U7017 , P3_ADD_552_U54 , P3_U2399 );
nand NAND2_5209 ( P3_U7018 , P3_EBX_REG_6_ , P3_U3253 );
nand NAND2_5210 ( P3_U7019 , P3_INSTQUEUE_REG_0__7_ , P3_U2408 );
nand NAND2_5211 ( P3_U7020 , P3_ADD_552_U53 , P3_U2399 );
nand NAND2_5212 ( P3_U7021 , P3_EBX_REG_7_ , P3_U3253 );
nand NAND2_5213 ( P3_U7022 , P3_U2605 , P3_U2408 );
nand NAND2_5214 ( P3_U7023 , P3_ADD_552_U52 , P3_U2399 );
nand NAND2_5215 ( P3_U7024 , P3_EBX_REG_8_ , P3_U3253 );
nand NAND2_5216 ( P3_U7025 , P3_U2606 , P3_U2408 );
nand NAND2_5217 ( P3_U7026 , P3_ADD_552_U51 , P3_U2399 );
nand NAND2_5218 ( P3_U7027 , P3_EBX_REG_9_ , P3_U3253 );
nand NAND2_5219 ( P3_U7028 , P3_U2607 , P3_U2408 );
nand NAND2_5220 ( P3_U7029 , P3_ADD_552_U81 , P3_U2399 );
nand NAND2_5221 ( P3_U7030 , P3_EBX_REG_10_ , P3_U3253 );
nand NAND2_5222 ( P3_U7031 , P3_U2608 , P3_U2408 );
nand NAND2_5223 ( P3_U7032 , P3_ADD_552_U80 , P3_U2399 );
nand NAND2_5224 ( P3_U7033 , P3_EBX_REG_11_ , P3_U3253 );
nand NAND2_5225 ( P3_U7034 , P3_U2609 , P3_U2408 );
nand NAND2_5226 ( P3_U7035 , P3_ADD_552_U79 , P3_U2399 );
nand NAND2_5227 ( P3_U7036 , P3_EBX_REG_12_ , P3_U3253 );
nand NAND2_5228 ( P3_U7037 , P3_U2610 , P3_U2408 );
nand NAND2_5229 ( P3_U7038 , P3_ADD_552_U78 , P3_U2399 );
nand NAND2_5230 ( P3_U7039 , P3_EBX_REG_13_ , P3_U3253 );
nand NAND2_5231 ( P3_U7040 , P3_U2611 , P3_U2408 );
nand NAND2_5232 ( P3_U7041 , P3_ADD_552_U77 , P3_U2399 );
nand NAND2_5233 ( P3_U7042 , P3_EBX_REG_14_ , P3_U3253 );
nand NAND2_5234 ( P3_U7043 , P3_U2612 , P3_U2408 );
nand NAND2_5235 ( P3_U7044 , P3_ADD_552_U76 , P3_U2399 );
nand NAND2_5236 ( P3_U7045 , P3_EBX_REG_15_ , P3_U3253 );
nand NAND2_5237 ( P3_U7046 , P3_U3062 , P3_U2408 );
nand NAND2_5238 ( P3_U7047 , P3_ADD_552_U75 , P3_U2399 );
nand NAND2_5239 ( P3_U7048 , P3_EBX_REG_16_ , P3_U3253 );
nand NAND2_5240 ( P3_U7049 , P3_U3063 , P3_U2408 );
nand NAND2_5241 ( P3_U7050 , P3_ADD_552_U74 , P3_U2399 );
nand NAND2_5242 ( P3_U7051 , P3_EBX_REG_17_ , P3_U3253 );
nand NAND2_5243 ( P3_U7052 , P3_U3064 , P3_U2408 );
nand NAND2_5244 ( P3_U7053 , P3_ADD_552_U73 , P3_U2399 );
nand NAND2_5245 ( P3_U7054 , P3_EBX_REG_18_ , P3_U3253 );
nand NAND2_5246 ( P3_U7055 , P3_U3065 , P3_U2408 );
nand NAND2_5247 ( P3_U7056 , P3_ADD_552_U72 , P3_U2399 );
nand NAND2_5248 ( P3_U7057 , P3_EBX_REG_19_ , P3_U3253 );
nand NAND2_5249 ( P3_U7058 , P3_U3066 , P3_U2408 );
nand NAND2_5250 ( P3_U7059 , P3_ADD_552_U70 , P3_U2399 );
nand NAND2_5251 ( P3_U7060 , P3_EBX_REG_20_ , P3_U3253 );
nand NAND2_5252 ( P3_U7061 , P3_U3067 , P3_U2408 );
nand NAND2_5253 ( P3_U7062 , P3_ADD_552_U69 , P3_U2399 );
nand NAND2_5254 ( P3_U7063 , P3_EBX_REG_21_ , P3_U3253 );
nand NAND2_5255 ( P3_U7064 , P3_U3068 , P3_U2408 );
nand NAND2_5256 ( P3_U7065 , P3_ADD_552_U68 , P3_U2399 );
nand NAND2_5257 ( P3_U7066 , P3_EBX_REG_22_ , P3_U3253 );
nand NAND2_5258 ( P3_U7067 , P3_ADD_402_1132_U25 , P3_U2408 );
nand NAND2_5259 ( P3_U7068 , P3_ADD_552_U67 , P3_U2399 );
nand NAND2_5260 ( P3_U7069 , P3_EBX_REG_23_ , P3_U3253 );
nand NAND2_5261 ( P3_U7070 , P3_ADD_402_1132_U24 , P3_U2408 );
nand NAND2_5262 ( P3_U7071 , P3_ADD_552_U66 , P3_U2399 );
nand NAND2_5263 ( P3_U7072 , P3_EBX_REG_24_ , P3_U3253 );
nand NAND2_5264 ( P3_U7073 , P3_ADD_402_1132_U23 , P3_U2408 );
nand NAND2_5265 ( P3_U7074 , P3_ADD_552_U65 , P3_U2399 );
nand NAND2_5266 ( P3_U7075 , P3_EBX_REG_25_ , P3_U3253 );
nand NAND2_5267 ( P3_U7076 , P3_ADD_402_1132_U22 , P3_U2408 );
nand NAND2_5268 ( P3_U7077 , P3_ADD_552_U64 , P3_U2399 );
nand NAND2_5269 ( P3_U7078 , P3_EBX_REG_26_ , P3_U3253 );
nand NAND2_5270 ( P3_U7079 , P3_ADD_402_1132_U21 , P3_U2408 );
nand NAND2_5271 ( P3_U7080 , P3_ADD_552_U63 , P3_U2399 );
nand NAND2_5272 ( P3_U7081 , P3_EBX_REG_27_ , P3_U3253 );
nand NAND2_5273 ( P3_U7082 , P3_ADD_402_1132_U20 , P3_U2408 );
nand NAND2_5274 ( P3_U7083 , P3_ADD_552_U62 , P3_U2399 );
nand NAND2_5275 ( P3_U7084 , P3_EBX_REG_28_ , P3_U3253 );
nand NAND2_5276 ( P3_U7085 , P3_ADD_402_1132_U19 , P3_U2408 );
nand NAND2_5277 ( P3_U7086 , P3_ADD_552_U61 , P3_U2399 );
nand NAND2_5278 ( P3_U7087 , P3_EBX_REG_29_ , P3_U3253 );
nand NAND2_5279 ( P3_U7088 , P3_ADD_402_1132_U18 , P3_U2408 );
nand NAND2_5280 ( P3_U7089 , P3_ADD_552_U59 , P3_U2399 );
nand NAND2_5281 ( P3_U7090 , P3_EBX_REG_30_ , P3_U3253 );
nand NAND2_5282 ( P3_U7091 , P3_ADD_552_U58 , P3_U2399 );
nand NAND2_5283 ( P3_U7092 , P3_EBX_REG_31_ , P3_U3253 );
nand NAND2_5284 ( P3_U7093 , P3_U5488 , P3_U5491 );
not NOT1_5285 ( P3_U7094 , P3_U3260 );
not NOT1_5286 ( P3_U7095 , P3_U3257 );
or OR2_5287 ( P3_U7096 , P3_STATEBS16_REG , U209 );
nand NAND2_5288 ( P3_U7097 , P3_EBX_REG_0_ , P3_U2602 );
nand NAND2_5289 ( P3_U7098 , P3_REIP_REG_0_ , P3_U2601 );
nand NAND2_5290 ( P3_U7099 , P3_EBX_REG_0_ , P3_U7910 );
nand NAND2_5291 ( P3_U7100 , P3_ADD_505_U5 , P3_U2455 );
nand NAND2_5292 ( P3_U7101 , P3_ADD_486_U5 , P3_U2454 );
nand NAND2_5293 ( P3_U7102 , P3_REIP_REG_0_ , P3_U2405 );
nand NAND2_5294 ( P3_U7103 , P3_U2403 , P3_PHYADDRPOINTER_REG_0_ );
nand NAND2_5295 ( P3_U7104 , P3_PHYADDRPOINTER_REG_0_ , P3_U4319 );
nand NAND2_5296 ( P3_U7105 , P3_U2401 , P3_PHYADDRPOINTER_REG_0_ );
nand NAND2_5297 ( P3_U7106 , P3_U7094 , P3_REIP_REG_0_ );
nand NAND2_5298 ( P3_U7107 , P3_SUB_414_U50 , P3_U2602 );
nand NAND2_5299 ( P3_U7108 , P3_ADD_467_U4 , P3_U2601 );
nand NAND2_5300 ( P3_U7109 , P3_EBX_REG_1_ , P3_U7910 );
nand NAND2_5301 ( P3_U7110 , P3_ADD_505_U17 , P3_U2455 );
nand NAND2_5302 ( P3_U7111 , P3_ADD_486_U17 , P3_U2454 );
nand NAND2_5303 ( P3_U7112 , P3_ADD_430_U4 , P3_U2405 );
nand NAND2_5304 ( P3_U7113 , P3_U2403 , P3_ADD_318_U4 );
nand NAND2_5305 ( P3_U7114 , P3_SUB_320_U50 , P3_U4319 );
nand NAND2_5306 ( P3_U7115 , P3_U2401 , P3_PHYADDRPOINTER_REG_1_ );
nand NAND2_5307 ( P3_U7116 , P3_U7094 , P3_REIP_REG_1_ );
nand NAND2_5308 ( P3_U7117 , P3_SUB_414_U17 , P3_U2602 );
nand NAND2_5309 ( P3_U7118 , P3_ADD_467_U71 , P3_U2601 );
nand NAND2_5310 ( P3_U7119 , P3_EBX_REG_2_ , P3_U7910 );
nand NAND2_5311 ( P3_U7120 , P3_ADD_505_U16 , P3_U2455 );
nand NAND2_5312 ( P3_U7121 , P3_ADD_486_U16 , P3_U2454 );
nand NAND2_5313 ( P3_U7122 , P3_ADD_430_U71 , P3_U2405 );
nand NAND2_5314 ( P3_U7123 , P3_U2403 , P3_ADD_318_U71 );
nand NAND2_5315 ( P3_U7124 , P3_SUB_320_U17 , P3_U4319 );
nand NAND2_5316 ( P3_U7125 , P3_U2401 , P3_PHYADDRPOINTER_REG_2_ );
nand NAND2_5317 ( P3_U7126 , P3_U7094 , P3_REIP_REG_2_ );
nand NAND2_5318 ( P3_U7127 , P3_SUB_414_U59 , P3_U2602 );
nand NAND2_5319 ( P3_U7128 , P3_ADD_467_U68 , P3_U2601 );
nand NAND2_5320 ( P3_U7129 , P3_EBX_REG_3_ , P3_U7910 );
nand NAND2_5321 ( P3_U7130 , P3_ADD_505_U15 , P3_U2455 );
nand NAND2_5322 ( P3_U7131 , P3_ADD_486_U15 , P3_U2454 );
nand NAND2_5323 ( P3_U7132 , P3_ADD_430_U68 , P3_U2405 );
nand NAND2_5324 ( P3_U7133 , P3_U2403 , P3_ADD_318_U68 );
nand NAND2_5325 ( P3_U7134 , P3_SUB_320_U59 , P3_U4319 );
nand NAND2_5326 ( P3_U7135 , P3_U2401 , P3_PHYADDRPOINTER_REG_3_ );
nand NAND2_5327 ( P3_U7136 , P3_U7094 , P3_REIP_REG_3_ );
nand NAND2_5328 ( P3_U7137 , P3_SUB_414_U18 , P3_U2602 );
nand NAND2_5329 ( P3_U7138 , P3_ADD_467_U67 , P3_U2601 );
nand NAND2_5330 ( P3_U7139 , P3_EBX_REG_4_ , P3_U7910 );
nand NAND2_5331 ( P3_U7140 , P3_ADD_505_U14 , P3_U2455 );
nand NAND2_5332 ( P3_U7141 , P3_ADD_486_U14 , P3_U2454 );
nand NAND2_5333 ( P3_U7142 , P3_ADD_430_U67 , P3_U2405 );
nand NAND2_5334 ( P3_U7143 , P3_U2403 , P3_ADD_318_U67 );
nand NAND2_5335 ( P3_U7144 , P3_SUB_320_U18 , P3_U4319 );
nand NAND2_5336 ( P3_U7145 , P3_U2401 , P3_PHYADDRPOINTER_REG_4_ );
nand NAND2_5337 ( P3_U7146 , P3_U7094 , P3_REIP_REG_4_ );
nand NAND2_5338 ( P3_U7147 , P3_SUB_414_U57 , P3_U2602 );
nand NAND2_5339 ( P3_U7148 , P3_ADD_467_U66 , P3_U2601 );
nand NAND2_5340 ( P3_U7149 , P3_EBX_REG_5_ , P3_U7910 );
nand NAND2_5341 ( P3_U7150 , P3_ADD_505_U6 , P3_U2455 );
nand NAND2_5342 ( P3_U7151 , P3_ADD_486_U6 , P3_U2454 );
nand NAND2_5343 ( P3_U7152 , P3_ADD_430_U66 , P3_U2405 );
nand NAND2_5344 ( P3_U7153 , P3_U2403 , P3_ADD_318_U66 );
nand NAND2_5345 ( P3_U7154 , P3_SUB_320_U57 , P3_U4319 );
nand NAND2_5346 ( P3_U7155 , P3_U2401 , P3_PHYADDRPOINTER_REG_5_ );
nand NAND2_5347 ( P3_U7156 , P3_U7094 , P3_REIP_REG_5_ );
nand NAND2_5348 ( P3_U7157 , P3_SUB_414_U19 , P3_U2602 );
nand NAND2_5349 ( P3_U7158 , P3_ADD_467_U65 , P3_U2601 );
nand NAND2_5350 ( P3_U7159 , P3_EBX_REG_6_ , P3_U7910 );
nand NAND2_5351 ( P3_U7160 , P3_ADD_430_U65 , P3_U2405 );
nand NAND2_5352 ( P3_U7161 , P3_U2403 , P3_ADD_318_U65 );
nand NAND2_5353 ( P3_U7162 , P3_SUB_320_U19 , P3_U4319 );
nand NAND2_5354 ( P3_U7163 , P3_U2401 , P3_PHYADDRPOINTER_REG_6_ );
nand NAND2_5355 ( P3_U7164 , P3_U7094 , P3_REIP_REG_6_ );
nand NAND2_5356 ( P3_U7165 , P3_SUB_414_U55 , P3_U2602 );
nand NAND2_5357 ( P3_U7166 , P3_ADD_467_U64 , P3_U2601 );
nand NAND2_5358 ( P3_U7167 , P3_EBX_REG_7_ , P3_U7910 );
nand NAND2_5359 ( P3_U7168 , P3_ADD_430_U64 , P3_U2405 );
nand NAND2_5360 ( P3_U7169 , P3_U2403 , P3_ADD_318_U64 );
nand NAND2_5361 ( P3_U7170 , P3_SUB_320_U55 , P3_U4319 );
nand NAND2_5362 ( P3_U7171 , P3_U2401 , P3_PHYADDRPOINTER_REG_7_ );
nand NAND2_5363 ( P3_U7172 , P3_U7094 , P3_REIP_REG_7_ );
nand NAND2_5364 ( P3_U7173 , P3_SUB_414_U20 , P3_U2602 );
nand NAND2_5365 ( P3_U7174 , P3_ADD_467_U63 , P3_U2601 );
nand NAND2_5366 ( P3_U7175 , P3_EBX_REG_8_ , P3_U7910 );
nand NAND2_5367 ( P3_U7176 , P3_ADD_430_U63 , P3_U2405 );
nand NAND2_5368 ( P3_U7177 , P3_U2403 , P3_ADD_318_U63 );
nand NAND2_5369 ( P3_U7178 , P3_SUB_320_U20 , P3_U4319 );
nand NAND2_5370 ( P3_U7179 , P3_U2401 , P3_PHYADDRPOINTER_REG_8_ );
nand NAND2_5371 ( P3_U7180 , P3_U7094 , P3_REIP_REG_8_ );
nand NAND2_5372 ( P3_U7181 , P3_SUB_414_U53 , P3_U2602 );
nand NAND2_5373 ( P3_U7182 , P3_ADD_467_U62 , P3_U2601 );
nand NAND2_5374 ( P3_U7183 , P3_EBX_REG_9_ , P3_U7910 );
nand NAND2_5375 ( P3_U7184 , P3_ADD_430_U62 , P3_U2405 );
nand NAND2_5376 ( P3_U7185 , P3_U2403 , P3_ADD_318_U62 );
nand NAND2_5377 ( P3_U7186 , P3_SUB_320_U53 , P3_U4319 );
nand NAND2_5378 ( P3_U7187 , P3_U2401 , P3_PHYADDRPOINTER_REG_9_ );
nand NAND2_5379 ( P3_U7188 , P3_U7094 , P3_REIP_REG_9_ );
nand NAND2_5380 ( P3_U7189 , P3_SUB_414_U6 , P3_U2602 );
nand NAND2_5381 ( P3_U7190 , P3_ADD_467_U91 , P3_U2601 );
nand NAND2_5382 ( P3_U7191 , P3_EBX_REG_10_ , P3_U7910 );
nand NAND2_5383 ( P3_U7192 , P3_ADD_430_U91 , P3_U2405 );
nand NAND2_5384 ( P3_U7193 , P3_U2403 , P3_ADD_318_U91 );
nand NAND2_5385 ( P3_U7194 , P3_SUB_320_U6 , P3_U4319 );
nand NAND2_5386 ( P3_U7195 , P3_U2401 , P3_PHYADDRPOINTER_REG_10_ );
nand NAND2_5387 ( P3_U7196 , P3_U7094 , P3_REIP_REG_10_ );
nand NAND2_5388 ( P3_U7197 , P3_SUB_414_U82 , P3_U2602 );
nand NAND2_5389 ( P3_U7198 , P3_ADD_467_U90 , P3_U2601 );
nand NAND2_5390 ( P3_U7199 , P3_EBX_REG_11_ , P3_U7910 );
nand NAND2_5391 ( P3_U7200 , P3_ADD_430_U90 , P3_U2405 );
nand NAND2_5392 ( P3_U7201 , P3_U2403 , P3_ADD_318_U90 );
nand NAND2_5393 ( P3_U7202 , P3_SUB_320_U82 , P3_U4319 );
nand NAND2_5394 ( P3_U7203 , P3_U2401 , P3_PHYADDRPOINTER_REG_11_ );
nand NAND2_5395 ( P3_U7204 , P3_U7094 , P3_REIP_REG_11_ );
nand NAND2_5396 ( P3_U7205 , P3_SUB_414_U7 , P3_U2602 );
nand NAND2_5397 ( P3_U7206 , P3_ADD_467_U89 , P3_U2601 );
nand NAND2_5398 ( P3_U7207 , P3_EBX_REG_12_ , P3_U7910 );
nand NAND2_5399 ( P3_U7208 , P3_ADD_430_U89 , P3_U2405 );
nand NAND2_5400 ( P3_U7209 , P3_U2403 , P3_ADD_318_U89 );
nand NAND2_5401 ( P3_U7210 , P3_SUB_320_U7 , P3_U4319 );
nand NAND2_5402 ( P3_U7211 , P3_U2401 , P3_PHYADDRPOINTER_REG_12_ );
nand NAND2_5403 ( P3_U7212 , P3_U7094 , P3_REIP_REG_12_ );
nand NAND2_5404 ( P3_U7213 , P3_SUB_414_U80 , P3_U2602 );
nand NAND2_5405 ( P3_U7214 , P3_ADD_467_U88 , P3_U2601 );
nand NAND2_5406 ( P3_U7215 , P3_EBX_REG_13_ , P3_U7910 );
nand NAND2_5407 ( P3_U7216 , P3_ADD_430_U88 , P3_U2405 );
nand NAND2_5408 ( P3_U7217 , P3_U2403 , P3_ADD_318_U88 );
nand NAND2_5409 ( P3_U7218 , P3_SUB_320_U80 , P3_U4319 );
nand NAND2_5410 ( P3_U7219 , P3_U2401 , P3_PHYADDRPOINTER_REG_13_ );
nand NAND2_5411 ( P3_U7220 , P3_U7094 , P3_REIP_REG_13_ );
nand NAND2_5412 ( P3_U7221 , P3_SUB_414_U8 , P3_U2602 );
nand NAND2_5413 ( P3_U7222 , P3_ADD_467_U87 , P3_U2601 );
nand NAND2_5414 ( P3_U7223 , P3_EBX_REG_14_ , P3_U7910 );
nand NAND2_5415 ( P3_U7224 , P3_ADD_430_U87 , P3_U2405 );
nand NAND2_5416 ( P3_U7225 , P3_U2403 , P3_ADD_318_U87 );
nand NAND2_5417 ( P3_U7226 , P3_SUB_320_U8 , P3_U4319 );
nand NAND2_5418 ( P3_U7227 , P3_U2401 , P3_PHYADDRPOINTER_REG_14_ );
nand NAND2_5419 ( P3_U7228 , P3_U7094 , P3_REIP_REG_14_ );
nand NAND2_5420 ( P3_U7229 , P3_SUB_414_U78 , P3_U2602 );
nand NAND2_5421 ( P3_U7230 , P3_ADD_467_U86 , P3_U2601 );
nand NAND2_5422 ( P3_U7231 , P3_EBX_REG_15_ , P3_U7910 );
nand NAND2_5423 ( P3_U7232 , P3_ADD_430_U86 , P3_U2405 );
nand NAND2_5424 ( P3_U7233 , P3_U2403 , P3_ADD_318_U86 );
nand NAND2_5425 ( P3_U7234 , P3_SUB_320_U78 , P3_U4319 );
nand NAND2_5426 ( P3_U7235 , P3_U2401 , P3_PHYADDRPOINTER_REG_15_ );
nand NAND2_5427 ( P3_U7236 , P3_U7094 , P3_REIP_REG_15_ );
nand NAND2_5428 ( P3_U7237 , P3_SUB_414_U9 , P3_U2602 );
nand NAND2_5429 ( P3_U7238 , P3_ADD_467_U85 , P3_U2601 );
nand NAND2_5430 ( P3_U7239 , P3_EBX_REG_16_ , P3_U7910 );
nand NAND2_5431 ( P3_U7240 , P3_ADD_430_U85 , P3_U2405 );
nand NAND2_5432 ( P3_U7241 , P3_U2403 , P3_ADD_318_U85 );
nand NAND2_5433 ( P3_U7242 , P3_SUB_320_U9 , P3_U4319 );
nand NAND2_5434 ( P3_U7243 , P3_U2401 , P3_PHYADDRPOINTER_REG_16_ );
nand NAND2_5435 ( P3_U7244 , P3_U7094 , P3_REIP_REG_16_ );
nand NAND2_5436 ( P3_U7245 , P3_SUB_414_U76 , P3_U2602 );
nand NAND2_5437 ( P3_U7246 , P3_ADD_467_U84 , P3_U2601 );
nand NAND2_5438 ( P3_U7247 , P3_EBX_REG_17_ , P3_U7910 );
nand NAND2_5439 ( P3_U7248 , P3_ADD_430_U84 , P3_U2405 );
nand NAND2_5440 ( P3_U7249 , P3_U2403 , P3_ADD_318_U84 );
nand NAND2_5441 ( P3_U7250 , P3_SUB_320_U76 , P3_U4319 );
nand NAND2_5442 ( P3_U7251 , P3_U2401 , P3_PHYADDRPOINTER_REG_17_ );
nand NAND2_5443 ( P3_U7252 , P3_U7094 , P3_REIP_REG_17_ );
nand NAND2_5444 ( P3_U7253 , P3_SUB_414_U10 , P3_U2602 );
nand NAND2_5445 ( P3_U7254 , P3_ADD_467_U83 , P3_U2601 );
nand NAND2_5446 ( P3_U7255 , P3_EBX_REG_18_ , P3_U7910 );
nand NAND2_5447 ( P3_U7256 , P3_ADD_430_U83 , P3_U2405 );
nand NAND2_5448 ( P3_U7257 , P3_U2403 , P3_ADD_318_U83 );
nand NAND2_5449 ( P3_U7258 , P3_SUB_320_U10 , P3_U4319 );
nand NAND2_5450 ( P3_U7259 , P3_U2401 , P3_PHYADDRPOINTER_REG_18_ );
nand NAND2_5451 ( P3_U7260 , P3_U7094 , P3_REIP_REG_18_ );
nand NAND2_5452 ( P3_U7261 , P3_SUB_414_U74 , P3_U2602 );
nand NAND2_5453 ( P3_U7262 , P3_ADD_467_U82 , P3_U2601 );
nand NAND2_5454 ( P3_U7263 , P3_EBX_REG_19_ , P3_U7910 );
nand NAND2_5455 ( P3_U7264 , P3_ADD_430_U82 , P3_U2405 );
nand NAND2_5456 ( P3_U7265 , P3_U2403 , P3_ADD_318_U82 );
nand NAND2_5457 ( P3_U7266 , P3_SUB_320_U74 , P3_U4319 );
nand NAND2_5458 ( P3_U7267 , P3_U2401 , P3_PHYADDRPOINTER_REG_19_ );
nand NAND2_5459 ( P3_U7268 , P3_U7094 , P3_REIP_REG_19_ );
nand NAND2_5460 ( P3_U7269 , P3_SUB_414_U11 , P3_U2602 );
nand NAND2_5461 ( P3_U7270 , P3_ADD_467_U81 , P3_U2601 );
nand NAND2_5462 ( P3_U7271 , P3_EBX_REG_20_ , P3_U7910 );
nand NAND2_5463 ( P3_U7272 , P3_ADD_430_U81 , P3_U2405 );
nand NAND2_5464 ( P3_U7273 , P3_U2403 , P3_ADD_318_U81 );
nand NAND2_5465 ( P3_U7274 , P3_SUB_320_U11 , P3_U4319 );
nand NAND2_5466 ( P3_U7275 , P3_U2401 , P3_PHYADDRPOINTER_REG_20_ );
nand NAND2_5467 ( P3_U7276 , P3_U7094 , P3_REIP_REG_20_ );
nand NAND2_5468 ( P3_U7277 , P3_SUB_414_U70 , P3_U2602 );
nand NAND2_5469 ( P3_U7278 , P3_ADD_467_U80 , P3_U2601 );
nand NAND2_5470 ( P3_U7279 , P3_EBX_REG_21_ , P3_U7910 );
nand NAND2_5471 ( P3_U7280 , P3_ADD_430_U80 , P3_U2405 );
nand NAND2_5472 ( P3_U7281 , P3_U2403 , P3_ADD_318_U80 );
nand NAND2_5473 ( P3_U7282 , P3_SUB_320_U70 , P3_U4319 );
nand NAND2_5474 ( P3_U7283 , P3_U2401 , P3_PHYADDRPOINTER_REG_21_ );
nand NAND2_5475 ( P3_U7284 , P3_U7094 , P3_REIP_REG_21_ );
nand NAND2_5476 ( P3_U7285 , P3_SUB_414_U12 , P3_U2602 );
nand NAND2_5477 ( P3_U7286 , P3_ADD_467_U79 , P3_U2601 );
nand NAND2_5478 ( P3_U7287 , P3_EBX_REG_22_ , P3_U7910 );
nand NAND2_5479 ( P3_U7288 , P3_ADD_430_U79 , P3_U2405 );
nand NAND2_5480 ( P3_U7289 , P3_U2403 , P3_ADD_318_U79 );
nand NAND2_5481 ( P3_U7290 , P3_SUB_320_U12 , P3_U4319 );
nand NAND2_5482 ( P3_U7291 , P3_U2401 , P3_PHYADDRPOINTER_REG_22_ );
nand NAND2_5483 ( P3_U7292 , P3_U7094 , P3_REIP_REG_22_ );
nand NAND2_5484 ( P3_U7293 , P3_SUB_414_U68 , P3_U2602 );
nand NAND2_5485 ( P3_U7294 , P3_ADD_467_U78 , P3_U2601 );
nand NAND2_5486 ( P3_U7295 , P3_EBX_REG_23_ , P3_U7910 );
nand NAND2_5487 ( P3_U7296 , P3_ADD_430_U78 , P3_U2405 );
nand NAND2_5488 ( P3_U7297 , P3_U2403 , P3_ADD_318_U78 );
nand NAND2_5489 ( P3_U7298 , P3_SUB_320_U68 , P3_U4319 );
nand NAND2_5490 ( P3_U7299 , P3_U2401 , P3_PHYADDRPOINTER_REG_23_ );
nand NAND2_5491 ( P3_U7300 , P3_U7094 , P3_REIP_REG_23_ );
nand NAND2_5492 ( P3_U7301 , P3_SUB_414_U13 , P3_U2602 );
nand NAND2_5493 ( P3_U7302 , P3_ADD_467_U77 , P3_U2601 );
nand NAND2_5494 ( P3_U7303 , P3_EBX_REG_24_ , P3_U7910 );
nand NAND2_5495 ( P3_U7304 , P3_ADD_430_U77 , P3_U2405 );
nand NAND2_5496 ( P3_U7305 , P3_U2403 , P3_ADD_318_U77 );
nand NAND2_5497 ( P3_U7306 , P3_SUB_320_U13 , P3_U4319 );
nand NAND2_5498 ( P3_U7307 , P3_U2401 , P3_PHYADDRPOINTER_REG_24_ );
nand NAND2_5499 ( P3_U7308 , P3_U7094 , P3_REIP_REG_24_ );
nand NAND2_5500 ( P3_U7309 , P3_SUB_414_U66 , P3_U2602 );
nand NAND2_5501 ( P3_U7310 , P3_ADD_467_U76 , P3_U2601 );
nand NAND2_5502 ( P3_U7311 , P3_EBX_REG_25_ , P3_U7910 );
nand NAND2_5503 ( P3_U7312 , P3_ADD_430_U76 , P3_U2405 );
nand NAND2_5504 ( P3_U7313 , P3_U2403 , P3_ADD_318_U76 );
nand NAND2_5505 ( P3_U7314 , P3_SUB_320_U66 , P3_U4319 );
nand NAND2_5506 ( P3_U7315 , P3_U2401 , P3_PHYADDRPOINTER_REG_25_ );
nand NAND2_5507 ( P3_U7316 , P3_U7094 , P3_REIP_REG_25_ );
nand NAND2_5508 ( P3_U7317 , P3_SUB_414_U14 , P3_U2602 );
nand NAND2_5509 ( P3_U7318 , P3_ADD_467_U75 , P3_U2601 );
nand NAND2_5510 ( P3_U7319 , P3_EBX_REG_26_ , P3_U7910 );
nand NAND2_5511 ( P3_U7320 , P3_ADD_430_U75 , P3_U2405 );
nand NAND2_5512 ( P3_U7321 , P3_U2403 , P3_ADD_318_U75 );
nand NAND2_5513 ( P3_U7322 , P3_SUB_320_U14 , P3_U4319 );
nand NAND2_5514 ( P3_U7323 , P3_U2401 , P3_PHYADDRPOINTER_REG_26_ );
nand NAND2_5515 ( P3_U7324 , P3_U7094 , P3_REIP_REG_26_ );
nand NAND2_5516 ( P3_U7325 , P3_SUB_414_U64 , P3_U2602 );
nand NAND2_5517 ( P3_U7326 , P3_ADD_467_U74 , P3_U2601 );
nand NAND2_5518 ( P3_U7327 , P3_EBX_REG_27_ , P3_U7910 );
nand NAND2_5519 ( P3_U7328 , P3_ADD_430_U74 , P3_U2405 );
nand NAND2_5520 ( P3_U7329 , P3_U2403 , P3_ADD_318_U74 );
nand NAND2_5521 ( P3_U7330 , P3_SUB_320_U64 , P3_U4319 );
nand NAND2_5522 ( P3_U7331 , P3_U2401 , P3_PHYADDRPOINTER_REG_27_ );
nand NAND2_5523 ( P3_U7332 , P3_U7094 , P3_REIP_REG_27_ );
nand NAND2_5524 ( P3_U7333 , P3_SUB_414_U15 , P3_U2602 );
nand NAND2_5525 ( P3_U7334 , P3_ADD_467_U73 , P3_U2601 );
nand NAND2_5526 ( P3_U7335 , P3_EBX_REG_28_ , P3_U7910 );
nand NAND2_5527 ( P3_U7336 , P3_ADD_430_U73 , P3_U2405 );
nand NAND2_5528 ( P3_U7337 , P3_U2403 , P3_ADD_318_U73 );
nand NAND2_5529 ( P3_U7338 , P3_SUB_320_U15 , P3_U4319 );
nand NAND2_5530 ( P3_U7339 , P3_U2401 , P3_PHYADDRPOINTER_REG_28_ );
nand NAND2_5531 ( P3_U7340 , P3_U7094 , P3_REIP_REG_28_ );
nand NAND2_5532 ( P3_U7341 , P3_SUB_414_U16 , P3_U2602 );
nand NAND2_5533 ( P3_U7342 , P3_ADD_467_U72 , P3_U2601 );
nand NAND2_5534 ( P3_U7343 , P3_EBX_REG_29_ , P3_U7910 );
nand NAND2_5535 ( P3_U7344 , P3_ADD_430_U72 , P3_U2405 );
nand NAND2_5536 ( P3_U7345 , P3_U2403 , P3_ADD_318_U72 );
nand NAND2_5537 ( P3_U7346 , P3_SUB_320_U16 , P3_U4319 );
nand NAND2_5538 ( P3_U7347 , P3_U2401 , P3_PHYADDRPOINTER_REG_29_ );
nand NAND2_5539 ( P3_U7348 , P3_U7094 , P3_REIP_REG_29_ );
nand NAND2_5540 ( P3_U7349 , P3_SUB_414_U62 , P3_U2602 );
nand NAND2_5541 ( P3_U7350 , P3_ADD_467_U70 , P3_U2601 );
nand NAND2_5542 ( P3_U7351 , P3_EBX_REG_30_ , P3_U7910 );
nand NAND2_5543 ( P3_U7352 , P3_ADD_430_U70 , P3_U2405 );
nand NAND2_5544 ( P3_U7353 , P3_U2403 , P3_ADD_318_U70 );
nand NAND2_5545 ( P3_U7354 , P3_SUB_320_U62 , P3_U4319 );
nand NAND2_5546 ( P3_U7355 , P3_U2401 , P3_PHYADDRPOINTER_REG_30_ );
nand NAND2_5547 ( P3_U7356 , P3_U7094 , P3_REIP_REG_30_ );
nand NAND2_5548 ( P3_U7357 , P3_U4135 , P3_U2603 );
nand NAND2_5549 ( P3_U7358 , P3_SUB_414_U51 , P3_U2602 );
nand NAND2_5550 ( P3_U7359 , P3_ADD_467_U69 , P3_U2601 );
nand NAND2_5551 ( P3_U7360 , P3_EBX_REG_31_ , P3_U7910 );
nand NAND2_5552 ( P3_U7361 , P3_ADD_430_U69 , P3_U2405 );
nand NAND2_5553 ( P3_U7362 , P3_U2403 , P3_ADD_318_U69 );
not NOT1_5554 ( P3_U7363 , P3_U7362 );
nand NAND2_5555 ( P3_U7364 , P3_U2401 , P3_PHYADDRPOINTER_REG_31_ );
nand NAND2_5556 ( P3_U7365 , P3_U7094 , P3_REIP_REG_31_ );
nand NAND2_5557 ( P3_U7366 , P3_DATAWIDTH_REG_1_ , P3_DATAWIDTH_REG_0_ );
or OR2_5558 ( P3_U7367 , P3_REIP_REG_1_ , P3_REIP_REG_0_ );
not NOT1_5559 ( P3_U7368 , P3_U4285 );
nand NAND2_5560 ( P3_U7369 , P3_FLUSH_REG , P3_U4285 );
nand NAND2_5561 ( P3_U7370 , P3_U4623 , P3_U2390 );
nand NAND2_5562 ( P3_U7371 , P3_U2453 , P3_U2630 );
nand NAND2_5563 ( P3_U7372 , P3_U3123 , P3_U7371 );
nand NAND2_5564 ( P3_U7373 , P3_U7372 , P3_U3121 );
not NOT1_5565 ( P3_U7374 , P3_U4287 );
nand NAND2_5566 ( P3_U7375 , P3_U4296 , P3_U2631 );
nand NAND2_5567 ( P3_U7376 , P3_U3112 , P3_U3118 );
nand NAND3_5568 ( P3_U7377 , P3_STATE2_REG_2_ , P3_U7919 , P3_U4150 );
nand NAND2_5569 ( P3_U7378 , P3_STATE2_REG_0_ , P3_U7377 );
nand NAND2_5570 ( P3_U7379 , P3_U3125 , P3_U7378 );
nand NAND2_5571 ( P3_U7380 , P3_U2390 , P3_U2604 );
nand NAND2_5572 ( P3_U7381 , P3_CODEFETCH_REG , P3_U7380 );
nand NAND2_5573 ( P3_U7382 , P3_U4347 , P3_STATE2_REG_0_ );
nand NAND2_5574 ( P3_U7383 , P3_ADS_N_REG , P3_STATE_REG_0_ );
not NOT1_5575 ( P3_U7384 , P3_U4288 );
nand NAND3_5576 ( P3_U7385 , P3_STATE2_REG_2_ , P3_U3111 , P3_U3114 );
nand NAND2_5577 ( P3_U7386 , P3_U4488 , P3_STATE2_REG_2_ );
nand NAND2_5578 ( P3_U7387 , P3_U2542 , P3_INSTQUEUE_REG_15__7_ );
nand NAND2_5579 ( P3_U7388 , P3_U2541 , P3_INSTQUEUE_REG_14__7_ );
nand NAND2_5580 ( P3_U7389 , P3_U2540 , P3_INSTQUEUE_REG_13__7_ );
nand NAND2_5581 ( P3_U7390 , P3_U2539 , P3_INSTQUEUE_REG_12__7_ );
nand NAND2_5582 ( P3_U7391 , P3_U2537 , P3_INSTQUEUE_REG_11__7_ );
nand NAND2_5583 ( P3_U7392 , P3_U2536 , P3_INSTQUEUE_REG_10__7_ );
nand NAND2_5584 ( P3_U7393 , P3_U2535 , P3_INSTQUEUE_REG_9__7_ );
nand NAND2_5585 ( P3_U7394 , P3_U2534 , P3_INSTQUEUE_REG_8__7_ );
nand NAND2_5586 ( P3_U7395 , P3_U2532 , P3_INSTQUEUE_REG_7__7_ );
nand NAND2_5587 ( P3_U7396 , P3_U2531 , P3_INSTQUEUE_REG_6__7_ );
nand NAND2_5588 ( P3_U7397 , P3_U2530 , P3_INSTQUEUE_REG_5__7_ );
nand NAND2_5589 ( P3_U7398 , P3_U2529 , P3_INSTQUEUE_REG_4__7_ );
nand NAND2_5590 ( P3_U7399 , P3_U2527 , P3_INSTQUEUE_REG_3__7_ );
nand NAND2_5591 ( P3_U7400 , P3_U2525 , P3_INSTQUEUE_REG_2__7_ );
nand NAND2_5592 ( P3_U7401 , P3_U2523 , P3_INSTQUEUE_REG_1__7_ );
nand NAND2_5593 ( P3_U7402 , P3_U2521 , P3_INSTQUEUE_REG_0__7_ );
nand NAND2_5594 ( P3_U7403 , P3_U2542 , P3_INSTQUEUE_REG_15__6_ );
nand NAND2_5595 ( P3_U7404 , P3_U2541 , P3_INSTQUEUE_REG_14__6_ );
nand NAND2_5596 ( P3_U7405 , P3_U2540 , P3_INSTQUEUE_REG_13__6_ );
nand NAND2_5597 ( P3_U7406 , P3_U2539 , P3_INSTQUEUE_REG_12__6_ );
nand NAND2_5598 ( P3_U7407 , P3_U2537 , P3_INSTQUEUE_REG_11__6_ );
nand NAND2_5599 ( P3_U7408 , P3_U2536 , P3_INSTQUEUE_REG_10__6_ );
nand NAND2_5600 ( P3_U7409 , P3_U2535 , P3_INSTQUEUE_REG_9__6_ );
nand NAND2_5601 ( P3_U7410 , P3_U2534 , P3_INSTQUEUE_REG_8__6_ );
nand NAND2_5602 ( P3_U7411 , P3_U2532 , P3_INSTQUEUE_REG_7__6_ );
nand NAND2_5603 ( P3_U7412 , P3_U2531 , P3_INSTQUEUE_REG_6__6_ );
nand NAND2_5604 ( P3_U7413 , P3_U2530 , P3_INSTQUEUE_REG_5__6_ );
nand NAND2_5605 ( P3_U7414 , P3_U2529 , P3_INSTQUEUE_REG_4__6_ );
nand NAND2_5606 ( P3_U7415 , P3_U2527 , P3_INSTQUEUE_REG_3__6_ );
nand NAND2_5607 ( P3_U7416 , P3_U2525 , P3_INSTQUEUE_REG_2__6_ );
nand NAND2_5608 ( P3_U7417 , P3_U2523 , P3_INSTQUEUE_REG_1__6_ );
nand NAND2_5609 ( P3_U7418 , P3_U2521 , P3_INSTQUEUE_REG_0__6_ );
nand NAND2_5610 ( P3_U7419 , P3_U2542 , P3_INSTQUEUE_REG_15__5_ );
nand NAND2_5611 ( P3_U7420 , P3_U2541 , P3_INSTQUEUE_REG_14__5_ );
nand NAND2_5612 ( P3_U7421 , P3_U2540 , P3_INSTQUEUE_REG_13__5_ );
nand NAND2_5613 ( P3_U7422 , P3_U2539 , P3_INSTQUEUE_REG_12__5_ );
nand NAND2_5614 ( P3_U7423 , P3_U2537 , P3_INSTQUEUE_REG_11__5_ );
nand NAND2_5615 ( P3_U7424 , P3_U2536 , P3_INSTQUEUE_REG_10__5_ );
nand NAND2_5616 ( P3_U7425 , P3_U2535 , P3_INSTQUEUE_REG_9__5_ );
nand NAND2_5617 ( P3_U7426 , P3_U2534 , P3_INSTQUEUE_REG_8__5_ );
nand NAND2_5618 ( P3_U7427 , P3_U2532 , P3_INSTQUEUE_REG_7__5_ );
nand NAND2_5619 ( P3_U7428 , P3_U2531 , P3_INSTQUEUE_REG_6__5_ );
nand NAND2_5620 ( P3_U7429 , P3_U2530 , P3_INSTQUEUE_REG_5__5_ );
nand NAND2_5621 ( P3_U7430 , P3_U2529 , P3_INSTQUEUE_REG_4__5_ );
nand NAND2_5622 ( P3_U7431 , P3_U2527 , P3_INSTQUEUE_REG_3__5_ );
nand NAND2_5623 ( P3_U7432 , P3_U2525 , P3_INSTQUEUE_REG_2__5_ );
nand NAND2_5624 ( P3_U7433 , P3_U2523 , P3_INSTQUEUE_REG_1__5_ );
nand NAND2_5625 ( P3_U7434 , P3_U2521 , P3_INSTQUEUE_REG_0__5_ );
nand NAND2_5626 ( P3_U7435 , P3_U2542 , P3_INSTQUEUE_REG_15__4_ );
nand NAND2_5627 ( P3_U7436 , P3_U2541 , P3_INSTQUEUE_REG_14__4_ );
nand NAND2_5628 ( P3_U7437 , P3_U2540 , P3_INSTQUEUE_REG_13__4_ );
nand NAND2_5629 ( P3_U7438 , P3_U2539 , P3_INSTQUEUE_REG_12__4_ );
nand NAND2_5630 ( P3_U7439 , P3_U2537 , P3_INSTQUEUE_REG_11__4_ );
nand NAND2_5631 ( P3_U7440 , P3_U2536 , P3_INSTQUEUE_REG_10__4_ );
nand NAND2_5632 ( P3_U7441 , P3_U2535 , P3_INSTQUEUE_REG_9__4_ );
nand NAND2_5633 ( P3_U7442 , P3_U2534 , P3_INSTQUEUE_REG_8__4_ );
nand NAND2_5634 ( P3_U7443 , P3_U2532 , P3_INSTQUEUE_REG_7__4_ );
nand NAND2_5635 ( P3_U7444 , P3_U2531 , P3_INSTQUEUE_REG_6__4_ );
nand NAND2_5636 ( P3_U7445 , P3_U2530 , P3_INSTQUEUE_REG_5__4_ );
nand NAND2_5637 ( P3_U7446 , P3_U2529 , P3_INSTQUEUE_REG_4__4_ );
nand NAND2_5638 ( P3_U7447 , P3_U2527 , P3_INSTQUEUE_REG_3__4_ );
nand NAND2_5639 ( P3_U7448 , P3_U2525 , P3_INSTQUEUE_REG_2__4_ );
nand NAND2_5640 ( P3_U7449 , P3_U2523 , P3_INSTQUEUE_REG_1__4_ );
nand NAND2_5641 ( P3_U7450 , P3_U2521 , P3_INSTQUEUE_REG_0__4_ );
nand NAND2_5642 ( P3_U7451 , P3_U2542 , P3_INSTQUEUE_REG_15__3_ );
nand NAND2_5643 ( P3_U7452 , P3_U2541 , P3_INSTQUEUE_REG_14__3_ );
nand NAND2_5644 ( P3_U7453 , P3_U2540 , P3_INSTQUEUE_REG_13__3_ );
nand NAND2_5645 ( P3_U7454 , P3_U2539 , P3_INSTQUEUE_REG_12__3_ );
nand NAND2_5646 ( P3_U7455 , P3_U2537 , P3_INSTQUEUE_REG_11__3_ );
nand NAND2_5647 ( P3_U7456 , P3_U2536 , P3_INSTQUEUE_REG_10__3_ );
nand NAND2_5648 ( P3_U7457 , P3_U2535 , P3_INSTQUEUE_REG_9__3_ );
nand NAND2_5649 ( P3_U7458 , P3_U2534 , P3_INSTQUEUE_REG_8__3_ );
nand NAND2_5650 ( P3_U7459 , P3_U2532 , P3_INSTQUEUE_REG_7__3_ );
nand NAND2_5651 ( P3_U7460 , P3_U2531 , P3_INSTQUEUE_REG_6__3_ );
nand NAND2_5652 ( P3_U7461 , P3_U2530 , P3_INSTQUEUE_REG_5__3_ );
nand NAND2_5653 ( P3_U7462 , P3_U2529 , P3_INSTQUEUE_REG_4__3_ );
nand NAND2_5654 ( P3_U7463 , P3_U2527 , P3_INSTQUEUE_REG_3__3_ );
nand NAND2_5655 ( P3_U7464 , P3_U2525 , P3_INSTQUEUE_REG_2__3_ );
nand NAND2_5656 ( P3_U7465 , P3_U2523 , P3_INSTQUEUE_REG_1__3_ );
nand NAND2_5657 ( P3_U7466 , P3_U2521 , P3_INSTQUEUE_REG_0__3_ );
nand NAND2_5658 ( P3_U7467 , P3_U2542 , P3_INSTQUEUE_REG_15__2_ );
nand NAND2_5659 ( P3_U7468 , P3_U2541 , P3_INSTQUEUE_REG_14__2_ );
nand NAND2_5660 ( P3_U7469 , P3_U2540 , P3_INSTQUEUE_REG_13__2_ );
nand NAND2_5661 ( P3_U7470 , P3_U2539 , P3_INSTQUEUE_REG_12__2_ );
nand NAND2_5662 ( P3_U7471 , P3_U2537 , P3_INSTQUEUE_REG_11__2_ );
nand NAND2_5663 ( P3_U7472 , P3_U2536 , P3_INSTQUEUE_REG_10__2_ );
nand NAND2_5664 ( P3_U7473 , P3_U2535 , P3_INSTQUEUE_REG_9__2_ );
nand NAND2_5665 ( P3_U7474 , P3_U2534 , P3_INSTQUEUE_REG_8__2_ );
nand NAND2_5666 ( P3_U7475 , P3_U2532 , P3_INSTQUEUE_REG_7__2_ );
nand NAND2_5667 ( P3_U7476 , P3_U2531 , P3_INSTQUEUE_REG_6__2_ );
nand NAND2_5668 ( P3_U7477 , P3_U2530 , P3_INSTQUEUE_REG_5__2_ );
nand NAND2_5669 ( P3_U7478 , P3_U2529 , P3_INSTQUEUE_REG_4__2_ );
nand NAND2_5670 ( P3_U7479 , P3_U2527 , P3_INSTQUEUE_REG_3__2_ );
nand NAND2_5671 ( P3_U7480 , P3_U2525 , P3_INSTQUEUE_REG_2__2_ );
nand NAND2_5672 ( P3_U7481 , P3_U2523 , P3_INSTQUEUE_REG_1__2_ );
nand NAND2_5673 ( P3_U7482 , P3_U2521 , P3_INSTQUEUE_REG_0__2_ );
nand NAND2_5674 ( P3_U7483 , P3_U2542 , P3_INSTQUEUE_REG_15__1_ );
nand NAND2_5675 ( P3_U7484 , P3_U2541 , P3_INSTQUEUE_REG_14__1_ );
nand NAND2_5676 ( P3_U7485 , P3_U2540 , P3_INSTQUEUE_REG_13__1_ );
nand NAND2_5677 ( P3_U7486 , P3_U2539 , P3_INSTQUEUE_REG_12__1_ );
nand NAND2_5678 ( P3_U7487 , P3_U2537 , P3_INSTQUEUE_REG_11__1_ );
nand NAND2_5679 ( P3_U7488 , P3_U2536 , P3_INSTQUEUE_REG_10__1_ );
nand NAND2_5680 ( P3_U7489 , P3_U2535 , P3_INSTQUEUE_REG_9__1_ );
nand NAND2_5681 ( P3_U7490 , P3_U2534 , P3_INSTQUEUE_REG_8__1_ );
nand NAND2_5682 ( P3_U7491 , P3_U2532 , P3_INSTQUEUE_REG_7__1_ );
nand NAND2_5683 ( P3_U7492 , P3_U2531 , P3_INSTQUEUE_REG_6__1_ );
nand NAND2_5684 ( P3_U7493 , P3_U2530 , P3_INSTQUEUE_REG_5__1_ );
nand NAND2_5685 ( P3_U7494 , P3_U2529 , P3_INSTQUEUE_REG_4__1_ );
nand NAND2_5686 ( P3_U7495 , P3_U2527 , P3_INSTQUEUE_REG_3__1_ );
nand NAND2_5687 ( P3_U7496 , P3_U2525 , P3_INSTQUEUE_REG_2__1_ );
nand NAND2_5688 ( P3_U7497 , P3_U2523 , P3_INSTQUEUE_REG_1__1_ );
nand NAND2_5689 ( P3_U7498 , P3_U2521 , P3_INSTQUEUE_REG_0__1_ );
nand NAND2_5690 ( P3_U7499 , P3_U2542 , P3_INSTQUEUE_REG_15__0_ );
nand NAND2_5691 ( P3_U7500 , P3_U2541 , P3_INSTQUEUE_REG_14__0_ );
nand NAND2_5692 ( P3_U7501 , P3_U2540 , P3_INSTQUEUE_REG_13__0_ );
nand NAND2_5693 ( P3_U7502 , P3_U2539 , P3_INSTQUEUE_REG_12__0_ );
nand NAND2_5694 ( P3_U7503 , P3_U2537 , P3_INSTQUEUE_REG_11__0_ );
nand NAND2_5695 ( P3_U7504 , P3_U2536 , P3_INSTQUEUE_REG_10__0_ );
nand NAND2_5696 ( P3_U7505 , P3_U2535 , P3_INSTQUEUE_REG_9__0_ );
nand NAND2_5697 ( P3_U7506 , P3_U2534 , P3_INSTQUEUE_REG_8__0_ );
nand NAND2_5698 ( P3_U7507 , P3_U2532 , P3_INSTQUEUE_REG_7__0_ );
nand NAND2_5699 ( P3_U7508 , P3_U2531 , P3_INSTQUEUE_REG_6__0_ );
nand NAND2_5700 ( P3_U7509 , P3_U2530 , P3_INSTQUEUE_REG_5__0_ );
nand NAND2_5701 ( P3_U7510 , P3_U2529 , P3_INSTQUEUE_REG_4__0_ );
nand NAND2_5702 ( P3_U7511 , P3_U2527 , P3_INSTQUEUE_REG_3__0_ );
nand NAND2_5703 ( P3_U7512 , P3_U2525 , P3_INSTQUEUE_REG_2__0_ );
nand NAND2_5704 ( P3_U7513 , P3_U2523 , P3_INSTQUEUE_REG_1__0_ );
nand NAND2_5705 ( P3_U7514 , P3_U2521 , P3_INSTQUEUE_REG_0__0_ );
nand NAND2_5706 ( P3_U7515 , P3_U4470 , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_5707 ( P3_U7516 , P3_U3266 );
nand NAND2_5708 ( P3_U7517 , P3_U2562 , P3_INSTQUEUE_REG_0__7_ );
nand NAND2_5709 ( P3_U7518 , P3_U2561 , P3_INSTQUEUE_REG_1__7_ );
nand NAND2_5710 ( P3_U7519 , P3_U2560 , P3_INSTQUEUE_REG_2__7_ );
nand NAND2_5711 ( P3_U7520 , P3_U2559 , P3_INSTQUEUE_REG_3__7_ );
nand NAND2_5712 ( P3_U7521 , P3_U2557 , P3_INSTQUEUE_REG_4__7_ );
nand NAND2_5713 ( P3_U7522 , P3_U2556 , P3_INSTQUEUE_REG_5__7_ );
nand NAND2_5714 ( P3_U7523 , P3_U2555 , P3_INSTQUEUE_REG_6__7_ );
nand NAND2_5715 ( P3_U7524 , P3_U2554 , P3_INSTQUEUE_REG_7__7_ );
nand NAND2_5716 ( P3_U7525 , P3_U2552 , P3_INSTQUEUE_REG_8__7_ );
nand NAND2_5717 ( P3_U7526 , P3_U2551 , P3_INSTQUEUE_REG_9__7_ );
nand NAND2_5718 ( P3_U7527 , P3_U2550 , P3_INSTQUEUE_REG_10__7_ );
nand NAND2_5719 ( P3_U7528 , P3_U2549 , P3_INSTQUEUE_REG_11__7_ );
nand NAND2_5720 ( P3_U7529 , P3_U2547 , P3_INSTQUEUE_REG_12__7_ );
nand NAND2_5721 ( P3_U7530 , P3_U2546 , P3_INSTQUEUE_REG_13__7_ );
nand NAND2_5722 ( P3_U7531 , P3_U2545 , P3_INSTQUEUE_REG_14__7_ );
nand NAND2_5723 ( P3_U7532 , P3_U2544 , P3_INSTQUEUE_REG_15__7_ );
nand NAND2_5724 ( P3_U7533 , P3_U2562 , P3_INSTQUEUE_REG_0__6_ );
nand NAND2_5725 ( P3_U7534 , P3_U2561 , P3_INSTQUEUE_REG_1__6_ );
nand NAND2_5726 ( P3_U7535 , P3_U2560 , P3_INSTQUEUE_REG_2__6_ );
nand NAND2_5727 ( P3_U7536 , P3_U2559 , P3_INSTQUEUE_REG_3__6_ );
nand NAND2_5728 ( P3_U7537 , P3_U2557 , P3_INSTQUEUE_REG_4__6_ );
nand NAND2_5729 ( P3_U7538 , P3_U2556 , P3_INSTQUEUE_REG_5__6_ );
nand NAND2_5730 ( P3_U7539 , P3_U2555 , P3_INSTQUEUE_REG_6__6_ );
nand NAND2_5731 ( P3_U7540 , P3_U2554 , P3_INSTQUEUE_REG_7__6_ );
nand NAND2_5732 ( P3_U7541 , P3_U2552 , P3_INSTQUEUE_REG_8__6_ );
nand NAND2_5733 ( P3_U7542 , P3_U2551 , P3_INSTQUEUE_REG_9__6_ );
nand NAND2_5734 ( P3_U7543 , P3_U2550 , P3_INSTQUEUE_REG_10__6_ );
nand NAND2_5735 ( P3_U7544 , P3_U2549 , P3_INSTQUEUE_REG_11__6_ );
nand NAND2_5736 ( P3_U7545 , P3_U2547 , P3_INSTQUEUE_REG_12__6_ );
nand NAND2_5737 ( P3_U7546 , P3_U2546 , P3_INSTQUEUE_REG_13__6_ );
nand NAND2_5738 ( P3_U7547 , P3_U2545 , P3_INSTQUEUE_REG_14__6_ );
nand NAND2_5739 ( P3_U7548 , P3_U2544 , P3_INSTQUEUE_REG_15__6_ );
nand NAND2_5740 ( P3_U7549 , P3_U2562 , P3_INSTQUEUE_REG_0__5_ );
nand NAND2_5741 ( P3_U7550 , P3_U2561 , P3_INSTQUEUE_REG_1__5_ );
nand NAND2_5742 ( P3_U7551 , P3_U2560 , P3_INSTQUEUE_REG_2__5_ );
nand NAND2_5743 ( P3_U7552 , P3_U2559 , P3_INSTQUEUE_REG_3__5_ );
nand NAND2_5744 ( P3_U7553 , P3_U2557 , P3_INSTQUEUE_REG_4__5_ );
nand NAND2_5745 ( P3_U7554 , P3_U2556 , P3_INSTQUEUE_REG_5__5_ );
nand NAND2_5746 ( P3_U7555 , P3_U2555 , P3_INSTQUEUE_REG_6__5_ );
nand NAND2_5747 ( P3_U7556 , P3_U2554 , P3_INSTQUEUE_REG_7__5_ );
nand NAND2_5748 ( P3_U7557 , P3_U2552 , P3_INSTQUEUE_REG_8__5_ );
nand NAND2_5749 ( P3_U7558 , P3_U2551 , P3_INSTQUEUE_REG_9__5_ );
nand NAND2_5750 ( P3_U7559 , P3_U2550 , P3_INSTQUEUE_REG_10__5_ );
nand NAND2_5751 ( P3_U7560 , P3_U2549 , P3_INSTQUEUE_REG_11__5_ );
nand NAND2_5752 ( P3_U7561 , P3_U2547 , P3_INSTQUEUE_REG_12__5_ );
nand NAND2_5753 ( P3_U7562 , P3_U2546 , P3_INSTQUEUE_REG_13__5_ );
nand NAND2_5754 ( P3_U7563 , P3_U2545 , P3_INSTQUEUE_REG_14__5_ );
nand NAND2_5755 ( P3_U7564 , P3_U2544 , P3_INSTQUEUE_REG_15__5_ );
nand NAND2_5756 ( P3_U7565 , P3_U2562 , P3_INSTQUEUE_REG_0__4_ );
nand NAND2_5757 ( P3_U7566 , P3_U2561 , P3_INSTQUEUE_REG_1__4_ );
nand NAND2_5758 ( P3_U7567 , P3_U2560 , P3_INSTQUEUE_REG_2__4_ );
nand NAND2_5759 ( P3_U7568 , P3_U2559 , P3_INSTQUEUE_REG_3__4_ );
nand NAND2_5760 ( P3_U7569 , P3_U2557 , P3_INSTQUEUE_REG_4__4_ );
nand NAND2_5761 ( P3_U7570 , P3_U2556 , P3_INSTQUEUE_REG_5__4_ );
nand NAND2_5762 ( P3_U7571 , P3_U2555 , P3_INSTQUEUE_REG_6__4_ );
nand NAND2_5763 ( P3_U7572 , P3_U2554 , P3_INSTQUEUE_REG_7__4_ );
nand NAND2_5764 ( P3_U7573 , P3_U2552 , P3_INSTQUEUE_REG_8__4_ );
nand NAND2_5765 ( P3_U7574 , P3_U2551 , P3_INSTQUEUE_REG_9__4_ );
nand NAND2_5766 ( P3_U7575 , P3_U2550 , P3_INSTQUEUE_REG_10__4_ );
nand NAND2_5767 ( P3_U7576 , P3_U2549 , P3_INSTQUEUE_REG_11__4_ );
nand NAND2_5768 ( P3_U7577 , P3_U2547 , P3_INSTQUEUE_REG_12__4_ );
nand NAND2_5769 ( P3_U7578 , P3_U2546 , P3_INSTQUEUE_REG_13__4_ );
nand NAND2_5770 ( P3_U7579 , P3_U2545 , P3_INSTQUEUE_REG_14__4_ );
nand NAND2_5771 ( P3_U7580 , P3_U2544 , P3_INSTQUEUE_REG_15__4_ );
nand NAND2_5772 ( P3_U7581 , P3_U2562 , P3_INSTQUEUE_REG_0__3_ );
nand NAND2_5773 ( P3_U7582 , P3_U2561 , P3_INSTQUEUE_REG_1__3_ );
nand NAND2_5774 ( P3_U7583 , P3_U2560 , P3_INSTQUEUE_REG_2__3_ );
nand NAND2_5775 ( P3_U7584 , P3_U2559 , P3_INSTQUEUE_REG_3__3_ );
nand NAND2_5776 ( P3_U7585 , P3_U2557 , P3_INSTQUEUE_REG_4__3_ );
nand NAND2_5777 ( P3_U7586 , P3_U2556 , P3_INSTQUEUE_REG_5__3_ );
nand NAND2_5778 ( P3_U7587 , P3_U2555 , P3_INSTQUEUE_REG_6__3_ );
nand NAND2_5779 ( P3_U7588 , P3_U2554 , P3_INSTQUEUE_REG_7__3_ );
nand NAND2_5780 ( P3_U7589 , P3_U2552 , P3_INSTQUEUE_REG_8__3_ );
nand NAND2_5781 ( P3_U7590 , P3_U2551 , P3_INSTQUEUE_REG_9__3_ );
nand NAND2_5782 ( P3_U7591 , P3_U2550 , P3_INSTQUEUE_REG_10__3_ );
nand NAND2_5783 ( P3_U7592 , P3_U2549 , P3_INSTQUEUE_REG_11__3_ );
nand NAND2_5784 ( P3_U7593 , P3_U2547 , P3_INSTQUEUE_REG_12__3_ );
nand NAND2_5785 ( P3_U7594 , P3_U2546 , P3_INSTQUEUE_REG_13__3_ );
nand NAND2_5786 ( P3_U7595 , P3_U2545 , P3_INSTQUEUE_REG_14__3_ );
nand NAND2_5787 ( P3_U7596 , P3_U2544 , P3_INSTQUEUE_REG_15__3_ );
nand NAND2_5788 ( P3_U7597 , P3_U2562 , P3_INSTQUEUE_REG_0__2_ );
nand NAND2_5789 ( P3_U7598 , P3_U2561 , P3_INSTQUEUE_REG_1__2_ );
nand NAND2_5790 ( P3_U7599 , P3_U2560 , P3_INSTQUEUE_REG_2__2_ );
nand NAND2_5791 ( P3_U7600 , P3_U2559 , P3_INSTQUEUE_REG_3__2_ );
nand NAND2_5792 ( P3_U7601 , P3_U2557 , P3_INSTQUEUE_REG_4__2_ );
nand NAND2_5793 ( P3_U7602 , P3_U2556 , P3_INSTQUEUE_REG_5__2_ );
nand NAND2_5794 ( P3_U7603 , P3_U2555 , P3_INSTQUEUE_REG_6__2_ );
nand NAND2_5795 ( P3_U7604 , P3_U2554 , P3_INSTQUEUE_REG_7__2_ );
nand NAND2_5796 ( P3_U7605 , P3_U2552 , P3_INSTQUEUE_REG_8__2_ );
nand NAND2_5797 ( P3_U7606 , P3_U2551 , P3_INSTQUEUE_REG_9__2_ );
nand NAND2_5798 ( P3_U7607 , P3_U2550 , P3_INSTQUEUE_REG_10__2_ );
nand NAND2_5799 ( P3_U7608 , P3_U2549 , P3_INSTQUEUE_REG_11__2_ );
nand NAND2_5800 ( P3_U7609 , P3_U2547 , P3_INSTQUEUE_REG_12__2_ );
nand NAND2_5801 ( P3_U7610 , P3_U2546 , P3_INSTQUEUE_REG_13__2_ );
nand NAND2_5802 ( P3_U7611 , P3_U2545 , P3_INSTQUEUE_REG_14__2_ );
nand NAND2_5803 ( P3_U7612 , P3_U2544 , P3_INSTQUEUE_REG_15__2_ );
nand NAND2_5804 ( P3_U7613 , P3_U2562 , P3_INSTQUEUE_REG_0__1_ );
nand NAND2_5805 ( P3_U7614 , P3_U2561 , P3_INSTQUEUE_REG_1__1_ );
nand NAND2_5806 ( P3_U7615 , P3_U2560 , P3_INSTQUEUE_REG_2__1_ );
nand NAND2_5807 ( P3_U7616 , P3_U2559 , P3_INSTQUEUE_REG_3__1_ );
nand NAND2_5808 ( P3_U7617 , P3_U2557 , P3_INSTQUEUE_REG_4__1_ );
nand NAND2_5809 ( P3_U7618 , P3_U2556 , P3_INSTQUEUE_REG_5__1_ );
nand NAND2_5810 ( P3_U7619 , P3_U2555 , P3_INSTQUEUE_REG_6__1_ );
nand NAND2_5811 ( P3_U7620 , P3_U2554 , P3_INSTQUEUE_REG_7__1_ );
nand NAND2_5812 ( P3_U7621 , P3_U2552 , P3_INSTQUEUE_REG_8__1_ );
nand NAND2_5813 ( P3_U7622 , P3_U2551 , P3_INSTQUEUE_REG_9__1_ );
nand NAND2_5814 ( P3_U7623 , P3_U2550 , P3_INSTQUEUE_REG_10__1_ );
nand NAND2_5815 ( P3_U7624 , P3_U2549 , P3_INSTQUEUE_REG_11__1_ );
nand NAND2_5816 ( P3_U7625 , P3_U2547 , P3_INSTQUEUE_REG_12__1_ );
nand NAND2_5817 ( P3_U7626 , P3_U2546 , P3_INSTQUEUE_REG_13__1_ );
nand NAND2_5818 ( P3_U7627 , P3_U2545 , P3_INSTQUEUE_REG_14__1_ );
nand NAND2_5819 ( P3_U7628 , P3_U2544 , P3_INSTQUEUE_REG_15__1_ );
nand NAND2_5820 ( P3_U7629 , P3_U2562 , P3_INSTQUEUE_REG_0__0_ );
nand NAND2_5821 ( P3_U7630 , P3_U2561 , P3_INSTQUEUE_REG_1__0_ );
nand NAND2_5822 ( P3_U7631 , P3_U2560 , P3_INSTQUEUE_REG_2__0_ );
nand NAND2_5823 ( P3_U7632 , P3_U2559 , P3_INSTQUEUE_REG_3__0_ );
nand NAND2_5824 ( P3_U7633 , P3_U2557 , P3_INSTQUEUE_REG_4__0_ );
nand NAND2_5825 ( P3_U7634 , P3_U2556 , P3_INSTQUEUE_REG_5__0_ );
nand NAND2_5826 ( P3_U7635 , P3_U2555 , P3_INSTQUEUE_REG_6__0_ );
nand NAND2_5827 ( P3_U7636 , P3_U2554 , P3_INSTQUEUE_REG_7__0_ );
nand NAND2_5828 ( P3_U7637 , P3_U2552 , P3_INSTQUEUE_REG_8__0_ );
nand NAND2_5829 ( P3_U7638 , P3_U2551 , P3_INSTQUEUE_REG_9__0_ );
nand NAND2_5830 ( P3_U7639 , P3_U2550 , P3_INSTQUEUE_REG_10__0_ );
nand NAND2_5831 ( P3_U7640 , P3_U2549 , P3_INSTQUEUE_REG_11__0_ );
nand NAND2_5832 ( P3_U7641 , P3_U2547 , P3_INSTQUEUE_REG_12__0_ );
nand NAND2_5833 ( P3_U7642 , P3_U2546 , P3_INSTQUEUE_REG_13__0_ );
nand NAND2_5834 ( P3_U7643 , P3_U2545 , P3_INSTQUEUE_REG_14__0_ );
nand NAND2_5835 ( P3_U7644 , P3_U2544 , P3_INSTQUEUE_REG_15__0_ );
not NOT1_5836 ( P3_U7645 , P3_U4289 );
nand NAND2_5837 ( P3_U7646 , P3_U2582 , P3_INSTQUEUE_REG_8__7_ );
nand NAND2_5838 ( P3_U7647 , P3_U2581 , P3_INSTQUEUE_REG_9__7_ );
nand NAND2_5839 ( P3_U7648 , P3_U2580 , P3_INSTQUEUE_REG_10__7_ );
nand NAND2_5840 ( P3_U7649 , P3_U2579 , P3_INSTQUEUE_REG_11__7_ );
nand NAND2_5841 ( P3_U7650 , P3_U2577 , P3_INSTQUEUE_REG_12__7_ );
nand NAND2_5842 ( P3_U7651 , P3_U2576 , P3_INSTQUEUE_REG_13__7_ );
nand NAND2_5843 ( P3_U7652 , P3_U2575 , P3_INSTQUEUE_REG_14__7_ );
nand NAND2_5844 ( P3_U7653 , P3_U2574 , P3_INSTQUEUE_REG_15__7_ );
nand NAND2_5845 ( P3_U7654 , P3_U2572 , P3_INSTQUEUE_REG_0__7_ );
nand NAND2_5846 ( P3_U7655 , P3_U2571 , P3_INSTQUEUE_REG_1__7_ );
nand NAND2_5847 ( P3_U7656 , P3_U2570 , P3_INSTQUEUE_REG_2__7_ );
nand NAND2_5848 ( P3_U7657 , P3_U2569 , P3_INSTQUEUE_REG_3__7_ );
nand NAND2_5849 ( P3_U7658 , P3_U2567 , P3_INSTQUEUE_REG_4__7_ );
nand NAND2_5850 ( P3_U7659 , P3_U2566 , P3_INSTQUEUE_REG_5__7_ );
nand NAND2_5851 ( P3_U7660 , P3_U2565 , P3_INSTQUEUE_REG_6__7_ );
nand NAND2_5852 ( P3_U7661 , P3_U2564 , P3_INSTQUEUE_REG_7__7_ );
nand NAND2_5853 ( P3_U7662 , P3_U2582 , P3_INSTQUEUE_REG_8__6_ );
nand NAND2_5854 ( P3_U7663 , P3_U2581 , P3_INSTQUEUE_REG_9__6_ );
nand NAND2_5855 ( P3_U7664 , P3_U2580 , P3_INSTQUEUE_REG_10__6_ );
nand NAND2_5856 ( P3_U7665 , P3_U2579 , P3_INSTQUEUE_REG_11__6_ );
nand NAND2_5857 ( P3_U7666 , P3_U2577 , P3_INSTQUEUE_REG_12__6_ );
nand NAND2_5858 ( P3_U7667 , P3_U2576 , P3_INSTQUEUE_REG_13__6_ );
nand NAND2_5859 ( P3_U7668 , P3_U2575 , P3_INSTQUEUE_REG_14__6_ );
nand NAND2_5860 ( P3_U7669 , P3_U2574 , P3_INSTQUEUE_REG_15__6_ );
nand NAND2_5861 ( P3_U7670 , P3_U2572 , P3_INSTQUEUE_REG_0__6_ );
nand NAND2_5862 ( P3_U7671 , P3_U2571 , P3_INSTQUEUE_REG_1__6_ );
nand NAND2_5863 ( P3_U7672 , P3_U2570 , P3_INSTQUEUE_REG_2__6_ );
nand NAND2_5864 ( P3_U7673 , P3_U2569 , P3_INSTQUEUE_REG_3__6_ );
nand NAND2_5865 ( P3_U7674 , P3_U2567 , P3_INSTQUEUE_REG_4__6_ );
nand NAND2_5866 ( P3_U7675 , P3_U2566 , P3_INSTQUEUE_REG_5__6_ );
nand NAND2_5867 ( P3_U7676 , P3_U2565 , P3_INSTQUEUE_REG_6__6_ );
nand NAND2_5868 ( P3_U7677 , P3_U2564 , P3_INSTQUEUE_REG_7__6_ );
nand NAND2_5869 ( P3_U7678 , P3_U2582 , P3_INSTQUEUE_REG_8__5_ );
nand NAND2_5870 ( P3_U7679 , P3_U2581 , P3_INSTQUEUE_REG_9__5_ );
nand NAND2_5871 ( P3_U7680 , P3_U2580 , P3_INSTQUEUE_REG_10__5_ );
nand NAND2_5872 ( P3_U7681 , P3_U2579 , P3_INSTQUEUE_REG_11__5_ );
nand NAND2_5873 ( P3_U7682 , P3_U2577 , P3_INSTQUEUE_REG_12__5_ );
nand NAND2_5874 ( P3_U7683 , P3_U2576 , P3_INSTQUEUE_REG_13__5_ );
nand NAND2_5875 ( P3_U7684 , P3_U2575 , P3_INSTQUEUE_REG_14__5_ );
nand NAND2_5876 ( P3_U7685 , P3_U2574 , P3_INSTQUEUE_REG_15__5_ );
nand NAND2_5877 ( P3_U7686 , P3_U2572 , P3_INSTQUEUE_REG_0__5_ );
nand NAND2_5878 ( P3_U7687 , P3_U2571 , P3_INSTQUEUE_REG_1__5_ );
nand NAND2_5879 ( P3_U7688 , P3_U2570 , P3_INSTQUEUE_REG_2__5_ );
nand NAND2_5880 ( P3_U7689 , P3_U2569 , P3_INSTQUEUE_REG_3__5_ );
nand NAND2_5881 ( P3_U7690 , P3_U2567 , P3_INSTQUEUE_REG_4__5_ );
nand NAND2_5882 ( P3_U7691 , P3_U2566 , P3_INSTQUEUE_REG_5__5_ );
nand NAND2_5883 ( P3_U7692 , P3_U2565 , P3_INSTQUEUE_REG_6__5_ );
nand NAND2_5884 ( P3_U7693 , P3_U2564 , P3_INSTQUEUE_REG_7__5_ );
nand NAND2_5885 ( P3_U7694 , P3_U2582 , P3_INSTQUEUE_REG_8__4_ );
nand NAND2_5886 ( P3_U7695 , P3_U2581 , P3_INSTQUEUE_REG_9__4_ );
nand NAND2_5887 ( P3_U7696 , P3_U2580 , P3_INSTQUEUE_REG_10__4_ );
nand NAND2_5888 ( P3_U7697 , P3_U2579 , P3_INSTQUEUE_REG_11__4_ );
nand NAND2_5889 ( P3_U7698 , P3_U2577 , P3_INSTQUEUE_REG_12__4_ );
nand NAND2_5890 ( P3_U7699 , P3_U2576 , P3_INSTQUEUE_REG_13__4_ );
nand NAND2_5891 ( P3_U7700 , P3_U2575 , P3_INSTQUEUE_REG_14__4_ );
nand NAND2_5892 ( P3_U7701 , P3_U2574 , P3_INSTQUEUE_REG_15__4_ );
nand NAND2_5893 ( P3_U7702 , P3_U2572 , P3_INSTQUEUE_REG_0__4_ );
nand NAND2_5894 ( P3_U7703 , P3_U2571 , P3_INSTQUEUE_REG_1__4_ );
nand NAND2_5895 ( P3_U7704 , P3_U2570 , P3_INSTQUEUE_REG_2__4_ );
nand NAND2_5896 ( P3_U7705 , P3_U2569 , P3_INSTQUEUE_REG_3__4_ );
nand NAND2_5897 ( P3_U7706 , P3_U2567 , P3_INSTQUEUE_REG_4__4_ );
nand NAND2_5898 ( P3_U7707 , P3_U2566 , P3_INSTQUEUE_REG_5__4_ );
nand NAND2_5899 ( P3_U7708 , P3_U2565 , P3_INSTQUEUE_REG_6__4_ );
nand NAND2_5900 ( P3_U7709 , P3_U2564 , P3_INSTQUEUE_REG_7__4_ );
nand NAND2_5901 ( P3_U7710 , P3_U2582 , P3_INSTQUEUE_REG_8__3_ );
nand NAND2_5902 ( P3_U7711 , P3_U2581 , P3_INSTQUEUE_REG_9__3_ );
nand NAND2_5903 ( P3_U7712 , P3_U2580 , P3_INSTQUEUE_REG_10__3_ );
nand NAND2_5904 ( P3_U7713 , P3_U2579 , P3_INSTQUEUE_REG_11__3_ );
nand NAND2_5905 ( P3_U7714 , P3_U2577 , P3_INSTQUEUE_REG_12__3_ );
nand NAND2_5906 ( P3_U7715 , P3_U2576 , P3_INSTQUEUE_REG_13__3_ );
nand NAND2_5907 ( P3_U7716 , P3_U2575 , P3_INSTQUEUE_REG_14__3_ );
nand NAND2_5908 ( P3_U7717 , P3_U2574 , P3_INSTQUEUE_REG_15__3_ );
nand NAND2_5909 ( P3_U7718 , P3_U2572 , P3_INSTQUEUE_REG_0__3_ );
nand NAND2_5910 ( P3_U7719 , P3_U2571 , P3_INSTQUEUE_REG_1__3_ );
nand NAND2_5911 ( P3_U7720 , P3_U2570 , P3_INSTQUEUE_REG_2__3_ );
nand NAND2_5912 ( P3_U7721 , P3_U2569 , P3_INSTQUEUE_REG_3__3_ );
nand NAND2_5913 ( P3_U7722 , P3_U2567 , P3_INSTQUEUE_REG_4__3_ );
nand NAND2_5914 ( P3_U7723 , P3_U2566 , P3_INSTQUEUE_REG_5__3_ );
nand NAND2_5915 ( P3_U7724 , P3_U2565 , P3_INSTQUEUE_REG_6__3_ );
nand NAND2_5916 ( P3_U7725 , P3_U2564 , P3_INSTQUEUE_REG_7__3_ );
nand NAND2_5917 ( P3_U7726 , P3_U2582 , P3_INSTQUEUE_REG_8__2_ );
nand NAND2_5918 ( P3_U7727 , P3_U2581 , P3_INSTQUEUE_REG_9__2_ );
nand NAND2_5919 ( P3_U7728 , P3_U2580 , P3_INSTQUEUE_REG_10__2_ );
nand NAND2_5920 ( P3_U7729 , P3_U2579 , P3_INSTQUEUE_REG_11__2_ );
nand NAND2_5921 ( P3_U7730 , P3_U2577 , P3_INSTQUEUE_REG_12__2_ );
nand NAND2_5922 ( P3_U7731 , P3_U2576 , P3_INSTQUEUE_REG_13__2_ );
nand NAND2_5923 ( P3_U7732 , P3_U2575 , P3_INSTQUEUE_REG_14__2_ );
nand NAND2_5924 ( P3_U7733 , P3_U2574 , P3_INSTQUEUE_REG_15__2_ );
nand NAND2_5925 ( P3_U7734 , P3_U2572 , P3_INSTQUEUE_REG_0__2_ );
nand NAND2_5926 ( P3_U7735 , P3_U2571 , P3_INSTQUEUE_REG_1__2_ );
nand NAND2_5927 ( P3_U7736 , P3_U2570 , P3_INSTQUEUE_REG_2__2_ );
nand NAND2_5928 ( P3_U7737 , P3_U2569 , P3_INSTQUEUE_REG_3__2_ );
nand NAND2_5929 ( P3_U7738 , P3_U2567 , P3_INSTQUEUE_REG_4__2_ );
nand NAND2_5930 ( P3_U7739 , P3_U2566 , P3_INSTQUEUE_REG_5__2_ );
nand NAND2_5931 ( P3_U7740 , P3_U2565 , P3_INSTQUEUE_REG_6__2_ );
nand NAND2_5932 ( P3_U7741 , P3_U2564 , P3_INSTQUEUE_REG_7__2_ );
nand NAND2_5933 ( P3_U7742 , P3_U2582 , P3_INSTQUEUE_REG_8__1_ );
nand NAND2_5934 ( P3_U7743 , P3_U2581 , P3_INSTQUEUE_REG_9__1_ );
nand NAND2_5935 ( P3_U7744 , P3_U2580 , P3_INSTQUEUE_REG_10__1_ );
nand NAND2_5936 ( P3_U7745 , P3_U2579 , P3_INSTQUEUE_REG_11__1_ );
nand NAND2_5937 ( P3_U7746 , P3_U2577 , P3_INSTQUEUE_REG_12__1_ );
nand NAND2_5938 ( P3_U7747 , P3_U2576 , P3_INSTQUEUE_REG_13__1_ );
nand NAND2_5939 ( P3_U7748 , P3_U2575 , P3_INSTQUEUE_REG_14__1_ );
nand NAND2_5940 ( P3_U7749 , P3_U2574 , P3_INSTQUEUE_REG_15__1_ );
nand NAND2_5941 ( P3_U7750 , P3_U2572 , P3_INSTQUEUE_REG_0__1_ );
nand NAND2_5942 ( P3_U7751 , P3_U2571 , P3_INSTQUEUE_REG_1__1_ );
nand NAND2_5943 ( P3_U7752 , P3_U2570 , P3_INSTQUEUE_REG_2__1_ );
nand NAND2_5944 ( P3_U7753 , P3_U2569 , P3_INSTQUEUE_REG_3__1_ );
nand NAND2_5945 ( P3_U7754 , P3_U2567 , P3_INSTQUEUE_REG_4__1_ );
nand NAND2_5946 ( P3_U7755 , P3_U2566 , P3_INSTQUEUE_REG_5__1_ );
nand NAND2_5947 ( P3_U7756 , P3_U2565 , P3_INSTQUEUE_REG_6__1_ );
nand NAND2_5948 ( P3_U7757 , P3_U2564 , P3_INSTQUEUE_REG_7__1_ );
nand NAND2_5949 ( P3_U7758 , P3_U2582 , P3_INSTQUEUE_REG_8__0_ );
nand NAND2_5950 ( P3_U7759 , P3_U2581 , P3_INSTQUEUE_REG_9__0_ );
nand NAND2_5951 ( P3_U7760 , P3_U2580 , P3_INSTQUEUE_REG_10__0_ );
nand NAND2_5952 ( P3_U7761 , P3_U2579 , P3_INSTQUEUE_REG_11__0_ );
nand NAND2_5953 ( P3_U7762 , P3_U2577 , P3_INSTQUEUE_REG_12__0_ );
nand NAND2_5954 ( P3_U7763 , P3_U2576 , P3_INSTQUEUE_REG_13__0_ );
nand NAND2_5955 ( P3_U7764 , P3_U2575 , P3_INSTQUEUE_REG_14__0_ );
nand NAND2_5956 ( P3_U7765 , P3_U2574 , P3_INSTQUEUE_REG_15__0_ );
nand NAND2_5957 ( P3_U7766 , P3_U2572 , P3_INSTQUEUE_REG_0__0_ );
nand NAND2_5958 ( P3_U7767 , P3_U2571 , P3_INSTQUEUE_REG_1__0_ );
nand NAND2_5959 ( P3_U7768 , P3_U2570 , P3_INSTQUEUE_REG_2__0_ );
nand NAND2_5960 ( P3_U7769 , P3_U2569 , P3_INSTQUEUE_REG_3__0_ );
nand NAND2_5961 ( P3_U7770 , P3_U2567 , P3_INSTQUEUE_REG_4__0_ );
nand NAND2_5962 ( P3_U7771 , P3_U2566 , P3_INSTQUEUE_REG_5__0_ );
nand NAND2_5963 ( P3_U7772 , P3_U2565 , P3_INSTQUEUE_REG_6__0_ );
nand NAND2_5964 ( P3_U7773 , P3_U2564 , P3_INSTQUEUE_REG_7__0_ );
nand NAND2_5965 ( P3_U7774 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_U3097 );
not NOT1_5966 ( P3_U7775 , P3_U3268 );
nand NAND2_5967 ( P3_U7776 , P3_U2600 , P3_INSTQUEUE_REG_8__7_ );
nand NAND2_5968 ( P3_U7777 , P3_U2599 , P3_INSTQUEUE_REG_9__7_ );
nand NAND2_5969 ( P3_U7778 , P3_U2598 , P3_INSTQUEUE_REG_10__7_ );
nand NAND2_5970 ( P3_U7779 , P3_U2597 , P3_INSTQUEUE_REG_11__7_ );
nand NAND2_5971 ( P3_U7780 , P3_U2595 , P3_INSTQUEUE_REG_12__7_ );
nand NAND2_5972 ( P3_U7781 , P3_U2594 , P3_INSTQUEUE_REG_13__7_ );
nand NAND2_5973 ( P3_U7782 , P3_U2593 , P3_INSTQUEUE_REG_14__7_ );
nand NAND2_5974 ( P3_U7783 , P3_U2592 , P3_INSTQUEUE_REG_15__7_ );
nand NAND2_5975 ( P3_U7784 , P3_U2591 , P3_INSTQUEUE_REG_0__7_ );
nand NAND2_5976 ( P3_U7785 , P3_U2590 , P3_INSTQUEUE_REG_1__7_ );
nand NAND2_5977 ( P3_U7786 , P3_U2589 , P3_INSTQUEUE_REG_2__7_ );
nand NAND2_5978 ( P3_U7787 , P3_U2588 , P3_INSTQUEUE_REG_3__7_ );
nand NAND2_5979 ( P3_U7788 , P3_U2586 , P3_INSTQUEUE_REG_4__7_ );
nand NAND2_5980 ( P3_U7789 , P3_U2585 , P3_INSTQUEUE_REG_5__7_ );
nand NAND2_5981 ( P3_U7790 , P3_U2584 , P3_INSTQUEUE_REG_6__7_ );
nand NAND2_5982 ( P3_U7791 , P3_U2583 , P3_INSTQUEUE_REG_7__7_ );
nand NAND2_5983 ( P3_U7792 , P3_U2600 , P3_INSTQUEUE_REG_8__6_ );
nand NAND2_5984 ( P3_U7793 , P3_U2599 , P3_INSTQUEUE_REG_9__6_ );
nand NAND2_5985 ( P3_U7794 , P3_U2598 , P3_INSTQUEUE_REG_10__6_ );
nand NAND2_5986 ( P3_U7795 , P3_U2597 , P3_INSTQUEUE_REG_11__6_ );
nand NAND2_5987 ( P3_U7796 , P3_U2595 , P3_INSTQUEUE_REG_12__6_ );
nand NAND2_5988 ( P3_U7797 , P3_U2594 , P3_INSTQUEUE_REG_13__6_ );
nand NAND2_5989 ( P3_U7798 , P3_U2593 , P3_INSTQUEUE_REG_14__6_ );
nand NAND2_5990 ( P3_U7799 , P3_U2592 , P3_INSTQUEUE_REG_15__6_ );
nand NAND2_5991 ( P3_U7800 , P3_U2591 , P3_INSTQUEUE_REG_0__6_ );
nand NAND2_5992 ( P3_U7801 , P3_U2590 , P3_INSTQUEUE_REG_1__6_ );
nand NAND2_5993 ( P3_U7802 , P3_U2589 , P3_INSTQUEUE_REG_2__6_ );
nand NAND2_5994 ( P3_U7803 , P3_U2588 , P3_INSTQUEUE_REG_3__6_ );
nand NAND2_5995 ( P3_U7804 , P3_U2586 , P3_INSTQUEUE_REG_4__6_ );
nand NAND2_5996 ( P3_U7805 , P3_U2585 , P3_INSTQUEUE_REG_5__6_ );
nand NAND2_5997 ( P3_U7806 , P3_U2584 , P3_INSTQUEUE_REG_6__6_ );
nand NAND2_5998 ( P3_U7807 , P3_U2583 , P3_INSTQUEUE_REG_7__6_ );
nand NAND2_5999 ( P3_U7808 , P3_U2600 , P3_INSTQUEUE_REG_8__5_ );
nand NAND2_6000 ( P3_U7809 , P3_U2599 , P3_INSTQUEUE_REG_9__5_ );
nand NAND2_6001 ( P3_U7810 , P3_U2598 , P3_INSTQUEUE_REG_10__5_ );
nand NAND2_6002 ( P3_U7811 , P3_U2597 , P3_INSTQUEUE_REG_11__5_ );
nand NAND2_6003 ( P3_U7812 , P3_U2595 , P3_INSTQUEUE_REG_12__5_ );
nand NAND2_6004 ( P3_U7813 , P3_U2594 , P3_INSTQUEUE_REG_13__5_ );
nand NAND2_6005 ( P3_U7814 , P3_U2593 , P3_INSTQUEUE_REG_14__5_ );
nand NAND2_6006 ( P3_U7815 , P3_U2592 , P3_INSTQUEUE_REG_15__5_ );
nand NAND2_6007 ( P3_U7816 , P3_U2591 , P3_INSTQUEUE_REG_0__5_ );
nand NAND2_6008 ( P3_U7817 , P3_U2590 , P3_INSTQUEUE_REG_1__5_ );
nand NAND2_6009 ( P3_U7818 , P3_U2589 , P3_INSTQUEUE_REG_2__5_ );
nand NAND2_6010 ( P3_U7819 , P3_U2588 , P3_INSTQUEUE_REG_3__5_ );
nand NAND2_6011 ( P3_U7820 , P3_U2586 , P3_INSTQUEUE_REG_4__5_ );
nand NAND2_6012 ( P3_U7821 , P3_U2585 , P3_INSTQUEUE_REG_5__5_ );
nand NAND2_6013 ( P3_U7822 , P3_U2584 , P3_INSTQUEUE_REG_6__5_ );
nand NAND2_6014 ( P3_U7823 , P3_U2583 , P3_INSTQUEUE_REG_7__5_ );
nand NAND2_6015 ( P3_U7824 , P3_U2600 , P3_INSTQUEUE_REG_8__4_ );
nand NAND2_6016 ( P3_U7825 , P3_U2599 , P3_INSTQUEUE_REG_9__4_ );
nand NAND2_6017 ( P3_U7826 , P3_U2598 , P3_INSTQUEUE_REG_10__4_ );
nand NAND2_6018 ( P3_U7827 , P3_U2597 , P3_INSTQUEUE_REG_11__4_ );
nand NAND2_6019 ( P3_U7828 , P3_U2595 , P3_INSTQUEUE_REG_12__4_ );
nand NAND2_6020 ( P3_U7829 , P3_U2594 , P3_INSTQUEUE_REG_13__4_ );
nand NAND2_6021 ( P3_U7830 , P3_U2593 , P3_INSTQUEUE_REG_14__4_ );
nand NAND2_6022 ( P3_U7831 , P3_U2592 , P3_INSTQUEUE_REG_15__4_ );
nand NAND2_6023 ( P3_U7832 , P3_U2591 , P3_INSTQUEUE_REG_0__4_ );
nand NAND2_6024 ( P3_U7833 , P3_U2590 , P3_INSTQUEUE_REG_1__4_ );
nand NAND2_6025 ( P3_U7834 , P3_U2589 , P3_INSTQUEUE_REG_2__4_ );
nand NAND2_6026 ( P3_U7835 , P3_U2588 , P3_INSTQUEUE_REG_3__4_ );
nand NAND2_6027 ( P3_U7836 , P3_U2586 , P3_INSTQUEUE_REG_4__4_ );
nand NAND2_6028 ( P3_U7837 , P3_U2585 , P3_INSTQUEUE_REG_5__4_ );
nand NAND2_6029 ( P3_U7838 , P3_U2584 , P3_INSTQUEUE_REG_6__4_ );
nand NAND2_6030 ( P3_U7839 , P3_U2583 , P3_INSTQUEUE_REG_7__4_ );
nand NAND2_6031 ( P3_U7840 , P3_U2600 , P3_INSTQUEUE_REG_8__3_ );
nand NAND2_6032 ( P3_U7841 , P3_U2599 , P3_INSTQUEUE_REG_9__3_ );
nand NAND2_6033 ( P3_U7842 , P3_U2598 , P3_INSTQUEUE_REG_10__3_ );
nand NAND2_6034 ( P3_U7843 , P3_U2597 , P3_INSTQUEUE_REG_11__3_ );
nand NAND2_6035 ( P3_U7844 , P3_U2595 , P3_INSTQUEUE_REG_12__3_ );
nand NAND2_6036 ( P3_U7845 , P3_U2594 , P3_INSTQUEUE_REG_13__3_ );
nand NAND2_6037 ( P3_U7846 , P3_U2593 , P3_INSTQUEUE_REG_14__3_ );
nand NAND2_6038 ( P3_U7847 , P3_U2592 , P3_INSTQUEUE_REG_15__3_ );
nand NAND2_6039 ( P3_U7848 , P3_U2591 , P3_INSTQUEUE_REG_0__3_ );
nand NAND2_6040 ( P3_U7849 , P3_U2590 , P3_INSTQUEUE_REG_1__3_ );
nand NAND2_6041 ( P3_U7850 , P3_U2589 , P3_INSTQUEUE_REG_2__3_ );
nand NAND2_6042 ( P3_U7851 , P3_U2588 , P3_INSTQUEUE_REG_3__3_ );
nand NAND2_6043 ( P3_U7852 , P3_U2586 , P3_INSTQUEUE_REG_4__3_ );
nand NAND2_6044 ( P3_U7853 , P3_U2585 , P3_INSTQUEUE_REG_5__3_ );
nand NAND2_6045 ( P3_U7854 , P3_U2584 , P3_INSTQUEUE_REG_6__3_ );
nand NAND2_6046 ( P3_U7855 , P3_U2583 , P3_INSTQUEUE_REG_7__3_ );
nand NAND2_6047 ( P3_U7856 , P3_U2600 , P3_INSTQUEUE_REG_8__2_ );
nand NAND2_6048 ( P3_U7857 , P3_U2599 , P3_INSTQUEUE_REG_9__2_ );
nand NAND2_6049 ( P3_U7858 , P3_U2598 , P3_INSTQUEUE_REG_10__2_ );
nand NAND2_6050 ( P3_U7859 , P3_U2597 , P3_INSTQUEUE_REG_11__2_ );
nand NAND2_6051 ( P3_U7860 , P3_U2595 , P3_INSTQUEUE_REG_12__2_ );
nand NAND2_6052 ( P3_U7861 , P3_U2594 , P3_INSTQUEUE_REG_13__2_ );
nand NAND2_6053 ( P3_U7862 , P3_U2593 , P3_INSTQUEUE_REG_14__2_ );
nand NAND2_6054 ( P3_U7863 , P3_U2592 , P3_INSTQUEUE_REG_15__2_ );
nand NAND2_6055 ( P3_U7864 , P3_U2591 , P3_INSTQUEUE_REG_0__2_ );
nand NAND2_6056 ( P3_U7865 , P3_U2590 , P3_INSTQUEUE_REG_1__2_ );
nand NAND2_6057 ( P3_U7866 , P3_U2589 , P3_INSTQUEUE_REG_2__2_ );
nand NAND2_6058 ( P3_U7867 , P3_U2588 , P3_INSTQUEUE_REG_3__2_ );
nand NAND2_6059 ( P3_U7868 , P3_U2586 , P3_INSTQUEUE_REG_4__2_ );
nand NAND2_6060 ( P3_U7869 , P3_U2585 , P3_INSTQUEUE_REG_5__2_ );
nand NAND2_6061 ( P3_U7870 , P3_U2584 , P3_INSTQUEUE_REG_6__2_ );
nand NAND2_6062 ( P3_U7871 , P3_U2583 , P3_INSTQUEUE_REG_7__2_ );
nand NAND2_6063 ( P3_U7872 , P3_U2600 , P3_INSTQUEUE_REG_8__1_ );
nand NAND2_6064 ( P3_U7873 , P3_U2599 , P3_INSTQUEUE_REG_9__1_ );
nand NAND2_6065 ( P3_U7874 , P3_U2598 , P3_INSTQUEUE_REG_10__1_ );
nand NAND2_6066 ( P3_U7875 , P3_U2597 , P3_INSTQUEUE_REG_11__1_ );
nand NAND2_6067 ( P3_U7876 , P3_U2595 , P3_INSTQUEUE_REG_12__1_ );
nand NAND2_6068 ( P3_U7877 , P3_U2594 , P3_INSTQUEUE_REG_13__1_ );
nand NAND2_6069 ( P3_U7878 , P3_U2593 , P3_INSTQUEUE_REG_14__1_ );
nand NAND2_6070 ( P3_U7879 , P3_U2592 , P3_INSTQUEUE_REG_15__1_ );
nand NAND2_6071 ( P3_U7880 , P3_U2591 , P3_INSTQUEUE_REG_0__1_ );
nand NAND2_6072 ( P3_U7881 , P3_U2590 , P3_INSTQUEUE_REG_1__1_ );
nand NAND2_6073 ( P3_U7882 , P3_U2589 , P3_INSTQUEUE_REG_2__1_ );
nand NAND2_6074 ( P3_U7883 , P3_U2588 , P3_INSTQUEUE_REG_3__1_ );
nand NAND2_6075 ( P3_U7884 , P3_U2586 , P3_INSTQUEUE_REG_4__1_ );
nand NAND2_6076 ( P3_U7885 , P3_U2585 , P3_INSTQUEUE_REG_5__1_ );
nand NAND2_6077 ( P3_U7886 , P3_U2584 , P3_INSTQUEUE_REG_6__1_ );
nand NAND2_6078 ( P3_U7887 , P3_U2583 , P3_INSTQUEUE_REG_7__1_ );
nand NAND2_6079 ( P3_U7888 , P3_U2600 , P3_INSTQUEUE_REG_8__0_ );
nand NAND2_6080 ( P3_U7889 , P3_U2599 , P3_INSTQUEUE_REG_9__0_ );
nand NAND2_6081 ( P3_U7890 , P3_U2598 , P3_INSTQUEUE_REG_10__0_ );
nand NAND2_6082 ( P3_U7891 , P3_U2597 , P3_INSTQUEUE_REG_11__0_ );
nand NAND2_6083 ( P3_U7892 , P3_U2595 , P3_INSTQUEUE_REG_12__0_ );
nand NAND2_6084 ( P3_U7893 , P3_U2594 , P3_INSTQUEUE_REG_13__0_ );
nand NAND2_6085 ( P3_U7894 , P3_U2593 , P3_INSTQUEUE_REG_14__0_ );
nand NAND2_6086 ( P3_U7895 , P3_U2592 , P3_INSTQUEUE_REG_15__0_ );
nand NAND2_6087 ( P3_U7896 , P3_U2591 , P3_INSTQUEUE_REG_0__0_ );
nand NAND2_6088 ( P3_U7897 , P3_U2590 , P3_INSTQUEUE_REG_1__0_ );
nand NAND2_6089 ( P3_U7898 , P3_U2589 , P3_INSTQUEUE_REG_2__0_ );
nand NAND2_6090 ( P3_U7899 , P3_U2588 , P3_INSTQUEUE_REG_3__0_ );
nand NAND2_6091 ( P3_U7900 , P3_U2586 , P3_INSTQUEUE_REG_4__0_ );
nand NAND2_6092 ( P3_U7901 , P3_U2585 , P3_INSTQUEUE_REG_5__0_ );
nand NAND2_6093 ( P3_U7902 , P3_U2584 , P3_INSTQUEUE_REG_6__0_ );
nand NAND2_6094 ( P3_U7903 , P3_U2583 , P3_INSTQUEUE_REG_7__0_ );
nand NAND2_6095 ( P3_U7904 , P3_STATE_REG_0_ , P3_U4292 );
or OR2_6096 ( P3_U7905 , U209 , P3_STATE2_REG_2_ );
nand NAND2_6097 ( P3_U7906 , P3_U3939 , P3_U6397 );
nand NAND2_6098 ( P3_U7907 , P3_U4134 , P3_U2603 );
nand NAND2_6099 ( P3_U7908 , P3_U2404 , P3_U3256 );
nand NAND2_6100 ( P3_U7909 , P3_U2392 , P3_U7096 );
nand NAND3_6101 ( P3_U7910 , P3_U7908 , P3_U4317 , P3_U7909 );
not NOT1_6102 ( P3_U7911 , P3_U3086 );
nand NAND2_6103 ( P3_U7912 , P3_U7911 , P3_U3088 );
nand NAND3_6104 ( P3_U7913 , P3_U4449 , P3_STATE_REG_1_ , P3_U4446 );
nand NAND2_6105 ( P3_U7914 , P3_STATE_REG_2_ , P3_U7904 );
nand NAND2_6106 ( P3_U7915 , P3_STATE_REG_1_ , P3_U4446 );
nand NAND2_6107 ( P3_U7916 , P3_U4505 , P3_U3106 );
nand NAND2_6108 ( P3_U7917 , P3_U4488 , P3_U4522 );
nand NAND2_6109 ( P3_U7918 , P3_U3208 , P3_U3219 );
nand NAND2_6110 ( P3_U7919 , P3_U7376 , P3_U3105 );
nand NAND2_6111 ( P3_U7920 , P3_BE_N_REG_3_ , P3_U3077 );
nand NAND2_6112 ( P3_U7921 , P3_BYTEENABLE_REG_3_ , P3_U4308 );
nand NAND2_6113 ( P3_U7922 , P3_BE_N_REG_2_ , P3_U3077 );
nand NAND2_6114 ( P3_U7923 , P3_BYTEENABLE_REG_2_ , P3_U4308 );
nand NAND2_6115 ( P3_U7924 , P3_BE_N_REG_1_ , P3_U3077 );
nand NAND2_6116 ( P3_U7925 , P3_BYTEENABLE_REG_1_ , P3_U4308 );
nand NAND2_6117 ( P3_U7926 , P3_BE_N_REG_0_ , P3_U3077 );
nand NAND2_6118 ( P3_U7927 , P3_BYTEENABLE_REG_0_ , P3_U4308 );
nand NAND3_6119 ( P3_U7928 , P3_STATE_REG_0_ , P3_REQUESTPENDING_REG , P3_U3079 );
nand NAND2_6120 ( P3_U7929 , P3_STATE_REG_2_ , P3_U3086 );
nand NAND2_6121 ( P3_U7930 , P3_U7929 , P3_U7928 );
nand NAND3_6122 ( P3_U7931 , P3_U7914 , P3_U4449 , P3_STATE_REG_1_ );
nand NAND2_6123 ( P3_U7932 , P3_U7930 , P3_U3076 );
nand NAND3_6124 ( P3_U7933 , P3_STATE_REG_0_ , P3_U3087 , P3_STATE_REG_2_ );
nand NAND2_6125 ( P3_U7934 , P3_U4459 , P3_U3079 );
or OR2_6126 ( P3_U7935 , P3_STATE_REG_0_ , P3_STATE_REG_1_ );
nand NAND2_6127 ( P3_U7936 , P3_STATE_REG_0_ , P3_U4346 );
not NOT1_6128 ( P3_U7937 , P3_U3278 );
nand NAND2_6129 ( P3_U7938 , P3_U7937 , P3_DATAWIDTH_REG_0_ );
nand NAND2_6130 ( P3_U7939 , P3_U3279 , P3_U3278 );
nand NAND2_6131 ( P3_U7940 , P3_U3278 , P3_U4464 );
nand NAND2_6132 ( P3_U7941 , P3_U7937 , P3_DATAWIDTH_REG_1_ );
nand NAND2_6133 ( P3_U7942 , P3_U4505 , P3_U3211 );
nand NAND2_6134 ( P3_U7943 , P3_U3104 , P3_U3214 );
nand NAND2_6135 ( P3_U7944 , P3_U4505 , P3_U3213 );
nand NAND2_6136 ( P3_U7945 , P3_U3104 , P3_U3210 );
nand NAND2_6137 ( P3_U7946 , P3_U4539 , P3_U4618 );
nand NAND2_6138 ( P3_U7947 , P3_U4620 , P3_U3101 );
nand NAND2_6139 ( P3_U7948 , P3_U4281 , P3_U4617 );
nand NAND2_6140 ( P3_U7949 , P3_U4622 , P3_U4624 );
nand NAND2_6141 ( P3_U7950 , P3_U4505 , P3_U3237 );
nand NAND2_6142 ( P3_U7951 , P3_U3104 , P3_U3238 );
nand NAND2_6143 ( P3_U7952 , P3_STATE2_REG_0_ , P3_U4627 );
nand NAND2_6144 ( P3_U7953 , P3_U4628 , P3_U3121 );
nand NAND2_6145 ( P3_U7954 , P3_STATE2_REG_3_ , P3_U3122 );
nand NAND2_6146 ( P3_U7955 , P3_U2453 , P3_U4630 );
or OR2_6147 ( P3_U7956 , P3_STATEBS16_REG , P3_STATE2_REG_0_ );
nand NAND2_6148 ( P3_U7957 , P3_STATE2_REG_0_ , P3_U7905 );
nand NAND2_6149 ( P3_U7958 , P3_STATE2_REG_0_ , P3_U4638 );
nand NAND3_6150 ( P3_U7959 , P3_U4637 , P3_U4629 , P3_U3121 );
nand NAND2_6151 ( P3_U7960 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_U3130 );
nand NAND2_6152 ( P3_U7961 , P3_U4648 , P3_U3131 );
not NOT1_6153 ( P3_U7962 , P3_U3269 );
nand NAND2_6154 ( P3_U7963 , P3_U7962 , P3_U4653 );
nand NAND2_6155 ( P3_U7964 , P3_U3269 , P3_U3138 );
not NOT1_6156 ( P3_U7965 , P3_U3270 );
nand NAND2_6157 ( P3_U7966 , P3_U7965 , P3_U4657 );
nand NAND2_6158 ( P3_U7967 , P3_U3270 , P3_U3140 );
not NOT1_6159 ( P3_U7968 , P3_U3271 );
nand NAND2_6160 ( P3_U7969 , P3_U3109 , P3_U3101 );
nand NAND2_6161 ( P3_U7970 , P3_U4539 , P3_U5483 );
nand NAND2_6162 ( P3_U7971 , P3_U3283 , P3_U4283 );
nand NAND2_6163 ( P3_U7972 , P3_U5499 , P3_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_6164 ( P3_U7973 , P3_U3218 , P3_U3107 );
nand NAND2_6165 ( P3_U7974 , P3_U4573 , P3_U4590 );
nand NAND2_6166 ( P3_U7975 , P3_U4539 , P3_U5512 );
nand NAND2_6167 ( P3_U7976 , P3_U5515 , P3_U3101 );
nand NAND3_6168 ( P3_U7977 , P3_U4556 , P3_U5517 , P3_U3110 );
nand NAND3_6169 ( P3_U7978 , P3_U5513 , P3_U3107 , P3_U4590 );
nand NAND2_6170 ( P3_U7979 , P3_U5499 , P3_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_6171 ( P3_U7980 , P3_U5546 , P3_U4283 );
nand NAND3_6172 ( P3_U7981 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_U3221 , P3_U3094 );
nand NAND3_6173 ( P3_U7982 , P3_U5531 , P3_U3097 , P3_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_6174 ( P3_U7983 , P3_INSTADDRPOINTER_REG_1_ , P3_U4284 );
nand NAND2_6175 ( P3_U7984 , P3_SUB_580_U6 , P3_INSTADDRPOINTER_REG_31_ );
not NOT1_6176 ( P3_U7985 , P3_U3287 );
nand NAND2_6177 ( P3_U7986 , P3_INSTADDRPOINTER_REG_0_ , P3_U4284 );
nand NAND2_6178 ( P3_U7987 , P3_INSTADDRPOINTER_REG_0_ , P3_INSTADDRPOINTER_REG_31_ );
not NOT1_6179 ( P3_U7988 , P3_U3286 );
nand NAND2_6180 ( P3_U7989 , P3_U5499 , P3_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_6181 ( P3_U7990 , P3_U5557 , P3_U4283 );
nand NAND2_6182 ( P3_U7991 , P3_U5499 , P3_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_6183 ( P3_U7992 , P3_U5570 , P3_U4283 );
nand NAND2_6184 ( P3_U7993 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_U3221 );
nand NAND2_6185 ( P3_U7994 , P3_U5571 , P3_U3093 );
nand NAND2_6186 ( P3_U7995 , P3_U5499 , P3_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_6187 ( P3_U7996 , P3_U5577 , P3_U4283 );
nand NAND2_6188 ( P3_U7997 , P3_U7968 , P3_U4647 );
nand NAND2_6189 ( P3_U7998 , P3_U3271 , P3_U3143 );
nand NAND2_6190 ( P3_U7999 , P3_U7998 , P3_U7997 );
nand NAND2_6191 ( P3_U8000 , P3_U5622 , P3_U3104 );
nand NAND2_6192 ( P3_U8001 , P3_U4505 , P3_U5619 );
nand NAND2_6193 ( P3_U8002 , P3_BYTEENABLE_REG_3_ , P3_U3261 );
nand NAND2_6194 ( P3_U8003 , P3_U3291 , P3_U4307 );
or OR2_6195 ( P3_U8004 , P3_DATAWIDTH_REG_0_ , P3_DATAWIDTH_REG_1_ );
nand NAND2_6196 ( P3_U8005 , P3_DATAWIDTH_REG_0_ , P3_U3240 );
nand NAND2_6197 ( P3_U8006 , P3_U8005 , P3_U8004 );
nand NAND2_6198 ( P3_U8007 , P3_U8006 , P3_U3081 );
nand NAND2_6199 ( P3_U8008 , P3_REIP_REG_0_ , P3_REIP_REG_1_ );
nand NAND2_6200 ( P3_U8009 , P3_U8008 , P3_U8007 );
nand NAND2_6201 ( P3_U8010 , P3_BYTEENABLE_REG_2_ , P3_U3261 );
nand NAND2_6202 ( P3_U8011 , P3_U8009 , P3_U4307 );
nand NAND2_6203 ( P3_U8012 , P3_BYTEENABLE_REG_1_ , P3_U3261 );
nand NAND2_6204 ( P3_U8013 , P3_U4307 , P3_REIP_REG_1_ );
nand NAND2_6205 ( P3_U8014 , P3_BYTEENABLE_REG_0_ , P3_U3261 );
nand NAND2_6206 ( P3_U8015 , P3_U4307 , P3_U7367 );
nand NAND2_6207 ( P3_U8016 , P3_U4308 , P3_U3264 );
nand NAND2_6208 ( P3_U8017 , P3_W_R_N_REG , P3_U3077 );
nand NAND2_6209 ( P3_U8018 , P3_U7368 , P3_U4617 );
nand NAND2_6210 ( P3_U8019 , P3_MORE_REG , P3_U4285 );
nand NAND2_6211 ( P3_U8020 , P3_U7937 , P3_STATEBS16_REG );
nand NAND2_6212 ( P3_U8021 , BS16 , P3_U3278 );
nand NAND2_6213 ( P3_U8022 , P3_U7374 , P3_REQUESTPENDING_REG );
nand NAND2_6214 ( P3_U8023 , P3_U7379 , P3_U4287 );
nand NAND2_6215 ( P3_U8024 , P3_U4308 , P3_U3263 );
nand NAND2_6216 ( P3_U8025 , P3_D_C_N_REG , P3_U3077 );
nand NAND2_6217 ( P3_U8026 , P3_M_IO_N_REG , P3_U3077 );
nand NAND2_6218 ( P3_U8027 , P3_MEMORYFETCH_REG , P3_U4308 );
nand NAND2_6219 ( P3_U8028 , P3_U7384 , P3_READREQUEST_REG );
nand NAND2_6220 ( P3_U8029 , P3_U7385 , P3_U4288 );
nand NAND2_6221 ( P3_U8030 , P3_U7384 , P3_MEMORYFETCH_REG );
nand NAND2_6222 ( P3_U8031 , P3_U7386 , P3_U4288 );
nand NAND2_6223 ( P3_U8032 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_U3097 );
nand NAND2_6224 ( P3_U8033 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_U3094 );
not NOT1_6225 ( P3_U8034 , P3_U3272 );
nand NAND2_6226 ( P3_U8035 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_U4289 );
nand NAND2_6227 ( P3_U8036 , P3_U7645 , P3_U3100 );
not NOT1_6228 ( P3_U8037 , P3_U3273 );
nand NAND2_6229 ( P3_U8038 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_U3207 );
nand NAND3_6230 ( P3_U8039 , P3_U3287 , P3_U3286 , P3_FLUSH_REG );
nand NAND2_6231 ( P3_U8040 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_U3207 );
nand NAND3_6232 ( P3_U8041 , P3_U3286 , P3_U7985 , P3_FLUSH_REG );
nand NAND2_6233 ( P3_U8042 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_U3207 );
nand NAND2_6234 ( P3_U8043 , P3_U7988 , P3_FLUSH_REG );
nand NAND2_6235 ( P3_U8044 , P3_U3303 , P3_U4290 );
nand NAND2_6236 ( P3_U8045 , P3_U5496 , P3_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_6237 ( P3_U8046 , P3_U5496 , P3_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_6238 ( P3_U8047 , P3_U5542 , P3_U4290 );
nand NAND2_6239 ( P3_U8048 , P3_U5496 , P3_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_6240 ( P3_U8049 , P3_U5553 , P3_U4290 );
nand NAND2_6241 ( P3_U8050 , P3_U5496 , P3_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_6242 ( P3_U8051 , P3_U5566 , P3_U4290 );
nand NAND2_6243 ( P3_U8052 , P3_U5496 , P3_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_6244 ( P3_U8053 , P3_U5573 , P3_U4290 );
nand NAND2_6245 ( P1_ADD_515_U170 , P1_ADD_515_U94 , P1_ADD_515_U7 );
nand NAND2_6246 ( P1_ADD_515_U169 , P1_INSTADDRPOINTER_REG_3_ , P1_ADD_515_U6 );
nand NAND2_6247 ( P1_ADD_515_U168 , P1_ADD_515_U122 , P1_ADD_515_U92 );
nand NAND2_6248 ( P1_ADD_515_U167 , P1_INSTADDRPOINTER_REG_31_ , P1_ADD_515_U93 );
nand NAND2_6249 ( P1_ADD_515_U166 , P1_ADD_515_U101 , P1_ADD_515_U21 );
nand NAND2_6250 ( P1_ADD_515_U165 , P1_INSTADDRPOINTER_REG_10_ , P1_ADD_515_U20 );
nand NAND2_6251 ( P1_ADD_515_U164 , P1_ADD_515_U110 , P1_ADD_515_U39 );
nand NAND2_6252 ( P1_ADD_515_U163 , P1_INSTADDRPOINTER_REG_19_ , P1_ADD_515_U38 );
nand NAND2_6253 ( P1_ADD_515_U162 , P1_ADD_515_U114 , P1_ADD_515_U47 );
nand NAND2_6254 ( P1_ADD_515_U161 , P1_INSTADDRPOINTER_REG_23_ , P1_ADD_515_U46 );
nand NAND2_6255 ( P1_ADD_515_U160 , P1_ADD_515_U99 , P1_ADD_515_U17 );
nand NAND2_6256 ( P1_ADD_515_U159 , P1_INSTADDRPOINTER_REG_8_ , P1_ADD_515_U16 );
nand NAND2_6257 ( P1_ADD_515_U158 , P1_ADD_515_U96 , P1_ADD_515_U11 );
nand NAND2_6258 ( P1_ADD_515_U157 , P1_INSTADDRPOINTER_REG_5_ , P1_ADD_515_U10 );
nand NAND2_6259 ( P1_ADD_515_U156 , P1_ADD_515_U105 , P1_ADD_515_U29 );
nand NAND2_6260 ( P1_ADD_515_U155 , P1_INSTADDRPOINTER_REG_14_ , P1_ADD_515_U28 );
nand NAND2_6261 ( P1_ADD_515_U154 , P1_ADD_515_U118 , P1_ADD_515_U55 );
nand NAND2_6262 ( P1_ADD_515_U153 , P1_INSTADDRPOINTER_REG_27_ , P1_ADD_515_U54 );
nand NAND2_6263 ( P1_ADD_515_U152 , P1_ADD_515_U95 , P1_ADD_515_U9 );
nand NAND2_6264 ( P1_ADD_515_U151 , P1_INSTADDRPOINTER_REG_4_ , P1_ADD_515_U8 );
nand NAND2_6265 ( P1_ADD_515_U150 , P1_ADD_515_U106 , P1_ADD_515_U31 );
nand NAND2_6266 ( P1_ADD_515_U149 , P1_INSTADDRPOINTER_REG_15_ , P1_ADD_515_U30 );
nand NAND2_6267 ( P1_ADD_515_U148 , P1_ADD_515_U117 , P1_ADD_515_U53 );
nand NAND2_6268 ( P1_ADD_515_U147 , P1_INSTADDRPOINTER_REG_26_ , P1_ADD_515_U52 );
nand NAND2_6269 ( P1_ADD_515_U146 , P1_ADD_515_U102 , P1_ADD_515_U23 );
nand NAND2_6270 ( P1_ADD_515_U145 , P1_INSTADDRPOINTER_REG_11_ , P1_ADD_515_U22 );
nand NAND2_6271 ( P1_ADD_515_U144 , P1_ADD_515_U109 , P1_ADD_515_U37 );
nand NAND2_6272 ( P1_ADD_515_U143 , P1_INSTADDRPOINTER_REG_18_ , P1_ADD_515_U36 );
nand NAND2_6273 ( P1_ADD_515_U142 , P1_ADD_515_U113 , P1_ADD_515_U45 );
nand NAND2_6274 ( P1_ADD_515_U141 , P1_INSTADDRPOINTER_REG_22_ , P1_ADD_515_U44 );
nand NAND2_6275 ( P1_ADD_515_U140 , P1_ADD_515_U100 , P1_ADD_515_U19 );
nand NAND2_6276 ( P1_ADD_515_U139 , P1_INSTADDRPOINTER_REG_9_ , P1_ADD_515_U18 );
nand NAND2_6277 ( P1_ADD_515_U138 , P1_ADD_515_U104 , P1_ADD_515_U27 );
nand NAND2_6278 ( P1_ADD_515_U137 , P1_INSTADDRPOINTER_REG_13_ , P1_ADD_515_U26 );
nand NAND2_6279 ( P1_ADD_515_U136 , P1_ADD_515_U111 , P1_ADD_515_U41 );
nand NAND2_6280 ( P1_ADD_515_U135 , P1_INSTADDRPOINTER_REG_20_ , P1_ADD_515_U40 );
nand NAND2_6281 ( P1_ADD_515_U134 , P1_INSTADDRPOINTER_REG_1_ , P1_ADD_515_U5 );
nand NAND2_6282 ( P1_ADD_515_U133 , P1_INSTADDRPOINTER_REG_2_ , P1_ADD_515_U4 );
nand NAND2_6283 ( P1_ADD_515_U132 , P1_ADD_515_U108 , P1_ADD_515_U35 );
nand NAND2_6284 ( P1_ADD_515_U131 , P1_INSTADDRPOINTER_REG_17_ , P1_ADD_515_U34 );
nand NAND2_6285 ( P1_ADD_515_U130 , P1_ADD_515_U115 , P1_ADD_515_U49 );
nand NAND2_6286 ( P1_ADD_515_U129 , P1_INSTADDRPOINTER_REG_24_ , P1_ADD_515_U48 );
nand NAND2_6287 ( P1_ADD_515_U128 , P1_ADD_515_U120 , P1_ADD_515_U59 );
nand NAND2_6288 ( P1_ADD_515_U127 , P1_INSTADDRPOINTER_REG_29_ , P1_ADD_515_U58 );
nand NAND2_6289 ( P1_ADD_515_U126 , P1_ADD_515_U121 , P1_ADD_515_U60 );
nand NAND2_6290 ( P1_ADD_515_U125 , P1_INSTADDRPOINTER_REG_30_ , P1_ADD_515_U61 );
nand NAND2_6291 ( P1_ADD_515_U124 , P1_ADD_515_U97 , P1_ADD_515_U12 );
nand NAND2_6292 ( P1_ADD_515_U123 , P1_INSTADDRPOINTER_REG_6_ , P1_ADD_515_U13 );
not NOT1_6293 ( P1_ADD_515_U122 , P1_ADD_515_U93 );
not NOT1_6294 ( P1_ADD_515_U121 , P1_ADD_515_U61 );
not NOT1_6295 ( P1_ADD_515_U120 , P1_ADD_515_U58 );
not NOT1_6296 ( P1_ADD_515_U119 , P1_ADD_515_U56 );
not NOT1_6297 ( P1_ADD_515_U118 , P1_ADD_515_U54 );
not NOT1_6298 ( P1_ADD_515_U117 , P1_ADD_515_U52 );
not NOT1_6299 ( P1_ADD_515_U116 , P1_ADD_515_U50 );
not NOT1_6300 ( P1_ADD_515_U115 , P1_ADD_515_U48 );
not NOT1_6301 ( P1_ADD_515_U114 , P1_ADD_515_U46 );
not NOT1_6302 ( P1_ADD_515_U113 , P1_ADD_515_U44 );
not NOT1_6303 ( P1_ADD_515_U112 , P1_ADD_515_U42 );
not NOT1_6304 ( P1_ADD_515_U111 , P1_ADD_515_U40 );
not NOT1_6305 ( P1_ADD_515_U110 , P1_ADD_515_U38 );
not NOT1_6306 ( P1_ADD_515_U109 , P1_ADD_515_U36 );
not NOT1_6307 ( P1_ADD_515_U108 , P1_ADD_515_U34 );
not NOT1_6308 ( P1_ADD_515_U107 , P1_ADD_515_U32 );
not NOT1_6309 ( P1_ADD_515_U106 , P1_ADD_515_U30 );
not NOT1_6310 ( P1_ADD_515_U105 , P1_ADD_515_U28 );
not NOT1_6311 ( P1_ADD_515_U104 , P1_ADD_515_U26 );
not NOT1_6312 ( P1_ADD_515_U103 , P1_ADD_515_U24 );
not NOT1_6313 ( P1_ADD_515_U102 , P1_ADD_515_U22 );
not NOT1_6314 ( P1_ADD_515_U101 , P1_ADD_515_U20 );
not NOT1_6315 ( P1_ADD_515_U100 , P1_ADD_515_U18 );
not NOT1_6316 ( P1_ADD_515_U99 , P1_ADD_515_U16 );
not NOT1_6317 ( P1_ADD_515_U98 , P1_ADD_515_U14 );
not NOT1_6318 ( P1_ADD_515_U97 , P1_ADD_515_U13 );
not NOT1_6319 ( P1_ADD_515_U96 , P1_ADD_515_U10 );
not NOT1_6320 ( P1_ADD_515_U95 , P1_ADD_515_U8 );
not NOT1_6321 ( P1_ADD_515_U94 , P1_ADD_515_U6 );
nand NAND2_6322 ( P1_ADD_515_U93 , P1_ADD_515_U121 , P1_INSTADDRPOINTER_REG_30_ );
not NOT1_6323 ( P1_ADD_515_U92 , P1_INSTADDRPOINTER_REG_31_ );
nand NAND2_6324 ( P1_ADD_515_U91 , P1_ADD_515_U182 , P1_ADD_515_U181 );
nand NAND2_6325 ( P1_ADD_515_U90 , P1_ADD_515_U180 , P1_ADD_515_U179 );
nand NAND2_6326 ( P1_ADD_515_U89 , P1_ADD_515_U178 , P1_ADD_515_U177 );
nand NAND2_6327 ( P1_ADD_515_U88 , P1_ADD_515_U176 , P1_ADD_515_U175 );
nand NAND2_6328 ( P1_ADD_515_U87 , P1_ADD_515_U174 , P1_ADD_515_U173 );
nand NAND2_6329 ( P1_ADD_515_U86 , P1_ADD_515_U172 , P1_ADD_515_U171 );
nand NAND2_6330 ( P1_ADD_515_U85 , P1_ADD_515_U170 , P1_ADD_515_U169 );
nand NAND2_6331 ( P1_ADD_515_U84 , P1_ADD_515_U168 , P1_ADD_515_U167 );
nand NAND2_6332 ( P1_ADD_515_U83 , P1_ADD_515_U166 , P1_ADD_515_U165 );
nand NAND2_6333 ( P1_ADD_515_U82 , P1_ADD_515_U164 , P1_ADD_515_U163 );
nand NAND2_6334 ( P1_ADD_515_U81 , P1_ADD_515_U162 , P1_ADD_515_U161 );
nand NAND2_6335 ( P1_ADD_515_U80 , P1_ADD_515_U160 , P1_ADD_515_U159 );
nand NAND2_6336 ( P1_ADD_515_U79 , P1_ADD_515_U158 , P1_ADD_515_U157 );
nand NAND2_6337 ( P1_ADD_515_U78 , P1_ADD_515_U156 , P1_ADD_515_U155 );
nand NAND2_6338 ( P1_ADD_515_U77 , P1_ADD_515_U154 , P1_ADD_515_U153 );
nand NAND2_6339 ( P1_ADD_515_U76 , P1_ADD_515_U152 , P1_ADD_515_U151 );
nand NAND2_6340 ( P1_ADD_515_U75 , P1_ADD_515_U150 , P1_ADD_515_U149 );
nand NAND2_6341 ( P1_ADD_515_U74 , P1_ADD_515_U148 , P1_ADD_515_U147 );
nand NAND2_6342 ( P1_ADD_515_U73 , P1_ADD_515_U146 , P1_ADD_515_U145 );
nand NAND2_6343 ( P1_ADD_515_U72 , P1_ADD_515_U144 , P1_ADD_515_U143 );
nand NAND2_6344 ( P1_ADD_515_U71 , P1_ADD_515_U142 , P1_ADD_515_U141 );
nand NAND2_6345 ( P1_ADD_515_U70 , P1_ADD_515_U140 , P1_ADD_515_U139 );
nand NAND2_6346 ( P1_ADD_515_U69 , P1_ADD_515_U138 , P1_ADD_515_U137 );
nand NAND2_6347 ( P1_ADD_515_U68 , P1_ADD_515_U136 , P1_ADD_515_U135 );
nand NAND2_6348 ( P1_ADD_515_U67 , P1_ADD_515_U134 , P1_ADD_515_U133 );
nand NAND2_6349 ( P1_ADD_515_U66 , P1_ADD_515_U132 , P1_ADD_515_U131 );
nand NAND2_6350 ( P1_ADD_515_U65 , P1_ADD_515_U130 , P1_ADD_515_U129 );
nand NAND2_6351 ( P1_ADD_515_U64 , P1_ADD_515_U128 , P1_ADD_515_U127 );
nand NAND2_6352 ( P1_ADD_515_U63 , P1_ADD_515_U126 , P1_ADD_515_U125 );
nand NAND2_6353 ( P1_ADD_515_U62 , P1_ADD_515_U124 , P1_ADD_515_U123 );
nand NAND2_6354 ( P1_ADD_515_U61 , P1_INSTADDRPOINTER_REG_29_ , P1_ADD_515_U120 );
not NOT1_6355 ( P1_ADD_515_U60 , P1_INSTADDRPOINTER_REG_30_ );
not NOT1_6356 ( P1_ADD_515_U59 , P1_INSTADDRPOINTER_REG_29_ );
nand NAND2_6357 ( P1_ADD_515_U58 , P1_INSTADDRPOINTER_REG_28_ , P1_ADD_515_U119 );
not NOT1_6358 ( P1_ADD_515_U57 , P1_INSTADDRPOINTER_REG_28_ );
nand NAND2_6359 ( P1_ADD_515_U56 , P1_INSTADDRPOINTER_REG_27_ , P1_ADD_515_U118 );
not NOT1_6360 ( P1_ADD_515_U55 , P1_INSTADDRPOINTER_REG_27_ );
nand NAND2_6361 ( P1_ADD_515_U54 , P1_INSTADDRPOINTER_REG_26_ , P1_ADD_515_U117 );
not NOT1_6362 ( P1_ADD_515_U53 , P1_INSTADDRPOINTER_REG_26_ );
nand NAND2_6363 ( P1_ADD_515_U52 , P1_INSTADDRPOINTER_REG_25_ , P1_ADD_515_U116 );
not NOT1_6364 ( P1_ADD_515_U51 , P1_INSTADDRPOINTER_REG_25_ );
nand NAND2_6365 ( P1_ADD_515_U50 , P1_INSTADDRPOINTER_REG_24_ , P1_ADD_515_U115 );
not NOT1_6366 ( P1_ADD_515_U49 , P1_INSTADDRPOINTER_REG_24_ );
nand NAND2_6367 ( P1_ADD_515_U48 , P1_INSTADDRPOINTER_REG_23_ , P1_ADD_515_U114 );
not NOT1_6368 ( P1_ADD_515_U47 , P1_INSTADDRPOINTER_REG_23_ );
nand NAND2_6369 ( P1_ADD_515_U46 , P1_INSTADDRPOINTER_REG_22_ , P1_ADD_515_U113 );
not NOT1_6370 ( P1_ADD_515_U45 , P1_INSTADDRPOINTER_REG_22_ );
nand NAND2_6371 ( P1_ADD_515_U44 , P1_INSTADDRPOINTER_REG_21_ , P1_ADD_515_U112 );
not NOT1_6372 ( P1_ADD_515_U43 , P1_INSTADDRPOINTER_REG_21_ );
nand NAND2_6373 ( P1_ADD_515_U42 , P1_INSTADDRPOINTER_REG_20_ , P1_ADD_515_U111 );
not NOT1_6374 ( P1_ADD_515_U41 , P1_INSTADDRPOINTER_REG_20_ );
nand NAND2_6375 ( P1_ADD_515_U40 , P1_INSTADDRPOINTER_REG_19_ , P1_ADD_515_U110 );
not NOT1_6376 ( P1_ADD_515_U39 , P1_INSTADDRPOINTER_REG_19_ );
nand NAND2_6377 ( P1_ADD_515_U38 , P1_INSTADDRPOINTER_REG_18_ , P1_ADD_515_U109 );
not NOT1_6378 ( P1_ADD_515_U37 , P1_INSTADDRPOINTER_REG_18_ );
nand NAND2_6379 ( P1_ADD_515_U36 , P1_INSTADDRPOINTER_REG_17_ , P1_ADD_515_U108 );
not NOT1_6380 ( P1_ADD_515_U35 , P1_INSTADDRPOINTER_REG_17_ );
nand NAND2_6381 ( P1_ADD_515_U34 , P1_INSTADDRPOINTER_REG_16_ , P1_ADD_515_U107 );
not NOT1_6382 ( P1_ADD_515_U33 , P1_INSTADDRPOINTER_REG_16_ );
nand NAND2_6383 ( P1_ADD_515_U32 , P1_INSTADDRPOINTER_REG_15_ , P1_ADD_515_U106 );
not NOT1_6384 ( P1_ADD_515_U31 , P1_INSTADDRPOINTER_REG_15_ );
nand NAND2_6385 ( P1_ADD_515_U30 , P1_INSTADDRPOINTER_REG_14_ , P1_ADD_515_U105 );
not NOT1_6386 ( P1_ADD_515_U29 , P1_INSTADDRPOINTER_REG_14_ );
nand NAND2_6387 ( P1_ADD_515_U28 , P1_INSTADDRPOINTER_REG_13_ , P1_ADD_515_U104 );
not NOT1_6388 ( P1_ADD_515_U27 , P1_INSTADDRPOINTER_REG_13_ );
nand NAND2_6389 ( P1_ADD_515_U26 , P1_INSTADDRPOINTER_REG_12_ , P1_ADD_515_U103 );
not NOT1_6390 ( P1_ADD_515_U25 , P1_INSTADDRPOINTER_REG_12_ );
nand NAND2_6391 ( P1_ADD_515_U24 , P1_INSTADDRPOINTER_REG_11_ , P1_ADD_515_U102 );
not NOT1_6392 ( P1_ADD_515_U23 , P1_INSTADDRPOINTER_REG_11_ );
nand NAND2_6393 ( P1_ADD_515_U22 , P1_INSTADDRPOINTER_REG_10_ , P1_ADD_515_U101 );
not NOT1_6394 ( P1_ADD_515_U21 , P1_INSTADDRPOINTER_REG_10_ );
nand NAND2_6395 ( P1_ADD_515_U20 , P1_INSTADDRPOINTER_REG_9_ , P1_ADD_515_U100 );
not NOT1_6396 ( P1_ADD_515_U19 , P1_INSTADDRPOINTER_REG_9_ );
nand NAND2_6397 ( P1_ADD_515_U18 , P1_INSTADDRPOINTER_REG_8_ , P1_ADD_515_U99 );
not NOT1_6398 ( P1_ADD_515_U17 , P1_INSTADDRPOINTER_REG_8_ );
nand NAND2_6399 ( P1_ADD_515_U16 , P1_INSTADDRPOINTER_REG_7_ , P1_ADD_515_U98 );
not NOT1_6400 ( P1_ADD_515_U15 , P1_INSTADDRPOINTER_REG_7_ );
nand NAND2_6401 ( P1_ADD_515_U14 , P1_ADD_515_U97 , P1_INSTADDRPOINTER_REG_6_ );
nand NAND2_6402 ( P1_ADD_515_U13 , P1_INSTADDRPOINTER_REG_5_ , P1_ADD_515_U96 );
not NOT1_6403 ( P1_ADD_515_U12 , P1_INSTADDRPOINTER_REG_6_ );
not NOT1_6404 ( P1_ADD_515_U11 , P1_INSTADDRPOINTER_REG_5_ );
nand NAND2_6405 ( P1_ADD_515_U10 , P1_INSTADDRPOINTER_REG_4_ , P1_ADD_515_U95 );
not NOT1_6406 ( P1_ADD_515_U9 , P1_INSTADDRPOINTER_REG_4_ );
nand NAND2_6407 ( P1_ADD_515_U8 , P1_INSTADDRPOINTER_REG_3_ , P1_ADD_515_U94 );
not NOT1_6408 ( P1_ADD_515_U7 , P1_INSTADDRPOINTER_REG_3_ );
nand NAND2_6409 ( P1_ADD_515_U6 , P1_INSTADDRPOINTER_REG_2_ , P1_INSTADDRPOINTER_REG_1_ );
not NOT1_6410 ( P1_ADD_515_U5 , P1_INSTADDRPOINTER_REG_2_ );
not NOT1_6411 ( P1_ADD_515_U4 , P1_INSTADDRPOINTER_REG_1_ );
nor nor_6412 ( P1_GTE_485_U7 , P1_R2238_U19 , P1_R2238_U20 , P1_R2238_U22 , P1_R2238_U21 );
nor nor_6413 ( P1_GTE_485_U6 , P1_R2238_U6 , P1_GTE_485_U7 );
nand NAND2_6414 ( P1_ADD_405_U186 , P1_ADD_405_U110 , P1_ADD_405_U33 );
nand NAND2_6415 ( P1_ADD_405_U185 , P1_INSTADDRPOINTER_REG_16_ , P1_ADD_405_U32 );
nand NAND2_6416 ( P1_ADD_405_U184 , P1_ADD_405_U119 , P1_ADD_405_U51 );
nand NAND2_6417 ( P1_ADD_405_U183 , P1_INSTADDRPOINTER_REG_25_ , P1_ADD_405_U50 );
nand NAND2_6418 ( P1_ADD_405_U182 , P1_ADD_405_U101 , P1_ADD_405_U15 );
nand NAND2_6419 ( P1_ADD_405_U181 , P1_INSTADDRPOINTER_REG_7_ , P1_ADD_405_U14 );
nand NAND2_6420 ( P1_ADD_405_U180 , P1_ADD_405_U106 , P1_ADD_405_U25 );
nand NAND2_6421 ( P1_ADD_405_U179 , P1_INSTADDRPOINTER_REG_12_ , P1_ADD_405_U24 );
nand NAND2_6422 ( P1_ADD_405_U178 , P1_ADD_405_U115 , P1_ADD_405_U43 );
nand NAND2_6423 ( P1_ADD_405_U177 , P1_INSTADDRPOINTER_REG_21_ , P1_ADD_405_U42 );
nand NAND2_6424 ( P1_ADD_405_U176 , P1_ADD_405_U122 , P1_ADD_405_U57 );
nand NAND2_6425 ( P1_ADD_405_U175 , P1_INSTADDRPOINTER_REG_28_ , P1_ADD_405_U56 );
nand NAND2_6426 ( P1_ADD_405_U174 , P1_INSTADDRPOINTER_REG_0_ , P1_ADD_405_U6 );
nand NAND2_6427 ( P1_ADD_405_U173 , P1_INSTADDRPOINTER_REG_1_ , P1_ADD_405_U4 );
and AND3_6428 ( P2_U2352 , P2_U2617 , P2_U3300 , P2_U7873 );
and AND2_6429 ( P2_U2353 , P2_U4343 , P2_U2439 );
and AND3_6430 ( P2_U2354 , P2_U7861 , P2_U7873 , P2_STATE2_REG_0_ );
and AND2_6431 ( P2_U2355 , P2_U2447 , P2_U7861 );
and AND2_6432 ( P2_U2356 , P2_STATE2_REG_0_ , P2_U3253 );
and AND2_6433 ( P2_U2357 , P2_U3712 , P2_U2458 );
and AND2_6434 ( P2_U2358 , P2_U4431 , P2_STATE2_REG_0_ );
and AND2_6435 ( P2_U2359 , P2_U4411 , P2_U3265 );
nor nor_6436 ( P2_U2360 , U211 , P2_STATEBS16_REG );
and AND2_6437 ( P2_U2361 , P2_R2238_U6 , P2_U2356 );
and AND2_6438 ( P2_U2362 , P2_U2398 , P2_U4443 );
and AND2_6439 ( P2_U2363 , P2_STATE2_REG_2_ , P2_U3535 );
and AND2_6440 ( P2_U2364 , P2_STATE2_REG_2_ , P2_U3546 );
and AND2_6441 ( P2_U2365 , P2_U4443 , P2_STATE2_REG_3_ );
and AND2_6442 ( P2_U2366 , P2_STATE2_REG_1_ , P2_U3546 );
and AND2_6443 ( P2_U2367 , P2_U2364 , P2_U4417 );
and AND2_6444 ( P2_U2368 , P2_U2363 , P2_U4420 );
and AND2_6445 ( P2_U2369 , P2_U2364 , P2_U4428 );
and AND2_6446 ( P2_U2370 , P2_U2447 , P2_U3537 );
and AND2_6447 ( P2_U2371 , P2_U3990 , P2_U3537 );
and AND2_6448 ( P2_U2372 , P2_U3989 , P2_U3537 );
and AND2_6449 ( P2_U2373 , P2_U4419 , P2_U3537 );
and AND2_6450 ( P2_U2374 , P2_U4468 , P2_STATE2_REG_0_ );
and AND2_6451 ( P2_U2375 , P2_U4441 , P2_U3521 );
and AND2_6452 ( P2_U2376 , P2_U3873 , P2_U2436 );
and AND2_6453 ( P2_U2377 , P2_U2367 , P2_U4411 );
and AND2_6454 ( P2_U2378 , P2_STATE2_REG_3_ , P2_U3546 );
and AND2_6455 ( P2_U2379 , P2_U4440 , P2_U7865 );
and AND2_6456 ( P2_U2380 , P2_U4441 , P2_U7865 );
and AND2_6457 ( P2_U2381 , P2_U3535 , P2_U3270 );
and AND2_6458 ( P2_U2382 , P2_U2366 , P2_U3647 );
and AND2_6459 ( P2_U2383 , P2_U2366 , P2_U3528 );
and AND2_6460 ( P2_U2384 , P2_U2368 , P2_U4417 );
and AND2_6461 ( P2_U2385 , P2_U2368 , P2_U4428 );
and AND2_6462 ( P2_U2386 , P2_U2363 , P2_U4436 );
and AND2_6463 ( P2_U2387 , P2_U5940 , P2_U3537 );
and AND2_6464 ( P2_U2388 , P2_U2363 , P2_U5675 );
and AND2_6465 ( P2_U2389 , P2_U2363 , P2_U5677 );
and AND2_6466 ( P2_U2390 , P2_U2363 , P2_U5679 );
and AND2_6467 ( P2_U2391 , P2_U2369 , P2_U3545 );
and AND2_6468 ( P2_U2392 , P2_U6571 , P2_U2369 );
and AND2_6469 ( P2_U2393 , P2_U4440 , P2_U3521 );
and AND2_6470 ( P2_U2394 , P2_U4442 , P2_U2616 );
and AND2_6471 ( P2_U2395 , P2_U4442 , P2_U7873 );
and AND2_6472 ( P2_U2396 , P2_U3541 , P2_U3284 );
and AND2_6473 ( P2_U2397 , P2_U4441 , P2_U4601 );
and AND2_6474 ( P2_U2398 , P2_U4430 , P2_STATEBS16_REG );
and AND2_6475 ( P2_U2399 , U314 , P2_U4443 );
and AND2_6476 ( P2_U2400 , U303 , P2_U4443 );
and AND2_6477 ( P2_U2401 , U292 , P2_U4443 );
and AND2_6478 ( P2_U2402 , U289 , P2_U4443 );
and AND2_6479 ( P2_U2403 , U288 , P2_U4443 );
and AND2_6480 ( P2_U2404 , U287 , P2_U4443 );
and AND2_6481 ( P2_U2405 , U286 , P2_U4443 );
and AND2_6482 ( P2_U2406 , U285 , P2_U4443 );
and AND2_6483 ( P2_U2407 , U298 , P2_U2362 );
and AND2_6484 ( P2_U2408 , U307 , P2_U2362 );
and AND2_6485 ( P2_U2409 , U297 , P2_U2362 );
and AND2_6486 ( P2_U2410 , U306 , P2_U2362 );
and AND2_6487 ( P2_U2411 , U296 , P2_U2362 );
and AND2_6488 ( P2_U2412 , U305 , P2_U2362 );
and AND2_6489 ( P2_U2413 , U295 , P2_U2362 );
and AND2_6490 ( P2_U2414 , U304 , P2_U2362 );
and AND2_6491 ( P2_U2415 , U294 , P2_U2362 );
and AND2_6492 ( P2_U2416 , U302 , P2_U2362 );
and AND2_6493 ( P2_U2417 , U293 , P2_U2362 );
and AND2_6494 ( P2_U2418 , U301 , P2_U2362 );
and AND2_6495 ( P2_U2419 , U291 , P2_U2362 );
and AND2_6496 ( P2_U2420 , U300 , P2_U2362 );
and AND2_6497 ( P2_U2421 , U290 , P2_U2362 );
and AND2_6498 ( P2_U2422 , U299 , P2_U2362 );
and AND2_6499 ( P2_U2423 , P2_U2365 , P2_U3255 );
and AND2_6500 ( P2_U2424 , P2_U2365 , P2_U3278 );
and AND2_6501 ( P2_U2425 , P2_U2365 , P2_U3521 );
and AND2_6502 ( P2_U2426 , P2_U2365 , P2_U3279 );
and AND2_6503 ( P2_U2427 , P2_U2375 , P2_U3279 );
and AND2_6504 ( P2_U2428 , P2_U2365 , P2_U2616 );
and AND2_6505 ( P2_U2429 , P2_U2365 , P2_U2617 );
and AND2_6506 ( P2_U2430 , P2_STATE2_REG_0_ , P2_U3541 );
and AND2_6507 ( P2_U2431 , P2_U2365 , P2_U3253 );
and AND2_6508 ( P2_U2432 , P2_U2365 , P2_U3280 );
and AND2_6509 ( P2_U2433 , P2_U2375 , P2_U3295 );
and AND2_6510 ( P2_U2434 , P2_U2375 , P2_U7869 );
and AND2_6511 ( P2_U2435 , P2_U2356 , P2_U3541 );
and AND2_6512 ( P2_U2436 , P2_U7859 , P2_U7867 );
and AND2_6513 ( P2_U2437 , P2_U2364 , P2_U7871 );
and AND2_6514 ( P2_U2438 , P2_U7859 , P2_U3278 );
and AND2_6515 ( P2_U2439 , P2_U4339 , P2_U3521 );
and AND2_6516 ( P2_U2440 , P2_U3580 , P2_U3428 );
and AND2_6517 ( P2_U2441 , P2_U4647 , P2_U3580 );
and AND2_6518 ( P2_U2442 , P2_U8067 , P2_U3428 );
and AND2_6519 ( P2_U2443 , P2_U4647 , P2_U8067 );
and AND2_6520 ( P2_U2444 , P2_U3243 , P2_U3307 );
and AND2_6521 ( P2_U2445 , P2_U4650 , P2_U3307 );
and AND2_6522 ( P2_U2446 , P2_R2088_U6 , P2_U4424 );
and AND2_6523 ( P2_U2447 , P2_STATE2_REG_0_ , P2_U2616 );
and AND2_6524 ( P2_U2448 , P2_STATE2_REG_2_ , P2_STATE2_REG_1_ );
and AND2_6525 ( P2_U2449 , P2_U3278 , P2_U3521 );
and AND2_6526 ( P2_U2450 , P2_U2354 , P2_U7871 );
and AND3_6527 ( P2_U2451 , P2_U4601 , P2_U2457 , P2_U2438 );
and AND3_6528 ( P2_U2452 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_U3272 , P2_INSTQUEUERD_ADDR_REG_2_ );
and AND3_6529 ( P2_U2453 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_U3271 , P2_INSTQUEUERD_ADDR_REG_2_ );
and AND3_6530 ( P2_U2454 , P2_U3271 , P2_U3272 , P2_INSTQUEUERD_ADDR_REG_2_ );
and AND3_6531 ( P2_U2455 , P2_U3276 , P2_U3272 , P2_INSTQUEUERD_ADDR_REG_1_ );
and AND3_6532 ( P2_U2456 , P2_U3276 , P2_U3271 , P2_INSTQUEUERD_ADDR_REG_0_ );
and AND2_6533 ( P2_U2457 , P2_U3521 , P2_U3255 );
and AND3_6534 ( P2_U2458 , P2_U2617 , P2_U3279 , P2_U7863 );
and AND3_6535 ( P2_U2459 , P2_U8053 , P2_U8052 , P2_U4393 );
and AND2_6536 ( P2_U2460 , P2_R2182_U40 , P2_U3317 );
and AND2_6537 ( P2_U2461 , P2_U3579 , P2_U3426 );
and AND2_6538 ( P2_U2462 , P2_R2182_U76 , P2_R2182_U40 );
and AND2_6539 ( P2_U2463 , P2_U4637 , P2_U2462 );
and AND2_6540 ( P2_U2464 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_INSTQUEUEWR_ADDR_REG_3_ );
and AND2_6541 ( P2_U2465 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_U3309 );
and AND2_6542 ( P2_U2466 , P2_R2099_U96 , P2_R2099_U95 );
and AND2_6543 ( P2_U2467 , P2_R2099_U5 , P2_R2099_U94 );
and AND2_6544 ( P2_U2468 , P2_U3320 , P2_U4657 );
and AND2_6545 ( P2_U2469 , P2_U4633 , P2_U2462 );
and AND2_6546 ( P2_U2470 , P2_R2099_U5 , P2_U3323 );
and AND2_6547 ( P2_U2471 , P2_U3339 , P2_U4715 );
and AND2_6548 ( P2_U2472 , P2_U4634 , P2_U2462 );
and AND2_6549 ( P2_U2473 , P2_R2099_U94 , P2_U3324 );
and AND2_6550 ( P2_U2474 , P2_U3354 , P2_U4774 );
and AND2_6551 ( P2_U2475 , P2_U4635 , P2_R2182_U69 );
nor nor_6552 ( P2_U2476 , P2_R2182_U69 , P2_R2182_U68 );
and AND2_6553 ( P2_U2477 , P2_U2476 , P2_U2462 );
nor nor_6554 ( P2_U2478 , P2_INSTQUEUEWR_ADDR_REG_0_ , P2_INSTQUEUEWR_ADDR_REG_1_ );
nor nor_6555 ( P2_U2479 , P2_R2099_U94 , P2_R2099_U5 );
and AND2_6556 ( P2_U2480 , P2_U3366 , P2_U4831 );
and AND2_6557 ( P2_U2481 , P2_U8064 , P2_U3426 );
and AND2_6558 ( P2_U2482 , P2_U4638 , P2_U4637 );
and AND2_6559 ( P2_U2483 , P2_R2099_U95 , P2_U3322 );
and AND2_6560 ( P2_U2484 , P2_U3379 , P2_U4889 );
and AND2_6561 ( P2_U2485 , P2_U4638 , P2_U4633 );
and AND2_6562 ( P2_U2486 , P2_U3391 , P2_U4946 );
and AND2_6563 ( P2_U2487 , P2_U4638 , P2_U4634 );
and AND2_6564 ( P2_U2488 , P2_U3402 , P2_U5004 );
and AND2_6565 ( P2_U2489 , P2_U4638 , P2_U2476 );
and AND2_6566 ( P2_U2490 , P2_U3414 , P2_U5061 );
and AND2_6567 ( P2_U2491 , P2_U4640 , P2_U3579 );
and AND2_6568 ( P2_U2492 , P2_R2099_U96 , P2_U3321 );
and AND2_6569 ( P2_U2493 , P2_U3427 , P2_U3425 );
and AND2_6570 ( P2_U2494 , P2_U4633 , P2_U2460 );
and AND2_6571 ( P2_U2495 , P2_U3440 , P2_U5174 );
and AND2_6572 ( P2_U2496 , P2_U4634 , P2_U2460 );
and AND2_6573 ( P2_U2497 , P2_U3451 , P2_U5232 );
and AND2_6574 ( P2_U2498 , P2_U2476 , P2_U2460 );
and AND2_6575 ( P2_U2499 , P2_U3463 , P2_U5289 );
and AND2_6576 ( P2_U2500 , P2_U4640 , P2_U8064 );
nor nor_6577 ( P2_U2501 , P2_R2182_U40 , P2_R2182_U76 );
and AND2_6578 ( P2_U2502 , P2_U2501 , P2_U4637 );
nor nor_6579 ( P2_U2503 , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_INSTQUEUEWR_ADDR_REG_2_ );
nor nor_6580 ( P2_U2504 , P2_R2099_U95 , P2_R2099_U96 );
and AND2_6581 ( P2_U2505 , P2_U3474 , P2_U5347 );
and AND2_6582 ( P2_U2506 , P2_U2501 , P2_U4633 );
and AND2_6583 ( P2_U2507 , P2_U3486 , P2_U5404 );
and AND2_6584 ( P2_U2508 , P2_U2501 , P2_U4634 );
and AND2_6585 ( P2_U2509 , P2_U3497 , P2_U5462 );
and AND2_6586 ( P2_U2510 , P2_U2501 , P2_U2476 );
and AND2_6587 ( P2_U2511 , P2_U3509 , P2_U5519 );
and AND3_6588 ( P2_U2512 , P2_U8069 , P2_U8068 , P2_U3869 );
and AND2_6589 ( P2_U2513 , P2_U5580 , P2_U5579 );
and AND3_6590 ( P2_U2514 , P2_U3881 , P2_U7896 , P2_U3882 );
and AND2_6591 ( P2_U2515 , P2_U8082 , P2_U8100 );
and AND2_6592 ( P2_U2516 , P2_U5616 , P2_INSTQUEUERD_ADDR_REG_0_ );
and AND2_6593 ( P2_U2517 , P2_U2515 , P2_U2516 );
and AND2_6594 ( P2_U2518 , P2_U5616 , P2_U3272 );
and AND2_6595 ( P2_U2519 , P2_U2515 , P2_U2518 );
and AND2_6596 ( P2_U2520 , P2_U8082 , P2_U3582 );
and AND2_6597 ( P2_U2521 , P2_U2520 , P2_U2516 );
and AND2_6598 ( P2_U2522 , P2_U2520 , P2_U2518 );
and AND2_6599 ( P2_U2523 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_U3530 );
and AND2_6600 ( P2_U2524 , P2_U2515 , P2_U2523 );
and AND2_6601 ( P2_U2525 , P2_U3272 , P2_U3530 );
and AND2_6602 ( P2_U2526 , P2_U2515 , P2_U2525 );
and AND2_6603 ( P2_U2527 , P2_U2520 , P2_U2523 );
and AND2_6604 ( P2_U2528 , P2_U2520 , P2_U2525 );
and AND2_6605 ( P2_U2529 , P2_U3582 , P2_U3581 );
and AND2_6606 ( P2_U2530 , P2_U2525 , P2_U2529 );
and AND2_6607 ( P2_U2531 , P2_U2523 , P2_U2529 );
and AND2_6608 ( P2_U2532 , P2_U8100 , P2_U3581 );
and AND2_6609 ( P2_U2533 , P2_U2525 , P2_U2532 );
and AND2_6610 ( P2_U2534 , P2_U2523 , P2_U2532 );
and AND2_6611 ( P2_U2535 , P2_U2529 , P2_U2518 );
and AND2_6612 ( P2_U2536 , P2_U2529 , P2_U2516 );
and AND2_6613 ( P2_U2537 , P2_U2518 , P2_U2532 );
and AND2_6614 ( P2_U2538 , P2_U2516 , P2_U2532 );
nor nor_6615 ( P2_U2539 , P2_R2147_U8 , P2_R2147_U4 );
nor nor_6616 ( P2_U2540 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_R2147_U9 );
and AND2_6617 ( P2_U2541 , P2_U2539 , P2_U2540 );
and AND2_6618 ( P2_U2542 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_U3529 );
and AND2_6619 ( P2_U2543 , P2_U2539 , P2_U2542 );
and AND2_6620 ( P2_U2544 , P2_R2147_U4 , P2_U3526 );
and AND2_6621 ( P2_U2545 , P2_U2544 , P2_U2540 );
and AND2_6622 ( P2_U2546 , P2_U2544 , P2_U2542 );
and AND2_6623 ( P2_U2547 , P2_R2147_U9 , P2_U3532 );
and AND2_6624 ( P2_U2548 , P2_U2539 , P2_U2547 );
and AND2_6625 ( P2_U2549 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_R2147_U9 );
and AND2_6626 ( P2_U2550 , P2_U2539 , P2_U2549 );
and AND2_6627 ( P2_U2551 , P2_U2544 , P2_U2547 );
and AND2_6628 ( P2_U2552 , P2_U2544 , P2_U2549 );
and AND2_6629 ( P2_U2553 , P2_R2147_U8 , P2_U3531 );
and AND2_6630 ( P2_U2554 , P2_U2540 , P2_U2553 );
and AND2_6631 ( P2_U2555 , P2_U2542 , P2_U2553 );
and AND2_6632 ( P2_U2556 , P2_R2147_U4 , P2_R2147_U8 );
and AND2_6633 ( P2_U2557 , P2_U2540 , P2_U2556 );
and AND2_6634 ( P2_U2558 , P2_U2542 , P2_U2556 );
and AND2_6635 ( P2_U2559 , P2_U2553 , P2_U2547 );
and AND2_6636 ( P2_U2560 , P2_U2553 , P2_U2549 );
and AND2_6637 ( P2_U2561 , P2_U2547 , P2_U2556 );
and AND2_6638 ( P2_U2562 , P2_U2549 , P2_U2556 );
and AND2_6639 ( P2_U2563 , P2_U8100 , P2_U3272 );
and AND2_6640 ( P2_U2564 , P2_U4409 , P2_U3583 );
and AND2_6641 ( P2_U2565 , P2_U2564 , P2_U2563 );
and AND2_6642 ( P2_U2566 , P2_U8100 , P2_INSTQUEUERD_ADDR_REG_0_ );
and AND2_6643 ( P2_U2567 , P2_U2564 , P2_U2566 );
and AND2_6644 ( P2_U2568 , P2_U3582 , P2_U3272 );
and AND2_6645 ( P2_U2569 , P2_U2564 , P2_U2568 );
and AND2_6646 ( P2_U2570 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_U3582 );
and AND2_6647 ( P2_U2571 , P2_U2564 , P2_U2570 );
and AND2_6648 ( P2_U2572 , P2_U3583 , P2_U3553 );
and AND2_6649 ( P2_U2573 , P2_U2572 , P2_U2563 );
and AND2_6650 ( P2_U2574 , P2_U2572 , P2_U2566 );
and AND2_6651 ( P2_U2575 , P2_U2572 , P2_U2568 );
and AND2_6652 ( P2_U2576 , P2_U2572 , P2_U2570 );
and AND2_6653 ( P2_U2577 , P2_U4409 , P2_U8149 );
and AND2_6654 ( P2_U2578 , P2_U2577 , P2_U2563 );
and AND2_6655 ( P2_U2579 , P2_U2577 , P2_U2566 );
and AND2_6656 ( P2_U2580 , P2_U2577 , P2_U2568 );
and AND2_6657 ( P2_U2581 , P2_U2577 , P2_U2570 );
and AND2_6658 ( P2_U2582 , P2_U8149 , P2_U3553 );
and AND2_6659 ( P2_U2583 , P2_U2563 , P2_U2582 );
and AND2_6660 ( P2_U2584 , P2_U2566 , P2_U2582 );
and AND2_6661 ( P2_U2585 , P2_U2568 , P2_U2582 );
and AND2_6662 ( P2_U2586 , P2_U2570 , P2_U2582 );
and AND2_6663 ( P2_U2587 , P2_EBX_REG_31_ , P2_U2391 );
and AND2_6664 ( P2_U2588 , P2_U2377 , P2_U2360 );
and AND4_6665 ( P2_U2589 , P2_U7581 , P2_U3550 , P2_U4457 , P2_U3549 );
and AND2_6666 ( P2_U2590 , P2_U5590 , P2_U2436 );
nand NAND2_6667 ( P2_U2591 , P2_U4274 , P2_U4273 );
nand NAND2_6668 ( P2_U2592 , P2_U4272 , P2_U4271 );
nand NAND2_6669 ( P2_U2593 , P2_U4270 , P2_U4269 );
nand NAND2_6670 ( P2_U2594 , P2_U4268 , P2_U4267 );
nand NAND2_6671 ( P2_U2595 , P2_U4266 , P2_U4265 );
nand NAND2_6672 ( P2_U2596 , P2_U4264 , P2_U4263 );
nand NAND2_6673 ( P2_U2597 , P2_U4262 , P2_U4261 );
nand NAND2_6674 ( P2_U2598 , P2_U4260 , P2_U4259 );
nand NAND4_6675 ( P2_U2599 , P2_U4258 , P2_U4257 , P2_U4256 , P2_U4255 );
nand NAND4_6676 ( P2_U2600 , P2_U4254 , P2_U4253 , P2_U4252 , P2_U4251 );
nand NAND4_6677 ( P2_U2601 , P2_U4250 , P2_U4249 , P2_U4248 , P2_U4247 );
nand NAND4_6678 ( P2_U2602 , P2_U4246 , P2_U4245 , P2_U4244 , P2_U4243 );
nand NAND4_6679 ( P2_U2603 , P2_U4242 , P2_U4241 , P2_U4240 , P2_U4239 );
nand NAND4_6680 ( P2_U2604 , P2_U4238 , P2_U4237 , P2_U4236 , P2_U4235 );
nand NAND4_6681 ( P2_U2605 , P2_U4234 , P2_U4233 , P2_U4232 , P2_U4231 );
nand NAND4_6682 ( P2_U2606 , P2_U4230 , P2_U4229 , P2_U4228 , P2_U4227 );
nand NAND4_6683 ( P2_U2607 , P2_U4226 , P2_U4225 , P2_U4224 , P2_U4223 );
nand NAND4_6684 ( P2_U2608 , P2_U4222 , P2_U4221 , P2_U4220 , P2_U4219 );
nand NAND4_6685 ( P2_U2609 , P2_U4218 , P2_U4217 , P2_U4216 , P2_U4215 );
nand NAND4_6686 ( P2_U2610 , P2_U4214 , P2_U4213 , P2_U4212 , P2_U4211 );
nand NAND4_6687 ( P2_U2611 , P2_U4210 , P2_U4209 , P2_U4208 , P2_U4207 );
nand NAND4_6688 ( P2_U2612 , P2_U4206 , P2_U4205 , P2_U4204 , P2_U4203 );
nand NAND4_6689 ( P2_U2613 , P2_U4202 , P2_U4201 , P2_U4200 , P2_U4199 );
nand NAND4_6690 ( P2_U2614 , P2_U4198 , P2_U4197 , P2_U4196 , P2_U4195 );
and AND2_6691 ( P2_U2615 , P2_INSTQUEUERD_ADDR_REG_4_ , P2_U3519 );
nand NAND2_6692 ( P2_U2616 , P2_U3706 , P2_U3705 );
nand NAND2_6693 ( P2_U2617 , P2_U3694 , P2_U3693 );
nand NAND2_6694 ( P2_U2618 , P2_U4350 , P2_U7453 );
nand NAND2_6695 ( P2_U2619 , P2_U4351 , P2_U7456 );
nand NAND2_6696 ( P2_U2620 , P2_U4353 , P2_U7462 );
nand NAND2_6697 ( P2_U2621 , P2_U4354 , P2_U7465 );
nand NAND2_6698 ( P2_U2622 , P2_U4355 , P2_U7468 );
nand NAND2_6699 ( P2_U2623 , P2_U4356 , P2_U7471 );
nand NAND2_6700 ( P2_U2624 , P2_U4357 , P2_U7474 );
nand NAND2_6701 ( P2_U2625 , P2_U4358 , P2_U7477 );
nand NAND2_6702 ( P2_U2626 , P2_U4359 , P2_U7480 );
nand NAND2_6703 ( P2_U2627 , P2_U4360 , P2_U7483 );
nand NAND2_6704 ( P2_U2628 , P2_U4361 , P2_U7486 );
nand NAND2_6705 ( P2_U2629 , P2_U4362 , P2_U7489 );
nand NAND2_6706 ( P2_U2630 , P2_U4364 , P2_U7495 );
nand NAND2_6707 ( P2_U2631 , P2_U4365 , P2_U7498 );
nand NAND2_6708 ( P2_U2632 , P2_U4366 , P2_U7501 );
nand NAND2_6709 ( P2_U2633 , P2_U4367 , P2_U7504 );
nand NAND3_6710 ( P2_U2634 , P2_U7508 , P2_U7507 , P2_U4368 );
nand NAND3_6711 ( P2_U2635 , P2_U7512 , P2_U7511 , P2_U4369 );
nand NAND3_6712 ( P2_U2636 , P2_U7516 , P2_U7515 , P2_U4370 );
nand NAND3_6713 ( P2_U2637 , P2_U7520 , P2_U7519 , P2_U4371 );
nand NAND3_6714 ( P2_U2638 , P2_U7524 , P2_U7523 , P2_U4372 );
nand NAND3_6715 ( P2_U2639 , P2_U7528 , P2_U7527 , P2_U4373 );
nand NAND3_6716 ( P2_U2640 , P2_U7434 , P2_U7433 , P2_U4344 );
nand NAND3_6717 ( P2_U2641 , P2_U7438 , P2_U7437 , P2_U4345 );
nand NAND2_6718 ( P2_U2642 , P2_U4346 , P2_U7441 );
nand NAND2_6719 ( P2_U2643 , P2_U4347 , P2_U7444 );
nand NAND2_6720 ( P2_U2644 , P2_U4348 , P2_U7447 );
nand NAND2_6721 ( P2_U2645 , P2_U4349 , P2_U7450 );
nand NAND2_6722 ( P2_U2646 , P2_U4352 , P2_U7459 );
nand NAND2_6723 ( P2_U2647 , P2_U4363 , P2_U7492 );
nand NAND2_6724 ( P2_U2648 , P2_U4374 , P2_U7531 );
nand NAND3_6725 ( P2_U2649 , P2_U7534 , P2_U3300 , P2_U4375 );
and AND2_6726 ( P2_U2650 , P2_U2352 , P2_U3242 );
and AND2_6727 ( P2_U2651 , P2_U2352 , P2_U7217 );
and AND2_6728 ( P2_U2652 , P2_U2352 , P2_U7251 );
and AND2_6729 ( P2_U2653 , P2_U2352 , P2_U7285 );
nand NAND2_6730 ( P2_U2654 , P2_U7423 , P2_U7422 );
nand NAND2_6731 ( P2_U2655 , P2_U4338 , P2_U7424 );
nand NAND2_6732 ( P2_U2656 , P2_U4340 , P2_U7427 );
nand NAND2_6733 ( P2_U2657 , P2_U4342 , P2_U7429 );
and AND2_6734 ( P2_U2658 , P2_U2354 , P2_U2598 );
and AND2_6735 ( P2_U2659 , P2_U2354 , P2_U2597 );
and AND2_6736 ( P2_U2660 , P2_U2354 , P2_U2596 );
and AND2_6737 ( P2_U2661 , P2_U2354 , P2_U2595 );
and AND2_6738 ( P2_U2662 , P2_U2354 , P2_U2594 );
and AND2_6739 ( P2_U2663 , P2_U2354 , P2_U2593 );
and AND2_6740 ( P2_U2664 , P2_U2354 , P2_U2592 );
and AND2_6741 ( P2_U2665 , P2_U2354 , P2_U2591 );
and AND2_6742 ( P2_U2666 , P2_U2614 , P2_U2355 );
and AND2_6743 ( P2_U2667 , P2_U2613 , P2_U2355 );
and AND2_6744 ( P2_U2668 , P2_U2612 , P2_U2355 );
and AND2_6745 ( P2_U2669 , P2_U2611 , P2_U2355 );
and AND2_6746 ( P2_U2670 , P2_U2610 , P2_U2355 );
and AND2_6747 ( P2_U2671 , P2_U2609 , P2_U2355 );
and AND2_6748 ( P2_U2672 , P2_U2608 , P2_U2355 );
and AND2_6749 ( P2_U2673 , P2_U2607 , P2_U2355 );
and AND2_6750 ( P2_U2674 , P2_INSTQUEUE_REG_0__7_ , P2_U2355 );
and AND2_6751 ( P2_U2675 , P2_INSTQUEUE_REG_0__6_ , P2_U2355 );
and AND2_6752 ( P2_U2676 , P2_INSTQUEUE_REG_0__5_ , P2_U2355 );
and AND2_6753 ( P2_U2677 , P2_INSTQUEUE_REG_0__4_ , P2_U2355 );
and AND2_6754 ( P2_U2678 , P2_INSTQUEUE_REG_0__3_ , P2_U2355 );
and AND2_6755 ( P2_U2679 , P2_INSTQUEUE_REG_0__2_ , P2_U2355 );
and AND2_6756 ( P2_U2680 , P2_INSTQUEUE_REG_0__1_ , P2_U2355 );
nand NAND2_6757 ( P2_U2681 , P2_U7166 , P2_U4275 );
and AND2_6758 ( P2_U2682 , P2_U2355 , P2_ADD_402_1132_U18 );
and AND2_6759 ( P2_U2683 , P2_ADD_402_1132_U19 , P2_U2355 );
and AND2_6760 ( P2_U2684 , P2_ADD_402_1132_U24 , P2_U2355 );
and AND2_6761 ( P2_U2685 , P2_ADD_402_1132_U22 , P2_U2355 );
and AND2_6762 ( P2_U2686 , P2_ADD_402_1132_U21 , P2_U2355 );
and AND2_6763 ( P2_U2687 , P2_ADD_402_1132_U25 , P2_U2355 );
and AND2_6764 ( P2_U2688 , P2_ADD_402_1132_U20 , P2_U2355 );
nand NAND2_6765 ( P2_U2689 , P2_U7142 , P2_U7141 );
nand NAND2_6766 ( P2_U2690 , P2_U7144 , P2_U7143 );
nand NAND2_6767 ( P2_U2691 , P2_U7146 , P2_U7145 );
nand NAND2_6768 ( P2_U2692 , P2_U7148 , P2_U7147 );
nand NAND2_6769 ( P2_U2693 , P2_U7153 , P2_U7152 );
nand NAND2_6770 ( P2_U2694 , P2_U7155 , P2_U7154 );
nand NAND2_6771 ( P2_U2695 , P2_U7157 , P2_U7156 );
nand NAND2_6772 ( P2_U2696 , P2_U7159 , P2_U7158 );
nand NAND2_6773 ( P1_ADD_405_U172 , P1_ADD_405_U97 , P1_ADD_405_U7 );
and AND2_6774 ( P2_U2698 , P2_INSTQUEUERD_ADDR_REG_4_ , P2_U3554 );
nand NAND3_6775 ( P2_U2699 , P2_U7139 , P2_U7140 , P2_U7138 );
nand NAND3_6776 ( P2_U2700 , P2_U7150 , P2_U7151 , P2_U7149 );
nand NAND3_6777 ( P2_U2701 , P2_U7161 , P2_U7162 , P2_U7160 );
nand NAND3_6778 ( P2_U2702 , P2_U7164 , P2_U7165 , P2_U7163 );
nand NAND2_6779 ( P2_U2703 , P2_U7727 , P2_U7726 );
nand NAND2_6780 ( P2_U2704 , P2_U7729 , P2_U7728 );
nand NAND2_6781 ( P2_U2705 , P2_U4390 , P2_U7730 );
nand NAND3_6782 ( P2_U2706 , P2_U7732 , P2_U7733 , P2_U3550 );
nand NAND2_6783 ( P2_U2707 , P2_U4391 , P2_U7734 );
and AND2_6784 ( P2_U2708 , P2_R2219_U25 , P2_U7723 );
and AND2_6785 ( P2_U2709 , P2_R2219_U26 , P2_U7723 );
and AND2_6786 ( P2_U2710 , P2_R2219_U27 , P2_U7723 );
nand NAND2_6787 ( P2_U2711 , P2_STATE2_REG_0_ , P2_U7724 );
nand NAND3_6788 ( P2_U2712 , P2_U7871 , P2_STATE2_REG_0_ , P2_U4407 );
nand NAND2_6789 ( P2_U2713 , P2_STATE2_REG_0_ , P2_U7725 );
nand NAND3_6790 ( P2_U2714 , P2_U7871 , P2_STATE2_REG_0_ , P2_U4408 );
nand NAND2_6791 ( P2_U2715 , P2_U2356 , P2_U2616 );
nand NAND4_6792 ( P2_U2716 , P2_U7620 , P2_U7619 , P2_U7618 , P2_U7617 );
nand NAND4_6793 ( P2_U2717 , P2_U7624 , P2_U7623 , P2_U7622 , P2_U7621 );
nand NAND4_6794 ( P2_U2718 , P2_U7632 , P2_U7631 , P2_U7630 , P2_U7629 );
nand NAND4_6795 ( P2_U2719 , P2_U7636 , P2_U7635 , P2_U7634 , P2_U7633 );
nand NAND4_6796 ( P2_U2720 , P2_U7640 , P2_U7639 , P2_U7638 , P2_U7637 );
nand NAND4_6797 ( P2_U2721 , P2_U7644 , P2_U7643 , P2_U7642 , P2_U7641 );
nand NAND4_6798 ( P2_U2722 , P2_U7648 , P2_U7647 , P2_U7646 , P2_U7645 );
nand NAND4_6799 ( P2_U2723 , P2_U7652 , P2_U7651 , P2_U7650 , P2_U7649 );
nand NAND4_6800 ( P2_U2724 , P2_U7656 , P2_U7655 , P2_U7654 , P2_U7653 );
nand NAND4_6801 ( P2_U2725 , P2_U7660 , P2_U7659 , P2_U7658 , P2_U7657 );
nand NAND4_6802 ( P2_U2726 , P2_U7664 , P2_U7663 , P2_U7662 , P2_U7661 );
nand NAND4_6803 ( P2_U2727 , P2_U7668 , P2_U7667 , P2_U7666 , P2_U7665 );
nand NAND4_6804 ( P2_U2728 , P2_U7676 , P2_U7675 , P2_U7674 , P2_U7673 );
nand NAND4_6805 ( P2_U2729 , P2_U7680 , P2_U7679 , P2_U7678 , P2_U7677 );
nand NAND4_6806 ( P2_U2730 , P2_U7684 , P2_U7683 , P2_U7682 , P2_U7681 );
nand NAND4_6807 ( P2_U2731 , P2_U7688 , P2_U7687 , P2_U7686 , P2_U7685 );
nand NAND4_6808 ( P2_U2732 , P2_U7692 , P2_U7691 , P2_U7690 , P2_U7689 );
nand NAND4_6809 ( P2_U2733 , P2_U7696 , P2_U7695 , P2_U7694 , P2_U7693 );
nand NAND4_6810 ( P2_U2734 , P2_U7700 , P2_U7699 , P2_U7698 , P2_U7697 );
nand NAND4_6811 ( P2_U2735 , P2_U7704 , P2_U7703 , P2_U7702 , P2_U7701 );
nand NAND4_6812 ( P2_U2736 , P2_U7708 , P2_U7707 , P2_U7706 , P2_U7705 );
nand NAND4_6813 ( P2_U2737 , P2_U7712 , P2_U7711 , P2_U7710 , P2_U7709 );
nand NAND4_6814 ( P2_U2738 , P2_U7596 , P2_U7595 , P2_U7594 , P2_U7593 );
nand NAND4_6815 ( P2_U2739 , P2_U7600 , P2_U7599 , P2_U7598 , P2_U7597 );
nand NAND4_6816 ( P2_U2740 , P2_U7604 , P2_U7603 , P2_U7602 , P2_U7601 );
nand NAND4_6817 ( P2_U2741 , P2_U7608 , P2_U7607 , P2_U7606 , P2_U7605 );
nand NAND4_6818 ( P2_U2742 , P2_U7612 , P2_U7611 , P2_U7610 , P2_U7609 );
nand NAND4_6819 ( P2_U2743 , P2_U7616 , P2_U7615 , P2_U7614 , P2_U7613 );
nand NAND4_6820 ( P2_U2744 , P2_U7628 , P2_U7627 , P2_U7626 , P2_U7625 );
nand NAND4_6821 ( P2_U2745 , P2_U7672 , P2_U7671 , P2_U7670 , P2_U7669 );
nand NAND4_6822 ( P2_U2746 , P2_U7716 , P2_U7715 , P2_U7714 , P2_U7713 );
nand NAND5_6823 ( P2_U2747 , P2_U7886 , P2_U7721 , P2_U4389 , P2_U4388 , P2_U7717 );
nand NAND2_6824 ( P2_U2748 , P2_U7583 , P2_U7582 );
nand NAND2_6825 ( P2_U2749 , P2_U4380 , P2_U7584 );
nand NAND2_6826 ( P2_U2750 , P2_U4382 , P2_U7588 );
and AND2_6827 ( P2_U2751 , P2_U7888 , P2_U7737 );
and AND3_6828 ( P2_U2752 , P2_U3280 , P2_INSTQUEUERD_ADDR_REG_4_ , P2_U7873 );
nand NAND2_6829 ( P2_U2753 , P2_U3286 , P2_U7572 );
nand NAND2_6830 ( P2_U2754 , P2_U3286 , P2_U7573 );
nand NAND2_6831 ( P2_U2755 , P2_U3286 , P2_U7574 );
nand NAND2_6832 ( P2_U2756 , P2_U3286 , P2_U7575 );
nand NAND2_6833 ( P2_U2757 , P2_U3286 , P2_U7576 );
and AND2_6834 ( P2_U2758 , P2_U4428 , P2_U3242 );
and AND2_6835 ( P2_U2759 , P2_U4428 , P2_U7217 );
and AND2_6836 ( P2_U2760 , P2_U4428 , P2_U7251 );
nand NAND2_6837 ( P2_U2761 , P2_U7563 , P2_U7562 );
nand NAND2_6838 ( P2_U2762 , P2_U7565 , P2_U7564 );
nand NAND2_6839 ( P2_U2763 , P2_U7567 , P2_U7566 );
nand NAND2_6840 ( P2_U2764 , P2_U7569 , P2_U7568 );
nand NAND2_6841 ( P2_U2765 , P2_U7571 , P2_U7570 );
nand NAND2_6842 ( P2_U2766 , P2_U4447 , P2_U7539 );
nand NAND2_6843 ( P2_U2767 , P2_U4447 , P2_U7540 );
nand NAND2_6844 ( P2_U2768 , P2_U4447 , P2_U7541 );
nand NAND2_6845 ( P2_U2769 , P2_U4447 , P2_U7542 );
nand NAND2_6846 ( P2_U2770 , P2_U4447 , P2_U7543 );
nand NAND2_6847 ( P2_U2771 , P2_U4447 , P2_U7544 );
nand NAND2_6848 ( P2_U2772 , P2_U4447 , P2_U7545 );
nand NAND2_6849 ( P2_U2773 , P2_U4447 , P2_U7546 );
nand NAND2_6850 ( P2_U2774 , P2_U4447 , P2_U7547 );
nand NAND2_6851 ( P2_U2775 , P2_U4447 , P2_U7548 );
nand NAND2_6852 ( P2_U2776 , P2_U4447 , P2_U7549 );
nand NAND2_6853 ( P2_U2777 , P2_U4447 , P2_U7550 );
nand NAND2_6854 ( P2_U2778 , P2_U4447 , P2_U7551 );
nand NAND2_6855 ( P2_U2779 , P2_U4447 , P2_U7552 );
nand NAND2_6856 ( P2_U2780 , P2_U4447 , P2_U7553 );
nand NAND2_6857 ( P2_U2781 , P2_U4447 , P2_U7554 );
nand NAND2_6858 ( P2_U2782 , P2_U4447 , P2_U7555 );
nand NAND2_6859 ( P2_U2783 , P2_U4447 , P2_U7556 );
nand NAND2_6860 ( P2_U2784 , P2_U4447 , P2_U7557 );
nand NAND2_6861 ( P2_U2785 , P2_U4447 , P2_U7558 );
nand NAND2_6862 ( P2_U2786 , P2_U4447 , P2_U7559 );
nand NAND2_6863 ( P2_U2787 , P2_U4447 , P2_U7560 );
nand NAND2_6864 ( P2_U2788 , P2_U4447 , P2_U7537 );
nand NAND2_6865 ( P2_U2789 , P2_U4447 , P2_U7538 );
and AND2_6866 ( P2_U2790 , P2_U3242 , P2_R2267_U63 );
and AND2_6867 ( P2_U2791 , P2_U3242 , P2_R2267_U16 );
and AND2_6868 ( P2_U2792 , P2_U3242 , P2_R2267_U15 );
and AND2_6869 ( P2_U2793 , P2_U3242 , P2_R2267_U67 );
and AND2_6870 ( P2_U2794 , P2_U3242 , P2_R2267_U14 );
and AND2_6871 ( P2_U2795 , P2_U3242 , P2_R2267_U69 );
and AND2_6872 ( P2_U2796 , P2_U3242 , P2_R2267_U13 );
and AND2_6873 ( P2_U2797 , P2_U3242 , P2_R2267_U71 );
and AND2_6874 ( P2_U2798 , P2_U3242 , P2_R2267_U12 );
and AND2_6875 ( P2_U2799 , P2_U3242 , P2_R2267_U73 );
and AND2_6876 ( P2_U2800 , P2_U3242 , P2_R2267_U11 );
and AND2_6877 ( P2_U2801 , P2_U3242 , P2_R2267_U75 );
and AND2_6878 ( P2_U2802 , P2_U3242 , P2_R2267_U10 );
and AND2_6879 ( P2_U2803 , P2_U3242 , P2_R2267_U79 );
and AND2_6880 ( P2_U2804 , P2_U3242 , P2_R2267_U9 );
and AND2_6881 ( P2_U2805 , P2_U3242 , P2_R2267_U81 );
and AND2_6882 ( P2_U2806 , P2_U3242 , P2_R2267_U8 );
and AND2_6883 ( P2_U2807 , P2_U3242 , P2_R2267_U83 );
and AND2_6884 ( P2_U2808 , P2_U3242 , P2_R2267_U7 );
and AND2_6885 ( P2_U2809 , P2_U3242 , P2_R2267_U85 );
and AND2_6886 ( P2_U2810 , P2_U3242 , P2_R2267_U6 );
and AND2_6887 ( P2_U2811 , P2_U3242 , P2_R2267_U87 );
and AND2_6888 ( P2_U2812 , P2_U3242 , P2_R2267_U20 );
and AND2_6889 ( P2_U2813 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3519 );
nand NAND2_6890 ( P2_U2814 , P2_U4190 , P2_U6861 );
nand NAND2_6891 ( P2_U2815 , P2_U7917 , P2_U6856 );
nand NAND2_6892 ( P2_U2816 , P2_U6855 , P2_U6854 );
nand NAND3_6893 ( P2_U2817 , P2_U8140 , P2_U8139 , P2_U4463 );
nand NAND3_6894 ( P2_U2818 , P2_U8136 , P2_U8135 , P2_U4463 );
nand NAND2_6895 ( P2_U2819 , P2_U6840 , P2_U6839 );
nand NAND3_6896 ( P2_U2820 , P2_U8128 , P2_U8127 , P2_U3548 );
nand NAND3_6897 ( P2_U2821 , P2_U3548 , P2_U4452 , P2_U6837 );
nand NAND2_6898 ( P2_U2822 , P2_U4398 , P2_U6836 );
nand NAND3_6899 ( P2_U2823 , P2_U8124 , P2_U8123 , P2_U4452 );
nand NAND5_6900 ( P2_U2824 , P2_U6827 , P2_U6829 , P2_U4168 , P2_U6830 , P2_U6828 );
nand NAND5_6901 ( P2_U2825 , P2_U6819 , P2_U6821 , P2_U4166 , P2_U6822 , P2_U6820 );
nand NAND5_6902 ( P2_U2826 , P2_U6811 , P2_U6813 , P2_U4164 , P2_U6814 , P2_U6812 );
nand NAND5_6903 ( P2_U2827 , P2_U6803 , P2_U6805 , P2_U4162 , P2_U6806 , P2_U6804 );
nand NAND5_6904 ( P2_U2828 , P2_U6795 , P2_U6797 , P2_U4160 , P2_U6798 , P2_U6796 );
nand NAND5_6905 ( P2_U2829 , P2_U6787 , P2_U6789 , P2_U4158 , P2_U6790 , P2_U6788 );
nand NAND5_6906 ( P2_U2830 , P2_U6779 , P2_U6781 , P2_U6782 , P2_U4156 , P2_U6780 );
nand NAND2_6907 ( P2_U2831 , P2_U6772 , P2_U4152 );
nand NAND2_6908 ( P2_U2832 , P2_U6764 , P2_U4149 );
nand NAND5_6909 ( P2_U2833 , P2_U6755 , P2_U6757 , P2_U6758 , P2_U6756 , P2_U4148 );
nand NAND2_6910 ( P2_U2834 , P2_U4146 , P2_U4144 );
nand NAND2_6911 ( P2_U2835 , P2_U4143 , P2_U4141 );
nand NAND2_6912 ( P2_U2836 , P2_U4140 , P2_U4138 );
nand NAND2_6913 ( P2_U2837 , P2_U4136 , P2_U4134 );
nand NAND2_6914 ( P2_U2838 , P2_U4132 , P2_U4130 );
nand NAND2_6915 ( P2_U2839 , P2_U4128 , P2_U4126 );
nand NAND2_6916 ( P2_U2840 , P2_U4124 , P2_U4122 );
nand NAND5_6917 ( P2_U2841 , P2_U6693 , P2_U4118 , P2_U6692 , P2_U6696 , P2_U4119 );
nand NAND5_6918 ( P2_U2842 , P2_U6685 , P2_U4115 , P2_U6684 , P2_U6688 , P2_U4116 );
nand NAND5_6919 ( P2_U2843 , P2_U6677 , P2_U4112 , P2_U6676 , P2_U6680 , P2_U4113 );
nand NAND5_6920 ( P2_U2844 , P2_U6670 , P2_U6669 , P2_U4109 , P2_U6672 , P2_U4110 );
nand NAND5_6921 ( P2_U2845 , P2_U6662 , P2_U6661 , P2_U4106 , P2_U6664 , P2_U4107 );
nand NAND5_6922 ( P2_U2846 , P2_U6654 , P2_U6653 , P2_U4103 , P2_U6656 , P2_U4104 );
nand NAND5_6923 ( P2_U2847 , P2_U6646 , P2_U6645 , P2_U4100 , P2_U6648 , P2_U4101 );
nand NAND5_6924 ( P2_U2848 , P2_U6638 , P2_U6637 , P2_U4097 , P2_U6640 , P2_U4098 );
nand NAND5_6925 ( P2_U2849 , P2_U6630 , P2_U6629 , P2_U4094 , P2_U6632 , P2_U4095 );
nand NAND2_6926 ( P2_U2850 , P2_U4093 , P2_U4091 );
nand NAND2_6927 ( P2_U2851 , P2_U4089 , P2_U4087 );
nand NAND4_6928 ( P2_U2852 , P2_U6602 , P2_U4082 , P2_U6606 , P2_U4084 );
nand NAND4_6929 ( P2_U2853 , P2_U6593 , P2_U4078 , P2_U6597 , P2_U4080 );
nand NAND4_6930 ( P2_U2854 , P2_U6584 , P2_U4074 , P2_U6588 , P2_U4076 );
nand NAND4_6931 ( P2_U2855 , P2_U6575 , P2_U4070 , P2_U6579 , P2_U4072 );
nand NAND2_6932 ( P2_U2856 , P2_U6565 , P2_U6564 );
nand NAND3_6933 ( P2_U2857 , P2_U6562 , P2_U6563 , P2_U6561 );
nand NAND3_6934 ( P2_U2858 , P2_U6559 , P2_U6560 , P2_U6558 );
nand NAND3_6935 ( P2_U2859 , P2_U6556 , P2_U6557 , P2_U6555 );
nand NAND3_6936 ( P2_U2860 , P2_U6553 , P2_U6554 , P2_U6552 );
nand NAND3_6937 ( P2_U2861 , P2_U6550 , P2_U6551 , P2_U6549 );
nand NAND3_6938 ( P2_U2862 , P2_U6547 , P2_U6548 , P2_U6546 );
nand NAND3_6939 ( P2_U2863 , P2_U6544 , P2_U6545 , P2_U6543 );
nand NAND3_6940 ( P2_U2864 , P2_U6541 , P2_U6542 , P2_U6540 );
nand NAND3_6941 ( P2_U2865 , P2_U6538 , P2_U6539 , P2_U6537 );
nand NAND3_6942 ( P2_U2866 , P2_U6535 , P2_U6536 , P2_U6534 );
nand NAND3_6943 ( P2_U2867 , P2_U6532 , P2_U6533 , P2_U6531 );
nand NAND3_6944 ( P2_U2868 , P2_U6529 , P2_U6530 , P2_U6528 );
nand NAND3_6945 ( P2_U2869 , P2_U6526 , P2_U6527 , P2_U6525 );
nand NAND3_6946 ( P2_U2870 , P2_U6523 , P2_U6524 , P2_U6522 );
nand NAND3_6947 ( P2_U2871 , P2_U6520 , P2_U6521 , P2_U6519 );
nand NAND3_6948 ( P2_U2872 , P2_U6517 , P2_U6518 , P2_U6516 );
nand NAND3_6949 ( P2_U2873 , P2_U6514 , P2_U6515 , P2_U6513 );
nand NAND3_6950 ( P2_U2874 , P2_U6511 , P2_U6512 , P2_U6510 );
nand NAND3_6951 ( P2_U2875 , P2_U6508 , P2_U6509 , P2_U6507 );
nand NAND3_6952 ( P2_U2876 , P2_U6505 , P2_U6506 , P2_U6504 );
nand NAND3_6953 ( P2_U2877 , P2_U6502 , P2_U6503 , P2_U6501 );
nand NAND3_6954 ( P2_U2878 , P2_U6499 , P2_U6500 , P2_U6498 );
nand NAND3_6955 ( P2_U2879 , P2_U6496 , P2_U6497 , P2_U6495 );
nand NAND3_6956 ( P2_U2880 , P2_U6493 , P2_U6492 , P2_U6494 );
nand NAND3_6957 ( P2_U2881 , P2_U6490 , P2_U6489 , P2_U6491 );
nand NAND3_6958 ( P2_U2882 , P2_U6487 , P2_U6486 , P2_U6488 );
nand NAND3_6959 ( P2_U2883 , P2_U6484 , P2_U6483 , P2_U6485 );
nand NAND3_6960 ( P2_U2884 , P2_U6481 , P2_U6480 , P2_U6482 );
nand NAND3_6961 ( P2_U2885 , P2_U6478 , P2_U6477 , P2_U6479 );
nand NAND3_6962 ( P2_U2886 , P2_U6475 , P2_U6474 , P2_U6476 );
nand NAND3_6963 ( P2_U2887 , P2_U6472 , P2_U6471 , P2_U6473 );
nand NAND3_6964 ( P2_U2888 , P2_U6468 , P2_U6466 , P2_U6467 );
nand NAND5_6965 ( P2_U2889 , P2_U6462 , P2_U6461 , P2_U6465 , P2_U6464 , P2_U6463 );
nand NAND5_6966 ( P2_U2890 , P2_U6457 , P2_U6456 , P2_U6460 , P2_U6459 , P2_U6458 );
nand NAND5_6967 ( P2_U2891 , P2_U6452 , P2_U6451 , P2_U6455 , P2_U6454 , P2_U6453 );
nand NAND5_6968 ( P2_U2892 , P2_U6447 , P2_U6446 , P2_U6450 , P2_U6449 , P2_U6448 );
nand NAND5_6969 ( P2_U2893 , P2_U6442 , P2_U6441 , P2_U6445 , P2_U6444 , P2_U6443 );
nand NAND5_6970 ( P2_U2894 , P2_U6437 , P2_U6436 , P2_U6440 , P2_U6439 , P2_U6438 );
nand NAND5_6971 ( P2_U2895 , P2_U6432 , P2_U6431 , P2_U6435 , P2_U6434 , P2_U6433 );
nand NAND5_6972 ( P2_U2896 , P2_U6427 , P2_U6426 , P2_U6430 , P2_U6429 , P2_U6428 );
nand NAND5_6973 ( P2_U2897 , P2_U6422 , P2_U6421 , P2_U6425 , P2_U6424 , P2_U6423 );
nand NAND5_6974 ( P2_U2898 , P2_U6417 , P2_U6416 , P2_U6420 , P2_U6419 , P2_U6418 );
nand NAND5_6975 ( P2_U2899 , P2_U6412 , P2_U6411 , P2_U6415 , P2_U6414 , P2_U6413 );
nand NAND5_6976 ( P2_U2900 , P2_U6407 , P2_U6406 , P2_U6410 , P2_U6409 , P2_U6408 );
nand NAND5_6977 ( P2_U2901 , P2_U6402 , P2_U6401 , P2_U6405 , P2_U6404 , P2_U6403 );
nand NAND5_6978 ( P2_U2902 , P2_U6397 , P2_U6396 , P2_U6400 , P2_U6399 , P2_U6398 );
nand NAND5_6979 ( P2_U2903 , P2_U6392 , P2_U6391 , P2_U6395 , P2_U6394 , P2_U6393 );
nand NAND4_6980 ( P2_U2904 , P2_U6390 , P2_U6387 , P2_U6389 , P2_U6388 );
nand NAND4_6981 ( P2_U2905 , P2_U6386 , P2_U6383 , P2_U6385 , P2_U6384 );
nand NAND4_6982 ( P2_U2906 , P2_U6382 , P2_U6379 , P2_U6381 , P2_U6380 );
nand NAND4_6983 ( P2_U2907 , P2_U6378 , P2_U6375 , P2_U6377 , P2_U6376 );
nand NAND4_6984 ( P2_U2908 , P2_U6374 , P2_U6371 , P2_U6373 , P2_U6372 );
nand NAND4_6985 ( P2_U2909 , P2_U6370 , P2_U6367 , P2_U6369 , P2_U6368 );
nand NAND3_6986 ( P2_U2910 , P2_U4068 , P2_U6363 , P2_U6364 );
nand NAND3_6987 ( P2_U2911 , P2_U4067 , P2_U6359 , P2_U6360 );
nand NAND3_6988 ( P2_U2912 , P2_U4066 , P2_U6355 , P2_U6356 );
nand NAND3_6989 ( P2_U2913 , P2_U6352 , P2_U6351 , P2_U4065 );
nand NAND3_6990 ( P2_U2914 , P2_U6348 , P2_U6347 , P2_U4064 );
nand NAND3_6991 ( P2_U2915 , P2_U6344 , P2_U6343 , P2_U4063 );
nand NAND3_6992 ( P2_U2916 , P2_U6340 , P2_U6339 , P2_U4062 );
nand NAND3_6993 ( P2_U2917 , P2_U6336 , P2_U6335 , P2_U4061 );
nand NAND3_6994 ( P2_U2918 , P2_U6332 , P2_U6331 , P2_U4060 );
nand NAND3_6995 ( P2_U2919 , P2_U6328 , P2_U6327 , P2_U4059 );
and AND2_6996 ( P2_U2920 , P2_DATAO_REG_31_ , P2_U6232 );
nand NAND3_6997 ( P2_U2921 , P2_U6324 , P2_U6323 , P2_U6325 );
nand NAND3_6998 ( P2_U2922 , P2_U6321 , P2_U6320 , P2_U6322 );
nand NAND3_6999 ( P2_U2923 , P2_U6318 , P2_U6317 , P2_U6319 );
nand NAND3_7000 ( P2_U2924 , P2_U6315 , P2_U6314 , P2_U6316 );
nand NAND3_7001 ( P2_U2925 , P2_U6312 , P2_U6311 , P2_U6313 );
nand NAND3_7002 ( P2_U2926 , P2_U6309 , P2_U6308 , P2_U6310 );
nand NAND3_7003 ( P2_U2927 , P2_U6306 , P2_U6305 , P2_U6307 );
nand NAND3_7004 ( P2_U2928 , P2_U6303 , P2_U6302 , P2_U6304 );
nand NAND3_7005 ( P2_U2929 , P2_U6300 , P2_U6299 , P2_U6301 );
nand NAND3_7006 ( P2_U2930 , P2_U6297 , P2_U6296 , P2_U6298 );
nand NAND3_7007 ( P2_U2931 , P2_U6294 , P2_U6293 , P2_U6295 );
nand NAND3_7008 ( P2_U2932 , P2_U6291 , P2_U6290 , P2_U6292 );
nand NAND3_7009 ( P2_U2933 , P2_U6288 , P2_U6287 , P2_U6289 );
nand NAND3_7010 ( P2_U2934 , P2_U6285 , P2_U6284 , P2_U6286 );
nand NAND3_7011 ( P2_U2935 , P2_U6282 , P2_U6281 , P2_U6283 );
nand NAND3_7012 ( P2_U2936 , P2_U6279 , P2_U6278 , P2_U6280 );
nand NAND3_7013 ( P2_U2937 , P2_U6276 , P2_U6275 , P2_U6277 );
nand NAND3_7014 ( P2_U2938 , P2_U6273 , P2_U6272 , P2_U6274 );
nand NAND3_7015 ( P2_U2939 , P2_U6270 , P2_U6269 , P2_U6271 );
nand NAND3_7016 ( P2_U2940 , P2_U6267 , P2_U6266 , P2_U6268 );
nand NAND3_7017 ( P2_U2941 , P2_U6264 , P2_U6263 , P2_U6265 );
nand NAND3_7018 ( P2_U2942 , P2_U6261 , P2_U6260 , P2_U6262 );
nand NAND3_7019 ( P2_U2943 , P2_U6258 , P2_U6257 , P2_U6259 );
nand NAND3_7020 ( P2_U2944 , P2_U6255 , P2_U6254 , P2_U6256 );
nand NAND3_7021 ( P2_U2945 , P2_U6252 , P2_U6251 , P2_U6253 );
nand NAND3_7022 ( P2_U2946 , P2_U6249 , P2_U6248 , P2_U6250 );
nand NAND3_7023 ( P2_U2947 , P2_U6246 , P2_U6245 , P2_U6247 );
nand NAND3_7024 ( P2_U2948 , P2_U6243 , P2_U6242 , P2_U6244 );
nand NAND3_7025 ( P2_U2949 , P2_U6240 , P2_U6239 , P2_U6241 );
nand NAND3_7026 ( P2_U2950 , P2_U6237 , P2_U6236 , P2_U6238 );
nand NAND3_7027 ( P2_U2951 , P2_U6234 , P2_U6233 , P2_U6235 );
nand NAND3_7028 ( P2_U2952 , P2_U6225 , P2_U6224 , P2_U6226 );
nand NAND3_7029 ( P2_U2953 , P2_U6222 , P2_U6221 , P2_U6223 );
nand NAND3_7030 ( P2_U2954 , P2_U6219 , P2_U6218 , P2_U6220 );
nand NAND3_7031 ( P2_U2955 , P2_U6216 , P2_U6215 , P2_U6217 );
nand NAND3_7032 ( P2_U2956 , P2_U6213 , P2_U6212 , P2_U6214 );
nand NAND3_7033 ( P2_U2957 , P2_U6210 , P2_U6209 , P2_U6211 );
nand NAND3_7034 ( P2_U2958 , P2_U6207 , P2_U6206 , P2_U6208 );
nand NAND3_7035 ( P2_U2959 , P2_U6204 , P2_U6203 , P2_U6205 );
nand NAND3_7036 ( P2_U2960 , P2_U6201 , P2_U6200 , P2_U6202 );
nand NAND3_7037 ( P2_U2961 , P2_U6198 , P2_U6197 , P2_U6199 );
nand NAND3_7038 ( P2_U2962 , P2_U6195 , P2_U6194 , P2_U6196 );
nand NAND3_7039 ( P2_U2963 , P2_U6192 , P2_U6191 , P2_U6193 );
nand NAND3_7040 ( P2_U2964 , P2_U6189 , P2_U6188 , P2_U6190 );
nand NAND3_7041 ( P2_U2965 , P2_U6186 , P2_U6185 , P2_U6187 );
nand NAND3_7042 ( P2_U2966 , P2_U6183 , P2_U6182 , P2_U6184 );
nand NAND3_7043 ( P2_U2967 , P2_U6180 , P2_U6179 , P2_U6181 );
nand NAND3_7044 ( P2_U2968 , P2_U6177 , P2_U6176 , P2_U6178 );
nand NAND3_7045 ( P2_U2969 , P2_U6174 , P2_U6173 , P2_U6175 );
nand NAND3_7046 ( P2_U2970 , P2_U6171 , P2_U6170 , P2_U6172 );
nand NAND3_7047 ( P2_U2971 , P2_U6168 , P2_U6167 , P2_U6169 );
nand NAND3_7048 ( P2_U2972 , P2_U6165 , P2_U6164 , P2_U6166 );
nand NAND3_7049 ( P2_U2973 , P2_U6162 , P2_U6161 , P2_U6163 );
nand NAND3_7050 ( P2_U2974 , P2_U6159 , P2_U6158 , P2_U6160 );
nand NAND3_7051 ( P2_U2975 , P2_U6156 , P2_U6155 , P2_U6157 );
nand NAND3_7052 ( P2_U2976 , P2_U6153 , P2_U6152 , P2_U6154 );
nand NAND3_7053 ( P2_U2977 , P2_U6150 , P2_U6149 , P2_U6151 );
nand NAND3_7054 ( P2_U2978 , P2_U6147 , P2_U6146 , P2_U6148 );
nand NAND3_7055 ( P2_U2979 , P2_U6144 , P2_U6143 , P2_U6145 );
nand NAND3_7056 ( P2_U2980 , P2_U6141 , P2_U6140 , P2_U6142 );
nand NAND3_7057 ( P2_U2981 , P2_U6138 , P2_U6137 , P2_U6139 );
nand NAND3_7058 ( P2_U2982 , P2_U6135 , P2_U6134 , P2_U6136 );
nand NAND2_7059 ( P2_U2983 , P2_U4054 , P2_U4053 );
nand NAND2_7060 ( P2_U2984 , P2_U4052 , P2_U4051 );
nand NAND2_7061 ( P2_U2985 , P2_U4050 , P2_U4049 );
nand NAND2_7062 ( P2_U2986 , P2_U4048 , P2_U4047 );
nand NAND2_7063 ( P2_U2987 , P2_U4046 , P2_U4045 );
nand NAND2_7064 ( P2_U2988 , P2_U4044 , P2_U4043 );
nand NAND2_7065 ( P2_U2989 , P2_U4042 , P2_U4041 );
nand NAND2_7066 ( P2_U2990 , P2_U4040 , P2_U4039 );
nand NAND2_7067 ( P2_U2991 , P2_U4038 , P2_U4037 );
nand NAND2_7068 ( P2_U2992 , P2_U4036 , P2_U4035 );
nand NAND2_7069 ( P2_U2993 , P2_U4034 , P2_U4033 );
nand NAND2_7070 ( P2_U2994 , P2_U4032 , P2_U4031 );
nand NAND2_7071 ( P2_U2995 , P2_U4030 , P2_U4029 );
nand NAND2_7072 ( P2_U2996 , P2_U4028 , P2_U4027 );
nand NAND2_7073 ( P2_U2997 , P2_U4026 , P2_U4025 );
nand NAND2_7074 ( P2_U2998 , P2_U4024 , P2_U4023 );
nand NAND2_7075 ( P2_U2999 , P2_U4022 , P2_U4021 );
nand NAND2_7076 ( P2_U3000 , P2_U4020 , P2_U4019 );
nand NAND2_7077 ( P2_U3001 , P2_U4018 , P2_U4017 );
nand NAND2_7078 ( P2_U3002 , P2_U4016 , P2_U4015 );
nand NAND2_7079 ( P2_U3003 , P2_U4014 , P2_U4013 );
nand NAND2_7080 ( P2_U3004 , P2_U4012 , P2_U4011 );
nand NAND2_7081 ( P2_U3005 , P2_U4010 , P2_U4009 );
nand NAND2_7082 ( P2_U3006 , P2_U4008 , P2_U4007 );
nand NAND2_7083 ( P2_U3007 , P2_U4006 , P2_U4005 );
nand NAND2_7084 ( P2_U3008 , P2_U4004 , P2_U4003 );
nand NAND2_7085 ( P2_U3009 , P2_U4002 , P2_U4001 );
nand NAND2_7086 ( P2_U3010 , P2_U4000 , P2_U3999 );
nand NAND2_7087 ( P2_U3011 , P2_U3998 , P2_U3997 );
nand NAND2_7088 ( P2_U3012 , P2_U3996 , P2_U3995 );
nand NAND2_7089 ( P2_U3013 , P2_U3994 , P2_U3993 );
nand NAND2_7090 ( P2_U3014 , P2_U3992 , P2_U3991 );
nand NAND5_7091 ( P2_U3015 , P2_U5933 , P2_U5932 , P2_U3988 , P2_U3987 , P2_U5928 );
nand NAND5_7092 ( P2_U3016 , P2_U5925 , P2_U5924 , P2_U3986 , P2_U3985 , P2_U5920 );
nand NAND4_7093 ( P2_U3017 , P2_U5917 , P2_U5916 , P2_U3984 , P2_U3983 );
nand NAND5_7094 ( P2_U3018 , P2_U5909 , P2_U5908 , P2_U3982 , P2_U3981 , P2_U3980 );
nand NAND5_7095 ( P2_U3019 , P2_U5901 , P2_U5900 , P2_U3979 , P2_U3978 , P2_U3977 );
nand NAND5_7096 ( P2_U3020 , P2_U5893 , P2_U5892 , P2_U3976 , P2_U3975 , P2_U3974 );
nand NAND5_7097 ( P2_U3021 , P2_U5885 , P2_U5884 , P2_U3973 , P2_U3972 , P2_U3971 );
nand NAND5_7098 ( P2_U3022 , P2_U5877 , P2_U5876 , P2_U3970 , P2_U3969 , P2_U3968 );
nand NAND5_7099 ( P2_U3023 , P2_U5869 , P2_U5868 , P2_U3967 , P2_U3966 , P2_U3965 );
nand NAND5_7100 ( P2_U3024 , P2_U5861 , P2_U5860 , P2_U3964 , P2_U3963 , P2_U3962 );
nand NAND5_7101 ( P2_U3025 , P2_U5853 , P2_U5852 , P2_U3961 , P2_U3960 , P2_U3959 );
nand NAND5_7102 ( P2_U3026 , P2_U5845 , P2_U5844 , P2_U3958 , P2_U3957 , P2_U3956 );
nand NAND5_7103 ( P2_U3027 , P2_U5837 , P2_U5836 , P2_U3955 , P2_U3954 , P2_U3953 );
nand NAND5_7104 ( P2_U3028 , P2_U5829 , P2_U5828 , P2_U3952 , P2_U3951 , P2_U3950 );
nand NAND5_7105 ( P2_U3029 , P2_U5821 , P2_U5820 , P2_U3949 , P2_U3948 , P2_U3947 );
nand NAND5_7106 ( P2_U3030 , P2_U5813 , P2_U5812 , P2_U3946 , P2_U3945 , P2_U3944 );
nand NAND5_7107 ( P2_U3031 , P2_U5805 , P2_U5804 , P2_U3943 , P2_U3942 , P2_U3941 );
nand NAND5_7108 ( P2_U3032 , P2_U5797 , P2_U5796 , P2_U3940 , P2_U3939 , P2_U3938 );
nand NAND5_7109 ( P2_U3033 , P2_U5789 , P2_U5788 , P2_U3937 , P2_U3936 , P2_U3935 );
nand NAND5_7110 ( P2_U3034 , P2_U5781 , P2_U5780 , P2_U3934 , P2_U3933 , P2_U3932 );
nand NAND5_7111 ( P2_U3035 , P2_U5773 , P2_U5772 , P2_U3931 , P2_U3930 , P2_U3929 );
nand NAND5_7112 ( P2_U3036 , P2_U5765 , P2_U5764 , P2_U3928 , P2_U3927 , P2_U3926 );
nand NAND5_7113 ( P2_U3037 , P2_U5757 , P2_U5756 , P2_U3925 , P2_U3924 , P2_U3923 );
nand NAND5_7114 ( P2_U3038 , P2_U5749 , P2_U5748 , P2_U3922 , P2_U3921 , P2_U3920 );
nand NAND5_7115 ( P2_U3039 , P2_U5741 , P2_U5740 , P2_U3919 , P2_U3918 , P2_U3917 );
nand NAND5_7116 ( P2_U3040 , P2_U5733 , P2_U5732 , P2_U3916 , P2_U3915 , P2_U3914 );
nand NAND5_7117 ( P2_U3041 , P2_U5725 , P2_U5724 , P2_U3913 , P2_U3912 , P2_U3911 );
nand NAND5_7118 ( P2_U3042 , P2_U5717 , P2_U5716 , P2_U3910 , P2_U3909 , P2_U3908 );
nand NAND5_7119 ( P2_U3043 , P2_U5709 , P2_U5708 , P2_U3907 , P2_U3906 , P2_U3905 );
nand NAND5_7120 ( P2_U3044 , P2_U5701 , P2_U5700 , P2_U3904 , P2_U3903 , P2_U3902 );
nand NAND5_7121 ( P2_U3045 , P2_U5693 , P2_U5692 , P2_U3901 , P2_U3900 , P2_U3899 );
nand NAND5_7122 ( P2_U3046 , P2_U5685 , P2_U5684 , P2_U3898 , P2_U3897 , P2_U3896 );
and AND2_7123 ( P2_U3047 , P2_INSTQUEUEWR_ADDR_REG_4_ , P2_U5643 );
nand NAND3_7124 ( P2_U3048 , P2_U5570 , P2_U5569 , P2_U3865 );
nand NAND3_7125 ( P2_U3049 , P2_U5565 , P2_U5564 , P2_U3864 );
nand NAND3_7126 ( P2_U3050 , P2_U5560 , P2_U5559 , P2_U3863 );
nand NAND3_7127 ( P2_U3051 , P2_U5555 , P2_U5554 , P2_U3862 );
nand NAND3_7128 ( P2_U3052 , P2_U5550 , P2_U5549 , P2_U3861 );
nand NAND3_7129 ( P2_U3053 , P2_U5545 , P2_U5544 , P2_U3860 );
nand NAND3_7130 ( P2_U3054 , P2_U5540 , P2_U5539 , P2_U3859 );
nand NAND3_7131 ( P2_U3055 , P2_U5535 , P2_U5534 , P2_U3858 );
nand NAND3_7132 ( P2_U3056 , P2_U5513 , P2_U5512 , P2_U3856 );
nand NAND3_7133 ( P2_U3057 , P2_U5508 , P2_U5507 , P2_U3855 );
nand NAND3_7134 ( P2_U3058 , P2_U5503 , P2_U5502 , P2_U3854 );
nand NAND3_7135 ( P2_U3059 , P2_U5498 , P2_U5497 , P2_U3853 );
nand NAND3_7136 ( P2_U3060 , P2_U5493 , P2_U5492 , P2_U3852 );
nand NAND3_7137 ( P2_U3061 , P2_U5488 , P2_U5487 , P2_U3851 );
nand NAND3_7138 ( P2_U3062 , P2_U5483 , P2_U5482 , P2_U3850 );
nand NAND3_7139 ( P2_U3063 , P2_U5478 , P2_U5477 , P2_U3849 );
nand NAND3_7140 ( P2_U3064 , P2_U5455 , P2_U5454 , P2_U3847 );
nand NAND3_7141 ( P2_U3065 , P2_U5450 , P2_U5449 , P2_U3846 );
nand NAND3_7142 ( P2_U3066 , P2_U5445 , P2_U5444 , P2_U3845 );
nand NAND3_7143 ( P2_U3067 , P2_U5440 , P2_U5439 , P2_U3844 );
nand NAND3_7144 ( P2_U3068 , P2_U5435 , P2_U5434 , P2_U3843 );
nand NAND3_7145 ( P2_U3069 , P2_U5430 , P2_U5429 , P2_U3842 );
nand NAND3_7146 ( P2_U3070 , P2_U5425 , P2_U5424 , P2_U3841 );
nand NAND3_7147 ( P2_U3071 , P2_U5420 , P2_U5419 , P2_U3840 );
nand NAND3_7148 ( P2_U3072 , P2_U5398 , P2_U5397 , P2_U3838 );
nand NAND3_7149 ( P2_U3073 , P2_U5393 , P2_U5392 , P2_U3837 );
nand NAND3_7150 ( P2_U3074 , P2_U5388 , P2_U5387 , P2_U3836 );
nand NAND3_7151 ( P2_U3075 , P2_U5383 , P2_U5382 , P2_U3835 );
nand NAND3_7152 ( P2_U3076 , P2_U5378 , P2_U5377 , P2_U3834 );
nand NAND3_7153 ( P2_U3077 , P2_U5373 , P2_U5372 , P2_U3833 );
nand NAND3_7154 ( P2_U3078 , P2_U5368 , P2_U5367 , P2_U3832 );
nand NAND3_7155 ( P2_U3079 , P2_U5363 , P2_U5362 , P2_U3831 );
nand NAND3_7156 ( P2_U3080 , P2_U5340 , P2_U5339 , P2_U3829 );
nand NAND3_7157 ( P2_U3081 , P2_U5335 , P2_U5334 , P2_U3828 );
nand NAND3_7158 ( P2_U3082 , P2_U5330 , P2_U5329 , P2_U3827 );
nand NAND3_7159 ( P2_U3083 , P2_U5325 , P2_U5324 , P2_U3826 );
nand NAND3_7160 ( P2_U3084 , P2_U5320 , P2_U5319 , P2_U3825 );
nand NAND3_7161 ( P2_U3085 , P2_U5315 , P2_U5314 , P2_U3824 );
nand NAND3_7162 ( P2_U3086 , P2_U5310 , P2_U5309 , P2_U3823 );
nand NAND3_7163 ( P2_U3087 , P2_U5305 , P2_U5304 , P2_U3822 );
nand NAND3_7164 ( P2_U3088 , P2_U5283 , P2_U5282 , P2_U3820 );
nand NAND3_7165 ( P2_U3089 , P2_U5278 , P2_U5277 , P2_U3819 );
nand NAND3_7166 ( P2_U3090 , P2_U5273 , P2_U5272 , P2_U3818 );
nand NAND3_7167 ( P2_U3091 , P2_U5268 , P2_U5267 , P2_U3817 );
nand NAND3_7168 ( P2_U3092 , P2_U5263 , P2_U5262 , P2_U3816 );
nand NAND3_7169 ( P2_U3093 , P2_U5258 , P2_U5257 , P2_U3815 );
nand NAND3_7170 ( P2_U3094 , P2_U5253 , P2_U5252 , P2_U3814 );
nand NAND3_7171 ( P2_U3095 , P2_U5248 , P2_U5247 , P2_U3813 );
nand NAND3_7172 ( P2_U3096 , P2_U5225 , P2_U5224 , P2_U3811 );
nand NAND3_7173 ( P2_U3097 , P2_U5220 , P2_U5219 , P2_U3810 );
nand NAND3_7174 ( P2_U3098 , P2_U5215 , P2_U5214 , P2_U3809 );
nand NAND3_7175 ( P2_U3099 , P2_U5210 , P2_U5209 , P2_U3808 );
nand NAND3_7176 ( P2_U3100 , P2_U5205 , P2_U5204 , P2_U3807 );
nand NAND3_7177 ( P2_U3101 , P2_U5200 , P2_U5199 , P2_U3806 );
nand NAND3_7178 ( P2_U3102 , P2_U5195 , P2_U5194 , P2_U3805 );
nand NAND3_7179 ( P2_U3103 , P2_U5190 , P2_U5189 , P2_U3804 );
nand NAND3_7180 ( P2_U3104 , P2_U5168 , P2_U5167 , P2_U3802 );
nand NAND3_7181 ( P2_U3105 , P2_U5163 , P2_U5162 , P2_U3801 );
nand NAND3_7182 ( P2_U3106 , P2_U5158 , P2_U5157 , P2_U3800 );
nand NAND3_7183 ( P2_U3107 , P2_U5153 , P2_U5152 , P2_U3799 );
nand NAND3_7184 ( P2_U3108 , P2_U5148 , P2_U5147 , P2_U3798 );
nand NAND3_7185 ( P2_U3109 , P2_U5143 , P2_U5142 , P2_U3797 );
nand NAND3_7186 ( P2_U3110 , P2_U5138 , P2_U5137 , P2_U3796 );
nand NAND3_7187 ( P2_U3111 , P2_U5133 , P2_U5132 , P2_U3795 );
nand NAND3_7188 ( P2_U3112 , P2_U5112 , P2_U5111 , P2_U3793 );
nand NAND3_7189 ( P2_U3113 , P2_U5107 , P2_U5106 , P2_U3792 );
nand NAND3_7190 ( P2_U3114 , P2_U5102 , P2_U5101 , P2_U3791 );
nand NAND3_7191 ( P2_U3115 , P2_U5097 , P2_U5096 , P2_U3790 );
nand NAND3_7192 ( P2_U3116 , P2_U5092 , P2_U5091 , P2_U3789 );
nand NAND3_7193 ( P2_U3117 , P2_U5087 , P2_U5086 , P2_U3788 );
nand NAND3_7194 ( P2_U3118 , P2_U5082 , P2_U5081 , P2_U3787 );
nand NAND3_7195 ( P2_U3119 , P2_U5077 , P2_U5076 , P2_U3786 );
nand NAND3_7196 ( P2_U3120 , P2_U5055 , P2_U5054 , P2_U3784 );
nand NAND3_7197 ( P2_U3121 , P2_U5050 , P2_U5049 , P2_U3783 );
nand NAND3_7198 ( P2_U3122 , P2_U5045 , P2_U5044 , P2_U3782 );
nand NAND3_7199 ( P2_U3123 , P2_U5040 , P2_U5039 , P2_U3781 );
nand NAND3_7200 ( P2_U3124 , P2_U5035 , P2_U5034 , P2_U3780 );
nand NAND3_7201 ( P2_U3125 , P2_U5030 , P2_U5029 , P2_U3779 );
nand NAND3_7202 ( P2_U3126 , P2_U5025 , P2_U5024 , P2_U3778 );
nand NAND3_7203 ( P2_U3127 , P2_U5020 , P2_U5019 , P2_U3777 );
nand NAND3_7204 ( P2_U3128 , P2_U4997 , P2_U4996 , P2_U3775 );
nand NAND3_7205 ( P2_U3129 , P2_U4992 , P2_U4991 , P2_U3774 );
nand NAND3_7206 ( P2_U3130 , P2_U4987 , P2_U4986 , P2_U3773 );
nand NAND3_7207 ( P2_U3131 , P2_U4982 , P2_U4981 , P2_U3772 );
nand NAND3_7208 ( P2_U3132 , P2_U4977 , P2_U4976 , P2_U3771 );
nand NAND3_7209 ( P2_U3133 , P2_U4972 , P2_U4971 , P2_U3770 );
nand NAND3_7210 ( P2_U3134 , P2_U4967 , P2_U4966 , P2_U3769 );
nand NAND3_7211 ( P2_U3135 , P2_U4962 , P2_U4961 , P2_U3768 );
nand NAND3_7212 ( P2_U3136 , P2_U4940 , P2_U4939 , P2_U3766 );
nand NAND3_7213 ( P2_U3137 , P2_U4935 , P2_U4934 , P2_U3765 );
nand NAND3_7214 ( P2_U3138 , P2_U4930 , P2_U4929 , P2_U3764 );
nand NAND3_7215 ( P2_U3139 , P2_U4925 , P2_U4924 , P2_U3763 );
nand NAND3_7216 ( P2_U3140 , P2_U4920 , P2_U4919 , P2_U3762 );
nand NAND3_7217 ( P2_U3141 , P2_U4915 , P2_U4914 , P2_U3761 );
nand NAND3_7218 ( P2_U3142 , P2_U4910 , P2_U4909 , P2_U3760 );
nand NAND3_7219 ( P2_U3143 , P2_U4905 , P2_U4904 , P2_U3759 );
nand NAND3_7220 ( P2_U3144 , P2_U4882 , P2_U4881 , P2_U3757 );
nand NAND3_7221 ( P2_U3145 , P2_U4877 , P2_U4876 , P2_U3756 );
nand NAND3_7222 ( P2_U3146 , P2_U4872 , P2_U4871 , P2_U3755 );
nand NAND3_7223 ( P2_U3147 , P2_U4867 , P2_U4866 , P2_U3754 );
nand NAND3_7224 ( P2_U3148 , P2_U4862 , P2_U4861 , P2_U3753 );
nand NAND3_7225 ( P2_U3149 , P2_U4857 , P2_U4856 , P2_U3752 );
nand NAND3_7226 ( P2_U3150 , P2_U4852 , P2_U4851 , P2_U3751 );
nand NAND3_7227 ( P2_U3151 , P2_U4847 , P2_U4846 , P2_U3750 );
nand NAND3_7228 ( P2_U3152 , P2_U4825 , P2_U4824 , P2_U3748 );
nand NAND3_7229 ( P2_U3153 , P2_U4820 , P2_U4819 , P2_U3747 );
nand NAND3_7230 ( P2_U3154 , P2_U4815 , P2_U4814 , P2_U3746 );
nand NAND3_7231 ( P2_U3155 , P2_U4810 , P2_U4809 , P2_U3745 );
nand NAND3_7232 ( P2_U3156 , P2_U4805 , P2_U4804 , P2_U3744 );
nand NAND3_7233 ( P2_U3157 , P2_U4800 , P2_U4799 , P2_U3743 );
nand NAND3_7234 ( P2_U3158 , P2_U4795 , P2_U4794 , P2_U3742 );
nand NAND3_7235 ( P2_U3159 , P2_U4790 , P2_U4789 , P2_U3741 );
nand NAND3_7236 ( P2_U3160 , P2_U4766 , P2_U4765 , P2_U3739 );
nand NAND3_7237 ( P2_U3161 , P2_U4761 , P2_U4760 , P2_U3738 );
nand NAND3_7238 ( P2_U3162 , P2_U4756 , P2_U4755 , P2_U3737 );
nand NAND3_7239 ( P2_U3163 , P2_U4751 , P2_U4750 , P2_U3736 );
nand NAND3_7240 ( P2_U3164 , P2_U4746 , P2_U4745 , P2_U3735 );
nand NAND3_7241 ( P2_U3165 , P2_U4741 , P2_U4740 , P2_U3734 );
nand NAND3_7242 ( P2_U3166 , P2_U4736 , P2_U4735 , P2_U3733 );
nand NAND3_7243 ( P2_U3167 , P2_U4731 , P2_U4730 , P2_U3732 );
nand NAND3_7244 ( P2_U3168 , P2_U4708 , P2_U4707 , P2_U3730 );
nand NAND3_7245 ( P2_U3169 , P2_U4703 , P2_U4702 , P2_U3729 );
nand NAND3_7246 ( P2_U3170 , P2_U4698 , P2_U4697 , P2_U3728 );
nand NAND3_7247 ( P2_U3171 , P2_U4693 , P2_U4692 , P2_U3727 );
nand NAND3_7248 ( P2_U3172 , P2_U4688 , P2_U4687 , P2_U3726 );
nand NAND3_7249 ( P2_U3173 , P2_U4683 , P2_U4682 , P2_U3725 );
nand NAND3_7250 ( P2_U3174 , P2_U4678 , P2_U4677 , P2_U3724 );
nand NAND3_7251 ( P2_U3175 , P2_U4673 , P2_U4672 , P2_U3723 );
nand NAND3_7252 ( P2_U3176 , P2_U8061 , P2_U8060 , P2_U3721 );
nand NAND4_7253 ( P2_U3177 , P2_U4629 , P2_U4628 , P2_U4627 , P2_U4454 );
nand NAND2_7254 ( P2_U3178 , P2_U3716 , P2_U4625 );
and AND2_7255 ( P2_U3179 , P2_DATAWIDTH_REG_31_ , P2_U7917 );
and AND2_7256 ( P2_U3180 , P2_DATAWIDTH_REG_30_ , P2_U7917 );
and AND2_7257 ( P2_U3181 , P2_DATAWIDTH_REG_29_ , P2_U7917 );
and AND2_7258 ( P2_U3182 , P2_DATAWIDTH_REG_28_ , P2_U7917 );
and AND2_7259 ( P2_U3183 , P2_DATAWIDTH_REG_27_ , P2_U7917 );
and AND2_7260 ( P2_U3184 , P2_DATAWIDTH_REG_26_ , P2_U7917 );
and AND2_7261 ( P2_U3185 , P2_DATAWIDTH_REG_25_ , P2_U7917 );
and AND2_7262 ( P2_U3186 , P2_DATAWIDTH_REG_24_ , P2_U7917 );
and AND2_7263 ( P2_U3187 , P2_DATAWIDTH_REG_23_ , P2_U7917 );
and AND2_7264 ( P2_U3188 , P2_DATAWIDTH_REG_22_ , P2_U7917 );
and AND2_7265 ( P2_U3189 , P2_DATAWIDTH_REG_21_ , P2_U7917 );
and AND2_7266 ( P2_U3190 , P2_DATAWIDTH_REG_20_ , P2_U7917 );
and AND2_7267 ( P2_U3191 , P2_DATAWIDTH_REG_19_ , P2_U7917 );
and AND2_7268 ( P2_U3192 , P2_DATAWIDTH_REG_18_ , P2_U7917 );
and AND2_7269 ( P2_U3193 , P2_DATAWIDTH_REG_17_ , P2_U7917 );
and AND2_7270 ( P2_U3194 , P2_DATAWIDTH_REG_16_ , P2_U7917 );
and AND2_7271 ( P2_U3195 , P2_DATAWIDTH_REG_15_ , P2_U7917 );
and AND2_7272 ( P2_U3196 , P2_DATAWIDTH_REG_14_ , P2_U7917 );
and AND2_7273 ( P2_U3197 , P2_DATAWIDTH_REG_13_ , P2_U7917 );
and AND2_7274 ( P2_U3198 , P2_DATAWIDTH_REG_12_ , P2_U7917 );
and AND2_7275 ( P2_U3199 , P2_DATAWIDTH_REG_11_ , P2_U7917 );
and AND2_7276 ( P2_U3200 , P2_DATAWIDTH_REG_10_ , P2_U7917 );
and AND2_7277 ( P2_U3201 , P2_DATAWIDTH_REG_9_ , P2_U7917 );
and AND2_7278 ( P2_U3202 , P2_DATAWIDTH_REG_8_ , P2_U7917 );
and AND2_7279 ( P2_U3203 , P2_DATAWIDTH_REG_7_ , P2_U7917 );
and AND2_7280 ( P2_U3204 , P2_DATAWIDTH_REG_6_ , P2_U7917 );
and AND2_7281 ( P2_U3205 , P2_DATAWIDTH_REG_5_ , P2_U7917 );
and AND2_7282 ( P2_U3206 , P2_DATAWIDTH_REG_4_ , P2_U7917 );
and AND2_7283 ( P2_U3207 , P2_DATAWIDTH_REG_3_ , P2_U7917 );
and AND2_7284 ( P2_U3208 , P2_DATAWIDTH_REG_2_ , P2_U7917 );
nand NAND3_7285 ( P2_U3209 , P2_U7914 , P2_U7913 , P2_U4588 );
nand NAND3_7286 ( P2_U3210 , P2_U7912 , P2_U7911 , P2_U3691 );
nand NAND2_7287 ( P2_U3211 , P2_U3690 , P2_U4579 );
nand NAND3_7288 ( P2_U3212 , P2_U4566 , P2_U4565 , P2_U4567 );
nand NAND3_7289 ( P2_U3213 , P2_U4563 , P2_U4562 , P2_U4564 );
nand NAND3_7290 ( P2_U3214 , P2_U4560 , P2_U4559 , P2_U4561 );
nand NAND3_7291 ( P2_U3215 , P2_U4557 , P2_U4556 , P2_U4558 );
nand NAND3_7292 ( P2_U3216 , P2_U4554 , P2_U4553 , P2_U4555 );
nand NAND3_7293 ( P2_U3217 , P2_U4551 , P2_U4550 , P2_U4552 );
nand NAND3_7294 ( P2_U3218 , P2_U4548 , P2_U4547 , P2_U4549 );
nand NAND3_7295 ( P2_U3219 , P2_U4545 , P2_U4544 , P2_U4546 );
nand NAND3_7296 ( P2_U3220 , P2_U4542 , P2_U4541 , P2_U4543 );
nand NAND3_7297 ( P2_U3221 , P2_U4539 , P2_U4538 , P2_U4540 );
nand NAND3_7298 ( P2_U3222 , P2_U4536 , P2_U4535 , P2_U4537 );
nand NAND3_7299 ( P2_U3223 , P2_U4533 , P2_U4532 , P2_U4534 );
nand NAND3_7300 ( P2_U3224 , P2_U4530 , P2_U4529 , P2_U4531 );
nand NAND3_7301 ( P2_U3225 , P2_U4527 , P2_U4526 , P2_U4528 );
nand NAND3_7302 ( P2_U3226 , P2_U4524 , P2_U4523 , P2_U4525 );
nand NAND3_7303 ( P2_U3227 , P2_U4521 , P2_U4520 , P2_U4522 );
nand NAND3_7304 ( P2_U3228 , P2_U4518 , P2_U4517 , P2_U4519 );
nand NAND3_7305 ( P2_U3229 , P2_U4515 , P2_U4514 , P2_U4516 );
nand NAND3_7306 ( P2_U3230 , P2_U4512 , P2_U4511 , P2_U4513 );
nand NAND3_7307 ( P2_U3231 , P2_U4509 , P2_U4508 , P2_U4510 );
nand NAND3_7308 ( P2_U3232 , P2_U4506 , P2_U4505 , P2_U4507 );
nand NAND3_7309 ( P2_U3233 , P2_U4503 , P2_U4502 , P2_U4504 );
nand NAND3_7310 ( P2_U3234 , P2_U4500 , P2_U4499 , P2_U4501 );
nand NAND3_7311 ( P2_U3235 , P2_U4497 , P2_U4496 , P2_U4498 );
nand NAND3_7312 ( P2_U3236 , P2_U4494 , P2_U4493 , P2_U4495 );
nand NAND3_7313 ( P2_U3237 , P2_U4491 , P2_U4490 , P2_U4492 );
nand NAND3_7314 ( P2_U3238 , P2_U4488 , P2_U4487 , P2_U4489 );
nand NAND3_7315 ( P2_U3239 , P2_U4485 , P2_U4484 , P2_U4486 );
nand NAND3_7316 ( P2_U3240 , P2_U4482 , P2_U4481 , P2_U4483 );
nand NAND3_7317 ( P2_U3241 , P2_U4479 , P2_U4478 , P2_U4480 );
nand NAND4_7318 ( P2_U3242 , P2_U4194 , P2_U4193 , P2_U4192 , P2_U4191 );
nand NAND2_7319 ( P2_U3243 , P2_U3349 , P2_U3335 );
not NOT1_7320 ( P2_U3244 , P2_STATE_REG_2_ );
nand NAND2_7321 ( P2_U3245 , P2_U2440 , P2_U3243 );
nand NAND2_7322 ( P2_U3246 , P2_U2440 , P2_U4650 );
nand NAND2_7323 ( P2_U3247 , P2_U2442 , P2_U3243 );
nand NAND2_7324 ( P2_U3248 , P2_U2442 , P2_U4650 );
nand NAND2_7325 ( P2_U3249 , P2_U2441 , P2_U3243 );
nand NAND2_7326 ( P2_U3250 , P2_U2441 , P2_U4650 );
nand NAND2_7327 ( P2_U3251 , P2_U2443 , P2_U3243 );
nand NAND2_7328 ( P2_U3252 , P2_U2443 , P2_U4650 );
nand NAND2_7329 ( P2_U3253 , P2_U3708 , P2_U3707 );
nand NAND2_7330 ( P2_U3254 , P2_U2590 , P2_U4429 );
nand NAND2_7331 ( P2_U3255 , P2_U3696 , P2_U3695 );
not NOT1_7332 ( P2_U3256 , P2_REQUESTPENDING_REG );
nand NAND4_7333 ( P2_U3257 , P2_U8051 , P2_U8050 , P2_U4609 , P2_U4608 );
not NOT1_7334 ( P2_U3258 , P2_STATE_REG_1_ );
nand NAND2_7335 ( P2_U3259 , P2_STATE_REG_1_ , P2_U3266 );
nand NAND2_7336 ( P2_U3260 , P2_U4439 , P2_U3244 );
nand NAND2_7337 ( P2_U3261 , P2_U4439 , P2_STATE_REG_2_ );
nand NAND2_7338 ( P2_U3262 , P2_STATE_REG_1_ , P2_U3244 );
or OR2_7339 ( P2_U3263 , P2_STATE_REG_2_ , P2_STATE_REG_1_ );
not NOT1_7340 ( P2_U3264 , HOLD );
not NOT1_7341 ( P2_U3265 , U211 );
not NOT1_7342 ( P2_U3266 , P2_STATE_REG_0_ );
nand NAND2_7343 ( P2_U3267 , P2_REQUESTPENDING_REG , P2_U3264 );
or OR2_7344 ( P2_U3268 , HOLD , P2_REQUESTPENDING_REG );
not NOT1_7345 ( P2_U3269 , P2_STATE2_REG_1_ );
not NOT1_7346 ( P2_U3270 , P2_STATE2_REG_2_ );
not NOT1_7347 ( P2_U3271 , P2_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_7348 ( P2_U3272 , P2_INSTQUEUERD_ADDR_REG_0_ );
not NOT1_7349 ( P2_U3273 , P2_INSTQUEUERD_ADDR_REG_3_ );
nand NAND3_7350 ( P2_U3274 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_U3276 , P2_INSTQUEUERD_ADDR_REG_0_ );
or OR3_7351 ( P2_U3275 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_INSTQUEUERD_ADDR_REG_1_ , P2_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_7352 ( P2_U3276 , P2_INSTQUEUERD_ADDR_REG_2_ );
nand NAND3_7353 ( P2_U3277 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_INSTQUEUERD_ADDR_REG_1_ , P2_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_7354 ( P2_U3278 , P2_U3700 , P2_U3699 );
nand NAND2_7355 ( P2_U3279 , P2_U3702 , P2_U3701 );
nand NAND2_7356 ( P2_U3280 , P2_U3704 , P2_U3703 );
nand NAND3_7357 ( P2_U3281 , P2_U7861 , P2_U7863 , P2_U7859 );
nand NAND3_7358 ( P2_U3282 , P2_U2457 , P2_U7869 , P2_U4476 );
nand NAND2_7359 ( P2_U3283 , P2_U3253 , P2_U7873 );
not NOT1_7360 ( P2_U3284 , P2_STATE2_REG_0_ );
nand NAND2_7361 ( P2_U3285 , P2_U4424 , P2_U3709 );
nand NAND2_7362 ( P2_U3286 , P2_U3253 , P2_U2616 );
not NOT1_7363 ( P2_U3287 , P2_GTE_370_U6 );
nand NAND3_7364 ( P2_U3288 , P2_U2457 , P2_U7859 , P2_U2458 );
nand NAND2_7365 ( P2_U3289 , P2_U2616 , P2_U7871 );
nand NAND2_7366 ( P2_U3290 , P2_U4595 , P2_U3266 );
nand NAND2_7367 ( P2_U3291 , P2_U3713 , P2_U2459 );
not NOT1_7368 ( P2_U3292 , P2_R2243_U8 );
nand NAND2_7369 ( P2_U3293 , P2_U2357 , P2_U3280 );
nand NAND2_7370 ( P2_U3294 , P2_U7871 , P2_U7873 );
nand NAND2_7371 ( P2_U3295 , P2_U7861 , P2_U2617 );
nand NAND2_7372 ( P2_U3296 , P2_U2451 , P2_U4428 );
not NOT1_7373 ( P2_U3297 , P2_R2167_U6 );
nand NAND5_7374 ( P2_U3298 , P2_U7894 , P2_U4444 , P2_LT_563_U6 , P2_U4614 , P2_U4610 );
nand NAND2_7375 ( P2_U3299 , P2_STATE2_REG_0_ , P2_U4619 );
not NOT1_7376 ( P2_U3300 , P2_STATE2_REG_3_ );
nand NAND2_7377 ( P2_U3301 , P2_STATE2_REG_0_ , P2_U3270 );
not NOT1_7378 ( P2_U3302 , P2_STATEBS16_REG );
or OR2_7379 ( P2_U3303 , P2_STATE2_REG_3_ , P2_STATE2_REG_1_ );
nand NAND2_7380 ( P2_U3304 , P2_STATE2_REG_2_ , P2_U3269 );
nand NAND2_7381 ( P2_U3305 , P2_STATE2_REG_3_ , P2_R2167_U6 );
nand NAND2_7382 ( P2_U3306 , P2_U4656 , P2_U3284 );
not NOT1_7383 ( P2_U3307 , P2_INSTQUEUEWR_ADDR_REG_0_ );
not NOT1_7384 ( P2_U3308 , P2_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_7385 ( P2_U3309 , P2_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_7386 ( P2_U3310 , P2_INSTQUEUEWR_ADDR_REG_2_ );
nand NAND2_7387 ( P2_U3311 , P2_INSTQUEUEWR_ADDR_REG_1_ , P2_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_7388 ( P2_U3312 , P2_U4642 , P2_U2464 );
or OR2_7389 ( P2_U3313 , P2_STATE2_REG_3_ , P2_STATE2_REG_2_ );
not NOT1_7390 ( P2_U3314 , P2_R2182_U69 );
not NOT1_7391 ( P2_U3315 , P2_R2182_U68 );
not NOT1_7392 ( P2_U3316 , P2_R2182_U40 );
not NOT1_7393 ( P2_U3317 , P2_R2182_U76 );
nand NAND2_7394 ( P2_U3318 , P2_R2182_U68 , P2_R2182_U69 );
nand NAND2_7395 ( P2_U3319 , P2_U3352 , P2_U3314 );
nand NAND2_7396 ( P2_U3320 , P2_U4636 , P2_U2461 );
not NOT1_7397 ( P2_U3321 , P2_R2099_U95 );
not NOT1_7398 ( P2_U3322 , P2_R2099_U96 );
not NOT1_7399 ( P2_U3323 , P2_R2099_U94 );
not NOT1_7400 ( P2_U3324 , P2_R2099_U5 );
nand NAND2_7401 ( P2_U3325 , P2_U3312 , P2_U4651 );
nand NAND2_7402 ( P2_U3326 , P2_U3570 , P2_U3312 );
not NOT1_7403 ( P2_U3327 , P2_INSTQUEUE_REG_15__7_ );
not NOT1_7404 ( P2_U3328 , P2_INSTQUEUE_REG_15__6_ );
not NOT1_7405 ( P2_U3329 , P2_INSTQUEUE_REG_15__5_ );
not NOT1_7406 ( P2_U3330 , P2_INSTQUEUE_REG_15__4_ );
not NOT1_7407 ( P2_U3331 , P2_INSTQUEUE_REG_15__3_ );
not NOT1_7408 ( P2_U3332 , P2_INSTQUEUE_REG_15__2_ );
not NOT1_7409 ( P2_U3333 , P2_INSTQUEUE_REG_15__1_ );
not NOT1_7410 ( P2_U3334 , P2_INSTQUEUE_REG_15__0_ );
nand NAND2_7411 ( P2_U3335 , P2_INSTQUEUEWR_ADDR_REG_1_ , P2_U3307 );
nand NAND2_7412 ( P2_U3336 , P2_U4649 , P2_U2464 );
nand NAND2_7413 ( P2_U3337 , P2_R2182_U68 , P2_U3314 );
nand NAND2_7414 ( P2_U3338 , P2_R2182_U69 , P2_U3352 );
nand NAND2_7415 ( P2_U3339 , P2_U4709 , P2_U2461 );
nand NAND2_7416 ( P2_U3340 , P2_U3569 , P2_U3336 );
not NOT1_7417 ( P2_U3341 , P2_INSTQUEUE_REG_14__7_ );
not NOT1_7418 ( P2_U3342 , P2_INSTQUEUE_REG_14__6_ );
not NOT1_7419 ( P2_U3343 , P2_INSTQUEUE_REG_14__5_ );
not NOT1_7420 ( P2_U3344 , P2_INSTQUEUE_REG_14__4_ );
not NOT1_7421 ( P2_U3345 , P2_INSTQUEUE_REG_14__3_ );
not NOT1_7422 ( P2_U3346 , P2_INSTQUEUE_REG_14__2_ );
not NOT1_7423 ( P2_U3347 , P2_INSTQUEUE_REG_14__1_ );
not NOT1_7424 ( P2_U3348 , P2_INSTQUEUE_REG_14__0_ );
nand NAND2_7425 ( P2_U3349 , P2_INSTQUEUEWR_ADDR_REG_0_ , P2_U3308 );
nand NAND2_7426 ( P2_U3350 , P2_U4648 , P2_U2464 );
nand NAND2_7427 ( P2_U3351 , P2_R2182_U69 , P2_U3315 );
nand NAND2_7428 ( P2_U3352 , P2_U3337 , P2_U3351 );
nand NAND2_7429 ( P2_U3353 , P2_U4635 , P2_U3314 );
nand NAND2_7430 ( P2_U3354 , P2_U4767 , P2_U2461 );
nand NAND2_7431 ( P2_U3355 , P2_U3350 , P2_U4770 );
nand NAND2_7432 ( P2_U3356 , P2_U3568 , P2_U3350 );
not NOT1_7433 ( P2_U3357 , P2_INSTQUEUE_REG_13__7_ );
not NOT1_7434 ( P2_U3358 , P2_INSTQUEUE_REG_13__6_ );
not NOT1_7435 ( P2_U3359 , P2_INSTQUEUE_REG_13__5_ );
not NOT1_7436 ( P2_U3360 , P2_INSTQUEUE_REG_13__4_ );
not NOT1_7437 ( P2_U3361 , P2_INSTQUEUE_REG_13__3_ );
not NOT1_7438 ( P2_U3362 , P2_INSTQUEUE_REG_13__2_ );
not NOT1_7439 ( P2_U3363 , P2_INSTQUEUE_REG_13__1_ );
not NOT1_7440 ( P2_U3364 , P2_INSTQUEUE_REG_13__0_ );
nand NAND2_7441 ( P2_U3365 , P2_U2478 , P2_U2464 );
nand NAND2_7442 ( P2_U3366 , P2_U2475 , P2_U2461 );
nand NAND2_7443 ( P2_U3367 , P2_U3567 , P2_U3365 );
not NOT1_7444 ( P2_U3368 , P2_INSTQUEUE_REG_12__7_ );
not NOT1_7445 ( P2_U3369 , P2_INSTQUEUE_REG_12__6_ );
not NOT1_7446 ( P2_U3370 , P2_INSTQUEUE_REG_12__5_ );
not NOT1_7447 ( P2_U3371 , P2_INSTQUEUE_REG_12__4_ );
not NOT1_7448 ( P2_U3372 , P2_INSTQUEUE_REG_12__3_ );
not NOT1_7449 ( P2_U3373 , P2_INSTQUEUE_REG_12__2_ );
not NOT1_7450 ( P2_U3374 , P2_INSTQUEUE_REG_12__1_ );
not NOT1_7451 ( P2_U3375 , P2_INSTQUEUE_REG_12__0_ );
nand NAND2_7452 ( P2_U3376 , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_U3310 );
nand NAND2_7453 ( P2_U3377 , P2_U4645 , P2_U4642 );
nand NAND2_7454 ( P2_U3378 , P2_R2182_U76 , P2_U3316 );
nand NAND2_7455 ( P2_U3379 , P2_U2481 , P2_U4636 );
nand NAND2_7456 ( P2_U3380 , P2_U3377 , P2_U4885 );
nand NAND2_7457 ( P2_U3381 , P2_U3566 , P2_U3377 );
not NOT1_7458 ( P2_U3382 , P2_INSTQUEUE_REG_11__7_ );
not NOT1_7459 ( P2_U3383 , P2_INSTQUEUE_REG_11__6_ );
not NOT1_7460 ( P2_U3384 , P2_INSTQUEUE_REG_11__5_ );
not NOT1_7461 ( P2_U3385 , P2_INSTQUEUE_REG_11__4_ );
not NOT1_7462 ( P2_U3386 , P2_INSTQUEUE_REG_11__3_ );
not NOT1_7463 ( P2_U3387 , P2_INSTQUEUE_REG_11__2_ );
not NOT1_7464 ( P2_U3388 , P2_INSTQUEUE_REG_11__1_ );
not NOT1_7465 ( P2_U3389 , P2_INSTQUEUE_REG_11__0_ );
nand NAND2_7466 ( P2_U3390 , P2_U4645 , P2_U4649 );
nand NAND2_7467 ( P2_U3391 , P2_U2481 , P2_U4709 );
nand NAND2_7468 ( P2_U3392 , P2_U3565 , P2_U3390 );
not NOT1_7469 ( P2_U3393 , P2_INSTQUEUE_REG_10__7_ );
not NOT1_7470 ( P2_U3394 , P2_INSTQUEUE_REG_10__6_ );
not NOT1_7471 ( P2_U3395 , P2_INSTQUEUE_REG_10__5_ );
not NOT1_7472 ( P2_U3396 , P2_INSTQUEUE_REG_10__4_ );
not NOT1_7473 ( P2_U3397 , P2_INSTQUEUE_REG_10__3_ );
not NOT1_7474 ( P2_U3398 , P2_INSTQUEUE_REG_10__2_ );
not NOT1_7475 ( P2_U3399 , P2_INSTQUEUE_REG_10__1_ );
not NOT1_7476 ( P2_U3400 , P2_INSTQUEUE_REG_10__0_ );
nand NAND2_7477 ( P2_U3401 , P2_U4645 , P2_U4648 );
nand NAND2_7478 ( P2_U3402 , P2_U2481 , P2_U4767 );
nand NAND2_7479 ( P2_U3403 , P2_U3401 , P2_U5000 );
nand NAND2_7480 ( P2_U3404 , P2_U3564 , P2_U3401 );
not NOT1_7481 ( P2_U3405 , P2_INSTQUEUE_REG_9__7_ );
not NOT1_7482 ( P2_U3406 , P2_INSTQUEUE_REG_9__6_ );
not NOT1_7483 ( P2_U3407 , P2_INSTQUEUE_REG_9__5_ );
not NOT1_7484 ( P2_U3408 , P2_INSTQUEUE_REG_9__4_ );
not NOT1_7485 ( P2_U3409 , P2_INSTQUEUE_REG_9__3_ );
not NOT1_7486 ( P2_U3410 , P2_INSTQUEUE_REG_9__2_ );
not NOT1_7487 ( P2_U3411 , P2_INSTQUEUE_REG_9__1_ );
not NOT1_7488 ( P2_U3412 , P2_INSTQUEUE_REG_9__0_ );
nand NAND2_7489 ( P2_U3413 , P2_U4645 , P2_U2478 );
nand NAND2_7490 ( P2_U3414 , P2_U2481 , P2_U2475 );
nand NAND2_7491 ( P2_U3415 , P2_U3563 , P2_U3413 );
not NOT1_7492 ( P2_U3416 , P2_INSTQUEUE_REG_8__7_ );
not NOT1_7493 ( P2_U3417 , P2_INSTQUEUE_REG_8__6_ );
not NOT1_7494 ( P2_U3418 , P2_INSTQUEUE_REG_8__5_ );
not NOT1_7495 ( P2_U3419 , P2_INSTQUEUE_REG_8__4_ );
not NOT1_7496 ( P2_U3420 , P2_INSTQUEUE_REG_8__3_ );
not NOT1_7497 ( P2_U3421 , P2_INSTQUEUE_REG_8__2_ );
not NOT1_7498 ( P2_U3422 , P2_INSTQUEUE_REG_8__1_ );
not NOT1_7499 ( P2_U3423 , P2_INSTQUEUE_REG_8__0_ );
nand NAND2_7500 ( P2_U3424 , P2_U2465 , P2_U4642 );
nand NAND2_7501 ( P2_U3425 , P2_U2460 , P2_U4637 );
nand NAND3_7502 ( P2_U3426 , P2_U3378 , P2_U4639 , P2_U3425 );
nand NAND2_7503 ( P2_U3427 , P2_U2491 , P2_U4636 );
nand NAND3_7504 ( P2_U3428 , P2_U3376 , P2_U4646 , P2_U3424 );
nand NAND2_7505 ( P2_U3429 , P2_U3424 , P2_U5114 );
nand NAND2_7506 ( P2_U3430 , P2_U3562 , P2_U3424 );
not NOT1_7507 ( P2_U3431 , P2_INSTQUEUE_REG_7__7_ );
not NOT1_7508 ( P2_U3432 , P2_INSTQUEUE_REG_7__6_ );
not NOT1_7509 ( P2_U3433 , P2_INSTQUEUE_REG_7__5_ );
not NOT1_7510 ( P2_U3434 , P2_INSTQUEUE_REG_7__4_ );
not NOT1_7511 ( P2_U3435 , P2_INSTQUEUE_REG_7__3_ );
not NOT1_7512 ( P2_U3436 , P2_INSTQUEUE_REG_7__2_ );
not NOT1_7513 ( P2_U3437 , P2_INSTQUEUE_REG_7__1_ );
not NOT1_7514 ( P2_U3438 , P2_INSTQUEUE_REG_7__0_ );
nand NAND2_7515 ( P2_U3439 , P2_U4649 , P2_U2465 );
nand NAND2_7516 ( P2_U3440 , P2_U2491 , P2_U4709 );
nand NAND2_7517 ( P2_U3441 , P2_U3561 , P2_U3439 );
not NOT1_7518 ( P2_U3442 , P2_INSTQUEUE_REG_6__7_ );
not NOT1_7519 ( P2_U3443 , P2_INSTQUEUE_REG_6__6_ );
not NOT1_7520 ( P2_U3444 , P2_INSTQUEUE_REG_6__5_ );
not NOT1_7521 ( P2_U3445 , P2_INSTQUEUE_REG_6__4_ );
not NOT1_7522 ( P2_U3446 , P2_INSTQUEUE_REG_6__3_ );
not NOT1_7523 ( P2_U3447 , P2_INSTQUEUE_REG_6__2_ );
not NOT1_7524 ( P2_U3448 , P2_INSTQUEUE_REG_6__1_ );
not NOT1_7525 ( P2_U3449 , P2_INSTQUEUE_REG_6__0_ );
nand NAND2_7526 ( P2_U3450 , P2_U4648 , P2_U2465 );
nand NAND2_7527 ( P2_U3451 , P2_U2491 , P2_U4767 );
nand NAND2_7528 ( P2_U3452 , P2_U3450 , P2_U5228 );
nand NAND2_7529 ( P2_U3453 , P2_U3560 , P2_U3450 );
not NOT1_7530 ( P2_U3454 , P2_INSTQUEUE_REG_5__7_ );
not NOT1_7531 ( P2_U3455 , P2_INSTQUEUE_REG_5__6_ );
not NOT1_7532 ( P2_U3456 , P2_INSTQUEUE_REG_5__5_ );
not NOT1_7533 ( P2_U3457 , P2_INSTQUEUE_REG_5__4_ );
not NOT1_7534 ( P2_U3458 , P2_INSTQUEUE_REG_5__3_ );
not NOT1_7535 ( P2_U3459 , P2_INSTQUEUE_REG_5__2_ );
not NOT1_7536 ( P2_U3460 , P2_INSTQUEUE_REG_5__1_ );
not NOT1_7537 ( P2_U3461 , P2_INSTQUEUE_REG_5__0_ );
nand NAND2_7538 ( P2_U3462 , P2_U2478 , P2_U2465 );
nand NAND2_7539 ( P2_U3463 , P2_U2491 , P2_U2475 );
nand NAND2_7540 ( P2_U3464 , P2_U3559 , P2_U3462 );
not NOT1_7541 ( P2_U3465 , P2_INSTQUEUE_REG_4__7_ );
not NOT1_7542 ( P2_U3466 , P2_INSTQUEUE_REG_4__6_ );
not NOT1_7543 ( P2_U3467 , P2_INSTQUEUE_REG_4__5_ );
not NOT1_7544 ( P2_U3468 , P2_INSTQUEUE_REG_4__4_ );
not NOT1_7545 ( P2_U3469 , P2_INSTQUEUE_REG_4__3_ );
not NOT1_7546 ( P2_U3470 , P2_INSTQUEUE_REG_4__2_ );
not NOT1_7547 ( P2_U3471 , P2_INSTQUEUE_REG_4__1_ );
not NOT1_7548 ( P2_U3472 , P2_INSTQUEUE_REG_4__0_ );
nand NAND2_7549 ( P2_U3473 , P2_U2503 , P2_U4642 );
nand NAND2_7550 ( P2_U3474 , P2_U2500 , P2_U4636 );
nand NAND2_7551 ( P2_U3475 , P2_U3473 , P2_U5343 );
nand NAND2_7552 ( P2_U3476 , P2_U3558 , P2_U3473 );
not NOT1_7553 ( P2_U3477 , P2_INSTQUEUE_REG_3__7_ );
not NOT1_7554 ( P2_U3478 , P2_INSTQUEUE_REG_3__6_ );
not NOT1_7555 ( P2_U3479 , P2_INSTQUEUE_REG_3__5_ );
not NOT1_7556 ( P2_U3480 , P2_INSTQUEUE_REG_3__4_ );
not NOT1_7557 ( P2_U3481 , P2_INSTQUEUE_REG_3__3_ );
not NOT1_7558 ( P2_U3482 , P2_INSTQUEUE_REG_3__2_ );
not NOT1_7559 ( P2_U3483 , P2_INSTQUEUE_REG_3__1_ );
not NOT1_7560 ( P2_U3484 , P2_INSTQUEUE_REG_3__0_ );
nand NAND2_7561 ( P2_U3485 , P2_U2503 , P2_U4649 );
nand NAND2_7562 ( P2_U3486 , P2_U2500 , P2_U4709 );
nand NAND2_7563 ( P2_U3487 , P2_U3557 , P2_U3485 );
not NOT1_7564 ( P2_U3488 , P2_INSTQUEUE_REG_2__7_ );
not NOT1_7565 ( P2_U3489 , P2_INSTQUEUE_REG_2__6_ );
not NOT1_7566 ( P2_U3490 , P2_INSTQUEUE_REG_2__5_ );
not NOT1_7567 ( P2_U3491 , P2_INSTQUEUE_REG_2__4_ );
not NOT1_7568 ( P2_U3492 , P2_INSTQUEUE_REG_2__3_ );
not NOT1_7569 ( P2_U3493 , P2_INSTQUEUE_REG_2__2_ );
not NOT1_7570 ( P2_U3494 , P2_INSTQUEUE_REG_2__1_ );
not NOT1_7571 ( P2_U3495 , P2_INSTQUEUE_REG_2__0_ );
nand NAND2_7572 ( P2_U3496 , P2_U2503 , P2_U4648 );
nand NAND2_7573 ( P2_U3497 , P2_U2500 , P2_U4767 );
nand NAND2_7574 ( P2_U3498 , P2_U3496 , P2_U5458 );
nand NAND2_7575 ( P2_U3499 , P2_U3556 , P2_U3496 );
not NOT1_7576 ( P2_U3500 , P2_INSTQUEUE_REG_1__7_ );
not NOT1_7577 ( P2_U3501 , P2_INSTQUEUE_REG_1__6_ );
not NOT1_7578 ( P2_U3502 , P2_INSTQUEUE_REG_1__5_ );
not NOT1_7579 ( P2_U3503 , P2_INSTQUEUE_REG_1__4_ );
not NOT1_7580 ( P2_U3504 , P2_INSTQUEUE_REG_1__3_ );
not NOT1_7581 ( P2_U3505 , P2_INSTQUEUE_REG_1__2_ );
not NOT1_7582 ( P2_U3506 , P2_INSTQUEUE_REG_1__1_ );
not NOT1_7583 ( P2_U3507 , P2_INSTQUEUE_REG_1__0_ );
nand NAND2_7584 ( P2_U3508 , P2_U2503 , P2_U2478 );
nand NAND2_7585 ( P2_U3509 , P2_U2500 , P2_U2475 );
nand NAND2_7586 ( P2_U3510 , P2_U3555 , P2_U3508 );
not NOT1_7587 ( P2_U3511 , P2_INSTQUEUE_REG_0__7_ );
not NOT1_7588 ( P2_U3512 , P2_INSTQUEUE_REG_0__6_ );
not NOT1_7589 ( P2_U3513 , P2_INSTQUEUE_REG_0__5_ );
not NOT1_7590 ( P2_U3514 , P2_INSTQUEUE_REG_0__4_ );
not NOT1_7591 ( P2_U3515 , P2_INSTQUEUE_REG_0__3_ );
not NOT1_7592 ( P2_U3516 , P2_INSTQUEUE_REG_0__2_ );
not NOT1_7593 ( P2_U3517 , P2_INSTQUEUE_REG_0__1_ );
not NOT1_7594 ( P2_U3518 , P2_INSTQUEUE_REG_0__0_ );
not NOT1_7595 ( P2_U3519 , P2_FLUSH_REG );
not NOT1_7596 ( P2_U3520 , P2_R2088_U6 );
nand NAND2_7597 ( P2_U3521 , P2_U3698 , P2_U3697 );
nand NAND2_7598 ( P2_U3522 , P2_U2451 , P2_U4429 );
nand NAND2_7599 ( P2_U3523 , P2_U4475 , P2_U4427 );
nand NAND2_7600 ( P2_U3524 , P2_U4429 , P2_U4475 );
nand NAND4_7601 ( P2_U3525 , P2_U7865 , P2_U7863 , P2_U3279 , P2_U7869 );
not NOT1_7602 ( P2_U3526 , P2_R2147_U8 );
nand NAND2_7603 ( P2_U3527 , P2_U3283 , P2_U3289 );
not NOT1_7604 ( P2_U3528 , P2_U3647 );
not NOT1_7605 ( P2_U3529 , P2_R2147_U9 );
nand NAND2_7606 ( P2_U3530 , P2_U3274 , P2_U5615 );
not NOT1_7607 ( P2_U3531 , P2_R2147_U4 );
not NOT1_7608 ( P2_U3532 , P2_INSTQUEUERD_ADDR_REG_0_ );
nand NAND3_7609 ( P2_U3533 , P2_U4455 , P2_U3306 , P2_U5642 );
nand NAND2_7610 ( P2_U3534 , P2_U4430 , P2_U3269 );
nand NAND2_7611 ( P2_U3535 , P2_U5672 , P2_U5671 );
nand NAND2_7612 ( P2_U3536 , P2_STATE2_REG_0_ , P2_U7873 );
nand NAND2_7613 ( P2_U3537 , P2_U5937 , P2_U5936 );
nand NAND2_7614 ( P2_U3538 , P2_U4055 , P2_U2446 );
nand NAND2_7615 ( P2_U3539 , P2_U4056 , P2_U2357 );
nand NAND2_7616 ( P2_U3540 , P2_STATE2_REG_2_ , P2_U3284 );
nand NAND2_7617 ( P2_U3541 , P2_U6231 , P2_U6230 );
nand NAND2_7618 ( P2_U3542 , P2_U2374 , P2_U6326 );
nand NAND2_7619 ( P2_U3543 , P2_U2374 , P2_U6470 );
not NOT1_7620 ( P2_U3544 , P2_EBX_REG_31_ );
or OR2_7621 ( P2_U3545 , P2_STATEBS16_REG , U211 );
nand NAND2_7622 ( P2_U3546 , P2_U4069 , P2_U4462 );
nand NAND4_7623 ( P2_U3547 , P2_U4181 , P2_U4177 , P2_U4174 , P2_U4171 );
nand NAND2_7624 ( P2_U3548 , P2_U4438 , P2_REIP_REG_1_ );
nand NAND2_7625 ( P2_U3549 , P2_U2356 , P2_U4420 );
nand NAND2_7626 ( P2_U3550 , P2_U4427 , P2_STATE2_REG_0_ );
not NOT1_7627 ( P2_U3551 , P2_CODEFETCH_REG );
not NOT1_7628 ( P2_U3552 , P2_READREQUEST_REG );
nand NAND2_7629 ( P2_U3553 , P2_U4405 , P2_U3275 );
nand NAND2_7630 ( P2_U3554 , P2_U4415 , P2_U3576 );
nand NAND2_7631 ( P2_U3555 , P2_U2504 , P2_U2479 );
nand NAND2_7632 ( P2_U3556 , P2_U2504 , P2_U2473 );
nand NAND2_7633 ( P2_U3557 , P2_U2504 , P2_U2470 );
nand NAND2_7634 ( P2_U3558 , P2_U2504 , P2_U2467 );
nand NAND2_7635 ( P2_U3559 , P2_U2492 , P2_U2479 );
nand NAND2_7636 ( P2_U3560 , P2_U2492 , P2_U2473 );
nand NAND2_7637 ( P2_U3561 , P2_U2492 , P2_U2470 );
nand NAND2_7638 ( P2_U3562 , P2_U2492 , P2_U2467 );
nand NAND2_7639 ( P2_U3563 , P2_U2483 , P2_U2479 );
nand NAND2_7640 ( P2_U3564 , P2_U2483 , P2_U2473 );
nand NAND2_7641 ( P2_U3565 , P2_U2483 , P2_U2470 );
nand NAND2_7642 ( P2_U3566 , P2_U2483 , P2_U2467 );
nand NAND2_7643 ( P2_U3567 , P2_U2479 , P2_U2466 );
nand NAND2_7644 ( P2_U3568 , P2_U2473 , P2_U2466 );
nand NAND2_7645 ( P2_U3569 , P2_U2470 , P2_U2466 );
nand NAND2_7646 ( P2_U3570 , P2_U2466 , P2_U2467 );
nand NAND2_7647 ( P2_U3571 , P2_U7865 , P2_U3300 );
not NOT1_7648 ( P2_U3572 , P2_U3242 );
or OR2_7649 ( P2_U3573 , P2_STATE2_REG_0_ , P2_STATE2_REG_1_ );
nand NAND3_7650 ( P2_U3574 , P2_U5571 , P2_U3295 , P2_U3521 );
nand NAND2_7651 ( P2_U3575 , P2_U4419 , P2_U7871 );
nand NAND2_7652 ( P2_U3576 , P2_U4419 , P2_U3279 );
nand NAND2_7653 ( P2_U3577 , P2_U4424 , P2_U6845 );
nand NAND2_7654 ( P2_U3578 , P2_U2590 , P2_U4428 );
nand NAND2_7655 ( P2_U3579 , P2_U8063 , P2_U8062 );
nand NAND2_7656 ( P2_U3580 , P2_U8066 , P2_U8065 );
nand NAND2_7657 ( P2_U3581 , P2_U8081 , P2_U8080 );
nand NAND2_7658 ( P2_U3582 , P2_U8099 , P2_U8098 );
nand NAND2_7659 ( P2_U3583 , P2_U8148 , P2_U8147 );
nand NAND2_7660 ( P2_U3584 , P2_U8151 , P2_U8150 );
nand NAND2_7661 ( P2_U3585 , P2_U7900 , P2_U7899 );
nand NAND2_7662 ( P2_U3586 , P2_U7902 , P2_U7901 );
nand NAND2_7663 ( P2_U3587 , P2_U7904 , P2_U7903 );
nand NAND2_7664 ( P2_U3588 , P2_U7906 , P2_U7905 );
nand NAND2_7665 ( P2_U3589 , P2_U7916 , P2_U7915 );
and AND2_7666 ( P2_U3590 , P2_U3263 , P2_U4401 );
nand NAND2_7667 ( P2_U3591 , P2_U7919 , P2_U7918 );
nand NAND2_7668 ( P2_U3592 , P2_U7921 , P2_U7920 );
nand NAND2_7669 ( P2_U3593 , P2_U8059 , P2_U8058 );
and AND2_7670 ( P2_U3594 , P2_U3866 , P2_U4434 );
nand NAND2_7671 ( P2_U3595 , P2_U8073 , P2_U8072 );
nand NAND2_7672 ( P2_U3596 , P2_U8084 , P2_U8083 );
nand NAND2_7673 ( P2_U3597 , P2_U8086 , P2_U8085 );
nand NAND2_7674 ( P2_U3598 , P2_U8089 , P2_U8088 );
nand NAND2_7675 ( P2_U3599 , P2_U8094 , P2_U8093 );
nand NAND2_7676 ( P2_U3600 , P2_U8102 , P2_U8101 );
nand NAND2_7677 ( P2_U3601 , P2_U8104 , P2_U8103 );
nand NAND2_7678 ( P2_U3602 , P2_U8106 , P2_U8105 );
nand NAND2_7679 ( P2_U3603 , P2_U8111 , P2_U8110 );
nand NAND2_7680 ( P2_U3604 , P2_U8113 , P2_U8112 );
nand NAND2_7681 ( P2_U3605 , P2_U8115 , P2_U8114 );
nor nor_7682 ( P2_U3606 , P2_REIP_REG_1_ , P2_DATAWIDTH_REG_1_ );
and AND2_7683 ( P2_U3607 , P2_U4183 , P2_U7898 );
nand NAND2_7684 ( P2_U3608 , P2_U8130 , P2_U8129 );
nand NAND2_7685 ( P2_U3609 , P2_U8134 , P2_U8133 );
nand NAND2_7686 ( P2_U3610 , P2_U8138 , P2_U8137 );
nand NAND2_7687 ( P2_U3611 , P2_U8142 , P2_U8141 );
nand NAND2_7688 ( P2_U3612 , P2_U8144 , P2_U8143 );
nand NAND2_7689 ( P2_U3613 , P2_U8282 , P2_U8281 );
nand NAND2_7690 ( P2_U3614 , P2_U8284 , P2_U8283 );
nand NAND2_7691 ( P2_U3615 , P2_U8286 , P2_U8285 );
and AND2_7692 ( P2_U3616 , P2_U4434 , P2_R2147_U7 );
nand NAND2_7693 ( P2_U3617 , P2_U8288 , P2_U8287 );
nand NAND2_7694 ( P2_U3618 , P2_U8290 , P2_U8289 );
nand NAND2_7695 ( P2_U3619 , P2_U8292 , P2_U8291 );
nand NAND2_7696 ( P2_U3620 , P2_U8294 , P2_U8293 );
nand NAND2_7697 ( P2_U3621 , P2_U8296 , P2_U8295 );
nand NAND2_7698 ( P2_U3622 , P2_U8298 , P2_U8297 );
nand NAND2_7699 ( P2_U3623 , P2_U8300 , P2_U8299 );
nand NAND2_7700 ( P2_U3624 , P2_U8302 , P2_U8301 );
nand NAND2_7701 ( P2_U3625 , P2_U8304 , P2_U8303 );
nand NAND2_7702 ( P2_U3626 , P2_U8306 , P2_U8305 );
nand NAND2_7703 ( P2_U3627 , P2_U8308 , P2_U8307 );
nand NAND2_7704 ( P2_U3628 , P2_U8310 , P2_U8309 );
nand NAND2_7705 ( P2_U3629 , P2_U8312 , P2_U8311 );
nand NAND2_7706 ( P2_U3630 , P2_U8314 , P2_U8313 );
nand NAND2_7707 ( P2_U3631 , P2_U8316 , P2_U8315 );
nand NAND2_7708 ( P2_U3632 , P2_U8318 , P2_U8317 );
nand NAND2_7709 ( P2_U3633 , P2_U8320 , P2_U8319 );
nand NAND2_7710 ( P2_U3634 , P2_U8322 , P2_U8321 );
nand NAND2_7711 ( P2_U3635 , P2_U8324 , P2_U8323 );
nand NAND2_7712 ( P2_U3636 , P2_U8326 , P2_U8325 );
nand NAND2_7713 ( P2_U3637 , P2_U8328 , P2_U8327 );
nand NAND2_7714 ( P2_U3638 , P2_U8330 , P2_U8329 );
nand NAND2_7715 ( P2_U3639 , P2_U8332 , P2_U8331 );
nand NAND2_7716 ( P2_U3640 , P2_U8334 , P2_U8333 );
nand NAND2_7717 ( P2_U3641 , P2_U8336 , P2_U8335 );
nand NAND2_7718 ( P2_U3642 , P2_U8338 , P2_U8337 );
nand NAND2_7719 ( P2_U3643 , P2_U8340 , P2_U8339 );
nand NAND2_7720 ( P2_U3644 , P2_U8342 , P2_U8341 );
nand NAND2_7721 ( P2_U3645 , P2_U8344 , P2_U8343 );
nand NAND2_7722 ( P2_U3646 , P2_U8346 , P2_U8345 );
nand NAND2_7723 ( P2_U3647 , P2_U8350 , P2_U8349 );
nand NAND2_7724 ( P2_U3648 , P2_U8352 , P2_U8351 );
nand NAND2_7725 ( P2_U3649 , P2_U8354 , P2_U8353 );
nand NAND2_7726 ( P2_U3650 , P2_U8356 , P2_U8355 );
nand NAND2_7727 ( P2_U3651 , P2_U8358 , P2_U8357 );
nand NAND2_7728 ( P2_U3652 , P2_U8360 , P2_U8359 );
nand NAND2_7729 ( P2_U3653 , P2_U8362 , P2_U8361 );
nand NAND2_7730 ( P2_U3654 , P2_U8364 , P2_U8363 );
nand NAND2_7731 ( P2_U3655 , P2_U8366 , P2_U8365 );
nand NAND2_7732 ( P2_U3656 , P2_U8368 , P2_U8367 );
nand NAND2_7733 ( P2_U3657 , P2_U8370 , P2_U8369 );
nand NAND2_7734 ( P2_U3658 , P2_U8372 , P2_U8371 );
nand NAND2_7735 ( P2_U3659 , P2_U8374 , P2_U8373 );
nand NAND2_7736 ( P2_U3660 , P2_U8376 , P2_U8375 );
nand NAND2_7737 ( P2_U3661 , P2_U8378 , P2_U8377 );
nand NAND2_7738 ( P2_U3662 , P2_U8380 , P2_U8379 );
nand NAND2_7739 ( P2_U3663 , P2_U8382 , P2_U8381 );
nand NAND2_7740 ( P2_U3664 , P2_U8384 , P2_U8383 );
nand NAND2_7741 ( P2_U3665 , P2_U8386 , P2_U8385 );
nand NAND2_7742 ( P2_U3666 , P2_U8388 , P2_U8387 );
nand NAND2_7743 ( P2_U3667 , P2_U8390 , P2_U8389 );
nand NAND2_7744 ( P2_U3668 , P2_U8392 , P2_U8391 );
nand NAND2_7745 ( P2_U3669 , P2_U8394 , P2_U8393 );
nand NAND2_7746 ( P2_U3670 , P2_U8396 , P2_U8395 );
nand NAND2_7747 ( P2_U3671 , P2_U8398 , P2_U8397 );
nand NAND2_7748 ( P2_U3672 , P2_U8400 , P2_U8399 );
nand NAND2_7749 ( P2_U3673 , P2_U8402 , P2_U8401 );
nand NAND2_7750 ( P2_U3674 , P2_U8404 , P2_U8403 );
nand NAND2_7751 ( P2_U3675 , P2_U8406 , P2_U8405 );
nand NAND2_7752 ( P2_U3676 , P2_U8408 , P2_U8407 );
nand NAND2_7753 ( P2_U3677 , P2_U8410 , P2_U8409 );
nand NAND2_7754 ( P2_U3678 , P2_U8412 , P2_U8411 );
nand NAND2_7755 ( P2_U3679 , P2_U8414 , P2_U8413 );
nand NAND2_7756 ( P2_U3680 , P2_U8416 , P2_U8415 );
nand NAND2_7757 ( P2_U3681 , P2_U8418 , P2_U8417 );
nand NAND2_7758 ( P2_U3682 , P2_U8420 , P2_U8419 );
nand NAND2_7759 ( P2_U3683 , P2_U8422 , P2_U8421 );
nand NAND2_7760 ( P2_U3684 , P2_U8424 , P2_U8423 );
nand NAND2_7761 ( P2_U3685 , P2_U8426 , P2_U8425 );
nand NAND2_7762 ( P2_U3686 , P2_U8428 , P2_U8427 );
nand NAND2_7763 ( P2_U3687 , P2_U8430 , P2_U8429 );
nand NAND2_7764 ( P2_U3688 , P2_U8432 , P2_U8431 );
nand NAND2_7765 ( P2_U3689 , P2_U8434 , P2_U8433 );
and AND2_7766 ( P2_U3690 , P2_U4578 , P2_U3261 );
and AND2_7767 ( P2_U3691 , P2_U4583 , P2_U3260 );
and AND2_7768 ( P2_U3692 , P2_REQUESTPENDING_REG , P2_STATE_REG_0_ );
and AND4_7769 ( P2_U3693 , P2_U7799 , P2_U7783 , P2_U7767 , P2_U7751 );
and AND4_7770 ( P2_U3694 , P2_U7868 , P2_U7847 , P2_U7831 , P2_U7815 );
and AND4_7771 ( P2_U3695 , P2_U7798 , P2_U7782 , P2_U7766 , P2_U7750 );
and AND4_7772 ( P2_U3696 , P2_U7866 , P2_U7846 , P2_U7830 , P2_U7814 );
and AND4_7773 ( P2_U3697 , P2_U7797 , P2_U7781 , P2_U7765 , P2_U7749 );
and AND4_7774 ( P2_U3698 , P2_U7864 , P2_U7845 , P2_U7829 , P2_U7813 );
and AND4_7775 ( P2_U3699 , P2_U7796 , P2_U7780 , P2_U7764 , P2_U7748 );
and AND4_7776 ( P2_U3700 , P2_U7862 , P2_U7844 , P2_U7828 , P2_U7812 );
and AND4_7777 ( P2_U3701 , P2_U7795 , P2_U7779 , P2_U7763 , P2_U7747 );
and AND4_7778 ( P2_U3702 , P2_U7860 , P2_U7843 , P2_U7827 , P2_U7811 );
and AND4_7779 ( P2_U3703 , P2_U7794 , P2_U7778 , P2_U7762 , P2_U7746 );
and AND4_7780 ( P2_U3704 , P2_U7858 , P2_U7842 , P2_U7826 , P2_U7810 );
and AND4_7781 ( P2_U3705 , P2_U7801 , P2_U7785 , P2_U7769 , P2_U7753 );
and AND4_7782 ( P2_U3706 , P2_U7872 , P2_U7849 , P2_U7833 , P2_U7817 );
and AND4_7783 ( P2_U3707 , P2_U7800 , P2_U7784 , P2_U7768 , P2_U7752 );
and AND4_7784 ( P2_U3708 , P2_U7870 , P2_U7848 , P2_U7832 , P2_U7816 );
and AND2_7785 ( P2_U3709 , P2_U3710 , P2_U4417 );
and AND2_7786 ( P2_U3710 , P2_STATE2_REG_0_ , P2_U4595 );
and AND2_7787 ( P2_U3711 , P2_U2360 , P2_U3266 );
and AND2_7788 ( P2_U3712 , P2_U3521 , P2_U7867 );
and AND2_7789 ( P2_U3713 , P2_U4599 , P2_U4598 );
and AND2_7790 ( P2_U3714 , P2_STATE2_REG_2_ , P2_U3573 );
and AND2_7791 ( P2_U3715 , P2_U3714 , P2_U4618 );
and AND2_7792 ( P2_U3716 , P2_U4624 , P2_U3304 );
and AND2_7793 ( P2_U3717 , P2_U4466 , P2_U3265 );
and AND2_7794 ( P2_U3718 , P2_STATE2_REG_3_ , P2_U3269 );
nor nor_7795 ( P2_U3719 , P2_STATE2_REG_2_ , P2_STATE2_REG_1_ );
and AND2_7796 ( P2_U3720 , P2_U4465 , P2_U4453 );
and AND2_7797 ( P2_U3721 , P2_U3720 , P2_U4632 );
and AND3_7798 ( P2_U3722 , P2_U4661 , P2_U4662 , P2_U4443 );
and AND3_7799 ( P2_U3723 , P2_U4670 , P2_U4669 , P2_U4671 );
and AND3_7800 ( P2_U3724 , P2_U4675 , P2_U4674 , P2_U4676 );
and AND3_7801 ( P2_U3725 , P2_U4680 , P2_U4679 , P2_U4681 );
and AND3_7802 ( P2_U3726 , P2_U4685 , P2_U4684 , P2_U4686 );
and AND3_7803 ( P2_U3727 , P2_U4690 , P2_U4689 , P2_U4691 );
and AND3_7804 ( P2_U3728 , P2_U4695 , P2_U4694 , P2_U4696 );
and AND3_7805 ( P2_U3729 , P2_U4700 , P2_U4699 , P2_U4701 );
and AND3_7806 ( P2_U3730 , P2_U4705 , P2_U4704 , P2_U4706 );
and AND3_7807 ( P2_U3731 , P2_U4719 , P2_U4720 , P2_U4443 );
and AND3_7808 ( P2_U3732 , P2_U4728 , P2_U4727 , P2_U4729 );
and AND3_7809 ( P2_U3733 , P2_U4733 , P2_U4732 , P2_U4734 );
and AND3_7810 ( P2_U3734 , P2_U4738 , P2_U4737 , P2_U4739 );
and AND3_7811 ( P2_U3735 , P2_U4743 , P2_U4742 , P2_U4744 );
and AND3_7812 ( P2_U3736 , P2_U4748 , P2_U4747 , P2_U4749 );
and AND3_7813 ( P2_U3737 , P2_U4753 , P2_U4752 , P2_U4754 );
and AND3_7814 ( P2_U3738 , P2_U4758 , P2_U4757 , P2_U4759 );
and AND3_7815 ( P2_U3739 , P2_U4763 , P2_U4762 , P2_U4764 );
and AND3_7816 ( P2_U3740 , P2_U4778 , P2_U4779 , P2_U4443 );
and AND3_7817 ( P2_U3741 , P2_U4787 , P2_U4786 , P2_U4788 );
and AND3_7818 ( P2_U3742 , P2_U4792 , P2_U4791 , P2_U4793 );
and AND3_7819 ( P2_U3743 , P2_U4797 , P2_U4796 , P2_U4798 );
and AND3_7820 ( P2_U3744 , P2_U4802 , P2_U4801 , P2_U4803 );
and AND3_7821 ( P2_U3745 , P2_U4807 , P2_U4806 , P2_U4808 );
and AND3_7822 ( P2_U3746 , P2_U4812 , P2_U4811 , P2_U4813 );
and AND3_7823 ( P2_U3747 , P2_U4817 , P2_U4816 , P2_U4818 );
and AND3_7824 ( P2_U3748 , P2_U4822 , P2_U4821 , P2_U4823 );
and AND3_7825 ( P2_U3749 , P2_U4835 , P2_U4836 , P2_U4443 );
and AND3_7826 ( P2_U3750 , P2_U4844 , P2_U4843 , P2_U4845 );
and AND3_7827 ( P2_U3751 , P2_U4849 , P2_U4848 , P2_U4850 );
and AND3_7828 ( P2_U3752 , P2_U4854 , P2_U4853 , P2_U4855 );
and AND3_7829 ( P2_U3753 , P2_U4859 , P2_U4858 , P2_U4860 );
and AND3_7830 ( P2_U3754 , P2_U4864 , P2_U4863 , P2_U4865 );
and AND3_7831 ( P2_U3755 , P2_U4869 , P2_U4868 , P2_U4870 );
and AND3_7832 ( P2_U3756 , P2_U4874 , P2_U4873 , P2_U4875 );
and AND3_7833 ( P2_U3757 , P2_U4879 , P2_U4878 , P2_U4880 );
and AND3_7834 ( P2_U3758 , P2_U4893 , P2_U4894 , P2_U4443 );
and AND3_7835 ( P2_U3759 , P2_U4902 , P2_U4901 , P2_U4903 );
and AND3_7836 ( P2_U3760 , P2_U4907 , P2_U4906 , P2_U4908 );
and AND3_7837 ( P2_U3761 , P2_U4912 , P2_U4911 , P2_U4913 );
and AND3_7838 ( P2_U3762 , P2_U4917 , P2_U4916 , P2_U4918 );
and AND3_7839 ( P2_U3763 , P2_U4922 , P2_U4921 , P2_U4923 );
and AND3_7840 ( P2_U3764 , P2_U4927 , P2_U4926 , P2_U4928 );
and AND3_7841 ( P2_U3765 , P2_U4932 , P2_U4931 , P2_U4933 );
and AND3_7842 ( P2_U3766 , P2_U4937 , P2_U4936 , P2_U4938 );
and AND3_7843 ( P2_U3767 , P2_U4950 , P2_U4951 , P2_U4443 );
and AND3_7844 ( P2_U3768 , P2_U4959 , P2_U4958 , P2_U4960 );
and AND3_7845 ( P2_U3769 , P2_U4964 , P2_U4963 , P2_U4965 );
and AND3_7846 ( P2_U3770 , P2_U4969 , P2_U4968 , P2_U4970 );
and AND3_7847 ( P2_U3771 , P2_U4974 , P2_U4973 , P2_U4975 );
and AND3_7848 ( P2_U3772 , P2_U4979 , P2_U4978 , P2_U4980 );
and AND3_7849 ( P2_U3773 , P2_U4984 , P2_U4983 , P2_U4985 );
and AND3_7850 ( P2_U3774 , P2_U4989 , P2_U4988 , P2_U4990 );
and AND3_7851 ( P2_U3775 , P2_U4994 , P2_U4993 , P2_U4995 );
and AND3_7852 ( P2_U3776 , P2_U5008 , P2_U5009 , P2_U4443 );
and AND3_7853 ( P2_U3777 , P2_U5017 , P2_U5016 , P2_U5018 );
and AND3_7854 ( P2_U3778 , P2_U5022 , P2_U5021 , P2_U5023 );
and AND3_7855 ( P2_U3779 , P2_U5027 , P2_U5026 , P2_U5028 );
and AND3_7856 ( P2_U3780 , P2_U5032 , P2_U5031 , P2_U5033 );
and AND3_7857 ( P2_U3781 , P2_U5037 , P2_U5036 , P2_U5038 );
and AND3_7858 ( P2_U3782 , P2_U5042 , P2_U5041 , P2_U5043 );
and AND3_7859 ( P2_U3783 , P2_U5047 , P2_U5046 , P2_U5048 );
and AND3_7860 ( P2_U3784 , P2_U5052 , P2_U5051 , P2_U5053 );
and AND3_7861 ( P2_U3785 , P2_U5065 , P2_U5066 , P2_U4443 );
and AND3_7862 ( P2_U3786 , P2_U5074 , P2_U5073 , P2_U5075 );
and AND3_7863 ( P2_U3787 , P2_U5079 , P2_U5078 , P2_U5080 );
and AND3_7864 ( P2_U3788 , P2_U5084 , P2_U5083 , P2_U5085 );
and AND3_7865 ( P2_U3789 , P2_U5089 , P2_U5088 , P2_U5090 );
and AND3_7866 ( P2_U3790 , P2_U5094 , P2_U5093 , P2_U5095 );
and AND3_7867 ( P2_U3791 , P2_U5099 , P2_U5098 , P2_U5100 );
and AND3_7868 ( P2_U3792 , P2_U5104 , P2_U5103 , P2_U5105 );
and AND3_7869 ( P2_U3793 , P2_U5109 , P2_U5108 , P2_U5110 );
and AND3_7870 ( P2_U3794 , P2_U5121 , P2_U5122 , P2_U4443 );
and AND3_7871 ( P2_U3795 , P2_U5130 , P2_U5129 , P2_U5131 );
and AND3_7872 ( P2_U3796 , P2_U5135 , P2_U5134 , P2_U5136 );
and AND3_7873 ( P2_U3797 , P2_U5140 , P2_U5139 , P2_U5141 );
and AND3_7874 ( P2_U3798 , P2_U5145 , P2_U5144 , P2_U5146 );
and AND3_7875 ( P2_U3799 , P2_U5150 , P2_U5149 , P2_U5151 );
and AND3_7876 ( P2_U3800 , P2_U5155 , P2_U5154 , P2_U5156 );
and AND3_7877 ( P2_U3801 , P2_U5160 , P2_U5159 , P2_U5161 );
and AND3_7878 ( P2_U3802 , P2_U5165 , P2_U5164 , P2_U5166 );
and AND3_7879 ( P2_U3803 , P2_U5178 , P2_U5179 , P2_U4443 );
and AND3_7880 ( P2_U3804 , P2_U5187 , P2_U5186 , P2_U5188 );
and AND3_7881 ( P2_U3805 , P2_U5192 , P2_U5191 , P2_U5193 );
and AND3_7882 ( P2_U3806 , P2_U5197 , P2_U5196 , P2_U5198 );
and AND3_7883 ( P2_U3807 , P2_U5202 , P2_U5201 , P2_U5203 );
and AND3_7884 ( P2_U3808 , P2_U5207 , P2_U5206 , P2_U5208 );
and AND3_7885 ( P2_U3809 , P2_U5212 , P2_U5211 , P2_U5213 );
and AND3_7886 ( P2_U3810 , P2_U5217 , P2_U5216 , P2_U5218 );
and AND3_7887 ( P2_U3811 , P2_U5222 , P2_U5221 , P2_U5223 );
and AND3_7888 ( P2_U3812 , P2_U5236 , P2_U5237 , P2_U4443 );
and AND3_7889 ( P2_U3813 , P2_U5245 , P2_U5244 , P2_U5246 );
and AND3_7890 ( P2_U3814 , P2_U5250 , P2_U5249 , P2_U5251 );
and AND3_7891 ( P2_U3815 , P2_U5255 , P2_U5254 , P2_U5256 );
and AND3_7892 ( P2_U3816 , P2_U5260 , P2_U5259 , P2_U5261 );
and AND3_7893 ( P2_U3817 , P2_U5265 , P2_U5264 , P2_U5266 );
and AND3_7894 ( P2_U3818 , P2_U5270 , P2_U5269 , P2_U5271 );
and AND3_7895 ( P2_U3819 , P2_U5275 , P2_U5274 , P2_U5276 );
and AND3_7896 ( P2_U3820 , P2_U5280 , P2_U5279 , P2_U5281 );
and AND3_7897 ( P2_U3821 , P2_U5293 , P2_U5294 , P2_U4443 );
and AND3_7898 ( P2_U3822 , P2_U5302 , P2_U5301 , P2_U5303 );
and AND3_7899 ( P2_U3823 , P2_U5307 , P2_U5306 , P2_U5308 );
and AND3_7900 ( P2_U3824 , P2_U5312 , P2_U5311 , P2_U5313 );
and AND3_7901 ( P2_U3825 , P2_U5317 , P2_U5316 , P2_U5318 );
and AND3_7902 ( P2_U3826 , P2_U5322 , P2_U5321 , P2_U5323 );
and AND3_7903 ( P2_U3827 , P2_U5327 , P2_U5326 , P2_U5328 );
and AND3_7904 ( P2_U3828 , P2_U5332 , P2_U5331 , P2_U5333 );
and AND3_7905 ( P2_U3829 , P2_U5337 , P2_U5336 , P2_U5338 );
and AND3_7906 ( P2_U3830 , P2_U5351 , P2_U5352 , P2_U4443 );
and AND3_7907 ( P2_U3831 , P2_U5360 , P2_U5359 , P2_U5361 );
and AND3_7908 ( P2_U3832 , P2_U5365 , P2_U5364 , P2_U5366 );
and AND3_7909 ( P2_U3833 , P2_U5370 , P2_U5369 , P2_U5371 );
and AND3_7910 ( P2_U3834 , P2_U5375 , P2_U5374 , P2_U5376 );
and AND3_7911 ( P2_U3835 , P2_U5380 , P2_U5379 , P2_U5381 );
and AND3_7912 ( P2_U3836 , P2_U5385 , P2_U5384 , P2_U5386 );
and AND3_7913 ( P2_U3837 , P2_U5390 , P2_U5389 , P2_U5391 );
and AND3_7914 ( P2_U3838 , P2_U5395 , P2_U5394 , P2_U5396 );
and AND3_7915 ( P2_U3839 , P2_U5408 , P2_U5409 , P2_U4443 );
and AND3_7916 ( P2_U3840 , P2_U5417 , P2_U5416 , P2_U5418 );
and AND3_7917 ( P2_U3841 , P2_U5422 , P2_U5421 , P2_U5423 );
and AND3_7918 ( P2_U3842 , P2_U5427 , P2_U5426 , P2_U5428 );
and AND3_7919 ( P2_U3843 , P2_U5432 , P2_U5431 , P2_U5433 );
and AND3_7920 ( P2_U3844 , P2_U5437 , P2_U5436 , P2_U5438 );
and AND3_7921 ( P2_U3845 , P2_U5442 , P2_U5441 , P2_U5443 );
and AND3_7922 ( P2_U3846 , P2_U5447 , P2_U5446 , P2_U5448 );
and AND3_7923 ( P2_U3847 , P2_U5452 , P2_U5451 , P2_U5453 );
and AND3_7924 ( P2_U3848 , P2_U5466 , P2_U5467 , P2_U4443 );
and AND3_7925 ( P2_U3849 , P2_U5475 , P2_U5474 , P2_U5476 );
and AND3_7926 ( P2_U3850 , P2_U5480 , P2_U5479 , P2_U5481 );
and AND3_7927 ( P2_U3851 , P2_U5485 , P2_U5484 , P2_U5486 );
and AND3_7928 ( P2_U3852 , P2_U5490 , P2_U5489 , P2_U5491 );
and AND3_7929 ( P2_U3853 , P2_U5495 , P2_U5494 , P2_U5496 );
and AND3_7930 ( P2_U3854 , P2_U5500 , P2_U5499 , P2_U5501 );
and AND3_7931 ( P2_U3855 , P2_U5505 , P2_U5504 , P2_U5506 );
and AND3_7932 ( P2_U3856 , P2_U5510 , P2_U5509 , P2_U5511 );
and AND3_7933 ( P2_U3857 , P2_U5523 , P2_U5524 , P2_U4443 );
and AND3_7934 ( P2_U3858 , P2_U5532 , P2_U5531 , P2_U5533 );
and AND3_7935 ( P2_U3859 , P2_U5537 , P2_U5536 , P2_U5538 );
and AND3_7936 ( P2_U3860 , P2_U5542 , P2_U5541 , P2_U5543 );
and AND3_7937 ( P2_U3861 , P2_U5547 , P2_U5546 , P2_U5548 );
and AND3_7938 ( P2_U3862 , P2_U5552 , P2_U5551 , P2_U5553 );
and AND3_7939 ( P2_U3863 , P2_U5557 , P2_U5556 , P2_U5558 );
and AND3_7940 ( P2_U3864 , P2_U5562 , P2_U5561 , P2_U5563 );
and AND3_7941 ( P2_U3865 , P2_U5567 , P2_U5566 , P2_U5568 );
and AND2_7942 ( P2_U3866 , P2_R2147_U7 , P2_U4466 );
and AND2_7943 ( P2_U3867 , P2_FLUSH_REG , P2_STATE2_REG_0_ );
and AND2_7944 ( P2_U3868 , P2_U5573 , P2_U5571 );
and AND2_7945 ( P2_U3869 , P2_U3868 , P2_U5576 );
and AND2_7946 ( P2_U3870 , P2_U4460 , P2_U4456 );
and AND4_7947 ( P2_U3871 , P2_U8071 , P2_U8070 , P2_U3870 , P2_U2512 );
and AND2_7948 ( P2_U3872 , P2_U5583 , P2_U4455 );
and AND2_7949 ( P2_U3873 , P2_U3521 , P2_U7869 );
and AND2_7950 ( P2_U3874 , P2_U7861 , P2_U3278 );
and AND2_7951 ( P2_U3875 , P2_U3874 , P2_U4429 );
and AND2_7952 ( P2_U3876 , P2_U4429 , P2_U3279 );
and AND2_7953 ( P2_U3877 , P2_U7859 , P2_U5593 );
and AND2_7954 ( P2_U3878 , P2_U7863 , P2_U3521 );
and AND3_7955 ( P2_U3879 , P2_U5587 , P2_U5588 , P2_U3281 );
and AND2_7956 ( P2_U3880 , P2_U5599 , P2_U3254 );
and AND3_7957 ( P2_U3881 , P2_U5601 , P2_U5600 , P2_U3880 );
and AND2_7958 ( P2_U3882 , P2_U7897 , P2_U5602 );
and AND2_7959 ( P2_U3883 , P2_U5608 , P2_U5607 );
and AND2_7960 ( P2_U3884 , P2_U3883 , P2_U5609 );
and AND2_7961 ( P2_U3885 , P2_U4396 , P2_U5617 );
and AND2_7962 ( P2_U3886 , P2_U4601 , P2_U2449 );
and AND2_7963 ( P2_U3887 , P2_U3582 , P2_U7859 );
and AND2_7964 ( P2_U3888 , P2_U5627 , P2_U5626 );
and AND2_7965 ( P2_U3889 , P2_U7859 , P2_U3272 );
and AND2_7966 ( P2_U3890 , P2_U5635 , P2_U5634 );
and AND2_7967 ( P2_U3891 , P2_U5649 , P2_U5650 );
and AND2_7968 ( P2_U3892 , P2_U5653 , P2_U5654 );
and AND2_7969 ( P2_U3893 , P2_U5658 , P2_U5659 );
and AND3_7970 ( P2_U3894 , P2_U4460 , P2_U5668 , P2_U4456 );
and AND2_7971 ( P2_U3895 , P2_U5674 , P2_U3578 );
and AND2_7972 ( P2_U3896 , P2_U5681 , P2_U5680 );
and AND2_7973 ( P2_U3897 , P2_U5683 , P2_U5682 );
and AND2_7974 ( P2_U3898 , P2_U5687 , P2_U5686 );
and AND2_7975 ( P2_U3899 , P2_U5689 , P2_U5688 );
and AND2_7976 ( P2_U3900 , P2_U5691 , P2_U5690 );
and AND2_7977 ( P2_U3901 , P2_U5695 , P2_U5694 );
and AND2_7978 ( P2_U3902 , P2_U5697 , P2_U5696 );
and AND2_7979 ( P2_U3903 , P2_U5699 , P2_U5698 );
and AND2_7980 ( P2_U3904 , P2_U5703 , P2_U5702 );
and AND2_7981 ( P2_U3905 , P2_U5705 , P2_U5704 );
and AND2_7982 ( P2_U3906 , P2_U5707 , P2_U5706 );
and AND2_7983 ( P2_U3907 , P2_U5711 , P2_U5710 );
and AND2_7984 ( P2_U3908 , P2_U5713 , P2_U5712 );
and AND2_7985 ( P2_U3909 , P2_U5715 , P2_U5714 );
and AND2_7986 ( P2_U3910 , P2_U5719 , P2_U5718 );
and AND2_7987 ( P2_U3911 , P2_U5721 , P2_U5720 );
and AND2_7988 ( P2_U3912 , P2_U5723 , P2_U5722 );
and AND2_7989 ( P2_U3913 , P2_U5727 , P2_U5726 );
and AND2_7990 ( P2_U3914 , P2_U5729 , P2_U5728 );
and AND2_7991 ( P2_U3915 , P2_U5731 , P2_U5730 );
and AND2_7992 ( P2_U3916 , P2_U5735 , P2_U5734 );
and AND2_7993 ( P2_U3917 , P2_U5737 , P2_U5736 );
and AND2_7994 ( P2_U3918 , P2_U5739 , P2_U5738 );
and AND2_7995 ( P2_U3919 , P2_U5743 , P2_U5742 );
and AND2_7996 ( P2_U3920 , P2_U5745 , P2_U5744 );
and AND2_7997 ( P2_U3921 , P2_U5747 , P2_U5746 );
and AND2_7998 ( P2_U3922 , P2_U5751 , P2_U5750 );
and AND2_7999 ( P2_U3923 , P2_U5753 , P2_U5752 );
and AND2_8000 ( P2_U3924 , P2_U5755 , P2_U5754 );
and AND2_8001 ( P2_U3925 , P2_U5759 , P2_U5758 );
and AND2_8002 ( P2_U3926 , P2_U5761 , P2_U5760 );
and AND2_8003 ( P2_U3927 , P2_U5763 , P2_U5762 );
and AND2_8004 ( P2_U3928 , P2_U5767 , P2_U5766 );
and AND2_8005 ( P2_U3929 , P2_U5769 , P2_U5768 );
and AND2_8006 ( P2_U3930 , P2_U5771 , P2_U5770 );
and AND2_8007 ( P2_U3931 , P2_U5775 , P2_U5774 );
and AND2_8008 ( P2_U3932 , P2_U5777 , P2_U5776 );
and AND2_8009 ( P2_U3933 , P2_U5779 , P2_U5778 );
and AND2_8010 ( P2_U3934 , P2_U5783 , P2_U5782 );
and AND2_8011 ( P2_U3935 , P2_U5785 , P2_U5784 );
and AND2_8012 ( P2_U3936 , P2_U5787 , P2_U5786 );
and AND2_8013 ( P2_U3937 , P2_U5791 , P2_U5790 );
and AND2_8014 ( P2_U3938 , P2_U5793 , P2_U5792 );
and AND2_8015 ( P2_U3939 , P2_U5795 , P2_U5794 );
and AND2_8016 ( P2_U3940 , P2_U5799 , P2_U5798 );
and AND2_8017 ( P2_U3941 , P2_U5801 , P2_U5800 );
and AND2_8018 ( P2_U3942 , P2_U5803 , P2_U5802 );
and AND2_8019 ( P2_U3943 , P2_U5807 , P2_U5806 );
and AND2_8020 ( P2_U3944 , P2_U5809 , P2_U5808 );
and AND2_8021 ( P2_U3945 , P2_U5811 , P2_U5810 );
and AND2_8022 ( P2_U3946 , P2_U5815 , P2_U5814 );
and AND2_8023 ( P2_U3947 , P2_U5817 , P2_U5816 );
and AND2_8024 ( P2_U3948 , P2_U5819 , P2_U5818 );
and AND2_8025 ( P2_U3949 , P2_U5823 , P2_U5822 );
and AND2_8026 ( P2_U3950 , P2_U5825 , P2_U5824 );
and AND2_8027 ( P2_U3951 , P2_U5827 , P2_U5826 );
and AND2_8028 ( P2_U3952 , P2_U5831 , P2_U5830 );
and AND2_8029 ( P2_U3953 , P2_U5833 , P2_U5832 );
and AND2_8030 ( P2_U3954 , P2_U5835 , P2_U5834 );
and AND2_8031 ( P2_U3955 , P2_U5839 , P2_U5838 );
and AND2_8032 ( P2_U3956 , P2_U5841 , P2_U5840 );
and AND2_8033 ( P2_U3957 , P2_U5843 , P2_U5842 );
and AND2_8034 ( P2_U3958 , P2_U5847 , P2_U5846 );
and AND2_8035 ( P2_U3959 , P2_U5849 , P2_U5848 );
and AND2_8036 ( P2_U3960 , P2_U5851 , P2_U5850 );
and AND2_8037 ( P2_U3961 , P2_U5855 , P2_U5854 );
and AND2_8038 ( P2_U3962 , P2_U5857 , P2_U5856 );
and AND2_8039 ( P2_U3963 , P2_U5859 , P2_U5858 );
and AND2_8040 ( P2_U3964 , P2_U5863 , P2_U5862 );
and AND2_8041 ( P2_U3965 , P2_U5865 , P2_U5864 );
and AND2_8042 ( P2_U3966 , P2_U5867 , P2_U5866 );
and AND2_8043 ( P2_U3967 , P2_U5871 , P2_U5870 );
and AND2_8044 ( P2_U3968 , P2_U5873 , P2_U5872 );
and AND2_8045 ( P2_U3969 , P2_U5875 , P2_U5874 );
and AND2_8046 ( P2_U3970 , P2_U5879 , P2_U5878 );
and AND2_8047 ( P2_U3971 , P2_U5881 , P2_U5880 );
and AND2_8048 ( P2_U3972 , P2_U5883 , P2_U5882 );
and AND2_8049 ( P2_U3973 , P2_U5887 , P2_U5886 );
and AND2_8050 ( P2_U3974 , P2_U5889 , P2_U5888 );
and AND2_8051 ( P2_U3975 , P2_U5891 , P2_U5890 );
and AND2_8052 ( P2_U3976 , P2_U5895 , P2_U5894 );
and AND2_8053 ( P2_U3977 , P2_U5897 , P2_U5896 );
and AND2_8054 ( P2_U3978 , P2_U5899 , P2_U5898 );
and AND2_8055 ( P2_U3979 , P2_U5903 , P2_U5902 );
and AND2_8056 ( P2_U3980 , P2_U5905 , P2_U5904 );
and AND2_8057 ( P2_U3981 , P2_U5907 , P2_U5906 );
and AND2_8058 ( P2_U3982 , P2_U5911 , P2_U5910 );
and AND4_8059 ( P2_U3983 , P2_U5915 , P2_U5914 , P2_U5913 , P2_U5912 );
and AND2_8060 ( P2_U3984 , P2_U5919 , P2_U5918 );
and AND3_8061 ( P2_U3985 , P2_U5923 , P2_U5922 , P2_U5921 );
and AND2_8062 ( P2_U3986 , P2_U5927 , P2_U5926 );
and AND3_8063 ( P2_U3987 , P2_U5931 , P2_U5930 , P2_U5929 );
and AND2_8064 ( P2_U3988 , P2_U5935 , P2_U5934 );
and AND2_8065 ( P2_U3989 , P2_STATE2_REG_1_ , P2_STATEBS16_REG );
nor nor_8066 ( P2_U3990 , P2_STATE2_REG_2_ , P2_STATE2_REG_1_ );
and AND3_8067 ( P2_U3991 , P2_U5942 , P2_U5941 , P2_U5943 );
and AND3_8068 ( P2_U3992 , P2_U5945 , P2_U5944 , P2_U5946 );
and AND3_8069 ( P2_U3993 , P2_U5948 , P2_U5947 , P2_U5949 );
and AND3_8070 ( P2_U3994 , P2_U5951 , P2_U5950 , P2_U5952 );
and AND3_8071 ( P2_U3995 , P2_U5954 , P2_U5953 , P2_U5955 );
and AND3_8072 ( P2_U3996 , P2_U5957 , P2_U5956 , P2_U5958 );
and AND3_8073 ( P2_U3997 , P2_U5960 , P2_U5959 , P2_U5961 );
and AND3_8074 ( P2_U3998 , P2_U5963 , P2_U5962 , P2_U5964 );
and AND3_8075 ( P2_U3999 , P2_U5966 , P2_U5965 , P2_U5967 );
and AND3_8076 ( P2_U4000 , P2_U5969 , P2_U5968 , P2_U5970 );
and AND3_8077 ( P2_U4001 , P2_U5972 , P2_U5971 , P2_U5973 );
and AND3_8078 ( P2_U4002 , P2_U5975 , P2_U5974 , P2_U5976 );
and AND3_8079 ( P2_U4003 , P2_U5978 , P2_U5977 , P2_U5979 );
and AND3_8080 ( P2_U4004 , P2_U5981 , P2_U5980 , P2_U5982 );
and AND3_8081 ( P2_U4005 , P2_U5984 , P2_U5983 , P2_U5985 );
and AND3_8082 ( P2_U4006 , P2_U5987 , P2_U5986 , P2_U5988 );
and AND3_8083 ( P2_U4007 , P2_U5990 , P2_U5989 , P2_U5991 );
and AND3_8084 ( P2_U4008 , P2_U5993 , P2_U5992 , P2_U5994 );
and AND3_8085 ( P2_U4009 , P2_U5996 , P2_U5995 , P2_U5997 );
and AND3_8086 ( P2_U4010 , P2_U5999 , P2_U5998 , P2_U6000 );
and AND3_8087 ( P2_U4011 , P2_U6002 , P2_U6001 , P2_U6003 );
and AND3_8088 ( P2_U4012 , P2_U6005 , P2_U6004 , P2_U6006 );
and AND3_8089 ( P2_U4013 , P2_U6008 , P2_U6007 , P2_U6009 );
and AND3_8090 ( P2_U4014 , P2_U6011 , P2_U6010 , P2_U6012 );
and AND3_8091 ( P2_U4015 , P2_U6014 , P2_U6013 , P2_U6015 );
and AND3_8092 ( P2_U4016 , P2_U6017 , P2_U6016 , P2_U6018 );
and AND3_8093 ( P2_U4017 , P2_U6020 , P2_U6019 , P2_U6021 );
and AND3_8094 ( P2_U4018 , P2_U6023 , P2_U6022 , P2_U6024 );
and AND3_8095 ( P2_U4019 , P2_U6026 , P2_U6025 , P2_U6027 );
and AND3_8096 ( P2_U4020 , P2_U6029 , P2_U6028 , P2_U6030 );
and AND3_8097 ( P2_U4021 , P2_U6032 , P2_U6031 , P2_U6033 );
and AND3_8098 ( P2_U4022 , P2_U6035 , P2_U6034 , P2_U6036 );
and AND3_8099 ( P2_U4023 , P2_U6038 , P2_U6037 , P2_U6039 );
and AND3_8100 ( P2_U4024 , P2_U6041 , P2_U6040 , P2_U6042 );
and AND3_8101 ( P2_U4025 , P2_U6044 , P2_U6043 , P2_U6045 );
and AND3_8102 ( P2_U4026 , P2_U6047 , P2_U6046 , P2_U6048 );
and AND3_8103 ( P2_U4027 , P2_U6050 , P2_U6049 , P2_U6051 );
and AND3_8104 ( P2_U4028 , P2_U6053 , P2_U6052 , P2_U6054 );
and AND3_8105 ( P2_U4029 , P2_U6056 , P2_U6055 , P2_U6057 );
and AND3_8106 ( P2_U4030 , P2_U6059 , P2_U6058 , P2_U6060 );
and AND3_8107 ( P2_U4031 , P2_U6062 , P2_U6061 , P2_U6063 );
and AND3_8108 ( P2_U4032 , P2_U6065 , P2_U6064 , P2_U6066 );
and AND3_8109 ( P2_U4033 , P2_U6068 , P2_U6067 , P2_U6069 );
and AND3_8110 ( P2_U4034 , P2_U6071 , P2_U6070 , P2_U6072 );
and AND3_8111 ( P2_U4035 , P2_U6074 , P2_U6073 , P2_U6075 );
and AND3_8112 ( P2_U4036 , P2_U6077 , P2_U6076 , P2_U6078 );
and AND3_8113 ( P2_U4037 , P2_U6080 , P2_U6079 , P2_U6081 );
and AND3_8114 ( P2_U4038 , P2_U6083 , P2_U6082 , P2_U6084 );
and AND3_8115 ( P2_U4039 , P2_U6086 , P2_U6085 , P2_U6087 );
and AND3_8116 ( P2_U4040 , P2_U6089 , P2_U6088 , P2_U6090 );
and AND3_8117 ( P2_U4041 , P2_U6092 , P2_U6091 , P2_U6093 );
and AND3_8118 ( P2_U4042 , P2_U6095 , P2_U6094 , P2_U6096 );
and AND3_8119 ( P2_U4043 , P2_U6098 , P2_U6097 , P2_U6099 );
and AND3_8120 ( P2_U4044 , P2_U6101 , P2_U6100 , P2_U6102 );
and AND3_8121 ( P2_U4045 , P2_U6104 , P2_U6103 , P2_U6105 );
and AND3_8122 ( P2_U4046 , P2_U6107 , P2_U6106 , P2_U6108 );
and AND3_8123 ( P2_U4047 , P2_U6110 , P2_U6109 , P2_U6111 );
and AND3_8124 ( P2_U4048 , P2_U6113 , P2_U6112 , P2_U6114 );
and AND3_8125 ( P2_U4049 , P2_U6116 , P2_U6115 , P2_U6117 );
and AND3_8126 ( P2_U4050 , P2_U6119 , P2_U6118 , P2_U6120 );
and AND3_8127 ( P2_U4051 , P2_U6122 , P2_U6121 , P2_U6123 );
and AND3_8128 ( P2_U4052 , P2_U6126 , P2_U6124 , P2_U6125 );
and AND3_8129 ( P2_U4053 , P2_U6128 , P2_U6127 , P2_U6129 );
and AND3_8130 ( P2_U4054 , P2_U6131 , P2_U6130 , P2_U6132 );
and AND3_8131 ( P2_U4055 , P2_U4468 , P2_U6133 , P2_U2356 );
and AND3_8132 ( P2_U4056 , P2_U3280 , P2_STATE2_REG_0_ , P2_U7871 );
and AND2_8133 ( P2_U4057 , P2_U2616 , P2_U4468 );
and AND2_8134 ( P2_U4058 , P2_U2374 , P2_U4417 );
and AND2_8135 ( P2_U4059 , P2_U6330 , P2_U6329 );
and AND2_8136 ( P2_U4060 , P2_U6334 , P2_U6333 );
and AND2_8137 ( P2_U4061 , P2_U6338 , P2_U6337 );
and AND2_8138 ( P2_U4062 , P2_U6342 , P2_U6341 );
and AND2_8139 ( P2_U4063 , P2_U6346 , P2_U6345 );
and AND2_8140 ( P2_U4064 , P2_U6350 , P2_U6349 );
and AND2_8141 ( P2_U4065 , P2_U6354 , P2_U6353 );
and AND2_8142 ( P2_U4066 , P2_U6358 , P2_U6357 );
and AND2_8143 ( P2_U4067 , P2_U6362 , P2_U6361 );
and AND2_8144 ( P2_U4068 , P2_U6366 , P2_U6365 );
and AND3_8145 ( P2_U4069 , P2_U4454 , P2_U4453 , P2_U6569 );
and AND3_8146 ( P2_U4070 , P2_U6574 , P2_U6573 , P2_U4071 );
and AND2_8147 ( P2_U4071 , P2_U6577 , P2_U6576 );
and AND2_8148 ( P2_U4072 , P2_U4073 , P2_U6578 );
and AND2_8149 ( P2_U4073 , P2_U6581 , P2_U6580 );
and AND3_8150 ( P2_U4074 , P2_U6583 , P2_U6582 , P2_U4075 );
and AND2_8151 ( P2_U4075 , P2_U6586 , P2_U6585 );
and AND2_8152 ( P2_U4076 , P2_U4077 , P2_U6587 );
and AND2_8153 ( P2_U4077 , P2_U6590 , P2_U6589 );
and AND3_8154 ( P2_U4078 , P2_U6592 , P2_U6591 , P2_U4079 );
and AND2_8155 ( P2_U4079 , P2_U6595 , P2_U6594 );
and AND2_8156 ( P2_U4080 , P2_U4081 , P2_U6596 );
and AND2_8157 ( P2_U4081 , P2_U6599 , P2_U6598 );
and AND3_8158 ( P2_U4082 , P2_U6601 , P2_U6600 , P2_U4083 );
and AND2_8159 ( P2_U4083 , P2_U6604 , P2_U6603 );
and AND2_8160 ( P2_U4084 , P2_U4085 , P2_U6605 );
and AND2_8161 ( P2_U4085 , P2_U6608 , P2_U6607 );
and AND3_8162 ( P2_U4086 , P2_U6609 , P2_U4446 , P2_U6610 );
and AND2_8163 ( P2_U4087 , P2_U4088 , P2_U6615 );
and AND2_8164 ( P2_U4088 , P2_U6617 , P2_U6616 );
and AND5_8165 ( P2_U4089 , P2_U6612 , P2_U6611 , P2_U4086 , P2_U6613 , P2_U6614 );
and AND3_8166 ( P2_U4090 , P2_U6618 , P2_U4446 , P2_U6619 );
and AND2_8167 ( P2_U4091 , P2_U4092 , P2_U6624 );
and AND2_8168 ( P2_U4092 , P2_U6626 , P2_U6625 );
and AND5_8169 ( P2_U4093 , P2_U6621 , P2_U6620 , P2_U4090 , P2_U6622 , P2_U6623 );
and AND3_8170 ( P2_U4094 , P2_U6627 , P2_U4446 , P2_U6628 );
and AND2_8171 ( P2_U4095 , P2_U4096 , P2_U6631 );
and AND2_8172 ( P2_U4096 , P2_U6634 , P2_U6633 );
and AND3_8173 ( P2_U4097 , P2_U6635 , P2_U4446 , P2_U6636 );
and AND2_8174 ( P2_U4098 , P2_U4099 , P2_U6639 );
and AND2_8175 ( P2_U4099 , P2_U6642 , P2_U6641 );
and AND3_8176 ( P2_U4100 , P2_U6643 , P2_U4446 , P2_U6644 );
and AND2_8177 ( P2_U4101 , P2_U4102 , P2_U6647 );
and AND2_8178 ( P2_U4102 , P2_U6650 , P2_U6649 );
and AND3_8179 ( P2_U4103 , P2_U6651 , P2_U4446 , P2_U6652 );
and AND2_8180 ( P2_U4104 , P2_U4105 , P2_U6655 );
and AND2_8181 ( P2_U4105 , P2_U6658 , P2_U6657 );
and AND3_8182 ( P2_U4106 , P2_U6659 , P2_U4446 , P2_U6660 );
and AND2_8183 ( P2_U4107 , P2_U4108 , P2_U6663 );
and AND2_8184 ( P2_U4108 , P2_U6666 , P2_U6665 );
and AND3_8185 ( P2_U4109 , P2_U6667 , P2_U4446 , P2_U6668 );
and AND2_8186 ( P2_U4110 , P2_U4111 , P2_U6671 );
and AND2_8187 ( P2_U4111 , P2_U6674 , P2_U6673 );
and AND3_8188 ( P2_U4112 , P2_U6675 , P2_U4446 , P2_U6678 );
and AND2_8189 ( P2_U4113 , P2_U4114 , P2_U6679 );
and AND2_8190 ( P2_U4114 , P2_U6682 , P2_U6681 );
and AND3_8191 ( P2_U4115 , P2_U6683 , P2_U4446 , P2_U6686 );
and AND2_8192 ( P2_U4116 , P2_U4117 , P2_U6687 );
and AND2_8193 ( P2_U4117 , P2_U6690 , P2_U6689 );
and AND3_8194 ( P2_U4118 , P2_U6691 , P2_U4446 , P2_U6694 );
and AND2_8195 ( P2_U4119 , P2_U4120 , P2_U6695 );
and AND2_8196 ( P2_U4120 , P2_U6698 , P2_U6697 );
and AND2_8197 ( P2_U4121 , P2_U6699 , P2_U4446 );
and AND2_8198 ( P2_U4122 , P2_U4123 , P2_U6703 );
and AND2_8199 ( P2_U4123 , P2_U6706 , P2_U6705 );
and AND5_8200 ( P2_U4124 , P2_U4121 , P2_U6701 , P2_U6702 , P2_U6700 , P2_U6704 );
and AND2_8201 ( P2_U4125 , P2_U6707 , P2_U4446 );
and AND2_8202 ( P2_U4126 , P2_U4127 , P2_U6711 );
and AND2_8203 ( P2_U4127 , P2_U6714 , P2_U6713 );
and AND5_8204 ( P2_U4128 , P2_U4125 , P2_U6709 , P2_U6710 , P2_U6708 , P2_U6712 );
and AND2_8205 ( P2_U4129 , P2_U6715 , P2_U4446 );
and AND2_8206 ( P2_U4130 , P2_U4131 , P2_U6719 );
and AND2_8207 ( P2_U4131 , P2_U6722 , P2_U6721 );
and AND5_8208 ( P2_U4132 , P2_U4129 , P2_U6717 , P2_U6718 , P2_U6716 , P2_U6720 );
and AND2_8209 ( P2_U4133 , P2_U6723 , P2_U4446 );
and AND2_8210 ( P2_U4134 , P2_U4135 , P2_U6727 );
and AND2_8211 ( P2_U4135 , P2_U6730 , P2_U6729 );
and AND5_8212 ( P2_U4136 , P2_U4133 , P2_U6725 , P2_U6726 , P2_U6724 , P2_U6728 );
and AND2_8213 ( P2_U4137 , P2_U6731 , P2_U4446 );
and AND2_8214 ( P2_U4138 , P2_U4139 , P2_U6735 );
and AND2_8215 ( P2_U4139 , P2_U6738 , P2_U6737 );
and AND5_8216 ( P2_U4140 , P2_U4137 , P2_U6733 , P2_U6734 , P2_U6732 , P2_U6736 );
and AND2_8217 ( P2_U4141 , P2_U4142 , P2_U6743 );
and AND2_8218 ( P2_U4142 , P2_U6746 , P2_U6745 );
and AND5_8219 ( P2_U4143 , P2_U6739 , P2_U6741 , P2_U6742 , P2_U6740 , P2_U6744 );
and AND2_8220 ( P2_U4144 , P2_U4145 , P2_U6751 );
and AND2_8221 ( P2_U4145 , P2_U6754 , P2_U6753 );
and AND5_8222 ( P2_U4146 , P2_U6747 , P2_U6749 , P2_U6750 , P2_U6748 , P2_U6752 );
and AND2_8223 ( P2_U4147 , P2_U6762 , P2_U6761 );
and AND3_8224 ( P2_U4148 , P2_U4147 , P2_U6759 , P2_U6760 );
and AND5_8225 ( P2_U4149 , P2_U6763 , P2_U6765 , P2_U6766 , P2_U6768 , P2_U4150 );
and AND2_8226 ( P2_U4150 , P2_U4151 , P2_U6767 );
and AND2_8227 ( P2_U4151 , P2_U6770 , P2_U6769 );
and AND5_8228 ( P2_U4152 , P2_U6771 , P2_U6773 , P2_U6774 , P2_U6776 , P2_U4153 );
and AND2_8229 ( P2_U4153 , P2_U4154 , P2_U6775 );
and AND2_8230 ( P2_U4154 , P2_U6778 , P2_U6777 );
and AND2_8231 ( P2_U4155 , P2_U6786 , P2_U6785 );
and AND3_8232 ( P2_U4156 , P2_U4155 , P2_U6783 , P2_U6784 );
and AND2_8233 ( P2_U4157 , P2_U6794 , P2_U6793 );
and AND3_8234 ( P2_U4158 , P2_U4157 , P2_U6791 , P2_U6792 );
and AND2_8235 ( P2_U4159 , P2_U6802 , P2_U6801 );
and AND3_8236 ( P2_U4160 , P2_U4159 , P2_U6799 , P2_U6800 );
and AND2_8237 ( P2_U4161 , P2_U6810 , P2_U6809 );
and AND3_8238 ( P2_U4162 , P2_U4161 , P2_U6807 , P2_U6808 );
and AND2_8239 ( P2_U4163 , P2_U6818 , P2_U6817 );
and AND3_8240 ( P2_U4164 , P2_U4163 , P2_U6815 , P2_U6816 );
and AND2_8241 ( P2_U4165 , P2_U6826 , P2_U6825 );
and AND3_8242 ( P2_U4166 , P2_U4165 , P2_U6823 , P2_U6824 );
and AND2_8243 ( P2_U4167 , P2_U6834 , P2_U6833 );
and AND3_8244 ( P2_U4168 , P2_U4167 , P2_U6831 , P2_U6832 );
nor nor_8245 ( P2_U4169 , P2_DATAWIDTH_REG_2_ , P2_DATAWIDTH_REG_3_ , P2_DATAWIDTH_REG_4_ , P2_DATAWIDTH_REG_5_ );
nor nor_8246 ( P2_U4170 , P2_DATAWIDTH_REG_6_ , P2_DATAWIDTH_REG_7_ , P2_DATAWIDTH_REG_8_ , P2_DATAWIDTH_REG_9_ );
and AND2_8247 ( P2_U4171 , P2_U4170 , P2_U4169 );
nor nor_8248 ( P2_U4172 , P2_DATAWIDTH_REG_10_ , P2_DATAWIDTH_REG_11_ , P2_DATAWIDTH_REG_12_ , P2_DATAWIDTH_REG_13_ );
nor nor_8249 ( P2_U4173 , P2_DATAWIDTH_REG_14_ , P2_DATAWIDTH_REG_15_ , P2_DATAWIDTH_REG_16_ , P2_DATAWIDTH_REG_17_ );
and AND2_8250 ( P2_U4174 , P2_U4173 , P2_U4172 );
nor nor_8251 ( P2_U4175 , P2_DATAWIDTH_REG_18_ , P2_DATAWIDTH_REG_19_ , P2_DATAWIDTH_REG_20_ , P2_DATAWIDTH_REG_21_ );
nor nor_8252 ( P2_U4176 , P2_DATAWIDTH_REG_22_ , P2_DATAWIDTH_REG_23_ , P2_DATAWIDTH_REG_24_ , P2_DATAWIDTH_REG_25_ );
and AND2_8253 ( P2_U4177 , P2_U4176 , P2_U4175 );
nor nor_8254 ( P2_U4178 , P2_DATAWIDTH_REG_26_ , P2_DATAWIDTH_REG_27_ );
nor nor_8255 ( P2_U4179 , P2_DATAWIDTH_REG_28_ , P2_DATAWIDTH_REG_29_ );
nor nor_8256 ( P2_U4180 , P2_DATAWIDTH_REG_30_ , P2_DATAWIDTH_REG_31_ );
and AND4_8257 ( P2_U4181 , P2_U4180 , P2_U6835 , P2_U4179 , P2_U4178 );
nor nor_8258 ( P2_U4182 , P2_DATAWIDTH_REG_1_ , P2_REIP_REG_0_ , P2_DATAWIDTH_REG_0_ );
nor nor_8259 ( P2_U4183 , P2_REIP_REG_1_ , P2_DATAWIDTH_REG_1_ );
and AND2_8260 ( P2_U4184 , P2_U6844 , P2_U7873 );
and AND2_8261 ( P2_U4185 , P2_U6848 , P2_U3301 );
and AND2_8262 ( P2_U4186 , P2_U4185 , P2_U6849 );
and AND2_8263 ( P2_U4187 , P2_STATE2_REG_1_ , P2_U3265 );
and AND3_8264 ( P2_U4188 , P2_U6842 , P2_U3313 , P2_U6841 );
and AND2_8265 ( P2_U4189 , P2_U2374 , P2_U3253 );
and AND2_8266 ( P2_U4190 , P2_U6860 , P2_U3534 );
and AND4_8267 ( P2_U4191 , P2_U6865 , P2_U6864 , P2_U6863 , P2_U6862 );
and AND4_8268 ( P2_U4192 , P2_U6869 , P2_U6868 , P2_U6867 , P2_U6866 );
and AND4_8269 ( P2_U4193 , P2_U6873 , P2_U6872 , P2_U6871 , P2_U6870 );
and AND4_8270 ( P2_U4194 , P2_U6877 , P2_U6876 , P2_U6875 , P2_U6874 );
and AND4_8271 ( P2_U4195 , P2_U6881 , P2_U6880 , P2_U6879 , P2_U6878 );
and AND4_8272 ( P2_U4196 , P2_U6885 , P2_U6884 , P2_U6883 , P2_U6882 );
and AND4_8273 ( P2_U4197 , P2_U6889 , P2_U6888 , P2_U6887 , P2_U6886 );
and AND4_8274 ( P2_U4198 , P2_U6893 , P2_U6892 , P2_U6891 , P2_U6890 );
and AND4_8275 ( P2_U4199 , P2_U6897 , P2_U6896 , P2_U6895 , P2_U6894 );
and AND4_8276 ( P2_U4200 , P2_U6901 , P2_U6900 , P2_U6899 , P2_U6898 );
and AND4_8277 ( P2_U4201 , P2_U6905 , P2_U6904 , P2_U6903 , P2_U6902 );
and AND4_8278 ( P2_U4202 , P2_U6909 , P2_U6908 , P2_U6907 , P2_U6906 );
and AND4_8279 ( P2_U4203 , P2_U6913 , P2_U6912 , P2_U6911 , P2_U6910 );
and AND4_8280 ( P2_U4204 , P2_U6917 , P2_U6916 , P2_U6915 , P2_U6914 );
and AND4_8281 ( P2_U4205 , P2_U6921 , P2_U6920 , P2_U6919 , P2_U6918 );
and AND4_8282 ( P2_U4206 , P2_U6925 , P2_U6924 , P2_U6923 , P2_U6922 );
and AND4_8283 ( P2_U4207 , P2_U6929 , P2_U6928 , P2_U6927 , P2_U6926 );
and AND4_8284 ( P2_U4208 , P2_U6933 , P2_U6932 , P2_U6931 , P2_U6930 );
and AND4_8285 ( P2_U4209 , P2_U6937 , P2_U6936 , P2_U6935 , P2_U6934 );
and AND4_8286 ( P2_U4210 , P2_U6941 , P2_U6940 , P2_U6939 , P2_U6938 );
and AND4_8287 ( P2_U4211 , P2_U6945 , P2_U6944 , P2_U6943 , P2_U6942 );
and AND4_8288 ( P2_U4212 , P2_U6949 , P2_U6948 , P2_U6947 , P2_U6946 );
and AND4_8289 ( P2_U4213 , P2_U6953 , P2_U6952 , P2_U6951 , P2_U6950 );
and AND4_8290 ( P2_U4214 , P2_U6957 , P2_U6956 , P2_U6955 , P2_U6954 );
and AND4_8291 ( P2_U4215 , P2_U6961 , P2_U6960 , P2_U6959 , P2_U6958 );
and AND4_8292 ( P2_U4216 , P2_U6965 , P2_U6964 , P2_U6963 , P2_U6962 );
and AND4_8293 ( P2_U4217 , P2_U6969 , P2_U6968 , P2_U6967 , P2_U6966 );
and AND4_8294 ( P2_U4218 , P2_U6973 , P2_U6972 , P2_U6971 , P2_U6970 );
and AND4_8295 ( P2_U4219 , P2_U6977 , P2_U6976 , P2_U6975 , P2_U6974 );
and AND4_8296 ( P2_U4220 , P2_U6981 , P2_U6980 , P2_U6979 , P2_U6978 );
and AND4_8297 ( P2_U4221 , P2_U6985 , P2_U6984 , P2_U6983 , P2_U6982 );
and AND4_8298 ( P2_U4222 , P2_U6989 , P2_U6988 , P2_U6987 , P2_U6986 );
and AND4_8299 ( P2_U4223 , P2_U6993 , P2_U6992 , P2_U6991 , P2_U6990 );
and AND4_8300 ( P2_U4224 , P2_U6997 , P2_U6996 , P2_U6995 , P2_U6994 );
and AND4_8301 ( P2_U4225 , P2_U7001 , P2_U7000 , P2_U6999 , P2_U6998 );
and AND4_8302 ( P2_U4226 , P2_U7005 , P2_U7004 , P2_U7003 , P2_U7002 );
and AND4_8303 ( P2_U4227 , P2_U7011 , P2_U7010 , P2_U7009 , P2_U7008 );
and AND4_8304 ( P2_U4228 , P2_U7015 , P2_U7014 , P2_U7013 , P2_U7012 );
and AND4_8305 ( P2_U4229 , P2_U7019 , P2_U7018 , P2_U7017 , P2_U7016 );
and AND4_8306 ( P2_U4230 , P2_U7023 , P2_U7022 , P2_U7021 , P2_U7020 );
and AND4_8307 ( P2_U4231 , P2_U7027 , P2_U7026 , P2_U7025 , P2_U7024 );
and AND4_8308 ( P2_U4232 , P2_U7031 , P2_U7030 , P2_U7029 , P2_U7028 );
and AND4_8309 ( P2_U4233 , P2_U7035 , P2_U7034 , P2_U7033 , P2_U7032 );
and AND4_8310 ( P2_U4234 , P2_U7039 , P2_U7038 , P2_U7037 , P2_U7036 );
and AND4_8311 ( P2_U4235 , P2_U7043 , P2_U7042 , P2_U7041 , P2_U7040 );
and AND4_8312 ( P2_U4236 , P2_U7047 , P2_U7046 , P2_U7045 , P2_U7044 );
and AND4_8313 ( P2_U4237 , P2_U7051 , P2_U7050 , P2_U7049 , P2_U7048 );
and AND4_8314 ( P2_U4238 , P2_U7055 , P2_U7054 , P2_U7053 , P2_U7052 );
and AND4_8315 ( P2_U4239 , P2_U7059 , P2_U7058 , P2_U7057 , P2_U7056 );
and AND4_8316 ( P2_U4240 , P2_U7063 , P2_U7062 , P2_U7061 , P2_U7060 );
and AND4_8317 ( P2_U4241 , P2_U7067 , P2_U7066 , P2_U7065 , P2_U7064 );
and AND4_8318 ( P2_U4242 , P2_U7071 , P2_U7070 , P2_U7069 , P2_U7068 );
and AND4_8319 ( P2_U4243 , P2_U7075 , P2_U7074 , P2_U7073 , P2_U7072 );
and AND4_8320 ( P2_U4244 , P2_U7079 , P2_U7078 , P2_U7077 , P2_U7076 );
and AND4_8321 ( P2_U4245 , P2_U7083 , P2_U7082 , P2_U7081 , P2_U7080 );
and AND4_8322 ( P2_U4246 , P2_U7087 , P2_U7086 , P2_U7085 , P2_U7084 );
and AND4_8323 ( P2_U4247 , P2_U7091 , P2_U7090 , P2_U7089 , P2_U7088 );
and AND4_8324 ( P2_U4248 , P2_U7095 , P2_U7094 , P2_U7093 , P2_U7092 );
and AND4_8325 ( P2_U4249 , P2_U7099 , P2_U7098 , P2_U7097 , P2_U7096 );
and AND4_8326 ( P2_U4250 , P2_U7103 , P2_U7102 , P2_U7101 , P2_U7100 );
and AND4_8327 ( P2_U4251 , P2_U7107 , P2_U7106 , P2_U7105 , P2_U7104 );
and AND4_8328 ( P2_U4252 , P2_U7111 , P2_U7110 , P2_U7109 , P2_U7108 );
and AND4_8329 ( P2_U4253 , P2_U7115 , P2_U7114 , P2_U7113 , P2_U7112 );
and AND4_8330 ( P2_U4254 , P2_U7119 , P2_U7118 , P2_U7117 , P2_U7116 );
and AND4_8331 ( P2_U4255 , P2_U7123 , P2_U7122 , P2_U7121 , P2_U7120 );
and AND4_8332 ( P2_U4256 , P2_U7127 , P2_U7126 , P2_U7125 , P2_U7124 );
and AND4_8333 ( P2_U4257 , P2_U7131 , P2_U7130 , P2_U7129 , P2_U7128 );
and AND4_8334 ( P2_U4258 , P2_U7135 , P2_U7134 , P2_U7133 , P2_U7132 );
and AND4_8335 ( P2_U4259 , P2_U7802 , P2_U7786 , P2_U7770 , P2_U7754 );
and AND4_8336 ( P2_U4260 , P2_U7874 , P2_U7850 , P2_U7834 , P2_U7818 );
and AND4_8337 ( P2_U4261 , P2_U7803 , P2_U7787 , P2_U7771 , P2_U7755 );
and AND4_8338 ( P2_U4262 , P2_U7875 , P2_U7851 , P2_U7835 , P2_U7819 );
and AND4_8339 ( P2_U4263 , P2_U7804 , P2_U7788 , P2_U7772 , P2_U7756 );
and AND4_8340 ( P2_U4264 , P2_U7876 , P2_U7852 , P2_U7836 , P2_U7820 );
and AND4_8341 ( P2_U4265 , P2_U7805 , P2_U7789 , P2_U7773 , P2_U7757 );
and AND4_8342 ( P2_U4266 , P2_U7877 , P2_U7853 , P2_U7837 , P2_U7821 );
and AND4_8343 ( P2_U4267 , P2_U7806 , P2_U7790 , P2_U7774 , P2_U7758 );
and AND4_8344 ( P2_U4268 , P2_U7878 , P2_U7854 , P2_U7838 , P2_U7822 );
and AND4_8345 ( P2_U4269 , P2_U7807 , P2_U7791 , P2_U7775 , P2_U7759 );
and AND4_8346 ( P2_U4270 , P2_U7879 , P2_U7855 , P2_U7839 , P2_U7823 );
and AND4_8347 ( P2_U4271 , P2_U7808 , P2_U7792 , P2_U7776 , P2_U7760 );
and AND4_8348 ( P2_U4272 , P2_U7880 , P2_U7856 , P2_U7840 , P2_U7824 );
and AND4_8349 ( P2_U4273 , P2_U7809 , P2_U7793 , P2_U7777 , P2_U7761 );
and AND4_8350 ( P2_U4274 , P2_U7881 , P2_U7857 , P2_U7841 , P2_U7825 );
and AND2_8351 ( P2_U4275 , P2_U7861 , P2_U4276 );
and AND3_8352 ( P2_U4276 , P2_STATE2_REG_2_ , P2_U3300 , P2_STATE2_REG_0_ );
and AND4_8353 ( P2_U4277 , P2_U7170 , P2_U7169 , P2_U7168 , P2_U7167 );
and AND4_8354 ( P2_U4278 , P2_U7174 , P2_U7173 , P2_U7172 , P2_U7171 );
and AND4_8355 ( P2_U4279 , P2_U7178 , P2_U7177 , P2_U7176 , P2_U7175 );
and AND4_8356 ( P2_U4280 , P2_U7182 , P2_U7181 , P2_U7180 , P2_U7179 );
and AND4_8357 ( P2_U4281 , P2_U7187 , P2_U7186 , P2_U7185 , P2_U7184 );
and AND4_8358 ( P2_U4282 , P2_U7191 , P2_U7190 , P2_U7189 , P2_U7188 );
and AND4_8359 ( P2_U4283 , P2_U7195 , P2_U7194 , P2_U7193 , P2_U7192 );
and AND4_8360 ( P2_U4284 , P2_U7199 , P2_U7198 , P2_U7197 , P2_U7196 );
and AND4_8361 ( P2_U4285 , P2_U7204 , P2_U7203 , P2_U7202 , P2_U7201 );
and AND4_8362 ( P2_U4286 , P2_U7208 , P2_U7207 , P2_U7206 , P2_U7205 );
and AND4_8363 ( P2_U4287 , P2_U7212 , P2_U7211 , P2_U7210 , P2_U7209 );
and AND4_8364 ( P2_U4288 , P2_U7216 , P2_U7215 , P2_U7214 , P2_U7213 );
and AND4_8365 ( P2_U4289 , P2_U7221 , P2_U7220 , P2_U7219 , P2_U7218 );
and AND4_8366 ( P2_U4290 , P2_U7225 , P2_U7224 , P2_U7223 , P2_U7222 );
and AND4_8367 ( P2_U4291 , P2_U7229 , P2_U7228 , P2_U7227 , P2_U7226 );
and AND4_8368 ( P2_U4292 , P2_U7233 , P2_U7232 , P2_U7231 , P2_U7230 );
and AND4_8369 ( P2_U4293 , P2_U7238 , P2_U7237 , P2_U7236 , P2_U7235 );
and AND4_8370 ( P2_U4294 , P2_U7242 , P2_U7241 , P2_U7240 , P2_U7239 );
and AND4_8371 ( P2_U4295 , P2_U7246 , P2_U7245 , P2_U7244 , P2_U7243 );
and AND4_8372 ( P2_U4296 , P2_U7250 , P2_U7249 , P2_U7248 , P2_U7247 );
and AND4_8373 ( P2_U4297 , P2_U7255 , P2_U7254 , P2_U7253 , P2_U7252 );
and AND4_8374 ( P2_U4298 , P2_U7259 , P2_U7258 , P2_U7257 , P2_U7256 );
and AND4_8375 ( P2_U4299 , P2_U7263 , P2_U7262 , P2_U7261 , P2_U7260 );
and AND4_8376 ( P2_U4300 , P2_U7267 , P2_U7266 , P2_U7265 , P2_U7264 );
and AND4_8377 ( P2_U4301 , P2_U7272 , P2_U7271 , P2_U7270 , P2_U7269 );
and AND4_8378 ( P2_U4302 , P2_U7276 , P2_U7275 , P2_U7274 , P2_U7273 );
and AND4_8379 ( P2_U4303 , P2_U7280 , P2_U7279 , P2_U7278 , P2_U7277 );
and AND4_8380 ( P2_U4304 , P2_U7284 , P2_U7283 , P2_U7282 , P2_U7281 );
and AND4_8381 ( P2_U4305 , P2_U7289 , P2_U7288 , P2_U7287 , P2_U7286 );
and AND4_8382 ( P2_U4306 , P2_U7293 , P2_U7292 , P2_U7291 , P2_U7290 );
and AND4_8383 ( P2_U4307 , P2_U7297 , P2_U7296 , P2_U7295 , P2_U7294 );
and AND4_8384 ( P2_U4308 , P2_U7301 , P2_U7300 , P2_U7299 , P2_U7298 );
and AND4_8385 ( P2_U4309 , P2_U7306 , P2_U7305 , P2_U7304 , P2_U7303 );
and AND4_8386 ( P2_U4310 , P2_U7310 , P2_U7309 , P2_U7308 , P2_U7307 );
and AND4_8387 ( P2_U4311 , P2_U7314 , P2_U7313 , P2_U7312 , P2_U7311 );
and AND4_8388 ( P2_U4312 , P2_U7318 , P2_U7317 , P2_U7316 , P2_U7315 );
and AND4_8389 ( P2_U4313 , P2_U7323 , P2_U7322 , P2_U7321 , P2_U7320 );
and AND4_8390 ( P2_U4314 , P2_U7327 , P2_U7326 , P2_U7325 , P2_U7324 );
and AND4_8391 ( P2_U4315 , P2_U7331 , P2_U7330 , P2_U7329 , P2_U7328 );
and AND4_8392 ( P2_U4316 , P2_U7335 , P2_U7334 , P2_U7333 , P2_U7332 );
and AND4_8393 ( P2_U4317 , P2_U7340 , P2_U7339 , P2_U7338 , P2_U7337 );
and AND4_8394 ( P2_U4318 , P2_U7344 , P2_U7343 , P2_U7342 , P2_U7341 );
and AND4_8395 ( P2_U4319 , P2_U7348 , P2_U7347 , P2_U7346 , P2_U7345 );
and AND4_8396 ( P2_U4320 , P2_U7352 , P2_U7351 , P2_U7350 , P2_U7349 );
and AND4_8397 ( P2_U4321 , P2_U7357 , P2_U7356 , P2_U7355 , P2_U7354 );
and AND4_8398 ( P2_U4322 , P2_U7361 , P2_U7360 , P2_U7359 , P2_U7358 );
and AND4_8399 ( P2_U4323 , P2_U7365 , P2_U7364 , P2_U7363 , P2_U7362 );
and AND4_8400 ( P2_U4324 , P2_U7369 , P2_U7368 , P2_U7367 , P2_U7366 );
and AND4_8401 ( P2_U4325 , P2_U7374 , P2_U7373 , P2_U7372 , P2_U7371 );
and AND4_8402 ( P2_U4326 , P2_U7378 , P2_U7377 , P2_U7376 , P2_U7375 );
and AND4_8403 ( P2_U4327 , P2_U7382 , P2_U7381 , P2_U7380 , P2_U7379 );
and AND4_8404 ( P2_U4328 , P2_U7386 , P2_U7385 , P2_U7384 , P2_U7383 );
and AND4_8405 ( P2_U4329 , P2_U7391 , P2_U7390 , P2_U7389 , P2_U7388 );
and AND4_8406 ( P2_U4330 , P2_U7395 , P2_U7394 , P2_U7393 , P2_U7392 );
and AND4_8407 ( P2_U4331 , P2_U7399 , P2_U7398 , P2_U7397 , P2_U7396 );
and AND4_8408 ( P2_U4332 , P2_U7403 , P2_U7402 , P2_U7401 , P2_U7400 );
and AND4_8409 ( P2_U4333 , P2_U7408 , P2_U7407 , P2_U7406 , P2_U7405 );
and AND4_8410 ( P2_U4334 , P2_U7412 , P2_U7411 , P2_U7410 , P2_U7409 );
and AND4_8411 ( P2_U4335 , P2_U7416 , P2_U7415 , P2_U7414 , P2_U7413 );
and AND4_8412 ( P2_U4336 , P2_U7420 , P2_U7419 , P2_U7418 , P2_U7417 );
and AND2_8413 ( P2_U4337 , P2_U2616 , P2_U3300 );
and AND2_8414 ( P2_U4338 , P2_U7425 , P2_U4413 );
and AND2_8415 ( P2_U4339 , P2_U4595 , P2_U3300 );
and AND3_8416 ( P2_U4340 , P2_U7426 , P2_U4414 , P2_U7428 );
and AND2_8417 ( P2_U4341 , P2_U7430 , P2_U3571 );
and AND2_8418 ( P2_U4342 , P2_U4413 , P2_U4341 );
and AND2_8419 ( P2_U4343 , P2_U7869 , P2_U7873 );
and AND2_8420 ( P2_U4344 , P2_U7436 , P2_U7435 );
and AND2_8421 ( P2_U4345 , P2_U7440 , P2_U7439 );
and AND2_8422 ( P2_U4346 , P2_U7442 , P2_U7443 );
and AND2_8423 ( P2_U4347 , P2_U7445 , P2_U7446 );
and AND2_8424 ( P2_U4348 , P2_U7448 , P2_U7449 );
and AND2_8425 ( P2_U4349 , P2_U7451 , P2_U7452 );
and AND2_8426 ( P2_U4350 , P2_U7454 , P2_U7455 );
and AND2_8427 ( P2_U4351 , P2_U7457 , P2_U7458 );
and AND2_8428 ( P2_U4352 , P2_U7460 , P2_U7461 );
and AND2_8429 ( P2_U4353 , P2_U7463 , P2_U7464 );
and AND2_8430 ( P2_U4354 , P2_U7466 , P2_U7467 );
and AND2_8431 ( P2_U4355 , P2_U7469 , P2_U7470 );
and AND2_8432 ( P2_U4356 , P2_U7472 , P2_U7473 );
and AND2_8433 ( P2_U4357 , P2_U7475 , P2_U7476 );
and AND2_8434 ( P2_U4358 , P2_U7478 , P2_U7479 );
and AND2_8435 ( P2_U4359 , P2_U7481 , P2_U7482 );
and AND2_8436 ( P2_U4360 , P2_U7484 , P2_U7485 );
and AND2_8437 ( P2_U4361 , P2_U7487 , P2_U7488 );
and AND2_8438 ( P2_U4362 , P2_U7490 , P2_U7491 );
and AND2_8439 ( P2_U4363 , P2_U7493 , P2_U7494 );
and AND2_8440 ( P2_U4364 , P2_U7496 , P2_U7497 );
and AND2_8441 ( P2_U4365 , P2_U7499 , P2_U7500 );
and AND2_8442 ( P2_U4366 , P2_U7502 , P2_U7503 );
and AND2_8443 ( P2_U4367 , P2_U7505 , P2_U7506 );
and AND2_8444 ( P2_U4368 , P2_U7510 , P2_U7509 );
and AND2_8445 ( P2_U4369 , P2_U7514 , P2_U7513 );
and AND2_8446 ( P2_U4370 , P2_U7518 , P2_U7517 );
and AND2_8447 ( P2_U4371 , P2_U7522 , P2_U7521 );
and AND2_8448 ( P2_U4372 , P2_U7526 , P2_U7525 );
and AND2_8449 ( P2_U4373 , P2_U7530 , P2_U7529 );
and AND2_8450 ( P2_U4374 , P2_U7532 , P2_U7533 );
and AND2_8451 ( P2_U4375 , P2_U7536 , P2_U7535 );
and AND2_8452 ( P2_U4376 , P2_U3255 , P2_U6845 );
and AND2_8453 ( P2_U4377 , P2_U7863 , P2_U3255 );
and AND2_8454 ( P2_U4378 , P2_U2356 , P2_U7873 );
and AND3_8455 ( P2_U4379 , P2_U7579 , P2_U7580 , P2_U7578 );
and AND2_8456 ( P2_U4380 , P2_U7585 , P2_U3269 );
and AND2_8457 ( P2_U4381 , P2_U2356 , P2_U4595 );
and AND5_8458 ( P2_U4382 , P2_U3577 , P2_U3539 , P2_U4472 , P2_U7587 , P2_U7586 );
and AND2_8459 ( P2_U4383 , P2_U7579 , P2_U4422 );
and AND2_8460 ( P2_U4384 , P2_U4383 , P2_U7578 );
and AND2_8461 ( P2_U4385 , P2_U7580 , P2_U4458 );
and AND2_8462 ( P2_U4386 , P2_U7590 , P2_U7589 );
and AND2_8463 ( P2_U4387 , P2_STATE2_REG_0_ , P2_U7736 );
and AND4_8464 ( P2_U4388 , P2_U3573 , P2_U4458 , P2_U4457 , P2_U3549 );
and AND2_8465 ( P2_U4389 , P2_U7719 , P2_U7718 );
and AND2_8466 ( P2_U4390 , P2_U7731 , P2_U3536 );
and AND2_8467 ( P2_U4391 , P2_U7735 , P2_U3536 );
and AND2_8468 ( P2_U4392 , P2_U7908 , P2_U7907 );
and AND2_8469 ( P2_U4393 , P2_U8055 , P2_U8054 );
nand NAND2_8470 ( P2_U4394 , P2_U3872 , P2_U5582 );
and AND2_8471 ( P2_U4395 , P2_U8079 , P2_U8078 );
and AND2_8472 ( P2_U4396 , P2_U8092 , P2_U8091 );
and AND2_8473 ( P2_U4397 , P2_U8120 , P2_U8119 );
and AND2_8474 ( P2_U4398 , P2_U8126 , P2_U8125 );
and AND2_8475 ( P2_U4399 , P2_U8132 , P2_U8131 );
nand NAND2_8476 ( P2_U4400 , P2_U2374 , P2_U3291 );
not NOT1_8477 ( P2_U4401 , BS16 );
nand NAND2_8478 ( P2_U4402 , P2_U4462 , P2_U4188 );
nand NAND2_8479 ( P2_U4403 , P2_U3534 , P2_U4462 );
and AND2_8480 ( P2_U4404 , P2_U8146 , P2_U8145 );
nand NAND2_8481 ( P2_U4405 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_U7006 );
nand NAND2_8482 ( P2_U4406 , P2_U2513 , P2_U3871 );
not NOT1_8483 ( P2_U4407 , P2_R2219_U29 );
not NOT1_8484 ( P2_U4408 , P2_R2219_U8 );
not NOT1_8485 ( P2_U4409 , P2_U3553 );
nand NAND2_8486 ( P2_U4410 , HOLD , P2_U3265 );
not NOT1_8487 ( P2_U4411 , P2_U3290 );
not NOT1_8488 ( P2_U4412 , P2_U3571 );
nand NAND2_8489 ( P2_U4413 , P2_U4337 , P2_U4601 );
nand NAND3_8490 ( P2_U4414 , P2_U2616 , P2_U3300 , P2_U7869 );
nand NAND2_8491 ( P2_U4415 , P2_U2447 , P2_U3279 );
not NOT1_8492 ( P2_U4416 , P2_U3576 );
not NOT1_8493 ( P2_U4417 , P2_U3283 );
not NOT1_8494 ( P2_U4418 , P2_U3550 );
not NOT1_8495 ( P2_U4419 , P2_U3536 );
not NOT1_8496 ( P2_U4420 , P2_U3288 );
not NOT1_8497 ( P2_U4421 , P2_U3539 );
nand NAND3_8498 ( P2_U4422 , P2_U2376 , P2_U3278 , P2_U2450 );
not NOT1_8499 ( P2_U4423 , P2_U3577 );
not NOT1_8500 ( P2_U4424 , P2_U3282 );
not NOT1_8501 ( P2_U4425 , P2_U3285 );
not NOT1_8502 ( P2_U4426 , P2_U3549 );
not NOT1_8503 ( P2_U4427 , P2_U3289 );
not NOT1_8504 ( P2_U4428 , P2_U3286 );
not NOT1_8505 ( P2_U4429 , P2_U3294 );
not NOT1_8506 ( P2_U4430 , P2_U3313 );
not NOT1_8507 ( P2_U4431 , P2_U3578 );
not NOT1_8508 ( P2_U4432 , P2_U3254 );
not NOT1_8509 ( P2_U4433 , P2_U3523 );
not NOT1_8510 ( P2_U4434 , P2_U3524 );
not NOT1_8511 ( P2_U4435 , P2_U3296 );
not NOT1_8512 ( P2_U4436 , P2_U3522 );
nand NAND2_8513 ( P2_U4437 , P2_U3875 , P2_U2376 );
not NOT1_8514 ( P2_U4438 , P2_U3547 );
not NOT1_8515 ( P2_U4439 , P2_U3259 );
not NOT1_8516 ( P2_U4440 , P2_U3543 );
not NOT1_8517 ( P2_U4441 , P2_U3542 );
not NOT1_8518 ( P2_U4442 , P2_U3538 );
not NOT1_8519 ( P2_U4443 , P2_U3306 );
not NOT1_8520 ( P2_U4444 , P2_LT_563_1260_U6 );
nand NAND2_8521 ( P2_U4445 , P2_U4430 , P2_U3302 );
nand NAND2_8522 ( P2_U4446 , P2_U4461 , P2_U3546 );
nand NAND2_8523 ( P2_U4447 , P2_R2219_U7 , P2_U2617 );
nand NAND2_8524 ( P2_U4448 , P2_U2367 , P2_U3290 );
not NOT1_8525 ( P2_U4449 , P2_U3261 );
not NOT1_8526 ( P2_U4450 , P2_U3260 );
not NOT1_8527 ( P2_U4451 , P2_U3425 );
nand NAND2_8528 ( P2_U4452 , P2_U4182 , P2_U4438 );
nand NAND2_8529 ( P2_U4453 , P2_U3718 , P2_U4474 );
nand NAND4_8530 ( P2_U4454 , P2_STATE2_REG_1_ , P2_U3302 , P2_U3270 , P2_U3284 );
nand NAND2_8531 ( P2_U4455 , P2_U3867 , P2_U2448 );
nand NAND2_8532 ( P2_U4456 , P2_U2446 , P2_U2359 );
nand NAND2_8533 ( P2_U4457 , P2_U2356 , P2_U3280 );
nand NAND2_8534 ( P2_U4458 , P2_U4378 , P2_U7577 );
not NOT1_8535 ( P2_U4459 , P2_U3575 );
nand NAND2_8536 ( P2_U4460 , P2_U2438 , P2_U3295 );
not NOT1_8537 ( P2_U4461 , P2_U3534 );
nand NAND2_8538 ( P2_U4462 , P2_U2374 , P2_U6568 );
nand NAND2_8539 ( P2_U4463 , P2_U4574 , P2_U3266 );
nand NAND2_8540 ( P2_U4464 , P2_U2448 , P2_U3292 );
nand NAND2_8541 ( P2_U4465 , P2_U4474 , U211 );
not NOT1_8542 ( P2_U4466 , P2_U3303 );
not NOT1_8543 ( P2_U4467 , P2_U3540 );
not NOT1_8544 ( P2_U4468 , P2_U3304 );
not NOT1_8545 ( P2_U4469 , P2_U3305 );
nand NAND2_8546 ( P2_U4470 , P2_U3876 , P2_U2376 );
not NOT1_8547 ( P2_U4471 , P2_U3573 );
nand NAND3_8548 ( P2_U4472 , P2_U2376 , P2_U7871 , P2_U4416 );
not NOT1_8549 ( P2_U4473 , P2_U3262 );
not NOT1_8550 ( P2_U4474 , P2_U3301 );
not NOT1_8551 ( P2_U4475 , P2_U3293 );
not NOT1_8552 ( P2_U4476 , P2_U3281 );
not NOT1_8553 ( P2_U4477 , P2_U3548 );
nand NAND2_8554 ( P2_U4478 , P2_REIP_REG_31_ , P2_U4450 );
nand NAND2_8555 ( P2_U4479 , P2_REIP_REG_30_ , P2_U4449 );
nand NAND2_8556 ( P2_U4480 , P2_ADDRESS_REG_29_ , P2_U3259 );
nand NAND2_8557 ( P2_U4481 , P2_REIP_REG_30_ , P2_U4450 );
nand NAND2_8558 ( P2_U4482 , P2_REIP_REG_29_ , P2_U4449 );
nand NAND2_8559 ( P2_U4483 , P2_ADDRESS_REG_28_ , P2_U3259 );
nand NAND2_8560 ( P2_U4484 , P2_REIP_REG_29_ , P2_U4450 );
nand NAND2_8561 ( P2_U4485 , P2_REIP_REG_28_ , P2_U4449 );
nand NAND2_8562 ( P2_U4486 , P2_ADDRESS_REG_27_ , P2_U3259 );
nand NAND2_8563 ( P2_U4487 , P2_REIP_REG_28_ , P2_U4450 );
nand NAND2_8564 ( P2_U4488 , P2_REIP_REG_27_ , P2_U4449 );
nand NAND2_8565 ( P2_U4489 , P2_ADDRESS_REG_26_ , P2_U3259 );
nand NAND2_8566 ( P2_U4490 , P2_REIP_REG_27_ , P2_U4450 );
nand NAND2_8567 ( P2_U4491 , P2_REIP_REG_26_ , P2_U4449 );
nand NAND2_8568 ( P2_U4492 , P2_ADDRESS_REG_25_ , P2_U3259 );
nand NAND2_8569 ( P2_U4493 , P2_REIP_REG_26_ , P2_U4450 );
nand NAND2_8570 ( P2_U4494 , P2_REIP_REG_25_ , P2_U4449 );
nand NAND2_8571 ( P2_U4495 , P2_ADDRESS_REG_24_ , P2_U3259 );
nand NAND2_8572 ( P2_U4496 , P2_REIP_REG_25_ , P2_U4450 );
nand NAND2_8573 ( P2_U4497 , P2_REIP_REG_24_ , P2_U4449 );
nand NAND2_8574 ( P2_U4498 , P2_ADDRESS_REG_23_ , P2_U3259 );
nand NAND2_8575 ( P2_U4499 , P2_REIP_REG_24_ , P2_U4450 );
nand NAND2_8576 ( P2_U4500 , P2_REIP_REG_23_ , P2_U4449 );
nand NAND2_8577 ( P2_U4501 , P2_ADDRESS_REG_22_ , P2_U3259 );
nand NAND2_8578 ( P2_U4502 , P2_REIP_REG_23_ , P2_U4450 );
nand NAND2_8579 ( P2_U4503 , P2_REIP_REG_22_ , P2_U4449 );
nand NAND2_8580 ( P2_U4504 , P2_ADDRESS_REG_21_ , P2_U3259 );
nand NAND2_8581 ( P2_U4505 , P2_REIP_REG_22_ , P2_U4450 );
nand NAND2_8582 ( P2_U4506 , P2_REIP_REG_21_ , P2_U4449 );
nand NAND2_8583 ( P2_U4507 , P2_ADDRESS_REG_20_ , P2_U3259 );
nand NAND2_8584 ( P2_U4508 , P2_REIP_REG_21_ , P2_U4450 );
nand NAND2_8585 ( P2_U4509 , P2_REIP_REG_20_ , P2_U4449 );
nand NAND2_8586 ( P2_U4510 , P2_ADDRESS_REG_19_ , P2_U3259 );
nand NAND2_8587 ( P2_U4511 , P2_REIP_REG_20_ , P2_U4450 );
nand NAND2_8588 ( P2_U4512 , P2_REIP_REG_19_ , P2_U4449 );
nand NAND2_8589 ( P2_U4513 , P2_ADDRESS_REG_18_ , P2_U3259 );
nand NAND2_8590 ( P2_U4514 , P2_REIP_REG_19_ , P2_U4450 );
nand NAND2_8591 ( P2_U4515 , P2_REIP_REG_18_ , P2_U4449 );
nand NAND2_8592 ( P2_U4516 , P2_ADDRESS_REG_17_ , P2_U3259 );
nand NAND2_8593 ( P2_U4517 , P2_REIP_REG_18_ , P2_U4450 );
nand NAND2_8594 ( P2_U4518 , P2_REIP_REG_17_ , P2_U4449 );
nand NAND2_8595 ( P2_U4519 , P2_ADDRESS_REG_16_ , P2_U3259 );
nand NAND2_8596 ( P2_U4520 , P2_REIP_REG_17_ , P2_U4450 );
nand NAND2_8597 ( P2_U4521 , P2_REIP_REG_16_ , P2_U4449 );
nand NAND2_8598 ( P2_U4522 , P2_ADDRESS_REG_15_ , P2_U3259 );
nand NAND2_8599 ( P2_U4523 , P2_REIP_REG_16_ , P2_U4450 );
nand NAND2_8600 ( P2_U4524 , P2_REIP_REG_15_ , P2_U4449 );
nand NAND2_8601 ( P2_U4525 , P2_ADDRESS_REG_14_ , P2_U3259 );
nand NAND2_8602 ( P2_U4526 , P2_REIP_REG_15_ , P2_U4450 );
nand NAND2_8603 ( P2_U4527 , P2_REIP_REG_14_ , P2_U4449 );
nand NAND2_8604 ( P2_U4528 , P2_ADDRESS_REG_13_ , P2_U3259 );
nand NAND2_8605 ( P2_U4529 , P2_REIP_REG_14_ , P2_U4450 );
nand NAND2_8606 ( P2_U4530 , P2_REIP_REG_13_ , P2_U4449 );
nand NAND2_8607 ( P2_U4531 , P2_ADDRESS_REG_12_ , P2_U3259 );
nand NAND2_8608 ( P2_U4532 , P2_REIP_REG_13_ , P2_U4450 );
nand NAND2_8609 ( P2_U4533 , P2_REIP_REG_12_ , P2_U4449 );
nand NAND2_8610 ( P2_U4534 , P2_ADDRESS_REG_11_ , P2_U3259 );
nand NAND2_8611 ( P2_U4535 , P2_REIP_REG_12_ , P2_U4450 );
nand NAND2_8612 ( P2_U4536 , P2_REIP_REG_11_ , P2_U4449 );
nand NAND2_8613 ( P2_U4537 , P2_ADDRESS_REG_10_ , P2_U3259 );
nand NAND2_8614 ( P2_U4538 , P2_REIP_REG_11_ , P2_U4450 );
nand NAND2_8615 ( P2_U4539 , P2_REIP_REG_10_ , P2_U4449 );
nand NAND2_8616 ( P2_U4540 , P2_ADDRESS_REG_9_ , P2_U3259 );
nand NAND2_8617 ( P2_U4541 , P2_REIP_REG_10_ , P2_U4450 );
nand NAND2_8618 ( P2_U4542 , P2_REIP_REG_9_ , P2_U4449 );
nand NAND2_8619 ( P2_U4543 , P2_ADDRESS_REG_8_ , P2_U3259 );
nand NAND2_8620 ( P2_U4544 , P2_REIP_REG_9_ , P2_U4450 );
nand NAND2_8621 ( P2_U4545 , P2_REIP_REG_8_ , P2_U4449 );
nand NAND2_8622 ( P2_U4546 , P2_ADDRESS_REG_7_ , P2_U3259 );
nand NAND2_8623 ( P2_U4547 , P2_REIP_REG_8_ , P2_U4450 );
nand NAND2_8624 ( P2_U4548 , P2_REIP_REG_7_ , P2_U4449 );
nand NAND2_8625 ( P2_U4549 , P2_ADDRESS_REG_6_ , P2_U3259 );
nand NAND2_8626 ( P2_U4550 , P2_REIP_REG_7_ , P2_U4450 );
nand NAND2_8627 ( P2_U4551 , P2_REIP_REG_6_ , P2_U4449 );
nand NAND2_8628 ( P2_U4552 , P2_ADDRESS_REG_5_ , P2_U3259 );
nand NAND2_8629 ( P2_U4553 , P2_REIP_REG_6_ , P2_U4450 );
nand NAND2_8630 ( P2_U4554 , P2_REIP_REG_5_ , P2_U4449 );
nand NAND2_8631 ( P2_U4555 , P2_ADDRESS_REG_4_ , P2_U3259 );
nand NAND2_8632 ( P2_U4556 , P2_REIP_REG_5_ , P2_U4450 );
nand NAND2_8633 ( P2_U4557 , P2_REIP_REG_4_ , P2_U4449 );
nand NAND2_8634 ( P2_U4558 , P2_ADDRESS_REG_3_ , P2_U3259 );
nand NAND2_8635 ( P2_U4559 , P2_REIP_REG_4_ , P2_U4450 );
nand NAND2_8636 ( P2_U4560 , P2_REIP_REG_3_ , P2_U4449 );
nand NAND2_8637 ( P2_U4561 , P2_ADDRESS_REG_2_ , P2_U3259 );
nand NAND2_8638 ( P2_U4562 , P2_REIP_REG_3_ , P2_U4450 );
nand NAND2_8639 ( P2_U4563 , P2_REIP_REG_2_ , P2_U4449 );
nand NAND2_8640 ( P2_U4564 , P2_ADDRESS_REG_1_ , P2_U3259 );
nand NAND2_8641 ( P2_U4565 , P2_REIP_REG_2_ , P2_U4450 );
nand NAND2_8642 ( P2_U4566 , P2_REIP_REG_1_ , P2_U4449 );
nand NAND2_8643 ( P2_U4567 , P2_ADDRESS_REG_0_ , P2_U3259 );
not NOT1_8644 ( P2_U4568 , P2_U3267 );
nand NAND2_8645 ( P2_U4569 , P2_U4568 , P2_U3265 );
nand NAND2_8646 ( P2_U4570 , NA , P2_U4473 );
not NOT1_8647 ( P2_U4571 , P2_U3268 );
nand NAND2_8648 ( P2_U4572 , P2_U4571 , P2_U3265 );
nand NAND2_8649 ( P2_U4573 , P2_U4392 , P2_U7891 );
not NOT1_8650 ( P2_U4574 , P2_U3263 );
nand NAND3_8651 ( P2_U4575 , HOLD , P2_U3256 , P2_U4574 );
nand NAND3_8652 ( P2_U4576 , P2_STATE_REG_1_ , P2_U3268 , U211 );
nand NAND2_8653 ( P2_U4577 , P2_U4576 , P2_U4575 );
nand NAND3_8654 ( P2_U4578 , P2_STATE_REG_0_ , P2_U4570 , P2_U4577 );
nand NAND2_8655 ( P2_U4579 , P2_STATE_REG_2_ , P2_U4573 );
nand NAND2_8656 ( P2_U4580 , P2_STATE_REG_0_ , P2_U4410 );
nand NAND2_8657 ( P2_U4581 , P2_U4580 , P2_STATE_REG_2_ );
nand NAND3_8658 ( P2_U4582 , P2_U7910 , P2_U7909 , P2_U7892 );
nand NAND2_8659 ( P2_U4583 , U211 , P2_U4439 );
nand NAND2_8660 ( P2_U4584 , P2_U3692 , P2_U7893 );
nand NAND2_8661 ( P2_U4585 , P2_STATE_REG_2_ , P2_U3267 );
nand NAND2_8662 ( P2_U4586 , NA , P2_U3266 );
nand NAND2_8663 ( P2_U4587 , P2_U4586 , P2_U4585 );
nand NAND2_8664 ( P2_U4588 , P2_U4587 , P2_U3258 );
nand NAND2_8665 ( P2_U4589 , P2_U4401 , P2_U3263 );
not NOT1_8666 ( P2_U4590 , P2_U3277 );
nand NAND2_8667 ( P2_U4591 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_8668 ( P2_U4592 , P2_U3274 );
not NOT1_8669 ( P2_U4593 , P2_U3275 );
nand NAND2_8670 ( P2_U4594 , P2_STATE_REG_2_ , P2_U3258 );
nand NAND2_8671 ( P2_U4595 , P2_U3262 , P2_U4594 );
not NOT1_8672 ( P2_U4596 , P2_U3527 );
nand NAND2_8673 ( P2_U4597 , P2_U3294 , P2_U3286 );
nand NAND2_8674 ( P2_U4598 , P2_U4597 , P2_U3265 );
nand NAND2_8675 ( P2_U4599 , P2_U2359 , P2_U3527 );
not NOT1_8676 ( P2_U4600 , P2_U3291 );
not NOT1_8677 ( P2_U4601 , P2_U3295 );
nand NAND2_8678 ( P2_U4602 , P2_U4424 , P2_U3253 );
nand NAND2_8679 ( P2_U4603 , P2_U3524 , P2_U4602 );
nand NAND2_8680 ( P2_U4604 , P2_U3523 , P2_U3522 );
nand NAND2_8681 ( P2_U4605 , P2_R2243_U8 , P2_U4428 );
nand NAND2_8682 ( P2_U4606 , P2_U4417 , P2_U3287 );
nand NAND2_8683 ( P2_U4607 , P2_U4606 , P2_U4605 );
nand NAND2_8684 ( P2_U4608 , P2_U4420 , P2_U4607 );
nand NAND2_8685 ( P2_U4609 , P2_U4603 , P2_U3520 );
not NOT1_8686 ( P2_U4610 , P2_U3257 );
nand NAND2_8687 ( P2_U4611 , P2_U4428 , P2_U3292 );
nand NAND2_8688 ( P2_U4612 , P2_GTE_370_U6 , P2_U4417 );
nand NAND2_8689 ( P2_U4613 , P2_U4612 , P2_U4611 );
nand NAND2_8690 ( P2_U4614 , P2_U4420 , P2_U4613 );
or OR2_8691 ( P2_U4615 , P2_MORE_REG , P2_FLUSH_REG );
not NOT1_8692 ( P2_U4616 , P2_U3298 );
nand NAND2_8693 ( P2_U4617 , P2_U4616 , P2_U3269 );
nand NAND2_8694 ( P2_U4618 , P2_U3711 , P2_U4425 );
nand NAND3_8695 ( P2_U4619 , P2_U8057 , P2_U8056 , P2_U3715 );
not NOT1_8696 ( P2_U4620 , P2_U3299 );
nand NAND2_8697 ( P2_U4621 , P2_U4474 , P2_U3265 );
nand NAND2_8698 ( P2_U4622 , P2_STATEBS16_REG , P2_U3284 );
nand NAND2_8699 ( P2_U4623 , P2_U4622 , P2_U4621 );
nand NAND2_8700 ( P2_U4624 , P2_STATE2_REG_1_ , P2_U4623 );
nand NAND2_8701 ( P2_U4625 , P2_STATE2_REG_2_ , P2_U3299 );
nand NAND2_8702 ( P2_U4626 , P2_U4619 , P2_U4465 );
nand NAND2_8703 ( P2_U4627 , P2_U3717 , P2_U4620 );
nand NAND2_8704 ( P2_U4628 , P2_STATE2_REG_1_ , P2_U4626 );
nand NAND2_8705 ( P2_U4629 , P2_U2374 , P2_U4619 );
nand NAND2_8706 ( P2_U4630 , P2_U3719 , P2_U4469 );
nand NAND2_8707 ( P2_U4631 , P2_U4619 , P2_U4464 );
nand NAND2_8708 ( P2_U4632 , P2_U2374 , P2_U3298 );
not NOT1_8709 ( P2_U4633 , P2_U3337 );
not NOT1_8710 ( P2_U4634 , P2_U3351 );
not NOT1_8711 ( P2_U4635 , P2_U3352 );
not NOT1_8712 ( P2_U4636 , P2_U3319 );
not NOT1_8713 ( P2_U4637 , P2_U3318 );
not NOT1_8714 ( P2_U4638 , P2_U3378 );
nand NAND2_8715 ( P2_U4639 , P2_R2182_U76 , P2_U3318 );
not NOT1_8716 ( P2_U4640 , P2_U3426 );
not NOT1_8717 ( P2_U4641 , P2_U3320 );
not NOT1_8718 ( P2_U4642 , P2_U3311 );
not NOT1_8719 ( P2_U4643 , P2_U3312 );
not NOT1_8720 ( P2_U4644 , P2_U3424 );
not NOT1_8721 ( P2_U4645 , P2_U3376 );
nand NAND2_8722 ( P2_U4646 , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_U3311 );
not NOT1_8723 ( P2_U4647 , P2_U3428 );
not NOT1_8724 ( P2_U4648 , P2_U3349 );
not NOT1_8725 ( P2_U4649 , P2_U3335 );
not NOT1_8726 ( P2_U4650 , P2_U3243 );
nand NAND2_8727 ( P2_U4651 , P2_U2440 , P2_U2444 );
not NOT1_8728 ( P2_U4652 , P2_U3325 );
not NOT1_8729 ( P2_U4653 , P2_U3570 );
not NOT1_8730 ( P2_U4654 , P2_U3326 );
nand NAND2_8731 ( P2_U4655 , P2_STATE2_REG_1_ , P2_U3270 );
nand NAND3_8732 ( P2_U4656 , P2_U4655 , P2_U3304 , P2_U3305 );
nand NAND2_8733 ( P2_U4657 , P2_U4637 , P2_U2462 );
nand NAND2_8734 ( P2_U4658 , P2_U2468 , P2_U2362 );
nand NAND2_8735 ( P2_U4659 , P2_U4445 , P2_U4658 );
nand NAND2_8736 ( P2_U4660 , P2_U4652 , P2_U4659 );
nand NAND2_8737 ( P2_U4661 , P2_U4654 , P2_STATE2_REG_2_ );
nand NAND2_8738 ( P2_U4662 , P2_STATE2_REG_3_ , P2_U3312 );
nand NAND2_8739 ( P2_U4663 , P2_U4660 , P2_U3722 );
nand NAND2_8740 ( P2_U4664 , P2_U2468 , P2_U2398 );
nand NAND2_8741 ( P2_U4665 , P2_U4445 , P2_U4664 );
nand NAND2_8742 ( P2_U4666 , P2_U4665 , P2_U3325 );
nand NAND2_8743 ( P2_U4667 , P2_STATE2_REG_2_ , P2_U3326 );
nand NAND2_8744 ( P2_U4668 , P2_U4667 , P2_U4666 );
nand NAND2_8745 ( P2_U4669 , P2_U2425 , P2_U4643 );
nand NAND2_8746 ( P2_U4670 , P2_U2422 , P2_U2463 );
nand NAND2_8747 ( P2_U4671 , P2_U2421 , P2_U4641 );
nand NAND2_8748 ( P2_U4672 , P2_U2406 , P2_U4668 );
nand NAND2_8749 ( P2_U4673 , P2_INSTQUEUE_REG_15__7_ , P2_U4663 );
nand NAND2_8750 ( P2_U4674 , P2_U2426 , P2_U4643 );
nand NAND2_8751 ( P2_U4675 , P2_U2420 , P2_U2463 );
nand NAND2_8752 ( P2_U4676 , P2_U2419 , P2_U4641 );
nand NAND2_8753 ( P2_U4677 , P2_U2405 , P2_U4668 );
nand NAND2_8754 ( P2_U4678 , P2_INSTQUEUE_REG_15__6_ , P2_U4663 );
nand NAND2_8755 ( P2_U4679 , P2_U2429 , P2_U4643 );
nand NAND2_8756 ( P2_U4680 , P2_U2418 , P2_U2463 );
nand NAND2_8757 ( P2_U4681 , P2_U2417 , P2_U4641 );
nand NAND2_8758 ( P2_U4682 , P2_U2404 , P2_U4668 );
nand NAND2_8759 ( P2_U4683 , P2_INSTQUEUE_REG_15__5_ , P2_U4663 );
nand NAND2_8760 ( P2_U4684 , P2_U2424 , P2_U4643 );
nand NAND2_8761 ( P2_U4685 , P2_U2416 , P2_U2463 );
nand NAND2_8762 ( P2_U4686 , P2_U2415 , P2_U4641 );
nand NAND2_8763 ( P2_U4687 , P2_U2403 , P2_U4668 );
nand NAND2_8764 ( P2_U4688 , P2_INSTQUEUE_REG_15__4_ , P2_U4663 );
nand NAND2_8765 ( P2_U4689 , P2_U2423 , P2_U4643 );
nand NAND2_8766 ( P2_U4690 , P2_U2414 , P2_U2463 );
nand NAND2_8767 ( P2_U4691 , P2_U2413 , P2_U4641 );
nand NAND2_8768 ( P2_U4692 , P2_U2402 , P2_U4668 );
nand NAND2_8769 ( P2_U4693 , P2_INSTQUEUE_REG_15__3_ , P2_U4663 );
nand NAND2_8770 ( P2_U4694 , P2_U2432 , P2_U4643 );
nand NAND2_8771 ( P2_U4695 , P2_U2412 , P2_U2463 );
nand NAND2_8772 ( P2_U4696 , P2_U2411 , P2_U4641 );
nand NAND2_8773 ( P2_U4697 , P2_U2401 , P2_U4668 );
nand NAND2_8774 ( P2_U4698 , P2_INSTQUEUE_REG_15__2_ , P2_U4663 );
nand NAND2_8775 ( P2_U4699 , P2_U2428 , P2_U4643 );
nand NAND2_8776 ( P2_U4700 , P2_U2410 , P2_U2463 );
nand NAND2_8777 ( P2_U4701 , P2_U2409 , P2_U4641 );
nand NAND2_8778 ( P2_U4702 , P2_U2400 , P2_U4668 );
nand NAND2_8779 ( P2_U4703 , P2_INSTQUEUE_REG_15__1_ , P2_U4663 );
nand NAND2_8780 ( P2_U4704 , P2_U2431 , P2_U4643 );
nand NAND2_8781 ( P2_U4705 , P2_U2408 , P2_U2463 );
nand NAND2_8782 ( P2_U4706 , P2_U2407 , P2_U4641 );
nand NAND2_8783 ( P2_U4707 , P2_U2399 , P2_U4668 );
nand NAND2_8784 ( P2_U4708 , P2_INSTQUEUE_REG_15__0_ , P2_U4663 );
not NOT1_8785 ( P2_U4709 , P2_U3338 );
not NOT1_8786 ( P2_U4710 , P2_U3339 );
not NOT1_8787 ( P2_U4711 , P2_U3336 );
not NOT1_8788 ( P2_U4712 , P2_U3245 );
not NOT1_8789 ( P2_U4713 , P2_U3569 );
not NOT1_8790 ( P2_U4714 , P2_U3340 );
nand NAND2_8791 ( P2_U4715 , P2_U4633 , P2_U2462 );
nand NAND2_8792 ( P2_U4716 , P2_U2471 , P2_U2362 );
nand NAND2_8793 ( P2_U4717 , P2_U4445 , P2_U4716 );
nand NAND2_8794 ( P2_U4718 , P2_U4717 , P2_U3245 );
nand NAND2_8795 ( P2_U4719 , P2_U4714 , P2_STATE2_REG_2_ );
nand NAND2_8796 ( P2_U4720 , P2_STATE2_REG_3_ , P2_U3336 );
nand NAND2_8797 ( P2_U4721 , P2_U4718 , P2_U3731 );
nand NAND2_8798 ( P2_U4722 , P2_U2471 , P2_U2398 );
nand NAND2_8799 ( P2_U4723 , P2_U4445 , P2_U4722 );
nand NAND2_8800 ( P2_U4724 , P2_U4723 , P2_U4712 );
nand NAND2_8801 ( P2_U4725 , P2_STATE2_REG_2_ , P2_U3340 );
nand NAND2_8802 ( P2_U4726 , P2_U4725 , P2_U4724 );
nand NAND2_8803 ( P2_U4727 , P2_U4711 , P2_U2425 );
nand NAND2_8804 ( P2_U4728 , P2_U2469 , P2_U2422 );
nand NAND2_8805 ( P2_U4729 , P2_U4710 , P2_U2421 );
nand NAND2_8806 ( P2_U4730 , P2_U2406 , P2_U4726 );
nand NAND2_8807 ( P2_U4731 , P2_INSTQUEUE_REG_14__7_ , P2_U4721 );
nand NAND2_8808 ( P2_U4732 , P2_U4711 , P2_U2426 );
nand NAND2_8809 ( P2_U4733 , P2_U2469 , P2_U2420 );
nand NAND2_8810 ( P2_U4734 , P2_U4710 , P2_U2419 );
nand NAND2_8811 ( P2_U4735 , P2_U2405 , P2_U4726 );
nand NAND2_8812 ( P2_U4736 , P2_INSTQUEUE_REG_14__6_ , P2_U4721 );
nand NAND2_8813 ( P2_U4737 , P2_U4711 , P2_U2429 );
nand NAND2_8814 ( P2_U4738 , P2_U2469 , P2_U2418 );
nand NAND2_8815 ( P2_U4739 , P2_U4710 , P2_U2417 );
nand NAND2_8816 ( P2_U4740 , P2_U2404 , P2_U4726 );
nand NAND2_8817 ( P2_U4741 , P2_INSTQUEUE_REG_14__5_ , P2_U4721 );
nand NAND2_8818 ( P2_U4742 , P2_U4711 , P2_U2424 );
nand NAND2_8819 ( P2_U4743 , P2_U2469 , P2_U2416 );
nand NAND2_8820 ( P2_U4744 , P2_U4710 , P2_U2415 );
nand NAND2_8821 ( P2_U4745 , P2_U2403 , P2_U4726 );
nand NAND2_8822 ( P2_U4746 , P2_INSTQUEUE_REG_14__4_ , P2_U4721 );
nand NAND2_8823 ( P2_U4747 , P2_U4711 , P2_U2423 );
nand NAND2_8824 ( P2_U4748 , P2_U2469 , P2_U2414 );
nand NAND2_8825 ( P2_U4749 , P2_U4710 , P2_U2413 );
nand NAND2_8826 ( P2_U4750 , P2_U2402 , P2_U4726 );
nand NAND2_8827 ( P2_U4751 , P2_INSTQUEUE_REG_14__3_ , P2_U4721 );
nand NAND2_8828 ( P2_U4752 , P2_U4711 , P2_U2432 );
nand NAND2_8829 ( P2_U4753 , P2_U2469 , P2_U2412 );
nand NAND2_8830 ( P2_U4754 , P2_U4710 , P2_U2411 );
nand NAND2_8831 ( P2_U4755 , P2_U2401 , P2_U4726 );
nand NAND2_8832 ( P2_U4756 , P2_INSTQUEUE_REG_14__2_ , P2_U4721 );
nand NAND2_8833 ( P2_U4757 , P2_U4711 , P2_U2428 );
nand NAND2_8834 ( P2_U4758 , P2_U2469 , P2_U2410 );
nand NAND2_8835 ( P2_U4759 , P2_U4710 , P2_U2409 );
nand NAND2_8836 ( P2_U4760 , P2_U2400 , P2_U4726 );
nand NAND2_8837 ( P2_U4761 , P2_INSTQUEUE_REG_14__1_ , P2_U4721 );
nand NAND2_8838 ( P2_U4762 , P2_U4711 , P2_U2431 );
nand NAND2_8839 ( P2_U4763 , P2_U2469 , P2_U2408 );
nand NAND2_8840 ( P2_U4764 , P2_U4710 , P2_U2407 );
nand NAND2_8841 ( P2_U4765 , P2_U2399 , P2_U4726 );
nand NAND2_8842 ( P2_U4766 , P2_INSTQUEUE_REG_14__0_ , P2_U4721 );
not NOT1_8843 ( P2_U4767 , P2_U3353 );
not NOT1_8844 ( P2_U4768 , P2_U3354 );
not NOT1_8845 ( P2_U4769 , P2_U3350 );
nand NAND2_8846 ( P2_U4770 , P2_U2445 , P2_U2440 );
not NOT1_8847 ( P2_U4771 , P2_U3355 );
not NOT1_8848 ( P2_U4772 , P2_U3568 );
not NOT1_8849 ( P2_U4773 , P2_U3356 );
nand NAND2_8850 ( P2_U4774 , P2_U4634 , P2_U2462 );
nand NAND2_8851 ( P2_U4775 , P2_U2474 , P2_U2362 );
nand NAND2_8852 ( P2_U4776 , P2_U4445 , P2_U4775 );
nand NAND2_8853 ( P2_U4777 , P2_U4771 , P2_U4776 );
nand NAND2_8854 ( P2_U4778 , P2_U4773 , P2_STATE2_REG_2_ );
nand NAND2_8855 ( P2_U4779 , P2_STATE2_REG_3_ , P2_U3350 );
nand NAND2_8856 ( P2_U4780 , P2_U4777 , P2_U3740 );
nand NAND2_8857 ( P2_U4781 , P2_U2474 , P2_U2398 );
nand NAND2_8858 ( P2_U4782 , P2_U4445 , P2_U4781 );
nand NAND2_8859 ( P2_U4783 , P2_U4782 , P2_U3355 );
nand NAND2_8860 ( P2_U4784 , P2_STATE2_REG_2_ , P2_U3356 );
nand NAND2_8861 ( P2_U4785 , P2_U4784 , P2_U4783 );
nand NAND2_8862 ( P2_U4786 , P2_U4769 , P2_U2425 );
nand NAND2_8863 ( P2_U4787 , P2_U2472 , P2_U2422 );
nand NAND2_8864 ( P2_U4788 , P2_U4768 , P2_U2421 );
nand NAND2_8865 ( P2_U4789 , P2_U2406 , P2_U4785 );
nand NAND2_8866 ( P2_U4790 , P2_INSTQUEUE_REG_13__7_ , P2_U4780 );
nand NAND2_8867 ( P2_U4791 , P2_U4769 , P2_U2426 );
nand NAND2_8868 ( P2_U4792 , P2_U2472 , P2_U2420 );
nand NAND2_8869 ( P2_U4793 , P2_U4768 , P2_U2419 );
nand NAND2_8870 ( P2_U4794 , P2_U2405 , P2_U4785 );
nand NAND2_8871 ( P2_U4795 , P2_INSTQUEUE_REG_13__6_ , P2_U4780 );
nand NAND2_8872 ( P2_U4796 , P2_U4769 , P2_U2429 );
nand NAND2_8873 ( P2_U4797 , P2_U2472 , P2_U2418 );
nand NAND2_8874 ( P2_U4798 , P2_U4768 , P2_U2417 );
nand NAND2_8875 ( P2_U4799 , P2_U2404 , P2_U4785 );
nand NAND2_8876 ( P2_U4800 , P2_INSTQUEUE_REG_13__5_ , P2_U4780 );
nand NAND2_8877 ( P2_U4801 , P2_U4769 , P2_U2424 );
nand NAND2_8878 ( P2_U4802 , P2_U2472 , P2_U2416 );
nand NAND2_8879 ( P2_U4803 , P2_U4768 , P2_U2415 );
nand NAND2_8880 ( P2_U4804 , P2_U2403 , P2_U4785 );
nand NAND2_8881 ( P2_U4805 , P2_INSTQUEUE_REG_13__4_ , P2_U4780 );
nand NAND2_8882 ( P2_U4806 , P2_U4769 , P2_U2423 );
nand NAND2_8883 ( P2_U4807 , P2_U2472 , P2_U2414 );
nand NAND2_8884 ( P2_U4808 , P2_U4768 , P2_U2413 );
nand NAND2_8885 ( P2_U4809 , P2_U2402 , P2_U4785 );
nand NAND2_8886 ( P2_U4810 , P2_INSTQUEUE_REG_13__3_ , P2_U4780 );
nand NAND2_8887 ( P2_U4811 , P2_U4769 , P2_U2432 );
nand NAND2_8888 ( P2_U4812 , P2_U2472 , P2_U2412 );
nand NAND2_8889 ( P2_U4813 , P2_U4768 , P2_U2411 );
nand NAND2_8890 ( P2_U4814 , P2_U2401 , P2_U4785 );
nand NAND2_8891 ( P2_U4815 , P2_INSTQUEUE_REG_13__2_ , P2_U4780 );
nand NAND2_8892 ( P2_U4816 , P2_U4769 , P2_U2428 );
nand NAND2_8893 ( P2_U4817 , P2_U2472 , P2_U2410 );
nand NAND2_8894 ( P2_U4818 , P2_U4768 , P2_U2409 );
nand NAND2_8895 ( P2_U4819 , P2_U2400 , P2_U4785 );
nand NAND2_8896 ( P2_U4820 , P2_INSTQUEUE_REG_13__1_ , P2_U4780 );
nand NAND2_8897 ( P2_U4821 , P2_U4769 , P2_U2431 );
nand NAND2_8898 ( P2_U4822 , P2_U2472 , P2_U2408 );
nand NAND2_8899 ( P2_U4823 , P2_U4768 , P2_U2407 );
nand NAND2_8900 ( P2_U4824 , P2_U2399 , P2_U4785 );
nand NAND2_8901 ( P2_U4825 , P2_INSTQUEUE_REG_13__0_ , P2_U4780 );
not NOT1_8902 ( P2_U4826 , P2_U3366 );
not NOT1_8903 ( P2_U4827 , P2_U3365 );
not NOT1_8904 ( P2_U4828 , P2_U3246 );
not NOT1_8905 ( P2_U4829 , P2_U3567 );
not NOT1_8906 ( P2_U4830 , P2_U3367 );
nand NAND2_8907 ( P2_U4831 , P2_U2476 , P2_U2462 );
nand NAND2_8908 ( P2_U4832 , P2_U2480 , P2_U2362 );
nand NAND2_8909 ( P2_U4833 , P2_U4445 , P2_U4832 );
nand NAND2_8910 ( P2_U4834 , P2_U4833 , P2_U3246 );
nand NAND2_8911 ( P2_U4835 , P2_U4830 , P2_STATE2_REG_2_ );
nand NAND2_8912 ( P2_U4836 , P2_STATE2_REG_3_ , P2_U3365 );
nand NAND2_8913 ( P2_U4837 , P2_U4834 , P2_U3749 );
nand NAND2_8914 ( P2_U4838 , P2_U2480 , P2_U2398 );
nand NAND2_8915 ( P2_U4839 , P2_U4445 , P2_U4838 );
nand NAND2_8916 ( P2_U4840 , P2_U4839 , P2_U4828 );
nand NAND2_8917 ( P2_U4841 , P2_STATE2_REG_2_ , P2_U3367 );
nand NAND2_8918 ( P2_U4842 , P2_U4841 , P2_U4840 );
nand NAND2_8919 ( P2_U4843 , P2_U4827 , P2_U2425 );
nand NAND2_8920 ( P2_U4844 , P2_U2477 , P2_U2422 );
nand NAND2_8921 ( P2_U4845 , P2_U4826 , P2_U2421 );
nand NAND2_8922 ( P2_U4846 , P2_U2406 , P2_U4842 );
nand NAND2_8923 ( P2_U4847 , P2_INSTQUEUE_REG_12__7_ , P2_U4837 );
nand NAND2_8924 ( P2_U4848 , P2_U4827 , P2_U2426 );
nand NAND2_8925 ( P2_U4849 , P2_U2477 , P2_U2420 );
nand NAND2_8926 ( P2_U4850 , P2_U4826 , P2_U2419 );
nand NAND2_8927 ( P2_U4851 , P2_U2405 , P2_U4842 );
nand NAND2_8928 ( P2_U4852 , P2_INSTQUEUE_REG_12__6_ , P2_U4837 );
nand NAND2_8929 ( P2_U4853 , P2_U4827 , P2_U2429 );
nand NAND2_8930 ( P2_U4854 , P2_U2477 , P2_U2418 );
nand NAND2_8931 ( P2_U4855 , P2_U4826 , P2_U2417 );
nand NAND2_8932 ( P2_U4856 , P2_U2404 , P2_U4842 );
nand NAND2_8933 ( P2_U4857 , P2_INSTQUEUE_REG_12__5_ , P2_U4837 );
nand NAND2_8934 ( P2_U4858 , P2_U4827 , P2_U2424 );
nand NAND2_8935 ( P2_U4859 , P2_U2477 , P2_U2416 );
nand NAND2_8936 ( P2_U4860 , P2_U4826 , P2_U2415 );
nand NAND2_8937 ( P2_U4861 , P2_U2403 , P2_U4842 );
nand NAND2_8938 ( P2_U4862 , P2_INSTQUEUE_REG_12__4_ , P2_U4837 );
nand NAND2_8939 ( P2_U4863 , P2_U4827 , P2_U2423 );
nand NAND2_8940 ( P2_U4864 , P2_U2477 , P2_U2414 );
nand NAND2_8941 ( P2_U4865 , P2_U4826 , P2_U2413 );
nand NAND2_8942 ( P2_U4866 , P2_U2402 , P2_U4842 );
nand NAND2_8943 ( P2_U4867 , P2_INSTQUEUE_REG_12__3_ , P2_U4837 );
nand NAND2_8944 ( P2_U4868 , P2_U4827 , P2_U2432 );
nand NAND2_8945 ( P2_U4869 , P2_U2477 , P2_U2412 );
nand NAND2_8946 ( P2_U4870 , P2_U4826 , P2_U2411 );
nand NAND2_8947 ( P2_U4871 , P2_U2401 , P2_U4842 );
nand NAND2_8948 ( P2_U4872 , P2_INSTQUEUE_REG_12__2_ , P2_U4837 );
nand NAND2_8949 ( P2_U4873 , P2_U4827 , P2_U2428 );
nand NAND2_8950 ( P2_U4874 , P2_U2477 , P2_U2410 );
nand NAND2_8951 ( P2_U4875 , P2_U4826 , P2_U2409 );
nand NAND2_8952 ( P2_U4876 , P2_U2400 , P2_U4842 );
nand NAND2_8953 ( P2_U4877 , P2_INSTQUEUE_REG_12__1_ , P2_U4837 );
nand NAND2_8954 ( P2_U4878 , P2_U4827 , P2_U2431 );
nand NAND2_8955 ( P2_U4879 , P2_U2477 , P2_U2408 );
nand NAND2_8956 ( P2_U4880 , P2_U4826 , P2_U2407 );
nand NAND2_8957 ( P2_U4881 , P2_U2399 , P2_U4842 );
nand NAND2_8958 ( P2_U4882 , P2_INSTQUEUE_REG_12__0_ , P2_U4837 );
not NOT1_8959 ( P2_U4883 , P2_U3379 );
not NOT1_8960 ( P2_U4884 , P2_U3377 );
nand NAND2_8961 ( P2_U4885 , P2_U2442 , P2_U2444 );
not NOT1_8962 ( P2_U4886 , P2_U3380 );
not NOT1_8963 ( P2_U4887 , P2_U3566 );
not NOT1_8964 ( P2_U4888 , P2_U3381 );
nand NAND2_8965 ( P2_U4889 , P2_U4638 , P2_U4637 );
nand NAND2_8966 ( P2_U4890 , P2_U2484 , P2_U2362 );
nand NAND2_8967 ( P2_U4891 , P2_U4445 , P2_U4890 );
nand NAND2_8968 ( P2_U4892 , P2_U4886 , P2_U4891 );
nand NAND2_8969 ( P2_U4893 , P2_U4888 , P2_STATE2_REG_2_ );
nand NAND2_8970 ( P2_U4894 , P2_STATE2_REG_3_ , P2_U3377 );
nand NAND2_8971 ( P2_U4895 , P2_U4892 , P2_U3758 );
nand NAND2_8972 ( P2_U4896 , P2_U2484 , P2_U2398 );
nand NAND2_8973 ( P2_U4897 , P2_U4445 , P2_U4896 );
nand NAND2_8974 ( P2_U4898 , P2_U4897 , P2_U3380 );
nand NAND2_8975 ( P2_U4899 , P2_STATE2_REG_2_ , P2_U3381 );
nand NAND2_8976 ( P2_U4900 , P2_U4899 , P2_U4898 );
nand NAND2_8977 ( P2_U4901 , P2_U4884 , P2_U2425 );
nand NAND2_8978 ( P2_U4902 , P2_U2482 , P2_U2422 );
nand NAND2_8979 ( P2_U4903 , P2_U4883 , P2_U2421 );
nand NAND2_8980 ( P2_U4904 , P2_U2406 , P2_U4900 );
nand NAND2_8981 ( P2_U4905 , P2_INSTQUEUE_REG_11__7_ , P2_U4895 );
nand NAND2_8982 ( P2_U4906 , P2_U4884 , P2_U2426 );
nand NAND2_8983 ( P2_U4907 , P2_U2482 , P2_U2420 );
nand NAND2_8984 ( P2_U4908 , P2_U4883 , P2_U2419 );
nand NAND2_8985 ( P2_U4909 , P2_U2405 , P2_U4900 );
nand NAND2_8986 ( P2_U4910 , P2_INSTQUEUE_REG_11__6_ , P2_U4895 );
nand NAND2_8987 ( P2_U4911 , P2_U4884 , P2_U2429 );
nand NAND2_8988 ( P2_U4912 , P2_U2482 , P2_U2418 );
nand NAND2_8989 ( P2_U4913 , P2_U4883 , P2_U2417 );
nand NAND2_8990 ( P2_U4914 , P2_U2404 , P2_U4900 );
nand NAND2_8991 ( P2_U4915 , P2_INSTQUEUE_REG_11__5_ , P2_U4895 );
nand NAND2_8992 ( P2_U4916 , P2_U4884 , P2_U2424 );
nand NAND2_8993 ( P2_U4917 , P2_U2482 , P2_U2416 );
nand NAND2_8994 ( P2_U4918 , P2_U4883 , P2_U2415 );
nand NAND2_8995 ( P2_U4919 , P2_U2403 , P2_U4900 );
nand NAND2_8996 ( P2_U4920 , P2_INSTQUEUE_REG_11__4_ , P2_U4895 );
nand NAND2_8997 ( P2_U4921 , P2_U4884 , P2_U2423 );
nand NAND2_8998 ( P2_U4922 , P2_U2482 , P2_U2414 );
nand NAND2_8999 ( P2_U4923 , P2_U4883 , P2_U2413 );
nand NAND2_9000 ( P2_U4924 , P2_U2402 , P2_U4900 );
nand NAND2_9001 ( P2_U4925 , P2_INSTQUEUE_REG_11__3_ , P2_U4895 );
nand NAND2_9002 ( P2_U4926 , P2_U4884 , P2_U2432 );
nand NAND2_9003 ( P2_U4927 , P2_U2482 , P2_U2412 );
nand NAND2_9004 ( P2_U4928 , P2_U4883 , P2_U2411 );
nand NAND2_9005 ( P2_U4929 , P2_U2401 , P2_U4900 );
nand NAND2_9006 ( P2_U4930 , P2_INSTQUEUE_REG_11__2_ , P2_U4895 );
nand NAND2_9007 ( P2_U4931 , P2_U4884 , P2_U2428 );
nand NAND2_9008 ( P2_U4932 , P2_U2482 , P2_U2410 );
nand NAND2_9009 ( P2_U4933 , P2_U4883 , P2_U2409 );
nand NAND2_9010 ( P2_U4934 , P2_U2400 , P2_U4900 );
nand NAND2_9011 ( P2_U4935 , P2_INSTQUEUE_REG_11__1_ , P2_U4895 );
nand NAND2_9012 ( P2_U4936 , P2_U4884 , P2_U2431 );
nand NAND2_9013 ( P2_U4937 , P2_U2482 , P2_U2408 );
nand NAND2_9014 ( P2_U4938 , P2_U4883 , P2_U2407 );
nand NAND2_9015 ( P2_U4939 , P2_U2399 , P2_U4900 );
nand NAND2_9016 ( P2_U4940 , P2_INSTQUEUE_REG_11__0_ , P2_U4895 );
not NOT1_9017 ( P2_U4941 , P2_U3391 );
not NOT1_9018 ( P2_U4942 , P2_U3390 );
not NOT1_9019 ( P2_U4943 , P2_U3247 );
not NOT1_9020 ( P2_U4944 , P2_U3565 );
not NOT1_9021 ( P2_U4945 , P2_U3392 );
nand NAND2_9022 ( P2_U4946 , P2_U4638 , P2_U4633 );
nand NAND2_9023 ( P2_U4947 , P2_U2486 , P2_U2362 );
nand NAND2_9024 ( P2_U4948 , P2_U4445 , P2_U4947 );
nand NAND2_9025 ( P2_U4949 , P2_U4948 , P2_U3247 );
nand NAND2_9026 ( P2_U4950 , P2_U4945 , P2_STATE2_REG_2_ );
nand NAND2_9027 ( P2_U4951 , P2_STATE2_REG_3_ , P2_U3390 );
nand NAND2_9028 ( P2_U4952 , P2_U4949 , P2_U3767 );
nand NAND2_9029 ( P2_U4953 , P2_U2486 , P2_U2398 );
nand NAND2_9030 ( P2_U4954 , P2_U4445 , P2_U4953 );
nand NAND2_9031 ( P2_U4955 , P2_U4954 , P2_U4943 );
nand NAND2_9032 ( P2_U4956 , P2_STATE2_REG_2_ , P2_U3392 );
nand NAND2_9033 ( P2_U4957 , P2_U4956 , P2_U4955 );
nand NAND2_9034 ( P2_U4958 , P2_U4942 , P2_U2425 );
nand NAND2_9035 ( P2_U4959 , P2_U2485 , P2_U2422 );
nand NAND2_9036 ( P2_U4960 , P2_U4941 , P2_U2421 );
nand NAND2_9037 ( P2_U4961 , P2_U2406 , P2_U4957 );
nand NAND2_9038 ( P2_U4962 , P2_INSTQUEUE_REG_10__7_ , P2_U4952 );
nand NAND2_9039 ( P2_U4963 , P2_U4942 , P2_U2426 );
nand NAND2_9040 ( P2_U4964 , P2_U2485 , P2_U2420 );
nand NAND2_9041 ( P2_U4965 , P2_U4941 , P2_U2419 );
nand NAND2_9042 ( P2_U4966 , P2_U2405 , P2_U4957 );
nand NAND2_9043 ( P2_U4967 , P2_INSTQUEUE_REG_10__6_ , P2_U4952 );
nand NAND2_9044 ( P2_U4968 , P2_U4942 , P2_U2429 );
nand NAND2_9045 ( P2_U4969 , P2_U2485 , P2_U2418 );
nand NAND2_9046 ( P2_U4970 , P2_U4941 , P2_U2417 );
nand NAND2_9047 ( P2_U4971 , P2_U2404 , P2_U4957 );
nand NAND2_9048 ( P2_U4972 , P2_INSTQUEUE_REG_10__5_ , P2_U4952 );
nand NAND2_9049 ( P2_U4973 , P2_U4942 , P2_U2424 );
nand NAND2_9050 ( P2_U4974 , P2_U2485 , P2_U2416 );
nand NAND2_9051 ( P2_U4975 , P2_U4941 , P2_U2415 );
nand NAND2_9052 ( P2_U4976 , P2_U2403 , P2_U4957 );
nand NAND2_9053 ( P2_U4977 , P2_INSTQUEUE_REG_10__4_ , P2_U4952 );
nand NAND2_9054 ( P2_U4978 , P2_U4942 , P2_U2423 );
nand NAND2_9055 ( P2_U4979 , P2_U2485 , P2_U2414 );
nand NAND2_9056 ( P2_U4980 , P2_U4941 , P2_U2413 );
nand NAND2_9057 ( P2_U4981 , P2_U2402 , P2_U4957 );
nand NAND2_9058 ( P2_U4982 , P2_INSTQUEUE_REG_10__3_ , P2_U4952 );
nand NAND2_9059 ( P2_U4983 , P2_U4942 , P2_U2432 );
nand NAND2_9060 ( P2_U4984 , P2_U2485 , P2_U2412 );
nand NAND2_9061 ( P2_U4985 , P2_U4941 , P2_U2411 );
nand NAND2_9062 ( P2_U4986 , P2_U2401 , P2_U4957 );
nand NAND2_9063 ( P2_U4987 , P2_INSTQUEUE_REG_10__2_ , P2_U4952 );
nand NAND2_9064 ( P2_U4988 , P2_U4942 , P2_U2428 );
nand NAND2_9065 ( P2_U4989 , P2_U2485 , P2_U2410 );
nand NAND2_9066 ( P2_U4990 , P2_U4941 , P2_U2409 );
nand NAND2_9067 ( P2_U4991 , P2_U2400 , P2_U4957 );
nand NAND2_9068 ( P2_U4992 , P2_INSTQUEUE_REG_10__1_ , P2_U4952 );
nand NAND2_9069 ( P2_U4993 , P2_U4942 , P2_U2431 );
nand NAND2_9070 ( P2_U4994 , P2_U2485 , P2_U2408 );
nand NAND2_9071 ( P2_U4995 , P2_U4941 , P2_U2407 );
nand NAND2_9072 ( P2_U4996 , P2_U2399 , P2_U4957 );
nand NAND2_9073 ( P2_U4997 , P2_INSTQUEUE_REG_10__0_ , P2_U4952 );
not NOT1_9074 ( P2_U4998 , P2_U3402 );
not NOT1_9075 ( P2_U4999 , P2_U3401 );
nand NAND2_9076 ( P2_U5000 , P2_U2442 , P2_U2445 );
not NOT1_9077 ( P2_U5001 , P2_U3403 );
not NOT1_9078 ( P2_U5002 , P2_U3564 );
not NOT1_9079 ( P2_U5003 , P2_U3404 );
nand NAND2_9080 ( P2_U5004 , P2_U4638 , P2_U4634 );
nand NAND2_9081 ( P2_U5005 , P2_U2488 , P2_U2362 );
nand NAND2_9082 ( P2_U5006 , P2_U4445 , P2_U5005 );
nand NAND2_9083 ( P2_U5007 , P2_U5001 , P2_U5006 );
nand NAND2_9084 ( P2_U5008 , P2_U5003 , P2_STATE2_REG_2_ );
nand NAND2_9085 ( P2_U5009 , P2_STATE2_REG_3_ , P2_U3401 );
nand NAND2_9086 ( P2_U5010 , P2_U5007 , P2_U3776 );
nand NAND2_9087 ( P2_U5011 , P2_U2488 , P2_U2398 );
nand NAND2_9088 ( P2_U5012 , P2_U4445 , P2_U5011 );
nand NAND2_9089 ( P2_U5013 , P2_U5012 , P2_U3403 );
nand NAND2_9090 ( P2_U5014 , P2_STATE2_REG_2_ , P2_U3404 );
nand NAND2_9091 ( P2_U5015 , P2_U5014 , P2_U5013 );
nand NAND2_9092 ( P2_U5016 , P2_U4999 , P2_U2425 );
nand NAND2_9093 ( P2_U5017 , P2_U2487 , P2_U2422 );
nand NAND2_9094 ( P2_U5018 , P2_U4998 , P2_U2421 );
nand NAND2_9095 ( P2_U5019 , P2_U2406 , P2_U5015 );
nand NAND2_9096 ( P2_U5020 , P2_INSTQUEUE_REG_9__7_ , P2_U5010 );
nand NAND2_9097 ( P2_U5021 , P2_U4999 , P2_U2426 );
nand NAND2_9098 ( P2_U5022 , P2_U2487 , P2_U2420 );
nand NAND2_9099 ( P2_U5023 , P2_U4998 , P2_U2419 );
nand NAND2_9100 ( P2_U5024 , P2_U2405 , P2_U5015 );
nand NAND2_9101 ( P2_U5025 , P2_INSTQUEUE_REG_9__6_ , P2_U5010 );
nand NAND2_9102 ( P2_U5026 , P2_U4999 , P2_U2429 );
nand NAND2_9103 ( P2_U5027 , P2_U2487 , P2_U2418 );
nand NAND2_9104 ( P2_U5028 , P2_U4998 , P2_U2417 );
nand NAND2_9105 ( P2_U5029 , P2_U2404 , P2_U5015 );
nand NAND2_9106 ( P2_U5030 , P2_INSTQUEUE_REG_9__5_ , P2_U5010 );
nand NAND2_9107 ( P2_U5031 , P2_U4999 , P2_U2424 );
nand NAND2_9108 ( P2_U5032 , P2_U2487 , P2_U2416 );
nand NAND2_9109 ( P2_U5033 , P2_U4998 , P2_U2415 );
nand NAND2_9110 ( P2_U5034 , P2_U2403 , P2_U5015 );
nand NAND2_9111 ( P2_U5035 , P2_INSTQUEUE_REG_9__4_ , P2_U5010 );
nand NAND2_9112 ( P2_U5036 , P2_U4999 , P2_U2423 );
nand NAND2_9113 ( P2_U5037 , P2_U2487 , P2_U2414 );
nand NAND2_9114 ( P2_U5038 , P2_U4998 , P2_U2413 );
nand NAND2_9115 ( P2_U5039 , P2_U2402 , P2_U5015 );
nand NAND2_9116 ( P2_U5040 , P2_INSTQUEUE_REG_9__3_ , P2_U5010 );
nand NAND2_9117 ( P2_U5041 , P2_U4999 , P2_U2432 );
nand NAND2_9118 ( P2_U5042 , P2_U2487 , P2_U2412 );
nand NAND2_9119 ( P2_U5043 , P2_U4998 , P2_U2411 );
nand NAND2_9120 ( P2_U5044 , P2_U2401 , P2_U5015 );
nand NAND2_9121 ( P2_U5045 , P2_INSTQUEUE_REG_9__2_ , P2_U5010 );
nand NAND2_9122 ( P2_U5046 , P2_U4999 , P2_U2428 );
nand NAND2_9123 ( P2_U5047 , P2_U2487 , P2_U2410 );
nand NAND2_9124 ( P2_U5048 , P2_U4998 , P2_U2409 );
nand NAND2_9125 ( P2_U5049 , P2_U2400 , P2_U5015 );
nand NAND2_9126 ( P2_U5050 , P2_INSTQUEUE_REG_9__1_ , P2_U5010 );
nand NAND2_9127 ( P2_U5051 , P2_U4999 , P2_U2431 );
nand NAND2_9128 ( P2_U5052 , P2_U2487 , P2_U2408 );
nand NAND2_9129 ( P2_U5053 , P2_U4998 , P2_U2407 );
nand NAND2_9130 ( P2_U5054 , P2_U2399 , P2_U5015 );
nand NAND2_9131 ( P2_U5055 , P2_INSTQUEUE_REG_9__0_ , P2_U5010 );
not NOT1_9132 ( P2_U5056 , P2_U3414 );
not NOT1_9133 ( P2_U5057 , P2_U3413 );
not NOT1_9134 ( P2_U5058 , P2_U3248 );
not NOT1_9135 ( P2_U5059 , P2_U3563 );
not NOT1_9136 ( P2_U5060 , P2_U3415 );
nand NAND2_9137 ( P2_U5061 , P2_U4638 , P2_U2476 );
nand NAND2_9138 ( P2_U5062 , P2_U2490 , P2_U2362 );
nand NAND2_9139 ( P2_U5063 , P2_U4445 , P2_U5062 );
nand NAND2_9140 ( P2_U5064 , P2_U5063 , P2_U3248 );
nand NAND2_9141 ( P2_U5065 , P2_U5060 , P2_STATE2_REG_2_ );
nand NAND2_9142 ( P2_U5066 , P2_STATE2_REG_3_ , P2_U3413 );
nand NAND2_9143 ( P2_U5067 , P2_U5064 , P2_U3785 );
nand NAND2_9144 ( P2_U5068 , P2_U2490 , P2_U2398 );
nand NAND2_9145 ( P2_U5069 , P2_U4445 , P2_U5068 );
nand NAND2_9146 ( P2_U5070 , P2_U5069 , P2_U5058 );
nand NAND2_9147 ( P2_U5071 , P2_STATE2_REG_2_ , P2_U3415 );
nand NAND2_9148 ( P2_U5072 , P2_U5071 , P2_U5070 );
nand NAND2_9149 ( P2_U5073 , P2_U5057 , P2_U2425 );
nand NAND2_9150 ( P2_U5074 , P2_U2489 , P2_U2422 );
nand NAND2_9151 ( P2_U5075 , P2_U5056 , P2_U2421 );
nand NAND2_9152 ( P2_U5076 , P2_U2406 , P2_U5072 );
nand NAND2_9153 ( P2_U5077 , P2_INSTQUEUE_REG_8__7_ , P2_U5067 );
nand NAND2_9154 ( P2_U5078 , P2_U5057 , P2_U2426 );
nand NAND2_9155 ( P2_U5079 , P2_U2489 , P2_U2420 );
nand NAND2_9156 ( P2_U5080 , P2_U5056 , P2_U2419 );
nand NAND2_9157 ( P2_U5081 , P2_U2405 , P2_U5072 );
nand NAND2_9158 ( P2_U5082 , P2_INSTQUEUE_REG_8__6_ , P2_U5067 );
nand NAND2_9159 ( P2_U5083 , P2_U5057 , P2_U2429 );
nand NAND2_9160 ( P2_U5084 , P2_U2489 , P2_U2418 );
nand NAND2_9161 ( P2_U5085 , P2_U5056 , P2_U2417 );
nand NAND2_9162 ( P2_U5086 , P2_U2404 , P2_U5072 );
nand NAND2_9163 ( P2_U5087 , P2_INSTQUEUE_REG_8__5_ , P2_U5067 );
nand NAND2_9164 ( P2_U5088 , P2_U5057 , P2_U2424 );
nand NAND2_9165 ( P2_U5089 , P2_U2489 , P2_U2416 );
nand NAND2_9166 ( P2_U5090 , P2_U5056 , P2_U2415 );
nand NAND2_9167 ( P2_U5091 , P2_U2403 , P2_U5072 );
nand NAND2_9168 ( P2_U5092 , P2_INSTQUEUE_REG_8__4_ , P2_U5067 );
nand NAND2_9169 ( P2_U5093 , P2_U5057 , P2_U2423 );
nand NAND2_9170 ( P2_U5094 , P2_U2489 , P2_U2414 );
nand NAND2_9171 ( P2_U5095 , P2_U5056 , P2_U2413 );
nand NAND2_9172 ( P2_U5096 , P2_U2402 , P2_U5072 );
nand NAND2_9173 ( P2_U5097 , P2_INSTQUEUE_REG_8__3_ , P2_U5067 );
nand NAND2_9174 ( P2_U5098 , P2_U5057 , P2_U2432 );
nand NAND2_9175 ( P2_U5099 , P2_U2489 , P2_U2412 );
nand NAND2_9176 ( P2_U5100 , P2_U5056 , P2_U2411 );
nand NAND2_9177 ( P2_U5101 , P2_U2401 , P2_U5072 );
nand NAND2_9178 ( P2_U5102 , P2_INSTQUEUE_REG_8__2_ , P2_U5067 );
nand NAND2_9179 ( P2_U5103 , P2_U5057 , P2_U2428 );
nand NAND2_9180 ( P2_U5104 , P2_U2489 , P2_U2410 );
nand NAND2_9181 ( P2_U5105 , P2_U5056 , P2_U2409 );
nand NAND2_9182 ( P2_U5106 , P2_U2400 , P2_U5072 );
nand NAND2_9183 ( P2_U5107 , P2_INSTQUEUE_REG_8__1_ , P2_U5067 );
nand NAND2_9184 ( P2_U5108 , P2_U5057 , P2_U2431 );
nand NAND2_9185 ( P2_U5109 , P2_U2489 , P2_U2408 );
nand NAND2_9186 ( P2_U5110 , P2_U5056 , P2_U2407 );
nand NAND2_9187 ( P2_U5111 , P2_U2399 , P2_U5072 );
nand NAND2_9188 ( P2_U5112 , P2_INSTQUEUE_REG_8__0_ , P2_U5067 );
not NOT1_9189 ( P2_U5113 , P2_U3427 );
nand NAND2_9190 ( P2_U5114 , P2_U2441 , P2_U2444 );
not NOT1_9191 ( P2_U5115 , P2_U3429 );
not NOT1_9192 ( P2_U5116 , P2_U3562 );
not NOT1_9193 ( P2_U5117 , P2_U3430 );
nand NAND2_9194 ( P2_U5118 , P2_U2493 , P2_U2362 );
nand NAND2_9195 ( P2_U5119 , P2_U4445 , P2_U5118 );
nand NAND2_9196 ( P2_U5120 , P2_U5115 , P2_U5119 );
nand NAND2_9197 ( P2_U5121 , P2_U5117 , P2_STATE2_REG_2_ );
nand NAND2_9198 ( P2_U5122 , P2_STATE2_REG_3_ , P2_U3424 );
nand NAND2_9199 ( P2_U5123 , P2_U5120 , P2_U3794 );
nand NAND2_9200 ( P2_U5124 , P2_U2493 , P2_U2398 );
nand NAND2_9201 ( P2_U5125 , P2_U4445 , P2_U5124 );
nand NAND2_9202 ( P2_U5126 , P2_U5125 , P2_U3429 );
nand NAND2_9203 ( P2_U5127 , P2_STATE2_REG_2_ , P2_U3430 );
nand NAND2_9204 ( P2_U5128 , P2_U5127 , P2_U5126 );
nand NAND2_9205 ( P2_U5129 , P2_U4644 , P2_U2425 );
nand NAND2_9206 ( P2_U5130 , P2_U4451 , P2_U2422 );
nand NAND2_9207 ( P2_U5131 , P2_U5113 , P2_U2421 );
nand NAND2_9208 ( P2_U5132 , P2_U2406 , P2_U5128 );
nand NAND2_9209 ( P2_U5133 , P2_INSTQUEUE_REG_7__7_ , P2_U5123 );
nand NAND2_9210 ( P2_U5134 , P2_U4644 , P2_U2426 );
nand NAND2_9211 ( P2_U5135 , P2_U4451 , P2_U2420 );
nand NAND2_9212 ( P2_U5136 , P2_U5113 , P2_U2419 );
nand NAND2_9213 ( P2_U5137 , P2_U2405 , P2_U5128 );
nand NAND2_9214 ( P2_U5138 , P2_INSTQUEUE_REG_7__6_ , P2_U5123 );
nand NAND2_9215 ( P2_U5139 , P2_U4644 , P2_U2429 );
nand NAND2_9216 ( P2_U5140 , P2_U4451 , P2_U2418 );
nand NAND2_9217 ( P2_U5141 , P2_U5113 , P2_U2417 );
nand NAND2_9218 ( P2_U5142 , P2_U2404 , P2_U5128 );
nand NAND2_9219 ( P2_U5143 , P2_INSTQUEUE_REG_7__5_ , P2_U5123 );
nand NAND2_9220 ( P2_U5144 , P2_U4644 , P2_U2424 );
nand NAND2_9221 ( P2_U5145 , P2_U4451 , P2_U2416 );
nand NAND2_9222 ( P2_U5146 , P2_U5113 , P2_U2415 );
nand NAND2_9223 ( P2_U5147 , P2_U2403 , P2_U5128 );
nand NAND2_9224 ( P2_U5148 , P2_INSTQUEUE_REG_7__4_ , P2_U5123 );
nand NAND2_9225 ( P2_U5149 , P2_U4644 , P2_U2423 );
nand NAND2_9226 ( P2_U5150 , P2_U4451 , P2_U2414 );
nand NAND2_9227 ( P2_U5151 , P2_U5113 , P2_U2413 );
nand NAND2_9228 ( P2_U5152 , P2_U2402 , P2_U5128 );
nand NAND2_9229 ( P2_U5153 , P2_INSTQUEUE_REG_7__3_ , P2_U5123 );
nand NAND2_9230 ( P2_U5154 , P2_U4644 , P2_U2432 );
nand NAND2_9231 ( P2_U5155 , P2_U4451 , P2_U2412 );
nand NAND2_9232 ( P2_U5156 , P2_U5113 , P2_U2411 );
nand NAND2_9233 ( P2_U5157 , P2_U2401 , P2_U5128 );
nand NAND2_9234 ( P2_U5158 , P2_INSTQUEUE_REG_7__2_ , P2_U5123 );
nand NAND2_9235 ( P2_U5159 , P2_U4644 , P2_U2428 );
nand NAND2_9236 ( P2_U5160 , P2_U4451 , P2_U2410 );
nand NAND2_9237 ( P2_U5161 , P2_U5113 , P2_U2409 );
nand NAND2_9238 ( P2_U5162 , P2_U2400 , P2_U5128 );
nand NAND2_9239 ( P2_U5163 , P2_INSTQUEUE_REG_7__1_ , P2_U5123 );
nand NAND2_9240 ( P2_U5164 , P2_U4644 , P2_U2431 );
nand NAND2_9241 ( P2_U5165 , P2_U4451 , P2_U2408 );
nand NAND2_9242 ( P2_U5166 , P2_U5113 , P2_U2407 );
nand NAND2_9243 ( P2_U5167 , P2_U2399 , P2_U5128 );
nand NAND2_9244 ( P2_U5168 , P2_INSTQUEUE_REG_7__0_ , P2_U5123 );
not NOT1_9245 ( P2_U5169 , P2_U3440 );
not NOT1_9246 ( P2_U5170 , P2_U3439 );
not NOT1_9247 ( P2_U5171 , P2_U3249 );
not NOT1_9248 ( P2_U5172 , P2_U3561 );
not NOT1_9249 ( P2_U5173 , P2_U3441 );
nand NAND2_9250 ( P2_U5174 , P2_U4633 , P2_U2460 );
nand NAND2_9251 ( P2_U5175 , P2_U2495 , P2_U2362 );
nand NAND2_9252 ( P2_U5176 , P2_U4445 , P2_U5175 );
nand NAND2_9253 ( P2_U5177 , P2_U5176 , P2_U3249 );
nand NAND2_9254 ( P2_U5178 , P2_U5173 , P2_STATE2_REG_2_ );
nand NAND2_9255 ( P2_U5179 , P2_STATE2_REG_3_ , P2_U3439 );
nand NAND2_9256 ( P2_U5180 , P2_U5177 , P2_U3803 );
nand NAND2_9257 ( P2_U5181 , P2_U2495 , P2_U2398 );
nand NAND2_9258 ( P2_U5182 , P2_U4445 , P2_U5181 );
nand NAND2_9259 ( P2_U5183 , P2_U5182 , P2_U5171 );
nand NAND2_9260 ( P2_U5184 , P2_STATE2_REG_2_ , P2_U3441 );
nand NAND2_9261 ( P2_U5185 , P2_U5184 , P2_U5183 );
nand NAND2_9262 ( P2_U5186 , P2_U5170 , P2_U2425 );
nand NAND2_9263 ( P2_U5187 , P2_U2494 , P2_U2422 );
nand NAND2_9264 ( P2_U5188 , P2_U5169 , P2_U2421 );
nand NAND2_9265 ( P2_U5189 , P2_U2406 , P2_U5185 );
nand NAND2_9266 ( P2_U5190 , P2_INSTQUEUE_REG_6__7_ , P2_U5180 );
nand NAND2_9267 ( P2_U5191 , P2_U5170 , P2_U2426 );
nand NAND2_9268 ( P2_U5192 , P2_U2494 , P2_U2420 );
nand NAND2_9269 ( P2_U5193 , P2_U5169 , P2_U2419 );
nand NAND2_9270 ( P2_U5194 , P2_U2405 , P2_U5185 );
nand NAND2_9271 ( P2_U5195 , P2_INSTQUEUE_REG_6__6_ , P2_U5180 );
nand NAND2_9272 ( P2_U5196 , P2_U5170 , P2_U2429 );
nand NAND2_9273 ( P2_U5197 , P2_U2494 , P2_U2418 );
nand NAND2_9274 ( P2_U5198 , P2_U5169 , P2_U2417 );
nand NAND2_9275 ( P2_U5199 , P2_U2404 , P2_U5185 );
nand NAND2_9276 ( P2_U5200 , P2_INSTQUEUE_REG_6__5_ , P2_U5180 );
nand NAND2_9277 ( P2_U5201 , P2_U5170 , P2_U2424 );
nand NAND2_9278 ( P2_U5202 , P2_U2494 , P2_U2416 );
nand NAND2_9279 ( P2_U5203 , P2_U5169 , P2_U2415 );
nand NAND2_9280 ( P2_U5204 , P2_U2403 , P2_U5185 );
nand NAND2_9281 ( P2_U5205 , P2_INSTQUEUE_REG_6__4_ , P2_U5180 );
nand NAND2_9282 ( P2_U5206 , P2_U5170 , P2_U2423 );
nand NAND2_9283 ( P2_U5207 , P2_U2494 , P2_U2414 );
nand NAND2_9284 ( P2_U5208 , P2_U5169 , P2_U2413 );
nand NAND2_9285 ( P2_U5209 , P2_U2402 , P2_U5185 );
nand NAND2_9286 ( P2_U5210 , P2_INSTQUEUE_REG_6__3_ , P2_U5180 );
nand NAND2_9287 ( P2_U5211 , P2_U5170 , P2_U2432 );
nand NAND2_9288 ( P2_U5212 , P2_U2494 , P2_U2412 );
nand NAND2_9289 ( P2_U5213 , P2_U5169 , P2_U2411 );
nand NAND2_9290 ( P2_U5214 , P2_U2401 , P2_U5185 );
nand NAND2_9291 ( P2_U5215 , P2_INSTQUEUE_REG_6__2_ , P2_U5180 );
nand NAND2_9292 ( P2_U5216 , P2_U5170 , P2_U2428 );
nand NAND2_9293 ( P2_U5217 , P2_U2494 , P2_U2410 );
nand NAND2_9294 ( P2_U5218 , P2_U5169 , P2_U2409 );
nand NAND2_9295 ( P2_U5219 , P2_U2400 , P2_U5185 );
nand NAND2_9296 ( P2_U5220 , P2_INSTQUEUE_REG_6__1_ , P2_U5180 );
nand NAND2_9297 ( P2_U5221 , P2_U5170 , P2_U2431 );
nand NAND2_9298 ( P2_U5222 , P2_U2494 , P2_U2408 );
nand NAND2_9299 ( P2_U5223 , P2_U5169 , P2_U2407 );
nand NAND2_9300 ( P2_U5224 , P2_U2399 , P2_U5185 );
nand NAND2_9301 ( P2_U5225 , P2_INSTQUEUE_REG_6__0_ , P2_U5180 );
not NOT1_9302 ( P2_U5226 , P2_U3451 );
not NOT1_9303 ( P2_U5227 , P2_U3450 );
nand NAND2_9304 ( P2_U5228 , P2_U2441 , P2_U2445 );
not NOT1_9305 ( P2_U5229 , P2_U3452 );
not NOT1_9306 ( P2_U5230 , P2_U3560 );
not NOT1_9307 ( P2_U5231 , P2_U3453 );
nand NAND2_9308 ( P2_U5232 , P2_U4634 , P2_U2460 );
nand NAND2_9309 ( P2_U5233 , P2_U2497 , P2_U2362 );
nand NAND2_9310 ( P2_U5234 , P2_U4445 , P2_U5233 );
nand NAND2_9311 ( P2_U5235 , P2_U5229 , P2_U5234 );
nand NAND2_9312 ( P2_U5236 , P2_U5231 , P2_STATE2_REG_2_ );
nand NAND2_9313 ( P2_U5237 , P2_STATE2_REG_3_ , P2_U3450 );
nand NAND2_9314 ( P2_U5238 , P2_U5235 , P2_U3812 );
nand NAND2_9315 ( P2_U5239 , P2_U2497 , P2_U2398 );
nand NAND2_9316 ( P2_U5240 , P2_U4445 , P2_U5239 );
nand NAND2_9317 ( P2_U5241 , P2_U5240 , P2_U3452 );
nand NAND2_9318 ( P2_U5242 , P2_STATE2_REG_2_ , P2_U3453 );
nand NAND2_9319 ( P2_U5243 , P2_U5242 , P2_U5241 );
nand NAND2_9320 ( P2_U5244 , P2_U5227 , P2_U2425 );
nand NAND2_9321 ( P2_U5245 , P2_U2496 , P2_U2422 );
nand NAND2_9322 ( P2_U5246 , P2_U5226 , P2_U2421 );
nand NAND2_9323 ( P2_U5247 , P2_U2406 , P2_U5243 );
nand NAND2_9324 ( P2_U5248 , P2_INSTQUEUE_REG_5__7_ , P2_U5238 );
nand NAND2_9325 ( P2_U5249 , P2_U5227 , P2_U2426 );
nand NAND2_9326 ( P2_U5250 , P2_U2496 , P2_U2420 );
nand NAND2_9327 ( P2_U5251 , P2_U5226 , P2_U2419 );
nand NAND2_9328 ( P2_U5252 , P2_U2405 , P2_U5243 );
nand NAND2_9329 ( P2_U5253 , P2_INSTQUEUE_REG_5__6_ , P2_U5238 );
nand NAND2_9330 ( P2_U5254 , P2_U5227 , P2_U2429 );
nand NAND2_9331 ( P2_U5255 , P2_U2496 , P2_U2418 );
nand NAND2_9332 ( P2_U5256 , P2_U5226 , P2_U2417 );
nand NAND2_9333 ( P2_U5257 , P2_U2404 , P2_U5243 );
nand NAND2_9334 ( P2_U5258 , P2_INSTQUEUE_REG_5__5_ , P2_U5238 );
nand NAND2_9335 ( P2_U5259 , P2_U5227 , P2_U2424 );
nand NAND2_9336 ( P2_U5260 , P2_U2496 , P2_U2416 );
nand NAND2_9337 ( P2_U5261 , P2_U5226 , P2_U2415 );
nand NAND2_9338 ( P2_U5262 , P2_U2403 , P2_U5243 );
nand NAND2_9339 ( P2_U5263 , P2_INSTQUEUE_REG_5__4_ , P2_U5238 );
nand NAND2_9340 ( P2_U5264 , P2_U5227 , P2_U2423 );
nand NAND2_9341 ( P2_U5265 , P2_U2496 , P2_U2414 );
nand NAND2_9342 ( P2_U5266 , P2_U5226 , P2_U2413 );
nand NAND2_9343 ( P2_U5267 , P2_U2402 , P2_U5243 );
nand NAND2_9344 ( P2_U5268 , P2_INSTQUEUE_REG_5__3_ , P2_U5238 );
nand NAND2_9345 ( P2_U5269 , P2_U5227 , P2_U2432 );
nand NAND2_9346 ( P2_U5270 , P2_U2496 , P2_U2412 );
nand NAND2_9347 ( P2_U5271 , P2_U5226 , P2_U2411 );
nand NAND2_9348 ( P2_U5272 , P2_U2401 , P2_U5243 );
nand NAND2_9349 ( P2_U5273 , P2_INSTQUEUE_REG_5__2_ , P2_U5238 );
nand NAND2_9350 ( P2_U5274 , P2_U5227 , P2_U2428 );
nand NAND2_9351 ( P2_U5275 , P2_U2496 , P2_U2410 );
nand NAND2_9352 ( P2_U5276 , P2_U5226 , P2_U2409 );
nand NAND2_9353 ( P2_U5277 , P2_U2400 , P2_U5243 );
nand NAND2_9354 ( P2_U5278 , P2_INSTQUEUE_REG_5__1_ , P2_U5238 );
nand NAND2_9355 ( P2_U5279 , P2_U5227 , P2_U2431 );
nand NAND2_9356 ( P2_U5280 , P2_U2496 , P2_U2408 );
nand NAND2_9357 ( P2_U5281 , P2_U5226 , P2_U2407 );
nand NAND2_9358 ( P2_U5282 , P2_U2399 , P2_U5243 );
nand NAND2_9359 ( P2_U5283 , P2_INSTQUEUE_REG_5__0_ , P2_U5238 );
not NOT1_9360 ( P2_U5284 , P2_U3463 );
not NOT1_9361 ( P2_U5285 , P2_U3462 );
not NOT1_9362 ( P2_U5286 , P2_U3250 );
not NOT1_9363 ( P2_U5287 , P2_U3559 );
not NOT1_9364 ( P2_U5288 , P2_U3464 );
nand NAND2_9365 ( P2_U5289 , P2_U2476 , P2_U2460 );
nand NAND2_9366 ( P2_U5290 , P2_U2499 , P2_U2362 );
nand NAND2_9367 ( P2_U5291 , P2_U4445 , P2_U5290 );
nand NAND2_9368 ( P2_U5292 , P2_U5291 , P2_U3250 );
nand NAND2_9369 ( P2_U5293 , P2_U5288 , P2_STATE2_REG_2_ );
nand NAND2_9370 ( P2_U5294 , P2_STATE2_REG_3_ , P2_U3462 );
nand NAND2_9371 ( P2_U5295 , P2_U5292 , P2_U3821 );
nand NAND2_9372 ( P2_U5296 , P2_U2499 , P2_U2398 );
nand NAND2_9373 ( P2_U5297 , P2_U4445 , P2_U5296 );
nand NAND2_9374 ( P2_U5298 , P2_U5297 , P2_U5286 );
nand NAND2_9375 ( P2_U5299 , P2_STATE2_REG_2_ , P2_U3464 );
nand NAND2_9376 ( P2_U5300 , P2_U5299 , P2_U5298 );
nand NAND2_9377 ( P2_U5301 , P2_U5285 , P2_U2425 );
nand NAND2_9378 ( P2_U5302 , P2_U2498 , P2_U2422 );
nand NAND2_9379 ( P2_U5303 , P2_U5284 , P2_U2421 );
nand NAND2_9380 ( P2_U5304 , P2_U2406 , P2_U5300 );
nand NAND2_9381 ( P2_U5305 , P2_INSTQUEUE_REG_4__7_ , P2_U5295 );
nand NAND2_9382 ( P2_U5306 , P2_U5285 , P2_U2426 );
nand NAND2_9383 ( P2_U5307 , P2_U2498 , P2_U2420 );
nand NAND2_9384 ( P2_U5308 , P2_U5284 , P2_U2419 );
nand NAND2_9385 ( P2_U5309 , P2_U2405 , P2_U5300 );
nand NAND2_9386 ( P2_U5310 , P2_INSTQUEUE_REG_4__6_ , P2_U5295 );
nand NAND2_9387 ( P2_U5311 , P2_U5285 , P2_U2429 );
nand NAND2_9388 ( P2_U5312 , P2_U2498 , P2_U2418 );
nand NAND2_9389 ( P2_U5313 , P2_U5284 , P2_U2417 );
nand NAND2_9390 ( P2_U5314 , P2_U2404 , P2_U5300 );
nand NAND2_9391 ( P2_U5315 , P2_INSTQUEUE_REG_4__5_ , P2_U5295 );
nand NAND2_9392 ( P2_U5316 , P2_U5285 , P2_U2424 );
nand NAND2_9393 ( P2_U5317 , P2_U2498 , P2_U2416 );
nand NAND2_9394 ( P2_U5318 , P2_U5284 , P2_U2415 );
nand NAND2_9395 ( P2_U5319 , P2_U2403 , P2_U5300 );
nand NAND2_9396 ( P2_U5320 , P2_INSTQUEUE_REG_4__4_ , P2_U5295 );
nand NAND2_9397 ( P2_U5321 , P2_U5285 , P2_U2423 );
nand NAND2_9398 ( P2_U5322 , P2_U2498 , P2_U2414 );
nand NAND2_9399 ( P2_U5323 , P2_U5284 , P2_U2413 );
nand NAND2_9400 ( P2_U5324 , P2_U2402 , P2_U5300 );
nand NAND2_9401 ( P2_U5325 , P2_INSTQUEUE_REG_4__3_ , P2_U5295 );
nand NAND2_9402 ( P2_U5326 , P2_U5285 , P2_U2432 );
nand NAND2_9403 ( P2_U5327 , P2_U2498 , P2_U2412 );
nand NAND2_9404 ( P2_U5328 , P2_U5284 , P2_U2411 );
nand NAND2_9405 ( P2_U5329 , P2_U2401 , P2_U5300 );
nand NAND2_9406 ( P2_U5330 , P2_INSTQUEUE_REG_4__2_ , P2_U5295 );
nand NAND2_9407 ( P2_U5331 , P2_U5285 , P2_U2428 );
nand NAND2_9408 ( P2_U5332 , P2_U2498 , P2_U2410 );
nand NAND2_9409 ( P2_U5333 , P2_U5284 , P2_U2409 );
nand NAND2_9410 ( P2_U5334 , P2_U2400 , P2_U5300 );
nand NAND2_9411 ( P2_U5335 , P2_INSTQUEUE_REG_4__1_ , P2_U5295 );
nand NAND2_9412 ( P2_U5336 , P2_U5285 , P2_U2431 );
nand NAND2_9413 ( P2_U5337 , P2_U2498 , P2_U2408 );
nand NAND2_9414 ( P2_U5338 , P2_U5284 , P2_U2407 );
nand NAND2_9415 ( P2_U5339 , P2_U2399 , P2_U5300 );
nand NAND2_9416 ( P2_U5340 , P2_INSTQUEUE_REG_4__0_ , P2_U5295 );
not NOT1_9417 ( P2_U5341 , P2_U3474 );
not NOT1_9418 ( P2_U5342 , P2_U3473 );
nand NAND2_9419 ( P2_U5343 , P2_U2443 , P2_U2444 );
not NOT1_9420 ( P2_U5344 , P2_U3475 );
not NOT1_9421 ( P2_U5345 , P2_U3558 );
not NOT1_9422 ( P2_U5346 , P2_U3476 );
nand NAND2_9423 ( P2_U5347 , P2_U2501 , P2_U4637 );
nand NAND2_9424 ( P2_U5348 , P2_U2505 , P2_U2362 );
nand NAND2_9425 ( P2_U5349 , P2_U4445 , P2_U5348 );
nand NAND2_9426 ( P2_U5350 , P2_U5344 , P2_U5349 );
nand NAND2_9427 ( P2_U5351 , P2_U5346 , P2_STATE2_REG_2_ );
nand NAND2_9428 ( P2_U5352 , P2_STATE2_REG_3_ , P2_U3473 );
nand NAND2_9429 ( P2_U5353 , P2_U5350 , P2_U3830 );
nand NAND2_9430 ( P2_U5354 , P2_U2505 , P2_U2398 );
nand NAND2_9431 ( P2_U5355 , P2_U4445 , P2_U5354 );
nand NAND2_9432 ( P2_U5356 , P2_U5355 , P2_U3475 );
nand NAND2_9433 ( P2_U5357 , P2_STATE2_REG_2_ , P2_U3476 );
nand NAND2_9434 ( P2_U5358 , P2_U5357 , P2_U5356 );
nand NAND2_9435 ( P2_U5359 , P2_U5342 , P2_U2425 );
nand NAND2_9436 ( P2_U5360 , P2_U2502 , P2_U2422 );
nand NAND2_9437 ( P2_U5361 , P2_U5341 , P2_U2421 );
nand NAND2_9438 ( P2_U5362 , P2_U2406 , P2_U5358 );
nand NAND2_9439 ( P2_U5363 , P2_INSTQUEUE_REG_3__7_ , P2_U5353 );
nand NAND2_9440 ( P2_U5364 , P2_U5342 , P2_U2426 );
nand NAND2_9441 ( P2_U5365 , P2_U2502 , P2_U2420 );
nand NAND2_9442 ( P2_U5366 , P2_U5341 , P2_U2419 );
nand NAND2_9443 ( P2_U5367 , P2_U2405 , P2_U5358 );
nand NAND2_9444 ( P2_U5368 , P2_INSTQUEUE_REG_3__6_ , P2_U5353 );
nand NAND2_9445 ( P2_U5369 , P2_U5342 , P2_U2429 );
nand NAND2_9446 ( P2_U5370 , P2_U2502 , P2_U2418 );
nand NAND2_9447 ( P2_U5371 , P2_U5341 , P2_U2417 );
nand NAND2_9448 ( P2_U5372 , P2_U2404 , P2_U5358 );
nand NAND2_9449 ( P2_U5373 , P2_INSTQUEUE_REG_3__5_ , P2_U5353 );
nand NAND2_9450 ( P2_U5374 , P2_U5342 , P2_U2424 );
nand NAND2_9451 ( P2_U5375 , P2_U2502 , P2_U2416 );
nand NAND2_9452 ( P2_U5376 , P2_U5341 , P2_U2415 );
nand NAND2_9453 ( P2_U5377 , P2_U2403 , P2_U5358 );
nand NAND2_9454 ( P2_U5378 , P2_INSTQUEUE_REG_3__4_ , P2_U5353 );
nand NAND2_9455 ( P2_U5379 , P2_U5342 , P2_U2423 );
nand NAND2_9456 ( P2_U5380 , P2_U2502 , P2_U2414 );
nand NAND2_9457 ( P2_U5381 , P2_U5341 , P2_U2413 );
nand NAND2_9458 ( P2_U5382 , P2_U2402 , P2_U5358 );
nand NAND2_9459 ( P2_U5383 , P2_INSTQUEUE_REG_3__3_ , P2_U5353 );
nand NAND2_9460 ( P2_U5384 , P2_U5342 , P2_U2432 );
nand NAND2_9461 ( P2_U5385 , P2_U2502 , P2_U2412 );
nand NAND2_9462 ( P2_U5386 , P2_U5341 , P2_U2411 );
nand NAND2_9463 ( P2_U5387 , P2_U2401 , P2_U5358 );
nand NAND2_9464 ( P2_U5388 , P2_INSTQUEUE_REG_3__2_ , P2_U5353 );
nand NAND2_9465 ( P2_U5389 , P2_U5342 , P2_U2428 );
nand NAND2_9466 ( P2_U5390 , P2_U2502 , P2_U2410 );
nand NAND2_9467 ( P2_U5391 , P2_U5341 , P2_U2409 );
nand NAND2_9468 ( P2_U5392 , P2_U2400 , P2_U5358 );
nand NAND2_9469 ( P2_U5393 , P2_INSTQUEUE_REG_3__1_ , P2_U5353 );
nand NAND2_9470 ( P2_U5394 , P2_U5342 , P2_U2431 );
nand NAND2_9471 ( P2_U5395 , P2_U2502 , P2_U2408 );
nand NAND2_9472 ( P2_U5396 , P2_U5341 , P2_U2407 );
nand NAND2_9473 ( P2_U5397 , P2_U2399 , P2_U5358 );
nand NAND2_9474 ( P2_U5398 , P2_INSTQUEUE_REG_3__0_ , P2_U5353 );
not NOT1_9475 ( P2_U5399 , P2_U3486 );
not NOT1_9476 ( P2_U5400 , P2_U3485 );
not NOT1_9477 ( P2_U5401 , P2_U3251 );
not NOT1_9478 ( P2_U5402 , P2_U3557 );
not NOT1_9479 ( P2_U5403 , P2_U3487 );
nand NAND2_9480 ( P2_U5404 , P2_U2501 , P2_U4633 );
nand NAND2_9481 ( P2_U5405 , P2_U2507 , P2_U2362 );
nand NAND2_9482 ( P2_U5406 , P2_U4445 , P2_U5405 );
nand NAND2_9483 ( P2_U5407 , P2_U5406 , P2_U3251 );
nand NAND2_9484 ( P2_U5408 , P2_U5403 , P2_STATE2_REG_2_ );
nand NAND2_9485 ( P2_U5409 , P2_STATE2_REG_3_ , P2_U3485 );
nand NAND2_9486 ( P2_U5410 , P2_U5407 , P2_U3839 );
nand NAND2_9487 ( P2_U5411 , P2_U2507 , P2_U2398 );
nand NAND2_9488 ( P2_U5412 , P2_U4445 , P2_U5411 );
nand NAND2_9489 ( P2_U5413 , P2_U5412 , P2_U5401 );
nand NAND2_9490 ( P2_U5414 , P2_STATE2_REG_2_ , P2_U3487 );
nand NAND2_9491 ( P2_U5415 , P2_U5414 , P2_U5413 );
nand NAND2_9492 ( P2_U5416 , P2_U5400 , P2_U2425 );
nand NAND2_9493 ( P2_U5417 , P2_U2506 , P2_U2422 );
nand NAND2_9494 ( P2_U5418 , P2_U5399 , P2_U2421 );
nand NAND2_9495 ( P2_U5419 , P2_U2406 , P2_U5415 );
nand NAND2_9496 ( P2_U5420 , P2_INSTQUEUE_REG_2__7_ , P2_U5410 );
nand NAND2_9497 ( P2_U5421 , P2_U5400 , P2_U2426 );
nand NAND2_9498 ( P2_U5422 , P2_U2506 , P2_U2420 );
nand NAND2_9499 ( P2_U5423 , P2_U5399 , P2_U2419 );
nand NAND2_9500 ( P2_U5424 , P2_U2405 , P2_U5415 );
nand NAND2_9501 ( P2_U5425 , P2_INSTQUEUE_REG_2__6_ , P2_U5410 );
nand NAND2_9502 ( P2_U5426 , P2_U5400 , P2_U2429 );
nand NAND2_9503 ( P2_U5427 , P2_U2506 , P2_U2418 );
nand NAND2_9504 ( P2_U5428 , P2_U5399 , P2_U2417 );
nand NAND2_9505 ( P2_U5429 , P2_U2404 , P2_U5415 );
nand NAND2_9506 ( P2_U5430 , P2_INSTQUEUE_REG_2__5_ , P2_U5410 );
nand NAND2_9507 ( P2_U5431 , P2_U5400 , P2_U2424 );
nand NAND2_9508 ( P2_U5432 , P2_U2506 , P2_U2416 );
nand NAND2_9509 ( P2_U5433 , P2_U5399 , P2_U2415 );
nand NAND2_9510 ( P2_U5434 , P2_U2403 , P2_U5415 );
nand NAND2_9511 ( P2_U5435 , P2_INSTQUEUE_REG_2__4_ , P2_U5410 );
nand NAND2_9512 ( P2_U5436 , P2_U5400 , P2_U2423 );
nand NAND2_9513 ( P2_U5437 , P2_U2506 , P2_U2414 );
nand NAND2_9514 ( P2_U5438 , P2_U5399 , P2_U2413 );
nand NAND2_9515 ( P2_U5439 , P2_U2402 , P2_U5415 );
nand NAND2_9516 ( P2_U5440 , P2_INSTQUEUE_REG_2__3_ , P2_U5410 );
nand NAND2_9517 ( P2_U5441 , P2_U5400 , P2_U2432 );
nand NAND2_9518 ( P2_U5442 , P2_U2506 , P2_U2412 );
nand NAND2_9519 ( P2_U5443 , P2_U5399 , P2_U2411 );
nand NAND2_9520 ( P2_U5444 , P2_U2401 , P2_U5415 );
nand NAND2_9521 ( P2_U5445 , P2_INSTQUEUE_REG_2__2_ , P2_U5410 );
nand NAND2_9522 ( P2_U5446 , P2_U5400 , P2_U2428 );
nand NAND2_9523 ( P2_U5447 , P2_U2506 , P2_U2410 );
nand NAND2_9524 ( P2_U5448 , P2_U5399 , P2_U2409 );
nand NAND2_9525 ( P2_U5449 , P2_U2400 , P2_U5415 );
nand NAND2_9526 ( P2_U5450 , P2_INSTQUEUE_REG_2__1_ , P2_U5410 );
nand NAND2_9527 ( P2_U5451 , P2_U5400 , P2_U2431 );
nand NAND2_9528 ( P2_U5452 , P2_U2506 , P2_U2408 );
nand NAND2_9529 ( P2_U5453 , P2_U5399 , P2_U2407 );
nand NAND2_9530 ( P2_U5454 , P2_U2399 , P2_U5415 );
nand NAND2_9531 ( P2_U5455 , P2_INSTQUEUE_REG_2__0_ , P2_U5410 );
not NOT1_9532 ( P2_U5456 , P2_U3497 );
not NOT1_9533 ( P2_U5457 , P2_U3496 );
nand NAND2_9534 ( P2_U5458 , P2_U2443 , P2_U2445 );
not NOT1_9535 ( P2_U5459 , P2_U3498 );
not NOT1_9536 ( P2_U5460 , P2_U3556 );
not NOT1_9537 ( P2_U5461 , P2_U3499 );
nand NAND2_9538 ( P2_U5462 , P2_U2501 , P2_U4634 );
nand NAND2_9539 ( P2_U5463 , P2_U2509 , P2_U2362 );
nand NAND2_9540 ( P2_U5464 , P2_U4445 , P2_U5463 );
nand NAND2_9541 ( P2_U5465 , P2_U5459 , P2_U5464 );
nand NAND2_9542 ( P2_U5466 , P2_U5461 , P2_STATE2_REG_2_ );
nand NAND2_9543 ( P2_U5467 , P2_STATE2_REG_3_ , P2_U3496 );
nand NAND2_9544 ( P2_U5468 , P2_U5465 , P2_U3848 );
nand NAND2_9545 ( P2_U5469 , P2_U2509 , P2_U2398 );
nand NAND2_9546 ( P2_U5470 , P2_U4445 , P2_U5469 );
nand NAND2_9547 ( P2_U5471 , P2_U5470 , P2_U3498 );
nand NAND2_9548 ( P2_U5472 , P2_STATE2_REG_2_ , P2_U3499 );
nand NAND2_9549 ( P2_U5473 , P2_U5472 , P2_U5471 );
nand NAND2_9550 ( P2_U5474 , P2_U5457 , P2_U2425 );
nand NAND2_9551 ( P2_U5475 , P2_U2508 , P2_U2422 );
nand NAND2_9552 ( P2_U5476 , P2_U5456 , P2_U2421 );
nand NAND2_9553 ( P2_U5477 , P2_U2406 , P2_U5473 );
nand NAND2_9554 ( P2_U5478 , P2_INSTQUEUE_REG_1__7_ , P2_U5468 );
nand NAND2_9555 ( P2_U5479 , P2_U5457 , P2_U2426 );
nand NAND2_9556 ( P2_U5480 , P2_U2508 , P2_U2420 );
nand NAND2_9557 ( P2_U5481 , P2_U5456 , P2_U2419 );
nand NAND2_9558 ( P2_U5482 , P2_U2405 , P2_U5473 );
nand NAND2_9559 ( P2_U5483 , P2_INSTQUEUE_REG_1__6_ , P2_U5468 );
nand NAND2_9560 ( P2_U5484 , P2_U5457 , P2_U2429 );
nand NAND2_9561 ( P2_U5485 , P2_U2508 , P2_U2418 );
nand NAND2_9562 ( P2_U5486 , P2_U5456 , P2_U2417 );
nand NAND2_9563 ( P2_U5487 , P2_U2404 , P2_U5473 );
nand NAND2_9564 ( P2_U5488 , P2_INSTQUEUE_REG_1__5_ , P2_U5468 );
nand NAND2_9565 ( P2_U5489 , P2_U5457 , P2_U2424 );
nand NAND2_9566 ( P2_U5490 , P2_U2508 , P2_U2416 );
nand NAND2_9567 ( P2_U5491 , P2_U5456 , P2_U2415 );
nand NAND2_9568 ( P2_U5492 , P2_U2403 , P2_U5473 );
nand NAND2_9569 ( P2_U5493 , P2_INSTQUEUE_REG_1__4_ , P2_U5468 );
nand NAND2_9570 ( P2_U5494 , P2_U5457 , P2_U2423 );
nand NAND2_9571 ( P2_U5495 , P2_U2508 , P2_U2414 );
nand NAND2_9572 ( P2_U5496 , P2_U5456 , P2_U2413 );
nand NAND2_9573 ( P2_U5497 , P2_U2402 , P2_U5473 );
nand NAND2_9574 ( P2_U5498 , P2_INSTQUEUE_REG_1__3_ , P2_U5468 );
nand NAND2_9575 ( P2_U5499 , P2_U5457 , P2_U2432 );
nand NAND2_9576 ( P2_U5500 , P2_U2508 , P2_U2412 );
nand NAND2_9577 ( P2_U5501 , P2_U5456 , P2_U2411 );
nand NAND2_9578 ( P2_U5502 , P2_U2401 , P2_U5473 );
nand NAND2_9579 ( P2_U5503 , P2_INSTQUEUE_REG_1__2_ , P2_U5468 );
nand NAND2_9580 ( P2_U5504 , P2_U5457 , P2_U2428 );
nand NAND2_9581 ( P2_U5505 , P2_U2508 , P2_U2410 );
nand NAND2_9582 ( P2_U5506 , P2_U5456 , P2_U2409 );
nand NAND2_9583 ( P2_U5507 , P2_U2400 , P2_U5473 );
nand NAND2_9584 ( P2_U5508 , P2_INSTQUEUE_REG_1__1_ , P2_U5468 );
nand NAND2_9585 ( P2_U5509 , P2_U5457 , P2_U2431 );
nand NAND2_9586 ( P2_U5510 , P2_U2508 , P2_U2408 );
nand NAND2_9587 ( P2_U5511 , P2_U5456 , P2_U2407 );
nand NAND2_9588 ( P2_U5512 , P2_U2399 , P2_U5473 );
nand NAND2_9589 ( P2_U5513 , P2_INSTQUEUE_REG_1__0_ , P2_U5468 );
not NOT1_9590 ( P2_U5514 , P2_U3509 );
not NOT1_9591 ( P2_U5515 , P2_U3508 );
not NOT1_9592 ( P2_U5516 , P2_U3252 );
not NOT1_9593 ( P2_U5517 , P2_U3555 );
not NOT1_9594 ( P2_U5518 , P2_U3510 );
nand NAND2_9595 ( P2_U5519 , P2_U2501 , P2_U2476 );
nand NAND2_9596 ( P2_U5520 , P2_U2511 , P2_U2362 );
nand NAND2_9597 ( P2_U5521 , P2_U4445 , P2_U5520 );
nand NAND2_9598 ( P2_U5522 , P2_U5521 , P2_U3252 );
nand NAND2_9599 ( P2_U5523 , P2_U5518 , P2_STATE2_REG_2_ );
nand NAND2_9600 ( P2_U5524 , P2_STATE2_REG_3_ , P2_U3508 );
nand NAND2_9601 ( P2_U5525 , P2_U5522 , P2_U3857 );
nand NAND2_9602 ( P2_U5526 , P2_U2511 , P2_U2398 );
nand NAND2_9603 ( P2_U5527 , P2_U4445 , P2_U5526 );
nand NAND2_9604 ( P2_U5528 , P2_U5527 , P2_U5516 );
nand NAND2_9605 ( P2_U5529 , P2_STATE2_REG_2_ , P2_U3510 );
nand NAND2_9606 ( P2_U5530 , P2_U5529 , P2_U5528 );
nand NAND2_9607 ( P2_U5531 , P2_U5515 , P2_U2425 );
nand NAND2_9608 ( P2_U5532 , P2_U2510 , P2_U2422 );
nand NAND2_9609 ( P2_U5533 , P2_U5514 , P2_U2421 );
nand NAND2_9610 ( P2_U5534 , P2_U2406 , P2_U5530 );
nand NAND2_9611 ( P2_U5535 , P2_INSTQUEUE_REG_0__7_ , P2_U5525 );
nand NAND2_9612 ( P2_U5536 , P2_U5515 , P2_U2426 );
nand NAND2_9613 ( P2_U5537 , P2_U2510 , P2_U2420 );
nand NAND2_9614 ( P2_U5538 , P2_U5514 , P2_U2419 );
nand NAND2_9615 ( P2_U5539 , P2_U2405 , P2_U5530 );
nand NAND2_9616 ( P2_U5540 , P2_INSTQUEUE_REG_0__6_ , P2_U5525 );
nand NAND2_9617 ( P2_U5541 , P2_U5515 , P2_U2429 );
nand NAND2_9618 ( P2_U5542 , P2_U2510 , P2_U2418 );
nand NAND2_9619 ( P2_U5543 , P2_U5514 , P2_U2417 );
nand NAND2_9620 ( P2_U5544 , P2_U2404 , P2_U5530 );
nand NAND2_9621 ( P2_U5545 , P2_INSTQUEUE_REG_0__5_ , P2_U5525 );
nand NAND2_9622 ( P2_U5546 , P2_U5515 , P2_U2424 );
nand NAND2_9623 ( P2_U5547 , P2_U2510 , P2_U2416 );
nand NAND2_9624 ( P2_U5548 , P2_U5514 , P2_U2415 );
nand NAND2_9625 ( P2_U5549 , P2_U2403 , P2_U5530 );
nand NAND2_9626 ( P2_U5550 , P2_INSTQUEUE_REG_0__4_ , P2_U5525 );
nand NAND2_9627 ( P2_U5551 , P2_U5515 , P2_U2423 );
nand NAND2_9628 ( P2_U5552 , P2_U2510 , P2_U2414 );
nand NAND2_9629 ( P2_U5553 , P2_U5514 , P2_U2413 );
nand NAND2_9630 ( P2_U5554 , P2_U2402 , P2_U5530 );
nand NAND2_9631 ( P2_U5555 , P2_INSTQUEUE_REG_0__3_ , P2_U5525 );
nand NAND2_9632 ( P2_U5556 , P2_U5515 , P2_U2432 );
nand NAND2_9633 ( P2_U5557 , P2_U2510 , P2_U2412 );
nand NAND2_9634 ( P2_U5558 , P2_U5514 , P2_U2411 );
nand NAND2_9635 ( P2_U5559 , P2_U2401 , P2_U5530 );
nand NAND2_9636 ( P2_U5560 , P2_INSTQUEUE_REG_0__2_ , P2_U5525 );
nand NAND2_9637 ( P2_U5561 , P2_U5515 , P2_U2428 );
nand NAND2_9638 ( P2_U5562 , P2_U2510 , P2_U2410 );
nand NAND2_9639 ( P2_U5563 , P2_U5514 , P2_U2409 );
nand NAND2_9640 ( P2_U5564 , P2_U2400 , P2_U5530 );
nand NAND2_9641 ( P2_U5565 , P2_INSTQUEUE_REG_0__1_ , P2_U5525 );
nand NAND2_9642 ( P2_U5566 , P2_U5515 , P2_U2431 );
nand NAND2_9643 ( P2_U5567 , P2_U2510 , P2_U2408 );
nand NAND2_9644 ( P2_U5568 , P2_U5514 , P2_U2407 );
nand NAND2_9645 ( P2_U5569 , P2_U2399 , P2_U5530 );
nand NAND2_9646 ( P2_U5570 , P2_INSTQUEUE_REG_0__0_ , P2_U5525 );
nand NAND2_9647 ( P2_U5571 , P2_U3279 , P2_U7869 );
not NOT1_9648 ( P2_U5572 , P2_U3574 );
nand NAND3_9649 ( P2_U5573 , P2_U7863 , P2_U2617 , P2_U7861 );
nand NAND4_9650 ( P2_U5574 , P2_U7895 , P2_U3521 , P2_U3255 , P2_U3289 );
nand NAND2_9651 ( P2_U5575 , P2_U2357 , P2_U7871 );
nand NAND2_9652 ( P2_U5576 , P2_U4417 , P2_U3574 );
nand NAND2_9653 ( P2_U5577 , P2_U4428 , P2_U4424 );
nand NAND2_9654 ( P2_U5578 , P2_U3524 , P2_U5577 );
nand NAND3_9655 ( P2_U5579 , P2_U5578 , P2_U3265 , P2_R2088_U6 );
nand NAND2_9656 ( P2_U5580 , P2_U4436 , P2_R2167_U6 );
not NOT1_9657 ( P2_U5581 , P2_U4406 );
nand NAND2_9658 ( P2_U5582 , P2_U2374 , P2_U4406 );
nand NAND2_9659 ( P2_U5583 , P2_STATE2_REG_3_ , P2_U3284 );
not NOT1_9660 ( P2_U5584 , P2_U4394 );
nand NAND2_9661 ( P2_U5585 , P2_U4591 , P2_U3276 );
nand NAND3_9662 ( P2_U5586 , P2_U2617 , P2_U3295 , P2_U3878 );
nand NAND2_9663 ( P2_U5587 , P2_U3295 , P2_U3255 );
nand NAND2_9664 ( P2_U5588 , P2_U7865 , P2_U3278 );
nand NAND3_9665 ( P2_U5589 , P2_U8075 , P2_U8074 , P2_U3879 );
not NOT1_9666 ( P2_U5590 , P2_U3525 );
nand NAND2_9667 ( P2_U5591 , P2_U7738 , P2_U3278 );
nand NAND4_9668 ( P2_U5592 , P2_U3521 , P2_U5591 , P2_U5573 , P2_U5571 );
nand NAND2_9669 ( P2_U5593 , P2_U4417 , P2_U3574 );
nand NAND2_9670 ( P2_U5594 , P2_U5592 , P2_U2616 );
nand NAND2_9671 ( P2_U5595 , P2_U3877 , P2_U5594 );
nand NAND2_9672 ( P2_U5596 , P2_U3295 , P2_U7873 );
nand NAND2_9673 ( P2_U5597 , P2_U3279 , P2_U7871 );
nand NAND2_9674 ( P2_U5598 , P2_U2617 , P2_U3521 );
nand NAND2_9675 ( P2_U5599 , P2_U4427 , P2_U5598 );
nand NAND2_9676 ( P2_U5600 , P2_U5597 , P2_U3280 );
nand NAND2_9677 ( P2_U5601 , P2_U2436 , P2_U7884 );
nand NAND2_9678 ( P2_U5602 , P2_U3527 , P2_U3278 );
nand NAND2_9679 ( P2_U5603 , P2_U2514 , P2_U3288 );
nand NAND3_9680 ( P2_U5604 , P2_U8077 , P2_U8076 , P2_U4470 );
nand NAND2_9681 ( P2_U5605 , P2_U3296 , P2_U3522 );
nand NAND2_9682 ( P2_U5606 , P2_U3578 , P2_U4437 );
nand NAND2_9683 ( P2_U5607 , P2_U4395 , P2_U5605 );
nand NAND2_9684 ( P2_U5608 , P2_U3581 , P2_U5606 );
nand NAND2_9685 ( P2_U5609 , P2_R2147_U8 , P2_U5604 );
nand NAND2_9686 ( P2_U5610 , P2_R2099_U95 , P2_U5603 );
nand NAND2_9687 ( P2_U5611 , P2_U3884 , P2_U5610 );
nand NAND2_9688 ( P2_U5612 , P2_R2182_U76 , P2_U4469 );
nand NAND2_9689 ( P2_U5613 , P2_U4466 , P2_U5611 );
nand NAND2_9690 ( P2_U5614 , P2_U5613 , P2_U5612 );
nand NAND2_9691 ( P2_U5615 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_U4591 );
not NOT1_9692 ( P2_U5616 , P2_U3530 );
nand NAND2_9693 ( P2_U5617 , P2_R2147_U9 , P2_U5604 );
nand NAND2_9694 ( P2_U5618 , P2_R2099_U96 , P2_U5603 );
nand NAND2_9695 ( P2_U5619 , P2_U3885 , P2_U5618 );
nand NAND3_9696 ( P2_U5620 , P2_U3598 , P2_U3597 , P2_STATE2_REG_1_ );
nand NAND2_9697 ( P2_U5621 , P2_R2182_U40 , P2_U4469 );
nand NAND2_9698 ( P2_U5622 , P2_U4466 , P2_U5619 );
nand NAND3_9699 ( P2_U5623 , P2_U5621 , P2_U5622 , P2_U5620 );
nand NAND3_9700 ( P2_U5624 , P2_U2449 , P2_U7861 , P2_U4429 );
nand NAND2_9701 ( P2_U5625 , P2_U7882 , P2_U5624 );
nand NAND2_9702 ( P2_U5626 , P2_U3887 , P2_U8097 );
nand NAND2_9703 ( P2_U5627 , P2_R2147_U4 , P2_U5604 );
nand NAND2_9704 ( P2_U5628 , P2_R2099_U5 , P2_U5603 );
nand NAND2_9705 ( P2_U5629 , P2_U3888 , P2_U5628 );
nand NAND3_9706 ( P2_U5630 , P2_STATE2_REG_1_ , P2_U8090 , P2_U3597 );
nand NAND2_9707 ( P2_U5631 , P2_R2182_U68 , P2_U4469 );
nand NAND2_9708 ( P2_U5632 , P2_U4466 , P2_U5629 );
nand NAND3_9709 ( P2_U5633 , P2_U5631 , P2_U5632 , P2_U5630 );
nand NAND2_9710 ( P2_U5634 , P2_U3889 , P2_U8097 );
nand NAND2_9711 ( P2_U5635 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_U5604 );
nand NAND2_9712 ( P2_U5636 , P2_R2099_U94 , P2_U5603 );
nand NAND2_9713 ( P2_U5637 , P2_U3890 , P2_U5636 );
nand NAND2_9714 ( P2_U5638 , P2_R2182_U69 , P2_U4469 );
nand NAND2_9715 ( P2_U5639 , P2_U4466 , P2_U5637 );
nand NAND2_9716 ( P2_U5640 , P2_U8087 , P2_STATE2_REG_1_ );
nand NAND3_9717 ( P2_U5641 , P2_U5639 , P2_U5638 , P2_U5640 );
nand NAND3_9718 ( P2_U5642 , P2_U2448 , P2_STATE2_REG_0_ , P2_R2243_U8 );
not NOT1_9719 ( P2_U5643 , P2_U3533 );
nand NAND2_9720 ( P2_U5644 , P2_U4445 , P2_U3303 );
nand NAND2_9721 ( P2_U5645 , P2_U4636 , P2_U3579 );
nand NAND2_9722 ( P2_U5646 , P2_U3426 , P2_U5645 );
nand NAND2_9723 ( P2_U5647 , P2_U3427 , P2_U5646 );
nand NAND2_9724 ( P2_U5648 , P2_U2398 , P2_U5647 );
nand NAND2_9725 ( P2_U5649 , P2_R2182_U76 , P2_U5644 );
nand NAND2_9726 ( P2_U5650 , P2_R2096_U75 , P2_STATE2_REG_3_ );
nand NAND2_9727 ( P2_U5651 , P2_U3891 , P2_U5648 );
nand NAND2_9728 ( P2_U5652 , P2_U2398 , P2_U8109 );
nand NAND2_9729 ( P2_U5653 , P2_R2182_U40 , P2_U5644 );
nand NAND2_9730 ( P2_U5654 , P2_R2096_U77 , P2_STATE2_REG_3_ );
nand NAND2_9731 ( P2_U5655 , P2_U3892 , P2_U5652 );
nand NAND2_9732 ( P2_U5656 , P2_U3338 , P2_U3353 );
nand NAND2_9733 ( P2_U5657 , P2_U2398 , P2_U5656 );
nand NAND2_9734 ( P2_U5658 , P2_R2182_U68 , P2_U5644 );
nand NAND2_9735 ( P2_U5659 , P2_R2096_U51 , P2_STATE2_REG_3_ );
nand NAND2_9736 ( P2_U5660 , P2_U3893 , P2_U5657 );
nand NAND2_9737 ( P2_U5661 , P2_U3313 , P2_U3303 );
nand NAND2_9738 ( P2_U5662 , P2_R2182_U69 , P2_U5661 );
nand NAND2_9739 ( P2_U5663 , P2_R2096_U68 , P2_STATE2_REG_3_ );
nand NAND3_9740 ( P2_U5664 , P2_U5662 , P2_U5663 , P2_U4464 );
nand NAND2_9741 ( P2_U5665 , P2_U2616 , P2_U3292 );
nand NAND2_9742 ( P2_U5666 , P2_GTE_370_U6 , P2_U4417 );
nand NAND2_9743 ( P2_U5667 , P2_U5666 , P2_U5665 );
nand NAND4_9744 ( P2_U5668 , P2_U8122 , P2_U8121 , P2_U3265 , P2_R2088_U6 );
nand NAND2_9745 ( P2_U5669 , P2_U4420 , P2_U5667 );
nand NAND4_9746 ( P2_U5670 , P2_U2512 , P2_U3894 , P2_U4397 , P2_U5669 );
nand NAND2_9747 ( P2_U5671 , P2_U2374 , P2_U5670 );
nand NAND2_9748 ( P2_U5672 , P2_U4461 , P2_U3284 );
not NOT1_9749 ( P2_U5673 , P2_U3535 );
nand NAND2_9750 ( P2_U5674 , P2_U4427 , P2_U4420 );
nand NAND2_9751 ( P2_U5675 , P2_U3895 , P2_U2514 );
nand NAND2_9752 ( P2_U5676 , P2_U4417 , P2_U4424 );
nand NAND4_9753 ( P2_U5677 , P2_U5676 , P2_U4470 , P2_U4437 , P2_U3524 );
nand NAND2_9754 ( P2_U5678 , P2_U4428 , P2_U4424 );
nand NAND3_9755 ( P2_U5679 , P2_U3296 , P2_U5678 , P2_U3523 );
nand NAND2_9756 ( P2_U5680 , P2_U2390 , P2_R2096_U68 );
nand NAND2_9757 ( P2_U5681 , P2_U2389 , P2_R2099_U94 );
nand NAND2_9758 ( P2_U5682 , P2_R2027_U5 , P2_U2388 );
nand NAND2_9759 ( P2_U5683 , P2_ADD_394_U4 , P2_U2386 );
nand NAND2_9760 ( P2_U5684 , P2_R2278_U83 , P2_U2385 );
nand NAND2_9761 ( P2_U5685 , P2_ADD_371_1212_U68 , P2_U2384 );
nand NAND2_9762 ( P2_U5686 , P2_REIP_REG_0_ , P2_U2381 );
nand NAND2_9763 ( P2_U5687 , P2_U5673 , P2_INSTADDRPOINTER_REG_0_ );
nand NAND2_9764 ( P2_U5688 , P2_U2390 , P2_R2096_U51 );
nand NAND2_9765 ( P2_U5689 , P2_U2389 , P2_R2099_U5 );
nand NAND2_9766 ( P2_U5690 , P2_R2027_U85 , P2_U2388 );
nand NAND2_9767 ( P2_U5691 , P2_ADD_394_U85 , P2_U2386 );
nand NAND2_9768 ( P2_U5692 , P2_R2278_U6 , P2_U2385 );
nand NAND2_9769 ( P2_U5693 , P2_ADD_371_1212_U25 , P2_U2384 );
nand NAND2_9770 ( P2_U5694 , P2_U2381 , P2_REIP_REG_1_ );
nand NAND2_9771 ( P2_U5695 , P2_U5673 , P2_INSTADDRPOINTER_REG_1_ );
nand NAND2_9772 ( P2_U5696 , P2_U2390 , P2_R2096_U77 );
nand NAND2_9773 ( P2_U5697 , P2_U2389 , P2_R2099_U96 );
nand NAND2_9774 ( P2_U5698 , P2_R2027_U74 , P2_U2388 );
nand NAND2_9775 ( P2_U5699 , P2_ADD_394_U5 , P2_U2386 );
nand NAND2_9776 ( P2_U5700 , P2_R2278_U92 , P2_U2385 );
nand NAND2_9777 ( P2_U5701 , P2_ADD_371_1212_U79 , P2_U2384 );
nand NAND2_9778 ( P2_U5702 , P2_U2381 , P2_REIP_REG_2_ );
nand NAND2_9779 ( P2_U5703 , P2_INSTADDRPOINTER_REG_2_ , P2_U5673 );
nand NAND2_9780 ( P2_U5704 , P2_U2390 , P2_R2096_U75 );
nand NAND2_9781 ( P2_U5705 , P2_U2389 , P2_R2099_U95 );
nand NAND2_9782 ( P2_U5706 , P2_R2027_U71 , P2_U2388 );
nand NAND2_9783 ( P2_U5707 , P2_ADD_394_U95 , P2_U2386 );
nand NAND2_9784 ( P2_U5708 , P2_R2278_U90 , P2_U2385 );
nand NAND2_9785 ( P2_U5709 , P2_ADD_371_1212_U84 , P2_U2384 );
nand NAND2_9786 ( P2_U5710 , P2_U2381 , P2_REIP_REG_3_ );
nand NAND2_9787 ( P2_U5711 , P2_INSTADDRPOINTER_REG_3_ , P2_U5673 );
nand NAND2_9788 ( P2_U5712 , P2_R2096_U74 , P2_U2390 );
nand NAND2_9789 ( P2_U5713 , P2_R2099_U98 , P2_U2389 );
nand NAND2_9790 ( P2_U5714 , P2_R2027_U70 , P2_U2388 );
nand NAND2_9791 ( P2_U5715 , P2_ADD_394_U76 , P2_U2386 );
nand NAND2_9792 ( P2_U5716 , P2_R2278_U89 , P2_U2385 );
nand NAND2_9793 ( P2_U5717 , P2_ADD_371_1212_U80 , P2_U2384 );
nand NAND2_9794 ( P2_U5718 , P2_U2381 , P2_REIP_REG_4_ );
nand NAND2_9795 ( P2_U5719 , P2_INSTADDRPOINTER_REG_4_ , P2_U5673 );
nand NAND2_9796 ( P2_U5720 , P2_R2096_U73 , P2_U2390 );
nand NAND2_9797 ( P2_U5721 , P2_R2099_U71 , P2_U2389 );
nand NAND2_9798 ( P2_U5722 , P2_R2027_U69 , P2_U2388 );
nand NAND2_9799 ( P2_U5723 , P2_ADD_394_U79 , P2_U2386 );
nand NAND2_9800 ( P2_U5724 , P2_R2278_U88 , P2_U2385 );
nand NAND2_9801 ( P2_U5725 , P2_ADD_371_1212_U81 , P2_U2384 );
nand NAND2_9802 ( P2_U5726 , P2_U2381 , P2_REIP_REG_5_ );
nand NAND2_9803 ( P2_U5727 , P2_INSTADDRPOINTER_REG_5_ , P2_U5673 );
nand NAND2_9804 ( P2_U5728 , P2_R2096_U72 , P2_U2390 );
nand NAND2_9805 ( P2_U5729 , P2_R2099_U70 , P2_U2389 );
nand NAND2_9806 ( P2_U5730 , P2_R2027_U68 , P2_U2388 );
nand NAND2_9807 ( P2_U5731 , P2_ADD_394_U63 , P2_U2386 );
nand NAND2_9808 ( P2_U5732 , P2_R2278_U87 , P2_U2385 );
nand NAND2_9809 ( P2_U5733 , P2_ADD_371_1212_U78 , P2_U2384 );
nand NAND2_9810 ( P2_U5734 , P2_U2381 , P2_REIP_REG_6_ );
nand NAND2_9811 ( P2_U5735 , P2_INSTADDRPOINTER_REG_6_ , P2_U5673 );
nand NAND2_9812 ( P2_U5736 , P2_R2096_U71 , P2_U2390 );
nand NAND2_9813 ( P2_U5737 , P2_R2099_U69 , P2_U2389 );
nand NAND2_9814 ( P2_U5738 , P2_R2027_U67 , P2_U2388 );
nand NAND2_9815 ( P2_U5739 , P2_ADD_394_U89 , P2_U2386 );
nand NAND2_9816 ( P2_U5740 , P2_R2278_U86 , P2_U2385 );
nand NAND2_9817 ( P2_U5741 , P2_ADD_371_1212_U85 , P2_U2384 );
nand NAND2_9818 ( P2_U5742 , P2_U2381 , P2_REIP_REG_7_ );
nand NAND2_9819 ( P2_U5743 , P2_INSTADDRPOINTER_REG_7_ , P2_U5673 );
nand NAND2_9820 ( P2_U5744 , P2_R2096_U70 , P2_U2390 );
nand NAND2_9821 ( P2_U5745 , P2_R2099_U68 , P2_U2389 );
nand NAND2_9822 ( P2_U5746 , P2_R2027_U66 , P2_U2388 );
nand NAND2_9823 ( P2_U5747 , P2_ADD_394_U80 , P2_U2386 );
nand NAND2_9824 ( P2_U5748 , P2_R2278_U85 , P2_U2385 );
nand NAND2_9825 ( P2_U5749 , P2_ADD_371_1212_U82 , P2_U2384 );
nand NAND2_9826 ( P2_U5750 , P2_U2381 , P2_REIP_REG_8_ );
nand NAND2_9827 ( P2_U5751 , P2_INSTADDRPOINTER_REG_8_ , P2_U5673 );
nand NAND2_9828 ( P2_U5752 , P2_R2096_U69 , P2_U2390 );
nand NAND2_9829 ( P2_U5753 , P2_R2099_U67 , P2_U2389 );
nand NAND2_9830 ( P2_U5754 , P2_R2027_U65 , P2_U2388 );
nand NAND2_9831 ( P2_U5755 , P2_ADD_394_U70 , P2_U2386 );
nand NAND2_9832 ( P2_U5756 , P2_R2278_U84 , P2_U2385 );
nand NAND2_9833 ( P2_U5757 , P2_ADD_371_1212_U118 , P2_U2384 );
nand NAND2_9834 ( P2_U5758 , P2_U2381 , P2_REIP_REG_9_ );
nand NAND2_9835 ( P2_U5759 , P2_INSTADDRPOINTER_REG_9_ , P2_U5673 );
nand NAND2_9836 ( P2_U5760 , P2_R2096_U97 , P2_U2390 );
nand NAND2_9837 ( P2_U5761 , P2_R2099_U93 , P2_U2389 );
nand NAND2_9838 ( P2_U5762 , P2_R2027_U95 , P2_U2388 );
nand NAND2_9839 ( P2_U5763 , P2_ADD_394_U83 , P2_U2386 );
nand NAND2_9840 ( P2_U5764 , P2_R2278_U112 , P2_U2385 );
nand NAND2_9841 ( P2_U5765 , P2_ADD_371_1212_U13 , P2_U2384 );
nand NAND2_9842 ( P2_U5766 , P2_U2381 , P2_REIP_REG_10_ );
nand NAND2_9843 ( P2_U5767 , P2_INSTADDRPOINTER_REG_10_ , P2_U5673 );
nand NAND2_9844 ( P2_U5768 , P2_R2096_U96 , P2_U2390 );
nand NAND2_9845 ( P2_U5769 , P2_R2099_U92 , P2_U2389 );
nand NAND2_9846 ( P2_U5770 , P2_R2027_U94 , P2_U2388 );
nand NAND2_9847 ( P2_U5771 , P2_ADD_394_U73 , P2_U2386 );
nand NAND2_9848 ( P2_U5772 , P2_R2278_U111 , P2_U2385 );
nand NAND2_9849 ( P2_U5773 , P2_ADD_371_1212_U14 , P2_U2384 );
nand NAND2_9850 ( P2_U5774 , P2_U2381 , P2_REIP_REG_11_ );
nand NAND2_9851 ( P2_U5775 , P2_INSTADDRPOINTER_REG_11_ , P2_U5673 );
nand NAND2_9852 ( P2_U5776 , P2_R2096_U95 , P2_U2390 );
nand NAND2_9853 ( P2_U5777 , P2_R2099_U91 , P2_U2389 );
nand NAND2_9854 ( P2_U5778 , P2_R2027_U93 , P2_U2388 );
nand NAND2_9855 ( P2_U5779 , P2_ADD_394_U88 , P2_U2386 );
nand NAND2_9856 ( P2_U5780 , P2_R2278_U110 , P2_U2385 );
nand NAND2_9857 ( P2_U5781 , P2_ADD_371_1212_U76 , P2_U2384 );
nand NAND2_9858 ( P2_U5782 , P2_U2381 , P2_REIP_REG_12_ );
nand NAND2_9859 ( P2_U5783 , P2_INSTADDRPOINTER_REG_12_ , P2_U5673 );
nand NAND2_9860 ( P2_U5784 , P2_R2096_U94 , P2_U2390 );
nand NAND2_9861 ( P2_U5785 , P2_R2099_U90 , P2_U2389 );
nand NAND2_9862 ( P2_U5786 , P2_R2027_U92 , P2_U2388 );
nand NAND2_9863 ( P2_U5787 , P2_ADD_394_U69 , P2_U2386 );
nand NAND2_9864 ( P2_U5788 , P2_R2278_U109 , P2_U2385 );
nand NAND2_9865 ( P2_U5789 , P2_ADD_371_1212_U15 , P2_U2384 );
nand NAND2_9866 ( P2_U5790 , P2_U2381 , P2_REIP_REG_13_ );
nand NAND2_9867 ( P2_U5791 , P2_INSTADDRPOINTER_REG_13_ , P2_U5673 );
nand NAND2_9868 ( P2_U5792 , P2_R2096_U93 , P2_U2390 );
nand NAND2_9869 ( P2_U5793 , P2_R2099_U89 , P2_U2389 );
nand NAND2_9870 ( P2_U5794 , P2_R2027_U91 , P2_U2388 );
nand NAND2_9871 ( P2_U5795 , P2_ADD_394_U78 , P2_U2386 );
nand NAND2_9872 ( P2_U5796 , P2_R2278_U108 , P2_U2385 );
nand NAND2_9873 ( P2_U5797 , P2_ADD_371_1212_U16 , P2_U2384 );
nand NAND2_9874 ( P2_U5798 , P2_U2381 , P2_REIP_REG_14_ );
nand NAND2_9875 ( P2_U5799 , P2_INSTADDRPOINTER_REG_14_ , P2_U5673 );
nand NAND2_9876 ( P2_U5800 , P2_R2096_U92 , P2_U2390 );
nand NAND2_9877 ( P2_U5801 , P2_R2099_U88 , P2_U2389 );
nand NAND2_9878 ( P2_U5802 , P2_R2027_U90 , P2_U2388 );
nand NAND2_9879 ( P2_U5803 , P2_ADD_394_U75 , P2_U2386 );
nand NAND2_9880 ( P2_U5804 , P2_R2278_U107 , P2_U2385 );
nand NAND2_9881 ( P2_U5805 , P2_ADD_371_1212_U73 , P2_U2384 );
nand NAND2_9882 ( P2_U5806 , P2_U2381 , P2_REIP_REG_15_ );
nand NAND2_9883 ( P2_U5807 , P2_INSTADDRPOINTER_REG_15_ , P2_U5673 );
nand NAND2_9884 ( P2_U5808 , P2_R2096_U91 , P2_U2390 );
nand NAND2_9885 ( P2_U5809 , P2_R2099_U87 , P2_U2389 );
nand NAND2_9886 ( P2_U5810 , P2_R2027_U89 , P2_U2388 );
nand NAND2_9887 ( P2_U5811 , P2_ADD_394_U91 , P2_U2386 );
nand NAND2_9888 ( P2_U5812 , P2_R2278_U106 , P2_U2385 );
nand NAND2_9889 ( P2_U5813 , P2_ADD_371_1212_U17 , P2_U2384 );
nand NAND2_9890 ( P2_U5814 , P2_U2381 , P2_REIP_REG_16_ );
nand NAND2_9891 ( P2_U5815 , P2_INSTADDRPOINTER_REG_16_ , P2_U5673 );
nand NAND2_9892 ( P2_U5816 , P2_R2096_U90 , P2_U2390 );
nand NAND2_9893 ( P2_U5817 , P2_R2099_U86 , P2_U2389 );
nand NAND2_9894 ( P2_U5818 , P2_R2027_U88 , P2_U2388 );
nand NAND2_9895 ( P2_U5819 , P2_ADD_394_U67 , P2_U2386 );
nand NAND2_9896 ( P2_U5820 , P2_R2278_U105 , P2_U2385 );
nand NAND2_9897 ( P2_U5821 , P2_ADD_371_1212_U71 , P2_U2384 );
nand NAND2_9898 ( P2_U5822 , P2_U2381 , P2_REIP_REG_17_ );
nand NAND2_9899 ( P2_U5823 , P2_INSTADDRPOINTER_REG_17_ , P2_U5673 );
nand NAND2_9900 ( P2_U5824 , P2_R2096_U89 , P2_U2390 );
nand NAND2_9901 ( P2_U5825 , P2_R2099_U85 , P2_U2389 );
nand NAND2_9902 ( P2_U5826 , P2_R2027_U87 , P2_U2388 );
nand NAND2_9903 ( P2_U5827 , P2_ADD_394_U72 , P2_U2386 );
nand NAND2_9904 ( P2_U5828 , P2_R2278_U104 , P2_U2385 );
nand NAND2_9905 ( P2_U5829 , P2_ADD_371_1212_U72 , P2_U2384 );
nand NAND2_9906 ( P2_U5830 , P2_U2381 , P2_REIP_REG_18_ );
nand NAND2_9907 ( P2_U5831 , P2_INSTADDRPOINTER_REG_18_ , P2_U5673 );
nand NAND2_9908 ( P2_U5832 , P2_R2096_U88 , P2_U2390 );
nand NAND2_9909 ( P2_U5833 , P2_R2099_U84 , P2_U2389 );
nand NAND2_9910 ( P2_U5834 , P2_R2027_U86 , P2_U2388 );
nand NAND2_9911 ( P2_U5835 , P2_ADD_394_U82 , P2_U2386 );
nand NAND2_9912 ( P2_U5836 , P2_R2278_U103 , P2_U2385 );
nand NAND2_9913 ( P2_U5837 , P2_ADD_371_1212_U18 , P2_U2384 );
nand NAND2_9914 ( P2_U5838 , P2_U2381 , P2_REIP_REG_19_ );
nand NAND2_9915 ( P2_U5839 , P2_INSTADDRPOINTER_REG_19_ , P2_U5673 );
nand NAND2_9916 ( P2_U5840 , P2_R2096_U87 , P2_U2390 );
nand NAND2_9917 ( P2_U5841 , P2_R2099_U83 , P2_U2389 );
nand NAND2_9918 ( P2_U5842 , P2_R2027_U84 , P2_U2388 );
nand NAND2_9919 ( P2_U5843 , P2_ADD_394_U68 , P2_U2386 );
nand NAND2_9920 ( P2_U5844 , P2_R2278_U102 , P2_U2385 );
nand NAND2_9921 ( P2_U5845 , P2_ADD_371_1212_U19 , P2_U2384 );
nand NAND2_9922 ( P2_U5846 , P2_U2381 , P2_REIP_REG_20_ );
nand NAND2_9923 ( P2_U5847 , P2_INSTADDRPOINTER_REG_20_ , P2_U5673 );
nand NAND2_9924 ( P2_U5848 , P2_R2096_U86 , P2_U2390 );
nand NAND2_9925 ( P2_U5849 , P2_R2099_U82 , P2_U2389 );
nand NAND2_9926 ( P2_U5850 , P2_R2027_U83 , P2_U2388 );
nand NAND2_9927 ( P2_U5851 , P2_ADD_394_U87 , P2_U2386 );
nand NAND2_9928 ( P2_U5852 , P2_R2278_U101 , P2_U2385 );
nand NAND2_9929 ( P2_U5853 , P2_ADD_371_1212_U75 , P2_U2384 );
nand NAND2_9930 ( P2_U5854 , P2_U2381 , P2_REIP_REG_21_ );
nand NAND2_9931 ( P2_U5855 , P2_INSTADDRPOINTER_REG_21_ , P2_U5673 );
nand NAND2_9932 ( P2_U5856 , P2_R2096_U85 , P2_U2390 );
nand NAND2_9933 ( P2_U5857 , P2_R2099_U81 , P2_U2389 );
nand NAND2_9934 ( P2_U5858 , P2_R2027_U82 , P2_U2388 );
nand NAND2_9935 ( P2_U5859 , P2_ADD_394_U71 , P2_U2386 );
nand NAND2_9936 ( P2_U5860 , P2_R2278_U100 , P2_U2385 );
nand NAND2_9937 ( P2_U5861 , P2_ADD_371_1212_U20 , P2_U2384 );
nand NAND2_9938 ( P2_U5862 , P2_U2381 , P2_REIP_REG_22_ );
nand NAND2_9939 ( P2_U5863 , P2_INSTADDRPOINTER_REG_22_ , P2_U5673 );
nand NAND2_9940 ( P2_U5864 , P2_R2096_U84 , P2_U2390 );
nand NAND2_9941 ( P2_U5865 , P2_R2099_U80 , P2_U2389 );
nand NAND2_9942 ( P2_U5866 , P2_R2027_U81 , P2_U2388 );
nand NAND2_9943 ( P2_U5867 , P2_ADD_394_U81 , P2_U2386 );
nand NAND2_9944 ( P2_U5868 , P2_R2278_U99 , P2_U2385 );
nand NAND2_9945 ( P2_U5869 , P2_ADD_371_1212_U21 , P2_U2384 );
nand NAND2_9946 ( P2_U5870 , P2_U2381 , P2_REIP_REG_23_ );
nand NAND2_9947 ( P2_U5871 , P2_INSTADDRPOINTER_REG_23_ , P2_U5673 );
nand NAND2_9948 ( P2_U5872 , P2_R2096_U83 , P2_U2390 );
nand NAND2_9949 ( P2_U5873 , P2_R2099_U79 , P2_U2389 );
nand NAND2_9950 ( P2_U5874 , P2_R2027_U80 , P2_U2388 );
nand NAND2_9951 ( P2_U5875 , P2_ADD_394_U66 , P2_U2386 );
nand NAND2_9952 ( P2_U5876 , P2_R2278_U98 , P2_U2385 );
nand NAND2_9953 ( P2_U5877 , P2_ADD_371_1212_U70 , P2_U2384 );
nand NAND2_9954 ( P2_U5878 , P2_U2381 , P2_REIP_REG_24_ );
nand NAND2_9955 ( P2_U5879 , P2_INSTADDRPOINTER_REG_24_ , P2_U5673 );
nand NAND2_9956 ( P2_U5880 , P2_R2096_U82 , P2_U2390 );
nand NAND2_9957 ( P2_U5881 , P2_R2099_U78 , P2_U2389 );
nand NAND2_9958 ( P2_U5882 , P2_R2027_U79 , P2_U2388 );
nand NAND2_9959 ( P2_U5883 , P2_ADD_394_U90 , P2_U2386 );
nand NAND2_9960 ( P2_U5884 , P2_R2278_U97 , P2_U2385 );
nand NAND2_9961 ( P2_U5885 , P2_ADD_371_1212_U77 , P2_U2384 );
nand NAND2_9962 ( P2_U5886 , P2_U2381 , P2_REIP_REG_25_ );
nand NAND2_9963 ( P2_U5887 , P2_INSTADDRPOINTER_REG_25_ , P2_U5673 );
nand NAND2_9964 ( P2_U5888 , P2_R2096_U81 , P2_U2390 );
nand NAND2_9965 ( P2_U5889 , P2_R2099_U77 , P2_U2389 );
nand NAND2_9966 ( P2_U5890 , P2_R2027_U78 , P2_U2388 );
nand NAND2_9967 ( P2_U5891 , P2_ADD_394_U74 , P2_U2386 );
nand NAND2_9968 ( P2_U5892 , P2_R2278_U96 , P2_U2385 );
nand NAND2_9969 ( P2_U5893 , P2_ADD_371_1212_U22 , P2_U2384 );
nand NAND2_9970 ( P2_U5894 , P2_U2381 , P2_REIP_REG_26_ );
nand NAND2_9971 ( P2_U5895 , P2_INSTADDRPOINTER_REG_26_ , P2_U5673 );
nand NAND2_9972 ( P2_U5896 , P2_R2096_U80 , P2_U2390 );
nand NAND2_9973 ( P2_U5897 , P2_R2099_U76 , P2_U2389 );
nand NAND2_9974 ( P2_U5898 , P2_R2027_U77 , P2_U2388 );
nand NAND2_9975 ( P2_U5899 , P2_ADD_394_U77 , P2_U2386 );
nand NAND2_9976 ( P2_U5900 , P2_R2278_U95 , P2_U2385 );
nand NAND2_9977 ( P2_U5901 , P2_ADD_371_1212_U74 , P2_U2384 );
nand NAND2_9978 ( P2_U5902 , P2_U2381 , P2_REIP_REG_27_ );
nand NAND2_9979 ( P2_U5903 , P2_INSTADDRPOINTER_REG_27_ , P2_U5673 );
nand NAND2_9980 ( P2_U5904 , P2_R2096_U79 , P2_U2390 );
nand NAND2_9981 ( P2_U5905 , P2_R2099_U75 , P2_U2389 );
nand NAND2_9982 ( P2_U5906 , P2_R2027_U76 , P2_U2388 );
nand NAND2_9983 ( P2_U5907 , P2_ADD_394_U86 , P2_U2386 );
nand NAND2_9984 ( P2_U5908 , P2_R2278_U94 , P2_U2385 );
nand NAND2_9985 ( P2_U5909 , P2_ADD_371_1212_U23 , P2_U2384 );
nand NAND2_9986 ( P2_U5910 , P2_U2381 , P2_REIP_REG_28_ );
nand NAND2_9987 ( P2_U5911 , P2_INSTADDRPOINTER_REG_28_ , P2_U5673 );
nand NAND2_9988 ( P2_U5912 , P2_R2096_U78 , P2_U2390 );
nand NAND2_9989 ( P2_U5913 , P2_R2099_U74 , P2_U2389 );
nand NAND2_9990 ( P2_U5914 , P2_R2027_U75 , P2_U2388 );
nand NAND2_9991 ( P2_U5915 , P2_ADD_394_U65 , P2_U2386 );
nand NAND2_9992 ( P2_U5916 , P2_R2278_U93 , P2_U2385 );
nand NAND2_9993 ( P2_U5917 , P2_ADD_371_1212_U24 , P2_U2384 );
nand NAND2_9994 ( P2_U5918 , P2_U2381 , P2_REIP_REG_29_ );
nand NAND2_9995 ( P2_U5919 , P2_INSTADDRPOINTER_REG_29_ , P2_U5673 );
nand NAND2_9996 ( P2_U5920 , P2_R2096_U76 , P2_U2390 );
nand NAND2_9997 ( P2_U5921 , P2_R2099_U73 , P2_U2389 );
nand NAND2_9998 ( P2_U5922 , P2_R2027_U73 , P2_U2388 );
nand NAND2_9999 ( P2_U5923 , P2_ADD_394_U64 , P2_U2386 );
nand NAND2_10000 ( P2_U5924 , P2_R2278_U91 , P2_U2385 );
nand NAND2_10001 ( P2_U5925 , P2_ADD_371_1212_U69 , P2_U2384 );
nand NAND2_10002 ( P2_U5926 , P2_U2381 , P2_REIP_REG_30_ );
nand NAND2_10003 ( P2_U5927 , P2_INSTADDRPOINTER_REG_30_ , P2_U5673 );
nand NAND2_10004 ( P2_U5928 , P2_R2096_U50 , P2_U2390 );
nand NAND2_10005 ( P2_U5929 , P2_R2099_U72 , P2_U2389 );
nand NAND2_10006 ( P2_U5930 , P2_R2027_U72 , P2_U2388 );
nand NAND2_10007 ( P2_U5931 , P2_ADD_394_U84 , P2_U2386 );
nand NAND2_10008 ( P2_U5932 , P2_R2278_U5 , P2_U2385 );
nand NAND2_10009 ( P2_U5933 , P2_ADD_371_1212_U83 , P2_U2384 );
nand NAND2_10010 ( P2_U5934 , P2_U2381 , P2_REIP_REG_31_ );
nand NAND2_10011 ( P2_U5935 , P2_INSTADDRPOINTER_REG_31_ , P2_U5673 );
nand NAND3_10012 ( P2_U5936 , P2_U4420 , P2_U2374 , P2_U4613 );
nand NAND2_10013 ( P2_U5937 , P2_U5661 , P2_U3284 );
not NOT1_10014 ( P2_U5938 , P2_U3537 );
nand NAND2_10015 ( P2_U5939 , P2_STATE2_REG_1_ , P2_U3302 );
nand NAND2_10016 ( P2_U5940 , P2_U3540 , P2_U5939 );
nand NAND2_10017 ( P2_U5941 , P2_PHYADDRPOINTER_REG_0_ , P2_U2387 );
nand NAND2_10018 ( P2_U5942 , P2_U2373 , P2_ADD_371_1212_U68 );
nand NAND2_10019 ( P2_U5943 , P2_U2372 , P2_R2099_U94 );
nand NAND2_10020 ( P2_U5944 , P2_U2371 , P2_REIP_REG_0_ );
nand NAND2_10021 ( P2_U5945 , P2_U2370 , P2_R2278_U83 );
nand NAND2_10022 ( P2_U5946 , P2_PHYADDRPOINTER_REG_0_ , P2_U5938 );
nand NAND2_10023 ( P2_U5947 , P2_R2337_U4 , P2_U2387 );
nand NAND2_10024 ( P2_U5948 , P2_U2373 , P2_ADD_371_1212_U25 );
nand NAND2_10025 ( P2_U5949 , P2_U2372 , P2_R2099_U5 );
nand NAND2_10026 ( P2_U5950 , P2_U2371 , P2_REIP_REG_1_ );
nand NAND2_10027 ( P2_U5951 , P2_U2370 , P2_R2278_U6 );
nand NAND2_10028 ( P2_U5952 , P2_PHYADDRPOINTER_REG_1_ , P2_U5938 );
nand NAND2_10029 ( P2_U5953 , P2_R2337_U70 , P2_U2387 );
nand NAND2_10030 ( P2_U5954 , P2_U2373 , P2_ADD_371_1212_U79 );
nand NAND2_10031 ( P2_U5955 , P2_U2372 , P2_R2099_U96 );
nand NAND2_10032 ( P2_U5956 , P2_U2371 , P2_REIP_REG_2_ );
nand NAND2_10033 ( P2_U5957 , P2_U2370 , P2_R2278_U92 );
nand NAND2_10034 ( P2_U5958 , P2_PHYADDRPOINTER_REG_2_ , P2_U5938 );
nand NAND2_10035 ( P2_U5959 , P2_R2337_U67 , P2_U2387 );
nand NAND2_10036 ( P2_U5960 , P2_U2373 , P2_ADD_371_1212_U84 );
nand NAND2_10037 ( P2_U5961 , P2_U2372 , P2_R2099_U95 );
nand NAND2_10038 ( P2_U5962 , P2_U2371 , P2_REIP_REG_3_ );
nand NAND2_10039 ( P2_U5963 , P2_U2370 , P2_R2278_U90 );
nand NAND2_10040 ( P2_U5964 , P2_PHYADDRPOINTER_REG_3_ , P2_U5938 );
nand NAND2_10041 ( P2_U5965 , P2_R2337_U66 , P2_U2387 );
nand NAND2_10042 ( P2_U5966 , P2_U2373 , P2_ADD_371_1212_U80 );
nand NAND2_10043 ( P2_U5967 , P2_U2372 , P2_R2099_U98 );
nand NAND2_10044 ( P2_U5968 , P2_U2371 , P2_REIP_REG_4_ );
nand NAND2_10045 ( P2_U5969 , P2_U2370 , P2_R2278_U89 );
nand NAND2_10046 ( P2_U5970 , P2_PHYADDRPOINTER_REG_4_ , P2_U5938 );
nand NAND2_10047 ( P2_U5971 , P2_R2337_U65 , P2_U2387 );
nand NAND2_10048 ( P2_U5972 , P2_U2373 , P2_ADD_371_1212_U81 );
nand NAND2_10049 ( P2_U5973 , P2_U2372 , P2_R2099_U71 );
nand NAND2_10050 ( P2_U5974 , P2_U2371 , P2_REIP_REG_5_ );
nand NAND2_10051 ( P2_U5975 , P2_U2370 , P2_R2278_U88 );
nand NAND2_10052 ( P2_U5976 , P2_PHYADDRPOINTER_REG_5_ , P2_U5938 );
nand NAND2_10053 ( P2_U5977 , P2_R2337_U64 , P2_U2387 );
nand NAND2_10054 ( P2_U5978 , P2_U2373 , P2_ADD_371_1212_U78 );
nand NAND2_10055 ( P2_U5979 , P2_U2372 , P2_R2099_U70 );
nand NAND2_10056 ( P2_U5980 , P2_U2371 , P2_REIP_REG_6_ );
nand NAND2_10057 ( P2_U5981 , P2_U2370 , P2_R2278_U87 );
nand NAND2_10058 ( P2_U5982 , P2_PHYADDRPOINTER_REG_6_ , P2_U5938 );
nand NAND2_10059 ( P2_U5983 , P2_R2337_U63 , P2_U2387 );
nand NAND2_10060 ( P2_U5984 , P2_U2373 , P2_ADD_371_1212_U85 );
nand NAND2_10061 ( P2_U5985 , P2_U2372 , P2_R2099_U69 );
nand NAND2_10062 ( P2_U5986 , P2_U2371 , P2_REIP_REG_7_ );
nand NAND2_10063 ( P2_U5987 , P2_U2370 , P2_R2278_U86 );
nand NAND2_10064 ( P2_U5988 , P2_PHYADDRPOINTER_REG_7_ , P2_U5938 );
nand NAND2_10065 ( P2_U5989 , P2_R2337_U62 , P2_U2387 );
nand NAND2_10066 ( P2_U5990 , P2_U2373 , P2_ADD_371_1212_U82 );
nand NAND2_10067 ( P2_U5991 , P2_U2372 , P2_R2099_U68 );
nand NAND2_10068 ( P2_U5992 , P2_U2371 , P2_REIP_REG_8_ );
nand NAND2_10069 ( P2_U5993 , P2_U2370 , P2_R2278_U85 );
nand NAND2_10070 ( P2_U5994 , P2_PHYADDRPOINTER_REG_8_ , P2_U5938 );
nand NAND2_10071 ( P2_U5995 , P2_R2337_U61 , P2_U2387 );
nand NAND2_10072 ( P2_U5996 , P2_U2373 , P2_ADD_371_1212_U118 );
nand NAND2_10073 ( P2_U5997 , P2_U2372 , P2_R2099_U67 );
nand NAND2_10074 ( P2_U5998 , P2_U2371 , P2_REIP_REG_9_ );
nand NAND2_10075 ( P2_U5999 , P2_U2370 , P2_R2278_U84 );
nand NAND2_10076 ( P2_U6000 , P2_PHYADDRPOINTER_REG_9_ , P2_U5938 );
nand NAND2_10077 ( P2_U6001 , P2_R2337_U90 , P2_U2387 );
nand NAND2_10078 ( P2_U6002 , P2_U2373 , P2_ADD_371_1212_U13 );
nand NAND2_10079 ( P2_U6003 , P2_U2372 , P2_R2099_U93 );
nand NAND2_10080 ( P2_U6004 , P2_U2371 , P2_REIP_REG_10_ );
nand NAND2_10081 ( P2_U6005 , P2_U2370 , P2_R2278_U112 );
nand NAND2_10082 ( P2_U6006 , P2_PHYADDRPOINTER_REG_10_ , P2_U5938 );
nand NAND2_10083 ( P2_U6007 , P2_R2337_U89 , P2_U2387 );
nand NAND2_10084 ( P2_U6008 , P2_U2373 , P2_ADD_371_1212_U14 );
nand NAND2_10085 ( P2_U6009 , P2_U2372 , P2_R2099_U92 );
nand NAND2_10086 ( P2_U6010 , P2_U2371 , P2_REIP_REG_11_ );
nand NAND2_10087 ( P2_U6011 , P2_U2370 , P2_R2278_U111 );
nand NAND2_10088 ( P2_U6012 , P2_PHYADDRPOINTER_REG_11_ , P2_U5938 );
nand NAND2_10089 ( P2_U6013 , P2_R2337_U88 , P2_U2387 );
nand NAND2_10090 ( P2_U6014 , P2_U2373 , P2_ADD_371_1212_U76 );
nand NAND2_10091 ( P2_U6015 , P2_U2372 , P2_R2099_U91 );
nand NAND2_10092 ( P2_U6016 , P2_U2371 , P2_REIP_REG_12_ );
nand NAND2_10093 ( P2_U6017 , P2_U2370 , P2_R2278_U110 );
nand NAND2_10094 ( P2_U6018 , P2_PHYADDRPOINTER_REG_12_ , P2_U5938 );
nand NAND2_10095 ( P2_U6019 , P2_R2337_U87 , P2_U2387 );
nand NAND2_10096 ( P2_U6020 , P2_U2373 , P2_ADD_371_1212_U15 );
nand NAND2_10097 ( P2_U6021 , P2_U2372 , P2_R2099_U90 );
nand NAND2_10098 ( P2_U6022 , P2_U2371 , P2_REIP_REG_13_ );
nand NAND2_10099 ( P2_U6023 , P2_U2370 , P2_R2278_U109 );
nand NAND2_10100 ( P2_U6024 , P2_PHYADDRPOINTER_REG_13_ , P2_U5938 );
nand NAND2_10101 ( P2_U6025 , P2_R2337_U86 , P2_U2387 );
nand NAND2_10102 ( P2_U6026 , P2_U2373 , P2_ADD_371_1212_U16 );
nand NAND2_10103 ( P2_U6027 , P2_U2372 , P2_R2099_U89 );
nand NAND2_10104 ( P2_U6028 , P2_U2371 , P2_REIP_REG_14_ );
nand NAND2_10105 ( P2_U6029 , P2_U2370 , P2_R2278_U108 );
nand NAND2_10106 ( P2_U6030 , P2_PHYADDRPOINTER_REG_14_ , P2_U5938 );
nand NAND2_10107 ( P2_U6031 , P2_R2337_U85 , P2_U2387 );
nand NAND2_10108 ( P2_U6032 , P2_U2373 , P2_ADD_371_1212_U73 );
nand NAND2_10109 ( P2_U6033 , P2_U2372 , P2_R2099_U88 );
nand NAND2_10110 ( P2_U6034 , P2_U2371 , P2_REIP_REG_15_ );
nand NAND2_10111 ( P2_U6035 , P2_U2370 , P2_R2278_U107 );
nand NAND2_10112 ( P2_U6036 , P2_PHYADDRPOINTER_REG_15_ , P2_U5938 );
nand NAND2_10113 ( P2_U6037 , P2_R2337_U84 , P2_U2387 );
nand NAND2_10114 ( P2_U6038 , P2_U2373 , P2_ADD_371_1212_U17 );
nand NAND2_10115 ( P2_U6039 , P2_U2372 , P2_R2099_U87 );
nand NAND2_10116 ( P2_U6040 , P2_U2371 , P2_REIP_REG_16_ );
nand NAND2_10117 ( P2_U6041 , P2_U2370 , P2_R2278_U106 );
nand NAND2_10118 ( P2_U6042 , P2_PHYADDRPOINTER_REG_16_ , P2_U5938 );
nand NAND2_10119 ( P2_U6043 , P2_R2337_U83 , P2_U2387 );
nand NAND2_10120 ( P2_U6044 , P2_U2373 , P2_ADD_371_1212_U71 );
nand NAND2_10121 ( P2_U6045 , P2_U2372 , P2_R2099_U86 );
nand NAND2_10122 ( P2_U6046 , P2_U2371 , P2_REIP_REG_17_ );
nand NAND2_10123 ( P2_U6047 , P2_U2370 , P2_R2278_U105 );
nand NAND2_10124 ( P2_U6048 , P2_PHYADDRPOINTER_REG_17_ , P2_U5938 );
nand NAND2_10125 ( P2_U6049 , P2_R2337_U82 , P2_U2387 );
nand NAND2_10126 ( P2_U6050 , P2_U2373 , P2_ADD_371_1212_U72 );
nand NAND2_10127 ( P2_U6051 , P2_U2372 , P2_R2099_U85 );
nand NAND2_10128 ( P2_U6052 , P2_U2371 , P2_REIP_REG_18_ );
nand NAND2_10129 ( P2_U6053 , P2_U2370 , P2_R2278_U104 );
nand NAND2_10130 ( P2_U6054 , P2_PHYADDRPOINTER_REG_18_ , P2_U5938 );
nand NAND2_10131 ( P2_U6055 , P2_R2337_U81 , P2_U2387 );
nand NAND2_10132 ( P2_U6056 , P2_U2373 , P2_ADD_371_1212_U18 );
nand NAND2_10133 ( P2_U6057 , P2_U2372 , P2_R2099_U84 );
nand NAND2_10134 ( P2_U6058 , P2_U2371 , P2_REIP_REG_19_ );
nand NAND2_10135 ( P2_U6059 , P2_U2370 , P2_R2278_U103 );
nand NAND2_10136 ( P2_U6060 , P2_PHYADDRPOINTER_REG_19_ , P2_U5938 );
nand NAND2_10137 ( P2_U6061 , P2_R2337_U80 , P2_U2387 );
nand NAND2_10138 ( P2_U6062 , P2_U2373 , P2_ADD_371_1212_U19 );
nand NAND2_10139 ( P2_U6063 , P2_U2372 , P2_R2099_U83 );
nand NAND2_10140 ( P2_U6064 , P2_U2371 , P2_REIP_REG_20_ );
nand NAND2_10141 ( P2_U6065 , P2_U2370 , P2_R2278_U102 );
nand NAND2_10142 ( P2_U6066 , P2_PHYADDRPOINTER_REG_20_ , P2_U5938 );
nand NAND2_10143 ( P2_U6067 , P2_R2337_U79 , P2_U2387 );
nand NAND2_10144 ( P2_U6068 , P2_U2373 , P2_ADD_371_1212_U75 );
nand NAND2_10145 ( P2_U6069 , P2_U2372 , P2_R2099_U82 );
nand NAND2_10146 ( P2_U6070 , P2_U2371 , P2_REIP_REG_21_ );
nand NAND2_10147 ( P2_U6071 , P2_U2370 , P2_R2278_U101 );
nand NAND2_10148 ( P2_U6072 , P2_PHYADDRPOINTER_REG_21_ , P2_U5938 );
nand NAND2_10149 ( P2_U6073 , P2_R2337_U78 , P2_U2387 );
nand NAND2_10150 ( P2_U6074 , P2_U2373 , P2_ADD_371_1212_U20 );
nand NAND2_10151 ( P2_U6075 , P2_U2372 , P2_R2099_U81 );
nand NAND2_10152 ( P2_U6076 , P2_U2371 , P2_REIP_REG_22_ );
nand NAND2_10153 ( P2_U6077 , P2_U2370 , P2_R2278_U100 );
nand NAND2_10154 ( P2_U6078 , P2_PHYADDRPOINTER_REG_22_ , P2_U5938 );
nand NAND2_10155 ( P2_U6079 , P2_R2337_U77 , P2_U2387 );
nand NAND2_10156 ( P2_U6080 , P2_U2373 , P2_ADD_371_1212_U21 );
nand NAND2_10157 ( P2_U6081 , P2_U2372 , P2_R2099_U80 );
nand NAND2_10158 ( P2_U6082 , P2_U2371 , P2_REIP_REG_23_ );
nand NAND2_10159 ( P2_U6083 , P2_U2370 , P2_R2278_U99 );
nand NAND2_10160 ( P2_U6084 , P2_PHYADDRPOINTER_REG_23_ , P2_U5938 );
nand NAND2_10161 ( P2_U6085 , P2_R2337_U76 , P2_U2387 );
nand NAND2_10162 ( P2_U6086 , P2_U2373 , P2_ADD_371_1212_U70 );
nand NAND2_10163 ( P2_U6087 , P2_U2372 , P2_R2099_U79 );
nand NAND2_10164 ( P2_U6088 , P2_U2371 , P2_REIP_REG_24_ );
nand NAND2_10165 ( P2_U6089 , P2_U2370 , P2_R2278_U98 );
nand NAND2_10166 ( P2_U6090 , P2_PHYADDRPOINTER_REG_24_ , P2_U5938 );
nand NAND2_10167 ( P2_U6091 , P2_R2337_U75 , P2_U2387 );
nand NAND2_10168 ( P2_U6092 , P2_U2373 , P2_ADD_371_1212_U77 );
nand NAND2_10169 ( P2_U6093 , P2_U2372 , P2_R2099_U78 );
nand NAND2_10170 ( P2_U6094 , P2_U2371 , P2_REIP_REG_25_ );
nand NAND2_10171 ( P2_U6095 , P2_U2370 , P2_R2278_U97 );
nand NAND2_10172 ( P2_U6096 , P2_PHYADDRPOINTER_REG_25_ , P2_U5938 );
nand NAND2_10173 ( P2_U6097 , P2_R2337_U74 , P2_U2387 );
nand NAND2_10174 ( P2_U6098 , P2_U2373 , P2_ADD_371_1212_U22 );
nand NAND2_10175 ( P2_U6099 , P2_U2372 , P2_R2099_U77 );
nand NAND2_10176 ( P2_U6100 , P2_U2371 , P2_REIP_REG_26_ );
nand NAND2_10177 ( P2_U6101 , P2_U2370 , P2_R2278_U96 );
nand NAND2_10178 ( P2_U6102 , P2_PHYADDRPOINTER_REG_26_ , P2_U5938 );
nand NAND2_10179 ( P2_U6103 , P2_R2337_U73 , P2_U2387 );
nand NAND2_10180 ( P2_U6104 , P2_U2373 , P2_ADD_371_1212_U74 );
nand NAND2_10181 ( P2_U6105 , P2_U2372 , P2_R2099_U76 );
nand NAND2_10182 ( P2_U6106 , P2_U2371 , P2_REIP_REG_27_ );
nand NAND2_10183 ( P2_U6107 , P2_U2370 , P2_R2278_U95 );
nand NAND2_10184 ( P2_U6108 , P2_PHYADDRPOINTER_REG_27_ , P2_U5938 );
nand NAND2_10185 ( P2_U6109 , P2_R2337_U72 , P2_U2387 );
nand NAND2_10186 ( P2_U6110 , P2_U2373 , P2_ADD_371_1212_U23 );
nand NAND2_10187 ( P2_U6111 , P2_U2372 , P2_R2099_U75 );
nand NAND2_10188 ( P2_U6112 , P2_U2371 , P2_REIP_REG_28_ );
nand NAND2_10189 ( P2_U6113 , P2_U2370 , P2_R2278_U94 );
nand NAND2_10190 ( P2_U6114 , P2_PHYADDRPOINTER_REG_28_ , P2_U5938 );
nand NAND2_10191 ( P2_U6115 , P2_R2337_U71 , P2_U2387 );
nand NAND2_10192 ( P2_U6116 , P2_U2373 , P2_ADD_371_1212_U24 );
nand NAND2_10193 ( P2_U6117 , P2_U2372 , P2_R2099_U74 );
nand NAND2_10194 ( P2_U6118 , P2_U2371 , P2_REIP_REG_29_ );
nand NAND2_10195 ( P2_U6119 , P2_U2370 , P2_R2278_U93 );
nand NAND2_10196 ( P2_U6120 , P2_PHYADDRPOINTER_REG_29_ , P2_U5938 );
nand NAND2_10197 ( P2_U6121 , P2_R2337_U69 , P2_U2387 );
nand NAND2_10198 ( P2_U6122 , P2_U2373 , P2_ADD_371_1212_U69 );
nand NAND2_10199 ( P2_U6123 , P2_U2372 , P2_R2099_U73 );
nand NAND2_10200 ( P2_U6124 , P2_U2371 , P2_REIP_REG_30_ );
nand NAND2_10201 ( P2_U6125 , P2_U2370 , P2_R2278_U91 );
nand NAND2_10202 ( P2_U6126 , P2_PHYADDRPOINTER_REG_30_ , P2_U5938 );
nand NAND2_10203 ( P2_U6127 , P2_R2337_U68 , P2_U2387 );
nand NAND2_10204 ( P2_U6128 , P2_U2373 , P2_ADD_371_1212_U83 );
nand NAND2_10205 ( P2_U6129 , P2_U2372 , P2_R2099_U72 );
nand NAND2_10206 ( P2_U6130 , P2_U2371 , P2_REIP_REG_31_ );
nand NAND2_10207 ( P2_U6131 , P2_U2370 , P2_R2278_U5 );
nand NAND2_10208 ( P2_U6132 , P2_PHYADDRPOINTER_REG_31_ , P2_U5938 );
nand NAND2_10209 ( P2_U6133 , U211 , P2_U2616 );
nand NAND2_10210 ( P2_U6134 , P2_EAX_REG_15_ , P2_U2395 );
nand NAND2_10211 ( P2_U6135 , U308 , P2_U2394 );
nand NAND2_10212 ( P2_U6136 , P2_LWORD_REG_15_ , P2_U3538 );
nand NAND2_10213 ( P2_U6137 , P2_EAX_REG_14_ , P2_U2395 );
nand NAND2_10214 ( P2_U6138 , U309 , P2_U2394 );
nand NAND2_10215 ( P2_U6139 , P2_LWORD_REG_14_ , P2_U3538 );
nand NAND2_10216 ( P2_U6140 , P2_EAX_REG_13_ , P2_U2395 );
nand NAND2_10217 ( P2_U6141 , U310 , P2_U2394 );
nand NAND2_10218 ( P2_U6142 , P2_LWORD_REG_13_ , P2_U3538 );
nand NAND2_10219 ( P2_U6143 , P2_EAX_REG_12_ , P2_U2395 );
nand NAND2_10220 ( P2_U6144 , U311 , P2_U2394 );
nand NAND2_10221 ( P2_U6145 , P2_LWORD_REG_12_ , P2_U3538 );
nand NAND2_10222 ( P2_U6146 , P2_EAX_REG_11_ , P2_U2395 );
nand NAND2_10223 ( P2_U6147 , U312 , P2_U2394 );
nand NAND2_10224 ( P2_U6148 , P2_LWORD_REG_11_ , P2_U3538 );
nand NAND2_10225 ( P2_U6149 , P2_EAX_REG_10_ , P2_U2395 );
nand NAND2_10226 ( P2_U6150 , U313 , P2_U2394 );
nand NAND2_10227 ( P2_U6151 , P2_LWORD_REG_10_ , P2_U3538 );
nand NAND2_10228 ( P2_U6152 , P2_EAX_REG_9_ , P2_U2395 );
nand NAND2_10229 ( P2_U6153 , U283 , P2_U2394 );
nand NAND2_10230 ( P2_U6154 , P2_LWORD_REG_9_ , P2_U3538 );
nand NAND2_10231 ( P2_U6155 , P2_EAX_REG_8_ , P2_U2395 );
nand NAND2_10232 ( P2_U6156 , U284 , P2_U2394 );
nand NAND2_10233 ( P2_U6157 , P2_LWORD_REG_8_ , P2_U3538 );
nand NAND2_10234 ( P2_U6158 , P2_EAX_REG_7_ , P2_U2395 );
nand NAND2_10235 ( P2_U6159 , P2_U2394 , U285 );
nand NAND2_10236 ( P2_U6160 , P2_LWORD_REG_7_ , P2_U3538 );
nand NAND2_10237 ( P2_U6161 , P2_EAX_REG_6_ , P2_U2395 );
nand NAND2_10238 ( P2_U6162 , P2_U2394 , U286 );
nand NAND2_10239 ( P2_U6163 , P2_LWORD_REG_6_ , P2_U3538 );
nand NAND2_10240 ( P2_U6164 , P2_EAX_REG_5_ , P2_U2395 );
nand NAND2_10241 ( P2_U6165 , P2_U2394 , U287 );
nand NAND2_10242 ( P2_U6166 , P2_LWORD_REG_5_ , P2_U3538 );
nand NAND2_10243 ( P2_U6167 , P2_EAX_REG_4_ , P2_U2395 );
nand NAND2_10244 ( P2_U6168 , P2_U2394 , U288 );
nand NAND2_10245 ( P2_U6169 , P2_LWORD_REG_4_ , P2_U3538 );
nand NAND2_10246 ( P2_U6170 , P2_EAX_REG_3_ , P2_U2395 );
nand NAND2_10247 ( P2_U6171 , P2_U2394 , U289 );
nand NAND2_10248 ( P2_U6172 , P2_LWORD_REG_3_ , P2_U3538 );
nand NAND2_10249 ( P2_U6173 , P2_EAX_REG_2_ , P2_U2395 );
nand NAND2_10250 ( P2_U6174 , P2_U2394 , U292 );
nand NAND2_10251 ( P2_U6175 , P2_LWORD_REG_2_ , P2_U3538 );
nand NAND2_10252 ( P2_U6176 , P2_EAX_REG_1_ , P2_U2395 );
nand NAND2_10253 ( P2_U6177 , P2_U2394 , U303 );
nand NAND2_10254 ( P2_U6178 , P2_LWORD_REG_1_ , P2_U3538 );
nand NAND2_10255 ( P2_U6179 , P2_EAX_REG_0_ , P2_U2395 );
nand NAND2_10256 ( P2_U6180 , P2_U2394 , U314 );
nand NAND2_10257 ( P2_U6181 , P2_LWORD_REG_0_ , P2_U3538 );
nand NAND2_10258 ( P2_U6182 , P2_EAX_REG_30_ , P2_U2395 );
nand NAND2_10259 ( P2_U6183 , U309 , P2_U2394 );
nand NAND2_10260 ( P2_U6184 , P2_UWORD_REG_14_ , P2_U3538 );
nand NAND2_10261 ( P2_U6185 , P2_EAX_REG_29_ , P2_U2395 );
nand NAND2_10262 ( P2_U6186 , U310 , P2_U2394 );
nand NAND2_10263 ( P2_U6187 , P2_UWORD_REG_13_ , P2_U3538 );
nand NAND2_10264 ( P2_U6188 , P2_EAX_REG_28_ , P2_U2395 );
nand NAND2_10265 ( P2_U6189 , U311 , P2_U2394 );
nand NAND2_10266 ( P2_U6190 , P2_UWORD_REG_12_ , P2_U3538 );
nand NAND2_10267 ( P2_U6191 , P2_EAX_REG_27_ , P2_U2395 );
nand NAND2_10268 ( P2_U6192 , U312 , P2_U2394 );
nand NAND2_10269 ( P2_U6193 , P2_UWORD_REG_11_ , P2_U3538 );
nand NAND2_10270 ( P2_U6194 , P2_EAX_REG_26_ , P2_U2395 );
nand NAND2_10271 ( P2_U6195 , U313 , P2_U2394 );
nand NAND2_10272 ( P2_U6196 , P2_UWORD_REG_10_ , P2_U3538 );
nand NAND2_10273 ( P2_U6197 , P2_EAX_REG_25_ , P2_U2395 );
nand NAND2_10274 ( P2_U6198 , U283 , P2_U2394 );
nand NAND2_10275 ( P2_U6199 , P2_UWORD_REG_9_ , P2_U3538 );
nand NAND2_10276 ( P2_U6200 , P2_EAX_REG_24_ , P2_U2395 );
nand NAND2_10277 ( P2_U6201 , U284 , P2_U2394 );
nand NAND2_10278 ( P2_U6202 , P2_UWORD_REG_8_ , P2_U3538 );
nand NAND2_10279 ( P2_U6203 , P2_EAX_REG_23_ , P2_U2395 );
nand NAND2_10280 ( P2_U6204 , P2_U2394 , U285 );
nand NAND2_10281 ( P2_U6205 , P2_UWORD_REG_7_ , P2_U3538 );
nand NAND2_10282 ( P2_U6206 , P2_EAX_REG_22_ , P2_U2395 );
nand NAND2_10283 ( P2_U6207 , P2_U2394 , U286 );
nand NAND2_10284 ( P2_U6208 , P2_UWORD_REG_6_ , P2_U3538 );
nand NAND2_10285 ( P2_U6209 , P2_EAX_REG_21_ , P2_U2395 );
nand NAND2_10286 ( P2_U6210 , P2_U2394 , U287 );
nand NAND2_10287 ( P2_U6211 , P2_UWORD_REG_5_ , P2_U3538 );
nand NAND2_10288 ( P2_U6212 , P2_EAX_REG_20_ , P2_U2395 );
nand NAND2_10289 ( P2_U6213 , P2_U2394 , U288 );
nand NAND2_10290 ( P2_U6214 , P2_UWORD_REG_4_ , P2_U3538 );
nand NAND2_10291 ( P2_U6215 , P2_EAX_REG_19_ , P2_U2395 );
nand NAND2_10292 ( P2_U6216 , P2_U2394 , U289 );
nand NAND2_10293 ( P2_U6217 , P2_UWORD_REG_3_ , P2_U3538 );
nand NAND2_10294 ( P2_U6218 , P2_EAX_REG_18_ , P2_U2395 );
nand NAND2_10295 ( P2_U6219 , P2_U2394 , U292 );
nand NAND2_10296 ( P2_U6220 , P2_UWORD_REG_2_ , P2_U3538 );
nand NAND2_10297 ( P2_U6221 , P2_EAX_REG_17_ , P2_U2395 );
nand NAND2_10298 ( P2_U6222 , P2_U2394 , U303 );
nand NAND2_10299 ( P2_U6223 , P2_UWORD_REG_1_ , P2_U3538 );
nand NAND2_10300 ( P2_U6224 , P2_EAX_REG_16_ , P2_U2395 );
nand NAND2_10301 ( P2_U6225 , P2_U2394 , U314 );
nand NAND2_10302 ( P2_U6226 , P2_UWORD_REG_0_ , P2_U3538 );
nand NAND3_10303 ( P2_U6227 , P2_U4057 , P2_U4421 , P2_R2167_U6 );
nand NAND2_10304 ( P2_U6228 , P2_U4058 , P2_U2446 );
nand NAND2_10305 ( P2_U6229 , P2_U6228 , P2_U6227 );
nand NAND2_10306 ( P2_U6230 , P2_U4411 , P2_U6229 );
nand NAND2_10307 ( P2_U6231 , P2_U4467 , P2_STATE2_REG_1_ );
not NOT1_10308 ( P2_U6232 , P2_U3541 );
nand NAND2_10309 ( P2_U6233 , P2_U2430 , P2_EAX_REG_0_ );
nand NAND2_10310 ( P2_U6234 , P2_U2396 , P2_LWORD_REG_0_ );
nand NAND2_10311 ( P2_U6235 , P2_DATAO_REG_0_ , P2_U6232 );
nand NAND2_10312 ( P2_U6236 , P2_U2430 , P2_EAX_REG_1_ );
nand NAND2_10313 ( P2_U6237 , P2_U2396 , P2_LWORD_REG_1_ );
nand NAND2_10314 ( P2_U6238 , P2_DATAO_REG_1_ , P2_U6232 );
nand NAND2_10315 ( P2_U6239 , P2_U2430 , P2_EAX_REG_2_ );
nand NAND2_10316 ( P2_U6240 , P2_U2396 , P2_LWORD_REG_2_ );
nand NAND2_10317 ( P2_U6241 , P2_DATAO_REG_2_ , P2_U6232 );
nand NAND2_10318 ( P2_U6242 , P2_U2430 , P2_EAX_REG_3_ );
nand NAND2_10319 ( P2_U6243 , P2_U2396 , P2_LWORD_REG_3_ );
nand NAND2_10320 ( P2_U6244 , P2_DATAO_REG_3_ , P2_U6232 );
nand NAND2_10321 ( P2_U6245 , P2_U2430 , P2_EAX_REG_4_ );
nand NAND2_10322 ( P2_U6246 , P2_U2396 , P2_LWORD_REG_4_ );
nand NAND2_10323 ( P2_U6247 , P2_DATAO_REG_4_ , P2_U6232 );
nand NAND2_10324 ( P2_U6248 , P2_U2430 , P2_EAX_REG_5_ );
nand NAND2_10325 ( P2_U6249 , P2_U2396 , P2_LWORD_REG_5_ );
nand NAND2_10326 ( P2_U6250 , P2_DATAO_REG_5_ , P2_U6232 );
nand NAND2_10327 ( P2_U6251 , P2_U2430 , P2_EAX_REG_6_ );
nand NAND2_10328 ( P2_U6252 , P2_U2396 , P2_LWORD_REG_6_ );
nand NAND2_10329 ( P2_U6253 , P2_DATAO_REG_6_ , P2_U6232 );
nand NAND2_10330 ( P2_U6254 , P2_U2430 , P2_EAX_REG_7_ );
nand NAND2_10331 ( P2_U6255 , P2_U2396 , P2_LWORD_REG_7_ );
nand NAND2_10332 ( P2_U6256 , P2_DATAO_REG_7_ , P2_U6232 );
nand NAND2_10333 ( P2_U6257 , P2_U2430 , P2_EAX_REG_8_ );
nand NAND2_10334 ( P2_U6258 , P2_U2396 , P2_LWORD_REG_8_ );
nand NAND2_10335 ( P2_U6259 , P2_DATAO_REG_8_ , P2_U6232 );
nand NAND2_10336 ( P2_U6260 , P2_U2430 , P2_EAX_REG_9_ );
nand NAND2_10337 ( P2_U6261 , P2_U2396 , P2_LWORD_REG_9_ );
nand NAND2_10338 ( P2_U6262 , P2_DATAO_REG_9_ , P2_U6232 );
nand NAND2_10339 ( P2_U6263 , P2_U2430 , P2_EAX_REG_10_ );
nand NAND2_10340 ( P2_U6264 , P2_U2396 , P2_LWORD_REG_10_ );
nand NAND2_10341 ( P2_U6265 , P2_DATAO_REG_10_ , P2_U6232 );
nand NAND2_10342 ( P2_U6266 , P2_U2430 , P2_EAX_REG_11_ );
nand NAND2_10343 ( P2_U6267 , P2_U2396 , P2_LWORD_REG_11_ );
nand NAND2_10344 ( P2_U6268 , P2_DATAO_REG_11_ , P2_U6232 );
nand NAND2_10345 ( P2_U6269 , P2_U2430 , P2_EAX_REG_12_ );
nand NAND2_10346 ( P2_U6270 , P2_U2396 , P2_LWORD_REG_12_ );
nand NAND2_10347 ( P2_U6271 , P2_DATAO_REG_12_ , P2_U6232 );
nand NAND2_10348 ( P2_U6272 , P2_U2430 , P2_EAX_REG_13_ );
nand NAND2_10349 ( P2_U6273 , P2_U2396 , P2_LWORD_REG_13_ );
nand NAND2_10350 ( P2_U6274 , P2_DATAO_REG_13_ , P2_U6232 );
nand NAND2_10351 ( P2_U6275 , P2_U2430 , P2_EAX_REG_14_ );
nand NAND2_10352 ( P2_U6276 , P2_U2396 , P2_LWORD_REG_14_ );
nand NAND2_10353 ( P2_U6277 , P2_DATAO_REG_14_ , P2_U6232 );
nand NAND2_10354 ( P2_U6278 , P2_U2430 , P2_EAX_REG_15_ );
nand NAND2_10355 ( P2_U6279 , P2_U2396 , P2_LWORD_REG_15_ );
nand NAND2_10356 ( P2_U6280 , P2_DATAO_REG_15_ , P2_U6232 );
nand NAND2_10357 ( P2_U6281 , P2_U2435 , P2_EAX_REG_16_ );
nand NAND2_10358 ( P2_U6282 , P2_U2396 , P2_UWORD_REG_0_ );
nand NAND2_10359 ( P2_U6283 , P2_DATAO_REG_16_ , P2_U6232 );
nand NAND2_10360 ( P2_U6284 , P2_U2435 , P2_EAX_REG_17_ );
nand NAND2_10361 ( P2_U6285 , P2_U2396 , P2_UWORD_REG_1_ );
nand NAND2_10362 ( P2_U6286 , P2_DATAO_REG_17_ , P2_U6232 );
nand NAND2_10363 ( P2_U6287 , P2_U2435 , P2_EAX_REG_18_ );
nand NAND2_10364 ( P2_U6288 , P2_U2396 , P2_UWORD_REG_2_ );
nand NAND2_10365 ( P2_U6289 , P2_DATAO_REG_18_ , P2_U6232 );
nand NAND2_10366 ( P2_U6290 , P2_U2435 , P2_EAX_REG_19_ );
nand NAND2_10367 ( P2_U6291 , P2_U2396 , P2_UWORD_REG_3_ );
nand NAND2_10368 ( P2_U6292 , P2_DATAO_REG_19_ , P2_U6232 );
nand NAND2_10369 ( P2_U6293 , P2_U2435 , P2_EAX_REG_20_ );
nand NAND2_10370 ( P2_U6294 , P2_U2396 , P2_UWORD_REG_4_ );
nand NAND2_10371 ( P2_U6295 , P2_DATAO_REG_20_ , P2_U6232 );
nand NAND2_10372 ( P2_U6296 , P2_U2435 , P2_EAX_REG_21_ );
nand NAND2_10373 ( P2_U6297 , P2_U2396 , P2_UWORD_REG_5_ );
nand NAND2_10374 ( P2_U6298 , P2_DATAO_REG_21_ , P2_U6232 );
nand NAND2_10375 ( P2_U6299 , P2_U2435 , P2_EAX_REG_22_ );
nand NAND2_10376 ( P2_U6300 , P2_U2396 , P2_UWORD_REG_6_ );
nand NAND2_10377 ( P2_U6301 , P2_DATAO_REG_22_ , P2_U6232 );
nand NAND2_10378 ( P2_U6302 , P2_U2435 , P2_EAX_REG_23_ );
nand NAND2_10379 ( P2_U6303 , P2_U2396 , P2_UWORD_REG_7_ );
nand NAND2_10380 ( P2_U6304 , P2_DATAO_REG_23_ , P2_U6232 );
nand NAND2_10381 ( P2_U6305 , P2_U2435 , P2_EAX_REG_24_ );
nand NAND2_10382 ( P2_U6306 , P2_U2396 , P2_UWORD_REG_8_ );
nand NAND2_10383 ( P2_U6307 , P2_DATAO_REG_24_ , P2_U6232 );
nand NAND2_10384 ( P2_U6308 , P2_U2435 , P2_EAX_REG_25_ );
nand NAND2_10385 ( P2_U6309 , P2_U2396 , P2_UWORD_REG_9_ );
nand NAND2_10386 ( P2_U6310 , P2_DATAO_REG_25_ , P2_U6232 );
nand NAND2_10387 ( P2_U6311 , P2_U2435 , P2_EAX_REG_26_ );
nand NAND2_10388 ( P2_U6312 , P2_U2396 , P2_UWORD_REG_10_ );
nand NAND2_10389 ( P2_U6313 , P2_DATAO_REG_26_ , P2_U6232 );
nand NAND2_10390 ( P2_U6314 , P2_U2435 , P2_EAX_REG_27_ );
nand NAND2_10391 ( P2_U6315 , P2_U2396 , P2_UWORD_REG_11_ );
nand NAND2_10392 ( P2_U6316 , P2_DATAO_REG_27_ , P2_U6232 );
nand NAND2_10393 ( P2_U6317 , P2_U2435 , P2_EAX_REG_28_ );
nand NAND2_10394 ( P2_U6318 , P2_U2396 , P2_UWORD_REG_12_ );
nand NAND2_10395 ( P2_U6319 , P2_DATAO_REG_28_ , P2_U6232 );
nand NAND2_10396 ( P2_U6320 , P2_U2435 , P2_EAX_REG_29_ );
nand NAND2_10397 ( P2_U6321 , P2_U2396 , P2_UWORD_REG_13_ );
nand NAND2_10398 ( P2_U6322 , P2_DATAO_REG_29_ , P2_U6232 );
nand NAND2_10399 ( P2_U6323 , P2_U2435 , P2_EAX_REG_30_ );
nand NAND2_10400 ( P2_U6324 , P2_U2396 , P2_UWORD_REG_14_ );
nand NAND2_10401 ( P2_U6325 , P2_DATAO_REG_30_ , P2_U6232 );
nand NAND2_10402 ( P2_U6326 , P2_U2513 , P2_U3254 );
nand NAND2_10403 ( P2_U6327 , P2_U2433 , U314 );
nand NAND2_10404 ( P2_U6328 , P2_ADD_391_1196_U87 , P2_U2397 );
nand NAND2_10405 ( P2_U6329 , P2_U2380 , P2_R2096_U68 );
nand NAND2_10406 ( P2_U6330 , P2_EAX_REG_0_ , P2_U3542 );
nand NAND2_10407 ( P2_U6331 , P2_U2433 , U303 );
nand NAND2_10408 ( P2_U6332 , P2_ADD_391_1196_U12 , P2_U2397 );
nand NAND2_10409 ( P2_U6333 , P2_U2380 , P2_R2096_U51 );
nand NAND2_10410 ( P2_U6334 , P2_EAX_REG_1_ , P2_U3542 );
nand NAND2_10411 ( P2_U6335 , P2_U2433 , U292 );
nand NAND2_10412 ( P2_U6336 , P2_ADD_391_1196_U92 , P2_U2397 );
nand NAND2_10413 ( P2_U6337 , P2_U2380 , P2_R2096_U77 );
nand NAND2_10414 ( P2_U6338 , P2_EAX_REG_2_ , P2_U3542 );
nand NAND2_10415 ( P2_U6339 , P2_U2433 , U289 );
nand NAND2_10416 ( P2_U6340 , P2_ADD_391_1196_U91 , P2_U2397 );
nand NAND2_10417 ( P2_U6341 , P2_U2380 , P2_R2096_U75 );
nand NAND2_10418 ( P2_U6342 , P2_EAX_REG_3_ , P2_U3542 );
nand NAND2_10419 ( P2_U6343 , P2_U2433 , U288 );
nand NAND2_10420 ( P2_U6344 , P2_ADD_391_1196_U90 , P2_U2397 );
nand NAND2_10421 ( P2_U6345 , P2_U2380 , P2_R2096_U74 );
nand NAND2_10422 ( P2_U6346 , P2_EAX_REG_4_ , P2_U3542 );
nand NAND2_10423 ( P2_U6347 , P2_U2433 , U287 );
nand NAND2_10424 ( P2_U6348 , P2_ADD_391_1196_U9 , P2_U2397 );
nand NAND2_10425 ( P2_U6349 , P2_U2380 , P2_R2096_U73 );
nand NAND2_10426 ( P2_U6350 , P2_EAX_REG_5_ , P2_U3542 );
nand NAND2_10427 ( P2_U6351 , P2_U2433 , U286 );
nand NAND2_10428 ( P2_U6352 , P2_ADD_391_1196_U89 , P2_U2397 );
nand NAND2_10429 ( P2_U6353 , P2_U2380 , P2_R2096_U72 );
nand NAND2_10430 ( P2_U6354 , P2_EAX_REG_6_ , P2_U3542 );
nand NAND2_10431 ( P2_U6355 , P2_U2433 , U285 );
nand NAND2_10432 ( P2_U6356 , P2_ADD_391_1196_U10 , P2_U2397 );
nand NAND2_10433 ( P2_U6357 , P2_U2380 , P2_R2096_U71 );
nand NAND2_10434 ( P2_U6358 , P2_EAX_REG_7_ , P2_U3542 );
nand NAND2_10435 ( P2_U6359 , P2_U2433 , U284 );
nand NAND2_10436 ( P2_U6360 , P2_ADD_391_1196_U88 , P2_U2397 );
nand NAND2_10437 ( P2_U6361 , P2_U2380 , P2_R2096_U70 );
nand NAND2_10438 ( P2_U6362 , P2_EAX_REG_8_ , P2_U3542 );
nand NAND2_10439 ( P2_U6363 , P2_U2433 , U283 );
nand NAND2_10440 ( P2_U6364 , P2_ADD_391_1196_U11 , P2_U2397 );
nand NAND2_10441 ( P2_U6365 , P2_U2380 , P2_R2096_U69 );
nand NAND2_10442 ( P2_U6366 , P2_EAX_REG_9_ , P2_U3542 );
nand NAND2_10443 ( P2_U6367 , P2_U2433 , U313 );
nand NAND2_10444 ( P2_U6368 , P2_ADD_391_1196_U109 , P2_U2397 );
nand NAND2_10445 ( P2_U6369 , P2_U2380 , P2_R2096_U97 );
nand NAND2_10446 ( P2_U6370 , P2_EAX_REG_10_ , P2_U3542 );
nand NAND2_10447 ( P2_U6371 , P2_U2433 , U312 );
nand NAND2_10448 ( P2_U6372 , P2_ADD_391_1196_U5 , P2_U2397 );
nand NAND2_10449 ( P2_U6373 , P2_U2380 , P2_R2096_U96 );
nand NAND2_10450 ( P2_U6374 , P2_EAX_REG_11_ , P2_U3542 );
nand NAND2_10451 ( P2_U6375 , P2_U2433 , U311 );
nand NAND2_10452 ( P2_U6376 , P2_ADD_391_1196_U108 , P2_U2397 );
nand NAND2_10453 ( P2_U6377 , P2_U2380 , P2_R2096_U95 );
nand NAND2_10454 ( P2_U6378 , P2_EAX_REG_12_ , P2_U3542 );
nand NAND2_10455 ( P2_U6379 , P2_U2433 , U310 );
nand NAND2_10456 ( P2_U6380 , P2_ADD_391_1196_U6 , P2_U2397 );
nand NAND2_10457 ( P2_U6381 , P2_U2380 , P2_R2096_U94 );
nand NAND2_10458 ( P2_U6382 , P2_EAX_REG_13_ , P2_U3542 );
nand NAND2_10459 ( P2_U6383 , P2_U2433 , U309 );
nand NAND2_10460 ( P2_U6384 , P2_ADD_391_1196_U107 , P2_U2397 );
nand NAND2_10461 ( P2_U6385 , P2_U2380 , P2_R2096_U93 );
nand NAND2_10462 ( P2_U6386 , P2_EAX_REG_14_ , P2_U3542 );
nand NAND2_10463 ( P2_U6387 , P2_U2433 , U308 );
nand NAND2_10464 ( P2_U6388 , P2_ADD_391_1196_U7 , P2_U2397 );
nand NAND2_10465 ( P2_U6389 , P2_U2380 , P2_R2096_U92 );
nand NAND2_10466 ( P2_U6390 , P2_EAX_REG_15_ , P2_U3542 );
nand NAND2_10467 ( P2_U6391 , P2_U2434 , U314 );
nand NAND2_10468 ( P2_U6392 , P2_U2427 , U307 );
nand NAND2_10469 ( P2_U6393 , P2_ADD_391_1196_U106 , P2_U2397 );
nand NAND2_10470 ( P2_U6394 , P2_U2380 , P2_R2096_U91 );
nand NAND2_10471 ( P2_U6395 , P2_EAX_REG_16_ , P2_U3542 );
nand NAND2_10472 ( P2_U6396 , P2_U2434 , U303 );
nand NAND2_10473 ( P2_U6397 , P2_U2427 , U306 );
nand NAND2_10474 ( P2_U6398 , P2_ADD_391_1196_U105 , P2_U2397 );
nand NAND2_10475 ( P2_U6399 , P2_U2380 , P2_R2096_U90 );
nand NAND2_10476 ( P2_U6400 , P2_EAX_REG_17_ , P2_U3542 );
nand NAND2_10477 ( P2_U6401 , P2_U2434 , U292 );
nand NAND2_10478 ( P2_U6402 , P2_U2427 , U305 );
nand NAND2_10479 ( P2_U6403 , P2_ADD_391_1196_U104 , P2_U2397 );
nand NAND2_10480 ( P2_U6404 , P2_U2380 , P2_R2096_U89 );
nand NAND2_10481 ( P2_U6405 , P2_EAX_REG_18_ , P2_U3542 );
nand NAND2_10482 ( P2_U6406 , P2_U2434 , U289 );
nand NAND2_10483 ( P2_U6407 , P2_U2427 , U304 );
nand NAND2_10484 ( P2_U6408 , P2_ADD_391_1196_U103 , P2_U2397 );
nand NAND2_10485 ( P2_U6409 , P2_U2380 , P2_R2096_U88 );
nand NAND2_10486 ( P2_U6410 , P2_EAX_REG_19_ , P2_U3542 );
nand NAND2_10487 ( P2_U6411 , P2_U2434 , U288 );
nand NAND2_10488 ( P2_U6412 , P2_U2427 , U302 );
nand NAND2_10489 ( P2_U6413 , P2_ADD_391_1196_U102 , P2_U2397 );
nand NAND2_10490 ( P2_U6414 , P2_U2380 , P2_R2096_U87 );
nand NAND2_10491 ( P2_U6415 , P2_EAX_REG_20_ , P2_U3542 );
nand NAND2_10492 ( P2_U6416 , P2_U2434 , U287 );
nand NAND2_10493 ( P2_U6417 , P2_U2427 , U301 );
nand NAND2_10494 ( P2_U6418 , P2_ADD_391_1196_U101 , P2_U2397 );
nand NAND2_10495 ( P2_U6419 , P2_U2380 , P2_R2096_U86 );
nand NAND2_10496 ( P2_U6420 , P2_EAX_REG_21_ , P2_U3542 );
nand NAND2_10497 ( P2_U6421 , P2_U2434 , U286 );
nand NAND2_10498 ( P2_U6422 , P2_U2427 , U300 );
nand NAND2_10499 ( P2_U6423 , P2_ADD_391_1196_U100 , P2_U2397 );
nand NAND2_10500 ( P2_U6424 , P2_U2380 , P2_R2096_U85 );
nand NAND2_10501 ( P2_U6425 , P2_EAX_REG_22_ , P2_U3542 );
nand NAND2_10502 ( P2_U6426 , P2_U2434 , U285 );
nand NAND2_10503 ( P2_U6427 , P2_U2427 , U299 );
nand NAND2_10504 ( P2_U6428 , P2_ADD_391_1196_U99 , P2_U2397 );
nand NAND2_10505 ( P2_U6429 , P2_U2380 , P2_R2096_U84 );
nand NAND2_10506 ( P2_U6430 , P2_EAX_REG_23_ , P2_U3542 );
nand NAND2_10507 ( P2_U6431 , P2_U2434 , U284 );
nand NAND2_10508 ( P2_U6432 , P2_U2427 , U298 );
nand NAND2_10509 ( P2_U6433 , P2_ADD_391_1196_U98 , P2_U2397 );
nand NAND2_10510 ( P2_U6434 , P2_U2380 , P2_R2096_U83 );
nand NAND2_10511 ( P2_U6435 , P2_EAX_REG_24_ , P2_U3542 );
nand NAND2_10512 ( P2_U6436 , P2_U2434 , U283 );
nand NAND2_10513 ( P2_U6437 , P2_U2427 , U297 );
nand NAND2_10514 ( P2_U6438 , P2_ADD_391_1196_U97 , P2_U2397 );
nand NAND2_10515 ( P2_U6439 , P2_U2380 , P2_R2096_U82 );
nand NAND2_10516 ( P2_U6440 , P2_EAX_REG_25_ , P2_U3542 );
nand NAND2_10517 ( P2_U6441 , P2_U2434 , U313 );
nand NAND2_10518 ( P2_U6442 , P2_U2427 , U296 );
nand NAND2_10519 ( P2_U6443 , P2_ADD_391_1196_U96 , P2_U2397 );
nand NAND2_10520 ( P2_U6444 , P2_U2380 , P2_R2096_U81 );
nand NAND2_10521 ( P2_U6445 , P2_EAX_REG_26_ , P2_U3542 );
nand NAND2_10522 ( P2_U6446 , P2_U2434 , U312 );
nand NAND2_10523 ( P2_U6447 , P2_U2427 , U295 );
nand NAND2_10524 ( P2_U6448 , P2_ADD_391_1196_U95 , P2_U2397 );
nand NAND2_10525 ( P2_U6449 , P2_U2380 , P2_R2096_U80 );
nand NAND2_10526 ( P2_U6450 , P2_EAX_REG_27_ , P2_U3542 );
nand NAND2_10527 ( P2_U6451 , P2_U2434 , U311 );
nand NAND2_10528 ( P2_U6452 , P2_U2427 , U294 );
nand NAND2_10529 ( P2_U6453 , P2_ADD_391_1196_U94 , P2_U2397 );
nand NAND2_10530 ( P2_U6454 , P2_U2380 , P2_R2096_U79 );
nand NAND2_10531 ( P2_U6455 , P2_EAX_REG_28_ , P2_U3542 );
nand NAND2_10532 ( P2_U6456 , P2_U2434 , U310 );
nand NAND2_10533 ( P2_U6457 , P2_U2427 , U293 );
nand NAND2_10534 ( P2_U6458 , P2_ADD_391_1196_U93 , P2_U2397 );
nand NAND2_10535 ( P2_U6459 , P2_U2380 , P2_R2096_U78 );
nand NAND2_10536 ( P2_U6460 , P2_EAX_REG_29_ , P2_U3542 );
nand NAND2_10537 ( P2_U6461 , P2_U2434 , U309 );
nand NAND2_10538 ( P2_U6462 , P2_U2427 , U291 );
nand NAND2_10539 ( P2_U6463 , P2_ADD_391_1196_U8 , P2_U2397 );
nand NAND2_10540 ( P2_U6464 , P2_U2380 , P2_R2096_U76 );
nand NAND2_10541 ( P2_U6465 , P2_EAX_REG_30_ , P2_U3542 );
nand NAND2_10542 ( P2_U6466 , P2_U2427 , U290 );
nand NAND2_10543 ( P2_U6467 , P2_U2380 , P2_R2096_U50 );
nand NAND2_10544 ( P2_U6468 , P2_EAX_REG_31_ , P2_U3542 );
nand NAND2_10545 ( P2_U6469 , P2_U4435 , P2_U3297 );
nand NAND2_10546 ( P2_U6470 , P2_U3578 , P2_U6469 );
nand NAND2_10547 ( P2_U6471 , P2_U2393 , P2_R2182_U69 );
nand NAND2_10548 ( P2_U6472 , P2_U2379 , P2_R2099_U94 );
nand NAND2_10549 ( P2_U6473 , P2_EBX_REG_0_ , P2_U3543 );
nand NAND2_10550 ( P2_U6474 , P2_U2393 , P2_R2182_U68 );
nand NAND2_10551 ( P2_U6475 , P2_U2379 , P2_R2099_U5 );
nand NAND2_10552 ( P2_U6476 , P2_EBX_REG_1_ , P2_U3543 );
nand NAND2_10553 ( P2_U6477 , P2_U2393 , P2_R2182_U40 );
nand NAND2_10554 ( P2_U6478 , P2_U2379 , P2_R2099_U96 );
nand NAND2_10555 ( P2_U6479 , P2_EBX_REG_2_ , P2_U3543 );
nand NAND2_10556 ( P2_U6480 , P2_U2393 , P2_R2182_U76 );
nand NAND2_10557 ( P2_U6481 , P2_U2379 , P2_R2099_U95 );
nand NAND2_10558 ( P2_U6482 , P2_EBX_REG_3_ , P2_U3543 );
nand NAND2_10559 ( P2_U6483 , P2_R2182_U75 , P2_U2393 );
nand NAND2_10560 ( P2_U6484 , P2_U2379 , P2_R2099_U98 );
nand NAND2_10561 ( P2_U6485 , P2_EBX_REG_4_ , P2_U3543 );
nand NAND2_10562 ( P2_U6486 , P2_R2182_U74 , P2_U2393 );
nand NAND2_10563 ( P2_U6487 , P2_U2379 , P2_R2099_U71 );
nand NAND2_10564 ( P2_U6488 , P2_EBX_REG_5_ , P2_U3543 );
nand NAND2_10565 ( P2_U6489 , P2_R2182_U73 , P2_U2393 );
nand NAND2_10566 ( P2_U6490 , P2_U2379 , P2_R2099_U70 );
nand NAND2_10567 ( P2_U6491 , P2_EBX_REG_6_ , P2_U3543 );
nand NAND2_10568 ( P2_U6492 , P2_R2182_U72 , P2_U2393 );
nand NAND2_10569 ( P2_U6493 , P2_U2379 , P2_R2099_U69 );
nand NAND2_10570 ( P2_U6494 , P2_EBX_REG_7_ , P2_U3543 );
nand NAND2_10571 ( P2_U6495 , P2_R2182_U71 , P2_U2393 );
nand NAND2_10572 ( P2_U6496 , P2_U2379 , P2_R2099_U68 );
nand NAND2_10573 ( P2_U6497 , P2_EBX_REG_8_ , P2_U3543 );
nand NAND2_10574 ( P2_U6498 , P2_R2182_U70 , P2_U2393 );
nand NAND2_10575 ( P2_U6499 , P2_U2379 , P2_R2099_U67 );
nand NAND2_10576 ( P2_U6500 , P2_EBX_REG_9_ , P2_U3543 );
nand NAND2_10577 ( P2_U6501 , P2_R2182_U96 , P2_U2393 );
nand NAND2_10578 ( P2_U6502 , P2_U2379 , P2_R2099_U93 );
nand NAND2_10579 ( P2_U6503 , P2_EBX_REG_10_ , P2_U3543 );
nand NAND2_10580 ( P2_U6504 , P2_R2182_U95 , P2_U2393 );
nand NAND2_10581 ( P2_U6505 , P2_U2379 , P2_R2099_U92 );
nand NAND2_10582 ( P2_U6506 , P2_EBX_REG_11_ , P2_U3543 );
nand NAND2_10583 ( P2_U6507 , P2_R2182_U94 , P2_U2393 );
nand NAND2_10584 ( P2_U6508 , P2_U2379 , P2_R2099_U91 );
nand NAND2_10585 ( P2_U6509 , P2_EBX_REG_12_ , P2_U3543 );
nand NAND2_10586 ( P2_U6510 , P2_R2182_U93 , P2_U2393 );
nand NAND2_10587 ( P2_U6511 , P2_U2379 , P2_R2099_U90 );
nand NAND2_10588 ( P2_U6512 , P2_EBX_REG_13_ , P2_U3543 );
nand NAND2_10589 ( P2_U6513 , P2_R2182_U92 , P2_U2393 );
nand NAND2_10590 ( P2_U6514 , P2_U2379 , P2_R2099_U89 );
nand NAND2_10591 ( P2_U6515 , P2_EBX_REG_14_ , P2_U3543 );
nand NAND2_10592 ( P2_U6516 , P2_R2182_U91 , P2_U2393 );
nand NAND2_10593 ( P2_U6517 , P2_U2379 , P2_R2099_U88 );
nand NAND2_10594 ( P2_U6518 , P2_EBX_REG_15_ , P2_U3543 );
nand NAND2_10595 ( P2_U6519 , P2_R2182_U90 , P2_U2393 );
nand NAND2_10596 ( P2_U6520 , P2_U2379 , P2_R2099_U87 );
nand NAND2_10597 ( P2_U6521 , P2_EBX_REG_16_ , P2_U3543 );
nand NAND2_10598 ( P2_U6522 , P2_R2182_U89 , P2_U2393 );
nand NAND2_10599 ( P2_U6523 , P2_U2379 , P2_R2099_U86 );
nand NAND2_10600 ( P2_U6524 , P2_EBX_REG_17_ , P2_U3543 );
nand NAND2_10601 ( P2_U6525 , P2_R2182_U88 , P2_U2393 );
nand NAND2_10602 ( P2_U6526 , P2_U2379 , P2_R2099_U85 );
nand NAND2_10603 ( P2_U6527 , P2_EBX_REG_18_ , P2_U3543 );
nand NAND2_10604 ( P2_U6528 , P2_R2182_U87 , P2_U2393 );
nand NAND2_10605 ( P2_U6529 , P2_U2379 , P2_R2099_U84 );
nand NAND2_10606 ( P2_U6530 , P2_EBX_REG_19_ , P2_U3543 );
nand NAND2_10607 ( P2_U6531 , P2_R2182_U86 , P2_U2393 );
nand NAND2_10608 ( P2_U6532 , P2_U2379 , P2_R2099_U83 );
nand NAND2_10609 ( P2_U6533 , P2_EBX_REG_20_ , P2_U3543 );
nand NAND2_10610 ( P2_U6534 , P2_R2182_U85 , P2_U2393 );
nand NAND2_10611 ( P2_U6535 , P2_U2379 , P2_R2099_U82 );
nand NAND2_10612 ( P2_U6536 , P2_EBX_REG_21_ , P2_U3543 );
nand NAND2_10613 ( P2_U6537 , P2_R2182_U84 , P2_U2393 );
nand NAND2_10614 ( P2_U6538 , P2_U2379 , P2_R2099_U81 );
nand NAND2_10615 ( P2_U6539 , P2_EBX_REG_22_ , P2_U3543 );
nand NAND2_10616 ( P2_U6540 , P2_R2182_U83 , P2_U2393 );
nand NAND2_10617 ( P2_U6541 , P2_U2379 , P2_R2099_U80 );
nand NAND2_10618 ( P2_U6542 , P2_EBX_REG_23_ , P2_U3543 );
nand NAND2_10619 ( P2_U6543 , P2_R2182_U82 , P2_U2393 );
nand NAND2_10620 ( P2_U6544 , P2_U2379 , P2_R2099_U79 );
nand NAND2_10621 ( P2_U6545 , P2_EBX_REG_24_ , P2_U3543 );
nand NAND2_10622 ( P2_U6546 , P2_R2182_U81 , P2_U2393 );
nand NAND2_10623 ( P2_U6547 , P2_U2379 , P2_R2099_U78 );
nand NAND2_10624 ( P2_U6548 , P2_EBX_REG_25_ , P2_U3543 );
nand NAND2_10625 ( P2_U6549 , P2_R2182_U80 , P2_U2393 );
nand NAND2_10626 ( P2_U6550 , P2_U2379 , P2_R2099_U77 );
nand NAND2_10627 ( P2_U6551 , P2_EBX_REG_26_ , P2_U3543 );
nand NAND2_10628 ( P2_U6552 , P2_R2182_U79 , P2_U2393 );
nand NAND2_10629 ( P2_U6553 , P2_U2379 , P2_R2099_U76 );
nand NAND2_10630 ( P2_U6554 , P2_EBX_REG_27_ , P2_U3543 );
nand NAND2_10631 ( P2_U6555 , P2_R2182_U78 , P2_U2393 );
nand NAND2_10632 ( P2_U6556 , P2_U2379 , P2_R2099_U75 );
nand NAND2_10633 ( P2_U6557 , P2_EBX_REG_28_ , P2_U3543 );
nand NAND2_10634 ( P2_U6558 , P2_R2182_U77 , P2_U2393 );
nand NAND2_10635 ( P2_U6559 , P2_U2379 , P2_R2099_U74 );
nand NAND2_10636 ( P2_U6560 , P2_EBX_REG_29_ , P2_U3543 );
nand NAND2_10637 ( P2_U6561 , P2_R2182_U41 , P2_U2393 );
nand NAND2_10638 ( P2_U6562 , P2_U2379 , P2_R2099_U73 );
nand NAND2_10639 ( P2_U6563 , P2_EBX_REG_30_ , P2_U3543 );
nand NAND2_10640 ( P2_U6564 , P2_U2379 , P2_R2099_U72 );
nand NAND2_10641 ( P2_U6565 , P2_EBX_REG_31_ , P2_U3543 );
nand NAND2_10642 ( P2_U6566 , P2_R2088_U6 , P2_U4603 );
nand NAND2_10643 ( P2_U6567 , P2_U4433 , P2_R2167_U6 );
nand NAND2_10644 ( P2_U6568 , P2_U6567 , P2_U6566 );
nand NAND2_10645 ( P2_U6569 , P2_U4461 , P2_U3284 );
not NOT1_10646 ( P2_U6570 , P2_U3546 );
not NOT1_10647 ( P2_U6571 , P2_U3545 );
or OR2_10648 ( P2_U6572 , P2_STATEBS16_REG , U211 );
nand NAND2_10649 ( P2_U6573 , P2_R2267_U21 , P2_U2587 );
nand NAND2_10650 ( P2_U6574 , P2_U2588 , P2_R2096_U68 );
nand NAND2_10651 ( P2_U6575 , P2_EBX_REG_0_ , P2_U7743 );
nand NAND2_10652 ( P2_U6576 , P2_U2437 , P2_R2182_U69 );
nand NAND2_10653 ( P2_U6577 , P2_U2392 , P2_R2099_U94 );
nand NAND2_10654 ( P2_U6578 , P2_U2383 , P2_PHYADDRPOINTER_REG_0_ );
nand NAND2_10655 ( P2_U6579 , P2_U2382 , P2_U3683 );
nand NAND2_10656 ( P2_U6580 , P2_U2378 , P2_PHYADDRPOINTER_REG_0_ );
nand NAND2_10657 ( P2_U6581 , P2_U6570 , P2_REIP_REG_0_ );
nand NAND2_10658 ( P2_U6582 , P2_R2267_U43 , P2_U2587 );
nand NAND2_10659 ( P2_U6583 , P2_U2588 , P2_R2096_U51 );
nand NAND2_10660 ( P2_U6584 , P2_EBX_REG_1_ , P2_U7743 );
nand NAND2_10661 ( P2_U6585 , P2_U2437 , P2_R2182_U68 );
nand NAND2_10662 ( P2_U6586 , P2_U2392 , P2_R2099_U5 );
nand NAND2_10663 ( P2_U6587 , P2_U2383 , P2_R2337_U4 );
nand NAND2_10664 ( P2_U6588 , P2_U2382 , P2_R1957_U49 );
nand NAND2_10665 ( P2_U6589 , P2_U2378 , P2_PHYADDRPOINTER_REG_1_ );
nand NAND2_10666 ( P2_U6590 , P2_U6570 , P2_REIP_REG_1_ );
nand NAND2_10667 ( P2_U6591 , P2_R2267_U65 , P2_U2587 );
nand NAND2_10668 ( P2_U6592 , P2_U2588 , P2_R2096_U77 );
nand NAND2_10669 ( P2_U6593 , P2_EBX_REG_2_ , P2_U7743 );
nand NAND2_10670 ( P2_U6594 , P2_U2437 , P2_R2182_U40 );
nand NAND2_10671 ( P2_U6595 , P2_U2392 , P2_R2099_U96 );
nand NAND2_10672 ( P2_U6596 , P2_U2383 , P2_R2337_U70 );
nand NAND2_10673 ( P2_U6597 , P2_R1957_U17 , P2_U2382 );
nand NAND2_10674 ( P2_U6598 , P2_U2378 , P2_PHYADDRPOINTER_REG_2_ );
nand NAND2_10675 ( P2_U6599 , P2_U6570 , P2_REIP_REG_2_ );
nand NAND2_10676 ( P2_U6600 , P2_R2267_U17 , P2_U2587 );
nand NAND2_10677 ( P2_U6601 , P2_U2588 , P2_R2096_U75 );
nand NAND2_10678 ( P2_U6602 , P2_EBX_REG_3_ , P2_U7743 );
nand NAND2_10679 ( P2_U6603 , P2_U2437 , P2_R2182_U76 );
nand NAND2_10680 ( P2_U6604 , P2_U2392 , P2_R2099_U95 );
nand NAND2_10681 ( P2_U6605 , P2_U2383 , P2_R2337_U67 );
nand NAND2_10682 ( P2_U6606 , P2_R1957_U59 , P2_U2382 );
nand NAND2_10683 ( P2_U6607 , P2_U2378 , P2_PHYADDRPOINTER_REG_3_ );
nand NAND2_10684 ( P2_U6608 , P2_U6570 , P2_REIP_REG_3_ );
nand NAND2_10685 ( P2_U6609 , P2_R2267_U60 , P2_U2587 );
nand NAND2_10686 ( P2_U6610 , P2_U2588 , P2_R2096_U74 );
nand NAND2_10687 ( P2_U6611 , P2_EBX_REG_4_ , P2_U7743 );
nand NAND2_10688 ( P2_U6612 , P2_U2437 , P2_R2182_U75 );
nand NAND2_10689 ( P2_U6613 , P2_U2392 , P2_R2099_U98 );
nand NAND2_10690 ( P2_U6614 , P2_U2383 , P2_R2337_U66 );
nand NAND2_10691 ( P2_U6615 , P2_R1957_U18 , P2_U2382 );
nand NAND2_10692 ( P2_U6616 , P2_U2378 , P2_PHYADDRPOINTER_REG_4_ );
nand NAND2_10693 ( P2_U6617 , P2_U6570 , P2_REIP_REG_4_ );
nand NAND2_10694 ( P2_U6618 , P2_R2267_U18 , P2_U2587 );
nand NAND2_10695 ( P2_U6619 , P2_U2588 , P2_R2096_U73 );
nand NAND2_10696 ( P2_U6620 , P2_EBX_REG_5_ , P2_U7743 );
nand NAND2_10697 ( P2_U6621 , P2_U2437 , P2_R2182_U74 );
nand NAND2_10698 ( P2_U6622 , P2_U2392 , P2_R2099_U71 );
nand NAND2_10699 ( P2_U6623 , P2_U2383 , P2_R2337_U65 );
nand NAND2_10700 ( P2_U6624 , P2_R1957_U57 , P2_U2382 );
nand NAND2_10701 ( P2_U6625 , P2_U2378 , P2_PHYADDRPOINTER_REG_5_ );
nand NAND2_10702 ( P2_U6626 , P2_U6570 , P2_REIP_REG_5_ );
nand NAND2_10703 ( P2_U6627 , P2_R2267_U58 , P2_U2587 );
nand NAND2_10704 ( P2_U6628 , P2_U2588 , P2_R2096_U72 );
nand NAND2_10705 ( P2_U6629 , P2_EBX_REG_6_ , P2_U7743 );
nand NAND2_10706 ( P2_U6630 , P2_U2392 , P2_R2099_U70 );
nand NAND2_10707 ( P2_U6631 , P2_U2383 , P2_R2337_U64 );
nand NAND2_10708 ( P2_U6632 , P2_R1957_U19 , P2_U2382 );
nand NAND2_10709 ( P2_U6633 , P2_U2378 , P2_PHYADDRPOINTER_REG_6_ );
nand NAND2_10710 ( P2_U6634 , P2_U6570 , P2_REIP_REG_6_ );
nand NAND2_10711 ( P2_U6635 , P2_R2267_U19 , P2_U2587 );
nand NAND2_10712 ( P2_U6636 , P2_U2588 , P2_R2096_U71 );
nand NAND2_10713 ( P2_U6637 , P2_EBX_REG_7_ , P2_U7743 );
nand NAND2_10714 ( P2_U6638 , P2_U2392 , P2_R2099_U69 );
nand NAND2_10715 ( P2_U6639 , P2_U2383 , P2_R2337_U63 );
nand NAND2_10716 ( P2_U6640 , P2_R1957_U55 , P2_U2382 );
nand NAND2_10717 ( P2_U6641 , P2_U2378 , P2_PHYADDRPOINTER_REG_7_ );
nand NAND2_10718 ( P2_U6642 , P2_U6570 , P2_REIP_REG_7_ );
nand NAND2_10719 ( P2_U6643 , P2_R2267_U56 , P2_U2587 );
nand NAND2_10720 ( P2_U6644 , P2_U2588 , P2_R2096_U70 );
nand NAND2_10721 ( P2_U6645 , P2_EBX_REG_8_ , P2_U7743 );
nand NAND2_10722 ( P2_U6646 , P2_U2392 , P2_R2099_U68 );
nand NAND2_10723 ( P2_U6647 , P2_U2383 , P2_R2337_U62 );
nand NAND2_10724 ( P2_U6648 , P2_R1957_U20 , P2_U2382 );
nand NAND2_10725 ( P2_U6649 , P2_U2378 , P2_PHYADDRPOINTER_REG_8_ );
nand NAND2_10726 ( P2_U6650 , P2_U6570 , P2_REIP_REG_8_ );
nand NAND2_10727 ( P2_U6651 , P2_R2267_U20 , P2_U2587 );
nand NAND2_10728 ( P2_U6652 , P2_U2588 , P2_R2096_U69 );
nand NAND2_10729 ( P2_U6653 , P2_EBX_REG_9_ , P2_U7743 );
nand NAND2_10730 ( P2_U6654 , P2_U2392 , P2_R2099_U67 );
nand NAND2_10731 ( P2_U6655 , P2_U2383 , P2_R2337_U61 );
nand NAND2_10732 ( P2_U6656 , P2_R1957_U53 , P2_U2382 );
nand NAND2_10733 ( P2_U6657 , P2_U2378 , P2_PHYADDRPOINTER_REG_9_ );
nand NAND2_10734 ( P2_U6658 , P2_U6570 , P2_REIP_REG_9_ );
nand NAND2_10735 ( P2_U6659 , P2_R2267_U87 , P2_U2587 );
nand NAND2_10736 ( P2_U6660 , P2_U2588 , P2_R2096_U97 );
nand NAND2_10737 ( P2_U6661 , P2_EBX_REG_10_ , P2_U7743 );
nand NAND2_10738 ( P2_U6662 , P2_U2392 , P2_R2099_U93 );
nand NAND2_10739 ( P2_U6663 , P2_U2383 , P2_R2337_U90 );
nand NAND2_10740 ( P2_U6664 , P2_R1957_U6 , P2_U2382 );
nand NAND2_10741 ( P2_U6665 , P2_U2378 , P2_PHYADDRPOINTER_REG_10_ );
nand NAND2_10742 ( P2_U6666 , P2_U6570 , P2_REIP_REG_10_ );
nand NAND2_10743 ( P2_U6667 , P2_R2267_U6 , P2_U2587 );
nand NAND2_10744 ( P2_U6668 , P2_U2588 , P2_R2096_U96 );
nand NAND2_10745 ( P2_U6669 , P2_EBX_REG_11_ , P2_U7743 );
nand NAND2_10746 ( P2_U6670 , P2_U2392 , P2_R2099_U92 );
nand NAND2_10747 ( P2_U6671 , P2_U2383 , P2_R2337_U89 );
nand NAND2_10748 ( P2_U6672 , P2_R1957_U82 , P2_U2382 );
nand NAND2_10749 ( P2_U6673 , P2_U2378 , P2_PHYADDRPOINTER_REG_11_ );
nand NAND2_10750 ( P2_U6674 , P2_U6570 , P2_REIP_REG_11_ );
nand NAND2_10751 ( P2_U6675 , P2_R2267_U85 , P2_U2587 );
nand NAND2_10752 ( P2_U6676 , P2_U2588 , P2_R2096_U95 );
nand NAND2_10753 ( P2_U6677 , P2_EBX_REG_12_ , P2_U7743 );
nand NAND2_10754 ( P2_U6678 , P2_U2392 , P2_R2099_U91 );
nand NAND2_10755 ( P2_U6679 , P2_U2383 , P2_R2337_U88 );
nand NAND2_10756 ( P2_U6680 , P2_R1957_U7 , P2_U2382 );
nand NAND2_10757 ( P2_U6681 , P2_U2378 , P2_PHYADDRPOINTER_REG_12_ );
nand NAND2_10758 ( P2_U6682 , P2_U6570 , P2_REIP_REG_12_ );
nand NAND2_10759 ( P2_U6683 , P2_R2267_U7 , P2_U2587 );
nand NAND2_10760 ( P2_U6684 , P2_U2588 , P2_R2096_U94 );
nand NAND2_10761 ( P2_U6685 , P2_EBX_REG_13_ , P2_U7743 );
nand NAND2_10762 ( P2_U6686 , P2_U2392 , P2_R2099_U90 );
nand NAND2_10763 ( P2_U6687 , P2_U2383 , P2_R2337_U87 );
nand NAND2_10764 ( P2_U6688 , P2_R1957_U80 , P2_U2382 );
nand NAND2_10765 ( P2_U6689 , P2_U2378 , P2_PHYADDRPOINTER_REG_13_ );
nand NAND2_10766 ( P2_U6690 , P2_U6570 , P2_REIP_REG_13_ );
nand NAND2_10767 ( P2_U6691 , P2_R2267_U83 , P2_U2587 );
nand NAND2_10768 ( P2_U6692 , P2_U2588 , P2_R2096_U93 );
nand NAND2_10769 ( P2_U6693 , P2_EBX_REG_14_ , P2_U7743 );
nand NAND2_10770 ( P2_U6694 , P2_U2392 , P2_R2099_U89 );
nand NAND2_10771 ( P2_U6695 , P2_U2383 , P2_R2337_U86 );
nand NAND2_10772 ( P2_U6696 , P2_R1957_U8 , P2_U2382 );
nand NAND2_10773 ( P2_U6697 , P2_U2378 , P2_PHYADDRPOINTER_REG_14_ );
nand NAND2_10774 ( P2_U6698 , P2_U6570 , P2_REIP_REG_14_ );
nand NAND2_10775 ( P2_U6699 , P2_R2267_U8 , P2_U2587 );
nand NAND2_10776 ( P2_U6700 , P2_U2588 , P2_R2096_U92 );
nand NAND2_10777 ( P2_U6701 , P2_EBX_REG_15_ , P2_U7743 );
nand NAND2_10778 ( P2_U6702 , P2_U2392 , P2_R2099_U88 );
nand NAND2_10779 ( P2_U6703 , P2_U2383 , P2_R2337_U85 );
nand NAND2_10780 ( P2_U6704 , P2_R1957_U78 , P2_U2382 );
nand NAND2_10781 ( P2_U6705 , P2_U2378 , P2_PHYADDRPOINTER_REG_15_ );
nand NAND2_10782 ( P2_U6706 , P2_U6570 , P2_REIP_REG_15_ );
nand NAND2_10783 ( P2_U6707 , P2_R2267_U81 , P2_U2587 );
nand NAND2_10784 ( P2_U6708 , P2_U2588 , P2_R2096_U91 );
nand NAND2_10785 ( P2_U6709 , P2_EBX_REG_16_ , P2_U7743 );
nand NAND2_10786 ( P2_U6710 , P2_U2392 , P2_R2099_U87 );
nand NAND2_10787 ( P2_U6711 , P2_U2383 , P2_R2337_U84 );
nand NAND2_10788 ( P2_U6712 , P2_R1957_U9 , P2_U2382 );
nand NAND2_10789 ( P2_U6713 , P2_U2378 , P2_PHYADDRPOINTER_REG_16_ );
nand NAND2_10790 ( P2_U6714 , P2_U6570 , P2_REIP_REG_16_ );
nand NAND2_10791 ( P2_U6715 , P2_R2267_U9 , P2_U2587 );
nand NAND2_10792 ( P2_U6716 , P2_U2588 , P2_R2096_U90 );
nand NAND2_10793 ( P2_U6717 , P2_EBX_REG_17_ , P2_U7743 );
nand NAND2_10794 ( P2_U6718 , P2_U2392 , P2_R2099_U86 );
nand NAND2_10795 ( P2_U6719 , P2_U2383 , P2_R2337_U83 );
nand NAND2_10796 ( P2_U6720 , P2_R1957_U76 , P2_U2382 );
nand NAND2_10797 ( P2_U6721 , P2_U2378 , P2_PHYADDRPOINTER_REG_17_ );
nand NAND2_10798 ( P2_U6722 , P2_U6570 , P2_REIP_REG_17_ );
nand NAND2_10799 ( P2_U6723 , P2_R2267_U79 , P2_U2587 );
nand NAND2_10800 ( P2_U6724 , P2_U2588 , P2_R2096_U89 );
nand NAND2_10801 ( P2_U6725 , P2_EBX_REG_18_ , P2_U7743 );
nand NAND2_10802 ( P2_U6726 , P2_U2392 , P2_R2099_U85 );
nand NAND2_10803 ( P2_U6727 , P2_U2383 , P2_R2337_U82 );
nand NAND2_10804 ( P2_U6728 , P2_R1957_U10 , P2_U2382 );
nand NAND2_10805 ( P2_U6729 , P2_U2378 , P2_PHYADDRPOINTER_REG_18_ );
nand NAND2_10806 ( P2_U6730 , P2_U6570 , P2_REIP_REG_18_ );
nand NAND2_10807 ( P2_U6731 , P2_R2267_U10 , P2_U2587 );
nand NAND2_10808 ( P2_U6732 , P2_U2588 , P2_R2096_U88 );
nand NAND2_10809 ( P2_U6733 , P2_EBX_REG_19_ , P2_U7743 );
nand NAND2_10810 ( P2_U6734 , P2_U2392 , P2_R2099_U84 );
nand NAND2_10811 ( P2_U6735 , P2_U2383 , P2_R2337_U81 );
nand NAND2_10812 ( P2_U6736 , P2_R1957_U74 , P2_U2382 );
nand NAND2_10813 ( P2_U6737 , P2_U2378 , P2_PHYADDRPOINTER_REG_19_ );
nand NAND2_10814 ( P2_U6738 , P2_U6570 , P2_REIP_REG_19_ );
nand NAND2_10815 ( P2_U6739 , P2_R2267_U75 , P2_U2587 );
nand NAND2_10816 ( P2_U6740 , P2_U2588 , P2_R2096_U87 );
nand NAND2_10817 ( P2_U6741 , P2_EBX_REG_20_ , P2_U7743 );
nand NAND2_10818 ( P2_U6742 , P2_U2392 , P2_R2099_U83 );
nand NAND2_10819 ( P2_U6743 , P2_U2383 , P2_R2337_U80 );
nand NAND2_10820 ( P2_U6744 , P2_R1957_U11 , P2_U2382 );
nand NAND2_10821 ( P2_U6745 , P2_U2378 , P2_PHYADDRPOINTER_REG_20_ );
nand NAND2_10822 ( P2_U6746 , P2_U6570 , P2_REIP_REG_20_ );
nand NAND2_10823 ( P2_U6747 , P2_R2267_U11 , P2_U2587 );
nand NAND2_10824 ( P2_U6748 , P2_U2588 , P2_R2096_U86 );
nand NAND2_10825 ( P2_U6749 , P2_EBX_REG_21_ , P2_U7743 );
nand NAND2_10826 ( P2_U6750 , P2_U2392 , P2_R2099_U82 );
nand NAND2_10827 ( P2_U6751 , P2_U2383 , P2_R2337_U79 );
nand NAND2_10828 ( P2_U6752 , P2_R1957_U70 , P2_U2382 );
nand NAND2_10829 ( P2_U6753 , P2_U2378 , P2_PHYADDRPOINTER_REG_21_ );
nand NAND2_10830 ( P2_U6754 , P2_U6570 , P2_REIP_REG_21_ );
nand NAND2_10831 ( P2_U6755 , P2_R2267_U73 , P2_U2587 );
nand NAND2_10832 ( P2_U6756 , P2_U2588 , P2_R2096_U85 );
nand NAND2_10833 ( P2_U6757 , P2_EBX_REG_22_ , P2_U7743 );
nand NAND2_10834 ( P2_U6758 , P2_U2392 , P2_R2099_U81 );
nand NAND2_10835 ( P2_U6759 , P2_U2383 , P2_R2337_U78 );
nand NAND2_10836 ( P2_U6760 , P2_R1957_U12 , P2_U2382 );
nand NAND2_10837 ( P2_U6761 , P2_U2378 , P2_PHYADDRPOINTER_REG_22_ );
nand NAND2_10838 ( P2_U6762 , P2_U6570 , P2_REIP_REG_22_ );
nand NAND2_10839 ( P2_U6763 , P2_R2267_U12 , P2_U2587 );
nand NAND2_10840 ( P2_U6764 , P2_U2588 , P2_R2096_U84 );
nand NAND2_10841 ( P2_U6765 , P2_EBX_REG_23_ , P2_U7743 );
nand NAND2_10842 ( P2_U6766 , P2_U2392 , P2_R2099_U80 );
nand NAND2_10843 ( P2_U6767 , P2_U2383 , P2_R2337_U77 );
nand NAND2_10844 ( P2_U6768 , P2_R1957_U68 , P2_U2382 );
nand NAND2_10845 ( P2_U6769 , P2_U2378 , P2_PHYADDRPOINTER_REG_23_ );
nand NAND2_10846 ( P2_U6770 , P2_U6570 , P2_REIP_REG_23_ );
nand NAND2_10847 ( P2_U6771 , P2_R2267_U71 , P2_U2587 );
nand NAND2_10848 ( P2_U6772 , P2_U2588 , P2_R2096_U83 );
nand NAND2_10849 ( P2_U6773 , P2_EBX_REG_24_ , P2_U7743 );
nand NAND2_10850 ( P2_U6774 , P2_U2392 , P2_R2099_U79 );
nand NAND2_10851 ( P2_U6775 , P2_U2383 , P2_R2337_U76 );
nand NAND2_10852 ( P2_U6776 , P2_R1957_U13 , P2_U2382 );
nand NAND2_10853 ( P2_U6777 , P2_U2378 , P2_PHYADDRPOINTER_REG_24_ );
nand NAND2_10854 ( P2_U6778 , P2_U6570 , P2_REIP_REG_24_ );
nand NAND2_10855 ( P2_U6779 , P2_R2267_U13 , P2_U2587 );
nand NAND2_10856 ( P2_U6780 , P2_U2588 , P2_R2096_U82 );
nand NAND2_10857 ( P2_U6781 , P2_EBX_REG_25_ , P2_U7743 );
nand NAND2_10858 ( P2_U6782 , P2_U2392 , P2_R2099_U78 );
nand NAND2_10859 ( P2_U6783 , P2_U2383 , P2_R2337_U75 );
nand NAND2_10860 ( P2_U6784 , P2_R1957_U66 , P2_U2382 );
nand NAND2_10861 ( P2_U6785 , P2_U2378 , P2_PHYADDRPOINTER_REG_25_ );
nand NAND2_10862 ( P2_U6786 , P2_U6570 , P2_REIP_REG_25_ );
nand NAND2_10863 ( P2_U6787 , P2_R2267_U69 , P2_U2587 );
nand NAND2_10864 ( P2_U6788 , P2_U2588 , P2_R2096_U81 );
nand NAND2_10865 ( P2_U6789 , P2_EBX_REG_26_ , P2_U7743 );
nand NAND2_10866 ( P2_U6790 , P2_U2392 , P2_R2099_U77 );
nand NAND2_10867 ( P2_U6791 , P2_U2383 , P2_R2337_U74 );
nand NAND2_10868 ( P2_U6792 , P2_R1957_U14 , P2_U2382 );
nand NAND2_10869 ( P2_U6793 , P2_U2378 , P2_PHYADDRPOINTER_REG_26_ );
nand NAND2_10870 ( P2_U6794 , P2_U6570 , P2_REIP_REG_26_ );
nand NAND2_10871 ( P2_U6795 , P2_R2267_U14 , P2_U2587 );
nand NAND2_10872 ( P2_U6796 , P2_U2588 , P2_R2096_U80 );
nand NAND2_10873 ( P2_U6797 , P2_EBX_REG_27_ , P2_U7743 );
nand NAND2_10874 ( P2_U6798 , P2_U2392 , P2_R2099_U76 );
nand NAND2_10875 ( P2_U6799 , P2_U2383 , P2_R2337_U73 );
nand NAND2_10876 ( P2_U6800 , P2_R1957_U64 , P2_U2382 );
nand NAND2_10877 ( P2_U6801 , P2_U2378 , P2_PHYADDRPOINTER_REG_27_ );
nand NAND2_10878 ( P2_U6802 , P2_U6570 , P2_REIP_REG_27_ );
nand NAND2_10879 ( P2_U6803 , P2_R2267_U67 , P2_U2587 );
nand NAND2_10880 ( P2_U6804 , P2_U2588 , P2_R2096_U79 );
nand NAND2_10881 ( P2_U6805 , P2_EBX_REG_28_ , P2_U7743 );
nand NAND2_10882 ( P2_U6806 , P2_U2392 , P2_R2099_U75 );
nand NAND2_10883 ( P2_U6807 , P2_U2383 , P2_R2337_U72 );
nand NAND2_10884 ( P2_U6808 , P2_R1957_U15 , P2_U2382 );
nand NAND2_10885 ( P2_U6809 , P2_U2378 , P2_PHYADDRPOINTER_REG_28_ );
nand NAND2_10886 ( P2_U6810 , P2_U6570 , P2_REIP_REG_28_ );
nand NAND2_10887 ( P2_U6811 , P2_R2267_U15 , P2_U2587 );
nand NAND2_10888 ( P2_U6812 , P2_U2588 , P2_R2096_U78 );
nand NAND2_10889 ( P2_U6813 , P2_EBX_REG_29_ , P2_U7743 );
nand NAND2_10890 ( P2_U6814 , P2_U2392 , P2_R2099_U74 );
nand NAND2_10891 ( P2_U6815 , P2_U2383 , P2_R2337_U71 );
nand NAND2_10892 ( P2_U6816 , P2_R1957_U16 , P2_U2382 );
nand NAND2_10893 ( P2_U6817 , P2_U2378 , P2_PHYADDRPOINTER_REG_29_ );
nand NAND2_10894 ( P2_U6818 , P2_U6570 , P2_REIP_REG_29_ );
nand NAND2_10895 ( P2_U6819 , P2_R2267_U16 , P2_U2587 );
nand NAND2_10896 ( P2_U6820 , P2_U2588 , P2_R2096_U76 );
nand NAND2_10897 ( P2_U6821 , P2_EBX_REG_30_ , P2_U7743 );
nand NAND2_10898 ( P2_U6822 , P2_U2392 , P2_R2099_U73 );
nand NAND2_10899 ( P2_U6823 , P2_U2383 , P2_R2337_U69 );
nand NAND2_10900 ( P2_U6824 , P2_R1957_U62 , P2_U2382 );
nand NAND2_10901 ( P2_U6825 , P2_U2378 , P2_PHYADDRPOINTER_REG_30_ );
nand NAND2_10902 ( P2_U6826 , P2_U6570 , P2_REIP_REG_30_ );
nand NAND2_10903 ( P2_U6827 , P2_R2267_U63 , P2_U2587 );
nand NAND2_10904 ( P2_U6828 , P2_U2588 , P2_R2096_U50 );
nand NAND2_10905 ( P2_U6829 , P2_EBX_REG_31_ , P2_U7743 );
nand NAND2_10906 ( P2_U6830 , P2_U2392 , P2_R2099_U72 );
nand NAND2_10907 ( P2_U6831 , P2_U2383 , P2_R2337_U68 );
nand NAND2_10908 ( P2_U6832 , P2_R1957_U50 , P2_U2382 );
nand NAND2_10909 ( P2_U6833 , P2_U2378 , P2_PHYADDRPOINTER_REG_31_ );
nand NAND2_10910 ( P2_U6834 , P2_U6570 , P2_REIP_REG_31_ );
nand NAND2_10911 ( P2_U6835 , P2_DATAWIDTH_REG_1_ , P2_DATAWIDTH_REG_0_ );
nand NAND2_10912 ( P2_U6836 , P2_U4477 , P2_REIP_REG_0_ );
nand NAND2_10913 ( P2_U6837 , P2_BYTEENABLE_REG_1_ , P2_U3547 );
not NOT1_10914 ( P2_U6838 , P2_U4400 );
nand NAND3_10915 ( P2_U6839 , P2_U4426 , P2_U4468 , P2_U4399 );
nand NAND2_10916 ( P2_U6840 , P2_FLUSH_REG , P2_U4400 );
nand NAND2_10917 ( P2_U6841 , P2_U4187 , P2_U4467 );
nand NAND2_10918 ( P2_U6842 , P2_U4466 , P2_U3284 );
not NOT1_10919 ( P2_U6843 , P2_U4402 );
nand NAND2_10920 ( P2_U6844 , P2_U4411 , P2_STATEBS16_REG );
not NOT1_10921 ( P2_U6845 , P2_U2715 );
nand NAND2_10922 ( P2_U6846 , P2_U2715 , P2_U3536 );
nand NAND2_10923 ( P2_U6847 , P2_U4411 , P2_U3265 );
nand NAND2_10924 ( P2_U6848 , P2_U4184 , P2_U2356 );
nand NAND2_10925 ( P2_U6849 , P2_U4418 , P2_U6847 );
nand NAND2_10926 ( P2_U6850 , U211 , P2_U6846 );
or OR2_10927 ( P2_U6851 , P2_STATE2_REG_2_ , P2_STATE2_REG_1_ );
nand NAND3_10928 ( P2_U6852 , P2_U6851 , P2_U6850 , P2_U4186 );
nand NAND2_10929 ( P2_U6853 , P2_U2374 , P2_U2459 );
nand NAND2_10930 ( P2_U6854 , P2_CODEFETCH_REG , P2_U6853 );
nand NAND2_10931 ( P2_U6855 , P2_U4461 , P2_STATE2_REG_0_ );
nand NAND2_10932 ( P2_U6856 , P2_ADS_N_REG , P2_STATE_REG_0_ );
not NOT1_10933 ( P2_U6857 , P2_U4403 );
nand NAND3_10934 ( P2_U6858 , P2_STATE2_REG_2_ , P2_U3286 , P2_U3294 );
nand NAND3_10935 ( P2_U6859 , P2_U4421 , P2_U4468 , P2_U4404 );
nand NAND2_10936 ( P2_U6860 , P2_U4189 , P2_U2446 );
nand NAND2_10937 ( P2_U6861 , P2_MEMORYFETCH_REG , P2_U6859 );
nand NAND2_10938 ( P2_U6862 , P2_U2538 , P2_INSTQUEUE_REG_8__7_ );
nand NAND2_10939 ( P2_U6863 , P2_U2537 , P2_INSTQUEUE_REG_9__7_ );
nand NAND2_10940 ( P2_U6864 , P2_U2536 , P2_INSTQUEUE_REG_10__7_ );
nand NAND2_10941 ( P2_U6865 , P2_U2535 , P2_INSTQUEUE_REG_11__7_ );
nand NAND2_10942 ( P2_U6866 , P2_U2534 , P2_INSTQUEUE_REG_12__7_ );
nand NAND2_10943 ( P2_U6867 , P2_U2533 , P2_INSTQUEUE_REG_13__7_ );
nand NAND2_10944 ( P2_U6868 , P2_U2531 , P2_INSTQUEUE_REG_14__7_ );
nand NAND2_10945 ( P2_U6869 , P2_U2530 , P2_INSTQUEUE_REG_15__7_ );
nand NAND2_10946 ( P2_U6870 , P2_U2528 , P2_INSTQUEUE_REG_7__7_ );
nand NAND2_10947 ( P2_U6871 , P2_U2527 , P2_INSTQUEUE_REG_6__7_ );
nand NAND2_10948 ( P2_U6872 , P2_U2526 , P2_INSTQUEUE_REG_5__7_ );
nand NAND2_10949 ( P2_U6873 , P2_U2524 , P2_INSTQUEUE_REG_4__7_ );
nand NAND2_10950 ( P2_U6874 , P2_U2522 , P2_INSTQUEUE_REG_3__7_ );
nand NAND2_10951 ( P2_U6875 , P2_U2521 , P2_INSTQUEUE_REG_2__7_ );
nand NAND2_10952 ( P2_U6876 , P2_U2519 , P2_INSTQUEUE_REG_1__7_ );
nand NAND2_10953 ( P2_U6877 , P2_U2517 , P2_INSTQUEUE_REG_0__7_ );
nand NAND2_10954 ( P2_U6878 , P2_U2562 , P2_INSTQUEUE_REG_15__7_ );
nand NAND2_10955 ( P2_U6879 , P2_U2561 , P2_INSTQUEUE_REG_14__7_ );
nand NAND2_10956 ( P2_U6880 , P2_U2560 , P2_INSTQUEUE_REG_13__7_ );
nand NAND2_10957 ( P2_U6881 , P2_U2559 , P2_INSTQUEUE_REG_12__7_ );
nand NAND2_10958 ( P2_U6882 , P2_U2558 , P2_INSTQUEUE_REG_11__7_ );
nand NAND2_10959 ( P2_U6883 , P2_U2557 , P2_INSTQUEUE_REG_10__7_ );
nand NAND2_10960 ( P2_U6884 , P2_U2555 , P2_INSTQUEUE_REG_9__7_ );
nand NAND2_10961 ( P2_U6885 , P2_U2554 , P2_INSTQUEUE_REG_8__7_ );
nand NAND2_10962 ( P2_U6886 , P2_U2552 , P2_INSTQUEUE_REG_7__7_ );
nand NAND2_10963 ( P2_U6887 , P2_U2551 , P2_INSTQUEUE_REG_6__7_ );
nand NAND2_10964 ( P2_U6888 , P2_U2550 , P2_INSTQUEUE_REG_5__7_ );
nand NAND2_10965 ( P2_U6889 , P2_U2548 , P2_INSTQUEUE_REG_4__7_ );
nand NAND2_10966 ( P2_U6890 , P2_U2546 , P2_INSTQUEUE_REG_3__7_ );
nand NAND2_10967 ( P2_U6891 , P2_U2545 , P2_INSTQUEUE_REG_2__7_ );
nand NAND2_10968 ( P2_U6892 , P2_U2543 , P2_INSTQUEUE_REG_1__7_ );
nand NAND2_10969 ( P2_U6893 , P2_U2541 , P2_INSTQUEUE_REG_0__7_ );
nand NAND2_10970 ( P2_U6894 , P2_U2562 , P2_INSTQUEUE_REG_15__6_ );
nand NAND2_10971 ( P2_U6895 , P2_U2561 , P2_INSTQUEUE_REG_14__6_ );
nand NAND2_10972 ( P2_U6896 , P2_U2560 , P2_INSTQUEUE_REG_13__6_ );
nand NAND2_10973 ( P2_U6897 , P2_U2559 , P2_INSTQUEUE_REG_12__6_ );
nand NAND2_10974 ( P2_U6898 , P2_U2558 , P2_INSTQUEUE_REG_11__6_ );
nand NAND2_10975 ( P2_U6899 , P2_U2557 , P2_INSTQUEUE_REG_10__6_ );
nand NAND2_10976 ( P2_U6900 , P2_U2555 , P2_INSTQUEUE_REG_9__6_ );
nand NAND2_10977 ( P2_U6901 , P2_U2554 , P2_INSTQUEUE_REG_8__6_ );
nand NAND2_10978 ( P2_U6902 , P2_U2552 , P2_INSTQUEUE_REG_7__6_ );
nand NAND2_10979 ( P2_U6903 , P2_U2551 , P2_INSTQUEUE_REG_6__6_ );
nand NAND2_10980 ( P2_U6904 , P2_U2550 , P2_INSTQUEUE_REG_5__6_ );
nand NAND2_10981 ( P2_U6905 , P2_U2548 , P2_INSTQUEUE_REG_4__6_ );
nand NAND2_10982 ( P2_U6906 , P2_U2546 , P2_INSTQUEUE_REG_3__6_ );
nand NAND2_10983 ( P2_U6907 , P2_U2545 , P2_INSTQUEUE_REG_2__6_ );
nand NAND2_10984 ( P2_U6908 , P2_U2543 , P2_INSTQUEUE_REG_1__6_ );
nand NAND2_10985 ( P2_U6909 , P2_U2541 , P2_INSTQUEUE_REG_0__6_ );
nand NAND2_10986 ( P2_U6910 , P2_U2562 , P2_INSTQUEUE_REG_15__5_ );
nand NAND2_10987 ( P2_U6911 , P2_U2561 , P2_INSTQUEUE_REG_14__5_ );
nand NAND2_10988 ( P2_U6912 , P2_U2560 , P2_INSTQUEUE_REG_13__5_ );
nand NAND2_10989 ( P2_U6913 , P2_U2559 , P2_INSTQUEUE_REG_12__5_ );
nand NAND2_10990 ( P2_U6914 , P2_U2558 , P2_INSTQUEUE_REG_11__5_ );
nand NAND2_10991 ( P2_U6915 , P2_U2557 , P2_INSTQUEUE_REG_10__5_ );
nand NAND2_10992 ( P2_U6916 , P2_U2555 , P2_INSTQUEUE_REG_9__5_ );
nand NAND2_10993 ( P2_U6917 , P2_U2554 , P2_INSTQUEUE_REG_8__5_ );
nand NAND2_10994 ( P2_U6918 , P2_U2552 , P2_INSTQUEUE_REG_7__5_ );
nand NAND2_10995 ( P2_U6919 , P2_U2551 , P2_INSTQUEUE_REG_6__5_ );
nand NAND2_10996 ( P2_U6920 , P2_U2550 , P2_INSTQUEUE_REG_5__5_ );
nand NAND2_10997 ( P2_U6921 , P2_U2548 , P2_INSTQUEUE_REG_4__5_ );
nand NAND2_10998 ( P2_U6922 , P2_U2546 , P2_INSTQUEUE_REG_3__5_ );
nand NAND2_10999 ( P2_U6923 , P2_U2545 , P2_INSTQUEUE_REG_2__5_ );
nand NAND2_11000 ( P2_U6924 , P2_U2543 , P2_INSTQUEUE_REG_1__5_ );
nand NAND2_11001 ( P2_U6925 , P2_U2541 , P2_INSTQUEUE_REG_0__5_ );
nand NAND2_11002 ( P2_U6926 , P2_U2562 , P2_INSTQUEUE_REG_15__4_ );
nand NAND2_11003 ( P2_U6927 , P2_U2561 , P2_INSTQUEUE_REG_14__4_ );
nand NAND2_11004 ( P2_U6928 , P2_U2560 , P2_INSTQUEUE_REG_13__4_ );
nand NAND2_11005 ( P2_U6929 , P2_U2559 , P2_INSTQUEUE_REG_12__4_ );
nand NAND2_11006 ( P2_U6930 , P2_U2558 , P2_INSTQUEUE_REG_11__4_ );
nand NAND2_11007 ( P2_U6931 , P2_U2557 , P2_INSTQUEUE_REG_10__4_ );
nand NAND2_11008 ( P2_U6932 , P2_U2555 , P2_INSTQUEUE_REG_9__4_ );
nand NAND2_11009 ( P2_U6933 , P2_U2554 , P2_INSTQUEUE_REG_8__4_ );
nand NAND2_11010 ( P2_U6934 , P2_U2552 , P2_INSTQUEUE_REG_7__4_ );
nand NAND2_11011 ( P2_U6935 , P2_U2551 , P2_INSTQUEUE_REG_6__4_ );
nand NAND2_11012 ( P2_U6936 , P2_U2550 , P2_INSTQUEUE_REG_5__4_ );
nand NAND2_11013 ( P2_U6937 , P2_U2548 , P2_INSTQUEUE_REG_4__4_ );
nand NAND2_11014 ( P2_U6938 , P2_U2546 , P2_INSTQUEUE_REG_3__4_ );
nand NAND2_11015 ( P2_U6939 , P2_U2545 , P2_INSTQUEUE_REG_2__4_ );
nand NAND2_11016 ( P2_U6940 , P2_U2543 , P2_INSTQUEUE_REG_1__4_ );
nand NAND2_11017 ( P2_U6941 , P2_U2541 , P2_INSTQUEUE_REG_0__4_ );
nand NAND2_11018 ( P2_U6942 , P2_U2562 , P2_INSTQUEUE_REG_15__3_ );
nand NAND2_11019 ( P2_U6943 , P2_U2561 , P2_INSTQUEUE_REG_14__3_ );
nand NAND2_11020 ( P2_U6944 , P2_U2560 , P2_INSTQUEUE_REG_13__3_ );
nand NAND2_11021 ( P2_U6945 , P2_U2559 , P2_INSTQUEUE_REG_12__3_ );
nand NAND2_11022 ( P2_U6946 , P2_U2558 , P2_INSTQUEUE_REG_11__3_ );
nand NAND2_11023 ( P2_U6947 , P2_U2557 , P2_INSTQUEUE_REG_10__3_ );
nand NAND2_11024 ( P2_U6948 , P2_U2555 , P2_INSTQUEUE_REG_9__3_ );
nand NAND2_11025 ( P2_U6949 , P2_U2554 , P2_INSTQUEUE_REG_8__3_ );
nand NAND2_11026 ( P2_U6950 , P2_U2552 , P2_INSTQUEUE_REG_7__3_ );
nand NAND2_11027 ( P2_U6951 , P2_U2551 , P2_INSTQUEUE_REG_6__3_ );
nand NAND2_11028 ( P2_U6952 , P2_U2550 , P2_INSTQUEUE_REG_5__3_ );
nand NAND2_11029 ( P2_U6953 , P2_U2548 , P2_INSTQUEUE_REG_4__3_ );
nand NAND2_11030 ( P2_U6954 , P2_U2546 , P2_INSTQUEUE_REG_3__3_ );
nand NAND2_11031 ( P2_U6955 , P2_U2545 , P2_INSTQUEUE_REG_2__3_ );
nand NAND2_11032 ( P2_U6956 , P2_U2543 , P2_INSTQUEUE_REG_1__3_ );
nand NAND2_11033 ( P2_U6957 , P2_U2541 , P2_INSTQUEUE_REG_0__3_ );
nand NAND2_11034 ( P2_U6958 , P2_U2562 , P2_INSTQUEUE_REG_15__2_ );
nand NAND2_11035 ( P2_U6959 , P2_U2561 , P2_INSTQUEUE_REG_14__2_ );
nand NAND2_11036 ( P2_U6960 , P2_U2560 , P2_INSTQUEUE_REG_13__2_ );
nand NAND2_11037 ( P2_U6961 , P2_U2559 , P2_INSTQUEUE_REG_12__2_ );
nand NAND2_11038 ( P2_U6962 , P2_U2558 , P2_INSTQUEUE_REG_11__2_ );
nand NAND2_11039 ( P2_U6963 , P2_U2557 , P2_INSTQUEUE_REG_10__2_ );
nand NAND2_11040 ( P2_U6964 , P2_U2555 , P2_INSTQUEUE_REG_9__2_ );
nand NAND2_11041 ( P2_U6965 , P2_U2554 , P2_INSTQUEUE_REG_8__2_ );
nand NAND2_11042 ( P2_U6966 , P2_U2552 , P2_INSTQUEUE_REG_7__2_ );
nand NAND2_11043 ( P2_U6967 , P2_U2551 , P2_INSTQUEUE_REG_6__2_ );
nand NAND2_11044 ( P2_U6968 , P2_U2550 , P2_INSTQUEUE_REG_5__2_ );
nand NAND2_11045 ( P2_U6969 , P2_U2548 , P2_INSTQUEUE_REG_4__2_ );
nand NAND2_11046 ( P2_U6970 , P2_U2546 , P2_INSTQUEUE_REG_3__2_ );
nand NAND2_11047 ( P2_U6971 , P2_U2545 , P2_INSTQUEUE_REG_2__2_ );
nand NAND2_11048 ( P2_U6972 , P2_U2543 , P2_INSTQUEUE_REG_1__2_ );
nand NAND2_11049 ( P2_U6973 , P2_U2541 , P2_INSTQUEUE_REG_0__2_ );
nand NAND2_11050 ( P2_U6974 , P2_U2562 , P2_INSTQUEUE_REG_15__1_ );
nand NAND2_11051 ( P2_U6975 , P2_U2561 , P2_INSTQUEUE_REG_14__1_ );
nand NAND2_11052 ( P2_U6976 , P2_U2560 , P2_INSTQUEUE_REG_13__1_ );
nand NAND2_11053 ( P2_U6977 , P2_U2559 , P2_INSTQUEUE_REG_12__1_ );
nand NAND2_11054 ( P2_U6978 , P2_U2558 , P2_INSTQUEUE_REG_11__1_ );
nand NAND2_11055 ( P2_U6979 , P2_U2557 , P2_INSTQUEUE_REG_10__1_ );
nand NAND2_11056 ( P2_U6980 , P2_U2555 , P2_INSTQUEUE_REG_9__1_ );
nand NAND2_11057 ( P2_U6981 , P2_U2554 , P2_INSTQUEUE_REG_8__1_ );
nand NAND2_11058 ( P2_U6982 , P2_U2552 , P2_INSTQUEUE_REG_7__1_ );
nand NAND2_11059 ( P2_U6983 , P2_U2551 , P2_INSTQUEUE_REG_6__1_ );
nand NAND2_11060 ( P2_U6984 , P2_U2550 , P2_INSTQUEUE_REG_5__1_ );
nand NAND2_11061 ( P2_U6985 , P2_U2548 , P2_INSTQUEUE_REG_4__1_ );
nand NAND2_11062 ( P2_U6986 , P2_U2546 , P2_INSTQUEUE_REG_3__1_ );
nand NAND2_11063 ( P2_U6987 , P2_U2545 , P2_INSTQUEUE_REG_2__1_ );
nand NAND2_11064 ( P2_U6988 , P2_U2543 , P2_INSTQUEUE_REG_1__1_ );
nand NAND2_11065 ( P2_U6989 , P2_U2541 , P2_INSTQUEUE_REG_0__1_ );
nand NAND2_11066 ( P2_U6990 , P2_U2562 , P2_INSTQUEUE_REG_15__0_ );
nand NAND2_11067 ( P2_U6991 , P2_U2561 , P2_INSTQUEUE_REG_14__0_ );
nand NAND2_11068 ( P2_U6992 , P2_U2560 , P2_INSTQUEUE_REG_13__0_ );
nand NAND2_11069 ( P2_U6993 , P2_U2559 , P2_INSTQUEUE_REG_12__0_ );
nand NAND2_11070 ( P2_U6994 , P2_U2558 , P2_INSTQUEUE_REG_11__0_ );
nand NAND2_11071 ( P2_U6995 , P2_U2557 , P2_INSTQUEUE_REG_10__0_ );
nand NAND2_11072 ( P2_U6996 , P2_U2555 , P2_INSTQUEUE_REG_9__0_ );
nand NAND2_11073 ( P2_U6997 , P2_U2554 , P2_INSTQUEUE_REG_8__0_ );
nand NAND2_11074 ( P2_U6998 , P2_U2552 , P2_INSTQUEUE_REG_7__0_ );
nand NAND2_11075 ( P2_U6999 , P2_U2551 , P2_INSTQUEUE_REG_6__0_ );
nand NAND2_11076 ( P2_U7000 , P2_U2550 , P2_INSTQUEUE_REG_5__0_ );
nand NAND2_11077 ( P2_U7001 , P2_U2548 , P2_INSTQUEUE_REG_4__0_ );
nand NAND2_11078 ( P2_U7002 , P2_U2546 , P2_INSTQUEUE_REG_3__0_ );
nand NAND2_11079 ( P2_U7003 , P2_U2545 , P2_INSTQUEUE_REG_2__0_ );
nand NAND2_11080 ( P2_U7004 , P2_U2543 , P2_INSTQUEUE_REG_1__0_ );
nand NAND2_11081 ( P2_U7005 , P2_U2541 , P2_INSTQUEUE_REG_0__0_ );
or OR2_11082 ( P2_U7006 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_11083 ( P2_U7007 , P2_U4405 );
nand NAND2_11084 ( P2_U7008 , P2_U2586 , P2_INSTQUEUE_REG_0__7_ );
nand NAND2_11085 ( P2_U7009 , P2_U2585 , P2_INSTQUEUE_REG_1__7_ );
nand NAND2_11086 ( P2_U7010 , P2_U2584 , P2_INSTQUEUE_REG_2__7_ );
nand NAND2_11087 ( P2_U7011 , P2_U2583 , P2_INSTQUEUE_REG_3__7_ );
nand NAND2_11088 ( P2_U7012 , P2_U2581 , P2_INSTQUEUE_REG_4__7_ );
nand NAND2_11089 ( P2_U7013 , P2_U2580 , P2_INSTQUEUE_REG_5__7_ );
nand NAND2_11090 ( P2_U7014 , P2_U2579 , P2_INSTQUEUE_REG_6__7_ );
nand NAND2_11091 ( P2_U7015 , P2_U2578 , P2_INSTQUEUE_REG_7__7_ );
nand NAND2_11092 ( P2_U7016 , P2_U2576 , P2_INSTQUEUE_REG_8__7_ );
nand NAND2_11093 ( P2_U7017 , P2_U2575 , P2_INSTQUEUE_REG_9__7_ );
nand NAND2_11094 ( P2_U7018 , P2_U2574 , P2_INSTQUEUE_REG_10__7_ );
nand NAND2_11095 ( P2_U7019 , P2_U2573 , P2_INSTQUEUE_REG_11__7_ );
nand NAND2_11096 ( P2_U7020 , P2_U2571 , P2_INSTQUEUE_REG_12__7_ );
nand NAND2_11097 ( P2_U7021 , P2_U2569 , P2_INSTQUEUE_REG_13__7_ );
nand NAND2_11098 ( P2_U7022 , P2_U2567 , P2_INSTQUEUE_REG_14__7_ );
nand NAND2_11099 ( P2_U7023 , P2_U2565 , P2_INSTQUEUE_REG_15__7_ );
nand NAND2_11100 ( P2_U7024 , P2_U2586 , P2_INSTQUEUE_REG_0__6_ );
nand NAND2_11101 ( P2_U7025 , P2_U2585 , P2_INSTQUEUE_REG_1__6_ );
nand NAND2_11102 ( P2_U7026 , P2_U2584 , P2_INSTQUEUE_REG_2__6_ );
nand NAND2_11103 ( P2_U7027 , P2_U2583 , P2_INSTQUEUE_REG_3__6_ );
nand NAND2_11104 ( P2_U7028 , P2_U2581 , P2_INSTQUEUE_REG_4__6_ );
nand NAND2_11105 ( P2_U7029 , P2_U2580 , P2_INSTQUEUE_REG_5__6_ );
nand NAND2_11106 ( P2_U7030 , P2_U2579 , P2_INSTQUEUE_REG_6__6_ );
nand NAND2_11107 ( P2_U7031 , P2_U2578 , P2_INSTQUEUE_REG_7__6_ );
nand NAND2_11108 ( P2_U7032 , P2_U2576 , P2_INSTQUEUE_REG_8__6_ );
nand NAND2_11109 ( P2_U7033 , P2_U2575 , P2_INSTQUEUE_REG_9__6_ );
nand NAND2_11110 ( P2_U7034 , P2_U2574 , P2_INSTQUEUE_REG_10__6_ );
nand NAND2_11111 ( P2_U7035 , P2_U2573 , P2_INSTQUEUE_REG_11__6_ );
nand NAND2_11112 ( P2_U7036 , P2_U2571 , P2_INSTQUEUE_REG_12__6_ );
nand NAND2_11113 ( P2_U7037 , P2_U2569 , P2_INSTQUEUE_REG_13__6_ );
nand NAND2_11114 ( P2_U7038 , P2_U2567 , P2_INSTQUEUE_REG_14__6_ );
nand NAND2_11115 ( P2_U7039 , P2_U2565 , P2_INSTQUEUE_REG_15__6_ );
nand NAND2_11116 ( P2_U7040 , P2_U2586 , P2_INSTQUEUE_REG_0__5_ );
nand NAND2_11117 ( P2_U7041 , P2_U2585 , P2_INSTQUEUE_REG_1__5_ );
nand NAND2_11118 ( P2_U7042 , P2_U2584 , P2_INSTQUEUE_REG_2__5_ );
nand NAND2_11119 ( P2_U7043 , P2_U2583 , P2_INSTQUEUE_REG_3__5_ );
nand NAND2_11120 ( P2_U7044 , P2_U2581 , P2_INSTQUEUE_REG_4__5_ );
nand NAND2_11121 ( P2_U7045 , P2_U2580 , P2_INSTQUEUE_REG_5__5_ );
nand NAND2_11122 ( P2_U7046 , P2_U2579 , P2_INSTQUEUE_REG_6__5_ );
nand NAND2_11123 ( P2_U7047 , P2_U2578 , P2_INSTQUEUE_REG_7__5_ );
nand NAND2_11124 ( P2_U7048 , P2_U2576 , P2_INSTQUEUE_REG_8__5_ );
nand NAND2_11125 ( P2_U7049 , P2_U2575 , P2_INSTQUEUE_REG_9__5_ );
nand NAND2_11126 ( P2_U7050 , P2_U2574 , P2_INSTQUEUE_REG_10__5_ );
nand NAND2_11127 ( P2_U7051 , P2_U2573 , P2_INSTQUEUE_REG_11__5_ );
nand NAND2_11128 ( P2_U7052 , P2_U2571 , P2_INSTQUEUE_REG_12__5_ );
nand NAND2_11129 ( P2_U7053 , P2_U2569 , P2_INSTQUEUE_REG_13__5_ );
nand NAND2_11130 ( P2_U7054 , P2_U2567 , P2_INSTQUEUE_REG_14__5_ );
nand NAND2_11131 ( P2_U7055 , P2_U2565 , P2_INSTQUEUE_REG_15__5_ );
nand NAND2_11132 ( P2_U7056 , P2_U2586 , P2_INSTQUEUE_REG_0__4_ );
nand NAND2_11133 ( P2_U7057 , P2_U2585 , P2_INSTQUEUE_REG_1__4_ );
nand NAND2_11134 ( P2_U7058 , P2_U2584 , P2_INSTQUEUE_REG_2__4_ );
nand NAND2_11135 ( P2_U7059 , P2_U2583 , P2_INSTQUEUE_REG_3__4_ );
nand NAND2_11136 ( P2_U7060 , P2_U2581 , P2_INSTQUEUE_REG_4__4_ );
nand NAND2_11137 ( P2_U7061 , P2_U2580 , P2_INSTQUEUE_REG_5__4_ );
nand NAND2_11138 ( P2_U7062 , P2_U2579 , P2_INSTQUEUE_REG_6__4_ );
nand NAND2_11139 ( P2_U7063 , P2_U2578 , P2_INSTQUEUE_REG_7__4_ );
nand NAND2_11140 ( P2_U7064 , P2_U2576 , P2_INSTQUEUE_REG_8__4_ );
nand NAND2_11141 ( P2_U7065 , P2_U2575 , P2_INSTQUEUE_REG_9__4_ );
nand NAND2_11142 ( P2_U7066 , P2_U2574 , P2_INSTQUEUE_REG_10__4_ );
nand NAND2_11143 ( P2_U7067 , P2_U2573 , P2_INSTQUEUE_REG_11__4_ );
nand NAND2_11144 ( P2_U7068 , P2_U2571 , P2_INSTQUEUE_REG_12__4_ );
nand NAND2_11145 ( P2_U7069 , P2_U2569 , P2_INSTQUEUE_REG_13__4_ );
nand NAND2_11146 ( P2_U7070 , P2_U2567 , P2_INSTQUEUE_REG_14__4_ );
nand NAND2_11147 ( P2_U7071 , P2_U2565 , P2_INSTQUEUE_REG_15__4_ );
nand NAND2_11148 ( P2_U7072 , P2_U2586 , P2_INSTQUEUE_REG_0__3_ );
nand NAND2_11149 ( P2_U7073 , P2_U2585 , P2_INSTQUEUE_REG_1__3_ );
nand NAND2_11150 ( P2_U7074 , P2_U2584 , P2_INSTQUEUE_REG_2__3_ );
nand NAND2_11151 ( P2_U7075 , P2_U2583 , P2_INSTQUEUE_REG_3__3_ );
nand NAND2_11152 ( P2_U7076 , P2_U2581 , P2_INSTQUEUE_REG_4__3_ );
nand NAND2_11153 ( P2_U7077 , P2_U2580 , P2_INSTQUEUE_REG_5__3_ );
nand NAND2_11154 ( P2_U7078 , P2_U2579 , P2_INSTQUEUE_REG_6__3_ );
nand NAND2_11155 ( P2_U7079 , P2_U2578 , P2_INSTQUEUE_REG_7__3_ );
nand NAND2_11156 ( P2_U7080 , P2_U2576 , P2_INSTQUEUE_REG_8__3_ );
nand NAND2_11157 ( P2_U7081 , P2_U2575 , P2_INSTQUEUE_REG_9__3_ );
nand NAND2_11158 ( P2_U7082 , P2_U2574 , P2_INSTQUEUE_REG_10__3_ );
nand NAND2_11159 ( P2_U7083 , P2_U2573 , P2_INSTQUEUE_REG_11__3_ );
nand NAND2_11160 ( P2_U7084 , P2_U2571 , P2_INSTQUEUE_REG_12__3_ );
nand NAND2_11161 ( P2_U7085 , P2_U2569 , P2_INSTQUEUE_REG_13__3_ );
nand NAND2_11162 ( P2_U7086 , P2_U2567 , P2_INSTQUEUE_REG_14__3_ );
nand NAND2_11163 ( P2_U7087 , P2_U2565 , P2_INSTQUEUE_REG_15__3_ );
nand NAND2_11164 ( P2_U7088 , P2_U2586 , P2_INSTQUEUE_REG_0__2_ );
nand NAND2_11165 ( P2_U7089 , P2_U2585 , P2_INSTQUEUE_REG_1__2_ );
nand NAND2_11166 ( P2_U7090 , P2_U2584 , P2_INSTQUEUE_REG_2__2_ );
nand NAND2_11167 ( P2_U7091 , P2_U2583 , P2_INSTQUEUE_REG_3__2_ );
nand NAND2_11168 ( P2_U7092 , P2_U2581 , P2_INSTQUEUE_REG_4__2_ );
nand NAND2_11169 ( P2_U7093 , P2_U2580 , P2_INSTQUEUE_REG_5__2_ );
nand NAND2_11170 ( P2_U7094 , P2_U2579 , P2_INSTQUEUE_REG_6__2_ );
nand NAND2_11171 ( P2_U7095 , P2_U2578 , P2_INSTQUEUE_REG_7__2_ );
nand NAND2_11172 ( P2_U7096 , P2_U2576 , P2_INSTQUEUE_REG_8__2_ );
nand NAND2_11173 ( P2_U7097 , P2_U2575 , P2_INSTQUEUE_REG_9__2_ );
nand NAND2_11174 ( P2_U7098 , P2_U2574 , P2_INSTQUEUE_REG_10__2_ );
nand NAND2_11175 ( P2_U7099 , P2_U2573 , P2_INSTQUEUE_REG_11__2_ );
nand NAND2_11176 ( P2_U7100 , P2_U2571 , P2_INSTQUEUE_REG_12__2_ );
nand NAND2_11177 ( P2_U7101 , P2_U2569 , P2_INSTQUEUE_REG_13__2_ );
nand NAND2_11178 ( P2_U7102 , P2_U2567 , P2_INSTQUEUE_REG_14__2_ );
nand NAND2_11179 ( P2_U7103 , P2_U2565 , P2_INSTQUEUE_REG_15__2_ );
nand NAND2_11180 ( P2_U7104 , P2_U2586 , P2_INSTQUEUE_REG_0__1_ );
nand NAND2_11181 ( P2_U7105 , P2_U2585 , P2_INSTQUEUE_REG_1__1_ );
nand NAND2_11182 ( P2_U7106 , P2_U2584 , P2_INSTQUEUE_REG_2__1_ );
nand NAND2_11183 ( P2_U7107 , P2_U2583 , P2_INSTQUEUE_REG_3__1_ );
nand NAND2_11184 ( P2_U7108 , P2_U2581 , P2_INSTQUEUE_REG_4__1_ );
nand NAND2_11185 ( P2_U7109 , P2_U2580 , P2_INSTQUEUE_REG_5__1_ );
nand NAND2_11186 ( P2_U7110 , P2_U2579 , P2_INSTQUEUE_REG_6__1_ );
nand NAND2_11187 ( P2_U7111 , P2_U2578 , P2_INSTQUEUE_REG_7__1_ );
nand NAND2_11188 ( P2_U7112 , P2_U2576 , P2_INSTQUEUE_REG_8__1_ );
nand NAND2_11189 ( P2_U7113 , P2_U2575 , P2_INSTQUEUE_REG_9__1_ );
nand NAND2_11190 ( P2_U7114 , P2_U2574 , P2_INSTQUEUE_REG_10__1_ );
nand NAND2_11191 ( P2_U7115 , P2_U2573 , P2_INSTQUEUE_REG_11__1_ );
nand NAND2_11192 ( P2_U7116 , P2_U2571 , P2_INSTQUEUE_REG_12__1_ );
nand NAND2_11193 ( P2_U7117 , P2_U2569 , P2_INSTQUEUE_REG_13__1_ );
nand NAND2_11194 ( P2_U7118 , P2_U2567 , P2_INSTQUEUE_REG_14__1_ );
nand NAND2_11195 ( P2_U7119 , P2_U2565 , P2_INSTQUEUE_REG_15__1_ );
nand NAND2_11196 ( P2_U7120 , P2_U2586 , P2_INSTQUEUE_REG_0__0_ );
nand NAND2_11197 ( P2_U7121 , P2_U2585 , P2_INSTQUEUE_REG_1__0_ );
nand NAND2_11198 ( P2_U7122 , P2_U2584 , P2_INSTQUEUE_REG_2__0_ );
nand NAND2_11199 ( P2_U7123 , P2_U2583 , P2_INSTQUEUE_REG_3__0_ );
nand NAND2_11200 ( P2_U7124 , P2_U2581 , P2_INSTQUEUE_REG_4__0_ );
nand NAND2_11201 ( P2_U7125 , P2_U2580 , P2_INSTQUEUE_REG_5__0_ );
nand NAND2_11202 ( P2_U7126 , P2_U2579 , P2_INSTQUEUE_REG_6__0_ );
nand NAND2_11203 ( P2_U7127 , P2_U2578 , P2_INSTQUEUE_REG_7__0_ );
nand NAND2_11204 ( P2_U7128 , P2_U2576 , P2_INSTQUEUE_REG_8__0_ );
nand NAND2_11205 ( P2_U7129 , P2_U2575 , P2_INSTQUEUE_REG_9__0_ );
nand NAND2_11206 ( P2_U7130 , P2_U2574 , P2_INSTQUEUE_REG_10__0_ );
nand NAND2_11207 ( P2_U7131 , P2_U2573 , P2_INSTQUEUE_REG_11__0_ );
nand NAND2_11208 ( P2_U7132 , P2_U2571 , P2_INSTQUEUE_REG_12__0_ );
nand NAND2_11209 ( P2_U7133 , P2_U2569 , P2_INSTQUEUE_REG_13__0_ );
nand NAND2_11210 ( P2_U7134 , P2_U2567 , P2_INSTQUEUE_REG_14__0_ );
nand NAND2_11211 ( P2_U7135 , P2_U2565 , P2_INSTQUEUE_REG_15__0_ );
not NOT1_11212 ( P2_U7136 , P2_U3554 );
nand NAND2_11213 ( P2_U7137 , P2_U7136 , P2_U3300 );
nand NAND2_11214 ( P2_U7138 , P2_U4467 , P2_R2099_U95 );
nand NAND2_11215 ( P2_U7139 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U7137 );
nand NAND2_11216 ( P2_U7140 , P2_U4430 , P2_U3428 );
nand NAND2_11217 ( P2_U7141 , P2_ADD_402_1132_U23 , P2_U2355 );
nand NAND2_11218 ( P2_U7142 , P2_U2354 , P2_U2606 );
nand NAND2_11219 ( P2_U7143 , P2_U2605 , P2_U2355 );
nand NAND2_11220 ( P2_U7144 , P2_U2354 , P2_U2605 );
nand NAND2_11221 ( P2_U7145 , P2_U2604 , P2_U2355 );
nand NAND2_11222 ( P2_U7146 , P2_U2354 , P2_U2604 );
nand NAND2_11223 ( P2_U7147 , P2_U2603 , P2_U2355 );
nand NAND2_11224 ( P2_U7148 , P2_U2354 , P2_U2603 );
nand NAND2_11225 ( P2_U7149 , P2_U4467 , P2_R2099_U96 );
nand NAND2_11226 ( P2_U7150 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_U7137 );
nand NAND2_11227 ( P2_U7151 , P2_U4430 , P2_U3580 );
nand NAND2_11228 ( P2_U7152 , P2_U2602 , P2_U2355 );
nand NAND2_11229 ( P2_U7153 , P2_U2354 , P2_U2602 );
nand NAND2_11230 ( P2_U7154 , P2_U2601 , P2_U2355 );
nand NAND2_11231 ( P2_U7155 , P2_U2354 , P2_U2601 );
nand NAND2_11232 ( P2_U7156 , P2_U2600 , P2_U2355 );
nand NAND2_11233 ( P2_U7157 , P2_U2354 , P2_U2600 );
nand NAND2_11234 ( P2_U7158 , P2_U2599 , P2_U2355 );
nand NAND2_11235 ( P2_U7159 , P2_U2354 , P2_U2599 );
nand NAND2_11236 ( P2_U7160 , P2_U4467 , P2_R2099_U5 );
nand NAND2_11237 ( P2_U7161 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_U7137 );
nand NAND2_11238 ( P2_U7162 , P2_U4430 , P2_U3243 );
nand NAND2_11239 ( P2_U7163 , P2_U4467 , P2_R2099_U94 );
nand NAND2_11240 ( P2_U7164 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_U7137 );
nand NAND2_11241 ( P2_U7165 , P2_U4430 , P2_U3307 );
nand NAND2_11242 ( P2_U7166 , P2_INSTQUEUE_REG_0__0_ , P2_U2355 );
nand NAND2_11243 ( P2_U7167 , P2_U5517 , P2_INSTQUEUE_REG_0__7_ );
nand NAND2_11244 ( P2_U7168 , P2_U5460 , P2_INSTQUEUE_REG_1__7_ );
nand NAND2_11245 ( P2_U7169 , P2_U5402 , P2_INSTQUEUE_REG_2__7_ );
nand NAND2_11246 ( P2_U7170 , P2_U5345 , P2_INSTQUEUE_REG_3__7_ );
nand NAND2_11247 ( P2_U7171 , P2_U5287 , P2_INSTQUEUE_REG_4__7_ );
nand NAND2_11248 ( P2_U7172 , P2_U5230 , P2_INSTQUEUE_REG_5__7_ );
nand NAND2_11249 ( P2_U7173 , P2_U5172 , P2_INSTQUEUE_REG_6__7_ );
nand NAND2_11250 ( P2_U7174 , P2_U5116 , P2_INSTQUEUE_REG_7__7_ );
nand NAND2_11251 ( P2_U7175 , P2_U5059 , P2_INSTQUEUE_REG_8__7_ );
nand NAND2_11252 ( P2_U7176 , P2_U5002 , P2_INSTQUEUE_REG_9__7_ );
nand NAND2_11253 ( P2_U7177 , P2_U4944 , P2_INSTQUEUE_REG_10__7_ );
nand NAND2_11254 ( P2_U7178 , P2_U4887 , P2_INSTQUEUE_REG_11__7_ );
nand NAND2_11255 ( P2_U7179 , P2_U4829 , P2_INSTQUEUE_REG_12__7_ );
nand NAND2_11256 ( P2_U7180 , P2_U4772 , P2_INSTQUEUE_REG_13__7_ );
nand NAND2_11257 ( P2_U7181 , P2_U4713 , P2_INSTQUEUE_REG_14__7_ );
nand NAND2_11258 ( P2_U7182 , P2_U4653 , P2_INSTQUEUE_REG_15__7_ );
nand NAND4_11259 ( P2_U7183 , P2_U4280 , P2_U4279 , P2_U4278 , P2_U4277 );
nand NAND2_11260 ( P2_U7184 , P2_U5517 , P2_INSTQUEUE_REG_0__6_ );
nand NAND2_11261 ( P2_U7185 , P2_U5460 , P2_INSTQUEUE_REG_1__6_ );
nand NAND2_11262 ( P2_U7186 , P2_U5402 , P2_INSTQUEUE_REG_2__6_ );
nand NAND2_11263 ( P2_U7187 , P2_U5345 , P2_INSTQUEUE_REG_3__6_ );
nand NAND2_11264 ( P2_U7188 , P2_U5287 , P2_INSTQUEUE_REG_4__6_ );
nand NAND2_11265 ( P2_U7189 , P2_U5230 , P2_INSTQUEUE_REG_5__6_ );
nand NAND2_11266 ( P2_U7190 , P2_U5172 , P2_INSTQUEUE_REG_6__6_ );
nand NAND2_11267 ( P2_U7191 , P2_U5116 , P2_INSTQUEUE_REG_7__6_ );
nand NAND2_11268 ( P2_U7192 , P2_U5059 , P2_INSTQUEUE_REG_8__6_ );
nand NAND2_11269 ( P2_U7193 , P2_U5002 , P2_INSTQUEUE_REG_9__6_ );
nand NAND2_11270 ( P2_U7194 , P2_U4944 , P2_INSTQUEUE_REG_10__6_ );
nand NAND2_11271 ( P2_U7195 , P2_U4887 , P2_INSTQUEUE_REG_11__6_ );
nand NAND2_11272 ( P2_U7196 , P2_U4829 , P2_INSTQUEUE_REG_12__6_ );
nand NAND2_11273 ( P2_U7197 , P2_U4772 , P2_INSTQUEUE_REG_13__6_ );
nand NAND2_11274 ( P2_U7198 , P2_U4713 , P2_INSTQUEUE_REG_14__6_ );
nand NAND2_11275 ( P2_U7199 , P2_U4653 , P2_INSTQUEUE_REG_15__6_ );
nand NAND4_11276 ( P2_U7200 , P2_U4284 , P2_U4283 , P2_U4282 , P2_U4281 );
nand NAND2_11277 ( P2_U7201 , P2_U2538 , P2_INSTQUEUE_REG_8__6_ );
nand NAND2_11278 ( P2_U7202 , P2_U2537 , P2_INSTQUEUE_REG_9__6_ );
nand NAND2_11279 ( P2_U7203 , P2_U2536 , P2_INSTQUEUE_REG_10__6_ );
nand NAND2_11280 ( P2_U7204 , P2_U2535 , P2_INSTQUEUE_REG_11__6_ );
nand NAND2_11281 ( P2_U7205 , P2_U2534 , P2_INSTQUEUE_REG_12__6_ );
nand NAND2_11282 ( P2_U7206 , P2_U2533 , P2_INSTQUEUE_REG_13__6_ );
nand NAND2_11283 ( P2_U7207 , P2_U2531 , P2_INSTQUEUE_REG_14__6_ );
nand NAND2_11284 ( P2_U7208 , P2_U2530 , P2_INSTQUEUE_REG_15__6_ );
nand NAND2_11285 ( P2_U7209 , P2_U2528 , P2_INSTQUEUE_REG_7__6_ );
nand NAND2_11286 ( P2_U7210 , P2_U2527 , P2_INSTQUEUE_REG_6__6_ );
nand NAND2_11287 ( P2_U7211 , P2_U2526 , P2_INSTQUEUE_REG_5__6_ );
nand NAND2_11288 ( P2_U7212 , P2_U2524 , P2_INSTQUEUE_REG_4__6_ );
nand NAND2_11289 ( P2_U7213 , P2_U2522 , P2_INSTQUEUE_REG_3__6_ );
nand NAND2_11290 ( P2_U7214 , P2_U2521 , P2_INSTQUEUE_REG_2__6_ );
nand NAND2_11291 ( P2_U7215 , P2_U2519 , P2_INSTQUEUE_REG_1__6_ );
nand NAND2_11292 ( P2_U7216 , P2_U2517 , P2_INSTQUEUE_REG_0__6_ );
nand NAND4_11293 ( P2_U7217 , P2_U4288 , P2_U4287 , P2_U4286 , P2_U4285 );
nand NAND2_11294 ( P2_U7218 , P2_U5517 , P2_INSTQUEUE_REG_0__5_ );
nand NAND2_11295 ( P2_U7219 , P2_U5460 , P2_INSTQUEUE_REG_1__5_ );
nand NAND2_11296 ( P2_U7220 , P2_U5402 , P2_INSTQUEUE_REG_2__5_ );
nand NAND2_11297 ( P2_U7221 , P2_U5345 , P2_INSTQUEUE_REG_3__5_ );
nand NAND2_11298 ( P2_U7222 , P2_U5287 , P2_INSTQUEUE_REG_4__5_ );
nand NAND2_11299 ( P2_U7223 , P2_U5230 , P2_INSTQUEUE_REG_5__5_ );
nand NAND2_11300 ( P2_U7224 , P2_U5172 , P2_INSTQUEUE_REG_6__5_ );
nand NAND2_11301 ( P2_U7225 , P2_U5116 , P2_INSTQUEUE_REG_7__5_ );
nand NAND2_11302 ( P2_U7226 , P2_U5059 , P2_INSTQUEUE_REG_8__5_ );
nand NAND2_11303 ( P2_U7227 , P2_U5002 , P2_INSTQUEUE_REG_9__5_ );
nand NAND2_11304 ( P2_U7228 , P2_U4944 , P2_INSTQUEUE_REG_10__5_ );
nand NAND2_11305 ( P2_U7229 , P2_U4887 , P2_INSTQUEUE_REG_11__5_ );
nand NAND2_11306 ( P2_U7230 , P2_U4829 , P2_INSTQUEUE_REG_12__5_ );
nand NAND2_11307 ( P2_U7231 , P2_U4772 , P2_INSTQUEUE_REG_13__5_ );
nand NAND2_11308 ( P2_U7232 , P2_U4713 , P2_INSTQUEUE_REG_14__5_ );
nand NAND2_11309 ( P2_U7233 , P2_U4653 , P2_INSTQUEUE_REG_15__5_ );
nand NAND4_11310 ( P2_U7234 , P2_U4292 , P2_U4291 , P2_U4290 , P2_U4289 );
nand NAND2_11311 ( P2_U7235 , P2_U2538 , P2_INSTQUEUE_REG_8__5_ );
nand NAND2_11312 ( P2_U7236 , P2_U2537 , P2_INSTQUEUE_REG_9__5_ );
nand NAND2_11313 ( P2_U7237 , P2_U2536 , P2_INSTQUEUE_REG_10__5_ );
nand NAND2_11314 ( P2_U7238 , P2_U2535 , P2_INSTQUEUE_REG_11__5_ );
nand NAND2_11315 ( P2_U7239 , P2_U2534 , P2_INSTQUEUE_REG_12__5_ );
nand NAND2_11316 ( P2_U7240 , P2_U2533 , P2_INSTQUEUE_REG_13__5_ );
nand NAND2_11317 ( P2_U7241 , P2_U2531 , P2_INSTQUEUE_REG_14__5_ );
nand NAND2_11318 ( P2_U7242 , P2_U2530 , P2_INSTQUEUE_REG_15__5_ );
nand NAND2_11319 ( P2_U7243 , P2_U2528 , P2_INSTQUEUE_REG_7__5_ );
nand NAND2_11320 ( P2_U7244 , P2_U2527 , P2_INSTQUEUE_REG_6__5_ );
nand NAND2_11321 ( P2_U7245 , P2_U2526 , P2_INSTQUEUE_REG_5__5_ );
nand NAND2_11322 ( P2_U7246 , P2_U2524 , P2_INSTQUEUE_REG_4__5_ );
nand NAND2_11323 ( P2_U7247 , P2_U2522 , P2_INSTQUEUE_REG_3__5_ );
nand NAND2_11324 ( P2_U7248 , P2_U2521 , P2_INSTQUEUE_REG_2__5_ );
nand NAND2_11325 ( P2_U7249 , P2_U2519 , P2_INSTQUEUE_REG_1__5_ );
nand NAND2_11326 ( P2_U7250 , P2_U2517 , P2_INSTQUEUE_REG_0__5_ );
nand NAND4_11327 ( P2_U7251 , P2_U4296 , P2_U4295 , P2_U4294 , P2_U4293 );
nand NAND2_11328 ( P2_U7252 , P2_U5517 , P2_INSTQUEUE_REG_0__4_ );
nand NAND2_11329 ( P2_U7253 , P2_U5460 , P2_INSTQUEUE_REG_1__4_ );
nand NAND2_11330 ( P2_U7254 , P2_U5402 , P2_INSTQUEUE_REG_2__4_ );
nand NAND2_11331 ( P2_U7255 , P2_U5345 , P2_INSTQUEUE_REG_3__4_ );
nand NAND2_11332 ( P2_U7256 , P2_U5287 , P2_INSTQUEUE_REG_4__4_ );
nand NAND2_11333 ( P2_U7257 , P2_U5230 , P2_INSTQUEUE_REG_5__4_ );
nand NAND2_11334 ( P2_U7258 , P2_U5172 , P2_INSTQUEUE_REG_6__4_ );
nand NAND2_11335 ( P2_U7259 , P2_U5116 , P2_INSTQUEUE_REG_7__4_ );
nand NAND2_11336 ( P2_U7260 , P2_U5059 , P2_INSTQUEUE_REG_8__4_ );
nand NAND2_11337 ( P2_U7261 , P2_U5002 , P2_INSTQUEUE_REG_9__4_ );
nand NAND2_11338 ( P2_U7262 , P2_U4944 , P2_INSTQUEUE_REG_10__4_ );
nand NAND2_11339 ( P2_U7263 , P2_U4887 , P2_INSTQUEUE_REG_11__4_ );
nand NAND2_11340 ( P2_U7264 , P2_U4829 , P2_INSTQUEUE_REG_12__4_ );
nand NAND2_11341 ( P2_U7265 , P2_U4772 , P2_INSTQUEUE_REG_13__4_ );
nand NAND2_11342 ( P2_U7266 , P2_U4713 , P2_INSTQUEUE_REG_14__4_ );
nand NAND2_11343 ( P2_U7267 , P2_U4653 , P2_INSTQUEUE_REG_15__4_ );
nand NAND4_11344 ( P2_U7268 , P2_U4300 , P2_U4299 , P2_U4298 , P2_U4297 );
nand NAND2_11345 ( P2_U7269 , P2_U2538 , P2_INSTQUEUE_REG_8__4_ );
nand NAND2_11346 ( P2_U7270 , P2_U2537 , P2_INSTQUEUE_REG_9__4_ );
nand NAND2_11347 ( P2_U7271 , P2_U2536 , P2_INSTQUEUE_REG_10__4_ );
nand NAND2_11348 ( P2_U7272 , P2_U2535 , P2_INSTQUEUE_REG_11__4_ );
nand NAND2_11349 ( P2_U7273 , P2_U2534 , P2_INSTQUEUE_REG_12__4_ );
nand NAND2_11350 ( P2_U7274 , P2_U2533 , P2_INSTQUEUE_REG_13__4_ );
nand NAND2_11351 ( P2_U7275 , P2_U2531 , P2_INSTQUEUE_REG_14__4_ );
nand NAND2_11352 ( P2_U7276 , P2_U2530 , P2_INSTQUEUE_REG_15__4_ );
nand NAND2_11353 ( P2_U7277 , P2_U2528 , P2_INSTQUEUE_REG_7__4_ );
nand NAND2_11354 ( P2_U7278 , P2_U2527 , P2_INSTQUEUE_REG_6__4_ );
nand NAND2_11355 ( P2_U7279 , P2_U2526 , P2_INSTQUEUE_REG_5__4_ );
nand NAND2_11356 ( P2_U7280 , P2_U2524 , P2_INSTQUEUE_REG_4__4_ );
nand NAND2_11357 ( P2_U7281 , P2_U2522 , P2_INSTQUEUE_REG_3__4_ );
nand NAND2_11358 ( P2_U7282 , P2_U2521 , P2_INSTQUEUE_REG_2__4_ );
nand NAND2_11359 ( P2_U7283 , P2_U2519 , P2_INSTQUEUE_REG_1__4_ );
nand NAND2_11360 ( P2_U7284 , P2_U2517 , P2_INSTQUEUE_REG_0__4_ );
nand NAND4_11361 ( P2_U7285 , P2_U4304 , P2_U4303 , P2_U4302 , P2_U4301 );
nand NAND2_11362 ( P2_U7286 , P2_U5517 , P2_INSTQUEUE_REG_0__3_ );
nand NAND2_11363 ( P2_U7287 , P2_U5460 , P2_INSTQUEUE_REG_1__3_ );
nand NAND2_11364 ( P2_U7288 , P2_U5402 , P2_INSTQUEUE_REG_2__3_ );
nand NAND2_11365 ( P2_U7289 , P2_U5345 , P2_INSTQUEUE_REG_3__3_ );
nand NAND2_11366 ( P2_U7290 , P2_U5287 , P2_INSTQUEUE_REG_4__3_ );
nand NAND2_11367 ( P2_U7291 , P2_U5230 , P2_INSTQUEUE_REG_5__3_ );
nand NAND2_11368 ( P2_U7292 , P2_U5172 , P2_INSTQUEUE_REG_6__3_ );
nand NAND2_11369 ( P2_U7293 , P2_U5116 , P2_INSTQUEUE_REG_7__3_ );
nand NAND2_11370 ( P2_U7294 , P2_U5059 , P2_INSTQUEUE_REG_8__3_ );
nand NAND2_11371 ( P2_U7295 , P2_U5002 , P2_INSTQUEUE_REG_9__3_ );
nand NAND2_11372 ( P2_U7296 , P2_U4944 , P2_INSTQUEUE_REG_10__3_ );
nand NAND2_11373 ( P2_U7297 , P2_U4887 , P2_INSTQUEUE_REG_11__3_ );
nand NAND2_11374 ( P2_U7298 , P2_U4829 , P2_INSTQUEUE_REG_12__3_ );
nand NAND2_11375 ( P2_U7299 , P2_U4772 , P2_INSTQUEUE_REG_13__3_ );
nand NAND2_11376 ( P2_U7300 , P2_U4713 , P2_INSTQUEUE_REG_14__3_ );
nand NAND2_11377 ( P2_U7301 , P2_U4653 , P2_INSTQUEUE_REG_15__3_ );
nand NAND4_11378 ( P2_U7302 , P2_U4308 , P2_U4307 , P2_U4306 , P2_U4305 );
nand NAND2_11379 ( P2_U7303 , P2_U2538 , P2_INSTQUEUE_REG_8__3_ );
nand NAND2_11380 ( P2_U7304 , P2_U2537 , P2_INSTQUEUE_REG_9__3_ );
nand NAND2_11381 ( P2_U7305 , P2_U2536 , P2_INSTQUEUE_REG_10__3_ );
nand NAND2_11382 ( P2_U7306 , P2_U2535 , P2_INSTQUEUE_REG_11__3_ );
nand NAND2_11383 ( P2_U7307 , P2_U2534 , P2_INSTQUEUE_REG_12__3_ );
nand NAND2_11384 ( P2_U7308 , P2_U2533 , P2_INSTQUEUE_REG_13__3_ );
nand NAND2_11385 ( P2_U7309 , P2_U2531 , P2_INSTQUEUE_REG_14__3_ );
nand NAND2_11386 ( P2_U7310 , P2_U2530 , P2_INSTQUEUE_REG_15__3_ );
nand NAND2_11387 ( P2_U7311 , P2_U2528 , P2_INSTQUEUE_REG_7__3_ );
nand NAND2_11388 ( P2_U7312 , P2_U2527 , P2_INSTQUEUE_REG_6__3_ );
nand NAND2_11389 ( P2_U7313 , P2_U2526 , P2_INSTQUEUE_REG_5__3_ );
nand NAND2_11390 ( P2_U7314 , P2_U2524 , P2_INSTQUEUE_REG_4__3_ );
nand NAND2_11391 ( P2_U7315 , P2_U2522 , P2_INSTQUEUE_REG_3__3_ );
nand NAND2_11392 ( P2_U7316 , P2_U2521 , P2_INSTQUEUE_REG_2__3_ );
nand NAND2_11393 ( P2_U7317 , P2_U2519 , P2_INSTQUEUE_REG_1__3_ );
nand NAND2_11394 ( P2_U7318 , P2_U2517 , P2_INSTQUEUE_REG_0__3_ );
nand NAND4_11395 ( P2_U7319 , P2_U4312 , P2_U4311 , P2_U4310 , P2_U4309 );
nand NAND2_11396 ( P2_U7320 , P2_U5517 , P2_INSTQUEUE_REG_0__2_ );
nand NAND2_11397 ( P2_U7321 , P2_U5460 , P2_INSTQUEUE_REG_1__2_ );
nand NAND2_11398 ( P2_U7322 , P2_U5402 , P2_INSTQUEUE_REG_2__2_ );
nand NAND2_11399 ( P2_U7323 , P2_U5345 , P2_INSTQUEUE_REG_3__2_ );
nand NAND2_11400 ( P2_U7324 , P2_U5287 , P2_INSTQUEUE_REG_4__2_ );
nand NAND2_11401 ( P2_U7325 , P2_U5230 , P2_INSTQUEUE_REG_5__2_ );
nand NAND2_11402 ( P2_U7326 , P2_U5172 , P2_INSTQUEUE_REG_6__2_ );
nand NAND2_11403 ( P2_U7327 , P2_U5116 , P2_INSTQUEUE_REG_7__2_ );
nand NAND2_11404 ( P2_U7328 , P2_U5059 , P2_INSTQUEUE_REG_8__2_ );
nand NAND2_11405 ( P2_U7329 , P2_U5002 , P2_INSTQUEUE_REG_9__2_ );
nand NAND2_11406 ( P2_U7330 , P2_U4944 , P2_INSTQUEUE_REG_10__2_ );
nand NAND2_11407 ( P2_U7331 , P2_U4887 , P2_INSTQUEUE_REG_11__2_ );
nand NAND2_11408 ( P2_U7332 , P2_U4829 , P2_INSTQUEUE_REG_12__2_ );
nand NAND2_11409 ( P2_U7333 , P2_U4772 , P2_INSTQUEUE_REG_13__2_ );
nand NAND2_11410 ( P2_U7334 , P2_U4713 , P2_INSTQUEUE_REG_14__2_ );
nand NAND2_11411 ( P2_U7335 , P2_U4653 , P2_INSTQUEUE_REG_15__2_ );
nand NAND4_11412 ( P2_U7336 , P2_U4316 , P2_U4315 , P2_U4314 , P2_U4313 );
nand NAND2_11413 ( P2_U7337 , P2_U2538 , P2_INSTQUEUE_REG_8__2_ );
nand NAND2_11414 ( P2_U7338 , P2_U2537 , P2_INSTQUEUE_REG_9__2_ );
nand NAND2_11415 ( P2_U7339 , P2_U2536 , P2_INSTQUEUE_REG_10__2_ );
nand NAND2_11416 ( P2_U7340 , P2_U2535 , P2_INSTQUEUE_REG_11__2_ );
nand NAND2_11417 ( P2_U7341 , P2_U2534 , P2_INSTQUEUE_REG_12__2_ );
nand NAND2_11418 ( P2_U7342 , P2_U2533 , P2_INSTQUEUE_REG_13__2_ );
nand NAND2_11419 ( P2_U7343 , P2_U2531 , P2_INSTQUEUE_REG_14__2_ );
nand NAND2_11420 ( P2_U7344 , P2_U2530 , P2_INSTQUEUE_REG_15__2_ );
nand NAND2_11421 ( P2_U7345 , P2_U2528 , P2_INSTQUEUE_REG_7__2_ );
nand NAND2_11422 ( P2_U7346 , P2_U2527 , P2_INSTQUEUE_REG_6__2_ );
nand NAND2_11423 ( P2_U7347 , P2_U2526 , P2_INSTQUEUE_REG_5__2_ );
nand NAND2_11424 ( P2_U7348 , P2_U2524 , P2_INSTQUEUE_REG_4__2_ );
nand NAND2_11425 ( P2_U7349 , P2_U2522 , P2_INSTQUEUE_REG_3__2_ );
nand NAND2_11426 ( P2_U7350 , P2_U2521 , P2_INSTQUEUE_REG_2__2_ );
nand NAND2_11427 ( P2_U7351 , P2_U2519 , P2_INSTQUEUE_REG_1__2_ );
nand NAND2_11428 ( P2_U7352 , P2_U2517 , P2_INSTQUEUE_REG_0__2_ );
nand NAND4_11429 ( P2_U7353 , P2_U4320 , P2_U4319 , P2_U4318 , P2_U4317 );
nand NAND2_11430 ( P2_U7354 , P2_U5517 , P2_INSTQUEUE_REG_0__1_ );
nand NAND2_11431 ( P2_U7355 , P2_U5460 , P2_INSTQUEUE_REG_1__1_ );
nand NAND2_11432 ( P2_U7356 , P2_U5402 , P2_INSTQUEUE_REG_2__1_ );
nand NAND2_11433 ( P2_U7357 , P2_U5345 , P2_INSTQUEUE_REG_3__1_ );
nand NAND2_11434 ( P2_U7358 , P2_U5287 , P2_INSTQUEUE_REG_4__1_ );
nand NAND2_11435 ( P2_U7359 , P2_U5230 , P2_INSTQUEUE_REG_5__1_ );
nand NAND2_11436 ( P2_U7360 , P2_U5172 , P2_INSTQUEUE_REG_6__1_ );
nand NAND2_11437 ( P2_U7361 , P2_U5116 , P2_INSTQUEUE_REG_7__1_ );
nand NAND2_11438 ( P2_U7362 , P2_U5059 , P2_INSTQUEUE_REG_8__1_ );
nand NAND2_11439 ( P2_U7363 , P2_U5002 , P2_INSTQUEUE_REG_9__1_ );
nand NAND2_11440 ( P2_U7364 , P2_U4944 , P2_INSTQUEUE_REG_10__1_ );
nand NAND2_11441 ( P2_U7365 , P2_U4887 , P2_INSTQUEUE_REG_11__1_ );
nand NAND2_11442 ( P2_U7366 , P2_U4829 , P2_INSTQUEUE_REG_12__1_ );
nand NAND2_11443 ( P2_U7367 , P2_U4772 , P2_INSTQUEUE_REG_13__1_ );
nand NAND2_11444 ( P2_U7368 , P2_U4713 , P2_INSTQUEUE_REG_14__1_ );
nand NAND2_11445 ( P2_U7369 , P2_U4653 , P2_INSTQUEUE_REG_15__1_ );
nand NAND4_11446 ( P2_U7370 , P2_U4324 , P2_U4323 , P2_U4322 , P2_U4321 );
nand NAND2_11447 ( P2_U7371 , P2_U2538 , P2_INSTQUEUE_REG_8__1_ );
nand NAND2_11448 ( P2_U7372 , P2_U2537 , P2_INSTQUEUE_REG_9__1_ );
nand NAND2_11449 ( P2_U7373 , P2_U2536 , P2_INSTQUEUE_REG_10__1_ );
nand NAND2_11450 ( P2_U7374 , P2_U2535 , P2_INSTQUEUE_REG_11__1_ );
nand NAND2_11451 ( P2_U7375 , P2_U2534 , P2_INSTQUEUE_REG_12__1_ );
nand NAND2_11452 ( P2_U7376 , P2_U2533 , P2_INSTQUEUE_REG_13__1_ );
nand NAND2_11453 ( P2_U7377 , P2_U2531 , P2_INSTQUEUE_REG_14__1_ );
nand NAND2_11454 ( P2_U7378 , P2_U2530 , P2_INSTQUEUE_REG_15__1_ );
nand NAND2_11455 ( P2_U7379 , P2_U2528 , P2_INSTQUEUE_REG_7__1_ );
nand NAND2_11456 ( P2_U7380 , P2_U2527 , P2_INSTQUEUE_REG_6__1_ );
nand NAND2_11457 ( P2_U7381 , P2_U2526 , P2_INSTQUEUE_REG_5__1_ );
nand NAND2_11458 ( P2_U7382 , P2_U2524 , P2_INSTQUEUE_REG_4__1_ );
nand NAND2_11459 ( P2_U7383 , P2_U2522 , P2_INSTQUEUE_REG_3__1_ );
nand NAND2_11460 ( P2_U7384 , P2_U2521 , P2_INSTQUEUE_REG_2__1_ );
nand NAND2_11461 ( P2_U7385 , P2_U2519 , P2_INSTQUEUE_REG_1__1_ );
nand NAND2_11462 ( P2_U7386 , P2_U2517 , P2_INSTQUEUE_REG_0__1_ );
nand NAND4_11463 ( P2_U7387 , P2_U4328 , P2_U4327 , P2_U4326 , P2_U4325 );
nand NAND2_11464 ( P2_U7388 , P2_U5517 , P2_INSTQUEUE_REG_0__0_ );
nand NAND2_11465 ( P2_U7389 , P2_U5460 , P2_INSTQUEUE_REG_1__0_ );
nand NAND2_11466 ( P2_U7390 , P2_U5402 , P2_INSTQUEUE_REG_2__0_ );
nand NAND2_11467 ( P2_U7391 , P2_U5345 , P2_INSTQUEUE_REG_3__0_ );
nand NAND2_11468 ( P2_U7392 , P2_U5287 , P2_INSTQUEUE_REG_4__0_ );
nand NAND2_11469 ( P2_U7393 , P2_U5230 , P2_INSTQUEUE_REG_5__0_ );
nand NAND2_11470 ( P2_U7394 , P2_U5172 , P2_INSTQUEUE_REG_6__0_ );
nand NAND2_11471 ( P2_U7395 , P2_U5116 , P2_INSTQUEUE_REG_7__0_ );
nand NAND2_11472 ( P2_U7396 , P2_U5059 , P2_INSTQUEUE_REG_8__0_ );
nand NAND2_11473 ( P2_U7397 , P2_U5002 , P2_INSTQUEUE_REG_9__0_ );
nand NAND2_11474 ( P2_U7398 , P2_U4944 , P2_INSTQUEUE_REG_10__0_ );
nand NAND2_11475 ( P2_U7399 , P2_U4887 , P2_INSTQUEUE_REG_11__0_ );
nand NAND2_11476 ( P2_U7400 , P2_U4829 , P2_INSTQUEUE_REG_12__0_ );
nand NAND2_11477 ( P2_U7401 , P2_U4772 , P2_INSTQUEUE_REG_13__0_ );
nand NAND2_11478 ( P2_U7402 , P2_U4713 , P2_INSTQUEUE_REG_14__0_ );
nand NAND2_11479 ( P2_U7403 , P2_U4653 , P2_INSTQUEUE_REG_15__0_ );
nand NAND4_11480 ( P2_U7404 , P2_U4332 , P2_U4331 , P2_U4330 , P2_U4329 );
nand NAND2_11481 ( P2_U7405 , P2_U2538 , P2_INSTQUEUE_REG_8__0_ );
nand NAND2_11482 ( P2_U7406 , P2_U2537 , P2_INSTQUEUE_REG_9__0_ );
nand NAND2_11483 ( P2_U7407 , P2_U2536 , P2_INSTQUEUE_REG_10__0_ );
nand NAND2_11484 ( P2_U7408 , P2_U2535 , P2_INSTQUEUE_REG_11__0_ );
nand NAND2_11485 ( P2_U7409 , P2_U2534 , P2_INSTQUEUE_REG_12__0_ );
nand NAND2_11486 ( P2_U7410 , P2_U2533 , P2_INSTQUEUE_REG_13__0_ );
nand NAND2_11487 ( P2_U7411 , P2_U2531 , P2_INSTQUEUE_REG_14__0_ );
nand NAND2_11488 ( P2_U7412 , P2_U2530 , P2_INSTQUEUE_REG_15__0_ );
nand NAND2_11489 ( P2_U7413 , P2_U2528 , P2_INSTQUEUE_REG_7__0_ );
nand NAND2_11490 ( P2_U7414 , P2_U2527 , P2_INSTQUEUE_REG_6__0_ );
nand NAND2_11491 ( P2_U7415 , P2_U2526 , P2_INSTQUEUE_REG_5__0_ );
nand NAND2_11492 ( P2_U7416 , P2_U2524 , P2_INSTQUEUE_REG_4__0_ );
nand NAND2_11493 ( P2_U7417 , P2_U2522 , P2_INSTQUEUE_REG_3__0_ );
nand NAND2_11494 ( P2_U7418 , P2_U2521 , P2_INSTQUEUE_REG_2__0_ );
nand NAND2_11495 ( P2_U7419 , P2_U2519 , P2_INSTQUEUE_REG_1__0_ );
nand NAND2_11496 ( P2_U7420 , P2_U2517 , P2_INSTQUEUE_REG_0__0_ );
nand NAND4_11497 ( P2_U7421 , P2_U4336 , P2_U4335 , P2_U4334 , P2_U4333 );
nand NAND2_11498 ( P2_U7422 , P2_U2352 , P2_U7319 );
nand NAND2_11499 ( P2_U7423 , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_STATE2_REG_3_ );
nand NAND2_11500 ( P2_U7424 , P2_U2352 , P2_U7353 );
nand NAND2_11501 ( P2_U7425 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_STATE2_REG_3_ );
nand NAND2_11502 ( P2_U7426 , P2_U2439 , P2_U3295 );
nand NAND2_11503 ( P2_U7427 , P2_U2352 , P2_U7387 );
nand NAND2_11504 ( P2_U7428 , P2_INSTQUEUEWR_ADDR_REG_1_ , P2_STATE2_REG_3_ );
nand NAND2_11505 ( P2_U7429 , P2_U2352 , P2_U7421 );
nand NAND2_11506 ( P2_U7430 , P2_INSTQUEUEWR_ADDR_REG_0_ , P2_STATE2_REG_3_ );
nand NAND2_11507 ( P2_U7431 , P2_U2439 , P2_U3279 );
nand NAND3_11508 ( P2_U7432 , P2_U4414 , P2_U7431 , P2_U4413 );
nand NAND2_11509 ( P2_U7433 , P2_INSTADDRPOINTER_REG_9_ , P2_U7432 );
nand NAND2_11510 ( P2_U7434 , P2_U2353 , P2_REIP_REG_9_ );
nand NAND2_11511 ( P2_U7435 , P2_U4412 , P2_EAX_REG_9_ );
nand NAND2_11512 ( P2_U7436 , P2_U2352 , P2_U2608 );
nand NAND2_11513 ( P2_U7437 , P2_INSTADDRPOINTER_REG_8_ , P2_U7432 );
nand NAND2_11514 ( P2_U7438 , P2_U2353 , P2_REIP_REG_8_ );
nand NAND2_11515 ( P2_U7439 , P2_U4412 , P2_EAX_REG_8_ );
nand NAND2_11516 ( P2_U7440 , P2_U2352 , P2_U2607 );
nand NAND2_11517 ( P2_U7441 , P2_INSTADDRPOINTER_REG_7_ , P2_U7432 );
nand NAND2_11518 ( P2_U7442 , P2_U2353 , P2_REIP_REG_7_ );
nand NAND2_11519 ( P2_U7443 , P2_U4412 , P2_EAX_REG_7_ );
nand NAND2_11520 ( P2_U7444 , P2_INSTADDRPOINTER_REG_6_ , P2_U7432 );
nand NAND2_11521 ( P2_U7445 , P2_U2353 , P2_REIP_REG_6_ );
nand NAND2_11522 ( P2_U7446 , P2_U4412 , P2_EAX_REG_6_ );
nand NAND2_11523 ( P2_U7447 , P2_INSTADDRPOINTER_REG_5_ , P2_U7432 );
nand NAND2_11524 ( P2_U7448 , P2_U2353 , P2_REIP_REG_5_ );
nand NAND2_11525 ( P2_U7449 , P2_U4412 , P2_EAX_REG_5_ );
nand NAND2_11526 ( P2_U7450 , P2_INSTADDRPOINTER_REG_4_ , P2_U7432 );
nand NAND2_11527 ( P2_U7451 , P2_U2353 , P2_REIP_REG_4_ );
nand NAND2_11528 ( P2_U7452 , P2_U4412 , P2_EAX_REG_4_ );
nand NAND2_11529 ( P2_U7453 , P2_INSTADDRPOINTER_REG_31_ , P2_U7432 );
nand NAND2_11530 ( P2_U7454 , P2_U2353 , P2_REIP_REG_31_ );
nand NAND2_11531 ( P2_U7455 , P2_U4412 , P2_EAX_REG_31_ );
nand NAND2_11532 ( P2_U7456 , P2_INSTADDRPOINTER_REG_30_ , P2_U7432 );
nand NAND2_11533 ( P2_U7457 , P2_U2353 , P2_REIP_REG_30_ );
nand NAND2_11534 ( P2_U7458 , P2_U4412 , P2_EAX_REG_30_ );
nand NAND2_11535 ( P2_U7459 , P2_INSTADDRPOINTER_REG_3_ , P2_U7432 );
nand NAND2_11536 ( P2_U7460 , P2_U2353 , P2_REIP_REG_3_ );
nand NAND2_11537 ( P2_U7461 , P2_U4412 , P2_EAX_REG_3_ );
nand NAND2_11538 ( P2_U7462 , P2_INSTADDRPOINTER_REG_29_ , P2_U7432 );
nand NAND2_11539 ( P2_U7463 , P2_U2353 , P2_REIP_REG_29_ );
nand NAND2_11540 ( P2_U7464 , P2_U4412 , P2_EAX_REG_29_ );
nand NAND2_11541 ( P2_U7465 , P2_INSTADDRPOINTER_REG_28_ , P2_U7432 );
nand NAND2_11542 ( P2_U7466 , P2_U2353 , P2_REIP_REG_28_ );
nand NAND2_11543 ( P2_U7467 , P2_U4412 , P2_EAX_REG_28_ );
nand NAND2_11544 ( P2_U7468 , P2_INSTADDRPOINTER_REG_27_ , P2_U7432 );
nand NAND2_11545 ( P2_U7469 , P2_U2353 , P2_REIP_REG_27_ );
nand NAND2_11546 ( P2_U7470 , P2_U4412 , P2_EAX_REG_27_ );
nand NAND2_11547 ( P2_U7471 , P2_INSTADDRPOINTER_REG_26_ , P2_U7432 );
nand NAND2_11548 ( P2_U7472 , P2_U2353 , P2_REIP_REG_26_ );
nand NAND2_11549 ( P2_U7473 , P2_U4412 , P2_EAX_REG_26_ );
nand NAND2_11550 ( P2_U7474 , P2_INSTADDRPOINTER_REG_25_ , P2_U7432 );
nand NAND2_11551 ( P2_U7475 , P2_U2353 , P2_REIP_REG_25_ );
nand NAND2_11552 ( P2_U7476 , P2_U4412 , P2_EAX_REG_25_ );
nand NAND2_11553 ( P2_U7477 , P2_INSTADDRPOINTER_REG_24_ , P2_U7432 );
nand NAND2_11554 ( P2_U7478 , P2_U2353 , P2_REIP_REG_24_ );
nand NAND2_11555 ( P2_U7479 , P2_U4412 , P2_EAX_REG_24_ );
nand NAND2_11556 ( P2_U7480 , P2_INSTADDRPOINTER_REG_23_ , P2_U7432 );
nand NAND2_11557 ( P2_U7481 , P2_U2353 , P2_REIP_REG_23_ );
nand NAND2_11558 ( P2_U7482 , P2_U4412 , P2_EAX_REG_23_ );
nand NAND2_11559 ( P2_U7483 , P2_INSTADDRPOINTER_REG_22_ , P2_U7432 );
nand NAND2_11560 ( P2_U7484 , P2_U2353 , P2_REIP_REG_22_ );
nand NAND2_11561 ( P2_U7485 , P2_U4412 , P2_EAX_REG_22_ );
nand NAND2_11562 ( P2_U7486 , P2_INSTADDRPOINTER_REG_21_ , P2_U7432 );
nand NAND2_11563 ( P2_U7487 , P2_U2353 , P2_REIP_REG_21_ );
nand NAND2_11564 ( P2_U7488 , P2_U4412 , P2_EAX_REG_21_ );
nand NAND2_11565 ( P2_U7489 , P2_INSTADDRPOINTER_REG_20_ , P2_U7432 );
nand NAND2_11566 ( P2_U7490 , P2_U2353 , P2_REIP_REG_20_ );
nand NAND2_11567 ( P2_U7491 , P2_U4412 , P2_EAX_REG_20_ );
nand NAND2_11568 ( P2_U7492 , P2_INSTADDRPOINTER_REG_2_ , P2_U7432 );
nand NAND2_11569 ( P2_U7493 , P2_U2353 , P2_REIP_REG_2_ );
nand NAND2_11570 ( P2_U7494 , P2_U4412 , P2_EAX_REG_2_ );
nand NAND2_11571 ( P2_U7495 , P2_INSTADDRPOINTER_REG_19_ , P2_U7432 );
nand NAND2_11572 ( P2_U7496 , P2_U2353 , P2_REIP_REG_19_ );
nand NAND2_11573 ( P2_U7497 , P2_U4412 , P2_EAX_REG_19_ );
nand NAND2_11574 ( P2_U7498 , P2_INSTADDRPOINTER_REG_18_ , P2_U7432 );
nand NAND2_11575 ( P2_U7499 , P2_U2353 , P2_REIP_REG_18_ );
nand NAND2_11576 ( P2_U7500 , P2_U4412 , P2_EAX_REG_18_ );
nand NAND2_11577 ( P2_U7501 , P2_INSTADDRPOINTER_REG_17_ , P2_U7432 );
nand NAND2_11578 ( P2_U7502 , P2_U2353 , P2_REIP_REG_17_ );
nand NAND2_11579 ( P2_U7503 , P2_U4412 , P2_EAX_REG_17_ );
nand NAND2_11580 ( P2_U7504 , P2_INSTADDRPOINTER_REG_16_ , P2_U7432 );
nand NAND2_11581 ( P2_U7505 , P2_U2353 , P2_REIP_REG_16_ );
nand NAND2_11582 ( P2_U7506 , P2_U4412 , P2_EAX_REG_16_ );
nand NAND2_11583 ( P2_U7507 , P2_INSTADDRPOINTER_REG_15_ , P2_U7432 );
nand NAND2_11584 ( P2_U7508 , P2_U2353 , P2_REIP_REG_15_ );
nand NAND2_11585 ( P2_U7509 , P2_U4412 , P2_EAX_REG_15_ );
nand NAND2_11586 ( P2_U7510 , P2_U2352 , P2_U2614 );
nand NAND2_11587 ( P2_U7511 , P2_INSTADDRPOINTER_REG_14_ , P2_U7432 );
nand NAND2_11588 ( P2_U7512 , P2_U2353 , P2_REIP_REG_14_ );
nand NAND2_11589 ( P2_U7513 , P2_U4412 , P2_EAX_REG_14_ );
nand NAND2_11590 ( P2_U7514 , P2_U2352 , P2_U2613 );
nand NAND2_11591 ( P2_U7515 , P2_INSTADDRPOINTER_REG_13_ , P2_U7432 );
nand NAND2_11592 ( P2_U7516 , P2_U2353 , P2_REIP_REG_13_ );
nand NAND2_11593 ( P2_U7517 , P2_U4412 , P2_EAX_REG_13_ );
nand NAND2_11594 ( P2_U7518 , P2_U2352 , P2_U2612 );
nand NAND2_11595 ( P2_U7519 , P2_INSTADDRPOINTER_REG_12_ , P2_U7432 );
nand NAND2_11596 ( P2_U7520 , P2_U2353 , P2_REIP_REG_12_ );
nand NAND2_11597 ( P2_U7521 , P2_U4412 , P2_EAX_REG_12_ );
nand NAND2_11598 ( P2_U7522 , P2_U2352 , P2_U2611 );
nand NAND2_11599 ( P2_U7523 , P2_INSTADDRPOINTER_REG_11_ , P2_U7432 );
nand NAND2_11600 ( P2_U7524 , P2_U2353 , P2_REIP_REG_11_ );
nand NAND2_11601 ( P2_U7525 , P2_U4412 , P2_EAX_REG_11_ );
nand NAND2_11602 ( P2_U7526 , P2_U2352 , P2_U2610 );
nand NAND2_11603 ( P2_U7527 , P2_INSTADDRPOINTER_REG_10_ , P2_U7432 );
nand NAND2_11604 ( P2_U7528 , P2_U2353 , P2_REIP_REG_10_ );
nand NAND2_11605 ( P2_U7529 , P2_U4412 , P2_EAX_REG_10_ );
nand NAND2_11606 ( P2_U7530 , P2_U2352 , P2_U2609 );
nand NAND2_11607 ( P2_U7531 , P2_INSTADDRPOINTER_REG_1_ , P2_U7432 );
nand NAND2_11608 ( P2_U7532 , P2_U2353 , P2_REIP_REG_1_ );
nand NAND2_11609 ( P2_U7533 , P2_U4412 , P2_EAX_REG_1_ );
nand NAND2_11610 ( P2_U7534 , P2_INSTADDRPOINTER_REG_0_ , P2_U7432 );
nand NAND2_11611 ( P2_U7535 , P2_U2353 , P2_REIP_REG_0_ );
nand NAND2_11612 ( P2_U7536 , P2_U4412 , P2_EAX_REG_0_ );
nand NAND2_11613 ( P2_U7537 , P2_EBX_REG_9_ , P2_U7869 );
nand NAND2_11614 ( P2_U7538 , P2_EBX_REG_8_ , P2_U7869 );
nand NAND2_11615 ( P2_U7539 , P2_EBX_REG_31_ , P2_U7869 );
nand NAND2_11616 ( P2_U7540 , P2_EBX_REG_30_ , P2_U7869 );
nand NAND2_11617 ( P2_U7541 , P2_EBX_REG_29_ , P2_U7869 );
nand NAND2_11618 ( P2_U7542 , P2_EBX_REG_28_ , P2_U7869 );
nand NAND2_11619 ( P2_U7543 , P2_EBX_REG_27_ , P2_U7869 );
nand NAND2_11620 ( P2_U7544 , P2_EBX_REG_26_ , P2_U7869 );
nand NAND2_11621 ( P2_U7545 , P2_EBX_REG_25_ , P2_U7869 );
nand NAND2_11622 ( P2_U7546 , P2_EBX_REG_24_ , P2_U7869 );
nand NAND2_11623 ( P2_U7547 , P2_EBX_REG_23_ , P2_U7869 );
nand NAND2_11624 ( P2_U7548 , P2_EBX_REG_22_ , P2_U7869 );
nand NAND2_11625 ( P2_U7549 , P2_EBX_REG_21_ , P2_U7869 );
nand NAND2_11626 ( P2_U7550 , P2_EBX_REG_20_ , P2_U7869 );
nand NAND2_11627 ( P2_U7551 , P2_EBX_REG_19_ , P2_U7869 );
nand NAND2_11628 ( P2_U7552 , P2_EBX_REG_18_ , P2_U7869 );
nand NAND2_11629 ( P2_U7553 , P2_EBX_REG_17_ , P2_U7869 );
nand NAND2_11630 ( P2_U7554 , P2_EBX_REG_16_ , P2_U7869 );
nand NAND2_11631 ( P2_U7555 , P2_EBX_REG_15_ , P2_U7869 );
nand NAND2_11632 ( P2_U7556 , P2_EBX_REG_14_ , P2_U7869 );
nand NAND2_11633 ( P2_U7557 , P2_EBX_REG_13_ , P2_U7869 );
nand NAND2_11634 ( P2_U7558 , P2_EBX_REG_12_ , P2_U7869 );
nand NAND2_11635 ( P2_U7559 , P2_EBX_REG_11_ , P2_U7869 );
nand NAND2_11636 ( P2_U7560 , P2_EBX_REG_10_ , P2_U7869 );
nand NAND2_11637 ( P2_U7561 , P2_U4596 , P2_U3294 );
nand NAND2_11638 ( P2_U7562 , P2_U4428 , P2_U7285 );
nand NAND2_11639 ( P2_U7563 , P2_INSTQUEUERD_ADDR_REG_4_ , P2_U7561 );
nand NAND2_11640 ( P2_U7564 , P2_U4428 , P2_U7319 );
nand NAND2_11641 ( P2_U7565 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U7561 );
nand NAND2_11642 ( P2_U7566 , P2_U4428 , P2_U7353 );
nand NAND2_11643 ( P2_U7567 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_U7561 );
nand NAND2_11644 ( P2_U7568 , P2_U4428 , P2_U7387 );
nand NAND2_11645 ( P2_U7569 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_U7561 );
nand NAND2_11646 ( P2_U7570 , P2_U4428 , P2_U7421 );
nand NAND2_11647 ( P2_U7571 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_U7561 );
nand NAND2_11648 ( P2_U7572 , P2_INSTQUEUEWR_ADDR_REG_4_ , P2_U7561 );
nand NAND2_11649 ( P2_U7573 , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_U7561 );
nand NAND2_11650 ( P2_U7574 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_U7561 );
nand NAND2_11651 ( P2_U7575 , P2_INSTQUEUEWR_ADDR_REG_1_ , P2_U7561 );
nand NAND2_11652 ( P2_U7576 , P2_INSTQUEUEWR_ADDR_REG_0_ , P2_U7561 );
nand NAND2_11653 ( P2_U7577 , P2_U4377 , P2_U5572 );
nand NAND2_11654 ( P2_U7578 , P2_STATE2_REG_0_ , P2_U4432 );
nand NAND2_11655 ( P2_U7579 , P2_U2617 , P2_U2450 );
nand NAND2_11656 ( P2_U7580 , P2_U4376 , P2_U5592 );
nand NAND3_11657 ( P2_U7581 , P2_U3525 , P2_U6845 , P2_U7867 );
nand NAND2_11658 ( P2_U7582 , P2_U4471 , P2_INSTQUEUEWR_ADDR_REG_3_ );
nand NAND2_11659 ( P2_U7583 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U7890 );
nand NAND2_11660 ( P2_U7584 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_U7890 );
nand NAND2_11661 ( P2_U7585 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_U3284 );
nand NAND2_11662 ( P2_U7586 , P2_U4381 , P2_U4424 );
nand NAND2_11663 ( P2_U7587 , P2_U4471 , P2_INSTQUEUEWR_ADDR_REG_1_ );
nand NAND2_11664 ( P2_U7588 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_U7890 );
nand NAND2_11665 ( P2_U7589 , P2_U2590 , P2_U6845 );
nand NAND2_11666 ( P2_U7590 , P2_U4471 , P2_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND3_11667 ( P2_U7591 , P2_U2376 , P2_U7871 , P2_U4416 );
nand NAND4_11668 ( P2_U7592 , P2_U7591 , P2_U3285 , P2_U4422 , P2_U3539 );
nand NAND2_11669 ( P2_U7593 , P2_INSTADDRPOINTER_REG_9_ , P2_U7592 );
nand NAND2_11670 ( P2_U7594 , P2_PHYADDRPOINTER_REG_9_ , P2_STATE2_REG_1_ );
nand NAND2_11671 ( P2_U7595 , P2_U4423 , P2_REIP_REG_9_ );
nand NAND2_11672 ( P2_U7596 , P2_U2358 , P2_EBX_REG_9_ );
nand NAND2_11673 ( P2_U7597 , P2_INSTADDRPOINTER_REG_8_ , P2_U7592 );
nand NAND2_11674 ( P2_U7598 , P2_PHYADDRPOINTER_REG_8_ , P2_STATE2_REG_1_ );
nand NAND2_11675 ( P2_U7599 , P2_U4423 , P2_REIP_REG_8_ );
nand NAND2_11676 ( P2_U7600 , P2_U2358 , P2_EBX_REG_8_ );
nand NAND2_11677 ( P2_U7601 , P2_INSTADDRPOINTER_REG_7_ , P2_U7592 );
nand NAND2_11678 ( P2_U7602 , P2_PHYADDRPOINTER_REG_7_ , P2_STATE2_REG_1_ );
nand NAND2_11679 ( P2_U7603 , P2_U4423 , P2_REIP_REG_7_ );
nand NAND2_11680 ( P2_U7604 , P2_U2358 , P2_EBX_REG_7_ );
nand NAND2_11681 ( P2_U7605 , P2_INSTADDRPOINTER_REG_6_ , P2_U7592 );
nand NAND2_11682 ( P2_U7606 , P2_PHYADDRPOINTER_REG_6_ , P2_STATE2_REG_1_ );
nand NAND2_11683 ( P2_U7607 , P2_U4423 , P2_REIP_REG_6_ );
nand NAND2_11684 ( P2_U7608 , P2_U2358 , P2_EBX_REG_6_ );
nand NAND2_11685 ( P2_U7609 , P2_INSTADDRPOINTER_REG_5_ , P2_U7592 );
nand NAND2_11686 ( P2_U7610 , P2_PHYADDRPOINTER_REG_5_ , P2_STATE2_REG_1_ );
nand NAND2_11687 ( P2_U7611 , P2_U4423 , P2_REIP_REG_5_ );
nand NAND2_11688 ( P2_U7612 , P2_U2358 , P2_EBX_REG_5_ );
nand NAND2_11689 ( P2_U7613 , P2_INSTADDRPOINTER_REG_4_ , P2_U7592 );
nand NAND2_11690 ( P2_U7614 , P2_PHYADDRPOINTER_REG_4_ , P2_STATE2_REG_1_ );
nand NAND2_11691 ( P2_U7615 , P2_U4423 , P2_REIP_REG_4_ );
nand NAND2_11692 ( P2_U7616 , P2_U2358 , P2_EBX_REG_4_ );
nand NAND2_11693 ( P2_U7617 , P2_INSTADDRPOINTER_REG_31_ , P2_U7592 );
nand NAND2_11694 ( P2_U7618 , P2_PHYADDRPOINTER_REG_31_ , P2_STATE2_REG_1_ );
nand NAND2_11695 ( P2_U7619 , P2_U4423 , P2_REIP_REG_31_ );
nand NAND2_11696 ( P2_U7620 , P2_U2358 , P2_EBX_REG_31_ );
nand NAND2_11697 ( P2_U7621 , P2_INSTADDRPOINTER_REG_30_ , P2_U7592 );
nand NAND2_11698 ( P2_U7622 , P2_PHYADDRPOINTER_REG_30_ , P2_STATE2_REG_1_ );
nand NAND2_11699 ( P2_U7623 , P2_U4423 , P2_REIP_REG_30_ );
nand NAND2_11700 ( P2_U7624 , P2_U2358 , P2_EBX_REG_30_ );
nand NAND2_11701 ( P2_U7625 , P2_INSTADDRPOINTER_REG_3_ , P2_U7592 );
nand NAND2_11702 ( P2_U7626 , P2_PHYADDRPOINTER_REG_3_ , P2_STATE2_REG_1_ );
nand NAND2_11703 ( P2_U7627 , P2_U4423 , P2_REIP_REG_3_ );
nand NAND2_11704 ( P2_U7628 , P2_U2358 , P2_EBX_REG_3_ );
nand NAND2_11705 ( P2_U7629 , P2_INSTADDRPOINTER_REG_29_ , P2_U7592 );
nand NAND2_11706 ( P2_U7630 , P2_PHYADDRPOINTER_REG_29_ , P2_STATE2_REG_1_ );
nand NAND2_11707 ( P2_U7631 , P2_U4423 , P2_REIP_REG_29_ );
nand NAND2_11708 ( P2_U7632 , P2_U2358 , P2_EBX_REG_29_ );
nand NAND2_11709 ( P2_U7633 , P2_INSTADDRPOINTER_REG_28_ , P2_U7592 );
nand NAND2_11710 ( P2_U7634 , P2_PHYADDRPOINTER_REG_28_ , P2_STATE2_REG_1_ );
nand NAND2_11711 ( P2_U7635 , P2_U4423 , P2_REIP_REG_28_ );
nand NAND2_11712 ( P2_U7636 , P2_U2358 , P2_EBX_REG_28_ );
nand NAND2_11713 ( P2_U7637 , P2_INSTADDRPOINTER_REG_27_ , P2_U7592 );
nand NAND2_11714 ( P2_U7638 , P2_PHYADDRPOINTER_REG_27_ , P2_STATE2_REG_1_ );
nand NAND2_11715 ( P2_U7639 , P2_U4423 , P2_REIP_REG_27_ );
nand NAND2_11716 ( P2_U7640 , P2_U2358 , P2_EBX_REG_27_ );
nand NAND2_11717 ( P2_U7641 , P2_INSTADDRPOINTER_REG_26_ , P2_U7592 );
nand NAND2_11718 ( P2_U7642 , P2_PHYADDRPOINTER_REG_26_ , P2_STATE2_REG_1_ );
nand NAND2_11719 ( P2_U7643 , P2_U4423 , P2_REIP_REG_26_ );
nand NAND2_11720 ( P2_U7644 , P2_U2358 , P2_EBX_REG_26_ );
nand NAND2_11721 ( P2_U7645 , P2_INSTADDRPOINTER_REG_25_ , P2_U7592 );
nand NAND2_11722 ( P2_U7646 , P2_PHYADDRPOINTER_REG_25_ , P2_STATE2_REG_1_ );
nand NAND2_11723 ( P2_U7647 , P2_U4423 , P2_REIP_REG_25_ );
nand NAND2_11724 ( P2_U7648 , P2_U2358 , P2_EBX_REG_25_ );
nand NAND2_11725 ( P2_U7649 , P2_INSTADDRPOINTER_REG_24_ , P2_U7592 );
nand NAND2_11726 ( P2_U7650 , P2_PHYADDRPOINTER_REG_24_ , P2_STATE2_REG_1_ );
nand NAND2_11727 ( P2_U7651 , P2_U4423 , P2_REIP_REG_24_ );
nand NAND2_11728 ( P2_U7652 , P2_U2358 , P2_EBX_REG_24_ );
nand NAND2_11729 ( P2_U7653 , P2_INSTADDRPOINTER_REG_23_ , P2_U7592 );
nand NAND2_11730 ( P2_U7654 , P2_PHYADDRPOINTER_REG_23_ , P2_STATE2_REG_1_ );
nand NAND2_11731 ( P2_U7655 , P2_U4423 , P2_REIP_REG_23_ );
nand NAND2_11732 ( P2_U7656 , P2_U2358 , P2_EBX_REG_23_ );
nand NAND2_11733 ( P2_U7657 , P2_INSTADDRPOINTER_REG_22_ , P2_U7592 );
nand NAND2_11734 ( P2_U7658 , P2_PHYADDRPOINTER_REG_22_ , P2_STATE2_REG_1_ );
nand NAND2_11735 ( P2_U7659 , P2_U4423 , P2_REIP_REG_22_ );
nand NAND2_11736 ( P2_U7660 , P2_U2358 , P2_EBX_REG_22_ );
nand NAND2_11737 ( P2_U7661 , P2_INSTADDRPOINTER_REG_21_ , P2_U7592 );
nand NAND2_11738 ( P2_U7662 , P2_PHYADDRPOINTER_REG_21_ , P2_STATE2_REG_1_ );
nand NAND2_11739 ( P2_U7663 , P2_U4423 , P2_REIP_REG_21_ );
nand NAND2_11740 ( P2_U7664 , P2_U2358 , P2_EBX_REG_21_ );
nand NAND2_11741 ( P2_U7665 , P2_INSTADDRPOINTER_REG_20_ , P2_U7592 );
nand NAND2_11742 ( P2_U7666 , P2_PHYADDRPOINTER_REG_20_ , P2_STATE2_REG_1_ );
nand NAND2_11743 ( P2_U7667 , P2_U4423 , P2_REIP_REG_20_ );
nand NAND2_11744 ( P2_U7668 , P2_U2358 , P2_EBX_REG_20_ );
nand NAND2_11745 ( P2_U7669 , P2_INSTADDRPOINTER_REG_2_ , P2_U7592 );
nand NAND2_11746 ( P2_U7670 , P2_PHYADDRPOINTER_REG_2_ , P2_STATE2_REG_1_ );
nand NAND2_11747 ( P2_U7671 , P2_U4423 , P2_REIP_REG_2_ );
nand NAND2_11748 ( P2_U7672 , P2_U2358 , P2_EBX_REG_2_ );
nand NAND2_11749 ( P2_U7673 , P2_INSTADDRPOINTER_REG_19_ , P2_U7592 );
nand NAND2_11750 ( P2_U7674 , P2_PHYADDRPOINTER_REG_19_ , P2_STATE2_REG_1_ );
nand NAND2_11751 ( P2_U7675 , P2_U4423 , P2_REIP_REG_19_ );
nand NAND2_11752 ( P2_U7676 , P2_U2358 , P2_EBX_REG_19_ );
nand NAND2_11753 ( P2_U7677 , P2_INSTADDRPOINTER_REG_18_ , P2_U7592 );
nand NAND2_11754 ( P2_U7678 , P2_PHYADDRPOINTER_REG_18_ , P2_STATE2_REG_1_ );
nand NAND2_11755 ( P2_U7679 , P2_U4423 , P2_REIP_REG_18_ );
nand NAND2_11756 ( P2_U7680 , P2_U2358 , P2_EBX_REG_18_ );
nand NAND2_11757 ( P2_U7681 , P2_INSTADDRPOINTER_REG_17_ , P2_U7592 );
nand NAND2_11758 ( P2_U7682 , P2_PHYADDRPOINTER_REG_17_ , P2_STATE2_REG_1_ );
nand NAND2_11759 ( P2_U7683 , P2_U4423 , P2_REIP_REG_17_ );
nand NAND2_11760 ( P2_U7684 , P2_U2358 , P2_EBX_REG_17_ );
nand NAND2_11761 ( P2_U7685 , P2_INSTADDRPOINTER_REG_16_ , P2_U7592 );
nand NAND2_11762 ( P2_U7686 , P2_PHYADDRPOINTER_REG_16_ , P2_STATE2_REG_1_ );
nand NAND2_11763 ( P2_U7687 , P2_U4423 , P2_REIP_REG_16_ );
nand NAND2_11764 ( P2_U7688 , P2_U2358 , P2_EBX_REG_16_ );
nand NAND2_11765 ( P2_U7689 , P2_INSTADDRPOINTER_REG_15_ , P2_U7592 );
nand NAND2_11766 ( P2_U7690 , P2_PHYADDRPOINTER_REG_15_ , P2_STATE2_REG_1_ );
nand NAND2_11767 ( P2_U7691 , P2_U4423 , P2_REIP_REG_15_ );
nand NAND2_11768 ( P2_U7692 , P2_U2358 , P2_EBX_REG_15_ );
nand NAND2_11769 ( P2_U7693 , P2_INSTADDRPOINTER_REG_14_ , P2_U7592 );
nand NAND2_11770 ( P2_U7694 , P2_PHYADDRPOINTER_REG_14_ , P2_STATE2_REG_1_ );
nand NAND2_11771 ( P2_U7695 , P2_U4423 , P2_REIP_REG_14_ );
nand NAND2_11772 ( P2_U7696 , P2_U2358 , P2_EBX_REG_14_ );
nand NAND2_11773 ( P2_U7697 , P2_INSTADDRPOINTER_REG_13_ , P2_U7592 );
nand NAND2_11774 ( P2_U7698 , P2_PHYADDRPOINTER_REG_13_ , P2_STATE2_REG_1_ );
nand NAND2_11775 ( P2_U7699 , P2_U4423 , P2_REIP_REG_13_ );
nand NAND2_11776 ( P2_U7700 , P2_U2358 , P2_EBX_REG_13_ );
nand NAND2_11777 ( P2_U7701 , P2_INSTADDRPOINTER_REG_12_ , P2_U7592 );
nand NAND2_11778 ( P2_U7702 , P2_PHYADDRPOINTER_REG_12_ , P2_STATE2_REG_1_ );
nand NAND2_11779 ( P2_U7703 , P2_U4423 , P2_REIP_REG_12_ );
nand NAND2_11780 ( P2_U7704 , P2_U2358 , P2_EBX_REG_12_ );
nand NAND2_11781 ( P2_U7705 , P2_INSTADDRPOINTER_REG_11_ , P2_U7592 );
nand NAND2_11782 ( P2_U7706 , P2_PHYADDRPOINTER_REG_11_ , P2_STATE2_REG_1_ );
nand NAND2_11783 ( P2_U7707 , P2_U4423 , P2_REIP_REG_11_ );
nand NAND2_11784 ( P2_U7708 , P2_U2358 , P2_EBX_REG_11_ );
nand NAND2_11785 ( P2_U7709 , P2_INSTADDRPOINTER_REG_10_ , P2_U7592 );
nand NAND2_11786 ( P2_U7710 , P2_PHYADDRPOINTER_REG_10_ , P2_STATE2_REG_1_ );
nand NAND2_11787 ( P2_U7711 , P2_U4423 , P2_REIP_REG_10_ );
nand NAND2_11788 ( P2_U7712 , P2_U2358 , P2_EBX_REG_10_ );
nand NAND2_11789 ( P2_U7713 , P2_INSTADDRPOINTER_REG_1_ , P2_U7592 );
nand NAND2_11790 ( P2_U7714 , P2_PHYADDRPOINTER_REG_1_ , P2_STATE2_REG_1_ );
nand NAND2_11791 ( P2_U7715 , P2_U4423 , P2_REIP_REG_1_ );
nand NAND2_11792 ( P2_U7716 , P2_U2358 , P2_EBX_REG_1_ );
nand NAND2_11793 ( P2_U7717 , P2_U4387 , P2_U7885 );
nand NAND2_11794 ( P2_U7718 , P2_INSTADDRPOINTER_REG_0_ , P2_U7739 );
nand NAND2_11795 ( P2_U7719 , P2_PHYADDRPOINTER_REG_0_ , P2_STATE2_REG_1_ );
nand NAND2_11796 ( P2_U7720 , P2_U4423 , P2_REIP_REG_0_ );
nand NAND2_11797 ( P2_U7721 , P2_U2358 , P2_EBX_REG_0_ );
nand NAND2_11798 ( P2_U7722 , P2_U7720 , P2_U3575 );
nand NAND2_11799 ( P2_U7723 , P2_U3550 , P2_U3536 );
nand NAND2_11800 ( P2_U7724 , P2_R2219_U28 , P2_U7723 );
nand NAND2_11801 ( P2_U7725 , P2_R2219_U30 , P2_U7723 );
nand NAND2_11802 ( P2_U7726 , P2_R2238_U19 , P2_U2356 );
nand NAND2_11803 ( P2_U7727 , P2_INSTQUEUERD_ADDR_REG_4_ , P2_U3284 );
nand NAND2_11804 ( P2_U7728 , P2_R2238_U20 , P2_U2356 );
nand NAND2_11805 ( P2_U7729 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3284 );
nand NAND2_11806 ( P2_U7730 , P2_R2238_U21 , P2_U2356 );
nand NAND2_11807 ( P2_U7731 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_U3284 );
nand NAND2_11808 ( P2_U7732 , P2_R2238_U22 , P2_U2356 );
nand NAND2_11809 ( P2_U7733 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_U3284 );
nand NAND2_11810 ( P2_U7734 , P2_R2238_U7 , P2_U2356 );
nand NAND2_11811 ( P2_U7735 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_U3284 );
nand NAND3_11812 ( P2_U7736 , P2_U3295 , P2_U7873 , P2_U3525 );
nand NAND4_11813 ( P2_U7737 , P2_U7590 , P2_U7589 , P2_U4422 , P2_U3272 );
nand NAND2_11814 ( P2_U7738 , P2_U7861 , P2_U2617 );
nand NAND4_11815 ( P2_U7739 , P2_U7591 , P2_U3285 , P2_U4422 , P2_U3539 );
nand NAND4_11816 ( P2_U7740 , P2_U3521 , P2_U7744 , P2_U5573 , P2_U5571 );
nand NAND2_11817 ( P2_U7741 , P2_U2391 , P2_U3544 );
nand NAND2_11818 ( P2_U7742 , P2_U2377 , P2_U6572 );
nand NAND3_11819 ( P2_U7743 , P2_U7741 , P2_U4448 , P2_U7742 );
nand NAND2_11820 ( P2_U7744 , P2_U7745 , P2_U3278 );
nand NAND2_11821 ( P2_U7745 , P2_U7861 , P2_U2617 );
nand NAND3_11822 ( P2_U7746 , P2_U8003 , P2_U8002 , P2_U4592 );
nand NAND3_11823 ( P2_U7747 , P2_U7971 , P2_U7970 , P2_U4592 );
nand NAND3_11824 ( P2_U7748 , P2_U7955 , P2_U7954 , P2_U4592 );
nand NAND3_11825 ( P2_U7749 , P2_U8035 , P2_U8034 , P2_U4592 );
nand NAND3_11826 ( P2_U7750 , P2_U8019 , P2_U8018 , P2_U4592 );
nand NAND3_11827 ( P2_U7751 , P2_U7987 , P2_U7986 , P2_U4592 );
nand NAND3_11828 ( P2_U7752 , P2_U7939 , P2_U7938 , P2_U4592 );
nand NAND3_11829 ( P2_U7753 , P2_U7923 , P2_U7922 , P2_U4592 );
nand NAND3_11830 ( P2_U7754 , P2_U8154 , P2_U8153 , P2_U4592 );
nand NAND3_11831 ( P2_U7755 , P2_U8170 , P2_U8169 , P2_U4592 );
nand NAND3_11832 ( P2_U7756 , P2_U8186 , P2_U8185 , P2_U4592 );
nand NAND3_11833 ( P2_U7757 , P2_U8202 , P2_U8201 , P2_U4592 );
nand NAND3_11834 ( P2_U7758 , P2_U8218 , P2_U8217 , P2_U4592 );
nand NAND3_11835 ( P2_U7759 , P2_U8234 , P2_U8233 , P2_U4592 );
nand NAND3_11836 ( P2_U7760 , P2_U8250 , P2_U8249 , P2_U4592 );
nand NAND3_11837 ( P2_U7761 , P2_U8266 , P2_U8265 , P2_U4592 );
nand NAND3_11838 ( P2_U7762 , P2_U8005 , P2_U8004 , P2_U4593 );
nand NAND3_11839 ( P2_U7763 , P2_U7973 , P2_U7972 , P2_U4593 );
nand NAND3_11840 ( P2_U7764 , P2_U7957 , P2_U7956 , P2_U4593 );
nand NAND3_11841 ( P2_U7765 , P2_U8037 , P2_U8036 , P2_U4593 );
nand NAND3_11842 ( P2_U7766 , P2_U8021 , P2_U8020 , P2_U4593 );
nand NAND3_11843 ( P2_U7767 , P2_U7989 , P2_U7988 , P2_U4593 );
nand NAND3_11844 ( P2_U7768 , P2_U7941 , P2_U7940 , P2_U4593 );
nand NAND3_11845 ( P2_U7769 , P2_U7925 , P2_U7924 , P2_U4593 );
nand NAND3_11846 ( P2_U7770 , P2_U8156 , P2_U8155 , P2_U4593 );
nand NAND3_11847 ( P2_U7771 , P2_U8172 , P2_U8171 , P2_U4593 );
nand NAND3_11848 ( P2_U7772 , P2_U8188 , P2_U8187 , P2_U4593 );
nand NAND3_11849 ( P2_U7773 , P2_U8204 , P2_U8203 , P2_U4593 );
nand NAND3_11850 ( P2_U7774 , P2_U8220 , P2_U8219 , P2_U4593 );
nand NAND3_11851 ( P2_U7775 , P2_U8236 , P2_U8235 , P2_U4593 );
nand NAND3_11852 ( P2_U7776 , P2_U8252 , P2_U8251 , P2_U4593 );
nand NAND3_11853 ( P2_U7777 , P2_U8268 , P2_U8267 , P2_U4593 );
nand NAND3_11854 ( P2_U7778 , P2_U8007 , P2_U8006 , P2_U2456 );
nand NAND3_11855 ( P2_U7779 , P2_U7975 , P2_U7974 , P2_U2456 );
nand NAND3_11856 ( P2_U7780 , P2_U7959 , P2_U7958 , P2_U2456 );
nand NAND3_11857 ( P2_U7781 , P2_U8039 , P2_U8038 , P2_U2456 );
nand NAND3_11858 ( P2_U7782 , P2_U8023 , P2_U8022 , P2_U2456 );
nand NAND3_11859 ( P2_U7783 , P2_U7991 , P2_U7990 , P2_U2456 );
nand NAND3_11860 ( P2_U7784 , P2_U7943 , P2_U7942 , P2_U2456 );
nand NAND3_11861 ( P2_U7785 , P2_U7927 , P2_U7926 , P2_U2456 );
nand NAND3_11862 ( P2_U7786 , P2_U8158 , P2_U8157 , P2_U2456 );
nand NAND3_11863 ( P2_U7787 , P2_U8174 , P2_U8173 , P2_U2456 );
nand NAND3_11864 ( P2_U7788 , P2_U8190 , P2_U8189 , P2_U2456 );
nand NAND3_11865 ( P2_U7789 , P2_U8206 , P2_U8205 , P2_U2456 );
nand NAND3_11866 ( P2_U7790 , P2_U8222 , P2_U8221 , P2_U2456 );
nand NAND3_11867 ( P2_U7791 , P2_U8238 , P2_U8237 , P2_U2456 );
nand NAND3_11868 ( P2_U7792 , P2_U8254 , P2_U8253 , P2_U2456 );
nand NAND3_11869 ( P2_U7793 , P2_U8270 , P2_U8269 , P2_U2456 );
nand NAND3_11870 ( P2_U7794 , P2_U8009 , P2_U8008 , P2_U2454 );
nand NAND3_11871 ( P2_U7795 , P2_U7977 , P2_U7976 , P2_U2454 );
nand NAND3_11872 ( P2_U7796 , P2_U7961 , P2_U7960 , P2_U2454 );
nand NAND3_11873 ( P2_U7797 , P2_U8041 , P2_U8040 , P2_U2454 );
nand NAND3_11874 ( P2_U7798 , P2_U8025 , P2_U8024 , P2_U2454 );
nand NAND3_11875 ( P2_U7799 , P2_U7993 , P2_U7992 , P2_U2454 );
nand NAND3_11876 ( P2_U7800 , P2_U7945 , P2_U7944 , P2_U2454 );
nand NAND3_11877 ( P2_U7801 , P2_U7929 , P2_U7928 , P2_U2454 );
nand NAND3_11878 ( P2_U7802 , P2_U8160 , P2_U8159 , P2_U2454 );
nand NAND3_11879 ( P2_U7803 , P2_U8176 , P2_U8175 , P2_U2454 );
nand NAND3_11880 ( P2_U7804 , P2_U8192 , P2_U8191 , P2_U2454 );
nand NAND3_11881 ( P2_U7805 , P2_U8208 , P2_U8207 , P2_U2454 );
nand NAND3_11882 ( P2_U7806 , P2_U8224 , P2_U8223 , P2_U2454 );
nand NAND3_11883 ( P2_U7807 , P2_U8240 , P2_U8239 , P2_U2454 );
nand NAND3_11884 ( P2_U7808 , P2_U8256 , P2_U8255 , P2_U2454 );
nand NAND3_11885 ( P2_U7809 , P2_U8272 , P2_U8271 , P2_U2454 );
nand NAND3_11886 ( P2_U7810 , P2_U8011 , P2_U8010 , P2_U4590 );
nand NAND3_11887 ( P2_U7811 , P2_U7979 , P2_U7978 , P2_U4590 );
nand NAND3_11888 ( P2_U7812 , P2_U7963 , P2_U7962 , P2_U4590 );
nand NAND3_11889 ( P2_U7813 , P2_U8043 , P2_U8042 , P2_U4590 );
nand NAND3_11890 ( P2_U7814 , P2_U8027 , P2_U8026 , P2_U4590 );
nand NAND3_11891 ( P2_U7815 , P2_U7995 , P2_U7994 , P2_U4590 );
nand NAND3_11892 ( P2_U7816 , P2_U7947 , P2_U7946 , P2_U4590 );
nand NAND3_11893 ( P2_U7817 , P2_U7931 , P2_U7930 , P2_U4590 );
nand NAND3_11894 ( P2_U7818 , P2_U8162 , P2_U8161 , P2_U4590 );
nand NAND3_11895 ( P2_U7819 , P2_U8178 , P2_U8177 , P2_U4590 );
nand NAND3_11896 ( P2_U7820 , P2_U8194 , P2_U8193 , P2_U4590 );
nand NAND3_11897 ( P2_U7821 , P2_U8210 , P2_U8209 , P2_U4590 );
nand NAND3_11898 ( P2_U7822 , P2_U8226 , P2_U8225 , P2_U4590 );
nand NAND3_11899 ( P2_U7823 , P2_U8242 , P2_U8241 , P2_U4590 );
nand NAND3_11900 ( P2_U7824 , P2_U8258 , P2_U8257 , P2_U4590 );
nand NAND3_11901 ( P2_U7825 , P2_U8274 , P2_U8273 , P2_U4590 );
nand NAND3_11902 ( P2_U7826 , P2_U8013 , P2_U8012 , P2_U2453 );
nand NAND3_11903 ( P2_U7827 , P2_U7981 , P2_U7980 , P2_U2453 );
nand NAND3_11904 ( P2_U7828 , P2_U7965 , P2_U7964 , P2_U2453 );
nand NAND3_11905 ( P2_U7829 , P2_U8045 , P2_U8044 , P2_U2453 );
nand NAND3_11906 ( P2_U7830 , P2_U8029 , P2_U8028 , P2_U2453 );
nand NAND3_11907 ( P2_U7831 , P2_U7997 , P2_U7996 , P2_U2453 );
nand NAND3_11908 ( P2_U7832 , P2_U7949 , P2_U7948 , P2_U2453 );
nand NAND3_11909 ( P2_U7833 , P2_U7933 , P2_U7932 , P2_U2453 );
nand NAND3_11910 ( P2_U7834 , P2_U8164 , P2_U8163 , P2_U2453 );
nand NAND3_11911 ( P2_U7835 , P2_U8180 , P2_U8179 , P2_U2453 );
nand NAND3_11912 ( P2_U7836 , P2_U8196 , P2_U8195 , P2_U2453 );
nand NAND3_11913 ( P2_U7837 , P2_U8212 , P2_U8211 , P2_U2453 );
nand NAND3_11914 ( P2_U7838 , P2_U8228 , P2_U8227 , P2_U2453 );
nand NAND3_11915 ( P2_U7839 , P2_U8244 , P2_U8243 , P2_U2453 );
nand NAND3_11916 ( P2_U7840 , P2_U8260 , P2_U8259 , P2_U2453 );
nand NAND3_11917 ( P2_U7841 , P2_U8276 , P2_U8275 , P2_U2453 );
nand NAND3_11918 ( P2_U7842 , P2_U8015 , P2_U8014 , P2_U2452 );
nand NAND3_11919 ( P2_U7843 , P2_U7983 , P2_U7982 , P2_U2452 );
nand NAND3_11920 ( P2_U7844 , P2_U7967 , P2_U7966 , P2_U2452 );
nand NAND3_11921 ( P2_U7845 , P2_U8047 , P2_U8046 , P2_U2452 );
nand NAND3_11922 ( P2_U7846 , P2_U8031 , P2_U8030 , P2_U2452 );
nand NAND3_11923 ( P2_U7847 , P2_U7999 , P2_U7998 , P2_U2452 );
nand NAND3_11924 ( P2_U7848 , P2_U7951 , P2_U7950 , P2_U2452 );
nand NAND3_11925 ( P2_U7849 , P2_U7935 , P2_U7934 , P2_U2452 );
nand NAND3_11926 ( P2_U7850 , P2_U8166 , P2_U8165 , P2_U2452 );
nand NAND3_11927 ( P2_U7851 , P2_U8182 , P2_U8181 , P2_U2452 );
nand NAND3_11928 ( P2_U7852 , P2_U8198 , P2_U8197 , P2_U2452 );
nand NAND3_11929 ( P2_U7853 , P2_U8214 , P2_U8213 , P2_U2452 );
nand NAND3_11930 ( P2_U7854 , P2_U8230 , P2_U8229 , P2_U2452 );
nand NAND3_11931 ( P2_U7855 , P2_U8246 , P2_U8245 , P2_U2452 );
nand NAND3_11932 ( P2_U7856 , P2_U8262 , P2_U8261 , P2_U2452 );
nand NAND3_11933 ( P2_U7857 , P2_U8278 , P2_U8277 , P2_U2452 );
nand NAND3_11934 ( P2_U7858 , P2_U8017 , P2_U8016 , P2_U2455 );
not NOT1_11935 ( P2_U7859 , P2_U3280 );
nand NAND3_11936 ( P2_U7860 , P2_U7985 , P2_U7984 , P2_U2455 );
not NOT1_11937 ( P2_U7861 , P2_U3279 );
nand NAND3_11938 ( P2_U7862 , P2_U7969 , P2_U7968 , P2_U2455 );
not NOT1_11939 ( P2_U7863 , P2_U3278 );
nand NAND3_11940 ( P2_U7864 , P2_U8049 , P2_U8048 , P2_U2455 );
not NOT1_11941 ( P2_U7865 , P2_U3521 );
nand NAND3_11942 ( P2_U7866 , P2_U8033 , P2_U8032 , P2_U2455 );
not NOT1_11943 ( P2_U7867 , P2_U3255 );
nand NAND3_11944 ( P2_U7868 , P2_U8001 , P2_U8000 , P2_U2455 );
not NOT1_11945 ( P2_U7869 , P2_U2617 );
nand NAND3_11946 ( P2_U7870 , P2_U7953 , P2_U7952 , P2_U2455 );
not NOT1_11947 ( P2_U7871 , P2_U3253 );
nand NAND3_11948 ( P2_U7872 , P2_U7937 , P2_U7936 , P2_U2455 );
not NOT1_11949 ( P2_U7873 , P2_U2616 );
nand NAND3_11950 ( P2_U7874 , P2_U8168 , P2_U8167 , P2_U2455 );
nand NAND3_11951 ( P2_U7875 , P2_U8184 , P2_U8183 , P2_U2455 );
nand NAND3_11952 ( P2_U7876 , P2_U8200 , P2_U8199 , P2_U2455 );
nand NAND3_11953 ( P2_U7877 , P2_U8216 , P2_U8215 , P2_U2455 );
nand NAND3_11954 ( P2_U7878 , P2_U8232 , P2_U8231 , P2_U2455 );
nand NAND3_11955 ( P2_U7879 , P2_U8248 , P2_U8247 , P2_U2455 );
nand NAND3_11956 ( P2_U7880 , P2_U8264 , P2_U8263 , P2_U2455 );
nand NAND3_11957 ( P2_U7881 , P2_U8280 , P2_U8279 , P2_U2455 );
nand NAND2_11958 ( P2_U7882 , P2_U5590 , P2_U4428 );
nand NAND2_11959 ( P2_U7883 , P2_U5596 , P2_U3525 );
nand NAND2_11960 ( P2_U7884 , P2_U4596 , P2_U7883 );
nand NAND3_11961 ( P2_U7885 , P2_U8348 , P2_U8347 , P2_U3253 );
nand NAND2_11962 ( P2_U7886 , P2_U7722 , P2_U5589 );
nand NAND2_11963 ( P2_U7887 , P2_U4459 , P2_U5589 );
nand NAND5_11964 ( P2_U7888 , P2_U4386 , P2_U7887 , P2_U2589 , P2_U4385 , P2_U4384 );
nand NAND2_11965 ( P2_U7889 , P2_U4459 , P2_U5589 );
nand NAND4_11966 ( P2_U7890 , P2_U7889 , P2_U4458 , P2_U2589 , P2_U4379 );
nand NAND3_11967 ( P2_U7891 , P2_U4572 , P2_STATE_REG_1_ , P2_U4569 );
nand NAND3_11968 ( P2_U7892 , P2_REQUESTPENDING_REG , P2_U3244 , P2_STATE_REG_0_ );
nand NAND2_11969 ( P2_U7893 , P2_STATE_REG_1_ , P2_U4569 );
nand NAND2_11970 ( P2_U7894 , P2_U4600 , P2_U4615 );
nand NAND2_11971 ( P2_U7895 , P2_U7863 , P2_U7871 );
nand NAND2_11972 ( P2_U7896 , P2_U3255 , P2_U5595 );
nand NAND2_11973 ( P2_U7897 , P2_U4429 , P2_U5589 );
nand NAND2_11974 ( P2_U7898 , P2_REIP_REG_0_ , P2_DATAWIDTH_REG_0_ );
nand NAND2_11975 ( P2_U7899 , P2_BE_N_REG_3_ , P2_U3259 );
nand NAND2_11976 ( P2_U7900 , P2_BYTEENABLE_REG_3_ , P2_U4439 );
nand NAND2_11977 ( P2_U7901 , P2_BE_N_REG_2_ , P2_U3259 );
nand NAND2_11978 ( P2_U7902 , P2_BYTEENABLE_REG_2_ , P2_U4439 );
nand NAND2_11979 ( P2_U7903 , P2_BE_N_REG_1_ , P2_U3259 );
nand NAND2_11980 ( P2_U7904 , P2_BYTEENABLE_REG_1_ , P2_U4439 );
nand NAND2_11981 ( P2_U7905 , P2_BE_N_REG_0_ , P2_U3259 );
nand NAND2_11982 ( P2_U7906 , P2_BYTEENABLE_REG_0_ , P2_U4439 );
nand NAND3_11983 ( P2_U7907 , P2_U3268 , P2_U3267 , P2_STATE_REG_0_ );
or OR2_11984 ( P2_U7908 , NA , P2_STATE_REG_0_ );
nand NAND2_11985 ( P2_U7909 , P2_STATE_REG_2_ , P2_U3266 );
nand NAND2_11986 ( P2_U7910 , P2_U4568 , P2_STATE_REG_0_ );
nand NAND3_11987 ( P2_U7911 , P2_U4581 , P2_U4572 , P2_STATE_REG_1_ );
nand NAND2_11988 ( P2_U7912 , P2_U4582 , P2_U3258 );
nand NAND3_11989 ( P2_U7913 , P2_STATE_REG_0_ , P2_U3267 , P2_STATE_REG_2_ );
nand NAND2_11990 ( P2_U7914 , P2_U4584 , P2_U3244 );
or OR2_11991 ( P2_U7915 , P2_STATE_REG_0_ , P2_STATE_REG_1_ );
nand NAND2_11992 ( P2_U7916 , P2_STATE_REG_0_ , P2_U4473 );
not NOT1_11993 ( P2_U7917 , P2_U3589 );
nand NAND2_11994 ( P2_U7918 , P2_U7917 , P2_DATAWIDTH_REG_0_ );
nand NAND2_11995 ( P2_U7919 , P2_U3590 , P2_U3589 );
nand NAND2_11996 ( P2_U7920 , P2_U3589 , P2_U4589 );
nand NAND2_11997 ( P2_U7921 , P2_U7917 , P2_DATAWIDTH_REG_1_ );
nand NAND2_11998 ( P2_U7922 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3388 );
or OR2_11999 ( P2_U7923 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_3__1_ );
or OR2_12000 ( P2_U7924 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_0__1_ );
nand NAND2_12001 ( P2_U7925 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3422 );
or OR2_12002 ( P2_U7926 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_1__1_ );
nand NAND2_12003 ( P2_U7927 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3411 );
nand NAND2_12004 ( P2_U7928 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3374 );
or OR2_12005 ( P2_U7929 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_4__1_ );
nand NAND2_12006 ( P2_U7930 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3333 );
or OR2_12007 ( P2_U7931 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_7__1_ );
nand NAND2_12008 ( P2_U7932 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3363 );
or OR2_12009 ( P2_U7933 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_5__1_ );
nand NAND2_12010 ( P2_U7934 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3347 );
or OR2_12011 ( P2_U7935 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_6__1_ );
nand NAND2_12012 ( P2_U7936 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3399 );
or OR2_12013 ( P2_U7937 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_2__1_ );
nand NAND2_12014 ( P2_U7938 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3389 );
or OR2_12015 ( P2_U7939 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_3__0_ );
or OR2_12016 ( P2_U7940 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_0__0_ );
nand NAND2_12017 ( P2_U7941 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3423 );
or OR2_12018 ( P2_U7942 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_1__0_ );
nand NAND2_12019 ( P2_U7943 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3412 );
nand NAND2_12020 ( P2_U7944 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3375 );
or OR2_12021 ( P2_U7945 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_4__0_ );
nand NAND2_12022 ( P2_U7946 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3334 );
or OR2_12023 ( P2_U7947 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_7__0_ );
nand NAND2_12024 ( P2_U7948 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3364 );
or OR2_12025 ( P2_U7949 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_5__0_ );
nand NAND2_12026 ( P2_U7950 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3348 );
or OR2_12027 ( P2_U7951 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_6__0_ );
nand NAND2_12028 ( P2_U7952 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3400 );
or OR2_12029 ( P2_U7953 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_2__0_ );
nand NAND2_12030 ( P2_U7954 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3385 );
or OR2_12031 ( P2_U7955 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_3__4_ );
or OR2_12032 ( P2_U7956 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_0__4_ );
nand NAND2_12033 ( P2_U7957 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3419 );
or OR2_12034 ( P2_U7958 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_1__4_ );
nand NAND2_12035 ( P2_U7959 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3408 );
nand NAND2_12036 ( P2_U7960 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3371 );
or OR2_12037 ( P2_U7961 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_4__4_ );
nand NAND2_12038 ( P2_U7962 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3330 );
or OR2_12039 ( P2_U7963 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_7__4_ );
nand NAND2_12040 ( P2_U7964 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3360 );
or OR2_12041 ( P2_U7965 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_5__4_ );
nand NAND2_12042 ( P2_U7966 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3344 );
or OR2_12043 ( P2_U7967 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_6__4_ );
nand NAND2_12044 ( P2_U7968 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3396 );
or OR2_12045 ( P2_U7969 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_2__4_ );
nand NAND2_12046 ( P2_U7970 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3383 );
or OR2_12047 ( P2_U7971 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_3__6_ );
or OR2_12048 ( P2_U7972 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_0__6_ );
nand NAND2_12049 ( P2_U7973 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3417 );
or OR2_12050 ( P2_U7974 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_1__6_ );
nand NAND2_12051 ( P2_U7975 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3406 );
nand NAND2_12052 ( P2_U7976 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3369 );
or OR2_12053 ( P2_U7977 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_4__6_ );
nand NAND2_12054 ( P2_U7978 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3328 );
or OR2_12055 ( P2_U7979 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_7__6_ );
nand NAND2_12056 ( P2_U7980 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3358 );
or OR2_12057 ( P2_U7981 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_5__6_ );
nand NAND2_12058 ( P2_U7982 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3342 );
or OR2_12059 ( P2_U7983 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_6__6_ );
nand NAND2_12060 ( P2_U7984 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3394 );
or OR2_12061 ( P2_U7985 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_2__6_ );
nand NAND2_12062 ( P2_U7986 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3384 );
or OR2_12063 ( P2_U7987 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_3__5_ );
or OR2_12064 ( P2_U7988 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_0__5_ );
nand NAND2_12065 ( P2_U7989 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3418 );
or OR2_12066 ( P2_U7990 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_1__5_ );
nand NAND2_12067 ( P2_U7991 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3407 );
nand NAND2_12068 ( P2_U7992 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3370 );
or OR2_12069 ( P2_U7993 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_4__5_ );
nand NAND2_12070 ( P2_U7994 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3329 );
or OR2_12071 ( P2_U7995 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_7__5_ );
nand NAND2_12072 ( P2_U7996 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3359 );
or OR2_12073 ( P2_U7997 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_5__5_ );
nand NAND2_12074 ( P2_U7998 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3343 );
or OR2_12075 ( P2_U7999 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_6__5_ );
nand NAND2_12076 ( P2_U8000 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3395 );
or OR2_12077 ( P2_U8001 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_2__5_ );
nand NAND2_12078 ( P2_U8002 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3387 );
or OR2_12079 ( P2_U8003 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_3__2_ );
or OR2_12080 ( P2_U8004 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_0__2_ );
nand NAND2_12081 ( P2_U8005 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3421 );
or OR2_12082 ( P2_U8006 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_1__2_ );
nand NAND2_12083 ( P2_U8007 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3410 );
nand NAND2_12084 ( P2_U8008 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3373 );
or OR2_12085 ( P2_U8009 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_4__2_ );
nand NAND2_12086 ( P2_U8010 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3332 );
or OR2_12087 ( P2_U8011 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_7__2_ );
nand NAND2_12088 ( P2_U8012 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3362 );
or OR2_12089 ( P2_U8013 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_5__2_ );
nand NAND2_12090 ( P2_U8014 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3346 );
or OR2_12091 ( P2_U8015 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_6__2_ );
nand NAND2_12092 ( P2_U8016 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3398 );
or OR2_12093 ( P2_U8017 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_2__2_ );
nand NAND2_12094 ( P2_U8018 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3386 );
or OR2_12095 ( P2_U8019 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_3__3_ );
or OR2_12096 ( P2_U8020 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_0__3_ );
nand NAND2_12097 ( P2_U8021 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3420 );
or OR2_12098 ( P2_U8022 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_1__3_ );
nand NAND2_12099 ( P2_U8023 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3409 );
nand NAND2_12100 ( P2_U8024 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3372 );
or OR2_12101 ( P2_U8025 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_4__3_ );
nand NAND2_12102 ( P2_U8026 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3331 );
or OR2_12103 ( P2_U8027 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_7__3_ );
nand NAND2_12104 ( P2_U8028 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3361 );
or OR2_12105 ( P2_U8029 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_5__3_ );
nand NAND2_12106 ( P2_U8030 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3345 );
or OR2_12107 ( P2_U8031 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_6__3_ );
nand NAND2_12108 ( P2_U8032 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3397 );
or OR2_12109 ( P2_U8033 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_2__3_ );
nand NAND2_12110 ( P2_U8034 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3382 );
or OR2_12111 ( P2_U8035 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_3__7_ );
or OR2_12112 ( P2_U8036 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_0__7_ );
nand NAND2_12113 ( P2_U8037 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3416 );
or OR2_12114 ( P2_U8038 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_1__7_ );
nand NAND2_12115 ( P2_U8039 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3405 );
nand NAND2_12116 ( P2_U8040 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3368 );
or OR2_12117 ( P2_U8041 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_4__7_ );
nand NAND2_12118 ( P2_U8042 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3327 );
or OR2_12119 ( P2_U8043 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_7__7_ );
nand NAND2_12120 ( P2_U8044 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3357 );
or OR2_12121 ( P2_U8045 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_5__7_ );
nand NAND2_12122 ( P2_U8046 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3341 );
or OR2_12123 ( P2_U8047 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_6__7_ );
nand NAND2_12124 ( P2_U8048 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3393 );
or OR2_12125 ( P2_U8049 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUE_REG_2__7_ );
nand NAND2_12126 ( P2_U8050 , P2_R2167_U6 , P2_U4435 );
nand NAND2_12127 ( P2_U8051 , P2_U4604 , P2_U3297 );
nand NAND2_12128 ( P2_U8052 , P2_U7871 , P2_U3293 );
nand NAND2_12129 ( P2_U8053 , P2_U3253 , P2_U3282 );
nand NAND2_12130 ( P2_U8054 , P2_U4427 , P2_U3297 );
nand NAND2_12131 ( P2_U8055 , P2_U3289 , P2_U3520 );
or OR2_12132 ( P2_U8056 , U211 , P2_STATE2_REG_0_ );
nand NAND2_12133 ( P2_U8057 , P2_STATE2_REG_0_ , P2_U4617 );
nand NAND2_12134 ( P2_U8058 , P2_STATE2_REG_3_ , P2_U3299 );
nand NAND2_12135 ( P2_U8059 , P2_U2448 , P2_U4620 );
nand NAND2_12136 ( P2_U8060 , P2_STATE2_REG_0_ , P2_U4631 );
nand NAND3_12137 ( P2_U8061 , P2_U4630 , P2_U4619 , P2_U3284 );
nand NAND2_12138 ( P2_U8062 , P2_R2182_U40 , P2_U3318 );
nand NAND2_12139 ( P2_U8063 , P2_U4637 , P2_U3316 );
not NOT1_12140 ( P2_U8064 , P2_U3579 );
nand NAND2_12141 ( P2_U8065 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_U3311 );
nand NAND2_12142 ( P2_U8066 , P2_U4642 , P2_U3310 );
not NOT1_12143 ( P2_U8067 , P2_U3580 );
nand NAND2_12144 ( P2_U8068 , P2_U7859 , P2_U5574 );
nand NAND2_12145 ( P2_U8069 , P2_U3280 , P2_U5575 );
nand NAND2_12146 ( P2_U8070 , P2_U4435 , P2_U3297 );
nand NAND3_12147 ( P2_U8071 , P2_U4433 , P2_U2359 , P2_R2167_U6 );
nand NAND2_12148 ( P2_U8072 , P2_U3594 , P2_U4394 );
nand NAND2_12149 ( P2_U8073 , P2_U5584 , P2_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_12150 ( P2_U8074 , P2_U3280 , P2_U5586 );
nand NAND3_12151 ( P2_U8075 , P2_U2617 , P2_U3279 , P2_U7859 );
nand NAND2_12152 ( P2_U8076 , P2_U4424 , P2_U3253 );
nand NAND2_12153 ( P2_U8077 , P2_U4475 , P2_U7871 );
nand NAND2_12154 ( P2_U8078 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U5585 );
nand NAND3_12155 ( P2_U8079 , P2_U4591 , P2_U3276 , P2_U3273 );
nand NAND2_12156 ( P2_U8080 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3277 );
nand NAND2_12157 ( P2_U8081 , P2_U4590 , P2_U3273 );
not NOT1_12158 ( P2_U8082 , P2_U3581 );
nand NAND2_12159 ( P2_U8083 , P2_U5584 , P2_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_12160 ( P2_U8084 , P2_U5614 , P2_U4394 );
nand NAND2_12161 ( P2_U8085 , P2_INSTADDRPOINTER_REG_0_ , P2_U3528 );
nand NAND2_12162 ( P2_U8086 , P2_U3647 , P2_U3683 );
not NOT1_12163 ( P2_U8087 , P2_U3597 );
nand NAND2_12164 ( P2_U8088 , P2_INSTADDRPOINTER_REG_1_ , P2_U3528 );
nand NAND2_12165 ( P2_U8089 , P2_R1957_U49 , P2_U3647 );
not NOT1_12166 ( P2_U8090 , P2_U3598 );
nand NAND2_12167 ( P2_U8091 , P2_U5616 , P2_U5605 );
nand NAND2_12168 ( P2_U8092 , P2_U3530 , P2_U5606 );
nand NAND2_12169 ( P2_U8093 , P2_U5584 , P2_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_12170 ( P2_U8094 , P2_U5623 , P2_U4394 );
nand NAND3_12171 ( P2_U8095 , P2_U3886 , P2_U4597 , P2_U3255 );
nand NAND3_12172 ( P2_U8096 , P2_U7869 , P2_U5625 , P2_U7867 );
nand NAND2_12173 ( P2_U8097 , P2_U8096 , P2_U8095 );
nand NAND2_12174 ( P2_U8098 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_U3271 );
nand NAND2_12175 ( P2_U8099 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_U3272 );
not NOT1_12176 ( P2_U8100 , P2_U3582 );
nand NAND2_12177 ( P2_U8101 , P2_U5584 , P2_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_12178 ( P2_U8102 , P2_U5633 , P2_U4394 );
nand NAND2_12179 ( P2_U8103 , P2_U5584 , P2_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_12180 ( P2_U8104 , P2_U5641 , P2_U4394 );
nand NAND2_12181 ( P2_U8105 , P2_U5643 , P2_INSTQUEUEWR_ADDR_REG_3_ );
nand NAND2_12182 ( P2_U8106 , P2_U5651 , P2_U3533 );
nand NAND2_12183 ( P2_U8107 , P2_U8064 , P2_U4636 );
nand NAND2_12184 ( P2_U8108 , P2_U3579 , P2_U3319 );
nand NAND2_12185 ( P2_U8109 , P2_U8108 , P2_U8107 );
nand NAND2_12186 ( P2_U8110 , P2_U5643 , P2_INSTQUEUEWR_ADDR_REG_2_ );
nand NAND2_12187 ( P2_U8111 , P2_U5655 , P2_U3533 );
nand NAND2_12188 ( P2_U8112 , P2_U5643 , P2_INSTQUEUEWR_ADDR_REG_1_ );
nand NAND2_12189 ( P2_U8113 , P2_U5660 , P2_U3533 );
nand NAND2_12190 ( P2_U8114 , P2_U5643 , P2_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_12191 ( P2_U8115 , P2_U5664 , P2_U3533 );
nand NAND3_12192 ( P2_U8116 , P2_U2359 , P2_U3280 , P2_U2616 );
nand NAND2_12193 ( P2_U8117 , P2_U2438 , P2_U7873 );
nand NAND2_12194 ( P2_U8118 , P2_U8117 , P2_U8116 );
nand NAND3_12195 ( P2_U8119 , P2_U3253 , P2_U3278 , P2_U3297 );
nand NAND2_12196 ( P2_U8120 , P2_U8118 , P2_R2167_U6 );
nand NAND2_12197 ( P2_U8121 , P2_U7859 , P2_U7873 );
nand NAND2_12198 ( P2_U8122 , P2_U2616 , P2_U3282 );
nand NAND2_12199 ( P2_U8123 , P2_BYTEENABLE_REG_3_ , P2_U3547 );
nand NAND2_12200 ( P2_U8124 , P2_U3606 , P2_U4438 );
nand NAND2_12201 ( P2_U8125 , P2_BYTEENABLE_REG_2_ , P2_U3547 );
nand NAND2_12202 ( P2_U8126 , P2_U3607 , P2_U4438 );
nand NAND2_12203 ( P2_U8127 , P2_BYTEENABLE_REG_0_ , P2_U3547 );
nand NAND2_12204 ( P2_U8128 , P2_U4438 , P2_REIP_REG_0_ );
nand NAND2_12205 ( P2_U8129 , P2_U4439 , P2_U3552 );
nand NAND2_12206 ( P2_U8130 , P2_W_R_N_REG , P2_U3259 );
nand NAND2_12207 ( P2_U8131 , P2_U3287 , P2_U7873 );
nand NAND2_12208 ( P2_U8132 , P2_R2243_U8 , P2_U2616 );
nand NAND2_12209 ( P2_U8133 , P2_U6838 , P2_U3257 );
nand NAND2_12210 ( P2_U8134 , P2_MORE_REG , P2_U4400 );
nand NAND2_12211 ( P2_U8135 , P2_U7917 , P2_STATEBS16_REG );
nand NAND2_12212 ( P2_U8136 , BS16 , P2_U3589 );
nand NAND2_12213 ( P2_U8137 , P2_U6843 , P2_REQUESTPENDING_REG );
nand NAND2_12214 ( P2_U8138 , P2_U6852 , P2_U4402 );
nand NAND2_12215 ( P2_U8139 , P2_U4439 , P2_U3551 );
nand NAND2_12216 ( P2_U8140 , P2_D_C_N_REG , P2_U3259 );
nand NAND2_12217 ( P2_U8141 , P2_M_IO_N_REG , P2_U3259 );
nand NAND2_12218 ( P2_U8142 , P2_MEMORYFETCH_REG , P2_U4439 );
nand NAND2_12219 ( P2_U8143 , P2_U6857 , P2_READREQUEST_REG );
nand NAND2_12220 ( P2_U8144 , P2_U6858 , P2_U4403 );
nand NAND2_12221 ( P2_U8145 , P2_U7873 , P2_U3520 );
nand NAND2_12222 ( P2_U8146 , P2_U2616 , P2_U3297 );
nand NAND2_12223 ( P2_U8147 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U4405 );
nand NAND2_12224 ( P2_U8148 , P2_U7007 , P2_U3273 );
not NOT1_12225 ( P2_U8149 , P2_U3583 );
nand NAND2_12226 ( P2_U8150 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_U3273 );
nand NAND2_12227 ( P2_U8151 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_U3276 );
not NOT1_12228 ( P2_U8152 , P2_U3584 );
nand NAND2_12229 ( P2_U8153 , P2_U3584 , P2_U3327 );
nand NAND2_12230 ( P2_U8154 , P2_U8152 , P2_U3431 );
nand NAND2_12231 ( P2_U8155 , P2_U3584 , P2_U3368 );
nand NAND2_12232 ( P2_U8156 , P2_U8152 , P2_U3465 );
nand NAND2_12233 ( P2_U8157 , P2_U3584 , P2_U3357 );
nand NAND2_12234 ( P2_U8158 , P2_U8152 , P2_U3454 );
nand NAND2_12235 ( P2_U8159 , P2_U3584 , P2_U3416 );
nand NAND2_12236 ( P2_U8160 , P2_U8152 , P2_U3511 );
nand NAND2_12237 ( P2_U8161 , P2_U3584 , P2_U3382 );
nand NAND2_12238 ( P2_U8162 , P2_U8152 , P2_U3477 );
nand NAND2_12239 ( P2_U8163 , P2_U3584 , P2_U3405 );
nand NAND2_12240 ( P2_U8164 , P2_U8152 , P2_U3500 );
nand NAND2_12241 ( P2_U8165 , P2_U3584 , P2_U3393 );
nand NAND2_12242 ( P2_U8166 , P2_U8152 , P2_U3488 );
nand NAND2_12243 ( P2_U8167 , P2_U3584 , P2_U3341 );
nand NAND2_12244 ( P2_U8168 , P2_U8152 , P2_U3442 );
nand NAND2_12245 ( P2_U8169 , P2_U3584 , P2_U3328 );
nand NAND2_12246 ( P2_U8170 , P2_U8152 , P2_U3432 );
nand NAND2_12247 ( P2_U8171 , P2_U3584 , P2_U3369 );
nand NAND2_12248 ( P2_U8172 , P2_U8152 , P2_U3466 );
nand NAND2_12249 ( P2_U8173 , P2_U3584 , P2_U3358 );
nand NAND2_12250 ( P2_U8174 , P2_U8152 , P2_U3455 );
nand NAND2_12251 ( P2_U8175 , P2_U3584 , P2_U3417 );
nand NAND2_12252 ( P2_U8176 , P2_U8152 , P2_U3512 );
nand NAND2_12253 ( P2_U8177 , P2_U3584 , P2_U3383 );
nand NAND2_12254 ( P2_U8178 , P2_U8152 , P2_U3478 );
nand NAND2_12255 ( P2_U8179 , P2_U3584 , P2_U3406 );
nand NAND2_12256 ( P2_U8180 , P2_U8152 , P2_U3501 );
nand NAND2_12257 ( P2_U8181 , P2_U3584 , P2_U3394 );
nand NAND2_12258 ( P2_U8182 , P2_U8152 , P2_U3489 );
nand NAND2_12259 ( P2_U8183 , P2_U3584 , P2_U3342 );
nand NAND2_12260 ( P2_U8184 , P2_U8152 , P2_U3443 );
nand NAND2_12261 ( P2_U8185 , P2_U3584 , P2_U3329 );
nand NAND2_12262 ( P2_U8186 , P2_U8152 , P2_U3433 );
nand NAND2_12263 ( P2_U8187 , P2_U3584 , P2_U3370 );
nand NAND2_12264 ( P2_U8188 , P2_U8152 , P2_U3467 );
nand NAND2_12265 ( P2_U8189 , P2_U3584 , P2_U3359 );
nand NAND2_12266 ( P2_U8190 , P2_U8152 , P2_U3456 );
nand NAND2_12267 ( P2_U8191 , P2_U3584 , P2_U3418 );
nand NAND2_12268 ( P2_U8192 , P2_U8152 , P2_U3513 );
nand NAND2_12269 ( P2_U8193 , P2_U3584 , P2_U3384 );
nand NAND2_12270 ( P2_U8194 , P2_U8152 , P2_U3479 );
nand NAND2_12271 ( P2_U8195 , P2_U3584 , P2_U3407 );
nand NAND2_12272 ( P2_U8196 , P2_U8152 , P2_U3502 );
nand NAND2_12273 ( P2_U8197 , P2_U3584 , P2_U3395 );
nand NAND2_12274 ( P2_U8198 , P2_U8152 , P2_U3490 );
nand NAND2_12275 ( P2_U8199 , P2_U3584 , P2_U3343 );
nand NAND2_12276 ( P2_U8200 , P2_U8152 , P2_U3444 );
nand NAND2_12277 ( P2_U8201 , P2_U3584 , P2_U3330 );
nand NAND2_12278 ( P2_U8202 , P2_U8152 , P2_U3434 );
nand NAND2_12279 ( P2_U8203 , P2_U3584 , P2_U3371 );
nand NAND2_12280 ( P2_U8204 , P2_U8152 , P2_U3468 );
nand NAND2_12281 ( P2_U8205 , P2_U3584 , P2_U3360 );
nand NAND2_12282 ( P2_U8206 , P2_U8152 , P2_U3457 );
nand NAND2_12283 ( P2_U8207 , P2_U3584 , P2_U3419 );
nand NAND2_12284 ( P2_U8208 , P2_U8152 , P2_U3514 );
nand NAND2_12285 ( P2_U8209 , P2_U3584 , P2_U3385 );
nand NAND2_12286 ( P2_U8210 , P2_U8152 , P2_U3480 );
nand NAND2_12287 ( P2_U8211 , P2_U3584 , P2_U3408 );
nand NAND2_12288 ( P2_U8212 , P2_U8152 , P2_U3503 );
nand NAND2_12289 ( P2_U8213 , P2_U3584 , P2_U3396 );
nand NAND2_12290 ( P2_U8214 , P2_U8152 , P2_U3491 );
nand NAND2_12291 ( P2_U8215 , P2_U3584 , P2_U3344 );
nand NAND2_12292 ( P2_U8216 , P2_U8152 , P2_U3445 );
nand NAND2_12293 ( P2_U8217 , P2_U3584 , P2_U3331 );
nand NAND2_12294 ( P2_U8218 , P2_U8152 , P2_U3435 );
nand NAND2_12295 ( P2_U8219 , P2_U3584 , P2_U3372 );
nand NAND2_12296 ( P2_U8220 , P2_U8152 , P2_U3469 );
nand NAND2_12297 ( P2_U8221 , P2_U3584 , P2_U3361 );
nand NAND2_12298 ( P2_U8222 , P2_U8152 , P2_U3458 );
nand NAND2_12299 ( P2_U8223 , P2_U3584 , P2_U3420 );
nand NAND2_12300 ( P2_U8224 , P2_U8152 , P2_U3515 );
nand NAND2_12301 ( P2_U8225 , P2_U3584 , P2_U3386 );
nand NAND2_12302 ( P2_U8226 , P2_U8152 , P2_U3481 );
nand NAND2_12303 ( P2_U8227 , P2_U3584 , P2_U3409 );
nand NAND2_12304 ( P2_U8228 , P2_U8152 , P2_U3504 );
nand NAND2_12305 ( P2_U8229 , P2_U3584 , P2_U3397 );
nand NAND2_12306 ( P2_U8230 , P2_U8152 , P2_U3492 );
nand NAND2_12307 ( P2_U8231 , P2_U3584 , P2_U3345 );
nand NAND2_12308 ( P2_U8232 , P2_U8152 , P2_U3446 );
nand NAND2_12309 ( P2_U8233 , P2_U3584 , P2_U3332 );
nand NAND2_12310 ( P2_U8234 , P2_U8152 , P2_U3436 );
nand NAND2_12311 ( P2_U8235 , P2_U3584 , P2_U3373 );
nand NAND2_12312 ( P2_U8236 , P2_U8152 , P2_U3470 );
nand NAND2_12313 ( P2_U8237 , P2_U3584 , P2_U3362 );
nand NAND2_12314 ( P2_U8238 , P2_U8152 , P2_U3459 );
nand NAND2_12315 ( P2_U8239 , P2_U3584 , P2_U3421 );
nand NAND2_12316 ( P2_U8240 , P2_U8152 , P2_U3516 );
nand NAND2_12317 ( P2_U8241 , P2_U3584 , P2_U3387 );
nand NAND2_12318 ( P2_U8242 , P2_U8152 , P2_U3482 );
nand NAND2_12319 ( P2_U8243 , P2_U3584 , P2_U3410 );
nand NAND2_12320 ( P2_U8244 , P2_U8152 , P2_U3505 );
nand NAND2_12321 ( P2_U8245 , P2_U3584 , P2_U3398 );
nand NAND2_12322 ( P2_U8246 , P2_U8152 , P2_U3493 );
nand NAND2_12323 ( P2_U8247 , P2_U3584 , P2_U3346 );
nand NAND2_12324 ( P2_U8248 , P2_U8152 , P2_U3447 );
nand NAND2_12325 ( P2_U8249 , P2_U3584 , P2_U3333 );
nand NAND2_12326 ( P2_U8250 , P2_U8152 , P2_U3437 );
nand NAND2_12327 ( P2_U8251 , P2_U3584 , P2_U3374 );
nand NAND2_12328 ( P2_U8252 , P2_U8152 , P2_U3471 );
nand NAND2_12329 ( P2_U8253 , P2_U3584 , P2_U3363 );
nand NAND2_12330 ( P2_U8254 , P2_U8152 , P2_U3460 );
nand NAND2_12331 ( P2_U8255 , P2_U3584 , P2_U3422 );
nand NAND2_12332 ( P2_U8256 , P2_U8152 , P2_U3517 );
nand NAND2_12333 ( P2_U8257 , P2_U3584 , P2_U3388 );
nand NAND2_12334 ( P2_U8258 , P2_U8152 , P2_U3483 );
nand NAND2_12335 ( P2_U8259 , P2_U3584 , P2_U3411 );
nand NAND2_12336 ( P2_U8260 , P2_U8152 , P2_U3506 );
nand NAND2_12337 ( P2_U8261 , P2_U3584 , P2_U3399 );
nand NAND2_12338 ( P2_U8262 , P2_U8152 , P2_U3494 );
nand NAND2_12339 ( P2_U8263 , P2_U3584 , P2_U3347 );
nand NAND2_12340 ( P2_U8264 , P2_U8152 , P2_U3448 );
nand NAND2_12341 ( P2_U8265 , P2_U3584 , P2_U3334 );
nand NAND2_12342 ( P2_U8266 , P2_U8152 , P2_U3438 );
nand NAND2_12343 ( P2_U8267 , P2_U3584 , P2_U3375 );
nand NAND2_12344 ( P2_U8268 , P2_U8152 , P2_U3472 );
nand NAND2_12345 ( P2_U8269 , P2_U3584 , P2_U3364 );
nand NAND2_12346 ( P2_U8270 , P2_U8152 , P2_U3461 );
nand NAND2_12347 ( P2_U8271 , P2_U3584 , P2_U3423 );
nand NAND2_12348 ( P2_U8272 , P2_U8152 , P2_U3518 );
nand NAND2_12349 ( P2_U8273 , P2_U3584 , P2_U3389 );
nand NAND2_12350 ( P2_U8274 , P2_U8152 , P2_U3484 );
nand NAND2_12351 ( P2_U8275 , P2_U3584 , P2_U3412 );
nand NAND2_12352 ( P2_U8276 , P2_U8152 , P2_U3507 );
nand NAND2_12353 ( P2_U8277 , P2_U3584 , P2_U3400 );
nand NAND2_12354 ( P2_U8278 , P2_U8152 , P2_U3495 );
nand NAND2_12355 ( P2_U8279 , P2_U3584 , P2_U3348 );
nand NAND2_12356 ( P2_U8280 , P2_U8152 , P2_U3449 );
nand NAND2_12357 ( P2_U8281 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_U3519 );
nand NAND3_12358 ( P2_U8282 , P2_U3598 , P2_U3597 , P2_FLUSH_REG );
nand NAND2_12359 ( P2_U8283 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_U3519 );
nand NAND3_12360 ( P2_U8284 , P2_U3597 , P2_U8090 , P2_FLUSH_REG );
nand NAND2_12361 ( P2_U8285 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_U3519 );
nand NAND2_12362 ( P2_U8286 , P2_U8087 , P2_FLUSH_REG );
nand NAND2_12363 ( P2_U8287 , P2_U3616 , P2_U4406 );
nand NAND2_12364 ( P2_U8288 , P2_U5581 , P2_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_12365 ( P2_U8289 , P2_U5581 , P2_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_12366 ( P2_U8290 , P2_U5611 , P2_U4406 );
nand NAND2_12367 ( P2_U8291 , P2_U5581 , P2_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_12368 ( P2_U8292 , P2_U5619 , P2_U4406 );
nand NAND2_12369 ( P2_U8293 , P2_U5581 , P2_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_12370 ( P2_U8294 , P2_U5629 , P2_U4406 );
nand NAND2_12371 ( P2_U8295 , P2_U5581 , P2_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_12372 ( P2_U8296 , P2_U5637 , P2_U4406 );
nand NAND2_12373 ( P2_U8297 , P2_U3242 , P2_U7873 );
nand NAND2_12374 ( P2_U8298 , P2_U2616 , P2_U7183 );
nand NAND2_12375 ( P2_U8299 , P2_U7217 , P2_U7873 );
nand NAND2_12376 ( P2_U8300 , P2_U2616 , P2_U7200 );
nand NAND2_12377 ( P2_U8301 , P2_U7251 , P2_U7873 );
nand NAND2_12378 ( P2_U8302 , P2_U2616 , P2_U7234 );
nand NAND2_12379 ( P2_U8303 , P2_U7285 , P2_U7873 );
nand NAND2_12380 ( P2_U8304 , P2_U2616 , P2_U7268 );
nand NAND2_12381 ( P2_U8305 , P2_U7319 , P2_U7873 );
nand NAND2_12382 ( P2_U8306 , P2_U2616 , P2_U7302 );
nand NAND2_12383 ( P2_U8307 , P2_U7353 , P2_U7873 );
nand NAND2_12384 ( P2_U8308 , P2_U2616 , P2_U7336 );
nand NAND2_12385 ( P2_U8309 , P2_U7387 , P2_U7873 );
nand NAND2_12386 ( P2_U8310 , P2_U2616 , P2_U7370 );
nand NAND2_12387 ( P2_U8311 , P2_U7421 , P2_U7873 );
nand NAND2_12388 ( P2_U8312 , P2_U2616 , P2_U7404 );
nand NAND2_12389 ( P2_U8313 , P2_R2256_U5 , P2_U3572 );
nand NAND2_12390 ( P2_U8314 , P2_U3242 , P2_R2267_U56 );
nand NAND2_12391 ( P2_U8315 , P2_R2256_U17 , P2_U3572 );
nand NAND2_12392 ( P2_U8316 , P2_U3242 , P2_R2267_U19 );
nand NAND2_12393 ( P2_U8317 , P2_R2256_U18 , P2_U3572 );
nand NAND2_12394 ( P2_U8318 , P2_U3242 , P2_R2267_U58 );
nand NAND2_12395 ( P2_U8319 , P2_R2256_U19 , P2_U3572 );
nand NAND2_12396 ( P2_U8320 , P2_U3242 , P2_R2267_U18 );
nand NAND2_12397 ( P2_U8321 , P2_R2256_U20 , P2_U3572 );
nand NAND2_12398 ( P2_U8322 , P2_U3242 , P2_R2267_U60 );
nand NAND2_12399 ( P2_U8323 , P2_R2256_U26 , P2_U3572 );
nand NAND2_12400 ( P2_U8324 , P2_U3242 , P2_R2267_U17 );
nand NAND2_12401 ( P2_U8325 , P2_R2256_U22 , P2_U3572 );
nand NAND2_12402 ( P2_U8326 , P2_U3242 , P2_R2267_U65 );
nand NAND2_12403 ( P2_U8327 , P2_R2256_U4 , P2_U3572 );
nand NAND2_12404 ( P2_U8328 , P2_U3242 , P2_R2267_U43 );
nand NAND2_12405 ( P2_U8329 , P2_R2256_U21 , P2_U3572 );
nand NAND2_12406 ( P2_U8330 , P2_U3242 , P2_R2267_U21 );
nand NAND2_12407 ( P2_U8331 , P2_R2219_U24 , P2_U2617 );
nand NAND2_12408 ( P2_U8332 , P2_EBX_REG_7_ , P2_U7869 );
nand NAND2_12409 ( P2_U8333 , P2_R2219_U25 , P2_U2617 );
nand NAND2_12410 ( P2_U8334 , P2_EBX_REG_6_ , P2_U7869 );
nand NAND2_12411 ( P2_U8335 , P2_R2219_U26 , P2_U2617 );
nand NAND2_12412 ( P2_U8336 , P2_EBX_REG_5_ , P2_U7869 );
nand NAND2_12413 ( P2_U8337 , P2_R2219_U27 , P2_U2617 );
nand NAND2_12414 ( P2_U8338 , P2_EBX_REG_4_ , P2_U7869 );
nand NAND2_12415 ( P2_U8339 , P2_R2219_U28 , P2_U2617 );
nand NAND2_12416 ( P2_U8340 , P2_EBX_REG_3_ , P2_U7869 );
nand NAND2_12417 ( P2_U8341 , P2_R2219_U29 , P2_U2617 );
nand NAND2_12418 ( P2_U8342 , P2_EBX_REG_2_ , P2_U7869 );
nand NAND2_12419 ( P2_U8343 , P2_R2219_U30 , P2_U2617 );
nand NAND2_12420 ( P2_U8344 , P2_EBX_REG_1_ , P2_U7869 );
nand NAND2_12421 ( P2_U8345 , P2_R2219_U8 , P2_U2617 );
nand NAND2_12422 ( P2_U8346 , P2_EBX_REG_0_ , P2_U7869 );
nand NAND2_12423 ( P2_U8347 , P2_U3255 , P2_U7740 );
nand NAND2_12424 ( P2_U8348 , P2_U7867 , P2_U3525 );
nand NAND2_12425 ( P2_U8349 , P2_R2337_U68 , P2_U3284 );
nand NAND2_12426 ( P2_U8350 , P2_INSTADDRPOINTER_REG_31_ , P2_STATE2_REG_0_ );
nand NAND2_12427 ( P2_U8351 , P2_R2238_U6 , P2_U3283 );
nand NAND2_12428 ( P2_U8352 , P2_SUB_450_U6 , P2_U4417 );
nand NAND2_12429 ( P2_U8353 , P2_R2238_U19 , P2_U3283 );
nand NAND2_12430 ( P2_U8354 , P2_SUB_450_U17 , P2_U4417 );
nand NAND2_12431 ( P2_U8355 , P2_R2238_U20 , P2_U3283 );
nand NAND2_12432 ( P2_U8356 , P2_SUB_450_U18 , P2_U4417 );
nand NAND2_12433 ( P2_U8357 , P2_R2238_U21 , P2_U3283 );
nand NAND2_12434 ( P2_U8358 , P2_SUB_450_U19 , P2_U4417 );
nand NAND2_12435 ( P2_U8359 , P2_R2238_U22 , P2_U3283 );
nand NAND2_12436 ( P2_U8360 , P2_SUB_450_U20 , P2_U4417 );
nand NAND2_12437 ( P2_U8361 , P2_R2337_U61 , P2_U3284 );
nand NAND2_12438 ( P2_U8362 , P2_INSTADDRPOINTER_REG_9_ , P2_STATE2_REG_0_ );
nand NAND2_12439 ( P2_U8363 , P2_R2337_U62 , P2_U3284 );
nand NAND2_12440 ( P2_U8364 , P2_INSTADDRPOINTER_REG_8_ , P2_STATE2_REG_0_ );
nand NAND2_12441 ( P2_U8365 , P2_R2337_U63 , P2_U3284 );
nand NAND2_12442 ( P2_U8366 , P2_INSTADDRPOINTER_REG_7_ , P2_STATE2_REG_0_ );
nand NAND2_12443 ( P2_U8367 , P2_R2337_U64 , P2_U3284 );
nand NAND2_12444 ( P2_U8368 , P2_INSTADDRPOINTER_REG_6_ , P2_STATE2_REG_0_ );
nand NAND2_12445 ( P2_U8369 , P2_R2337_U65 , P2_U3284 );
nand NAND2_12446 ( P2_U8370 , P2_INSTADDRPOINTER_REG_5_ , P2_STATE2_REG_0_ );
nand NAND2_12447 ( P2_U8371 , P2_R2337_U66 , P2_U3284 );
nand NAND2_12448 ( P2_U8372 , P2_INSTADDRPOINTER_REG_4_ , P2_STATE2_REG_0_ );
nand NAND2_12449 ( P2_U8373 , P2_R2337_U69 , P2_U3284 );
nand NAND2_12450 ( P2_U8374 , P2_INSTADDRPOINTER_REG_30_ , P2_STATE2_REG_0_ );
nand NAND2_12451 ( P2_U8375 , P2_R2337_U67 , P2_U3284 );
nand NAND2_12452 ( P2_U8376 , P2_INSTADDRPOINTER_REG_3_ , P2_STATE2_REG_0_ );
nand NAND2_12453 ( P2_U8377 , P2_R2337_U71 , P2_U3284 );
nand NAND2_12454 ( P2_U8378 , P2_INSTADDRPOINTER_REG_29_ , P2_STATE2_REG_0_ );
nand NAND2_12455 ( P2_U8379 , P2_R2337_U72 , P2_U3284 );
nand NAND2_12456 ( P2_U8380 , P2_INSTADDRPOINTER_REG_28_ , P2_STATE2_REG_0_ );
nand NAND2_12457 ( P2_U8381 , P2_R2337_U73 , P2_U3284 );
nand NAND2_12458 ( P2_U8382 , P2_INSTADDRPOINTER_REG_27_ , P2_STATE2_REG_0_ );
nand NAND2_12459 ( P2_U8383 , P2_R2337_U74 , P2_U3284 );
nand NAND2_12460 ( P2_U8384 , P2_INSTADDRPOINTER_REG_26_ , P2_STATE2_REG_0_ );
nand NAND2_12461 ( P2_U8385 , P2_R2337_U75 , P2_U3284 );
nand NAND2_12462 ( P2_U8386 , P2_INSTADDRPOINTER_REG_25_ , P2_STATE2_REG_0_ );
nand NAND2_12463 ( P2_U8387 , P2_R2337_U76 , P2_U3284 );
nand NAND2_12464 ( P2_U8388 , P2_INSTADDRPOINTER_REG_24_ , P2_STATE2_REG_0_ );
nand NAND2_12465 ( P2_U8389 , P2_R2337_U77 , P2_U3284 );
nand NAND2_12466 ( P2_U8390 , P2_INSTADDRPOINTER_REG_23_ , P2_STATE2_REG_0_ );
nand NAND2_12467 ( P2_U8391 , P2_R2337_U78 , P2_U3284 );
nand NAND2_12468 ( P2_U8392 , P2_INSTADDRPOINTER_REG_22_ , P2_STATE2_REG_0_ );
nand NAND2_12469 ( P2_U8393 , P2_R2337_U79 , P2_U3284 );
nand NAND2_12470 ( P2_U8394 , P2_INSTADDRPOINTER_REG_21_ , P2_STATE2_REG_0_ );
nand NAND2_12471 ( P2_U8395 , P2_R2337_U80 , P2_U3284 );
nand NAND2_12472 ( P2_U8396 , P2_INSTADDRPOINTER_REG_20_ , P2_STATE2_REG_0_ );
nand NAND2_12473 ( P2_U8397 , P2_R2337_U70 , P2_U3284 );
nand NAND2_12474 ( P2_U8398 , P2_INSTADDRPOINTER_REG_2_ , P2_STATE2_REG_0_ );
nand NAND2_12475 ( P2_U8399 , P2_R2337_U81 , P2_U3284 );
nand NAND2_12476 ( P2_U8400 , P2_INSTADDRPOINTER_REG_19_ , P2_STATE2_REG_0_ );
nand NAND2_12477 ( P2_U8401 , P2_R2337_U82 , P2_U3284 );
nand NAND2_12478 ( P2_U8402 , P2_INSTADDRPOINTER_REG_18_ , P2_STATE2_REG_0_ );
nand NAND2_12479 ( P2_U8403 , P2_R2337_U83 , P2_U3284 );
nand NAND2_12480 ( P2_U8404 , P2_INSTADDRPOINTER_REG_17_ , P2_STATE2_REG_0_ );
nand NAND2_12481 ( P2_U8405 , P2_R2337_U84 , P2_U3284 );
nand NAND2_12482 ( P2_U8406 , P2_INSTADDRPOINTER_REG_16_ , P2_STATE2_REG_0_ );
nand NAND2_12483 ( P2_U8407 , P2_R2337_U85 , P2_U3284 );
nand NAND2_12484 ( P2_U8408 , P2_INSTADDRPOINTER_REG_15_ , P2_STATE2_REG_0_ );
nand NAND2_12485 ( P2_U8409 , P2_R2337_U86 , P2_U3284 );
nand NAND2_12486 ( P2_U8410 , P2_INSTADDRPOINTER_REG_14_ , P2_STATE2_REG_0_ );
nand NAND2_12487 ( P2_U8411 , P2_R2337_U87 , P2_U3284 );
nand NAND2_12488 ( P2_U8412 , P2_INSTADDRPOINTER_REG_13_ , P2_STATE2_REG_0_ );
nand NAND2_12489 ( P2_U8413 , P2_R2337_U88 , P2_U3284 );
nand NAND2_12490 ( P2_U8414 , P2_INSTADDRPOINTER_REG_12_ , P2_STATE2_REG_0_ );
nand NAND2_12491 ( P2_U8415 , P2_R2337_U89 , P2_U3284 );
nand NAND2_12492 ( P2_U8416 , P2_INSTADDRPOINTER_REG_11_ , P2_STATE2_REG_0_ );
nand NAND2_12493 ( P2_U8417 , P2_R2337_U90 , P2_U3284 );
nand NAND2_12494 ( P2_U8418 , P2_INSTADDRPOINTER_REG_10_ , P2_STATE2_REG_0_ );
nand NAND2_12495 ( P2_U8419 , P2_R2337_U4 , P2_U3284 );
nand NAND2_12496 ( P2_U8420 , P2_INSTADDRPOINTER_REG_1_ , P2_STATE2_REG_0_ );
nand NAND2_12497 ( P2_U8421 , P2_PHYADDRPOINTER_REG_0_ , P2_U3284 );
nand NAND2_12498 ( P2_U8422 , P2_INSTADDRPOINTER_REG_0_ , P2_STATE2_REG_0_ );
nand NAND2_12499 ( P2_U8423 , P2_R2238_U6 , P2_U3269 );
nand NAND2_12500 ( P2_U8424 , P2_U2615 , P2_STATE2_REG_1_ );
nand NAND2_12501 ( P2_U8425 , P2_R2238_U19 , P2_U3269 );
nand NAND2_12502 ( P2_U8426 , P2_U2615 , P2_STATE2_REG_1_ );
nand NAND2_12503 ( P2_U8427 , P2_R2238_U20 , P2_U3269 );
nand NAND2_12504 ( P2_U8428 , P2_SUB_589_U8 , P2_STATE2_REG_1_ );
nand NAND2_12505 ( P2_U8429 , P2_R2238_U21 , P2_U3269 );
nand NAND2_12506 ( P2_U8430 , P2_SUB_589_U9 , P2_STATE2_REG_1_ );
nand NAND2_12507 ( P2_U8431 , P2_R2238_U22 , P2_U3269 );
nand NAND2_12508 ( P2_U8432 , P2_SUB_589_U6 , P2_STATE2_REG_1_ );
nand NAND2_12509 ( P2_U8433 , P2_R2238_U7 , P2_U3269 );
nand NAND2_12510 ( P2_U8434 , P2_SUB_589_U7 , P2_STATE2_REG_1_ );
nand NAND2_12511 ( P1_ADD_405_U171 , P1_INSTADDRPOINTER_REG_3_ , P1_ADD_405_U94 );
nand NAND2_12512 ( P1_ADD_405_U170 , P1_ADD_405_U126 , P1_ADD_405_U92 );
nand NAND2_12513 ( P1_ADD_405_U169 , P1_INSTADDRPOINTER_REG_31_ , P1_ADD_405_U93 );
nand NAND2_12514 ( P1_ADD_405_U168 , P1_ADD_405_U104 , P1_ADD_405_U21 );
nand NAND2_12515 ( P1_ADD_405_U167 , P1_INSTADDRPOINTER_REG_10_ , P1_ADD_405_U20 );
nand NAND2_12516 ( P1_ADD_405_U166 , P1_ADD_405_U113 , P1_ADD_405_U39 );
nand NAND2_12517 ( P1_ADD_405_U165 , P1_INSTADDRPOINTER_REG_19_ , P1_ADD_405_U38 );
nand NAND2_12518 ( P1_ADD_405_U164 , P1_ADD_405_U117 , P1_ADD_405_U47 );
nand NAND2_12519 ( P1_ADD_405_U163 , P1_INSTADDRPOINTER_REG_23_ , P1_ADD_405_U46 );
nand NAND2_12520 ( P1_ADD_405_U162 , P1_ADD_405_U102 , P1_ADD_405_U17 );
nand NAND2_12521 ( P1_ADD_405_U161 , P1_INSTADDRPOINTER_REG_8_ , P1_ADD_405_U16 );
nand NAND2_12522 ( P1_ADD_405_U160 , P1_ADD_405_U99 , P1_ADD_405_U11 );
nand NAND2_12523 ( P1_ADD_405_U159 , P1_INSTADDRPOINTER_REG_5_ , P1_ADD_405_U10 );
nand NAND2_12524 ( P1_ADD_405_U158 , P1_ADD_405_U108 , P1_ADD_405_U29 );
nand NAND2_12525 ( P1_ADD_405_U157 , P1_INSTADDRPOINTER_REG_14_ , P1_ADD_405_U28 );
nand NAND2_12526 ( P1_ADD_405_U156 , P1_ADD_405_U121 , P1_ADD_405_U55 );
nand NAND2_12527 ( P1_ADD_405_U155 , P1_INSTADDRPOINTER_REG_27_ , P1_ADD_405_U54 );
nand NAND2_12528 ( P1_ADD_405_U154 , P1_ADD_405_U98 , P1_ADD_405_U9 );
nand NAND2_12529 ( P1_ADD_405_U153 , P1_INSTADDRPOINTER_REG_4_ , P1_ADD_405_U8 );
nand NAND2_12530 ( P1_ADD_405_U152 , P1_ADD_405_U109 , P1_ADD_405_U31 );
nand NAND2_12531 ( P1_ADD_405_U151 , P1_INSTADDRPOINTER_REG_15_ , P1_ADD_405_U30 );
nand NAND2_12532 ( P1_ADD_405_U150 , P1_ADD_405_U120 , P1_ADD_405_U53 );
nand NAND2_12533 ( P1_ADD_405_U149 , P1_INSTADDRPOINTER_REG_26_ , P1_ADD_405_U52 );
nand NAND2_12534 ( P1_ADD_405_U148 , P1_ADD_405_U105 , P1_ADD_405_U23 );
nand NAND2_12535 ( P1_ADD_405_U147 , P1_INSTADDRPOINTER_REG_11_ , P1_ADD_405_U22 );
nand NAND2_12536 ( P1_ADD_405_U146 , P1_ADD_405_U112 , P1_ADD_405_U37 );
nand NAND2_12537 ( P1_ADD_405_U145 , P1_INSTADDRPOINTER_REG_18_ , P1_ADD_405_U36 );
nand NAND2_12538 ( P1_ADD_405_U144 , P1_ADD_405_U116 , P1_ADD_405_U45 );
nand NAND2_12539 ( P1_ADD_405_U143 , P1_INSTADDRPOINTER_REG_22_ , P1_ADD_405_U44 );
nand NAND2_12540 ( P1_ADD_405_U142 , P1_ADD_405_U103 , P1_ADD_405_U19 );
nand NAND2_12541 ( P1_ADD_405_U141 , P1_INSTADDRPOINTER_REG_9_ , P1_ADD_405_U18 );
nand NAND2_12542 ( P1_ADD_405_U140 , P1_ADD_405_U107 , P1_ADD_405_U27 );
nand NAND2_12543 ( P1_ADD_405_U139 , P1_INSTADDRPOINTER_REG_13_ , P1_ADD_405_U26 );
nand NAND2_12544 ( P1_ADD_405_U138 , P1_ADD_405_U114 , P1_ADD_405_U41 );
nand NAND2_12545 ( P1_ADD_405_U137 , P1_INSTADDRPOINTER_REG_20_ , P1_ADD_405_U40 );
nand NAND2_12546 ( P1_ADD_405_U136 , P1_ADD_405_U111 , P1_ADD_405_U35 );
nand NAND2_12547 ( P1_ADD_405_U135 , P1_INSTADDRPOINTER_REG_17_ , P1_ADD_405_U34 );
nand NAND2_12548 ( P1_ADD_405_U134 , P1_ADD_405_U118 , P1_ADD_405_U49 );
nand NAND2_12549 ( P1_ADD_405_U133 , P1_INSTADDRPOINTER_REG_24_ , P1_ADD_405_U48 );
nand NAND2_12550 ( P1_ADD_405_U132 , P1_ADD_405_U123 , P1_ADD_405_U59 );
nand NAND2_12551 ( P1_ADD_405_U131 , P1_INSTADDRPOINTER_REG_29_ , P1_ADD_405_U58 );
nand NAND2_12552 ( P1_ADD_405_U130 , P1_ADD_405_U124 , P1_ADD_405_U60 );
nand NAND2_12553 ( P1_ADD_405_U129 , P1_INSTADDRPOINTER_REG_30_ , P1_ADD_405_U61 );
nand NAND2_12554 ( P1_ADD_405_U128 , P1_ADD_405_U100 , P1_ADD_405_U12 );
nand NAND2_12555 ( P1_ADD_405_U127 , P1_INSTADDRPOINTER_REG_6_ , P1_ADD_405_U13 );
not NOT1_12556 ( P1_ADD_405_U126 , P1_ADD_405_U93 );
nand NAND3_12557 ( P1_ADD_405_U125 , P1_INSTADDRPOINTER_REG_1_ , P1_INSTADDRPOINTER_REG_0_ , P1_INSTADDRPOINTER_REG_2_ );
not NOT1_12558 ( P1_ADD_405_U124 , P1_ADD_405_U61 );
not NOT1_12559 ( P1_ADD_405_U123 , P1_ADD_405_U58 );
not NOT1_12560 ( P1_ADD_405_U122 , P1_ADD_405_U56 );
not NOT1_12561 ( P1_ADD_405_U121 , P1_ADD_405_U54 );
not NOT1_12562 ( P1_ADD_405_U120 , P1_ADD_405_U52 );
not NOT1_12563 ( P1_ADD_405_U119 , P1_ADD_405_U50 );
not NOT1_12564 ( P1_ADD_405_U118 , P1_ADD_405_U48 );
not NOT1_12565 ( P1_ADD_405_U117 , P1_ADD_405_U46 );
not NOT1_12566 ( P1_ADD_405_U116 , P1_ADD_405_U44 );
not NOT1_12567 ( P1_ADD_405_U115 , P1_ADD_405_U42 );
nor nor_12568 ( P1_U2352 , P1_STATEBS16_REG , P1_STATE2_REG_2_ );
and AND2_12569 ( P1_U2353 , P1_U4231 , P1_STATE2_REG_2_ );
and AND2_12570 ( P1_U2354 , P1_U4265 , P1_U4477 );
and AND2_12571 ( P1_U2355 , P1_U3234 , P1_U2450 );
and AND2_12572 ( P1_U2356 , P1_R2238_U6 , P1_U4192 );
and AND3_12573 ( P1_U2357 , P1_U5959 , P1_U3865 , P1_R2167_U17 );
and AND2_12574 ( P1_U2358 , P1_U2388 , P1_U4224 );
and AND2_12575 ( P1_U2359 , P1_STATE2_REG_2_ , P1_U3431 );
and AND2_12576 ( P1_U2360 , P1_STATE2_REG_2_ , P1_U3414 );
and AND2_12577 ( P1_U2361 , P1_U4224 , P1_STATE2_REG_3_ );
and AND2_12578 ( P1_U2362 , P1_U2359 , P1_U4208 );
and AND2_12579 ( P1_U2363 , P1_U2359 , P1_U4210 );
and AND2_12580 ( P1_U2364 , P1_U3864 , P1_U3416 );
and AND2_12581 ( P1_U2365 , P1_U4261 , P1_U3416 );
and AND3_12582 ( P1_U2366 , P1_U3431 , P1_STATE2_REG_1_ , P1_U3430 );
and AND3_12583 ( P1_U2367 , P1_STATE2_REG_1_ , P1_U3431 , P1_R2337_U69 );
and AND2_12584 ( P1_U2368 , P1_U4235 , P1_STATE2_REG_0_ );
and AND2_12585 ( P1_U2369 , P1_U2362 , P1_U4497 );
and AND2_12586 ( P1_U2370 , P1_U3414 , P1_U3263 );
and AND2_12587 ( P1_U2371 , P1_U4222 , P1_U4449 );
and AND2_12588 ( P1_U2372 , P1_STATE2_REG_0_ , P1_U3416 );
and AND2_12589 ( P1_U2373 , P1_STATE2_REG_3_ , P1_U3431 );
and AND2_12590 ( P1_U2374 , P1_U2360 , P1_U4214 );
and AND2_12591 ( P1_U2375 , P1_U2360 , P1_U4216 );
and AND2_12592 ( P1_U2376 , P1_U5798 , P1_U3416 );
and AND2_12593 ( P1_U2377 , P1_U3762 , P1_U3414 );
and AND2_12594 ( P1_U2378 , P1_U2360 , P1_U5569 );
and AND2_12595 ( P1_U2379 , P1_U2363 , P1_U3280 );
and AND2_12596 ( P1_U2380 , P1_U2360 , P1_U7608 );
and AND2_12597 ( P1_U2381 , P1_U2357 , P1_U3271 );
and AND2_12598 ( P1_U2382 , P1_U2357 , P1_U4477 );
and AND2_12599 ( P1_U2383 , P1_U4222 , P1_U3391 );
and AND2_12600 ( P1_U2384 , P1_STATE2_REG_0_ , P1_U3417 );
and AND2_12601 ( P1_U2385 , P1_U3417 , P1_U3294 );
and AND2_12602 ( P1_U2386 , P1_U4223 , P1_U3423 );
and AND2_12603 ( P1_U2387 , P1_U3884 , P1_U4223 );
and AND2_12604 ( P1_U2388 , P1_STATEBS16_REG , P1_U4209 );
and AND2_12605 ( P1_U2389 , P1_U2452 , P1_U7494 );
and AND2_12606 ( P1_U2390 , U346 , P1_U4224 );
and AND2_12607 ( P1_U2391 , U335 , P1_U4224 );
and AND2_12608 ( P1_U2392 , U324 , P1_U4224 );
and AND2_12609 ( P1_U2393 , U321 , P1_U4224 );
and AND2_12610 ( P1_U2394 , U320 , P1_U4224 );
and AND2_12611 ( P1_U2395 , U319 , P1_U4224 );
and AND2_12612 ( P1_U2396 , U318 , P1_U4224 );
and AND2_12613 ( P1_U2397 , U317 , P1_U4224 );
and AND2_12614 ( P1_U2398 , U330 , P1_U2358 );
and AND2_12615 ( P1_U2399 , U339 , P1_U2358 );
and AND2_12616 ( P1_U2400 , U329 , P1_U2358 );
and AND2_12617 ( P1_U2401 , U338 , P1_U2358 );
and AND2_12618 ( P1_U2402 , U328 , P1_U2358 );
and AND2_12619 ( P1_U2403 , U337 , P1_U2358 );
and AND2_12620 ( P1_U2404 , U327 , P1_U2358 );
and AND2_12621 ( P1_U2405 , U336 , P1_U2358 );
and AND2_12622 ( P1_U2406 , U326 , P1_U2358 );
and AND2_12623 ( P1_U2407 , U334 , P1_U2358 );
and AND2_12624 ( P1_U2408 , U325 , P1_U2358 );
and AND2_12625 ( P1_U2409 , U333 , P1_U2358 );
and AND2_12626 ( P1_U2410 , U323 , P1_U2358 );
and AND2_12627 ( P1_U2411 , U332 , P1_U2358 );
and AND2_12628 ( P1_U2412 , U322 , P1_U2358 );
and AND2_12629 ( P1_U2413 , U331 , P1_U2358 );
and AND2_12630 ( P1_U2414 , P1_U2361 , P1_U3271 );
and AND2_12631 ( P1_U2415 , P1_U2361 , P1_U3391 );
and AND2_12632 ( P1_U2416 , P1_U2361 , P1_U3277 );
and AND2_12633 ( P1_U2417 , P1_U2361 , P1_U3284 );
and AND2_12634 ( P1_U2418 , P1_U2361 , P1_U3283 );
and AND2_12635 ( P1_U2419 , P1_U2361 , P1_U3278 );
and AND2_12636 ( P1_U2420 , P1_U2361 , P1_U4173 );
and AND2_12637 ( P1_U2421 , P1_U2361 , P1_U4171 );
and AND2_12638 ( P1_U2422 , P1_U4223 , P1_U5461 );
and AND2_12639 ( P1_U2423 , P1_U4223 , P1_U4231 );
and AND2_12640 ( P1_U2424 , P1_U2384 , P1_U3284 );
and AND2_12641 ( P1_U2425 , P1_U2368 , P1_U2448 );
and AND2_12642 ( P1_U2426 , P1_U3889 , P1_U3431 );
nor nor_12643 ( P1_U2427 , P1_STATE2_REG_1_ , P1_STATE2_REG_3_ );
and AND2_12644 ( P1_U2428 , P1_STATE2_REG_2_ , P1_STATE2_REG_1_ );
and AND2_12645 ( P1_U2429 , P1_U6366 , P1_U3431 );
and AND2_12646 ( P1_U2430 , P1_STATE2_REG_1_ , P1_U3387 );
and AND2_12647 ( P1_U2431 , P1_U4199 , P1_U7494 );
and AND2_12648 ( P1_U2432 , P1_U3455 , P1_U3360 );
and AND2_12649 ( P1_U2433 , P1_U4540 , P1_U3455 );
and AND2_12650 ( P1_U2434 , P1_U7696 , P1_U3360 );
and AND2_12651 ( P1_U2435 , P1_U4540 , P1_U7696 );
and AND2_12652 ( P1_U2436 , P1_U3235 , P1_U3301 );
and AND2_12653 ( P1_U2437 , P1_U4543 , P1_U3301 );
and AND2_12654 ( P1_U2438 , P1_R2182_U42 , P1_R2182_U25 );
and AND2_12655 ( P1_U2439 , P1_R2182_U42 , P1_U3316 );
and AND2_12656 ( P1_U2440 , P1_R2182_U25 , P1_U3317 );
nor nor_12657 ( P1_U2441 , P1_R2182_U42 , P1_R2182_U25 );
and AND2_12658 ( P1_U2442 , P1_R2182_U33 , P1_R2182_U34 );
and AND2_12659 ( P1_U2443 , P1_R2182_U33 , P1_U3318 );
and AND2_12660 ( P1_U2444 , P1_R2182_U34 , P1_U3319 );
nor nor_12661 ( P1_U2445 , P1_R2182_U33 , P1_R2182_U34 );
and AND2_12662 ( P1_U2446 , P1_STATE2_REG_1_ , P1_U3471 );
and AND2_12663 ( P1_U2447 , P1_U3577 , P1_U2452 );
and AND2_12664 ( P1_U2448 , P1_R2167_U17 , P1_U3284 );
and AND2_12665 ( P1_U2449 , P1_U4494 , P1_U3271 );
and AND2_12666 ( P1_U2450 , P1_STATE2_REG_0_ , P1_U4400 );
and AND2_12667 ( P1_U2451 , P1_U4251 , P1_STATE2_REG_0_ );
and AND4_12668 ( P1_U2452 , P1_U4400 , P1_U3277 , P1_U3391 , P1_U4173 );
and AND4_12669 ( P1_U2453 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_12670 ( P1_U2454 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3266 );
and AND4_12671 ( P1_U2455 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3266 );
and AND2_12672 ( P1_U2456 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_U3265 );
and AND4_12673 ( P1_U2457 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3265 );
and AND2_12674 ( P1_U2458 , P1_U3507 , P1_U4378 );
and AND4_12675 ( P1_U2459 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3264 );
and AND3_12676 ( P1_U2460 , P1_U3264 , P1_U3266 , P1_INSTQUEUERD_ADDR_REG_1_ );
and AND2_12677 ( P1_U2461 , P1_U3506 , P1_U3505 );
and AND3_12678 ( P1_U2462 , P1_U3264 , P1_U3265 , P1_INSTQUEUERD_ADDR_REG_0_ );
and AND2_12679 ( P1_U2463 , P1_U3504 , P1_U3503 );
and AND2_12680 ( P1_U2464 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_U4380 );
and AND2_12681 ( P1_U2465 , P1_U3502 , P1_U3501 );
and AND2_12682 ( P1_U2466 , P1_U3500 , P1_U3499 );
and AND3_12683 ( P1_U2467 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3270 , P1_U4378 );
and AND2_12684 ( P1_U2468 , P1_U3498 , P1_U3497 );
nor nor_12685 ( P1_U2469 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND3_12686 ( P1_U2470 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3266 , P1_U2469 );
and AND3_12687 ( P1_U2471 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_U3265 , P1_U2469 );
and AND2_12688 ( P1_U2472 , P1_U4380 , P1_U3270 );
and AND3_12689 ( P1_U2473 , P1_U7680 , P1_U7679 , P1_U3406 );
and AND2_12690 ( P1_U2474 , P1_R2144_U49 , P1_U3312 );
and AND2_12691 ( P1_U2475 , P1_U3454 , P1_U3358 );
and AND2_12692 ( P1_U2476 , P1_R2144_U8 , P1_R2144_U49 );
and AND2_12693 ( P1_U2477 , P1_U4528 , P1_U2476 );
and AND2_12694 ( P1_U2478 , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_INSTQUEUEWR_ADDR_REG_3_ );
and AND2_12695 ( P1_U2479 , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_U3303 );
and AND2_12696 ( P1_U2480 , P1_U3315 , P1_U4548 );
and AND2_12697 ( P1_U2481 , P1_U4524 , P1_U2476 );
and AND2_12698 ( P1_U2482 , P1_U3327 , P1_U4606 );
and AND2_12699 ( P1_U2483 , P1_U4525 , P1_U2476 );
and AND2_12700 ( P1_U2484 , P1_U3334 , P1_U4665 );
and AND2_12701 ( P1_U2485 , P1_U4526 , P1_R2144_U43 );
nor nor_12702 ( P1_U2486 , P1_R2144_U43 , P1_R2144_U50 );
and AND2_12703 ( P1_U2487 , P1_U2486 , P1_U2476 );
nor nor_12704 ( P1_U2488 , P1_INSTQUEUEWR_ADDR_REG_0_ , P1_INSTQUEUEWR_ADDR_REG_1_ );
and AND2_12705 ( P1_U2489 , P1_U3338 , P1_U4722 );
and AND2_12706 ( P1_U2490 , P1_U7693 , P1_U3358 );
and AND2_12707 ( P1_U2491 , P1_U4529 , P1_U4528 );
and AND2_12708 ( P1_U2492 , P1_U3343 , P1_U4780 );
and AND2_12709 ( P1_U2493 , P1_U4529 , P1_U4524 );
and AND2_12710 ( P1_U2494 , P1_U3347 , P1_U4837 );
and AND2_12711 ( P1_U2495 , P1_U4529 , P1_U4525 );
and AND2_12712 ( P1_U2496 , P1_U3350 , P1_U4895 );
and AND2_12713 ( P1_U2497 , P1_U4529 , P1_U2486 );
and AND2_12714 ( P1_U2498 , P1_U3354 , P1_U4952 );
and AND2_12715 ( P1_U2499 , P1_U4531 , P1_U3454 );
and AND2_12716 ( P1_U2500 , P1_U3359 , P1_U3357 );
and AND2_12717 ( P1_U2501 , P1_U4524 , P1_U2474 );
and AND2_12718 ( P1_U2502 , P1_U3364 , P1_U5065 );
and AND2_12719 ( P1_U2503 , P1_U4525 , P1_U2474 );
and AND2_12720 ( P1_U2504 , P1_U3367 , P1_U5123 );
and AND2_12721 ( P1_U2505 , P1_U2486 , P1_U2474 );
and AND2_12722 ( P1_U2506 , P1_U3371 , P1_U5180 );
and AND2_12723 ( P1_U2507 , P1_U4531 , P1_U7693 );
nor nor_12724 ( P1_U2508 , P1_R2144_U49 , P1_R2144_U8 );
and AND2_12725 ( P1_U2509 , P1_U2508 , P1_U4528 );
nor nor_12726 ( P1_U2510 , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_INSTQUEUEWR_ADDR_REG_2_ );
and AND2_12727 ( P1_U2511 , P1_U3374 , P1_U5238 );
and AND2_12728 ( P1_U2512 , P1_U2508 , P1_U4524 );
and AND2_12729 ( P1_U2513 , P1_U3378 , P1_U5295 );
and AND2_12730 ( P1_U2514 , P1_U2508 , P1_U4525 );
and AND2_12731 ( P1_U2515 , P1_U3381 , P1_U5353 );
and AND2_12732 ( P1_U2516 , P1_U2508 , P1_U2486 );
and AND2_12733 ( P1_U2517 , P1_U3385 , P1_U5410 );
and AND3_12734 ( P1_U2518 , P1_U7700 , P1_U7699 , P1_U5468 );
and AND2_12735 ( P1_U2519 , P1_U3744 , P1_U5499 );
and AND2_12736 ( P1_U2520 , P1_U4219 , P1_U3446 );
and AND2_12737 ( P1_U2521 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_U3402 );
and AND2_12738 ( P1_U2522 , P1_U5483 , P1_U5511 );
and AND2_12739 ( P1_U2523 , P1_U2522 , P1_U2521 );
and AND2_12740 ( P1_U2524 , P1_U3266 , P1_U3402 );
and AND2_12741 ( P1_U2525 , P1_U2522 , P1_U2524 );
and AND2_12742 ( P1_U2526 , P1_U5519 , P1_INSTQUEUERD_ADDR_REG_0_ );
and AND2_12743 ( P1_U2527 , P1_U2522 , P1_U2526 );
and AND2_12744 ( P1_U2528 , P1_U5519 , P1_U3266 );
and AND2_12745 ( P1_U2529 , P1_U2522 , P1_U2528 );
and AND2_12746 ( P1_U2530 , P1_U5483 , P1_U3401 );
and AND2_12747 ( P1_U2531 , P1_U2530 , P1_U2521 );
and AND2_12748 ( P1_U2532 , P1_U2530 , P1_U2524 );
and AND2_12749 ( P1_U2533 , P1_U2530 , P1_U2526 );
and AND2_12750 ( P1_U2534 , P1_U2530 , P1_U2528 );
and AND2_12751 ( P1_U2535 , P1_U5511 , P1_U3438 );
and AND2_12752 ( P1_U2536 , P1_U2535 , P1_U2521 );
and AND2_12753 ( P1_U2537 , P1_U2535 , P1_U2524 );
and AND2_12754 ( P1_U2538 , P1_U2535 , P1_U2526 );
and AND2_12755 ( P1_U2539 , P1_U2535 , P1_U2528 );
and AND2_12756 ( P1_U2540 , P1_U3438 , P1_U3401 );
and AND2_12757 ( P1_U2541 , P1_U2521 , P1_U2540 );
and AND2_12758 ( P1_U2542 , P1_U2524 , P1_U2540 );
and AND2_12759 ( P1_U2543 , P1_U2526 , P1_U2540 );
and AND2_12760 ( P1_U2544 , P1_U2528 , P1_U2540 );
and AND2_12761 ( P1_U2545 , P1_U5480 , P1_U7720 );
and AND2_12762 ( P1_U2546 , P1_U2545 , P1_U2454 );
and AND2_12763 ( P1_U2547 , P1_U2545 , P1_U3498 );
and AND2_12764 ( P1_U2548 , P1_U2545 , P1_U4378 );
and AND2_12765 ( P1_U2549 , P1_U2545 , P1_U2456 );
and AND2_12766 ( P1_U2550 , P1_U5480 , P1_U3456 );
and AND2_12767 ( P1_U2551 , P1_U2550 , P1_U2454 );
and AND2_12768 ( P1_U2552 , P1_U2550 , P1_U3498 );
and AND2_12769 ( P1_U2553 , P1_U2550 , P1_U4378 );
and AND2_12770 ( P1_U2554 , P1_U2550 , P1_U2456 );
and AND2_12771 ( P1_U2555 , P1_U7720 , P1_U3442 );
and AND2_12772 ( P1_U2556 , P1_U2555 , P1_U2454 );
and AND2_12773 ( P1_U2557 , P1_U2555 , P1_U3498 );
and AND2_12774 ( P1_U2558 , P1_U2555 , P1_U4378 );
and AND2_12775 ( P1_U2559 , P1_U2555 , P1_U2456 );
and AND2_12776 ( P1_U2560 , P1_U3456 , P1_U3442 );
and AND2_12777 ( P1_U2561 , P1_U2560 , P1_U2454 );
and AND2_12778 ( P1_U2562 , P1_U2560 , P1_U3498 );
and AND2_12779 ( P1_U2563 , P1_U2560 , P1_U4378 );
and AND2_12780 ( P1_U2564 , P1_U2560 , P1_U2456 );
and AND2_12781 ( P1_U2565 , P1_U7065 , P1_U4379 );
and AND2_12782 ( P1_U2566 , P1_U7065 , P1_U2460 );
and AND2_12783 ( P1_U2567 , P1_U7065 , P1_U2462 );
and AND2_12784 ( P1_U2568 , P1_U7065 , P1_U4380 );
and AND2_12785 ( P1_U2569 , P1_U7065 , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_12786 ( P1_U2570 , P1_U2569 , P1_U3498 );
and AND2_12787 ( P1_U2571 , P1_U2569 , P1_U2454 );
and AND2_12788 ( P1_U2572 , P1_U2569 , P1_U2456 );
and AND2_12789 ( P1_U2573 , P1_U2569 , P1_U4378 );
and AND2_12790 ( P1_U2574 , P1_U4379 , P1_U3445 );
and AND2_12791 ( P1_U2575 , P1_U2460 , P1_U3445 );
and AND2_12792 ( P1_U2576 , P1_U2462 , P1_U3445 );
and AND2_12793 ( P1_U2577 , P1_U4380 , P1_U3445 );
and AND2_12794 ( P1_U2578 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3445 );
and AND2_12795 ( P1_U2579 , P1_U2578 , P1_U3498 );
and AND2_12796 ( P1_U2580 , P1_U2578 , P1_U2454 );
and AND2_12797 ( P1_U2581 , P1_U2578 , P1_U2456 );
and AND2_12798 ( P1_U2582 , P1_U2578 , P1_U4378 );
and AND2_12799 ( P1_U2583 , P1_U7790 , P1_U4184 );
and AND2_12800 ( P1_U2584 , P1_U2583 , P1_U2524 );
and AND2_12801 ( P1_U2585 , P1_U2583 , P1_U2521 );
and AND2_12802 ( P1_U2586 , P1_U2583 , P1_U2528 );
and AND2_12803 ( P1_U2587 , P1_U2583 , P1_U2526 );
and AND2_12804 ( P1_U2588 , P1_U7790 , P1_U3452 );
and AND2_12805 ( P1_U2589 , P1_U2588 , P1_U2524 );
and AND2_12806 ( P1_U2590 , P1_U2588 , P1_U2521 );
and AND2_12807 ( P1_U2591 , P1_U2588 , P1_U2528 );
and AND2_12808 ( P1_U2592 , P1_U2588 , P1_U2526 );
and AND2_12809 ( P1_U2593 , P1_U4184 , P1_U3457 );
and AND2_12810 ( P1_U2594 , P1_U2593 , P1_U2524 );
and AND2_12811 ( P1_U2595 , P1_U2593 , P1_U2521 );
and AND2_12812 ( P1_U2596 , P1_U2593 , P1_U2528 );
and AND2_12813 ( P1_U2597 , P1_U2593 , P1_U2526 );
and AND2_12814 ( P1_U2598 , P1_U3457 , P1_U3452 );
and AND2_12815 ( P1_U2599 , P1_U2598 , P1_U2524 );
and AND2_12816 ( P1_U2600 , P1_U2598 , P1_U2521 );
and AND2_12817 ( P1_U2601 , P1_U2598 , P1_U2528 );
and AND2_12818 ( P1_U2602 , P1_U2598 , P1_U2526 );
and AND2_12819 ( P1_U2603 , P1_STATE2_REG_0_ , P1_U3389 );
and AND2_12820 ( P1_U2604 , P1_EBX_REG_31_ , P1_U2379 );
and AND5_12821 ( P1_U2605 , P1_U3533 , P1_U2607 , P1_U3532 , P1_U3531 , P1_U3530 );
and AND2_12822 ( P1_U2606 , P1_U7504 , P1_U3427 );
and AND2_12823 ( P1_U2607 , P1_U7672 , P1_U7671 );
and AND2_12824 ( P1_U2608 , P1_U7787 , P1_U7786 );
nand NAND3_12825 ( P1_U2609 , P1_U6853 , P1_U6854 , P1_U6855 );
nand NAND2_12826 ( P1_U2610 , P1_U6856 , P1_U4026 );
nand NAND3_12827 ( P1_U2611 , P1_U6841 , P1_U6842 , P1_U6843 );
nand NAND3_12828 ( P1_U2612 , P1_U6844 , P1_U6845 , P1_U6846 );
nand NAND3_12829 ( P1_U2613 , P1_U6847 , P1_U6848 , P1_U6849 );
nand NAND2_12830 ( P1_U2614 , P1_U6756 , P1_U4005 );
nand NAND2_12831 ( P1_U2615 , P1_U6753 , P1_U4004 );
nand NAND3_12832 ( P1_U2616 , P1_U6850 , P1_U6851 , P1_U6852 );
nand NAND2_12833 ( P1_U2617 , P1_U6750 , P1_U4003 );
nand NAND2_12834 ( P1_U2618 , P1_U6747 , P1_U4002 );
not NOT1_12835 ( P1_ADD_405_U114 , P1_ADD_405_U40 );
and AND2_12836 ( P1_U2620 , P1_R2144_U145 , P1_U6746 );
and AND2_12837 ( P1_U2621 , P1_R2144_U145 , P1_U6746 );
and AND2_12838 ( P1_U2622 , P1_R2144_U145 , P1_U6746 );
and AND2_12839 ( P1_U2623 , P1_R2144_U145 , P1_U6746 );
and AND2_12840 ( P1_U2624 , P1_R2144_U145 , P1_U6746 );
and AND2_12841 ( P1_U2625 , P1_R2144_U145 , P1_U6746 );
and AND2_12842 ( P1_U2626 , P1_R2144_U145 , P1_U6746 );
and AND2_12843 ( P1_U2627 , P1_R2144_U145 , P1_U6746 );
and AND2_12844 ( P1_U2628 , P1_R2144_U145 , P1_U6746 );
and AND2_12845 ( P1_U2629 , P1_R2144_U145 , P1_U6746 );
and AND2_12846 ( P1_U2630 , P1_R2144_U145 , P1_U6746 );
and AND2_12847 ( P1_U2631 , P1_R2144_U145 , P1_U6746 );
and AND2_12848 ( P1_U2632 , P1_R2144_U145 , P1_U6746 );
and AND2_12849 ( P1_U2633 , P1_R2144_U145 , P1_U6746 );
and AND2_12850 ( P1_U2634 , P1_R2144_U11 , P1_U6746 );
and AND2_12851 ( P1_U2635 , P1_R2144_U37 , P1_U6746 );
and AND2_12852 ( P1_U2636 , P1_R2144_U38 , P1_U6746 );
and AND2_12853 ( P1_U2637 , P1_R2144_U39 , P1_U6746 );
and AND2_12854 ( P1_U2638 , P1_R2144_U40 , P1_U6746 );
and AND2_12855 ( P1_U2639 , P1_R2144_U41 , P1_U6746 );
and AND2_12856 ( P1_U2640 , P1_R2144_U42 , P1_U6746 );
and AND2_12857 ( P1_U2641 , P1_R2144_U30 , P1_U6746 );
and AND2_12858 ( P1_U2642 , P1_R2144_U80 , P1_U6746 );
and AND2_12859 ( P1_U2643 , P1_R2144_U10 , P1_U6746 );
and AND2_12860 ( P1_U2644 , P1_R2144_U9 , P1_U6746 );
and AND2_12861 ( P1_U2645 , P1_R2144_U45 , P1_U6746 );
and AND2_12862 ( P1_U2646 , P1_R2144_U47 , P1_U6746 );
and AND2_12863 ( P1_U2647 , P1_R2144_U8 , P1_U6746 );
nand NAND2_12864 ( P1_U2648 , P1_U3440 , P1_U6869 );
and AND2_12865 ( P1_U2649 , P1_R2144_U50 , P1_U6746 );
and AND2_12866 ( P1_U2650 , P1_STATE2_REG_2_ , P1_U6870 );
nand NAND3_12867 ( P1_U2651 , P1_U6769 , P1_U6768 , P1_U6770 );
nand NAND2_12868 ( P1_U2652 , P1_U6771 , P1_U4009 );
nand NAND2_12869 ( P1_U2653 , P1_U6780 , P1_U4011 );
nand NAND2_12870 ( P1_U2654 , P1_U6784 , P1_U4012 );
nand NAND2_12871 ( P1_U2655 , P1_U6788 , P1_U4013 );
nand NAND2_12872 ( P1_U2656 , P1_U6792 , P1_U4014 );
nand NAND2_12873 ( P1_U2657 , P1_U6796 , P1_U4015 );
nand NAND2_12874 ( P1_U2658 , P1_U6800 , P1_U4016 );
nand NAND2_12875 ( P1_U2659 , P1_U6804 , P1_U4017 );
nand NAND2_12876 ( P1_U2660 , P1_U6808 , P1_U4018 );
nand NAND2_12877 ( P1_U2661 , P1_U6812 , P1_U4019 );
nand NAND2_12878 ( P1_U2662 , P1_U6816 , P1_U4020 );
nand NAND2_12879 ( P1_U2663 , P1_U6825 , P1_U4022 );
nand NAND2_12880 ( P1_U2664 , P1_U6829 , P1_U4023 );
nand NAND2_12881 ( P1_U2665 , P1_U6833 , P1_U4024 );
nand NAND2_12882 ( P1_U2666 , P1_U6837 , P1_U4025 );
nand NAND2_12883 ( P1_U2667 , P1_U6759 , P1_U4006 );
nand NAND4_12884 ( P1_U2668 , P1_U6767 , P1_U6766 , P1_U4008 , P1_U6763 );
nand NAND4_12885 ( P1_U2669 , P1_U6779 , P1_U6778 , P1_U4010 , P1_U6775 );
nand NAND4_12886 ( P1_U2670 , P1_U6824 , P1_U6823 , P1_U4021 , P1_U6820 );
nand NAND4_12887 ( P1_U2671 , P1_U6863 , P1_U6862 , P1_U4027 , P1_U6859 );
nand NAND5_12888 ( P1_U2672 , P1_U6866 , P1_U6864 , P1_U6865 , P1_U6868 , P1_U6867 );
nand NAND2_12889 ( P1_U2673 , P1_U7458 , P1_U7457 );
nand NAND2_12890 ( P1_U2674 , P1_U7460 , P1_U7459 );
nand NAND2_12891 ( P1_U2675 , P1_U4168 , P1_U7463 );
nand NAND2_12892 ( P1_U2676 , P1_U4169 , P1_U7466 );
nand NAND3_12893 ( P1_U2677 , P1_U7794 , P1_U7793 , P1_U7467 );
nand NAND2_12894 ( P1_U2678 , P1_U7456 , P1_U3284 );
nand NAND2_12895 ( P1_U2679 , P1_U7405 , P1_U7404 );
nand NAND2_12896 ( P1_U2680 , P1_U7407 , P1_U7406 );
nand NAND2_12897 ( P1_U2681 , P1_U7411 , P1_U7410 );
nand NAND2_12898 ( P1_U2682 , P1_U7413 , P1_U7412 );
nand NAND2_12899 ( P1_U2683 , P1_U7415 , P1_U7414 );
nand NAND2_12900 ( P1_U2684 , P1_U7417 , P1_U7416 );
nand NAND2_12901 ( P1_U2685 , P1_U7419 , P1_U7418 );
nand NAND2_12902 ( P1_U2686 , P1_U7421 , P1_U7420 );
nand NAND2_12903 ( P1_U2687 , P1_U7423 , P1_U7422 );
nand NAND2_12904 ( P1_U2688 , P1_U7425 , P1_U7424 );
nand NAND2_12905 ( P1_U2689 , P1_U7427 , P1_U7426 );
nand NAND2_12906 ( P1_U2690 , P1_U7429 , P1_U7428 );
nand NAND2_12907 ( P1_U2691 , P1_U7433 , P1_U7432 );
nand NAND2_12908 ( P1_U2692 , P1_U7435 , P1_U7434 );
nand NAND2_12909 ( P1_U2693 , P1_U7437 , P1_U7436 );
nand NAND2_12910 ( P1_U2694 , P1_U7439 , P1_U7438 );
nand NAND2_12911 ( P1_U2695 , P1_U7441 , P1_U7440 );
nand NAND2_12912 ( P1_U2696 , P1_U7443 , P1_U7442 );
nand NAND2_12913 ( P1_U2697 , P1_U7445 , P1_U7444 );
nand NAND2_12914 ( P1_U2698 , P1_U7447 , P1_U7446 );
nand NAND2_12915 ( P1_U2699 , P1_U7449 , P1_U7448 );
nand NAND2_12916 ( P1_U2700 , P1_U7451 , P1_U7450 );
nand NAND2_12917 ( P1_U2701 , P1_U7393 , P1_U7392 );
nand NAND2_12918 ( P1_U2702 , P1_U7395 , P1_U7394 );
nand NAND2_12919 ( P1_U2703 , P1_U7397 , P1_U7396 );
nand NAND2_12920 ( P1_U2704 , P1_U7399 , P1_U7398 );
nand NAND2_12921 ( P1_U2705 , P1_U7401 , P1_U7400 );
nand NAND2_12922 ( P1_U2706 , P1_U7403 , P1_U7402 );
nand NAND2_12923 ( P1_U2707 , P1_U7409 , P1_U7408 );
nand NAND2_12924 ( P1_U2708 , P1_U7431 , P1_U7430 );
nand NAND2_12925 ( P1_U2709 , P1_U7453 , P1_U7452 );
nand NAND2_12926 ( P1_U2710 , P1_U7455 , P1_U7454 );
nand NAND2_12927 ( P1_U2711 , P1_U7377 , P1_U7376 );
nand NAND2_12928 ( P1_U2712 , P1_U7379 , P1_U7378 );
nand NAND2_12929 ( P1_U2713 , P1_U4165 , P1_U4239 );
nand NAND4_12930 ( P1_U2714 , P1_U7386 , P1_U7385 , P1_U4166 , P1_U3434 );
nand NAND2_12931 ( P1_U2715 , P1_U4239 , P1_U4167 );
nand NAND2_12932 ( P1_U2716 , P1_U7365 , P1_U7364 );
nand NAND2_12933 ( P1_U2717 , P1_U7367 , P1_U7366 );
nand NAND2_12934 ( P1_U2718 , P1_U4161 , P1_U7368 );
nand NAND2_12935 ( P1_U2719 , P1_U4162 , P1_U7370 );
nand NAND2_12936 ( P1_U2720 , P1_U4163 , P1_U7372 );
nand NAND2_12937 ( P1_U2721 , P1_U4164 , P1_U7374 );
nand NAND2_12938 ( P1_U2722 , P1_U4159 , P1_U4192 );
and AND2_12939 ( P1_U2723 , P1_U7236 , P1_U7083 );
and AND2_12940 ( P1_U2724 , P1_U7253 , P1_U7083 );
and AND2_12941 ( P1_U2725 , P1_U7270 , P1_U7083 );
and AND2_12942 ( P1_U2726 , P1_U7620 , P1_U7083 );
and AND2_12943 ( P1_U2727 , P1_U7302 , P1_U7083 );
and AND2_12944 ( P1_U2728 , P1_U7319 , P1_U7083 );
and AND2_12945 ( P1_U2729 , P1_U7336 , P1_U7083 );
and AND2_12946 ( P1_U2730 , P1_U7353 , P1_U7083 );
nand NAND2_12947 ( P1_U2731 , P1_U2606 , P1_U7354 );
and AND2_12948 ( P1_U2732 , P1_U7083 , P1_U7082 );
and AND2_12949 ( P1_U2733 , P1_U7114 , P1_U7083 );
and AND2_12950 ( P1_U2734 , P1_U7131 , P1_U7083 );
and AND2_12951 ( P1_U2735 , P1_U7618 , P1_U7083 );
and AND2_12952 ( P1_U2736 , P1_U7163 , P1_U7083 );
and AND2_12953 ( P1_U2737 , P1_U7180 , P1_U7083 );
and AND2_12954 ( P1_U2738 , P1_U7197 , P1_U7083 );
and AND2_12955 ( P1_U2739 , P1_U7214 , P1_U7083 );
and AND2_12956 ( P1_U2740 , P1_INSTQUEUERD_ADDR_REG_4_ , P1_U7063 );
nand NAND2_12957 ( P1_U2741 , P1_U4078 , P1_U7096 );
and AND2_12958 ( P1_U2742 , P1_U7492 , P1_U7491 );
and AND2_12959 ( P1_U2743 , P1_U7506 , P1_U7470 );
and AND2_12960 ( P1_U2744 , P1_U7479 , P1_U7478 );
nand NAND2_12961 ( P1_U2745 , P1_U7048 , P1_U7047 );
nand NAND2_12962 ( P1_U2746 , P1_U7050 , P1_U7049 );
nand NAND2_12963 ( P1_U2747 , P1_U7052 , P1_U7051 );
nand NAND2_12964 ( P1_U2748 , P1_U7616 , P1_U7053 );
nand NAND2_12965 ( P1_U2749 , P1_U7055 , P1_U7054 );
nand NAND2_12966 ( P1_U2750 , P1_U7057 , P1_U7056 );
nand NAND2_12967 ( P1_U2751 , P1_U4061 , P1_U7058 );
nand NAND3_12968 ( P1_U2752 , P1_U4062 , P1_U7060 , P1_U7061 );
and AND2_12969 ( P1_U2753 , P1_U6957 , P1_U6909 );
and AND2_12970 ( P1_U2754 , P1_U6974 , P1_U6909 );
and AND2_12971 ( P1_U2755 , P1_U6991 , P1_U6909 );
and AND2_12972 ( P1_U2756 , P1_U7615 , P1_U6909 );
and AND2_12973 ( P1_U2757 , P1_U7023 , P1_U6909 );
and AND2_12974 ( P1_U2758 , P1_U7040 , P1_U6909 );
and AND2_12975 ( P1_U2759 , P1_U6909 , P1_U6908 );
and AND2_12976 ( P1_U2760 , P1_U6926 , P1_U6909 );
nand NAND2_12977 ( P1_U2761 , P1_U6928 , P1_U6927 );
nand NAND2_12978 ( P1_U2762 , P1_U6930 , P1_U6929 );
nand NAND2_12979 ( P1_U2763 , P1_U6932 , P1_U6931 );
nand NAND2_12980 ( P1_U2764 , P1_U6934 , P1_U6933 );
nand NAND3_12981 ( P1_U2765 , P1_U6936 , P1_U6935 , P1_U6937 );
nand NAND3_12982 ( P1_U2766 , P1_U6939 , P1_U6938 , P1_U6940 );
nand NAND3_12983 ( P1_U2767 , P1_U7043 , P1_U7041 , P1_U7042 );
nand NAND3_12984 ( P1_U2768 , P1_U7046 , P1_U7044 , P1_U7045 );
and AND2_12985 ( P1_U2769 , P1_R2144_U145 , P1_U4159 );
and AND2_12986 ( P1_U2770 , P1_U4159 , P1_R2144_U145 );
and AND2_12987 ( P1_U2771 , P1_U4159 , P1_R2144_U145 );
and AND2_12988 ( P1_U2772 , P1_U4159 , P1_R2144_U145 );
and AND2_12989 ( P1_U2773 , P1_U4159 , P1_R2144_U145 );
and AND2_12990 ( P1_U2774 , P1_U4159 , P1_R2144_U145 );
and AND2_12991 ( P1_U2775 , P1_U4159 , P1_R2144_U145 );
and AND2_12992 ( P1_U2776 , P1_U4159 , P1_R2144_U145 );
and AND2_12993 ( P1_U2777 , P1_U4159 , P1_R2144_U145 );
and AND2_12994 ( P1_U2778 , P1_U4159 , P1_R2144_U145 );
and AND2_12995 ( P1_U2779 , P1_U4159 , P1_R2144_U145 );
and AND2_12996 ( P1_U2780 , P1_U4159 , P1_R2144_U145 );
and AND2_12997 ( P1_U2781 , P1_U4159 , P1_R2144_U145 );
and AND2_12998 ( P1_U2782 , P1_U4159 , P1_R2144_U145 );
and AND2_12999 ( P1_U2783 , P1_U4159 , P1_R2144_U145 );
and AND2_13000 ( P1_U2784 , P1_U4159 , P1_R2144_U11 );
and AND2_13001 ( P1_U2785 , P1_U4159 , P1_R2144_U37 );
and AND2_13002 ( P1_U2786 , P1_U4159 , P1_R2144_U38 );
and AND2_13003 ( P1_U2787 , P1_U4159 , P1_R2144_U39 );
and AND2_13004 ( P1_U2788 , P1_U4159 , P1_R2144_U40 );
and AND2_13005 ( P1_U2789 , P1_U4159 , P1_R2144_U41 );
and AND2_13006 ( P1_U2790 , P1_U4159 , P1_R2144_U42 );
and AND2_13007 ( P1_U2791 , P1_U4159 , P1_R2144_U30 );
nand NAND2_13008 ( P1_U2792 , P1_U6872 , P1_U6871 );
nand NAND2_13009 ( P1_U2793 , P1_U6874 , P1_U6873 );
nand NAND2_13010 ( P1_U2794 , P1_U6876 , P1_U6875 );
nand NAND2_13011 ( P1_U2795 , P1_U6878 , P1_U6877 );
nand NAND2_13012 ( P1_U2796 , P1_U6880 , P1_U6879 );
nand NAND2_13013 ( P1_U2797 , P1_U6882 , P1_U6881 );
nand NAND3_13014 ( P1_U2798 , P1_U6884 , P1_U6885 , P1_U6883 );
nand NAND3_13015 ( P1_U2799 , P1_U4028 , P1_U6887 , P1_U6886 );
nand NAND3_13016 ( P1_U2800 , P1_U6890 , P1_U6891 , P1_U6889 );
nand NAND3_13017 ( P1_U2801 , P1_U6617 , P1_U3432 , P1_U7498 );
nand NAND2_13018 ( P1_U2802 , P1_U7650 , P1_U6613 );
nand NAND2_13019 ( P1_U2803 , P1_U6612 , P1_U6611 );
nand NAND3_13020 ( P1_U2804 , P1_U7769 , P1_U7768 , P1_U4243 );
nand NAND3_13021 ( P1_U2805 , P1_U7765 , P1_U7764 , P1_U4243 );
nand NAND2_13022 ( P1_U2806 , P1_U6601 , P1_U4248 );
nand NAND3_13023 ( P1_U2807 , P1_U7757 , P1_U7756 , P1_U4240 );
nand NAND3_13024 ( P1_U2808 , P1_U7747 , P1_U7746 , P1_U4240 );
nand NAND5_13025 ( P1_U2809 , P1_U6593 , P1_U3948 , P1_U3949 , P1_U6591 , P1_U6595 );
nand NAND5_13026 ( P1_U2810 , P1_U6586 , P1_U3946 , P1_U3947 , P1_U6584 , P1_U6588 );
nand NAND5_13027 ( P1_U2811 , P1_U6579 , P1_U3944 , P1_U3945 , P1_U6577 , P1_U6581 );
nand NAND5_13028 ( P1_U2812 , P1_U6572 , P1_U3942 , P1_U3943 , P1_U6570 , P1_U6574 );
nand NAND5_13029 ( P1_U2813 , P1_U6565 , P1_U3940 , P1_U3941 , P1_U6563 , P1_U6567 );
nand NAND5_13030 ( P1_U2814 , P1_U6558 , P1_U3938 , P1_U3939 , P1_U6556 , P1_U6560 );
nand NAND5_13031 ( P1_U2815 , P1_U6551 , P1_U3936 , P1_U3937 , P1_U6549 , P1_U6553 );
nand NAND5_13032 ( P1_U2816 , P1_U6544 , P1_U3934 , P1_U3935 , P1_U6542 , P1_U6546 );
nand NAND5_13033 ( P1_U2817 , P1_U6537 , P1_U3932 , P1_U3933 , P1_U6535 , P1_U6539 );
nand NAND5_13034 ( P1_U2818 , P1_U6530 , P1_U3930 , P1_U3931 , P1_U6528 , P1_U6532 );
nand NAND5_13035 ( P1_U2819 , P1_U6523 , P1_U3928 , P1_U3929 , P1_U6521 , P1_U6525 );
nand NAND5_13036 ( P1_U2820 , P1_U6516 , P1_U3926 , P1_U3927 , P1_U6514 , P1_U6518 );
nand NAND5_13037 ( P1_U2821 , P1_U3924 , P1_U6509 , P1_U3925 , P1_U6507 , P1_U6511 );
nand NAND5_13038 ( P1_U2822 , P1_U3922 , P1_U6502 , P1_U3923 , P1_U6500 , P1_U6504 );
nand NAND5_13039 ( P1_U2823 , P1_U3920 , P1_U6495 , P1_U3921 , P1_U6493 , P1_U6497 );
nand NAND5_13040 ( P1_U2824 , P1_U6488 , P1_U6487 , P1_U3919 , P1_U3918 , P1_U6490 );
nand NAND5_13041 ( P1_U2825 , P1_U6481 , P1_U6480 , P1_U3917 , P1_U3916 , P1_U6483 );
nand NAND5_13042 ( P1_U2826 , P1_U3915 , P1_U6474 , P1_U3914 , P1_U6473 , P1_U6476 );
nand NAND5_13043 ( P1_U2827 , P1_U3913 , P1_U6467 , P1_U3912 , P1_U6466 , P1_U6469 );
nand NAND5_13044 ( P1_U2828 , P1_U3911 , P1_U6460 , P1_U3910 , P1_U6459 , P1_U6462 );
nand NAND5_13045 ( P1_U2829 , P1_U3909 , P1_U6453 , P1_U3908 , P1_U6452 , P1_U6455 );
nand NAND5_13046 ( P1_U2830 , P1_U3907 , P1_U6446 , P1_U3906 , P1_U6445 , P1_U6448 );
nand NAND5_13047 ( P1_U2831 , P1_U3905 , P1_U6439 , P1_U3904 , P1_U6438 , P1_U6441 );
nand NAND5_13048 ( P1_U2832 , P1_U3903 , P1_U6432 , P1_U3902 , P1_U6431 , P1_U6434 );
nand NAND5_13049 ( P1_U2833 , P1_U3901 , P1_U6425 , P1_U3900 , P1_U6424 , P1_U6427 );
nand NAND5_13050 ( P1_U2834 , P1_U3899 , P1_U6418 , P1_U3898 , P1_U6417 , P1_U6420 );
nand NAND4_13051 ( P1_U2835 , P1_U3896 , P1_U6409 , P1_U6410 , P1_U3897 );
nand NAND5_13052 ( P1_U2836 , P1_U3894 , P1_U6401 , P1_U3895 , P1_U6403 , P1_U6402 );
nand NAND4_13053 ( P1_U2837 , P1_U6393 , P1_U6392 , P1_U6394 , P1_U3893 );
nand NAND4_13054 ( P1_U2838 , P1_U6385 , P1_U6384 , P1_U6386 , P1_U3892 );
nand NAND4_13055 ( P1_U2839 , P1_U6377 , P1_U6376 , P1_U6378 , P1_U3891 );
nand NAND4_13056 ( P1_U2840 , P1_U6369 , P1_U6368 , P1_U6370 , P1_U3890 );
nand NAND2_13057 ( P1_U2841 , P1_U6359 , P1_U6358 );
nand NAND3_13058 ( P1_U2842 , P1_U6356 , P1_U6357 , P1_U6355 );
nand NAND3_13059 ( P1_U2843 , P1_U6353 , P1_U6354 , P1_U6352 );
nand NAND3_13060 ( P1_U2844 , P1_U6350 , P1_U6351 , P1_U6349 );
nand NAND3_13061 ( P1_U2845 , P1_U6347 , P1_U6348 , P1_U6346 );
nand NAND3_13062 ( P1_U2846 , P1_U6344 , P1_U6345 , P1_U6343 );
nand NAND3_13063 ( P1_U2847 , P1_U6341 , P1_U6342 , P1_U6340 );
nand NAND3_13064 ( P1_U2848 , P1_U6338 , P1_U6339 , P1_U6337 );
nand NAND3_13065 ( P1_U2849 , P1_U6335 , P1_U6336 , P1_U6334 );
nand NAND3_13066 ( P1_U2850 , P1_U6332 , P1_U6333 , P1_U6331 );
nand NAND3_13067 ( P1_U2851 , P1_U6329 , P1_U6330 , P1_U6328 );
nand NAND3_13068 ( P1_U2852 , P1_U6326 , P1_U6327 , P1_U6325 );
nand NAND3_13069 ( P1_U2853 , P1_U6323 , P1_U6324 , P1_U6322 );
nand NAND3_13070 ( P1_U2854 , P1_U6320 , P1_U6321 , P1_U6319 );
nand NAND3_13071 ( P1_U2855 , P1_U6317 , P1_U6318 , P1_U6316 );
nand NAND3_13072 ( P1_U2856 , P1_U6314 , P1_U6315 , P1_U6313 );
nand NAND3_13073 ( P1_U2857 , P1_U6311 , P1_U6312 , P1_U6310 );
nand NAND3_13074 ( P1_U2858 , P1_U6308 , P1_U6309 , P1_U6307 );
nand NAND3_13075 ( P1_U2859 , P1_U6305 , P1_U6306 , P1_U6304 );
nand NAND3_13076 ( P1_U2860 , P1_U6302 , P1_U6303 , P1_U6301 );
nand NAND3_13077 ( P1_U2861 , P1_U6299 , P1_U6300 , P1_U6298 );
nand NAND3_13078 ( P1_U2862 , P1_U6296 , P1_U6297 , P1_U6295 );
nand NAND3_13079 ( P1_U2863 , P1_U6293 , P1_U6294 , P1_U6292 );
nand NAND3_13080 ( P1_U2864 , P1_U6290 , P1_U6291 , P1_U6289 );
nand NAND3_13081 ( P1_U2865 , P1_U6287 , P1_U6288 , P1_U6286 );
nand NAND3_13082 ( P1_U2866 , P1_U6284 , P1_U6285 , P1_U6283 );
nand NAND3_13083 ( P1_U2867 , P1_U6281 , P1_U6282 , P1_U6280 );
nand NAND3_13084 ( P1_U2868 , P1_U6278 , P1_U6279 , P1_U6277 );
nand NAND3_13085 ( P1_U2869 , P1_U6275 , P1_U6276 , P1_U6274 );
nand NAND3_13086 ( P1_U2870 , P1_U6272 , P1_U6273 , P1_U6271 );
nand NAND3_13087 ( P1_U2871 , P1_U6269 , P1_U6270 , P1_U6268 );
nand NAND3_13088 ( P1_U2872 , P1_U6266 , P1_U6265 , P1_U6267 );
nand NAND2_13089 ( P1_U2873 , P1_U4176 , P1_U6262 );
nand NAND4_13090 ( P1_U2874 , P1_U6259 , P1_U6258 , P1_U6261 , P1_U6260 );
nand NAND4_13091 ( P1_U2875 , P1_U6255 , P1_U6254 , P1_U6257 , P1_U6256 );
nand NAND4_13092 ( P1_U2876 , P1_U6251 , P1_U6250 , P1_U6253 , P1_U6252 );
nand NAND4_13093 ( P1_U2877 , P1_U6247 , P1_U6246 , P1_U6249 , P1_U6248 );
nand NAND4_13094 ( P1_U2878 , P1_U6243 , P1_U6242 , P1_U6245 , P1_U6244 );
nand NAND4_13095 ( P1_U2879 , P1_U6239 , P1_U6238 , P1_U6241 , P1_U6240 );
nand NAND4_13096 ( P1_U2880 , P1_U6235 , P1_U6234 , P1_U6237 , P1_U6236 );
nand NAND4_13097 ( P1_U2881 , P1_U6231 , P1_U6230 , P1_U6233 , P1_U6232 );
nand NAND4_13098 ( P1_U2882 , P1_U6227 , P1_U6226 , P1_U6229 , P1_U6228 );
nand NAND4_13099 ( P1_U2883 , P1_U6223 , P1_U6222 , P1_U6225 , P1_U6224 );
nand NAND4_13100 ( P1_U2884 , P1_U6219 , P1_U6218 , P1_U6221 , P1_U6220 );
nand NAND4_13101 ( P1_U2885 , P1_U6215 , P1_U6214 , P1_U6217 , P1_U6216 );
nand NAND4_13102 ( P1_U2886 , P1_U6211 , P1_U6210 , P1_U6213 , P1_U6212 );
nand NAND4_13103 ( P1_U2887 , P1_U6207 , P1_U6206 , P1_U6209 , P1_U6208 );
nand NAND4_13104 ( P1_U2888 , P1_U6203 , P1_U6202 , P1_U6205 , P1_U6204 );
nand NAND3_13105 ( P1_U2889 , P1_U6201 , P1_U6199 , P1_U6200 );
nand NAND3_13106 ( P1_U2890 , P1_U6198 , P1_U6196 , P1_U6197 );
nand NAND3_13107 ( P1_U2891 , P1_U6195 , P1_U6193 , P1_U6194 );
nand NAND3_13108 ( P1_U2892 , P1_U6192 , P1_U6190 , P1_U6191 );
nand NAND3_13109 ( P1_U2893 , P1_U6189 , P1_U6187 , P1_U6188 );
nand NAND3_13110 ( P1_U2894 , P1_U6186 , P1_U6184 , P1_U6185 );
nand NAND3_13111 ( P1_U2895 , P1_U6183 , P1_U6181 , P1_U6182 );
nand NAND3_13112 ( P1_U2896 , P1_U6180 , P1_U6178 , P1_U6179 );
nand NAND3_13113 ( P1_U2897 , P1_U6177 , P1_U6175 , P1_U6176 );
nand NAND3_13114 ( P1_U2898 , P1_U6174 , P1_U6172 , P1_U6173 );
nand NAND3_13115 ( P1_U2899 , P1_U6171 , P1_U6169 , P1_U6170 );
nand NAND3_13116 ( P1_U2900 , P1_U6168 , P1_U6166 , P1_U6167 );
nand NAND3_13117 ( P1_U2901 , P1_U6165 , P1_U6163 , P1_U6164 );
nand NAND3_13118 ( P1_U2902 , P1_U6162 , P1_U6160 , P1_U6161 );
nand NAND3_13119 ( P1_U2903 , P1_U6158 , P1_U6157 , P1_U6159 );
nand NAND3_13120 ( P1_U2904 , P1_U6155 , P1_U6154 , P1_U6156 );
and AND2_13121 ( P1_U2905 , P1_DATAO_REG_31_ , P1_U6055 );
nand NAND2_13122 ( P1_U2906 , P1_U3882 , P1_U6146 );
nand NAND2_13123 ( P1_U2907 , P1_U3881 , P1_U6143 );
nand NAND2_13124 ( P1_U2908 , P1_U3880 , P1_U6140 );
nand NAND2_13125 ( P1_U2909 , P1_U3879 , P1_U6137 );
nand NAND2_13126 ( P1_U2910 , P1_U3878 , P1_U6134 );
nand NAND2_13127 ( P1_U2911 , P1_U3877 , P1_U6131 );
nand NAND2_13128 ( P1_U2912 , P1_U3876 , P1_U6128 );
nand NAND2_13129 ( P1_U2913 , P1_U3875 , P1_U6125 );
nand NAND2_13130 ( P1_U2914 , P1_U3874 , P1_U6122 );
nand NAND2_13131 ( P1_U2915 , P1_U3873 , P1_U6119 );
nand NAND2_13132 ( P1_U2916 , P1_U3872 , P1_U6116 );
nand NAND2_13133 ( P1_U2917 , P1_U3871 , P1_U6113 );
nand NAND2_13134 ( P1_U2918 , P1_U3870 , P1_U6110 );
nand NAND2_13135 ( P1_U2919 , P1_U3869 , P1_U6107 );
nand NAND2_13136 ( P1_U2920 , P1_U3868 , P1_U6104 );
nand NAND3_13137 ( P1_U2921 , P1_U6102 , P1_U6101 , P1_U6103 );
nand NAND3_13138 ( P1_U2922 , P1_U6099 , P1_U6098 , P1_U6100 );
nand NAND3_13139 ( P1_U2923 , P1_U6096 , P1_U6095 , P1_U6097 );
nand NAND3_13140 ( P1_U2924 , P1_U6093 , P1_U6092 , P1_U6094 );
nand NAND3_13141 ( P1_U2925 , P1_U6090 , P1_U6089 , P1_U6091 );
nand NAND3_13142 ( P1_U2926 , P1_U6087 , P1_U6086 , P1_U6088 );
nand NAND3_13143 ( P1_U2927 , P1_U6084 , P1_U6083 , P1_U6085 );
nand NAND3_13144 ( P1_U2928 , P1_U6081 , P1_U6080 , P1_U6082 );
nand NAND3_13145 ( P1_U2929 , P1_U6078 , P1_U6077 , P1_U6079 );
nand NAND3_13146 ( P1_U2930 , P1_U6075 , P1_U6074 , P1_U6076 );
nand NAND3_13147 ( P1_U2931 , P1_U6072 , P1_U6071 , P1_U6073 );
nand NAND3_13148 ( P1_U2932 , P1_U6069 , P1_U6068 , P1_U6070 );
nand NAND3_13149 ( P1_U2933 , P1_U6066 , P1_U6065 , P1_U6067 );
nand NAND3_13150 ( P1_U2934 , P1_U6063 , P1_U6062 , P1_U6064 );
nand NAND3_13151 ( P1_U2935 , P1_U6060 , P1_U6059 , P1_U6061 );
nand NAND3_13152 ( P1_U2936 , P1_U6057 , P1_U6056 , P1_U6058 );
nand NAND2_13153 ( P1_U2937 , P1_U7540 , P1_U7542 );
nand NAND2_13154 ( P1_U2938 , P1_U7539 , P1_U7544 );
nand NAND2_13155 ( P1_U2939 , P1_U7538 , P1_U7546 );
nand NAND2_13156 ( P1_U2940 , P1_U7537 , P1_U7548 );
nand NAND2_13157 ( P1_U2941 , P1_U7536 , P1_U7550 );
nand NAND2_13158 ( P1_U2942 , P1_U7535 , P1_U7552 );
nand NAND2_13159 ( P1_U2943 , P1_U7534 , P1_U7554 );
nand NAND2_13160 ( P1_U2944 , P1_U7533 , P1_U7556 );
nand NAND2_13161 ( P1_U2945 , P1_U7532 , P1_U7558 );
nand NAND2_13162 ( P1_U2946 , P1_U7531 , P1_U7560 );
nand NAND2_13163 ( P1_U2947 , P1_U7530 , P1_U7562 );
nand NAND2_13164 ( P1_U2948 , P1_U7529 , P1_U7564 );
nand NAND2_13165 ( P1_U2949 , P1_U7528 , P1_U7566 );
nand NAND2_13166 ( P1_U2950 , P1_U7527 , P1_U7568 );
nand NAND2_13167 ( P1_U2951 , P1_U7526 , P1_U7570 );
nand NAND2_13168 ( P1_U2952 , P1_U7525 , P1_U7572 );
nand NAND2_13169 ( P1_U2953 , P1_U7524 , P1_U7574 );
nand NAND2_13170 ( P1_U2954 , P1_U7523 , P1_U7576 );
nand NAND2_13171 ( P1_U2955 , P1_U7522 , P1_U7578 );
nand NAND2_13172 ( P1_U2956 , P1_U7521 , P1_U7580 );
nand NAND2_13173 ( P1_U2957 , P1_U7520 , P1_U7582 );
nand NAND2_13174 ( P1_U2958 , P1_U7519 , P1_U7584 );
nand NAND2_13175 ( P1_U2959 , P1_U7518 , P1_U7586 );
nand NAND2_13176 ( P1_U2960 , P1_U7517 , P1_U7588 );
nand NAND2_13177 ( P1_U2961 , P1_U7516 , P1_U7590 );
nand NAND2_13178 ( P1_U2962 , P1_U7515 , P1_U7592 );
nand NAND2_13179 ( P1_U2963 , P1_U7514 , P1_U7594 );
nand NAND2_13180 ( P1_U2964 , P1_U7513 , P1_U7596 );
nand NAND2_13181 ( P1_U2965 , P1_U7512 , P1_U7598 );
nand NAND2_13182 ( P1_U2966 , P1_U7511 , P1_U7600 );
nand NAND2_13183 ( P1_U2967 , P1_U7510 , P1_U7602 );
nand NAND5_13184 ( P1_U2968 , P1_U5956 , P1_U5954 , P1_U5958 , P1_U5955 , P1_U5957 );
nand NAND5_13185 ( P1_U2969 , P1_U5951 , P1_U5949 , P1_U5953 , P1_U5950 , P1_U5952 );
nand NAND5_13186 ( P1_U2970 , P1_U5946 , P1_U5944 , P1_U5948 , P1_U5945 , P1_U5947 );
nand NAND5_13187 ( P1_U2971 , P1_U5941 , P1_U5939 , P1_U5943 , P1_U5940 , P1_U5942 );
nand NAND5_13188 ( P1_U2972 , P1_U5936 , P1_U5934 , P1_U5938 , P1_U5935 , P1_U5937 );
nand NAND5_13189 ( P1_U2973 , P1_U5931 , P1_U5929 , P1_U5933 , P1_U5930 , P1_U5932 );
nand NAND5_13190 ( P1_U2974 , P1_U5926 , P1_U5924 , P1_U5928 , P1_U5925 , P1_U5927 );
nand NAND5_13191 ( P1_U2975 , P1_U5921 , P1_U5919 , P1_U5923 , P1_U5920 , P1_U5922 );
nand NAND5_13192 ( P1_U2976 , P1_U5916 , P1_U5914 , P1_U5918 , P1_U5915 , P1_U5917 );
nand NAND5_13193 ( P1_U2977 , P1_U5911 , P1_U5909 , P1_U5913 , P1_U5910 , P1_U5912 );
nand NAND5_13194 ( P1_U2978 , P1_U5906 , P1_U5904 , P1_U5908 , P1_U5905 , P1_U5907 );
nand NAND5_13195 ( P1_U2979 , P1_U5901 , P1_U5899 , P1_U5903 , P1_U5900 , P1_U5902 );
nand NAND5_13196 ( P1_U2980 , P1_U5896 , P1_U5894 , P1_U5898 , P1_U5895 , P1_U5897 );
nand NAND5_13197 ( P1_U2981 , P1_U5891 , P1_U5889 , P1_U5893 , P1_U5890 , P1_U5892 );
nand NAND5_13198 ( P1_U2982 , P1_U5886 , P1_U5884 , P1_U5888 , P1_U5885 , P1_U5887 );
nand NAND5_13199 ( P1_U2983 , P1_U5881 , P1_U5879 , P1_U5883 , P1_U5880 , P1_U5882 );
nand NAND5_13200 ( P1_U2984 , P1_U5876 , P1_U5874 , P1_U5878 , P1_U5875 , P1_U5877 );
nand NAND5_13201 ( P1_U2985 , P1_U5871 , P1_U5869 , P1_U5873 , P1_U5870 , P1_U5872 );
nand NAND5_13202 ( P1_U2986 , P1_U5866 , P1_U5864 , P1_U5868 , P1_U5865 , P1_U5867 );
nand NAND5_13203 ( P1_U2987 , P1_U5861 , P1_U5859 , P1_U5863 , P1_U5860 , P1_U5862 );
nand NAND5_13204 ( P1_U2988 , P1_U5856 , P1_U5854 , P1_U5858 , P1_U5855 , P1_U5857 );
nand NAND5_13205 ( P1_U2989 , P1_U5851 , P1_U5849 , P1_U5853 , P1_U5850 , P1_U5852 );
nand NAND5_13206 ( P1_U2990 , P1_U5846 , P1_U5844 , P1_U5848 , P1_U5845 , P1_U5847 );
nand NAND5_13207 ( P1_U2991 , P1_U5841 , P1_U5839 , P1_U5843 , P1_U5840 , P1_U5842 );
nand NAND5_13208 ( P1_U2992 , P1_U5836 , P1_U5834 , P1_U5835 , P1_U5838 , P1_U5837 );
nand NAND5_13209 ( P1_U2993 , P1_U5831 , P1_U5829 , P1_U5830 , P1_U5833 , P1_U5832 );
nand NAND5_13210 ( P1_U2994 , P1_U5826 , P1_U5824 , P1_U5825 , P1_U5828 , P1_U5827 );
nand NAND5_13211 ( P1_U2995 , P1_U5821 , P1_U5819 , P1_U5820 , P1_U5823 , P1_U5822 );
nand NAND5_13212 ( P1_U2996 , P1_U5816 , P1_U5814 , P1_U5815 , P1_U5818 , P1_U5817 );
nand NAND5_13213 ( P1_U2997 , P1_U5811 , P1_U5809 , P1_U5810 , P1_U5813 , P1_U5812 );
nand NAND5_13214 ( P1_U2998 , P1_U5805 , P1_U5804 , P1_U5806 , P1_U5808 , P1_U5807 );
nand NAND5_13215 ( P1_U2999 , P1_U5800 , P1_U5799 , P1_U5801 , P1_U5803 , P1_U5802 );
nand NAND4_13216 ( P1_U3000 , P1_U3861 , P1_U3859 , P1_U5787 , P1_U5789 );
nand NAND4_13217 ( P1_U3001 , P1_U3858 , P1_U3856 , P1_U5780 , P1_U5782 );
nand NAND4_13218 ( P1_U3002 , P1_U3855 , P1_U3853 , P1_U5773 , P1_U5775 );
nand NAND4_13219 ( P1_U3003 , P1_U3852 , P1_U3850 , P1_U5766 , P1_U5768 );
nand NAND4_13220 ( P1_U3004 , P1_U3849 , P1_U3847 , P1_U5759 , P1_U5761 );
nand NAND4_13221 ( P1_U3005 , P1_U3846 , P1_U3844 , P1_U5752 , P1_U5754 );
nand NAND4_13222 ( P1_U3006 , P1_U3843 , P1_U3841 , P1_U5745 , P1_U5747 );
nand NAND4_13223 ( P1_U3007 , P1_U3840 , P1_U3838 , P1_U5738 , P1_U5740 );
nand NAND4_13224 ( P1_U3008 , P1_U3837 , P1_U3835 , P1_U5731 , P1_U5733 );
nand NAND4_13225 ( P1_U3009 , P1_U3834 , P1_U3832 , P1_U5724 , P1_U5726 );
nand NAND4_13226 ( P1_U3010 , P1_U3831 , P1_U3829 , P1_U5717 , P1_U5719 );
nand NAND4_13227 ( P1_U3011 , P1_U3828 , P1_U3826 , P1_U5710 , P1_U5712 );
nand NAND4_13228 ( P1_U3012 , P1_U3825 , P1_U3823 , P1_U5703 , P1_U5705 );
nand NAND4_13229 ( P1_U3013 , P1_U3822 , P1_U3820 , P1_U5696 , P1_U5698 );
nand NAND4_13230 ( P1_U3014 , P1_U3819 , P1_U3817 , P1_U5689 , P1_U5691 );
nand NAND4_13231 ( P1_U3015 , P1_U3816 , P1_U3814 , P1_U5682 , P1_U5684 );
nand NAND4_13232 ( P1_U3016 , P1_U3813 , P1_U3811 , P1_U5675 , P1_U5677 );
nand NAND4_13233 ( P1_U3017 , P1_U3810 , P1_U3808 , P1_U5668 , P1_U5670 );
nand NAND4_13234 ( P1_U3018 , P1_U3807 , P1_U3805 , P1_U5661 , P1_U5663 );
nand NAND3_13235 ( P1_U3019 , P1_U3802 , P1_U3804 , P1_U5656 );
nand NAND3_13236 ( P1_U3020 , P1_U3799 , P1_U3801 , P1_U5649 );
nand NAND3_13237 ( P1_U3021 , P1_U3796 , P1_U3798 , P1_U5642 );
nand NAND3_13238 ( P1_U3022 , P1_U3793 , P1_U3795 , P1_U5635 );
nand NAND3_13239 ( P1_U3023 , P1_U3790 , P1_U3792 , P1_U5628 );
nand NAND3_13240 ( P1_U3024 , P1_U3787 , P1_U3789 , P1_U5621 );
nand NAND3_13241 ( P1_U3025 , P1_U3784 , P1_U3786 , P1_U5614 );
nand NAND3_13242 ( P1_U3026 , P1_U3781 , P1_U3783 , P1_U5607 );
nand NAND3_13243 ( P1_U3027 , P1_U3778 , P1_U3780 , P1_U5600 );
nand NAND2_13244 ( P1_U3028 , P1_U3775 , P1_U3776 );
nand NAND3_13245 ( P1_U3029 , P1_U3772 , P1_U3771 , P1_U3774 );
nand NAND3_13246 ( P1_U3030 , P1_U3768 , P1_U3767 , P1_U3770 );
nand NAND3_13247 ( P1_U3031 , P1_U3764 , P1_U3763 , P1_U3766 );
and AND2_13248 ( P1_U3032 , P1_INSTQUEUEWR_ADDR_REG_4_ , P1_U5537 );
nand NAND3_13249 ( P1_U3033 , P1_U5460 , P1_U5459 , P1_U3730 );
nand NAND3_13250 ( P1_U3034 , P1_U5455 , P1_U5454 , P1_U3729 );
nand NAND3_13251 ( P1_U3035 , P1_U5450 , P1_U5449 , P1_U3728 );
nand NAND3_13252 ( P1_U3036 , P1_U5445 , P1_U5444 , P1_U3727 );
nand NAND3_13253 ( P1_U3037 , P1_U7612 , P1_U5440 , P1_U3726 );
nand NAND3_13254 ( P1_U3038 , P1_U5436 , P1_U5435 , P1_U3725 );
nand NAND3_13255 ( P1_U3039 , P1_U5431 , P1_U5430 , P1_U3724 );
nand NAND3_13256 ( P1_U3040 , P1_U5426 , P1_U5425 , P1_U3723 );
nand NAND3_13257 ( P1_U3041 , P1_U5404 , P1_U5403 , P1_U3721 );
nand NAND3_13258 ( P1_U3042 , P1_U5399 , P1_U5398 , P1_U3720 );
nand NAND3_13259 ( P1_U3043 , P1_U5394 , P1_U5393 , P1_U3719 );
nand NAND3_13260 ( P1_U3044 , P1_U5389 , P1_U5388 , P1_U3718 );
nand NAND3_13261 ( P1_U3045 , P1_U5384 , P1_U5383 , P1_U3717 );
nand NAND3_13262 ( P1_U3046 , P1_U5379 , P1_U5378 , P1_U3716 );
nand NAND3_13263 ( P1_U3047 , P1_U5374 , P1_U5373 , P1_U3715 );
nand NAND3_13264 ( P1_U3048 , P1_U5369 , P1_U5368 , P1_U3714 );
nand NAND3_13265 ( P1_U3049 , P1_U5346 , P1_U5345 , P1_U3712 );
nand NAND3_13266 ( P1_U3050 , P1_U5341 , P1_U5340 , P1_U3711 );
nand NAND3_13267 ( P1_U3051 , P1_U5336 , P1_U5335 , P1_U3710 );
nand NAND3_13268 ( P1_U3052 , P1_U5331 , P1_U5330 , P1_U3709 );
nand NAND3_13269 ( P1_U3053 , P1_U5326 , P1_U5325 , P1_U3708 );
nand NAND3_13270 ( P1_U3054 , P1_U5321 , P1_U5320 , P1_U3707 );
nand NAND3_13271 ( P1_U3055 , P1_U5316 , P1_U5315 , P1_U3706 );
nand NAND3_13272 ( P1_U3056 , P1_U5311 , P1_U5310 , P1_U3705 );
nand NAND3_13273 ( P1_U3057 , P1_U5289 , P1_U5288 , P1_U3703 );
nand NAND3_13274 ( P1_U3058 , P1_U5284 , P1_U5283 , P1_U3702 );
nand NAND3_13275 ( P1_U3059 , P1_U5279 , P1_U5278 , P1_U3701 );
nand NAND3_13276 ( P1_U3060 , P1_U5274 , P1_U5273 , P1_U3700 );
nand NAND3_13277 ( P1_U3061 , P1_U5269 , P1_U5268 , P1_U3699 );
nand NAND3_13278 ( P1_U3062 , P1_U5264 , P1_U5263 , P1_U3698 );
nand NAND3_13279 ( P1_U3063 , P1_U5259 , P1_U5258 , P1_U3697 );
nand NAND3_13280 ( P1_U3064 , P1_U5254 , P1_U5253 , P1_U3696 );
nand NAND3_13281 ( P1_U3065 , P1_U5231 , P1_U5230 , P1_U3694 );
nand NAND3_13282 ( P1_U3066 , P1_U5226 , P1_U5225 , P1_U3693 );
nand NAND3_13283 ( P1_U3067 , P1_U5221 , P1_U5220 , P1_U3692 );
nand NAND3_13284 ( P1_U3068 , P1_U5216 , P1_U5215 , P1_U3691 );
nand NAND3_13285 ( P1_U3069 , P1_U5211 , P1_U5210 , P1_U3690 );
nand NAND3_13286 ( P1_U3070 , P1_U5206 , P1_U5205 , P1_U3689 );
nand NAND3_13287 ( P1_U3071 , P1_U5201 , P1_U5200 , P1_U3688 );
nand NAND3_13288 ( P1_U3072 , P1_U5196 , P1_U5195 , P1_U3687 );
nand NAND3_13289 ( P1_U3073 , P1_U5174 , P1_U5173 , P1_U3685 );
nand NAND3_13290 ( P1_U3074 , P1_U5169 , P1_U5168 , P1_U3684 );
nand NAND3_13291 ( P1_U3075 , P1_U5164 , P1_U5163 , P1_U3683 );
nand NAND3_13292 ( P1_U3076 , P1_U5159 , P1_U5158 , P1_U3682 );
nand NAND3_13293 ( P1_U3077 , P1_U5154 , P1_U5153 , P1_U3681 );
nand NAND3_13294 ( P1_U3078 , P1_U5149 , P1_U5148 , P1_U3680 );
nand NAND3_13295 ( P1_U3079 , P1_U5144 , P1_U5143 , P1_U3679 );
nand NAND3_13296 ( P1_U3080 , P1_U5139 , P1_U5138 , P1_U3678 );
nand NAND3_13297 ( P1_U3081 , P1_U5116 , P1_U5115 , P1_U3676 );
nand NAND3_13298 ( P1_U3082 , P1_U5111 , P1_U5110 , P1_U3675 );
nand NAND3_13299 ( P1_U3083 , P1_U5106 , P1_U5105 , P1_U3674 );
nand NAND3_13300 ( P1_U3084 , P1_U5101 , P1_U5100 , P1_U3673 );
nand NAND3_13301 ( P1_U3085 , P1_U5096 , P1_U5095 , P1_U3672 );
nand NAND3_13302 ( P1_U3086 , P1_U5091 , P1_U5090 , P1_U3671 );
nand NAND3_13303 ( P1_U3087 , P1_U5086 , P1_U5085 , P1_U3670 );
nand NAND3_13304 ( P1_U3088 , P1_U5081 , P1_U5080 , P1_U3669 );
nand NAND3_13305 ( P1_U3089 , P1_U5059 , P1_U5058 , P1_U3667 );
nand NAND3_13306 ( P1_U3090 , P1_U5054 , P1_U5053 , P1_U3666 );
nand NAND3_13307 ( P1_U3091 , P1_U5049 , P1_U5048 , P1_U3665 );
nand NAND3_13308 ( P1_U3092 , P1_U5044 , P1_U5043 , P1_U3664 );
nand NAND3_13309 ( P1_U3093 , P1_U5039 , P1_U5038 , P1_U3663 );
nand NAND3_13310 ( P1_U3094 , P1_U5034 , P1_U5033 , P1_U3662 );
nand NAND3_13311 ( P1_U3095 , P1_U5029 , P1_U5028 , P1_U3661 );
nand NAND3_13312 ( P1_U3096 , P1_U5024 , P1_U5023 , P1_U3660 );
nand NAND3_13313 ( P1_U3097 , P1_U5003 , P1_U5002 , P1_U3658 );
nand NAND3_13314 ( P1_U3098 , P1_U4998 , P1_U4997 , P1_U3657 );
nand NAND3_13315 ( P1_U3099 , P1_U4993 , P1_U4992 , P1_U3656 );
nand NAND3_13316 ( P1_U3100 , P1_U4988 , P1_U4987 , P1_U3655 );
nand NAND3_13317 ( P1_U3101 , P1_U4983 , P1_U4982 , P1_U3654 );
nand NAND3_13318 ( P1_U3102 , P1_U4978 , P1_U4977 , P1_U3653 );
nand NAND3_13319 ( P1_U3103 , P1_U4973 , P1_U4972 , P1_U3652 );
nand NAND3_13320 ( P1_U3104 , P1_U4968 , P1_U4967 , P1_U3651 );
nand NAND3_13321 ( P1_U3105 , P1_U4946 , P1_U4945 , P1_U3649 );
nand NAND3_13322 ( P1_U3106 , P1_U4941 , P1_U4940 , P1_U3648 );
nand NAND3_13323 ( P1_U3107 , P1_U4936 , P1_U4935 , P1_U3647 );
nand NAND3_13324 ( P1_U3108 , P1_U4931 , P1_U4930 , P1_U3646 );
nand NAND3_13325 ( P1_U3109 , P1_U4926 , P1_U4925 , P1_U3645 );
nand NAND3_13326 ( P1_U3110 , P1_U4921 , P1_U4920 , P1_U3644 );
nand NAND3_13327 ( P1_U3111 , P1_U4916 , P1_U4915 , P1_U3643 );
nand NAND3_13328 ( P1_U3112 , P1_U4911 , P1_U4910 , P1_U3642 );
nand NAND3_13329 ( P1_U3113 , P1_U4888 , P1_U4887 , P1_U3640 );
nand NAND3_13330 ( P1_U3114 , P1_U4883 , P1_U4882 , P1_U3639 );
nand NAND3_13331 ( P1_U3115 , P1_U4878 , P1_U4877 , P1_U3638 );
nand NAND3_13332 ( P1_U3116 , P1_U4873 , P1_U4872 , P1_U3637 );
nand NAND3_13333 ( P1_U3117 , P1_U4868 , P1_U4867 , P1_U3636 );
nand NAND3_13334 ( P1_U3118 , P1_U4863 , P1_U4862 , P1_U3635 );
nand NAND3_13335 ( P1_U3119 , P1_U4858 , P1_U4857 , P1_U3634 );
nand NAND3_13336 ( P1_U3120 , P1_U4853 , P1_U4852 , P1_U3633 );
nand NAND3_13337 ( P1_U3121 , P1_U4831 , P1_U4830 , P1_U3631 );
nand NAND3_13338 ( P1_U3122 , P1_U4826 , P1_U4825 , P1_U3630 );
nand NAND3_13339 ( P1_U3123 , P1_U4821 , P1_U4820 , P1_U3629 );
nand NAND3_13340 ( P1_U3124 , P1_U4816 , P1_U4815 , P1_U3628 );
nand NAND3_13341 ( P1_U3125 , P1_U4811 , P1_U4810 , P1_U3627 );
nand NAND3_13342 ( P1_U3126 , P1_U4806 , P1_U4805 , P1_U3626 );
nand NAND3_13343 ( P1_U3127 , P1_U4801 , P1_U4800 , P1_U3625 );
nand NAND3_13344 ( P1_U3128 , P1_U4796 , P1_U4795 , P1_U3624 );
nand NAND3_13345 ( P1_U3129 , P1_U4773 , P1_U4772 , P1_U3622 );
nand NAND3_13346 ( P1_U3130 , P1_U4768 , P1_U4767 , P1_U3621 );
nand NAND3_13347 ( P1_U3131 , P1_U4763 , P1_U4762 , P1_U3620 );
nand NAND3_13348 ( P1_U3132 , P1_U4758 , P1_U4757 , P1_U3619 );
nand NAND3_13349 ( P1_U3133 , P1_U4753 , P1_U4752 , P1_U3618 );
nand NAND3_13350 ( P1_U3134 , P1_U4748 , P1_U4747 , P1_U3617 );
nand NAND3_13351 ( P1_U3135 , P1_U4743 , P1_U4742 , P1_U3616 );
nand NAND3_13352 ( P1_U3136 , P1_U4738 , P1_U4737 , P1_U3615 );
nand NAND3_13353 ( P1_U3137 , P1_U4716 , P1_U4715 , P1_U3613 );
nand NAND3_13354 ( P1_U3138 , P1_U4711 , P1_U4710 , P1_U3612 );
nand NAND3_13355 ( P1_U3139 , P1_U4706 , P1_U4705 , P1_U3611 );
nand NAND3_13356 ( P1_U3140 , P1_U4701 , P1_U4700 , P1_U3610 );
nand NAND3_13357 ( P1_U3141 , P1_U4696 , P1_U4695 , P1_U3609 );
nand NAND3_13358 ( P1_U3142 , P1_U4691 , P1_U4690 , P1_U3608 );
nand NAND3_13359 ( P1_U3143 , P1_U4686 , P1_U4685 , P1_U3607 );
nand NAND3_13360 ( P1_U3144 , P1_U4681 , P1_U4680 , P1_U3606 );
nand NAND3_13361 ( P1_U3145 , P1_U4657 , P1_U4656 , P1_U3604 );
nand NAND3_13362 ( P1_U3146 , P1_U4652 , P1_U4651 , P1_U3603 );
nand NAND3_13363 ( P1_U3147 , P1_U4647 , P1_U4646 , P1_U3602 );
nand NAND3_13364 ( P1_U3148 , P1_U4642 , P1_U4641 , P1_U3601 );
nand NAND3_13365 ( P1_U3149 , P1_U4637 , P1_U4636 , P1_U3600 );
nand NAND3_13366 ( P1_U3150 , P1_U4632 , P1_U4631 , P1_U3599 );
nand NAND3_13367 ( P1_U3151 , P1_U4627 , P1_U4626 , P1_U3598 );
nand NAND3_13368 ( P1_U3152 , P1_U4622 , P1_U4621 , P1_U3597 );
nand NAND3_13369 ( P1_U3153 , P1_U4599 , P1_U4598 , P1_U3595 );
nand NAND3_13370 ( P1_U3154 , P1_U4594 , P1_U4593 , P1_U3594 );
nand NAND3_13371 ( P1_U3155 , P1_U4589 , P1_U4588 , P1_U3593 );
nand NAND3_13372 ( P1_U3156 , P1_U4584 , P1_U4583 , P1_U3592 );
nand NAND3_13373 ( P1_U3157 , P1_U4579 , P1_U4578 , P1_U3591 );
nand NAND3_13374 ( P1_U3158 , P1_U4574 , P1_U4573 , P1_U3590 );
nand NAND3_13375 ( P1_U3159 , P1_U4569 , P1_U4568 , P1_U3589 );
nand NAND3_13376 ( P1_U3160 , P1_U4564 , P1_U4563 , P1_U3588 );
nand NAND3_13377 ( P1_U3161 , P1_U7690 , P1_U7689 , P1_U3586 );
nand NAND4_13378 ( P1_U3162 , P1_U4520 , P1_U4519 , P1_U4518 , P1_U4244 );
nand NAND2_13379 ( P1_U3163 , P1_U3582 , P1_U4516 );
and AND2_13380 ( P1_U3164 , P1_DATAWIDTH_REG_31_ , P1_U7650 );
and AND2_13381 ( P1_U3165 , P1_DATAWIDTH_REG_30_ , P1_U7650 );
and AND2_13382 ( P1_U3166 , P1_DATAWIDTH_REG_29_ , P1_U7650 );
and AND2_13383 ( P1_U3167 , P1_DATAWIDTH_REG_28_ , P1_U7650 );
and AND2_13384 ( P1_U3168 , P1_DATAWIDTH_REG_27_ , P1_U7650 );
and AND2_13385 ( P1_U3169 , P1_DATAWIDTH_REG_26_ , P1_U7650 );
and AND2_13386 ( P1_U3170 , P1_DATAWIDTH_REG_25_ , P1_U7650 );
and AND2_13387 ( P1_U3171 , P1_DATAWIDTH_REG_24_ , P1_U7650 );
and AND2_13388 ( P1_U3172 , P1_DATAWIDTH_REG_23_ , P1_U7650 );
and AND2_13389 ( P1_U3173 , P1_DATAWIDTH_REG_22_ , P1_U7650 );
and AND2_13390 ( P1_U3174 , P1_DATAWIDTH_REG_21_ , P1_U7650 );
and AND2_13391 ( P1_U3175 , P1_DATAWIDTH_REG_20_ , P1_U7650 );
and AND2_13392 ( P1_U3176 , P1_DATAWIDTH_REG_19_ , P1_U7650 );
and AND2_13393 ( P1_U3177 , P1_DATAWIDTH_REG_18_ , P1_U7650 );
and AND2_13394 ( P1_U3178 , P1_DATAWIDTH_REG_17_ , P1_U7650 );
and AND2_13395 ( P1_U3179 , P1_DATAWIDTH_REG_16_ , P1_U7650 );
and AND2_13396 ( P1_U3180 , P1_DATAWIDTH_REG_15_ , P1_U7650 );
and AND2_13397 ( P1_U3181 , P1_DATAWIDTH_REG_14_ , P1_U7650 );
and AND2_13398 ( P1_U3182 , P1_DATAWIDTH_REG_13_ , P1_U7650 );
and AND2_13399 ( P1_U3183 , P1_DATAWIDTH_REG_12_ , P1_U7650 );
and AND2_13400 ( P1_U3184 , P1_DATAWIDTH_REG_11_ , P1_U7650 );
and AND2_13401 ( P1_U3185 , P1_DATAWIDTH_REG_10_ , P1_U7650 );
and AND2_13402 ( P1_U3186 , P1_DATAWIDTH_REG_9_ , P1_U7650 );
and AND2_13403 ( P1_U3187 , P1_DATAWIDTH_REG_8_ , P1_U7650 );
and AND2_13404 ( P1_U3188 , P1_DATAWIDTH_REG_7_ , P1_U7650 );
and AND2_13405 ( P1_U3189 , P1_DATAWIDTH_REG_6_ , P1_U7650 );
and AND2_13406 ( P1_U3190 , P1_DATAWIDTH_REG_5_ , P1_U7650 );
and AND2_13407 ( P1_U3191 , P1_DATAWIDTH_REG_4_ , P1_U7650 );
and AND2_13408 ( P1_U3192 , P1_DATAWIDTH_REG_3_ , P1_U7650 );
and AND2_13409 ( P1_U3193 , P1_DATAWIDTH_REG_2_ , P1_U7650 );
nand NAND3_13410 ( P1_U3194 , P1_U7647 , P1_U7646 , P1_U4375 );
nand NAND3_13411 ( P1_U3195 , P1_U7645 , P1_U7644 , P1_U3495 );
nand NAND2_13412 ( P1_U3196 , P1_U3494 , P1_U4369 );
nand NAND3_13413 ( P1_U3197 , P1_U4355 , P1_U4354 , P1_U4356 );
nand NAND3_13414 ( P1_U3198 , P1_U4352 , P1_U4351 , P1_U4353 );
nand NAND3_13415 ( P1_U3199 , P1_U4349 , P1_U4348 , P1_U4350 );
nand NAND3_13416 ( P1_U3200 , P1_U4346 , P1_U4345 , P1_U4347 );
nand NAND3_13417 ( P1_U3201 , P1_U4343 , P1_U4342 , P1_U4344 );
nand NAND3_13418 ( P1_U3202 , P1_U4340 , P1_U4339 , P1_U4341 );
nand NAND3_13419 ( P1_U3203 , P1_U4337 , P1_U4336 , P1_U4338 );
nand NAND3_13420 ( P1_U3204 , P1_U4334 , P1_U4333 , P1_U4335 );
nand NAND3_13421 ( P1_U3205 , P1_U4331 , P1_U4330 , P1_U4332 );
nand NAND3_13422 ( P1_U3206 , P1_U4328 , P1_U4327 , P1_U4329 );
nand NAND3_13423 ( P1_U3207 , P1_U4325 , P1_U4324 , P1_U4326 );
nand NAND3_13424 ( P1_U3208 , P1_U4322 , P1_U4321 , P1_U4323 );
nand NAND3_13425 ( P1_U3209 , P1_U4319 , P1_U4318 , P1_U4320 );
nand NAND3_13426 ( P1_U3210 , P1_U4316 , P1_U4315 , P1_U4317 );
nand NAND3_13427 ( P1_U3211 , P1_U4313 , P1_U4312 , P1_U4314 );
nand NAND3_13428 ( P1_U3212 , P1_U4310 , P1_U4309 , P1_U4311 );
nand NAND3_13429 ( P1_U3213 , P1_U4307 , P1_U4306 , P1_U4308 );
nand NAND3_13430 ( P1_U3214 , P1_U4304 , P1_U4303 , P1_U4305 );
nand NAND3_13431 ( P1_U3215 , P1_U4301 , P1_U4300 , P1_U4302 );
nand NAND3_13432 ( P1_U3216 , P1_U4298 , P1_U4297 , P1_U4299 );
nand NAND3_13433 ( P1_U3217 , P1_U4295 , P1_U4294 , P1_U4296 );
nand NAND3_13434 ( P1_U3218 , P1_U4292 , P1_U4291 , P1_U4293 );
nand NAND3_13435 ( P1_U3219 , P1_U4289 , P1_U4288 , P1_U4290 );
nand NAND3_13436 ( P1_U3220 , P1_U4286 , P1_U4285 , P1_U4287 );
nand NAND3_13437 ( P1_U3221 , P1_U4283 , P1_U4282 , P1_U4284 );
nand NAND3_13438 ( P1_U3222 , P1_U4280 , P1_U4279 , P1_U4281 );
nand NAND3_13439 ( P1_U3223 , P1_U4277 , P1_U4276 , P1_U4278 );
nand NAND3_13440 ( P1_U3224 , P1_U4274 , P1_U4273 , P1_U4275 );
nand NAND3_13441 ( P1_U3225 , P1_U4271 , P1_U4270 , P1_U4272 );
nand NAND3_13442 ( P1_U3226 , P1_U4268 , P1_U4267 , P1_U4269 );
nand NAND4_13443 ( P1_U3227 , P1_U4001 , P1_U4000 , P1_U3999 , P1_U3998 );
nand NAND4_13444 ( P1_U3228 , P1_U3997 , P1_U3996 , P1_U3995 , P1_U3994 );
nand NAND4_13445 ( P1_U3229 , P1_U3993 , P1_U3992 , P1_U3991 , P1_U3990 );
nand NAND4_13446 ( P1_U3230 , P1_U3989 , P1_U3988 , P1_U3987 , P1_U3986 );
nand NAND4_13447 ( P1_U3231 , P1_U3985 , P1_U3984 , P1_U3983 , P1_U3982 );
nand NAND4_13448 ( P1_U3232 , P1_U3981 , P1_U3980 , P1_U3979 , P1_U3978 );
nand NAND4_13449 ( P1_U3233 , P1_U3977 , P1_U3976 , P1_U3975 , P1_U3974 );
nand NAND4_13450 ( P1_U3234 , P1_U3973 , P1_U3972 , P1_U3971 , P1_U3970 );
nand NAND2_13451 ( P1_U3235 , P1_U3329 , P1_U3323 );
nand NAND2_13452 ( P1_U3236 , P1_U2432 , P1_U3235 );
nand NAND2_13453 ( P1_U3237 , P1_U2432 , P1_U4543 );
nand NAND2_13454 ( P1_U3238 , P1_U2434 , P1_U3235 );
nand NAND2_13455 ( P1_U3239 , P1_U2434 , P1_U4543 );
nand NAND2_13456 ( P1_U3240 , P1_U2433 , P1_U3235 );
nand NAND2_13457 ( P1_U3241 , P1_U2433 , P1_U4543 );
nand NAND2_13458 ( P1_U3242 , P1_U2435 , P1_U3235 );
nand NAND2_13459 ( P1_U3243 , P1_U2435 , P1_U4543 );
nand NAND3_13460 ( P1_U3244 , P1_U3391 , P1_U3394 , P1_U5463 );
nand NAND2_13461 ( P1_U3245 , P1_U7086 , P1_U5464 );
nand NAND4_13462 ( P1_U3246 , P1_U7792 , P1_U7791 , P1_U4158 , P1_U4156 );
not NOT1_13463 ( P1_U3247 , P1_REQUESTPENDING_REG );
not NOT1_13464 ( P1_U3248 , P1_STATE_REG_1_ );
nand NAND2_13465 ( P1_U3249 , P1_STATE_REG_1_ , P1_U3258 );
nand NAND2_13466 ( P1_U3250 , P1_U4221 , P1_U3251 );
not NOT1_13467 ( P1_U3251 , P1_STATE_REG_2_ );
nand NAND2_13468 ( P1_U3252 , P1_STATE_REG_2_ , P1_U4221 );
not NOT1_13469 ( P1_U3253 , P1_REIP_REG_1_ );
nand NAND2_13470 ( P1_U3254 , P1_STATE_REG_1_ , P1_U3251 );
or OR2_13471 ( P1_U3255 , P1_STATE_REG_1_ , P1_STATE_REG_2_ );
not NOT1_13472 ( P1_U3256 , HOLD );
not NOT1_13473 ( P1_U3257 , U210 );
not NOT1_13474 ( P1_U3258 , P1_STATE_REG_0_ );
nand NAND2_13475 ( P1_U3259 , P1_STATE_REG_0_ , P1_U3260 );
nand NAND2_13476 ( P1_U3260 , P1_REQUESTPENDING_REG , P1_U3256 );
or OR2_13477 ( P1_U3261 , HOLD , P1_REQUESTPENDING_REG );
not NOT1_13478 ( P1_U3262 , P1_STATE2_REG_1_ );
not NOT1_13479 ( P1_U3263 , P1_STATE2_REG_2_ );
not NOT1_13480 ( P1_U3264 , P1_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_13481 ( P1_U3265 , P1_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_13482 ( P1_U3266 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND4_13483 ( P1_U3267 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3270 );
or OR3_13484 ( P1_U3268 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ );
or OR2_13485 ( P1_U3269 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_0_ );
not NOT1_13486 ( P1_U3270 , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND4_13487 ( P1_U3271 , P1_U3567 , P1_U3566 , P1_U3565 , P1_U3564 );
nand NAND2_13488 ( P1_U3272 , P1_U4496 , P1_U3258 );
not NOT1_13489 ( P1_U3273 , P1_R2167_U17 );
nand NAND2_13490 ( P1_U3274 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3270 );
nand NAND2_13491 ( P1_U3275 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ );
nand NAND4_13492 ( P1_U3276 , P1_U3519 , P1_U3518 , P1_U3517 , P1_U3516 );
nand NAND5_13493 ( P1_U3277 , P1_U3539 , P1_U4170 , P1_U3538 , P1_U3537 , P1_U3536 );
nand NAND4_13494 ( P1_U3278 , P1_U3557 , P1_U3556 , P1_U3555 , P1_U3554 );
nand NAND2_13495 ( P1_U3279 , P1_U3559 , P1_U3558 );
or OR2_13496 ( P1_U3280 , P1_STATEBS16_REG , U210 );
nand NAND2_13497 ( P1_U3281 , P1_R2167_U17 , P1_U4497 );
nand NAND2_13498 ( P1_U3282 , P1_U4477 , P1_U3284 );
nand NAND4_13499 ( P1_U3283 , P1_U3511 , P1_U3510 , P1_U3509 , P1_U3508 );
nand NAND4_13500 ( P1_U3284 , P1_U3563 , P1_U3562 , P1_U3561 , P1_U3560 );
nand NAND2_13501 ( P1_U3285 , P1_U2473 , P1_U4501 );
nand NAND2_13502 ( P1_U3286 , P1_U2389 , P1_U3283 );
nand NAND2_13503 ( P1_U3287 , P1_U4494 , P1_U4477 );
nand NAND2_13504 ( P1_U3288 , P1_U4249 , P1_U2447 );
nand NAND4_13505 ( P1_U3289 , P1_U4460 , P1_U3391 , P1_U4173 , P1_U3278 );
nand NAND2_13506 ( P1_U3290 , P1_U3271 , P1_U3283 );
nand NAND2_13507 ( P1_U3291 , P1_U4190 , P1_U3284 );
nand NAND2_13508 ( P1_U3292 , P1_U4256 , P1_U2431 );
nand NAND5_13509 ( P1_U3293 , P1_U4178 , P1_U4509 , P1_U7626 , P1_U4225 , P1_LT_563_U6 );
not NOT1_13510 ( P1_U3294 , P1_STATE2_REG_0_ );
nand NAND2_13511 ( P1_U3295 , P1_STATE2_REG_0_ , P1_U7604 );
not NOT1_13512 ( P1_U3296 , P1_STATE2_REG_3_ );
nand NAND2_13513 ( P1_U3297 , P1_STATE2_REG_2_ , P1_U3262 );
or OR2_13514 ( P1_U3298 , P1_STATE2_REG_2_ , P1_STATE2_REG_1_ );
nand NAND2_13515 ( P1_U3299 , P1_STATE2_REG_3_ , P1_R2167_U17 );
nand NAND2_13516 ( P1_U3300 , P1_U4547 , P1_U3294 );
not NOT1_13517 ( P1_U3301 , P1_INSTQUEUEWR_ADDR_REG_0_ );
not NOT1_13518 ( P1_U3302 , P1_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_13519 ( P1_U3303 , P1_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_13520 ( P1_U3304 , P1_INSTQUEUEWR_ADDR_REG_2_ );
nand NAND2_13521 ( P1_U3305 , P1_INSTQUEUEWR_ADDR_REG_1_ , P1_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_13522 ( P1_U3306 , P1_U4533 , P1_U2478 );
or OR2_13523 ( P1_U3307 , P1_STATE2_REG_2_ , P1_STATE2_REG_3_ );
not NOT1_13524 ( P1_U3308 , P1_STATEBS16_REG );
not NOT1_13525 ( P1_U3309 , P1_R2144_U43 );
not NOT1_13526 ( P1_U3310 , P1_R2144_U50 );
not NOT1_13527 ( P1_U3311 , P1_R2144_U49 );
not NOT1_13528 ( P1_U3312 , P1_R2144_U8 );
nand NAND2_13529 ( P1_U3313 , P1_R2144_U50 , P1_R2144_U43 );
nand NAND2_13530 ( P1_U3314 , P1_U3332 , P1_U3309 );
nand NAND2_13531 ( P1_U3315 , P1_U4527 , P1_U2475 );
not NOT1_13532 ( P1_U3316 , P1_R2182_U25 );
not NOT1_13533 ( P1_U3317 , P1_R2182_U42 );
not NOT1_13534 ( P1_U3318 , P1_R2182_U34 );
not NOT1_13535 ( P1_U3319 , P1_R2182_U33 );
nand NAND2_13536 ( P1_U3320 , P1_U4209 , P1_U3308 );
nand NAND2_13537 ( P1_U3321 , P1_U3306 , P1_U4535 );
nand NAND2_13538 ( P1_U3322 , P1_U3306 , P1_U4544 );
nand NAND2_13539 ( P1_U3323 , P1_INSTQUEUEWR_ADDR_REG_1_ , P1_U3301 );
nand NAND2_13540 ( P1_U3324 , P1_U4542 , P1_U2478 );
nand NAND2_13541 ( P1_U3325 , P1_R2144_U50 , P1_U3309 );
nand NAND2_13542 ( P1_U3326 , P1_R2144_U43 , P1_U3332 );
nand NAND2_13543 ( P1_U3327 , P1_U4600 , P1_U2475 );
nand NAND2_13544 ( P1_U3328 , P1_U3324 , P1_U4603 );
nand NAND2_13545 ( P1_U3329 , P1_INSTQUEUEWR_ADDR_REG_0_ , P1_U3302 );
nand NAND2_13546 ( P1_U3330 , P1_U4541 , P1_U2478 );
nand NAND2_13547 ( P1_U3331 , P1_R2144_U43 , P1_U3310 );
nand NAND2_13548 ( P1_U3332 , P1_U3325 , P1_U3331 );
nand NAND2_13549 ( P1_U3333 , P1_U4526 , P1_U3309 );
nand NAND2_13550 ( P1_U3334 , P1_U4658 , P1_U2475 );
nand NAND2_13551 ( P1_U3335 , P1_U3330 , P1_U4661 );
nand NAND2_13552 ( P1_U3336 , P1_U3330 , P1_U4663 );
nand NAND2_13553 ( P1_U3337 , P1_U2488 , P1_U2478 );
nand NAND2_13554 ( P1_U3338 , P1_U2485 , P1_U2475 );
nand NAND2_13555 ( P1_U3339 , P1_U3337 , P1_U4719 );
nand NAND2_13556 ( P1_U3340 , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_U3304 );
nand NAND2_13557 ( P1_U3341 , P1_U4538 , P1_U4533 );
nand NAND2_13558 ( P1_U3342 , P1_R2144_U8 , P1_U3311 );
nand NAND2_13559 ( P1_U3343 , P1_U2490 , P1_U4527 );
nand NAND2_13560 ( P1_U3344 , P1_U3341 , P1_U4776 );
nand NAND2_13561 ( P1_U3345 , P1_U3341 , P1_U4778 );
nand NAND2_13562 ( P1_U3346 , P1_U4538 , P1_U4542 );
nand NAND2_13563 ( P1_U3347 , P1_U2490 , P1_U4600 );
nand NAND2_13564 ( P1_U3348 , P1_U3346 , P1_U4834 );
nand NAND2_13565 ( P1_U3349 , P1_U4538 , P1_U4541 );
nand NAND2_13566 ( P1_U3350 , P1_U2490 , P1_U4658 );
nand NAND2_13567 ( P1_U3351 , P1_U3349 , P1_U4891 );
nand NAND2_13568 ( P1_U3352 , P1_U3349 , P1_U4893 );
nand NAND2_13569 ( P1_U3353 , P1_U4538 , P1_U2488 );
nand NAND2_13570 ( P1_U3354 , P1_U2490 , P1_U2485 );
nand NAND2_13571 ( P1_U3355 , P1_U3353 , P1_U4949 );
nand NAND2_13572 ( P1_U3356 , P1_U2479 , P1_U4533 );
nand NAND2_13573 ( P1_U3357 , P1_U2474 , P1_U4528 );
nand NAND3_13574 ( P1_U3358 , P1_U3342 , P1_U4530 , P1_U3357 );
nand NAND2_13575 ( P1_U3359 , P1_U2499 , P1_U4527 );
nand NAND3_13576 ( P1_U3360 , P1_U3340 , P1_U4539 , P1_U3356 );
nand NAND2_13577 ( P1_U3361 , P1_U3356 , P1_U5005 );
nand NAND2_13578 ( P1_U3362 , P1_U3356 , P1_U5007 );
nand NAND2_13579 ( P1_U3363 , P1_U4542 , P1_U2479 );
nand NAND2_13580 ( P1_U3364 , P1_U2499 , P1_U4600 );
nand NAND2_13581 ( P1_U3365 , P1_U3363 , P1_U5062 );
nand NAND2_13582 ( P1_U3366 , P1_U4541 , P1_U2479 );
nand NAND2_13583 ( P1_U3367 , P1_U2499 , P1_U4658 );
nand NAND2_13584 ( P1_U3368 , P1_U3366 , P1_U5119 );
nand NAND2_13585 ( P1_U3369 , P1_U3366 , P1_U5121 );
nand NAND2_13586 ( P1_U3370 , P1_U2488 , P1_U2479 );
nand NAND2_13587 ( P1_U3371 , P1_U2499 , P1_U2485 );
nand NAND2_13588 ( P1_U3372 , P1_U3370 , P1_U5177 );
nand NAND2_13589 ( P1_U3373 , P1_U2510 , P1_U4533 );
nand NAND2_13590 ( P1_U3374 , P1_U2507 , P1_U4527 );
nand NAND2_13591 ( P1_U3375 , P1_U3373 , P1_U5234 );
nand NAND2_13592 ( P1_U3376 , P1_U3373 , P1_U5236 );
nand NAND2_13593 ( P1_U3377 , P1_U2510 , P1_U4542 );
nand NAND2_13594 ( P1_U3378 , P1_U2507 , P1_U4600 );
nand NAND2_13595 ( P1_U3379 , P1_U3377 , P1_U5292 );
nand NAND2_13596 ( P1_U3380 , P1_U2510 , P1_U4541 );
nand NAND2_13597 ( P1_U3381 , P1_U2507 , P1_U4658 );
nand NAND2_13598 ( P1_U3382 , P1_U3380 , P1_U5349 );
nand NAND2_13599 ( P1_U3383 , P1_U3380 , P1_U5351 );
nand NAND2_13600 ( P1_U3384 , P1_U2510 , P1_U2488 );
nand NAND2_13601 ( P1_U3385 , P1_U2507 , P1_U2485 );
nand NAND2_13602 ( P1_U3386 , P1_U3384 , P1_U5407 );
not NOT1_13603 ( P1_U3387 , P1_FLUSH_REG );
not NOT1_13604 ( P1_U3388 , P1_GTE_485_U6 );
nand NAND2_13605 ( P1_U3389 , P1_U3284 , P1_U3278 );
nand NAND2_13606 ( P1_U3390 , P1_U3284 , P1_U3271 );
nand NAND4_13607 ( P1_U3391 , P1_U3515 , P1_U3514 , P1_U3513 , P1_U3512 );
nand NAND3_13608 ( P1_U3392 , P1_U5490 , P1_U5489 , P1_U7628 );
nand NAND2_13609 ( P1_U3393 , P1_U4399 , P1_U3284 );
nand NAND2_13610 ( P1_U3394 , P1_U2605 , P1_U3277 );
nand NAND3_13611 ( P1_U3395 , P1_U4399 , P1_U7494 , P1_U4494 );
nand NAND2_13612 ( P1_U3396 , P1_U3741 , P1_U4247 );
nand NAND5_13613 ( P1_U3397 , P1_U7494 , P1_U4477 , P1_U2605 , P1_U4494 , P1_U4399 );
nand NAND5_13614 ( P1_U3398 , P1_U2605 , P1_U4460 , P1_U4171 , P1_U4449 , P1_U4400 );
nand NAND3_13615 ( P1_U3399 , P1_U4199 , P1_U4477 , P1_U4234 );
nand NAND2_13616 ( P1_U3400 , P1_U2449 , P1_U2447 );
nand NAND2_13617 ( P1_U3401 , P1_U3444 , P1_U5510 );
nand NAND2_13618 ( P1_U3402 , P1_U3269 , P1_U3275 );
not NOT1_13619 ( P1_U3403 , P1_LT_589_U6 );
nand NAND3_13620 ( P1_U3404 , P1_U4242 , P1_U3300 , P1_U5536 );
nand NAND3_13621 ( P1_U3405 , P1_STATE2_REG_0_ , P1_U3278 , P1_U3284 );
nand NAND2_13622 ( P1_U3406 , P1_U3271 , P1_U3273 );
nand NAND2_13623 ( P1_U3407 , P1_U3277 , P1_U3391 );
nand NAND2_13624 ( P1_U3408 , P1_U2427 , P1_U3294 );
nand NAND2_13625 ( P1_U3409 , P1_U4460 , P1_U3391 );
nand NAND2_13626 ( P1_U3410 , P1_U4253 , P1_U3278 );
nand NAND2_13627 ( P1_U3411 , P1_U4190 , P1_U2452 );
nand NAND2_13628 ( P1_U3412 , P1_STATE2_REG_2_ , P1_U3271 );
not NOT1_13629 ( P1_U3413 , P1_REIP_REG_0_ );
nand NAND2_13630 ( P1_U3414 , P1_U3756 , P1_U5562 );
nand NAND2_13631 ( P1_U3415 , P1_U4400 , P1_U4173 );
nand NAND2_13632 ( P1_U3416 , P1_U3863 , P1_U4248 );
nand NAND2_13633 ( P1_U3417 , P1_U6054 , P1_U6053 );
nand NAND2_13634 ( P1_U3418 , P1_STATE2_REG_0_ , P1_U4494 );
nand NAND2_13635 ( P1_U3419 , P1_U4399 , P1_U7494 );
nand NAND2_13636 ( P1_U3420 , P1_U4206 , P1_U4477 );
nand NAND2_13637 ( P1_U3421 , P1_U4194 , P1_U2431 );
nand NAND2_13638 ( P1_U3422 , P1_U4210 , P1_STATE2_REG_0_ );
nand NAND2_13639 ( P1_U3423 , P1_U4503 , P1_U3391 );
nand NAND2_13640 ( P1_U3424 , P1_U4235 , P1_U6153 );
nand NAND2_13641 ( P1_U3425 , P1_STATE2_REG_0_ , P1_U4216 );
nand NAND2_13642 ( P1_U3426 , P1_U4235 , P1_U6264 );
nand NAND4_13643 ( P1_U3427 , P1_STATE2_REG_0_ , P1_U4249 , P1_U3886 , P1_U2452 );
nand NAND2_13644 ( P1_U3428 , P1_U3866 , P1_U2447 );
not NOT1_13645 ( P1_U3429 , P1_EBX_REG_31_ );
not NOT1_13646 ( P1_U3430 , P1_R2337_U69 );
nand NAND2_13647 ( P1_U3431 , P1_U4228 , P1_U3887 );
nand NAND2_13648 ( P1_U3432 , P1_U4209 , P1_U3262 );
nand NAND4_13649 ( P1_U3433 , P1_U3962 , P1_U3958 , P1_U3955 , P1_U3952 );
nand NAND2_13650 ( P1_U3434 , P1_U4206 , P1_U3271 );
not NOT1_13651 ( P1_U3435 , P1_CODEFETCH_REG );
not NOT1_13652 ( P1_U3436 , P1_READREQUEST_REG );
nand NAND2_13653 ( P1_U3437 , P1_U2447 , P1_U4498 );
nand NAND2_13654 ( P1_U3438 , P1_U3267 , P1_U5482 );
nand NAND2_13655 ( P1_U3439 , P1_U4449 , P1_STATE2_REG_2_ );
nand NAND2_13656 ( P1_U3440 , P1_STATEBS16_REG , P1_U3263 );
not NOT1_13657 ( P1_U3441 , P1_U3234 );
nand NAND2_13658 ( P1_U3442 , P1_U5479 , P1_U5478 );
nand NAND2_13659 ( P1_U3443 , P1_U2450 , P1_U3441 );
nand NAND3_13660 ( P1_U3444 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3264 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_13661 ( P1_U3445 , P1_U3274 , P1_U7064 );
nand NAND2_13662 ( P1_U3446 , P1_U4197 , P1_U4234 );
nand NAND3_13663 ( P1_U3447 , P1_U4231 , P1_U4400 , P1_U4250 );
nand NAND3_13664 ( P1_U3448 , P1_U4231 , P1_U3278 , P1_U4250 );
nand NAND2_13665 ( P1_U3449 , P1_U4477 , P1_U4496 );
nand NAND4_13666 ( P1_U3450 , P1_U4074 , P1_U7093 , P1_U4075 , P1_U4077 );
nand NAND2_13667 ( P1_U3451 , P1_U4254 , P1_U4266 );
nand NAND2_13668 ( P1_U3452 , P1_U4183 , P1_U3268 );
nand NAND2_13669 ( P1_U3453 , P1_STATE2_REG_0_ , P1_U2605 );
nand NAND2_13670 ( P1_U3454 , P1_U7692 , P1_U7691 );
nand NAND2_13671 ( P1_U3455 , P1_U7695 , P1_U7694 );
nand NAND2_13672 ( P1_U3456 , P1_U7719 , P1_U7718 );
nand NAND2_13673 ( P1_U3457 , P1_U7789 , P1_U7788 );
nand NAND2_13674 ( P1_U3458 , P1_U7634 , P1_U7633 );
nand NAND2_13675 ( P1_U3459 , P1_U7636 , P1_U7635 );
nand NAND2_13676 ( P1_U3460 , P1_U7638 , P1_U7637 );
nand NAND2_13677 ( P1_U3461 , P1_U7640 , P1_U7639 );
nand NAND2_13678 ( P1_U3462 , P1_U7649 , P1_U7648 );
and AND2_13679 ( P1_U3463 , P1_U3255 , P1_U4179 );
nand NAND2_13680 ( P1_U3464 , P1_U7652 , P1_U7651 );
nand NAND2_13681 ( P1_U3465 , P1_U7654 , P1_U7653 );
nand NAND2_13682 ( P1_U3466 , P1_U7686 , P1_U7685 );
and AND3_13683 ( P1_U3467 , P1_U2427 , P1_U4215 , P1_R2182_U24 );
nand NAND2_13684 ( P1_U3468 , P1_U7702 , P1_U7701 );
nand NAND2_13685 ( P1_U3469 , P1_U7709 , P1_U7708 );
nand NAND2_13686 ( P1_U3470 , P1_U7711 , P1_U7710 );
nand NAND2_13687 ( P1_U3471 , P1_U7714 , P1_U7713 );
nand NAND2_13688 ( P1_U3472 , P1_U7722 , P1_U7721 );
nand NAND2_13689 ( P1_U3473 , P1_U7724 , P1_U7723 );
nand NAND2_13690 ( P1_U3474 , P1_U7728 , P1_U7727 );
nand NAND2_13691 ( P1_U3475 , P1_U7730 , P1_U7729 );
nand NAND2_13692 ( P1_U3476 , P1_U7735 , P1_U7734 );
nand NAND2_13693 ( P1_U3477 , P1_U7737 , P1_U7736 );
nand NAND2_13694 ( P1_U3478 , P1_U7739 , P1_U7738 );
and AND2_13695 ( P1_U3479 , P1_R2358_U22 , P1_U4449 );
nor nor_13696 ( P1_U3480 , P1_DATAWIDTH_REG_1_ , P1_REIP_REG_1_ );
nand NAND2_13697 ( P1_U3481 , P1_U7755 , P1_U7754 );
nand NAND2_13698 ( P1_U3482 , P1_U7759 , P1_U7758 );
nand NAND2_13699 ( P1_U3483 , P1_U7761 , P1_U7760 );
nand NAND2_13700 ( P1_U3484 , P1_U7763 , P1_U7762 );
nand NAND2_13701 ( P1_U3485 , P1_U7767 , P1_U7766 );
nand NAND2_13702 ( P1_U3486 , P1_U7771 , P1_U7770 );
nand NAND2_13703 ( P1_U3487 , P1_U7773 , P1_U7772 );
and AND2_13704 ( P1_U3488 , P1_R2182_U24 , P1_U4215 );
nand NAND2_13705 ( P1_U3489 , P1_U7775 , P1_U7774 );
nand NAND2_13706 ( P1_U3490 , P1_U7777 , P1_U7776 );
nand NAND2_13707 ( P1_U3491 , P1_U7779 , P1_U7778 );
nand NAND2_13708 ( P1_U3492 , P1_U7781 , P1_U7780 );
nand NAND2_13709 ( P1_U3493 , P1_U7783 , P1_U7782 );
and AND2_13710 ( P1_U3494 , P1_U4368 , P1_U3252 );
and AND2_13711 ( P1_U3495 , P1_U4370 , P1_U3250 );
and AND2_13712 ( P1_U3496 , P1_REQUESTPENDING_REG , P1_STATE_REG_0_ );
nor nor_13713 ( P1_U3497 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_INSTQUEUERD_ADDR_REG_3_ );
and AND2_13714 ( P1_U3498 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ );
nor nor_13715 ( P1_U3499 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_3_ );
and AND2_13716 ( P1_U3500 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_2_ );
nor nor_13717 ( P1_U3501 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_3_ );
and AND2_13718 ( P1_U3502 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ );
nor nor_13719 ( P1_U3503 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_13720 ( P1_U3504 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_0_ );
nor nor_13721 ( P1_U3505 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_13722 ( P1_U3506 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_1_ );
and AND2_13723 ( P1_U3507 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND4_13724 ( P1_U3508 , P1_U4386 , P1_U4385 , P1_U4384 , P1_U4383 );
and AND4_13725 ( P1_U3509 , P1_U4390 , P1_U4389 , P1_U4388 , P1_U4387 );
and AND4_13726 ( P1_U3510 , P1_U4394 , P1_U4393 , P1_U4392 , P1_U4391 );
and AND4_13727 ( P1_U3511 , P1_U4398 , P1_U4397 , P1_U4396 , P1_U4395 );
and AND4_13728 ( P1_U3512 , P1_U4436 , P1_U4435 , P1_U4434 , P1_U4433 );
and AND4_13729 ( P1_U3513 , P1_U4440 , P1_U4439 , P1_U4438 , P1_U4437 );
and AND4_13730 ( P1_U3514 , P1_U4444 , P1_U4443 , P1_U4442 , P1_U4441 );
and AND4_13731 ( P1_U3515 , P1_U4448 , P1_U4447 , P1_U4446 , P1_U4445 );
and AND4_13732 ( P1_U3516 , P1_U4419 , P1_U4418 , P1_U4417 , P1_U4416 );
and AND4_13733 ( P1_U3517 , P1_U4423 , P1_U4422 , P1_U4421 , P1_U4420 );
and AND4_13734 ( P1_U3518 , P1_U4427 , P1_U4426 , P1_U4425 , P1_U4424 );
and AND4_13735 ( P1_U3519 , P1_U4431 , P1_U4430 , P1_U4429 , P1_U4428 );
nor nor_13736 ( P1_U3520 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_3_ );
and AND2_13737 ( P1_U3521 , P1_INSTQUEUE_REG_5__5_ , P1_INSTQUEUERD_ADDR_REG_0_ );
nor nor_13738 ( P1_U3522 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_3_ );
and AND2_13739 ( P1_U3523 , P1_INSTQUEUE_REG_6__5_ , P1_INSTQUEUERD_ADDR_REG_1_ );
and AND2_13740 ( P1_U3524 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUE_REG_8__5_ );
nor nor_13741 ( P1_U3525 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_13742 ( P1_U3526 , P1_INSTQUEUE_REG_10__5_ , P1_INSTQUEUERD_ADDR_REG_3_ );
and AND2_13743 ( P1_U3527 , P1_INSTQUEUE_REG_12__5_ , P1_INSTQUEUERD_ADDR_REG_3_ );
nor nor_13744 ( P1_U3528 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_13745 ( P1_U3529 , P1_INSTQUEUE_REG_9__5_ , P1_INSTQUEUERD_ADDR_REG_0_ );
and AND4_13746 ( P1_U3530 , P1_U4404 , P1_U4403 , P1_U4402 , P1_U4401 );
and AND4_13747 ( P1_U3531 , P1_U4408 , P1_U4407 , P1_U4406 , P1_U4405 );
and AND4_13748 ( P1_U3532 , P1_U4412 , P1_U4411 , P1_U4410 , P1_U4409 );
and AND2_13749 ( P1_U3533 , P1_U4414 , P1_U4413 );
nor nor_13750 ( P1_U3534 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_INSTQUEUERD_ADDR_REG_3_ );
and AND2_13751 ( P1_U3535 , P1_INSTQUEUE_REG_3__6_ , P1_INSTQUEUERD_ADDR_REG_0_ );
and AND4_13752 ( P1_U3536 , P1_U4453 , P1_U4452 , P1_U4451 , P1_U4450 );
and AND3_13753 ( P1_U3537 , P1_U4455 , P1_U4454 , P1_U4456 );
and AND3_13754 ( P1_U3538 , P1_U4458 , P1_U4457 , P1_U4459 );
and AND4_13755 ( P1_U3539 , P1_U7678 , P1_U7677 , P1_U7676 , P1_U7675 );
nor nor_13756 ( P1_U3540 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_INSTQUEUERD_ADDR_REG_3_ );
and AND2_13757 ( P1_U3541 , P1_INSTQUEUE_REG_1__4_ , P1_INSTQUEUERD_ADDR_REG_0_ );
nor nor_13758 ( P1_U3542 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ );
and AND2_13759 ( P1_U3543 , P1_INSTQUEUE_REG_4__4_ , P1_INSTQUEUERD_ADDR_REG_2_ );
nor nor_13760 ( P1_U3544 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ );
and AND2_13761 ( P1_U3545 , P1_INSTQUEUE_REG_12__4_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_13762 ( P1_U3546 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_13763 ( P1_U3547 , P1_INSTQUEUE_REG_13__4_ , P1_INSTQUEUERD_ADDR_REG_3_ );
nor nor_13764 ( P1_U3548 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_3_ );
and AND2_13765 ( P1_U3549 , P1_INSTQUEUE_REG_6__4_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_13766 ( P1_U3550 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_13767 ( P1_U3551 , P1_INSTQUEUE_REG_14__4_ , P1_INSTQUEUERD_ADDR_REG_3_ );
nor nor_13768 ( P1_U3552 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ );
and AND2_13769 ( P1_U3553 , P1_INSTQUEUE_REG_9__4_ , P1_INSTQUEUERD_ADDR_REG_3_ );
and AND4_13770 ( P1_U3554 , P1_U7658 , P1_U7657 , P1_U7656 , P1_U7655 );
and AND4_13771 ( P1_U3555 , P1_U7662 , P1_U7661 , P1_U7660 , P1_U7659 );
and AND4_13772 ( P1_U3556 , P1_U7666 , P1_U7665 , P1_U7664 , P1_U7663 );
and AND4_13773 ( P1_U3557 , P1_U7670 , P1_U7669 , P1_U7668 , P1_U7667 );
and AND3_13774 ( P1_U3558 , P1_U3391 , P1_U3283 , P1_U7494 );
and AND3_13775 ( P1_U3559 , P1_U4460 , P1_U2605 , P1_U4400 );
and AND4_13776 ( P1_U3560 , P1_U4481 , P1_U4480 , P1_U4479 , P1_U4478 );
and AND4_13777 ( P1_U3561 , P1_U4485 , P1_U4484 , P1_U4483 , P1_U4482 );
and AND4_13778 ( P1_U3562 , P1_U4489 , P1_U4488 , P1_U4487 , P1_U4486 );
and AND4_13779 ( P1_U3563 , P1_U4493 , P1_U4492 , P1_U4491 , P1_U4490 );
and AND4_13780 ( P1_U3564 , P1_U4464 , P1_U4463 , P1_U4462 , P1_U4461 );
and AND4_13781 ( P1_U3565 , P1_U4468 , P1_U4467 , P1_U4466 , P1_U4465 );
and AND4_13782 ( P1_U3566 , P1_U4472 , P1_U4471 , P1_U4470 , P1_U4469 );
and AND4_13783 ( P1_U3567 , P1_U4476 , P1_U4475 , P1_U4474 , P1_U4473 );
and AND2_13784 ( P1_U3568 , P1_U4377 , P1_U4208 );
and AND4_13785 ( P1_U3569 , P1_U4419 , P1_U4418 , P1_U4417 , P1_U4416 );
and AND4_13786 ( P1_U3570 , P1_U4423 , P1_U4422 , P1_U4421 , P1_U4420 );
and AND4_13787 ( P1_U3571 , P1_U4427 , P1_U4426 , P1_U4425 , P1_U4424 );
and AND4_13788 ( P1_U3572 , P1_U4431 , P1_U4430 , P1_U4429 , P1_U4428 );
and AND4_13789 ( P1_U3573 , P1_U4404 , P1_U4403 , P1_U4402 , P1_U4401 );
and AND4_13790 ( P1_U3574 , P1_U4408 , P1_U4407 , P1_U4406 , P1_U4405 );
and AND4_13791 ( P1_U3575 , P1_U4412 , P1_U4411 , P1_U4410 , P1_U4409 );
and AND2_13792 ( P1_U3576 , P1_U4414 , P1_U4413 );
and AND2_13793 ( P1_U3577 , P1_U4399 , P1_U4171 );
and AND2_13794 ( P1_U3578 , P1_U4249 , P1_U3283 );
and AND4_13795 ( P1_U3579 , P1_U3284 , P1_U3283 , P1_U4400 , P1_U7494 );
and AND2_13796 ( P1_U3580 , P1_U4217 , P1_U3400 );
and AND2_13797 ( P1_U3581 , P1_STATE2_REG_2_ , P1_U7603 );
and AND2_13798 ( P1_U3582 , P1_U4515 , P1_U3297 );
and AND2_13799 ( P1_U3583 , P1_U2427 , P1_U3257 );
and AND2_13800 ( P1_U3584 , P1_STATE2_REG_3_ , P1_STATE2_REG_0_ );
and AND2_13801 ( P1_U3585 , P1_U4246 , P1_U4241 );
and AND2_13802 ( P1_U3586 , P1_U3585 , P1_U4523 );
and AND3_13803 ( P1_U3587 , P1_U4552 , P1_U4553 , P1_U4224 );
and AND3_13804 ( P1_U3588 , P1_U4561 , P1_U4560 , P1_U4562 );
and AND3_13805 ( P1_U3589 , P1_U4566 , P1_U4565 , P1_U4567 );
and AND3_13806 ( P1_U3590 , P1_U4571 , P1_U4570 , P1_U4572 );
and AND3_13807 ( P1_U3591 , P1_U4576 , P1_U4575 , P1_U4577 );
and AND3_13808 ( P1_U3592 , P1_U4581 , P1_U4580 , P1_U4582 );
and AND3_13809 ( P1_U3593 , P1_U4586 , P1_U4585 , P1_U4587 );
and AND3_13810 ( P1_U3594 , P1_U4591 , P1_U4590 , P1_U4592 );
and AND3_13811 ( P1_U3595 , P1_U4596 , P1_U4595 , P1_U4597 );
and AND3_13812 ( P1_U3596 , P1_U4610 , P1_U4611 , P1_U4224 );
and AND3_13813 ( P1_U3597 , P1_U4619 , P1_U4618 , P1_U4620 );
and AND3_13814 ( P1_U3598 , P1_U4624 , P1_U4623 , P1_U4625 );
and AND3_13815 ( P1_U3599 , P1_U4629 , P1_U4628 , P1_U4630 );
and AND3_13816 ( P1_U3600 , P1_U4634 , P1_U4633 , P1_U4635 );
and AND3_13817 ( P1_U3601 , P1_U4639 , P1_U4638 , P1_U4640 );
and AND3_13818 ( P1_U3602 , P1_U4644 , P1_U4643 , P1_U4645 );
and AND3_13819 ( P1_U3603 , P1_U4649 , P1_U4648 , P1_U4650 );
and AND3_13820 ( P1_U3604 , P1_U4654 , P1_U4653 , P1_U4655 );
and AND3_13821 ( P1_U3605 , P1_U4669 , P1_U4670 , P1_U4224 );
and AND3_13822 ( P1_U3606 , P1_U4678 , P1_U4677 , P1_U4679 );
and AND3_13823 ( P1_U3607 , P1_U4683 , P1_U4682 , P1_U4684 );
and AND3_13824 ( P1_U3608 , P1_U4688 , P1_U4687 , P1_U4689 );
and AND3_13825 ( P1_U3609 , P1_U4693 , P1_U4692 , P1_U4694 );
and AND3_13826 ( P1_U3610 , P1_U4698 , P1_U4697 , P1_U4699 );
and AND3_13827 ( P1_U3611 , P1_U4703 , P1_U4702 , P1_U4704 );
and AND3_13828 ( P1_U3612 , P1_U4708 , P1_U4707 , P1_U4709 );
and AND3_13829 ( P1_U3613 , P1_U4713 , P1_U4712 , P1_U4714 );
and AND3_13830 ( P1_U3614 , P1_U4726 , P1_U4727 , P1_U4224 );
and AND3_13831 ( P1_U3615 , P1_U4735 , P1_U4734 , P1_U4736 );
and AND3_13832 ( P1_U3616 , P1_U4740 , P1_U4739 , P1_U4741 );
and AND3_13833 ( P1_U3617 , P1_U4745 , P1_U4744 , P1_U4746 );
and AND3_13834 ( P1_U3618 , P1_U4750 , P1_U4749 , P1_U4751 );
and AND3_13835 ( P1_U3619 , P1_U4755 , P1_U4754 , P1_U4756 );
and AND3_13836 ( P1_U3620 , P1_U4760 , P1_U4759 , P1_U4761 );
and AND3_13837 ( P1_U3621 , P1_U4765 , P1_U4764 , P1_U4766 );
and AND3_13838 ( P1_U3622 , P1_U4770 , P1_U4769 , P1_U4771 );
and AND3_13839 ( P1_U3623 , P1_U4784 , P1_U4785 , P1_U4224 );
and AND3_13840 ( P1_U3624 , P1_U4793 , P1_U4792 , P1_U4794 );
and AND3_13841 ( P1_U3625 , P1_U4798 , P1_U4797 , P1_U4799 );
and AND3_13842 ( P1_U3626 , P1_U4803 , P1_U4802 , P1_U4804 );
and AND3_13843 ( P1_U3627 , P1_U4808 , P1_U4807 , P1_U4809 );
and AND3_13844 ( P1_U3628 , P1_U4813 , P1_U4812 , P1_U4814 );
and AND3_13845 ( P1_U3629 , P1_U4818 , P1_U4817 , P1_U4819 );
and AND3_13846 ( P1_U3630 , P1_U4823 , P1_U4822 , P1_U4824 );
and AND3_13847 ( P1_U3631 , P1_U4828 , P1_U4827 , P1_U4829 );
and AND3_13848 ( P1_U3632 , P1_U4841 , P1_U4842 , P1_U4224 );
and AND3_13849 ( P1_U3633 , P1_U4850 , P1_U4849 , P1_U4851 );
and AND3_13850 ( P1_U3634 , P1_U4855 , P1_U4854 , P1_U4856 );
and AND3_13851 ( P1_U3635 , P1_U4860 , P1_U4859 , P1_U4861 );
and AND3_13852 ( P1_U3636 , P1_U4865 , P1_U4864 , P1_U4866 );
and AND3_13853 ( P1_U3637 , P1_U4870 , P1_U4869 , P1_U4871 );
and AND3_13854 ( P1_U3638 , P1_U4875 , P1_U4874 , P1_U4876 );
and AND3_13855 ( P1_U3639 , P1_U4880 , P1_U4879 , P1_U4881 );
and AND3_13856 ( P1_U3640 , P1_U4885 , P1_U4884 , P1_U4886 );
and AND3_13857 ( P1_U3641 , P1_U4899 , P1_U4900 , P1_U4224 );
and AND3_13858 ( P1_U3642 , P1_U4908 , P1_U4907 , P1_U4909 );
and AND3_13859 ( P1_U3643 , P1_U4913 , P1_U4912 , P1_U4914 );
and AND3_13860 ( P1_U3644 , P1_U4918 , P1_U4917 , P1_U4919 );
and AND3_13861 ( P1_U3645 , P1_U4923 , P1_U4922 , P1_U4924 );
and AND3_13862 ( P1_U3646 , P1_U4928 , P1_U4927 , P1_U4929 );
and AND3_13863 ( P1_U3647 , P1_U4933 , P1_U4932 , P1_U4934 );
and AND3_13864 ( P1_U3648 , P1_U4938 , P1_U4937 , P1_U4939 );
and AND3_13865 ( P1_U3649 , P1_U4943 , P1_U4942 , P1_U4944 );
and AND3_13866 ( P1_U3650 , P1_U4956 , P1_U4957 , P1_U4224 );
and AND3_13867 ( P1_U3651 , P1_U4965 , P1_U4964 , P1_U4966 );
and AND3_13868 ( P1_U3652 , P1_U4970 , P1_U4969 , P1_U4971 );
and AND3_13869 ( P1_U3653 , P1_U4975 , P1_U4974 , P1_U4976 );
and AND3_13870 ( P1_U3654 , P1_U4980 , P1_U4979 , P1_U4981 );
and AND3_13871 ( P1_U3655 , P1_U4985 , P1_U4984 , P1_U4986 );
and AND3_13872 ( P1_U3656 , P1_U4990 , P1_U4989 , P1_U4991 );
and AND3_13873 ( P1_U3657 , P1_U4995 , P1_U4994 , P1_U4996 );
and AND3_13874 ( P1_U3658 , P1_U5000 , P1_U4999 , P1_U5001 );
and AND3_13875 ( P1_U3659 , P1_U5012 , P1_U5013 , P1_U4224 );
and AND3_13876 ( P1_U3660 , P1_U5021 , P1_U5020 , P1_U5022 );
and AND3_13877 ( P1_U3661 , P1_U5026 , P1_U5025 , P1_U5027 );
and AND3_13878 ( P1_U3662 , P1_U5031 , P1_U5030 , P1_U5032 );
and AND3_13879 ( P1_U3663 , P1_U5036 , P1_U5035 , P1_U5037 );
and AND3_13880 ( P1_U3664 , P1_U5041 , P1_U5040 , P1_U5042 );
and AND3_13881 ( P1_U3665 , P1_U5046 , P1_U5045 , P1_U5047 );
and AND3_13882 ( P1_U3666 , P1_U5051 , P1_U5050 , P1_U5052 );
and AND3_13883 ( P1_U3667 , P1_U5056 , P1_U5055 , P1_U5057 );
and AND3_13884 ( P1_U3668 , P1_U5069 , P1_U5070 , P1_U4224 );
and AND3_13885 ( P1_U3669 , P1_U5078 , P1_U5077 , P1_U5079 );
and AND3_13886 ( P1_U3670 , P1_U5083 , P1_U5082 , P1_U5084 );
and AND3_13887 ( P1_U3671 , P1_U5088 , P1_U5087 , P1_U5089 );
and AND3_13888 ( P1_U3672 , P1_U5093 , P1_U5092 , P1_U5094 );
and AND3_13889 ( P1_U3673 , P1_U5098 , P1_U5097 , P1_U5099 );
and AND3_13890 ( P1_U3674 , P1_U5103 , P1_U5102 , P1_U5104 );
and AND3_13891 ( P1_U3675 , P1_U5108 , P1_U5107 , P1_U5109 );
and AND3_13892 ( P1_U3676 , P1_U5113 , P1_U5112 , P1_U5114 );
and AND3_13893 ( P1_U3677 , P1_U5127 , P1_U5128 , P1_U4224 );
and AND3_13894 ( P1_U3678 , P1_U5136 , P1_U5135 , P1_U5137 );
and AND3_13895 ( P1_U3679 , P1_U5141 , P1_U5140 , P1_U5142 );
and AND3_13896 ( P1_U3680 , P1_U5146 , P1_U5145 , P1_U5147 );
and AND3_13897 ( P1_U3681 , P1_U5151 , P1_U5150 , P1_U5152 );
and AND3_13898 ( P1_U3682 , P1_U5156 , P1_U5155 , P1_U5157 );
and AND3_13899 ( P1_U3683 , P1_U5161 , P1_U5160 , P1_U5162 );
and AND3_13900 ( P1_U3684 , P1_U5166 , P1_U5165 , P1_U5167 );
and AND3_13901 ( P1_U3685 , P1_U5171 , P1_U5170 , P1_U5172 );
and AND3_13902 ( P1_U3686 , P1_U5184 , P1_U5185 , P1_U4224 );
and AND3_13903 ( P1_U3687 , P1_U5193 , P1_U5192 , P1_U5194 );
and AND3_13904 ( P1_U3688 , P1_U5198 , P1_U5197 , P1_U5199 );
and AND3_13905 ( P1_U3689 , P1_U5203 , P1_U5202 , P1_U5204 );
and AND3_13906 ( P1_U3690 , P1_U5208 , P1_U5207 , P1_U5209 );
and AND3_13907 ( P1_U3691 , P1_U5213 , P1_U5212 , P1_U5214 );
and AND3_13908 ( P1_U3692 , P1_U5218 , P1_U5217 , P1_U5219 );
and AND3_13909 ( P1_U3693 , P1_U5223 , P1_U5222 , P1_U5224 );
and AND3_13910 ( P1_U3694 , P1_U5228 , P1_U5227 , P1_U5229 );
and AND3_13911 ( P1_U3695 , P1_U5242 , P1_U5243 , P1_U4224 );
and AND3_13912 ( P1_U3696 , P1_U5251 , P1_U5250 , P1_U5252 );
and AND3_13913 ( P1_U3697 , P1_U5256 , P1_U5255 , P1_U5257 );
and AND3_13914 ( P1_U3698 , P1_U5261 , P1_U5260 , P1_U5262 );
and AND3_13915 ( P1_U3699 , P1_U5266 , P1_U5265 , P1_U5267 );
and AND3_13916 ( P1_U3700 , P1_U5271 , P1_U5270 , P1_U5272 );
and AND3_13917 ( P1_U3701 , P1_U5276 , P1_U5275 , P1_U5277 );
and AND3_13918 ( P1_U3702 , P1_U5281 , P1_U5280 , P1_U5282 );
and AND3_13919 ( P1_U3703 , P1_U5286 , P1_U5285 , P1_U5287 );
and AND3_13920 ( P1_U3704 , P1_U5299 , P1_U5300 , P1_U4224 );
and AND3_13921 ( P1_U3705 , P1_U5308 , P1_U5307 , P1_U5309 );
and AND3_13922 ( P1_U3706 , P1_U5313 , P1_U5312 , P1_U5314 );
and AND3_13923 ( P1_U3707 , P1_U5318 , P1_U5317 , P1_U5319 );
and AND3_13924 ( P1_U3708 , P1_U5323 , P1_U5322 , P1_U5324 );
and AND3_13925 ( P1_U3709 , P1_U5328 , P1_U5327 , P1_U5329 );
and AND3_13926 ( P1_U3710 , P1_U5333 , P1_U5332 , P1_U5334 );
and AND3_13927 ( P1_U3711 , P1_U5338 , P1_U5337 , P1_U5339 );
and AND3_13928 ( P1_U3712 , P1_U5343 , P1_U5342 , P1_U5344 );
and AND3_13929 ( P1_U3713 , P1_U5357 , P1_U5358 , P1_U4224 );
and AND3_13930 ( P1_U3714 , P1_U5366 , P1_U5365 , P1_U5367 );
and AND3_13931 ( P1_U3715 , P1_U5371 , P1_U5370 , P1_U5372 );
and AND3_13932 ( P1_U3716 , P1_U5376 , P1_U5375 , P1_U5377 );
and AND3_13933 ( P1_U3717 , P1_U5381 , P1_U5380 , P1_U5382 );
and AND3_13934 ( P1_U3718 , P1_U5386 , P1_U5385 , P1_U5387 );
and AND3_13935 ( P1_U3719 , P1_U5391 , P1_U5390 , P1_U5392 );
and AND3_13936 ( P1_U3720 , P1_U5396 , P1_U5395 , P1_U5397 );
and AND3_13937 ( P1_U3721 , P1_U5401 , P1_U5400 , P1_U5402 );
and AND3_13938 ( P1_U3722 , P1_U5414 , P1_U5415 , P1_U4224 );
and AND3_13939 ( P1_U3723 , P1_U5423 , P1_U5422 , P1_U5424 );
and AND3_13940 ( P1_U3724 , P1_U5428 , P1_U5427 , P1_U5429 );
and AND3_13941 ( P1_U3725 , P1_U5433 , P1_U5432 , P1_U5434 );
and AND3_13942 ( P1_U3726 , P1_U5438 , P1_U5437 , P1_U5439 );
and AND3_13943 ( P1_U3727 , P1_U5442 , P1_U5441 , P1_U5443 );
and AND3_13944 ( P1_U3728 , P1_U5447 , P1_U5446 , P1_U5448 );
and AND3_13945 ( P1_U3729 , P1_U5452 , P1_U5451 , P1_U5453 );
and AND3_13946 ( P1_U3730 , P1_U5457 , P1_U5456 , P1_U5458 );
and AND2_13947 ( P1_U3731 , P1_FLUSH_REG , P1_STATE2_REG_0_ );
and AND2_13948 ( P1_U3732 , P1_U4494 , P1_U4399 );
and AND2_13949 ( P1_U3733 , P1_U4497 , P1_U3257 );
and AND2_13950 ( P1_U3734 , P1_U4210 , P1_U3257 );
and AND2_13951 ( P1_U3735 , P1_U7496 , P1_U4217 );
and AND2_13952 ( P1_U3736 , P1_U5471 , P1_U5472 );
and AND2_13953 ( P1_U3737 , P1_U3736 , P1_U5470 );
and AND2_13954 ( P1_U3738 , P1_U3737 , P1_U2518 );
and AND2_13955 ( P1_U3739 , P1_U5475 , P1_U4242 );
and AND2_13956 ( P1_U3740 , P1_U5486 , P1_U5485 );
and AND2_13957 ( P1_U3741 , P1_U4449 , P1_U4400 );
and AND2_13958 ( P1_U3742 , P1_U5496 , P1_U3393 );
and AND2_13959 ( P1_U3743 , P1_U5498 , P1_U5497 );
and AND4_13960 ( P1_U3744 , P1_U5500 , P1_U7627 , P1_U3742 , P1_U3743 );
and AND2_13961 ( P1_U3745 , P1_U4263 , P1_U3397 );
and AND5_13962 ( P1_U3746 , P1_U3411 , P1_U3288 , P1_U3745 , P1_U2520 , P1_U3279 );
and AND2_13963 ( P1_U3747 , P1_U3748 , P1_U5502 );
and AND2_13964 ( P1_U3748 , P1_U5505 , P1_U5504 );
and AND3_13965 ( P1_U3749 , P1_U7717 , P1_U7716 , P1_U5513 );
and AND2_13966 ( P1_U3750 , P1_U5524 , P1_U5522 );
and AND2_13967 ( P1_U3751 , P1_U5543 , P1_U5544 );
and AND2_13968 ( P1_U3752 , P1_U5547 , P1_U5548 );
and AND2_13969 ( P1_U3753 , P1_U5552 , P1_U5553 );
and AND2_13970 ( P1_U3754 , P1_U5558 , P1_U3257 );
and AND2_13971 ( P1_U3755 , P1_U3284 , P1_U3407 );
and AND2_13972 ( P1_U3756 , P1_U5563 , P1_U5561 );
and AND3_13973 ( P1_U3757 , P1_U3398 , P1_U3399 , P1_U5567 );
and AND3_13974 ( P1_U3758 , P1_U2520 , P1_U5568 , P1_U3757 );
and AND2_13975 ( P1_U3759 , P1_U4186 , P1_U3284 );
and AND3_13976 ( P1_U3760 , P1_U3288 , P1_U4217 , P1_U3448 );
and AND2_13977 ( P1_U3761 , P1_U5566 , P1_U7507 );
and AND2_13978 ( P1_U3762 , P1_U7508 , P1_STATE2_REG_2_ );
and AND2_13979 ( P1_U3763 , P1_U5571 , P1_U5570 );
and AND2_13980 ( P1_U3764 , P1_U5573 , P1_U5572 );
and AND2_13981 ( P1_U3765 , P1_U5575 , P1_U5576 );
and AND2_13982 ( P1_U3766 , P1_U3765 , P1_U5574 );
and AND2_13983 ( P1_U3767 , P1_U5578 , P1_U5577 );
and AND2_13984 ( P1_U3768 , P1_U5580 , P1_U5579 );
and AND2_13985 ( P1_U3769 , P1_U5582 , P1_U5583 );
and AND2_13986 ( P1_U3770 , P1_U3769 , P1_U5581 );
and AND2_13987 ( P1_U3771 , P1_U5585 , P1_U5584 );
and AND2_13988 ( P1_U3772 , P1_U5587 , P1_U5586 );
and AND2_13989 ( P1_U3773 , P1_U5589 , P1_U5590 );
and AND2_13990 ( P1_U3774 , P1_U3773 , P1_U5588 );
and AND3_13991 ( P1_U3775 , P1_U5592 , P1_U5591 , P1_U5594 );
and AND3_13992 ( P1_U3776 , P1_U3777 , P1_U5595 , P1_U5593 );
and AND2_13993 ( P1_U3777 , P1_U5596 , P1_U5597 );
and AND3_13994 ( P1_U3778 , P1_U5599 , P1_U5598 , P1_U5601 );
and AND2_13995 ( P1_U3779 , P1_U5603 , P1_U5604 );
and AND2_13996 ( P1_U3780 , P1_U3779 , P1_U5602 );
and AND3_13997 ( P1_U3781 , P1_U5606 , P1_U5605 , P1_U5608 );
and AND2_13998 ( P1_U3782 , P1_U5610 , P1_U5611 );
and AND2_13999 ( P1_U3783 , P1_U3782 , P1_U5609 );
and AND3_14000 ( P1_U3784 , P1_U5613 , P1_U5612 , P1_U5615 );
and AND2_14001 ( P1_U3785 , P1_U5617 , P1_U5618 );
and AND2_14002 ( P1_U3786 , P1_U3785 , P1_U5616 );
and AND3_14003 ( P1_U3787 , P1_U5620 , P1_U5619 , P1_U5622 );
and AND2_14004 ( P1_U3788 , P1_U5624 , P1_U5625 );
and AND2_14005 ( P1_U3789 , P1_U3788 , P1_U5623 );
and AND3_14006 ( P1_U3790 , P1_U5627 , P1_U5626 , P1_U5629 );
and AND2_14007 ( P1_U3791 , P1_U5631 , P1_U5632 );
and AND2_14008 ( P1_U3792 , P1_U3791 , P1_U5630 );
and AND3_14009 ( P1_U3793 , P1_U5634 , P1_U5633 , P1_U5636 );
and AND2_14010 ( P1_U3794 , P1_U5638 , P1_U5639 );
and AND2_14011 ( P1_U3795 , P1_U3794 , P1_U5637 );
and AND3_14012 ( P1_U3796 , P1_U5641 , P1_U5640 , P1_U5643 );
and AND2_14013 ( P1_U3797 , P1_U5645 , P1_U5646 );
and AND2_14014 ( P1_U3798 , P1_U3797 , P1_U5644 );
and AND3_14015 ( P1_U3799 , P1_U5648 , P1_U5647 , P1_U5650 );
and AND2_14016 ( P1_U3800 , P1_U5652 , P1_U5653 );
and AND2_14017 ( P1_U3801 , P1_U3800 , P1_U5651 );
and AND3_14018 ( P1_U3802 , P1_U5655 , P1_U5654 , P1_U5657 );
and AND2_14019 ( P1_U3803 , P1_U5659 , P1_U5660 );
and AND2_14020 ( P1_U3804 , P1_U3803 , P1_U5658 );
and AND2_14021 ( P1_U3805 , P1_U5662 , P1_U5664 );
and AND2_14022 ( P1_U3806 , P1_U5666 , P1_U5667 );
and AND2_14023 ( P1_U3807 , P1_U3806 , P1_U5665 );
and AND2_14024 ( P1_U3808 , P1_U5669 , P1_U5671 );
and AND2_14025 ( P1_U3809 , P1_U5673 , P1_U5674 );
and AND2_14026 ( P1_U3810 , P1_U3809 , P1_U5672 );
and AND2_14027 ( P1_U3811 , P1_U5676 , P1_U5678 );
and AND2_14028 ( P1_U3812 , P1_U5680 , P1_U5681 );
and AND2_14029 ( P1_U3813 , P1_U3812 , P1_U5679 );
and AND2_14030 ( P1_U3814 , P1_U5683 , P1_U5685 );
and AND2_14031 ( P1_U3815 , P1_U5687 , P1_U5688 );
and AND2_14032 ( P1_U3816 , P1_U3815 , P1_U5686 );
and AND2_14033 ( P1_U3817 , P1_U5690 , P1_U5692 );
and AND2_14034 ( P1_U3818 , P1_U5694 , P1_U5695 );
and AND2_14035 ( P1_U3819 , P1_U3818 , P1_U5693 );
and AND2_14036 ( P1_U3820 , P1_U5697 , P1_U5699 );
and AND2_14037 ( P1_U3821 , P1_U5701 , P1_U5702 );
and AND2_14038 ( P1_U3822 , P1_U3821 , P1_U5700 );
and AND2_14039 ( P1_U3823 , P1_U5704 , P1_U5706 );
and AND2_14040 ( P1_U3824 , P1_U5708 , P1_U5709 );
and AND2_14041 ( P1_U3825 , P1_U3824 , P1_U5707 );
and AND2_14042 ( P1_U3826 , P1_U5711 , P1_U5713 );
and AND2_14043 ( P1_U3827 , P1_U5715 , P1_U5716 );
and AND2_14044 ( P1_U3828 , P1_U3827 , P1_U5714 );
and AND2_14045 ( P1_U3829 , P1_U5718 , P1_U5720 );
and AND2_14046 ( P1_U3830 , P1_U5722 , P1_U5723 );
and AND2_14047 ( P1_U3831 , P1_U3830 , P1_U5721 );
and AND2_14048 ( P1_U3832 , P1_U5725 , P1_U5727 );
and AND2_14049 ( P1_U3833 , P1_U5729 , P1_U5730 );
and AND2_14050 ( P1_U3834 , P1_U3833 , P1_U5728 );
and AND2_14051 ( P1_U3835 , P1_U5732 , P1_U5734 );
and AND2_14052 ( P1_U3836 , P1_U5736 , P1_U5737 );
and AND2_14053 ( P1_U3837 , P1_U3836 , P1_U5735 );
and AND2_14054 ( P1_U3838 , P1_U5739 , P1_U5741 );
and AND2_14055 ( P1_U3839 , P1_U5743 , P1_U5744 );
and AND2_14056 ( P1_U3840 , P1_U3839 , P1_U5742 );
and AND2_14057 ( P1_U3841 , P1_U5746 , P1_U5748 );
and AND2_14058 ( P1_U3842 , P1_U5750 , P1_U5751 );
and AND2_14059 ( P1_U3843 , P1_U3842 , P1_U5749 );
and AND2_14060 ( P1_U3844 , P1_U5753 , P1_U5755 );
and AND2_14061 ( P1_U3845 , P1_U5757 , P1_U5758 );
and AND2_14062 ( P1_U3846 , P1_U3845 , P1_U5756 );
and AND2_14063 ( P1_U3847 , P1_U5760 , P1_U5762 );
and AND2_14064 ( P1_U3848 , P1_U5764 , P1_U5765 );
and AND2_14065 ( P1_U3849 , P1_U3848 , P1_U5763 );
and AND2_14066 ( P1_U3850 , P1_U5767 , P1_U5769 );
and AND2_14067 ( P1_U3851 , P1_U5771 , P1_U5772 );
and AND2_14068 ( P1_U3852 , P1_U3851 , P1_U5770 );
and AND2_14069 ( P1_U3853 , P1_U5774 , P1_U5776 );
and AND2_14070 ( P1_U3854 , P1_U5778 , P1_U5779 );
and AND2_14071 ( P1_U3855 , P1_U3854 , P1_U5777 );
and AND2_14072 ( P1_U3856 , P1_U5781 , P1_U5783 );
and AND2_14073 ( P1_U3857 , P1_U5785 , P1_U5786 );
and AND2_14074 ( P1_U3858 , P1_U3857 , P1_U5784 );
and AND2_14075 ( P1_U3859 , P1_U5788 , P1_U5790 );
and AND2_14076 ( P1_U3860 , P1_U5792 , P1_U5793 );
and AND2_14077 ( P1_U3861 , P1_U3860 , P1_U5791 );
and AND3_14078 ( P1_U3862 , P1_U3283 , P1_U3262 , P1_U7494 );
and AND2_14079 ( P1_U3863 , P1_U5794 , P1_U3408 );
and AND2_14080 ( P1_U3864 , P1_STATE2_REG_1_ , P1_STATEBS16_REG );
and AND2_14081 ( P1_U3865 , P1_U2368 , P1_U3284 );
and AND2_14082 ( P1_U3866 , P1_U2449 , P1_STATE2_REG_0_ );
and AND2_14083 ( P1_U3867 , P1_U4208 , P1_U2368 );
and AND2_14084 ( P1_U3868 , P1_U6105 , P1_U6106 );
and AND2_14085 ( P1_U3869 , P1_U6108 , P1_U6109 );
and AND2_14086 ( P1_U3870 , P1_U6111 , P1_U6112 );
and AND2_14087 ( P1_U3871 , P1_U6114 , P1_U6115 );
and AND2_14088 ( P1_U3872 , P1_U6117 , P1_U6118 );
and AND2_14089 ( P1_U3873 , P1_U6120 , P1_U6121 );
and AND2_14090 ( P1_U3874 , P1_U6123 , P1_U6124 );
and AND2_14091 ( P1_U3875 , P1_U6126 , P1_U6127 );
and AND2_14092 ( P1_U3876 , P1_U6129 , P1_U6130 );
and AND2_14093 ( P1_U3877 , P1_U6132 , P1_U6133 );
and AND2_14094 ( P1_U3878 , P1_U6135 , P1_U6136 );
and AND2_14095 ( P1_U3879 , P1_U6138 , P1_U6139 );
and AND2_14096 ( P1_U3880 , P1_U6141 , P1_U6142 );
and AND2_14097 ( P1_U3881 , P1_U6144 , P1_U6145 );
and AND2_14098 ( P1_U3882 , P1_U6147 , P1_U6148 );
and AND2_14099 ( P1_U3883 , P1_U6151 , P1_U6150 );
and AND2_14100 ( P1_U3884 , P1_U2605 , P1_U3391 );
and AND3_14101 ( P1_U3885 , P1_STATE2_REG_0_ , P1_U3271 , P1_U7494 );
and AND2_14102 ( P1_U3886 , P1_U4399 , P1_U4171 );
and AND3_14103 ( P1_U3887 , P1_U4241 , P1_U4244 , P1_U6362 );
nor nor_14104 ( P1_U3888 , U210 , P1_STATEBS16_REG );
and AND2_14105 ( P1_U3889 , P1_U4494 , P1_U4186 );
and AND5_14106 ( P1_U3890 , P1_U6373 , P1_U6372 , P1_U6375 , P1_U6374 , P1_U6371 );
and AND5_14107 ( P1_U3891 , P1_U6381 , P1_U6380 , P1_U6383 , P1_U6382 , P1_U6379 );
and AND5_14108 ( P1_U3892 , P1_U6389 , P1_U6388 , P1_U6391 , P1_U6390 , P1_U6387 );
and AND5_14109 ( P1_U3893 , P1_U6397 , P1_U6396 , P1_U6399 , P1_U6398 , P1_U6395 );
and AND2_14110 ( P1_U3894 , P1_U6400 , P1_U4227 );
and AND4_14111 ( P1_U3895 , P1_U6405 , P1_U6404 , P1_U6407 , P1_U6406 );
and AND2_14112 ( P1_U3896 , P1_U6408 , P1_U4227 );
and AND5_14113 ( P1_U3897 , P1_U6413 , P1_U6412 , P1_U6415 , P1_U6414 , P1_U6411 );
and AND2_14114 ( P1_U3898 , P1_U6416 , P1_U4227 );
and AND3_14115 ( P1_U3899 , P1_U6422 , P1_U6419 , P1_U6421 );
and AND2_14116 ( P1_U3900 , P1_U6423 , P1_U4227 );
and AND3_14117 ( P1_U3901 , P1_U6429 , P1_U6426 , P1_U6428 );
and AND2_14118 ( P1_U3902 , P1_U6430 , P1_U4227 );
and AND3_14119 ( P1_U3903 , P1_U6436 , P1_U6433 , P1_U6435 );
and AND2_14120 ( P1_U3904 , P1_U6437 , P1_U4227 );
and AND3_14121 ( P1_U3905 , P1_U6443 , P1_U6440 , P1_U6442 );
and AND2_14122 ( P1_U3906 , P1_U6444 , P1_U4227 );
and AND3_14123 ( P1_U3907 , P1_U6450 , P1_U6447 , P1_U6449 );
and AND2_14124 ( P1_U3908 , P1_U6451 , P1_U4227 );
and AND3_14125 ( P1_U3909 , P1_U6457 , P1_U6454 , P1_U6456 );
and AND2_14126 ( P1_U3910 , P1_U6458 , P1_U4227 );
and AND3_14127 ( P1_U3911 , P1_U6464 , P1_U6461 , P1_U6463 );
and AND2_14128 ( P1_U3912 , P1_U6465 , P1_U4227 );
and AND3_14129 ( P1_U3913 , P1_U6471 , P1_U6468 , P1_U6470 );
and AND2_14130 ( P1_U3914 , P1_U6472 , P1_U4227 );
and AND3_14131 ( P1_U3915 , P1_U6478 , P1_U6475 , P1_U6477 );
and AND2_14132 ( P1_U3916 , P1_U6479 , P1_U4227 );
and AND3_14133 ( P1_U3917 , P1_U6485 , P1_U6482 , P1_U6484 );
and AND2_14134 ( P1_U3918 , P1_U6486 , P1_U4227 );
and AND3_14135 ( P1_U3919 , P1_U6492 , P1_U6489 , P1_U6491 );
and AND2_14136 ( P1_U3920 , P1_U4227 , P1_U6494 );
and AND3_14137 ( P1_U3921 , P1_U6499 , P1_U6496 , P1_U6498 );
and AND2_14138 ( P1_U3922 , P1_U4227 , P1_U6501 );
and AND3_14139 ( P1_U3923 , P1_U6506 , P1_U6503 , P1_U6505 );
and AND2_14140 ( P1_U3924 , P1_U4227 , P1_U6508 );
and AND3_14141 ( P1_U3925 , P1_U6513 , P1_U6510 , P1_U6512 );
and AND2_14142 ( P1_U3926 , P1_U6517 , P1_U6515 );
and AND2_14143 ( P1_U3927 , P1_U6519 , P1_U6520 );
and AND2_14144 ( P1_U3928 , P1_U6524 , P1_U6522 );
and AND2_14145 ( P1_U3929 , P1_U6526 , P1_U6527 );
and AND2_14146 ( P1_U3930 , P1_U6531 , P1_U6529 );
and AND2_14147 ( P1_U3931 , P1_U6533 , P1_U6534 );
and AND2_14148 ( P1_U3932 , P1_U6538 , P1_U6536 );
and AND2_14149 ( P1_U3933 , P1_U6540 , P1_U6541 );
and AND2_14150 ( P1_U3934 , P1_U6545 , P1_U6543 );
and AND2_14151 ( P1_U3935 , P1_U6547 , P1_U6548 );
and AND2_14152 ( P1_U3936 , P1_U6552 , P1_U6550 );
and AND2_14153 ( P1_U3937 , P1_U6554 , P1_U6555 );
and AND2_14154 ( P1_U3938 , P1_U6559 , P1_U6557 );
and AND2_14155 ( P1_U3939 , P1_U6561 , P1_U6562 );
and AND2_14156 ( P1_U3940 , P1_U6566 , P1_U6564 );
and AND2_14157 ( P1_U3941 , P1_U6568 , P1_U6569 );
and AND2_14158 ( P1_U3942 , P1_U6573 , P1_U6571 );
and AND2_14159 ( P1_U3943 , P1_U6575 , P1_U6576 );
and AND2_14160 ( P1_U3944 , P1_U6580 , P1_U6578 );
and AND2_14161 ( P1_U3945 , P1_U6582 , P1_U6583 );
and AND2_14162 ( P1_U3946 , P1_U6587 , P1_U6585 );
and AND2_14163 ( P1_U3947 , P1_U6589 , P1_U6590 );
and AND2_14164 ( P1_U3948 , P1_U6594 , P1_U6592 );
and AND2_14165 ( P1_U3949 , P1_U6596 , P1_U6597 );
nor nor_14166 ( P1_U3950 , P1_DATAWIDTH_REG_2_ , P1_DATAWIDTH_REG_3_ , P1_DATAWIDTH_REG_4_ , P1_DATAWIDTH_REG_5_ );
nor nor_14167 ( P1_U3951 , P1_DATAWIDTH_REG_6_ , P1_DATAWIDTH_REG_7_ , P1_DATAWIDTH_REG_8_ , P1_DATAWIDTH_REG_9_ );
and AND2_14168 ( P1_U3952 , P1_U3951 , P1_U3950 );
nor nor_14169 ( P1_U3953 , P1_DATAWIDTH_REG_10_ , P1_DATAWIDTH_REG_11_ , P1_DATAWIDTH_REG_12_ , P1_DATAWIDTH_REG_13_ );
nor nor_14170 ( P1_U3954 , P1_DATAWIDTH_REG_14_ , P1_DATAWIDTH_REG_15_ , P1_DATAWIDTH_REG_16_ , P1_DATAWIDTH_REG_17_ );
and AND2_14171 ( P1_U3955 , P1_U3954 , P1_U3953 );
nor nor_14172 ( P1_U3956 , P1_DATAWIDTH_REG_18_ , P1_DATAWIDTH_REG_19_ , P1_DATAWIDTH_REG_20_ , P1_DATAWIDTH_REG_21_ );
nor nor_14173 ( P1_U3957 , P1_DATAWIDTH_REG_22_ , P1_DATAWIDTH_REG_23_ , P1_DATAWIDTH_REG_24_ , P1_DATAWIDTH_REG_25_ );
and AND2_14174 ( P1_U3958 , P1_U3957 , P1_U3956 );
nor nor_14175 ( P1_U3959 , P1_DATAWIDTH_REG_26_ , P1_DATAWIDTH_REG_27_ );
nor nor_14176 ( P1_U3960 , P1_DATAWIDTH_REG_28_ , P1_DATAWIDTH_REG_29_ );
nor nor_14177 ( P1_U3961 , P1_DATAWIDTH_REG_30_ , P1_DATAWIDTH_REG_31_ );
and AND4_14178 ( P1_U3962 , P1_U3961 , P1_U6598 , P1_U3960 , P1_U3959 );
nor nor_14179 ( P1_U3963 , P1_REIP_REG_0_ , P1_DATAWIDTH_REG_0_ , P1_DATAWIDTH_REG_1_ );
and AND2_14180 ( P1_U3964 , P1_STATE2_REG_2_ , P1_U3257 );
and AND2_14181 ( P1_U3965 , P1_U6608 , P1_U3298 );
nor nor_14182 ( P1_U3966 , U210 , P1_STATE2_REG_0_ );
and AND3_14183 ( P1_U3967 , P1_U3307 , P1_U3408 , P1_U6602 );
and AND2_14184 ( P1_U3968 , P1_STATE2_REG_2_ , P1_U3287 );
and AND2_14185 ( P1_U3969 , P1_U4235 , P1_U4206 );
and AND4_14186 ( P1_U3970 , P1_U6621 , P1_U6620 , P1_U6619 , P1_U6618 );
and AND4_14187 ( P1_U3971 , P1_U6625 , P1_U6624 , P1_U6623 , P1_U6622 );
and AND4_14188 ( P1_U3972 , P1_U6629 , P1_U6628 , P1_U6627 , P1_U6626 );
and AND4_14189 ( P1_U3973 , P1_U6633 , P1_U6632 , P1_U6631 , P1_U6630 );
and AND4_14190 ( P1_U3974 , P1_U6637 , P1_U6636 , P1_U6635 , P1_U6634 );
and AND4_14191 ( P1_U3975 , P1_U6641 , P1_U6640 , P1_U6639 , P1_U6638 );
and AND4_14192 ( P1_U3976 , P1_U6645 , P1_U6644 , P1_U6643 , P1_U6642 );
and AND4_14193 ( P1_U3977 , P1_U6649 , P1_U6648 , P1_U6647 , P1_U6646 );
and AND4_14194 ( P1_U3978 , P1_U6653 , P1_U6652 , P1_U6651 , P1_U6650 );
and AND4_14195 ( P1_U3979 , P1_U6657 , P1_U6656 , P1_U6655 , P1_U6654 );
and AND4_14196 ( P1_U3980 , P1_U6661 , P1_U6660 , P1_U6659 , P1_U6658 );
and AND4_14197 ( P1_U3981 , P1_U6665 , P1_U6664 , P1_U6663 , P1_U6662 );
and AND4_14198 ( P1_U3982 , P1_U6669 , P1_U6668 , P1_U6667 , P1_U6666 );
and AND4_14199 ( P1_U3983 , P1_U6673 , P1_U6672 , P1_U6671 , P1_U6670 );
and AND4_14200 ( P1_U3984 , P1_U6677 , P1_U6676 , P1_U6675 , P1_U6674 );
and AND4_14201 ( P1_U3985 , P1_U7613 , P1_U6680 , P1_U6679 , P1_U6678 );
and AND4_14202 ( P1_U3986 , P1_U6684 , P1_U6683 , P1_U6682 , P1_U6681 );
and AND4_14203 ( P1_U3987 , P1_U6688 , P1_U6687 , P1_U6686 , P1_U6685 );
and AND4_14204 ( P1_U3988 , P1_U6692 , P1_U6691 , P1_U6690 , P1_U6689 );
and AND4_14205 ( P1_U3989 , P1_U6696 , P1_U6695 , P1_U6694 , P1_U6693 );
and AND4_14206 ( P1_U3990 , P1_U6700 , P1_U6699 , P1_U6698 , P1_U6697 );
and AND4_14207 ( P1_U3991 , P1_U6704 , P1_U6703 , P1_U6702 , P1_U6701 );
and AND4_14208 ( P1_U3992 , P1_U6708 , P1_U6707 , P1_U6706 , P1_U6705 );
and AND4_14209 ( P1_U3993 , P1_U6712 , P1_U6711 , P1_U6710 , P1_U6709 );
and AND4_14210 ( P1_U3994 , P1_U6716 , P1_U6715 , P1_U6714 , P1_U6713 );
and AND4_14211 ( P1_U3995 , P1_U6720 , P1_U6719 , P1_U6718 , P1_U6717 );
and AND4_14212 ( P1_U3996 , P1_U6724 , P1_U6723 , P1_U6722 , P1_U6721 );
and AND4_14213 ( P1_U3997 , P1_U6728 , P1_U6727 , P1_U6726 , P1_U6725 );
and AND4_14214 ( P1_U3998 , P1_U6732 , P1_U6731 , P1_U6730 , P1_U6729 );
and AND4_14215 ( P1_U3999 , P1_U6736 , P1_U6735 , P1_U6734 , P1_U6733 );
and AND4_14216 ( P1_U4000 , P1_U6740 , P1_U6739 , P1_U6738 , P1_U6737 );
and AND4_14217 ( P1_U4001 , P1_U6744 , P1_U6743 , P1_U6742 , P1_U6741 );
and AND2_14218 ( P1_U4002 , P1_U6749 , P1_U6748 );
and AND2_14219 ( P1_U4003 , P1_U6752 , P1_U6751 );
and AND2_14220 ( P1_U4004 , P1_U6755 , P1_U6754 );
and AND2_14221 ( P1_U4005 , P1_U6758 , P1_U6757 );
and AND2_14222 ( P1_U4006 , P1_U6760 , P1_U4007 );
and AND2_14223 ( P1_U4007 , P1_U6762 , P1_U6761 );
and AND2_14224 ( P1_U4008 , P1_U6764 , P1_U6765 );
and AND3_14225 ( P1_U4009 , P1_U6772 , P1_U6773 , P1_U6774 );
and AND2_14226 ( P1_U4010 , P1_U6776 , P1_U6777 );
and AND3_14227 ( P1_U4011 , P1_U6781 , P1_U6782 , P1_U6783 );
and AND3_14228 ( P1_U4012 , P1_U6785 , P1_U6786 , P1_U6787 );
and AND3_14229 ( P1_U4013 , P1_U6789 , P1_U6790 , P1_U6791 );
and AND3_14230 ( P1_U4014 , P1_U6793 , P1_U6794 , P1_U6795 );
and AND3_14231 ( P1_U4015 , P1_U6797 , P1_U6798 , P1_U6799 );
and AND3_14232 ( P1_U4016 , P1_U6801 , P1_U6802 , P1_U6803 );
and AND3_14233 ( P1_U4017 , P1_U6805 , P1_U6806 , P1_U6807 );
and AND3_14234 ( P1_U4018 , P1_U6809 , P1_U6810 , P1_U6811 );
and AND3_14235 ( P1_U4019 , P1_U6813 , P1_U6814 , P1_U6815 );
and AND3_14236 ( P1_U4020 , P1_U6817 , P1_U6818 , P1_U6819 );
and AND2_14237 ( P1_U4021 , P1_U6821 , P1_U6822 );
and AND3_14238 ( P1_U4022 , P1_U6826 , P1_U6827 , P1_U6828 );
and AND3_14239 ( P1_U4023 , P1_U6830 , P1_U6831 , P1_U6832 );
and AND3_14240 ( P1_U4024 , P1_U6834 , P1_U6835 , P1_U6836 );
and AND3_14241 ( P1_U4025 , P1_U6838 , P1_U6839 , P1_U6840 );
and AND2_14242 ( P1_U4026 , P1_U6858 , P1_U6857 );
and AND2_14243 ( P1_U4027 , P1_U6860 , P1_U6861 );
and AND3_14244 ( P1_U4028 , P1_U7494 , P1_U6888 , P1_U3283 );
and AND4_14245 ( P1_U4029 , P1_U6895 , P1_U6894 , P1_U6893 , P1_U6892 );
and AND4_14246 ( P1_U4030 , P1_U6899 , P1_U6898 , P1_U6897 , P1_U6896 );
and AND4_14247 ( P1_U4031 , P1_U6903 , P1_U6902 , P1_U6901 , P1_U6900 );
and AND4_14248 ( P1_U4032 , P1_U6907 , P1_U6906 , P1_U6905 , P1_U6904 );
and AND4_14249 ( P1_U4033 , P1_U6913 , P1_U6912 , P1_U6911 , P1_U6910 );
and AND4_14250 ( P1_U4034 , P1_U6917 , P1_U6916 , P1_U6915 , P1_U6914 );
and AND4_14251 ( P1_U4035 , P1_U6921 , P1_U6920 , P1_U6919 , P1_U6918 );
and AND4_14252 ( P1_U4036 , P1_U6925 , P1_U6924 , P1_U6923 , P1_U6922 );
and AND4_14253 ( P1_U4037 , P1_U6944 , P1_U6943 , P1_U6942 , P1_U6941 );
and AND4_14254 ( P1_U4038 , P1_U6948 , P1_U6947 , P1_U6946 , P1_U6945 );
and AND4_14255 ( P1_U4039 , P1_U6952 , P1_U6951 , P1_U6950 , P1_U6949 );
and AND4_14256 ( P1_U4040 , P1_U6956 , P1_U6955 , P1_U6954 , P1_U6953 );
and AND4_14257 ( P1_U4041 , P1_U6961 , P1_U6960 , P1_U6959 , P1_U6958 );
and AND4_14258 ( P1_U4042 , P1_U6965 , P1_U6964 , P1_U6963 , P1_U6962 );
and AND4_14259 ( P1_U4043 , P1_U6969 , P1_U6968 , P1_U6967 , P1_U6966 );
and AND4_14260 ( P1_U4044 , P1_U6973 , P1_U6972 , P1_U6971 , P1_U6970 );
and AND4_14261 ( P1_U4045 , P1_U6978 , P1_U6977 , P1_U6976 , P1_U6975 );
and AND4_14262 ( P1_U4046 , P1_U6982 , P1_U6981 , P1_U6980 , P1_U6979 );
and AND4_14263 ( P1_U4047 , P1_U6986 , P1_U6985 , P1_U6984 , P1_U6983 );
and AND4_14264 ( P1_U4048 , P1_U6990 , P1_U6989 , P1_U6988 , P1_U6987 );
and AND4_14265 ( P1_U4049 , P1_U6995 , P1_U6994 , P1_U6993 , P1_U6992 );
and AND4_14266 ( P1_U4050 , P1_U6999 , P1_U6998 , P1_U6997 , P1_U6996 );
and AND4_14267 ( P1_U4051 , P1_U7003 , P1_U7002 , P1_U7001 , P1_U7000 );
and AND4_14268 ( P1_U4052 , P1_U7614 , P1_U7006 , P1_U7005 , P1_U7004 );
and AND4_14269 ( P1_U4053 , P1_U7010 , P1_U7009 , P1_U7008 , P1_U7007 );
and AND4_14270 ( P1_U4054 , P1_U7014 , P1_U7013 , P1_U7012 , P1_U7011 );
and AND4_14271 ( P1_U4055 , P1_U7018 , P1_U7017 , P1_U7016 , P1_U7015 );
and AND4_14272 ( P1_U4056 , P1_U7022 , P1_U7021 , P1_U7020 , P1_U7019 );
and AND4_14273 ( P1_U4057 , P1_U7027 , P1_U7026 , P1_U7025 , P1_U7024 );
and AND4_14274 ( P1_U4058 , P1_U7031 , P1_U7030 , P1_U7029 , P1_U7028 );
and AND4_14275 ( P1_U4059 , P1_U7035 , P1_U7034 , P1_U7033 , P1_U7032 );
and AND4_14276 ( P1_U4060 , P1_U7039 , P1_U7038 , P1_U7037 , P1_U7036 );
and AND2_14277 ( P1_U4061 , P1_U7059 , P1_U3443 );
and AND2_14278 ( P1_U4062 , P1_STATE2_REG_0_ , P1_U7062 );
and AND4_14279 ( P1_U4063 , P1_U7069 , P1_U7068 , P1_U7067 , P1_U7066 );
and AND4_14280 ( P1_U4064 , P1_U7073 , P1_U7072 , P1_U7071 , P1_U7070 );
and AND4_14281 ( P1_U4065 , P1_U7077 , P1_U7076 , P1_U7075 , P1_U7074 );
and AND4_14282 ( P1_U4066 , P1_U7081 , P1_U7080 , P1_U7079 , P1_U7078 );
and AND2_14283 ( P1_U4067 , P1_U4256 , P1_STATE2_REG_0_ );
and AND4_14284 ( P1_U4068 , P1_U4405 , P1_U4404 , P1_U4403 , P1_U4401 );
and AND3_14285 ( P1_U4069 , P1_U4407 , P1_U4406 , P1_U4408 );
and AND4_14286 ( P1_U4070 , P1_U4412 , P1_U4411 , P1_U4410 , P1_U4409 );
and AND2_14287 ( P1_U4071 , P1_U4414 , P1_U4413 );
and AND2_14288 ( P1_U4072 , P1_U4400 , P1_U3391 );
and AND2_14289 ( P1_U4073 , P1_STATE2_REG_0_ , P1_U3284 );
and AND2_14290 ( P1_U4074 , P1_U7090 , P1_U7089 );
and AND3_14291 ( P1_U4075 , P1_U7472 , P1_U3434 , P1_U7473 );
and AND3_14292 ( P1_U4076 , P1_U7475 , P1_U7476 , P1_U7474 );
and AND3_14293 ( P1_U4077 , P1_U2606 , P1_U7477 , P1_U4076 );
and AND2_14294 ( P1_U4078 , P1_U7097 , P1_U7095 );
and AND4_14295 ( P1_U4079 , P1_U7101 , P1_U7100 , P1_U7099 , P1_U7098 );
and AND4_14296 ( P1_U4080 , P1_U7105 , P1_U7104 , P1_U7103 , P1_U7102 );
and AND4_14297 ( P1_U4081 , P1_U7109 , P1_U7108 , P1_U7107 , P1_U7106 );
and AND4_14298 ( P1_U4082 , P1_U7113 , P1_U7112 , P1_U7111 , P1_U7110 );
and AND4_14299 ( P1_U4083 , P1_U7118 , P1_U7117 , P1_U7116 , P1_U7115 );
and AND4_14300 ( P1_U4084 , P1_U7122 , P1_U7121 , P1_U7120 , P1_U7119 );
and AND4_14301 ( P1_U4085 , P1_U7126 , P1_U7125 , P1_U7124 , P1_U7123 );
and AND4_14302 ( P1_U4086 , P1_U7130 , P1_U7129 , P1_U7128 , P1_U7127 );
and AND4_14303 ( P1_U4087 , P1_U7135 , P1_U7134 , P1_U7133 , P1_U7132 );
and AND4_14304 ( P1_U4088 , P1_U7139 , P1_U7138 , P1_U7137 , P1_U7136 );
and AND4_14305 ( P1_U4089 , P1_U7143 , P1_U7142 , P1_U7141 , P1_U7140 );
and AND2_14306 ( P1_U4090 , P1_U7145 , P1_U7144 );
and AND3_14307 ( P1_U4091 , P1_U7617 , P1_U7146 , P1_U4090 );
and AND4_14308 ( P1_U4092 , P1_U7150 , P1_U7149 , P1_U7148 , P1_U7147 );
and AND4_14309 ( P1_U4093 , P1_U7154 , P1_U7153 , P1_U7152 , P1_U7151 );
and AND4_14310 ( P1_U4094 , P1_U7158 , P1_U7157 , P1_U7156 , P1_U7155 );
and AND4_14311 ( P1_U4095 , P1_U7162 , P1_U7161 , P1_U7160 , P1_U7159 );
and AND4_14312 ( P1_U4096 , P1_U7167 , P1_U7166 , P1_U7165 , P1_U7164 );
and AND4_14313 ( P1_U4097 , P1_U7171 , P1_U7170 , P1_U7169 , P1_U7168 );
and AND4_14314 ( P1_U4098 , P1_U7175 , P1_U7174 , P1_U7173 , P1_U7172 );
and AND4_14315 ( P1_U4099 , P1_U7179 , P1_U7178 , P1_U7177 , P1_U7176 );
and AND4_14316 ( P1_U4100 , P1_U7184 , P1_U7183 , P1_U7182 , P1_U7181 );
and AND4_14317 ( P1_U4101 , P1_U7188 , P1_U7187 , P1_U7186 , P1_U7185 );
and AND4_14318 ( P1_U4102 , P1_U7192 , P1_U7191 , P1_U7190 , P1_U7189 );
and AND4_14319 ( P1_U4103 , P1_U7196 , P1_U7195 , P1_U7194 , P1_U7193 );
and AND4_14320 ( P1_U4104 , P1_U7201 , P1_U7200 , P1_U7199 , P1_U7198 );
and AND4_14321 ( P1_U4105 , P1_U7205 , P1_U7204 , P1_U7203 , P1_U7202 );
and AND4_14322 ( P1_U4106 , P1_U7209 , P1_U7208 , P1_U7207 , P1_U7206 );
and AND4_14323 ( P1_U4107 , P1_U7213 , P1_U7212 , P1_U7211 , P1_U7210 );
and AND2_14324 ( P1_U4108 , P1_U7215 , P1_U3264 );
and AND2_14325 ( P1_U4109 , P1_U7216 , P1_U7215 );
and AND2_14326 ( P1_U4110 , P1_U7217 , P1_U3265 );
and AND2_14327 ( P1_U4111 , P1_U7089 , P1_U3427 );
and AND2_14328 ( P1_U4112 , P1_U7218 , P1_U7217 );
and AND3_14329 ( P1_U4113 , P1_U4112 , P1_U7472 , P1_U7473 );
and AND4_14330 ( P1_U4114 , P1_U7090 , P1_U3434 , P1_U4111 , P1_U4113 );
and AND4_14331 ( P1_U4115 , P1_U7486 , P1_U7480 , P1_U7476 , P1_U7474 );
and AND4_14332 ( P1_U4116 , P1_U7505 , P1_U7489 , P1_U7488 , P1_U7487 );
and AND2_14333 ( P1_U4117 , P1_U7090 , P1_U7089 );
and AND3_14334 ( P1_U4118 , P1_U7472 , P1_U3434 , P1_U7473 );
and AND3_14335 ( P1_U4119 , P1_U7475 , P1_U7476 , P1_U7474 );
and AND4_14336 ( P1_U4120 , P1_U2608 , P1_U7477 , P1_U2606 , P1_U4119 );
and AND4_14337 ( P1_U4121 , P1_U7223 , P1_U7222 , P1_U7221 , P1_U7220 );
and AND4_14338 ( P1_U4122 , P1_U7227 , P1_U7226 , P1_U7225 , P1_U7224 );
and AND4_14339 ( P1_U4123 , P1_U7231 , P1_U7230 , P1_U7229 , P1_U7228 );
and AND4_14340 ( P1_U4124 , P1_U7235 , P1_U7234 , P1_U7233 , P1_U7232 );
and AND4_14341 ( P1_U4125 , P1_U7240 , P1_U7239 , P1_U7238 , P1_U7237 );
and AND4_14342 ( P1_U4126 , P1_U7244 , P1_U7243 , P1_U7242 , P1_U7241 );
and AND4_14343 ( P1_U4127 , P1_U7248 , P1_U7247 , P1_U7246 , P1_U7245 );
and AND4_14344 ( P1_U4128 , P1_U7252 , P1_U7251 , P1_U7250 , P1_U7249 );
and AND4_14345 ( P1_U4129 , P1_U7257 , P1_U7256 , P1_U7255 , P1_U7254 );
and AND4_14346 ( P1_U4130 , P1_U7261 , P1_U7260 , P1_U7259 , P1_U7258 );
and AND4_14347 ( P1_U4131 , P1_U7265 , P1_U7264 , P1_U7263 , P1_U7262 );
and AND4_14348 ( P1_U4132 , P1_U7269 , P1_U7268 , P1_U7267 , P1_U7266 );
and AND4_14349 ( P1_U4133 , P1_U7274 , P1_U7273 , P1_U7272 , P1_U7271 );
and AND4_14350 ( P1_U4134 , P1_U7278 , P1_U7277 , P1_U7276 , P1_U7275 );
and AND4_14351 ( P1_U4135 , P1_U7282 , P1_U7281 , P1_U7280 , P1_U7279 );
and AND4_14352 ( P1_U4136 , P1_U7619 , P1_U7285 , P1_U7284 , P1_U7283 );
and AND4_14353 ( P1_U4137 , P1_U7289 , P1_U7288 , P1_U7287 , P1_U7286 );
and AND4_14354 ( P1_U4138 , P1_U7293 , P1_U7292 , P1_U7291 , P1_U7290 );
and AND4_14355 ( P1_U4139 , P1_U7297 , P1_U7296 , P1_U7295 , P1_U7294 );
and AND4_14356 ( P1_U4140 , P1_U7301 , P1_U7300 , P1_U7299 , P1_U7298 );
and AND4_14357 ( P1_U4141 , P1_U7306 , P1_U7305 , P1_U7304 , P1_U7303 );
and AND4_14358 ( P1_U4142 , P1_U7310 , P1_U7309 , P1_U7308 , P1_U7307 );
and AND4_14359 ( P1_U4143 , P1_U7314 , P1_U7313 , P1_U7312 , P1_U7311 );
and AND4_14360 ( P1_U4144 , P1_U7318 , P1_U7317 , P1_U7316 , P1_U7315 );
and AND4_14361 ( P1_U4145 , P1_U7323 , P1_U7322 , P1_U7321 , P1_U7320 );
and AND4_14362 ( P1_U4146 , P1_U7327 , P1_U7326 , P1_U7325 , P1_U7324 );
and AND4_14363 ( P1_U4147 , P1_U7331 , P1_U7330 , P1_U7329 , P1_U7328 );
and AND4_14364 ( P1_U4148 , P1_U7335 , P1_U7334 , P1_U7333 , P1_U7332 );
and AND4_14365 ( P1_U4149 , P1_U7340 , P1_U7339 , P1_U7338 , P1_U7337 );
and AND4_14366 ( P1_U4150 , P1_U7344 , P1_U7343 , P1_U7342 , P1_U7341 );
and AND4_14367 ( P1_U4151 , P1_U7348 , P1_U7347 , P1_U7346 , P1_U7345 );
and AND4_14368 ( P1_U4152 , P1_U7352 , P1_U7351 , P1_U7350 , P1_U7349 );
and AND2_14369 ( P1_U4153 , P1_U3284 , P1_U3419 );
and AND2_14370 ( P1_U4154 , P1_U3283 , P1_U3391 );
and AND3_14371 ( P1_U4155 , P1_U7357 , P1_U7358 , P1_U4263 );
and AND2_14372 ( P1_U4156 , P1_U4155 , P1_U7359 );
and AND2_14373 ( P1_U4157 , P1_STATE2_REG_0_ , P1_U2427 );
and AND2_14374 ( P1_U4158 , P1_U4157 , P1_U7360 );
and AND2_14375 ( P1_U4159 , P1_U3271 , P1_U4173 );
and AND2_14376 ( P1_U4160 , P1_STATE2_REG_0_ , P1_U4173 );
and AND2_14377 ( P1_U4161 , P1_U7369 , P1_STATE2_REG_0_ );
and AND2_14378 ( P1_U4162 , P1_U7371 , P1_U2603 );
and AND2_14379 ( P1_U4163 , P1_U7373 , P1_STATE2_REG_0_ );
and AND2_14380 ( P1_U4164 , P1_U7375 , P1_U2603 );
and AND2_14381 ( P1_U4165 , P1_U7382 , P1_U7383 );
and AND2_14382 ( P1_U4166 , P1_U3453 , P1_U7384 );
and AND3_14383 ( P1_U4167 , P1_U7389 , P1_U7388 , P1_U7387 );
and AND2_14384 ( P1_U4168 , P1_U7462 , P1_U7461 );
and AND2_14385 ( P1_U4169 , P1_U7465 , P1_U7464 );
and AND2_14386 ( P1_U4170 , P1_U7674 , P1_U7673 );
nand NAND4_14387 ( P1_U4171 , P1_U3572 , P1_U3571 , P1_U3570 , P1_U3569 );
nand NAND2_14388 ( P1_U4172 , P1_U3739 , P1_U5474 );
nand NAND5_14389 ( P1_U4173 , P1_U3576 , P1_U2607 , P1_U3575 , P1_U3574 , P1_U3573 );
not NOT1_14390 ( P1_U4174 , P1_INSTADDRPOINTER_REG_31_ );
and AND2_14391 ( P1_U4175 , P1_U7726 , P1_U7725 );
and AND2_14392 ( P1_U4176 , P1_U7745 , P1_U7744 );
nand NAND2_14393 ( P1_U4177 , P1_U2368 , P1_U3285 );
nand NAND2_14394 ( P1_U4178 , P1_U4508 , P1_U3391 );
not NOT1_14395 ( P1_U4179 , BS16 );
nand NAND2_14396 ( P1_U4180 , P1_U3967 , P1_U4228 );
nand NAND2_14397 ( P1_U4181 , P1_U4228 , P1_U3432 );
nand NAND3_14398 ( P1_U4182 , P1_U7698 , P1_U7697 , P1_U3738 );
nand NAND2_14399 ( P1_U4183 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3269 );
not NOT1_14400 ( P1_U4184 , P1_U3452 );
nand NAND2_14401 ( P1_U4185 , HOLD , P1_U3257 );
not NOT1_14402 ( P1_U4186 , P1_U3412 );
not NOT1_14403 ( P1_U4187 , P1_U3440 );
not NOT1_14404 ( P1_U4188 , P1_U3439 );
not NOT1_14405 ( P1_U4189 , P1_U3393 );
not NOT1_14406 ( P1_U4190 , P1_U3290 );
not NOT1_14407 ( P1_U4191 , P1_U3449 );
not NOT1_14408 ( P1_U4192 , P1_U3405 );
not NOT1_14409 ( P1_U4193 , P1_U3434 );
not NOT1_14410 ( P1_U4194 , P1_U3420 );
nand NAND2_14411 ( P1_U4195 , P1_U4265 , P1_U3271 );
nand NAND2_14412 ( P1_U4196 , P1_U4460 , P1_U2605 );
not NOT1_14413 ( P1_U4197 , P1_U3396 );
not NOT1_14414 ( P1_U4198 , P1_U3425 );
not NOT1_14415 ( P1_U4199 , P1_U3289 );
not NOT1_14416 ( P1_U4200 , P1_U3421 );
not NOT1_14417 ( P1_U4201 , P1_U3422 );
not NOT1_14418 ( P1_U4202 , P1_U3428 );
not NOT1_14419 ( P1_U4203 , P1_U3408 );
not NOT1_14420 ( P1_U4204 , P1_U3427 );
nand NAND3_14421 ( P1_U4205 , P1_U3885 , P1_U4189 , P1_U4197 );
not NOT1_14422 ( P1_U4206 , P1_U3418 );
not NOT1_14423 ( P1_U4207 , P1_U3443 );
not NOT1_14424 ( P1_U4208 , P1_U3282 );
not NOT1_14425 ( P1_U4209 , P1_U3307 );
not NOT1_14426 ( P1_U4210 , P1_U3390 );
not NOT1_14427 ( P1_U4211 , P1_U3446 );
not NOT1_14428 ( P1_U4212 , P1_U3447 );
not NOT1_14429 ( P1_U4213 , P1_U3448 );
not NOT1_14430 ( P1_U4214 , P1_U3400 );
not NOT1_14431 ( P1_U4215 , P1_U3288 );
not NOT1_14432 ( P1_U4216 , P1_U3292 );
nand NAND2_14433 ( P1_U4217 , P1_U3578 , P1_U2431 );
not NOT1_14434 ( P1_U4218 , P1_U3399 );
nand NAND2_14435 ( P1_U4219 , P1_U4449 , P1_U3271 );
not NOT1_14436 ( P1_U4220 , P1_U3433 );
not NOT1_14437 ( P1_U4221 , P1_U3249 );
not NOT1_14438 ( P1_U4222 , P1_U3426 );
not NOT1_14439 ( P1_U4223 , P1_U3424 );
not NOT1_14440 ( P1_U4224 , P1_U3300 );
not NOT1_14441 ( P1_U4225 , P1_LT_563_1260_U6 );
not NOT1_14442 ( P1_U4226 , P1_U3320 );
nand NAND2_14443 ( P1_U4227 , P1_U4255 , P1_U3431 );
nand NAND2_14444 ( P1_U4228 , P1_U4235 , P1_U7500 );
nand NAND2_14445 ( P1_U4229 , P1_U2362 , P1_U3272 );
nand NAND2_14446 ( P1_U4230 , P1_U2363 , P1_U4377 );
not NOT1_14447 ( P1_U4231 , P1_U3407 );
not NOT1_14448 ( P1_U4232 , P1_U3252 );
not NOT1_14449 ( P1_U4233 , P1_U3250 );
not NOT1_14450 ( P1_U4234 , P1_U3395 );
not NOT1_14451 ( P1_U4235 , P1_U3297 );
not NOT1_14452 ( P1_U4236 , P1_U3398 );
not NOT1_14453 ( P1_U4237 , P1_U4178 );
not NOT1_14454 ( P1_U4238 , P1_U3357 );
nand NAND2_14455 ( P1_U4239 , P1_U4477 , P1_U7381 );
nand NAND2_14456 ( P1_U4240 , P1_U3963 , P1_U4220 );
nand NAND2_14457 ( P1_U4241 , P1_U3584 , P1_U4261 );
nand NAND2_14458 ( P1_U4242 , P1_U3731 , P1_U2428 );
nand NAND2_14459 ( P1_U4243 , P1_U4364 , P1_U3258 );
nand NAND3_14460 ( P1_U4244 , P1_STATE2_REG_1_ , P1_U3294 , P1_U2352 );
nand NAND2_14461 ( P1_U4245 , P1_U2428 , P1_U3403 );
nand NAND3_14462 ( P1_U4246 , P1_STATE2_REG_0_ , P1_U3263 , U210 );
not NOT1_14463 ( P1_U4247 , P1_U3394 );
nand NAND4_14464 ( P1_U4248 , P1_U2451 , P1_U2353 , P1_U3862 , P1_U2448 );
not NOT1_14465 ( P1_U4249 , P1_U3287 );
not NOT1_14466 ( P1_U4250 , P1_U3397 );
not NOT1_14467 ( P1_U4251 , P1_U3415 );
not NOT1_14468 ( P1_U4252 , P1_U3299 );
not NOT1_14469 ( P1_U4253 , P1_U3409 );
not NOT1_14470 ( P1_U4254 , P1_U3419 );
not NOT1_14471 ( P1_U4255 , P1_U3432 );
not NOT1_14472 ( P1_U4256 , P1_U3291 );
not NOT1_14473 ( P1_U4257 , P1_U3389 );
not NOT1_14474 ( P1_U4258 , P1_U3254 );
not NOT1_14475 ( P1_U4259 , P1_U3281 );
not NOT1_14476 ( P1_U4260 , P1_U3406 );
not NOT1_14477 ( P1_U4261 , P1_U3298 );
not NOT1_14478 ( P1_U4262 , P1_U3286 );
nand NAND2_14479 ( P1_U4263 , P1_U4236 , P1_U4399 );
not NOT1_14480 ( P1_U4264 , P1_U3411 );
not NOT1_14481 ( P1_U4265 , P1_U3453 );
not NOT1_14482 ( P1_U4266 , P1_U3410 );
nand NAND2_14483 ( P1_U4267 , P1_REIP_REG_31_ , P1_U4233 );
nand NAND2_14484 ( P1_U4268 , P1_REIP_REG_30_ , P1_U4232 );
nand NAND2_14485 ( P1_U4269 , P1_ADDRESS_REG_29_ , P1_U3249 );
nand NAND2_14486 ( P1_U4270 , P1_REIP_REG_30_ , P1_U4233 );
nand NAND2_14487 ( P1_U4271 , P1_REIP_REG_29_ , P1_U4232 );
nand NAND2_14488 ( P1_U4272 , P1_ADDRESS_REG_28_ , P1_U3249 );
nand NAND2_14489 ( P1_U4273 , P1_REIP_REG_29_ , P1_U4233 );
nand NAND2_14490 ( P1_U4274 , P1_REIP_REG_28_ , P1_U4232 );
nand NAND2_14491 ( P1_U4275 , P1_ADDRESS_REG_27_ , P1_U3249 );
nand NAND2_14492 ( P1_U4276 , P1_REIP_REG_28_ , P1_U4233 );
nand NAND2_14493 ( P1_U4277 , P1_REIP_REG_27_ , P1_U4232 );
nand NAND2_14494 ( P1_U4278 , P1_ADDRESS_REG_26_ , P1_U3249 );
nand NAND2_14495 ( P1_U4279 , P1_REIP_REG_27_ , P1_U4233 );
nand NAND2_14496 ( P1_U4280 , P1_REIP_REG_26_ , P1_U4232 );
nand NAND2_14497 ( P1_U4281 , P1_ADDRESS_REG_25_ , P1_U3249 );
nand NAND2_14498 ( P1_U4282 , P1_REIP_REG_26_ , P1_U4233 );
nand NAND2_14499 ( P1_U4283 , P1_REIP_REG_25_ , P1_U4232 );
nand NAND2_14500 ( P1_U4284 , P1_ADDRESS_REG_24_ , P1_U3249 );
nand NAND2_14501 ( P1_U4285 , P1_REIP_REG_25_ , P1_U4233 );
nand NAND2_14502 ( P1_U4286 , P1_REIP_REG_24_ , P1_U4232 );
nand NAND2_14503 ( P1_U4287 , P1_ADDRESS_REG_23_ , P1_U3249 );
nand NAND2_14504 ( P1_U4288 , P1_REIP_REG_24_ , P1_U4233 );
nand NAND2_14505 ( P1_U4289 , P1_REIP_REG_23_ , P1_U4232 );
nand NAND2_14506 ( P1_U4290 , P1_ADDRESS_REG_22_ , P1_U3249 );
nand NAND2_14507 ( P1_U4291 , P1_REIP_REG_23_ , P1_U4233 );
nand NAND2_14508 ( P1_U4292 , P1_REIP_REG_22_ , P1_U4232 );
nand NAND2_14509 ( P1_U4293 , P1_ADDRESS_REG_21_ , P1_U3249 );
nand NAND2_14510 ( P1_U4294 , P1_REIP_REG_22_ , P1_U4233 );
nand NAND2_14511 ( P1_U4295 , P1_REIP_REG_21_ , P1_U4232 );
nand NAND2_14512 ( P1_U4296 , P1_ADDRESS_REG_20_ , P1_U3249 );
nand NAND2_14513 ( P1_U4297 , P1_REIP_REG_21_ , P1_U4233 );
nand NAND2_14514 ( P1_U4298 , P1_REIP_REG_20_ , P1_U4232 );
nand NAND2_14515 ( P1_U4299 , P1_ADDRESS_REG_19_ , P1_U3249 );
nand NAND2_14516 ( P1_U4300 , P1_REIP_REG_20_ , P1_U4233 );
nand NAND2_14517 ( P1_U4301 , P1_REIP_REG_19_ , P1_U4232 );
nand NAND2_14518 ( P1_U4302 , P1_ADDRESS_REG_18_ , P1_U3249 );
nand NAND2_14519 ( P1_U4303 , P1_REIP_REG_19_ , P1_U4233 );
nand NAND2_14520 ( P1_U4304 , P1_REIP_REG_18_ , P1_U4232 );
nand NAND2_14521 ( P1_U4305 , P1_ADDRESS_REG_17_ , P1_U3249 );
nand NAND2_14522 ( P1_U4306 , P1_REIP_REG_18_ , P1_U4233 );
nand NAND2_14523 ( P1_U4307 , P1_REIP_REG_17_ , P1_U4232 );
nand NAND2_14524 ( P1_U4308 , P1_ADDRESS_REG_16_ , P1_U3249 );
nand NAND2_14525 ( P1_U4309 , P1_REIP_REG_17_ , P1_U4233 );
nand NAND2_14526 ( P1_U4310 , P1_REIP_REG_16_ , P1_U4232 );
nand NAND2_14527 ( P1_U4311 , P1_ADDRESS_REG_15_ , P1_U3249 );
nand NAND2_14528 ( P1_U4312 , P1_REIP_REG_16_ , P1_U4233 );
nand NAND2_14529 ( P1_U4313 , P1_REIP_REG_15_ , P1_U4232 );
nand NAND2_14530 ( P1_U4314 , P1_ADDRESS_REG_14_ , P1_U3249 );
nand NAND2_14531 ( P1_U4315 , P1_REIP_REG_15_ , P1_U4233 );
nand NAND2_14532 ( P1_U4316 , P1_REIP_REG_14_ , P1_U4232 );
nand NAND2_14533 ( P1_U4317 , P1_ADDRESS_REG_13_ , P1_U3249 );
nand NAND2_14534 ( P1_U4318 , P1_REIP_REG_14_ , P1_U4233 );
nand NAND2_14535 ( P1_U4319 , P1_REIP_REG_13_ , P1_U4232 );
nand NAND2_14536 ( P1_U4320 , P1_ADDRESS_REG_12_ , P1_U3249 );
nand NAND2_14537 ( P1_U4321 , P1_REIP_REG_13_ , P1_U4233 );
nand NAND2_14538 ( P1_U4322 , P1_REIP_REG_12_ , P1_U4232 );
nand NAND2_14539 ( P1_U4323 , P1_ADDRESS_REG_11_ , P1_U3249 );
nand NAND2_14540 ( P1_U4324 , P1_REIP_REG_12_ , P1_U4233 );
nand NAND2_14541 ( P1_U4325 , P1_REIP_REG_11_ , P1_U4232 );
nand NAND2_14542 ( P1_U4326 , P1_ADDRESS_REG_10_ , P1_U3249 );
nand NAND2_14543 ( P1_U4327 , P1_REIP_REG_11_ , P1_U4233 );
nand NAND2_14544 ( P1_U4328 , P1_REIP_REG_10_ , P1_U4232 );
nand NAND2_14545 ( P1_U4329 , P1_ADDRESS_REG_9_ , P1_U3249 );
nand NAND2_14546 ( P1_U4330 , P1_REIP_REG_10_ , P1_U4233 );
nand NAND2_14547 ( P1_U4331 , P1_REIP_REG_9_ , P1_U4232 );
nand NAND2_14548 ( P1_U4332 , P1_ADDRESS_REG_8_ , P1_U3249 );
nand NAND2_14549 ( P1_U4333 , P1_REIP_REG_9_ , P1_U4233 );
nand NAND2_14550 ( P1_U4334 , P1_REIP_REG_8_ , P1_U4232 );
nand NAND2_14551 ( P1_U4335 , P1_ADDRESS_REG_7_ , P1_U3249 );
nand NAND2_14552 ( P1_U4336 , P1_REIP_REG_8_ , P1_U4233 );
nand NAND2_14553 ( P1_U4337 , P1_REIP_REG_7_ , P1_U4232 );
nand NAND2_14554 ( P1_U4338 , P1_ADDRESS_REG_6_ , P1_U3249 );
nand NAND2_14555 ( P1_U4339 , P1_REIP_REG_7_ , P1_U4233 );
nand NAND2_14556 ( P1_U4340 , P1_REIP_REG_6_ , P1_U4232 );
nand NAND2_14557 ( P1_U4341 , P1_ADDRESS_REG_5_ , P1_U3249 );
nand NAND2_14558 ( P1_U4342 , P1_REIP_REG_6_ , P1_U4233 );
nand NAND2_14559 ( P1_U4343 , P1_REIP_REG_5_ , P1_U4232 );
nand NAND2_14560 ( P1_U4344 , P1_ADDRESS_REG_4_ , P1_U3249 );
nand NAND2_14561 ( P1_U4345 , P1_REIP_REG_5_ , P1_U4233 );
nand NAND2_14562 ( P1_U4346 , P1_REIP_REG_4_ , P1_U4232 );
nand NAND2_14563 ( P1_U4347 , P1_ADDRESS_REG_3_ , P1_U3249 );
nand NAND2_14564 ( P1_U4348 , P1_REIP_REG_4_ , P1_U4233 );
nand NAND2_14565 ( P1_U4349 , P1_REIP_REG_3_ , P1_U4232 );
nand NAND2_14566 ( P1_U4350 , P1_ADDRESS_REG_2_ , P1_U3249 );
nand NAND2_14567 ( P1_U4351 , P1_REIP_REG_3_ , P1_U4233 );
nand NAND2_14568 ( P1_U4352 , P1_REIP_REG_2_ , P1_U4232 );
nand NAND2_14569 ( P1_U4353 , P1_ADDRESS_REG_1_ , P1_U3249 );
nand NAND2_14570 ( P1_U4354 , P1_REIP_REG_2_ , P1_U4233 );
nand NAND2_14571 ( P1_U4355 , P1_REIP_REG_1_ , P1_U4232 );
nand NAND2_14572 ( P1_U4356 , P1_ADDRESS_REG_0_ , P1_U3249 );
not NOT1_14573 ( P1_U4357 , P1_U3260 );
nand NAND2_14574 ( P1_U4358 , P1_U4357 , P1_U3257 );
nand NAND2_14575 ( P1_U4359 , NA , P1_U4258 );
not NOT1_14576 ( P1_U4360 , P1_U3261 );
nand NAND2_14577 ( P1_U4361 , P1_U4360 , P1_U3257 );
or OR2_14578 ( P1_U4362 , P1_STATE_REG_0_ , NA );
nand NAND3_14579 ( P1_U4363 , P1_U7622 , P1_U4362 , P1_U7623 );
not NOT1_14580 ( P1_U4364 , P1_U3255 );
nand NAND3_14581 ( P1_U4365 , HOLD , P1_U3247 , P1_U4364 );
nand NAND3_14582 ( P1_U4366 , P1_STATE_REG_1_ , P1_U3261 , U210 );
nand NAND2_14583 ( P1_U4367 , P1_U4366 , P1_U4365 );
nand NAND3_14584 ( P1_U4368 , P1_STATE_REG_0_ , P1_U4359 , P1_U4367 );
nand NAND2_14585 ( P1_U4369 , P1_STATE_REG_2_ , P1_U4363 );
nand NAND2_14586 ( P1_U4370 , U210 , P1_U4221 );
nand NAND2_14587 ( P1_U4371 , P1_U3496 , P1_U7625 );
nand NAND2_14588 ( P1_U4372 , P1_STATE_REG_2_ , P1_U3260 );
nand NAND2_14589 ( P1_U4373 , NA , P1_U3258 );
nand NAND2_14590 ( P1_U4374 , P1_U4373 , P1_U4372 );
nand NAND2_14591 ( P1_U4375 , P1_U4374 , P1_U3248 );
nand NAND2_14592 ( P1_U4376 , P1_U4179 , P1_U3255 );
not NOT1_14593 ( P1_U4377 , P1_U3280 );
not NOT1_14594 ( P1_U4378 , P1_U3269 );
not NOT1_14595 ( P1_U4379 , P1_U3444 );
not NOT1_14596 ( P1_U4380 , P1_U3268 );
not NOT1_14597 ( P1_U4381 , P1_U3274 );
not NOT1_14598 ( P1_U4382 , P1_U3267 );
nand NAND2_14599 ( P1_U4383 , P1_INSTQUEUE_REG_7__3_ , P1_U4382 );
nand NAND2_14600 ( P1_U4384 , P1_INSTQUEUE_REG_0__3_ , P1_U2472 );
nand NAND2_14601 ( P1_U4385 , P1_INSTQUEUE_REG_1__3_ , P1_U2471 );
nand NAND2_14602 ( P1_U4386 , P1_INSTQUEUE_REG_2__3_ , P1_U2470 );
nand NAND2_14603 ( P1_U4387 , P1_INSTQUEUE_REG_3__3_ , P1_U2468 );
nand NAND2_14604 ( P1_U4388 , P1_INSTQUEUE_REG_4__3_ , P1_U2467 );
nand NAND2_14605 ( P1_U4389 , P1_INSTQUEUE_REG_5__3_ , P1_U2466 );
nand NAND2_14606 ( P1_U4390 , P1_INSTQUEUE_REG_6__3_ , P1_U2465 );
nand NAND2_14607 ( P1_U4391 , P1_INSTQUEUE_REG_8__3_ , P1_U2464 );
nand NAND2_14608 ( P1_U4392 , P1_INSTQUEUE_REG_9__3_ , P1_U2463 );
nand NAND2_14609 ( P1_U4393 , P1_INSTQUEUE_REG_10__3_ , P1_U2461 );
nand NAND2_14610 ( P1_U4394 , P1_INSTQUEUE_REG_11__3_ , P1_U2459 );
nand NAND2_14611 ( P1_U4395 , P1_INSTQUEUE_REG_12__3_ , P1_U2458 );
nand NAND2_14612 ( P1_U4396 , P1_INSTQUEUE_REG_13__3_ , P1_U2457 );
nand NAND2_14613 ( P1_U4397 , P1_INSTQUEUE_REG_14__3_ , P1_U2455 );
nand NAND2_14614 ( P1_U4398 , P1_INSTQUEUE_REG_15__3_ , P1_U2453 );
not NOT1_14615 ( P1_U4399 , P1_U3283 );
not NOT1_14616 ( P1_U4400 , P1_U3278 );
nand NAND5_14617 ( P1_U4401 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3270 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUE_REG_7__5_ , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND3_14618 ( P1_U4402 , P1_INSTQUEUE_REG_0__5_ , P1_U3270 , P1_U4380 );
nand NAND4_14619 ( P1_U4403 , P1_INSTQUEUE_REG_1__5_ , P1_U2469 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_U3265 );
nand NAND4_14620 ( P1_U4404 , P1_INSTQUEUE_REG_2__5_ , P1_U2469 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3266 );
nand NAND4_14621 ( P1_U4405 , P1_INSTQUEUE_REG_4__5_ , P1_U4378 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3270 );
nand NAND3_14622 ( P1_U4406 , P1_U3520 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3521 );
nand NAND3_14623 ( P1_U4407 , P1_U3522 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3523 );
nand NAND2_14624 ( P1_U4408 , P1_U3524 , P1_U4380 );
nand NAND3_14625 ( P1_U4409 , P1_U3525 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3526 );
nand NAND5_14626 ( P1_U4410 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3264 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUE_REG_11__5_ , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND3_14627 ( P1_U4411 , P1_U4378 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3527 );
nand NAND5_14628 ( P1_U4412 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3265 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUE_REG_13__5_ , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_14629 ( P1_U4413 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3266 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUE_REG_14__5_ , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_14630 ( P1_U4414 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUE_REG_15__5_ , P1_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_14631 ( P1_U4415 , P1_U4173 );
nand NAND2_14632 ( P1_U4416 , P1_INSTQUEUE_REG_7__2_ , P1_U4382 );
nand NAND2_14633 ( P1_U4417 , P1_INSTQUEUE_REG_0__2_ , P1_U2472 );
nand NAND2_14634 ( P1_U4418 , P1_INSTQUEUE_REG_1__2_ , P1_U2471 );
nand NAND2_14635 ( P1_U4419 , P1_INSTQUEUE_REG_2__2_ , P1_U2470 );
nand NAND2_14636 ( P1_U4420 , P1_INSTQUEUE_REG_3__2_ , P1_U2468 );
nand NAND2_14637 ( P1_U4421 , P1_INSTQUEUE_REG_4__2_ , P1_U2467 );
nand NAND2_14638 ( P1_U4422 , P1_INSTQUEUE_REG_5__2_ , P1_U2466 );
nand NAND2_14639 ( P1_U4423 , P1_INSTQUEUE_REG_6__2_ , P1_U2465 );
nand NAND2_14640 ( P1_U4424 , P1_INSTQUEUE_REG_8__2_ , P1_U2464 );
nand NAND2_14641 ( P1_U4425 , P1_INSTQUEUE_REG_9__2_ , P1_U2463 );
nand NAND2_14642 ( P1_U4426 , P1_INSTQUEUE_REG_10__2_ , P1_U2461 );
nand NAND2_14643 ( P1_U4427 , P1_INSTQUEUE_REG_11__2_ , P1_U2459 );
nand NAND2_14644 ( P1_U4428 , P1_INSTQUEUE_REG_12__2_ , P1_U2458 );
nand NAND2_14645 ( P1_U4429 , P1_INSTQUEUE_REG_13__2_ , P1_U2457 );
nand NAND2_14646 ( P1_U4430 , P1_INSTQUEUE_REG_14__2_ , P1_U2455 );
nand NAND2_14647 ( P1_U4431 , P1_INSTQUEUE_REG_15__2_ , P1_U2453 );
not NOT1_14648 ( P1_U4432 , P1_U4171 );
nand NAND2_14649 ( P1_U4433 , P1_INSTQUEUE_REG_7__7_ , P1_U4382 );
nand NAND2_14650 ( P1_U4434 , P1_INSTQUEUE_REG_0__7_ , P1_U2472 );
nand NAND2_14651 ( P1_U4435 , P1_INSTQUEUE_REG_1__7_ , P1_U2471 );
nand NAND2_14652 ( P1_U4436 , P1_INSTQUEUE_REG_2__7_ , P1_U2470 );
nand NAND2_14653 ( P1_U4437 , P1_INSTQUEUE_REG_3__7_ , P1_U2468 );
nand NAND2_14654 ( P1_U4438 , P1_INSTQUEUE_REG_4__7_ , P1_U2467 );
nand NAND2_14655 ( P1_U4439 , P1_INSTQUEUE_REG_5__7_ , P1_U2466 );
nand NAND2_14656 ( P1_U4440 , P1_INSTQUEUE_REG_6__7_ , P1_U2465 );
nand NAND2_14657 ( P1_U4441 , P1_INSTQUEUE_REG_8__7_ , P1_U2464 );
nand NAND2_14658 ( P1_U4442 , P1_INSTQUEUE_REG_9__7_ , P1_U2463 );
nand NAND2_14659 ( P1_U4443 , P1_INSTQUEUE_REG_10__7_ , P1_U2461 );
nand NAND2_14660 ( P1_U4444 , P1_INSTQUEUE_REG_11__7_ , P1_U2459 );
nand NAND2_14661 ( P1_U4445 , P1_INSTQUEUE_REG_12__7_ , P1_U2458 );
nand NAND2_14662 ( P1_U4446 , P1_INSTQUEUE_REG_13__7_ , P1_U2457 );
nand NAND2_14663 ( P1_U4447 , P1_INSTQUEUE_REG_14__7_ , P1_U2455 );
nand NAND2_14664 ( P1_U4448 , P1_INSTQUEUE_REG_15__7_ , P1_U2453 );
not NOT1_14665 ( P1_U4449 , P1_U3391 );
nand NAND3_14666 ( P1_U4450 , P1_U3498 , P1_U4381 , P1_INSTQUEUE_REG_7__6_ );
nand NAND3_14667 ( P1_U4451 , P1_INSTQUEUE_REG_1__6_ , P1_U2469 , P1_U2456 );
nand NAND3_14668 ( P1_U4452 , P1_INSTQUEUE_REG_2__6_ , P1_U2469 , P1_U2454 );
nand NAND3_14669 ( P1_U4453 , P1_INSTQUEUE_REG_4__6_ , P1_U4378 , P1_U4381 );
nand NAND3_14670 ( P1_U4454 , P1_U2456 , P1_U4381 , P1_INSTQUEUE_REG_5__6_ );
nand NAND3_14671 ( P1_U4455 , P1_U2454 , P1_U4381 , P1_INSTQUEUE_REG_6__6_ );
nand NAND3_14672 ( P1_U4456 , P1_INSTQUEUE_REG_12__6_ , P1_U4378 , P1_U3507 );
nand NAND3_14673 ( P1_U4457 , P1_U3507 , P1_U2456 , P1_INSTQUEUE_REG_13__6_ );
nand NAND3_14674 ( P1_U4458 , P1_U3507 , P1_U2454 , P1_INSTQUEUE_REG_14__6_ );
nand NAND3_14675 ( P1_U4459 , P1_U3507 , P1_U3498 , P1_INSTQUEUE_REG_15__6_ );
not NOT1_14676 ( P1_U4460 , P1_U3277 );
nand NAND2_14677 ( P1_U4461 , P1_INSTQUEUE_REG_7__1_ , P1_U4382 );
nand NAND2_14678 ( P1_U4462 , P1_INSTQUEUE_REG_0__1_ , P1_U2472 );
nand NAND2_14679 ( P1_U4463 , P1_INSTQUEUE_REG_1__1_ , P1_U2471 );
nand NAND2_14680 ( P1_U4464 , P1_INSTQUEUE_REG_2__1_ , P1_U2470 );
nand NAND2_14681 ( P1_U4465 , P1_INSTQUEUE_REG_3__1_ , P1_U2468 );
nand NAND2_14682 ( P1_U4466 , P1_INSTQUEUE_REG_4__1_ , P1_U2467 );
nand NAND2_14683 ( P1_U4467 , P1_INSTQUEUE_REG_5__1_ , P1_U2466 );
nand NAND2_14684 ( P1_U4468 , P1_INSTQUEUE_REG_6__1_ , P1_U2465 );
nand NAND2_14685 ( P1_U4469 , P1_INSTQUEUE_REG_8__1_ , P1_U2464 );
nand NAND2_14686 ( P1_U4470 , P1_INSTQUEUE_REG_9__1_ , P1_U2463 );
nand NAND2_14687 ( P1_U4471 , P1_INSTQUEUE_REG_10__1_ , P1_U2461 );
nand NAND2_14688 ( P1_U4472 , P1_INSTQUEUE_REG_11__1_ , P1_U2459 );
nand NAND2_14689 ( P1_U4473 , P1_INSTQUEUE_REG_12__1_ , P1_U2458 );
nand NAND2_14690 ( P1_U4474 , P1_INSTQUEUE_REG_13__1_ , P1_U2457 );
nand NAND2_14691 ( P1_U4475 , P1_INSTQUEUE_REG_14__1_ , P1_U2455 );
nand NAND2_14692 ( P1_U4476 , P1_INSTQUEUE_REG_15__1_ , P1_U2453 );
not NOT1_14693 ( P1_U4477 , P1_U3271 );
nand NAND2_14694 ( P1_U4478 , P1_INSTQUEUE_REG_7__0_ , P1_U4382 );
nand NAND2_14695 ( P1_U4479 , P1_INSTQUEUE_REG_0__0_ , P1_U2472 );
nand NAND2_14696 ( P1_U4480 , P1_INSTQUEUE_REG_1__0_ , P1_U2471 );
nand NAND2_14697 ( P1_U4481 , P1_INSTQUEUE_REG_2__0_ , P1_U2470 );
nand NAND2_14698 ( P1_U4482 , P1_INSTQUEUE_REG_3__0_ , P1_U2468 );
nand NAND2_14699 ( P1_U4483 , P1_INSTQUEUE_REG_4__0_ , P1_U2467 );
nand NAND2_14700 ( P1_U4484 , P1_INSTQUEUE_REG_5__0_ , P1_U2466 );
nand NAND2_14701 ( P1_U4485 , P1_INSTQUEUE_REG_6__0_ , P1_U2465 );
nand NAND2_14702 ( P1_U4486 , P1_INSTQUEUE_REG_8__0_ , P1_U2464 );
nand NAND2_14703 ( P1_U4487 , P1_INSTQUEUE_REG_9__0_ , P1_U2463 );
nand NAND2_14704 ( P1_U4488 , P1_INSTQUEUE_REG_10__0_ , P1_U2461 );
nand NAND2_14705 ( P1_U4489 , P1_INSTQUEUE_REG_11__0_ , P1_U2459 );
nand NAND2_14706 ( P1_U4490 , P1_INSTQUEUE_REG_12__0_ , P1_U2458 );
nand NAND2_14707 ( P1_U4491 , P1_INSTQUEUE_REG_13__0_ , P1_U2457 );
nand NAND2_14708 ( P1_U4492 , P1_INSTQUEUE_REG_14__0_ , P1_U2455 );
nand NAND2_14709 ( P1_U4493 , P1_INSTQUEUE_REG_15__0_ , P1_U2453 );
not NOT1_14710 ( P1_U4494 , P1_U3284 );
nand NAND2_14711 ( P1_U4495 , P1_STATE_REG_2_ , P1_U3248 );
nand NAND2_14712 ( P1_U4496 , P1_U3254 , P1_U4495 );
not NOT1_14713 ( P1_U4497 , P1_U3272 );
nand NAND2_14714 ( P1_U4498 , P1_U4477 , P1_U3388 );
not NOT1_14715 ( P1_U4499 , P1_U3437 );
nand NAND3_14716 ( P1_U4500 , P1_U3272 , P1_U3390 , P1_U3287 );
nand NAND2_14717 ( P1_U4501 , P1_U4500 , P1_U3257 );
not NOT1_14718 ( P1_U4502 , P1_U3285 );
nand NAND2_14719 ( P1_U4503 , P1_U4460 , P1_U4173 );
nand NAND2_14720 ( P1_U4504 , P1_U4196 , P1_U3286 );
nand NAND2_14721 ( P1_U4505 , P1_U4504 , P1_U3579 );
nand NAND2_14722 ( P1_U4506 , P1_U3580 , P1_U4505 );
nand NAND2_14723 ( P1_U4507 , P1_U4215 , P1_U3388 );
nand NAND3_14724 ( P1_U4508 , P1_U7682 , P1_U7681 , P1_U4507 );
nand NAND2_14725 ( P1_U4509 , P1_U2448 , P1_U4262 );
or OR2_14726 ( P1_U4510 , P1_MORE_REG , P1_FLUSH_REG );
not NOT1_14727 ( P1_U4511 , P1_U3293 );
nand NAND2_14728 ( P1_U4512 , P1_U4511 , P1_U3262 );
nand NAND2_14729 ( P1_U4513 , P1_STATE2_REG_1_ , U210 );
not NOT1_14730 ( P1_U4514 , P1_U3295 );
nand NAND3_14731 ( P1_U4515 , P1_U7688 , P1_U7687 , P1_STATE2_REG_1_ );
nand NAND2_14732 ( P1_U4516 , P1_STATE2_REG_2_ , P1_U3295 );
nand NAND2_14733 ( P1_U4517 , P1_U7604 , P1_U4246 );
nand NAND2_14734 ( P1_U4518 , P1_U3583 , P1_U4514 );
nand NAND2_14735 ( P1_U4519 , P1_STATE2_REG_1_ , P1_U4517 );
nand NAND2_14736 ( P1_U4520 , P1_U2368 , P1_U7604 );
nand NAND2_14737 ( P1_U4521 , P1_U4252 , P1_U4261 );
nand NAND2_14738 ( P1_U4522 , P1_U7604 , P1_U4245 );
nand NAND2_14739 ( P1_U4523 , P1_U2368 , P1_U3293 );
not NOT1_14740 ( P1_U4524 , P1_U3325 );
not NOT1_14741 ( P1_U4525 , P1_U3331 );
not NOT1_14742 ( P1_U4526 , P1_U3332 );
not NOT1_14743 ( P1_U4527 , P1_U3314 );
not NOT1_14744 ( P1_U4528 , P1_U3313 );
not NOT1_14745 ( P1_U4529 , P1_U3342 );
nand NAND2_14746 ( P1_U4530 , P1_R2144_U8 , P1_U3313 );
not NOT1_14747 ( P1_U4531 , P1_U3358 );
not NOT1_14748 ( P1_U4532 , P1_U3315 );
not NOT1_14749 ( P1_U4533 , P1_U3305 );
not NOT1_14750 ( P1_U4534 , P1_U3306 );
nand NAND2_14751 ( P1_U4535 , P1_U2438 , P1_U2442 );
not NOT1_14752 ( P1_U4536 , P1_U3321 );
not NOT1_14753 ( P1_U4537 , P1_U3356 );
not NOT1_14754 ( P1_U4538 , P1_U3340 );
nand NAND2_14755 ( P1_U4539 , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_U3305 );
not NOT1_14756 ( P1_U4540 , P1_U3360 );
not NOT1_14757 ( P1_U4541 , P1_U3329 );
not NOT1_14758 ( P1_U4542 , P1_U3323 );
not NOT1_14759 ( P1_U4543 , P1_U3235 );
nand NAND2_14760 ( P1_U4544 , P1_U2432 , P1_U2436 );
not NOT1_14761 ( P1_U4545 , P1_U3322 );
nand NAND2_14762 ( P1_U4546 , P1_STATE2_REG_1_ , P1_U3263 );
nand NAND3_14763 ( P1_U4547 , P1_U4546 , P1_U3297 , P1_U3299 );
nand NAND2_14764 ( P1_U4548 , P1_U4528 , P1_U2476 );
nand NAND2_14765 ( P1_U4549 , P1_U2480 , P1_U2358 );
nand NAND2_14766 ( P1_U4550 , P1_U3320 , P1_U4549 );
nand NAND2_14767 ( P1_U4551 , P1_U4536 , P1_U4550 );
nand NAND2_14768 ( P1_U4552 , P1_STATE2_REG_3_ , P1_U3306 );
nand NAND2_14769 ( P1_U4553 , P1_U4545 , P1_STATE2_REG_2_ );
nand NAND2_14770 ( P1_U4554 , P1_U4551 , P1_U3587 );
nand NAND2_14771 ( P1_U4555 , P1_U2480 , P1_U2388 );
nand NAND2_14772 ( P1_U4556 , P1_U3320 , P1_U4555 );
nand NAND2_14773 ( P1_U4557 , P1_U4556 , P1_U3321 );
nand NAND2_14774 ( P1_U4558 , P1_STATE2_REG_2_ , P1_U3322 );
nand NAND2_14775 ( P1_U4559 , P1_U4558 , P1_U4557 );
nand NAND2_14776 ( P1_U4560 , P1_U2415 , P1_U4534 );
nand NAND2_14777 ( P1_U4561 , P1_U2413 , P1_U2477 );
nand NAND2_14778 ( P1_U4562 , P1_U2412 , P1_U4532 );
nand NAND2_14779 ( P1_U4563 , P1_U2397 , P1_U4559 );
nand NAND2_14780 ( P1_U4564 , P1_INSTQUEUE_REG_15__7_ , P1_U4554 );
nand NAND2_14781 ( P1_U4565 , P1_U2416 , P1_U4534 );
nand NAND2_14782 ( P1_U4566 , P1_U2411 , P1_U2477 );
nand NAND2_14783 ( P1_U4567 , P1_U2410 , P1_U4532 );
nand NAND2_14784 ( P1_U4568 , P1_U2396 , P1_U4559 );
nand NAND2_14785 ( P1_U4569 , P1_INSTQUEUE_REG_15__6_ , P1_U4554 );
nand NAND2_14786 ( P1_U4570 , P1_U2420 , P1_U4534 );
nand NAND2_14787 ( P1_U4571 , P1_U2409 , P1_U2477 );
nand NAND2_14788 ( P1_U4572 , P1_U2408 , P1_U4532 );
nand NAND2_14789 ( P1_U4573 , P1_U2395 , P1_U4559 );
nand NAND2_14790 ( P1_U4574 , P1_INSTQUEUE_REG_15__5_ , P1_U4554 );
nand NAND2_14791 ( P1_U4575 , P1_U2419 , P1_U4534 );
nand NAND2_14792 ( P1_U4576 , P1_U2407 , P1_U2477 );
nand NAND2_14793 ( P1_U4577 , P1_U2406 , P1_U4532 );
nand NAND2_14794 ( P1_U4578 , P1_U2394 , P1_U4559 );
nand NAND2_14795 ( P1_U4579 , P1_INSTQUEUE_REG_15__4_ , P1_U4554 );
nand NAND2_14796 ( P1_U4580 , P1_U2418 , P1_U4534 );
nand NAND2_14797 ( P1_U4581 , P1_U2405 , P1_U2477 );
nand NAND2_14798 ( P1_U4582 , P1_U2404 , P1_U4532 );
nand NAND2_14799 ( P1_U4583 , P1_U2393 , P1_U4559 );
nand NAND2_14800 ( P1_U4584 , P1_INSTQUEUE_REG_15__3_ , P1_U4554 );
nand NAND2_14801 ( P1_U4585 , P1_U2421 , P1_U4534 );
nand NAND2_14802 ( P1_U4586 , P1_U2403 , P1_U2477 );
nand NAND2_14803 ( P1_U4587 , P1_U2402 , P1_U4532 );
nand NAND2_14804 ( P1_U4588 , P1_U2392 , P1_U4559 );
nand NAND2_14805 ( P1_U4589 , P1_INSTQUEUE_REG_15__2_ , P1_U4554 );
nand NAND2_14806 ( P1_U4590 , P1_U2414 , P1_U4534 );
nand NAND2_14807 ( P1_U4591 , P1_U2401 , P1_U2477 );
nand NAND2_14808 ( P1_U4592 , P1_U2400 , P1_U4532 );
nand NAND2_14809 ( P1_U4593 , P1_U2391 , P1_U4559 );
nand NAND2_14810 ( P1_U4594 , P1_INSTQUEUE_REG_15__1_ , P1_U4554 );
nand NAND2_14811 ( P1_U4595 , P1_U2417 , P1_U4534 );
nand NAND2_14812 ( P1_U4596 , P1_U2399 , P1_U2477 );
nand NAND2_14813 ( P1_U4597 , P1_U2398 , P1_U4532 );
nand NAND2_14814 ( P1_U4598 , P1_U2390 , P1_U4559 );
nand NAND2_14815 ( P1_U4599 , P1_INSTQUEUE_REG_15__0_ , P1_U4554 );
not NOT1_14816 ( P1_U4600 , P1_U3326 );
not NOT1_14817 ( P1_U4601 , P1_U3327 );
not NOT1_14818 ( P1_U4602 , P1_U3324 );
nand NAND2_14819 ( P1_U4603 , P1_U2443 , P1_U2438 );
not NOT1_14820 ( P1_U4604 , P1_U3328 );
not NOT1_14821 ( P1_U4605 , P1_U3236 );
nand NAND2_14822 ( P1_U4606 , P1_U4524 , P1_U2476 );
nand NAND2_14823 ( P1_U4607 , P1_U2482 , P1_U2358 );
nand NAND2_14824 ( P1_U4608 , P1_U3320 , P1_U4607 );
nand NAND2_14825 ( P1_U4609 , P1_U4604 , P1_U4608 );
nand NAND2_14826 ( P1_U4610 , P1_STATE2_REG_3_ , P1_U3324 );
nand NAND2_14827 ( P1_U4611 , P1_STATE2_REG_2_ , P1_U3236 );
nand NAND2_14828 ( P1_U4612 , P1_U4609 , P1_U3596 );
nand NAND2_14829 ( P1_U4613 , P1_U2482 , P1_U2388 );
nand NAND2_14830 ( P1_U4614 , P1_U3320 , P1_U4613 );
nand NAND2_14831 ( P1_U4615 , P1_U4614 , P1_U3328 );
nand NAND2_14832 ( P1_U4616 , P1_STATE2_REG_2_ , P1_U4605 );
nand NAND2_14833 ( P1_U4617 , P1_U4616 , P1_U4615 );
nand NAND2_14834 ( P1_U4618 , P1_U4602 , P1_U2415 );
nand NAND2_14835 ( P1_U4619 , P1_U2481 , P1_U2413 );
nand NAND2_14836 ( P1_U4620 , P1_U4601 , P1_U2412 );
nand NAND2_14837 ( P1_U4621 , P1_U2397 , P1_U4617 );
nand NAND2_14838 ( P1_U4622 , P1_INSTQUEUE_REG_14__7_ , P1_U4612 );
nand NAND2_14839 ( P1_U4623 , P1_U4602 , P1_U2416 );
nand NAND2_14840 ( P1_U4624 , P1_U2481 , P1_U2411 );
nand NAND2_14841 ( P1_U4625 , P1_U4601 , P1_U2410 );
nand NAND2_14842 ( P1_U4626 , P1_U2396 , P1_U4617 );
nand NAND2_14843 ( P1_U4627 , P1_INSTQUEUE_REG_14__6_ , P1_U4612 );
nand NAND2_14844 ( P1_U4628 , P1_U4602 , P1_U2420 );
nand NAND2_14845 ( P1_U4629 , P1_U2481 , P1_U2409 );
nand NAND2_14846 ( P1_U4630 , P1_U4601 , P1_U2408 );
nand NAND2_14847 ( P1_U4631 , P1_U2395 , P1_U4617 );
nand NAND2_14848 ( P1_U4632 , P1_INSTQUEUE_REG_14__5_ , P1_U4612 );
nand NAND2_14849 ( P1_U4633 , P1_U4602 , P1_U2419 );
nand NAND2_14850 ( P1_U4634 , P1_U2481 , P1_U2407 );
nand NAND2_14851 ( P1_U4635 , P1_U4601 , P1_U2406 );
nand NAND2_14852 ( P1_U4636 , P1_U2394 , P1_U4617 );
nand NAND2_14853 ( P1_U4637 , P1_INSTQUEUE_REG_14__4_ , P1_U4612 );
nand NAND2_14854 ( P1_U4638 , P1_U4602 , P1_U2418 );
nand NAND2_14855 ( P1_U4639 , P1_U2481 , P1_U2405 );
nand NAND2_14856 ( P1_U4640 , P1_U4601 , P1_U2404 );
nand NAND2_14857 ( P1_U4641 , P1_U2393 , P1_U4617 );
nand NAND2_14858 ( P1_U4642 , P1_INSTQUEUE_REG_14__3_ , P1_U4612 );
nand NAND2_14859 ( P1_U4643 , P1_U4602 , P1_U2421 );
nand NAND2_14860 ( P1_U4644 , P1_U2481 , P1_U2403 );
nand NAND2_14861 ( P1_U4645 , P1_U4601 , P1_U2402 );
nand NAND2_14862 ( P1_U4646 , P1_U2392 , P1_U4617 );
nand NAND2_14863 ( P1_U4647 , P1_INSTQUEUE_REG_14__2_ , P1_U4612 );
nand NAND2_14864 ( P1_U4648 , P1_U4602 , P1_U2414 );
nand NAND2_14865 ( P1_U4649 , P1_U2481 , P1_U2401 );
nand NAND2_14866 ( P1_U4650 , P1_U4601 , P1_U2400 );
nand NAND2_14867 ( P1_U4651 , P1_U2391 , P1_U4617 );
nand NAND2_14868 ( P1_U4652 , P1_INSTQUEUE_REG_14__1_ , P1_U4612 );
nand NAND2_14869 ( P1_U4653 , P1_U4602 , P1_U2417 );
nand NAND2_14870 ( P1_U4654 , P1_U2481 , P1_U2399 );
nand NAND2_14871 ( P1_U4655 , P1_U4601 , P1_U2398 );
nand NAND2_14872 ( P1_U4656 , P1_U2390 , P1_U4617 );
nand NAND2_14873 ( P1_U4657 , P1_INSTQUEUE_REG_14__0_ , P1_U4612 );
not NOT1_14874 ( P1_U4658 , P1_U3333 );
not NOT1_14875 ( P1_U4659 , P1_U3334 );
not NOT1_14876 ( P1_U4660 , P1_U3330 );
nand NAND2_14877 ( P1_U4661 , P1_U2444 , P1_U2438 );
not NOT1_14878 ( P1_U4662 , P1_U3335 );
nand NAND2_14879 ( P1_U4663 , P1_U2437 , P1_U2432 );
not NOT1_14880 ( P1_U4664 , P1_U3336 );
nand NAND2_14881 ( P1_U4665 , P1_U4525 , P1_U2476 );
nand NAND2_14882 ( P1_U4666 , P1_U2484 , P1_U2358 );
nand NAND2_14883 ( P1_U4667 , P1_U3320 , P1_U4666 );
nand NAND2_14884 ( P1_U4668 , P1_U4662 , P1_U4667 );
nand NAND2_14885 ( P1_U4669 , P1_STATE2_REG_3_ , P1_U3330 );
nand NAND2_14886 ( P1_U4670 , P1_U4664 , P1_STATE2_REG_2_ );
nand NAND2_14887 ( P1_U4671 , P1_U4668 , P1_U3605 );
nand NAND2_14888 ( P1_U4672 , P1_U2484 , P1_U2388 );
nand NAND2_14889 ( P1_U4673 , P1_U3320 , P1_U4672 );
nand NAND2_14890 ( P1_U4674 , P1_U4673 , P1_U3335 );
nand NAND2_14891 ( P1_U4675 , P1_STATE2_REG_2_ , P1_U3336 );
nand NAND2_14892 ( P1_U4676 , P1_U4675 , P1_U4674 );
nand NAND2_14893 ( P1_U4677 , P1_U4660 , P1_U2415 );
nand NAND2_14894 ( P1_U4678 , P1_U2483 , P1_U2413 );
nand NAND2_14895 ( P1_U4679 , P1_U4659 , P1_U2412 );
nand NAND2_14896 ( P1_U4680 , P1_U2397 , P1_U4676 );
nand NAND2_14897 ( P1_U4681 , P1_INSTQUEUE_REG_13__7_ , P1_U4671 );
nand NAND2_14898 ( P1_U4682 , P1_U4660 , P1_U2416 );
nand NAND2_14899 ( P1_U4683 , P1_U2483 , P1_U2411 );
nand NAND2_14900 ( P1_U4684 , P1_U4659 , P1_U2410 );
nand NAND2_14901 ( P1_U4685 , P1_U2396 , P1_U4676 );
nand NAND2_14902 ( P1_U4686 , P1_INSTQUEUE_REG_13__6_ , P1_U4671 );
nand NAND2_14903 ( P1_U4687 , P1_U4660 , P1_U2420 );
nand NAND2_14904 ( P1_U4688 , P1_U2483 , P1_U2409 );
nand NAND2_14905 ( P1_U4689 , P1_U4659 , P1_U2408 );
nand NAND2_14906 ( P1_U4690 , P1_U2395 , P1_U4676 );
nand NAND2_14907 ( P1_U4691 , P1_INSTQUEUE_REG_13__5_ , P1_U4671 );
nand NAND2_14908 ( P1_U4692 , P1_U4660 , P1_U2419 );
nand NAND2_14909 ( P1_U4693 , P1_U2483 , P1_U2407 );
nand NAND2_14910 ( P1_U4694 , P1_U4659 , P1_U2406 );
nand NAND2_14911 ( P1_U4695 , P1_U2394 , P1_U4676 );
nand NAND2_14912 ( P1_U4696 , P1_INSTQUEUE_REG_13__4_ , P1_U4671 );
nand NAND2_14913 ( P1_U4697 , P1_U4660 , P1_U2418 );
nand NAND2_14914 ( P1_U4698 , P1_U2483 , P1_U2405 );
nand NAND2_14915 ( P1_U4699 , P1_U4659 , P1_U2404 );
nand NAND2_14916 ( P1_U4700 , P1_U2393 , P1_U4676 );
nand NAND2_14917 ( P1_U4701 , P1_INSTQUEUE_REG_13__3_ , P1_U4671 );
nand NAND2_14918 ( P1_U4702 , P1_U4660 , P1_U2421 );
nand NAND2_14919 ( P1_U4703 , P1_U2483 , P1_U2403 );
nand NAND2_14920 ( P1_U4704 , P1_U4659 , P1_U2402 );
nand NAND2_14921 ( P1_U4705 , P1_U2392 , P1_U4676 );
nand NAND2_14922 ( P1_U4706 , P1_INSTQUEUE_REG_13__2_ , P1_U4671 );
nand NAND2_14923 ( P1_U4707 , P1_U4660 , P1_U2414 );
nand NAND2_14924 ( P1_U4708 , P1_U2483 , P1_U2401 );
nand NAND2_14925 ( P1_U4709 , P1_U4659 , P1_U2400 );
nand NAND2_14926 ( P1_U4710 , P1_U2391 , P1_U4676 );
nand NAND2_14927 ( P1_U4711 , P1_INSTQUEUE_REG_13__1_ , P1_U4671 );
nand NAND2_14928 ( P1_U4712 , P1_U4660 , P1_U2417 );
nand NAND2_14929 ( P1_U4713 , P1_U2483 , P1_U2399 );
nand NAND2_14930 ( P1_U4714 , P1_U4659 , P1_U2398 );
nand NAND2_14931 ( P1_U4715 , P1_U2390 , P1_U4676 );
nand NAND2_14932 ( P1_U4716 , P1_INSTQUEUE_REG_13__0_ , P1_U4671 );
not NOT1_14933 ( P1_U4717 , P1_U3338 );
not NOT1_14934 ( P1_U4718 , P1_U3337 );
nand NAND2_14935 ( P1_U4719 , P1_U2445 , P1_U2438 );
not NOT1_14936 ( P1_U4720 , P1_U3339 );
not NOT1_14937 ( P1_U4721 , P1_U3237 );
nand NAND2_14938 ( P1_U4722 , P1_U2486 , P1_U2476 );
nand NAND2_14939 ( P1_U4723 , P1_U2489 , P1_U2358 );
nand NAND2_14940 ( P1_U4724 , P1_U3320 , P1_U4723 );
nand NAND2_14941 ( P1_U4725 , P1_U4720 , P1_U4724 );
nand NAND2_14942 ( P1_U4726 , P1_STATE2_REG_3_ , P1_U3337 );
nand NAND2_14943 ( P1_U4727 , P1_STATE2_REG_2_ , P1_U3237 );
nand NAND2_14944 ( P1_U4728 , P1_U4725 , P1_U3614 );
nand NAND2_14945 ( P1_U4729 , P1_U2489 , P1_U2388 );
nand NAND2_14946 ( P1_U4730 , P1_U3320 , P1_U4729 );
nand NAND2_14947 ( P1_U4731 , P1_U4730 , P1_U3339 );
nand NAND2_14948 ( P1_U4732 , P1_STATE2_REG_2_ , P1_U4721 );
nand NAND2_14949 ( P1_U4733 , P1_U4732 , P1_U4731 );
nand NAND2_14950 ( P1_U4734 , P1_U4718 , P1_U2415 );
nand NAND2_14951 ( P1_U4735 , P1_U2487 , P1_U2413 );
nand NAND2_14952 ( P1_U4736 , P1_U4717 , P1_U2412 );
nand NAND2_14953 ( P1_U4737 , P1_U2397 , P1_U4733 );
nand NAND2_14954 ( P1_U4738 , P1_INSTQUEUE_REG_12__7_ , P1_U4728 );
nand NAND2_14955 ( P1_U4739 , P1_U4718 , P1_U2416 );
nand NAND2_14956 ( P1_U4740 , P1_U2487 , P1_U2411 );
nand NAND2_14957 ( P1_U4741 , P1_U4717 , P1_U2410 );
nand NAND2_14958 ( P1_U4742 , P1_U2396 , P1_U4733 );
nand NAND2_14959 ( P1_U4743 , P1_INSTQUEUE_REG_12__6_ , P1_U4728 );
nand NAND2_14960 ( P1_U4744 , P1_U4718 , P1_U2420 );
nand NAND2_14961 ( P1_U4745 , P1_U2487 , P1_U2409 );
nand NAND2_14962 ( P1_U4746 , P1_U4717 , P1_U2408 );
nand NAND2_14963 ( P1_U4747 , P1_U2395 , P1_U4733 );
nand NAND2_14964 ( P1_U4748 , P1_INSTQUEUE_REG_12__5_ , P1_U4728 );
nand NAND2_14965 ( P1_U4749 , P1_U4718 , P1_U2419 );
nand NAND2_14966 ( P1_U4750 , P1_U2487 , P1_U2407 );
nand NAND2_14967 ( P1_U4751 , P1_U4717 , P1_U2406 );
nand NAND2_14968 ( P1_U4752 , P1_U2394 , P1_U4733 );
nand NAND2_14969 ( P1_U4753 , P1_INSTQUEUE_REG_12__4_ , P1_U4728 );
nand NAND2_14970 ( P1_U4754 , P1_U4718 , P1_U2418 );
nand NAND2_14971 ( P1_U4755 , P1_U2487 , P1_U2405 );
nand NAND2_14972 ( P1_U4756 , P1_U4717 , P1_U2404 );
nand NAND2_14973 ( P1_U4757 , P1_U2393 , P1_U4733 );
nand NAND2_14974 ( P1_U4758 , P1_INSTQUEUE_REG_12__3_ , P1_U4728 );
nand NAND2_14975 ( P1_U4759 , P1_U4718 , P1_U2421 );
nand NAND2_14976 ( P1_U4760 , P1_U2487 , P1_U2403 );
nand NAND2_14977 ( P1_U4761 , P1_U4717 , P1_U2402 );
nand NAND2_14978 ( P1_U4762 , P1_U2392 , P1_U4733 );
nand NAND2_14979 ( P1_U4763 , P1_INSTQUEUE_REG_12__2_ , P1_U4728 );
nand NAND2_14980 ( P1_U4764 , P1_U4718 , P1_U2414 );
nand NAND2_14981 ( P1_U4765 , P1_U2487 , P1_U2401 );
nand NAND2_14982 ( P1_U4766 , P1_U4717 , P1_U2400 );
nand NAND2_14983 ( P1_U4767 , P1_U2391 , P1_U4733 );
nand NAND2_14984 ( P1_U4768 , P1_INSTQUEUE_REG_12__1_ , P1_U4728 );
nand NAND2_14985 ( P1_U4769 , P1_U4718 , P1_U2417 );
nand NAND2_14986 ( P1_U4770 , P1_U2487 , P1_U2399 );
nand NAND2_14987 ( P1_U4771 , P1_U4717 , P1_U2398 );
nand NAND2_14988 ( P1_U4772 , P1_U2390 , P1_U4733 );
nand NAND2_14989 ( P1_U4773 , P1_INSTQUEUE_REG_12__0_ , P1_U4728 );
not NOT1_14990 ( P1_U4774 , P1_U3343 );
not NOT1_14991 ( P1_U4775 , P1_U3341 );
nand NAND2_14992 ( P1_U4776 , P1_U2440 , P1_U2442 );
not NOT1_14993 ( P1_U4777 , P1_U3344 );
nand NAND2_14994 ( P1_U4778 , P1_U2434 , P1_U2436 );
not NOT1_14995 ( P1_U4779 , P1_U3345 );
nand NAND2_14996 ( P1_U4780 , P1_U4529 , P1_U4528 );
nand NAND2_14997 ( P1_U4781 , P1_U2492 , P1_U2358 );
nand NAND2_14998 ( P1_U4782 , P1_U3320 , P1_U4781 );
nand NAND2_14999 ( P1_U4783 , P1_U4777 , P1_U4782 );
nand NAND2_15000 ( P1_U4784 , P1_STATE2_REG_3_ , P1_U3341 );
nand NAND2_15001 ( P1_U4785 , P1_U4779 , P1_STATE2_REG_2_ );
nand NAND2_15002 ( P1_U4786 , P1_U4783 , P1_U3623 );
nand NAND2_15003 ( P1_U4787 , P1_U2492 , P1_U2388 );
nand NAND2_15004 ( P1_U4788 , P1_U3320 , P1_U4787 );
nand NAND2_15005 ( P1_U4789 , P1_U4788 , P1_U3344 );
nand NAND2_15006 ( P1_U4790 , P1_STATE2_REG_2_ , P1_U3345 );
nand NAND2_15007 ( P1_U4791 , P1_U4790 , P1_U4789 );
nand NAND2_15008 ( P1_U4792 , P1_U4775 , P1_U2415 );
nand NAND2_15009 ( P1_U4793 , P1_U2491 , P1_U2413 );
nand NAND2_15010 ( P1_U4794 , P1_U4774 , P1_U2412 );
nand NAND2_15011 ( P1_U4795 , P1_U2397 , P1_U4791 );
nand NAND2_15012 ( P1_U4796 , P1_INSTQUEUE_REG_11__7_ , P1_U4786 );
nand NAND2_15013 ( P1_U4797 , P1_U4775 , P1_U2416 );
nand NAND2_15014 ( P1_U4798 , P1_U2491 , P1_U2411 );
nand NAND2_15015 ( P1_U4799 , P1_U4774 , P1_U2410 );
nand NAND2_15016 ( P1_U4800 , P1_U2396 , P1_U4791 );
nand NAND2_15017 ( P1_U4801 , P1_INSTQUEUE_REG_11__6_ , P1_U4786 );
nand NAND2_15018 ( P1_U4802 , P1_U4775 , P1_U2420 );
nand NAND2_15019 ( P1_U4803 , P1_U2491 , P1_U2409 );
nand NAND2_15020 ( P1_U4804 , P1_U4774 , P1_U2408 );
nand NAND2_15021 ( P1_U4805 , P1_U2395 , P1_U4791 );
nand NAND2_15022 ( P1_U4806 , P1_INSTQUEUE_REG_11__5_ , P1_U4786 );
nand NAND2_15023 ( P1_U4807 , P1_U4775 , P1_U2419 );
nand NAND2_15024 ( P1_U4808 , P1_U2491 , P1_U2407 );
nand NAND2_15025 ( P1_U4809 , P1_U4774 , P1_U2406 );
nand NAND2_15026 ( P1_U4810 , P1_U2394 , P1_U4791 );
nand NAND2_15027 ( P1_U4811 , P1_INSTQUEUE_REG_11__4_ , P1_U4786 );
nand NAND2_15028 ( P1_U4812 , P1_U4775 , P1_U2418 );
nand NAND2_15029 ( P1_U4813 , P1_U2491 , P1_U2405 );
nand NAND2_15030 ( P1_U4814 , P1_U4774 , P1_U2404 );
nand NAND2_15031 ( P1_U4815 , P1_U2393 , P1_U4791 );
nand NAND2_15032 ( P1_U4816 , P1_INSTQUEUE_REG_11__3_ , P1_U4786 );
nand NAND2_15033 ( P1_U4817 , P1_U4775 , P1_U2421 );
nand NAND2_15034 ( P1_U4818 , P1_U2491 , P1_U2403 );
nand NAND2_15035 ( P1_U4819 , P1_U4774 , P1_U2402 );
nand NAND2_15036 ( P1_U4820 , P1_U2392 , P1_U4791 );
nand NAND2_15037 ( P1_U4821 , P1_INSTQUEUE_REG_11__2_ , P1_U4786 );
nand NAND2_15038 ( P1_U4822 , P1_U4775 , P1_U2414 );
nand NAND2_15039 ( P1_U4823 , P1_U2491 , P1_U2401 );
nand NAND2_15040 ( P1_U4824 , P1_U4774 , P1_U2400 );
nand NAND2_15041 ( P1_U4825 , P1_U2391 , P1_U4791 );
nand NAND2_15042 ( P1_U4826 , P1_INSTQUEUE_REG_11__1_ , P1_U4786 );
nand NAND2_15043 ( P1_U4827 , P1_U4775 , P1_U2417 );
nand NAND2_15044 ( P1_U4828 , P1_U2491 , P1_U2399 );
nand NAND2_15045 ( P1_U4829 , P1_U4774 , P1_U2398 );
nand NAND2_15046 ( P1_U4830 , P1_U2390 , P1_U4791 );
nand NAND2_15047 ( P1_U4831 , P1_INSTQUEUE_REG_11__0_ , P1_U4786 );
not NOT1_15048 ( P1_U4832 , P1_U3347 );
not NOT1_15049 ( P1_U4833 , P1_U3346 );
nand NAND2_15050 ( P1_U4834 , P1_U2440 , P1_U2443 );
not NOT1_15051 ( P1_U4835 , P1_U3348 );
not NOT1_15052 ( P1_U4836 , P1_U3238 );
nand NAND2_15053 ( P1_U4837 , P1_U4529 , P1_U4524 );
nand NAND2_15054 ( P1_U4838 , P1_U2494 , P1_U2358 );
nand NAND2_15055 ( P1_U4839 , P1_U3320 , P1_U4838 );
nand NAND2_15056 ( P1_U4840 , P1_U4835 , P1_U4839 );
nand NAND2_15057 ( P1_U4841 , P1_STATE2_REG_3_ , P1_U3346 );
nand NAND2_15058 ( P1_U4842 , P1_STATE2_REG_2_ , P1_U3238 );
nand NAND2_15059 ( P1_U4843 , P1_U4840 , P1_U3632 );
nand NAND2_15060 ( P1_U4844 , P1_U2494 , P1_U2388 );
nand NAND2_15061 ( P1_U4845 , P1_U3320 , P1_U4844 );
nand NAND2_15062 ( P1_U4846 , P1_U4845 , P1_U3348 );
nand NAND2_15063 ( P1_U4847 , P1_STATE2_REG_2_ , P1_U4836 );
nand NAND2_15064 ( P1_U4848 , P1_U4847 , P1_U4846 );
nand NAND2_15065 ( P1_U4849 , P1_U4833 , P1_U2415 );
nand NAND2_15066 ( P1_U4850 , P1_U2493 , P1_U2413 );
nand NAND2_15067 ( P1_U4851 , P1_U4832 , P1_U2412 );
nand NAND2_15068 ( P1_U4852 , P1_U2397 , P1_U4848 );
nand NAND2_15069 ( P1_U4853 , P1_INSTQUEUE_REG_10__7_ , P1_U4843 );
nand NAND2_15070 ( P1_U4854 , P1_U4833 , P1_U2416 );
nand NAND2_15071 ( P1_U4855 , P1_U2493 , P1_U2411 );
nand NAND2_15072 ( P1_U4856 , P1_U4832 , P1_U2410 );
nand NAND2_15073 ( P1_U4857 , P1_U2396 , P1_U4848 );
nand NAND2_15074 ( P1_U4858 , P1_INSTQUEUE_REG_10__6_ , P1_U4843 );
nand NAND2_15075 ( P1_U4859 , P1_U4833 , P1_U2420 );
nand NAND2_15076 ( P1_U4860 , P1_U2493 , P1_U2409 );
nand NAND2_15077 ( P1_U4861 , P1_U4832 , P1_U2408 );
nand NAND2_15078 ( P1_U4862 , P1_U2395 , P1_U4848 );
nand NAND2_15079 ( P1_U4863 , P1_INSTQUEUE_REG_10__5_ , P1_U4843 );
nand NAND2_15080 ( P1_U4864 , P1_U4833 , P1_U2419 );
nand NAND2_15081 ( P1_U4865 , P1_U2493 , P1_U2407 );
nand NAND2_15082 ( P1_U4866 , P1_U4832 , P1_U2406 );
nand NAND2_15083 ( P1_U4867 , P1_U2394 , P1_U4848 );
nand NAND2_15084 ( P1_U4868 , P1_INSTQUEUE_REG_10__4_ , P1_U4843 );
nand NAND2_15085 ( P1_U4869 , P1_U4833 , P1_U2418 );
nand NAND2_15086 ( P1_U4870 , P1_U2493 , P1_U2405 );
nand NAND2_15087 ( P1_U4871 , P1_U4832 , P1_U2404 );
nand NAND2_15088 ( P1_U4872 , P1_U2393 , P1_U4848 );
nand NAND2_15089 ( P1_U4873 , P1_INSTQUEUE_REG_10__3_ , P1_U4843 );
nand NAND2_15090 ( P1_U4874 , P1_U4833 , P1_U2421 );
nand NAND2_15091 ( P1_U4875 , P1_U2493 , P1_U2403 );
nand NAND2_15092 ( P1_U4876 , P1_U4832 , P1_U2402 );
nand NAND2_15093 ( P1_U4877 , P1_U2392 , P1_U4848 );
nand NAND2_15094 ( P1_U4878 , P1_INSTQUEUE_REG_10__2_ , P1_U4843 );
nand NAND2_15095 ( P1_U4879 , P1_U4833 , P1_U2414 );
nand NAND2_15096 ( P1_U4880 , P1_U2493 , P1_U2401 );
nand NAND2_15097 ( P1_U4881 , P1_U4832 , P1_U2400 );
nand NAND2_15098 ( P1_U4882 , P1_U2391 , P1_U4848 );
nand NAND2_15099 ( P1_U4883 , P1_INSTQUEUE_REG_10__1_ , P1_U4843 );
nand NAND2_15100 ( P1_U4884 , P1_U4833 , P1_U2417 );
nand NAND2_15101 ( P1_U4885 , P1_U2493 , P1_U2399 );
nand NAND2_15102 ( P1_U4886 , P1_U4832 , P1_U2398 );
nand NAND2_15103 ( P1_U4887 , P1_U2390 , P1_U4848 );
nand NAND2_15104 ( P1_U4888 , P1_INSTQUEUE_REG_10__0_ , P1_U4843 );
not NOT1_15105 ( P1_U4889 , P1_U3350 );
not NOT1_15106 ( P1_U4890 , P1_U3349 );
nand NAND2_15107 ( P1_U4891 , P1_U2440 , P1_U2444 );
not NOT1_15108 ( P1_U4892 , P1_U3351 );
nand NAND2_15109 ( P1_U4893 , P1_U2434 , P1_U2437 );
not NOT1_15110 ( P1_U4894 , P1_U3352 );
nand NAND2_15111 ( P1_U4895 , P1_U4529 , P1_U4525 );
nand NAND2_15112 ( P1_U4896 , P1_U2496 , P1_U2358 );
nand NAND2_15113 ( P1_U4897 , P1_U3320 , P1_U4896 );
nand NAND2_15114 ( P1_U4898 , P1_U4892 , P1_U4897 );
nand NAND2_15115 ( P1_U4899 , P1_STATE2_REG_3_ , P1_U3349 );
nand NAND2_15116 ( P1_U4900 , P1_U4894 , P1_STATE2_REG_2_ );
nand NAND2_15117 ( P1_U4901 , P1_U4898 , P1_U3641 );
nand NAND2_15118 ( P1_U4902 , P1_U2496 , P1_U2388 );
nand NAND2_15119 ( P1_U4903 , P1_U3320 , P1_U4902 );
nand NAND2_15120 ( P1_U4904 , P1_U4903 , P1_U3351 );
nand NAND2_15121 ( P1_U4905 , P1_STATE2_REG_2_ , P1_U3352 );
nand NAND2_15122 ( P1_U4906 , P1_U4905 , P1_U4904 );
nand NAND2_15123 ( P1_U4907 , P1_U4890 , P1_U2415 );
nand NAND2_15124 ( P1_U4908 , P1_U2495 , P1_U2413 );
nand NAND2_15125 ( P1_U4909 , P1_U4889 , P1_U2412 );
nand NAND2_15126 ( P1_U4910 , P1_U2397 , P1_U4906 );
nand NAND2_15127 ( P1_U4911 , P1_INSTQUEUE_REG_9__7_ , P1_U4901 );
nand NAND2_15128 ( P1_U4912 , P1_U4890 , P1_U2416 );
nand NAND2_15129 ( P1_U4913 , P1_U2495 , P1_U2411 );
nand NAND2_15130 ( P1_U4914 , P1_U4889 , P1_U2410 );
nand NAND2_15131 ( P1_U4915 , P1_U2396 , P1_U4906 );
nand NAND2_15132 ( P1_U4916 , P1_INSTQUEUE_REG_9__6_ , P1_U4901 );
nand NAND2_15133 ( P1_U4917 , P1_U4890 , P1_U2420 );
nand NAND2_15134 ( P1_U4918 , P1_U2495 , P1_U2409 );
nand NAND2_15135 ( P1_U4919 , P1_U4889 , P1_U2408 );
nand NAND2_15136 ( P1_U4920 , P1_U2395 , P1_U4906 );
nand NAND2_15137 ( P1_U4921 , P1_INSTQUEUE_REG_9__5_ , P1_U4901 );
nand NAND2_15138 ( P1_U4922 , P1_U4890 , P1_U2419 );
nand NAND2_15139 ( P1_U4923 , P1_U2495 , P1_U2407 );
nand NAND2_15140 ( P1_U4924 , P1_U4889 , P1_U2406 );
nand NAND2_15141 ( P1_U4925 , P1_U2394 , P1_U4906 );
nand NAND2_15142 ( P1_U4926 , P1_INSTQUEUE_REG_9__4_ , P1_U4901 );
nand NAND2_15143 ( P1_U4927 , P1_U4890 , P1_U2418 );
nand NAND2_15144 ( P1_U4928 , P1_U2495 , P1_U2405 );
nand NAND2_15145 ( P1_U4929 , P1_U4889 , P1_U2404 );
nand NAND2_15146 ( P1_U4930 , P1_U2393 , P1_U4906 );
nand NAND2_15147 ( P1_U4931 , P1_INSTQUEUE_REG_9__3_ , P1_U4901 );
nand NAND2_15148 ( P1_U4932 , P1_U4890 , P1_U2421 );
nand NAND2_15149 ( P1_U4933 , P1_U2495 , P1_U2403 );
nand NAND2_15150 ( P1_U4934 , P1_U4889 , P1_U2402 );
nand NAND2_15151 ( P1_U4935 , P1_U2392 , P1_U4906 );
nand NAND2_15152 ( P1_U4936 , P1_INSTQUEUE_REG_9__2_ , P1_U4901 );
nand NAND2_15153 ( P1_U4937 , P1_U4890 , P1_U2414 );
nand NAND2_15154 ( P1_U4938 , P1_U2495 , P1_U2401 );
nand NAND2_15155 ( P1_U4939 , P1_U4889 , P1_U2400 );
nand NAND2_15156 ( P1_U4940 , P1_U2391 , P1_U4906 );
nand NAND2_15157 ( P1_U4941 , P1_INSTQUEUE_REG_9__1_ , P1_U4901 );
nand NAND2_15158 ( P1_U4942 , P1_U4890 , P1_U2417 );
nand NAND2_15159 ( P1_U4943 , P1_U2495 , P1_U2399 );
nand NAND2_15160 ( P1_U4944 , P1_U4889 , P1_U2398 );
nand NAND2_15161 ( P1_U4945 , P1_U2390 , P1_U4906 );
nand NAND2_15162 ( P1_U4946 , P1_INSTQUEUE_REG_9__0_ , P1_U4901 );
not NOT1_15163 ( P1_U4947 , P1_U3354 );
not NOT1_15164 ( P1_U4948 , P1_U3353 );
nand NAND2_15165 ( P1_U4949 , P1_U2440 , P1_U2445 );
not NOT1_15166 ( P1_U4950 , P1_U3355 );
not NOT1_15167 ( P1_U4951 , P1_U3239 );
nand NAND2_15168 ( P1_U4952 , P1_U4529 , P1_U2486 );
nand NAND2_15169 ( P1_U4953 , P1_U2498 , P1_U2358 );
nand NAND2_15170 ( P1_U4954 , P1_U3320 , P1_U4953 );
nand NAND2_15171 ( P1_U4955 , P1_U4950 , P1_U4954 );
nand NAND2_15172 ( P1_U4956 , P1_STATE2_REG_3_ , P1_U3353 );
nand NAND2_15173 ( P1_U4957 , P1_STATE2_REG_2_ , P1_U3239 );
nand NAND2_15174 ( P1_U4958 , P1_U4955 , P1_U3650 );
nand NAND2_15175 ( P1_U4959 , P1_U2498 , P1_U2388 );
nand NAND2_15176 ( P1_U4960 , P1_U3320 , P1_U4959 );
nand NAND2_15177 ( P1_U4961 , P1_U4960 , P1_U3355 );
nand NAND2_15178 ( P1_U4962 , P1_STATE2_REG_2_ , P1_U4951 );
nand NAND2_15179 ( P1_U4963 , P1_U4962 , P1_U4961 );
nand NAND2_15180 ( P1_U4964 , P1_U4948 , P1_U2415 );
nand NAND2_15181 ( P1_U4965 , P1_U2497 , P1_U2413 );
nand NAND2_15182 ( P1_U4966 , P1_U4947 , P1_U2412 );
nand NAND2_15183 ( P1_U4967 , P1_U2397 , P1_U4963 );
nand NAND2_15184 ( P1_U4968 , P1_INSTQUEUE_REG_8__7_ , P1_U4958 );
nand NAND2_15185 ( P1_U4969 , P1_U4948 , P1_U2416 );
nand NAND2_15186 ( P1_U4970 , P1_U2497 , P1_U2411 );
nand NAND2_15187 ( P1_U4971 , P1_U4947 , P1_U2410 );
nand NAND2_15188 ( P1_U4972 , P1_U2396 , P1_U4963 );
nand NAND2_15189 ( P1_U4973 , P1_INSTQUEUE_REG_8__6_ , P1_U4958 );
nand NAND2_15190 ( P1_U4974 , P1_U4948 , P1_U2420 );
nand NAND2_15191 ( P1_U4975 , P1_U2497 , P1_U2409 );
nand NAND2_15192 ( P1_U4976 , P1_U4947 , P1_U2408 );
nand NAND2_15193 ( P1_U4977 , P1_U2395 , P1_U4963 );
nand NAND2_15194 ( P1_U4978 , P1_INSTQUEUE_REG_8__5_ , P1_U4958 );
nand NAND2_15195 ( P1_U4979 , P1_U4948 , P1_U2419 );
nand NAND2_15196 ( P1_U4980 , P1_U2497 , P1_U2407 );
nand NAND2_15197 ( P1_U4981 , P1_U4947 , P1_U2406 );
nand NAND2_15198 ( P1_U4982 , P1_U2394 , P1_U4963 );
nand NAND2_15199 ( P1_U4983 , P1_INSTQUEUE_REG_8__4_ , P1_U4958 );
nand NAND2_15200 ( P1_U4984 , P1_U4948 , P1_U2418 );
nand NAND2_15201 ( P1_U4985 , P1_U2497 , P1_U2405 );
nand NAND2_15202 ( P1_U4986 , P1_U4947 , P1_U2404 );
nand NAND2_15203 ( P1_U4987 , P1_U2393 , P1_U4963 );
nand NAND2_15204 ( P1_U4988 , P1_INSTQUEUE_REG_8__3_ , P1_U4958 );
nand NAND2_15205 ( P1_U4989 , P1_U4948 , P1_U2421 );
nand NAND2_15206 ( P1_U4990 , P1_U2497 , P1_U2403 );
nand NAND2_15207 ( P1_U4991 , P1_U4947 , P1_U2402 );
nand NAND2_15208 ( P1_U4992 , P1_U2392 , P1_U4963 );
nand NAND2_15209 ( P1_U4993 , P1_INSTQUEUE_REG_8__2_ , P1_U4958 );
nand NAND2_15210 ( P1_U4994 , P1_U4948 , P1_U2414 );
nand NAND2_15211 ( P1_U4995 , P1_U2497 , P1_U2401 );
nand NAND2_15212 ( P1_U4996 , P1_U4947 , P1_U2400 );
nand NAND2_15213 ( P1_U4997 , P1_U2391 , P1_U4963 );
nand NAND2_15214 ( P1_U4998 , P1_INSTQUEUE_REG_8__1_ , P1_U4958 );
nand NAND2_15215 ( P1_U4999 , P1_U4948 , P1_U2417 );
nand NAND2_15216 ( P1_U5000 , P1_U2497 , P1_U2399 );
nand NAND2_15217 ( P1_U5001 , P1_U4947 , P1_U2398 );
nand NAND2_15218 ( P1_U5002 , P1_U2390 , P1_U4963 );
nand NAND2_15219 ( P1_U5003 , P1_INSTQUEUE_REG_8__0_ , P1_U4958 );
not NOT1_15220 ( P1_U5004 , P1_U3359 );
nand NAND2_15221 ( P1_U5005 , P1_U2439 , P1_U2442 );
not NOT1_15222 ( P1_U5006 , P1_U3361 );
nand NAND2_15223 ( P1_U5007 , P1_U2433 , P1_U2436 );
not NOT1_15224 ( P1_U5008 , P1_U3362 );
nand NAND2_15225 ( P1_U5009 , P1_U2500 , P1_U2358 );
nand NAND2_15226 ( P1_U5010 , P1_U3320 , P1_U5009 );
nand NAND2_15227 ( P1_U5011 , P1_U5006 , P1_U5010 );
nand NAND2_15228 ( P1_U5012 , P1_STATE2_REG_3_ , P1_U3356 );
nand NAND2_15229 ( P1_U5013 , P1_U5008 , P1_STATE2_REG_2_ );
nand NAND2_15230 ( P1_U5014 , P1_U5011 , P1_U3659 );
nand NAND2_15231 ( P1_U5015 , P1_U2500 , P1_U2388 );
nand NAND2_15232 ( P1_U5016 , P1_U3320 , P1_U5015 );
nand NAND2_15233 ( P1_U5017 , P1_U5016 , P1_U3361 );
nand NAND2_15234 ( P1_U5018 , P1_STATE2_REG_2_ , P1_U3362 );
nand NAND2_15235 ( P1_U5019 , P1_U5018 , P1_U5017 );
nand NAND2_15236 ( P1_U5020 , P1_U4537 , P1_U2415 );
nand NAND2_15237 ( P1_U5021 , P1_U4238 , P1_U2413 );
nand NAND2_15238 ( P1_U5022 , P1_U5004 , P1_U2412 );
nand NAND2_15239 ( P1_U5023 , P1_U2397 , P1_U5019 );
nand NAND2_15240 ( P1_U5024 , P1_INSTQUEUE_REG_7__7_ , P1_U5014 );
nand NAND2_15241 ( P1_U5025 , P1_U4537 , P1_U2416 );
nand NAND2_15242 ( P1_U5026 , P1_U4238 , P1_U2411 );
nand NAND2_15243 ( P1_U5027 , P1_U5004 , P1_U2410 );
nand NAND2_15244 ( P1_U5028 , P1_U2396 , P1_U5019 );
nand NAND2_15245 ( P1_U5029 , P1_INSTQUEUE_REG_7__6_ , P1_U5014 );
nand NAND2_15246 ( P1_U5030 , P1_U4537 , P1_U2420 );
nand NAND2_15247 ( P1_U5031 , P1_U4238 , P1_U2409 );
nand NAND2_15248 ( P1_U5032 , P1_U5004 , P1_U2408 );
nand NAND2_15249 ( P1_U5033 , P1_U2395 , P1_U5019 );
nand NAND2_15250 ( P1_U5034 , P1_INSTQUEUE_REG_7__5_ , P1_U5014 );
nand NAND2_15251 ( P1_U5035 , P1_U4537 , P1_U2419 );
nand NAND2_15252 ( P1_U5036 , P1_U4238 , P1_U2407 );
nand NAND2_15253 ( P1_U5037 , P1_U5004 , P1_U2406 );
nand NAND2_15254 ( P1_U5038 , P1_U2394 , P1_U5019 );
nand NAND2_15255 ( P1_U5039 , P1_INSTQUEUE_REG_7__4_ , P1_U5014 );
nand NAND2_15256 ( P1_U5040 , P1_U4537 , P1_U2418 );
nand NAND2_15257 ( P1_U5041 , P1_U4238 , P1_U2405 );
nand NAND2_15258 ( P1_U5042 , P1_U5004 , P1_U2404 );
nand NAND2_15259 ( P1_U5043 , P1_U2393 , P1_U5019 );
nand NAND2_15260 ( P1_U5044 , P1_INSTQUEUE_REG_7__3_ , P1_U5014 );
nand NAND2_15261 ( P1_U5045 , P1_U4537 , P1_U2421 );
nand NAND2_15262 ( P1_U5046 , P1_U4238 , P1_U2403 );
nand NAND2_15263 ( P1_U5047 , P1_U5004 , P1_U2402 );
nand NAND2_15264 ( P1_U5048 , P1_U2392 , P1_U5019 );
nand NAND2_15265 ( P1_U5049 , P1_INSTQUEUE_REG_7__2_ , P1_U5014 );
nand NAND2_15266 ( P1_U5050 , P1_U4537 , P1_U2414 );
nand NAND2_15267 ( P1_U5051 , P1_U4238 , P1_U2401 );
nand NAND2_15268 ( P1_U5052 , P1_U5004 , P1_U2400 );
nand NAND2_15269 ( P1_U5053 , P1_U2391 , P1_U5019 );
nand NAND2_15270 ( P1_U5054 , P1_INSTQUEUE_REG_7__1_ , P1_U5014 );
nand NAND2_15271 ( P1_U5055 , P1_U4537 , P1_U2417 );
nand NAND2_15272 ( P1_U5056 , P1_U4238 , P1_U2399 );
nand NAND2_15273 ( P1_U5057 , P1_U5004 , P1_U2398 );
nand NAND2_15274 ( P1_U5058 , P1_U2390 , P1_U5019 );
nand NAND2_15275 ( P1_U5059 , P1_INSTQUEUE_REG_7__0_ , P1_U5014 );
not NOT1_15276 ( P1_U5060 , P1_U3364 );
not NOT1_15277 ( P1_U5061 , P1_U3363 );
nand NAND2_15278 ( P1_U5062 , P1_U2439 , P1_U2443 );
not NOT1_15279 ( P1_U5063 , P1_U3365 );
not NOT1_15280 ( P1_U5064 , P1_U3240 );
nand NAND2_15281 ( P1_U5065 , P1_U4524 , P1_U2474 );
nand NAND2_15282 ( P1_U5066 , P1_U2502 , P1_U2358 );
nand NAND2_15283 ( P1_U5067 , P1_U3320 , P1_U5066 );
nand NAND2_15284 ( P1_U5068 , P1_U5063 , P1_U5067 );
nand NAND2_15285 ( P1_U5069 , P1_STATE2_REG_3_ , P1_U3363 );
nand NAND2_15286 ( P1_U5070 , P1_STATE2_REG_2_ , P1_U3240 );
nand NAND2_15287 ( P1_U5071 , P1_U5068 , P1_U3668 );
nand NAND2_15288 ( P1_U5072 , P1_U2502 , P1_U2388 );
nand NAND2_15289 ( P1_U5073 , P1_U3320 , P1_U5072 );
nand NAND2_15290 ( P1_U5074 , P1_U5073 , P1_U3365 );
nand NAND2_15291 ( P1_U5075 , P1_STATE2_REG_2_ , P1_U5064 );
nand NAND2_15292 ( P1_U5076 , P1_U5075 , P1_U5074 );
nand NAND2_15293 ( P1_U5077 , P1_U5061 , P1_U2415 );
nand NAND2_15294 ( P1_U5078 , P1_U2501 , P1_U2413 );
nand NAND2_15295 ( P1_U5079 , P1_U5060 , P1_U2412 );
nand NAND2_15296 ( P1_U5080 , P1_U2397 , P1_U5076 );
nand NAND2_15297 ( P1_U5081 , P1_INSTQUEUE_REG_6__7_ , P1_U5071 );
nand NAND2_15298 ( P1_U5082 , P1_U5061 , P1_U2416 );
nand NAND2_15299 ( P1_U5083 , P1_U2501 , P1_U2411 );
nand NAND2_15300 ( P1_U5084 , P1_U5060 , P1_U2410 );
nand NAND2_15301 ( P1_U5085 , P1_U2396 , P1_U5076 );
nand NAND2_15302 ( P1_U5086 , P1_INSTQUEUE_REG_6__6_ , P1_U5071 );
nand NAND2_15303 ( P1_U5087 , P1_U5061 , P1_U2420 );
nand NAND2_15304 ( P1_U5088 , P1_U2501 , P1_U2409 );
nand NAND2_15305 ( P1_U5089 , P1_U5060 , P1_U2408 );
nand NAND2_15306 ( P1_U5090 , P1_U2395 , P1_U5076 );
nand NAND2_15307 ( P1_U5091 , P1_INSTQUEUE_REG_6__5_ , P1_U5071 );
nand NAND2_15308 ( P1_U5092 , P1_U5061 , P1_U2419 );
nand NAND2_15309 ( P1_U5093 , P1_U2501 , P1_U2407 );
nand NAND2_15310 ( P1_U5094 , P1_U5060 , P1_U2406 );
nand NAND2_15311 ( P1_U5095 , P1_U2394 , P1_U5076 );
nand NAND2_15312 ( P1_U5096 , P1_INSTQUEUE_REG_6__4_ , P1_U5071 );
nand NAND2_15313 ( P1_U5097 , P1_U5061 , P1_U2418 );
nand NAND2_15314 ( P1_U5098 , P1_U2501 , P1_U2405 );
nand NAND2_15315 ( P1_U5099 , P1_U5060 , P1_U2404 );
nand NAND2_15316 ( P1_U5100 , P1_U2393 , P1_U5076 );
nand NAND2_15317 ( P1_U5101 , P1_INSTQUEUE_REG_6__3_ , P1_U5071 );
nand NAND2_15318 ( P1_U5102 , P1_U5061 , P1_U2421 );
nand NAND2_15319 ( P1_U5103 , P1_U2501 , P1_U2403 );
nand NAND2_15320 ( P1_U5104 , P1_U5060 , P1_U2402 );
nand NAND2_15321 ( P1_U5105 , P1_U2392 , P1_U5076 );
nand NAND2_15322 ( P1_U5106 , P1_INSTQUEUE_REG_6__2_ , P1_U5071 );
nand NAND2_15323 ( P1_U5107 , P1_U5061 , P1_U2414 );
nand NAND2_15324 ( P1_U5108 , P1_U2501 , P1_U2401 );
nand NAND2_15325 ( P1_U5109 , P1_U5060 , P1_U2400 );
nand NAND2_15326 ( P1_U5110 , P1_U2391 , P1_U5076 );
nand NAND2_15327 ( P1_U5111 , P1_INSTQUEUE_REG_6__1_ , P1_U5071 );
nand NAND2_15328 ( P1_U5112 , P1_U5061 , P1_U2417 );
nand NAND2_15329 ( P1_U5113 , P1_U2501 , P1_U2399 );
nand NAND2_15330 ( P1_U5114 , P1_U5060 , P1_U2398 );
nand NAND2_15331 ( P1_U5115 , P1_U2390 , P1_U5076 );
nand NAND2_15332 ( P1_U5116 , P1_INSTQUEUE_REG_6__0_ , P1_U5071 );
not NOT1_15333 ( P1_U5117 , P1_U3367 );
not NOT1_15334 ( P1_U5118 , P1_U3366 );
nand NAND2_15335 ( P1_U5119 , P1_U2439 , P1_U2444 );
not NOT1_15336 ( P1_U5120 , P1_U3368 );
nand NAND2_15337 ( P1_U5121 , P1_U2433 , P1_U2437 );
not NOT1_15338 ( P1_U5122 , P1_U3369 );
nand NAND2_15339 ( P1_U5123 , P1_U4525 , P1_U2474 );
nand NAND2_15340 ( P1_U5124 , P1_U2504 , P1_U2358 );
nand NAND2_15341 ( P1_U5125 , P1_U3320 , P1_U5124 );
nand NAND2_15342 ( P1_U5126 , P1_U5120 , P1_U5125 );
nand NAND2_15343 ( P1_U5127 , P1_STATE2_REG_3_ , P1_U3366 );
nand NAND2_15344 ( P1_U5128 , P1_U5122 , P1_STATE2_REG_2_ );
nand NAND2_15345 ( P1_U5129 , P1_U5126 , P1_U3677 );
nand NAND2_15346 ( P1_U5130 , P1_U2504 , P1_U2388 );
nand NAND2_15347 ( P1_U5131 , P1_U3320 , P1_U5130 );
nand NAND2_15348 ( P1_U5132 , P1_U5131 , P1_U3368 );
nand NAND2_15349 ( P1_U5133 , P1_STATE2_REG_2_ , P1_U3369 );
nand NAND2_15350 ( P1_U5134 , P1_U5133 , P1_U5132 );
nand NAND2_15351 ( P1_U5135 , P1_U5118 , P1_U2415 );
nand NAND2_15352 ( P1_U5136 , P1_U2503 , P1_U2413 );
nand NAND2_15353 ( P1_U5137 , P1_U5117 , P1_U2412 );
nand NAND2_15354 ( P1_U5138 , P1_U2397 , P1_U5134 );
nand NAND2_15355 ( P1_U5139 , P1_INSTQUEUE_REG_5__7_ , P1_U5129 );
nand NAND2_15356 ( P1_U5140 , P1_U5118 , P1_U2416 );
nand NAND2_15357 ( P1_U5141 , P1_U2503 , P1_U2411 );
nand NAND2_15358 ( P1_U5142 , P1_U5117 , P1_U2410 );
nand NAND2_15359 ( P1_U5143 , P1_U2396 , P1_U5134 );
nand NAND2_15360 ( P1_U5144 , P1_INSTQUEUE_REG_5__6_ , P1_U5129 );
nand NAND2_15361 ( P1_U5145 , P1_U5118 , P1_U2420 );
nand NAND2_15362 ( P1_U5146 , P1_U2503 , P1_U2409 );
nand NAND2_15363 ( P1_U5147 , P1_U5117 , P1_U2408 );
nand NAND2_15364 ( P1_U5148 , P1_U2395 , P1_U5134 );
nand NAND2_15365 ( P1_U5149 , P1_INSTQUEUE_REG_5__5_ , P1_U5129 );
nand NAND2_15366 ( P1_U5150 , P1_U5118 , P1_U2419 );
nand NAND2_15367 ( P1_U5151 , P1_U2503 , P1_U2407 );
nand NAND2_15368 ( P1_U5152 , P1_U5117 , P1_U2406 );
nand NAND2_15369 ( P1_U5153 , P1_U2394 , P1_U5134 );
nand NAND2_15370 ( P1_U5154 , P1_INSTQUEUE_REG_5__4_ , P1_U5129 );
nand NAND2_15371 ( P1_U5155 , P1_U5118 , P1_U2418 );
nand NAND2_15372 ( P1_U5156 , P1_U2503 , P1_U2405 );
nand NAND2_15373 ( P1_U5157 , P1_U5117 , P1_U2404 );
nand NAND2_15374 ( P1_U5158 , P1_U2393 , P1_U5134 );
nand NAND2_15375 ( P1_U5159 , P1_INSTQUEUE_REG_5__3_ , P1_U5129 );
nand NAND2_15376 ( P1_U5160 , P1_U5118 , P1_U2421 );
nand NAND2_15377 ( P1_U5161 , P1_U2503 , P1_U2403 );
nand NAND2_15378 ( P1_U5162 , P1_U5117 , P1_U2402 );
nand NAND2_15379 ( P1_U5163 , P1_U2392 , P1_U5134 );
nand NAND2_15380 ( P1_U5164 , P1_INSTQUEUE_REG_5__2_ , P1_U5129 );
nand NAND2_15381 ( P1_U5165 , P1_U5118 , P1_U2414 );
nand NAND2_15382 ( P1_U5166 , P1_U2503 , P1_U2401 );
nand NAND2_15383 ( P1_U5167 , P1_U5117 , P1_U2400 );
nand NAND2_15384 ( P1_U5168 , P1_U2391 , P1_U5134 );
nand NAND2_15385 ( P1_U5169 , P1_INSTQUEUE_REG_5__1_ , P1_U5129 );
nand NAND2_15386 ( P1_U5170 , P1_U5118 , P1_U2417 );
nand NAND2_15387 ( P1_U5171 , P1_U2503 , P1_U2399 );
nand NAND2_15388 ( P1_U5172 , P1_U5117 , P1_U2398 );
nand NAND2_15389 ( P1_U5173 , P1_U2390 , P1_U5134 );
nand NAND2_15390 ( P1_U5174 , P1_INSTQUEUE_REG_5__0_ , P1_U5129 );
not NOT1_15391 ( P1_U5175 , P1_U3371 );
not NOT1_15392 ( P1_U5176 , P1_U3370 );
nand NAND2_15393 ( P1_U5177 , P1_U2439 , P1_U2445 );
not NOT1_15394 ( P1_U5178 , P1_U3372 );
not NOT1_15395 ( P1_U5179 , P1_U3241 );
nand NAND2_15396 ( P1_U5180 , P1_U2486 , P1_U2474 );
nand NAND2_15397 ( P1_U5181 , P1_U2506 , P1_U2358 );
nand NAND2_15398 ( P1_U5182 , P1_U3320 , P1_U5181 );
nand NAND2_15399 ( P1_U5183 , P1_U5178 , P1_U5182 );
nand NAND2_15400 ( P1_U5184 , P1_STATE2_REG_3_ , P1_U3370 );
nand NAND2_15401 ( P1_U5185 , P1_STATE2_REG_2_ , P1_U3241 );
nand NAND2_15402 ( P1_U5186 , P1_U5183 , P1_U3686 );
nand NAND2_15403 ( P1_U5187 , P1_U2506 , P1_U2388 );
nand NAND2_15404 ( P1_U5188 , P1_U3320 , P1_U5187 );
nand NAND2_15405 ( P1_U5189 , P1_U5188 , P1_U3372 );
nand NAND2_15406 ( P1_U5190 , P1_STATE2_REG_2_ , P1_U5179 );
nand NAND2_15407 ( P1_U5191 , P1_U5190 , P1_U5189 );
nand NAND2_15408 ( P1_U5192 , P1_U5176 , P1_U2415 );
nand NAND2_15409 ( P1_U5193 , P1_U2505 , P1_U2413 );
nand NAND2_15410 ( P1_U5194 , P1_U5175 , P1_U2412 );
nand NAND2_15411 ( P1_U5195 , P1_U2397 , P1_U5191 );
nand NAND2_15412 ( P1_U5196 , P1_INSTQUEUE_REG_4__7_ , P1_U5186 );
nand NAND2_15413 ( P1_U5197 , P1_U5176 , P1_U2416 );
nand NAND2_15414 ( P1_U5198 , P1_U2505 , P1_U2411 );
nand NAND2_15415 ( P1_U5199 , P1_U5175 , P1_U2410 );
nand NAND2_15416 ( P1_U5200 , P1_U2396 , P1_U5191 );
nand NAND2_15417 ( P1_U5201 , P1_INSTQUEUE_REG_4__6_ , P1_U5186 );
nand NAND2_15418 ( P1_U5202 , P1_U5176 , P1_U2420 );
nand NAND2_15419 ( P1_U5203 , P1_U2505 , P1_U2409 );
nand NAND2_15420 ( P1_U5204 , P1_U5175 , P1_U2408 );
nand NAND2_15421 ( P1_U5205 , P1_U2395 , P1_U5191 );
nand NAND2_15422 ( P1_U5206 , P1_INSTQUEUE_REG_4__5_ , P1_U5186 );
nand NAND2_15423 ( P1_U5207 , P1_U5176 , P1_U2419 );
nand NAND2_15424 ( P1_U5208 , P1_U2505 , P1_U2407 );
nand NAND2_15425 ( P1_U5209 , P1_U5175 , P1_U2406 );
nand NAND2_15426 ( P1_U5210 , P1_U2394 , P1_U5191 );
nand NAND2_15427 ( P1_U5211 , P1_INSTQUEUE_REG_4__4_ , P1_U5186 );
nand NAND2_15428 ( P1_U5212 , P1_U5176 , P1_U2418 );
nand NAND2_15429 ( P1_U5213 , P1_U2505 , P1_U2405 );
nand NAND2_15430 ( P1_U5214 , P1_U5175 , P1_U2404 );
nand NAND2_15431 ( P1_U5215 , P1_U2393 , P1_U5191 );
nand NAND2_15432 ( P1_U5216 , P1_INSTQUEUE_REG_4__3_ , P1_U5186 );
nand NAND2_15433 ( P1_U5217 , P1_U5176 , P1_U2421 );
nand NAND2_15434 ( P1_U5218 , P1_U2505 , P1_U2403 );
nand NAND2_15435 ( P1_U5219 , P1_U5175 , P1_U2402 );
nand NAND2_15436 ( P1_U5220 , P1_U2392 , P1_U5191 );
nand NAND2_15437 ( P1_U5221 , P1_INSTQUEUE_REG_4__2_ , P1_U5186 );
nand NAND2_15438 ( P1_U5222 , P1_U5176 , P1_U2414 );
nand NAND2_15439 ( P1_U5223 , P1_U2505 , P1_U2401 );
nand NAND2_15440 ( P1_U5224 , P1_U5175 , P1_U2400 );
nand NAND2_15441 ( P1_U5225 , P1_U2391 , P1_U5191 );
nand NAND2_15442 ( P1_U5226 , P1_INSTQUEUE_REG_4__1_ , P1_U5186 );
nand NAND2_15443 ( P1_U5227 , P1_U5176 , P1_U2417 );
nand NAND2_15444 ( P1_U5228 , P1_U2505 , P1_U2399 );
nand NAND2_15445 ( P1_U5229 , P1_U5175 , P1_U2398 );
nand NAND2_15446 ( P1_U5230 , P1_U2390 , P1_U5191 );
nand NAND2_15447 ( P1_U5231 , P1_INSTQUEUE_REG_4__0_ , P1_U5186 );
not NOT1_15448 ( P1_U5232 , P1_U3374 );
not NOT1_15449 ( P1_U5233 , P1_U3373 );
nand NAND2_15450 ( P1_U5234 , P1_U2441 , P1_U2442 );
not NOT1_15451 ( P1_U5235 , P1_U3375 );
nand NAND2_15452 ( P1_U5236 , P1_U2435 , P1_U2436 );
not NOT1_15453 ( P1_U5237 , P1_U3376 );
nand NAND2_15454 ( P1_U5238 , P1_U2508 , P1_U4528 );
nand NAND2_15455 ( P1_U5239 , P1_U2511 , P1_U2358 );
nand NAND2_15456 ( P1_U5240 , P1_U3320 , P1_U5239 );
nand NAND2_15457 ( P1_U5241 , P1_U5235 , P1_U5240 );
nand NAND2_15458 ( P1_U5242 , P1_STATE2_REG_3_ , P1_U3373 );
nand NAND2_15459 ( P1_U5243 , P1_U5237 , P1_STATE2_REG_2_ );
nand NAND2_15460 ( P1_U5244 , P1_U5241 , P1_U3695 );
nand NAND2_15461 ( P1_U5245 , P1_U2511 , P1_U2388 );
nand NAND2_15462 ( P1_U5246 , P1_U3320 , P1_U5245 );
nand NAND2_15463 ( P1_U5247 , P1_U5246 , P1_U3375 );
nand NAND2_15464 ( P1_U5248 , P1_STATE2_REG_2_ , P1_U3376 );
nand NAND2_15465 ( P1_U5249 , P1_U5248 , P1_U5247 );
nand NAND2_15466 ( P1_U5250 , P1_U5233 , P1_U2415 );
nand NAND2_15467 ( P1_U5251 , P1_U2509 , P1_U2413 );
nand NAND2_15468 ( P1_U5252 , P1_U5232 , P1_U2412 );
nand NAND2_15469 ( P1_U5253 , P1_U2397 , P1_U5249 );
nand NAND2_15470 ( P1_U5254 , P1_INSTQUEUE_REG_3__7_ , P1_U5244 );
nand NAND2_15471 ( P1_U5255 , P1_U5233 , P1_U2416 );
nand NAND2_15472 ( P1_U5256 , P1_U2509 , P1_U2411 );
nand NAND2_15473 ( P1_U5257 , P1_U5232 , P1_U2410 );
nand NAND2_15474 ( P1_U5258 , P1_U2396 , P1_U5249 );
nand NAND2_15475 ( P1_U5259 , P1_INSTQUEUE_REG_3__6_ , P1_U5244 );
nand NAND2_15476 ( P1_U5260 , P1_U5233 , P1_U2420 );
nand NAND2_15477 ( P1_U5261 , P1_U2509 , P1_U2409 );
nand NAND2_15478 ( P1_U5262 , P1_U5232 , P1_U2408 );
nand NAND2_15479 ( P1_U5263 , P1_U2395 , P1_U5249 );
nand NAND2_15480 ( P1_U5264 , P1_INSTQUEUE_REG_3__5_ , P1_U5244 );
nand NAND2_15481 ( P1_U5265 , P1_U5233 , P1_U2419 );
nand NAND2_15482 ( P1_U5266 , P1_U2509 , P1_U2407 );
nand NAND2_15483 ( P1_U5267 , P1_U5232 , P1_U2406 );
nand NAND2_15484 ( P1_U5268 , P1_U2394 , P1_U5249 );
nand NAND2_15485 ( P1_U5269 , P1_INSTQUEUE_REG_3__4_ , P1_U5244 );
nand NAND2_15486 ( P1_U5270 , P1_U5233 , P1_U2418 );
nand NAND2_15487 ( P1_U5271 , P1_U2509 , P1_U2405 );
nand NAND2_15488 ( P1_U5272 , P1_U5232 , P1_U2404 );
nand NAND2_15489 ( P1_U5273 , P1_U2393 , P1_U5249 );
nand NAND2_15490 ( P1_U5274 , P1_INSTQUEUE_REG_3__3_ , P1_U5244 );
nand NAND2_15491 ( P1_U5275 , P1_U5233 , P1_U2421 );
nand NAND2_15492 ( P1_U5276 , P1_U2509 , P1_U2403 );
nand NAND2_15493 ( P1_U5277 , P1_U5232 , P1_U2402 );
nand NAND2_15494 ( P1_U5278 , P1_U2392 , P1_U5249 );
nand NAND2_15495 ( P1_U5279 , P1_INSTQUEUE_REG_3__2_ , P1_U5244 );
nand NAND2_15496 ( P1_U5280 , P1_U5233 , P1_U2414 );
nand NAND2_15497 ( P1_U5281 , P1_U2509 , P1_U2401 );
nand NAND2_15498 ( P1_U5282 , P1_U5232 , P1_U2400 );
nand NAND2_15499 ( P1_U5283 , P1_U2391 , P1_U5249 );
nand NAND2_15500 ( P1_U5284 , P1_INSTQUEUE_REG_3__1_ , P1_U5244 );
nand NAND2_15501 ( P1_U5285 , P1_U5233 , P1_U2417 );
nand NAND2_15502 ( P1_U5286 , P1_U2509 , P1_U2399 );
nand NAND2_15503 ( P1_U5287 , P1_U5232 , P1_U2398 );
nand NAND2_15504 ( P1_U5288 , P1_U2390 , P1_U5249 );
nand NAND2_15505 ( P1_U5289 , P1_INSTQUEUE_REG_3__0_ , P1_U5244 );
not NOT1_15506 ( P1_U5290 , P1_U3378 );
not NOT1_15507 ( P1_U5291 , P1_U3377 );
nand NAND2_15508 ( P1_U5292 , P1_U2441 , P1_U2443 );
not NOT1_15509 ( P1_U5293 , P1_U3379 );
not NOT1_15510 ( P1_U5294 , P1_U3242 );
nand NAND2_15511 ( P1_U5295 , P1_U2508 , P1_U4524 );
nand NAND2_15512 ( P1_U5296 , P1_U2513 , P1_U2358 );
nand NAND2_15513 ( P1_U5297 , P1_U3320 , P1_U5296 );
nand NAND2_15514 ( P1_U5298 , P1_U5293 , P1_U5297 );
nand NAND2_15515 ( P1_U5299 , P1_STATE2_REG_3_ , P1_U3377 );
nand NAND2_15516 ( P1_U5300 , P1_STATE2_REG_2_ , P1_U3242 );
nand NAND2_15517 ( P1_U5301 , P1_U5298 , P1_U3704 );
nand NAND2_15518 ( P1_U5302 , P1_U2513 , P1_U2388 );
nand NAND2_15519 ( P1_U5303 , P1_U3320 , P1_U5302 );
nand NAND2_15520 ( P1_U5304 , P1_U5303 , P1_U3379 );
nand NAND2_15521 ( P1_U5305 , P1_STATE2_REG_2_ , P1_U5294 );
nand NAND2_15522 ( P1_U5306 , P1_U5305 , P1_U5304 );
nand NAND2_15523 ( P1_U5307 , P1_U5291 , P1_U2415 );
nand NAND2_15524 ( P1_U5308 , P1_U2512 , P1_U2413 );
nand NAND2_15525 ( P1_U5309 , P1_U5290 , P1_U2412 );
nand NAND2_15526 ( P1_U5310 , P1_U2397 , P1_U5306 );
nand NAND2_15527 ( P1_U5311 , P1_INSTQUEUE_REG_2__7_ , P1_U5301 );
nand NAND2_15528 ( P1_U5312 , P1_U5291 , P1_U2416 );
nand NAND2_15529 ( P1_U5313 , P1_U2512 , P1_U2411 );
nand NAND2_15530 ( P1_U5314 , P1_U5290 , P1_U2410 );
nand NAND2_15531 ( P1_U5315 , P1_U2396 , P1_U5306 );
nand NAND2_15532 ( P1_U5316 , P1_INSTQUEUE_REG_2__6_ , P1_U5301 );
nand NAND2_15533 ( P1_U5317 , P1_U5291 , P1_U2420 );
nand NAND2_15534 ( P1_U5318 , P1_U2512 , P1_U2409 );
nand NAND2_15535 ( P1_U5319 , P1_U5290 , P1_U2408 );
nand NAND2_15536 ( P1_U5320 , P1_U2395 , P1_U5306 );
nand NAND2_15537 ( P1_U5321 , P1_INSTQUEUE_REG_2__5_ , P1_U5301 );
nand NAND2_15538 ( P1_U5322 , P1_U5291 , P1_U2419 );
nand NAND2_15539 ( P1_U5323 , P1_U2512 , P1_U2407 );
nand NAND2_15540 ( P1_U5324 , P1_U5290 , P1_U2406 );
nand NAND2_15541 ( P1_U5325 , P1_U2394 , P1_U5306 );
nand NAND2_15542 ( P1_U5326 , P1_INSTQUEUE_REG_2__4_ , P1_U5301 );
nand NAND2_15543 ( P1_U5327 , P1_U5291 , P1_U2418 );
nand NAND2_15544 ( P1_U5328 , P1_U2512 , P1_U2405 );
nand NAND2_15545 ( P1_U5329 , P1_U5290 , P1_U2404 );
nand NAND2_15546 ( P1_U5330 , P1_U2393 , P1_U5306 );
nand NAND2_15547 ( P1_U5331 , P1_INSTQUEUE_REG_2__3_ , P1_U5301 );
nand NAND2_15548 ( P1_U5332 , P1_U5291 , P1_U2421 );
nand NAND2_15549 ( P1_U5333 , P1_U2512 , P1_U2403 );
nand NAND2_15550 ( P1_U5334 , P1_U5290 , P1_U2402 );
nand NAND2_15551 ( P1_U5335 , P1_U2392 , P1_U5306 );
nand NAND2_15552 ( P1_U5336 , P1_INSTQUEUE_REG_2__2_ , P1_U5301 );
nand NAND2_15553 ( P1_U5337 , P1_U5291 , P1_U2414 );
nand NAND2_15554 ( P1_U5338 , P1_U2512 , P1_U2401 );
nand NAND2_15555 ( P1_U5339 , P1_U5290 , P1_U2400 );
nand NAND2_15556 ( P1_U5340 , P1_U2391 , P1_U5306 );
nand NAND2_15557 ( P1_U5341 , P1_INSTQUEUE_REG_2__1_ , P1_U5301 );
nand NAND2_15558 ( P1_U5342 , P1_U5291 , P1_U2417 );
nand NAND2_15559 ( P1_U5343 , P1_U2512 , P1_U2399 );
nand NAND2_15560 ( P1_U5344 , P1_U5290 , P1_U2398 );
nand NAND2_15561 ( P1_U5345 , P1_U2390 , P1_U5306 );
nand NAND2_15562 ( P1_U5346 , P1_INSTQUEUE_REG_2__0_ , P1_U5301 );
not NOT1_15563 ( P1_U5347 , P1_U3381 );
not NOT1_15564 ( P1_U5348 , P1_U3380 );
nand NAND2_15565 ( P1_U5349 , P1_U2441 , P1_U2444 );
not NOT1_15566 ( P1_U5350 , P1_U3382 );
nand NAND2_15567 ( P1_U5351 , P1_U2435 , P1_U2437 );
not NOT1_15568 ( P1_U5352 , P1_U3383 );
nand NAND2_15569 ( P1_U5353 , P1_U2508 , P1_U4525 );
nand NAND2_15570 ( P1_U5354 , P1_U2515 , P1_U2358 );
nand NAND2_15571 ( P1_U5355 , P1_U3320 , P1_U5354 );
nand NAND2_15572 ( P1_U5356 , P1_U5350 , P1_U5355 );
nand NAND2_15573 ( P1_U5357 , P1_STATE2_REG_3_ , P1_U3380 );
nand NAND2_15574 ( P1_U5358 , P1_U5352 , P1_STATE2_REG_2_ );
nand NAND2_15575 ( P1_U5359 , P1_U5356 , P1_U3713 );
nand NAND2_15576 ( P1_U5360 , P1_U2515 , P1_U2388 );
nand NAND2_15577 ( P1_U5361 , P1_U3320 , P1_U5360 );
nand NAND2_15578 ( P1_U5362 , P1_U5361 , P1_U3382 );
nand NAND2_15579 ( P1_U5363 , P1_STATE2_REG_2_ , P1_U3383 );
nand NAND2_15580 ( P1_U5364 , P1_U5363 , P1_U5362 );
nand NAND2_15581 ( P1_U5365 , P1_U5348 , P1_U2415 );
nand NAND2_15582 ( P1_U5366 , P1_U2514 , P1_U2413 );
nand NAND2_15583 ( P1_U5367 , P1_U5347 , P1_U2412 );
nand NAND2_15584 ( P1_U5368 , P1_U2397 , P1_U5364 );
nand NAND2_15585 ( P1_U5369 , P1_INSTQUEUE_REG_1__7_ , P1_U5359 );
nand NAND2_15586 ( P1_U5370 , P1_U5348 , P1_U2416 );
nand NAND2_15587 ( P1_U5371 , P1_U2514 , P1_U2411 );
nand NAND2_15588 ( P1_U5372 , P1_U5347 , P1_U2410 );
nand NAND2_15589 ( P1_U5373 , P1_U2396 , P1_U5364 );
nand NAND2_15590 ( P1_U5374 , P1_INSTQUEUE_REG_1__6_ , P1_U5359 );
nand NAND2_15591 ( P1_U5375 , P1_U5348 , P1_U2420 );
nand NAND2_15592 ( P1_U5376 , P1_U2514 , P1_U2409 );
nand NAND2_15593 ( P1_U5377 , P1_U5347 , P1_U2408 );
nand NAND2_15594 ( P1_U5378 , P1_U2395 , P1_U5364 );
nand NAND2_15595 ( P1_U5379 , P1_INSTQUEUE_REG_1__5_ , P1_U5359 );
nand NAND2_15596 ( P1_U5380 , P1_U5348 , P1_U2419 );
nand NAND2_15597 ( P1_U5381 , P1_U2514 , P1_U2407 );
nand NAND2_15598 ( P1_U5382 , P1_U5347 , P1_U2406 );
nand NAND2_15599 ( P1_U5383 , P1_U2394 , P1_U5364 );
nand NAND2_15600 ( P1_U5384 , P1_INSTQUEUE_REG_1__4_ , P1_U5359 );
nand NAND2_15601 ( P1_U5385 , P1_U5348 , P1_U2418 );
nand NAND2_15602 ( P1_U5386 , P1_U2514 , P1_U2405 );
nand NAND2_15603 ( P1_U5387 , P1_U5347 , P1_U2404 );
nand NAND2_15604 ( P1_U5388 , P1_U2393 , P1_U5364 );
nand NAND2_15605 ( P1_U5389 , P1_INSTQUEUE_REG_1__3_ , P1_U5359 );
nand NAND2_15606 ( P1_U5390 , P1_U5348 , P1_U2421 );
nand NAND2_15607 ( P1_U5391 , P1_U2514 , P1_U2403 );
nand NAND2_15608 ( P1_U5392 , P1_U5347 , P1_U2402 );
nand NAND2_15609 ( P1_U5393 , P1_U2392 , P1_U5364 );
nand NAND2_15610 ( P1_U5394 , P1_INSTQUEUE_REG_1__2_ , P1_U5359 );
nand NAND2_15611 ( P1_U5395 , P1_U5348 , P1_U2414 );
nand NAND2_15612 ( P1_U5396 , P1_U2514 , P1_U2401 );
nand NAND2_15613 ( P1_U5397 , P1_U5347 , P1_U2400 );
nand NAND2_15614 ( P1_U5398 , P1_U2391 , P1_U5364 );
nand NAND2_15615 ( P1_U5399 , P1_INSTQUEUE_REG_1__1_ , P1_U5359 );
nand NAND2_15616 ( P1_U5400 , P1_U5348 , P1_U2417 );
nand NAND2_15617 ( P1_U5401 , P1_U2514 , P1_U2399 );
nand NAND2_15618 ( P1_U5402 , P1_U5347 , P1_U2398 );
nand NAND2_15619 ( P1_U5403 , P1_U2390 , P1_U5364 );
nand NAND2_15620 ( P1_U5404 , P1_INSTQUEUE_REG_1__0_ , P1_U5359 );
not NOT1_15621 ( P1_U5405 , P1_U3385 );
not NOT1_15622 ( P1_U5406 , P1_U3384 );
nand NAND2_15623 ( P1_U5407 , P1_U2441 , P1_U2445 );
not NOT1_15624 ( P1_U5408 , P1_U3386 );
not NOT1_15625 ( P1_U5409 , P1_U3243 );
nand NAND2_15626 ( P1_U5410 , P1_U2508 , P1_U2486 );
nand NAND2_15627 ( P1_U5411 , P1_U2517 , P1_U2358 );
nand NAND2_15628 ( P1_U5412 , P1_U3320 , P1_U5411 );
nand NAND2_15629 ( P1_U5413 , P1_U5408 , P1_U5412 );
nand NAND2_15630 ( P1_U5414 , P1_STATE2_REG_3_ , P1_U3384 );
nand NAND2_15631 ( P1_U5415 , P1_STATE2_REG_2_ , P1_U3243 );
nand NAND2_15632 ( P1_U5416 , P1_U5413 , P1_U3722 );
nand NAND2_15633 ( P1_U5417 , P1_U2517 , P1_U2388 );
nand NAND2_15634 ( P1_U5418 , P1_U3320 , P1_U5417 );
nand NAND2_15635 ( P1_U5419 , P1_U5418 , P1_U3386 );
nand NAND2_15636 ( P1_U5420 , P1_STATE2_REG_2_ , P1_U5409 );
nand NAND2_15637 ( P1_U5421 , P1_U5420 , P1_U5419 );
nand NAND2_15638 ( P1_U5422 , P1_U5406 , P1_U2415 );
nand NAND2_15639 ( P1_U5423 , P1_U2516 , P1_U2413 );
nand NAND2_15640 ( P1_U5424 , P1_U5405 , P1_U2412 );
nand NAND2_15641 ( P1_U5425 , P1_U2397 , P1_U5421 );
nand NAND2_15642 ( P1_U5426 , P1_INSTQUEUE_REG_0__7_ , P1_U5416 );
nand NAND2_15643 ( P1_U5427 , P1_U5406 , P1_U2416 );
nand NAND2_15644 ( P1_U5428 , P1_U2516 , P1_U2411 );
nand NAND2_15645 ( P1_U5429 , P1_U5405 , P1_U2410 );
nand NAND2_15646 ( P1_U5430 , P1_U2396 , P1_U5421 );
nand NAND2_15647 ( P1_U5431 , P1_INSTQUEUE_REG_0__6_ , P1_U5416 );
nand NAND2_15648 ( P1_U5432 , P1_U5406 , P1_U2420 );
nand NAND2_15649 ( P1_U5433 , P1_U2516 , P1_U2409 );
nand NAND2_15650 ( P1_U5434 , P1_U5405 , P1_U2408 );
nand NAND2_15651 ( P1_U5435 , P1_U2395 , P1_U5421 );
nand NAND2_15652 ( P1_U5436 , P1_INSTQUEUE_REG_0__5_ , P1_U5416 );
nand NAND2_15653 ( P1_U5437 , P1_U5406 , P1_U2419 );
nand NAND2_15654 ( P1_U5438 , P1_U2516 , P1_U2407 );
nand NAND2_15655 ( P1_U5439 , P1_U5405 , P1_U2406 );
nand NAND2_15656 ( P1_U5440 , P1_U2394 , P1_U5421 );
nand NAND2_15657 ( P1_U5441 , P1_U5406 , P1_U2418 );
nand NAND2_15658 ( P1_U5442 , P1_U2516 , P1_U2405 );
nand NAND2_15659 ( P1_U5443 , P1_U5405 , P1_U2404 );
nand NAND2_15660 ( P1_U5444 , P1_U2393 , P1_U5421 );
nand NAND2_15661 ( P1_U5445 , P1_INSTQUEUE_REG_0__3_ , P1_U5416 );
nand NAND2_15662 ( P1_U5446 , P1_U5406 , P1_U2421 );
nand NAND2_15663 ( P1_U5447 , P1_U2516 , P1_U2403 );
nand NAND2_15664 ( P1_U5448 , P1_U5405 , P1_U2402 );
nand NAND2_15665 ( P1_U5449 , P1_U2392 , P1_U5421 );
nand NAND2_15666 ( P1_U5450 , P1_INSTQUEUE_REG_0__2_ , P1_U5416 );
nand NAND2_15667 ( P1_U5451 , P1_U5406 , P1_U2414 );
nand NAND2_15668 ( P1_U5452 , P1_U2516 , P1_U2401 );
nand NAND2_15669 ( P1_U5453 , P1_U5405 , P1_U2400 );
nand NAND2_15670 ( P1_U5454 , P1_U2391 , P1_U5421 );
nand NAND2_15671 ( P1_U5455 , P1_INSTQUEUE_REG_0__1_ , P1_U5416 );
nand NAND2_15672 ( P1_U5456 , P1_U5406 , P1_U2417 );
nand NAND2_15673 ( P1_U5457 , P1_U2516 , P1_U2399 );
nand NAND2_15674 ( P1_U5458 , P1_U5405 , P1_U2398 );
nand NAND2_15675 ( P1_U5459 , P1_U2390 , P1_U5421 );
nand NAND2_15676 ( P1_U5460 , P1_INSTQUEUE_REG_0__0_ , P1_U5416 );
not NOT1_15677 ( P1_U5461 , P1_U3423 );
nand NAND3_15678 ( P1_U5462 , P1_U3391 , P1_U3394 , P1_U4503 );
nand NAND3_15679 ( P1_U5463 , P1_U4400 , P1_U4173 , P1_U4460 );
not NOT1_15680 ( P1_U5464 , P1_U3244 );
nand NAND2_15681 ( P1_U5465 , P1_U4494 , P1_U3289 );
nand NAND3_15682 ( P1_U5466 , P1_U5465 , P1_U3283 , P1_U5464 );
nand NAND2_15683 ( P1_U5467 , P1_U3732 , P1_U2452 );
nand NAND2_15684 ( P1_U5468 , P1_U4208 , P1_U5462 );
nand NAND2_15685 ( P1_U5469 , P1_U3733 , P1_U7609 );
nand NAND3_15686 ( P1_U5470 , P1_U4215 , P1_U3257 , P1_GTE_485_U6 );
nand NAND2_15687 ( P1_U5471 , P1_U2449 , P1_U7494 );
nand NAND2_15688 ( P1_U5472 , P1_U4257 , P1_U4503 );
not NOT1_15689 ( P1_U5473 , P1_U4182 );
nand NAND2_15690 ( P1_U5474 , P1_U2368 , P1_U4182 );
nand NAND2_15691 ( P1_U5475 , P1_STATE2_REG_3_ , P1_U3294 );
not NOT1_15692 ( P1_U5476 , P1_U4172 );
nand NAND2_15693 ( P1_U5477 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_15694 ( P1_U5478 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_U5477 );
nand NAND2_15695 ( P1_U5479 , P1_U4381 , P1_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_15696 ( P1_U5480 , P1_U3442 );
nand NAND2_15697 ( P1_U5481 , P1_U3498 , P1_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_15698 ( P1_U5482 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_U5481 );
not NOT1_15699 ( P1_U5483 , P1_U3438 );
nand NAND2_15700 ( P1_U5484 , P1_U3275 , P1_U3264 );
nand NAND2_15701 ( P1_U5485 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_U5484 );
nand NAND2_15702 ( P1_U5486 , P1_U2469 , P1_U3275 );
nand NAND2_15703 ( P1_U5487 , P1_U4494 , P1_U3290 );
nand NAND2_15704 ( P1_U5488 , P1_U4400 , P1_U2605 );
nand NAND3_15705 ( P1_U5489 , P1_U7704 , P1_U7703 , P1_U7494 );
nand NAND2_15706 ( P1_U5490 , P1_U4449 , P1_U5488 );
nand NAND3_15707 ( P1_U5491 , P1_U4400 , P1_U3394 , P1_U3409 );
nand NAND2_15708 ( P1_U5492 , P1_U5491 , P1_U4171 );
nand NAND2_15709 ( P1_U5493 , P1_U7629 , P1_U5492 );
nand NAND2_15710 ( P1_U5494 , P1_U4460 , P1_U4171 );
nand NAND2_15711 ( P1_U5495 , P1_U3395 , P1_U5494 );
nand NAND2_15712 ( P1_U5496 , P1_U4208 , P1_U5462 );
nand NAND2_15713 ( P1_U5497 , P1_U4257 , P1_U4503 );
nand NAND2_15714 ( P1_U5498 , P1_U5495 , P1_U3271 );
nand NAND2_15715 ( P1_U5499 , P1_U4494 , P1_U7707 );
nand NAND2_15716 ( P1_U5500 , P1_U4190 , P1_U3244 );
nand NAND2_15717 ( P1_U5501 , P1_U3292 , P1_U4217 );
nand NAND2_15718 ( P1_U5502 , P1_U3740 , P1_U5501 );
nand NAND2_15719 ( P1_U5503 , P1_R2182_U25 , P1_U7509 );
nand NAND2_15720 ( P1_U5504 , P1_U4218 , P1_U3438 );
nand NAND2_15721 ( P1_U5505 , P1_U4214 , P1_U3442 );
nand NAND2_15722 ( P1_U5506 , P1_U5503 , P1_U3747 );
nand NAND2_15723 ( P1_U5507 , P1_U4252 , P1_U3438 );
nand NAND2_15724 ( P1_U5508 , P1_U2427 , P1_U5506 );
nand NAND2_15725 ( P1_U5509 , P1_U5508 , P1_U5507 );
nand NAND2_15726 ( P1_U5510 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3275 );
not NOT1_15727 ( P1_U5511 , P1_U3401 );
nand NAND2_15728 ( P1_U5512 , P1_R2182_U42 , P1_U7509 );
nand NAND2_15729 ( P1_U5513 , P1_U4214 , P1_U3456 );
nand NAND2_15730 ( P1_U5514 , P1_U3749 , P1_U5512 );
nand NAND2_15731 ( P1_U5515 , P1_U2446 , P1_U3470 );
nand NAND2_15732 ( P1_U5516 , P1_U4252 , P1_U3401 );
nand NAND2_15733 ( P1_U5517 , P1_U2427 , P1_U5514 );
nand NAND3_15734 ( P1_U5518 , P1_U5517 , P1_U5515 , P1_U5516 );
not NOT1_15735 ( P1_U5519 , P1_U3402 );
nand NAND2_15736 ( P1_U5520 , P1_U2431 , P1_U4249 );
nand NAND2_15737 ( P1_U5521 , P1_U3292 , P1_U5520 );
nand NAND2_15738 ( P1_U5522 , P1_U5519 , P1_U5521 );
nand NAND2_15739 ( P1_U5523 , P1_R2182_U33 , P1_U7509 );
nand NAND2_15740 ( P1_U5524 , P1_U4214 , P1_U3265 );
nand NAND2_15741 ( P1_U5525 , P1_U3750 , P1_U5523 );
nand NAND2_15742 ( P1_U5526 , P1_U7712 , P1_U2446 );
nand NAND2_15743 ( P1_U5527 , P1_U5519 , P1_U4252 );
nand NAND2_15744 ( P1_U5528 , P1_U2427 , P1_U5525 );
nand NAND3_15745 ( P1_U5529 , P1_U5528 , P1_U5526 , P1_U5527 );
nand NAND2_15746 ( P1_U5530 , P1_R2182_U34 , P1_U7509 );
nand NAND2_15747 ( P1_U5531 , P1_U4175 , P1_U5530 );
nand NAND2_15748 ( P1_U5532 , P1_U4252 , P1_U3266 );
nand NAND2_15749 ( P1_U5533 , P1_U2427 , P1_U5531 );
nand NAND2_15750 ( P1_U5534 , P1_U7715 , P1_STATE2_REG_1_ );
nand NAND3_15751 ( P1_U5535 , P1_U5533 , P1_U5534 , P1_U5532 );
nand NAND3_15752 ( P1_U5536 , P1_U2428 , P1_STATE2_REG_0_ , P1_LT_589_U6 );
not NOT1_15753 ( P1_U5537 , P1_U3404 );
nand NAND2_15754 ( P1_U5538 , P1_STATE2_REG_1_ , P1_U3296 );
nand NAND2_15755 ( P1_U5539 , P1_U4527 , P1_U3454 );
nand NAND2_15756 ( P1_U5540 , P1_U3358 , P1_U5539 );
nand NAND2_15757 ( P1_U5541 , P1_U3359 , P1_U5540 );
nand NAND2_15758 ( P1_U5542 , P1_U2388 , P1_U5541 );
nand NAND2_15759 ( P1_U5543 , P1_R2182_U25 , P1_U5538 );
nand NAND2_15760 ( P1_U5544 , P1_U4226 , P1_R2144_U8 );
nand NAND2_15761 ( P1_U5545 , P1_U3751 , P1_U5542 );
nand NAND2_15762 ( P1_U5546 , P1_U2388 , P1_U7733 );
nand NAND2_15763 ( P1_U5547 , P1_R2182_U42 , P1_U5538 );
nand NAND2_15764 ( P1_U5548 , P1_U4226 , P1_R2144_U49 );
nand NAND2_15765 ( P1_U5549 , P1_U3752 , P1_U5546 );
nand NAND2_15766 ( P1_U5550 , P1_U3326 , P1_U3333 );
nand NAND2_15767 ( P1_U5551 , P1_U2388 , P1_U5550 );
nand NAND2_15768 ( P1_U5552 , P1_R2182_U33 , P1_U5538 );
nand NAND2_15769 ( P1_U5553 , P1_U4226 , P1_R2144_U50 );
nand NAND2_15770 ( P1_U5554 , P1_U3753 , P1_U5551 );
nand NAND2_15771 ( P1_U5555 , P1_R2182_U34 , P1_U5538 );
nand NAND2_15772 ( P1_U5556 , P1_R2144_U43 , P1_U4209 );
nand NAND3_15773 ( P1_U5557 , P1_U5555 , P1_U5556 , P1_U4245 );
nand NAND2_15774 ( P1_U5558 , P1_U4477 , P1_U3272 );
nand NAND2_15775 ( P1_U5559 , P1_U4260 , P1_U2431 );
nand NAND4_15776 ( P1_U5560 , P1_U2518 , P1_U5559 , P1_U7743 , P1_U7742 );
nand NAND3_15777 ( P1_U5561 , P1_U4235 , P1_U4503 , P1_U4192 );
nand NAND2_15778 ( P1_U5562 , P1_U2368 , P1_U5560 );
nand NAND2_15779 ( P1_U5563 , P1_U4203 , P1_U3263 );
not NOT1_15780 ( P1_U5564 , P1_U3414 );
nand NAND2_15781 ( P1_U5565 , P1_U4262 , P1_U4208 );
nand NAND2_15782 ( P1_U5566 , P1_U4256 , P1_U2389 );
nand NAND2_15783 ( P1_U5567 , P1_U4266 , P1_U4250 );
nand NAND2_15784 ( P1_U5568 , P1_U4264 , P1_U4494 );
nand NAND2_15785 ( P1_U5569 , P1_U3758 , P1_U2519 );
nand NAND2_15786 ( P1_U5570 , P1_R2099_U86 , P1_U2380 );
nand NAND2_15787 ( P1_U5571 , P1_R2027_U5 , P1_U2378 );
nand NAND2_15788 ( P1_U5572 , P1_R2278_U99 , P1_U2377 );
nand NAND2_15789 ( P1_U5573 , P1_ADD_405_U4 , P1_U2375 );
nand NAND2_15790 ( P1_U5574 , P1_INSTADDRPOINTER_REG_0_ , P1_U2374 );
nand NAND2_15791 ( P1_U5575 , P1_REIP_REG_0_ , P1_U2370 );
nand NAND2_15792 ( P1_U5576 , P1_U5564 , P1_INSTADDRPOINTER_REG_0_ );
nand NAND2_15793 ( P1_U5577 , P1_R2099_U87 , P1_U2380 );
nand NAND2_15794 ( P1_U5578 , P1_R2027_U71 , P1_U2378 );
nand NAND2_15795 ( P1_U5579 , P1_R2278_U19 , P1_U2377 );
nand NAND2_15796 ( P1_U5580 , P1_ADD_405_U85 , P1_U2375 );
nand NAND2_15797 ( P1_U5581 , P1_ADD_515_U4 , P1_U2374 );
nand NAND2_15798 ( P1_U5582 , P1_U2370 , P1_REIP_REG_1_ );
nand NAND2_15799 ( P1_U5583 , P1_U5564 , P1_INSTADDRPOINTER_REG_1_ );
nand NAND2_15800 ( P1_U5584 , P1_R2099_U138 , P1_U2380 );
nand NAND2_15801 ( P1_U5585 , P1_R2027_U60 , P1_U2378 );
nand NAND2_15802 ( P1_U5586 , P1_R2278_U107 , P1_U2377 );
nand NAND2_15803 ( P1_U5587 , P1_ADD_405_U5 , P1_U2375 );
nand NAND2_15804 ( P1_U5588 , P1_ADD_515_U67 , P1_U2374 );
nand NAND2_15805 ( P1_U5589 , P1_U2370 , P1_REIP_REG_2_ );
nand NAND2_15806 ( P1_U5590 , P1_INSTADDRPOINTER_REG_2_ , P1_U5564 );
nand NAND2_15807 ( P1_U5591 , P1_R2099_U42 , P1_U2380 );
nand NAND2_15808 ( P1_U5592 , P1_R2027_U57 , P1_U2378 );
nand NAND2_15809 ( P1_U5593 , P1_R2278_U105 , P1_U2377 );
nand NAND2_15810 ( P1_U5594 , P1_ADD_405_U95 , P1_U2375 );
nand NAND2_15811 ( P1_U5595 , P1_ADD_515_U85 , P1_U2374 );
nand NAND2_15812 ( P1_U5596 , P1_U2370 , P1_REIP_REG_3_ );
nand NAND2_15813 ( P1_U5597 , P1_INSTADDRPOINTER_REG_3_ , P1_U5564 );
nand NAND2_15814 ( P1_U5598 , P1_R2099_U41 , P1_U2380 );
nand NAND2_15815 ( P1_U5599 , P1_R2027_U56 , P1_U2378 );
nand NAND2_15816 ( P1_U5600 , P1_R2278_U104 , P1_U2377 );
nand NAND2_15817 ( P1_U5601 , P1_ADD_405_U76 , P1_U2375 );
nand NAND2_15818 ( P1_U5602 , P1_ADD_515_U76 , P1_U2374 );
nand NAND2_15819 ( P1_U5603 , P1_U2370 , P1_REIP_REG_4_ );
nand NAND2_15820 ( P1_U5604 , P1_INSTADDRPOINTER_REG_4_ , P1_U5564 );
nand NAND2_15821 ( P1_U5605 , P1_R2099_U40 , P1_U2380 );
nand NAND2_15822 ( P1_U5606 , P1_R2027_U55 , P1_U2378 );
nand NAND2_15823 ( P1_U5607 , P1_R2278_U17 , P1_U2377 );
nand NAND2_15824 ( P1_U5608 , P1_ADD_405_U79 , P1_U2375 );
nand NAND2_15825 ( P1_U5609 , P1_ADD_515_U79 , P1_U2374 );
nand NAND2_15826 ( P1_U5610 , P1_U2370 , P1_REIP_REG_5_ );
nand NAND2_15827 ( P1_U5611 , P1_INSTADDRPOINTER_REG_5_ , P1_U5564 );
nand NAND2_15828 ( P1_U5612 , P1_R2099_U39 , P1_U2380 );
nand NAND2_15829 ( P1_U5613 , P1_R2027_U54 , P1_U2378 );
nand NAND2_15830 ( P1_U5614 , P1_R2278_U103 , P1_U2377 );
nand NAND2_15831 ( P1_U5615 , P1_ADD_405_U63 , P1_U2375 );
nand NAND2_15832 ( P1_U5616 , P1_ADD_515_U62 , P1_U2374 );
nand NAND2_15833 ( P1_U5617 , P1_U2370 , P1_REIP_REG_6_ );
nand NAND2_15834 ( P1_U5618 , P1_INSTADDRPOINTER_REG_6_ , P1_U5564 );
nand NAND2_15835 ( P1_U5619 , P1_R2099_U38 , P1_U2380 );
nand NAND2_15836 ( P1_U5620 , P1_R2027_U53 , P1_U2378 );
nand NAND2_15837 ( P1_U5621 , P1_R2278_U18 , P1_U2377 );
nand NAND2_15838 ( P1_U5622 , P1_ADD_405_U89 , P1_U2375 );
nand NAND2_15839 ( P1_U5623 , P1_ADD_515_U89 , P1_U2374 );
nand NAND2_15840 ( P1_U5624 , P1_U2370 , P1_REIP_REG_7_ );
nand NAND2_15841 ( P1_U5625 , P1_INSTADDRPOINTER_REG_7_ , P1_U5564 );
nand NAND2_15842 ( P1_U5626 , P1_R2099_U37 , P1_U2380 );
nand NAND2_15843 ( P1_U5627 , P1_R2027_U52 , P1_U2378 );
nand NAND2_15844 ( P1_U5628 , P1_R2278_U102 , P1_U2377 );
nand NAND2_15845 ( P1_U5629 , P1_ADD_405_U80 , P1_U2375 );
nand NAND2_15846 ( P1_U5630 , P1_ADD_515_U80 , P1_U2374 );
nand NAND2_15847 ( P1_U5631 , P1_U2370 , P1_REIP_REG_8_ );
nand NAND2_15848 ( P1_U5632 , P1_INSTADDRPOINTER_REG_8_ , P1_U5564 );
nand NAND2_15849 ( P1_U5633 , P1_R2099_U36 , P1_U2380 );
nand NAND2_15850 ( P1_U5634 , P1_R2027_U51 , P1_U2378 );
nand NAND2_15851 ( P1_U5635 , P1_R2278_U101 , P1_U2377 );
nand NAND2_15852 ( P1_U5636 , P1_ADD_405_U70 , P1_U2375 );
nand NAND2_15853 ( P1_U5637 , P1_ADD_515_U70 , P1_U2374 );
nand NAND2_15854 ( P1_U5638 , P1_U2370 , P1_REIP_REG_9_ );
nand NAND2_15855 ( P1_U5639 , P1_INSTADDRPOINTER_REG_9_ , P1_U5564 );
nand NAND2_15856 ( P1_U5640 , P1_R2099_U85 , P1_U2380 );
nand NAND2_15857 ( P1_U5641 , P1_R2027_U81 , P1_U2378 );
nand NAND2_15858 ( P1_U5642 , P1_R2278_U126 , P1_U2377 );
nand NAND2_15859 ( P1_U5643 , P1_ADD_405_U83 , P1_U2375 );
nand NAND2_15860 ( P1_U5644 , P1_ADD_515_U83 , P1_U2374 );
nand NAND2_15861 ( P1_U5645 , P1_U2370 , P1_REIP_REG_10_ );
nand NAND2_15862 ( P1_U5646 , P1_INSTADDRPOINTER_REG_10_ , P1_U5564 );
nand NAND2_15863 ( P1_U5647 , P1_R2099_U84 , P1_U2380 );
nand NAND2_15864 ( P1_U5648 , P1_R2027_U80 , P1_U2378 );
nand NAND2_15865 ( P1_U5649 , P1_R2278_U15 , P1_U2377 );
nand NAND2_15866 ( P1_U5650 , P1_ADD_405_U73 , P1_U2375 );
nand NAND2_15867 ( P1_U5651 , P1_ADD_515_U73 , P1_U2374 );
nand NAND2_15868 ( P1_U5652 , P1_U2370 , P1_REIP_REG_11_ );
nand NAND2_15869 ( P1_U5653 , P1_INSTADDRPOINTER_REG_11_ , P1_U5564 );
nand NAND2_15870 ( P1_U5654 , P1_R2099_U83 , P1_U2380 );
nand NAND2_15871 ( P1_U5655 , P1_R2027_U79 , P1_U2378 );
nand NAND2_15872 ( P1_U5656 , P1_R2278_U125 , P1_U2377 );
nand NAND2_15873 ( P1_U5657 , P1_ADD_405_U88 , P1_U2375 );
nand NAND2_15874 ( P1_U5658 , P1_ADD_515_U88 , P1_U2374 );
nand NAND2_15875 ( P1_U5659 , P1_U2370 , P1_REIP_REG_12_ );
nand NAND2_15876 ( P1_U5660 , P1_INSTADDRPOINTER_REG_12_ , P1_U5564 );
nand NAND2_15877 ( P1_U5661 , P1_R2099_U82 , P1_U2380 );
nand NAND2_15878 ( P1_U5662 , P1_R2027_U78 , P1_U2378 );
nand NAND2_15879 ( P1_U5663 , P1_R2278_U123 , P1_U2377 );
nand NAND2_15880 ( P1_U5664 , P1_ADD_405_U69 , P1_U2375 );
nand NAND2_15881 ( P1_U5665 , P1_ADD_515_U69 , P1_U2374 );
nand NAND2_15882 ( P1_U5666 , P1_U2370 , P1_REIP_REG_13_ );
nand NAND2_15883 ( P1_U5667 , P1_INSTADDRPOINTER_REG_13_ , P1_U5564 );
nand NAND2_15884 ( P1_U5668 , P1_R2099_U81 , P1_U2380 );
nand NAND2_15885 ( P1_U5669 , P1_R2027_U77 , P1_U2378 );
nand NAND2_15886 ( P1_U5670 , P1_R2278_U122 , P1_U2377 );
nand NAND2_15887 ( P1_U5671 , P1_ADD_405_U78 , P1_U2375 );
nand NAND2_15888 ( P1_U5672 , P1_ADD_515_U78 , P1_U2374 );
nand NAND2_15889 ( P1_U5673 , P1_U2370 , P1_REIP_REG_14_ );
nand NAND2_15890 ( P1_U5674 , P1_INSTADDRPOINTER_REG_14_ , P1_U5564 );
nand NAND2_15891 ( P1_U5675 , P1_R2099_U80 , P1_U2380 );
nand NAND2_15892 ( P1_U5676 , P1_R2027_U76 , P1_U2378 );
nand NAND2_15893 ( P1_U5677 , P1_R2278_U20 , P1_U2377 );
nand NAND2_15894 ( P1_U5678 , P1_ADD_405_U75 , P1_U2375 );
nand NAND2_15895 ( P1_U5679 , P1_ADD_515_U75 , P1_U2374 );
nand NAND2_15896 ( P1_U5680 , P1_U2370 , P1_REIP_REG_15_ );
nand NAND2_15897 ( P1_U5681 , P1_INSTADDRPOINTER_REG_15_ , P1_U5564 );
nand NAND2_15898 ( P1_U5682 , P1_R2099_U79 , P1_U2380 );
nand NAND2_15899 ( P1_U5683 , P1_R2027_U75 , P1_U2378 );
nand NAND2_15900 ( P1_U5684 , P1_R2278_U121 , P1_U2377 );
nand NAND2_15901 ( P1_U5685 , P1_ADD_405_U91 , P1_U2375 );
nand NAND2_15902 ( P1_U5686 , P1_ADD_515_U91 , P1_U2374 );
nand NAND2_15903 ( P1_U5687 , P1_U2370 , P1_REIP_REG_16_ );
nand NAND2_15904 ( P1_U5688 , P1_INSTADDRPOINTER_REG_16_ , P1_U5564 );
nand NAND2_15905 ( P1_U5689 , P1_R2099_U78 , P1_U2380 );
nand NAND2_15906 ( P1_U5690 , P1_R2027_U74 , P1_U2378 );
nand NAND2_15907 ( P1_U5691 , P1_R2278_U120 , P1_U2377 );
nand NAND2_15908 ( P1_U5692 , P1_ADD_405_U67 , P1_U2375 );
nand NAND2_15909 ( P1_U5693 , P1_ADD_515_U66 , P1_U2374 );
nand NAND2_15910 ( P1_U5694 , P1_U2370 , P1_REIP_REG_17_ );
nand NAND2_15911 ( P1_U5695 , P1_INSTADDRPOINTER_REG_17_ , P1_U5564 );
nand NAND2_15912 ( P1_U5696 , P1_R2099_U77 , P1_U2380 );
nand NAND2_15913 ( P1_U5697 , P1_R2027_U73 , P1_U2378 );
nand NAND2_15914 ( P1_U5698 , P1_R2278_U119 , P1_U2377 );
nand NAND2_15915 ( P1_U5699 , P1_ADD_405_U72 , P1_U2375 );
nand NAND2_15916 ( P1_U5700 , P1_ADD_515_U72 , P1_U2374 );
nand NAND2_15917 ( P1_U5701 , P1_U2370 , P1_REIP_REG_18_ );
nand NAND2_15918 ( P1_U5702 , P1_INSTADDRPOINTER_REG_18_ , P1_U5564 );
nand NAND2_15919 ( P1_U5703 , P1_R2099_U76 , P1_U2380 );
nand NAND2_15920 ( P1_U5704 , P1_R2027_U72 , P1_U2378 );
nand NAND2_15921 ( P1_U5705 , P1_R2278_U118 , P1_U2377 );
nand NAND2_15922 ( P1_U5706 , P1_ADD_405_U82 , P1_U2375 );
nand NAND2_15923 ( P1_U5707 , P1_ADD_515_U82 , P1_U2374 );
nand NAND2_15924 ( P1_U5708 , P1_U2370 , P1_REIP_REG_19_ );
nand NAND2_15925 ( P1_U5709 , P1_INSTADDRPOINTER_REG_19_ , P1_U5564 );
nand NAND2_15926 ( P1_U5710 , P1_R2099_U75 , P1_U2380 );
nand NAND2_15927 ( P1_U5711 , P1_R2027_U70 , P1_U2378 );
nand NAND2_15928 ( P1_U5712 , P1_R2278_U117 , P1_U2377 );
nand NAND2_15929 ( P1_U5713 , P1_ADD_405_U68 , P1_U2375 );
nand NAND2_15930 ( P1_U5714 , P1_ADD_515_U68 , P1_U2374 );
nand NAND2_15931 ( P1_U5715 , P1_U2370 , P1_REIP_REG_20_ );
nand NAND2_15932 ( P1_U5716 , P1_INSTADDRPOINTER_REG_20_ , P1_U5564 );
nand NAND2_15933 ( P1_U5717 , P1_R2099_U74 , P1_U2380 );
nand NAND2_15934 ( P1_U5718 , P1_R2027_U69 , P1_U2378 );
nand NAND2_15935 ( P1_U5719 , P1_R2278_U116 , P1_U2377 );
nand NAND2_15936 ( P1_U5720 , P1_ADD_405_U87 , P1_U2375 );
nand NAND2_15937 ( P1_U5721 , P1_ADD_515_U87 , P1_U2374 );
nand NAND2_15938 ( P1_U5722 , P1_U2370 , P1_REIP_REG_21_ );
nand NAND2_15939 ( P1_U5723 , P1_INSTADDRPOINTER_REG_21_ , P1_U5564 );
nand NAND2_15940 ( P1_U5724 , P1_R2099_U73 , P1_U2380 );
nand NAND2_15941 ( P1_U5725 , P1_R2027_U68 , P1_U2378 );
nand NAND2_15942 ( P1_U5726 , P1_R2278_U115 , P1_U2377 );
nand NAND2_15943 ( P1_U5727 , P1_ADD_405_U71 , P1_U2375 );
nand NAND2_15944 ( P1_U5728 , P1_ADD_515_U71 , P1_U2374 );
nand NAND2_15945 ( P1_U5729 , P1_U2370 , P1_REIP_REG_22_ );
nand NAND2_15946 ( P1_U5730 , P1_INSTADDRPOINTER_REG_22_ , P1_U5564 );
nand NAND2_15947 ( P1_U5731 , P1_R2099_U72 , P1_U2380 );
nand NAND2_15948 ( P1_U5732 , P1_R2027_U67 , P1_U2378 );
nand NAND2_15949 ( P1_U5733 , P1_R2278_U114 , P1_U2377 );
nand NAND2_15950 ( P1_U5734 , P1_ADD_405_U81 , P1_U2375 );
nand NAND2_15951 ( P1_U5735 , P1_ADD_515_U81 , P1_U2374 );
nand NAND2_15952 ( P1_U5736 , P1_U2370 , P1_REIP_REG_23_ );
nand NAND2_15953 ( P1_U5737 , P1_INSTADDRPOINTER_REG_23_ , P1_U5564 );
nand NAND2_15954 ( P1_U5738 , P1_R2099_U71 , P1_U2380 );
nand NAND2_15955 ( P1_U5739 , P1_R2027_U66 , P1_U2378 );
nand NAND2_15956 ( P1_U5740 , P1_R2278_U113 , P1_U2377 );
nand NAND2_15957 ( P1_U5741 , P1_ADD_405_U66 , P1_U2375 );
nand NAND2_15958 ( P1_U5742 , P1_ADD_515_U65 , P1_U2374 );
nand NAND2_15959 ( P1_U5743 , P1_U2370 , P1_REIP_REG_24_ );
nand NAND2_15960 ( P1_U5744 , P1_INSTADDRPOINTER_REG_24_ , P1_U5564 );
nand NAND2_15961 ( P1_U5745 , P1_R2099_U70 , P1_U2380 );
nand NAND2_15962 ( P1_U5746 , P1_R2027_U65 , P1_U2378 );
nand NAND2_15963 ( P1_U5747 , P1_R2278_U112 , P1_U2377 );
nand NAND2_15964 ( P1_U5748 , P1_ADD_405_U90 , P1_U2375 );
nand NAND2_15965 ( P1_U5749 , P1_ADD_515_U90 , P1_U2374 );
nand NAND2_15966 ( P1_U5750 , P1_U2370 , P1_REIP_REG_25_ );
nand NAND2_15967 ( P1_U5751 , P1_INSTADDRPOINTER_REG_25_ , P1_U5564 );
nand NAND2_15968 ( P1_U5752 , P1_R2099_U69 , P1_U2380 );
nand NAND2_15969 ( P1_U5753 , P1_R2027_U64 , P1_U2378 );
nand NAND2_15970 ( P1_U5754 , P1_R2278_U111 , P1_U2377 );
nand NAND2_15971 ( P1_U5755 , P1_ADD_405_U74 , P1_U2375 );
nand NAND2_15972 ( P1_U5756 , P1_ADD_515_U74 , P1_U2374 );
nand NAND2_15973 ( P1_U5757 , P1_U2370 , P1_REIP_REG_26_ );
nand NAND2_15974 ( P1_U5758 , P1_INSTADDRPOINTER_REG_26_ , P1_U5564 );
nand NAND2_15975 ( P1_U5759 , P1_R2099_U68 , P1_U2380 );
nand NAND2_15976 ( P1_U5760 , P1_R2027_U63 , P1_U2378 );
nand NAND2_15977 ( P1_U5761 , P1_R2278_U110 , P1_U2377 );
nand NAND2_15978 ( P1_U5762 , P1_ADD_405_U77 , P1_U2375 );
nand NAND2_15979 ( P1_U5763 , P1_ADD_515_U77 , P1_U2374 );
nand NAND2_15980 ( P1_U5764 , P1_U2370 , P1_REIP_REG_27_ );
nand NAND2_15981 ( P1_U5765 , P1_INSTADDRPOINTER_REG_27_ , P1_U5564 );
nand NAND2_15982 ( P1_U5766 , P1_R2099_U67 , P1_U2380 );
nand NAND2_15983 ( P1_U5767 , P1_R2027_U62 , P1_U2378 );
nand NAND2_15984 ( P1_U5768 , P1_R2278_U109 , P1_U2377 );
nand NAND2_15985 ( P1_U5769 , P1_ADD_405_U86 , P1_U2375 );
nand NAND2_15986 ( P1_U5770 , P1_ADD_515_U86 , P1_U2374 );
nand NAND2_15987 ( P1_U5771 , P1_U2370 , P1_REIP_REG_28_ );
nand NAND2_15988 ( P1_U5772 , P1_INSTADDRPOINTER_REG_28_ , P1_U5564 );
nand NAND2_15989 ( P1_U5773 , P1_R2099_U66 , P1_U2380 );
nand NAND2_15990 ( P1_U5774 , P1_R2027_U61 , P1_U2378 );
nand NAND2_15991 ( P1_U5775 , P1_R2278_U108 , P1_U2377 );
nand NAND2_15992 ( P1_U5776 , P1_ADD_405_U65 , P1_U2375 );
nand NAND2_15993 ( P1_U5777 , P1_ADD_515_U64 , P1_U2374 );
nand NAND2_15994 ( P1_U5778 , P1_U2370 , P1_REIP_REG_29_ );
nand NAND2_15995 ( P1_U5779 , P1_INSTADDRPOINTER_REG_29_ , P1_U5564 );
nand NAND2_15996 ( P1_U5780 , P1_R2099_U65 , P1_U2380 );
nand NAND2_15997 ( P1_U5781 , P1_R2027_U59 , P1_U2378 );
nand NAND2_15998 ( P1_U5782 , P1_R2278_U106 , P1_U2377 );
nand NAND2_15999 ( P1_U5783 , P1_ADD_405_U64 , P1_U2375 );
nand NAND2_16000 ( P1_U5784 , P1_ADD_515_U63 , P1_U2374 );
nand NAND2_16001 ( P1_U5785 , P1_U2370 , P1_REIP_REG_30_ );
nand NAND2_16002 ( P1_U5786 , P1_INSTADDRPOINTER_REG_30_ , P1_U5564 );
nand NAND2_16003 ( P1_U5787 , P1_R2099_U64 , P1_U2380 );
nand NAND2_16004 ( P1_U5788 , P1_R2027_U58 , P1_U2378 );
nand NAND2_16005 ( P1_U5789 , P1_R2278_U16 , P1_U2377 );
nand NAND2_16006 ( P1_U5790 , P1_ADD_405_U84 , P1_U2375 );
nand NAND2_16007 ( P1_U5791 , P1_ADD_515_U84 , P1_U2374 );
nand NAND2_16008 ( P1_U5792 , P1_U2370 , P1_REIP_REG_31_ );
nand NAND2_16009 ( P1_U5793 , P1_INSTADDRPOINTER_REG_31_ , P1_U5564 );
nand NAND2_16010 ( P1_U5794 , P1_U4209 , P1_U3294 );
not NOT1_16011 ( P1_U5795 , P1_U3416 );
nand NAND2_16012 ( P1_U5796 , P1_STATE2_REG_2_ , P1_U3294 );
nand NAND2_16013 ( P1_U5797 , P1_STATE2_REG_1_ , P1_U3308 );
nand NAND2_16014 ( P1_U5798 , P1_U5797 , P1_U5796 );
nand NAND2_16015 ( P1_U5799 , P1_PHYADDRPOINTER_REG_0_ , P1_U2376 );
nand NAND2_16016 ( P1_U5800 , P1_U2372 , P1_R2278_U99 );
nand NAND2_16017 ( P1_U5801 , P1_U2365 , P1_REIP_REG_0_ );
nand NAND2_16018 ( P1_U5802 , P1_R2358_U76 , P1_U2364 );
nand NAND2_16019 ( P1_U5803 , P1_PHYADDRPOINTER_REG_0_ , P1_U5795 );
nand NAND2_16020 ( P1_U5804 , P1_R2337_U4 , P1_U2376 );
nand NAND2_16021 ( P1_U5805 , P1_U2372 , P1_R2278_U19 );
nand NAND2_16022 ( P1_U5806 , P1_U2365 , P1_REIP_REG_1_ );
nand NAND2_16023 ( P1_U5807 , P1_R2358_U107 , P1_U2364 );
nand NAND2_16024 ( P1_U5808 , P1_PHYADDRPOINTER_REG_1_ , P1_U5795 );
nand NAND2_16025 ( P1_U5809 , P1_R2337_U71 , P1_U2376 );
nand NAND2_16026 ( P1_U5810 , P1_U2372 , P1_R2278_U107 );
nand NAND2_16027 ( P1_U5811 , P1_U2365 , P1_REIP_REG_2_ );
nand NAND2_16028 ( P1_U5812 , P1_R2358_U18 , P1_U2364 );
nand NAND2_16029 ( P1_U5813 , P1_PHYADDRPOINTER_REG_2_ , P1_U5795 );
nand NAND2_16030 ( P1_U5814 , P1_R2337_U68 , P1_U2376 );
nand NAND2_16031 ( P1_U5815 , P1_U2372 , P1_R2278_U105 );
nand NAND2_16032 ( P1_U5816 , P1_U2365 , P1_REIP_REG_3_ );
nand NAND2_16033 ( P1_U5817 , P1_R2358_U19 , P1_U2364 );
nand NAND2_16034 ( P1_U5818 , P1_PHYADDRPOINTER_REG_3_ , P1_U5795 );
nand NAND2_16035 ( P1_U5819 , P1_R2337_U67 , P1_U2376 );
nand NAND2_16036 ( P1_U5820 , P1_U2372 , P1_R2278_U104 );
nand NAND2_16037 ( P1_U5821 , P1_U2365 , P1_REIP_REG_4_ );
nand NAND2_16038 ( P1_U5822 , P1_R2358_U84 , P1_U2364 );
nand NAND2_16039 ( P1_U5823 , P1_PHYADDRPOINTER_REG_4_ , P1_U5795 );
nand NAND2_16040 ( P1_U5824 , P1_R2337_U66 , P1_U2376 );
nand NAND2_16041 ( P1_U5825 , P1_U2372 , P1_R2278_U17 );
nand NAND2_16042 ( P1_U5826 , P1_U2365 , P1_REIP_REG_5_ );
nand NAND2_16043 ( P1_U5827 , P1_R2358_U82 , P1_U2364 );
nand NAND2_16044 ( P1_U5828 , P1_PHYADDRPOINTER_REG_5_ , P1_U5795 );
nand NAND2_16045 ( P1_U5829 , P1_R2337_U65 , P1_U2376 );
nand NAND2_16046 ( P1_U5830 , P1_U2372 , P1_R2278_U103 );
nand NAND2_16047 ( P1_U5831 , P1_U2365 , P1_REIP_REG_6_ );
nand NAND2_16048 ( P1_U5832 , P1_R2358_U20 , P1_U2364 );
nand NAND2_16049 ( P1_U5833 , P1_PHYADDRPOINTER_REG_6_ , P1_U5795 );
nand NAND2_16050 ( P1_U5834 , P1_R2337_U64 , P1_U2376 );
nand NAND2_16051 ( P1_U5835 , P1_U2372 , P1_R2278_U18 );
nand NAND2_16052 ( P1_U5836 , P1_U2365 , P1_REIP_REG_7_ );
nand NAND2_16053 ( P1_U5837 , P1_R2358_U21 , P1_U2364 );
nand NAND2_16054 ( P1_U5838 , P1_PHYADDRPOINTER_REG_7_ , P1_U5795 );
nand NAND2_16055 ( P1_U5839 , P1_R2337_U63 , P1_U2376 );
nand NAND2_16056 ( P1_U5840 , P1_U2372 , P1_R2278_U102 );
nand NAND2_16057 ( P1_U5841 , P1_U2365 , P1_REIP_REG_8_ );
nand NAND2_16058 ( P1_U5842 , P1_R2358_U80 , P1_U2364 );
nand NAND2_16059 ( P1_U5843 , P1_PHYADDRPOINTER_REG_8_ , P1_U5795 );
nand NAND2_16060 ( P1_U5844 , P1_R2337_U62 , P1_U2376 );
nand NAND2_16061 ( P1_U5845 , P1_U2372 , P1_R2278_U101 );
nand NAND2_16062 ( P1_U5846 , P1_U2365 , P1_REIP_REG_9_ );
nand NAND2_16063 ( P1_U5847 , P1_R2358_U78 , P1_U2364 );
nand NAND2_16064 ( P1_U5848 , P1_PHYADDRPOINTER_REG_9_ , P1_U5795 );
nand NAND2_16065 ( P1_U5849 , P1_R2337_U91 , P1_U2376 );
nand NAND2_16066 ( P1_U5850 , P1_U2372 , P1_R2278_U126 );
nand NAND2_16067 ( P1_U5851 , P1_U2365 , P1_REIP_REG_10_ );
nand NAND2_16068 ( P1_U5852 , P1_R2358_U14 , P1_U2364 );
nand NAND2_16069 ( P1_U5853 , P1_PHYADDRPOINTER_REG_10_ , P1_U5795 );
nand NAND2_16070 ( P1_U5854 , P1_R2337_U90 , P1_U2376 );
nand NAND2_16071 ( P1_U5855 , P1_U2372 , P1_R2278_U15 );
nand NAND2_16072 ( P1_U5856 , P1_U2365 , P1_REIP_REG_11_ );
nand NAND2_16073 ( P1_U5857 , P1_R2358_U15 , P1_U2364 );
nand NAND2_16074 ( P1_U5858 , P1_PHYADDRPOINTER_REG_11_ , P1_U5795 );
nand NAND2_16075 ( P1_U5859 , P1_R2337_U89 , P1_U2376 );
nand NAND2_16076 ( P1_U5860 , P1_U2372 , P1_R2278_U125 );
nand NAND2_16077 ( P1_U5861 , P1_U2365 , P1_REIP_REG_12_ );
nand NAND2_16078 ( P1_U5862 , P1_R2358_U119 , P1_U2364 );
nand NAND2_16079 ( P1_U5863 , P1_PHYADDRPOINTER_REG_12_ , P1_U5795 );
nand NAND2_16080 ( P1_U5864 , P1_R2337_U88 , P1_U2376 );
nand NAND2_16081 ( P1_U5865 , P1_U2372 , P1_R2278_U123 );
nand NAND2_16082 ( P1_U5866 , P1_U2365 , P1_REIP_REG_13_ );
nand NAND2_16083 ( P1_U5867 , P1_R2358_U117 , P1_U2364 );
nand NAND2_16084 ( P1_U5868 , P1_PHYADDRPOINTER_REG_13_ , P1_U5795 );
nand NAND2_16085 ( P1_U5869 , P1_R2337_U87 , P1_U2376 );
nand NAND2_16086 ( P1_U5870 , P1_U2372 , P1_R2278_U122 );
nand NAND2_16087 ( P1_U5871 , P1_U2365 , P1_REIP_REG_14_ );
nand NAND2_16088 ( P1_U5872 , P1_R2358_U16 , P1_U2364 );
nand NAND2_16089 ( P1_U5873 , P1_PHYADDRPOINTER_REG_14_ , P1_U5795 );
nand NAND2_16090 ( P1_U5874 , P1_R2337_U86 , P1_U2376 );
nand NAND2_16091 ( P1_U5875 , P1_U2372 , P1_R2278_U20 );
nand NAND2_16092 ( P1_U5876 , P1_U2365 , P1_REIP_REG_15_ );
nand NAND2_16093 ( P1_U5877 , P1_R2358_U17 , P1_U2364 );
nand NAND2_16094 ( P1_U5878 , P1_PHYADDRPOINTER_REG_15_ , P1_U5795 );
nand NAND2_16095 ( P1_U5879 , P1_R2337_U85 , P1_U2376 );
nand NAND2_16096 ( P1_U5880 , P1_U2372 , P1_R2278_U121 );
nand NAND2_16097 ( P1_U5881 , P1_U2365 , P1_REIP_REG_16_ );
nand NAND2_16098 ( P1_U5882 , P1_R2358_U115 , P1_U2364 );
nand NAND2_16099 ( P1_U5883 , P1_PHYADDRPOINTER_REG_16_ , P1_U5795 );
nand NAND2_16100 ( P1_U5884 , P1_R2337_U84 , P1_U2376 );
nand NAND2_16101 ( P1_U5885 , P1_U2372 , P1_R2278_U120 );
nand NAND2_16102 ( P1_U5886 , P1_U2365 , P1_REIP_REG_17_ );
nand NAND2_16103 ( P1_U5887 , P1_R2358_U113 , P1_U2364 );
nand NAND2_16104 ( P1_U5888 , P1_PHYADDRPOINTER_REG_17_ , P1_U5795 );
nand NAND2_16105 ( P1_U5889 , P1_R2337_U83 , P1_U2376 );
nand NAND2_16106 ( P1_U5890 , P1_U2372 , P1_R2278_U119 );
nand NAND2_16107 ( P1_U5891 , P1_U2365 , P1_REIP_REG_18_ );
nand NAND2_16108 ( P1_U5892 , P1_R2358_U111 , P1_U2364 );
nand NAND2_16109 ( P1_U5893 , P1_PHYADDRPOINTER_REG_18_ , P1_U5795 );
nand NAND2_16110 ( P1_U5894 , P1_R2337_U82 , P1_U2376 );
nand NAND2_16111 ( P1_U5895 , P1_U2372 , P1_R2278_U118 );
nand NAND2_16112 ( P1_U5896 , P1_U2365 , P1_REIP_REG_19_ );
nand NAND2_16113 ( P1_U5897 , P1_R2358_U109 , P1_U2364 );
nand NAND2_16114 ( P1_U5898 , P1_PHYADDRPOINTER_REG_19_ , P1_U5795 );
nand NAND2_16115 ( P1_U5899 , P1_R2337_U81 , P1_U2376 );
nand NAND2_16116 ( P1_U5900 , P1_U2372 , P1_R2278_U117 );
nand NAND2_16117 ( P1_U5901 , P1_U2365 , P1_REIP_REG_20_ );
nand NAND2_16118 ( P1_U5902 , P1_R2358_U105 , P1_U2364 );
nand NAND2_16119 ( P1_U5903 , P1_PHYADDRPOINTER_REG_20_ , P1_U5795 );
nand NAND2_16120 ( P1_U5904 , P1_R2337_U80 , P1_U2376 );
nand NAND2_16121 ( P1_U5905 , P1_U2372 , P1_R2278_U116 );
nand NAND2_16122 ( P1_U5906 , P1_U2365 , P1_REIP_REG_21_ );
nand NAND2_16123 ( P1_U5907 , P1_R2358_U103 , P1_U2364 );
nand NAND2_16124 ( P1_U5908 , P1_PHYADDRPOINTER_REG_21_ , P1_U5795 );
nand NAND2_16125 ( P1_U5909 , P1_R2337_U79 , P1_U2376 );
nand NAND2_16126 ( P1_U5910 , P1_U2372 , P1_R2278_U115 );
nand NAND2_16127 ( P1_U5911 , P1_U2365 , P1_REIP_REG_22_ );
nand NAND2_16128 ( P1_U5912 , P1_R2358_U101 , P1_U2364 );
nand NAND2_16129 ( P1_U5913 , P1_PHYADDRPOINTER_REG_22_ , P1_U5795 );
nand NAND2_16130 ( P1_U5914 , P1_R2337_U78 , P1_U2376 );
nand NAND2_16131 ( P1_U5915 , P1_U2372 , P1_R2278_U114 );
nand NAND2_16132 ( P1_U5916 , P1_U2365 , P1_REIP_REG_23_ );
nand NAND2_16133 ( P1_U5917 , P1_R2358_U99 , P1_U2364 );
nand NAND2_16134 ( P1_U5918 , P1_PHYADDRPOINTER_REG_23_ , P1_U5795 );
nand NAND2_16135 ( P1_U5919 , P1_R2337_U77 , P1_U2376 );
nand NAND2_16136 ( P1_U5920 , P1_U2372 , P1_R2278_U113 );
nand NAND2_16137 ( P1_U5921 , P1_U2365 , P1_REIP_REG_24_ );
nand NAND2_16138 ( P1_U5922 , P1_R2358_U97 , P1_U2364 );
nand NAND2_16139 ( P1_U5923 , P1_PHYADDRPOINTER_REG_24_ , P1_U5795 );
nand NAND2_16140 ( P1_U5924 , P1_R2337_U76 , P1_U2376 );
nand NAND2_16141 ( P1_U5925 , P1_U2372 , P1_R2278_U112 );
nand NAND2_16142 ( P1_U5926 , P1_U2365 , P1_REIP_REG_25_ );
nand NAND2_16143 ( P1_U5927 , P1_R2358_U95 , P1_U2364 );
nand NAND2_16144 ( P1_U5928 , P1_PHYADDRPOINTER_REG_25_ , P1_U5795 );
nand NAND2_16145 ( P1_U5929 , P1_R2337_U75 , P1_U2376 );
nand NAND2_16146 ( P1_U5930 , P1_U2372 , P1_R2278_U111 );
nand NAND2_16147 ( P1_U5931 , P1_U2365 , P1_REIP_REG_26_ );
nand NAND2_16148 ( P1_U5932 , P1_R2358_U93 , P1_U2364 );
nand NAND2_16149 ( P1_U5933 , P1_PHYADDRPOINTER_REG_26_ , P1_U5795 );
nand NAND2_16150 ( P1_U5934 , P1_R2337_U74 , P1_U2376 );
nand NAND2_16151 ( P1_U5935 , P1_U2372 , P1_R2278_U110 );
nand NAND2_16152 ( P1_U5936 , P1_U2365 , P1_REIP_REG_27_ );
nand NAND2_16153 ( P1_U5937 , P1_R2358_U91 , P1_U2364 );
nand NAND2_16154 ( P1_U5938 , P1_PHYADDRPOINTER_REG_27_ , P1_U5795 );
nand NAND2_16155 ( P1_U5939 , P1_R2337_U73 , P1_U2376 );
nand NAND2_16156 ( P1_U5940 , P1_U2372 , P1_R2278_U109 );
nand NAND2_16157 ( P1_U5941 , P1_U2365 , P1_REIP_REG_28_ );
nand NAND2_16158 ( P1_U5942 , P1_R2358_U89 , P1_U2364 );
nand NAND2_16159 ( P1_U5943 , P1_PHYADDRPOINTER_REG_28_ , P1_U5795 );
nand NAND2_16160 ( P1_U5944 , P1_R2337_U72 , P1_U2376 );
nand NAND2_16161 ( P1_U5945 , P1_U2372 , P1_R2278_U108 );
nand NAND2_16162 ( P1_U5946 , P1_U2365 , P1_REIP_REG_29_ );
nand NAND2_16163 ( P1_U5947 , P1_R2358_U87 , P1_U2364 );
nand NAND2_16164 ( P1_U5948 , P1_PHYADDRPOINTER_REG_29_ , P1_U5795 );
nand NAND2_16165 ( P1_U5949 , P1_R2337_U70 , P1_U2376 );
nand NAND2_16166 ( P1_U5950 , P1_U2372 , P1_R2278_U106 );
nand NAND2_16167 ( P1_U5951 , P1_U2365 , P1_REIP_REG_30_ );
nand NAND2_16168 ( P1_U5952 , P1_R2358_U85 , P1_U2364 );
nand NAND2_16169 ( P1_U5953 , P1_PHYADDRPOINTER_REG_30_ , P1_U5795 );
nand NAND2_16170 ( P1_U5954 , P1_R2337_U69 , P1_U2376 );
nand NAND2_16171 ( P1_U5955 , P1_U2372 , P1_R2278_U16 );
nand NAND2_16172 ( P1_U5956 , P1_U2365 , P1_REIP_REG_31_ );
nand NAND2_16173 ( P1_U5957 , P1_R2358_U22 , P1_U2364 );
nand NAND2_16174 ( P1_U5958 , P1_PHYADDRPOINTER_REG_31_ , P1_U5795 );
nand NAND2_16175 ( P1_U5959 , U210 , P1_U3282 );
nand NAND2_16176 ( P1_U5960 , P1_EAX_REG_15_ , P1_U2382 );
nand NAND2_16177 ( P1_U5961 , U340 , P1_U2381 );
nand NAND2_16178 ( P1_U5962 , P1_U5961 , P1_U5960 );
nand NAND2_16179 ( P1_U5963 , P1_EAX_REG_14_ , P1_U2382 );
nand NAND2_16180 ( P1_U5964 , U341 , P1_U2381 );
nand NAND2_16181 ( P1_U5965 , P1_U5964 , P1_U5963 );
nand NAND2_16182 ( P1_U5966 , P1_EAX_REG_13_ , P1_U2382 );
nand NAND2_16183 ( P1_U5967 , U342 , P1_U2381 );
nand NAND2_16184 ( P1_U5968 , P1_U5967 , P1_U5966 );
nand NAND2_16185 ( P1_U5969 , P1_EAX_REG_12_ , P1_U2382 );
nand NAND2_16186 ( P1_U5970 , U343 , P1_U2381 );
nand NAND2_16187 ( P1_U5971 , P1_U5970 , P1_U5969 );
nand NAND2_16188 ( P1_U5972 , P1_EAX_REG_11_ , P1_U2382 );
nand NAND2_16189 ( P1_U5973 , U344 , P1_U2381 );
nand NAND2_16190 ( P1_U5974 , P1_U5973 , P1_U5972 );
nand NAND2_16191 ( P1_U5975 , P1_EAX_REG_10_ , P1_U2382 );
nand NAND2_16192 ( P1_U5976 , U345 , P1_U2381 );
nand NAND2_16193 ( P1_U5977 , P1_U5976 , P1_U5975 );
nand NAND2_16194 ( P1_U5978 , P1_EAX_REG_9_ , P1_U2382 );
nand NAND2_16195 ( P1_U5979 , U315 , P1_U2381 );
nand NAND2_16196 ( P1_U5980 , P1_U5979 , P1_U5978 );
nand NAND2_16197 ( P1_U5981 , P1_EAX_REG_8_ , P1_U2382 );
nand NAND2_16198 ( P1_U5982 , U316 , P1_U2381 );
nand NAND2_16199 ( P1_U5983 , P1_U5982 , P1_U5981 );
nand NAND2_16200 ( P1_U5984 , P1_EAX_REG_7_ , P1_U2382 );
nand NAND2_16201 ( P1_U5985 , P1_U2381 , U317 );
nand NAND2_16202 ( P1_U5986 , P1_U5985 , P1_U5984 );
nand NAND2_16203 ( P1_U5987 , P1_EAX_REG_6_ , P1_U2382 );
nand NAND2_16204 ( P1_U5988 , P1_U2381 , U318 );
nand NAND2_16205 ( P1_U5989 , P1_U5988 , P1_U5987 );
nand NAND2_16206 ( P1_U5990 , P1_EAX_REG_5_ , P1_U2382 );
nand NAND2_16207 ( P1_U5991 , P1_U2381 , U319 );
nand NAND2_16208 ( P1_U5992 , P1_U5991 , P1_U5990 );
nand NAND2_16209 ( P1_U5993 , P1_EAX_REG_4_ , P1_U2382 );
nand NAND2_16210 ( P1_U5994 , P1_U2381 , U320 );
nand NAND2_16211 ( P1_U5995 , P1_U5994 , P1_U5993 );
nand NAND2_16212 ( P1_U5996 , P1_EAX_REG_3_ , P1_U2382 );
nand NAND2_16213 ( P1_U5997 , P1_U2381 , U321 );
nand NAND2_16214 ( P1_U5998 , P1_U5997 , P1_U5996 );
nand NAND2_16215 ( P1_U5999 , P1_EAX_REG_2_ , P1_U2382 );
nand NAND2_16216 ( P1_U6000 , P1_U2381 , U324 );
nand NAND2_16217 ( P1_U6001 , P1_U6000 , P1_U5999 );
nand NAND2_16218 ( P1_U6002 , P1_EAX_REG_1_ , P1_U2382 );
nand NAND2_16219 ( P1_U6003 , P1_U2381 , U335 );
nand NAND2_16220 ( P1_U6004 , P1_U6003 , P1_U6002 );
nand NAND2_16221 ( P1_U6005 , P1_EAX_REG_0_ , P1_U2382 );
nand NAND2_16222 ( P1_U6006 , P1_U2381 , U346 );
nand NAND2_16223 ( P1_U6007 , P1_U6006 , P1_U6005 );
nand NAND2_16224 ( P1_U6008 , P1_EAX_REG_30_ , P1_U2382 );
nand NAND2_16225 ( P1_U6009 , U341 , P1_U2381 );
nand NAND2_16226 ( P1_U6010 , P1_U6009 , P1_U6008 );
nand NAND2_16227 ( P1_U6011 , P1_EAX_REG_29_ , P1_U2382 );
nand NAND2_16228 ( P1_U6012 , U342 , P1_U2381 );
nand NAND2_16229 ( P1_U6013 , P1_U6012 , P1_U6011 );
nand NAND2_16230 ( P1_U6014 , P1_EAX_REG_28_ , P1_U2382 );
nand NAND2_16231 ( P1_U6015 , U343 , P1_U2381 );
nand NAND2_16232 ( P1_U6016 , P1_U6015 , P1_U6014 );
nand NAND2_16233 ( P1_U6017 , P1_EAX_REG_27_ , P1_U2382 );
nand NAND2_16234 ( P1_U6018 , U344 , P1_U2381 );
nand NAND2_16235 ( P1_U6019 , P1_U6018 , P1_U6017 );
nand NAND2_16236 ( P1_U6020 , P1_EAX_REG_26_ , P1_U2382 );
nand NAND2_16237 ( P1_U6021 , U345 , P1_U2381 );
nand NAND2_16238 ( P1_U6022 , P1_U6021 , P1_U6020 );
nand NAND2_16239 ( P1_U6023 , P1_EAX_REG_25_ , P1_U2382 );
nand NAND2_16240 ( P1_U6024 , U315 , P1_U2381 );
nand NAND2_16241 ( P1_U6025 , P1_U6024 , P1_U6023 );
nand NAND2_16242 ( P1_U6026 , P1_EAX_REG_24_ , P1_U2382 );
nand NAND2_16243 ( P1_U6027 , U316 , P1_U2381 );
nand NAND2_16244 ( P1_U6028 , P1_U6027 , P1_U6026 );
nand NAND2_16245 ( P1_U6029 , P1_EAX_REG_23_ , P1_U2382 );
nand NAND2_16246 ( P1_U6030 , P1_U2381 , U317 );
nand NAND2_16247 ( P1_U6031 , P1_U6030 , P1_U6029 );
nand NAND2_16248 ( P1_U6032 , P1_EAX_REG_22_ , P1_U2382 );
nand NAND2_16249 ( P1_U6033 , P1_U2381 , U318 );
nand NAND2_16250 ( P1_U6034 , P1_U6033 , P1_U6032 );
nand NAND2_16251 ( P1_U6035 , P1_EAX_REG_21_ , P1_U2382 );
nand NAND2_16252 ( P1_U6036 , P1_U2381 , U319 );
nand NAND2_16253 ( P1_U6037 , P1_U6036 , P1_U6035 );
nand NAND2_16254 ( P1_U6038 , P1_EAX_REG_20_ , P1_U2382 );
nand NAND2_16255 ( P1_U6039 , P1_U2381 , U320 );
nand NAND2_16256 ( P1_U6040 , P1_U6039 , P1_U6038 );
nand NAND2_16257 ( P1_U6041 , P1_EAX_REG_19_ , P1_U2382 );
nand NAND2_16258 ( P1_U6042 , P1_U2381 , U321 );
nand NAND2_16259 ( P1_U6043 , P1_U6042 , P1_U6041 );
nand NAND2_16260 ( P1_U6044 , P1_EAX_REG_18_ , P1_U2382 );
nand NAND2_16261 ( P1_U6045 , P1_U2381 , U324 );
nand NAND2_16262 ( P1_U6046 , P1_U6045 , P1_U6044 );
nand NAND2_16263 ( P1_U6047 , P1_EAX_REG_17_ , P1_U2382 );
nand NAND2_16264 ( P1_U6048 , P1_U2381 , U335 );
nand NAND2_16265 ( P1_U6049 , P1_U6048 , P1_U6047 );
nand NAND2_16266 ( P1_U6050 , P1_EAX_REG_16_ , P1_U2382 );
nand NAND2_16267 ( P1_U6051 , P1_U2381 , U346 );
nand NAND2_16268 ( P1_U6052 , P1_U6051 , P1_U6050 );
nand NAND3_16269 ( P1_U6053 , P1_U4235 , P1_U7606 , P1_U4259 );
nand NAND2_16270 ( P1_U6054 , P1_U2428 , P1_U3294 );
not NOT1_16271 ( P1_U6055 , P1_U3417 );
nand NAND2_16272 ( P1_U6056 , P1_U2385 , P1_LWORD_REG_0_ );
nand NAND2_16273 ( P1_U6057 , P1_U2384 , P1_EAX_REG_0_ );
nand NAND2_16274 ( P1_U6058 , P1_DATAO_REG_0_ , P1_U6055 );
nand NAND2_16275 ( P1_U6059 , P1_U2385 , P1_LWORD_REG_1_ );
nand NAND2_16276 ( P1_U6060 , P1_U2384 , P1_EAX_REG_1_ );
nand NAND2_16277 ( P1_U6061 , P1_DATAO_REG_1_ , P1_U6055 );
nand NAND2_16278 ( P1_U6062 , P1_U2385 , P1_LWORD_REG_2_ );
nand NAND2_16279 ( P1_U6063 , P1_U2384 , P1_EAX_REG_2_ );
nand NAND2_16280 ( P1_U6064 , P1_DATAO_REG_2_ , P1_U6055 );
nand NAND2_16281 ( P1_U6065 , P1_U2385 , P1_LWORD_REG_3_ );
nand NAND2_16282 ( P1_U6066 , P1_U2384 , P1_EAX_REG_3_ );
nand NAND2_16283 ( P1_U6067 , P1_DATAO_REG_3_ , P1_U6055 );
nand NAND2_16284 ( P1_U6068 , P1_U2385 , P1_LWORD_REG_4_ );
nand NAND2_16285 ( P1_U6069 , P1_U2384 , P1_EAX_REG_4_ );
nand NAND2_16286 ( P1_U6070 , P1_DATAO_REG_4_ , P1_U6055 );
nand NAND2_16287 ( P1_U6071 , P1_U2385 , P1_LWORD_REG_5_ );
nand NAND2_16288 ( P1_U6072 , P1_U2384 , P1_EAX_REG_5_ );
nand NAND2_16289 ( P1_U6073 , P1_DATAO_REG_5_ , P1_U6055 );
nand NAND2_16290 ( P1_U6074 , P1_U2385 , P1_LWORD_REG_6_ );
nand NAND2_16291 ( P1_U6075 , P1_U2384 , P1_EAX_REG_6_ );
nand NAND2_16292 ( P1_U6076 , P1_DATAO_REG_6_ , P1_U6055 );
nand NAND2_16293 ( P1_U6077 , P1_U2385 , P1_LWORD_REG_7_ );
nand NAND2_16294 ( P1_U6078 , P1_U2384 , P1_EAX_REG_7_ );
nand NAND2_16295 ( P1_U6079 , P1_DATAO_REG_7_ , P1_U6055 );
nand NAND2_16296 ( P1_U6080 , P1_U2385 , P1_LWORD_REG_8_ );
nand NAND2_16297 ( P1_U6081 , P1_U2384 , P1_EAX_REG_8_ );
nand NAND2_16298 ( P1_U6082 , P1_DATAO_REG_8_ , P1_U6055 );
nand NAND2_16299 ( P1_U6083 , P1_U2385 , P1_LWORD_REG_9_ );
nand NAND2_16300 ( P1_U6084 , P1_U2384 , P1_EAX_REG_9_ );
nand NAND2_16301 ( P1_U6085 , P1_DATAO_REG_9_ , P1_U6055 );
nand NAND2_16302 ( P1_U6086 , P1_U2385 , P1_LWORD_REG_10_ );
nand NAND2_16303 ( P1_U6087 , P1_U2384 , P1_EAX_REG_10_ );
nand NAND2_16304 ( P1_U6088 , P1_DATAO_REG_10_ , P1_U6055 );
nand NAND2_16305 ( P1_U6089 , P1_U2385 , P1_LWORD_REG_11_ );
nand NAND2_16306 ( P1_U6090 , P1_U2384 , P1_EAX_REG_11_ );
nand NAND2_16307 ( P1_U6091 , P1_DATAO_REG_11_ , P1_U6055 );
nand NAND2_16308 ( P1_U6092 , P1_U2385 , P1_LWORD_REG_12_ );
nand NAND2_16309 ( P1_U6093 , P1_U2384 , P1_EAX_REG_12_ );
nand NAND2_16310 ( P1_U6094 , P1_DATAO_REG_12_ , P1_U6055 );
nand NAND2_16311 ( P1_U6095 , P1_U2385 , P1_LWORD_REG_13_ );
nand NAND2_16312 ( P1_U6096 , P1_U2384 , P1_EAX_REG_13_ );
nand NAND2_16313 ( P1_U6097 , P1_DATAO_REG_13_ , P1_U6055 );
nand NAND2_16314 ( P1_U6098 , P1_U2385 , P1_LWORD_REG_14_ );
nand NAND2_16315 ( P1_U6099 , P1_U2384 , P1_EAX_REG_14_ );
nand NAND2_16316 ( P1_U6100 , P1_DATAO_REG_14_ , P1_U6055 );
nand NAND2_16317 ( P1_U6101 , P1_U2385 , P1_LWORD_REG_15_ );
nand NAND2_16318 ( P1_U6102 , P1_U2384 , P1_EAX_REG_15_ );
nand NAND2_16319 ( P1_U6103 , P1_DATAO_REG_15_ , P1_U6055 );
nand NAND2_16320 ( P1_U6104 , P1_U2424 , P1_EAX_REG_16_ );
nand NAND2_16321 ( P1_U6105 , P1_U2385 , P1_UWORD_REG_0_ );
nand NAND2_16322 ( P1_U6106 , P1_DATAO_REG_16_ , P1_U6055 );
nand NAND2_16323 ( P1_U6107 , P1_U2424 , P1_EAX_REG_17_ );
nand NAND2_16324 ( P1_U6108 , P1_U2385 , P1_UWORD_REG_1_ );
nand NAND2_16325 ( P1_U6109 , P1_DATAO_REG_17_ , P1_U6055 );
nand NAND2_16326 ( P1_U6110 , P1_U2424 , P1_EAX_REG_18_ );
nand NAND2_16327 ( P1_U6111 , P1_U2385 , P1_UWORD_REG_2_ );
nand NAND2_16328 ( P1_U6112 , P1_DATAO_REG_18_ , P1_U6055 );
nand NAND2_16329 ( P1_U6113 , P1_U2424 , P1_EAX_REG_19_ );
nand NAND2_16330 ( P1_U6114 , P1_U2385 , P1_UWORD_REG_3_ );
nand NAND2_16331 ( P1_U6115 , P1_DATAO_REG_19_ , P1_U6055 );
nand NAND2_16332 ( P1_U6116 , P1_U2424 , P1_EAX_REG_20_ );
nand NAND2_16333 ( P1_U6117 , P1_U2385 , P1_UWORD_REG_4_ );
nand NAND2_16334 ( P1_U6118 , P1_DATAO_REG_20_ , P1_U6055 );
nand NAND2_16335 ( P1_U6119 , P1_U2424 , P1_EAX_REG_21_ );
nand NAND2_16336 ( P1_U6120 , P1_U2385 , P1_UWORD_REG_5_ );
nand NAND2_16337 ( P1_U6121 , P1_DATAO_REG_21_ , P1_U6055 );
nand NAND2_16338 ( P1_U6122 , P1_U2424 , P1_EAX_REG_22_ );
nand NAND2_16339 ( P1_U6123 , P1_U2385 , P1_UWORD_REG_6_ );
nand NAND2_16340 ( P1_U6124 , P1_DATAO_REG_22_ , P1_U6055 );
nand NAND2_16341 ( P1_U6125 , P1_U2424 , P1_EAX_REG_23_ );
nand NAND2_16342 ( P1_U6126 , P1_U2385 , P1_UWORD_REG_7_ );
nand NAND2_16343 ( P1_U6127 , P1_DATAO_REG_23_ , P1_U6055 );
nand NAND2_16344 ( P1_U6128 , P1_U2424 , P1_EAX_REG_24_ );
nand NAND2_16345 ( P1_U6129 , P1_U2385 , P1_UWORD_REG_8_ );
nand NAND2_16346 ( P1_U6130 , P1_DATAO_REG_24_ , P1_U6055 );
nand NAND2_16347 ( P1_U6131 , P1_U2424 , P1_EAX_REG_25_ );
nand NAND2_16348 ( P1_U6132 , P1_U2385 , P1_UWORD_REG_9_ );
nand NAND2_16349 ( P1_U6133 , P1_DATAO_REG_25_ , P1_U6055 );
nand NAND2_16350 ( P1_U6134 , P1_U2424 , P1_EAX_REG_26_ );
nand NAND2_16351 ( P1_U6135 , P1_U2385 , P1_UWORD_REG_10_ );
nand NAND2_16352 ( P1_U6136 , P1_DATAO_REG_26_ , P1_U6055 );
nand NAND2_16353 ( P1_U6137 , P1_U2424 , P1_EAX_REG_27_ );
nand NAND2_16354 ( P1_U6138 , P1_U2385 , P1_UWORD_REG_11_ );
nand NAND2_16355 ( P1_U6139 , P1_DATAO_REG_27_ , P1_U6055 );
nand NAND2_16356 ( P1_U6140 , P1_U2424 , P1_EAX_REG_28_ );
nand NAND2_16357 ( P1_U6141 , P1_U2385 , P1_UWORD_REG_12_ );
nand NAND2_16358 ( P1_U6142 , P1_DATAO_REG_28_ , P1_U6055 );
nand NAND2_16359 ( P1_U6143 , P1_U2424 , P1_EAX_REG_29_ );
nand NAND2_16360 ( P1_U6144 , P1_U2385 , P1_UWORD_REG_13_ );
nand NAND2_16361 ( P1_U6145 , P1_DATAO_REG_29_ , P1_U6055 );
nand NAND2_16362 ( P1_U6146 , P1_U2424 , P1_EAX_REG_30_ );
nand NAND2_16363 ( P1_U6147 , P1_U2385 , P1_UWORD_REG_14_ );
nand NAND2_16364 ( P1_U6148 , P1_DATAO_REG_30_ , P1_U6055 );
nand NAND3_16365 ( P1_U6149 , P1_U4194 , P1_U2447 , P1_GTE_485_U6 );
nand NAND3_16366 ( P1_U6150 , P1_U4254 , P1_U4197 , P1_U4194 );
nand NAND3_16367 ( P1_U6151 , P1_U4200 , P1_U3283 , P1_R2167_U17 );
nand NAND2_16368 ( P1_U6152 , P1_U7503 , P1_U3257 );
nand NAND2_16369 ( P1_U6153 , P1_U3883 , P1_U6152 );
nand NAND2_16370 ( P1_U6154 , P1_U2422 , U346 );
nand NAND2_16371 ( P1_U6155 , P1_U2386 , P1_R2358_U76 );
nand NAND2_16372 ( P1_U6156 , P1_EAX_REG_0_ , P1_U3424 );
nand NAND2_16373 ( P1_U6157 , P1_U2422 , U335 );
nand NAND2_16374 ( P1_U6158 , P1_U2386 , P1_R2358_U107 );
nand NAND2_16375 ( P1_U6159 , P1_EAX_REG_1_ , P1_U3424 );
nand NAND2_16376 ( P1_U6160 , P1_U2422 , U324 );
nand NAND2_16377 ( P1_U6161 , P1_U2386 , P1_R2358_U18 );
nand NAND2_16378 ( P1_U6162 , P1_EAX_REG_2_ , P1_U3424 );
nand NAND2_16379 ( P1_U6163 , P1_U2422 , U321 );
nand NAND2_16380 ( P1_U6164 , P1_U2386 , P1_R2358_U19 );
nand NAND2_16381 ( P1_U6165 , P1_EAX_REG_3_ , P1_U3424 );
nand NAND2_16382 ( P1_U6166 , P1_U2422 , U320 );
nand NAND2_16383 ( P1_U6167 , P1_U2386 , P1_R2358_U84 );
nand NAND2_16384 ( P1_U6168 , P1_EAX_REG_4_ , P1_U3424 );
nand NAND2_16385 ( P1_U6169 , P1_U2422 , U319 );
nand NAND2_16386 ( P1_U6170 , P1_U2386 , P1_R2358_U82 );
nand NAND2_16387 ( P1_U6171 , P1_EAX_REG_5_ , P1_U3424 );
nand NAND2_16388 ( P1_U6172 , P1_U2422 , U318 );
nand NAND2_16389 ( P1_U6173 , P1_U2386 , P1_R2358_U20 );
nand NAND2_16390 ( P1_U6174 , P1_EAX_REG_6_ , P1_U3424 );
nand NAND2_16391 ( P1_U6175 , P1_U2422 , U317 );
nand NAND2_16392 ( P1_U6176 , P1_U2386 , P1_R2358_U21 );
nand NAND2_16393 ( P1_U6177 , P1_EAX_REG_7_ , P1_U3424 );
nand NAND2_16394 ( P1_U6178 , P1_U2422 , U316 );
nand NAND2_16395 ( P1_U6179 , P1_U2386 , P1_R2358_U80 );
nand NAND2_16396 ( P1_U6180 , P1_EAX_REG_8_ , P1_U3424 );
nand NAND2_16397 ( P1_U6181 , P1_U2422 , U315 );
nand NAND2_16398 ( P1_U6182 , P1_U2386 , P1_R2358_U78 );
nand NAND2_16399 ( P1_U6183 , P1_EAX_REG_9_ , P1_U3424 );
nand NAND2_16400 ( P1_U6184 , P1_U2422 , U345 );
nand NAND2_16401 ( P1_U6185 , P1_U2386 , P1_R2358_U14 );
nand NAND2_16402 ( P1_U6186 , P1_EAX_REG_10_ , P1_U3424 );
nand NAND2_16403 ( P1_U6187 , P1_U2422 , U344 );
nand NAND2_16404 ( P1_U6188 , P1_U2386 , P1_R2358_U15 );
nand NAND2_16405 ( P1_U6189 , P1_EAX_REG_11_ , P1_U3424 );
nand NAND2_16406 ( P1_U6190 , P1_U2422 , U343 );
nand NAND2_16407 ( P1_U6191 , P1_U2386 , P1_R2358_U119 );
nand NAND2_16408 ( P1_U6192 , P1_EAX_REG_12_ , P1_U3424 );
nand NAND2_16409 ( P1_U6193 , P1_U2422 , U342 );
nand NAND2_16410 ( P1_U6194 , P1_U2386 , P1_R2358_U117 );
nand NAND2_16411 ( P1_U6195 , P1_EAX_REG_13_ , P1_U3424 );
nand NAND2_16412 ( P1_U6196 , P1_U2422 , U341 );
nand NAND2_16413 ( P1_U6197 , P1_U2386 , P1_R2358_U16 );
nand NAND2_16414 ( P1_U6198 , P1_EAX_REG_14_ , P1_U3424 );
nand NAND2_16415 ( P1_U6199 , P1_U2422 , U340 );
nand NAND2_16416 ( P1_U6200 , P1_U2386 , P1_R2358_U17 );
nand NAND2_16417 ( P1_U6201 , P1_EAX_REG_15_ , P1_U3424 );
nand NAND2_16418 ( P1_U6202 , P1_U2423 , U339 );
nand NAND2_16419 ( P1_U6203 , P1_U2387 , U346 );
nand NAND2_16420 ( P1_U6204 , P1_U2386 , P1_R2358_U115 );
nand NAND2_16421 ( P1_U6205 , P1_EAX_REG_16_ , P1_U3424 );
nand NAND2_16422 ( P1_U6206 , P1_U2423 , U338 );
nand NAND2_16423 ( P1_U6207 , P1_U2387 , U335 );
nand NAND2_16424 ( P1_U6208 , P1_U2386 , P1_R2358_U113 );
nand NAND2_16425 ( P1_U6209 , P1_EAX_REG_17_ , P1_U3424 );
nand NAND2_16426 ( P1_U6210 , P1_U2423 , U337 );
nand NAND2_16427 ( P1_U6211 , P1_U2387 , U324 );
nand NAND2_16428 ( P1_U6212 , P1_U2386 , P1_R2358_U111 );
nand NAND2_16429 ( P1_U6213 , P1_EAX_REG_18_ , P1_U3424 );
nand NAND2_16430 ( P1_U6214 , P1_U2423 , U336 );
nand NAND2_16431 ( P1_U6215 , P1_U2387 , U321 );
nand NAND2_16432 ( P1_U6216 , P1_U2386 , P1_R2358_U109 );
nand NAND2_16433 ( P1_U6217 , P1_EAX_REG_19_ , P1_U3424 );
nand NAND2_16434 ( P1_U6218 , P1_U2423 , U334 );
nand NAND2_16435 ( P1_U6219 , P1_U2387 , U320 );
nand NAND2_16436 ( P1_U6220 , P1_U2386 , P1_R2358_U105 );
nand NAND2_16437 ( P1_U6221 , P1_EAX_REG_20_ , P1_U3424 );
nand NAND2_16438 ( P1_U6222 , P1_U2423 , U333 );
nand NAND2_16439 ( P1_U6223 , P1_U2387 , U319 );
nand NAND2_16440 ( P1_U6224 , P1_U2386 , P1_R2358_U103 );
nand NAND2_16441 ( P1_U6225 , P1_EAX_REG_21_ , P1_U3424 );
nand NAND2_16442 ( P1_U6226 , P1_U2423 , U332 );
nand NAND2_16443 ( P1_U6227 , P1_U2387 , U318 );
nand NAND2_16444 ( P1_U6228 , P1_U2386 , P1_R2358_U101 );
nand NAND2_16445 ( P1_U6229 , P1_EAX_REG_22_ , P1_U3424 );
nand NAND2_16446 ( P1_U6230 , P1_U2423 , U331 );
nand NAND2_16447 ( P1_U6231 , P1_U2387 , U317 );
nand NAND2_16448 ( P1_U6232 , P1_U2386 , P1_R2358_U99 );
nand NAND2_16449 ( P1_U6233 , P1_EAX_REG_23_ , P1_U3424 );
nand NAND2_16450 ( P1_U6234 , P1_U2423 , U330 );
nand NAND2_16451 ( P1_U6235 , P1_U2387 , U316 );
nand NAND2_16452 ( P1_U6236 , P1_U2386 , P1_R2358_U97 );
nand NAND2_16453 ( P1_U6237 , P1_EAX_REG_24_ , P1_U3424 );
nand NAND2_16454 ( P1_U6238 , P1_U2423 , U329 );
nand NAND2_16455 ( P1_U6239 , P1_U2387 , U315 );
nand NAND2_16456 ( P1_U6240 , P1_U2386 , P1_R2358_U95 );
nand NAND2_16457 ( P1_U6241 , P1_EAX_REG_25_ , P1_U3424 );
nand NAND2_16458 ( P1_U6242 , P1_U2423 , U328 );
nand NAND2_16459 ( P1_U6243 , P1_U2387 , U345 );
nand NAND2_16460 ( P1_U6244 , P1_U2386 , P1_R2358_U93 );
nand NAND2_16461 ( P1_U6245 , P1_EAX_REG_26_ , P1_U3424 );
nand NAND2_16462 ( P1_U6246 , P1_U2423 , U327 );
nand NAND2_16463 ( P1_U6247 , P1_U2387 , U344 );
nand NAND2_16464 ( P1_U6248 , P1_U2386 , P1_R2358_U91 );
nand NAND2_16465 ( P1_U6249 , P1_EAX_REG_27_ , P1_U3424 );
nand NAND2_16466 ( P1_U6250 , P1_U2423 , U326 );
nand NAND2_16467 ( P1_U6251 , P1_U2387 , U343 );
nand NAND2_16468 ( P1_U6252 , P1_U2386 , P1_R2358_U89 );
nand NAND2_16469 ( P1_U6253 , P1_EAX_REG_28_ , P1_U3424 );
nand NAND2_16470 ( P1_U6254 , P1_U2423 , U325 );
nand NAND2_16471 ( P1_U6255 , P1_U2387 , U342 );
nand NAND2_16472 ( P1_U6256 , P1_U2386 , P1_R2358_U87 );
nand NAND2_16473 ( P1_U6257 , P1_EAX_REG_29_ , P1_U3424 );
nand NAND2_16474 ( P1_U6258 , P1_U2423 , U323 );
nand NAND2_16475 ( P1_U6259 , P1_U2387 , U341 );
nand NAND2_16476 ( P1_U6260 , P1_U2386 , P1_R2358_U85 );
nand NAND2_16477 ( P1_U6261 , P1_EAX_REG_30_ , P1_U3424 );
nand NAND2_16478 ( P1_U6262 , P1_U2423 , U322 );
nand NAND2_16479 ( P1_U6263 , P1_U4198 , P1_U3273 );
nand NAND2_16480 ( P1_U6264 , P1_U4205 , P1_U6263 );
nand NAND2_16481 ( P1_U6265 , P1_U2383 , P1_R2358_U76 );
nand NAND2_16482 ( P1_U6266 , P1_U2371 , P1_R2099_U86 );
nand NAND2_16483 ( P1_U6267 , P1_EBX_REG_0_ , P1_U3426 );
nand NAND2_16484 ( P1_U6268 , P1_U2383 , P1_R2358_U107 );
nand NAND2_16485 ( P1_U6269 , P1_U2371 , P1_R2099_U87 );
nand NAND2_16486 ( P1_U6270 , P1_EBX_REG_1_ , P1_U3426 );
nand NAND2_16487 ( P1_U6271 , P1_U2383 , P1_R2358_U18 );
nand NAND2_16488 ( P1_U6272 , P1_U2371 , P1_R2099_U138 );
nand NAND2_16489 ( P1_U6273 , P1_EBX_REG_2_ , P1_U3426 );
nand NAND2_16490 ( P1_U6274 , P1_U2383 , P1_R2358_U19 );
nand NAND2_16491 ( P1_U6275 , P1_U2371 , P1_R2099_U42 );
nand NAND2_16492 ( P1_U6276 , P1_EBX_REG_3_ , P1_U3426 );
nand NAND2_16493 ( P1_U6277 , P1_U2383 , P1_R2358_U84 );
nand NAND2_16494 ( P1_U6278 , P1_U2371 , P1_R2099_U41 );
nand NAND2_16495 ( P1_U6279 , P1_EBX_REG_4_ , P1_U3426 );
nand NAND2_16496 ( P1_U6280 , P1_U2383 , P1_R2358_U82 );
nand NAND2_16497 ( P1_U6281 , P1_U2371 , P1_R2099_U40 );
nand NAND2_16498 ( P1_U6282 , P1_EBX_REG_5_ , P1_U3426 );
nand NAND2_16499 ( P1_U6283 , P1_U2383 , P1_R2358_U20 );
nand NAND2_16500 ( P1_U6284 , P1_U2371 , P1_R2099_U39 );
nand NAND2_16501 ( P1_U6285 , P1_EBX_REG_6_ , P1_U3426 );
nand NAND2_16502 ( P1_U6286 , P1_U2383 , P1_R2358_U21 );
nand NAND2_16503 ( P1_U6287 , P1_U2371 , P1_R2099_U38 );
nand NAND2_16504 ( P1_U6288 , P1_EBX_REG_7_ , P1_U3426 );
nand NAND2_16505 ( P1_U6289 , P1_U2383 , P1_R2358_U80 );
nand NAND2_16506 ( P1_U6290 , P1_U2371 , P1_R2099_U37 );
nand NAND2_16507 ( P1_U6291 , P1_EBX_REG_8_ , P1_U3426 );
nand NAND2_16508 ( P1_U6292 , P1_U2383 , P1_R2358_U78 );
nand NAND2_16509 ( P1_U6293 , P1_U2371 , P1_R2099_U36 );
nand NAND2_16510 ( P1_U6294 , P1_EBX_REG_9_ , P1_U3426 );
nand NAND2_16511 ( P1_U6295 , P1_U2383 , P1_R2358_U14 );
nand NAND2_16512 ( P1_U6296 , P1_U2371 , P1_R2099_U85 );
nand NAND2_16513 ( P1_U6297 , P1_EBX_REG_10_ , P1_U3426 );
nand NAND2_16514 ( P1_U6298 , P1_U2383 , P1_R2358_U15 );
nand NAND2_16515 ( P1_U6299 , P1_U2371 , P1_R2099_U84 );
nand NAND2_16516 ( P1_U6300 , P1_EBX_REG_11_ , P1_U3426 );
nand NAND2_16517 ( P1_U6301 , P1_U2383 , P1_R2358_U119 );
nand NAND2_16518 ( P1_U6302 , P1_U2371 , P1_R2099_U83 );
nand NAND2_16519 ( P1_U6303 , P1_EBX_REG_12_ , P1_U3426 );
nand NAND2_16520 ( P1_U6304 , P1_U2383 , P1_R2358_U117 );
nand NAND2_16521 ( P1_U6305 , P1_U2371 , P1_R2099_U82 );
nand NAND2_16522 ( P1_U6306 , P1_EBX_REG_13_ , P1_U3426 );
nand NAND2_16523 ( P1_U6307 , P1_U2383 , P1_R2358_U16 );
nand NAND2_16524 ( P1_U6308 , P1_U2371 , P1_R2099_U81 );
nand NAND2_16525 ( P1_U6309 , P1_EBX_REG_14_ , P1_U3426 );
nand NAND2_16526 ( P1_U6310 , P1_U2383 , P1_R2358_U17 );
nand NAND2_16527 ( P1_U6311 , P1_U2371 , P1_R2099_U80 );
nand NAND2_16528 ( P1_U6312 , P1_EBX_REG_15_ , P1_U3426 );
nand NAND2_16529 ( P1_U6313 , P1_U2383 , P1_R2358_U115 );
nand NAND2_16530 ( P1_U6314 , P1_U2371 , P1_R2099_U79 );
nand NAND2_16531 ( P1_U6315 , P1_EBX_REG_16_ , P1_U3426 );
nand NAND2_16532 ( P1_U6316 , P1_U2383 , P1_R2358_U113 );
nand NAND2_16533 ( P1_U6317 , P1_U2371 , P1_R2099_U78 );
nand NAND2_16534 ( P1_U6318 , P1_EBX_REG_17_ , P1_U3426 );
nand NAND2_16535 ( P1_U6319 , P1_U2383 , P1_R2358_U111 );
nand NAND2_16536 ( P1_U6320 , P1_U2371 , P1_R2099_U77 );
nand NAND2_16537 ( P1_U6321 , P1_EBX_REG_18_ , P1_U3426 );
nand NAND2_16538 ( P1_U6322 , P1_U2383 , P1_R2358_U109 );
nand NAND2_16539 ( P1_U6323 , P1_U2371 , P1_R2099_U76 );
nand NAND2_16540 ( P1_U6324 , P1_EBX_REG_19_ , P1_U3426 );
nand NAND2_16541 ( P1_U6325 , P1_U2383 , P1_R2358_U105 );
nand NAND2_16542 ( P1_U6326 , P1_U2371 , P1_R2099_U75 );
nand NAND2_16543 ( P1_U6327 , P1_EBX_REG_20_ , P1_U3426 );
nand NAND2_16544 ( P1_U6328 , P1_U2383 , P1_R2358_U103 );
nand NAND2_16545 ( P1_U6329 , P1_U2371 , P1_R2099_U74 );
nand NAND2_16546 ( P1_U6330 , P1_EBX_REG_21_ , P1_U3426 );
nand NAND2_16547 ( P1_U6331 , P1_U2383 , P1_R2358_U101 );
nand NAND2_16548 ( P1_U6332 , P1_U2371 , P1_R2099_U73 );
nand NAND2_16549 ( P1_U6333 , P1_EBX_REG_22_ , P1_U3426 );
nand NAND2_16550 ( P1_U6334 , P1_U2383 , P1_R2358_U99 );
nand NAND2_16551 ( P1_U6335 , P1_U2371 , P1_R2099_U72 );
nand NAND2_16552 ( P1_U6336 , P1_EBX_REG_23_ , P1_U3426 );
nand NAND2_16553 ( P1_U6337 , P1_U2383 , P1_R2358_U97 );
nand NAND2_16554 ( P1_U6338 , P1_U2371 , P1_R2099_U71 );
nand NAND2_16555 ( P1_U6339 , P1_EBX_REG_24_ , P1_U3426 );
nand NAND2_16556 ( P1_U6340 , P1_U2383 , P1_R2358_U95 );
nand NAND2_16557 ( P1_U6341 , P1_U2371 , P1_R2099_U70 );
nand NAND2_16558 ( P1_U6342 , P1_EBX_REG_25_ , P1_U3426 );
nand NAND2_16559 ( P1_U6343 , P1_U2383 , P1_R2358_U93 );
nand NAND2_16560 ( P1_U6344 , P1_U2371 , P1_R2099_U69 );
nand NAND2_16561 ( P1_U6345 , P1_EBX_REG_26_ , P1_U3426 );
nand NAND2_16562 ( P1_U6346 , P1_U2383 , P1_R2358_U91 );
nand NAND2_16563 ( P1_U6347 , P1_U2371 , P1_R2099_U68 );
nand NAND2_16564 ( P1_U6348 , P1_EBX_REG_27_ , P1_U3426 );
nand NAND2_16565 ( P1_U6349 , P1_U2383 , P1_R2358_U89 );
nand NAND2_16566 ( P1_U6350 , P1_U2371 , P1_R2099_U67 );
nand NAND2_16567 ( P1_U6351 , P1_EBX_REG_28_ , P1_U3426 );
nand NAND2_16568 ( P1_U6352 , P1_U2383 , P1_R2358_U87 );
nand NAND2_16569 ( P1_U6353 , P1_U2371 , P1_R2099_U66 );
nand NAND2_16570 ( P1_U6354 , P1_EBX_REG_29_ , P1_U3426 );
nand NAND2_16571 ( P1_U6355 , P1_U2383 , P1_R2358_U85 );
nand NAND2_16572 ( P1_U6356 , P1_U2371 , P1_R2099_U65 );
nand NAND2_16573 ( P1_U6357 , P1_EBX_REG_30_ , P1_U3426 );
nand NAND2_16574 ( P1_U6358 , P1_U2371 , P1_R2099_U64 );
nand NAND2_16575 ( P1_U6359 , P1_EBX_REG_31_ , P1_U3426 );
nand NAND2_16576 ( P1_U6360 , P1_U4204 , P1_GTE_485_U6 );
nand NAND2_16577 ( P1_U6361 , P1_U4202 , P1_R2167_U17 );
nand NAND2_16578 ( P1_U6362 , P1_U4203 , P1_U3263 );
not NOT1_16579 ( P1_U6363 , P1_U3431 );
nand NAND2_16580 ( P1_U6364 , P1_U4249 , P1_STATE2_REG_2_ );
nand NAND2_16581 ( P1_U6365 , P1_R2337_U69 , P1_STATE2_REG_1_ );
nand NAND2_16582 ( P1_U6366 , P1_U6365 , P1_U6364 );
or OR2_16583 ( P1_U6367 , P1_STATEBS16_REG , U210 );
nand NAND2_16584 ( P1_U6368 , P1_U2604 , P1_R2099_U86 );
nand NAND2_16585 ( P1_U6369 , P1_REIP_REG_0_ , P1_U7485 );
nand NAND2_16586 ( P1_U6370 , P1_EBX_REG_0_ , P1_U7484 );
nand NAND2_16587 ( P1_U6371 , P1_U2429 , P1_R2358_U76 );
nand NAND2_16588 ( P1_U6372 , P1_U2426 , P1_R2182_U34 );
nand NAND2_16589 ( P1_U6373 , P1_U2373 , P1_PHYADDRPOINTER_REG_0_ );
nand NAND2_16590 ( P1_U6374 , P1_U2366 , P1_PHYADDRPOINTER_REG_0_ );
nand NAND2_16591 ( P1_U6375 , P1_U6363 , P1_REIP_REG_0_ );
nand NAND2_16592 ( P1_U6376 , P1_U2604 , P1_R2099_U87 );
nand NAND2_16593 ( P1_U6377 , P1_R2096_U4 , P1_U7485 );
nand NAND2_16594 ( P1_U6378 , P1_EBX_REG_1_ , P1_U7484 );
nand NAND2_16595 ( P1_U6379 , P1_U2429 , P1_R2358_U107 );
nand NAND2_16596 ( P1_U6380 , P1_U2426 , P1_R2182_U33 );
nand NAND2_16597 ( P1_U6381 , P1_U2373 , P1_PHYADDRPOINTER_REG_1_ );
nand NAND2_16598 ( P1_U6382 , P1_U2366 , P1_R2337_U4 );
nand NAND2_16599 ( P1_U6383 , P1_U6363 , P1_REIP_REG_1_ );
nand NAND2_16600 ( P1_U6384 , P1_U2604 , P1_R2099_U138 );
nand NAND2_16601 ( P1_U6385 , P1_R2096_U71 , P1_U7485 );
nand NAND2_16602 ( P1_U6386 , P1_EBX_REG_2_ , P1_U7484 );
nand NAND2_16603 ( P1_U6387 , P1_U2429 , P1_R2358_U18 );
nand NAND2_16604 ( P1_U6388 , P1_U2426 , P1_R2182_U42 );
nand NAND2_16605 ( P1_U6389 , P1_U2373 , P1_PHYADDRPOINTER_REG_2_ );
nand NAND2_16606 ( P1_U6390 , P1_U2366 , P1_R2337_U71 );
nand NAND2_16607 ( P1_U6391 , P1_U6363 , P1_REIP_REG_2_ );
nand NAND2_16608 ( P1_U6392 , P1_U2604 , P1_R2099_U42 );
nand NAND2_16609 ( P1_U6393 , P1_R2096_U68 , P1_U7485 );
nand NAND2_16610 ( P1_U6394 , P1_EBX_REG_3_ , P1_U7484 );
nand NAND2_16611 ( P1_U6395 , P1_U2429 , P1_R2358_U19 );
nand NAND2_16612 ( P1_U6396 , P1_U2426 , P1_R2182_U25 );
nand NAND2_16613 ( P1_U6397 , P1_U2373 , P1_PHYADDRPOINTER_REG_3_ );
nand NAND2_16614 ( P1_U6398 , P1_U2366 , P1_R2337_U68 );
nand NAND2_16615 ( P1_U6399 , P1_U6363 , P1_REIP_REG_3_ );
nand NAND2_16616 ( P1_U6400 , P1_U2604 , P1_R2099_U41 );
nand NAND2_16617 ( P1_U6401 , P1_R2096_U67 , P1_U7485 );
nand NAND2_16618 ( P1_U6402 , P1_EBX_REG_4_ , P1_U7484 );
nand NAND2_16619 ( P1_U6403 , P1_U2429 , P1_R2358_U84 );
nand NAND2_16620 ( P1_U6404 , P1_U2426 , P1_R2182_U24 );
nand NAND2_16621 ( P1_U6405 , P1_U2373 , P1_PHYADDRPOINTER_REG_4_ );
nand NAND2_16622 ( P1_U6406 , P1_U2366 , P1_R2337_U67 );
nand NAND2_16623 ( P1_U6407 , P1_U6363 , P1_REIP_REG_4_ );
nand NAND2_16624 ( P1_U6408 , P1_U2604 , P1_R2099_U40 );
nand NAND2_16625 ( P1_U6409 , P1_R2096_U66 , P1_U7485 );
nand NAND2_16626 ( P1_U6410 , P1_EBX_REG_5_ , P1_U7484 );
nand NAND2_16627 ( P1_U6411 , P1_U2429 , P1_R2358_U82 );
nand NAND2_16628 ( P1_U6412 , P1_R2182_U5 , P1_U2426 );
nand NAND2_16629 ( P1_U6413 , P1_U2373 , P1_PHYADDRPOINTER_REG_5_ );
nand NAND2_16630 ( P1_U6414 , P1_U2366 , P1_R2337_U66 );
nand NAND2_16631 ( P1_U6415 , P1_U6363 , P1_REIP_REG_5_ );
nand NAND2_16632 ( P1_U6416 , P1_U2604 , P1_R2099_U39 );
nand NAND2_16633 ( P1_U6417 , P1_R2096_U65 , P1_U7485 );
nand NAND2_16634 ( P1_U6418 , P1_EBX_REG_6_ , P1_U7484 );
nand NAND2_16635 ( P1_U6419 , P1_U2373 , P1_PHYADDRPOINTER_REG_6_ );
nand NAND2_16636 ( P1_U6420 , P1_U2367 , P1_R2358_U20 );
nand NAND2_16637 ( P1_U6421 , P1_U2366 , P1_R2337_U65 );
nand NAND2_16638 ( P1_U6422 , P1_U6363 , P1_REIP_REG_6_ );
nand NAND2_16639 ( P1_U6423 , P1_U2604 , P1_R2099_U38 );
nand NAND2_16640 ( P1_U6424 , P1_R2096_U64 , P1_U7485 );
nand NAND2_16641 ( P1_U6425 , P1_EBX_REG_7_ , P1_U7484 );
nand NAND2_16642 ( P1_U6426 , P1_U2373 , P1_PHYADDRPOINTER_REG_7_ );
nand NAND2_16643 ( P1_U6427 , P1_U2367 , P1_R2358_U21 );
nand NAND2_16644 ( P1_U6428 , P1_U2366 , P1_R2337_U64 );
nand NAND2_16645 ( P1_U6429 , P1_U6363 , P1_REIP_REG_7_ );
nand NAND2_16646 ( P1_U6430 , P1_U2604 , P1_R2099_U37 );
nand NAND2_16647 ( P1_U6431 , P1_R2096_U63 , P1_U7485 );
nand NAND2_16648 ( P1_U6432 , P1_EBX_REG_8_ , P1_U7484 );
nand NAND2_16649 ( P1_U6433 , P1_U2373 , P1_PHYADDRPOINTER_REG_8_ );
nand NAND2_16650 ( P1_U6434 , P1_U2367 , P1_R2358_U80 );
nand NAND2_16651 ( P1_U6435 , P1_U2366 , P1_R2337_U63 );
nand NAND2_16652 ( P1_U6436 , P1_U6363 , P1_REIP_REG_8_ );
nand NAND2_16653 ( P1_U6437 , P1_U2604 , P1_R2099_U36 );
nand NAND2_16654 ( P1_U6438 , P1_R2096_U62 , P1_U7485 );
nand NAND2_16655 ( P1_U6439 , P1_EBX_REG_9_ , P1_U7484 );
nand NAND2_16656 ( P1_U6440 , P1_U2373 , P1_PHYADDRPOINTER_REG_9_ );
nand NAND2_16657 ( P1_U6441 , P1_U2367 , P1_R2358_U78 );
nand NAND2_16658 ( P1_U6442 , P1_U2366 , P1_R2337_U62 );
nand NAND2_16659 ( P1_U6443 , P1_U6363 , P1_REIP_REG_9_ );
nand NAND2_16660 ( P1_U6444 , P1_U2604 , P1_R2099_U85 );
nand NAND2_16661 ( P1_U6445 , P1_R2096_U91 , P1_U7485 );
nand NAND2_16662 ( P1_U6446 , P1_EBX_REG_10_ , P1_U7484 );
nand NAND2_16663 ( P1_U6447 , P1_U2373 , P1_PHYADDRPOINTER_REG_10_ );
nand NAND2_16664 ( P1_U6448 , P1_U2367 , P1_R2358_U14 );
nand NAND2_16665 ( P1_U6449 , P1_U2366 , P1_R2337_U91 );
nand NAND2_16666 ( P1_U6450 , P1_U6363 , P1_REIP_REG_10_ );
nand NAND2_16667 ( P1_U6451 , P1_U2604 , P1_R2099_U84 );
nand NAND2_16668 ( P1_U6452 , P1_R2096_U90 , P1_U7485 );
nand NAND2_16669 ( P1_U6453 , P1_EBX_REG_11_ , P1_U7484 );
nand NAND2_16670 ( P1_U6454 , P1_U2373 , P1_PHYADDRPOINTER_REG_11_ );
nand NAND2_16671 ( P1_U6455 , P1_U2367 , P1_R2358_U15 );
nand NAND2_16672 ( P1_U6456 , P1_U2366 , P1_R2337_U90 );
nand NAND2_16673 ( P1_U6457 , P1_U6363 , P1_REIP_REG_11_ );
nand NAND2_16674 ( P1_U6458 , P1_U2604 , P1_R2099_U83 );
nand NAND2_16675 ( P1_U6459 , P1_R2096_U89 , P1_U7485 );
nand NAND2_16676 ( P1_U6460 , P1_EBX_REG_12_ , P1_U7484 );
nand NAND2_16677 ( P1_U6461 , P1_U2373 , P1_PHYADDRPOINTER_REG_12_ );
nand NAND2_16678 ( P1_U6462 , P1_U2367 , P1_R2358_U119 );
nand NAND2_16679 ( P1_U6463 , P1_U2366 , P1_R2337_U89 );
nand NAND2_16680 ( P1_U6464 , P1_U6363 , P1_REIP_REG_12_ );
nand NAND2_16681 ( P1_U6465 , P1_U2604 , P1_R2099_U82 );
nand NAND2_16682 ( P1_U6466 , P1_R2096_U88 , P1_U7485 );
nand NAND2_16683 ( P1_U6467 , P1_EBX_REG_13_ , P1_U7484 );
nand NAND2_16684 ( P1_U6468 , P1_U2373 , P1_PHYADDRPOINTER_REG_13_ );
nand NAND2_16685 ( P1_U6469 , P1_U2367 , P1_R2358_U117 );
nand NAND2_16686 ( P1_U6470 , P1_U2366 , P1_R2337_U88 );
nand NAND2_16687 ( P1_U6471 , P1_U6363 , P1_REIP_REG_13_ );
nand NAND2_16688 ( P1_U6472 , P1_U2604 , P1_R2099_U81 );
nand NAND2_16689 ( P1_U6473 , P1_R2096_U87 , P1_U7485 );
nand NAND2_16690 ( P1_U6474 , P1_EBX_REG_14_ , P1_U7484 );
nand NAND2_16691 ( P1_U6475 , P1_U2373 , P1_PHYADDRPOINTER_REG_14_ );
nand NAND2_16692 ( P1_U6476 , P1_U2367 , P1_R2358_U16 );
nand NAND2_16693 ( P1_U6477 , P1_U2366 , P1_R2337_U87 );
nand NAND2_16694 ( P1_U6478 , P1_U6363 , P1_REIP_REG_14_ );
nand NAND2_16695 ( P1_U6479 , P1_U2604 , P1_R2099_U80 );
nand NAND2_16696 ( P1_U6480 , P1_R2096_U86 , P1_U7485 );
nand NAND2_16697 ( P1_U6481 , P1_EBX_REG_15_ , P1_U7484 );
nand NAND2_16698 ( P1_U6482 , P1_U2373 , P1_PHYADDRPOINTER_REG_15_ );
nand NAND2_16699 ( P1_U6483 , P1_U2367 , P1_R2358_U17 );
nand NAND2_16700 ( P1_U6484 , P1_U2366 , P1_R2337_U86 );
nand NAND2_16701 ( P1_U6485 , P1_U6363 , P1_REIP_REG_15_ );
nand NAND2_16702 ( P1_U6486 , P1_U2604 , P1_R2099_U79 );
nand NAND2_16703 ( P1_U6487 , P1_R2096_U85 , P1_U7485 );
nand NAND2_16704 ( P1_U6488 , P1_EBX_REG_16_ , P1_U7484 );
nand NAND2_16705 ( P1_U6489 , P1_U2373 , P1_PHYADDRPOINTER_REG_16_ );
nand NAND2_16706 ( P1_U6490 , P1_U2367 , P1_R2358_U115 );
nand NAND2_16707 ( P1_U6491 , P1_U2366 , P1_R2337_U85 );
nand NAND2_16708 ( P1_U6492 , P1_U6363 , P1_REIP_REG_16_ );
nand NAND2_16709 ( P1_U6493 , P1_U2604 , P1_R2099_U78 );
nand NAND2_16710 ( P1_U6494 , P1_R2096_U84 , P1_U7485 );
nand NAND2_16711 ( P1_U6495 , P1_EBX_REG_17_ , P1_U7484 );
nand NAND2_16712 ( P1_U6496 , P1_U2373 , P1_PHYADDRPOINTER_REG_17_ );
nand NAND2_16713 ( P1_U6497 , P1_U2367 , P1_R2358_U113 );
nand NAND2_16714 ( P1_U6498 , P1_U2366 , P1_R2337_U84 );
nand NAND2_16715 ( P1_U6499 , P1_U6363 , P1_REIP_REG_17_ );
nand NAND2_16716 ( P1_U6500 , P1_U2604 , P1_R2099_U77 );
nand NAND2_16717 ( P1_U6501 , P1_R2096_U83 , P1_U7485 );
nand NAND2_16718 ( P1_U6502 , P1_EBX_REG_18_ , P1_U7484 );
nand NAND2_16719 ( P1_U6503 , P1_U2373 , P1_PHYADDRPOINTER_REG_18_ );
nand NAND2_16720 ( P1_U6504 , P1_U2367 , P1_R2358_U111 );
nand NAND2_16721 ( P1_U6505 , P1_U2366 , P1_R2337_U83 );
nand NAND2_16722 ( P1_U6506 , P1_U6363 , P1_REIP_REG_18_ );
nand NAND2_16723 ( P1_U6507 , P1_U2604 , P1_R2099_U76 );
nand NAND2_16724 ( P1_U6508 , P1_R2096_U82 , P1_U7485 );
nand NAND2_16725 ( P1_U6509 , P1_EBX_REG_19_ , P1_U7484 );
nand NAND2_16726 ( P1_U6510 , P1_U2373 , P1_PHYADDRPOINTER_REG_19_ );
nand NAND2_16727 ( P1_U6511 , P1_U2367 , P1_R2358_U109 );
nand NAND2_16728 ( P1_U6512 , P1_U2366 , P1_R2337_U82 );
nand NAND2_16729 ( P1_U6513 , P1_U6363 , P1_REIP_REG_19_ );
nand NAND2_16730 ( P1_U6514 , P1_U2604 , P1_R2099_U75 );
nand NAND2_16731 ( P1_U6515 , P1_R2096_U81 , P1_U7485 );
nand NAND2_16732 ( P1_U6516 , P1_EBX_REG_20_ , P1_U7484 );
nand NAND2_16733 ( P1_U6517 , P1_U2373 , P1_PHYADDRPOINTER_REG_20_ );
nand NAND2_16734 ( P1_U6518 , P1_U2367 , P1_R2358_U105 );
nand NAND2_16735 ( P1_U6519 , P1_U2366 , P1_R2337_U81 );
nand NAND2_16736 ( P1_U6520 , P1_U6363 , P1_REIP_REG_20_ );
nand NAND2_16737 ( P1_U6521 , P1_U2604 , P1_R2099_U74 );
nand NAND2_16738 ( P1_U6522 , P1_R2096_U80 , P1_U7485 );
nand NAND2_16739 ( P1_U6523 , P1_EBX_REG_21_ , P1_U7484 );
nand NAND2_16740 ( P1_U6524 , P1_U2373 , P1_PHYADDRPOINTER_REG_21_ );
nand NAND2_16741 ( P1_U6525 , P1_U2367 , P1_R2358_U103 );
nand NAND2_16742 ( P1_U6526 , P1_U2366 , P1_R2337_U80 );
nand NAND2_16743 ( P1_U6527 , P1_U6363 , P1_REIP_REG_21_ );
nand NAND2_16744 ( P1_U6528 , P1_U2604 , P1_R2099_U73 );
nand NAND2_16745 ( P1_U6529 , P1_R2096_U79 , P1_U7485 );
nand NAND2_16746 ( P1_U6530 , P1_EBX_REG_22_ , P1_U7484 );
nand NAND2_16747 ( P1_U6531 , P1_U2373 , P1_PHYADDRPOINTER_REG_22_ );
nand NAND2_16748 ( P1_U6532 , P1_U2367 , P1_R2358_U101 );
nand NAND2_16749 ( P1_U6533 , P1_U2366 , P1_R2337_U79 );
nand NAND2_16750 ( P1_U6534 , P1_U6363 , P1_REIP_REG_22_ );
nand NAND2_16751 ( P1_U6535 , P1_U2604 , P1_R2099_U72 );
nand NAND2_16752 ( P1_U6536 , P1_R2096_U78 , P1_U7485 );
nand NAND2_16753 ( P1_U6537 , P1_EBX_REG_23_ , P1_U7484 );
nand NAND2_16754 ( P1_U6538 , P1_U2373 , P1_PHYADDRPOINTER_REG_23_ );
nand NAND2_16755 ( P1_U6539 , P1_U2367 , P1_R2358_U99 );
nand NAND2_16756 ( P1_U6540 , P1_U2366 , P1_R2337_U78 );
nand NAND2_16757 ( P1_U6541 , P1_U6363 , P1_REIP_REG_23_ );
nand NAND2_16758 ( P1_U6542 , P1_U2604 , P1_R2099_U71 );
nand NAND2_16759 ( P1_U6543 , P1_R2096_U77 , P1_U7485 );
nand NAND2_16760 ( P1_U6544 , P1_EBX_REG_24_ , P1_U7484 );
nand NAND2_16761 ( P1_U6545 , P1_U2373 , P1_PHYADDRPOINTER_REG_24_ );
nand NAND2_16762 ( P1_U6546 , P1_U2367 , P1_R2358_U97 );
nand NAND2_16763 ( P1_U6547 , P1_U2366 , P1_R2337_U77 );
nand NAND2_16764 ( P1_U6548 , P1_U6363 , P1_REIP_REG_24_ );
nand NAND2_16765 ( P1_U6549 , P1_U2604 , P1_R2099_U70 );
nand NAND2_16766 ( P1_U6550 , P1_R2096_U76 , P1_U7485 );
nand NAND2_16767 ( P1_U6551 , P1_EBX_REG_25_ , P1_U7484 );
nand NAND2_16768 ( P1_U6552 , P1_U2373 , P1_PHYADDRPOINTER_REG_25_ );
nand NAND2_16769 ( P1_U6553 , P1_U2367 , P1_R2358_U95 );
nand NAND2_16770 ( P1_U6554 , P1_U2366 , P1_R2337_U76 );
nand NAND2_16771 ( P1_U6555 , P1_U6363 , P1_REIP_REG_25_ );
nand NAND2_16772 ( P1_U6556 , P1_U2604 , P1_R2099_U69 );
nand NAND2_16773 ( P1_U6557 , P1_R2096_U75 , P1_U7485 );
nand NAND2_16774 ( P1_U6558 , P1_EBX_REG_26_ , P1_U7484 );
nand NAND2_16775 ( P1_U6559 , P1_U2373 , P1_PHYADDRPOINTER_REG_26_ );
nand NAND2_16776 ( P1_U6560 , P1_U2367 , P1_R2358_U93 );
nand NAND2_16777 ( P1_U6561 , P1_U2366 , P1_R2337_U75 );
nand NAND2_16778 ( P1_U6562 , P1_U6363 , P1_REIP_REG_26_ );
nand NAND2_16779 ( P1_U6563 , P1_U2604 , P1_R2099_U68 );
nand NAND2_16780 ( P1_U6564 , P1_R2096_U74 , P1_U7485 );
nand NAND2_16781 ( P1_U6565 , P1_EBX_REG_27_ , P1_U7484 );
nand NAND2_16782 ( P1_U6566 , P1_U2373 , P1_PHYADDRPOINTER_REG_27_ );
nand NAND2_16783 ( P1_U6567 , P1_U2367 , P1_R2358_U91 );
nand NAND2_16784 ( P1_U6568 , P1_U2366 , P1_R2337_U74 );
nand NAND2_16785 ( P1_U6569 , P1_U6363 , P1_REIP_REG_27_ );
nand NAND2_16786 ( P1_U6570 , P1_U2604 , P1_R2099_U67 );
nand NAND2_16787 ( P1_U6571 , P1_R2096_U73 , P1_U7485 );
nand NAND2_16788 ( P1_U6572 , P1_EBX_REG_28_ , P1_U7484 );
nand NAND2_16789 ( P1_U6573 , P1_U2373 , P1_PHYADDRPOINTER_REG_28_ );
nand NAND2_16790 ( P1_U6574 , P1_U2367 , P1_R2358_U89 );
nand NAND2_16791 ( P1_U6575 , P1_U2366 , P1_R2337_U73 );
nand NAND2_16792 ( P1_U6576 , P1_U6363 , P1_REIP_REG_28_ );
nand NAND2_16793 ( P1_U6577 , P1_U2604 , P1_R2099_U66 );
nand NAND2_16794 ( P1_U6578 , P1_R2096_U72 , P1_U7485 );
nand NAND2_16795 ( P1_U6579 , P1_EBX_REG_29_ , P1_U7484 );
nand NAND2_16796 ( P1_U6580 , P1_U2373 , P1_PHYADDRPOINTER_REG_29_ );
nand NAND2_16797 ( P1_U6581 , P1_U2367 , P1_R2358_U87 );
nand NAND2_16798 ( P1_U6582 , P1_U2366 , P1_R2337_U72 );
nand NAND2_16799 ( P1_U6583 , P1_U6363 , P1_REIP_REG_29_ );
nand NAND2_16800 ( P1_U6584 , P1_U2604 , P1_R2099_U65 );
nand NAND2_16801 ( P1_U6585 , P1_R2096_U70 , P1_U7485 );
nand NAND2_16802 ( P1_U6586 , P1_EBX_REG_30_ , P1_U7484 );
nand NAND2_16803 ( P1_U6587 , P1_U2373 , P1_PHYADDRPOINTER_REG_30_ );
nand NAND2_16804 ( P1_U6588 , P1_U2367 , P1_R2358_U85 );
nand NAND2_16805 ( P1_U6589 , P1_U2366 , P1_R2337_U70 );
nand NAND2_16806 ( P1_U6590 , P1_U6363 , P1_REIP_REG_30_ );
nand NAND2_16807 ( P1_U6591 , P1_U2604 , P1_R2099_U64 );
nand NAND2_16808 ( P1_U6592 , P1_R2096_U69 , P1_U7485 );
nand NAND2_16809 ( P1_U6593 , P1_EBX_REG_31_ , P1_U7484 );
nand NAND2_16810 ( P1_U6594 , P1_U2373 , P1_PHYADDRPOINTER_REG_31_ );
nand NAND2_16811 ( P1_U6595 , P1_U2367 , P1_R2358_U22 );
nand NAND2_16812 ( P1_U6596 , P1_U2366 , P1_R2337_U69 );
nand NAND2_16813 ( P1_U6597 , P1_U6363 , P1_REIP_REG_31_ );
nand NAND2_16814 ( P1_U6598 , P1_DATAWIDTH_REG_1_ , P1_DATAWIDTH_REG_0_ );
or OR2_16815 ( P1_U6599 , P1_REIP_REG_1_ , P1_REIP_REG_0_ );
not NOT1_16816 ( P1_U6600 , P1_U4177 );
nand NAND2_16817 ( P1_U6601 , P1_FLUSH_REG , P1_U4177 );
nand NAND2_16818 ( P1_U6602 , P1_U3966 , P1_U2428 );
not NOT1_16819 ( P1_U6603 , P1_U4180 );
nand NAND2_16820 ( P1_U6604 , P1_STATEBS16_REG , P1_U4497 );
nand NAND2_16821 ( P1_U6605 , P1_U4208 , P1_U6604 );
nand NAND2_16822 ( P1_U6606 , P1_U3964 , P1_U6605 );
nand NAND2_16823 ( P1_U6607 , P1_STATE2_REG_0_ , P1_U6606 );
nand NAND2_16824 ( P1_U6608 , P1_U4193 , P1_U3272 );
nand NAND2_16825 ( P1_U6609 , P1_U3965 , P1_U6607 );
nand NAND2_16826 ( P1_U6610 , P1_U2368 , P1_U2473 );
nand NAND2_16827 ( P1_U6611 , P1_CODEFETCH_REG , P1_U6610 );
nand NAND2_16828 ( P1_U6612 , P1_U4255 , P1_STATE2_REG_0_ );
nand NAND2_16829 ( P1_U6613 , P1_ADS_N_REG , P1_STATE_REG_0_ );
not NOT1_16830 ( P1_U6614 , P1_U4181 );
nand NAND2_16831 ( P1_U6615 , P1_U3968 , P1_U3291 );
nand NAND3_16832 ( P1_U6616 , P1_U4499 , P1_U3969 , P1_U3406 );
nand NAND2_16833 ( P1_U6617 , P1_MEMORYFETCH_REG , P1_U6616 );
nand NAND2_16834 ( P1_U6618 , P1_U2544 , P1_INSTQUEUE_REG_15__7_ );
nand NAND2_16835 ( P1_U6619 , P1_U2543 , P1_INSTQUEUE_REG_14__7_ );
nand NAND2_16836 ( P1_U6620 , P1_U2542 , P1_INSTQUEUE_REG_13__7_ );
nand NAND2_16837 ( P1_U6621 , P1_U2541 , P1_INSTQUEUE_REG_12__7_ );
nand NAND2_16838 ( P1_U6622 , P1_U2539 , P1_INSTQUEUE_REG_11__7_ );
nand NAND2_16839 ( P1_U6623 , P1_U2538 , P1_INSTQUEUE_REG_10__7_ );
nand NAND2_16840 ( P1_U6624 , P1_U2537 , P1_INSTQUEUE_REG_9__7_ );
nand NAND2_16841 ( P1_U6625 , P1_U2536 , P1_INSTQUEUE_REG_8__7_ );
nand NAND2_16842 ( P1_U6626 , P1_U2534 , P1_INSTQUEUE_REG_7__7_ );
nand NAND2_16843 ( P1_U6627 , P1_U2533 , P1_INSTQUEUE_REG_6__7_ );
nand NAND2_16844 ( P1_U6628 , P1_U2532 , P1_INSTQUEUE_REG_5__7_ );
nand NAND2_16845 ( P1_U6629 , P1_U2531 , P1_INSTQUEUE_REG_4__7_ );
nand NAND2_16846 ( P1_U6630 , P1_U2529 , P1_INSTQUEUE_REG_3__7_ );
nand NAND2_16847 ( P1_U6631 , P1_U2527 , P1_INSTQUEUE_REG_2__7_ );
nand NAND2_16848 ( P1_U6632 , P1_U2525 , P1_INSTQUEUE_REG_1__7_ );
nand NAND2_16849 ( P1_U6633 , P1_U2523 , P1_INSTQUEUE_REG_0__7_ );
nand NAND2_16850 ( P1_U6634 , P1_U2544 , P1_INSTQUEUE_REG_15__6_ );
nand NAND2_16851 ( P1_U6635 , P1_U2543 , P1_INSTQUEUE_REG_14__6_ );
nand NAND2_16852 ( P1_U6636 , P1_U2542 , P1_INSTQUEUE_REG_13__6_ );
nand NAND2_16853 ( P1_U6637 , P1_U2541 , P1_INSTQUEUE_REG_12__6_ );
nand NAND2_16854 ( P1_U6638 , P1_U2539 , P1_INSTQUEUE_REG_11__6_ );
nand NAND2_16855 ( P1_U6639 , P1_U2538 , P1_INSTQUEUE_REG_10__6_ );
nand NAND2_16856 ( P1_U6640 , P1_U2537 , P1_INSTQUEUE_REG_9__6_ );
nand NAND2_16857 ( P1_U6641 , P1_U2536 , P1_INSTQUEUE_REG_8__6_ );
nand NAND2_16858 ( P1_U6642 , P1_U2534 , P1_INSTQUEUE_REG_7__6_ );
nand NAND2_16859 ( P1_U6643 , P1_U2533 , P1_INSTQUEUE_REG_6__6_ );
nand NAND2_16860 ( P1_U6644 , P1_U2532 , P1_INSTQUEUE_REG_5__6_ );
nand NAND2_16861 ( P1_U6645 , P1_U2531 , P1_INSTQUEUE_REG_4__6_ );
nand NAND2_16862 ( P1_U6646 , P1_U2529 , P1_INSTQUEUE_REG_3__6_ );
nand NAND2_16863 ( P1_U6647 , P1_U2527 , P1_INSTQUEUE_REG_2__6_ );
nand NAND2_16864 ( P1_U6648 , P1_U2525 , P1_INSTQUEUE_REG_1__6_ );
nand NAND2_16865 ( P1_U6649 , P1_U2523 , P1_INSTQUEUE_REG_0__6_ );
nand NAND2_16866 ( P1_U6650 , P1_U2544 , P1_INSTQUEUE_REG_15__5_ );
nand NAND2_16867 ( P1_U6651 , P1_U2543 , P1_INSTQUEUE_REG_14__5_ );
nand NAND2_16868 ( P1_U6652 , P1_U2542 , P1_INSTQUEUE_REG_13__5_ );
nand NAND2_16869 ( P1_U6653 , P1_U2541 , P1_INSTQUEUE_REG_12__5_ );
nand NAND2_16870 ( P1_U6654 , P1_U2539 , P1_INSTQUEUE_REG_11__5_ );
nand NAND2_16871 ( P1_U6655 , P1_U2538 , P1_INSTQUEUE_REG_10__5_ );
nand NAND2_16872 ( P1_U6656 , P1_U2537 , P1_INSTQUEUE_REG_9__5_ );
nand NAND2_16873 ( P1_U6657 , P1_U2536 , P1_INSTQUEUE_REG_8__5_ );
nand NAND2_16874 ( P1_U6658 , P1_U2534 , P1_INSTQUEUE_REG_7__5_ );
nand NAND2_16875 ( P1_U6659 , P1_U2533 , P1_INSTQUEUE_REG_6__5_ );
nand NAND2_16876 ( P1_U6660 , P1_U2532 , P1_INSTQUEUE_REG_5__5_ );
nand NAND2_16877 ( P1_U6661 , P1_U2531 , P1_INSTQUEUE_REG_4__5_ );
nand NAND2_16878 ( P1_U6662 , P1_U2529 , P1_INSTQUEUE_REG_3__5_ );
nand NAND2_16879 ( P1_U6663 , P1_U2527 , P1_INSTQUEUE_REG_2__5_ );
nand NAND2_16880 ( P1_U6664 , P1_U2525 , P1_INSTQUEUE_REG_1__5_ );
nand NAND2_16881 ( P1_U6665 , P1_U2523 , P1_INSTQUEUE_REG_0__5_ );
nand NAND2_16882 ( P1_U6666 , P1_U2544 , P1_INSTQUEUE_REG_15__4_ );
nand NAND2_16883 ( P1_U6667 , P1_U2543 , P1_INSTQUEUE_REG_14__4_ );
nand NAND2_16884 ( P1_U6668 , P1_U2542 , P1_INSTQUEUE_REG_13__4_ );
nand NAND2_16885 ( P1_U6669 , P1_U2541 , P1_INSTQUEUE_REG_12__4_ );
nand NAND2_16886 ( P1_U6670 , P1_U2539 , P1_INSTQUEUE_REG_11__4_ );
nand NAND2_16887 ( P1_U6671 , P1_U2538 , P1_INSTQUEUE_REG_10__4_ );
nand NAND2_16888 ( P1_U6672 , P1_U2537 , P1_INSTQUEUE_REG_9__4_ );
nand NAND2_16889 ( P1_U6673 , P1_U2536 , P1_INSTQUEUE_REG_8__4_ );
nand NAND2_16890 ( P1_U6674 , P1_U2534 , P1_INSTQUEUE_REG_7__4_ );
nand NAND2_16891 ( P1_U6675 , P1_U2533 , P1_INSTQUEUE_REG_6__4_ );
nand NAND2_16892 ( P1_U6676 , P1_U2532 , P1_INSTQUEUE_REG_5__4_ );
nand NAND2_16893 ( P1_U6677 , P1_U2531 , P1_INSTQUEUE_REG_4__4_ );
nand NAND2_16894 ( P1_U6678 , P1_U2529 , P1_INSTQUEUE_REG_3__4_ );
nand NAND2_16895 ( P1_U6679 , P1_U2527 , P1_INSTQUEUE_REG_2__4_ );
nand NAND2_16896 ( P1_U6680 , P1_U2525 , P1_INSTQUEUE_REG_1__4_ );
nand NAND2_16897 ( P1_U6681 , P1_U2544 , P1_INSTQUEUE_REG_15__3_ );
nand NAND2_16898 ( P1_U6682 , P1_U2543 , P1_INSTQUEUE_REG_14__3_ );
nand NAND2_16899 ( P1_U6683 , P1_U2542 , P1_INSTQUEUE_REG_13__3_ );
nand NAND2_16900 ( P1_U6684 , P1_U2541 , P1_INSTQUEUE_REG_12__3_ );
nand NAND2_16901 ( P1_U6685 , P1_U2539 , P1_INSTQUEUE_REG_11__3_ );
nand NAND2_16902 ( P1_U6686 , P1_U2538 , P1_INSTQUEUE_REG_10__3_ );
nand NAND2_16903 ( P1_U6687 , P1_U2537 , P1_INSTQUEUE_REG_9__3_ );
nand NAND2_16904 ( P1_U6688 , P1_U2536 , P1_INSTQUEUE_REG_8__3_ );
nand NAND2_16905 ( P1_U6689 , P1_U2534 , P1_INSTQUEUE_REG_7__3_ );
nand NAND2_16906 ( P1_U6690 , P1_U2533 , P1_INSTQUEUE_REG_6__3_ );
nand NAND2_16907 ( P1_U6691 , P1_U2532 , P1_INSTQUEUE_REG_5__3_ );
nand NAND2_16908 ( P1_U6692 , P1_U2531 , P1_INSTQUEUE_REG_4__3_ );
nand NAND2_16909 ( P1_U6693 , P1_U2529 , P1_INSTQUEUE_REG_3__3_ );
nand NAND2_16910 ( P1_U6694 , P1_U2527 , P1_INSTQUEUE_REG_2__3_ );
nand NAND2_16911 ( P1_U6695 , P1_U2525 , P1_INSTQUEUE_REG_1__3_ );
nand NAND2_16912 ( P1_U6696 , P1_U2523 , P1_INSTQUEUE_REG_0__3_ );
nand NAND2_16913 ( P1_U6697 , P1_U2544 , P1_INSTQUEUE_REG_15__2_ );
nand NAND2_16914 ( P1_U6698 , P1_U2543 , P1_INSTQUEUE_REG_14__2_ );
nand NAND2_16915 ( P1_U6699 , P1_U2542 , P1_INSTQUEUE_REG_13__2_ );
nand NAND2_16916 ( P1_U6700 , P1_U2541 , P1_INSTQUEUE_REG_12__2_ );
nand NAND2_16917 ( P1_U6701 , P1_U2539 , P1_INSTQUEUE_REG_11__2_ );
nand NAND2_16918 ( P1_U6702 , P1_U2538 , P1_INSTQUEUE_REG_10__2_ );
nand NAND2_16919 ( P1_U6703 , P1_U2537 , P1_INSTQUEUE_REG_9__2_ );
nand NAND2_16920 ( P1_U6704 , P1_U2536 , P1_INSTQUEUE_REG_8__2_ );
nand NAND2_16921 ( P1_U6705 , P1_U2534 , P1_INSTQUEUE_REG_7__2_ );
nand NAND2_16922 ( P1_U6706 , P1_U2533 , P1_INSTQUEUE_REG_6__2_ );
nand NAND2_16923 ( P1_U6707 , P1_U2532 , P1_INSTQUEUE_REG_5__2_ );
nand NAND2_16924 ( P1_U6708 , P1_U2531 , P1_INSTQUEUE_REG_4__2_ );
nand NAND2_16925 ( P1_U6709 , P1_U2529 , P1_INSTQUEUE_REG_3__2_ );
nand NAND2_16926 ( P1_U6710 , P1_U2527 , P1_INSTQUEUE_REG_2__2_ );
nand NAND2_16927 ( P1_U6711 , P1_U2525 , P1_INSTQUEUE_REG_1__2_ );
nand NAND2_16928 ( P1_U6712 , P1_U2523 , P1_INSTQUEUE_REG_0__2_ );
nand NAND2_16929 ( P1_U6713 , P1_U2544 , P1_INSTQUEUE_REG_15__1_ );
nand NAND2_16930 ( P1_U6714 , P1_U2543 , P1_INSTQUEUE_REG_14__1_ );
nand NAND2_16931 ( P1_U6715 , P1_U2542 , P1_INSTQUEUE_REG_13__1_ );
nand NAND2_16932 ( P1_U6716 , P1_U2541 , P1_INSTQUEUE_REG_12__1_ );
nand NAND2_16933 ( P1_U6717 , P1_U2539 , P1_INSTQUEUE_REG_11__1_ );
nand NAND2_16934 ( P1_U6718 , P1_U2538 , P1_INSTQUEUE_REG_10__1_ );
nand NAND2_16935 ( P1_U6719 , P1_U2537 , P1_INSTQUEUE_REG_9__1_ );
nand NAND2_16936 ( P1_U6720 , P1_U2536 , P1_INSTQUEUE_REG_8__1_ );
nand NAND2_16937 ( P1_U6721 , P1_U2534 , P1_INSTQUEUE_REG_7__1_ );
nand NAND2_16938 ( P1_U6722 , P1_U2533 , P1_INSTQUEUE_REG_6__1_ );
nand NAND2_16939 ( P1_U6723 , P1_U2532 , P1_INSTQUEUE_REG_5__1_ );
nand NAND2_16940 ( P1_U6724 , P1_U2531 , P1_INSTQUEUE_REG_4__1_ );
nand NAND2_16941 ( P1_U6725 , P1_U2529 , P1_INSTQUEUE_REG_3__1_ );
nand NAND2_16942 ( P1_U6726 , P1_U2527 , P1_INSTQUEUE_REG_2__1_ );
nand NAND2_16943 ( P1_U6727 , P1_U2525 , P1_INSTQUEUE_REG_1__1_ );
nand NAND2_16944 ( P1_U6728 , P1_U2523 , P1_INSTQUEUE_REG_0__1_ );
nand NAND2_16945 ( P1_U6729 , P1_U2544 , P1_INSTQUEUE_REG_15__0_ );
nand NAND2_16946 ( P1_U6730 , P1_U2543 , P1_INSTQUEUE_REG_14__0_ );
nand NAND2_16947 ( P1_U6731 , P1_U2542 , P1_INSTQUEUE_REG_13__0_ );
nand NAND2_16948 ( P1_U6732 , P1_U2541 , P1_INSTQUEUE_REG_12__0_ );
nand NAND2_16949 ( P1_U6733 , P1_U2539 , P1_INSTQUEUE_REG_11__0_ );
nand NAND2_16950 ( P1_U6734 , P1_U2538 , P1_INSTQUEUE_REG_10__0_ );
nand NAND2_16951 ( P1_U6735 , P1_U2537 , P1_INSTQUEUE_REG_9__0_ );
nand NAND2_16952 ( P1_U6736 , P1_U2536 , P1_INSTQUEUE_REG_8__0_ );
nand NAND2_16953 ( P1_U6737 , P1_U2534 , P1_INSTQUEUE_REG_7__0_ );
nand NAND2_16954 ( P1_U6738 , P1_U2533 , P1_INSTQUEUE_REG_6__0_ );
nand NAND2_16955 ( P1_U6739 , P1_U2532 , P1_INSTQUEUE_REG_5__0_ );
nand NAND2_16956 ( P1_U6740 , P1_U2531 , P1_INSTQUEUE_REG_4__0_ );
nand NAND2_16957 ( P1_U6741 , P1_U2529 , P1_INSTQUEUE_REG_3__0_ );
nand NAND2_16958 ( P1_U6742 , P1_U2527 , P1_INSTQUEUE_REG_2__0_ );
nand NAND2_16959 ( P1_U6743 , P1_U2525 , P1_INSTQUEUE_REG_1__0_ );
nand NAND2_16960 ( P1_U6744 , P1_U2523 , P1_INSTQUEUE_REG_0__0_ );
nand NAND2_16961 ( P1_U6745 , P1_U4460 , P1_STATE2_REG_2_ );
nand NAND2_16962 ( P1_U6746 , P1_U3412 , P1_U6745 );
nand NAND2_16963 ( P1_U6747 , P1_U4188 , P1_EAX_REG_9_ );
nand NAND2_16964 ( P1_U6748 , P1_U4187 , P1_PHYADDRPOINTER_REG_9_ );
nand NAND2_16965 ( P1_U6749 , P1_R2337_U62 , P1_U2352 );
nand NAND2_16966 ( P1_U6750 , P1_U4188 , P1_EAX_REG_8_ );
nand NAND2_16967 ( P1_U6751 , P1_U4187 , P1_PHYADDRPOINTER_REG_8_ );
nand NAND2_16968 ( P1_U6752 , P1_R2337_U63 , P1_U2352 );
nand NAND2_16969 ( P1_U6753 , P1_U4188 , P1_EAX_REG_7_ );
nand NAND2_16970 ( P1_U6754 , P1_U4187 , P1_PHYADDRPOINTER_REG_7_ );
nand NAND2_16971 ( P1_U6755 , P1_R2337_U64 , P1_U2352 );
nand NAND2_16972 ( P1_U6756 , P1_U4188 , P1_EAX_REG_6_ );
nand NAND2_16973 ( P1_U6757 , P1_U4187 , P1_PHYADDRPOINTER_REG_6_ );
nand NAND2_16974 ( P1_U6758 , P1_R2337_U65 , P1_U2352 );
nand NAND2_16975 ( P1_U6759 , P1_R2182_U5 , P1_U6746 );
nand NAND2_16976 ( P1_U6760 , P1_U4188 , P1_EAX_REG_5_ );
nand NAND2_16977 ( P1_U6761 , P1_U4187 , P1_PHYADDRPOINTER_REG_5_ );
nand NAND2_16978 ( P1_U6762 , P1_R2337_U66 , P1_U2352 );
nand NAND2_16979 ( P1_U6763 , P1_R2182_U24 , P1_U6746 );
nand NAND2_16980 ( P1_U6764 , P1_U4188 , P1_EAX_REG_4_ );
nand NAND2_16981 ( P1_U6765 , P1_U4187 , P1_PHYADDRPOINTER_REG_4_ );
nand NAND2_16982 ( P1_U6766 , P1_R2337_U67 , P1_U2352 );
nand NAND2_16983 ( P1_U6767 , P1_U2353 , P1_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_16984 ( P1_U6768 , P1_U4188 , P1_EAX_REG_31_ );
nand NAND2_16985 ( P1_U6769 , P1_U4187 , P1_PHYADDRPOINTER_REG_31_ );
nand NAND2_16986 ( P1_U6770 , P1_R2337_U69 , P1_U2352 );
nand NAND2_16987 ( P1_U6771 , P1_R2182_U26 , P1_U6746 );
nand NAND2_16988 ( P1_U6772 , P1_U4188 , P1_EAX_REG_30_ );
nand NAND2_16989 ( P1_U6773 , P1_U4187 , P1_PHYADDRPOINTER_REG_30_ );
nand NAND2_16990 ( P1_U6774 , P1_R2337_U70 , P1_U2352 );
nand NAND2_16991 ( P1_U6775 , P1_R2182_U25 , P1_U6746 );
nand NAND2_16992 ( P1_U6776 , P1_U4188 , P1_EAX_REG_3_ );
nand NAND2_16993 ( P1_U6777 , P1_U4187 , P1_PHYADDRPOINTER_REG_3_ );
nand NAND2_16994 ( P1_U6778 , P1_R2337_U68 , P1_U2352 );
nand NAND2_16995 ( P1_U6779 , P1_U2353 , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_16996 ( P1_U6780 , P1_R2182_U27 , P1_U6746 );
nand NAND2_16997 ( P1_U6781 , P1_U4188 , P1_EAX_REG_29_ );
nand NAND2_16998 ( P1_U6782 , P1_U4187 , P1_PHYADDRPOINTER_REG_29_ );
nand NAND2_16999 ( P1_U6783 , P1_R2337_U72 , P1_U2352 );
nand NAND2_17000 ( P1_U6784 , P1_R2182_U28 , P1_U6746 );
nand NAND2_17001 ( P1_U6785 , P1_U4188 , P1_EAX_REG_28_ );
nand NAND2_17002 ( P1_U6786 , P1_U4187 , P1_PHYADDRPOINTER_REG_28_ );
nand NAND2_17003 ( P1_U6787 , P1_R2337_U73 , P1_U2352 );
nand NAND2_17004 ( P1_U6788 , P1_R2182_U29 , P1_U6746 );
nand NAND2_17005 ( P1_U6789 , P1_U4188 , P1_EAX_REG_27_ );
nand NAND2_17006 ( P1_U6790 , P1_U4187 , P1_PHYADDRPOINTER_REG_27_ );
nand NAND2_17007 ( P1_U6791 , P1_R2337_U74 , P1_U2352 );
nand NAND2_17008 ( P1_U6792 , P1_R2182_U30 , P1_U6746 );
nand NAND2_17009 ( P1_U6793 , P1_U4188 , P1_EAX_REG_26_ );
nand NAND2_17010 ( P1_U6794 , P1_U4187 , P1_PHYADDRPOINTER_REG_26_ );
nand NAND2_17011 ( P1_U6795 , P1_R2337_U75 , P1_U2352 );
nand NAND2_17012 ( P1_U6796 , P1_R2182_U31 , P1_U6746 );
nand NAND2_17013 ( P1_U6797 , P1_U4188 , P1_EAX_REG_25_ );
nand NAND2_17014 ( P1_U6798 , P1_U4187 , P1_PHYADDRPOINTER_REG_25_ );
nand NAND2_17015 ( P1_U6799 , P1_R2337_U76 , P1_U2352 );
nand NAND2_17016 ( P1_U6800 , P1_R2182_U32 , P1_U6746 );
nand NAND2_17017 ( P1_U6801 , P1_U4188 , P1_EAX_REG_24_ );
nand NAND2_17018 ( P1_U6802 , P1_U4187 , P1_PHYADDRPOINTER_REG_24_ );
nand NAND2_17019 ( P1_U6803 , P1_R2337_U77 , P1_U2352 );
nand NAND2_17020 ( P1_U6804 , P1_R2182_U6 , P1_U6746 );
nand NAND2_17021 ( P1_U6805 , P1_U4188 , P1_EAX_REG_23_ );
nand NAND2_17022 ( P1_U6806 , P1_U4187 , P1_PHYADDRPOINTER_REG_23_ );
nand NAND2_17023 ( P1_U6807 , P1_R2337_U78 , P1_U2352 );
nand NAND2_17024 ( P1_U6808 , P1_U2724 , P1_U6746 );
nand NAND2_17025 ( P1_U6809 , P1_U4188 , P1_EAX_REG_22_ );
nand NAND2_17026 ( P1_U6810 , P1_U4187 , P1_PHYADDRPOINTER_REG_22_ );
nand NAND2_17027 ( P1_U6811 , P1_R2337_U79 , P1_U2352 );
nand NAND2_17028 ( P1_U6812 , P1_U2725 , P1_U6746 );
nand NAND2_17029 ( P1_U6813 , P1_U4188 , P1_EAX_REG_21_ );
nand NAND2_17030 ( P1_U6814 , P1_U4187 , P1_PHYADDRPOINTER_REG_21_ );
nand NAND2_17031 ( P1_U6815 , P1_R2337_U80 , P1_U2352 );
nand NAND2_17032 ( P1_U6816 , P1_U2726 , P1_U6746 );
nand NAND2_17033 ( P1_U6817 , P1_U4188 , P1_EAX_REG_20_ );
nand NAND2_17034 ( P1_U6818 , P1_U4187 , P1_PHYADDRPOINTER_REG_20_ );
nand NAND2_17035 ( P1_U6819 , P1_R2337_U81 , P1_U2352 );
nand NAND2_17036 ( P1_U6820 , P1_R2182_U42 , P1_U6746 );
nand NAND2_17037 ( P1_U6821 , P1_U4188 , P1_EAX_REG_2_ );
nand NAND2_17038 ( P1_U6822 , P1_U4187 , P1_PHYADDRPOINTER_REG_2_ );
nand NAND2_17039 ( P1_U6823 , P1_R2337_U71 , P1_U2352 );
nand NAND2_17040 ( P1_U6824 , P1_U2353 , P1_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_17041 ( P1_U6825 , P1_U2727 , P1_U6746 );
nand NAND2_17042 ( P1_U6826 , P1_U4188 , P1_EAX_REG_19_ );
nand NAND2_17043 ( P1_U6827 , P1_U4187 , P1_PHYADDRPOINTER_REG_19_ );
nand NAND2_17044 ( P1_U6828 , P1_R2337_U82 , P1_U2352 );
nand NAND2_17045 ( P1_U6829 , P1_U2728 , P1_U6746 );
nand NAND2_17046 ( P1_U6830 , P1_U4188 , P1_EAX_REG_18_ );
nand NAND2_17047 ( P1_U6831 , P1_U4187 , P1_PHYADDRPOINTER_REG_18_ );
nand NAND2_17048 ( P1_U6832 , P1_R2337_U83 , P1_U2352 );
nand NAND2_17049 ( P1_U6833 , P1_U2729 , P1_U6746 );
nand NAND2_17050 ( P1_U6834 , P1_U4188 , P1_EAX_REG_17_ );
nand NAND2_17051 ( P1_U6835 , P1_U4187 , P1_PHYADDRPOINTER_REG_17_ );
nand NAND2_17052 ( P1_U6836 , P1_R2337_U84 , P1_U2352 );
nand NAND2_17053 ( P1_U6837 , P1_U2730 , P1_U6746 );
nand NAND2_17054 ( P1_U6838 , P1_U4188 , P1_EAX_REG_16_ );
nand NAND2_17055 ( P1_U6839 , P1_U4187 , P1_PHYADDRPOINTER_REG_16_ );
nand NAND2_17056 ( P1_U6840 , P1_R2337_U85 , P1_U2352 );
nand NAND2_17057 ( P1_U6841 , P1_U4188 , P1_EAX_REG_15_ );
nand NAND2_17058 ( P1_U6842 , P1_U4187 , P1_PHYADDRPOINTER_REG_15_ );
nand NAND2_17059 ( P1_U6843 , P1_R2337_U86 , P1_U2352 );
nand NAND2_17060 ( P1_U6844 , P1_U4188 , P1_EAX_REG_14_ );
nand NAND2_17061 ( P1_U6845 , P1_U4187 , P1_PHYADDRPOINTER_REG_14_ );
nand NAND2_17062 ( P1_U6846 , P1_R2337_U87 , P1_U2352 );
nand NAND2_17063 ( P1_U6847 , P1_U4188 , P1_EAX_REG_13_ );
nand NAND2_17064 ( P1_U6848 , P1_U4187 , P1_PHYADDRPOINTER_REG_13_ );
nand NAND2_17065 ( P1_U6849 , P1_R2337_U88 , P1_U2352 );
nand NAND2_17066 ( P1_U6850 , P1_U4188 , P1_EAX_REG_12_ );
nand NAND2_17067 ( P1_U6851 , P1_U4187 , P1_PHYADDRPOINTER_REG_12_ );
nand NAND2_17068 ( P1_U6852 , P1_R2337_U89 , P1_U2352 );
nand NAND2_17069 ( P1_U6853 , P1_U4188 , P1_EAX_REG_11_ );
nand NAND2_17070 ( P1_U6854 , P1_U4187 , P1_PHYADDRPOINTER_REG_11_ );
nand NAND2_17071 ( P1_U6855 , P1_R2337_U90 , P1_U2352 );
nand NAND2_17072 ( P1_U6856 , P1_U4188 , P1_EAX_REG_10_ );
nand NAND2_17073 ( P1_U6857 , P1_U4187 , P1_PHYADDRPOINTER_REG_10_ );
nand NAND2_17074 ( P1_U6858 , P1_R2337_U91 , P1_U2352 );
nand NAND2_17075 ( P1_U6859 , P1_R2182_U33 , P1_U6746 );
nand NAND2_17076 ( P1_U6860 , P1_U4188 , P1_EAX_REG_1_ );
nand NAND2_17077 ( P1_U6861 , P1_U4187 , P1_PHYADDRPOINTER_REG_1_ );
nand NAND2_17078 ( P1_U6862 , P1_R2337_U4 , P1_U2352 );
nand NAND2_17079 ( P1_U6863 , P1_U2353 , P1_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_17080 ( P1_U6864 , P1_R2182_U34 , P1_U6746 );
nand NAND2_17081 ( P1_U6865 , P1_U4188 , P1_EAX_REG_0_ );
nand NAND2_17082 ( P1_U6866 , P1_U4187 , P1_PHYADDRPOINTER_REG_0_ );
nand NAND2_17083 ( P1_U6867 , P1_PHYADDRPOINTER_REG_0_ , P1_U2352 );
nand NAND2_17084 ( P1_U6868 , P1_U2353 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_17085 ( P1_U6869 , P1_R2144_U49 , P1_U6746 );
nand NAND3_17086 ( P1_U6870 , P1_U3439 , P1_U4460 , P1_U3309 );
nand NAND2_17087 ( P1_U6871 , P1_U4159 , P1_R2144_U80 );
nand NAND2_17088 ( P1_U6872 , P1_ADD_371_U6 , P1_U4208 );
nand NAND2_17089 ( P1_U6873 , P1_U4159 , P1_R2144_U10 );
nand NAND2_17090 ( P1_U6874 , P1_ADD_371_U21 , P1_U4208 );
nand NAND2_17091 ( P1_U6875 , P1_U4159 , P1_R2144_U9 );
nand NAND2_17092 ( P1_U6876 , P1_ADD_371_U17 , P1_U4208 );
nand NAND2_17093 ( P1_U6877 , P1_U4159 , P1_R2144_U45 );
nand NAND2_17094 ( P1_U6878 , P1_ADD_371_U19 , P1_U4208 );
nand NAND2_17095 ( P1_U6879 , P1_U4159 , P1_R2144_U47 );
nand NAND2_17096 ( P1_U6880 , P1_ADD_371_U18 , P1_U4208 );
nand NAND2_17097 ( P1_U6881 , P1_U4159 , P1_R2144_U8 );
nand NAND2_17098 ( P1_U6882 , P1_ADD_371_U24 , P1_U4208 );
nand NAND2_17099 ( P1_U6883 , P1_U4159 , P1_R2144_U49 );
nand NAND2_17100 ( P1_U6884 , P1_ADD_371_U5 , P1_U4208 );
nand NAND2_17101 ( P1_U6885 , P1_U4494 , P1_U3283 );
nand NAND2_17102 ( P1_U6886 , P1_U4159 , P1_R2144_U50 );
nand NAND2_17103 ( P1_U6887 , P1_ADD_371_U20 , P1_U4208 );
nand NAND2_17104 ( P1_U6888 , P1_U2605 , P1_U3284 );
nand NAND2_17105 ( P1_U6889 , P1_U4159 , P1_R2144_U43 );
nand NAND2_17106 ( P1_U6890 , P1_ADD_371_U4 , P1_U4208 );
nand NAND2_17107 ( P1_U6891 , P1_U4494 , P1_U3283 );
nand NAND2_17108 ( P1_U6892 , P1_U2564 , P1_INSTQUEUE_REG_15__1_ );
nand NAND2_17109 ( P1_U6893 , P1_U2563 , P1_INSTQUEUE_REG_14__1_ );
nand NAND2_17110 ( P1_U6894 , P1_U2562 , P1_INSTQUEUE_REG_13__1_ );
nand NAND2_17111 ( P1_U6895 , P1_U2561 , P1_INSTQUEUE_REG_12__1_ );
nand NAND2_17112 ( P1_U6896 , P1_U2559 , P1_INSTQUEUE_REG_11__1_ );
nand NAND2_17113 ( P1_U6897 , P1_U2558 , P1_INSTQUEUE_REG_10__1_ );
nand NAND2_17114 ( P1_U6898 , P1_U2557 , P1_INSTQUEUE_REG_9__1_ );
nand NAND2_17115 ( P1_U6899 , P1_U2556 , P1_INSTQUEUE_REG_8__1_ );
nand NAND2_17116 ( P1_U6900 , P1_U2554 , P1_INSTQUEUE_REG_7__1_ );
nand NAND2_17117 ( P1_U6901 , P1_U2553 , P1_INSTQUEUE_REG_6__1_ );
nand NAND2_17118 ( P1_U6902 , P1_U2552 , P1_INSTQUEUE_REG_5__1_ );
nand NAND2_17119 ( P1_U6903 , P1_U2551 , P1_INSTQUEUE_REG_4__1_ );
nand NAND2_17120 ( P1_U6904 , P1_U2549 , P1_INSTQUEUE_REG_3__1_ );
nand NAND2_17121 ( P1_U6905 , P1_U2548 , P1_INSTQUEUE_REG_2__1_ );
nand NAND2_17122 ( P1_U6906 , P1_U2547 , P1_INSTQUEUE_REG_1__1_ );
nand NAND2_17123 ( P1_U6907 , P1_U2546 , P1_INSTQUEUE_REG_0__1_ );
nand NAND4_17124 ( P1_U6908 , P1_U4032 , P1_U4031 , P1_U4030 , P1_U4029 );
nand NAND2_17125 ( P1_U6909 , P1_U3405 , P1_U3418 );
nand NAND2_17126 ( P1_U6910 , P1_U2564 , P1_INSTQUEUE_REG_15__0_ );
nand NAND2_17127 ( P1_U6911 , P1_U2563 , P1_INSTQUEUE_REG_14__0_ );
nand NAND2_17128 ( P1_U6912 , P1_U2562 , P1_INSTQUEUE_REG_13__0_ );
nand NAND2_17129 ( P1_U6913 , P1_U2561 , P1_INSTQUEUE_REG_12__0_ );
nand NAND2_17130 ( P1_U6914 , P1_U2559 , P1_INSTQUEUE_REG_11__0_ );
nand NAND2_17131 ( P1_U6915 , P1_U2558 , P1_INSTQUEUE_REG_10__0_ );
nand NAND2_17132 ( P1_U6916 , P1_U2557 , P1_INSTQUEUE_REG_9__0_ );
nand NAND2_17133 ( P1_U6917 , P1_U2556 , P1_INSTQUEUE_REG_8__0_ );
nand NAND2_17134 ( P1_U6918 , P1_U2554 , P1_INSTQUEUE_REG_7__0_ );
nand NAND2_17135 ( P1_U6919 , P1_U2553 , P1_INSTQUEUE_REG_6__0_ );
nand NAND2_17136 ( P1_U6920 , P1_U2552 , P1_INSTQUEUE_REG_5__0_ );
nand NAND2_17137 ( P1_U6921 , P1_U2551 , P1_INSTQUEUE_REG_4__0_ );
nand NAND2_17138 ( P1_U6922 , P1_U2549 , P1_INSTQUEUE_REG_3__0_ );
nand NAND2_17139 ( P1_U6923 , P1_U2548 , P1_INSTQUEUE_REG_2__0_ );
nand NAND2_17140 ( P1_U6924 , P1_U2547 , P1_INSTQUEUE_REG_1__0_ );
nand NAND2_17141 ( P1_U6925 , P1_U2546 , P1_INSTQUEUE_REG_0__0_ );
nand NAND4_17142 ( P1_U6926 , P1_U4036 , P1_U4035 , P1_U4034 , P1_U4033 );
nand NAND2_17143 ( P1_U6927 , P1_U4207 , P1_U3234 );
nand NAND2_17144 ( P1_U6928 , P1_U2355 , P1_SUB_357_U8 );
nand NAND2_17145 ( P1_U6929 , P1_U4207 , P1_U3233 );
nand NAND2_17146 ( P1_U6930 , P1_SUB_357_U6 , P1_U2355 );
nand NAND2_17147 ( P1_U6931 , P1_U4207 , P1_U3232 );
nand NAND2_17148 ( P1_U6932 , P1_SUB_357_U9 , P1_U2355 );
nand NAND2_17149 ( P1_U6933 , P1_U4207 , P1_U3231 );
nand NAND2_17150 ( P1_U6934 , P1_SUB_357_U13 , P1_U2355 );
nand NAND2_17151 ( P1_U6935 , P1_U4207 , P1_U3230 );
nand NAND2_17152 ( P1_U6936 , P1_SUB_357_U11 , P1_U2355 );
nand NAND2_17153 ( P1_U6937 , P1_R2182_U25 , P1_U3294 );
nand NAND2_17154 ( P1_U6938 , P1_U4207 , P1_U3229 );
nand NAND2_17155 ( P1_U6939 , P1_SUB_357_U12 , P1_U2355 );
nand NAND2_17156 ( P1_U6940 , P1_R2182_U42 , P1_U3294 );
nand NAND2_17157 ( P1_U6941 , P1_U2564 , P1_INSTQUEUE_REG_15__7_ );
nand NAND2_17158 ( P1_U6942 , P1_U2563 , P1_INSTQUEUE_REG_14__7_ );
nand NAND2_17159 ( P1_U6943 , P1_U2562 , P1_INSTQUEUE_REG_13__7_ );
nand NAND2_17160 ( P1_U6944 , P1_U2561 , P1_INSTQUEUE_REG_12__7_ );
nand NAND2_17161 ( P1_U6945 , P1_U2559 , P1_INSTQUEUE_REG_11__7_ );
nand NAND2_17162 ( P1_U6946 , P1_U2558 , P1_INSTQUEUE_REG_10__7_ );
nand NAND2_17163 ( P1_U6947 , P1_U2557 , P1_INSTQUEUE_REG_9__7_ );
nand NAND2_17164 ( P1_U6948 , P1_U2556 , P1_INSTQUEUE_REG_8__7_ );
nand NAND2_17165 ( P1_U6949 , P1_U2554 , P1_INSTQUEUE_REG_7__7_ );
nand NAND2_17166 ( P1_U6950 , P1_U2553 , P1_INSTQUEUE_REG_6__7_ );
nand NAND2_17167 ( P1_U6951 , P1_U2552 , P1_INSTQUEUE_REG_5__7_ );
nand NAND2_17168 ( P1_U6952 , P1_U2551 , P1_INSTQUEUE_REG_4__7_ );
nand NAND2_17169 ( P1_U6953 , P1_U2549 , P1_INSTQUEUE_REG_3__7_ );
nand NAND2_17170 ( P1_U6954 , P1_U2548 , P1_INSTQUEUE_REG_2__7_ );
nand NAND2_17171 ( P1_U6955 , P1_U2547 , P1_INSTQUEUE_REG_1__7_ );
nand NAND2_17172 ( P1_U6956 , P1_U2546 , P1_INSTQUEUE_REG_0__7_ );
nand NAND4_17173 ( P1_U6957 , P1_U4040 , P1_U4039 , P1_U4038 , P1_U4037 );
nand NAND2_17174 ( P1_U6958 , P1_U2564 , P1_INSTQUEUE_REG_15__6_ );
nand NAND2_17175 ( P1_U6959 , P1_U2563 , P1_INSTQUEUE_REG_14__6_ );
nand NAND2_17176 ( P1_U6960 , P1_U2562 , P1_INSTQUEUE_REG_13__6_ );
nand NAND2_17177 ( P1_U6961 , P1_U2561 , P1_INSTQUEUE_REG_12__6_ );
nand NAND2_17178 ( P1_U6962 , P1_U2559 , P1_INSTQUEUE_REG_11__6_ );
nand NAND2_17179 ( P1_U6963 , P1_U2558 , P1_INSTQUEUE_REG_10__6_ );
nand NAND2_17180 ( P1_U6964 , P1_U2557 , P1_INSTQUEUE_REG_9__6_ );
nand NAND2_17181 ( P1_U6965 , P1_U2556 , P1_INSTQUEUE_REG_8__6_ );
nand NAND2_17182 ( P1_U6966 , P1_U2554 , P1_INSTQUEUE_REG_7__6_ );
nand NAND2_17183 ( P1_U6967 , P1_U2553 , P1_INSTQUEUE_REG_6__6_ );
nand NAND2_17184 ( P1_U6968 , P1_U2552 , P1_INSTQUEUE_REG_5__6_ );
nand NAND2_17185 ( P1_U6969 , P1_U2551 , P1_INSTQUEUE_REG_4__6_ );
nand NAND2_17186 ( P1_U6970 , P1_U2549 , P1_INSTQUEUE_REG_3__6_ );
nand NAND2_17187 ( P1_U6971 , P1_U2548 , P1_INSTQUEUE_REG_2__6_ );
nand NAND2_17188 ( P1_U6972 , P1_U2547 , P1_INSTQUEUE_REG_1__6_ );
nand NAND2_17189 ( P1_U6973 , P1_U2546 , P1_INSTQUEUE_REG_0__6_ );
nand NAND4_17190 ( P1_U6974 , P1_U4044 , P1_U4043 , P1_U4042 , P1_U4041 );
nand NAND2_17191 ( P1_U6975 , P1_U2564 , P1_INSTQUEUE_REG_15__5_ );
nand NAND2_17192 ( P1_U6976 , P1_U2563 , P1_INSTQUEUE_REG_14__5_ );
nand NAND2_17193 ( P1_U6977 , P1_U2562 , P1_INSTQUEUE_REG_13__5_ );
nand NAND2_17194 ( P1_U6978 , P1_U2561 , P1_INSTQUEUE_REG_12__5_ );
nand NAND2_17195 ( P1_U6979 , P1_U2559 , P1_INSTQUEUE_REG_11__5_ );
nand NAND2_17196 ( P1_U6980 , P1_U2558 , P1_INSTQUEUE_REG_10__5_ );
nand NAND2_17197 ( P1_U6981 , P1_U2557 , P1_INSTQUEUE_REG_9__5_ );
nand NAND2_17198 ( P1_U6982 , P1_U2556 , P1_INSTQUEUE_REG_8__5_ );
nand NAND2_17199 ( P1_U6983 , P1_U2554 , P1_INSTQUEUE_REG_7__5_ );
nand NAND2_17200 ( P1_U6984 , P1_U2553 , P1_INSTQUEUE_REG_6__5_ );
nand NAND2_17201 ( P1_U6985 , P1_U2552 , P1_INSTQUEUE_REG_5__5_ );
nand NAND2_17202 ( P1_U6986 , P1_U2551 , P1_INSTQUEUE_REG_4__5_ );
nand NAND2_17203 ( P1_U6987 , P1_U2549 , P1_INSTQUEUE_REG_3__5_ );
nand NAND2_17204 ( P1_U6988 , P1_U2548 , P1_INSTQUEUE_REG_2__5_ );
nand NAND2_17205 ( P1_U6989 , P1_U2547 , P1_INSTQUEUE_REG_1__5_ );
nand NAND2_17206 ( P1_U6990 , P1_U2546 , P1_INSTQUEUE_REG_0__5_ );
nand NAND4_17207 ( P1_U6991 , P1_U4048 , P1_U4047 , P1_U4046 , P1_U4045 );
nand NAND2_17208 ( P1_U6992 , P1_U2564 , P1_INSTQUEUE_REG_15__4_ );
nand NAND2_17209 ( P1_U6993 , P1_U2563 , P1_INSTQUEUE_REG_14__4_ );
nand NAND2_17210 ( P1_U6994 , P1_U2562 , P1_INSTQUEUE_REG_13__4_ );
nand NAND2_17211 ( P1_U6995 , P1_U2561 , P1_INSTQUEUE_REG_12__4_ );
nand NAND2_17212 ( P1_U6996 , P1_U2559 , P1_INSTQUEUE_REG_11__4_ );
nand NAND2_17213 ( P1_U6997 , P1_U2558 , P1_INSTQUEUE_REG_10__4_ );
nand NAND2_17214 ( P1_U6998 , P1_U2557 , P1_INSTQUEUE_REG_9__4_ );
nand NAND2_17215 ( P1_U6999 , P1_U2556 , P1_INSTQUEUE_REG_8__4_ );
nand NAND2_17216 ( P1_U7000 , P1_U2554 , P1_INSTQUEUE_REG_7__4_ );
nand NAND2_17217 ( P1_U7001 , P1_U2553 , P1_INSTQUEUE_REG_6__4_ );
nand NAND2_17218 ( P1_U7002 , P1_U2552 , P1_INSTQUEUE_REG_5__4_ );
nand NAND2_17219 ( P1_U7003 , P1_U2551 , P1_INSTQUEUE_REG_4__4_ );
nand NAND2_17220 ( P1_U7004 , P1_U2549 , P1_INSTQUEUE_REG_3__4_ );
nand NAND2_17221 ( P1_U7005 , P1_U2548 , P1_INSTQUEUE_REG_2__4_ );
nand NAND2_17222 ( P1_U7006 , P1_U2547 , P1_INSTQUEUE_REG_1__4_ );
nand NAND2_17223 ( P1_U7007 , P1_U2564 , P1_INSTQUEUE_REG_15__3_ );
nand NAND2_17224 ( P1_U7008 , P1_U2563 , P1_INSTQUEUE_REG_14__3_ );
nand NAND2_17225 ( P1_U7009 , P1_U2562 , P1_INSTQUEUE_REG_13__3_ );
nand NAND2_17226 ( P1_U7010 , P1_U2561 , P1_INSTQUEUE_REG_12__3_ );
nand NAND2_17227 ( P1_U7011 , P1_U2559 , P1_INSTQUEUE_REG_11__3_ );
nand NAND2_17228 ( P1_U7012 , P1_U2558 , P1_INSTQUEUE_REG_10__3_ );
nand NAND2_17229 ( P1_U7013 , P1_U2557 , P1_INSTQUEUE_REG_9__3_ );
nand NAND2_17230 ( P1_U7014 , P1_U2556 , P1_INSTQUEUE_REG_8__3_ );
nand NAND2_17231 ( P1_U7015 , P1_U2554 , P1_INSTQUEUE_REG_7__3_ );
nand NAND2_17232 ( P1_U7016 , P1_U2553 , P1_INSTQUEUE_REG_6__3_ );
nand NAND2_17233 ( P1_U7017 , P1_U2552 , P1_INSTQUEUE_REG_5__3_ );
nand NAND2_17234 ( P1_U7018 , P1_U2551 , P1_INSTQUEUE_REG_4__3_ );
nand NAND2_17235 ( P1_U7019 , P1_U2549 , P1_INSTQUEUE_REG_3__3_ );
nand NAND2_17236 ( P1_U7020 , P1_U2548 , P1_INSTQUEUE_REG_2__3_ );
nand NAND2_17237 ( P1_U7021 , P1_U2547 , P1_INSTQUEUE_REG_1__3_ );
nand NAND2_17238 ( P1_U7022 , P1_U2546 , P1_INSTQUEUE_REG_0__3_ );
nand NAND4_17239 ( P1_U7023 , P1_U4056 , P1_U4055 , P1_U4054 , P1_U4053 );
nand NAND2_17240 ( P1_U7024 , P1_U2564 , P1_INSTQUEUE_REG_15__2_ );
nand NAND2_17241 ( P1_U7025 , P1_U2563 , P1_INSTQUEUE_REG_14__2_ );
nand NAND2_17242 ( P1_U7026 , P1_U2562 , P1_INSTQUEUE_REG_13__2_ );
nand NAND2_17243 ( P1_U7027 , P1_U2561 , P1_INSTQUEUE_REG_12__2_ );
nand NAND2_17244 ( P1_U7028 , P1_U2559 , P1_INSTQUEUE_REG_11__2_ );
nand NAND2_17245 ( P1_U7029 , P1_U2558 , P1_INSTQUEUE_REG_10__2_ );
nand NAND2_17246 ( P1_U7030 , P1_U2557 , P1_INSTQUEUE_REG_9__2_ );
nand NAND2_17247 ( P1_U7031 , P1_U2556 , P1_INSTQUEUE_REG_8__2_ );
nand NAND2_17248 ( P1_U7032 , P1_U2554 , P1_INSTQUEUE_REG_7__2_ );
nand NAND2_17249 ( P1_U7033 , P1_U2553 , P1_INSTQUEUE_REG_6__2_ );
nand NAND2_17250 ( P1_U7034 , P1_U2552 , P1_INSTQUEUE_REG_5__2_ );
nand NAND2_17251 ( P1_U7035 , P1_U2551 , P1_INSTQUEUE_REG_4__2_ );
nand NAND2_17252 ( P1_U7036 , P1_U2549 , P1_INSTQUEUE_REG_3__2_ );
nand NAND2_17253 ( P1_U7037 , P1_U2548 , P1_INSTQUEUE_REG_2__2_ );
nand NAND2_17254 ( P1_U7038 , P1_U2547 , P1_INSTQUEUE_REG_1__2_ );
nand NAND2_17255 ( P1_U7039 , P1_U2546 , P1_INSTQUEUE_REG_0__2_ );
nand NAND4_17256 ( P1_U7040 , P1_U4060 , P1_U4059 , P1_U4058 , P1_U4057 );
nand NAND2_17257 ( P1_U7041 , P1_U4207 , P1_U3228 );
nand NAND2_17258 ( P1_U7042 , P1_SUB_357_U7 , P1_U2355 );
nand NAND2_17259 ( P1_U7043 , P1_R2182_U33 , P1_U3294 );
nand NAND2_17260 ( P1_U7044 , P1_U4207 , P1_U3227 );
nand NAND2_17261 ( P1_U7045 , P1_SUB_357_U10 , P1_U2355 );
nand NAND2_17262 ( P1_U7046 , P1_R2182_U34 , P1_U3294 );
nand NAND2_17263 ( P1_U7047 , P1_U4206 , P1_U3234 );
nand NAND2_17264 ( P1_U7048 , P1_U4192 , P1_INSTQUEUE_REG_0__7_ );
nand NAND2_17265 ( P1_U7049 , P1_U4206 , P1_U3233 );
nand NAND2_17266 ( P1_U7050 , P1_U4192 , P1_INSTQUEUE_REG_0__6_ );
nand NAND2_17267 ( P1_U7051 , P1_U4206 , P1_U3232 );
nand NAND2_17268 ( P1_U7052 , P1_U4192 , P1_INSTQUEUE_REG_0__5_ );
nand NAND2_17269 ( P1_U7053 , P1_U4206 , P1_U3231 );
nand NAND2_17270 ( P1_U7054 , P1_U4206 , P1_U3230 );
nand NAND2_17271 ( P1_U7055 , P1_U4192 , P1_INSTQUEUE_REG_0__3_ );
nand NAND2_17272 ( P1_U7056 , P1_U4206 , P1_U3229 );
nand NAND2_17273 ( P1_U7057 , P1_U4192 , P1_INSTQUEUE_REG_0__2_ );
nand NAND2_17274 ( P1_U7058 , P1_U4206 , P1_U3228 );
nand NAND2_17275 ( P1_U7059 , P1_U4192 , P1_INSTQUEUE_REG_0__1_ );
nand NAND2_17276 ( P1_U7060 , P1_U4206 , P1_U3227 );
nand NAND2_17277 ( P1_U7061 , P1_U3234 , P1_U4400 );
nand NAND2_17278 ( P1_U7062 , P1_U4192 , P1_INSTQUEUE_REG_0__0_ );
nand NAND2_17279 ( P1_U7063 , P1_U3428 , P1_U3427 );
nand NAND2_17280 ( P1_U7064 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_U3264 );
not NOT1_17281 ( P1_U7065 , P1_U3445 );
nand NAND2_17282 ( P1_U7066 , P1_U2582 , P1_INSTQUEUE_REG_8__7_ );
nand NAND2_17283 ( P1_U7067 , P1_U2581 , P1_INSTQUEUE_REG_9__7_ );
nand NAND2_17284 ( P1_U7068 , P1_U2580 , P1_INSTQUEUE_REG_10__7_ );
nand NAND2_17285 ( P1_U7069 , P1_U2579 , P1_INSTQUEUE_REG_11__7_ );
nand NAND2_17286 ( P1_U7070 , P1_U2577 , P1_INSTQUEUE_REG_12__7_ );
nand NAND2_17287 ( P1_U7071 , P1_U2576 , P1_INSTQUEUE_REG_13__7_ );
nand NAND2_17288 ( P1_U7072 , P1_U2575 , P1_INSTQUEUE_REG_14__7_ );
nand NAND2_17289 ( P1_U7073 , P1_U2574 , P1_INSTQUEUE_REG_15__7_ );
nand NAND2_17290 ( P1_U7074 , P1_U2573 , P1_INSTQUEUE_REG_0__7_ );
nand NAND2_17291 ( P1_U7075 , P1_U2572 , P1_INSTQUEUE_REG_1__7_ );
nand NAND2_17292 ( P1_U7076 , P1_U2571 , P1_INSTQUEUE_REG_2__7_ );
nand NAND2_17293 ( P1_U7077 , P1_U2570 , P1_INSTQUEUE_REG_3__7_ );
nand NAND2_17294 ( P1_U7078 , P1_U2568 , P1_INSTQUEUE_REG_4__7_ );
nand NAND2_17295 ( P1_U7079 , P1_U2567 , P1_INSTQUEUE_REG_5__7_ );
nand NAND2_17296 ( P1_U7080 , P1_U2566 , P1_INSTQUEUE_REG_6__7_ );
nand NAND2_17297 ( P1_U7081 , P1_U2565 , P1_INSTQUEUE_REG_7__7_ );
nand NAND4_17298 ( P1_U7082 , P1_U4066 , P1_U4065 , P1_U4064 , P1_U4063 );
nand NAND2_17299 ( P1_U7083 , P1_U3425 , P1_U3421 );
nand NAND2_17300 ( P1_U7084 , P1_U4073 , P1_U4191 );
nand NAND2_17301 ( P1_U7085 , P1_U7084 , P1_U3422 );
nand NAND2_17302 ( P1_U7086 , P1_U4503 , P1_U3278 );
not NOT1_17303 ( P1_U7087 , P1_U3245 );
nand NAND4_17304 ( P1_U7088 , P1_U4400 , P1_U4503 , P1_U4154 , P1_U3394 );
nand NAND2_17305 ( P1_U7089 , P1_U4189 , P1_STATE2_REG_0_ );
nand NAND2_17306 ( P1_U7090 , P1_U4067 , P1_U3245 );
not NOT1_17307 ( P1_U7091 , P1_U3451 );
nand NAND3_17308 ( P1_U7092 , P1_U3451 , P1_U5492 , P1_U7629 );
nand NAND2_17309 ( P1_U7093 , P1_U4194 , P1_U7092 );
not NOT1_17310 ( P1_U7094 , P1_U3450 );
nand NAND2_17311 ( P1_U7095 , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_U3297 );
nand NAND2_17312 ( P1_U7096 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_U3450 );
nand NAND2_17313 ( P1_U7097 , P1_U4203 , P1_U3360 );
nand NAND2_17314 ( P1_U7098 , P1_U2582 , P1_INSTQUEUE_REG_8__6_ );
nand NAND2_17315 ( P1_U7099 , P1_U2581 , P1_INSTQUEUE_REG_9__6_ );
nand NAND2_17316 ( P1_U7100 , P1_U2580 , P1_INSTQUEUE_REG_10__6_ );
nand NAND2_17317 ( P1_U7101 , P1_U2579 , P1_INSTQUEUE_REG_11__6_ );
nand NAND2_17318 ( P1_U7102 , P1_U2577 , P1_INSTQUEUE_REG_12__6_ );
nand NAND2_17319 ( P1_U7103 , P1_U2576 , P1_INSTQUEUE_REG_13__6_ );
nand NAND2_17320 ( P1_U7104 , P1_U2575 , P1_INSTQUEUE_REG_14__6_ );
nand NAND2_17321 ( P1_U7105 , P1_U2574 , P1_INSTQUEUE_REG_15__6_ );
nand NAND2_17322 ( P1_U7106 , P1_U2573 , P1_INSTQUEUE_REG_0__6_ );
nand NAND2_17323 ( P1_U7107 , P1_U2572 , P1_INSTQUEUE_REG_1__6_ );
nand NAND2_17324 ( P1_U7108 , P1_U2571 , P1_INSTQUEUE_REG_2__6_ );
nand NAND2_17325 ( P1_U7109 , P1_U2570 , P1_INSTQUEUE_REG_3__6_ );
nand NAND2_17326 ( P1_U7110 , P1_U2568 , P1_INSTQUEUE_REG_4__6_ );
nand NAND2_17327 ( P1_U7111 , P1_U2567 , P1_INSTQUEUE_REG_5__6_ );
nand NAND2_17328 ( P1_U7112 , P1_U2566 , P1_INSTQUEUE_REG_6__6_ );
nand NAND2_17329 ( P1_U7113 , P1_U2565 , P1_INSTQUEUE_REG_7__6_ );
nand NAND4_17330 ( P1_U7114 , P1_U4082 , P1_U4081 , P1_U4080 , P1_U4079 );
nand NAND2_17331 ( P1_U7115 , P1_U2582 , P1_INSTQUEUE_REG_8__5_ );
nand NAND2_17332 ( P1_U7116 , P1_U2581 , P1_INSTQUEUE_REG_9__5_ );
nand NAND2_17333 ( P1_U7117 , P1_U2580 , P1_INSTQUEUE_REG_10__5_ );
nand NAND2_17334 ( P1_U7118 , P1_U2579 , P1_INSTQUEUE_REG_11__5_ );
nand NAND2_17335 ( P1_U7119 , P1_U2577 , P1_INSTQUEUE_REG_12__5_ );
nand NAND2_17336 ( P1_U7120 , P1_U2576 , P1_INSTQUEUE_REG_13__5_ );
nand NAND2_17337 ( P1_U7121 , P1_U2575 , P1_INSTQUEUE_REG_14__5_ );
nand NAND2_17338 ( P1_U7122 , P1_U2574 , P1_INSTQUEUE_REG_15__5_ );
nand NAND2_17339 ( P1_U7123 , P1_U2573 , P1_INSTQUEUE_REG_0__5_ );
nand NAND2_17340 ( P1_U7124 , P1_U2572 , P1_INSTQUEUE_REG_1__5_ );
nand NAND2_17341 ( P1_U7125 , P1_U2571 , P1_INSTQUEUE_REG_2__5_ );
nand NAND2_17342 ( P1_U7126 , P1_U2570 , P1_INSTQUEUE_REG_3__5_ );
nand NAND2_17343 ( P1_U7127 , P1_U2568 , P1_INSTQUEUE_REG_4__5_ );
nand NAND2_17344 ( P1_U7128 , P1_U2567 , P1_INSTQUEUE_REG_5__5_ );
nand NAND2_17345 ( P1_U7129 , P1_U2566 , P1_INSTQUEUE_REG_6__5_ );
nand NAND2_17346 ( P1_U7130 , P1_U2565 , P1_INSTQUEUE_REG_7__5_ );
nand NAND4_17347 ( P1_U7131 , P1_U4086 , P1_U4085 , P1_U4084 , P1_U4083 );
nand NAND2_17348 ( P1_U7132 , P1_U2582 , P1_INSTQUEUE_REG_8__4_ );
nand NAND2_17349 ( P1_U7133 , P1_U2581 , P1_INSTQUEUE_REG_9__4_ );
nand NAND2_17350 ( P1_U7134 , P1_U2580 , P1_INSTQUEUE_REG_10__4_ );
nand NAND2_17351 ( P1_U7135 , P1_U2579 , P1_INSTQUEUE_REG_11__4_ );
nand NAND2_17352 ( P1_U7136 , P1_U2577 , P1_INSTQUEUE_REG_12__4_ );
nand NAND2_17353 ( P1_U7137 , P1_U2576 , P1_INSTQUEUE_REG_13__4_ );
nand NAND2_17354 ( P1_U7138 , P1_U2575 , P1_INSTQUEUE_REG_14__4_ );
nand NAND2_17355 ( P1_U7139 , P1_U2574 , P1_INSTQUEUE_REG_15__4_ );
nand NAND2_17356 ( P1_U7140 , P1_U2572 , P1_INSTQUEUE_REG_1__4_ );
nand NAND2_17357 ( P1_U7141 , P1_U2571 , P1_INSTQUEUE_REG_2__4_ );
nand NAND2_17358 ( P1_U7142 , P1_U2570 , P1_INSTQUEUE_REG_3__4_ );
nand NAND2_17359 ( P1_U7143 , P1_U2568 , P1_INSTQUEUE_REG_4__4_ );
nand NAND2_17360 ( P1_U7144 , P1_U2567 , P1_INSTQUEUE_REG_5__4_ );
nand NAND2_17361 ( P1_U7145 , P1_U2566 , P1_INSTQUEUE_REG_6__4_ );
nand NAND2_17362 ( P1_U7146 , P1_U2565 , P1_INSTQUEUE_REG_7__4_ );
nand NAND2_17363 ( P1_U7147 , P1_U2582 , P1_INSTQUEUE_REG_8__3_ );
nand NAND2_17364 ( P1_U7148 , P1_U2581 , P1_INSTQUEUE_REG_9__3_ );
nand NAND2_17365 ( P1_U7149 , P1_U2580 , P1_INSTQUEUE_REG_10__3_ );
nand NAND2_17366 ( P1_U7150 , P1_U2579 , P1_INSTQUEUE_REG_11__3_ );
nand NAND2_17367 ( P1_U7151 , P1_U2577 , P1_INSTQUEUE_REG_12__3_ );
nand NAND2_17368 ( P1_U7152 , P1_U2576 , P1_INSTQUEUE_REG_13__3_ );
nand NAND2_17369 ( P1_U7153 , P1_U2575 , P1_INSTQUEUE_REG_14__3_ );
nand NAND2_17370 ( P1_U7154 , P1_U2574 , P1_INSTQUEUE_REG_15__3_ );
nand NAND2_17371 ( P1_U7155 , P1_U2573 , P1_INSTQUEUE_REG_0__3_ );
nand NAND2_17372 ( P1_U7156 , P1_U2572 , P1_INSTQUEUE_REG_1__3_ );
nand NAND2_17373 ( P1_U7157 , P1_U2571 , P1_INSTQUEUE_REG_2__3_ );
nand NAND2_17374 ( P1_U7158 , P1_U2570 , P1_INSTQUEUE_REG_3__3_ );
nand NAND2_17375 ( P1_U7159 , P1_U2568 , P1_INSTQUEUE_REG_4__3_ );
nand NAND2_17376 ( P1_U7160 , P1_U2567 , P1_INSTQUEUE_REG_5__3_ );
nand NAND2_17377 ( P1_U7161 , P1_U2566 , P1_INSTQUEUE_REG_6__3_ );
nand NAND2_17378 ( P1_U7162 , P1_U2565 , P1_INSTQUEUE_REG_7__3_ );
nand NAND4_17379 ( P1_U7163 , P1_U4095 , P1_U4094 , P1_U4093 , P1_U4092 );
nand NAND2_17380 ( P1_U7164 , P1_U2582 , P1_INSTQUEUE_REG_8__2_ );
nand NAND2_17381 ( P1_U7165 , P1_U2581 , P1_INSTQUEUE_REG_9__2_ );
nand NAND2_17382 ( P1_U7166 , P1_U2580 , P1_INSTQUEUE_REG_10__2_ );
nand NAND2_17383 ( P1_U7167 , P1_U2579 , P1_INSTQUEUE_REG_11__2_ );
nand NAND2_17384 ( P1_U7168 , P1_U2577 , P1_INSTQUEUE_REG_12__2_ );
nand NAND2_17385 ( P1_U7169 , P1_U2576 , P1_INSTQUEUE_REG_13__2_ );
nand NAND2_17386 ( P1_U7170 , P1_U2575 , P1_INSTQUEUE_REG_14__2_ );
nand NAND2_17387 ( P1_U7171 , P1_U2574 , P1_INSTQUEUE_REG_15__2_ );
nand NAND2_17388 ( P1_U7172 , P1_U2573 , P1_INSTQUEUE_REG_0__2_ );
nand NAND2_17389 ( P1_U7173 , P1_U2572 , P1_INSTQUEUE_REG_1__2_ );
nand NAND2_17390 ( P1_U7174 , P1_U2571 , P1_INSTQUEUE_REG_2__2_ );
nand NAND2_17391 ( P1_U7175 , P1_U2570 , P1_INSTQUEUE_REG_3__2_ );
nand NAND2_17392 ( P1_U7176 , P1_U2568 , P1_INSTQUEUE_REG_4__2_ );
nand NAND2_17393 ( P1_U7177 , P1_U2567 , P1_INSTQUEUE_REG_5__2_ );
nand NAND2_17394 ( P1_U7178 , P1_U2566 , P1_INSTQUEUE_REG_6__2_ );
nand NAND2_17395 ( P1_U7179 , P1_U2565 , P1_INSTQUEUE_REG_7__2_ );
nand NAND4_17396 ( P1_U7180 , P1_U4099 , P1_U4098 , P1_U4097 , P1_U4096 );
nand NAND2_17397 ( P1_U7181 , P1_U2582 , P1_INSTQUEUE_REG_8__1_ );
nand NAND2_17398 ( P1_U7182 , P1_U2581 , P1_INSTQUEUE_REG_9__1_ );
nand NAND2_17399 ( P1_U7183 , P1_U2580 , P1_INSTQUEUE_REG_10__1_ );
nand NAND2_17400 ( P1_U7184 , P1_U2579 , P1_INSTQUEUE_REG_11__1_ );
nand NAND2_17401 ( P1_U7185 , P1_U2577 , P1_INSTQUEUE_REG_12__1_ );
nand NAND2_17402 ( P1_U7186 , P1_U2576 , P1_INSTQUEUE_REG_13__1_ );
nand NAND2_17403 ( P1_U7187 , P1_U2575 , P1_INSTQUEUE_REG_14__1_ );
nand NAND2_17404 ( P1_U7188 , P1_U2574 , P1_INSTQUEUE_REG_15__1_ );
nand NAND2_17405 ( P1_U7189 , P1_U2573 , P1_INSTQUEUE_REG_0__1_ );
nand NAND2_17406 ( P1_U7190 , P1_U2572 , P1_INSTQUEUE_REG_1__1_ );
nand NAND2_17407 ( P1_U7191 , P1_U2571 , P1_INSTQUEUE_REG_2__1_ );
nand NAND2_17408 ( P1_U7192 , P1_U2570 , P1_INSTQUEUE_REG_3__1_ );
nand NAND2_17409 ( P1_U7193 , P1_U2568 , P1_INSTQUEUE_REG_4__1_ );
nand NAND2_17410 ( P1_U7194 , P1_U2567 , P1_INSTQUEUE_REG_5__1_ );
nand NAND2_17411 ( P1_U7195 , P1_U2566 , P1_INSTQUEUE_REG_6__1_ );
nand NAND2_17412 ( P1_U7196 , P1_U2565 , P1_INSTQUEUE_REG_7__1_ );
nand NAND4_17413 ( P1_U7197 , P1_U4103 , P1_U4102 , P1_U4101 , P1_U4100 );
nand NAND2_17414 ( P1_U7198 , P1_U2582 , P1_INSTQUEUE_REG_8__0_ );
nand NAND2_17415 ( P1_U7199 , P1_U2581 , P1_INSTQUEUE_REG_9__0_ );
nand NAND2_17416 ( P1_U7200 , P1_U2580 , P1_INSTQUEUE_REG_10__0_ );
nand NAND2_17417 ( P1_U7201 , P1_U2579 , P1_INSTQUEUE_REG_11__0_ );
nand NAND2_17418 ( P1_U7202 , P1_U2577 , P1_INSTQUEUE_REG_12__0_ );
nand NAND2_17419 ( P1_U7203 , P1_U2576 , P1_INSTQUEUE_REG_13__0_ );
nand NAND2_17420 ( P1_U7204 , P1_U2575 , P1_INSTQUEUE_REG_14__0_ );
nand NAND2_17421 ( P1_U7205 , P1_U2574 , P1_INSTQUEUE_REG_15__0_ );
nand NAND2_17422 ( P1_U7206 , P1_U2573 , P1_INSTQUEUE_REG_0__0_ );
nand NAND2_17423 ( P1_U7207 , P1_U2572 , P1_INSTQUEUE_REG_1__0_ );
nand NAND2_17424 ( P1_U7208 , P1_U2571 , P1_INSTQUEUE_REG_2__0_ );
nand NAND2_17425 ( P1_U7209 , P1_U2570 , P1_INSTQUEUE_REG_3__0_ );
nand NAND2_17426 ( P1_U7210 , P1_U2568 , P1_INSTQUEUE_REG_4__0_ );
nand NAND2_17427 ( P1_U7211 , P1_U2567 , P1_INSTQUEUE_REG_5__0_ );
nand NAND2_17428 ( P1_U7212 , P1_U2566 , P1_INSTQUEUE_REG_6__0_ );
nand NAND2_17429 ( P1_U7213 , P1_U2565 , P1_INSTQUEUE_REG_7__0_ );
nand NAND4_17430 ( P1_U7214 , P1_U4107 , P1_U4106 , P1_U4105 , P1_U4104 );
nand NAND2_17431 ( P1_U7215 , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_U3297 );
nand NAND2_17432 ( P1_U7216 , P1_U4203 , P1_U3455 );
nand NAND2_17433 ( P1_U7217 , P1_INSTQUEUEWR_ADDR_REG_1_ , P1_U3297 );
nand NAND2_17434 ( P1_U7218 , P1_U4203 , P1_U3235 );
not NOT1_17435 ( P1_U7219 , P1_U4183 );
nand NAND2_17436 ( P1_U7220 , P1_U2602 , P1_INSTQUEUE_REG_8__7_ );
nand NAND2_17437 ( P1_U7221 , P1_U2601 , P1_INSTQUEUE_REG_9__7_ );
nand NAND2_17438 ( P1_U7222 , P1_U2600 , P1_INSTQUEUE_REG_10__7_ );
nand NAND2_17439 ( P1_U7223 , P1_U2599 , P1_INSTQUEUE_REG_11__7_ );
nand NAND2_17440 ( P1_U7224 , P1_U2597 , P1_INSTQUEUE_REG_12__7_ );
nand NAND2_17441 ( P1_U7225 , P1_U2596 , P1_INSTQUEUE_REG_13__7_ );
nand NAND2_17442 ( P1_U7226 , P1_U2595 , P1_INSTQUEUE_REG_14__7_ );
nand NAND2_17443 ( P1_U7227 , P1_U2594 , P1_INSTQUEUE_REG_15__7_ );
nand NAND2_17444 ( P1_U7228 , P1_U2592 , P1_INSTQUEUE_REG_0__7_ );
nand NAND2_17445 ( P1_U7229 , P1_U2591 , P1_INSTQUEUE_REG_1__7_ );
nand NAND2_17446 ( P1_U7230 , P1_U2590 , P1_INSTQUEUE_REG_2__7_ );
nand NAND2_17447 ( P1_U7231 , P1_U2589 , P1_INSTQUEUE_REG_3__7_ );
nand NAND2_17448 ( P1_U7232 , P1_U2587 , P1_INSTQUEUE_REG_4__7_ );
nand NAND2_17449 ( P1_U7233 , P1_U2586 , P1_INSTQUEUE_REG_5__7_ );
nand NAND2_17450 ( P1_U7234 , P1_U2585 , P1_INSTQUEUE_REG_6__7_ );
nand NAND2_17451 ( P1_U7235 , P1_U2584 , P1_INSTQUEUE_REG_7__7_ );
nand NAND4_17452 ( P1_U7236 , P1_U4124 , P1_U4123 , P1_U4122 , P1_U4121 );
nand NAND2_17453 ( P1_U7237 , P1_U2602 , P1_INSTQUEUE_REG_8__6_ );
nand NAND2_17454 ( P1_U7238 , P1_U2601 , P1_INSTQUEUE_REG_9__6_ );
nand NAND2_17455 ( P1_U7239 , P1_U2600 , P1_INSTQUEUE_REG_10__6_ );
nand NAND2_17456 ( P1_U7240 , P1_U2599 , P1_INSTQUEUE_REG_11__6_ );
nand NAND2_17457 ( P1_U7241 , P1_U2597 , P1_INSTQUEUE_REG_12__6_ );
nand NAND2_17458 ( P1_U7242 , P1_U2596 , P1_INSTQUEUE_REG_13__6_ );
nand NAND2_17459 ( P1_U7243 , P1_U2595 , P1_INSTQUEUE_REG_14__6_ );
nand NAND2_17460 ( P1_U7244 , P1_U2594 , P1_INSTQUEUE_REG_15__6_ );
nand NAND2_17461 ( P1_U7245 , P1_U2592 , P1_INSTQUEUE_REG_0__6_ );
nand NAND2_17462 ( P1_U7246 , P1_U2591 , P1_INSTQUEUE_REG_1__6_ );
nand NAND2_17463 ( P1_U7247 , P1_U2590 , P1_INSTQUEUE_REG_2__6_ );
nand NAND2_17464 ( P1_U7248 , P1_U2589 , P1_INSTQUEUE_REG_3__6_ );
nand NAND2_17465 ( P1_U7249 , P1_U2587 , P1_INSTQUEUE_REG_4__6_ );
nand NAND2_17466 ( P1_U7250 , P1_U2586 , P1_INSTQUEUE_REG_5__6_ );
nand NAND2_17467 ( P1_U7251 , P1_U2585 , P1_INSTQUEUE_REG_6__6_ );
nand NAND2_17468 ( P1_U7252 , P1_U2584 , P1_INSTQUEUE_REG_7__6_ );
nand NAND4_17469 ( P1_U7253 , P1_U4128 , P1_U4127 , P1_U4126 , P1_U4125 );
nand NAND2_17470 ( P1_U7254 , P1_U2602 , P1_INSTQUEUE_REG_8__5_ );
nand NAND2_17471 ( P1_U7255 , P1_U2601 , P1_INSTQUEUE_REG_9__5_ );
nand NAND2_17472 ( P1_U7256 , P1_U2600 , P1_INSTQUEUE_REG_10__5_ );
nand NAND2_17473 ( P1_U7257 , P1_U2599 , P1_INSTQUEUE_REG_11__5_ );
nand NAND2_17474 ( P1_U7258 , P1_U2597 , P1_INSTQUEUE_REG_12__5_ );
nand NAND2_17475 ( P1_U7259 , P1_U2596 , P1_INSTQUEUE_REG_13__5_ );
nand NAND2_17476 ( P1_U7260 , P1_U2595 , P1_INSTQUEUE_REG_14__5_ );
nand NAND2_17477 ( P1_U7261 , P1_U2594 , P1_INSTQUEUE_REG_15__5_ );
nand NAND2_17478 ( P1_U7262 , P1_U2592 , P1_INSTQUEUE_REG_0__5_ );
nand NAND2_17479 ( P1_U7263 , P1_U2591 , P1_INSTQUEUE_REG_1__5_ );
nand NAND2_17480 ( P1_U7264 , P1_U2590 , P1_INSTQUEUE_REG_2__5_ );
nand NAND2_17481 ( P1_U7265 , P1_U2589 , P1_INSTQUEUE_REG_3__5_ );
nand NAND2_17482 ( P1_U7266 , P1_U2587 , P1_INSTQUEUE_REG_4__5_ );
nand NAND2_17483 ( P1_U7267 , P1_U2586 , P1_INSTQUEUE_REG_5__5_ );
nand NAND2_17484 ( P1_U7268 , P1_U2585 , P1_INSTQUEUE_REG_6__5_ );
nand NAND2_17485 ( P1_U7269 , P1_U2584 , P1_INSTQUEUE_REG_7__5_ );
nand NAND4_17486 ( P1_U7270 , P1_U4132 , P1_U4131 , P1_U4130 , P1_U4129 );
nand NAND2_17487 ( P1_U7271 , P1_U2602 , P1_INSTQUEUE_REG_8__4_ );
nand NAND2_17488 ( P1_U7272 , P1_U2601 , P1_INSTQUEUE_REG_9__4_ );
nand NAND2_17489 ( P1_U7273 , P1_U2600 , P1_INSTQUEUE_REG_10__4_ );
nand NAND2_17490 ( P1_U7274 , P1_U2599 , P1_INSTQUEUE_REG_11__4_ );
nand NAND2_17491 ( P1_U7275 , P1_U2597 , P1_INSTQUEUE_REG_12__4_ );
nand NAND2_17492 ( P1_U7276 , P1_U2596 , P1_INSTQUEUE_REG_13__4_ );
nand NAND2_17493 ( P1_U7277 , P1_U2595 , P1_INSTQUEUE_REG_14__4_ );
nand NAND2_17494 ( P1_U7278 , P1_U2594 , P1_INSTQUEUE_REG_15__4_ );
nand NAND2_17495 ( P1_U7279 , P1_U2591 , P1_INSTQUEUE_REG_1__4_ );
nand NAND2_17496 ( P1_U7280 , P1_U2590 , P1_INSTQUEUE_REG_2__4_ );
nand NAND2_17497 ( P1_U7281 , P1_U2589 , P1_INSTQUEUE_REG_3__4_ );
nand NAND2_17498 ( P1_U7282 , P1_U2587 , P1_INSTQUEUE_REG_4__4_ );
nand NAND2_17499 ( P1_U7283 , P1_U2586 , P1_INSTQUEUE_REG_5__4_ );
nand NAND2_17500 ( P1_U7284 , P1_U2585 , P1_INSTQUEUE_REG_6__4_ );
nand NAND2_17501 ( P1_U7285 , P1_U2584 , P1_INSTQUEUE_REG_7__4_ );
nand NAND2_17502 ( P1_U7286 , P1_U2602 , P1_INSTQUEUE_REG_8__3_ );
nand NAND2_17503 ( P1_U7287 , P1_U2601 , P1_INSTQUEUE_REG_9__3_ );
nand NAND2_17504 ( P1_U7288 , P1_U2600 , P1_INSTQUEUE_REG_10__3_ );
nand NAND2_17505 ( P1_U7289 , P1_U2599 , P1_INSTQUEUE_REG_11__3_ );
nand NAND2_17506 ( P1_U7290 , P1_U2597 , P1_INSTQUEUE_REG_12__3_ );
nand NAND2_17507 ( P1_U7291 , P1_U2596 , P1_INSTQUEUE_REG_13__3_ );
nand NAND2_17508 ( P1_U7292 , P1_U2595 , P1_INSTQUEUE_REG_14__3_ );
nand NAND2_17509 ( P1_U7293 , P1_U2594 , P1_INSTQUEUE_REG_15__3_ );
nand NAND2_17510 ( P1_U7294 , P1_U2592 , P1_INSTQUEUE_REG_0__3_ );
nand NAND2_17511 ( P1_U7295 , P1_U2591 , P1_INSTQUEUE_REG_1__3_ );
nand NAND2_17512 ( P1_U7296 , P1_U2590 , P1_INSTQUEUE_REG_2__3_ );
nand NAND2_17513 ( P1_U7297 , P1_U2589 , P1_INSTQUEUE_REG_3__3_ );
nand NAND2_17514 ( P1_U7298 , P1_U2587 , P1_INSTQUEUE_REG_4__3_ );
nand NAND2_17515 ( P1_U7299 , P1_U2586 , P1_INSTQUEUE_REG_5__3_ );
nand NAND2_17516 ( P1_U7300 , P1_U2585 , P1_INSTQUEUE_REG_6__3_ );
nand NAND2_17517 ( P1_U7301 , P1_U2584 , P1_INSTQUEUE_REG_7__3_ );
nand NAND4_17518 ( P1_U7302 , P1_U4140 , P1_U4139 , P1_U4138 , P1_U4137 );
nand NAND2_17519 ( P1_U7303 , P1_U2602 , P1_INSTQUEUE_REG_8__2_ );
nand NAND2_17520 ( P1_U7304 , P1_U2601 , P1_INSTQUEUE_REG_9__2_ );
nand NAND2_17521 ( P1_U7305 , P1_U2600 , P1_INSTQUEUE_REG_10__2_ );
nand NAND2_17522 ( P1_U7306 , P1_U2599 , P1_INSTQUEUE_REG_11__2_ );
nand NAND2_17523 ( P1_U7307 , P1_U2597 , P1_INSTQUEUE_REG_12__2_ );
nand NAND2_17524 ( P1_U7308 , P1_U2596 , P1_INSTQUEUE_REG_13__2_ );
nand NAND2_17525 ( P1_U7309 , P1_U2595 , P1_INSTQUEUE_REG_14__2_ );
nand NAND2_17526 ( P1_U7310 , P1_U2594 , P1_INSTQUEUE_REG_15__2_ );
nand NAND2_17527 ( P1_U7311 , P1_U2592 , P1_INSTQUEUE_REG_0__2_ );
nand NAND2_17528 ( P1_U7312 , P1_U2591 , P1_INSTQUEUE_REG_1__2_ );
nand NAND2_17529 ( P1_U7313 , P1_U2590 , P1_INSTQUEUE_REG_2__2_ );
nand NAND2_17530 ( P1_U7314 , P1_U2589 , P1_INSTQUEUE_REG_3__2_ );
nand NAND2_17531 ( P1_U7315 , P1_U2587 , P1_INSTQUEUE_REG_4__2_ );
nand NAND2_17532 ( P1_U7316 , P1_U2586 , P1_INSTQUEUE_REG_5__2_ );
nand NAND2_17533 ( P1_U7317 , P1_U2585 , P1_INSTQUEUE_REG_6__2_ );
nand NAND2_17534 ( P1_U7318 , P1_U2584 , P1_INSTQUEUE_REG_7__2_ );
nand NAND4_17535 ( P1_U7319 , P1_U4144 , P1_U4143 , P1_U4142 , P1_U4141 );
nand NAND2_17536 ( P1_U7320 , P1_U2602 , P1_INSTQUEUE_REG_8__1_ );
nand NAND2_17537 ( P1_U7321 , P1_U2601 , P1_INSTQUEUE_REG_9__1_ );
nand NAND2_17538 ( P1_U7322 , P1_U2600 , P1_INSTQUEUE_REG_10__1_ );
nand NAND2_17539 ( P1_U7323 , P1_U2599 , P1_INSTQUEUE_REG_11__1_ );
nand NAND2_17540 ( P1_U7324 , P1_U2597 , P1_INSTQUEUE_REG_12__1_ );
nand NAND2_17541 ( P1_U7325 , P1_U2596 , P1_INSTQUEUE_REG_13__1_ );
nand NAND2_17542 ( P1_U7326 , P1_U2595 , P1_INSTQUEUE_REG_14__1_ );
nand NAND2_17543 ( P1_U7327 , P1_U2594 , P1_INSTQUEUE_REG_15__1_ );
nand NAND2_17544 ( P1_U7328 , P1_U2592 , P1_INSTQUEUE_REG_0__1_ );
nand NAND2_17545 ( P1_U7329 , P1_U2591 , P1_INSTQUEUE_REG_1__1_ );
nand NAND2_17546 ( P1_U7330 , P1_U2590 , P1_INSTQUEUE_REG_2__1_ );
nand NAND2_17547 ( P1_U7331 , P1_U2589 , P1_INSTQUEUE_REG_3__1_ );
nand NAND2_17548 ( P1_U7332 , P1_U2587 , P1_INSTQUEUE_REG_4__1_ );
nand NAND2_17549 ( P1_U7333 , P1_U2586 , P1_INSTQUEUE_REG_5__1_ );
nand NAND2_17550 ( P1_U7334 , P1_U2585 , P1_INSTQUEUE_REG_6__1_ );
nand NAND2_17551 ( P1_U7335 , P1_U2584 , P1_INSTQUEUE_REG_7__1_ );
nand NAND4_17552 ( P1_U7336 , P1_U4148 , P1_U4147 , P1_U4146 , P1_U4145 );
nand NAND2_17553 ( P1_U7337 , P1_U2602 , P1_INSTQUEUE_REG_8__0_ );
nand NAND2_17554 ( P1_U7338 , P1_U2601 , P1_INSTQUEUE_REG_9__0_ );
nand NAND2_17555 ( P1_U7339 , P1_U2600 , P1_INSTQUEUE_REG_10__0_ );
nand NAND2_17556 ( P1_U7340 , P1_U2599 , P1_INSTQUEUE_REG_11__0_ );
nand NAND2_17557 ( P1_U7341 , P1_U2597 , P1_INSTQUEUE_REG_12__0_ );
nand NAND2_17558 ( P1_U7342 , P1_U2596 , P1_INSTQUEUE_REG_13__0_ );
nand NAND2_17559 ( P1_U7343 , P1_U2595 , P1_INSTQUEUE_REG_14__0_ );
nand NAND2_17560 ( P1_U7344 , P1_U2594 , P1_INSTQUEUE_REG_15__0_ );
nand NAND2_17561 ( P1_U7345 , P1_U2592 , P1_INSTQUEUE_REG_0__0_ );
nand NAND2_17562 ( P1_U7346 , P1_U2591 , P1_INSTQUEUE_REG_1__0_ );
nand NAND2_17563 ( P1_U7347 , P1_U2590 , P1_INSTQUEUE_REG_2__0_ );
nand NAND2_17564 ( P1_U7348 , P1_U2589 , P1_INSTQUEUE_REG_3__0_ );
nand NAND2_17565 ( P1_U7349 , P1_U2587 , P1_INSTQUEUE_REG_4__0_ );
nand NAND2_17566 ( P1_U7350 , P1_U2586 , P1_INSTQUEUE_REG_5__0_ );
nand NAND2_17567 ( P1_U7351 , P1_U2585 , P1_INSTQUEUE_REG_6__0_ );
nand NAND2_17568 ( P1_U7352 , P1_U2584 , P1_INSTQUEUE_REG_7__0_ );
nand NAND4_17569 ( P1_U7353 , P1_U4152 , P1_U4151 , P1_U4150 , P1_U4149 );
nand NAND3_17570 ( P1_U7354 , P1_U4231 , P1_U2354 , P1_U4234 );
nand NAND2_17571 ( P1_U7355 , P1_U4153 , P1_U7087 );
nand NAND2_17572 ( P1_U7356 , P1_U3396 , P1_U3410 );
nand NAND2_17573 ( P1_U7357 , P1_U4234 , P1_U7356 );
nand NAND2_17574 ( P1_U7358 , P1_U4190 , P1_U2452 );
nand NAND2_17575 ( P1_U7359 , P1_U7355 , P1_U3271 );
nand NAND2_17576 ( P1_U7360 , P1_U4208 , P1_U7088 );
nand NAND2_17577 ( P1_U7361 , P1_U4160 , P1_U4208 );
nand NAND2_17578 ( P1_U7362 , P1_U2451 , P1_U4210 );
nand NAND5_17579 ( P1_U7363 , P1_U3420 , P1_U3434 , P1_U4195 , P1_U7362 , P1_U7361 );
nand NAND2_17580 ( P1_U7364 , P1_R2238_U6 , P1_U7363 );
nand NAND2_17581 ( P1_U7365 , P1_SUB_450_U6 , P1_U2354 );
nand NAND2_17582 ( P1_U7366 , P1_R2238_U19 , P1_U7363 );
nand NAND2_17583 ( P1_U7367 , P1_SUB_450_U19 , P1_U2354 );
nand NAND2_17584 ( P1_U7368 , P1_R2238_U20 , P1_U7363 );
nand NAND2_17585 ( P1_U7369 , P1_SUB_450_U20 , P1_U2354 );
nand NAND2_17586 ( P1_U7370 , P1_R2238_U21 , P1_U7363 );
nand NAND2_17587 ( P1_U7371 , P1_SUB_450_U21 , P1_U2354 );
nand NAND2_17588 ( P1_U7372 , P1_R2238_U22 , P1_U7363 );
nand NAND2_17589 ( P1_U7373 , P1_SUB_450_U22 , P1_U2354 );
nand NAND2_17590 ( P1_U7374 , P1_R2238_U7 , P1_U7363 );
nand NAND2_17591 ( P1_U7375 , P1_SUB_450_U7 , P1_U2354 );
nand NAND2_17592 ( P1_U7376 , P1_R2238_U19 , P1_U4192 );
nand NAND2_17593 ( P1_U7377 , P1_INSTQUEUERD_ADDR_REG_4_ , P1_U3294 );
nand NAND2_17594 ( P1_U7378 , P1_R2238_U20 , P1_U4192 );
nand NAND2_17595 ( P1_U7379 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_U3294 );
nand NAND2_17596 ( P1_U7380 , P1_STATE2_REG_0_ , P1_U4173 );
nand NAND2_17597 ( P1_U7381 , P1_U3420 , P1_U7380 );
nand NAND2_17598 ( P1_U7382 , P1_R2238_U21 , P1_U4192 );
nand NAND2_17599 ( P1_U7383 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3294 );
nand NAND2_17600 ( P1_U7384 , P1_U2450 , P1_U3271 );
nand NAND2_17601 ( P1_U7385 , P1_R2238_U22 , P1_U4192 );
nand NAND2_17602 ( P1_U7386 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3294 );
nand NAND2_17603 ( P1_U7387 , P1_U2451 , P1_U3284 );
nand NAND2_17604 ( P1_U7388 , P1_R2238_U7 , P1_U4192 );
nand NAND2_17605 ( P1_U7389 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_U3294 );
nand NAND2_17606 ( P1_U7390 , P1_U3393 , P1_U3290 );
nand NAND2_17607 ( P1_U7391 , P1_U3284 , P1_U3449 );
nand NAND2_17608 ( P1_U7392 , P1_INSTADDRPOINTER_REG_9_ , P1_U7391 );
nand NAND2_17609 ( P1_U7393 , P1_EBX_REG_9_ , P1_U7390 );
nand NAND2_17610 ( P1_U7394 , P1_INSTADDRPOINTER_REG_8_ , P1_U7391 );
nand NAND2_17611 ( P1_U7395 , P1_EBX_REG_8_ , P1_U7390 );
nand NAND2_17612 ( P1_U7396 , P1_INSTADDRPOINTER_REG_7_ , P1_U7391 );
nand NAND2_17613 ( P1_U7397 , P1_EBX_REG_7_ , P1_U7390 );
nand NAND2_17614 ( P1_U7398 , P1_INSTADDRPOINTER_REG_6_ , P1_U7391 );
nand NAND2_17615 ( P1_U7399 , P1_EBX_REG_6_ , P1_U7390 );
nand NAND2_17616 ( P1_U7400 , P1_INSTADDRPOINTER_REG_5_ , P1_U7391 );
nand NAND2_17617 ( P1_U7401 , P1_EBX_REG_5_ , P1_U7390 );
nand NAND2_17618 ( P1_U7402 , P1_INSTADDRPOINTER_REG_4_ , P1_U7391 );
nand NAND2_17619 ( P1_U7403 , P1_EBX_REG_4_ , P1_U7390 );
nand NAND2_17620 ( P1_U7404 , P1_INSTADDRPOINTER_REG_31_ , P1_U7391 );
nand NAND2_17621 ( P1_U7405 , P1_EBX_REG_31_ , P1_U7390 );
nand NAND2_17622 ( P1_U7406 , P1_INSTADDRPOINTER_REG_30_ , P1_U7391 );
nand NAND2_17623 ( P1_U7407 , P1_EBX_REG_30_ , P1_U7390 );
nand NAND2_17624 ( P1_U7408 , P1_INSTADDRPOINTER_REG_3_ , P1_U7391 );
nand NAND2_17625 ( P1_U7409 , P1_EBX_REG_3_ , P1_U7390 );
nand NAND2_17626 ( P1_U7410 , P1_INSTADDRPOINTER_REG_29_ , P1_U7391 );
nand NAND2_17627 ( P1_U7411 , P1_EBX_REG_29_ , P1_U7390 );
nand NAND2_17628 ( P1_U7412 , P1_INSTADDRPOINTER_REG_28_ , P1_U7391 );
nand NAND2_17629 ( P1_U7413 , P1_EBX_REG_28_ , P1_U7390 );
nand NAND2_17630 ( P1_U7414 , P1_INSTADDRPOINTER_REG_27_ , P1_U7391 );
nand NAND2_17631 ( P1_U7415 , P1_EBX_REG_27_ , P1_U7390 );
nand NAND2_17632 ( P1_U7416 , P1_INSTADDRPOINTER_REG_26_ , P1_U7391 );
nand NAND2_17633 ( P1_U7417 , P1_EBX_REG_26_ , P1_U7390 );
nand NAND2_17634 ( P1_U7418 , P1_INSTADDRPOINTER_REG_25_ , P1_U7391 );
nand NAND2_17635 ( P1_U7419 , P1_EBX_REG_25_ , P1_U7390 );
nand NAND2_17636 ( P1_U7420 , P1_INSTADDRPOINTER_REG_24_ , P1_U7391 );
nand NAND2_17637 ( P1_U7421 , P1_EBX_REG_24_ , P1_U7390 );
nand NAND2_17638 ( P1_U7422 , P1_INSTADDRPOINTER_REG_23_ , P1_U7391 );
nand NAND2_17639 ( P1_U7423 , P1_EBX_REG_23_ , P1_U7390 );
nand NAND2_17640 ( P1_U7424 , P1_INSTADDRPOINTER_REG_22_ , P1_U7391 );
nand NAND2_17641 ( P1_U7425 , P1_EBX_REG_22_ , P1_U7390 );
nand NAND2_17642 ( P1_U7426 , P1_INSTADDRPOINTER_REG_21_ , P1_U7391 );
nand NAND2_17643 ( P1_U7427 , P1_EBX_REG_21_ , P1_U7390 );
nand NAND2_17644 ( P1_U7428 , P1_INSTADDRPOINTER_REG_20_ , P1_U7391 );
nand NAND2_17645 ( P1_U7429 , P1_EBX_REG_20_ , P1_U7390 );
nand NAND2_17646 ( P1_U7430 , P1_INSTADDRPOINTER_REG_2_ , P1_U7391 );
nand NAND2_17647 ( P1_U7431 , P1_EBX_REG_2_ , P1_U7390 );
nand NAND2_17648 ( P1_U7432 , P1_INSTADDRPOINTER_REG_19_ , P1_U7391 );
nand NAND2_17649 ( P1_U7433 , P1_EBX_REG_19_ , P1_U7390 );
nand NAND2_17650 ( P1_U7434 , P1_INSTADDRPOINTER_REG_18_ , P1_U7391 );
nand NAND2_17651 ( P1_U7435 , P1_EBX_REG_18_ , P1_U7390 );
nand NAND2_17652 ( P1_U7436 , P1_INSTADDRPOINTER_REG_17_ , P1_U7391 );
nand NAND2_17653 ( P1_U7437 , P1_EBX_REG_17_ , P1_U7390 );
nand NAND2_17654 ( P1_U7438 , P1_INSTADDRPOINTER_REG_16_ , P1_U7391 );
nand NAND2_17655 ( P1_U7439 , P1_EBX_REG_16_ , P1_U7390 );
nand NAND2_17656 ( P1_U7440 , P1_INSTADDRPOINTER_REG_15_ , P1_U7391 );
nand NAND2_17657 ( P1_U7441 , P1_EBX_REG_15_ , P1_U7390 );
nand NAND2_17658 ( P1_U7442 , P1_INSTADDRPOINTER_REG_14_ , P1_U7391 );
nand NAND2_17659 ( P1_U7443 , P1_EBX_REG_14_ , P1_U7390 );
nand NAND2_17660 ( P1_U7444 , P1_INSTADDRPOINTER_REG_13_ , P1_U7391 );
nand NAND2_17661 ( P1_U7445 , P1_EBX_REG_13_ , P1_U7390 );
nand NAND2_17662 ( P1_U7446 , P1_INSTADDRPOINTER_REG_12_ , P1_U7391 );
nand NAND2_17663 ( P1_U7447 , P1_EBX_REG_12_ , P1_U7390 );
nand NAND2_17664 ( P1_U7448 , P1_INSTADDRPOINTER_REG_11_ , P1_U7391 );
nand NAND2_17665 ( P1_U7449 , P1_EBX_REG_11_ , P1_U7390 );
nand NAND2_17666 ( P1_U7450 , P1_INSTADDRPOINTER_REG_10_ , P1_U7391 );
nand NAND2_17667 ( P1_U7451 , P1_EBX_REG_10_ , P1_U7390 );
nand NAND2_17668 ( P1_U7452 , P1_INSTADDRPOINTER_REG_1_ , P1_U7391 );
nand NAND2_17669 ( P1_U7453 , P1_EBX_REG_1_ , P1_U7390 );
nand NAND2_17670 ( P1_U7454 , P1_INSTADDRPOINTER_REG_0_ , P1_U7391 );
nand NAND2_17671 ( P1_U7455 , P1_EBX_REG_0_ , P1_U7390 );
nand NAND2_17672 ( P1_U7456 , P1_U4477 , P1_U4496 );
nand NAND2_17673 ( P1_U7457 , P1_U2430 , P1_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_17674 ( P1_U7458 , P1_U3489 , P1_U3262 );
nand NAND2_17675 ( P1_U7459 , P1_U2430 , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_17676 ( P1_U7460 , P1_U3490 , P1_U3262 );
nand NAND3_17677 ( P1_U7461 , P1_FLUSH_REG , P1_U2446 , P1_U3470 );
nand NAND2_17678 ( P1_U7462 , P1_U2430 , P1_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_17679 ( P1_U7463 , P1_U3491 , P1_U3262 );
nand NAND3_17680 ( P1_U7464 , P1_U2446 , P1_FLUSH_REG , P1_U7712 );
nand NAND2_17681 ( P1_U7465 , P1_U2430 , P1_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_17682 ( P1_U7466 , P1_U3492 , P1_U3262 );
nand NAND2_17683 ( P1_U7467 , P1_U2430 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_17684 ( P1_U7468 , P1_STATE_REG_0_ , P1_U4185 );
or OR2_17685 ( P1_U7469 , U210 , P1_STATE2_REG_2_ );
nand NAND2_17686 ( P1_U7470 , P1_U4110 , P1_U7218 );
nand NAND2_17687 ( P1_U7471 , P1_U7084 , P1_U3422 );
nand NAND2_17688 ( P1_U7472 , P1_U4211 , P1_STATE2_REG_0_ );
nand NAND2_17689 ( P1_U7473 , P1_U4212 , P1_STATE2_REG_0_ );
nand NAND2_17690 ( P1_U7474 , P1_U4213 , P1_STATE2_REG_0_ );
nand NAND2_17691 ( P1_U7475 , P1_U4236 , P1_STATE2_REG_0_ );
nand NAND2_17692 ( P1_U7476 , P1_U4264 , P1_STATE2_REG_0_ );
nand NAND2_17693 ( P1_U7477 , P1_STATE2_REG_0_ , P1_U7632 );
nand NAND2_17694 ( P1_U7478 , P1_U2608 , P1_U3266 );
nand NAND4_17695 ( P1_U7479 , P1_U4117 , P1_U7093 , P1_U4118 , P1_U4120 );
nand NAND2_17696 ( P1_U7480 , P1_STATE2_REG_0_ , P1_U7632 );
nand NAND2_17697 ( P1_U7481 , P1_U2379 , P1_U3429 );
nand NAND2_17698 ( P1_U7482 , P1_U2369 , P1_U6367 );
nand NAND2_17699 ( P1_U7483 , P1_U3888 , P1_U2369 );
nand NAND3_17700 ( P1_U7484 , P1_U7481 , P1_U4229 , P1_U7482 );
nand NAND2_17701 ( P1_U7485 , P1_U7483 , P1_U4230 );
nand NAND3_17702 ( P1_U7486 , P1_U5491 , P1_U4171 , P1_U4194 );
nand NAND2_17703 ( P1_U7487 , P1_U7091 , P1_U4194 );
nand NAND2_17704 ( P1_U7488 , P1_U4194 , P1_U3392 );
nand NAND2_17705 ( P1_U7489 , P1_U4236 , P1_STATE2_REG_0_ );
nand NAND3_17706 ( P1_U7490 , P1_U7785 , P1_U7784 , P1_U4072 );
nand NAND2_17707 ( P1_U7491 , P1_U4108 , P1_U7216 );
nand NAND2_17708 ( P1_U7492 , P1_U4109 , P1_U7094 );
not NOT1_17709 ( P1_U7493 , P1_U3279 );
not NOT1_17710 ( P1_U7494 , P1_U3276 );
nand NAND5_17711 ( P1_U7495 , P1_U4071 , P1_U2607 , P1_U4070 , P1_U4069 , P1_U4068 );
nand NAND2_17712 ( P1_U7496 , P1_U3734 , P1_U7493 );
nand NAND2_17713 ( P1_U7497 , P1_U3735 , P1_U5469 );
nand NAND2_17714 ( P1_U7498 , P1_U2425 , P1_U7493 );
nand NAND2_17715 ( P1_U7499 , P1_U2425 , P1_U7493 );
nand NAND3_17716 ( P1_U7500 , P1_U6361 , P1_U6360 , P1_U7499 );
nand NAND2_17717 ( P1_U7501 , P1_U7493 , P1_R2167_U17 );
nand NAND3_17718 ( P1_U7502 , P1_U7493 , P1_U4201 , P1_R2167_U17 );
nand NAND2_17719 ( P1_U7503 , P1_U7502 , P1_U6149 );
nand NAND2_17720 ( P1_U7504 , P1_U7493 , P1_U7085 );
nand NAND2_17721 ( P1_U7505 , P1_U7493 , P1_U7471 );
nand NAND3_17722 ( P1_U7506 , P1_U4116 , P1_U4115 , P1_U4114 );
nand NAND2_17723 ( P1_U7507 , P1_U3759 , P1_U7493 );
nand NAND3_17724 ( P1_U7508 , P1_U3761 , P1_U5565 , P1_U3760 );
nand NAND2_17725 ( P1_U7509 , P1_U3746 , P1_U2519 );
nand NAND2_17726 ( P1_U7510 , P1_U7493 , P1_U5962 );
nand NAND2_17727 ( P1_U7511 , P1_U7493 , P1_U5965 );
nand NAND2_17728 ( P1_U7512 , P1_U7493 , P1_U5968 );
nand NAND2_17729 ( P1_U7513 , P1_U7493 , P1_U5971 );
nand NAND2_17730 ( P1_U7514 , P1_U7493 , P1_U5974 );
nand NAND2_17731 ( P1_U7515 , P1_U7493 , P1_U5977 );
nand NAND2_17732 ( P1_U7516 , P1_U7493 , P1_U5980 );
nand NAND2_17733 ( P1_U7517 , P1_U7493 , P1_U5983 );
nand NAND2_17734 ( P1_U7518 , P1_U7493 , P1_U5986 );
nand NAND2_17735 ( P1_U7519 , P1_U7493 , P1_U5989 );
nand NAND2_17736 ( P1_U7520 , P1_U7493 , P1_U5992 );
nand NAND2_17737 ( P1_U7521 , P1_U7493 , P1_U5995 );
nand NAND2_17738 ( P1_U7522 , P1_U7493 , P1_U5998 );
nand NAND2_17739 ( P1_U7523 , P1_U7493 , P1_U6001 );
nand NAND2_17740 ( P1_U7524 , P1_U7493 , P1_U6004 );
nand NAND2_17741 ( P1_U7525 , P1_U7493 , P1_U6007 );
nand NAND2_17742 ( P1_U7526 , P1_U7493 , P1_U6010 );
nand NAND2_17743 ( P1_U7527 , P1_U7493 , P1_U6013 );
nand NAND2_17744 ( P1_U7528 , P1_U7493 , P1_U6016 );
nand NAND2_17745 ( P1_U7529 , P1_U7493 , P1_U6019 );
nand NAND2_17746 ( P1_U7530 , P1_U7493 , P1_U6022 );
nand NAND2_17747 ( P1_U7531 , P1_U7493 , P1_U6025 );
nand NAND2_17748 ( P1_U7532 , P1_U7493 , P1_U6028 );
nand NAND2_17749 ( P1_U7533 , P1_U7493 , P1_U6031 );
nand NAND2_17750 ( P1_U7534 , P1_U7493 , P1_U6034 );
nand NAND2_17751 ( P1_U7535 , P1_U7493 , P1_U6037 );
nand NAND2_17752 ( P1_U7536 , P1_U7493 , P1_U6040 );
nand NAND2_17753 ( P1_U7537 , P1_U7493 , P1_U6043 );
nand NAND2_17754 ( P1_U7538 , P1_U7493 , P1_U6046 );
nand NAND2_17755 ( P1_U7539 , P1_U7493 , P1_U6049 );
nand NAND2_17756 ( P1_U7540 , P1_U7493 , P1_U6052 );
nand NAND2_17757 ( P1_U7541 , P1_U2357 , P1_U7493 );
nand NAND2_17758 ( P1_U7542 , P1_UWORD_REG_0_ , P1_U7541 );
nand NAND2_17759 ( P1_U7543 , P1_U2357 , P1_U7493 );
nand NAND2_17760 ( P1_U7544 , P1_UWORD_REG_1_ , P1_U7543 );
nand NAND2_17761 ( P1_U7545 , P1_U2357 , P1_U7493 );
nand NAND2_17762 ( P1_U7546 , P1_UWORD_REG_2_ , P1_U7545 );
nand NAND2_17763 ( P1_U7547 , P1_U2357 , P1_U7493 );
nand NAND2_17764 ( P1_U7548 , P1_UWORD_REG_3_ , P1_U7547 );
nand NAND2_17765 ( P1_U7549 , P1_U2357 , P1_U7493 );
nand NAND2_17766 ( P1_U7550 , P1_UWORD_REG_4_ , P1_U7549 );
nand NAND2_17767 ( P1_U7551 , P1_U2357 , P1_U7493 );
nand NAND2_17768 ( P1_U7552 , P1_UWORD_REG_5_ , P1_U7551 );
nand NAND2_17769 ( P1_U7553 , P1_U2357 , P1_U7493 );
nand NAND2_17770 ( P1_U7554 , P1_UWORD_REG_6_ , P1_U7553 );
nand NAND2_17771 ( P1_U7555 , P1_U2357 , P1_U7493 );
nand NAND2_17772 ( P1_U7556 , P1_UWORD_REG_7_ , P1_U7555 );
nand NAND2_17773 ( P1_U7557 , P1_U2357 , P1_U7493 );
nand NAND2_17774 ( P1_U7558 , P1_UWORD_REG_8_ , P1_U7557 );
nand NAND2_17775 ( P1_U7559 , P1_U2357 , P1_U7493 );
nand NAND2_17776 ( P1_U7560 , P1_UWORD_REG_9_ , P1_U7559 );
nand NAND2_17777 ( P1_U7561 , P1_U2357 , P1_U7493 );
nand NAND2_17778 ( P1_U7562 , P1_UWORD_REG_10_ , P1_U7561 );
nand NAND2_17779 ( P1_U7563 , P1_U2357 , P1_U7493 );
nand NAND2_17780 ( P1_U7564 , P1_UWORD_REG_11_ , P1_U7563 );
nand NAND2_17781 ( P1_U7565 , P1_U2357 , P1_U7493 );
nand NAND2_17782 ( P1_U7566 , P1_UWORD_REG_12_ , P1_U7565 );
nand NAND2_17783 ( P1_U7567 , P1_U2357 , P1_U7493 );
nand NAND2_17784 ( P1_U7568 , P1_UWORD_REG_13_ , P1_U7567 );
nand NAND2_17785 ( P1_U7569 , P1_U2357 , P1_U7493 );
nand NAND2_17786 ( P1_U7570 , P1_UWORD_REG_14_ , P1_U7569 );
nand NAND2_17787 ( P1_U7571 , P1_U2357 , P1_U7493 );
nand NAND2_17788 ( P1_U7572 , P1_LWORD_REG_0_ , P1_U7571 );
nand NAND2_17789 ( P1_U7573 , P1_U2357 , P1_U7493 );
nand NAND2_17790 ( P1_U7574 , P1_LWORD_REG_1_ , P1_U7573 );
nand NAND2_17791 ( P1_U7575 , P1_U2357 , P1_U7493 );
nand NAND2_17792 ( P1_U7576 , P1_LWORD_REG_2_ , P1_U7575 );
nand NAND2_17793 ( P1_U7577 , P1_U2357 , P1_U7493 );
nand NAND2_17794 ( P1_U7578 , P1_LWORD_REG_3_ , P1_U7577 );
nand NAND2_17795 ( P1_U7579 , P1_U2357 , P1_U7493 );
nand NAND2_17796 ( P1_U7580 , P1_LWORD_REG_4_ , P1_U7579 );
nand NAND2_17797 ( P1_U7581 , P1_U2357 , P1_U7493 );
nand NAND2_17798 ( P1_U7582 , P1_LWORD_REG_5_ , P1_U7581 );
nand NAND2_17799 ( P1_U7583 , P1_U2357 , P1_U7493 );
nand NAND2_17800 ( P1_U7584 , P1_LWORD_REG_6_ , P1_U7583 );
nand NAND2_17801 ( P1_U7585 , P1_U2357 , P1_U7493 );
nand NAND2_17802 ( P1_U7586 , P1_LWORD_REG_7_ , P1_U7585 );
nand NAND2_17803 ( P1_U7587 , P1_U2357 , P1_U7493 );
nand NAND2_17804 ( P1_U7588 , P1_LWORD_REG_8_ , P1_U7587 );
nand NAND2_17805 ( P1_U7589 , P1_U2357 , P1_U7493 );
nand NAND2_17806 ( P1_U7590 , P1_LWORD_REG_9_ , P1_U7589 );
nand NAND2_17807 ( P1_U7591 , P1_U2357 , P1_U7493 );
nand NAND2_17808 ( P1_U7592 , P1_LWORD_REG_10_ , P1_U7591 );
nand NAND2_17809 ( P1_U7593 , P1_U2357 , P1_U7493 );
nand NAND2_17810 ( P1_U7594 , P1_LWORD_REG_11_ , P1_U7593 );
nand NAND2_17811 ( P1_U7595 , P1_U2357 , P1_U7493 );
nand NAND2_17812 ( P1_U7596 , P1_LWORD_REG_12_ , P1_U7595 );
nand NAND2_17813 ( P1_U7597 , P1_U2357 , P1_U7493 );
nand NAND2_17814 ( P1_U7598 , P1_LWORD_REG_13_ , P1_U7597 );
nand NAND2_17815 ( P1_U7599 , P1_U2357 , P1_U7493 );
nand NAND2_17816 ( P1_U7600 , P1_LWORD_REG_14_ , P1_U7599 );
nand NAND2_17817 ( P1_U7601 , P1_U2357 , P1_U7493 );
nand NAND2_17818 ( P1_U7602 , P1_LWORD_REG_15_ , P1_U7601 );
nand NAND3_17819 ( P1_U7603 , P1_U7493 , P1_U3568 , P1_U4259 );
nand NAND3_17820 ( P1_U7604 , P1_U7684 , P1_U7683 , P1_U3581 );
nand NAND2_17821 ( P1_U7605 , P1_U3867 , P1_U7493 );
nand NAND2_17822 ( P1_U7606 , P1_U7605 , P1_U3428 );
nand NAND2_17823 ( P1_U7607 , P1_U4208 , P1_U7493 );
nand NAND2_17824 ( P1_U7608 , P1_U7607 , P1_U3447 );
nand NAND2_17825 ( P1_U7609 , P1_U3279 , P1_U3400 );
nand NAND2_17826 ( P1_U7610 , P1_U3754 , P1_U7493 );
nand NAND2_17827 ( P1_U7611 , P1_U3755 , P1_U7610 );
nand NAND2_17828 ( P1_U7612 , P1_INSTQUEUE_REG_0__4_ , P1_U5416 );
nand NAND2_17829 ( P1_U7613 , P1_U2523 , P1_INSTQUEUE_REG_0__4_ );
nand NAND2_17830 ( P1_U7614 , P1_U2546 , P1_INSTQUEUE_REG_0__4_ );
nand NAND4_17831 ( P1_U7615 , P1_U4052 , P1_U4051 , P1_U4050 , P1_U4049 );
nand NAND2_17832 ( P1_U7616 , P1_U4192 , P1_INSTQUEUE_REG_0__4_ );
nand NAND2_17833 ( P1_U7617 , P1_U2573 , P1_INSTQUEUE_REG_0__4_ );
nand NAND4_17834 ( P1_U7618 , P1_U4091 , P1_U4089 , P1_U4088 , P1_U4087 );
nand NAND2_17835 ( P1_U7619 , P1_U2592 , P1_INSTQUEUE_REG_0__4_ );
nand NAND4_17836 ( P1_U7620 , P1_U4136 , P1_U4135 , P1_U4134 , P1_U4133 );
not NOT1_17837 ( P1_U7621 , P1_U3259 );
nand NAND2_17838 ( P1_U7622 , P1_U7621 , P1_U3261 );
nand NAND3_17839 ( P1_U7623 , P1_U4361 , P1_STATE_REG_1_ , P1_U4358 );
nand NAND2_17840 ( P1_U7624 , P1_STATE_REG_2_ , P1_U7468 );
nand NAND2_17841 ( P1_U7625 , P1_STATE_REG_1_ , P1_U4358 );
nand NAND2_17842 ( P1_U7626 , P1_U4502 , P1_U4510 );
nand NAND2_17843 ( P1_U7627 , P1_U5487 , P1_U4171 );
nand NAND2_17844 ( P1_U7628 , P1_U3283 , P1_U3289 );
not NOT1_17845 ( P1_U7629 , P1_U3392 );
nand NAND2_17846 ( P1_U7630 , P1_U4208 , P1_U7490 );
nand NAND2_17847 ( P1_U7631 , P1_U5487 , P1_U4171 );
nand NAND2_17848 ( P1_U7632 , P1_U7631 , P1_U7630 );
nand NAND2_17849 ( P1_U7633 , P1_BE_N_REG_3_ , P1_U3249 );
nand NAND2_17850 ( P1_U7634 , P1_BYTEENABLE_REG_3_ , P1_U4221 );
nand NAND2_17851 ( P1_U7635 , P1_BE_N_REG_2_ , P1_U3249 );
nand NAND2_17852 ( P1_U7636 , P1_BYTEENABLE_REG_2_ , P1_U4221 );
nand NAND2_17853 ( P1_U7637 , P1_BE_N_REG_1_ , P1_U3249 );
nand NAND2_17854 ( P1_U7638 , P1_BYTEENABLE_REG_1_ , P1_U4221 );
nand NAND2_17855 ( P1_U7639 , P1_BE_N_REG_0_ , P1_U3249 );
nand NAND2_17856 ( P1_U7640 , P1_BYTEENABLE_REG_0_ , P1_U4221 );
nand NAND3_17857 ( P1_U7641 , P1_STATE_REG_0_ , P1_REQUESTPENDING_REG , P1_U3251 );
nand NAND2_17858 ( P1_U7642 , P1_STATE_REG_2_ , P1_U3259 );
nand NAND2_17859 ( P1_U7643 , P1_U7642 , P1_U7641 );
nand NAND3_17860 ( P1_U7644 , P1_U7624 , P1_U4361 , P1_STATE_REG_1_ );
nand NAND2_17861 ( P1_U7645 , P1_U7643 , P1_U3248 );
nand NAND3_17862 ( P1_U7646 , P1_STATE_REG_0_ , P1_U3260 , P1_STATE_REG_2_ );
nand NAND2_17863 ( P1_U7647 , P1_U4371 , P1_U3251 );
or OR2_17864 ( P1_U7648 , P1_STATE_REG_0_ , P1_STATE_REG_1_ );
nand NAND2_17865 ( P1_U7649 , P1_STATE_REG_0_ , P1_U4258 );
not NOT1_17866 ( P1_U7650 , P1_U3462 );
nand NAND2_17867 ( P1_U7651 , P1_U7650 , P1_DATAWIDTH_REG_0_ );
nand NAND2_17868 ( P1_U7652 , P1_U3463 , P1_U3462 );
nand NAND2_17869 ( P1_U7653 , P1_U3462 , P1_U4376 );
nand NAND2_17870 ( P1_U7654 , P1_U7650 , P1_DATAWIDTH_REG_1_ );
nand NAND3_17871 ( P1_U7655 , P1_U3541 , P1_U3540 , P1_U3265 );
nand NAND5_17872 ( P1_U7656 , P1_INSTQUEUE_REG_7__4_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3270 , P1_INSTQUEUERD_ADDR_REG_1_ );
nand NAND5_17873 ( P1_U7657 , P1_INSTQUEUE_REG_5__4_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3270 , P1_U3265 );
nand NAND5_17874 ( P1_U7658 , P1_INSTQUEUE_REG_2__4_ , P1_U3270 , P1_U3264 , P1_U3266 , P1_INSTQUEUERD_ADDR_REG_1_ );
nand NAND3_17875 ( P1_U7659 , P1_U3543 , P1_U3542 , P1_U3270 );
nand NAND3_17876 ( P1_U7660 , P1_U3545 , P1_U3544 , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND3_17877 ( P1_U7661 , P1_U3547 , P1_U3546 , P1_U3265 );
nand NAND3_17878 ( P1_U7662 , P1_U3549 , P1_U3548 , P1_INSTQUEUERD_ADDR_REG_1_ );
nand NAND3_17879 ( P1_U7663 , P1_U3551 , P1_U3550 , P1_U3266 );
nand NAND5_17880 ( P1_U7664 , P1_INSTQUEUE_REG_15__4_ , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_INSTQUEUERD_ADDR_REG_2_ , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND5_17881 ( P1_U7665 , P1_INSTQUEUE_REG_0__4_ , P1_U3264 , P1_U3265 , P1_U3266 , P1_U3270 );
nand NAND5_17882 ( P1_U7666 , P1_INSTQUEUE_REG_8__4_ , P1_U3264 , P1_U3265 , P1_U3266 , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_17883 ( P1_U7667 , P1_INSTQUEUE_REG_10__4_ , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3264 , P1_U3266 );
nand NAND3_17884 ( P1_U7668 , P1_U3553 , P1_U3552 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND5_17885 ( P1_U7669 , P1_INSTQUEUE_REG_3__4_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3264 , P1_U3270 );
nand NAND5_17886 ( P1_U7670 , P1_INSTQUEUE_REG_11__4_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3264 , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_17887 ( P1_U7671 , P1_INSTQUEUE_REG_3__5_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3264 , P1_U3270 );
nand NAND3_17888 ( P1_U7672 , P1_U3529 , P1_U3528 , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND5_17889 ( P1_U7673 , P1_INSTQUEUE_REG_9__6_ , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_0_ , P1_U3264 , P1_U3265 );
nand NAND3_17890 ( P1_U7674 , P1_U3535 , P1_U3534 , P1_INSTQUEUERD_ADDR_REG_1_ );
nand NAND5_17891 ( P1_U7675 , P1_INSTQUEUE_REG_10__6_ , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3264 , P1_U3266 );
nand NAND5_17892 ( P1_U7676 , P1_INSTQUEUE_REG_11__6_ , P1_INSTQUEUERD_ADDR_REG_3_ , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3264 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND5_17893 ( P1_U7677 , P1_INSTQUEUE_REG_0__6_ , P1_U3264 , P1_U3265 , P1_U3266 , P1_U3270 );
nand NAND5_17894 ( P1_U7678 , P1_INSTQUEUE_REG_8__6_ , P1_U3264 , P1_U3265 , P1_U3266 , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_17895 ( P1_U7679 , P1_U4494 , P1_U3437 );
nand NAND2_17896 ( P1_U7680 , P1_U7501 , P1_U3284 );
nand NAND2_17897 ( P1_U7681 , P1_U4216 , P1_R2167_U17 );
nand NAND2_17898 ( P1_U7682 , P1_U4506 , P1_U3273 );
nand NAND2_17899 ( P1_U7683 , P1_STATE2_REG_0_ , P1_U4512 );
nand NAND2_17900 ( P1_U7684 , P1_U4513 , P1_U3294 );
nand NAND2_17901 ( P1_U7685 , P1_STATE2_REG_3_ , P1_U3295 );
nand NAND2_17902 ( P1_U7686 , P1_U2428 , P1_U4514 );
or OR2_17903 ( P1_U7687 , P1_STATEBS16_REG , P1_STATE2_REG_0_ );
nand NAND2_17904 ( P1_U7688 , P1_STATE2_REG_0_ , P1_U7469 );
nand NAND2_17905 ( P1_U7689 , P1_STATE2_REG_0_ , P1_U4522 );
nand NAND3_17906 ( P1_U7690 , P1_U7604 , P1_U4521 , P1_U3294 );
nand NAND2_17907 ( P1_U7691 , P1_R2144_U49 , P1_U3313 );
nand NAND2_17908 ( P1_U7692 , P1_U4528 , P1_U3311 );
not NOT1_17909 ( P1_U7693 , P1_U3454 );
nand NAND2_17910 ( P1_U7694 , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_U3305 );
nand NAND2_17911 ( P1_U7695 , P1_U4533 , P1_U3304 );
not NOT1_17912 ( P1_U7696 , P1_U3455 );
nand NAND2_17913 ( P1_U7697 , P1_U4216 , P1_U3273 );
nand NAND2_17914 ( P1_U7698 , P1_R2167_U17 , P1_U7497 );
nand NAND2_17915 ( P1_U7699 , P1_U4432 , P1_U5466 );
nand NAND2_17916 ( P1_U7700 , P1_U5467 , P1_U4171 );
nand NAND2_17917 ( P1_U7701 , P1_U3467 , P1_U4172 );
nand NAND2_17918 ( P1_U7702 , P1_U5476 , P1_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_17919 ( P1_U7703 , P1_U4460 , P1_U3278 );
nand NAND2_17920 ( P1_U7704 , P1_U4415 , P1_U3277 );
nand NAND2_17921 ( P1_U7705 , P1_U3271 , P1_U3415 );
nand NAND2_17922 ( P1_U7706 , P1_U4477 , P1_U5493 );
nand NAND2_17923 ( P1_U7707 , P1_U7706 , P1_U7705 );
nand NAND2_17924 ( P1_U7708 , P1_U5476 , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_17925 ( P1_U7709 , P1_U5509 , P1_U4172 );
nand NAND2_17926 ( P1_U7710 , P1_INSTADDRPOINTER_REG_1_ , P1_U4174 );
nand NAND2_17927 ( P1_U7711 , P1_SUB_580_U6 , P1_INSTADDRPOINTER_REG_31_ );
not NOT1_17928 ( P1_U7712 , P1_U3470 );
nand NAND2_17929 ( P1_U7713 , P1_INSTADDRPOINTER_REG_0_ , P1_U4174 );
nand NAND2_17930 ( P1_U7714 , P1_INSTADDRPOINTER_REG_0_ , P1_INSTADDRPOINTER_REG_31_ );
not NOT1_17931 ( P1_U7715 , P1_U3471 );
nand NAND2_17932 ( P1_U7716 , P1_U5511 , P1_U5501 );
nand NAND2_17933 ( P1_U7717 , P1_U4218 , P1_U3401 );
nand NAND2_17934 ( P1_U7718 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_U3264 );
nand NAND2_17935 ( P1_U7719 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_U3265 );
not NOT1_17936 ( P1_U7720 , P1_U3456 );
nand NAND2_17937 ( P1_U7721 , P1_U5476 , P1_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_17938 ( P1_U7722 , P1_U5518 , P1_U4172 );
nand NAND2_17939 ( P1_U7723 , P1_U5476 , P1_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_17940 ( P1_U7724 , P1_U5529 , P1_U4172 );
nand NAND2_17941 ( P1_U7725 , P1_U4214 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_17942 ( P1_U7726 , P1_U5521 , P1_U3266 );
nand NAND2_17943 ( P1_U7727 , P1_U5476 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_17944 ( P1_U7728 , P1_U5535 , P1_U4172 );
nand NAND2_17945 ( P1_U7729 , P1_U5537 , P1_INSTQUEUEWR_ADDR_REG_3_ );
nand NAND2_17946 ( P1_U7730 , P1_U5545 , P1_U3404 );
nand NAND2_17947 ( P1_U7731 , P1_U7693 , P1_U4527 );
nand NAND2_17948 ( P1_U7732 , P1_U3454 , P1_U3314 );
nand NAND2_17949 ( P1_U7733 , P1_U7732 , P1_U7731 );
nand NAND2_17950 ( P1_U7734 , P1_U5537 , P1_INSTQUEUEWR_ADDR_REG_2_ );
nand NAND2_17951 ( P1_U7735 , P1_U5549 , P1_U3404 );
nand NAND2_17952 ( P1_U7736 , P1_U5537 , P1_INSTQUEUEWR_ADDR_REG_1_ );
nand NAND2_17953 ( P1_U7737 , P1_U5554 , P1_U3404 );
nand NAND2_17954 ( P1_U7738 , P1_U5537 , P1_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_17955 ( P1_U7739 , P1_U5557 , P1_U3404 );
nand NAND2_17956 ( P1_U7740 , P1_U4477 , P1_U3388 );
nand NAND2_17957 ( P1_U7741 , P1_U3271 , P1_U3281 );
nand NAND4_17958 ( P1_U7742 , P1_U7741 , P1_U7740 , P1_U3257 , P1_U4171 );
nand NAND3_17959 ( P1_U7743 , P1_R2167_U17 , P1_U7611 , P1_U4432 );
nand NAND2_17960 ( P1_U7744 , P1_EAX_REG_31_ , P1_U3424 );
nand NAND2_17961 ( P1_U7745 , P1_U3479 , P1_U4223 );
nand NAND2_17962 ( P1_U7746 , P1_BYTEENABLE_REG_3_ , P1_U3433 );
nand NAND2_17963 ( P1_U7747 , P1_U3480 , P1_U4220 );
or OR2_17964 ( P1_U7748 , P1_DATAWIDTH_REG_0_ , P1_DATAWIDTH_REG_1_ );
nand NAND2_17965 ( P1_U7749 , P1_DATAWIDTH_REG_0_ , P1_U3413 );
nand NAND2_17966 ( P1_U7750 , P1_U7749 , P1_U7748 );
nand NAND2_17967 ( P1_U7751 , P1_U7750 , P1_U3253 );
nand NAND2_17968 ( P1_U7752 , P1_REIP_REG_0_ , P1_REIP_REG_1_ );
nand NAND2_17969 ( P1_U7753 , P1_U7752 , P1_U7751 );
nand NAND2_17970 ( P1_U7754 , P1_BYTEENABLE_REG_2_ , P1_U3433 );
nand NAND2_17971 ( P1_U7755 , P1_U7753 , P1_U4220 );
nand NAND2_17972 ( P1_U7756 , P1_BYTEENABLE_REG_1_ , P1_U3433 );
nand NAND2_17973 ( P1_U7757 , P1_U4220 , P1_REIP_REG_1_ );
nand NAND2_17974 ( P1_U7758 , P1_BYTEENABLE_REG_0_ , P1_U3433 );
nand NAND2_17975 ( P1_U7759 , P1_U4220 , P1_U6599 );
nand NAND2_17976 ( P1_U7760 , P1_U4221 , P1_U3436 );
nand NAND2_17977 ( P1_U7761 , P1_W_R_N_REG , P1_U3249 );
nand NAND2_17978 ( P1_U7762 , P1_MORE_REG , P1_U4177 );
nand NAND2_17979 ( P1_U7763 , P1_U4237 , P1_U6600 );
nand NAND2_17980 ( P1_U7764 , P1_U7650 , P1_STATEBS16_REG );
nand NAND2_17981 ( P1_U7765 , BS16 , P1_U3462 );
nand NAND2_17982 ( P1_U7766 , P1_U6603 , P1_REQUESTPENDING_REG );
nand NAND2_17983 ( P1_U7767 , P1_U6609 , P1_U4180 );
nand NAND2_17984 ( P1_U7768 , P1_U4221 , P1_U3435 );
nand NAND2_17985 ( P1_U7769 , P1_D_C_N_REG , P1_U3249 );
nand NAND2_17986 ( P1_U7770 , P1_M_IO_N_REG , P1_U3249 );
nand NAND2_17987 ( P1_U7771 , P1_MEMORYFETCH_REG , P1_U4221 );
nand NAND2_17988 ( P1_U7772 , P1_U6614 , P1_READREQUEST_REG );
nand NAND2_17989 ( P1_U7773 , P1_U6615 , P1_U4181 );
nand NAND2_17990 ( P1_U7774 , P1_U3488 , P1_U4182 );
nand NAND2_17991 ( P1_U7775 , P1_U5473 , P1_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_17992 ( P1_U7776 , P1_U5473 , P1_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_17993 ( P1_U7777 , P1_U5506 , P1_U4182 );
nand NAND2_17994 ( P1_U7778 , P1_U5473 , P1_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_17995 ( P1_U7779 , P1_U5514 , P1_U4182 );
nand NAND2_17996 ( P1_U7780 , P1_U5473 , P1_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_17997 ( P1_U7781 , P1_U5525 , P1_U4182 );
nand NAND2_17998 ( P1_U7782 , P1_U5473 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_17999 ( P1_U7783 , P1_U5531 , P1_U4182 );
nand NAND2_18000 ( P1_U7784 , P1_U2605 , P1_U3277 );
nand NAND2_18001 ( P1_U7785 , P1_U4460 , P1_U7495 );
nand NAND2_18002 ( P1_U7786 , P1_U4203 , P1_U3301 );
nand NAND2_18003 ( P1_U7787 , P1_INSTQUEUEWR_ADDR_REG_0_ , P1_U3297 );
nand NAND2_18004 ( P1_U7788 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_U4183 );
nand NAND2_18005 ( P1_U7789 , P1_U7219 , P1_U3270 );
not NOT1_18006 ( P1_U7790 , P1_U3457 );
nand NAND2_18007 ( P1_U7791 , P1_U3276 , P1_U3284 );
nand NAND2_18008 ( P1_U7792 , P1_U7707 , P1_U4494 );
nand NAND2_18009 ( P1_U7793 , P1_U3493 , P1_U3262 );
nand NAND3_18010 ( P1_U7794 , P1_FLUSH_REG , P1_U7715 , P1_STATE2_REG_1_ );
not NOT1_18011 ( P1_ADD_405_U113 , P1_ADD_405_U38 );
not NOT1_18012 ( P1_ADD_405_U112 , P1_ADD_405_U36 );
not NOT1_18013 ( P1_ADD_405_U111 , P1_ADD_405_U34 );
not NOT1_18014 ( P1_ADD_405_U110 , P1_ADD_405_U32 );
not NOT1_18015 ( P1_ADD_405_U109 , P1_ADD_405_U30 );
not NOT1_18016 ( P1_ADD_405_U108 , P1_ADD_405_U28 );
not NOT1_18017 ( P1_ADD_405_U107 , P1_ADD_405_U26 );
not NOT1_18018 ( P1_ADD_405_U106 , P1_ADD_405_U24 );
not NOT1_18019 ( P1_ADD_405_U105 , P1_ADD_405_U22 );
not NOT1_18020 ( P1_ADD_405_U104 , P1_ADD_405_U20 );
not NOT1_18021 ( P1_ADD_405_U103 , P1_ADD_405_U18 );
not NOT1_18022 ( P1_ADD_405_U102 , P1_ADD_405_U16 );
not NOT1_18023 ( P1_ADD_405_U101 , P1_ADD_405_U14 );
not NOT1_18024 ( P1_ADD_405_U100 , P1_ADD_405_U13 );
not NOT1_18025 ( P1_ADD_405_U99 , P1_ADD_405_U10 );
not NOT1_18026 ( P1_ADD_405_U98 , P1_ADD_405_U8 );
not NOT1_18027 ( P1_ADD_405_U97 , P1_ADD_405_U94 );
nand NAND2_18028 ( P1_ADD_405_U96 , P1_INSTADDRPOINTER_REG_1_ , P1_INSTADDRPOINTER_REG_0_ );
and AND2_18029 ( P1_ADD_405_U95 , P1_ADD_405_U172 , P1_ADD_405_U171 );
nand NAND2_18030 ( P1_ADD_405_U94 , P1_ADD_405_U62 , P1_ADD_405_U96 );
nand NAND2_18031 ( P1_ADD_405_U93 , P1_ADD_405_U124 , P1_INSTADDRPOINTER_REG_30_ );
not NOT1_18032 ( P1_ADD_405_U92 , P1_INSTADDRPOINTER_REG_31_ );
nand NAND2_18033 ( P1_ADD_405_U91 , P1_ADD_405_U186 , P1_ADD_405_U185 );
nand NAND2_18034 ( P1_ADD_405_U90 , P1_ADD_405_U184 , P1_ADD_405_U183 );
nand NAND2_18035 ( P1_ADD_405_U89 , P1_ADD_405_U182 , P1_ADD_405_U181 );
nand NAND2_18036 ( P1_ADD_405_U88 , P1_ADD_405_U180 , P1_ADD_405_U179 );
nand NAND2_18037 ( P1_ADD_405_U87 , P1_ADD_405_U178 , P1_ADD_405_U177 );
nand NAND2_18038 ( LT_782_120_U6 , P3_DATAO_REG_30_ , LT_782_120_U7 );
not NOT1_18039 ( LT_782_120_U7 , P3_DATAO_REG_31_ );
nand NAND2_18040 ( LT_782_U6 , P1_DATAO_REG_30_ , LT_782_U7 );
not NOT1_18041 ( LT_782_U7 , P1_DATAO_REG_31_ );
not NOT1_18042 ( LT_748_U6 , P2_ADDRESS_REG_29_ );
and AND2_18043 ( R170_U6 , P2_ADDRESS_REG_29_ , R170_U15 );
or OR4_18044 ( R170_U7 , P2_ADDRESS_REG_17_ , P2_ADDRESS_REG_9_ , P2_ADDRESS_REG_7_ , P2_ADDRESS_REG_22_ );
nor nor_18045 ( R170_U8 , R170_U7 , P2_ADDRESS_REG_10_ , P2_ADDRESS_REG_19_ , P2_ADDRESS_REG_25_ , P2_ADDRESS_REG_24_ );
or OR4_18046 ( R170_U9 , P2_ADDRESS_REG_16_ , P2_ADDRESS_REG_0_ , P2_ADDRESS_REG_18_ , P2_ADDRESS_REG_8_ );
nor nor_18047 ( R170_U10 , R170_U9 , P2_ADDRESS_REG_23_ , P2_ADDRESS_REG_1_ , P2_ADDRESS_REG_11_ );
or OR4_18048 ( R170_U11 , P2_ADDRESS_REG_26_ , P2_ADDRESS_REG_21_ , P2_ADDRESS_REG_28_ , P2_ADDRESS_REG_6_ );
nor nor_18049 ( R170_U12 , R170_U11 , P2_ADDRESS_REG_12_ , P2_ADDRESS_REG_14_ , P2_ADDRESS_REG_4_ );
or OR4_18050 ( R170_U13 , P2_ADDRESS_REG_13_ , P2_ADDRESS_REG_20_ , P2_ADDRESS_REG_3_ , P2_ADDRESS_REG_27_ );
nor nor_18051 ( R170_U14 , R170_U13 , P2_ADDRESS_REG_2_ , P2_ADDRESS_REG_5_ , P2_ADDRESS_REG_15_ );
nand NAND4_18052 ( R170_U15 , R170_U14 , R170_U12 , R170_U10 , R170_U8 );
and AND2_18053 ( R165_U6 , P1_ADDRESS_REG_29_ , R165_U15 );
or OR4_18054 ( R165_U7 , P1_ADDRESS_REG_17_ , P1_ADDRESS_REG_9_ , P1_ADDRESS_REG_7_ , P1_ADDRESS_REG_22_ );
nor nor_18055 ( R165_U8 , R165_U7 , P1_ADDRESS_REG_10_ , P1_ADDRESS_REG_19_ , P1_ADDRESS_REG_25_ , P1_ADDRESS_REG_24_ );
or OR4_18056 ( R165_U9 , P1_ADDRESS_REG_16_ , P1_ADDRESS_REG_0_ , P1_ADDRESS_REG_18_ , P1_ADDRESS_REG_8_ );
nor nor_18057 ( R165_U10 , R165_U9 , P1_ADDRESS_REG_23_ , P1_ADDRESS_REG_1_ , P1_ADDRESS_REG_11_ );
or OR4_18058 ( R165_U11 , P1_ADDRESS_REG_26_ , P1_ADDRESS_REG_21_ , P1_ADDRESS_REG_28_ , P1_ADDRESS_REG_6_ );
nor nor_18059 ( R165_U12 , R165_U11 , P1_ADDRESS_REG_12_ , P1_ADDRESS_REG_14_ , P1_ADDRESS_REG_4_ );
or OR4_18060 ( R165_U13 , P1_ADDRESS_REG_13_ , P1_ADDRESS_REG_20_ , P1_ADDRESS_REG_3_ , P1_ADDRESS_REG_27_ );
nor nor_18061 ( R165_U14 , R165_U13 , P1_ADDRESS_REG_2_ , P1_ADDRESS_REG_5_ , P1_ADDRESS_REG_15_ );
nand NAND4_18062 ( R165_U15 , R165_U14 , R165_U12 , R165_U10 , R165_U8 );
nand NAND2_18063 ( LT_782_119_U6 , P2_DATAO_REG_30_ , LT_782_119_U7 );
not NOT1_18064 ( LT_782_119_U7 , P2_DATAO_REG_31_ );
not NOT1_18065 ( P3_ADD_526_U5 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_18066 ( P3_ADD_526_U6 , P3_INSTADDRPOINTER_REG_2_ );
not NOT1_18067 ( P3_ADD_526_U7 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_18068 ( P3_ADD_526_U8 , P3_INSTADDRPOINTER_REG_4_ );
not NOT1_18069 ( P3_ADD_526_U9 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND3_18070 ( P3_ADD_526_U10 , P3_INSTADDRPOINTER_REG_2_ , P3_INSTADDRPOINTER_REG_0_ , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_18071 ( P3_ADD_526_U11 , P3_INSTADDRPOINTER_REG_6_ );
not NOT1_18072 ( P3_ADD_526_U12 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_18073 ( P3_ADD_526_U13 , P3_ADD_526_U82 , P3_ADD_526_U111 );
not NOT1_18074 ( P3_ADD_526_U14 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_18075 ( P3_ADD_526_U15 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_18076 ( P3_ADD_526_U16 , P3_ADD_526_U83 , P3_ADD_526_U112 );
nand NAND2_18077 ( P3_ADD_526_U17 , P3_ADD_526_U84 , P3_ADD_526_U118 );
not NOT1_18078 ( P3_ADD_526_U18 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_18079 ( P3_ADD_526_U19 , P3_INSTADDRPOINTER_REG_10_ );
not NOT1_18080 ( P3_ADD_526_U20 , P3_INSTADDRPOINTER_REG_12_ );
not NOT1_18081 ( P3_ADD_526_U21 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_18082 ( P3_ADD_526_U22 , P3_ADD_526_U85 , P3_ADD_526_U120 );
not NOT1_18083 ( P3_ADD_526_U23 , P3_INSTADDRPOINTER_REG_14_ );
not NOT1_18084 ( P3_ADD_526_U24 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_18085 ( P3_ADD_526_U25 , P3_ADD_526_U86 , P3_ADD_526_U113 );
not NOT1_18086 ( P3_ADD_526_U26 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_18087 ( P3_ADD_526_U27 , P3_ADD_526_U87 , P3_ADD_526_U119 );
not NOT1_18088 ( P3_ADD_526_U28 , P3_INSTADDRPOINTER_REG_16_ );
not NOT1_18089 ( P3_ADD_526_U29 , P3_INSTADDRPOINTER_REG_18_ );
not NOT1_18090 ( P3_ADD_526_U30 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_18091 ( P3_ADD_526_U31 , P3_ADD_526_U88 , P3_ADD_526_U124 );
not NOT1_18092 ( P3_ADD_526_U32 , P3_INSTADDRPOINTER_REG_20_ );
not NOT1_18093 ( P3_ADD_526_U33 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_18094 ( P3_ADD_526_U34 , P3_ADD_526_U89 , P3_ADD_526_U117 );
not NOT1_18095 ( P3_ADD_526_U35 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_18096 ( P3_ADD_526_U36 , P3_ADD_526_U90 , P3_ADD_526_U114 );
not NOT1_18097 ( P3_ADD_526_U37 , P3_INSTADDRPOINTER_REG_22_ );
not NOT1_18098 ( P3_ADD_526_U38 , P3_INSTADDRPOINTER_REG_24_ );
not NOT1_18099 ( P3_ADD_526_U39 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_18100 ( P3_ADD_526_U40 , P3_ADD_526_U91 , P3_ADD_526_U121 );
not NOT1_18101 ( P3_ADD_526_U41 , P3_INSTADDRPOINTER_REG_26_ );
not NOT1_18102 ( P3_ADD_526_U42 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_18103 ( P3_ADD_526_U43 , P3_ADD_526_U92 , P3_ADD_526_U115 );
not NOT1_18104 ( P3_ADD_526_U44 , P3_INSTADDRPOINTER_REG_27_ );
not NOT1_18105 ( P3_ADD_526_U45 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_18106 ( P3_ADD_526_U46 , P3_ADD_526_U93 , P3_ADD_526_U116 );
not NOT1_18107 ( P3_ADD_526_U47 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_18108 ( P3_ADD_526_U48 , P3_ADD_526_U94 , P3_ADD_526_U122 );
nand NAND2_18109 ( P3_ADD_526_U49 , P3_ADD_526_U123 , P3_INSTADDRPOINTER_REG_29_ );
not NOT1_18110 ( P3_ADD_526_U50 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_18111 ( P3_ADD_526_U51 , P3_ADD_526_U142 , P3_ADD_526_U141 );
nand NAND2_18112 ( P3_ADD_526_U52 , P3_ADD_526_U144 , P3_ADD_526_U143 );
nand NAND2_18113 ( P3_ADD_526_U53 , P3_ADD_526_U146 , P3_ADD_526_U145 );
nand NAND2_18114 ( P3_ADD_526_U54 , P3_ADD_526_U148 , P3_ADD_526_U147 );
nand NAND2_18115 ( P3_ADD_526_U55 , P3_ADD_526_U150 , P3_ADD_526_U149 );
nand NAND2_18116 ( P3_ADD_526_U56 , P3_ADD_526_U152 , P3_ADD_526_U151 );
nand NAND2_18117 ( P3_ADD_526_U57 , P3_ADD_526_U154 , P3_ADD_526_U153 );
nand NAND2_18118 ( P3_ADD_526_U58 , P3_ADD_526_U156 , P3_ADD_526_U155 );
nand NAND2_18119 ( P3_ADD_526_U59 , P3_ADD_526_U158 , P3_ADD_526_U157 );
nand NAND2_18120 ( P3_ADD_526_U60 , P3_ADD_526_U160 , P3_ADD_526_U159 );
nand NAND2_18121 ( P3_ADD_526_U61 , P3_ADD_526_U162 , P3_ADD_526_U161 );
nand NAND2_18122 ( P3_ADD_526_U62 , P3_ADD_526_U164 , P3_ADD_526_U163 );
nand NAND2_18123 ( P3_ADD_526_U63 , P3_ADD_526_U166 , P3_ADD_526_U165 );
nand NAND2_18124 ( P3_ADD_526_U64 , P3_ADD_526_U168 , P3_ADD_526_U167 );
nand NAND2_18125 ( P3_ADD_526_U65 , P3_ADD_526_U170 , P3_ADD_526_U169 );
nand NAND2_18126 ( P3_ADD_526_U66 , P3_ADD_526_U172 , P3_ADD_526_U171 );
nand NAND2_18127 ( P3_ADD_526_U67 , P3_ADD_526_U174 , P3_ADD_526_U173 );
nand NAND2_18128 ( P3_ADD_526_U68 , P3_ADD_526_U176 , P3_ADD_526_U175 );
nand NAND2_18129 ( P3_ADD_526_U69 , P3_ADD_526_U178 , P3_ADD_526_U177 );
nand NAND2_18130 ( P3_ADD_526_U70 , P3_ADD_526_U180 , P3_ADD_526_U179 );
nand NAND2_18131 ( P3_ADD_526_U71 , P3_ADD_526_U182 , P3_ADD_526_U181 );
nand NAND2_18132 ( P3_ADD_526_U72 , P3_ADD_526_U184 , P3_ADD_526_U183 );
nand NAND2_18133 ( P3_ADD_526_U73 , P3_ADD_526_U186 , P3_ADD_526_U185 );
nand NAND2_18134 ( P3_ADD_526_U74 , P3_ADD_526_U188 , P3_ADD_526_U187 );
nand NAND2_18135 ( P3_ADD_526_U75 , P3_ADD_526_U190 , P3_ADD_526_U189 );
nand NAND2_18136 ( P3_ADD_526_U76 , P3_ADD_526_U192 , P3_ADD_526_U191 );
nand NAND2_18137 ( P3_ADD_526_U77 , P3_ADD_526_U194 , P3_ADD_526_U193 );
nand NAND2_18138 ( P3_ADD_526_U78 , P3_ADD_526_U196 , P3_ADD_526_U195 );
nand NAND2_18139 ( P3_ADD_526_U79 , P3_ADD_526_U198 , P3_ADD_526_U197 );
nand NAND2_18140 ( P3_ADD_526_U80 , P3_ADD_526_U200 , P3_ADD_526_U199 );
nand NAND2_18141 ( P3_ADD_526_U81 , P3_ADD_526_U202 , P3_ADD_526_U201 );
and AND2_18142 ( P3_ADD_526_U82 , P3_INSTADDRPOINTER_REG_3_ , P3_INSTADDRPOINTER_REG_4_ );
and AND2_18143 ( P3_ADD_526_U83 , P3_INSTADDRPOINTER_REG_5_ , P3_INSTADDRPOINTER_REG_6_ );
and AND2_18144 ( P3_ADD_526_U84 , P3_INSTADDRPOINTER_REG_7_ , P3_INSTADDRPOINTER_REG_8_ );
and AND2_18145 ( P3_ADD_526_U85 , P3_INSTADDRPOINTER_REG_9_ , P3_INSTADDRPOINTER_REG_10_ );
and AND2_18146 ( P3_ADD_526_U86 , P3_INSTADDRPOINTER_REG_11_ , P3_INSTADDRPOINTER_REG_12_ );
and AND2_18147 ( P3_ADD_526_U87 , P3_INSTADDRPOINTER_REG_13_ , P3_INSTADDRPOINTER_REG_14_ );
and AND2_18148 ( P3_ADD_526_U88 , P3_INSTADDRPOINTER_REG_16_ , P3_INSTADDRPOINTER_REG_15_ );
and AND2_18149 ( P3_ADD_526_U89 , P3_INSTADDRPOINTER_REG_17_ , P3_INSTADDRPOINTER_REG_18_ );
and AND2_18150 ( P3_ADD_526_U90 , P3_INSTADDRPOINTER_REG_19_ , P3_INSTADDRPOINTER_REG_20_ );
and AND2_18151 ( P3_ADD_526_U91 , P3_INSTADDRPOINTER_REG_22_ , P3_INSTADDRPOINTER_REG_21_ );
and AND2_18152 ( P3_ADD_526_U92 , P3_INSTADDRPOINTER_REG_23_ , P3_INSTADDRPOINTER_REG_24_ );
and AND2_18153 ( P3_ADD_526_U93 , P3_INSTADDRPOINTER_REG_25_ , P3_INSTADDRPOINTER_REG_26_ );
and AND2_18154 ( P3_ADD_526_U94 , P3_INSTADDRPOINTER_REG_28_ , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_18155 ( P3_ADD_526_U95 , P3_ADD_526_U118 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_18156 ( P3_ADD_526_U96 , P3_ADD_526_U112 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_18157 ( P3_ADD_526_U97 , P3_ADD_526_U111 , P3_INSTADDRPOINTER_REG_3_ );
not NOT1_18158 ( P3_ADD_526_U98 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_18159 ( P3_ADD_526_U99 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_526_U128 );
nand NAND2_18160 ( P3_ADD_526_U100 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
nand NAND2_18161 ( P3_ADD_526_U101 , P3_ADD_526_U122 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_18162 ( P3_ADD_526_U102 , P3_ADD_526_U116 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_18163 ( P3_ADD_526_U103 , P3_ADD_526_U115 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_18164 ( P3_ADD_526_U104 , P3_ADD_526_U121 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_18165 ( P3_ADD_526_U105 , P3_ADD_526_U114 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_18166 ( P3_ADD_526_U106 , P3_ADD_526_U117 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_18167 ( P3_ADD_526_U107 , P3_ADD_526_U124 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_18168 ( P3_ADD_526_U108 , P3_ADD_526_U119 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_18169 ( P3_ADD_526_U109 , P3_ADD_526_U113 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_18170 ( P3_ADD_526_U110 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_526_U120 );
not NOT1_18171 ( P3_ADD_526_U111 , P3_ADD_526_U10 );
not NOT1_18172 ( P3_ADD_526_U112 , P3_ADD_526_U13 );
not NOT1_18173 ( P3_ADD_526_U113 , P3_ADD_526_U22 );
not NOT1_18174 ( P3_ADD_526_U114 , P3_ADD_526_U34 );
not NOT1_18175 ( P3_ADD_526_U115 , P3_ADD_526_U40 );
not NOT1_18176 ( P3_ADD_526_U116 , P3_ADD_526_U43 );
not NOT1_18177 ( P3_ADD_526_U117 , P3_ADD_526_U31 );
not NOT1_18178 ( P3_ADD_526_U118 , P3_ADD_526_U16 );
not NOT1_18179 ( P3_ADD_526_U119 , P3_ADD_526_U25 );
not NOT1_18180 ( P3_ADD_526_U120 , P3_ADD_526_U17 );
not NOT1_18181 ( P3_ADD_526_U121 , P3_ADD_526_U36 );
not NOT1_18182 ( P3_ADD_526_U122 , P3_ADD_526_U46 );
not NOT1_18183 ( P3_ADD_526_U123 , P3_ADD_526_U48 );
not NOT1_18184 ( P3_ADD_526_U124 , P3_ADD_526_U27 );
not NOT1_18185 ( P3_ADD_526_U125 , P3_ADD_526_U95 );
not NOT1_18186 ( P3_ADD_526_U126 , P3_ADD_526_U96 );
not NOT1_18187 ( P3_ADD_526_U127 , P3_ADD_526_U97 );
not NOT1_18188 ( P3_ADD_526_U128 , P3_ADD_526_U49 );
not NOT1_18189 ( P3_ADD_526_U129 , P3_ADD_526_U99 );
not NOT1_18190 ( P3_ADD_526_U130 , P3_ADD_526_U100 );
not NOT1_18191 ( P3_ADD_526_U131 , P3_ADD_526_U101 );
not NOT1_18192 ( P3_ADD_526_U132 , P3_ADD_526_U102 );
not NOT1_18193 ( P3_ADD_526_U133 , P3_ADD_526_U103 );
not NOT1_18194 ( P3_ADD_526_U134 , P3_ADD_526_U104 );
not NOT1_18195 ( P3_ADD_526_U135 , P3_ADD_526_U105 );
not NOT1_18196 ( P3_ADD_526_U136 , P3_ADD_526_U106 );
not NOT1_18197 ( P3_ADD_526_U137 , P3_ADD_526_U107 );
not NOT1_18198 ( P3_ADD_526_U138 , P3_ADD_526_U108 );
not NOT1_18199 ( P3_ADD_526_U139 , P3_ADD_526_U109 );
not NOT1_18200 ( P3_ADD_526_U140 , P3_ADD_526_U110 );
nand NAND2_18201 ( P3_ADD_526_U141 , P3_ADD_526_U120 , P3_ADD_526_U18 );
nand NAND2_18202 ( P3_ADD_526_U142 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_526_U17 );
nand NAND2_18203 ( P3_ADD_526_U143 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_526_U95 );
nand NAND2_18204 ( P3_ADD_526_U144 , P3_ADD_526_U125 , P3_ADD_526_U14 );
nand NAND2_18205 ( P3_ADD_526_U145 , P3_ADD_526_U118 , P3_ADD_526_U15 );
nand NAND2_18206 ( P3_ADD_526_U146 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_526_U16 );
nand NAND2_18207 ( P3_ADD_526_U147 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_526_U96 );
nand NAND2_18208 ( P3_ADD_526_U148 , P3_ADD_526_U126 , P3_ADD_526_U11 );
nand NAND2_18209 ( P3_ADD_526_U149 , P3_ADD_526_U112 , P3_ADD_526_U12 );
nand NAND2_18210 ( P3_ADD_526_U150 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_526_U13 );
nand NAND2_18211 ( P3_ADD_526_U151 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_526_U97 );
nand NAND2_18212 ( P3_ADD_526_U152 , P3_ADD_526_U127 , P3_ADD_526_U8 );
nand NAND2_18213 ( P3_ADD_526_U153 , P3_ADD_526_U111 , P3_ADD_526_U9 );
nand NAND2_18214 ( P3_ADD_526_U154 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_526_U10 );
nand NAND2_18215 ( P3_ADD_526_U155 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_526_U99 );
nand NAND2_18216 ( P3_ADD_526_U156 , P3_ADD_526_U129 , P3_ADD_526_U98 );
nand NAND2_18217 ( P3_ADD_526_U157 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_526_U49 );
nand NAND2_18218 ( P3_ADD_526_U158 , P3_ADD_526_U128 , P3_ADD_526_U50 );
nand NAND2_18219 ( P3_ADD_526_U159 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_526_U100 );
nand NAND2_18220 ( P3_ADD_526_U160 , P3_ADD_526_U130 , P3_ADD_526_U6 );
nand NAND2_18221 ( P3_ADD_526_U161 , P3_ADD_526_U123 , P3_ADD_526_U47 );
nand NAND2_18222 ( P3_ADD_526_U162 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_526_U48 );
nand NAND2_18223 ( P3_ADD_526_U163 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_526_U101 );
nand NAND2_18224 ( P3_ADD_526_U164 , P3_ADD_526_U131 , P3_ADD_526_U45 );
nand NAND2_18225 ( P3_ADD_526_U165 , P3_ADD_526_U122 , P3_ADD_526_U44 );
nand NAND2_18226 ( P3_ADD_526_U166 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_526_U46 );
nand NAND2_18227 ( P3_ADD_526_U167 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_526_U102 );
nand NAND2_18228 ( P3_ADD_526_U168 , P3_ADD_526_U132 , P3_ADD_526_U41 );
nand NAND2_18229 ( P3_ADD_526_U169 , P3_ADD_526_U116 , P3_ADD_526_U42 );
nand NAND2_18230 ( P3_ADD_526_U170 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_526_U43 );
nand NAND2_18231 ( P3_ADD_526_U171 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_526_U103 );
nand NAND2_18232 ( P3_ADD_526_U172 , P3_ADD_526_U133 , P3_ADD_526_U38 );
nand NAND2_18233 ( P3_ADD_526_U173 , P3_ADD_526_U115 , P3_ADD_526_U39 );
nand NAND2_18234 ( P3_ADD_526_U174 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_526_U40 );
nand NAND2_18235 ( P3_ADD_526_U175 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_526_U104 );
nand NAND2_18236 ( P3_ADD_526_U176 , P3_ADD_526_U134 , P3_ADD_526_U37 );
nand NAND2_18237 ( P3_ADD_526_U177 , P3_ADD_526_U121 , P3_ADD_526_U35 );
nand NAND2_18238 ( P3_ADD_526_U178 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_526_U36 );
nand NAND2_18239 ( P3_ADD_526_U179 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_526_U105 );
nand NAND2_18240 ( P3_ADD_526_U180 , P3_ADD_526_U135 , P3_ADD_526_U32 );
nand NAND2_18241 ( P3_ADD_526_U181 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_526_U7 );
nand NAND2_18242 ( P3_ADD_526_U182 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_526_U5 );
nand NAND2_18243 ( P3_ADD_526_U183 , P3_ADD_526_U114 , P3_ADD_526_U33 );
nand NAND2_18244 ( P3_ADD_526_U184 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_526_U34 );
nand NAND2_18245 ( P3_ADD_526_U185 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_526_U106 );
nand NAND2_18246 ( P3_ADD_526_U186 , P3_ADD_526_U136 , P3_ADD_526_U29 );
nand NAND2_18247 ( P3_ADD_526_U187 , P3_ADD_526_U117 , P3_ADD_526_U30 );
nand NAND2_18248 ( P3_ADD_526_U188 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_526_U31 );
nand NAND2_18249 ( P3_ADD_526_U189 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_526_U107 );
nand NAND2_18250 ( P3_ADD_526_U190 , P3_ADD_526_U137 , P3_ADD_526_U28 );
nand NAND2_18251 ( P3_ADD_526_U191 , P3_ADD_526_U124 , P3_ADD_526_U26 );
nand NAND2_18252 ( P3_ADD_526_U192 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_526_U27 );
nand NAND2_18253 ( P3_ADD_526_U193 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_526_U108 );
nand NAND2_18254 ( P3_ADD_526_U194 , P3_ADD_526_U138 , P3_ADD_526_U23 );
nand NAND2_18255 ( P3_ADD_526_U195 , P3_ADD_526_U119 , P3_ADD_526_U24 );
nand NAND2_18256 ( P3_ADD_526_U196 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_526_U25 );
nand NAND2_18257 ( P3_ADD_526_U197 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_526_U109 );
nand NAND2_18258 ( P3_ADD_526_U198 , P3_ADD_526_U139 , P3_ADD_526_U20 );
nand NAND2_18259 ( P3_ADD_526_U199 , P3_ADD_526_U113 , P3_ADD_526_U21 );
nand NAND2_18260 ( P3_ADD_526_U200 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_526_U22 );
nand NAND2_18261 ( P3_ADD_526_U201 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_526_U110 );
nand NAND2_18262 ( P3_ADD_526_U202 , P3_ADD_526_U140 , P3_ADD_526_U19 );
not NOT1_18263 ( P3_ADD_552_U5 , P3_EBX_REG_0_ );
not NOT1_18264 ( P3_ADD_552_U6 , P3_EBX_REG_2_ );
not NOT1_18265 ( P3_ADD_552_U7 , P3_EBX_REG_1_ );
not NOT1_18266 ( P3_ADD_552_U8 , P3_EBX_REG_4_ );
not NOT1_18267 ( P3_ADD_552_U9 , P3_EBX_REG_3_ );
nand NAND3_18268 ( P3_ADD_552_U10 , P3_EBX_REG_2_ , P3_EBX_REG_0_ , P3_EBX_REG_1_ );
not NOT1_18269 ( P3_ADD_552_U11 , P3_EBX_REG_6_ );
not NOT1_18270 ( P3_ADD_552_U12 , P3_EBX_REG_5_ );
nand NAND2_18271 ( P3_ADD_552_U13 , P3_ADD_552_U82 , P3_ADD_552_U111 );
not NOT1_18272 ( P3_ADD_552_U14 , P3_EBX_REG_8_ );
not NOT1_18273 ( P3_ADD_552_U15 , P3_EBX_REG_7_ );
nand NAND2_18274 ( P3_ADD_552_U16 , P3_ADD_552_U83 , P3_ADD_552_U112 );
nand NAND2_18275 ( P3_ADD_552_U17 , P3_ADD_552_U84 , P3_ADD_552_U118 );
not NOT1_18276 ( P3_ADD_552_U18 , P3_EBX_REG_9_ );
not NOT1_18277 ( P3_ADD_552_U19 , P3_EBX_REG_10_ );
not NOT1_18278 ( P3_ADD_552_U20 , P3_EBX_REG_12_ );
not NOT1_18279 ( P3_ADD_552_U21 , P3_EBX_REG_11_ );
nand NAND2_18280 ( P3_ADD_552_U22 , P3_ADD_552_U85 , P3_ADD_552_U120 );
not NOT1_18281 ( P3_ADD_552_U23 , P3_EBX_REG_14_ );
not NOT1_18282 ( P3_ADD_552_U24 , P3_EBX_REG_13_ );
nand NAND2_18283 ( P3_ADD_552_U25 , P3_ADD_552_U86 , P3_ADD_552_U113 );
not NOT1_18284 ( P3_ADD_552_U26 , P3_EBX_REG_15_ );
nand NAND2_18285 ( P3_ADD_552_U27 , P3_ADD_552_U87 , P3_ADD_552_U119 );
not NOT1_18286 ( P3_ADD_552_U28 , P3_EBX_REG_16_ );
not NOT1_18287 ( P3_ADD_552_U29 , P3_EBX_REG_18_ );
not NOT1_18288 ( P3_ADD_552_U30 , P3_EBX_REG_17_ );
nand NAND2_18289 ( P3_ADD_552_U31 , P3_ADD_552_U88 , P3_ADD_552_U124 );
not NOT1_18290 ( P3_ADD_552_U32 , P3_EBX_REG_20_ );
not NOT1_18291 ( P3_ADD_552_U33 , P3_EBX_REG_19_ );
nand NAND2_18292 ( P3_ADD_552_U34 , P3_ADD_552_U89 , P3_ADD_552_U117 );
not NOT1_18293 ( P3_ADD_552_U35 , P3_EBX_REG_21_ );
nand NAND2_18294 ( P3_ADD_552_U36 , P3_ADD_552_U90 , P3_ADD_552_U114 );
not NOT1_18295 ( P3_ADD_552_U37 , P3_EBX_REG_22_ );
not NOT1_18296 ( P3_ADD_552_U38 , P3_EBX_REG_24_ );
not NOT1_18297 ( P3_ADD_552_U39 , P3_EBX_REG_23_ );
nand NAND2_18298 ( P3_ADD_552_U40 , P3_ADD_552_U91 , P3_ADD_552_U121 );
not NOT1_18299 ( P3_ADD_552_U41 , P3_EBX_REG_26_ );
not NOT1_18300 ( P3_ADD_552_U42 , P3_EBX_REG_25_ );
nand NAND2_18301 ( P3_ADD_552_U43 , P3_ADD_552_U92 , P3_ADD_552_U115 );
not NOT1_18302 ( P3_ADD_552_U44 , P3_EBX_REG_27_ );
not NOT1_18303 ( P3_ADD_552_U45 , P3_EBX_REG_28_ );
nand NAND2_18304 ( P3_ADD_552_U46 , P3_ADD_552_U93 , P3_ADD_552_U116 );
not NOT1_18305 ( P3_ADD_552_U47 , P3_EBX_REG_29_ );
nand NAND2_18306 ( P3_ADD_552_U48 , P3_ADD_552_U94 , P3_ADD_552_U122 );
nand NAND2_18307 ( P3_ADD_552_U49 , P3_ADD_552_U123 , P3_EBX_REG_29_ );
not NOT1_18308 ( P3_ADD_552_U50 , P3_EBX_REG_30_ );
nand NAND2_18309 ( P3_ADD_552_U51 , P3_ADD_552_U142 , P3_ADD_552_U141 );
nand NAND2_18310 ( P3_ADD_552_U52 , P3_ADD_552_U144 , P3_ADD_552_U143 );
nand NAND2_18311 ( P3_ADD_552_U53 , P3_ADD_552_U146 , P3_ADD_552_U145 );
nand NAND2_18312 ( P3_ADD_552_U54 , P3_ADD_552_U148 , P3_ADD_552_U147 );
nand NAND2_18313 ( P3_ADD_552_U55 , P3_ADD_552_U150 , P3_ADD_552_U149 );
nand NAND2_18314 ( P3_ADD_552_U56 , P3_ADD_552_U152 , P3_ADD_552_U151 );
nand NAND2_18315 ( P3_ADD_552_U57 , P3_ADD_552_U154 , P3_ADD_552_U153 );
nand NAND2_18316 ( P3_ADD_552_U58 , P3_ADD_552_U156 , P3_ADD_552_U155 );
nand NAND2_18317 ( P3_ADD_552_U59 , P3_ADD_552_U158 , P3_ADD_552_U157 );
nand NAND2_18318 ( P3_ADD_552_U60 , P3_ADD_552_U160 , P3_ADD_552_U159 );
nand NAND2_18319 ( P3_ADD_552_U61 , P3_ADD_552_U162 , P3_ADD_552_U161 );
nand NAND2_18320 ( P3_ADD_552_U62 , P3_ADD_552_U164 , P3_ADD_552_U163 );
nand NAND2_18321 ( P3_ADD_552_U63 , P3_ADD_552_U166 , P3_ADD_552_U165 );
nand NAND2_18322 ( P3_ADD_552_U64 , P3_ADD_552_U168 , P3_ADD_552_U167 );
nand NAND2_18323 ( P3_ADD_552_U65 , P3_ADD_552_U170 , P3_ADD_552_U169 );
nand NAND2_18324 ( P3_ADD_552_U66 , P3_ADD_552_U172 , P3_ADD_552_U171 );
nand NAND2_18325 ( P3_ADD_552_U67 , P3_ADD_552_U174 , P3_ADD_552_U173 );
nand NAND2_18326 ( P3_ADD_552_U68 , P3_ADD_552_U176 , P3_ADD_552_U175 );
nand NAND2_18327 ( P3_ADD_552_U69 , P3_ADD_552_U178 , P3_ADD_552_U177 );
nand NAND2_18328 ( P3_ADD_552_U70 , P3_ADD_552_U180 , P3_ADD_552_U179 );
nand NAND2_18329 ( P3_ADD_552_U71 , P3_ADD_552_U182 , P3_ADD_552_U181 );
nand NAND2_18330 ( P3_ADD_552_U72 , P3_ADD_552_U184 , P3_ADD_552_U183 );
nand NAND2_18331 ( P3_ADD_552_U73 , P3_ADD_552_U186 , P3_ADD_552_U185 );
nand NAND2_18332 ( P3_ADD_552_U74 , P3_ADD_552_U188 , P3_ADD_552_U187 );
nand NAND2_18333 ( P3_ADD_552_U75 , P3_ADD_552_U190 , P3_ADD_552_U189 );
nand NAND2_18334 ( P3_ADD_552_U76 , P3_ADD_552_U192 , P3_ADD_552_U191 );
nand NAND2_18335 ( P3_ADD_552_U77 , P3_ADD_552_U194 , P3_ADD_552_U193 );
nand NAND2_18336 ( P3_ADD_552_U78 , P3_ADD_552_U196 , P3_ADD_552_U195 );
nand NAND2_18337 ( P3_ADD_552_U79 , P3_ADD_552_U198 , P3_ADD_552_U197 );
nand NAND2_18338 ( P3_ADD_552_U80 , P3_ADD_552_U200 , P3_ADD_552_U199 );
nand NAND2_18339 ( P3_ADD_552_U81 , P3_ADD_552_U202 , P3_ADD_552_U201 );
and AND2_18340 ( P3_ADD_552_U82 , P3_EBX_REG_3_ , P3_EBX_REG_4_ );
and AND2_18341 ( P3_ADD_552_U83 , P3_EBX_REG_5_ , P3_EBX_REG_6_ );
and AND2_18342 ( P3_ADD_552_U84 , P3_EBX_REG_7_ , P3_EBX_REG_8_ );
and AND2_18343 ( P3_ADD_552_U85 , P3_EBX_REG_9_ , P3_EBX_REG_10_ );
and AND2_18344 ( P3_ADD_552_U86 , P3_EBX_REG_11_ , P3_EBX_REG_12_ );
and AND2_18345 ( P3_ADD_552_U87 , P3_EBX_REG_13_ , P3_EBX_REG_14_ );
and AND2_18346 ( P3_ADD_552_U88 , P3_EBX_REG_16_ , P3_EBX_REG_15_ );
and AND2_18347 ( P3_ADD_552_U89 , P3_EBX_REG_17_ , P3_EBX_REG_18_ );
and AND2_18348 ( P3_ADD_552_U90 , P3_EBX_REG_19_ , P3_EBX_REG_20_ );
and AND2_18349 ( P3_ADD_552_U91 , P3_EBX_REG_22_ , P3_EBX_REG_21_ );
and AND2_18350 ( P3_ADD_552_U92 , P3_EBX_REG_23_ , P3_EBX_REG_24_ );
and AND2_18351 ( P3_ADD_552_U93 , P3_EBX_REG_25_ , P3_EBX_REG_26_ );
and AND2_18352 ( P3_ADD_552_U94 , P3_EBX_REG_28_ , P3_EBX_REG_27_ );
nand NAND2_18353 ( P3_ADD_552_U95 , P3_ADD_552_U118 , P3_EBX_REG_7_ );
nand NAND2_18354 ( P3_ADD_552_U96 , P3_ADD_552_U112 , P3_EBX_REG_5_ );
nand NAND2_18355 ( P3_ADD_552_U97 , P3_ADD_552_U111 , P3_EBX_REG_3_ );
not NOT1_18356 ( P3_ADD_552_U98 , P3_EBX_REG_31_ );
nand NAND2_18357 ( P3_ADD_552_U99 , P3_EBX_REG_30_ , P3_ADD_552_U128 );
nand NAND2_18358 ( P3_ADD_552_U100 , P3_EBX_REG_1_ , P3_EBX_REG_0_ );
nand NAND2_18359 ( P3_ADD_552_U101 , P3_ADD_552_U122 , P3_EBX_REG_27_ );
nand NAND2_18360 ( P3_ADD_552_U102 , P3_ADD_552_U116 , P3_EBX_REG_25_ );
nand NAND2_18361 ( P3_ADD_552_U103 , P3_ADD_552_U115 , P3_EBX_REG_23_ );
nand NAND2_18362 ( P3_ADD_552_U104 , P3_ADD_552_U121 , P3_EBX_REG_21_ );
nand NAND2_18363 ( P3_ADD_552_U105 , P3_ADD_552_U114 , P3_EBX_REG_19_ );
nand NAND2_18364 ( P3_ADD_552_U106 , P3_ADD_552_U117 , P3_EBX_REG_17_ );
nand NAND2_18365 ( P3_ADD_552_U107 , P3_ADD_552_U124 , P3_EBX_REG_15_ );
nand NAND2_18366 ( P3_ADD_552_U108 , P3_ADD_552_U119 , P3_EBX_REG_13_ );
nand NAND2_18367 ( P3_ADD_552_U109 , P3_ADD_552_U113 , P3_EBX_REG_11_ );
nand NAND2_18368 ( P3_ADD_552_U110 , P3_EBX_REG_9_ , P3_ADD_552_U120 );
not NOT1_18369 ( P3_ADD_552_U111 , P3_ADD_552_U10 );
not NOT1_18370 ( P3_ADD_552_U112 , P3_ADD_552_U13 );
not NOT1_18371 ( P3_ADD_552_U113 , P3_ADD_552_U22 );
not NOT1_18372 ( P3_ADD_552_U114 , P3_ADD_552_U34 );
not NOT1_18373 ( P3_ADD_552_U115 , P3_ADD_552_U40 );
not NOT1_18374 ( P3_ADD_552_U116 , P3_ADD_552_U43 );
not NOT1_18375 ( P3_ADD_552_U117 , P3_ADD_552_U31 );
not NOT1_18376 ( P3_ADD_552_U118 , P3_ADD_552_U16 );
not NOT1_18377 ( P3_ADD_552_U119 , P3_ADD_552_U25 );
not NOT1_18378 ( P3_ADD_552_U120 , P3_ADD_552_U17 );
not NOT1_18379 ( P3_ADD_552_U121 , P3_ADD_552_U36 );
not NOT1_18380 ( P3_ADD_552_U122 , P3_ADD_552_U46 );
not NOT1_18381 ( P3_ADD_552_U123 , P3_ADD_552_U48 );
not NOT1_18382 ( P3_ADD_552_U124 , P3_ADD_552_U27 );
not NOT1_18383 ( P3_ADD_552_U125 , P3_ADD_552_U95 );
not NOT1_18384 ( P3_ADD_552_U126 , P3_ADD_552_U96 );
not NOT1_18385 ( P3_ADD_552_U127 , P3_ADD_552_U97 );
not NOT1_18386 ( P3_ADD_552_U128 , P3_ADD_552_U49 );
not NOT1_18387 ( P3_ADD_552_U129 , P3_ADD_552_U99 );
not NOT1_18388 ( P3_ADD_552_U130 , P3_ADD_552_U100 );
not NOT1_18389 ( P3_ADD_552_U131 , P3_ADD_552_U101 );
not NOT1_18390 ( P3_ADD_552_U132 , P3_ADD_552_U102 );
not NOT1_18391 ( P3_ADD_552_U133 , P3_ADD_552_U103 );
not NOT1_18392 ( P3_ADD_552_U134 , P3_ADD_552_U104 );
not NOT1_18393 ( P3_ADD_552_U135 , P3_ADD_552_U105 );
not NOT1_18394 ( P3_ADD_552_U136 , P3_ADD_552_U106 );
not NOT1_18395 ( P3_ADD_552_U137 , P3_ADD_552_U107 );
not NOT1_18396 ( P3_ADD_552_U138 , P3_ADD_552_U108 );
not NOT1_18397 ( P3_ADD_552_U139 , P3_ADD_552_U109 );
not NOT1_18398 ( P3_ADD_552_U140 , P3_ADD_552_U110 );
nand NAND2_18399 ( P3_ADD_552_U141 , P3_ADD_552_U120 , P3_ADD_552_U18 );
nand NAND2_18400 ( P3_ADD_552_U142 , P3_EBX_REG_9_ , P3_ADD_552_U17 );
nand NAND2_18401 ( P3_ADD_552_U143 , P3_EBX_REG_8_ , P3_ADD_552_U95 );
nand NAND2_18402 ( P3_ADD_552_U144 , P3_ADD_552_U125 , P3_ADD_552_U14 );
nand NAND2_18403 ( P3_ADD_552_U145 , P3_ADD_552_U118 , P3_ADD_552_U15 );
nand NAND2_18404 ( P3_ADD_552_U146 , P3_EBX_REG_7_ , P3_ADD_552_U16 );
nand NAND2_18405 ( P3_ADD_552_U147 , P3_EBX_REG_6_ , P3_ADD_552_U96 );
nand NAND2_18406 ( P3_ADD_552_U148 , P3_ADD_552_U126 , P3_ADD_552_U11 );
nand NAND2_18407 ( P3_ADD_552_U149 , P3_ADD_552_U112 , P3_ADD_552_U12 );
nand NAND2_18408 ( P3_ADD_552_U150 , P3_EBX_REG_5_ , P3_ADD_552_U13 );
nand NAND2_18409 ( P3_ADD_552_U151 , P3_EBX_REG_4_ , P3_ADD_552_U97 );
nand NAND2_18410 ( P3_ADD_552_U152 , P3_ADD_552_U127 , P3_ADD_552_U8 );
nand NAND2_18411 ( P3_ADD_552_U153 , P3_ADD_552_U111 , P3_ADD_552_U9 );
nand NAND2_18412 ( P3_ADD_552_U154 , P3_EBX_REG_3_ , P3_ADD_552_U10 );
nand NAND2_18413 ( P3_ADD_552_U155 , P3_EBX_REG_31_ , P3_ADD_552_U99 );
nand NAND2_18414 ( P3_ADD_552_U156 , P3_ADD_552_U129 , P3_ADD_552_U98 );
nand NAND2_18415 ( P3_ADD_552_U157 , P3_EBX_REG_30_ , P3_ADD_552_U49 );
nand NAND2_18416 ( P3_ADD_552_U158 , P3_ADD_552_U128 , P3_ADD_552_U50 );
nand NAND2_18417 ( P3_ADD_552_U159 , P3_EBX_REG_2_ , P3_ADD_552_U100 );
nand NAND2_18418 ( P3_ADD_552_U160 , P3_ADD_552_U130 , P3_ADD_552_U6 );
nand NAND2_18419 ( P3_ADD_552_U161 , P3_ADD_552_U123 , P3_ADD_552_U47 );
nand NAND2_18420 ( P3_ADD_552_U162 , P3_EBX_REG_29_ , P3_ADD_552_U48 );
nand NAND2_18421 ( P3_ADD_552_U163 , P3_EBX_REG_28_ , P3_ADD_552_U101 );
nand NAND2_18422 ( P3_ADD_552_U164 , P3_ADD_552_U131 , P3_ADD_552_U45 );
nand NAND2_18423 ( P3_ADD_552_U165 , P3_ADD_552_U122 , P3_ADD_552_U44 );
nand NAND2_18424 ( P3_ADD_552_U166 , P3_EBX_REG_27_ , P3_ADD_552_U46 );
nand NAND2_18425 ( P3_ADD_552_U167 , P3_EBX_REG_26_ , P3_ADD_552_U102 );
nand NAND2_18426 ( P3_ADD_552_U168 , P3_ADD_552_U132 , P3_ADD_552_U41 );
nand NAND2_18427 ( P3_ADD_552_U169 , P3_ADD_552_U116 , P3_ADD_552_U42 );
nand NAND2_18428 ( P3_ADD_552_U170 , P3_EBX_REG_25_ , P3_ADD_552_U43 );
nand NAND2_18429 ( P3_ADD_552_U171 , P3_EBX_REG_24_ , P3_ADD_552_U103 );
nand NAND2_18430 ( P3_ADD_552_U172 , P3_ADD_552_U133 , P3_ADD_552_U38 );
nand NAND2_18431 ( P3_ADD_552_U173 , P3_ADD_552_U115 , P3_ADD_552_U39 );
nand NAND2_18432 ( P3_ADD_552_U174 , P3_EBX_REG_23_ , P3_ADD_552_U40 );
nand NAND2_18433 ( P3_ADD_552_U175 , P3_EBX_REG_22_ , P3_ADD_552_U104 );
nand NAND2_18434 ( P3_ADD_552_U176 , P3_ADD_552_U134 , P3_ADD_552_U37 );
nand NAND2_18435 ( P3_ADD_552_U177 , P3_ADD_552_U121 , P3_ADD_552_U35 );
nand NAND2_18436 ( P3_ADD_552_U178 , P3_EBX_REG_21_ , P3_ADD_552_U36 );
nand NAND2_18437 ( P3_ADD_552_U179 , P3_EBX_REG_20_ , P3_ADD_552_U105 );
nand NAND2_18438 ( P3_ADD_552_U180 , P3_ADD_552_U135 , P3_ADD_552_U32 );
nand NAND2_18439 ( P3_ADD_552_U181 , P3_EBX_REG_0_ , P3_ADD_552_U7 );
nand NAND2_18440 ( P3_ADD_552_U182 , P3_EBX_REG_1_ , P3_ADD_552_U5 );
nand NAND2_18441 ( P3_ADD_552_U183 , P3_ADD_552_U114 , P3_ADD_552_U33 );
nand NAND2_18442 ( P3_ADD_552_U184 , P3_EBX_REG_19_ , P3_ADD_552_U34 );
nand NAND2_18443 ( P3_ADD_552_U185 , P3_EBX_REG_18_ , P3_ADD_552_U106 );
nand NAND2_18444 ( P3_ADD_552_U186 , P3_ADD_552_U136 , P3_ADD_552_U29 );
nand NAND2_18445 ( P3_ADD_552_U187 , P3_ADD_552_U117 , P3_ADD_552_U30 );
nand NAND2_18446 ( P3_ADD_552_U188 , P3_EBX_REG_17_ , P3_ADD_552_U31 );
nand NAND2_18447 ( P3_ADD_552_U189 , P3_EBX_REG_16_ , P3_ADD_552_U107 );
nand NAND2_18448 ( P3_ADD_552_U190 , P3_ADD_552_U137 , P3_ADD_552_U28 );
nand NAND2_18449 ( P3_ADD_552_U191 , P3_ADD_552_U124 , P3_ADD_552_U26 );
nand NAND2_18450 ( P3_ADD_552_U192 , P3_EBX_REG_15_ , P3_ADD_552_U27 );
nand NAND2_18451 ( P3_ADD_552_U193 , P3_EBX_REG_14_ , P3_ADD_552_U108 );
nand NAND2_18452 ( P3_ADD_552_U194 , P3_ADD_552_U138 , P3_ADD_552_U23 );
nand NAND2_18453 ( P3_ADD_552_U195 , P3_ADD_552_U119 , P3_ADD_552_U24 );
nand NAND2_18454 ( P3_ADD_552_U196 , P3_EBX_REG_13_ , P3_ADD_552_U25 );
nand NAND2_18455 ( P3_ADD_552_U197 , P3_EBX_REG_12_ , P3_ADD_552_U109 );
nand NAND2_18456 ( P3_ADD_552_U198 , P3_ADD_552_U139 , P3_ADD_552_U20 );
nand NAND2_18457 ( P3_ADD_552_U199 , P3_ADD_552_U113 , P3_ADD_552_U21 );
nand NAND2_18458 ( P3_ADD_552_U200 , P3_EBX_REG_11_ , P3_ADD_552_U22 );
nand NAND2_18459 ( P3_ADD_552_U201 , P3_EBX_REG_10_ , P3_ADD_552_U110 );
nand NAND2_18460 ( P3_ADD_552_U202 , P3_ADD_552_U140 , P3_ADD_552_U19 );
not NOT1_18461 ( P3_ADD_546_U5 , P3_EAX_REG_0_ );
not NOT1_18462 ( P3_ADD_546_U6 , P3_EAX_REG_2_ );
not NOT1_18463 ( P3_ADD_546_U7 , P3_EAX_REG_1_ );
not NOT1_18464 ( P3_ADD_546_U8 , P3_EAX_REG_4_ );
not NOT1_18465 ( P3_ADD_546_U9 , P3_EAX_REG_3_ );
nand NAND3_18466 ( P3_ADD_546_U10 , P3_EAX_REG_2_ , P3_EAX_REG_0_ , P3_EAX_REG_1_ );
not NOT1_18467 ( P3_ADD_546_U11 , P3_EAX_REG_6_ );
not NOT1_18468 ( P3_ADD_546_U12 , P3_EAX_REG_5_ );
nand NAND2_18469 ( P3_ADD_546_U13 , P3_ADD_546_U82 , P3_ADD_546_U111 );
not NOT1_18470 ( P3_ADD_546_U14 , P3_EAX_REG_8_ );
not NOT1_18471 ( P3_ADD_546_U15 , P3_EAX_REG_7_ );
nand NAND2_18472 ( P3_ADD_546_U16 , P3_ADD_546_U83 , P3_ADD_546_U112 );
nand NAND2_18473 ( P3_ADD_546_U17 , P3_ADD_546_U84 , P3_ADD_546_U118 );
not NOT1_18474 ( P3_ADD_546_U18 , P3_EAX_REG_9_ );
not NOT1_18475 ( P3_ADD_546_U19 , P3_EAX_REG_10_ );
not NOT1_18476 ( P3_ADD_546_U20 , P3_EAX_REG_12_ );
not NOT1_18477 ( P3_ADD_546_U21 , P3_EAX_REG_11_ );
nand NAND2_18478 ( P3_ADD_546_U22 , P3_ADD_546_U85 , P3_ADD_546_U120 );
not NOT1_18479 ( P3_ADD_546_U23 , P3_EAX_REG_14_ );
not NOT1_18480 ( P3_ADD_546_U24 , P3_EAX_REG_13_ );
nand NAND2_18481 ( P3_ADD_546_U25 , P3_ADD_546_U86 , P3_ADD_546_U113 );
not NOT1_18482 ( P3_ADD_546_U26 , P3_EAX_REG_15_ );
nand NAND2_18483 ( P3_ADD_546_U27 , P3_ADD_546_U87 , P3_ADD_546_U119 );
not NOT1_18484 ( P3_ADD_546_U28 , P3_EAX_REG_16_ );
not NOT1_18485 ( P3_ADD_546_U29 , P3_EAX_REG_18_ );
not NOT1_18486 ( P3_ADD_546_U30 , P3_EAX_REG_17_ );
nand NAND2_18487 ( P3_ADD_546_U31 , P3_ADD_546_U88 , P3_ADD_546_U124 );
not NOT1_18488 ( P3_ADD_546_U32 , P3_EAX_REG_20_ );
not NOT1_18489 ( P3_ADD_546_U33 , P3_EAX_REG_19_ );
nand NAND2_18490 ( P3_ADD_546_U34 , P3_ADD_546_U89 , P3_ADD_546_U117 );
not NOT1_18491 ( P3_ADD_546_U35 , P3_EAX_REG_21_ );
nand NAND2_18492 ( P3_ADD_546_U36 , P3_ADD_546_U90 , P3_ADD_546_U114 );
not NOT1_18493 ( P3_ADD_546_U37 , P3_EAX_REG_22_ );
not NOT1_18494 ( P3_ADD_546_U38 , P3_EAX_REG_24_ );
not NOT1_18495 ( P3_ADD_546_U39 , P3_EAX_REG_23_ );
nand NAND2_18496 ( P3_ADD_546_U40 , P3_ADD_546_U91 , P3_ADD_546_U121 );
not NOT1_18497 ( P3_ADD_546_U41 , P3_EAX_REG_26_ );
not NOT1_18498 ( P3_ADD_546_U42 , P3_EAX_REG_25_ );
nand NAND2_18499 ( P3_ADD_546_U43 , P3_ADD_546_U92 , P3_ADD_546_U115 );
not NOT1_18500 ( P3_ADD_546_U44 , P3_EAX_REG_27_ );
not NOT1_18501 ( P3_ADD_546_U45 , P3_EAX_REG_28_ );
nand NAND2_18502 ( P3_ADD_546_U46 , P3_ADD_546_U93 , P3_ADD_546_U116 );
not NOT1_18503 ( P3_ADD_546_U47 , P3_EAX_REG_29_ );
nand NAND2_18504 ( P3_ADD_546_U48 , P3_ADD_546_U94 , P3_ADD_546_U122 );
nand NAND2_18505 ( P3_ADD_546_U49 , P3_ADD_546_U123 , P3_EAX_REG_29_ );
not NOT1_18506 ( P3_ADD_546_U50 , P3_EAX_REG_30_ );
nand NAND2_18507 ( P3_ADD_546_U51 , P3_ADD_546_U142 , P3_ADD_546_U141 );
nand NAND2_18508 ( P3_ADD_546_U52 , P3_ADD_546_U144 , P3_ADD_546_U143 );
nand NAND2_18509 ( P3_ADD_546_U53 , P3_ADD_546_U146 , P3_ADD_546_U145 );
nand NAND2_18510 ( P3_ADD_546_U54 , P3_ADD_546_U148 , P3_ADD_546_U147 );
nand NAND2_18511 ( P3_ADD_546_U55 , P3_ADD_546_U150 , P3_ADD_546_U149 );
nand NAND2_18512 ( P3_ADD_546_U56 , P3_ADD_546_U152 , P3_ADD_546_U151 );
nand NAND2_18513 ( P3_ADD_546_U57 , P3_ADD_546_U154 , P3_ADD_546_U153 );
nand NAND2_18514 ( P3_ADD_546_U58 , P3_ADD_546_U156 , P3_ADD_546_U155 );
nand NAND2_18515 ( P3_ADD_546_U59 , P3_ADD_546_U158 , P3_ADD_546_U157 );
nand NAND2_18516 ( P3_ADD_546_U60 , P3_ADD_546_U160 , P3_ADD_546_U159 );
nand NAND2_18517 ( P3_ADD_546_U61 , P3_ADD_546_U162 , P3_ADD_546_U161 );
nand NAND2_18518 ( P3_ADD_546_U62 , P3_ADD_546_U164 , P3_ADD_546_U163 );
nand NAND2_18519 ( P3_ADD_546_U63 , P3_ADD_546_U166 , P3_ADD_546_U165 );
nand NAND2_18520 ( P3_ADD_546_U64 , P3_ADD_546_U168 , P3_ADD_546_U167 );
nand NAND2_18521 ( P3_ADD_546_U65 , P3_ADD_546_U170 , P3_ADD_546_U169 );
nand NAND2_18522 ( P3_ADD_546_U66 , P3_ADD_546_U172 , P3_ADD_546_U171 );
nand NAND2_18523 ( P3_ADD_546_U67 , P3_ADD_546_U174 , P3_ADD_546_U173 );
nand NAND2_18524 ( P3_ADD_546_U68 , P3_ADD_546_U176 , P3_ADD_546_U175 );
nand NAND2_18525 ( P3_ADD_546_U69 , P3_ADD_546_U178 , P3_ADD_546_U177 );
nand NAND2_18526 ( P3_ADD_546_U70 , P3_ADD_546_U180 , P3_ADD_546_U179 );
nand NAND2_18527 ( P3_ADD_546_U71 , P3_ADD_546_U182 , P3_ADD_546_U181 );
nand NAND2_18528 ( P3_ADD_546_U72 , P3_ADD_546_U184 , P3_ADD_546_U183 );
nand NAND2_18529 ( P3_ADD_546_U73 , P3_ADD_546_U186 , P3_ADD_546_U185 );
nand NAND2_18530 ( P3_ADD_546_U74 , P3_ADD_546_U188 , P3_ADD_546_U187 );
nand NAND2_18531 ( P3_ADD_546_U75 , P3_ADD_546_U190 , P3_ADD_546_U189 );
nand NAND2_18532 ( P3_ADD_546_U76 , P3_ADD_546_U192 , P3_ADD_546_U191 );
nand NAND2_18533 ( P3_ADD_546_U77 , P3_ADD_546_U194 , P3_ADD_546_U193 );
nand NAND2_18534 ( P3_ADD_546_U78 , P3_ADD_546_U196 , P3_ADD_546_U195 );
nand NAND2_18535 ( P3_ADD_546_U79 , P3_ADD_546_U198 , P3_ADD_546_U197 );
nand NAND2_18536 ( P3_ADD_546_U80 , P3_ADD_546_U200 , P3_ADD_546_U199 );
nand NAND2_18537 ( P3_ADD_546_U81 , P3_ADD_546_U202 , P3_ADD_546_U201 );
and AND2_18538 ( P3_ADD_546_U82 , P3_EAX_REG_3_ , P3_EAX_REG_4_ );
and AND2_18539 ( P3_ADD_546_U83 , P3_EAX_REG_5_ , P3_EAX_REG_6_ );
and AND2_18540 ( P3_ADD_546_U84 , P3_EAX_REG_7_ , P3_EAX_REG_8_ );
and AND2_18541 ( P3_ADD_546_U85 , P3_EAX_REG_9_ , P3_EAX_REG_10_ );
and AND2_18542 ( P3_ADD_546_U86 , P3_EAX_REG_11_ , P3_EAX_REG_12_ );
and AND2_18543 ( P3_ADD_546_U87 , P3_EAX_REG_13_ , P3_EAX_REG_14_ );
and AND2_18544 ( P3_ADD_546_U88 , P3_EAX_REG_16_ , P3_EAX_REG_15_ );
and AND2_18545 ( P3_ADD_546_U89 , P3_EAX_REG_17_ , P3_EAX_REG_18_ );
and AND2_18546 ( P3_ADD_546_U90 , P3_EAX_REG_19_ , P3_EAX_REG_20_ );
and AND2_18547 ( P3_ADD_546_U91 , P3_EAX_REG_22_ , P3_EAX_REG_21_ );
and AND2_18548 ( P3_ADD_546_U92 , P3_EAX_REG_23_ , P3_EAX_REG_24_ );
and AND2_18549 ( P3_ADD_546_U93 , P3_EAX_REG_25_ , P3_EAX_REG_26_ );
and AND2_18550 ( P3_ADD_546_U94 , P3_EAX_REG_28_ , P3_EAX_REG_27_ );
nand NAND2_18551 ( P3_ADD_546_U95 , P3_ADD_546_U118 , P3_EAX_REG_7_ );
nand NAND2_18552 ( P3_ADD_546_U96 , P3_ADD_546_U112 , P3_EAX_REG_5_ );
nand NAND2_18553 ( P3_ADD_546_U97 , P3_ADD_546_U111 , P3_EAX_REG_3_ );
not NOT1_18554 ( P3_ADD_546_U98 , P3_EAX_REG_31_ );
nand NAND2_18555 ( P3_ADD_546_U99 , P3_EAX_REG_30_ , P3_ADD_546_U128 );
nand NAND2_18556 ( P3_ADD_546_U100 , P3_EAX_REG_1_ , P3_EAX_REG_0_ );
nand NAND2_18557 ( P3_ADD_546_U101 , P3_ADD_546_U122 , P3_EAX_REG_27_ );
nand NAND2_18558 ( P3_ADD_546_U102 , P3_ADD_546_U116 , P3_EAX_REG_25_ );
nand NAND2_18559 ( P3_ADD_546_U103 , P3_ADD_546_U115 , P3_EAX_REG_23_ );
nand NAND2_18560 ( P3_ADD_546_U104 , P3_ADD_546_U121 , P3_EAX_REG_21_ );
nand NAND2_18561 ( P3_ADD_546_U105 , P3_ADD_546_U114 , P3_EAX_REG_19_ );
nand NAND2_18562 ( P3_ADD_546_U106 , P3_ADD_546_U117 , P3_EAX_REG_17_ );
nand NAND2_18563 ( P3_ADD_546_U107 , P3_ADD_546_U124 , P3_EAX_REG_15_ );
nand NAND2_18564 ( P3_ADD_546_U108 , P3_ADD_546_U119 , P3_EAX_REG_13_ );
nand NAND2_18565 ( P3_ADD_546_U109 , P3_ADD_546_U113 , P3_EAX_REG_11_ );
nand NAND2_18566 ( P3_ADD_546_U110 , P3_EAX_REG_9_ , P3_ADD_546_U120 );
not NOT1_18567 ( P3_ADD_546_U111 , P3_ADD_546_U10 );
not NOT1_18568 ( P3_ADD_546_U112 , P3_ADD_546_U13 );
not NOT1_18569 ( P3_ADD_546_U113 , P3_ADD_546_U22 );
not NOT1_18570 ( P3_ADD_546_U114 , P3_ADD_546_U34 );
not NOT1_18571 ( P3_ADD_546_U115 , P3_ADD_546_U40 );
not NOT1_18572 ( P3_ADD_546_U116 , P3_ADD_546_U43 );
not NOT1_18573 ( P3_ADD_546_U117 , P3_ADD_546_U31 );
not NOT1_18574 ( P3_ADD_546_U118 , P3_ADD_546_U16 );
not NOT1_18575 ( P3_ADD_546_U119 , P3_ADD_546_U25 );
not NOT1_18576 ( P3_ADD_546_U120 , P3_ADD_546_U17 );
not NOT1_18577 ( P3_ADD_546_U121 , P3_ADD_546_U36 );
not NOT1_18578 ( P3_ADD_546_U122 , P3_ADD_546_U46 );
not NOT1_18579 ( P3_ADD_546_U123 , P3_ADD_546_U48 );
not NOT1_18580 ( P3_ADD_546_U124 , P3_ADD_546_U27 );
not NOT1_18581 ( P3_ADD_546_U125 , P3_ADD_546_U95 );
not NOT1_18582 ( P3_ADD_546_U126 , P3_ADD_546_U96 );
not NOT1_18583 ( P3_ADD_546_U127 , P3_ADD_546_U97 );
not NOT1_18584 ( P3_ADD_546_U128 , P3_ADD_546_U49 );
not NOT1_18585 ( P3_ADD_546_U129 , P3_ADD_546_U99 );
not NOT1_18586 ( P3_ADD_546_U130 , P3_ADD_546_U100 );
not NOT1_18587 ( P3_ADD_546_U131 , P3_ADD_546_U101 );
not NOT1_18588 ( P3_ADD_546_U132 , P3_ADD_546_U102 );
not NOT1_18589 ( P3_ADD_546_U133 , P3_ADD_546_U103 );
not NOT1_18590 ( P3_ADD_546_U134 , P3_ADD_546_U104 );
not NOT1_18591 ( P3_ADD_546_U135 , P3_ADD_546_U105 );
not NOT1_18592 ( P3_ADD_546_U136 , P3_ADD_546_U106 );
not NOT1_18593 ( P3_ADD_546_U137 , P3_ADD_546_U107 );
not NOT1_18594 ( P3_ADD_546_U138 , P3_ADD_546_U108 );
not NOT1_18595 ( P3_ADD_546_U139 , P3_ADD_546_U109 );
not NOT1_18596 ( P3_ADD_546_U140 , P3_ADD_546_U110 );
nand NAND2_18597 ( P3_ADD_546_U141 , P3_ADD_546_U120 , P3_ADD_546_U18 );
nand NAND2_18598 ( P3_ADD_546_U142 , P3_EAX_REG_9_ , P3_ADD_546_U17 );
nand NAND2_18599 ( P3_ADD_546_U143 , P3_EAX_REG_8_ , P3_ADD_546_U95 );
nand NAND2_18600 ( P3_ADD_546_U144 , P3_ADD_546_U125 , P3_ADD_546_U14 );
nand NAND2_18601 ( P3_ADD_546_U145 , P3_ADD_546_U118 , P3_ADD_546_U15 );
nand NAND2_18602 ( P3_ADD_546_U146 , P3_EAX_REG_7_ , P3_ADD_546_U16 );
nand NAND2_18603 ( P3_ADD_546_U147 , P3_EAX_REG_6_ , P3_ADD_546_U96 );
nand NAND2_18604 ( P3_ADD_546_U148 , P3_ADD_546_U126 , P3_ADD_546_U11 );
nand NAND2_18605 ( P3_ADD_546_U149 , P3_ADD_546_U112 , P3_ADD_546_U12 );
nand NAND2_18606 ( P3_ADD_546_U150 , P3_EAX_REG_5_ , P3_ADD_546_U13 );
nand NAND2_18607 ( P3_ADD_546_U151 , P3_EAX_REG_4_ , P3_ADD_546_U97 );
nand NAND2_18608 ( P3_ADD_546_U152 , P3_ADD_546_U127 , P3_ADD_546_U8 );
nand NAND2_18609 ( P3_ADD_546_U153 , P3_ADD_546_U111 , P3_ADD_546_U9 );
nand NAND2_18610 ( P3_ADD_546_U154 , P3_EAX_REG_3_ , P3_ADD_546_U10 );
nand NAND2_18611 ( P3_ADD_546_U155 , P3_EAX_REG_31_ , P3_ADD_546_U99 );
nand NAND2_18612 ( P3_ADD_546_U156 , P3_ADD_546_U129 , P3_ADD_546_U98 );
nand NAND2_18613 ( P3_ADD_546_U157 , P3_EAX_REG_30_ , P3_ADD_546_U49 );
nand NAND2_18614 ( P3_ADD_546_U158 , P3_ADD_546_U128 , P3_ADD_546_U50 );
nand NAND2_18615 ( P3_ADD_546_U159 , P3_EAX_REG_2_ , P3_ADD_546_U100 );
nand NAND2_18616 ( P3_ADD_546_U160 , P3_ADD_546_U130 , P3_ADD_546_U6 );
nand NAND2_18617 ( P3_ADD_546_U161 , P3_ADD_546_U123 , P3_ADD_546_U47 );
nand NAND2_18618 ( P3_ADD_546_U162 , P3_EAX_REG_29_ , P3_ADD_546_U48 );
nand NAND2_18619 ( P3_ADD_546_U163 , P3_EAX_REG_28_ , P3_ADD_546_U101 );
nand NAND2_18620 ( P3_ADD_546_U164 , P3_ADD_546_U131 , P3_ADD_546_U45 );
nand NAND2_18621 ( P3_ADD_546_U165 , P3_ADD_546_U122 , P3_ADD_546_U44 );
nand NAND2_18622 ( P3_ADD_546_U166 , P3_EAX_REG_27_ , P3_ADD_546_U46 );
nand NAND2_18623 ( P3_ADD_546_U167 , P3_EAX_REG_26_ , P3_ADD_546_U102 );
nand NAND2_18624 ( P3_ADD_546_U168 , P3_ADD_546_U132 , P3_ADD_546_U41 );
nand NAND2_18625 ( P3_ADD_546_U169 , P3_ADD_546_U116 , P3_ADD_546_U42 );
nand NAND2_18626 ( P3_ADD_546_U170 , P3_EAX_REG_25_ , P3_ADD_546_U43 );
nand NAND2_18627 ( P3_ADD_546_U171 , P3_EAX_REG_24_ , P3_ADD_546_U103 );
nand NAND2_18628 ( P3_ADD_546_U172 , P3_ADD_546_U133 , P3_ADD_546_U38 );
nand NAND2_18629 ( P3_ADD_546_U173 , P3_ADD_546_U115 , P3_ADD_546_U39 );
nand NAND2_18630 ( P3_ADD_546_U174 , P3_EAX_REG_23_ , P3_ADD_546_U40 );
nand NAND2_18631 ( P3_ADD_546_U175 , P3_EAX_REG_22_ , P3_ADD_546_U104 );
nand NAND2_18632 ( P3_ADD_546_U176 , P3_ADD_546_U134 , P3_ADD_546_U37 );
nand NAND2_18633 ( P3_ADD_546_U177 , P3_ADD_546_U121 , P3_ADD_546_U35 );
nand NAND2_18634 ( P3_ADD_546_U178 , P3_EAX_REG_21_ , P3_ADD_546_U36 );
nand NAND2_18635 ( P3_ADD_546_U179 , P3_EAX_REG_20_ , P3_ADD_546_U105 );
nand NAND2_18636 ( P3_ADD_546_U180 , P3_ADD_546_U135 , P3_ADD_546_U32 );
nand NAND2_18637 ( P3_ADD_546_U181 , P3_EAX_REG_0_ , P3_ADD_546_U7 );
nand NAND2_18638 ( P3_ADD_546_U182 , P3_EAX_REG_1_ , P3_ADD_546_U5 );
nand NAND2_18639 ( P3_ADD_546_U183 , P3_ADD_546_U114 , P3_ADD_546_U33 );
nand NAND2_18640 ( P3_ADD_546_U184 , P3_EAX_REG_19_ , P3_ADD_546_U34 );
nand NAND2_18641 ( P3_ADD_546_U185 , P3_EAX_REG_18_ , P3_ADD_546_U106 );
nand NAND2_18642 ( P3_ADD_546_U186 , P3_ADD_546_U136 , P3_ADD_546_U29 );
nand NAND2_18643 ( P3_ADD_546_U187 , P3_ADD_546_U117 , P3_ADD_546_U30 );
nand NAND2_18644 ( P3_ADD_546_U188 , P3_EAX_REG_17_ , P3_ADD_546_U31 );
nand NAND2_18645 ( P3_ADD_546_U189 , P3_EAX_REG_16_ , P3_ADD_546_U107 );
nand NAND2_18646 ( P3_ADD_546_U190 , P3_ADD_546_U137 , P3_ADD_546_U28 );
nand NAND2_18647 ( P3_ADD_546_U191 , P3_ADD_546_U124 , P3_ADD_546_U26 );
nand NAND2_18648 ( P3_ADD_546_U192 , P3_EAX_REG_15_ , P3_ADD_546_U27 );
nand NAND2_18649 ( P3_ADD_546_U193 , P3_EAX_REG_14_ , P3_ADD_546_U108 );
nand NAND2_18650 ( P3_ADD_546_U194 , P3_ADD_546_U138 , P3_ADD_546_U23 );
nand NAND2_18651 ( P3_ADD_546_U195 , P3_ADD_546_U119 , P3_ADD_546_U24 );
nand NAND2_18652 ( P3_ADD_546_U196 , P3_EAX_REG_13_ , P3_ADD_546_U25 );
nand NAND2_18653 ( P3_ADD_546_U197 , P3_EAX_REG_12_ , P3_ADD_546_U109 );
nand NAND2_18654 ( P3_ADD_546_U198 , P3_ADD_546_U139 , P3_ADD_546_U20 );
nand NAND2_18655 ( P3_ADD_546_U199 , P3_ADD_546_U113 , P3_ADD_546_U21 );
nand NAND2_18656 ( P3_ADD_546_U200 , P3_EAX_REG_11_ , P3_ADD_546_U22 );
nand NAND2_18657 ( P3_ADD_546_U201 , P3_EAX_REG_10_ , P3_ADD_546_U110 );
nand NAND2_18658 ( P3_ADD_546_U202 , P3_ADD_546_U140 , P3_ADD_546_U19 );
nor nor_18659 ( P3_GTE_401_U6 , P3_SUB_401_U6 , P3_GTE_401_U8 );
and AND2_18660 ( P3_GTE_401_U7 , P3_SUB_401_U21 , P3_GTE_401_U9 );
nor nor_18661 ( P3_GTE_401_U8 , P3_SUB_401_U19 , P3_SUB_401_U20 , P3_GTE_401_U7 );
or OR2_18662 ( P3_GTE_401_U9 , P3_SUB_401_U7 , P3_SUB_401_U22 );
not NOT1_18663 ( P3_ADD_391_1180_U4 , P3_U2613 );
not NOT1_18664 ( P3_ADD_391_1180_U5 , P3_U3069 );
nand NAND2_18665 ( P3_ADD_391_1180_U6 , P3_U3069 , P3_U2613 );
not NOT1_18666 ( P3_ADD_391_1180_U7 , P3_U2614 );
nand NAND2_18667 ( P3_ADD_391_1180_U8 , P3_U2614 , P3_ADD_391_1180_U28 );
not NOT1_18668 ( P3_ADD_391_1180_U9 , P3_U2615 );
nand NAND2_18669 ( P3_ADD_391_1180_U10 , P3_U2615 , P3_ADD_391_1180_U29 );
not NOT1_18670 ( P3_ADD_391_1180_U11 , P3_U2616 );
nand NAND2_18671 ( P3_ADD_391_1180_U12 , P3_U2616 , P3_ADD_391_1180_U30 );
not NOT1_18672 ( P3_ADD_391_1180_U13 , P3_U2617 );
nand NAND2_18673 ( P3_ADD_391_1180_U14 , P3_U2617 , P3_ADD_391_1180_U31 );
not NOT1_18674 ( P3_ADD_391_1180_U15 , P3_U2618 );
nand NAND2_18675 ( P3_ADD_391_1180_U16 , P3_U2618 , P3_ADD_391_1180_U32 );
not NOT1_18676 ( P3_ADD_391_1180_U17 , P3_U2619 );
nand NAND2_18677 ( P3_ADD_391_1180_U18 , P3_ADD_391_1180_U36 , P3_ADD_391_1180_U35 );
nand NAND2_18678 ( P3_ADD_391_1180_U19 , P3_ADD_391_1180_U38 , P3_ADD_391_1180_U37 );
nand NAND2_18679 ( P3_ADD_391_1180_U20 , P3_ADD_391_1180_U40 , P3_ADD_391_1180_U39 );
nand NAND2_18680 ( P3_ADD_391_1180_U21 , P3_ADD_391_1180_U42 , P3_ADD_391_1180_U41 );
nand NAND2_18681 ( P3_ADD_391_1180_U22 , P3_ADD_391_1180_U44 , P3_ADD_391_1180_U43 );
nand NAND2_18682 ( P3_ADD_391_1180_U23 , P3_ADD_391_1180_U46 , P3_ADD_391_1180_U45 );
nand NAND2_18683 ( P3_ADD_391_1180_U24 , P3_ADD_391_1180_U48 , P3_ADD_391_1180_U47 );
nand NAND2_18684 ( P3_ADD_391_1180_U25 , P3_ADD_391_1180_U50 , P3_ADD_391_1180_U49 );
not NOT1_18685 ( P3_ADD_391_1180_U26 , P3_U2620 );
nand NAND2_18686 ( P3_ADD_391_1180_U27 , P3_U2619 , P3_ADD_391_1180_U33 );
not NOT1_18687 ( P3_ADD_391_1180_U28 , P3_ADD_391_1180_U6 );
not NOT1_18688 ( P3_ADD_391_1180_U29 , P3_ADD_391_1180_U8 );
not NOT1_18689 ( P3_ADD_391_1180_U30 , P3_ADD_391_1180_U10 );
not NOT1_18690 ( P3_ADD_391_1180_U31 , P3_ADD_391_1180_U12 );
not NOT1_18691 ( P3_ADD_391_1180_U32 , P3_ADD_391_1180_U14 );
not NOT1_18692 ( P3_ADD_391_1180_U33 , P3_ADD_391_1180_U16 );
not NOT1_18693 ( P3_ADD_391_1180_U34 , P3_ADD_391_1180_U27 );
nand NAND2_18694 ( P3_ADD_391_1180_U35 , P3_U2620 , P3_ADD_391_1180_U27 );
nand NAND2_18695 ( P3_ADD_391_1180_U36 , P3_ADD_391_1180_U34 , P3_ADD_391_1180_U26 );
nand NAND2_18696 ( P3_ADD_391_1180_U37 , P3_U2619 , P3_ADD_391_1180_U16 );
nand NAND2_18697 ( P3_ADD_391_1180_U38 , P3_ADD_391_1180_U33 , P3_ADD_391_1180_U17 );
nand NAND2_18698 ( P3_ADD_391_1180_U39 , P3_U2618 , P3_ADD_391_1180_U14 );
nand NAND2_18699 ( P3_ADD_391_1180_U40 , P3_ADD_391_1180_U32 , P3_ADD_391_1180_U15 );
nand NAND2_18700 ( P3_ADD_391_1180_U41 , P3_U2617 , P3_ADD_391_1180_U12 );
nand NAND2_18701 ( P3_ADD_391_1180_U42 , P3_ADD_391_1180_U31 , P3_ADD_391_1180_U13 );
nand NAND2_18702 ( P3_ADD_391_1180_U43 , P3_U2616 , P3_ADD_391_1180_U10 );
nand NAND2_18703 ( P3_ADD_391_1180_U44 , P3_ADD_391_1180_U30 , P3_ADD_391_1180_U11 );
nand NAND2_18704 ( P3_ADD_391_1180_U45 , P3_U2615 , P3_ADD_391_1180_U8 );
nand NAND2_18705 ( P3_ADD_391_1180_U46 , P3_ADD_391_1180_U29 , P3_ADD_391_1180_U9 );
nand NAND2_18706 ( P3_ADD_391_1180_U47 , P3_U2614 , P3_ADD_391_1180_U6 );
nand NAND2_18707 ( P3_ADD_391_1180_U48 , P3_ADD_391_1180_U28 , P3_ADD_391_1180_U7 );
nand NAND2_18708 ( P3_ADD_391_1180_U49 , P3_U3069 , P3_ADD_391_1180_U4 );
nand NAND2_18709 ( P3_ADD_391_1180_U50 , P3_U2613 , P3_ADD_391_1180_U5 );
not NOT1_18710 ( P3_ADD_476_U4 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_18711 ( P3_ADD_476_U5 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_18712 ( P3_ADD_476_U6 , P3_INSTADDRPOINTER_REG_2_ , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_18713 ( P3_ADD_476_U7 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_18714 ( P3_ADD_476_U8 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_476_U94 );
not NOT1_18715 ( P3_ADD_476_U9 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_18716 ( P3_ADD_476_U10 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_476_U95 );
not NOT1_18717 ( P3_ADD_476_U11 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_18718 ( P3_ADD_476_U12 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_476_U96 );
not NOT1_18719 ( P3_ADD_476_U13 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_18720 ( P3_ADD_476_U14 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_476_U97 );
not NOT1_18721 ( P3_ADD_476_U15 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_18722 ( P3_ADD_476_U16 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_476_U98 );
not NOT1_18723 ( P3_ADD_476_U17 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_18724 ( P3_ADD_476_U18 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_18725 ( P3_ADD_476_U19 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_476_U99 );
nand NAND2_18726 ( P3_ADD_476_U20 , P3_ADD_476_U100 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_18727 ( P3_ADD_476_U21 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_18728 ( P3_ADD_476_U22 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_476_U101 );
not NOT1_18729 ( P3_ADD_476_U23 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_18730 ( P3_ADD_476_U24 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_476_U102 );
not NOT1_18731 ( P3_ADD_476_U25 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_18732 ( P3_ADD_476_U26 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_476_U103 );
not NOT1_18733 ( P3_ADD_476_U27 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_18734 ( P3_ADD_476_U28 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_476_U104 );
not NOT1_18735 ( P3_ADD_476_U29 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_18736 ( P3_ADD_476_U30 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_476_U105 );
not NOT1_18737 ( P3_ADD_476_U31 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_18738 ( P3_ADD_476_U32 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_476_U106 );
not NOT1_18739 ( P3_ADD_476_U33 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_18740 ( P3_ADD_476_U34 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_476_U107 );
not NOT1_18741 ( P3_ADD_476_U35 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_18742 ( P3_ADD_476_U36 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_476_U108 );
not NOT1_18743 ( P3_ADD_476_U37 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_18744 ( P3_ADD_476_U38 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_476_U109 );
not NOT1_18745 ( P3_ADD_476_U39 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_18746 ( P3_ADD_476_U40 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_476_U110 );
not NOT1_18747 ( P3_ADD_476_U41 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_18748 ( P3_ADD_476_U42 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_476_U111 );
not NOT1_18749 ( P3_ADD_476_U43 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_18750 ( P3_ADD_476_U44 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_476_U112 );
not NOT1_18751 ( P3_ADD_476_U45 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_18752 ( P3_ADD_476_U46 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_476_U113 );
not NOT1_18753 ( P3_ADD_476_U47 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_18754 ( P3_ADD_476_U48 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_476_U114 );
not NOT1_18755 ( P3_ADD_476_U49 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_18756 ( P3_ADD_476_U50 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_476_U115 );
not NOT1_18757 ( P3_ADD_476_U51 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_18758 ( P3_ADD_476_U52 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_476_U116 );
not NOT1_18759 ( P3_ADD_476_U53 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_18760 ( P3_ADD_476_U54 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_476_U117 );
not NOT1_18761 ( P3_ADD_476_U55 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_18762 ( P3_ADD_476_U56 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_476_U118 );
not NOT1_18763 ( P3_ADD_476_U57 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_18764 ( P3_ADD_476_U58 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_476_U119 );
not NOT1_18765 ( P3_ADD_476_U59 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_18766 ( P3_ADD_476_U60 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_476_U120 );
not NOT1_18767 ( P3_ADD_476_U61 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_18768 ( P3_ADD_476_U62 , P3_ADD_476_U124 , P3_ADD_476_U123 );
nand NAND2_18769 ( P3_ADD_476_U63 , P3_ADD_476_U126 , P3_ADD_476_U125 );
nand NAND2_18770 ( P3_ADD_476_U64 , P3_ADD_476_U128 , P3_ADD_476_U127 );
nand NAND2_18771 ( P3_ADD_476_U65 , P3_ADD_476_U130 , P3_ADD_476_U129 );
nand NAND2_18772 ( P3_ADD_476_U66 , P3_ADD_476_U132 , P3_ADD_476_U131 );
nand NAND2_18773 ( P3_ADD_476_U67 , P3_ADD_476_U134 , P3_ADD_476_U133 );
nand NAND2_18774 ( P3_ADD_476_U68 , P3_ADD_476_U136 , P3_ADD_476_U135 );
nand NAND2_18775 ( P3_ADD_476_U69 , P3_ADD_476_U138 , P3_ADD_476_U137 );
nand NAND2_18776 ( P3_ADD_476_U70 , P3_ADD_476_U140 , P3_ADD_476_U139 );
nand NAND2_18777 ( P3_ADD_476_U71 , P3_ADD_476_U142 , P3_ADD_476_U141 );
nand NAND2_18778 ( P3_ADD_476_U72 , P3_ADD_476_U144 , P3_ADD_476_U143 );
nand NAND2_18779 ( P3_ADD_476_U73 , P3_ADD_476_U146 , P3_ADD_476_U145 );
nand NAND2_18780 ( P3_ADD_476_U74 , P3_ADD_476_U148 , P3_ADD_476_U147 );
nand NAND2_18781 ( P3_ADD_476_U75 , P3_ADD_476_U150 , P3_ADD_476_U149 );
nand NAND2_18782 ( P3_ADD_476_U76 , P3_ADD_476_U152 , P3_ADD_476_U151 );
nand NAND2_18783 ( P3_ADD_476_U77 , P3_ADD_476_U154 , P3_ADD_476_U153 );
nand NAND2_18784 ( P3_ADD_476_U78 , P3_ADD_476_U156 , P3_ADD_476_U155 );
nand NAND2_18785 ( P3_ADD_476_U79 , P3_ADD_476_U158 , P3_ADD_476_U157 );
nand NAND2_18786 ( P3_ADD_476_U80 , P3_ADD_476_U160 , P3_ADD_476_U159 );
nand NAND2_18787 ( P3_ADD_476_U81 , P3_ADD_476_U162 , P3_ADD_476_U161 );
nand NAND2_18788 ( P3_ADD_476_U82 , P3_ADD_476_U164 , P3_ADD_476_U163 );
nand NAND2_18789 ( P3_ADD_476_U83 , P3_ADD_476_U166 , P3_ADD_476_U165 );
nand NAND2_18790 ( P3_ADD_476_U84 , P3_ADD_476_U168 , P3_ADD_476_U167 );
nand NAND2_18791 ( P3_ADD_476_U85 , P3_ADD_476_U170 , P3_ADD_476_U169 );
nand NAND2_18792 ( P3_ADD_476_U86 , P3_ADD_476_U172 , P3_ADD_476_U171 );
nand NAND2_18793 ( P3_ADD_476_U87 , P3_ADD_476_U174 , P3_ADD_476_U173 );
nand NAND2_18794 ( P3_ADD_476_U88 , P3_ADD_476_U176 , P3_ADD_476_U175 );
nand NAND2_18795 ( P3_ADD_476_U89 , P3_ADD_476_U178 , P3_ADD_476_U177 );
nand NAND2_18796 ( P3_ADD_476_U90 , P3_ADD_476_U180 , P3_ADD_476_U179 );
nand NAND2_18797 ( P3_ADD_476_U91 , P3_ADD_476_U182 , P3_ADD_476_U181 );
not NOT1_18798 ( P3_ADD_476_U92 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_18799 ( P3_ADD_476_U93 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_476_U121 );
not NOT1_18800 ( P3_ADD_476_U94 , P3_ADD_476_U6 );
not NOT1_18801 ( P3_ADD_476_U95 , P3_ADD_476_U8 );
not NOT1_18802 ( P3_ADD_476_U96 , P3_ADD_476_U10 );
not NOT1_18803 ( P3_ADD_476_U97 , P3_ADD_476_U12 );
not NOT1_18804 ( P3_ADD_476_U98 , P3_ADD_476_U14 );
not NOT1_18805 ( P3_ADD_476_U99 , P3_ADD_476_U16 );
not NOT1_18806 ( P3_ADD_476_U100 , P3_ADD_476_U19 );
not NOT1_18807 ( P3_ADD_476_U101 , P3_ADD_476_U20 );
not NOT1_18808 ( P3_ADD_476_U102 , P3_ADD_476_U22 );
not NOT1_18809 ( P3_ADD_476_U103 , P3_ADD_476_U24 );
not NOT1_18810 ( P3_ADD_476_U104 , P3_ADD_476_U26 );
not NOT1_18811 ( P3_ADD_476_U105 , P3_ADD_476_U28 );
not NOT1_18812 ( P3_ADD_476_U106 , P3_ADD_476_U30 );
not NOT1_18813 ( P3_ADD_476_U107 , P3_ADD_476_U32 );
not NOT1_18814 ( P3_ADD_476_U108 , P3_ADD_476_U34 );
not NOT1_18815 ( P3_ADD_476_U109 , P3_ADD_476_U36 );
not NOT1_18816 ( P3_ADD_476_U110 , P3_ADD_476_U38 );
not NOT1_18817 ( P3_ADD_476_U111 , P3_ADD_476_U40 );
not NOT1_18818 ( P3_ADD_476_U112 , P3_ADD_476_U42 );
not NOT1_18819 ( P3_ADD_476_U113 , P3_ADD_476_U44 );
not NOT1_18820 ( P3_ADD_476_U114 , P3_ADD_476_U46 );
not NOT1_18821 ( P3_ADD_476_U115 , P3_ADD_476_U48 );
not NOT1_18822 ( P3_ADD_476_U116 , P3_ADD_476_U50 );
not NOT1_18823 ( P3_ADD_476_U117 , P3_ADD_476_U52 );
not NOT1_18824 ( P3_ADD_476_U118 , P3_ADD_476_U54 );
not NOT1_18825 ( P3_ADD_476_U119 , P3_ADD_476_U56 );
not NOT1_18826 ( P3_ADD_476_U120 , P3_ADD_476_U58 );
not NOT1_18827 ( P3_ADD_476_U121 , P3_ADD_476_U60 );
not NOT1_18828 ( P3_ADD_476_U122 , P3_ADD_476_U93 );
nand NAND2_18829 ( P3_ADD_476_U123 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_476_U19 );
nand NAND2_18830 ( P3_ADD_476_U124 , P3_ADD_476_U100 , P3_ADD_476_U18 );
nand NAND2_18831 ( P3_ADD_476_U125 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_476_U16 );
nand NAND2_18832 ( P3_ADD_476_U126 , P3_ADD_476_U99 , P3_ADD_476_U17 );
nand NAND2_18833 ( P3_ADD_476_U127 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_476_U14 );
nand NAND2_18834 ( P3_ADD_476_U128 , P3_ADD_476_U98 , P3_ADD_476_U15 );
nand NAND2_18835 ( P3_ADD_476_U129 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_476_U12 );
nand NAND2_18836 ( P3_ADD_476_U130 , P3_ADD_476_U97 , P3_ADD_476_U13 );
nand NAND2_18837 ( P3_ADD_476_U131 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_476_U10 );
nand NAND2_18838 ( P3_ADD_476_U132 , P3_ADD_476_U96 , P3_ADD_476_U11 );
nand NAND2_18839 ( P3_ADD_476_U133 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_476_U8 );
nand NAND2_18840 ( P3_ADD_476_U134 , P3_ADD_476_U95 , P3_ADD_476_U9 );
nand NAND2_18841 ( P3_ADD_476_U135 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_476_U6 );
nand NAND2_18842 ( P3_ADD_476_U136 , P3_ADD_476_U94 , P3_ADD_476_U7 );
nand NAND2_18843 ( P3_ADD_476_U137 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_476_U93 );
nand NAND2_18844 ( P3_ADD_476_U138 , P3_ADD_476_U122 , P3_ADD_476_U92 );
nand NAND2_18845 ( P3_ADD_476_U139 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_476_U60 );
nand NAND2_18846 ( P3_ADD_476_U140 , P3_ADD_476_U121 , P3_ADD_476_U61 );
nand NAND2_18847 ( P3_ADD_476_U141 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_476_U4 );
nand NAND2_18848 ( P3_ADD_476_U142 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_476_U5 );
nand NAND2_18849 ( P3_ADD_476_U143 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_476_U58 );
nand NAND2_18850 ( P3_ADD_476_U144 , P3_ADD_476_U120 , P3_ADD_476_U59 );
nand NAND2_18851 ( P3_ADD_476_U145 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_476_U56 );
nand NAND2_18852 ( P3_ADD_476_U146 , P3_ADD_476_U119 , P3_ADD_476_U57 );
nand NAND2_18853 ( P3_ADD_476_U147 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_476_U54 );
nand NAND2_18854 ( P3_ADD_476_U148 , P3_ADD_476_U118 , P3_ADD_476_U55 );
nand NAND2_18855 ( P3_ADD_476_U149 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_476_U52 );
nand NAND2_18856 ( P3_ADD_476_U150 , P3_ADD_476_U117 , P3_ADD_476_U53 );
nand NAND2_18857 ( P3_ADD_476_U151 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_476_U50 );
nand NAND2_18858 ( P3_ADD_476_U152 , P3_ADD_476_U116 , P3_ADD_476_U51 );
nand NAND2_18859 ( P3_ADD_476_U153 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_476_U48 );
nand NAND2_18860 ( P3_ADD_476_U154 , P3_ADD_476_U115 , P3_ADD_476_U49 );
nand NAND2_18861 ( P3_ADD_476_U155 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_476_U46 );
nand NAND2_18862 ( P3_ADD_476_U156 , P3_ADD_476_U114 , P3_ADD_476_U47 );
nand NAND2_18863 ( P3_ADD_476_U157 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_476_U44 );
nand NAND2_18864 ( P3_ADD_476_U158 , P3_ADD_476_U113 , P3_ADD_476_U45 );
nand NAND2_18865 ( P3_ADD_476_U159 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_476_U42 );
nand NAND2_18866 ( P3_ADD_476_U160 , P3_ADD_476_U112 , P3_ADD_476_U43 );
nand NAND2_18867 ( P3_ADD_476_U161 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_476_U40 );
nand NAND2_18868 ( P3_ADD_476_U162 , P3_ADD_476_U111 , P3_ADD_476_U41 );
nand NAND2_18869 ( P3_ADD_476_U163 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_476_U38 );
nand NAND2_18870 ( P3_ADD_476_U164 , P3_ADD_476_U110 , P3_ADD_476_U39 );
nand NAND2_18871 ( P3_ADD_476_U165 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_476_U36 );
nand NAND2_18872 ( P3_ADD_476_U166 , P3_ADD_476_U109 , P3_ADD_476_U37 );
nand NAND2_18873 ( P3_ADD_476_U167 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_476_U34 );
nand NAND2_18874 ( P3_ADD_476_U168 , P3_ADD_476_U108 , P3_ADD_476_U35 );
nand NAND2_18875 ( P3_ADD_476_U169 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_476_U32 );
nand NAND2_18876 ( P3_ADD_476_U170 , P3_ADD_476_U107 , P3_ADD_476_U33 );
nand NAND2_18877 ( P3_ADD_476_U171 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_476_U30 );
nand NAND2_18878 ( P3_ADD_476_U172 , P3_ADD_476_U106 , P3_ADD_476_U31 );
nand NAND2_18879 ( P3_ADD_476_U173 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_476_U28 );
nand NAND2_18880 ( P3_ADD_476_U174 , P3_ADD_476_U105 , P3_ADD_476_U29 );
nand NAND2_18881 ( P3_ADD_476_U175 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_476_U26 );
nand NAND2_18882 ( P3_ADD_476_U176 , P3_ADD_476_U104 , P3_ADD_476_U27 );
nand NAND2_18883 ( P3_ADD_476_U177 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_476_U24 );
nand NAND2_18884 ( P3_ADD_476_U178 , P3_ADD_476_U103 , P3_ADD_476_U25 );
nand NAND2_18885 ( P3_ADD_476_U179 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_476_U22 );
nand NAND2_18886 ( P3_ADD_476_U180 , P3_ADD_476_U102 , P3_ADD_476_U23 );
nand NAND2_18887 ( P3_ADD_476_U181 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_476_U20 );
nand NAND2_18888 ( P3_ADD_476_U182 , P3_ADD_476_U101 , P3_ADD_476_U21 );
nor nor_18889 ( P3_GTE_390_U6 , P3_SUB_390_U6 , P3_GTE_390_U8 );
and AND2_18890 ( P3_GTE_390_U7 , P3_SUB_390_U21 , P3_GTE_390_U9 );
nor nor_18891 ( P3_GTE_390_U8 , P3_SUB_390_U19 , P3_SUB_390_U20 , P3_GTE_390_U7 );
or OR2_18892 ( P3_GTE_390_U9 , P3_SUB_390_U7 , P3_SUB_390_U22 );
not NOT1_18893 ( P3_ADD_531_U5 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_18894 ( P3_ADD_531_U6 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_18895 ( P3_ADD_531_U7 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_18896 ( P3_ADD_531_U8 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_18897 ( P3_ADD_531_U9 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_531_U98 );
not NOT1_18898 ( P3_ADD_531_U10 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_18899 ( P3_ADD_531_U11 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_531_U99 );
not NOT1_18900 ( P3_ADD_531_U12 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_18901 ( P3_ADD_531_U13 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_531_U100 );
not NOT1_18902 ( P3_ADD_531_U14 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_18903 ( P3_ADD_531_U15 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_531_U101 );
not NOT1_18904 ( P3_ADD_531_U16 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_18905 ( P3_ADD_531_U17 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_531_U102 );
not NOT1_18906 ( P3_ADD_531_U18 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_18907 ( P3_ADD_531_U19 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_531_U103 );
not NOT1_18908 ( P3_ADD_531_U20 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_18909 ( P3_ADD_531_U21 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_18910 ( P3_ADD_531_U22 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_531_U104 );
nand NAND2_18911 ( P3_ADD_531_U23 , P3_ADD_531_U105 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_18912 ( P3_ADD_531_U24 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_18913 ( P3_ADD_531_U25 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_531_U106 );
not NOT1_18914 ( P3_ADD_531_U26 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_18915 ( P3_ADD_531_U27 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_531_U107 );
not NOT1_18916 ( P3_ADD_531_U28 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_18917 ( P3_ADD_531_U29 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_531_U108 );
not NOT1_18918 ( P3_ADD_531_U30 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_18919 ( P3_ADD_531_U31 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_531_U109 );
not NOT1_18920 ( P3_ADD_531_U32 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_18921 ( P3_ADD_531_U33 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_531_U110 );
not NOT1_18922 ( P3_ADD_531_U34 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_18923 ( P3_ADD_531_U35 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_531_U111 );
not NOT1_18924 ( P3_ADD_531_U36 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_18925 ( P3_ADD_531_U37 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_531_U112 );
not NOT1_18926 ( P3_ADD_531_U38 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_18927 ( P3_ADD_531_U39 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_531_U113 );
not NOT1_18928 ( P3_ADD_531_U40 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_18929 ( P3_ADD_531_U41 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_531_U114 );
not NOT1_18930 ( P3_ADD_531_U42 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_18931 ( P3_ADD_531_U43 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_531_U115 );
not NOT1_18932 ( P3_ADD_531_U44 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_18933 ( P3_ADD_531_U45 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_531_U116 );
not NOT1_18934 ( P3_ADD_531_U46 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_18935 ( P3_ADD_531_U47 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_531_U117 );
not NOT1_18936 ( P3_ADD_531_U48 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_18937 ( P3_ADD_531_U49 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_531_U118 );
not NOT1_18938 ( P3_ADD_531_U50 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_18939 ( P3_ADD_531_U51 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_531_U119 );
not NOT1_18940 ( P3_ADD_531_U52 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_18941 ( P3_ADD_531_U53 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_531_U120 );
not NOT1_18942 ( P3_ADD_531_U54 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_18943 ( P3_ADD_531_U55 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_531_U121 );
not NOT1_18944 ( P3_ADD_531_U56 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_18945 ( P3_ADD_531_U57 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_531_U122 );
not NOT1_18946 ( P3_ADD_531_U58 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_18947 ( P3_ADD_531_U59 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_531_U123 );
not NOT1_18948 ( P3_ADD_531_U60 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_18949 ( P3_ADD_531_U61 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_531_U124 );
not NOT1_18950 ( P3_ADD_531_U62 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_18951 ( P3_ADD_531_U63 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_531_U125 );
not NOT1_18952 ( P3_ADD_531_U64 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_18953 ( P3_ADD_531_U65 , P3_ADD_531_U129 , P3_ADD_531_U128 );
nand NAND2_18954 ( P3_ADD_531_U66 , P3_ADD_531_U131 , P3_ADD_531_U130 );
nand NAND2_18955 ( P3_ADD_531_U67 , P3_ADD_531_U133 , P3_ADD_531_U132 );
nand NAND2_18956 ( P3_ADD_531_U68 , P3_ADD_531_U135 , P3_ADD_531_U134 );
nand NAND2_18957 ( P3_ADD_531_U69 , P3_ADD_531_U137 , P3_ADD_531_U136 );
nand NAND2_18958 ( P3_ADD_531_U70 , P3_ADD_531_U139 , P3_ADD_531_U138 );
nand NAND2_18959 ( P3_ADD_531_U71 , P3_ADD_531_U141 , P3_ADD_531_U140 );
nand NAND2_18960 ( P3_ADD_531_U72 , P3_ADD_531_U143 , P3_ADD_531_U142 );
nand NAND2_18961 ( P3_ADD_531_U73 , P3_ADD_531_U145 , P3_ADD_531_U144 );
nand NAND2_18962 ( P3_ADD_531_U74 , P3_ADD_531_U147 , P3_ADD_531_U146 );
nand NAND2_18963 ( P3_ADD_531_U75 , P3_ADD_531_U149 , P3_ADD_531_U148 );
nand NAND2_18964 ( P3_ADD_531_U76 , P3_ADD_531_U151 , P3_ADD_531_U150 );
nand NAND2_18965 ( P3_ADD_531_U77 , P3_ADD_531_U153 , P3_ADD_531_U152 );
nand NAND2_18966 ( P3_ADD_531_U78 , P3_ADD_531_U155 , P3_ADD_531_U154 );
nand NAND2_18967 ( P3_ADD_531_U79 , P3_ADD_531_U157 , P3_ADD_531_U156 );
nand NAND2_18968 ( P3_ADD_531_U80 , P3_ADD_531_U159 , P3_ADD_531_U158 );
nand NAND2_18969 ( P3_ADD_531_U81 , P3_ADD_531_U161 , P3_ADD_531_U160 );
nand NAND2_18970 ( P3_ADD_531_U82 , P3_ADD_531_U163 , P3_ADD_531_U162 );
nand NAND2_18971 ( P3_ADD_531_U83 , P3_ADD_531_U165 , P3_ADD_531_U164 );
nand NAND2_18972 ( P3_ADD_531_U84 , P3_ADD_531_U167 , P3_ADD_531_U166 );
nand NAND2_18973 ( P3_ADD_531_U85 , P3_ADD_531_U169 , P3_ADD_531_U168 );
nand NAND2_18974 ( P3_ADD_531_U86 , P3_ADD_531_U171 , P3_ADD_531_U170 );
nand NAND2_18975 ( P3_ADD_531_U87 , P3_ADD_531_U173 , P3_ADD_531_U172 );
nand NAND2_18976 ( P3_ADD_531_U88 , P3_ADD_531_U175 , P3_ADD_531_U174 );
nand NAND2_18977 ( P3_ADD_531_U89 , P3_ADD_531_U177 , P3_ADD_531_U176 );
nand NAND2_18978 ( P3_ADD_531_U90 , P3_ADD_531_U179 , P3_ADD_531_U178 );
nand NAND2_18979 ( P3_ADD_531_U91 , P3_ADD_531_U181 , P3_ADD_531_U180 );
nand NAND2_18980 ( P3_ADD_531_U92 , P3_ADD_531_U183 , P3_ADD_531_U182 );
nand NAND2_18981 ( P3_ADD_531_U93 , P3_ADD_531_U185 , P3_ADD_531_U184 );
nand NAND2_18982 ( P3_ADD_531_U94 , P3_ADD_531_U187 , P3_ADD_531_U186 );
nand NAND2_18983 ( P3_ADD_531_U95 , P3_ADD_531_U189 , P3_ADD_531_U188 );
not NOT1_18984 ( P3_ADD_531_U96 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_18985 ( P3_ADD_531_U97 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_531_U126 );
not NOT1_18986 ( P3_ADD_531_U98 , P3_ADD_531_U7 );
not NOT1_18987 ( P3_ADD_531_U99 , P3_ADD_531_U9 );
not NOT1_18988 ( P3_ADD_531_U100 , P3_ADD_531_U11 );
not NOT1_18989 ( P3_ADD_531_U101 , P3_ADD_531_U13 );
not NOT1_18990 ( P3_ADD_531_U102 , P3_ADD_531_U15 );
not NOT1_18991 ( P3_ADD_531_U103 , P3_ADD_531_U17 );
not NOT1_18992 ( P3_ADD_531_U104 , P3_ADD_531_U19 );
not NOT1_18993 ( P3_ADD_531_U105 , P3_ADD_531_U22 );
not NOT1_18994 ( P3_ADD_531_U106 , P3_ADD_531_U23 );
not NOT1_18995 ( P3_ADD_531_U107 , P3_ADD_531_U25 );
not NOT1_18996 ( P3_ADD_531_U108 , P3_ADD_531_U27 );
not NOT1_18997 ( P3_ADD_531_U109 , P3_ADD_531_U29 );
not NOT1_18998 ( P3_ADD_531_U110 , P3_ADD_531_U31 );
not NOT1_18999 ( P3_ADD_531_U111 , P3_ADD_531_U33 );
not NOT1_19000 ( P3_ADD_531_U112 , P3_ADD_531_U35 );
not NOT1_19001 ( P3_ADD_531_U113 , P3_ADD_531_U37 );
not NOT1_19002 ( P3_ADD_531_U114 , P3_ADD_531_U39 );
not NOT1_19003 ( P3_ADD_531_U115 , P3_ADD_531_U41 );
not NOT1_19004 ( P3_ADD_531_U116 , P3_ADD_531_U43 );
not NOT1_19005 ( P3_ADD_531_U117 , P3_ADD_531_U45 );
not NOT1_19006 ( P3_ADD_531_U118 , P3_ADD_531_U47 );
not NOT1_19007 ( P3_ADD_531_U119 , P3_ADD_531_U49 );
not NOT1_19008 ( P3_ADD_531_U120 , P3_ADD_531_U51 );
not NOT1_19009 ( P3_ADD_531_U121 , P3_ADD_531_U53 );
not NOT1_19010 ( P3_ADD_531_U122 , P3_ADD_531_U55 );
not NOT1_19011 ( P3_ADD_531_U123 , P3_ADD_531_U57 );
not NOT1_19012 ( P3_ADD_531_U124 , P3_ADD_531_U59 );
not NOT1_19013 ( P3_ADD_531_U125 , P3_ADD_531_U61 );
not NOT1_19014 ( P3_ADD_531_U126 , P3_ADD_531_U63 );
not NOT1_19015 ( P3_ADD_531_U127 , P3_ADD_531_U97 );
nand NAND2_19016 ( P3_ADD_531_U128 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_531_U22 );
nand NAND2_19017 ( P3_ADD_531_U129 , P3_ADD_531_U105 , P3_ADD_531_U21 );
nand NAND2_19018 ( P3_ADD_531_U130 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_531_U19 );
nand NAND2_19019 ( P3_ADD_531_U131 , P3_ADD_531_U104 , P3_ADD_531_U20 );
nand NAND2_19020 ( P3_ADD_531_U132 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_531_U17 );
nand NAND2_19021 ( P3_ADD_531_U133 , P3_ADD_531_U103 , P3_ADD_531_U18 );
nand NAND2_19022 ( P3_ADD_531_U134 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_531_U15 );
nand NAND2_19023 ( P3_ADD_531_U135 , P3_ADD_531_U102 , P3_ADD_531_U16 );
nand NAND2_19024 ( P3_ADD_531_U136 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_531_U13 );
nand NAND2_19025 ( P3_ADD_531_U137 , P3_ADD_531_U101 , P3_ADD_531_U14 );
nand NAND2_19026 ( P3_ADD_531_U138 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_531_U11 );
nand NAND2_19027 ( P3_ADD_531_U139 , P3_ADD_531_U100 , P3_ADD_531_U12 );
nand NAND2_19028 ( P3_ADD_531_U140 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_531_U9 );
nand NAND2_19029 ( P3_ADD_531_U141 , P3_ADD_531_U99 , P3_ADD_531_U10 );
nand NAND2_19030 ( P3_ADD_531_U142 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_531_U97 );
nand NAND2_19031 ( P3_ADD_531_U143 , P3_ADD_531_U127 , P3_ADD_531_U96 );
nand NAND2_19032 ( P3_ADD_531_U144 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_531_U63 );
nand NAND2_19033 ( P3_ADD_531_U145 , P3_ADD_531_U126 , P3_ADD_531_U64 );
nand NAND2_19034 ( P3_ADD_531_U146 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_531_U7 );
nand NAND2_19035 ( P3_ADD_531_U147 , P3_ADD_531_U98 , P3_ADD_531_U8 );
nand NAND2_19036 ( P3_ADD_531_U148 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_531_U61 );
nand NAND2_19037 ( P3_ADD_531_U149 , P3_ADD_531_U125 , P3_ADD_531_U62 );
nand NAND2_19038 ( P3_ADD_531_U150 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_531_U59 );
nand NAND2_19039 ( P3_ADD_531_U151 , P3_ADD_531_U124 , P3_ADD_531_U60 );
nand NAND2_19040 ( P3_ADD_531_U152 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_531_U57 );
nand NAND2_19041 ( P3_ADD_531_U153 , P3_ADD_531_U123 , P3_ADD_531_U58 );
nand NAND2_19042 ( P3_ADD_531_U154 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_531_U55 );
nand NAND2_19043 ( P3_ADD_531_U155 , P3_ADD_531_U122 , P3_ADD_531_U56 );
nand NAND2_19044 ( P3_ADD_531_U156 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_531_U53 );
nand NAND2_19045 ( P3_ADD_531_U157 , P3_ADD_531_U121 , P3_ADD_531_U54 );
nand NAND2_19046 ( P3_ADD_531_U158 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_531_U51 );
nand NAND2_19047 ( P3_ADD_531_U159 , P3_ADD_531_U120 , P3_ADD_531_U52 );
nand NAND2_19048 ( P3_ADD_531_U160 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_531_U49 );
nand NAND2_19049 ( P3_ADD_531_U161 , P3_ADD_531_U119 , P3_ADD_531_U50 );
nand NAND2_19050 ( P3_ADD_531_U162 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_531_U47 );
nand NAND2_19051 ( P3_ADD_531_U163 , P3_ADD_531_U118 , P3_ADD_531_U48 );
nand NAND2_19052 ( P3_ADD_531_U164 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_531_U45 );
nand NAND2_19053 ( P3_ADD_531_U165 , P3_ADD_531_U117 , P3_ADD_531_U46 );
nand NAND2_19054 ( P3_ADD_531_U166 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_531_U43 );
nand NAND2_19055 ( P3_ADD_531_U167 , P3_ADD_531_U116 , P3_ADD_531_U44 );
nand NAND2_19056 ( P3_ADD_531_U168 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_531_U5 );
nand NAND2_19057 ( P3_ADD_531_U169 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_531_U6 );
nand NAND2_19058 ( P3_ADD_531_U170 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_531_U41 );
nand NAND2_19059 ( P3_ADD_531_U171 , P3_ADD_531_U115 , P3_ADD_531_U42 );
nand NAND2_19060 ( P3_ADD_531_U172 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_531_U39 );
nand NAND2_19061 ( P3_ADD_531_U173 , P3_ADD_531_U114 , P3_ADD_531_U40 );
nand NAND2_19062 ( P3_ADD_531_U174 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_531_U37 );
nand NAND2_19063 ( P3_ADD_531_U175 , P3_ADD_531_U113 , P3_ADD_531_U38 );
nand NAND2_19064 ( P3_ADD_531_U176 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_531_U35 );
nand NAND2_19065 ( P3_ADD_531_U177 , P3_ADD_531_U112 , P3_ADD_531_U36 );
nand NAND2_19066 ( P3_ADD_531_U178 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_531_U33 );
nand NAND2_19067 ( P3_ADD_531_U179 , P3_ADD_531_U111 , P3_ADD_531_U34 );
nand NAND2_19068 ( P3_ADD_531_U180 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_531_U31 );
nand NAND2_19069 ( P3_ADD_531_U181 , P3_ADD_531_U110 , P3_ADD_531_U32 );
nand NAND2_19070 ( P3_ADD_531_U182 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_531_U29 );
nand NAND2_19071 ( P3_ADD_531_U183 , P3_ADD_531_U109 , P3_ADD_531_U30 );
nand NAND2_19072 ( P3_ADD_531_U184 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_531_U27 );
nand NAND2_19073 ( P3_ADD_531_U185 , P3_ADD_531_U108 , P3_ADD_531_U28 );
nand NAND2_19074 ( P3_ADD_531_U186 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_531_U25 );
nand NAND2_19075 ( P3_ADD_531_U187 , P3_ADD_531_U107 , P3_ADD_531_U26 );
nand NAND2_19076 ( P3_ADD_531_U188 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_531_U23 );
nand NAND2_19077 ( P3_ADD_531_U189 , P3_ADD_531_U106 , P3_ADD_531_U24 );
and AND2_19078 ( P3_SUB_320_U6 , P3_SUB_320_U126 , P3_SUB_320_U28 );
and AND2_19079 ( P3_SUB_320_U7 , P3_SUB_320_U124 , P3_SUB_320_U29 );
and AND2_19080 ( P3_SUB_320_U8 , P3_SUB_320_U122 , P3_SUB_320_U30 );
and AND2_19081 ( P3_SUB_320_U9 , P3_SUB_320_U120 , P3_SUB_320_U31 );
and AND2_19082 ( P3_SUB_320_U10 , P3_SUB_320_U118 , P3_SUB_320_U32 );
and AND2_19083 ( P3_SUB_320_U11 , P3_SUB_320_U116 , P3_SUB_320_U33 );
and AND2_19084 ( P3_SUB_320_U12 , P3_SUB_320_U114 , P3_SUB_320_U34 );
and AND2_19085 ( P3_SUB_320_U13 , P3_SUB_320_U112 , P3_SUB_320_U35 );
and AND2_19086 ( P3_SUB_320_U14 , P3_SUB_320_U110 , P3_SUB_320_U36 );
and AND2_19087 ( P3_SUB_320_U15 , P3_SUB_320_U108 , P3_SUB_320_U37 );
and AND2_19088 ( P3_SUB_320_U16 , P3_SUB_320_U106 , P3_SUB_320_U38 );
and AND2_19089 ( P3_SUB_320_U17 , P3_SUB_320_U105 , P3_SUB_320_U21 );
and AND2_19090 ( P3_SUB_320_U18 , P3_SUB_320_U92 , P3_SUB_320_U22 );
and AND2_19091 ( P3_SUB_320_U19 , P3_SUB_320_U90 , P3_SUB_320_U23 );
and AND2_19092 ( P3_SUB_320_U20 , P3_SUB_320_U88 , P3_SUB_320_U24 );
or OR3_19093 ( P3_SUB_320_U21 , P3_ADD_318_U4 , P3_PHYADDRPOINTER_REG_0_ , P3_ADD_318_U71 );
nand NAND3_19094 ( P3_SUB_320_U22 , P3_SUB_320_U27 , P3_SUB_320_U58 , P3_SUB_320_U83 );
nand NAND3_19095 ( P3_SUB_320_U23 , P3_SUB_320_U26 , P3_SUB_320_U56 , P3_SUB_320_U84 );
nand NAND3_19096 ( P3_SUB_320_U24 , P3_SUB_320_U25 , P3_SUB_320_U54 , P3_SUB_320_U85 );
not NOT1_19097 ( P3_SUB_320_U25 , P3_ADD_318_U63 );
not NOT1_19098 ( P3_SUB_320_U26 , P3_ADD_318_U65 );
not NOT1_19099 ( P3_SUB_320_U27 , P3_ADD_318_U67 );
nand NAND3_19100 ( P3_SUB_320_U28 , P3_SUB_320_U52 , P3_SUB_320_U49 , P3_SUB_320_U86 );
nand NAND3_19101 ( P3_SUB_320_U29 , P3_SUB_320_U48 , P3_SUB_320_U81 , P3_SUB_320_U93 );
nand NAND3_19102 ( P3_SUB_320_U30 , P3_SUB_320_U47 , P3_SUB_320_U79 , P3_SUB_320_U94 );
nand NAND3_19103 ( P3_SUB_320_U31 , P3_SUB_320_U46 , P3_SUB_320_U77 , P3_SUB_320_U95 );
nand NAND3_19104 ( P3_SUB_320_U32 , P3_SUB_320_U45 , P3_SUB_320_U75 , P3_SUB_320_U96 );
nand NAND3_19105 ( P3_SUB_320_U33 , P3_SUB_320_U44 , P3_SUB_320_U73 , P3_SUB_320_U97 );
nand NAND3_19106 ( P3_SUB_320_U34 , P3_SUB_320_U43 , P3_SUB_320_U69 , P3_SUB_320_U98 );
nand NAND3_19107 ( P3_SUB_320_U35 , P3_SUB_320_U42 , P3_SUB_320_U67 , P3_SUB_320_U99 );
nand NAND3_19108 ( P3_SUB_320_U36 , P3_SUB_320_U41 , P3_SUB_320_U65 , P3_SUB_320_U100 );
nand NAND3_19109 ( P3_SUB_320_U37 , P3_SUB_320_U40 , P3_SUB_320_U63 , P3_SUB_320_U101 );
nand NAND2_19110 ( P3_SUB_320_U38 , P3_SUB_320_U102 , P3_SUB_320_U39 );
not NOT1_19111 ( P3_SUB_320_U39 , P3_ADD_318_U72 );
not NOT1_19112 ( P3_SUB_320_U40 , P3_ADD_318_U73 );
not NOT1_19113 ( P3_SUB_320_U41 , P3_ADD_318_U75 );
not NOT1_19114 ( P3_SUB_320_U42 , P3_ADD_318_U77 );
not NOT1_19115 ( P3_SUB_320_U43 , P3_ADD_318_U79 );
not NOT1_19116 ( P3_SUB_320_U44 , P3_ADD_318_U81 );
not NOT1_19117 ( P3_SUB_320_U45 , P3_ADD_318_U83 );
not NOT1_19118 ( P3_SUB_320_U46 , P3_ADD_318_U85 );
not NOT1_19119 ( P3_SUB_320_U47 , P3_ADD_318_U87 );
not NOT1_19120 ( P3_SUB_320_U48 , P3_ADD_318_U89 );
not NOT1_19121 ( P3_SUB_320_U49 , P3_ADD_318_U91 );
nand NAND2_19122 ( P3_SUB_320_U50 , P3_SUB_320_U149 , P3_SUB_320_U148 );
nand NAND2_19123 ( P3_SUB_320_U51 , P3_SUB_320_U137 , P3_SUB_320_U136 );
not NOT1_19124 ( P3_SUB_320_U52 , P3_ADD_318_U62 );
and AND2_19125 ( P3_SUB_320_U53 , P3_SUB_320_U129 , P3_SUB_320_U128 );
not NOT1_19126 ( P3_SUB_320_U54 , P3_ADD_318_U64 );
and AND2_19127 ( P3_SUB_320_U55 , P3_SUB_320_U131 , P3_SUB_320_U130 );
not NOT1_19128 ( P3_SUB_320_U56 , P3_ADD_318_U66 );
and AND2_19129 ( P3_SUB_320_U57 , P3_SUB_320_U133 , P3_SUB_320_U132 );
not NOT1_19130 ( P3_SUB_320_U58 , P3_ADD_318_U68 );
and AND2_19131 ( P3_SUB_320_U59 , P3_SUB_320_U135 , P3_SUB_320_U134 );
not NOT1_19132 ( P3_SUB_320_U60 , P3_ADD_318_U69 );
not NOT1_19133 ( P3_SUB_320_U61 , P3_ADD_318_U70 );
and AND2_19134 ( P3_SUB_320_U62 , P3_SUB_320_U139 , P3_SUB_320_U138 );
not NOT1_19135 ( P3_SUB_320_U63 , P3_ADD_318_U74 );
and AND2_19136 ( P3_SUB_320_U64 , P3_SUB_320_U141 , P3_SUB_320_U140 );
not NOT1_19137 ( P3_SUB_320_U65 , P3_ADD_318_U76 );
and AND2_19138 ( P3_SUB_320_U66 , P3_SUB_320_U143 , P3_SUB_320_U142 );
not NOT1_19139 ( P3_SUB_320_U67 , P3_ADD_318_U78 );
and AND2_19140 ( P3_SUB_320_U68 , P3_SUB_320_U145 , P3_SUB_320_U144 );
not NOT1_19141 ( P3_SUB_320_U69 , P3_ADD_318_U80 );
and AND2_19142 ( P3_SUB_320_U70 , P3_SUB_320_U147 , P3_SUB_320_U146 );
not NOT1_19143 ( P3_SUB_320_U71 , P3_ADD_318_U4 );
not NOT1_19144 ( P3_SUB_320_U72 , P3_PHYADDRPOINTER_REG_0_ );
not NOT1_19145 ( P3_SUB_320_U73 , P3_ADD_318_U82 );
and AND2_19146 ( P3_SUB_320_U74 , P3_SUB_320_U151 , P3_SUB_320_U150 );
not NOT1_19147 ( P3_SUB_320_U75 , P3_ADD_318_U84 );
and AND2_19148 ( P3_SUB_320_U76 , P3_SUB_320_U153 , P3_SUB_320_U152 );
not NOT1_19149 ( P3_SUB_320_U77 , P3_ADD_318_U86 );
and AND2_19150 ( P3_SUB_320_U78 , P3_SUB_320_U155 , P3_SUB_320_U154 );
not NOT1_19151 ( P3_SUB_320_U79 , P3_ADD_318_U88 );
and AND2_19152 ( P3_SUB_320_U80 , P3_SUB_320_U157 , P3_SUB_320_U156 );
not NOT1_19153 ( P3_SUB_320_U81 , P3_ADD_318_U90 );
and AND2_19154 ( P3_SUB_320_U82 , P3_SUB_320_U159 , P3_SUB_320_U158 );
not NOT1_19155 ( P3_SUB_320_U83 , P3_SUB_320_U21 );
not NOT1_19156 ( P3_SUB_320_U84 , P3_SUB_320_U22 );
not NOT1_19157 ( P3_SUB_320_U85 , P3_SUB_320_U23 );
not NOT1_19158 ( P3_SUB_320_U86 , P3_SUB_320_U24 );
nand NAND2_19159 ( P3_SUB_320_U87 , P3_SUB_320_U85 , P3_SUB_320_U54 );
nand NAND2_19160 ( P3_SUB_320_U88 , P3_ADD_318_U63 , P3_SUB_320_U87 );
nand NAND2_19161 ( P3_SUB_320_U89 , P3_SUB_320_U84 , P3_SUB_320_U56 );
nand NAND2_19162 ( P3_SUB_320_U90 , P3_ADD_318_U65 , P3_SUB_320_U89 );
nand NAND2_19163 ( P3_SUB_320_U91 , P3_SUB_320_U83 , P3_SUB_320_U58 );
nand NAND2_19164 ( P3_SUB_320_U92 , P3_ADD_318_U67 , P3_SUB_320_U91 );
not NOT1_19165 ( P3_SUB_320_U93 , P3_SUB_320_U28 );
not NOT1_19166 ( P3_SUB_320_U94 , P3_SUB_320_U29 );
not NOT1_19167 ( P3_SUB_320_U95 , P3_SUB_320_U30 );
not NOT1_19168 ( P3_SUB_320_U96 , P3_SUB_320_U31 );
not NOT1_19169 ( P3_SUB_320_U97 , P3_SUB_320_U32 );
not NOT1_19170 ( P3_SUB_320_U98 , P3_SUB_320_U33 );
not NOT1_19171 ( P3_SUB_320_U99 , P3_SUB_320_U34 );
not NOT1_19172 ( P3_SUB_320_U100 , P3_SUB_320_U35 );
not NOT1_19173 ( P3_SUB_320_U101 , P3_SUB_320_U36 );
not NOT1_19174 ( P3_SUB_320_U102 , P3_SUB_320_U37 );
not NOT1_19175 ( P3_SUB_320_U103 , P3_SUB_320_U38 );
or OR2_19176 ( P3_SUB_320_U104 , P3_ADD_318_U4 , P3_PHYADDRPOINTER_REG_0_ );
nand NAND2_19177 ( P3_SUB_320_U105 , P3_ADD_318_U71 , P3_SUB_320_U104 );
nand NAND2_19178 ( P3_SUB_320_U106 , P3_ADD_318_U72 , P3_SUB_320_U37 );
nand NAND2_19179 ( P3_SUB_320_U107 , P3_SUB_320_U101 , P3_SUB_320_U63 );
nand NAND2_19180 ( P3_SUB_320_U108 , P3_ADD_318_U73 , P3_SUB_320_U107 );
nand NAND2_19181 ( P3_SUB_320_U109 , P3_SUB_320_U100 , P3_SUB_320_U65 );
nand NAND2_19182 ( P3_SUB_320_U110 , P3_ADD_318_U75 , P3_SUB_320_U109 );
nand NAND2_19183 ( P3_SUB_320_U111 , P3_SUB_320_U99 , P3_SUB_320_U67 );
nand NAND2_19184 ( P3_SUB_320_U112 , P3_ADD_318_U77 , P3_SUB_320_U111 );
nand NAND2_19185 ( P3_SUB_320_U113 , P3_SUB_320_U98 , P3_SUB_320_U69 );
nand NAND2_19186 ( P3_SUB_320_U114 , P3_ADD_318_U79 , P3_SUB_320_U113 );
nand NAND2_19187 ( P3_SUB_320_U115 , P3_SUB_320_U97 , P3_SUB_320_U73 );
nand NAND2_19188 ( P3_SUB_320_U116 , P3_ADD_318_U81 , P3_SUB_320_U115 );
nand NAND2_19189 ( P3_SUB_320_U117 , P3_SUB_320_U96 , P3_SUB_320_U75 );
nand NAND2_19190 ( P3_SUB_320_U118 , P3_ADD_318_U83 , P3_SUB_320_U117 );
nand NAND2_19191 ( P3_SUB_320_U119 , P3_SUB_320_U95 , P3_SUB_320_U77 );
nand NAND2_19192 ( P3_SUB_320_U120 , P3_ADD_318_U85 , P3_SUB_320_U119 );
nand NAND2_19193 ( P3_SUB_320_U121 , P3_SUB_320_U94 , P3_SUB_320_U79 );
nand NAND2_19194 ( P3_SUB_320_U122 , P3_ADD_318_U87 , P3_SUB_320_U121 );
nand NAND2_19195 ( P3_SUB_320_U123 , P3_SUB_320_U93 , P3_SUB_320_U81 );
nand NAND2_19196 ( P3_SUB_320_U124 , P3_ADD_318_U89 , P3_SUB_320_U123 );
nand NAND2_19197 ( P3_SUB_320_U125 , P3_SUB_320_U86 , P3_SUB_320_U52 );
nand NAND2_19198 ( P3_SUB_320_U126 , P3_ADD_318_U91 , P3_SUB_320_U125 );
nand NAND2_19199 ( P3_SUB_320_U127 , P3_SUB_320_U103 , P3_SUB_320_U61 );
nand NAND2_19200 ( P3_SUB_320_U128 , P3_ADD_318_U62 , P3_SUB_320_U24 );
nand NAND2_19201 ( P3_SUB_320_U129 , P3_SUB_320_U86 , P3_SUB_320_U52 );
nand NAND2_19202 ( P3_SUB_320_U130 , P3_ADD_318_U64 , P3_SUB_320_U23 );
nand NAND2_19203 ( P3_SUB_320_U131 , P3_SUB_320_U85 , P3_SUB_320_U54 );
nand NAND2_19204 ( P3_SUB_320_U132 , P3_ADD_318_U66 , P3_SUB_320_U22 );
nand NAND2_19205 ( P3_SUB_320_U133 , P3_SUB_320_U84 , P3_SUB_320_U56 );
nand NAND2_19206 ( P3_SUB_320_U134 , P3_ADD_318_U68 , P3_SUB_320_U21 );
nand NAND2_19207 ( P3_SUB_320_U135 , P3_SUB_320_U83 , P3_SUB_320_U58 );
nand NAND2_19208 ( P3_SUB_320_U136 , P3_SUB_320_U127 , P3_SUB_320_U60 );
nand NAND3_19209 ( P3_SUB_320_U137 , P3_SUB_320_U103 , P3_SUB_320_U61 , P3_ADD_318_U69 );
nand NAND2_19210 ( P3_SUB_320_U138 , P3_ADD_318_U70 , P3_SUB_320_U38 );
nand NAND2_19211 ( P3_SUB_320_U139 , P3_SUB_320_U103 , P3_SUB_320_U61 );
nand NAND2_19212 ( P3_SUB_320_U140 , P3_ADD_318_U74 , P3_SUB_320_U36 );
nand NAND2_19213 ( P3_SUB_320_U141 , P3_SUB_320_U101 , P3_SUB_320_U63 );
nand NAND2_19214 ( P3_SUB_320_U142 , P3_ADD_318_U76 , P3_SUB_320_U35 );
nand NAND2_19215 ( P3_SUB_320_U143 , P3_SUB_320_U100 , P3_SUB_320_U65 );
nand NAND2_19216 ( P3_SUB_320_U144 , P3_ADD_318_U78 , P3_SUB_320_U34 );
nand NAND2_19217 ( P3_SUB_320_U145 , P3_SUB_320_U99 , P3_SUB_320_U67 );
nand NAND2_19218 ( P3_SUB_320_U146 , P3_ADD_318_U80 , P3_SUB_320_U33 );
nand NAND2_19219 ( P3_SUB_320_U147 , P3_SUB_320_U98 , P3_SUB_320_U69 );
nand NAND2_19220 ( P3_SUB_320_U148 , P3_ADD_318_U4 , P3_SUB_320_U72 );
nand NAND2_19221 ( P3_SUB_320_U149 , P3_PHYADDRPOINTER_REG_0_ , P3_SUB_320_U71 );
nand NAND2_19222 ( P3_SUB_320_U150 , P3_ADD_318_U82 , P3_SUB_320_U32 );
nand NAND2_19223 ( P3_SUB_320_U151 , P3_SUB_320_U97 , P3_SUB_320_U73 );
nand NAND2_19224 ( P3_SUB_320_U152 , P3_ADD_318_U84 , P3_SUB_320_U31 );
nand NAND2_19225 ( P3_SUB_320_U153 , P3_SUB_320_U96 , P3_SUB_320_U75 );
nand NAND2_19226 ( P3_SUB_320_U154 , P3_ADD_318_U86 , P3_SUB_320_U30 );
nand NAND2_19227 ( P3_SUB_320_U155 , P3_SUB_320_U95 , P3_SUB_320_U77 );
nand NAND2_19228 ( P3_SUB_320_U156 , P3_ADD_318_U88 , P3_SUB_320_U29 );
nand NAND2_19229 ( P3_SUB_320_U157 , P3_SUB_320_U94 , P3_SUB_320_U79 );
nand NAND2_19230 ( P3_SUB_320_U158 , P3_ADD_318_U90 , P3_SUB_320_U28 );
nand NAND2_19231 ( P3_SUB_320_U159 , P3_SUB_320_U93 , P3_SUB_320_U81 );
not NOT1_19232 ( P3_ADD_505_U5 , P3_INSTQUEUERD_ADDR_REG_0_ );
and AND2_19233 ( P3_ADD_505_U6 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_ADD_505_U20 );
not NOT1_19234 ( P3_ADD_505_U7 , P3_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_19235 ( P3_ADD_505_U8 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_INSTQUEUERD_ADDR_REG_0_ );
not NOT1_19236 ( P3_ADD_505_U9 , P3_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_19237 ( P3_ADD_505_U10 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_ADD_505_U18 );
not NOT1_19238 ( P3_ADD_505_U11 , P3_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_19239 ( P3_ADD_505_U12 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_ADD_505_U19 );
not NOT1_19240 ( P3_ADD_505_U13 , P3_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_19241 ( P3_ADD_505_U14 , P3_ADD_505_U22 , P3_ADD_505_U21 );
nand NAND2_19242 ( P3_ADD_505_U15 , P3_ADD_505_U24 , P3_ADD_505_U23 );
nand NAND2_19243 ( P3_ADD_505_U16 , P3_ADD_505_U26 , P3_ADD_505_U25 );
nand NAND2_19244 ( P3_ADD_505_U17 , P3_ADD_505_U28 , P3_ADD_505_U27 );
not NOT1_19245 ( P3_ADD_505_U18 , P3_ADD_505_U8 );
not NOT1_19246 ( P3_ADD_505_U19 , P3_ADD_505_U10 );
not NOT1_19247 ( P3_ADD_505_U20 , P3_ADD_505_U12 );
nand NAND2_19248 ( P3_ADD_505_U21 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_ADD_505_U12 );
nand NAND2_19249 ( P3_ADD_505_U22 , P3_ADD_505_U20 , P3_ADD_505_U13 );
nand NAND2_19250 ( P3_ADD_505_U23 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_ADD_505_U10 );
nand NAND2_19251 ( P3_ADD_505_U24 , P3_ADD_505_U19 , P3_ADD_505_U11 );
nand NAND2_19252 ( P3_ADD_505_U25 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_ADD_505_U8 );
nand NAND2_19253 ( P3_ADD_505_U26 , P3_ADD_505_U18 , P3_ADD_505_U9 );
nand NAND2_19254 ( P3_ADD_505_U27 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_ADD_505_U5 );
nand NAND2_19255 ( P3_ADD_505_U28 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_ADD_505_U7 );
nor nor_19256 ( P3_GTE_485_U6 , P3_SUB_485_U6 , P3_GTE_485_U7 );
nor nor_19257 ( P3_GTE_485_U7 , P3_SUB_485_U16 , P3_SUB_485_U17 , P3_SUB_485_U19 , P3_SUB_485_U18 );
not NOT1_19258 ( P3_ADD_318_U4 , P3_PHYADDRPOINTER_REG_1_ );
not NOT1_19259 ( P3_ADD_318_U5 , P3_PHYADDRPOINTER_REG_2_ );
nand NAND2_19260 ( P3_ADD_318_U6 , P3_PHYADDRPOINTER_REG_2_ , P3_PHYADDRPOINTER_REG_1_ );
not NOT1_19261 ( P3_ADD_318_U7 , P3_PHYADDRPOINTER_REG_3_ );
nand NAND2_19262 ( P3_ADD_318_U8 , P3_PHYADDRPOINTER_REG_3_ , P3_ADD_318_U94 );
not NOT1_19263 ( P3_ADD_318_U9 , P3_PHYADDRPOINTER_REG_4_ );
nand NAND2_19264 ( P3_ADD_318_U10 , P3_PHYADDRPOINTER_REG_4_ , P3_ADD_318_U95 );
not NOT1_19265 ( P3_ADD_318_U11 , P3_PHYADDRPOINTER_REG_5_ );
nand NAND2_19266 ( P3_ADD_318_U12 , P3_PHYADDRPOINTER_REG_5_ , P3_ADD_318_U96 );
not NOT1_19267 ( P3_ADD_318_U13 , P3_PHYADDRPOINTER_REG_6_ );
nand NAND2_19268 ( P3_ADD_318_U14 , P3_PHYADDRPOINTER_REG_6_ , P3_ADD_318_U97 );
not NOT1_19269 ( P3_ADD_318_U15 , P3_PHYADDRPOINTER_REG_7_ );
nand NAND2_19270 ( P3_ADD_318_U16 , P3_PHYADDRPOINTER_REG_7_ , P3_ADD_318_U98 );
not NOT1_19271 ( P3_ADD_318_U17 , P3_PHYADDRPOINTER_REG_8_ );
not NOT1_19272 ( P3_ADD_318_U18 , P3_PHYADDRPOINTER_REG_9_ );
nand NAND2_19273 ( P3_ADD_318_U19 , P3_PHYADDRPOINTER_REG_8_ , P3_ADD_318_U99 );
nand NAND2_19274 ( P3_ADD_318_U20 , P3_ADD_318_U100 , P3_PHYADDRPOINTER_REG_9_ );
not NOT1_19275 ( P3_ADD_318_U21 , P3_PHYADDRPOINTER_REG_10_ );
nand NAND2_19276 ( P3_ADD_318_U22 , P3_PHYADDRPOINTER_REG_10_ , P3_ADD_318_U101 );
not NOT1_19277 ( P3_ADD_318_U23 , P3_PHYADDRPOINTER_REG_11_ );
nand NAND2_19278 ( P3_ADD_318_U24 , P3_PHYADDRPOINTER_REG_11_ , P3_ADD_318_U102 );
not NOT1_19279 ( P3_ADD_318_U25 , P3_PHYADDRPOINTER_REG_12_ );
nand NAND2_19280 ( P3_ADD_318_U26 , P3_PHYADDRPOINTER_REG_12_ , P3_ADD_318_U103 );
not NOT1_19281 ( P3_ADD_318_U27 , P3_PHYADDRPOINTER_REG_13_ );
nand NAND2_19282 ( P3_ADD_318_U28 , P3_PHYADDRPOINTER_REG_13_ , P3_ADD_318_U104 );
not NOT1_19283 ( P3_ADD_318_U29 , P3_PHYADDRPOINTER_REG_14_ );
nand NAND2_19284 ( P3_ADD_318_U30 , P3_PHYADDRPOINTER_REG_14_ , P3_ADD_318_U105 );
not NOT1_19285 ( P3_ADD_318_U31 , P3_PHYADDRPOINTER_REG_15_ );
nand NAND2_19286 ( P3_ADD_318_U32 , P3_PHYADDRPOINTER_REG_15_ , P3_ADD_318_U106 );
not NOT1_19287 ( P3_ADD_318_U33 , P3_PHYADDRPOINTER_REG_16_ );
nand NAND2_19288 ( P3_ADD_318_U34 , P3_PHYADDRPOINTER_REG_16_ , P3_ADD_318_U107 );
not NOT1_19289 ( P3_ADD_318_U35 , P3_PHYADDRPOINTER_REG_17_ );
nand NAND2_19290 ( P3_ADD_318_U36 , P3_PHYADDRPOINTER_REG_17_ , P3_ADD_318_U108 );
not NOT1_19291 ( P3_ADD_318_U37 , P3_PHYADDRPOINTER_REG_18_ );
nand NAND2_19292 ( P3_ADD_318_U38 , P3_PHYADDRPOINTER_REG_18_ , P3_ADD_318_U109 );
not NOT1_19293 ( P3_ADD_318_U39 , P3_PHYADDRPOINTER_REG_19_ );
nand NAND2_19294 ( P3_ADD_318_U40 , P3_PHYADDRPOINTER_REG_19_ , P3_ADD_318_U110 );
not NOT1_19295 ( P3_ADD_318_U41 , P3_PHYADDRPOINTER_REG_20_ );
nand NAND2_19296 ( P3_ADD_318_U42 , P3_PHYADDRPOINTER_REG_20_ , P3_ADD_318_U111 );
not NOT1_19297 ( P3_ADD_318_U43 , P3_PHYADDRPOINTER_REG_21_ );
nand NAND2_19298 ( P3_ADD_318_U44 , P3_PHYADDRPOINTER_REG_21_ , P3_ADD_318_U112 );
not NOT1_19299 ( P3_ADD_318_U45 , P3_PHYADDRPOINTER_REG_22_ );
nand NAND2_19300 ( P3_ADD_318_U46 , P3_PHYADDRPOINTER_REG_22_ , P3_ADD_318_U113 );
not NOT1_19301 ( P3_ADD_318_U47 , P3_PHYADDRPOINTER_REG_23_ );
nand NAND2_19302 ( P3_ADD_318_U48 , P3_PHYADDRPOINTER_REG_23_ , P3_ADD_318_U114 );
not NOT1_19303 ( P3_ADD_318_U49 , P3_PHYADDRPOINTER_REG_24_ );
nand NAND2_19304 ( P3_ADD_318_U50 , P3_PHYADDRPOINTER_REG_24_ , P3_ADD_318_U115 );
not NOT1_19305 ( P3_ADD_318_U51 , P3_PHYADDRPOINTER_REG_25_ );
nand NAND2_19306 ( P3_ADD_318_U52 , P3_PHYADDRPOINTER_REG_25_ , P3_ADD_318_U116 );
not NOT1_19307 ( P3_ADD_318_U53 , P3_PHYADDRPOINTER_REG_26_ );
nand NAND2_19308 ( P3_ADD_318_U54 , P3_PHYADDRPOINTER_REG_26_ , P3_ADD_318_U117 );
not NOT1_19309 ( P3_ADD_318_U55 , P3_PHYADDRPOINTER_REG_27_ );
nand NAND2_19310 ( P3_ADD_318_U56 , P3_PHYADDRPOINTER_REG_27_ , P3_ADD_318_U118 );
not NOT1_19311 ( P3_ADD_318_U57 , P3_PHYADDRPOINTER_REG_28_ );
nand NAND2_19312 ( P3_ADD_318_U58 , P3_PHYADDRPOINTER_REG_28_ , P3_ADD_318_U119 );
not NOT1_19313 ( P3_ADD_318_U59 , P3_PHYADDRPOINTER_REG_29_ );
nand NAND2_19314 ( P3_ADD_318_U60 , P3_PHYADDRPOINTER_REG_29_ , P3_ADD_318_U120 );
not NOT1_19315 ( P3_ADD_318_U61 , P3_PHYADDRPOINTER_REG_30_ );
nand NAND2_19316 ( P3_ADD_318_U62 , P3_ADD_318_U124 , P3_ADD_318_U123 );
nand NAND2_19317 ( P3_ADD_318_U63 , P3_ADD_318_U126 , P3_ADD_318_U125 );
nand NAND2_19318 ( P3_ADD_318_U64 , P3_ADD_318_U128 , P3_ADD_318_U127 );
nand NAND2_19319 ( P3_ADD_318_U65 , P3_ADD_318_U130 , P3_ADD_318_U129 );
nand NAND2_19320 ( P3_ADD_318_U66 , P3_ADD_318_U132 , P3_ADD_318_U131 );
nand NAND2_19321 ( P3_ADD_318_U67 , P3_ADD_318_U134 , P3_ADD_318_U133 );
nand NAND2_19322 ( P3_ADD_318_U68 , P3_ADD_318_U136 , P3_ADD_318_U135 );
nand NAND2_19323 ( P3_ADD_318_U69 , P3_ADD_318_U138 , P3_ADD_318_U137 );
nand NAND2_19324 ( P3_ADD_318_U70 , P3_ADD_318_U140 , P3_ADD_318_U139 );
nand NAND2_19325 ( P3_ADD_318_U71 , P3_ADD_318_U142 , P3_ADD_318_U141 );
nand NAND2_19326 ( P3_ADD_318_U72 , P3_ADD_318_U144 , P3_ADD_318_U143 );
nand NAND2_19327 ( P3_ADD_318_U73 , P3_ADD_318_U146 , P3_ADD_318_U145 );
nand NAND2_19328 ( P3_ADD_318_U74 , P3_ADD_318_U148 , P3_ADD_318_U147 );
nand NAND2_19329 ( P3_ADD_318_U75 , P3_ADD_318_U150 , P3_ADD_318_U149 );
nand NAND2_19330 ( P3_ADD_318_U76 , P3_ADD_318_U152 , P3_ADD_318_U151 );
nand NAND2_19331 ( P3_ADD_318_U77 , P3_ADD_318_U154 , P3_ADD_318_U153 );
nand NAND2_19332 ( P3_ADD_318_U78 , P3_ADD_318_U156 , P3_ADD_318_U155 );
nand NAND2_19333 ( P3_ADD_318_U79 , P3_ADD_318_U158 , P3_ADD_318_U157 );
nand NAND2_19334 ( P3_ADD_318_U80 , P3_ADD_318_U160 , P3_ADD_318_U159 );
nand NAND2_19335 ( P3_ADD_318_U81 , P3_ADD_318_U162 , P3_ADD_318_U161 );
nand NAND2_19336 ( P3_ADD_318_U82 , P3_ADD_318_U164 , P3_ADD_318_U163 );
nand NAND2_19337 ( P3_ADD_318_U83 , P3_ADD_318_U166 , P3_ADD_318_U165 );
nand NAND2_19338 ( P3_ADD_318_U84 , P3_ADD_318_U168 , P3_ADD_318_U167 );
nand NAND2_19339 ( P3_ADD_318_U85 , P3_ADD_318_U170 , P3_ADD_318_U169 );
nand NAND2_19340 ( P3_ADD_318_U86 , P3_ADD_318_U172 , P3_ADD_318_U171 );
nand NAND2_19341 ( P3_ADD_318_U87 , P3_ADD_318_U174 , P3_ADD_318_U173 );
nand NAND2_19342 ( P3_ADD_318_U88 , P3_ADD_318_U176 , P3_ADD_318_U175 );
nand NAND2_19343 ( P3_ADD_318_U89 , P3_ADD_318_U178 , P3_ADD_318_U177 );
nand NAND2_19344 ( P3_ADD_318_U90 , P3_ADD_318_U180 , P3_ADD_318_U179 );
nand NAND2_19345 ( P3_ADD_318_U91 , P3_ADD_318_U182 , P3_ADD_318_U181 );
not NOT1_19346 ( P3_ADD_318_U92 , P3_PHYADDRPOINTER_REG_31_ );
nand NAND2_19347 ( P3_ADD_318_U93 , P3_PHYADDRPOINTER_REG_30_ , P3_ADD_318_U121 );
not NOT1_19348 ( P3_ADD_318_U94 , P3_ADD_318_U6 );
not NOT1_19349 ( P3_ADD_318_U95 , P3_ADD_318_U8 );
not NOT1_19350 ( P3_ADD_318_U96 , P3_ADD_318_U10 );
not NOT1_19351 ( P3_ADD_318_U97 , P3_ADD_318_U12 );
not NOT1_19352 ( P3_ADD_318_U98 , P3_ADD_318_U14 );
not NOT1_19353 ( P3_ADD_318_U99 , P3_ADD_318_U16 );
not NOT1_19354 ( P3_ADD_318_U100 , P3_ADD_318_U19 );
not NOT1_19355 ( P3_ADD_318_U101 , P3_ADD_318_U20 );
not NOT1_19356 ( P3_ADD_318_U102 , P3_ADD_318_U22 );
not NOT1_19357 ( P3_ADD_318_U103 , P3_ADD_318_U24 );
not NOT1_19358 ( P3_ADD_318_U104 , P3_ADD_318_U26 );
not NOT1_19359 ( P3_ADD_318_U105 , P3_ADD_318_U28 );
not NOT1_19360 ( P3_ADD_318_U106 , P3_ADD_318_U30 );
not NOT1_19361 ( P3_ADD_318_U107 , P3_ADD_318_U32 );
not NOT1_19362 ( P3_ADD_318_U108 , P3_ADD_318_U34 );
not NOT1_19363 ( P3_ADD_318_U109 , P3_ADD_318_U36 );
not NOT1_19364 ( P3_ADD_318_U110 , P3_ADD_318_U38 );
not NOT1_19365 ( P3_ADD_318_U111 , P3_ADD_318_U40 );
not NOT1_19366 ( P3_ADD_318_U112 , P3_ADD_318_U42 );
not NOT1_19367 ( P3_ADD_318_U113 , P3_ADD_318_U44 );
not NOT1_19368 ( P3_ADD_318_U114 , P3_ADD_318_U46 );
not NOT1_19369 ( P3_ADD_318_U115 , P3_ADD_318_U48 );
not NOT1_19370 ( P3_ADD_318_U116 , P3_ADD_318_U50 );
not NOT1_19371 ( P3_ADD_318_U117 , P3_ADD_318_U52 );
not NOT1_19372 ( P3_ADD_318_U118 , P3_ADD_318_U54 );
not NOT1_19373 ( P3_ADD_318_U119 , P3_ADD_318_U56 );
not NOT1_19374 ( P3_ADD_318_U120 , P3_ADD_318_U58 );
not NOT1_19375 ( P3_ADD_318_U121 , P3_ADD_318_U60 );
not NOT1_19376 ( P3_ADD_318_U122 , P3_ADD_318_U93 );
nand NAND2_19377 ( P3_ADD_318_U123 , P3_PHYADDRPOINTER_REG_9_ , P3_ADD_318_U19 );
nand NAND2_19378 ( P3_ADD_318_U124 , P3_ADD_318_U100 , P3_ADD_318_U18 );
nand NAND2_19379 ( P3_ADD_318_U125 , P3_PHYADDRPOINTER_REG_8_ , P3_ADD_318_U16 );
nand NAND2_19380 ( P3_ADD_318_U126 , P3_ADD_318_U99 , P3_ADD_318_U17 );
nand NAND2_19381 ( P3_ADD_318_U127 , P3_PHYADDRPOINTER_REG_7_ , P3_ADD_318_U14 );
nand NAND2_19382 ( P3_ADD_318_U128 , P3_ADD_318_U98 , P3_ADD_318_U15 );
nand NAND2_19383 ( P3_ADD_318_U129 , P3_PHYADDRPOINTER_REG_6_ , P3_ADD_318_U12 );
nand NAND2_19384 ( P3_ADD_318_U130 , P3_ADD_318_U97 , P3_ADD_318_U13 );
nand NAND2_19385 ( P3_ADD_318_U131 , P3_PHYADDRPOINTER_REG_5_ , P3_ADD_318_U10 );
nand NAND2_19386 ( P3_ADD_318_U132 , P3_ADD_318_U96 , P3_ADD_318_U11 );
nand NAND2_19387 ( P3_ADD_318_U133 , P3_PHYADDRPOINTER_REG_4_ , P3_ADD_318_U8 );
nand NAND2_19388 ( P3_ADD_318_U134 , P3_ADD_318_U95 , P3_ADD_318_U9 );
nand NAND2_19389 ( P3_ADD_318_U135 , P3_PHYADDRPOINTER_REG_3_ , P3_ADD_318_U6 );
nand NAND2_19390 ( P3_ADD_318_U136 , P3_ADD_318_U94 , P3_ADD_318_U7 );
nand NAND2_19391 ( P3_ADD_318_U137 , P3_PHYADDRPOINTER_REG_31_ , P3_ADD_318_U93 );
nand NAND2_19392 ( P3_ADD_318_U138 , P3_ADD_318_U122 , P3_ADD_318_U92 );
nand NAND2_19393 ( P3_ADD_318_U139 , P3_PHYADDRPOINTER_REG_30_ , P3_ADD_318_U60 );
nand NAND2_19394 ( P3_ADD_318_U140 , P3_ADD_318_U121 , P3_ADD_318_U61 );
nand NAND2_19395 ( P3_ADD_318_U141 , P3_PHYADDRPOINTER_REG_2_ , P3_ADD_318_U4 );
nand NAND2_19396 ( P3_ADD_318_U142 , P3_PHYADDRPOINTER_REG_1_ , P3_ADD_318_U5 );
nand NAND2_19397 ( P3_ADD_318_U143 , P3_PHYADDRPOINTER_REG_29_ , P3_ADD_318_U58 );
nand NAND2_19398 ( P3_ADD_318_U144 , P3_ADD_318_U120 , P3_ADD_318_U59 );
nand NAND2_19399 ( P3_ADD_318_U145 , P3_PHYADDRPOINTER_REG_28_ , P3_ADD_318_U56 );
nand NAND2_19400 ( P3_ADD_318_U146 , P3_ADD_318_U119 , P3_ADD_318_U57 );
nand NAND2_19401 ( P3_ADD_318_U147 , P3_PHYADDRPOINTER_REG_27_ , P3_ADD_318_U54 );
nand NAND2_19402 ( P3_ADD_318_U148 , P3_ADD_318_U118 , P3_ADD_318_U55 );
nand NAND2_19403 ( P3_ADD_318_U149 , P3_PHYADDRPOINTER_REG_26_ , P3_ADD_318_U52 );
nand NAND2_19404 ( P3_ADD_318_U150 , P3_ADD_318_U117 , P3_ADD_318_U53 );
nand NAND2_19405 ( P3_ADD_318_U151 , P3_PHYADDRPOINTER_REG_25_ , P3_ADD_318_U50 );
nand NAND2_19406 ( P3_ADD_318_U152 , P3_ADD_318_U116 , P3_ADD_318_U51 );
nand NAND2_19407 ( P3_ADD_318_U153 , P3_PHYADDRPOINTER_REG_24_ , P3_ADD_318_U48 );
nand NAND2_19408 ( P3_ADD_318_U154 , P3_ADD_318_U115 , P3_ADD_318_U49 );
nand NAND2_19409 ( P3_ADD_318_U155 , P3_PHYADDRPOINTER_REG_23_ , P3_ADD_318_U46 );
nand NAND2_19410 ( P3_ADD_318_U156 , P3_ADD_318_U114 , P3_ADD_318_U47 );
nand NAND2_19411 ( P3_ADD_318_U157 , P3_PHYADDRPOINTER_REG_22_ , P3_ADD_318_U44 );
nand NAND2_19412 ( P3_ADD_318_U158 , P3_ADD_318_U113 , P3_ADD_318_U45 );
nand NAND2_19413 ( P3_ADD_318_U159 , P3_PHYADDRPOINTER_REG_21_ , P3_ADD_318_U42 );
nand NAND2_19414 ( P3_ADD_318_U160 , P3_ADD_318_U112 , P3_ADD_318_U43 );
nand NAND2_19415 ( P3_ADD_318_U161 , P3_PHYADDRPOINTER_REG_20_ , P3_ADD_318_U40 );
nand NAND2_19416 ( P3_ADD_318_U162 , P3_ADD_318_U111 , P3_ADD_318_U41 );
nand NAND2_19417 ( P3_ADD_318_U163 , P3_PHYADDRPOINTER_REG_19_ , P3_ADD_318_U38 );
nand NAND2_19418 ( P3_ADD_318_U164 , P3_ADD_318_U110 , P3_ADD_318_U39 );
nand NAND2_19419 ( P3_ADD_318_U165 , P3_PHYADDRPOINTER_REG_18_ , P3_ADD_318_U36 );
nand NAND2_19420 ( P3_ADD_318_U166 , P3_ADD_318_U109 , P3_ADD_318_U37 );
nand NAND2_19421 ( P3_ADD_318_U167 , P3_PHYADDRPOINTER_REG_17_ , P3_ADD_318_U34 );
nand NAND2_19422 ( P3_ADD_318_U168 , P3_ADD_318_U108 , P3_ADD_318_U35 );
nand NAND2_19423 ( P3_ADD_318_U169 , P3_PHYADDRPOINTER_REG_16_ , P3_ADD_318_U32 );
nand NAND2_19424 ( P3_ADD_318_U170 , P3_ADD_318_U107 , P3_ADD_318_U33 );
nand NAND2_19425 ( P3_ADD_318_U171 , P3_PHYADDRPOINTER_REG_15_ , P3_ADD_318_U30 );
nand NAND2_19426 ( P3_ADD_318_U172 , P3_ADD_318_U106 , P3_ADD_318_U31 );
nand NAND2_19427 ( P3_ADD_318_U173 , P3_PHYADDRPOINTER_REG_14_ , P3_ADD_318_U28 );
nand NAND2_19428 ( P3_ADD_318_U174 , P3_ADD_318_U105 , P3_ADD_318_U29 );
nand NAND2_19429 ( P3_ADD_318_U175 , P3_PHYADDRPOINTER_REG_13_ , P3_ADD_318_U26 );
nand NAND2_19430 ( P3_ADD_318_U176 , P3_ADD_318_U104 , P3_ADD_318_U27 );
nand NAND2_19431 ( P3_ADD_318_U177 , P3_PHYADDRPOINTER_REG_12_ , P3_ADD_318_U24 );
nand NAND2_19432 ( P3_ADD_318_U178 , P3_ADD_318_U103 , P3_ADD_318_U25 );
nand NAND2_19433 ( P3_ADD_318_U179 , P3_PHYADDRPOINTER_REG_11_ , P3_ADD_318_U22 );
nand NAND2_19434 ( P3_ADD_318_U180 , P3_ADD_318_U102 , P3_ADD_318_U23 );
nand NAND2_19435 ( P3_ADD_318_U181 , P3_PHYADDRPOINTER_REG_10_ , P3_ADD_318_U20 );
nand NAND2_19436 ( P3_ADD_318_U182 , P3_ADD_318_U101 , P3_ADD_318_U21 );
nand NAND2_19437 ( P3_SUB_370_U6 , P3_SUB_370_U45 , P3_SUB_370_U44 );
nand NAND2_19438 ( P3_SUB_370_U7 , P3_SUB_370_U9 , P3_SUB_370_U46 );
not NOT1_19439 ( P3_SUB_370_U8 , P3_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_19440 ( P3_SUB_370_U9 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_SUB_370_U18 );
not NOT1_19441 ( P3_SUB_370_U10 , P3_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_19442 ( P3_SUB_370_U11 , P3_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_19443 ( P3_SUB_370_U12 , P3_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_19444 ( P3_SUB_370_U13 , P3_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_19445 ( P3_SUB_370_U14 , P3_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_19446 ( P3_SUB_370_U15 , P3_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_19447 ( P3_SUB_370_U16 , P3_SUB_370_U41 , P3_SUB_370_U40 );
not NOT1_19448 ( P3_SUB_370_U17 , P3_INSTQUEUERD_ADDR_REG_4_ );
not NOT1_19449 ( P3_SUB_370_U18 , P3_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_19450 ( P3_SUB_370_U19 , P3_SUB_370_U51 , P3_SUB_370_U50 );
nand NAND2_19451 ( P3_SUB_370_U20 , P3_SUB_370_U56 , P3_SUB_370_U55 );
nand NAND2_19452 ( P3_SUB_370_U21 , P3_SUB_370_U61 , P3_SUB_370_U60 );
nand NAND2_19453 ( P3_SUB_370_U22 , P3_SUB_370_U66 , P3_SUB_370_U65 );
nand NAND2_19454 ( P3_SUB_370_U23 , P3_SUB_370_U48 , P3_SUB_370_U47 );
nand NAND2_19455 ( P3_SUB_370_U24 , P3_SUB_370_U53 , P3_SUB_370_U52 );
nand NAND2_19456 ( P3_SUB_370_U25 , P3_SUB_370_U58 , P3_SUB_370_U57 );
nand NAND2_19457 ( P3_SUB_370_U26 , P3_SUB_370_U63 , P3_SUB_370_U62 );
nand NAND2_19458 ( P3_SUB_370_U27 , P3_SUB_370_U37 , P3_SUB_370_U36 );
nand NAND2_19459 ( P3_SUB_370_U28 , P3_SUB_370_U33 , P3_SUB_370_U32 );
not NOT1_19460 ( P3_SUB_370_U29 , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_19461 ( P3_SUB_370_U30 , P3_SUB_370_U9 );
nand NAND2_19462 ( P3_SUB_370_U31 , P3_SUB_370_U30 , P3_SUB_370_U10 );
nand NAND2_19463 ( P3_SUB_370_U32 , P3_SUB_370_U31 , P3_SUB_370_U29 );
nand NAND2_19464 ( P3_SUB_370_U33 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_370_U9 );
not NOT1_19465 ( P3_SUB_370_U34 , P3_SUB_370_U28 );
nand NAND2_19466 ( P3_SUB_370_U35 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_370_U12 );
nand NAND2_19467 ( P3_SUB_370_U36 , P3_SUB_370_U35 , P3_SUB_370_U28 );
nand NAND2_19468 ( P3_SUB_370_U37 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_370_U11 );
not NOT1_19469 ( P3_SUB_370_U38 , P3_SUB_370_U27 );
nand NAND2_19470 ( P3_SUB_370_U39 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_370_U14 );
nand NAND2_19471 ( P3_SUB_370_U40 , P3_SUB_370_U39 , P3_SUB_370_U27 );
nand NAND2_19472 ( P3_SUB_370_U41 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_370_U13 );
not NOT1_19473 ( P3_SUB_370_U42 , P3_SUB_370_U16 );
nand NAND2_19474 ( P3_SUB_370_U43 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_370_U17 );
nand NAND2_19475 ( P3_SUB_370_U44 , P3_SUB_370_U42 , P3_SUB_370_U43 );
nand NAND2_19476 ( P3_SUB_370_U45 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_370_U15 );
nand NAND2_19477 ( P3_SUB_370_U46 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_SUB_370_U8 );
nand NAND2_19478 ( P3_SUB_370_U47 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_370_U15 );
nand NAND2_19479 ( P3_SUB_370_U48 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_370_U17 );
not NOT1_19480 ( P3_SUB_370_U49 , P3_SUB_370_U23 );
nand NAND2_19481 ( P3_SUB_370_U50 , P3_SUB_370_U49 , P3_SUB_370_U42 );
nand NAND2_19482 ( P3_SUB_370_U51 , P3_SUB_370_U23 , P3_SUB_370_U16 );
nand NAND2_19483 ( P3_SUB_370_U52 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_370_U14 );
nand NAND2_19484 ( P3_SUB_370_U53 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_370_U13 );
not NOT1_19485 ( P3_SUB_370_U54 , P3_SUB_370_U24 );
nand NAND2_19486 ( P3_SUB_370_U55 , P3_SUB_370_U38 , P3_SUB_370_U54 );
nand NAND2_19487 ( P3_SUB_370_U56 , P3_SUB_370_U24 , P3_SUB_370_U27 );
nand NAND2_19488 ( P3_SUB_370_U57 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_370_U12 );
nand NAND2_19489 ( P3_SUB_370_U58 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_370_U11 );
not NOT1_19490 ( P3_SUB_370_U59 , P3_SUB_370_U25 );
nand NAND2_19491 ( P3_SUB_370_U60 , P3_SUB_370_U34 , P3_SUB_370_U59 );
nand NAND2_19492 ( P3_SUB_370_U61 , P3_SUB_370_U25 , P3_SUB_370_U28 );
nand NAND2_19493 ( P3_SUB_370_U62 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_SUB_370_U10 );
nand NAND2_19494 ( P3_SUB_370_U63 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_370_U29 );
not NOT1_19495 ( P3_SUB_370_U64 , P3_SUB_370_U26 );
nand NAND2_19496 ( P3_SUB_370_U65 , P3_SUB_370_U64 , P3_SUB_370_U30 );
nand NAND2_19497 ( P3_SUB_370_U66 , P3_SUB_370_U26 , P3_SUB_370_U9 );
not NOT1_19498 ( P3_ADD_315_U4 , P3_PHYADDRPOINTER_REG_2_ );
not NOT1_19499 ( P3_ADD_315_U5 , P3_PHYADDRPOINTER_REG_3_ );
nand NAND2_19500 ( P3_ADD_315_U6 , P3_PHYADDRPOINTER_REG_3_ , P3_PHYADDRPOINTER_REG_2_ );
not NOT1_19501 ( P3_ADD_315_U7 , P3_PHYADDRPOINTER_REG_4_ );
nand NAND2_19502 ( P3_ADD_315_U8 , P3_PHYADDRPOINTER_REG_4_ , P3_ADD_315_U91 );
not NOT1_19503 ( P3_ADD_315_U9 , P3_PHYADDRPOINTER_REG_5_ );
nand NAND2_19504 ( P3_ADD_315_U10 , P3_PHYADDRPOINTER_REG_5_ , P3_ADD_315_U92 );
not NOT1_19505 ( P3_ADD_315_U11 , P3_PHYADDRPOINTER_REG_6_ );
nand NAND2_19506 ( P3_ADD_315_U12 , P3_PHYADDRPOINTER_REG_6_ , P3_ADD_315_U93 );
not NOT1_19507 ( P3_ADD_315_U13 , P3_PHYADDRPOINTER_REG_7_ );
nand NAND2_19508 ( P3_ADD_315_U14 , P3_PHYADDRPOINTER_REG_7_ , P3_ADD_315_U94 );
not NOT1_19509 ( P3_ADD_315_U15 , P3_PHYADDRPOINTER_REG_8_ );
not NOT1_19510 ( P3_ADD_315_U16 , P3_PHYADDRPOINTER_REG_9_ );
nand NAND2_19511 ( P3_ADD_315_U17 , P3_PHYADDRPOINTER_REG_8_ , P3_ADD_315_U95 );
nand NAND2_19512 ( P3_ADD_315_U18 , P3_ADD_315_U96 , P3_PHYADDRPOINTER_REG_9_ );
not NOT1_19513 ( P3_ADD_315_U19 , P3_PHYADDRPOINTER_REG_10_ );
nand NAND2_19514 ( P3_ADD_315_U20 , P3_PHYADDRPOINTER_REG_10_ , P3_ADD_315_U97 );
not NOT1_19515 ( P3_ADD_315_U21 , P3_PHYADDRPOINTER_REG_11_ );
nand NAND2_19516 ( P3_ADD_315_U22 , P3_PHYADDRPOINTER_REG_11_ , P3_ADD_315_U98 );
not NOT1_19517 ( P3_ADD_315_U23 , P3_PHYADDRPOINTER_REG_12_ );
nand NAND2_19518 ( P3_ADD_315_U24 , P3_PHYADDRPOINTER_REG_12_ , P3_ADD_315_U99 );
not NOT1_19519 ( P3_ADD_315_U25 , P3_PHYADDRPOINTER_REG_13_ );
nand NAND2_19520 ( P3_ADD_315_U26 , P3_PHYADDRPOINTER_REG_13_ , P3_ADD_315_U100 );
not NOT1_19521 ( P3_ADD_315_U27 , P3_PHYADDRPOINTER_REG_14_ );
nand NAND2_19522 ( P3_ADD_315_U28 , P3_PHYADDRPOINTER_REG_14_ , P3_ADD_315_U101 );
not NOT1_19523 ( P3_ADD_315_U29 , P3_PHYADDRPOINTER_REG_15_ );
nand NAND2_19524 ( P3_ADD_315_U30 , P3_PHYADDRPOINTER_REG_15_ , P3_ADD_315_U102 );
not NOT1_19525 ( P3_ADD_315_U31 , P3_PHYADDRPOINTER_REG_16_ );
nand NAND2_19526 ( P3_ADD_315_U32 , P3_PHYADDRPOINTER_REG_16_ , P3_ADD_315_U103 );
not NOT1_19527 ( P3_ADD_315_U33 , P3_PHYADDRPOINTER_REG_17_ );
nand NAND2_19528 ( P3_ADD_315_U34 , P3_PHYADDRPOINTER_REG_17_ , P3_ADD_315_U104 );
not NOT1_19529 ( P3_ADD_315_U35 , P3_PHYADDRPOINTER_REG_18_ );
nand NAND2_19530 ( P3_ADD_315_U36 , P3_PHYADDRPOINTER_REG_18_ , P3_ADD_315_U105 );
not NOT1_19531 ( P3_ADD_315_U37 , P3_PHYADDRPOINTER_REG_19_ );
nand NAND2_19532 ( P3_ADD_315_U38 , P3_PHYADDRPOINTER_REG_19_ , P3_ADD_315_U106 );
not NOT1_19533 ( P3_ADD_315_U39 , P3_PHYADDRPOINTER_REG_20_ );
nand NAND2_19534 ( P3_ADD_315_U40 , P3_PHYADDRPOINTER_REG_20_ , P3_ADD_315_U107 );
not NOT1_19535 ( P3_ADD_315_U41 , P3_PHYADDRPOINTER_REG_21_ );
nand NAND2_19536 ( P3_ADD_315_U42 , P3_PHYADDRPOINTER_REG_21_ , P3_ADD_315_U108 );
not NOT1_19537 ( P3_ADD_315_U43 , P3_PHYADDRPOINTER_REG_22_ );
nand NAND2_19538 ( P3_ADD_315_U44 , P3_PHYADDRPOINTER_REG_22_ , P3_ADD_315_U109 );
not NOT1_19539 ( P3_ADD_315_U45 , P3_PHYADDRPOINTER_REG_23_ );
nand NAND2_19540 ( P3_ADD_315_U46 , P3_PHYADDRPOINTER_REG_23_ , P3_ADD_315_U110 );
not NOT1_19541 ( P3_ADD_315_U47 , P3_PHYADDRPOINTER_REG_24_ );
nand NAND2_19542 ( P3_ADD_315_U48 , P3_PHYADDRPOINTER_REG_24_ , P3_ADD_315_U111 );
not NOT1_19543 ( P3_ADD_315_U49 , P3_PHYADDRPOINTER_REG_25_ );
nand NAND2_19544 ( P3_ADD_315_U50 , P3_PHYADDRPOINTER_REG_25_ , P3_ADD_315_U112 );
not NOT1_19545 ( P3_ADD_315_U51 , P3_PHYADDRPOINTER_REG_26_ );
nand NAND2_19546 ( P3_ADD_315_U52 , P3_PHYADDRPOINTER_REG_26_ , P3_ADD_315_U113 );
not NOT1_19547 ( P3_ADD_315_U53 , P3_PHYADDRPOINTER_REG_27_ );
nand NAND2_19548 ( P3_ADD_315_U54 , P3_PHYADDRPOINTER_REG_27_ , P3_ADD_315_U114 );
not NOT1_19549 ( P3_ADD_315_U55 , P3_PHYADDRPOINTER_REG_28_ );
nand NAND2_19550 ( P3_ADD_315_U56 , P3_PHYADDRPOINTER_REG_28_ , P3_ADD_315_U115 );
not NOT1_19551 ( P3_ADD_315_U57 , P3_PHYADDRPOINTER_REG_29_ );
nand NAND2_19552 ( P3_ADD_315_U58 , P3_PHYADDRPOINTER_REG_29_ , P3_ADD_315_U116 );
not NOT1_19553 ( P3_ADD_315_U59 , P3_PHYADDRPOINTER_REG_30_ );
nand NAND2_19554 ( P3_ADD_315_U60 , P3_ADD_315_U120 , P3_ADD_315_U119 );
nand NAND2_19555 ( P3_ADD_315_U61 , P3_ADD_315_U122 , P3_ADD_315_U121 );
nand NAND2_19556 ( P3_ADD_315_U62 , P3_ADD_315_U124 , P3_ADD_315_U123 );
nand NAND2_19557 ( P3_ADD_315_U63 , P3_ADD_315_U126 , P3_ADD_315_U125 );
nand NAND2_19558 ( P3_ADD_315_U64 , P3_ADD_315_U128 , P3_ADD_315_U127 );
nand NAND2_19559 ( P3_ADD_315_U65 , P3_ADD_315_U130 , P3_ADD_315_U129 );
nand NAND2_19560 ( P3_ADD_315_U66 , P3_ADD_315_U132 , P3_ADD_315_U131 );
nand NAND2_19561 ( P3_ADD_315_U67 , P3_ADD_315_U134 , P3_ADD_315_U133 );
nand NAND2_19562 ( P3_ADD_315_U68 , P3_ADD_315_U136 , P3_ADD_315_U135 );
nand NAND2_19563 ( P3_ADD_315_U69 , P3_ADD_315_U138 , P3_ADD_315_U137 );
nand NAND2_19564 ( P3_ADD_315_U70 , P3_ADD_315_U140 , P3_ADD_315_U139 );
nand NAND2_19565 ( P3_ADD_315_U71 , P3_ADD_315_U142 , P3_ADD_315_U141 );
nand NAND2_19566 ( P3_ADD_315_U72 , P3_ADD_315_U144 , P3_ADD_315_U143 );
nand NAND2_19567 ( P3_ADD_315_U73 , P3_ADD_315_U146 , P3_ADD_315_U145 );
nand NAND2_19568 ( P3_ADD_315_U74 , P3_ADD_315_U148 , P3_ADD_315_U147 );
nand NAND2_19569 ( P3_ADD_315_U75 , P3_ADD_315_U150 , P3_ADD_315_U149 );
nand NAND2_19570 ( P3_ADD_315_U76 , P3_ADD_315_U152 , P3_ADD_315_U151 );
nand NAND2_19571 ( P3_ADD_315_U77 , P3_ADD_315_U154 , P3_ADD_315_U153 );
nand NAND2_19572 ( P3_ADD_315_U78 , P3_ADD_315_U156 , P3_ADD_315_U155 );
nand NAND2_19573 ( P3_ADD_315_U79 , P3_ADD_315_U158 , P3_ADD_315_U157 );
nand NAND2_19574 ( P3_ADD_315_U80 , P3_ADD_315_U160 , P3_ADD_315_U159 );
nand NAND2_19575 ( P3_ADD_315_U81 , P3_ADD_315_U162 , P3_ADD_315_U161 );
nand NAND2_19576 ( P3_ADD_315_U82 , P3_ADD_315_U164 , P3_ADD_315_U163 );
nand NAND2_19577 ( P3_ADD_315_U83 , P3_ADD_315_U166 , P3_ADD_315_U165 );
nand NAND2_19578 ( P3_ADD_315_U84 , P3_ADD_315_U168 , P3_ADD_315_U167 );
nand NAND2_19579 ( P3_ADD_315_U85 , P3_ADD_315_U170 , P3_ADD_315_U169 );
nand NAND2_19580 ( P3_ADD_315_U86 , P3_ADD_315_U172 , P3_ADD_315_U171 );
nand NAND2_19581 ( P3_ADD_315_U87 , P3_ADD_315_U174 , P3_ADD_315_U173 );
nand NAND2_19582 ( P3_ADD_315_U88 , P3_ADD_315_U176 , P3_ADD_315_U175 );
not NOT1_19583 ( P3_ADD_315_U89 , P3_PHYADDRPOINTER_REG_31_ );
nand NAND2_19584 ( P3_ADD_315_U90 , P3_PHYADDRPOINTER_REG_30_ , P3_ADD_315_U117 );
not NOT1_19585 ( P3_ADD_315_U91 , P3_ADD_315_U6 );
not NOT1_19586 ( P3_ADD_315_U92 , P3_ADD_315_U8 );
not NOT1_19587 ( P3_ADD_315_U93 , P3_ADD_315_U10 );
not NOT1_19588 ( P3_ADD_315_U94 , P3_ADD_315_U12 );
not NOT1_19589 ( P3_ADD_315_U95 , P3_ADD_315_U14 );
not NOT1_19590 ( P3_ADD_315_U96 , P3_ADD_315_U17 );
not NOT1_19591 ( P3_ADD_315_U97 , P3_ADD_315_U18 );
not NOT1_19592 ( P3_ADD_315_U98 , P3_ADD_315_U20 );
not NOT1_19593 ( P3_ADD_315_U99 , P3_ADD_315_U22 );
not NOT1_19594 ( P3_ADD_315_U100 , P3_ADD_315_U24 );
not NOT1_19595 ( P3_ADD_315_U101 , P3_ADD_315_U26 );
not NOT1_19596 ( P3_ADD_315_U102 , P3_ADD_315_U28 );
not NOT1_19597 ( P3_ADD_315_U103 , P3_ADD_315_U30 );
not NOT1_19598 ( P3_ADD_315_U104 , P3_ADD_315_U32 );
not NOT1_19599 ( P3_ADD_315_U105 , P3_ADD_315_U34 );
not NOT1_19600 ( P3_ADD_315_U106 , P3_ADD_315_U36 );
not NOT1_19601 ( P3_ADD_315_U107 , P3_ADD_315_U38 );
not NOT1_19602 ( P3_ADD_315_U108 , P3_ADD_315_U40 );
not NOT1_19603 ( P3_ADD_315_U109 , P3_ADD_315_U42 );
not NOT1_19604 ( P3_ADD_315_U110 , P3_ADD_315_U44 );
not NOT1_19605 ( P3_ADD_315_U111 , P3_ADD_315_U46 );
not NOT1_19606 ( P3_ADD_315_U112 , P3_ADD_315_U48 );
not NOT1_19607 ( P3_ADD_315_U113 , P3_ADD_315_U50 );
not NOT1_19608 ( P3_ADD_315_U114 , P3_ADD_315_U52 );
not NOT1_19609 ( P3_ADD_315_U115 , P3_ADD_315_U54 );
not NOT1_19610 ( P3_ADD_315_U116 , P3_ADD_315_U56 );
not NOT1_19611 ( P3_ADD_315_U117 , P3_ADD_315_U58 );
not NOT1_19612 ( P3_ADD_315_U118 , P3_ADD_315_U90 );
nand NAND2_19613 ( P3_ADD_315_U119 , P3_PHYADDRPOINTER_REG_9_ , P3_ADD_315_U17 );
nand NAND2_19614 ( P3_ADD_315_U120 , P3_ADD_315_U96 , P3_ADD_315_U16 );
nand NAND2_19615 ( P3_ADD_315_U121 , P3_PHYADDRPOINTER_REG_8_ , P3_ADD_315_U14 );
nand NAND2_19616 ( P3_ADD_315_U122 , P3_ADD_315_U95 , P3_ADD_315_U15 );
nand NAND2_19617 ( P3_ADD_315_U123 , P3_PHYADDRPOINTER_REG_7_ , P3_ADD_315_U12 );
nand NAND2_19618 ( P3_ADD_315_U124 , P3_ADD_315_U94 , P3_ADD_315_U13 );
nand NAND2_19619 ( P3_ADD_315_U125 , P3_PHYADDRPOINTER_REG_6_ , P3_ADD_315_U10 );
nand NAND2_19620 ( P3_ADD_315_U126 , P3_ADD_315_U93 , P3_ADD_315_U11 );
nand NAND2_19621 ( P3_ADD_315_U127 , P3_PHYADDRPOINTER_REG_5_ , P3_ADD_315_U8 );
nand NAND2_19622 ( P3_ADD_315_U128 , P3_ADD_315_U92 , P3_ADD_315_U9 );
nand NAND2_19623 ( P3_ADD_315_U129 , P3_PHYADDRPOINTER_REG_4_ , P3_ADD_315_U6 );
nand NAND2_19624 ( P3_ADD_315_U130 , P3_ADD_315_U91 , P3_ADD_315_U7 );
nand NAND2_19625 ( P3_ADD_315_U131 , P3_PHYADDRPOINTER_REG_3_ , P3_ADD_315_U4 );
nand NAND2_19626 ( P3_ADD_315_U132 , P3_PHYADDRPOINTER_REG_2_ , P3_ADD_315_U5 );
nand NAND2_19627 ( P3_ADD_315_U133 , P3_PHYADDRPOINTER_REG_31_ , P3_ADD_315_U90 );
nand NAND2_19628 ( P3_ADD_315_U134 , P3_ADD_315_U118 , P3_ADD_315_U89 );
nand NAND2_19629 ( P3_ADD_315_U135 , P3_PHYADDRPOINTER_REG_30_ , P3_ADD_315_U58 );
nand NAND2_19630 ( P3_ADD_315_U136 , P3_ADD_315_U117 , P3_ADD_315_U59 );
nand NAND2_19631 ( P3_ADD_315_U137 , P3_PHYADDRPOINTER_REG_29_ , P3_ADD_315_U56 );
nand NAND2_19632 ( P3_ADD_315_U138 , P3_ADD_315_U116 , P3_ADD_315_U57 );
nand NAND2_19633 ( P3_ADD_315_U139 , P3_PHYADDRPOINTER_REG_28_ , P3_ADD_315_U54 );
nand NAND2_19634 ( P3_ADD_315_U140 , P3_ADD_315_U115 , P3_ADD_315_U55 );
nand NAND2_19635 ( P3_ADD_315_U141 , P3_PHYADDRPOINTER_REG_27_ , P3_ADD_315_U52 );
nand NAND2_19636 ( P3_ADD_315_U142 , P3_ADD_315_U114 , P3_ADD_315_U53 );
nand NAND2_19637 ( P3_ADD_315_U143 , P3_PHYADDRPOINTER_REG_26_ , P3_ADD_315_U50 );
nand NAND2_19638 ( P3_ADD_315_U144 , P3_ADD_315_U113 , P3_ADD_315_U51 );
nand NAND2_19639 ( P3_ADD_315_U145 , P3_PHYADDRPOINTER_REG_25_ , P3_ADD_315_U48 );
nand NAND2_19640 ( P3_ADD_315_U146 , P3_ADD_315_U112 , P3_ADD_315_U49 );
nand NAND2_19641 ( P3_ADD_315_U147 , P3_PHYADDRPOINTER_REG_24_ , P3_ADD_315_U46 );
nand NAND2_19642 ( P3_ADD_315_U148 , P3_ADD_315_U111 , P3_ADD_315_U47 );
nand NAND2_19643 ( P3_ADD_315_U149 , P3_PHYADDRPOINTER_REG_23_ , P3_ADD_315_U44 );
nand NAND2_19644 ( P3_ADD_315_U150 , P3_ADD_315_U110 , P3_ADD_315_U45 );
nand NAND2_19645 ( P3_ADD_315_U151 , P3_PHYADDRPOINTER_REG_22_ , P3_ADD_315_U42 );
nand NAND2_19646 ( P3_ADD_315_U152 , P3_ADD_315_U109 , P3_ADD_315_U43 );
nand NAND2_19647 ( P3_ADD_315_U153 , P3_PHYADDRPOINTER_REG_21_ , P3_ADD_315_U40 );
nand NAND2_19648 ( P3_ADD_315_U154 , P3_ADD_315_U108 , P3_ADD_315_U41 );
nand NAND2_19649 ( P3_ADD_315_U155 , P3_PHYADDRPOINTER_REG_20_ , P3_ADD_315_U38 );
nand NAND2_19650 ( P3_ADD_315_U156 , P3_ADD_315_U107 , P3_ADD_315_U39 );
nand NAND2_19651 ( P3_ADD_315_U157 , P3_PHYADDRPOINTER_REG_19_ , P3_ADD_315_U36 );
nand NAND2_19652 ( P3_ADD_315_U158 , P3_ADD_315_U106 , P3_ADD_315_U37 );
nand NAND2_19653 ( P3_ADD_315_U159 , P3_PHYADDRPOINTER_REG_18_ , P3_ADD_315_U34 );
nand NAND2_19654 ( P3_ADD_315_U160 , P3_ADD_315_U105 , P3_ADD_315_U35 );
nand NAND2_19655 ( P3_ADD_315_U161 , P3_PHYADDRPOINTER_REG_17_ , P3_ADD_315_U32 );
nand NAND2_19656 ( P3_ADD_315_U162 , P3_ADD_315_U104 , P3_ADD_315_U33 );
nand NAND2_19657 ( P3_ADD_315_U163 , P3_PHYADDRPOINTER_REG_16_ , P3_ADD_315_U30 );
nand NAND2_19658 ( P3_ADD_315_U164 , P3_ADD_315_U103 , P3_ADD_315_U31 );
nand NAND2_19659 ( P3_ADD_315_U165 , P3_PHYADDRPOINTER_REG_15_ , P3_ADD_315_U28 );
nand NAND2_19660 ( P3_ADD_315_U166 , P3_ADD_315_U102 , P3_ADD_315_U29 );
nand NAND2_19661 ( P3_ADD_315_U167 , P3_PHYADDRPOINTER_REG_14_ , P3_ADD_315_U26 );
nand NAND2_19662 ( P3_ADD_315_U168 , P3_ADD_315_U101 , P3_ADD_315_U27 );
nand NAND2_19663 ( P3_ADD_315_U169 , P3_PHYADDRPOINTER_REG_13_ , P3_ADD_315_U24 );
nand NAND2_19664 ( P3_ADD_315_U170 , P3_ADD_315_U100 , P3_ADD_315_U25 );
nand NAND2_19665 ( P3_ADD_315_U171 , P3_PHYADDRPOINTER_REG_12_ , P3_ADD_315_U22 );
nand NAND2_19666 ( P3_ADD_315_U172 , P3_ADD_315_U99 , P3_ADD_315_U23 );
nand NAND2_19667 ( P3_ADD_315_U173 , P3_PHYADDRPOINTER_REG_11_ , P3_ADD_315_U20 );
nand NAND2_19668 ( P3_ADD_315_U174 , P3_ADD_315_U98 , P3_ADD_315_U21 );
nand NAND2_19669 ( P3_ADD_315_U175 , P3_PHYADDRPOINTER_REG_10_ , P3_ADD_315_U18 );
nand NAND2_19670 ( P3_ADD_315_U176 , P3_ADD_315_U97 , P3_ADD_315_U19 );
nor nor_19671 ( P3_GTE_355_U6 , P3_SUB_355_U6 , P3_GTE_355_U8 );
and AND2_19672 ( P3_GTE_355_U7 , P3_SUB_355_U7 , P3_SUB_355_U22 );
nor nor_19673 ( P3_GTE_355_U8 , P3_SUB_355_U19 , P3_SUB_355_U20 , P3_GTE_355_U7 , P3_SUB_355_U21 );
and AND2_19674 ( P3_ADD_360_1242_U4 , P3_ADD_360_1242_U186 , P3_ADD_360_1242_U45 );
and AND2_19675 ( P3_ADD_360_1242_U5 , P3_ADD_360_1242_U184 , P3_ADD_360_1242_U46 );
and AND2_19676 ( P3_ADD_360_1242_U6 , P3_ADD_360_1242_U182 , P3_ADD_360_1242_U76 );
and AND2_19677 ( P3_ADD_360_1242_U7 , P3_ADD_360_1242_U181 , P3_ADD_360_1242_U50 );
and AND2_19678 ( P3_ADD_360_1242_U8 , P3_ADD_360_1242_U179 , P3_ADD_360_1242_U53 );
and AND2_19679 ( P3_ADD_360_1242_U9 , P3_ADD_360_1242_U177 , P3_ADD_360_1242_U56 );
and AND2_19680 ( P3_ADD_360_1242_U10 , P3_ADD_360_1242_U175 , P3_ADD_360_1242_U58 );
and AND2_19681 ( P3_ADD_360_1242_U11 , P3_ADD_360_1242_U174 , P3_ADD_360_1242_U60 );
and AND2_19682 ( P3_ADD_360_1242_U12 , P3_ADD_360_1242_U173 , P3_ADD_360_1242_U63 );
and AND2_19683 ( P3_ADD_360_1242_U13 , P3_ADD_360_1242_U171 , P3_ADD_360_1242_U66 );
and AND2_19684 ( P3_ADD_360_1242_U14 , P3_ADD_360_1242_U169 , P3_ADD_360_1242_U68 );
and AND2_19685 ( P3_ADD_360_1242_U15 , P3_ADD_360_1242_U168 , P3_ADD_360_1242_U71 );
and AND2_19686 ( P3_ADD_360_1242_U16 , P3_ADD_360_1242_U166 , P3_ADD_360_1242_U73 );
and AND2_19687 ( P3_ADD_360_1242_U17 , P3_ADD_360_1242_U153 , P3_ADD_360_1242_U152 );
and AND2_19688 ( P3_ADD_360_1242_U18 , P3_ADD_360_1242_U151 , P3_ADD_360_1242_U149 );
nand NAND3_19689 ( P3_ADD_360_1242_U19 , P3_ADD_360_1242_U248 , P3_ADD_360_1242_U247 , P3_ADD_360_1242_U192 );
not NOT1_19690 ( P3_ADD_360_1242_U20 , P3_ADD_360_U19 );
not NOT1_19691 ( P3_ADD_360_1242_U21 , P3_INSTADDRPOINTER_REG_4_ );
not NOT1_19692 ( P3_ADD_360_1242_U22 , P3_ADD_360_U20 );
not NOT1_19693 ( P3_ADD_360_1242_U23 , P3_INSTADDRPOINTER_REG_3_ );
not NOT1_19694 ( P3_ADD_360_1242_U24 , P3_U2621 );
not NOT1_19695 ( P3_ADD_360_1242_U25 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_19696 ( P3_ADD_360_1242_U26 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_19697 ( P3_ADD_360_1242_U27 , P3_INSTADDRPOINTER_REG_0_ , P3_U2621 );
not NOT1_19698 ( P3_ADD_360_1242_U28 , P3_ADD_360_U4 );
not NOT1_19699 ( P3_ADD_360_1242_U29 , P3_ADD_360_U21 );
not NOT1_19700 ( P3_ADD_360_1242_U30 , P3_INSTADDRPOINTER_REG_2_ );
not NOT1_19701 ( P3_ADD_360_1242_U31 , P3_INSTADDRPOINTER_REG_5_ );
not NOT1_19702 ( P3_ADD_360_1242_U32 , P3_ADD_360_U18 );
not NOT1_19703 ( P3_ADD_360_1242_U33 , P3_ADD_360_U17 );
not NOT1_19704 ( P3_ADD_360_1242_U34 , P3_INSTADDRPOINTER_REG_6_ );
not NOT1_19705 ( P3_ADD_360_1242_U35 , P3_INSTADDRPOINTER_REG_7_ );
not NOT1_19706 ( P3_ADD_360_1242_U36 , P3_ADD_360_U16 );
not NOT1_19707 ( P3_ADD_360_1242_U37 , P3_ADD_360_U5 );
not NOT1_19708 ( P3_ADD_360_1242_U38 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_19709 ( P3_ADD_360_1242_U39 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_19710 ( P3_ADD_360_1242_U40 , P3_ADD_360_1242_U131 , P3_ADD_360_1242_U130 );
nand NAND2_19711 ( P3_ADD_360_1242_U41 , P3_ADD_360_1242_U40 , P3_ADD_360_1242_U133 );
not NOT1_19712 ( P3_ADD_360_1242_U42 , P3_INSTADDRPOINTER_REG_10_ );
not NOT1_19713 ( P3_ADD_360_1242_U43 , P3_INSTADDRPOINTER_REG_11_ );
not NOT1_19714 ( P3_ADD_360_1242_U44 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_19715 ( P3_ADD_360_1242_U45 , P3_ADD_360_1242_U97 , P3_ADD_360_1242_U105 );
nand NAND2_19716 ( P3_ADD_360_1242_U46 , P3_ADD_360_1242_U98 , P3_ADD_360_1242_U119 );
not NOT1_19717 ( P3_ADD_360_1242_U47 , P3_INSTADDRPOINTER_REG_13_ );
not NOT1_19718 ( P3_ADD_360_1242_U48 , P3_INSTADDRPOINTER_REG_15_ );
not NOT1_19719 ( P3_ADD_360_1242_U49 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_19720 ( P3_ADD_360_1242_U50 , P3_ADD_360_1242_U154 , P3_ADD_360_1242_U99 );
not NOT1_19721 ( P3_ADD_360_1242_U51 , P3_INSTADDRPOINTER_REG_17_ );
not NOT1_19722 ( P3_ADD_360_1242_U52 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_19723 ( P3_ADD_360_1242_U53 , P3_ADD_360_1242_U100 , P3_ADD_360_1242_U156 );
not NOT1_19724 ( P3_ADD_360_1242_U54 , P3_INSTADDRPOINTER_REG_18_ );
not NOT1_19725 ( P3_ADD_360_1242_U55 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_19726 ( P3_ADD_360_1242_U56 , P3_ADD_360_1242_U101 , P3_ADD_360_1242_U157 );
not NOT1_19727 ( P3_ADD_360_1242_U57 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_19728 ( P3_ADD_360_1242_U58 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_360_1242_U158 );
not NOT1_19729 ( P3_ADD_360_1242_U59 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_19730 ( P3_ADD_360_1242_U60 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_360_1242_U159 );
not NOT1_19731 ( P3_ADD_360_1242_U61 , P3_INSTADDRPOINTER_REG_23_ );
not NOT1_19732 ( P3_ADD_360_1242_U62 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_19733 ( P3_ADD_360_1242_U63 , P3_ADD_360_1242_U102 , P3_ADD_360_1242_U160 );
not NOT1_19734 ( P3_ADD_360_1242_U64 , P3_INSTADDRPOINTER_REG_25_ );
not NOT1_19735 ( P3_ADD_360_1242_U65 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_19736 ( P3_ADD_360_1242_U66 , P3_ADD_360_1242_U103 , P3_ADD_360_1242_U161 );
not NOT1_19737 ( P3_ADD_360_1242_U67 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_19738 ( P3_ADD_360_1242_U68 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_360_1242_U162 );
not NOT1_19739 ( P3_ADD_360_1242_U69 , P3_INSTADDRPOINTER_REG_28_ );
not NOT1_19740 ( P3_ADD_360_1242_U70 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_19741 ( P3_ADD_360_1242_U71 , P3_ADD_360_1242_U104 , P3_ADD_360_1242_U163 );
not NOT1_19742 ( P3_ADD_360_1242_U72 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_19743 ( P3_ADD_360_1242_U73 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_360_1242_U164 );
not NOT1_19744 ( P3_ADD_360_1242_U74 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_19745 ( P3_ADD_360_1242_U75 , P3_ADD_360_U4 , P3_ADD_360_1242_U124 );
nand NAND2_19746 ( P3_ADD_360_1242_U76 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_360_1242_U154 );
nand NAND2_19747 ( P3_ADD_360_1242_U77 , P3_ADD_360_1242_U230 , P3_ADD_360_1242_U229 );
nand NAND2_19748 ( P3_ADD_360_1242_U78 , P3_ADD_360_1242_U239 , P3_ADD_360_1242_U238 );
nand NAND2_19749 ( P3_ADD_360_1242_U79 , P3_ADD_360_1242_U241 , P3_ADD_360_1242_U240 );
nand NAND2_19750 ( P3_ADD_360_1242_U80 , P3_ADD_360_1242_U243 , P3_ADD_360_1242_U242 );
nand NAND2_19751 ( P3_ADD_360_1242_U81 , P3_ADD_360_1242_U250 , P3_ADD_360_1242_U249 );
nand NAND2_19752 ( P3_ADD_360_1242_U82 , P3_ADD_360_1242_U252 , P3_ADD_360_1242_U251 );
nand NAND2_19753 ( P3_ADD_360_1242_U83 , P3_ADD_360_1242_U254 , P3_ADD_360_1242_U253 );
nand NAND2_19754 ( P3_ADD_360_1242_U84 , P3_ADD_360_1242_U256 , P3_ADD_360_1242_U255 );
nand NAND2_19755 ( P3_ADD_360_1242_U85 , P3_ADD_360_1242_U258 , P3_ADD_360_1242_U257 );
nand NAND2_19756 ( P3_ADD_360_1242_U86 , P3_ADD_360_1242_U201 , P3_ADD_360_1242_U200 );
nand NAND2_19757 ( P3_ADD_360_1242_U87 , P3_ADD_360_1242_U208 , P3_ADD_360_1242_U207 );
nand NAND2_19758 ( P3_ADD_360_1242_U88 , P3_ADD_360_1242_U215 , P3_ADD_360_1242_U214 );
nand NAND2_19759 ( P3_ADD_360_1242_U89 , P3_ADD_360_1242_U222 , P3_ADD_360_1242_U221 );
nand NAND2_19760 ( P3_ADD_360_1242_U90 , P3_ADD_360_1242_U228 , P3_ADD_360_1242_U227 );
nand NAND2_19761 ( P3_ADD_360_1242_U91 , P3_ADD_360_1242_U237 , P3_ADD_360_1242_U236 );
and AND2_19762 ( P3_ADD_360_1242_U92 , P3_ADD_360_U20 , P3_INSTADDRPOINTER_REG_3_ );
and AND2_19763 ( P3_ADD_360_1242_U93 , P3_ADD_360_1242_U133 , P3_ADD_360_1242_U123 );
and AND2_19764 ( P3_ADD_360_1242_U94 , P3_ADD_360_1242_U190 , P3_ADD_360_1242_U125 );
and AND3_19765 ( P3_ADD_360_1242_U95 , P3_ADD_360_1242_U224 , P3_ADD_360_1242_U223 , P3_ADD_360_1242_U135 );
and AND2_19766 ( P3_ADD_360_1242_U96 , P3_ADD_360_1242_U125 , P3_ADD_360_1242_U123 );
and AND2_19767 ( P3_ADD_360_1242_U97 , P3_INSTADDRPOINTER_REG_9_ , P3_INSTADDRPOINTER_REG_10_ );
and AND2_19768 ( P3_ADD_360_1242_U98 , P3_INSTADDRPOINTER_REG_12_ , P3_INSTADDRPOINTER_REG_11_ );
and AND3_19769 ( P3_ADD_360_1242_U99 , P3_INSTADDRPOINTER_REG_14_ , P3_INSTADDRPOINTER_REG_15_ , P3_INSTADDRPOINTER_REG_13_ );
and AND2_19770 ( P3_ADD_360_1242_U100 , P3_INSTADDRPOINTER_REG_17_ , P3_INSTADDRPOINTER_REG_16_ );
and AND2_19771 ( P3_ADD_360_1242_U101 , P3_INSTADDRPOINTER_REG_18_ , P3_INSTADDRPOINTER_REG_19_ );
and AND2_19772 ( P3_ADD_360_1242_U102 , P3_INSTADDRPOINTER_REG_23_ , P3_INSTADDRPOINTER_REG_22_ );
and AND2_19773 ( P3_ADD_360_1242_U103 , P3_INSTADDRPOINTER_REG_25_ , P3_INSTADDRPOINTER_REG_24_ );
and AND2_19774 ( P3_ADD_360_1242_U104 , P3_INSTADDRPOINTER_REG_28_ , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_19775 ( P3_ADD_360_1242_U105 , P3_ADD_360_1242_U147 , P3_ADD_360_1242_U146 );
and AND2_19776 ( P3_ADD_360_1242_U106 , P3_ADD_360_1242_U194 , P3_ADD_360_1242_U193 );
and AND2_19777 ( P3_ADD_360_1242_U107 , P3_ADD_360_1242_U196 , P3_ADD_360_1242_U195 );
nand NAND3_19778 ( P3_ADD_360_1242_U108 , P3_ADD_360_1242_U143 , P3_ADD_360_1242_U120 , P3_ADD_360_1242_U189 );
and AND2_19779 ( P3_ADD_360_1242_U109 , P3_ADD_360_1242_U203 , P3_ADD_360_1242_U202 );
nand NAND2_19780 ( P3_ADD_360_1242_U110 , P3_ADD_360_1242_U141 , P3_ADD_360_1242_U140 );
and AND2_19781 ( P3_ADD_360_1242_U111 , P3_ADD_360_1242_U210 , P3_ADD_360_1242_U209 );
nand NAND3_19782 ( P3_ADD_360_1242_U112 , P3_ADD_360_1242_U137 , P3_ADD_360_1242_U121 , P3_ADD_360_1242_U188 );
and AND2_19783 ( P3_ADD_360_1242_U113 , P3_ADD_360_1242_U217 , P3_ADD_360_1242_U216 );
nand NAND2_19784 ( P3_ADD_360_1242_U114 , P3_ADD_360_1242_U94 , P3_ADD_360_1242_U191 );
and AND2_19785 ( P3_ADD_360_1242_U115 , P3_ADD_360_1242_U226 , P3_ADD_360_1242_U225 );
not NOT1_19786 ( P3_ADD_360_1242_U116 , P3_INSTADDRPOINTER_REG_31_ );
and AND2_19787 ( P3_ADD_360_1242_U117 , P3_ADD_360_1242_U232 , P3_ADD_360_1242_U231 );
nand NAND2_19788 ( P3_ADD_360_1242_U118 , P3_ADD_360_1242_U75 , P3_ADD_360_1242_U127 );
not NOT1_19789 ( P3_ADD_360_1242_U119 , P3_ADD_360_1242_U45 );
nand NAND2_19790 ( P3_ADD_360_1242_U120 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_360_1242_U110 );
nand NAND2_19791 ( P3_ADD_360_1242_U121 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_360_1242_U114 );
not NOT1_19792 ( P3_ADD_360_1242_U122 , P3_ADD_360_1242_U75 );
or OR2_19793 ( P3_ADD_360_1242_U123 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_360_U19 );
not NOT1_19794 ( P3_ADD_360_1242_U124 , P3_ADD_360_1242_U27 );
nand NAND2_19795 ( P3_ADD_360_1242_U125 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_360_U19 );
nand NAND2_19796 ( P3_ADD_360_1242_U126 , P3_ADD_360_1242_U28 , P3_ADD_360_1242_U27 );
nand NAND2_19797 ( P3_ADD_360_1242_U127 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_360_1242_U126 );
not NOT1_19798 ( P3_ADD_360_1242_U128 , P3_ADD_360_1242_U118 );
or OR2_19799 ( P3_ADD_360_1242_U129 , P3_ADD_360_U21 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_19800 ( P3_ADD_360_1242_U130 , P3_ADD_360_1242_U129 , P3_ADD_360_1242_U118 );
nand NAND2_19801 ( P3_ADD_360_1242_U131 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_360_U21 );
not NOT1_19802 ( P3_ADD_360_1242_U132 , P3_ADD_360_1242_U40 );
or OR2_19803 ( P3_ADD_360_1242_U133 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_360_U20 );
not NOT1_19804 ( P3_ADD_360_1242_U134 , P3_ADD_360_1242_U41 );
nand NAND2_19805 ( P3_ADD_360_1242_U135 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_360_U20 );
not NOT1_19806 ( P3_ADD_360_1242_U136 , P3_ADD_360_1242_U114 );
nand NAND2_19807 ( P3_ADD_360_1242_U137 , P3_ADD_360_U18 , P3_ADD_360_1242_U114 );
not NOT1_19808 ( P3_ADD_360_1242_U138 , P3_ADD_360_1242_U112 );
or OR2_19809 ( P3_ADD_360_1242_U139 , P3_ADD_360_U17 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_19810 ( P3_ADD_360_1242_U140 , P3_ADD_360_1242_U139 , P3_ADD_360_1242_U112 );
nand NAND2_19811 ( P3_ADD_360_1242_U141 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_360_U17 );
not NOT1_19812 ( P3_ADD_360_1242_U142 , P3_ADD_360_1242_U110 );
nand NAND2_19813 ( P3_ADD_360_1242_U143 , P3_ADD_360_U16 , P3_ADD_360_1242_U110 );
not NOT1_19814 ( P3_ADD_360_1242_U144 , P3_ADD_360_1242_U108 );
or OR2_19815 ( P3_ADD_360_1242_U145 , P3_ADD_360_U5 , P3_INSTADDRPOINTER_REG_8_ );
nand NAND2_19816 ( P3_ADD_360_1242_U146 , P3_ADD_360_1242_U145 , P3_ADD_360_1242_U108 );
nand NAND2_19817 ( P3_ADD_360_1242_U147 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_360_U5 );
not NOT1_19818 ( P3_ADD_360_1242_U148 , P3_ADD_360_1242_U105 );
nand NAND2_19819 ( P3_ADD_360_1242_U149 , P3_ADD_360_1242_U95 , P3_ADD_360_1242_U41 );
nand NAND2_19820 ( P3_ADD_360_1242_U150 , P3_ADD_360_1242_U135 , P3_ADD_360_1242_U41 );
nand NAND2_19821 ( P3_ADD_360_1242_U151 , P3_ADD_360_1242_U96 , P3_ADD_360_1242_U150 );
nand NAND2_19822 ( P3_ADD_360_1242_U152 , P3_ADD_360_1242_U115 , P3_ADD_360_1242_U132 );
nand NAND2_19823 ( P3_ADD_360_1242_U153 , P3_ADD_360_1242_U134 , P3_ADD_360_1242_U135 );
not NOT1_19824 ( P3_ADD_360_1242_U154 , P3_ADD_360_1242_U46 );
not NOT1_19825 ( P3_ADD_360_1242_U155 , P3_ADD_360_1242_U76 );
not NOT1_19826 ( P3_ADD_360_1242_U156 , P3_ADD_360_1242_U50 );
not NOT1_19827 ( P3_ADD_360_1242_U157 , P3_ADD_360_1242_U53 );
not NOT1_19828 ( P3_ADD_360_1242_U158 , P3_ADD_360_1242_U56 );
not NOT1_19829 ( P3_ADD_360_1242_U159 , P3_ADD_360_1242_U58 );
not NOT1_19830 ( P3_ADD_360_1242_U160 , P3_ADD_360_1242_U60 );
not NOT1_19831 ( P3_ADD_360_1242_U161 , P3_ADD_360_1242_U63 );
not NOT1_19832 ( P3_ADD_360_1242_U162 , P3_ADD_360_1242_U66 );
not NOT1_19833 ( P3_ADD_360_1242_U163 , P3_ADD_360_1242_U68 );
not NOT1_19834 ( P3_ADD_360_1242_U164 , P3_ADD_360_1242_U71 );
not NOT1_19835 ( P3_ADD_360_1242_U165 , P3_ADD_360_1242_U73 );
nand NAND2_19836 ( P3_ADD_360_1242_U166 , P3_ADD_360_1242_U72 , P3_ADD_360_1242_U71 );
nand NAND2_19837 ( P3_ADD_360_1242_U167 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_360_1242_U163 );
nand NAND2_19838 ( P3_ADD_360_1242_U168 , P3_ADD_360_1242_U69 , P3_ADD_360_1242_U167 );
nand NAND2_19839 ( P3_ADD_360_1242_U169 , P3_ADD_360_1242_U67 , P3_ADD_360_1242_U66 );
nand NAND2_19840 ( P3_ADD_360_1242_U170 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_360_1242_U161 );
nand NAND2_19841 ( P3_ADD_360_1242_U171 , P3_ADD_360_1242_U64 , P3_ADD_360_1242_U170 );
nand NAND2_19842 ( P3_ADD_360_1242_U172 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_360_1242_U160 );
nand NAND2_19843 ( P3_ADD_360_1242_U173 , P3_ADD_360_1242_U61 , P3_ADD_360_1242_U172 );
nand NAND2_19844 ( P3_ADD_360_1242_U174 , P3_ADD_360_1242_U59 , P3_ADD_360_1242_U58 );
nand NAND2_19845 ( P3_ADD_360_1242_U175 , P3_ADD_360_1242_U57 , P3_ADD_360_1242_U56 );
nand NAND2_19846 ( P3_ADD_360_1242_U176 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_360_1242_U157 );
nand NAND2_19847 ( P3_ADD_360_1242_U177 , P3_ADD_360_1242_U55 , P3_ADD_360_1242_U176 );
nand NAND2_19848 ( P3_ADD_360_1242_U178 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_360_1242_U156 );
nand NAND2_19849 ( P3_ADD_360_1242_U179 , P3_ADD_360_1242_U51 , P3_ADD_360_1242_U178 );
nand NAND2_19850 ( P3_ADD_360_1242_U180 , P3_ADD_360_1242_U155 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_19851 ( P3_ADD_360_1242_U181 , P3_ADD_360_1242_U48 , P3_ADD_360_1242_U180 );
nand NAND2_19852 ( P3_ADD_360_1242_U182 , P3_ADD_360_1242_U47 , P3_ADD_360_1242_U46 );
nand NAND2_19853 ( P3_ADD_360_1242_U183 , P3_ADD_360_1242_U119 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_19854 ( P3_ADD_360_1242_U184 , P3_ADD_360_1242_U44 , P3_ADD_360_1242_U183 );
nand NAND2_19855 ( P3_ADD_360_1242_U185 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_360_1242_U105 );
nand NAND2_19856 ( P3_ADD_360_1242_U186 , P3_ADD_360_1242_U42 , P3_ADD_360_1242_U185 );
nand NAND2_19857 ( P3_ADD_360_1242_U187 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_360_1242_U165 );
nand NAND2_19858 ( P3_ADD_360_1242_U188 , P3_ADD_360_U18 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_19859 ( P3_ADD_360_1242_U189 , P3_ADD_360_U16 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_19860 ( P3_ADD_360_1242_U190 , P3_ADD_360_1242_U92 , P3_ADD_360_1242_U123 );
nand NAND2_19861 ( P3_ADD_360_1242_U191 , P3_ADD_360_1242_U93 , P3_ADD_360_1242_U40 );
nand NAND2_19862 ( P3_ADD_360_1242_U192 , P3_ADD_360_1242_U122 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_19863 ( P3_ADD_360_1242_U193 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_360_1242_U105 );
nand NAND2_19864 ( P3_ADD_360_1242_U194 , P3_ADD_360_1242_U148 , P3_ADD_360_1242_U39 );
nand NAND2_19865 ( P3_ADD_360_1242_U195 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_360_1242_U37 );
nand NAND2_19866 ( P3_ADD_360_1242_U196 , P3_ADD_360_U5 , P3_ADD_360_1242_U38 );
nand NAND2_19867 ( P3_ADD_360_1242_U197 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_360_1242_U37 );
nand NAND2_19868 ( P3_ADD_360_1242_U198 , P3_ADD_360_U5 , P3_ADD_360_1242_U38 );
nand NAND2_19869 ( P3_ADD_360_1242_U199 , P3_ADD_360_1242_U198 , P3_ADD_360_1242_U197 );
nand NAND2_19870 ( P3_ADD_360_1242_U200 , P3_ADD_360_1242_U107 , P3_ADD_360_1242_U108 );
nand NAND2_19871 ( P3_ADD_360_1242_U201 , P3_ADD_360_1242_U144 , P3_ADD_360_1242_U199 );
nand NAND2_19872 ( P3_ADD_360_1242_U202 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_360_1242_U36 );
nand NAND2_19873 ( P3_ADD_360_1242_U203 , P3_ADD_360_U16 , P3_ADD_360_1242_U35 );
nand NAND2_19874 ( P3_ADD_360_1242_U204 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_360_1242_U36 );
nand NAND2_19875 ( P3_ADD_360_1242_U205 , P3_ADD_360_U16 , P3_ADD_360_1242_U35 );
nand NAND2_19876 ( P3_ADD_360_1242_U206 , P3_ADD_360_1242_U205 , P3_ADD_360_1242_U204 );
nand NAND2_19877 ( P3_ADD_360_1242_U207 , P3_ADD_360_1242_U109 , P3_ADD_360_1242_U110 );
nand NAND2_19878 ( P3_ADD_360_1242_U208 , P3_ADD_360_1242_U142 , P3_ADD_360_1242_U206 );
nand NAND2_19879 ( P3_ADD_360_1242_U209 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_360_1242_U33 );
nand NAND2_19880 ( P3_ADD_360_1242_U210 , P3_ADD_360_U17 , P3_ADD_360_1242_U34 );
nand NAND2_19881 ( P3_ADD_360_1242_U211 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_360_1242_U33 );
nand NAND2_19882 ( P3_ADD_360_1242_U212 , P3_ADD_360_U17 , P3_ADD_360_1242_U34 );
nand NAND2_19883 ( P3_ADD_360_1242_U213 , P3_ADD_360_1242_U212 , P3_ADD_360_1242_U211 );
nand NAND2_19884 ( P3_ADD_360_1242_U214 , P3_ADD_360_1242_U111 , P3_ADD_360_1242_U112 );
nand NAND2_19885 ( P3_ADD_360_1242_U215 , P3_ADD_360_1242_U138 , P3_ADD_360_1242_U213 );
nand NAND2_19886 ( P3_ADD_360_1242_U216 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_360_1242_U32 );
nand NAND2_19887 ( P3_ADD_360_1242_U217 , P3_ADD_360_U18 , P3_ADD_360_1242_U31 );
nand NAND2_19888 ( P3_ADD_360_1242_U218 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_360_1242_U32 );
nand NAND2_19889 ( P3_ADD_360_1242_U219 , P3_ADD_360_U18 , P3_ADD_360_1242_U31 );
nand NAND2_19890 ( P3_ADD_360_1242_U220 , P3_ADD_360_1242_U219 , P3_ADD_360_1242_U218 );
nand NAND2_19891 ( P3_ADD_360_1242_U221 , P3_ADD_360_1242_U113 , P3_ADD_360_1242_U114 );
nand NAND2_19892 ( P3_ADD_360_1242_U222 , P3_ADD_360_1242_U136 , P3_ADD_360_1242_U220 );
nand NAND2_19893 ( P3_ADD_360_1242_U223 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_360_1242_U20 );
nand NAND2_19894 ( P3_ADD_360_1242_U224 , P3_ADD_360_U19 , P3_ADD_360_1242_U21 );
nand NAND2_19895 ( P3_ADD_360_1242_U225 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_360_1242_U22 );
nand NAND2_19896 ( P3_ADD_360_1242_U226 , P3_ADD_360_U20 , P3_ADD_360_1242_U23 );
nand NAND2_19897 ( P3_ADD_360_1242_U227 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_360_1242_U187 );
nand NAND3_19898 ( P3_ADD_360_1242_U228 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_360_1242_U165 , P3_ADD_360_1242_U116 );
nand NAND2_19899 ( P3_ADD_360_1242_U229 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_360_1242_U73 );
nand NAND2_19900 ( P3_ADD_360_1242_U230 , P3_ADD_360_1242_U165 , P3_ADD_360_1242_U74 );
nand NAND2_19901 ( P3_ADD_360_1242_U231 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_360_1242_U29 );
nand NAND2_19902 ( P3_ADD_360_1242_U232 , P3_ADD_360_U21 , P3_ADD_360_1242_U30 );
nand NAND2_19903 ( P3_ADD_360_1242_U233 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_360_1242_U29 );
nand NAND2_19904 ( P3_ADD_360_1242_U234 , P3_ADD_360_U21 , P3_ADD_360_1242_U30 );
nand NAND2_19905 ( P3_ADD_360_1242_U235 , P3_ADD_360_1242_U234 , P3_ADD_360_1242_U233 );
nand NAND2_19906 ( P3_ADD_360_1242_U236 , P3_ADD_360_1242_U117 , P3_ADD_360_1242_U118 );
nand NAND2_19907 ( P3_ADD_360_1242_U237 , P3_ADD_360_1242_U128 , P3_ADD_360_1242_U235 );
nand NAND2_19908 ( P3_ADD_360_1242_U238 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_360_1242_U68 );
nand NAND2_19909 ( P3_ADD_360_1242_U239 , P3_ADD_360_1242_U163 , P3_ADD_360_1242_U70 );
nand NAND2_19910 ( P3_ADD_360_1242_U240 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_360_1242_U63 );
nand NAND2_19911 ( P3_ADD_360_1242_U241 , P3_ADD_360_1242_U161 , P3_ADD_360_1242_U65 );
nand NAND2_19912 ( P3_ADD_360_1242_U242 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_360_1242_U60 );
nand NAND2_19913 ( P3_ADD_360_1242_U243 , P3_ADD_360_1242_U160 , P3_ADD_360_1242_U62 );
nand NAND2_19914 ( P3_ADD_360_1242_U244 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_360_1242_U27 );
nand NAND2_19915 ( P3_ADD_360_1242_U245 , P3_ADD_360_1242_U124 , P3_ADD_360_1242_U26 );
nand NAND2_19916 ( P3_ADD_360_1242_U246 , P3_ADD_360_1242_U245 , P3_ADD_360_1242_U244 );
nand NAND3_19917 ( P3_ADD_360_1242_U247 , P3_ADD_360_1242_U27 , P3_ADD_360_1242_U26 , P3_ADD_360_U4 );
nand NAND2_19918 ( P3_ADD_360_1242_U248 , P3_ADD_360_1242_U246 , P3_ADD_360_1242_U28 );
nand NAND2_19919 ( P3_ADD_360_1242_U249 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_360_1242_U53 );
nand NAND2_19920 ( P3_ADD_360_1242_U250 , P3_ADD_360_1242_U157 , P3_ADD_360_1242_U54 );
nand NAND2_19921 ( P3_ADD_360_1242_U251 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_360_1242_U50 );
nand NAND2_19922 ( P3_ADD_360_1242_U252 , P3_ADD_360_1242_U156 , P3_ADD_360_1242_U52 );
nand NAND2_19923 ( P3_ADD_360_1242_U253 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_360_1242_U76 );
nand NAND2_19924 ( P3_ADD_360_1242_U254 , P3_ADD_360_1242_U155 , P3_ADD_360_1242_U49 );
nand NAND2_19925 ( P3_ADD_360_1242_U255 , P3_ADD_360_1242_U119 , P3_ADD_360_1242_U43 );
nand NAND2_19926 ( P3_ADD_360_1242_U256 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_360_1242_U45 );
nand NAND2_19927 ( P3_ADD_360_1242_U257 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_360_1242_U24 );
nand NAND2_19928 ( P3_ADD_360_1242_U258 , P3_U2621 , P3_ADD_360_1242_U25 );
or OR2_19929 ( P3_LT_563_1260_U6 , P3_LT_563_1260_U7 , P3_U3304 );
nor nor_19930 ( P3_LT_563_1260_U7 , P3_SUB_563_U7 , P3_SUB_563_U6 );
not NOT1_19931 ( P3_SUB_589_U6 , P3_U3301 );
not NOT1_19932 ( P3_SUB_589_U7 , P3_U3302 );
not NOT1_19933 ( P3_SUB_589_U8 , P3_U2632 );
not NOT1_19934 ( P3_SUB_589_U9 , P3_U3300 );
not NOT1_19935 ( P3_ADD_467_U4 , P3_REIP_REG_1_ );
not NOT1_19936 ( P3_ADD_467_U5 , P3_REIP_REG_2_ );
nand NAND2_19937 ( P3_ADD_467_U6 , P3_REIP_REG_2_ , P3_REIP_REG_1_ );
not NOT1_19938 ( P3_ADD_467_U7 , P3_REIP_REG_3_ );
nand NAND2_19939 ( P3_ADD_467_U8 , P3_REIP_REG_3_ , P3_ADD_467_U94 );
not NOT1_19940 ( P3_ADD_467_U9 , P3_REIP_REG_4_ );
nand NAND2_19941 ( P3_ADD_467_U10 , P3_REIP_REG_4_ , P3_ADD_467_U95 );
not NOT1_19942 ( P3_ADD_467_U11 , P3_REIP_REG_5_ );
nand NAND2_19943 ( P3_ADD_467_U12 , P3_REIP_REG_5_ , P3_ADD_467_U96 );
not NOT1_19944 ( P3_ADD_467_U13 , P3_REIP_REG_6_ );
nand NAND2_19945 ( P3_ADD_467_U14 , P3_REIP_REG_6_ , P3_ADD_467_U97 );
not NOT1_19946 ( P3_ADD_467_U15 , P3_REIP_REG_7_ );
nand NAND2_19947 ( P3_ADD_467_U16 , P3_REIP_REG_7_ , P3_ADD_467_U98 );
not NOT1_19948 ( P3_ADD_467_U17 , P3_REIP_REG_8_ );
not NOT1_19949 ( P3_ADD_467_U18 , P3_REIP_REG_9_ );
nand NAND2_19950 ( P3_ADD_467_U19 , P3_REIP_REG_8_ , P3_ADD_467_U99 );
nand NAND2_19951 ( P3_ADD_467_U20 , P3_ADD_467_U100 , P3_REIP_REG_9_ );
not NOT1_19952 ( P3_ADD_467_U21 , P3_REIP_REG_10_ );
nand NAND2_19953 ( P3_ADD_467_U22 , P3_REIP_REG_10_ , P3_ADD_467_U101 );
not NOT1_19954 ( P3_ADD_467_U23 , P3_REIP_REG_11_ );
nand NAND2_19955 ( P3_ADD_467_U24 , P3_REIP_REG_11_ , P3_ADD_467_U102 );
not NOT1_19956 ( P3_ADD_467_U25 , P3_REIP_REG_12_ );
nand NAND2_19957 ( P3_ADD_467_U26 , P3_REIP_REG_12_ , P3_ADD_467_U103 );
not NOT1_19958 ( P3_ADD_467_U27 , P3_REIP_REG_13_ );
nand NAND2_19959 ( P3_ADD_467_U28 , P3_REIP_REG_13_ , P3_ADD_467_U104 );
not NOT1_19960 ( P3_ADD_467_U29 , P3_REIP_REG_14_ );
nand NAND2_19961 ( P3_ADD_467_U30 , P3_REIP_REG_14_ , P3_ADD_467_U105 );
not NOT1_19962 ( P3_ADD_467_U31 , P3_REIP_REG_15_ );
nand NAND2_19963 ( P3_ADD_467_U32 , P3_REIP_REG_15_ , P3_ADD_467_U106 );
not NOT1_19964 ( P3_ADD_467_U33 , P3_REIP_REG_16_ );
nand NAND2_19965 ( P3_ADD_467_U34 , P3_REIP_REG_16_ , P3_ADD_467_U107 );
not NOT1_19966 ( P3_ADD_467_U35 , P3_REIP_REG_17_ );
nand NAND2_19967 ( P3_ADD_467_U36 , P3_REIP_REG_17_ , P3_ADD_467_U108 );
not NOT1_19968 ( P3_ADD_467_U37 , P3_REIP_REG_18_ );
nand NAND2_19969 ( P3_ADD_467_U38 , P3_REIP_REG_18_ , P3_ADD_467_U109 );
not NOT1_19970 ( P3_ADD_467_U39 , P3_REIP_REG_19_ );
nand NAND2_19971 ( P3_ADD_467_U40 , P3_REIP_REG_19_ , P3_ADD_467_U110 );
not NOT1_19972 ( P3_ADD_467_U41 , P3_REIP_REG_20_ );
nand NAND2_19973 ( P3_ADD_467_U42 , P3_REIP_REG_20_ , P3_ADD_467_U111 );
not NOT1_19974 ( P3_ADD_467_U43 , P3_REIP_REG_21_ );
nand NAND2_19975 ( P3_ADD_467_U44 , P3_REIP_REG_21_ , P3_ADD_467_U112 );
not NOT1_19976 ( P3_ADD_467_U45 , P3_REIP_REG_22_ );
nand NAND2_19977 ( P3_ADD_467_U46 , P3_REIP_REG_22_ , P3_ADD_467_U113 );
not NOT1_19978 ( P3_ADD_467_U47 , P3_REIP_REG_23_ );
nand NAND2_19979 ( P3_ADD_467_U48 , P3_REIP_REG_23_ , P3_ADD_467_U114 );
not NOT1_19980 ( P3_ADD_467_U49 , P3_REIP_REG_24_ );
nand NAND2_19981 ( P3_ADD_467_U50 , P3_REIP_REG_24_ , P3_ADD_467_U115 );
not NOT1_19982 ( P3_ADD_467_U51 , P3_REIP_REG_25_ );
nand NAND2_19983 ( P3_ADD_467_U52 , P3_REIP_REG_25_ , P3_ADD_467_U116 );
not NOT1_19984 ( P3_ADD_467_U53 , P3_REIP_REG_26_ );
nand NAND2_19985 ( P3_ADD_467_U54 , P3_REIP_REG_26_ , P3_ADD_467_U117 );
not NOT1_19986 ( P3_ADD_467_U55 , P3_REIP_REG_27_ );
nand NAND2_19987 ( P3_ADD_467_U56 , P3_REIP_REG_27_ , P3_ADD_467_U118 );
not NOT1_19988 ( P3_ADD_467_U57 , P3_REIP_REG_28_ );
nand NAND2_19989 ( P3_ADD_467_U58 , P3_REIP_REG_28_ , P3_ADD_467_U119 );
not NOT1_19990 ( P3_ADD_467_U59 , P3_REIP_REG_29_ );
nand NAND2_19991 ( P3_ADD_467_U60 , P3_REIP_REG_29_ , P3_ADD_467_U120 );
not NOT1_19992 ( P3_ADD_467_U61 , P3_REIP_REG_30_ );
nand NAND2_19993 ( P3_ADD_467_U62 , P3_ADD_467_U124 , P3_ADD_467_U123 );
nand NAND2_19994 ( P3_ADD_467_U63 , P3_ADD_467_U126 , P3_ADD_467_U125 );
nand NAND2_19995 ( P3_ADD_467_U64 , P3_ADD_467_U128 , P3_ADD_467_U127 );
nand NAND2_19996 ( P3_ADD_467_U65 , P3_ADD_467_U130 , P3_ADD_467_U129 );
nand NAND2_19997 ( P3_ADD_467_U66 , P3_ADD_467_U132 , P3_ADD_467_U131 );
nand NAND2_19998 ( P3_ADD_467_U67 , P3_ADD_467_U134 , P3_ADD_467_U133 );
nand NAND2_19999 ( P3_ADD_467_U68 , P3_ADD_467_U136 , P3_ADD_467_U135 );
nand NAND2_20000 ( P3_ADD_467_U69 , P3_ADD_467_U138 , P3_ADD_467_U137 );
nand NAND2_20001 ( P3_ADD_467_U70 , P3_ADD_467_U140 , P3_ADD_467_U139 );
nand NAND2_20002 ( P3_ADD_467_U71 , P3_ADD_467_U142 , P3_ADD_467_U141 );
nand NAND2_20003 ( P3_ADD_467_U72 , P3_ADD_467_U144 , P3_ADD_467_U143 );
nand NAND2_20004 ( P3_ADD_467_U73 , P3_ADD_467_U146 , P3_ADD_467_U145 );
nand NAND2_20005 ( P3_ADD_467_U74 , P3_ADD_467_U148 , P3_ADD_467_U147 );
nand NAND2_20006 ( P3_ADD_467_U75 , P3_ADD_467_U150 , P3_ADD_467_U149 );
nand NAND2_20007 ( P3_ADD_467_U76 , P3_ADD_467_U152 , P3_ADD_467_U151 );
nand NAND2_20008 ( P3_ADD_467_U77 , P3_ADD_467_U154 , P3_ADD_467_U153 );
nand NAND2_20009 ( P3_ADD_467_U78 , P3_ADD_467_U156 , P3_ADD_467_U155 );
nand NAND2_20010 ( P3_ADD_467_U79 , P3_ADD_467_U158 , P3_ADD_467_U157 );
nand NAND2_20011 ( P3_ADD_467_U80 , P3_ADD_467_U160 , P3_ADD_467_U159 );
nand NAND2_20012 ( P3_ADD_467_U81 , P3_ADD_467_U162 , P3_ADD_467_U161 );
nand NAND2_20013 ( P3_ADD_467_U82 , P3_ADD_467_U164 , P3_ADD_467_U163 );
nand NAND2_20014 ( P3_ADD_467_U83 , P3_ADD_467_U166 , P3_ADD_467_U165 );
nand NAND2_20015 ( P3_ADD_467_U84 , P3_ADD_467_U168 , P3_ADD_467_U167 );
nand NAND2_20016 ( P3_ADD_467_U85 , P3_ADD_467_U170 , P3_ADD_467_U169 );
nand NAND2_20017 ( P3_ADD_467_U86 , P3_ADD_467_U172 , P3_ADD_467_U171 );
nand NAND2_20018 ( P3_ADD_467_U87 , P3_ADD_467_U174 , P3_ADD_467_U173 );
nand NAND2_20019 ( P3_ADD_467_U88 , P3_ADD_467_U176 , P3_ADD_467_U175 );
nand NAND2_20020 ( P3_ADD_467_U89 , P3_ADD_467_U178 , P3_ADD_467_U177 );
nand NAND2_20021 ( P3_ADD_467_U90 , P3_ADD_467_U180 , P3_ADD_467_U179 );
nand NAND2_20022 ( P3_ADD_467_U91 , P3_ADD_467_U182 , P3_ADD_467_U181 );
not NOT1_20023 ( P3_ADD_467_U92 , P3_REIP_REG_31_ );
nand NAND2_20024 ( P3_ADD_467_U93 , P3_REIP_REG_30_ , P3_ADD_467_U121 );
not NOT1_20025 ( P3_ADD_467_U94 , P3_ADD_467_U6 );
not NOT1_20026 ( P3_ADD_467_U95 , P3_ADD_467_U8 );
not NOT1_20027 ( P3_ADD_467_U96 , P3_ADD_467_U10 );
not NOT1_20028 ( P3_ADD_467_U97 , P3_ADD_467_U12 );
not NOT1_20029 ( P3_ADD_467_U98 , P3_ADD_467_U14 );
not NOT1_20030 ( P3_ADD_467_U99 , P3_ADD_467_U16 );
not NOT1_20031 ( P3_ADD_467_U100 , P3_ADD_467_U19 );
not NOT1_20032 ( P3_ADD_467_U101 , P3_ADD_467_U20 );
not NOT1_20033 ( P3_ADD_467_U102 , P3_ADD_467_U22 );
not NOT1_20034 ( P3_ADD_467_U103 , P3_ADD_467_U24 );
not NOT1_20035 ( P3_ADD_467_U104 , P3_ADD_467_U26 );
not NOT1_20036 ( P3_ADD_467_U105 , P3_ADD_467_U28 );
not NOT1_20037 ( P3_ADD_467_U106 , P3_ADD_467_U30 );
not NOT1_20038 ( P3_ADD_467_U107 , P3_ADD_467_U32 );
not NOT1_20039 ( P3_ADD_467_U108 , P3_ADD_467_U34 );
not NOT1_20040 ( P3_ADD_467_U109 , P3_ADD_467_U36 );
not NOT1_20041 ( P3_ADD_467_U110 , P3_ADD_467_U38 );
not NOT1_20042 ( P3_ADD_467_U111 , P3_ADD_467_U40 );
not NOT1_20043 ( P3_ADD_467_U112 , P3_ADD_467_U42 );
not NOT1_20044 ( P3_ADD_467_U113 , P3_ADD_467_U44 );
not NOT1_20045 ( P3_ADD_467_U114 , P3_ADD_467_U46 );
not NOT1_20046 ( P3_ADD_467_U115 , P3_ADD_467_U48 );
not NOT1_20047 ( P3_ADD_467_U116 , P3_ADD_467_U50 );
not NOT1_20048 ( P3_ADD_467_U117 , P3_ADD_467_U52 );
not NOT1_20049 ( P3_ADD_467_U118 , P3_ADD_467_U54 );
not NOT1_20050 ( P3_ADD_467_U119 , P3_ADD_467_U56 );
not NOT1_20051 ( P3_ADD_467_U120 , P3_ADD_467_U58 );
not NOT1_20052 ( P3_ADD_467_U121 , P3_ADD_467_U60 );
not NOT1_20053 ( P3_ADD_467_U122 , P3_ADD_467_U93 );
nand NAND2_20054 ( P3_ADD_467_U123 , P3_REIP_REG_9_ , P3_ADD_467_U19 );
nand NAND2_20055 ( P3_ADD_467_U124 , P3_ADD_467_U100 , P3_ADD_467_U18 );
nand NAND2_20056 ( P3_ADD_467_U125 , P3_REIP_REG_8_ , P3_ADD_467_U16 );
nand NAND2_20057 ( P3_ADD_467_U126 , P3_ADD_467_U99 , P3_ADD_467_U17 );
nand NAND2_20058 ( P3_ADD_467_U127 , P3_REIP_REG_7_ , P3_ADD_467_U14 );
nand NAND2_20059 ( P3_ADD_467_U128 , P3_ADD_467_U98 , P3_ADD_467_U15 );
nand NAND2_20060 ( P3_ADD_467_U129 , P3_REIP_REG_6_ , P3_ADD_467_U12 );
nand NAND2_20061 ( P3_ADD_467_U130 , P3_ADD_467_U97 , P3_ADD_467_U13 );
nand NAND2_20062 ( P3_ADD_467_U131 , P3_REIP_REG_5_ , P3_ADD_467_U10 );
nand NAND2_20063 ( P3_ADD_467_U132 , P3_ADD_467_U96 , P3_ADD_467_U11 );
nand NAND2_20064 ( P3_ADD_467_U133 , P3_REIP_REG_4_ , P3_ADD_467_U8 );
nand NAND2_20065 ( P3_ADD_467_U134 , P3_ADD_467_U95 , P3_ADD_467_U9 );
nand NAND2_20066 ( P3_ADD_467_U135 , P3_REIP_REG_3_ , P3_ADD_467_U6 );
nand NAND2_20067 ( P3_ADD_467_U136 , P3_ADD_467_U94 , P3_ADD_467_U7 );
nand NAND2_20068 ( P3_ADD_467_U137 , P3_REIP_REG_31_ , P3_ADD_467_U93 );
nand NAND2_20069 ( P3_ADD_467_U138 , P3_ADD_467_U122 , P3_ADD_467_U92 );
nand NAND2_20070 ( P3_ADD_467_U139 , P3_REIP_REG_30_ , P3_ADD_467_U60 );
nand NAND2_20071 ( P3_ADD_467_U140 , P3_ADD_467_U121 , P3_ADD_467_U61 );
nand NAND2_20072 ( P3_ADD_467_U141 , P3_REIP_REG_2_ , P3_ADD_467_U4 );
nand NAND2_20073 ( P3_ADD_467_U142 , P3_REIP_REG_1_ , P3_ADD_467_U5 );
nand NAND2_20074 ( P3_ADD_467_U143 , P3_REIP_REG_29_ , P3_ADD_467_U58 );
nand NAND2_20075 ( P3_ADD_467_U144 , P3_ADD_467_U120 , P3_ADD_467_U59 );
nand NAND2_20076 ( P3_ADD_467_U145 , P3_REIP_REG_28_ , P3_ADD_467_U56 );
nand NAND2_20077 ( P3_ADD_467_U146 , P3_ADD_467_U119 , P3_ADD_467_U57 );
nand NAND2_20078 ( P3_ADD_467_U147 , P3_REIP_REG_27_ , P3_ADD_467_U54 );
nand NAND2_20079 ( P3_ADD_467_U148 , P3_ADD_467_U118 , P3_ADD_467_U55 );
nand NAND2_20080 ( P3_ADD_467_U149 , P3_REIP_REG_26_ , P3_ADD_467_U52 );
nand NAND2_20081 ( P3_ADD_467_U150 , P3_ADD_467_U117 , P3_ADD_467_U53 );
nand NAND2_20082 ( P3_ADD_467_U151 , P3_REIP_REG_25_ , P3_ADD_467_U50 );
nand NAND2_20083 ( P3_ADD_467_U152 , P3_ADD_467_U116 , P3_ADD_467_U51 );
nand NAND2_20084 ( P3_ADD_467_U153 , P3_REIP_REG_24_ , P3_ADD_467_U48 );
nand NAND2_20085 ( P3_ADD_467_U154 , P3_ADD_467_U115 , P3_ADD_467_U49 );
nand NAND2_20086 ( P3_ADD_467_U155 , P3_REIP_REG_23_ , P3_ADD_467_U46 );
nand NAND2_20087 ( P3_ADD_467_U156 , P3_ADD_467_U114 , P3_ADD_467_U47 );
nand NAND2_20088 ( P3_ADD_467_U157 , P3_REIP_REG_22_ , P3_ADD_467_U44 );
nand NAND2_20089 ( P3_ADD_467_U158 , P3_ADD_467_U113 , P3_ADD_467_U45 );
nand NAND2_20090 ( P3_ADD_467_U159 , P3_REIP_REG_21_ , P3_ADD_467_U42 );
nand NAND2_20091 ( P3_ADD_467_U160 , P3_ADD_467_U112 , P3_ADD_467_U43 );
nand NAND2_20092 ( P3_ADD_467_U161 , P3_REIP_REG_20_ , P3_ADD_467_U40 );
nand NAND2_20093 ( P3_ADD_467_U162 , P3_ADD_467_U111 , P3_ADD_467_U41 );
nand NAND2_20094 ( P3_ADD_467_U163 , P3_REIP_REG_19_ , P3_ADD_467_U38 );
nand NAND2_20095 ( P3_ADD_467_U164 , P3_ADD_467_U110 , P3_ADD_467_U39 );
nand NAND2_20096 ( P3_ADD_467_U165 , P3_REIP_REG_18_ , P3_ADD_467_U36 );
nand NAND2_20097 ( P3_ADD_467_U166 , P3_ADD_467_U109 , P3_ADD_467_U37 );
nand NAND2_20098 ( P3_ADD_467_U167 , P3_REIP_REG_17_ , P3_ADD_467_U34 );
nand NAND2_20099 ( P3_ADD_467_U168 , P3_ADD_467_U108 , P3_ADD_467_U35 );
nand NAND2_20100 ( P3_ADD_467_U169 , P3_REIP_REG_16_ , P3_ADD_467_U32 );
nand NAND2_20101 ( P3_ADD_467_U170 , P3_ADD_467_U107 , P3_ADD_467_U33 );
nand NAND2_20102 ( P3_ADD_467_U171 , P3_REIP_REG_15_ , P3_ADD_467_U30 );
nand NAND2_20103 ( P3_ADD_467_U172 , P3_ADD_467_U106 , P3_ADD_467_U31 );
nand NAND2_20104 ( P3_ADD_467_U173 , P3_REIP_REG_14_ , P3_ADD_467_U28 );
nand NAND2_20105 ( P3_ADD_467_U174 , P3_ADD_467_U105 , P3_ADD_467_U29 );
nand NAND2_20106 ( P3_ADD_467_U175 , P3_REIP_REG_13_ , P3_ADD_467_U26 );
nand NAND2_20107 ( P3_ADD_467_U176 , P3_ADD_467_U104 , P3_ADD_467_U27 );
nand NAND2_20108 ( P3_ADD_467_U177 , P3_REIP_REG_12_ , P3_ADD_467_U24 );
nand NAND2_20109 ( P3_ADD_467_U178 , P3_ADD_467_U103 , P3_ADD_467_U25 );
nand NAND2_20110 ( P3_ADD_467_U179 , P3_REIP_REG_11_ , P3_ADD_467_U22 );
nand NAND2_20111 ( P3_ADD_467_U180 , P3_ADD_467_U102 , P3_ADD_467_U23 );
nand NAND2_20112 ( P3_ADD_467_U181 , P3_REIP_REG_10_ , P3_ADD_467_U20 );
nand NAND2_20113 ( P3_ADD_467_U182 , P3_ADD_467_U101 , P3_ADD_467_U21 );
not NOT1_20114 ( P3_ADD_430_U4 , P3_REIP_REG_1_ );
not NOT1_20115 ( P3_ADD_430_U5 , P3_REIP_REG_2_ );
nand NAND2_20116 ( P3_ADD_430_U6 , P3_REIP_REG_2_ , P3_REIP_REG_1_ );
not NOT1_20117 ( P3_ADD_430_U7 , P3_REIP_REG_3_ );
nand NAND2_20118 ( P3_ADD_430_U8 , P3_REIP_REG_3_ , P3_ADD_430_U94 );
not NOT1_20119 ( P3_ADD_430_U9 , P3_REIP_REG_4_ );
nand NAND2_20120 ( P3_ADD_430_U10 , P3_REIP_REG_4_ , P3_ADD_430_U95 );
not NOT1_20121 ( P3_ADD_430_U11 , P3_REIP_REG_5_ );
nand NAND2_20122 ( P3_ADD_430_U12 , P3_REIP_REG_5_ , P3_ADD_430_U96 );
not NOT1_20123 ( P3_ADD_430_U13 , P3_REIP_REG_6_ );
nand NAND2_20124 ( P3_ADD_430_U14 , P3_REIP_REG_6_ , P3_ADD_430_U97 );
not NOT1_20125 ( P3_ADD_430_U15 , P3_REIP_REG_7_ );
nand NAND2_20126 ( P3_ADD_430_U16 , P3_REIP_REG_7_ , P3_ADD_430_U98 );
not NOT1_20127 ( P3_ADD_430_U17 , P3_REIP_REG_8_ );
not NOT1_20128 ( P3_ADD_430_U18 , P3_REIP_REG_9_ );
nand NAND2_20129 ( P3_ADD_430_U19 , P3_REIP_REG_8_ , P3_ADD_430_U99 );
nand NAND2_20130 ( P3_ADD_430_U20 , P3_ADD_430_U100 , P3_REIP_REG_9_ );
not NOT1_20131 ( P3_ADD_430_U21 , P3_REIP_REG_10_ );
nand NAND2_20132 ( P3_ADD_430_U22 , P3_REIP_REG_10_ , P3_ADD_430_U101 );
not NOT1_20133 ( P3_ADD_430_U23 , P3_REIP_REG_11_ );
nand NAND2_20134 ( P3_ADD_430_U24 , P3_REIP_REG_11_ , P3_ADD_430_U102 );
not NOT1_20135 ( P3_ADD_430_U25 , P3_REIP_REG_12_ );
nand NAND2_20136 ( P3_ADD_430_U26 , P3_REIP_REG_12_ , P3_ADD_430_U103 );
not NOT1_20137 ( P3_ADD_430_U27 , P3_REIP_REG_13_ );
nand NAND2_20138 ( P3_ADD_430_U28 , P3_REIP_REG_13_ , P3_ADD_430_U104 );
not NOT1_20139 ( P3_ADD_430_U29 , P3_REIP_REG_14_ );
nand NAND2_20140 ( P3_ADD_430_U30 , P3_REIP_REG_14_ , P3_ADD_430_U105 );
not NOT1_20141 ( P3_ADD_430_U31 , P3_REIP_REG_15_ );
nand NAND2_20142 ( P3_ADD_430_U32 , P3_REIP_REG_15_ , P3_ADD_430_U106 );
not NOT1_20143 ( P3_ADD_430_U33 , P3_REIP_REG_16_ );
nand NAND2_20144 ( P3_ADD_430_U34 , P3_REIP_REG_16_ , P3_ADD_430_U107 );
not NOT1_20145 ( P3_ADD_430_U35 , P3_REIP_REG_17_ );
nand NAND2_20146 ( P3_ADD_430_U36 , P3_REIP_REG_17_ , P3_ADD_430_U108 );
not NOT1_20147 ( P3_ADD_430_U37 , P3_REIP_REG_18_ );
nand NAND2_20148 ( P3_ADD_430_U38 , P3_REIP_REG_18_ , P3_ADD_430_U109 );
not NOT1_20149 ( P3_ADD_430_U39 , P3_REIP_REG_19_ );
nand NAND2_20150 ( P3_ADD_430_U40 , P3_REIP_REG_19_ , P3_ADD_430_U110 );
not NOT1_20151 ( P3_ADD_430_U41 , P3_REIP_REG_20_ );
nand NAND2_20152 ( P3_ADD_430_U42 , P3_REIP_REG_20_ , P3_ADD_430_U111 );
not NOT1_20153 ( P3_ADD_430_U43 , P3_REIP_REG_21_ );
nand NAND2_20154 ( P3_ADD_430_U44 , P3_REIP_REG_21_ , P3_ADD_430_U112 );
not NOT1_20155 ( P3_ADD_430_U45 , P3_REIP_REG_22_ );
nand NAND2_20156 ( P3_ADD_430_U46 , P3_REIP_REG_22_ , P3_ADD_430_U113 );
not NOT1_20157 ( P3_ADD_430_U47 , P3_REIP_REG_23_ );
nand NAND2_20158 ( P3_ADD_430_U48 , P3_REIP_REG_23_ , P3_ADD_430_U114 );
not NOT1_20159 ( P3_ADD_430_U49 , P3_REIP_REG_24_ );
nand NAND2_20160 ( P3_ADD_430_U50 , P3_REIP_REG_24_ , P3_ADD_430_U115 );
not NOT1_20161 ( P3_ADD_430_U51 , P3_REIP_REG_25_ );
nand NAND2_20162 ( P3_ADD_430_U52 , P3_REIP_REG_25_ , P3_ADD_430_U116 );
not NOT1_20163 ( P3_ADD_430_U53 , P3_REIP_REG_26_ );
nand NAND2_20164 ( P3_ADD_430_U54 , P3_REIP_REG_26_ , P3_ADD_430_U117 );
not NOT1_20165 ( P3_ADD_430_U55 , P3_REIP_REG_27_ );
nand NAND2_20166 ( P3_ADD_430_U56 , P3_REIP_REG_27_ , P3_ADD_430_U118 );
not NOT1_20167 ( P3_ADD_430_U57 , P3_REIP_REG_28_ );
nand NAND2_20168 ( P3_ADD_430_U58 , P3_REIP_REG_28_ , P3_ADD_430_U119 );
not NOT1_20169 ( P3_ADD_430_U59 , P3_REIP_REG_29_ );
nand NAND2_20170 ( P3_ADD_430_U60 , P3_REIP_REG_29_ , P3_ADD_430_U120 );
not NOT1_20171 ( P3_ADD_430_U61 , P3_REIP_REG_30_ );
nand NAND2_20172 ( P3_ADD_430_U62 , P3_ADD_430_U124 , P3_ADD_430_U123 );
nand NAND2_20173 ( P3_ADD_430_U63 , P3_ADD_430_U126 , P3_ADD_430_U125 );
nand NAND2_20174 ( P3_ADD_430_U64 , P3_ADD_430_U128 , P3_ADD_430_U127 );
nand NAND2_20175 ( P3_ADD_430_U65 , P3_ADD_430_U130 , P3_ADD_430_U129 );
nand NAND2_20176 ( P3_ADD_430_U66 , P3_ADD_430_U132 , P3_ADD_430_U131 );
nand NAND2_20177 ( P3_ADD_430_U67 , P3_ADD_430_U134 , P3_ADD_430_U133 );
nand NAND2_20178 ( P3_ADD_430_U68 , P3_ADD_430_U136 , P3_ADD_430_U135 );
nand NAND2_20179 ( P3_ADD_430_U69 , P3_ADD_430_U138 , P3_ADD_430_U137 );
nand NAND2_20180 ( P3_ADD_430_U70 , P3_ADD_430_U140 , P3_ADD_430_U139 );
nand NAND2_20181 ( P3_ADD_430_U71 , P3_ADD_430_U142 , P3_ADD_430_U141 );
nand NAND2_20182 ( P3_ADD_430_U72 , P3_ADD_430_U144 , P3_ADD_430_U143 );
nand NAND2_20183 ( P3_ADD_430_U73 , P3_ADD_430_U146 , P3_ADD_430_U145 );
nand NAND2_20184 ( P3_ADD_430_U74 , P3_ADD_430_U148 , P3_ADD_430_U147 );
nand NAND2_20185 ( P3_ADD_430_U75 , P3_ADD_430_U150 , P3_ADD_430_U149 );
nand NAND2_20186 ( P3_ADD_430_U76 , P3_ADD_430_U152 , P3_ADD_430_U151 );
nand NAND2_20187 ( P3_ADD_430_U77 , P3_ADD_430_U154 , P3_ADD_430_U153 );
nand NAND2_20188 ( P3_ADD_430_U78 , P3_ADD_430_U156 , P3_ADD_430_U155 );
nand NAND2_20189 ( P3_ADD_430_U79 , P3_ADD_430_U158 , P3_ADD_430_U157 );
nand NAND2_20190 ( P3_ADD_430_U80 , P3_ADD_430_U160 , P3_ADD_430_U159 );
nand NAND2_20191 ( P3_ADD_430_U81 , P3_ADD_430_U162 , P3_ADD_430_U161 );
nand NAND2_20192 ( P3_ADD_430_U82 , P3_ADD_430_U164 , P3_ADD_430_U163 );
nand NAND2_20193 ( P3_ADD_430_U83 , P3_ADD_430_U166 , P3_ADD_430_U165 );
nand NAND2_20194 ( P3_ADD_430_U84 , P3_ADD_430_U168 , P3_ADD_430_U167 );
nand NAND2_20195 ( P3_ADD_430_U85 , P3_ADD_430_U170 , P3_ADD_430_U169 );
nand NAND2_20196 ( P3_ADD_430_U86 , P3_ADD_430_U172 , P3_ADD_430_U171 );
nand NAND2_20197 ( P3_ADD_430_U87 , P3_ADD_430_U174 , P3_ADD_430_U173 );
nand NAND2_20198 ( P3_ADD_430_U88 , P3_ADD_430_U176 , P3_ADD_430_U175 );
nand NAND2_20199 ( P3_ADD_430_U89 , P3_ADD_430_U178 , P3_ADD_430_U177 );
nand NAND2_20200 ( P3_ADD_430_U90 , P3_ADD_430_U180 , P3_ADD_430_U179 );
nand NAND2_20201 ( P3_ADD_430_U91 , P3_ADD_430_U182 , P3_ADD_430_U181 );
not NOT1_20202 ( P3_ADD_430_U92 , P3_REIP_REG_31_ );
nand NAND2_20203 ( P3_ADD_430_U93 , P3_REIP_REG_30_ , P3_ADD_430_U121 );
not NOT1_20204 ( P3_ADD_430_U94 , P3_ADD_430_U6 );
not NOT1_20205 ( P3_ADD_430_U95 , P3_ADD_430_U8 );
not NOT1_20206 ( P3_ADD_430_U96 , P3_ADD_430_U10 );
not NOT1_20207 ( P3_ADD_430_U97 , P3_ADD_430_U12 );
not NOT1_20208 ( P3_ADD_430_U98 , P3_ADD_430_U14 );
not NOT1_20209 ( P3_ADD_430_U99 , P3_ADD_430_U16 );
not NOT1_20210 ( P3_ADD_430_U100 , P3_ADD_430_U19 );
not NOT1_20211 ( P3_ADD_430_U101 , P3_ADD_430_U20 );
not NOT1_20212 ( P3_ADD_430_U102 , P3_ADD_430_U22 );
not NOT1_20213 ( P3_ADD_430_U103 , P3_ADD_430_U24 );
not NOT1_20214 ( P3_ADD_430_U104 , P3_ADD_430_U26 );
not NOT1_20215 ( P3_ADD_430_U105 , P3_ADD_430_U28 );
not NOT1_20216 ( P3_ADD_430_U106 , P3_ADD_430_U30 );
not NOT1_20217 ( P3_ADD_430_U107 , P3_ADD_430_U32 );
not NOT1_20218 ( P3_ADD_430_U108 , P3_ADD_430_U34 );
not NOT1_20219 ( P3_ADD_430_U109 , P3_ADD_430_U36 );
not NOT1_20220 ( P3_ADD_430_U110 , P3_ADD_430_U38 );
not NOT1_20221 ( P3_ADD_430_U111 , P3_ADD_430_U40 );
not NOT1_20222 ( P3_ADD_430_U112 , P3_ADD_430_U42 );
not NOT1_20223 ( P3_ADD_430_U113 , P3_ADD_430_U44 );
not NOT1_20224 ( P3_ADD_430_U114 , P3_ADD_430_U46 );
not NOT1_20225 ( P3_ADD_430_U115 , P3_ADD_430_U48 );
not NOT1_20226 ( P3_ADD_430_U116 , P3_ADD_430_U50 );
not NOT1_20227 ( P3_ADD_430_U117 , P3_ADD_430_U52 );
not NOT1_20228 ( P3_ADD_430_U118 , P3_ADD_430_U54 );
not NOT1_20229 ( P3_ADD_430_U119 , P3_ADD_430_U56 );
not NOT1_20230 ( P3_ADD_430_U120 , P3_ADD_430_U58 );
not NOT1_20231 ( P3_ADD_430_U121 , P3_ADD_430_U60 );
not NOT1_20232 ( P3_ADD_430_U122 , P3_ADD_430_U93 );
nand NAND2_20233 ( P3_ADD_430_U123 , P3_REIP_REG_9_ , P3_ADD_430_U19 );
nand NAND2_20234 ( P3_ADD_430_U124 , P3_ADD_430_U100 , P3_ADD_430_U18 );
nand NAND2_20235 ( P3_ADD_430_U125 , P3_REIP_REG_8_ , P3_ADD_430_U16 );
nand NAND2_20236 ( P3_ADD_430_U126 , P3_ADD_430_U99 , P3_ADD_430_U17 );
nand NAND2_20237 ( P3_ADD_430_U127 , P3_REIP_REG_7_ , P3_ADD_430_U14 );
nand NAND2_20238 ( P3_ADD_430_U128 , P3_ADD_430_U98 , P3_ADD_430_U15 );
nand NAND2_20239 ( P3_ADD_430_U129 , P3_REIP_REG_6_ , P3_ADD_430_U12 );
nand NAND2_20240 ( P3_ADD_430_U130 , P3_ADD_430_U97 , P3_ADD_430_U13 );
nand NAND2_20241 ( P3_ADD_430_U131 , P3_REIP_REG_5_ , P3_ADD_430_U10 );
nand NAND2_20242 ( P3_ADD_430_U132 , P3_ADD_430_U96 , P3_ADD_430_U11 );
nand NAND2_20243 ( P3_ADD_430_U133 , P3_REIP_REG_4_ , P3_ADD_430_U8 );
nand NAND2_20244 ( P3_ADD_430_U134 , P3_ADD_430_U95 , P3_ADD_430_U9 );
nand NAND2_20245 ( P3_ADD_430_U135 , P3_REIP_REG_3_ , P3_ADD_430_U6 );
nand NAND2_20246 ( P3_ADD_430_U136 , P3_ADD_430_U94 , P3_ADD_430_U7 );
nand NAND2_20247 ( P3_ADD_430_U137 , P3_REIP_REG_31_ , P3_ADD_430_U93 );
nand NAND2_20248 ( P3_ADD_430_U138 , P3_ADD_430_U122 , P3_ADD_430_U92 );
nand NAND2_20249 ( P3_ADD_430_U139 , P3_REIP_REG_30_ , P3_ADD_430_U60 );
nand NAND2_20250 ( P3_ADD_430_U140 , P3_ADD_430_U121 , P3_ADD_430_U61 );
nand NAND2_20251 ( P3_ADD_430_U141 , P3_REIP_REG_2_ , P3_ADD_430_U4 );
nand NAND2_20252 ( P3_ADD_430_U142 , P3_REIP_REG_1_ , P3_ADD_430_U5 );
nand NAND2_20253 ( P3_ADD_430_U143 , P3_REIP_REG_29_ , P3_ADD_430_U58 );
nand NAND2_20254 ( P3_ADD_430_U144 , P3_ADD_430_U120 , P3_ADD_430_U59 );
nand NAND2_20255 ( P3_ADD_430_U145 , P3_REIP_REG_28_ , P3_ADD_430_U56 );
nand NAND2_20256 ( P3_ADD_430_U146 , P3_ADD_430_U119 , P3_ADD_430_U57 );
nand NAND2_20257 ( P3_ADD_430_U147 , P3_REIP_REG_27_ , P3_ADD_430_U54 );
nand NAND2_20258 ( P3_ADD_430_U148 , P3_ADD_430_U118 , P3_ADD_430_U55 );
nand NAND2_20259 ( P3_ADD_430_U149 , P3_REIP_REG_26_ , P3_ADD_430_U52 );
nand NAND2_20260 ( P3_ADD_430_U150 , P3_ADD_430_U117 , P3_ADD_430_U53 );
nand NAND2_20261 ( P3_ADD_430_U151 , P3_REIP_REG_25_ , P3_ADD_430_U50 );
nand NAND2_20262 ( P3_ADD_430_U152 , P3_ADD_430_U116 , P3_ADD_430_U51 );
nand NAND2_20263 ( P3_ADD_430_U153 , P3_REIP_REG_24_ , P3_ADD_430_U48 );
nand NAND2_20264 ( P3_ADD_430_U154 , P3_ADD_430_U115 , P3_ADD_430_U49 );
nand NAND2_20265 ( P3_ADD_430_U155 , P3_REIP_REG_23_ , P3_ADD_430_U46 );
nand NAND2_20266 ( P3_ADD_430_U156 , P3_ADD_430_U114 , P3_ADD_430_U47 );
nand NAND2_20267 ( P3_ADD_430_U157 , P3_REIP_REG_22_ , P3_ADD_430_U44 );
nand NAND2_20268 ( P3_ADD_430_U158 , P3_ADD_430_U113 , P3_ADD_430_U45 );
nand NAND2_20269 ( P3_ADD_430_U159 , P3_REIP_REG_21_ , P3_ADD_430_U42 );
nand NAND2_20270 ( P3_ADD_430_U160 , P3_ADD_430_U112 , P3_ADD_430_U43 );
nand NAND2_20271 ( P3_ADD_430_U161 , P3_REIP_REG_20_ , P3_ADD_430_U40 );
nand NAND2_20272 ( P3_ADD_430_U162 , P3_ADD_430_U111 , P3_ADD_430_U41 );
nand NAND2_20273 ( P3_ADD_430_U163 , P3_REIP_REG_19_ , P3_ADD_430_U38 );
nand NAND2_20274 ( P3_ADD_430_U164 , P3_ADD_430_U110 , P3_ADD_430_U39 );
nand NAND2_20275 ( P3_ADD_430_U165 , P3_REIP_REG_18_ , P3_ADD_430_U36 );
nand NAND2_20276 ( P3_ADD_430_U166 , P3_ADD_430_U109 , P3_ADD_430_U37 );
nand NAND2_20277 ( P3_ADD_430_U167 , P3_REIP_REG_17_ , P3_ADD_430_U34 );
nand NAND2_20278 ( P3_ADD_430_U168 , P3_ADD_430_U108 , P3_ADD_430_U35 );
nand NAND2_20279 ( P3_ADD_430_U169 , P3_REIP_REG_16_ , P3_ADD_430_U32 );
nand NAND2_20280 ( P3_ADD_430_U170 , P3_ADD_430_U107 , P3_ADD_430_U33 );
nand NAND2_20281 ( P3_ADD_430_U171 , P3_REIP_REG_15_ , P3_ADD_430_U30 );
nand NAND2_20282 ( P3_ADD_430_U172 , P3_ADD_430_U106 , P3_ADD_430_U31 );
nand NAND2_20283 ( P3_ADD_430_U173 , P3_REIP_REG_14_ , P3_ADD_430_U28 );
nand NAND2_20284 ( P3_ADD_430_U174 , P3_ADD_430_U105 , P3_ADD_430_U29 );
nand NAND2_20285 ( P3_ADD_430_U175 , P3_REIP_REG_13_ , P3_ADD_430_U26 );
nand NAND2_20286 ( P3_ADD_430_U176 , P3_ADD_430_U104 , P3_ADD_430_U27 );
nand NAND2_20287 ( P3_ADD_430_U177 , P3_REIP_REG_12_ , P3_ADD_430_U24 );
nand NAND2_20288 ( P3_ADD_430_U178 , P3_ADD_430_U103 , P3_ADD_430_U25 );
nand NAND2_20289 ( P3_ADD_430_U179 , P3_REIP_REG_11_ , P3_ADD_430_U22 );
nand NAND2_20290 ( P3_ADD_430_U180 , P3_ADD_430_U102 , P3_ADD_430_U23 );
nand NAND2_20291 ( P3_ADD_430_U181 , P3_REIP_REG_10_ , P3_ADD_430_U20 );
nand NAND2_20292 ( P3_ADD_430_U182 , P3_ADD_430_U101 , P3_ADD_430_U21 );
not NOT1_20293 ( P3_ADD_380_U5 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_20294 ( P3_ADD_380_U6 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_20295 ( P3_ADD_380_U7 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_20296 ( P3_ADD_380_U8 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_20297 ( P3_ADD_380_U9 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_380_U98 );
not NOT1_20298 ( P3_ADD_380_U10 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_20299 ( P3_ADD_380_U11 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_380_U99 );
not NOT1_20300 ( P3_ADD_380_U12 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_20301 ( P3_ADD_380_U13 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_380_U100 );
not NOT1_20302 ( P3_ADD_380_U14 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_20303 ( P3_ADD_380_U15 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_380_U101 );
not NOT1_20304 ( P3_ADD_380_U16 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_20305 ( P3_ADD_380_U17 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_380_U102 );
not NOT1_20306 ( P3_ADD_380_U18 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_20307 ( P3_ADD_380_U19 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_380_U103 );
not NOT1_20308 ( P3_ADD_380_U20 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_20309 ( P3_ADD_380_U21 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_20310 ( P3_ADD_380_U22 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_380_U104 );
nand NAND2_20311 ( P3_ADD_380_U23 , P3_ADD_380_U105 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_20312 ( P3_ADD_380_U24 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_20313 ( P3_ADD_380_U25 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_380_U106 );
not NOT1_20314 ( P3_ADD_380_U26 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_20315 ( P3_ADD_380_U27 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_380_U107 );
not NOT1_20316 ( P3_ADD_380_U28 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_20317 ( P3_ADD_380_U29 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_380_U108 );
not NOT1_20318 ( P3_ADD_380_U30 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_20319 ( P3_ADD_380_U31 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_380_U109 );
not NOT1_20320 ( P3_ADD_380_U32 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_20321 ( P3_ADD_380_U33 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_380_U110 );
not NOT1_20322 ( P3_ADD_380_U34 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_20323 ( P3_ADD_380_U35 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_380_U111 );
not NOT1_20324 ( P3_ADD_380_U36 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_20325 ( P3_ADD_380_U37 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_380_U112 );
not NOT1_20326 ( P3_ADD_380_U38 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_20327 ( P3_ADD_380_U39 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_380_U113 );
not NOT1_20328 ( P3_ADD_380_U40 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_20329 ( P3_ADD_380_U41 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_380_U114 );
not NOT1_20330 ( P3_ADD_380_U42 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_20331 ( P3_ADD_380_U43 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_380_U115 );
not NOT1_20332 ( P3_ADD_380_U44 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_20333 ( P3_ADD_380_U45 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_380_U116 );
not NOT1_20334 ( P3_ADD_380_U46 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_20335 ( P3_ADD_380_U47 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_380_U117 );
not NOT1_20336 ( P3_ADD_380_U48 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_20337 ( P3_ADD_380_U49 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_380_U118 );
not NOT1_20338 ( P3_ADD_380_U50 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_20339 ( P3_ADD_380_U51 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_380_U119 );
not NOT1_20340 ( P3_ADD_380_U52 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_20341 ( P3_ADD_380_U53 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_380_U120 );
not NOT1_20342 ( P3_ADD_380_U54 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_20343 ( P3_ADD_380_U55 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_380_U121 );
not NOT1_20344 ( P3_ADD_380_U56 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_20345 ( P3_ADD_380_U57 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_380_U122 );
not NOT1_20346 ( P3_ADD_380_U58 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_20347 ( P3_ADD_380_U59 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_380_U123 );
not NOT1_20348 ( P3_ADD_380_U60 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_20349 ( P3_ADD_380_U61 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_380_U124 );
not NOT1_20350 ( P3_ADD_380_U62 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_20351 ( P3_ADD_380_U63 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_380_U125 );
not NOT1_20352 ( P3_ADD_380_U64 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_20353 ( P3_ADD_380_U65 , P3_ADD_380_U129 , P3_ADD_380_U128 );
nand NAND2_20354 ( P3_ADD_380_U66 , P3_ADD_380_U131 , P3_ADD_380_U130 );
nand NAND2_20355 ( P3_ADD_380_U67 , P3_ADD_380_U133 , P3_ADD_380_U132 );
nand NAND2_20356 ( P3_ADD_380_U68 , P3_ADD_380_U135 , P3_ADD_380_U134 );
nand NAND2_20357 ( P3_ADD_380_U69 , P3_ADD_380_U137 , P3_ADD_380_U136 );
nand NAND2_20358 ( P3_ADD_380_U70 , P3_ADD_380_U139 , P3_ADD_380_U138 );
nand NAND2_20359 ( P3_ADD_380_U71 , P3_ADD_380_U141 , P3_ADD_380_U140 );
nand NAND2_20360 ( P3_ADD_380_U72 , P3_ADD_380_U143 , P3_ADD_380_U142 );
nand NAND2_20361 ( P3_ADD_380_U73 , P3_ADD_380_U145 , P3_ADD_380_U144 );
nand NAND2_20362 ( P3_ADD_380_U74 , P3_ADD_380_U147 , P3_ADD_380_U146 );
nand NAND2_20363 ( P3_ADD_380_U75 , P3_ADD_380_U149 , P3_ADD_380_U148 );
nand NAND2_20364 ( P3_ADD_380_U76 , P3_ADD_380_U151 , P3_ADD_380_U150 );
nand NAND2_20365 ( P3_ADD_380_U77 , P3_ADD_380_U153 , P3_ADD_380_U152 );
nand NAND2_20366 ( P3_ADD_380_U78 , P3_ADD_380_U155 , P3_ADD_380_U154 );
nand NAND2_20367 ( P3_ADD_380_U79 , P3_ADD_380_U157 , P3_ADD_380_U156 );
nand NAND2_20368 ( P3_ADD_380_U80 , P3_ADD_380_U159 , P3_ADD_380_U158 );
nand NAND2_20369 ( P3_ADD_380_U81 , P3_ADD_380_U161 , P3_ADD_380_U160 );
nand NAND2_20370 ( P3_ADD_380_U82 , P3_ADD_380_U163 , P3_ADD_380_U162 );
nand NAND2_20371 ( P3_ADD_380_U83 , P3_ADD_380_U165 , P3_ADD_380_U164 );
nand NAND2_20372 ( P3_ADD_380_U84 , P3_ADD_380_U167 , P3_ADD_380_U166 );
nand NAND2_20373 ( P3_ADD_380_U85 , P3_ADD_380_U169 , P3_ADD_380_U168 );
nand NAND2_20374 ( P3_ADD_380_U86 , P3_ADD_380_U171 , P3_ADD_380_U170 );
nand NAND2_20375 ( P3_ADD_380_U87 , P3_ADD_380_U173 , P3_ADD_380_U172 );
nand NAND2_20376 ( P3_ADD_380_U88 , P3_ADD_380_U175 , P3_ADD_380_U174 );
nand NAND2_20377 ( P3_ADD_380_U89 , P3_ADD_380_U177 , P3_ADD_380_U176 );
nand NAND2_20378 ( P3_ADD_380_U90 , P3_ADD_380_U179 , P3_ADD_380_U178 );
nand NAND2_20379 ( P3_ADD_380_U91 , P3_ADD_380_U181 , P3_ADD_380_U180 );
nand NAND2_20380 ( P3_ADD_380_U92 , P3_ADD_380_U183 , P3_ADD_380_U182 );
nand NAND2_20381 ( P3_ADD_380_U93 , P3_ADD_380_U185 , P3_ADD_380_U184 );
nand NAND2_20382 ( P3_ADD_380_U94 , P3_ADD_380_U187 , P3_ADD_380_U186 );
nand NAND2_20383 ( P3_ADD_380_U95 , P3_ADD_380_U189 , P3_ADD_380_U188 );
not NOT1_20384 ( P3_ADD_380_U96 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_20385 ( P3_ADD_380_U97 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_380_U126 );
not NOT1_20386 ( P3_ADD_380_U98 , P3_ADD_380_U7 );
not NOT1_20387 ( P3_ADD_380_U99 , P3_ADD_380_U9 );
not NOT1_20388 ( P3_ADD_380_U100 , P3_ADD_380_U11 );
not NOT1_20389 ( P3_ADD_380_U101 , P3_ADD_380_U13 );
not NOT1_20390 ( P3_ADD_380_U102 , P3_ADD_380_U15 );
not NOT1_20391 ( P3_ADD_380_U103 , P3_ADD_380_U17 );
not NOT1_20392 ( P3_ADD_380_U104 , P3_ADD_380_U19 );
not NOT1_20393 ( P3_ADD_380_U105 , P3_ADD_380_U22 );
not NOT1_20394 ( P3_ADD_380_U106 , P3_ADD_380_U23 );
not NOT1_20395 ( P3_ADD_380_U107 , P3_ADD_380_U25 );
not NOT1_20396 ( P3_ADD_380_U108 , P3_ADD_380_U27 );
not NOT1_20397 ( P3_ADD_380_U109 , P3_ADD_380_U29 );
not NOT1_20398 ( P3_ADD_380_U110 , P3_ADD_380_U31 );
not NOT1_20399 ( P3_ADD_380_U111 , P3_ADD_380_U33 );
not NOT1_20400 ( P3_ADD_380_U112 , P3_ADD_380_U35 );
not NOT1_20401 ( P3_ADD_380_U113 , P3_ADD_380_U37 );
not NOT1_20402 ( P3_ADD_380_U114 , P3_ADD_380_U39 );
not NOT1_20403 ( P3_ADD_380_U115 , P3_ADD_380_U41 );
not NOT1_20404 ( P3_ADD_380_U116 , P3_ADD_380_U43 );
not NOT1_20405 ( P3_ADD_380_U117 , P3_ADD_380_U45 );
not NOT1_20406 ( P3_ADD_380_U118 , P3_ADD_380_U47 );
not NOT1_20407 ( P3_ADD_380_U119 , P3_ADD_380_U49 );
not NOT1_20408 ( P3_ADD_380_U120 , P3_ADD_380_U51 );
not NOT1_20409 ( P3_ADD_380_U121 , P3_ADD_380_U53 );
not NOT1_20410 ( P3_ADD_380_U122 , P3_ADD_380_U55 );
not NOT1_20411 ( P3_ADD_380_U123 , P3_ADD_380_U57 );
not NOT1_20412 ( P3_ADD_380_U124 , P3_ADD_380_U59 );
not NOT1_20413 ( P3_ADD_380_U125 , P3_ADD_380_U61 );
not NOT1_20414 ( P3_ADD_380_U126 , P3_ADD_380_U63 );
not NOT1_20415 ( P3_ADD_380_U127 , P3_ADD_380_U97 );
nand NAND2_20416 ( P3_ADD_380_U128 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_380_U22 );
nand NAND2_20417 ( P3_ADD_380_U129 , P3_ADD_380_U105 , P3_ADD_380_U21 );
nand NAND2_20418 ( P3_ADD_380_U130 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_380_U19 );
nand NAND2_20419 ( P3_ADD_380_U131 , P3_ADD_380_U104 , P3_ADD_380_U20 );
nand NAND2_20420 ( P3_ADD_380_U132 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_380_U17 );
nand NAND2_20421 ( P3_ADD_380_U133 , P3_ADD_380_U103 , P3_ADD_380_U18 );
nand NAND2_20422 ( P3_ADD_380_U134 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_380_U15 );
nand NAND2_20423 ( P3_ADD_380_U135 , P3_ADD_380_U102 , P3_ADD_380_U16 );
nand NAND2_20424 ( P3_ADD_380_U136 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_380_U13 );
nand NAND2_20425 ( P3_ADD_380_U137 , P3_ADD_380_U101 , P3_ADD_380_U14 );
nand NAND2_20426 ( P3_ADD_380_U138 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_380_U11 );
nand NAND2_20427 ( P3_ADD_380_U139 , P3_ADD_380_U100 , P3_ADD_380_U12 );
nand NAND2_20428 ( P3_ADD_380_U140 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_380_U9 );
nand NAND2_20429 ( P3_ADD_380_U141 , P3_ADD_380_U99 , P3_ADD_380_U10 );
nand NAND2_20430 ( P3_ADD_380_U142 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_380_U97 );
nand NAND2_20431 ( P3_ADD_380_U143 , P3_ADD_380_U127 , P3_ADD_380_U96 );
nand NAND2_20432 ( P3_ADD_380_U144 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_380_U63 );
nand NAND2_20433 ( P3_ADD_380_U145 , P3_ADD_380_U126 , P3_ADD_380_U64 );
nand NAND2_20434 ( P3_ADD_380_U146 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_380_U7 );
nand NAND2_20435 ( P3_ADD_380_U147 , P3_ADD_380_U98 , P3_ADD_380_U8 );
nand NAND2_20436 ( P3_ADD_380_U148 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_380_U61 );
nand NAND2_20437 ( P3_ADD_380_U149 , P3_ADD_380_U125 , P3_ADD_380_U62 );
nand NAND2_20438 ( P3_ADD_380_U150 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_380_U59 );
nand NAND2_20439 ( P3_ADD_380_U151 , P3_ADD_380_U124 , P3_ADD_380_U60 );
nand NAND2_20440 ( P3_ADD_380_U152 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_380_U57 );
nand NAND2_20441 ( P3_ADD_380_U153 , P3_ADD_380_U123 , P3_ADD_380_U58 );
nand NAND2_20442 ( P3_ADD_380_U154 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_380_U55 );
nand NAND2_20443 ( P3_ADD_380_U155 , P3_ADD_380_U122 , P3_ADD_380_U56 );
nand NAND2_20444 ( P3_ADD_380_U156 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_380_U53 );
nand NAND2_20445 ( P3_ADD_380_U157 , P3_ADD_380_U121 , P3_ADD_380_U54 );
nand NAND2_20446 ( P3_ADD_380_U158 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_380_U51 );
nand NAND2_20447 ( P3_ADD_380_U159 , P3_ADD_380_U120 , P3_ADD_380_U52 );
nand NAND2_20448 ( P3_ADD_380_U160 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_380_U49 );
nand NAND2_20449 ( P3_ADD_380_U161 , P3_ADD_380_U119 , P3_ADD_380_U50 );
nand NAND2_20450 ( P3_ADD_380_U162 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_380_U47 );
nand NAND2_20451 ( P3_ADD_380_U163 , P3_ADD_380_U118 , P3_ADD_380_U48 );
nand NAND2_20452 ( P3_ADD_380_U164 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_380_U45 );
nand NAND2_20453 ( P3_ADD_380_U165 , P3_ADD_380_U117 , P3_ADD_380_U46 );
nand NAND2_20454 ( P3_ADD_380_U166 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_380_U43 );
nand NAND2_20455 ( P3_ADD_380_U167 , P3_ADD_380_U116 , P3_ADD_380_U44 );
nand NAND2_20456 ( P3_ADD_380_U168 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_380_U5 );
nand NAND2_20457 ( P3_ADD_380_U169 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_380_U6 );
nand NAND2_20458 ( P3_ADD_380_U170 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_380_U41 );
nand NAND2_20459 ( P3_ADD_380_U171 , P3_ADD_380_U115 , P3_ADD_380_U42 );
nand NAND2_20460 ( P3_ADD_380_U172 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_380_U39 );
nand NAND2_20461 ( P3_ADD_380_U173 , P3_ADD_380_U114 , P3_ADD_380_U40 );
nand NAND2_20462 ( P3_ADD_380_U174 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_380_U37 );
nand NAND2_20463 ( P3_ADD_380_U175 , P3_ADD_380_U113 , P3_ADD_380_U38 );
nand NAND2_20464 ( P3_ADD_380_U176 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_380_U35 );
nand NAND2_20465 ( P3_ADD_380_U177 , P3_ADD_380_U112 , P3_ADD_380_U36 );
nand NAND2_20466 ( P3_ADD_380_U178 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_380_U33 );
nand NAND2_20467 ( P3_ADD_380_U179 , P3_ADD_380_U111 , P3_ADD_380_U34 );
nand NAND2_20468 ( P3_ADD_380_U180 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_380_U31 );
nand NAND2_20469 ( P3_ADD_380_U181 , P3_ADD_380_U110 , P3_ADD_380_U32 );
nand NAND2_20470 ( P3_ADD_380_U182 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_380_U29 );
nand NAND2_20471 ( P3_ADD_380_U183 , P3_ADD_380_U109 , P3_ADD_380_U30 );
nand NAND2_20472 ( P3_ADD_380_U184 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_380_U27 );
nand NAND2_20473 ( P3_ADD_380_U185 , P3_ADD_380_U108 , P3_ADD_380_U28 );
nand NAND2_20474 ( P3_ADD_380_U186 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_380_U25 );
nand NAND2_20475 ( P3_ADD_380_U187 , P3_ADD_380_U107 , P3_ADD_380_U26 );
nand NAND2_20476 ( P3_ADD_380_U188 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_380_U23 );
nand NAND2_20477 ( P3_ADD_380_U189 , P3_ADD_380_U106 , P3_ADD_380_U24 );
nor nor_20478 ( P3_GTE_370_U6 , P3_SUB_370_U6 , P3_GTE_370_U8 );
and AND2_20479 ( P3_GTE_370_U7 , P3_SUB_370_U21 , P3_GTE_370_U9 );
nor nor_20480 ( P3_GTE_370_U8 , P3_SUB_370_U19 , P3_GTE_370_U7 , P3_SUB_370_U20 );
or OR2_20481 ( P3_GTE_370_U9 , P3_SUB_370_U7 , P3_SUB_370_U22 );
not NOT1_20482 ( P3_ADD_344_U5 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_20483 ( P3_ADD_344_U6 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_20484 ( P3_ADD_344_U7 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_20485 ( P3_ADD_344_U8 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_20486 ( P3_ADD_344_U9 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_344_U98 );
not NOT1_20487 ( P3_ADD_344_U10 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_20488 ( P3_ADD_344_U11 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_344_U99 );
not NOT1_20489 ( P3_ADD_344_U12 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_20490 ( P3_ADD_344_U13 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_344_U100 );
not NOT1_20491 ( P3_ADD_344_U14 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_20492 ( P3_ADD_344_U15 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_344_U101 );
not NOT1_20493 ( P3_ADD_344_U16 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_20494 ( P3_ADD_344_U17 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_344_U102 );
not NOT1_20495 ( P3_ADD_344_U18 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_20496 ( P3_ADD_344_U19 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_344_U103 );
not NOT1_20497 ( P3_ADD_344_U20 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_20498 ( P3_ADD_344_U21 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_20499 ( P3_ADD_344_U22 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_344_U104 );
nand NAND2_20500 ( P3_ADD_344_U23 , P3_ADD_344_U105 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_20501 ( P3_ADD_344_U24 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_20502 ( P3_ADD_344_U25 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_344_U106 );
not NOT1_20503 ( P3_ADD_344_U26 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_20504 ( P3_ADD_344_U27 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_344_U107 );
not NOT1_20505 ( P3_ADD_344_U28 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_20506 ( P3_ADD_344_U29 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_344_U108 );
not NOT1_20507 ( P3_ADD_344_U30 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_20508 ( P3_ADD_344_U31 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_344_U109 );
not NOT1_20509 ( P3_ADD_344_U32 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_20510 ( P3_ADD_344_U33 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_344_U110 );
not NOT1_20511 ( P3_ADD_344_U34 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_20512 ( P3_ADD_344_U35 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_344_U111 );
not NOT1_20513 ( P3_ADD_344_U36 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_20514 ( P3_ADD_344_U37 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_344_U112 );
not NOT1_20515 ( P3_ADD_344_U38 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_20516 ( P3_ADD_344_U39 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_344_U113 );
not NOT1_20517 ( P3_ADD_344_U40 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_20518 ( P3_ADD_344_U41 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_344_U114 );
not NOT1_20519 ( P3_ADD_344_U42 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_20520 ( P3_ADD_344_U43 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_344_U115 );
not NOT1_20521 ( P3_ADD_344_U44 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_20522 ( P3_ADD_344_U45 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_344_U116 );
not NOT1_20523 ( P3_ADD_344_U46 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_20524 ( P3_ADD_344_U47 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_344_U117 );
not NOT1_20525 ( P3_ADD_344_U48 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_20526 ( P3_ADD_344_U49 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_344_U118 );
not NOT1_20527 ( P3_ADD_344_U50 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_20528 ( P3_ADD_344_U51 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_344_U119 );
not NOT1_20529 ( P3_ADD_344_U52 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_20530 ( P3_ADD_344_U53 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_344_U120 );
not NOT1_20531 ( P3_ADD_344_U54 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_20532 ( P3_ADD_344_U55 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_344_U121 );
not NOT1_20533 ( P3_ADD_344_U56 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_20534 ( P3_ADD_344_U57 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_344_U122 );
not NOT1_20535 ( P3_ADD_344_U58 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_20536 ( P3_ADD_344_U59 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_344_U123 );
not NOT1_20537 ( P3_ADD_344_U60 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_20538 ( P3_ADD_344_U61 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_344_U124 );
not NOT1_20539 ( P3_ADD_344_U62 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_20540 ( P3_ADD_344_U63 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_344_U125 );
not NOT1_20541 ( P3_ADD_344_U64 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_20542 ( P3_ADD_344_U65 , P3_ADD_344_U129 , P3_ADD_344_U128 );
nand NAND2_20543 ( P3_ADD_344_U66 , P3_ADD_344_U131 , P3_ADD_344_U130 );
nand NAND2_20544 ( P3_ADD_344_U67 , P3_ADD_344_U133 , P3_ADD_344_U132 );
nand NAND2_20545 ( P3_ADD_344_U68 , P3_ADD_344_U135 , P3_ADD_344_U134 );
nand NAND2_20546 ( P3_ADD_344_U69 , P3_ADD_344_U137 , P3_ADD_344_U136 );
nand NAND2_20547 ( P3_ADD_344_U70 , P3_ADD_344_U139 , P3_ADD_344_U138 );
nand NAND2_20548 ( P3_ADD_344_U71 , P3_ADD_344_U141 , P3_ADD_344_U140 );
nand NAND2_20549 ( P3_ADD_344_U72 , P3_ADD_344_U143 , P3_ADD_344_U142 );
nand NAND2_20550 ( P3_ADD_344_U73 , P3_ADD_344_U145 , P3_ADD_344_U144 );
nand NAND2_20551 ( P3_ADD_344_U74 , P3_ADD_344_U147 , P3_ADD_344_U146 );
nand NAND2_20552 ( P3_ADD_344_U75 , P3_ADD_344_U149 , P3_ADD_344_U148 );
nand NAND2_20553 ( P3_ADD_344_U76 , P3_ADD_344_U151 , P3_ADD_344_U150 );
nand NAND2_20554 ( P3_ADD_344_U77 , P3_ADD_344_U153 , P3_ADD_344_U152 );
nand NAND2_20555 ( P3_ADD_344_U78 , P3_ADD_344_U155 , P3_ADD_344_U154 );
nand NAND2_20556 ( P3_ADD_344_U79 , P3_ADD_344_U157 , P3_ADD_344_U156 );
nand NAND2_20557 ( P3_ADD_344_U80 , P3_ADD_344_U159 , P3_ADD_344_U158 );
nand NAND2_20558 ( P3_ADD_344_U81 , P3_ADD_344_U161 , P3_ADD_344_U160 );
nand NAND2_20559 ( P3_ADD_344_U82 , P3_ADD_344_U163 , P3_ADD_344_U162 );
nand NAND2_20560 ( P3_ADD_344_U83 , P3_ADD_344_U165 , P3_ADD_344_U164 );
nand NAND2_20561 ( P3_ADD_344_U84 , P3_ADD_344_U167 , P3_ADD_344_U166 );
nand NAND2_20562 ( P3_ADD_344_U85 , P3_ADD_344_U169 , P3_ADD_344_U168 );
nand NAND2_20563 ( P3_ADD_344_U86 , P3_ADD_344_U171 , P3_ADD_344_U170 );
nand NAND2_20564 ( P3_ADD_344_U87 , P3_ADD_344_U173 , P3_ADD_344_U172 );
nand NAND2_20565 ( P3_ADD_344_U88 , P3_ADD_344_U175 , P3_ADD_344_U174 );
nand NAND2_20566 ( P3_ADD_344_U89 , P3_ADD_344_U177 , P3_ADD_344_U176 );
nand NAND2_20567 ( P3_ADD_344_U90 , P3_ADD_344_U179 , P3_ADD_344_U178 );
nand NAND2_20568 ( P3_ADD_344_U91 , P3_ADD_344_U181 , P3_ADD_344_U180 );
nand NAND2_20569 ( P3_ADD_344_U92 , P3_ADD_344_U183 , P3_ADD_344_U182 );
nand NAND2_20570 ( P3_ADD_344_U93 , P3_ADD_344_U185 , P3_ADD_344_U184 );
nand NAND2_20571 ( P3_ADD_344_U94 , P3_ADD_344_U187 , P3_ADD_344_U186 );
nand NAND2_20572 ( P3_ADD_344_U95 , P3_ADD_344_U189 , P3_ADD_344_U188 );
not NOT1_20573 ( P3_ADD_344_U96 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_20574 ( P3_ADD_344_U97 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_344_U126 );
not NOT1_20575 ( P3_ADD_344_U98 , P3_ADD_344_U7 );
not NOT1_20576 ( P3_ADD_344_U99 , P3_ADD_344_U9 );
not NOT1_20577 ( P3_ADD_344_U100 , P3_ADD_344_U11 );
not NOT1_20578 ( P3_ADD_344_U101 , P3_ADD_344_U13 );
not NOT1_20579 ( P3_ADD_344_U102 , P3_ADD_344_U15 );
not NOT1_20580 ( P3_ADD_344_U103 , P3_ADD_344_U17 );
not NOT1_20581 ( P3_ADD_344_U104 , P3_ADD_344_U19 );
not NOT1_20582 ( P3_ADD_344_U105 , P3_ADD_344_U22 );
not NOT1_20583 ( P3_ADD_344_U106 , P3_ADD_344_U23 );
not NOT1_20584 ( P3_ADD_344_U107 , P3_ADD_344_U25 );
not NOT1_20585 ( P3_ADD_344_U108 , P3_ADD_344_U27 );
not NOT1_20586 ( P3_ADD_344_U109 , P3_ADD_344_U29 );
not NOT1_20587 ( P3_ADD_344_U110 , P3_ADD_344_U31 );
not NOT1_20588 ( P3_ADD_344_U111 , P3_ADD_344_U33 );
not NOT1_20589 ( P3_ADD_344_U112 , P3_ADD_344_U35 );
not NOT1_20590 ( P3_ADD_344_U113 , P3_ADD_344_U37 );
not NOT1_20591 ( P3_ADD_344_U114 , P3_ADD_344_U39 );
not NOT1_20592 ( P3_ADD_344_U115 , P3_ADD_344_U41 );
not NOT1_20593 ( P3_ADD_344_U116 , P3_ADD_344_U43 );
not NOT1_20594 ( P3_ADD_344_U117 , P3_ADD_344_U45 );
not NOT1_20595 ( P3_ADD_344_U118 , P3_ADD_344_U47 );
not NOT1_20596 ( P3_ADD_344_U119 , P3_ADD_344_U49 );
not NOT1_20597 ( P3_ADD_344_U120 , P3_ADD_344_U51 );
not NOT1_20598 ( P3_ADD_344_U121 , P3_ADD_344_U53 );
not NOT1_20599 ( P3_ADD_344_U122 , P3_ADD_344_U55 );
not NOT1_20600 ( P3_ADD_344_U123 , P3_ADD_344_U57 );
not NOT1_20601 ( P3_ADD_344_U124 , P3_ADD_344_U59 );
not NOT1_20602 ( P3_ADD_344_U125 , P3_ADD_344_U61 );
not NOT1_20603 ( P3_ADD_344_U126 , P3_ADD_344_U63 );
not NOT1_20604 ( P3_ADD_344_U127 , P3_ADD_344_U97 );
nand NAND2_20605 ( P3_ADD_344_U128 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_344_U22 );
nand NAND2_20606 ( P3_ADD_344_U129 , P3_ADD_344_U105 , P3_ADD_344_U21 );
nand NAND2_20607 ( P3_ADD_344_U130 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_344_U19 );
nand NAND2_20608 ( P3_ADD_344_U131 , P3_ADD_344_U104 , P3_ADD_344_U20 );
nand NAND2_20609 ( P3_ADD_344_U132 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_344_U17 );
nand NAND2_20610 ( P3_ADD_344_U133 , P3_ADD_344_U103 , P3_ADD_344_U18 );
nand NAND2_20611 ( P3_ADD_344_U134 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_344_U15 );
nand NAND2_20612 ( P3_ADD_344_U135 , P3_ADD_344_U102 , P3_ADD_344_U16 );
nand NAND2_20613 ( P3_ADD_344_U136 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_344_U13 );
nand NAND2_20614 ( P3_ADD_344_U137 , P3_ADD_344_U101 , P3_ADD_344_U14 );
nand NAND2_20615 ( P3_ADD_344_U138 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_344_U11 );
nand NAND2_20616 ( P3_ADD_344_U139 , P3_ADD_344_U100 , P3_ADD_344_U12 );
nand NAND2_20617 ( P3_ADD_344_U140 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_344_U9 );
nand NAND2_20618 ( P3_ADD_344_U141 , P3_ADD_344_U99 , P3_ADD_344_U10 );
nand NAND2_20619 ( P3_ADD_344_U142 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_344_U97 );
nand NAND2_20620 ( P3_ADD_344_U143 , P3_ADD_344_U127 , P3_ADD_344_U96 );
nand NAND2_20621 ( P3_ADD_344_U144 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_344_U63 );
nand NAND2_20622 ( P3_ADD_344_U145 , P3_ADD_344_U126 , P3_ADD_344_U64 );
nand NAND2_20623 ( P3_ADD_344_U146 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_344_U7 );
nand NAND2_20624 ( P3_ADD_344_U147 , P3_ADD_344_U98 , P3_ADD_344_U8 );
nand NAND2_20625 ( P3_ADD_344_U148 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_344_U61 );
nand NAND2_20626 ( P3_ADD_344_U149 , P3_ADD_344_U125 , P3_ADD_344_U62 );
nand NAND2_20627 ( P3_ADD_344_U150 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_344_U59 );
nand NAND2_20628 ( P3_ADD_344_U151 , P3_ADD_344_U124 , P3_ADD_344_U60 );
nand NAND2_20629 ( P3_ADD_344_U152 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_344_U57 );
nand NAND2_20630 ( P3_ADD_344_U153 , P3_ADD_344_U123 , P3_ADD_344_U58 );
nand NAND2_20631 ( P3_ADD_344_U154 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_344_U55 );
nand NAND2_20632 ( P3_ADD_344_U155 , P3_ADD_344_U122 , P3_ADD_344_U56 );
nand NAND2_20633 ( P3_ADD_344_U156 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_344_U53 );
nand NAND2_20634 ( P3_ADD_344_U157 , P3_ADD_344_U121 , P3_ADD_344_U54 );
nand NAND2_20635 ( P3_ADD_344_U158 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_344_U51 );
nand NAND2_20636 ( P3_ADD_344_U159 , P3_ADD_344_U120 , P3_ADD_344_U52 );
nand NAND2_20637 ( P3_ADD_344_U160 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_344_U49 );
nand NAND2_20638 ( P3_ADD_344_U161 , P3_ADD_344_U119 , P3_ADD_344_U50 );
nand NAND2_20639 ( P3_ADD_344_U162 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_344_U47 );
nand NAND2_20640 ( P3_ADD_344_U163 , P3_ADD_344_U118 , P3_ADD_344_U48 );
nand NAND2_20641 ( P3_ADD_344_U164 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_344_U45 );
nand NAND2_20642 ( P3_ADD_344_U165 , P3_ADD_344_U117 , P3_ADD_344_U46 );
nand NAND2_20643 ( P3_ADD_344_U166 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_344_U43 );
nand NAND2_20644 ( P3_ADD_344_U167 , P3_ADD_344_U116 , P3_ADD_344_U44 );
nand NAND2_20645 ( P3_ADD_344_U168 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_344_U5 );
nand NAND2_20646 ( P3_ADD_344_U169 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_344_U6 );
nand NAND2_20647 ( P3_ADD_344_U170 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_344_U41 );
nand NAND2_20648 ( P3_ADD_344_U171 , P3_ADD_344_U115 , P3_ADD_344_U42 );
nand NAND2_20649 ( P3_ADD_344_U172 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_344_U39 );
nand NAND2_20650 ( P3_ADD_344_U173 , P3_ADD_344_U114 , P3_ADD_344_U40 );
nand NAND2_20651 ( P3_ADD_344_U174 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_344_U37 );
nand NAND2_20652 ( P3_ADD_344_U175 , P3_ADD_344_U113 , P3_ADD_344_U38 );
nand NAND2_20653 ( P3_ADD_344_U176 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_344_U35 );
nand NAND2_20654 ( P3_ADD_344_U177 , P3_ADD_344_U112 , P3_ADD_344_U36 );
nand NAND2_20655 ( P3_ADD_344_U178 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_344_U33 );
nand NAND2_20656 ( P3_ADD_344_U179 , P3_ADD_344_U111 , P3_ADD_344_U34 );
nand NAND2_20657 ( P3_ADD_344_U180 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_344_U31 );
nand NAND2_20658 ( P3_ADD_344_U181 , P3_ADD_344_U110 , P3_ADD_344_U32 );
nand NAND2_20659 ( P3_ADD_344_U182 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_344_U29 );
nand NAND2_20660 ( P3_ADD_344_U183 , P3_ADD_344_U109 , P3_ADD_344_U30 );
nand NAND2_20661 ( P3_ADD_344_U184 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_344_U27 );
nand NAND2_20662 ( P3_ADD_344_U185 , P3_ADD_344_U108 , P3_ADD_344_U28 );
nand NAND2_20663 ( P3_ADD_344_U186 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_344_U25 );
nand NAND2_20664 ( P3_ADD_344_U187 , P3_ADD_344_U107 , P3_ADD_344_U26 );
nand NAND2_20665 ( P3_ADD_344_U188 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_344_U23 );
nand NAND2_20666 ( P3_ADD_344_U189 , P3_ADD_344_U106 , P3_ADD_344_U24 );
nand NAND2_20667 ( P3_LT_563_U6 , P3_LT_563_U27 , P3_LT_563_U28 );
not NOT1_20668 ( P3_LT_563_U7 , P3_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_20669 ( P3_LT_563_U8 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_LT_563_U15 );
not NOT1_20670 ( P3_LT_563_U9 , P3_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_20671 ( P3_LT_563_U10 , P3_U3306 );
not NOT1_20672 ( P3_LT_563_U11 , P3_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_20673 ( P3_LT_563_U12 , P3_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_20674 ( P3_LT_563_U13 , P3_U3305 );
not NOT1_20675 ( P3_LT_563_U14 , P3_U3304 );
not NOT1_20676 ( P3_LT_563_U15 , P3_U3308 );
not NOT1_20677 ( P3_LT_563_U16 , P3_LT_563_U8 );
nand NAND2_20678 ( P3_LT_563_U17 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_LT_563_U16 );
nand NAND2_20679 ( P3_LT_563_U18 , P3_U3307 , P3_LT_563_U17 );
nand NAND2_20680 ( P3_LT_563_U19 , P3_LT_563_U8 , P3_LT_563_U9 );
nand NAND2_20681 ( P3_LT_563_U20 , P3_U3306 , P3_LT_563_U11 );
nand NAND3_20682 ( P3_LT_563_U21 , P3_LT_563_U19 , P3_LT_563_U20 , P3_LT_563_U18 );
nand NAND2_20683 ( P3_LT_563_U22 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_LT_563_U10 );
nand NAND2_20684 ( P3_LT_563_U23 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_LT_563_U13 );
nand NAND3_20685 ( P3_LT_563_U24 , P3_LT_563_U22 , P3_LT_563_U23 , P3_LT_563_U21 );
nand NAND2_20686 ( P3_LT_563_U25 , P3_U3305 , P3_LT_563_U12 );
nand NAND2_20687 ( P3_LT_563_U26 , P3_U3304 , P3_LT_563_U7 );
nand NAND3_20688 ( P3_LT_563_U27 , P3_LT_563_U25 , P3_LT_563_U26 , P3_LT_563_U24 );
nand NAND2_20689 ( P3_LT_563_U28 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_LT_563_U14 );
not NOT1_20690 ( P3_ADD_339_U4 , P3_PHYADDRPOINTER_REG_1_ );
not NOT1_20691 ( P3_ADD_339_U5 , P3_PHYADDRPOINTER_REG_2_ );
nand NAND2_20692 ( P3_ADD_339_U6 , P3_PHYADDRPOINTER_REG_2_ , P3_PHYADDRPOINTER_REG_1_ );
not NOT1_20693 ( P3_ADD_339_U7 , P3_PHYADDRPOINTER_REG_3_ );
nand NAND2_20694 ( P3_ADD_339_U8 , P3_PHYADDRPOINTER_REG_3_ , P3_ADD_339_U94 );
not NOT1_20695 ( P3_ADD_339_U9 , P3_PHYADDRPOINTER_REG_4_ );
nand NAND2_20696 ( P3_ADD_339_U10 , P3_PHYADDRPOINTER_REG_4_ , P3_ADD_339_U95 );
not NOT1_20697 ( P3_ADD_339_U11 , P3_PHYADDRPOINTER_REG_5_ );
nand NAND2_20698 ( P3_ADD_339_U12 , P3_PHYADDRPOINTER_REG_5_ , P3_ADD_339_U96 );
not NOT1_20699 ( P3_ADD_339_U13 , P3_PHYADDRPOINTER_REG_6_ );
nand NAND2_20700 ( P3_ADD_339_U14 , P3_PHYADDRPOINTER_REG_6_ , P3_ADD_339_U97 );
not NOT1_20701 ( P3_ADD_339_U15 , P3_PHYADDRPOINTER_REG_7_ );
nand NAND2_20702 ( P3_ADD_339_U16 , P3_PHYADDRPOINTER_REG_7_ , P3_ADD_339_U98 );
not NOT1_20703 ( P3_ADD_339_U17 , P3_PHYADDRPOINTER_REG_8_ );
not NOT1_20704 ( P3_ADD_339_U18 , P3_PHYADDRPOINTER_REG_9_ );
nand NAND2_20705 ( P3_ADD_339_U19 , P3_PHYADDRPOINTER_REG_8_ , P3_ADD_339_U99 );
nand NAND2_20706 ( P3_ADD_339_U20 , P3_ADD_339_U100 , P3_PHYADDRPOINTER_REG_9_ );
not NOT1_20707 ( P3_ADD_339_U21 , P3_PHYADDRPOINTER_REG_10_ );
nand NAND2_20708 ( P3_ADD_339_U22 , P3_PHYADDRPOINTER_REG_10_ , P3_ADD_339_U101 );
not NOT1_20709 ( P3_ADD_339_U23 , P3_PHYADDRPOINTER_REG_11_ );
nand NAND2_20710 ( P3_ADD_339_U24 , P3_PHYADDRPOINTER_REG_11_ , P3_ADD_339_U102 );
not NOT1_20711 ( P3_ADD_339_U25 , P3_PHYADDRPOINTER_REG_12_ );
nand NAND2_20712 ( P3_ADD_339_U26 , P3_PHYADDRPOINTER_REG_12_ , P3_ADD_339_U103 );
not NOT1_20713 ( P3_ADD_339_U27 , P3_PHYADDRPOINTER_REG_13_ );
nand NAND2_20714 ( P3_ADD_339_U28 , P3_PHYADDRPOINTER_REG_13_ , P3_ADD_339_U104 );
not NOT1_20715 ( P3_ADD_339_U29 , P3_PHYADDRPOINTER_REG_14_ );
nand NAND2_20716 ( P3_ADD_339_U30 , P3_PHYADDRPOINTER_REG_14_ , P3_ADD_339_U105 );
not NOT1_20717 ( P3_ADD_339_U31 , P3_PHYADDRPOINTER_REG_15_ );
nand NAND2_20718 ( P3_ADD_339_U32 , P3_PHYADDRPOINTER_REG_15_ , P3_ADD_339_U106 );
not NOT1_20719 ( P3_ADD_339_U33 , P3_PHYADDRPOINTER_REG_16_ );
nand NAND2_20720 ( P3_ADD_339_U34 , P3_PHYADDRPOINTER_REG_16_ , P3_ADD_339_U107 );
not NOT1_20721 ( P3_ADD_339_U35 , P3_PHYADDRPOINTER_REG_17_ );
nand NAND2_20722 ( P3_ADD_339_U36 , P3_PHYADDRPOINTER_REG_17_ , P3_ADD_339_U108 );
not NOT1_20723 ( P3_ADD_339_U37 , P3_PHYADDRPOINTER_REG_18_ );
nand NAND2_20724 ( P3_ADD_339_U38 , P3_PHYADDRPOINTER_REG_18_ , P3_ADD_339_U109 );
not NOT1_20725 ( P3_ADD_339_U39 , P3_PHYADDRPOINTER_REG_19_ );
nand NAND2_20726 ( P3_ADD_339_U40 , P3_PHYADDRPOINTER_REG_19_ , P3_ADD_339_U110 );
not NOT1_20727 ( P3_ADD_339_U41 , P3_PHYADDRPOINTER_REG_20_ );
nand NAND2_20728 ( P3_ADD_339_U42 , P3_PHYADDRPOINTER_REG_20_ , P3_ADD_339_U111 );
not NOT1_20729 ( P3_ADD_339_U43 , P3_PHYADDRPOINTER_REG_21_ );
nand NAND2_20730 ( P3_ADD_339_U44 , P3_PHYADDRPOINTER_REG_21_ , P3_ADD_339_U112 );
not NOT1_20731 ( P3_ADD_339_U45 , P3_PHYADDRPOINTER_REG_22_ );
nand NAND2_20732 ( P3_ADD_339_U46 , P3_PHYADDRPOINTER_REG_22_ , P3_ADD_339_U113 );
not NOT1_20733 ( P3_ADD_339_U47 , P3_PHYADDRPOINTER_REG_23_ );
nand NAND2_20734 ( P3_ADD_339_U48 , P3_PHYADDRPOINTER_REG_23_ , P3_ADD_339_U114 );
not NOT1_20735 ( P3_ADD_339_U49 , P3_PHYADDRPOINTER_REG_24_ );
nand NAND2_20736 ( P3_ADD_339_U50 , P3_PHYADDRPOINTER_REG_24_ , P3_ADD_339_U115 );
not NOT1_20737 ( P3_ADD_339_U51 , P3_PHYADDRPOINTER_REG_25_ );
nand NAND2_20738 ( P3_ADD_339_U52 , P3_PHYADDRPOINTER_REG_25_ , P3_ADD_339_U116 );
not NOT1_20739 ( P3_ADD_339_U53 , P3_PHYADDRPOINTER_REG_26_ );
nand NAND2_20740 ( P3_ADD_339_U54 , P3_PHYADDRPOINTER_REG_26_ , P3_ADD_339_U117 );
not NOT1_20741 ( P3_ADD_339_U55 , P3_PHYADDRPOINTER_REG_27_ );
nand NAND2_20742 ( P3_ADD_339_U56 , P3_PHYADDRPOINTER_REG_27_ , P3_ADD_339_U118 );
not NOT1_20743 ( P3_ADD_339_U57 , P3_PHYADDRPOINTER_REG_28_ );
nand NAND2_20744 ( P3_ADD_339_U58 , P3_PHYADDRPOINTER_REG_28_ , P3_ADD_339_U119 );
not NOT1_20745 ( P3_ADD_339_U59 , P3_PHYADDRPOINTER_REG_29_ );
nand NAND2_20746 ( P3_ADD_339_U60 , P3_PHYADDRPOINTER_REG_29_ , P3_ADD_339_U120 );
not NOT1_20747 ( P3_ADD_339_U61 , P3_PHYADDRPOINTER_REG_30_ );
nand NAND2_20748 ( P3_ADD_339_U62 , P3_ADD_339_U124 , P3_ADD_339_U123 );
nand NAND2_20749 ( P3_ADD_339_U63 , P3_ADD_339_U126 , P3_ADD_339_U125 );
nand NAND2_20750 ( P3_ADD_339_U64 , P3_ADD_339_U128 , P3_ADD_339_U127 );
nand NAND2_20751 ( P3_ADD_339_U65 , P3_ADD_339_U130 , P3_ADD_339_U129 );
nand NAND2_20752 ( P3_ADD_339_U66 , P3_ADD_339_U132 , P3_ADD_339_U131 );
nand NAND2_20753 ( P3_ADD_339_U67 , P3_ADD_339_U134 , P3_ADD_339_U133 );
nand NAND2_20754 ( P3_ADD_339_U68 , P3_ADD_339_U136 , P3_ADD_339_U135 );
nand NAND2_20755 ( P3_ADD_339_U69 , P3_ADD_339_U138 , P3_ADD_339_U137 );
nand NAND2_20756 ( P3_ADD_339_U70 , P3_ADD_339_U140 , P3_ADD_339_U139 );
nand NAND2_20757 ( P3_ADD_339_U71 , P3_ADD_339_U142 , P3_ADD_339_U141 );
nand NAND2_20758 ( P3_ADD_339_U72 , P3_ADD_339_U144 , P3_ADD_339_U143 );
nand NAND2_20759 ( P3_ADD_339_U73 , P3_ADD_339_U146 , P3_ADD_339_U145 );
nand NAND2_20760 ( P3_ADD_339_U74 , P3_ADD_339_U148 , P3_ADD_339_U147 );
nand NAND2_20761 ( P3_ADD_339_U75 , P3_ADD_339_U150 , P3_ADD_339_U149 );
nand NAND2_20762 ( P3_ADD_339_U76 , P3_ADD_339_U152 , P3_ADD_339_U151 );
nand NAND2_20763 ( P3_ADD_339_U77 , P3_ADD_339_U154 , P3_ADD_339_U153 );
nand NAND2_20764 ( P3_ADD_339_U78 , P3_ADD_339_U156 , P3_ADD_339_U155 );
nand NAND2_20765 ( P3_ADD_339_U79 , P3_ADD_339_U158 , P3_ADD_339_U157 );
nand NAND2_20766 ( P3_ADD_339_U80 , P3_ADD_339_U160 , P3_ADD_339_U159 );
nand NAND2_20767 ( P3_ADD_339_U81 , P3_ADD_339_U162 , P3_ADD_339_U161 );
nand NAND2_20768 ( P3_ADD_339_U82 , P3_ADD_339_U164 , P3_ADD_339_U163 );
nand NAND2_20769 ( P3_ADD_339_U83 , P3_ADD_339_U166 , P3_ADD_339_U165 );
nand NAND2_20770 ( P3_ADD_339_U84 , P3_ADD_339_U168 , P3_ADD_339_U167 );
nand NAND2_20771 ( P3_ADD_339_U85 , P3_ADD_339_U170 , P3_ADD_339_U169 );
nand NAND2_20772 ( P3_ADD_339_U86 , P3_ADD_339_U172 , P3_ADD_339_U171 );
nand NAND2_20773 ( P3_ADD_339_U87 , P3_ADD_339_U174 , P3_ADD_339_U173 );
nand NAND2_20774 ( P3_ADD_339_U88 , P3_ADD_339_U176 , P3_ADD_339_U175 );
nand NAND2_20775 ( P3_ADD_339_U89 , P3_ADD_339_U178 , P3_ADD_339_U177 );
nand NAND2_20776 ( P3_ADD_339_U90 , P3_ADD_339_U180 , P3_ADD_339_U179 );
nand NAND2_20777 ( P3_ADD_339_U91 , P3_ADD_339_U182 , P3_ADD_339_U181 );
not NOT1_20778 ( P3_ADD_339_U92 , P3_PHYADDRPOINTER_REG_31_ );
nand NAND2_20779 ( P3_ADD_339_U93 , P3_PHYADDRPOINTER_REG_30_ , P3_ADD_339_U121 );
not NOT1_20780 ( P3_ADD_339_U94 , P3_ADD_339_U6 );
not NOT1_20781 ( P3_ADD_339_U95 , P3_ADD_339_U8 );
not NOT1_20782 ( P3_ADD_339_U96 , P3_ADD_339_U10 );
not NOT1_20783 ( P3_ADD_339_U97 , P3_ADD_339_U12 );
not NOT1_20784 ( P3_ADD_339_U98 , P3_ADD_339_U14 );
not NOT1_20785 ( P3_ADD_339_U99 , P3_ADD_339_U16 );
not NOT1_20786 ( P3_ADD_339_U100 , P3_ADD_339_U19 );
not NOT1_20787 ( P3_ADD_339_U101 , P3_ADD_339_U20 );
not NOT1_20788 ( P3_ADD_339_U102 , P3_ADD_339_U22 );
not NOT1_20789 ( P3_ADD_339_U103 , P3_ADD_339_U24 );
not NOT1_20790 ( P3_ADD_339_U104 , P3_ADD_339_U26 );
not NOT1_20791 ( P3_ADD_339_U105 , P3_ADD_339_U28 );
not NOT1_20792 ( P3_ADD_339_U106 , P3_ADD_339_U30 );
not NOT1_20793 ( P3_ADD_339_U107 , P3_ADD_339_U32 );
not NOT1_20794 ( P3_ADD_339_U108 , P3_ADD_339_U34 );
not NOT1_20795 ( P3_ADD_339_U109 , P3_ADD_339_U36 );
not NOT1_20796 ( P3_ADD_339_U110 , P3_ADD_339_U38 );
not NOT1_20797 ( P3_ADD_339_U111 , P3_ADD_339_U40 );
not NOT1_20798 ( P3_ADD_339_U112 , P3_ADD_339_U42 );
not NOT1_20799 ( P3_ADD_339_U113 , P3_ADD_339_U44 );
not NOT1_20800 ( P3_ADD_339_U114 , P3_ADD_339_U46 );
not NOT1_20801 ( P3_ADD_339_U115 , P3_ADD_339_U48 );
not NOT1_20802 ( P3_ADD_339_U116 , P3_ADD_339_U50 );
not NOT1_20803 ( P3_ADD_339_U117 , P3_ADD_339_U52 );
not NOT1_20804 ( P3_ADD_339_U118 , P3_ADD_339_U54 );
not NOT1_20805 ( P3_ADD_339_U119 , P3_ADD_339_U56 );
not NOT1_20806 ( P3_ADD_339_U120 , P3_ADD_339_U58 );
not NOT1_20807 ( P3_ADD_339_U121 , P3_ADD_339_U60 );
not NOT1_20808 ( P3_ADD_339_U122 , P3_ADD_339_U93 );
nand NAND2_20809 ( P3_ADD_339_U123 , P3_PHYADDRPOINTER_REG_9_ , P3_ADD_339_U19 );
nand NAND2_20810 ( P3_ADD_339_U124 , P3_ADD_339_U100 , P3_ADD_339_U18 );
nand NAND2_20811 ( P3_ADD_339_U125 , P3_PHYADDRPOINTER_REG_8_ , P3_ADD_339_U16 );
nand NAND2_20812 ( P3_ADD_339_U126 , P3_ADD_339_U99 , P3_ADD_339_U17 );
nand NAND2_20813 ( P3_ADD_339_U127 , P3_PHYADDRPOINTER_REG_7_ , P3_ADD_339_U14 );
nand NAND2_20814 ( P3_ADD_339_U128 , P3_ADD_339_U98 , P3_ADD_339_U15 );
nand NAND2_20815 ( P3_ADD_339_U129 , P3_PHYADDRPOINTER_REG_6_ , P3_ADD_339_U12 );
nand NAND2_20816 ( P3_ADD_339_U130 , P3_ADD_339_U97 , P3_ADD_339_U13 );
nand NAND2_20817 ( P3_ADD_339_U131 , P3_PHYADDRPOINTER_REG_5_ , P3_ADD_339_U10 );
nand NAND2_20818 ( P3_ADD_339_U132 , P3_ADD_339_U96 , P3_ADD_339_U11 );
nand NAND2_20819 ( P3_ADD_339_U133 , P3_PHYADDRPOINTER_REG_4_ , P3_ADD_339_U8 );
nand NAND2_20820 ( P3_ADD_339_U134 , P3_ADD_339_U95 , P3_ADD_339_U9 );
nand NAND2_20821 ( P3_ADD_339_U135 , P3_PHYADDRPOINTER_REG_3_ , P3_ADD_339_U6 );
nand NAND2_20822 ( P3_ADD_339_U136 , P3_ADD_339_U94 , P3_ADD_339_U7 );
nand NAND2_20823 ( P3_ADD_339_U137 , P3_PHYADDRPOINTER_REG_31_ , P3_ADD_339_U93 );
nand NAND2_20824 ( P3_ADD_339_U138 , P3_ADD_339_U122 , P3_ADD_339_U92 );
nand NAND2_20825 ( P3_ADD_339_U139 , P3_PHYADDRPOINTER_REG_30_ , P3_ADD_339_U60 );
nand NAND2_20826 ( P3_ADD_339_U140 , P3_ADD_339_U121 , P3_ADD_339_U61 );
nand NAND2_20827 ( P3_ADD_339_U141 , P3_PHYADDRPOINTER_REG_2_ , P3_ADD_339_U4 );
nand NAND2_20828 ( P3_ADD_339_U142 , P3_PHYADDRPOINTER_REG_1_ , P3_ADD_339_U5 );
nand NAND2_20829 ( P3_ADD_339_U143 , P3_PHYADDRPOINTER_REG_29_ , P3_ADD_339_U58 );
nand NAND2_20830 ( P3_ADD_339_U144 , P3_ADD_339_U120 , P3_ADD_339_U59 );
nand NAND2_20831 ( P3_ADD_339_U145 , P3_PHYADDRPOINTER_REG_28_ , P3_ADD_339_U56 );
nand NAND2_20832 ( P3_ADD_339_U146 , P3_ADD_339_U119 , P3_ADD_339_U57 );
nand NAND2_20833 ( P3_ADD_339_U147 , P3_PHYADDRPOINTER_REG_27_ , P3_ADD_339_U54 );
nand NAND2_20834 ( P3_ADD_339_U148 , P3_ADD_339_U118 , P3_ADD_339_U55 );
nand NAND2_20835 ( P3_ADD_339_U149 , P3_PHYADDRPOINTER_REG_26_ , P3_ADD_339_U52 );
nand NAND2_20836 ( P3_ADD_339_U150 , P3_ADD_339_U117 , P3_ADD_339_U53 );
nand NAND2_20837 ( P3_ADD_339_U151 , P3_PHYADDRPOINTER_REG_25_ , P3_ADD_339_U50 );
nand NAND2_20838 ( P3_ADD_339_U152 , P3_ADD_339_U116 , P3_ADD_339_U51 );
nand NAND2_20839 ( P3_ADD_339_U153 , P3_PHYADDRPOINTER_REG_24_ , P3_ADD_339_U48 );
nand NAND2_20840 ( P3_ADD_339_U154 , P3_ADD_339_U115 , P3_ADD_339_U49 );
nand NAND2_20841 ( P3_ADD_339_U155 , P3_PHYADDRPOINTER_REG_23_ , P3_ADD_339_U46 );
nand NAND2_20842 ( P3_ADD_339_U156 , P3_ADD_339_U114 , P3_ADD_339_U47 );
nand NAND2_20843 ( P3_ADD_339_U157 , P3_PHYADDRPOINTER_REG_22_ , P3_ADD_339_U44 );
nand NAND2_20844 ( P3_ADD_339_U158 , P3_ADD_339_U113 , P3_ADD_339_U45 );
nand NAND2_20845 ( P3_ADD_339_U159 , P3_PHYADDRPOINTER_REG_21_ , P3_ADD_339_U42 );
nand NAND2_20846 ( P3_ADD_339_U160 , P3_ADD_339_U112 , P3_ADD_339_U43 );
nand NAND2_20847 ( P3_ADD_339_U161 , P3_PHYADDRPOINTER_REG_20_ , P3_ADD_339_U40 );
nand NAND2_20848 ( P3_ADD_339_U162 , P3_ADD_339_U111 , P3_ADD_339_U41 );
nand NAND2_20849 ( P3_ADD_339_U163 , P3_PHYADDRPOINTER_REG_19_ , P3_ADD_339_U38 );
nand NAND2_20850 ( P3_ADD_339_U164 , P3_ADD_339_U110 , P3_ADD_339_U39 );
nand NAND2_20851 ( P3_ADD_339_U165 , P3_PHYADDRPOINTER_REG_18_ , P3_ADD_339_U36 );
nand NAND2_20852 ( P3_ADD_339_U166 , P3_ADD_339_U109 , P3_ADD_339_U37 );
nand NAND2_20853 ( P3_ADD_339_U167 , P3_PHYADDRPOINTER_REG_17_ , P3_ADD_339_U34 );
nand NAND2_20854 ( P3_ADD_339_U168 , P3_ADD_339_U108 , P3_ADD_339_U35 );
nand NAND2_20855 ( P3_ADD_339_U169 , P3_PHYADDRPOINTER_REG_16_ , P3_ADD_339_U32 );
nand NAND2_20856 ( P3_ADD_339_U170 , P3_ADD_339_U107 , P3_ADD_339_U33 );
nand NAND2_20857 ( P3_ADD_339_U171 , P3_PHYADDRPOINTER_REG_15_ , P3_ADD_339_U30 );
nand NAND2_20858 ( P3_ADD_339_U172 , P3_ADD_339_U106 , P3_ADD_339_U31 );
nand NAND2_20859 ( P3_ADD_339_U173 , P3_PHYADDRPOINTER_REG_14_ , P3_ADD_339_U28 );
nand NAND2_20860 ( P3_ADD_339_U174 , P3_ADD_339_U105 , P3_ADD_339_U29 );
nand NAND2_20861 ( P3_ADD_339_U175 , P3_PHYADDRPOINTER_REG_13_ , P3_ADD_339_U26 );
nand NAND2_20862 ( P3_ADD_339_U176 , P3_ADD_339_U104 , P3_ADD_339_U27 );
nand NAND2_20863 ( P3_ADD_339_U177 , P3_PHYADDRPOINTER_REG_12_ , P3_ADD_339_U24 );
nand NAND2_20864 ( P3_ADD_339_U178 , P3_ADD_339_U103 , P3_ADD_339_U25 );
nand NAND2_20865 ( P3_ADD_339_U179 , P3_PHYADDRPOINTER_REG_11_ , P3_ADD_339_U22 );
nand NAND2_20866 ( P3_ADD_339_U180 , P3_ADD_339_U102 , P3_ADD_339_U23 );
nand NAND2_20867 ( P3_ADD_339_U181 , P3_PHYADDRPOINTER_REG_10_ , P3_ADD_339_U20 );
nand NAND2_20868 ( P3_ADD_339_U182 , P3_ADD_339_U101 , P3_ADD_339_U21 );
not NOT1_20869 ( P3_ADD_360_U4 , P3_U2622 );
and AND2_20870 ( P3_ADD_360_U5 , P3_ADD_360_U22 , P3_ADD_360_U27 );
not NOT1_20871 ( P3_ADD_360_U6 , P3_U2623 );
nand NAND2_20872 ( P3_ADD_360_U7 , P3_U2623 , P3_U2622 );
not NOT1_20873 ( P3_ADD_360_U8 , P3_U2624 );
nand NAND2_20874 ( P3_ADD_360_U9 , P3_U2624 , P3_ADD_360_U24 );
not NOT1_20875 ( P3_ADD_360_U10 , P3_U2625 );
nand NAND2_20876 ( P3_ADD_360_U11 , P3_U2625 , P3_ADD_360_U25 );
not NOT1_20877 ( P3_ADD_360_U12 , P3_U2626 );
nand NAND2_20878 ( P3_ADD_360_U13 , P3_U2626 , P3_ADD_360_U26 );
not NOT1_20879 ( P3_ADD_360_U14 , P3_U2628 );
not NOT1_20880 ( P3_ADD_360_U15 , P3_U2627 );
nand NAND2_20881 ( P3_ADD_360_U16 , P3_ADD_360_U30 , P3_ADD_360_U29 );
nand NAND2_20882 ( P3_ADD_360_U17 , P3_ADD_360_U32 , P3_ADD_360_U31 );
nand NAND2_20883 ( P3_ADD_360_U18 , P3_ADD_360_U34 , P3_ADD_360_U33 );
nand NAND2_20884 ( P3_ADD_360_U19 , P3_ADD_360_U36 , P3_ADD_360_U35 );
nand NAND2_20885 ( P3_ADD_360_U20 , P3_ADD_360_U38 , P3_ADD_360_U37 );
nand NAND2_20886 ( P3_ADD_360_U21 , P3_ADD_360_U40 , P3_ADD_360_U39 );
and AND2_20887 ( P3_ADD_360_U22 , P3_U2628 , P3_U2627 );
nand NAND2_20888 ( P3_ADD_360_U23 , P3_U2627 , P3_ADD_360_U27 );
not NOT1_20889 ( P3_ADD_360_U24 , P3_ADD_360_U7 );
not NOT1_20890 ( P3_ADD_360_U25 , P3_ADD_360_U9 );
not NOT1_20891 ( P3_ADD_360_U26 , P3_ADD_360_U11 );
not NOT1_20892 ( P3_ADD_360_U27 , P3_ADD_360_U13 );
not NOT1_20893 ( P3_ADD_360_U28 , P3_ADD_360_U23 );
nand NAND2_20894 ( P3_ADD_360_U29 , P3_U2628 , P3_ADD_360_U23 );
nand NAND2_20895 ( P3_ADD_360_U30 , P3_ADD_360_U28 , P3_ADD_360_U14 );
nand NAND2_20896 ( P3_ADD_360_U31 , P3_U2627 , P3_ADD_360_U13 );
nand NAND2_20897 ( P3_ADD_360_U32 , P3_ADD_360_U27 , P3_ADD_360_U15 );
nand NAND2_20898 ( P3_ADD_360_U33 , P3_U2626 , P3_ADD_360_U11 );
nand NAND2_20899 ( P3_ADD_360_U34 , P3_ADD_360_U26 , P3_ADD_360_U12 );
nand NAND2_20900 ( P3_ADD_360_U35 , P3_U2625 , P3_ADD_360_U9 );
nand NAND2_20901 ( P3_ADD_360_U36 , P3_ADD_360_U25 , P3_ADD_360_U10 );
nand NAND2_20902 ( P3_ADD_360_U37 , P3_U2624 , P3_ADD_360_U7 );
nand NAND2_20903 ( P3_ADD_360_U38 , P3_ADD_360_U24 , P3_ADD_360_U8 );
nand NAND2_20904 ( P3_ADD_360_U39 , P3_U2623 , P3_ADD_360_U4 );
nand NAND2_20905 ( P3_ADD_360_U40 , P3_U2622 , P3_ADD_360_U6 );
not NOT1_20906 ( P3_LTE_597_U6 , P3_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_20907 ( P3_SUB_580_U6 , P3_SUB_580_U10 , P3_SUB_580_U9 );
not NOT1_20908 ( P3_SUB_580_U7 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_20909 ( P3_SUB_580_U8 , P3_INSTADDRPOINTER_REG_0_ );
nand NAND2_20910 ( P3_SUB_580_U9 , P3_INSTADDRPOINTER_REG_1_ , P3_SUB_580_U8 );
nand NAND2_20911 ( P3_SUB_580_U10 , P3_INSTADDRPOINTER_REG_0_ , P3_SUB_580_U7 );
or OR2_20912 ( P3_LT_589_U6 , P3_LT_589_U8 , P3_U2629 );
and AND2_20913 ( P3_LT_589_U7 , P3_SUB_589_U7 , P3_SUB_589_U6 );
nor nor_20914 ( P3_LT_589_U8 , P3_LT_589_U7 , P3_SUB_589_U8 , P3_SUB_589_U9 );
not NOT1_20915 ( P3_ADD_541_U4 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_20916 ( P3_ADD_541_U5 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_20917 ( P3_ADD_541_U6 , P3_INSTADDRPOINTER_REG_2_ , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_20918 ( P3_ADD_541_U7 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_20919 ( P3_ADD_541_U8 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_541_U94 );
not NOT1_20920 ( P3_ADD_541_U9 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_20921 ( P3_ADD_541_U10 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_541_U95 );
not NOT1_20922 ( P3_ADD_541_U11 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_20923 ( P3_ADD_541_U12 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_541_U96 );
not NOT1_20924 ( P3_ADD_541_U13 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_20925 ( P3_ADD_541_U14 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_541_U97 );
not NOT1_20926 ( P3_ADD_541_U15 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_20927 ( P3_ADD_541_U16 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_541_U98 );
not NOT1_20928 ( P3_ADD_541_U17 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_20929 ( P3_ADD_541_U18 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_20930 ( P3_ADD_541_U19 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_541_U99 );
nand NAND2_20931 ( P3_ADD_541_U20 , P3_ADD_541_U100 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_20932 ( P3_ADD_541_U21 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_20933 ( P3_ADD_541_U22 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_541_U101 );
not NOT1_20934 ( P3_ADD_541_U23 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_20935 ( P3_ADD_541_U24 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_541_U102 );
not NOT1_20936 ( P3_ADD_541_U25 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_20937 ( P3_ADD_541_U26 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_541_U103 );
not NOT1_20938 ( P3_ADD_541_U27 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_20939 ( P3_ADD_541_U28 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_541_U104 );
not NOT1_20940 ( P3_ADD_541_U29 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_20941 ( P3_ADD_541_U30 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_541_U105 );
not NOT1_20942 ( P3_ADD_541_U31 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_20943 ( P3_ADD_541_U32 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_541_U106 );
not NOT1_20944 ( P3_ADD_541_U33 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_20945 ( P3_ADD_541_U34 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_541_U107 );
not NOT1_20946 ( P3_ADD_541_U35 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_20947 ( P3_ADD_541_U36 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_541_U108 );
not NOT1_20948 ( P3_ADD_541_U37 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_20949 ( P3_ADD_541_U38 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_541_U109 );
not NOT1_20950 ( P3_ADD_541_U39 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_20951 ( P3_ADD_541_U40 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_541_U110 );
not NOT1_20952 ( P3_ADD_541_U41 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_20953 ( P3_ADD_541_U42 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_541_U111 );
not NOT1_20954 ( P3_ADD_541_U43 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_20955 ( P3_ADD_541_U44 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_541_U112 );
not NOT1_20956 ( P3_ADD_541_U45 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_20957 ( P3_ADD_541_U46 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_541_U113 );
not NOT1_20958 ( P3_ADD_541_U47 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_20959 ( P3_ADD_541_U48 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_541_U114 );
not NOT1_20960 ( P3_ADD_541_U49 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_20961 ( P3_ADD_541_U50 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_541_U115 );
not NOT1_20962 ( P3_ADD_541_U51 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_20963 ( P3_ADD_541_U52 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_541_U116 );
not NOT1_20964 ( P3_ADD_541_U53 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_20965 ( P3_ADD_541_U54 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_541_U117 );
not NOT1_20966 ( P3_ADD_541_U55 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_20967 ( P3_ADD_541_U56 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_541_U118 );
not NOT1_20968 ( P3_ADD_541_U57 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_20969 ( P3_ADD_541_U58 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_541_U119 );
not NOT1_20970 ( P3_ADD_541_U59 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_20971 ( P3_ADD_541_U60 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_541_U120 );
not NOT1_20972 ( P3_ADD_541_U61 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_20973 ( P3_ADD_541_U62 , P3_ADD_541_U124 , P3_ADD_541_U123 );
nand NAND2_20974 ( P3_ADD_541_U63 , P3_ADD_541_U126 , P3_ADD_541_U125 );
nand NAND2_20975 ( P3_ADD_541_U64 , P3_ADD_541_U128 , P3_ADD_541_U127 );
nand NAND2_20976 ( P3_ADD_541_U65 , P3_ADD_541_U130 , P3_ADD_541_U129 );
nand NAND2_20977 ( P3_ADD_541_U66 , P3_ADD_541_U132 , P3_ADD_541_U131 );
nand NAND2_20978 ( P3_ADD_541_U67 , P3_ADD_541_U134 , P3_ADD_541_U133 );
nand NAND2_20979 ( P3_ADD_541_U68 , P3_ADD_541_U136 , P3_ADD_541_U135 );
nand NAND2_20980 ( P3_ADD_541_U69 , P3_ADD_541_U138 , P3_ADD_541_U137 );
nand NAND2_20981 ( P3_ADD_541_U70 , P3_ADD_541_U140 , P3_ADD_541_U139 );
nand NAND2_20982 ( P3_ADD_541_U71 , P3_ADD_541_U142 , P3_ADD_541_U141 );
nand NAND2_20983 ( P3_ADD_541_U72 , P3_ADD_541_U144 , P3_ADD_541_U143 );
nand NAND2_20984 ( P3_ADD_541_U73 , P3_ADD_541_U146 , P3_ADD_541_U145 );
nand NAND2_20985 ( P3_ADD_541_U74 , P3_ADD_541_U148 , P3_ADD_541_U147 );
nand NAND2_20986 ( P3_ADD_541_U75 , P3_ADD_541_U150 , P3_ADD_541_U149 );
nand NAND2_20987 ( P3_ADD_541_U76 , P3_ADD_541_U152 , P3_ADD_541_U151 );
nand NAND2_20988 ( P3_ADD_541_U77 , P3_ADD_541_U154 , P3_ADD_541_U153 );
nand NAND2_20989 ( P3_ADD_541_U78 , P3_ADD_541_U156 , P3_ADD_541_U155 );
nand NAND2_20990 ( P3_ADD_541_U79 , P3_ADD_541_U158 , P3_ADD_541_U157 );
nand NAND2_20991 ( P3_ADD_541_U80 , P3_ADD_541_U160 , P3_ADD_541_U159 );
nand NAND2_20992 ( P3_ADD_541_U81 , P3_ADD_541_U162 , P3_ADD_541_U161 );
nand NAND2_20993 ( P3_ADD_541_U82 , P3_ADD_541_U164 , P3_ADD_541_U163 );
nand NAND2_20994 ( P3_ADD_541_U83 , P3_ADD_541_U166 , P3_ADD_541_U165 );
nand NAND2_20995 ( P3_ADD_541_U84 , P3_ADD_541_U168 , P3_ADD_541_U167 );
nand NAND2_20996 ( P3_ADD_541_U85 , P3_ADD_541_U170 , P3_ADD_541_U169 );
nand NAND2_20997 ( P3_ADD_541_U86 , P3_ADD_541_U172 , P3_ADD_541_U171 );
nand NAND2_20998 ( P3_ADD_541_U87 , P3_ADD_541_U174 , P3_ADD_541_U173 );
nand NAND2_20999 ( P3_ADD_541_U88 , P3_ADD_541_U176 , P3_ADD_541_U175 );
nand NAND2_21000 ( P3_ADD_541_U89 , P3_ADD_541_U178 , P3_ADD_541_U177 );
nand NAND2_21001 ( P3_ADD_541_U90 , P3_ADD_541_U180 , P3_ADD_541_U179 );
nand NAND2_21002 ( P3_ADD_541_U91 , P3_ADD_541_U182 , P3_ADD_541_U181 );
not NOT1_21003 ( P3_ADD_541_U92 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_21004 ( P3_ADD_541_U93 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_541_U121 );
not NOT1_21005 ( P3_ADD_541_U94 , P3_ADD_541_U6 );
not NOT1_21006 ( P3_ADD_541_U95 , P3_ADD_541_U8 );
not NOT1_21007 ( P3_ADD_541_U96 , P3_ADD_541_U10 );
not NOT1_21008 ( P3_ADD_541_U97 , P3_ADD_541_U12 );
not NOT1_21009 ( P3_ADD_541_U98 , P3_ADD_541_U14 );
not NOT1_21010 ( P3_ADD_541_U99 , P3_ADD_541_U16 );
not NOT1_21011 ( P3_ADD_541_U100 , P3_ADD_541_U19 );
not NOT1_21012 ( P3_ADD_541_U101 , P3_ADD_541_U20 );
not NOT1_21013 ( P3_ADD_541_U102 , P3_ADD_541_U22 );
not NOT1_21014 ( P3_ADD_541_U103 , P3_ADD_541_U24 );
not NOT1_21015 ( P3_ADD_541_U104 , P3_ADD_541_U26 );
not NOT1_21016 ( P3_ADD_541_U105 , P3_ADD_541_U28 );
not NOT1_21017 ( P3_ADD_541_U106 , P3_ADD_541_U30 );
not NOT1_21018 ( P3_ADD_541_U107 , P3_ADD_541_U32 );
not NOT1_21019 ( P3_ADD_541_U108 , P3_ADD_541_U34 );
not NOT1_21020 ( P3_ADD_541_U109 , P3_ADD_541_U36 );
not NOT1_21021 ( P3_ADD_541_U110 , P3_ADD_541_U38 );
not NOT1_21022 ( P3_ADD_541_U111 , P3_ADD_541_U40 );
not NOT1_21023 ( P3_ADD_541_U112 , P3_ADD_541_U42 );
not NOT1_21024 ( P3_ADD_541_U113 , P3_ADD_541_U44 );
not NOT1_21025 ( P3_ADD_541_U114 , P3_ADD_541_U46 );
not NOT1_21026 ( P3_ADD_541_U115 , P3_ADD_541_U48 );
not NOT1_21027 ( P3_ADD_541_U116 , P3_ADD_541_U50 );
not NOT1_21028 ( P3_ADD_541_U117 , P3_ADD_541_U52 );
not NOT1_21029 ( P3_ADD_541_U118 , P3_ADD_541_U54 );
not NOT1_21030 ( P3_ADD_541_U119 , P3_ADD_541_U56 );
not NOT1_21031 ( P3_ADD_541_U120 , P3_ADD_541_U58 );
not NOT1_21032 ( P3_ADD_541_U121 , P3_ADD_541_U60 );
not NOT1_21033 ( P3_ADD_541_U122 , P3_ADD_541_U93 );
nand NAND2_21034 ( P3_ADD_541_U123 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_541_U19 );
nand NAND2_21035 ( P3_ADD_541_U124 , P3_ADD_541_U100 , P3_ADD_541_U18 );
nand NAND2_21036 ( P3_ADD_541_U125 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_541_U16 );
nand NAND2_21037 ( P3_ADD_541_U126 , P3_ADD_541_U99 , P3_ADD_541_U17 );
nand NAND2_21038 ( P3_ADD_541_U127 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_541_U14 );
nand NAND2_21039 ( P3_ADD_541_U128 , P3_ADD_541_U98 , P3_ADD_541_U15 );
nand NAND2_21040 ( P3_ADD_541_U129 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_541_U12 );
nand NAND2_21041 ( P3_ADD_541_U130 , P3_ADD_541_U97 , P3_ADD_541_U13 );
nand NAND2_21042 ( P3_ADD_541_U131 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_541_U10 );
nand NAND2_21043 ( P3_ADD_541_U132 , P3_ADD_541_U96 , P3_ADD_541_U11 );
nand NAND2_21044 ( P3_ADD_541_U133 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_541_U8 );
nand NAND2_21045 ( P3_ADD_541_U134 , P3_ADD_541_U95 , P3_ADD_541_U9 );
nand NAND2_21046 ( P3_ADD_541_U135 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_541_U6 );
nand NAND2_21047 ( P3_ADD_541_U136 , P3_ADD_541_U94 , P3_ADD_541_U7 );
nand NAND2_21048 ( P3_ADD_541_U137 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_541_U93 );
nand NAND2_21049 ( P3_ADD_541_U138 , P3_ADD_541_U122 , P3_ADD_541_U92 );
nand NAND2_21050 ( P3_ADD_541_U139 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_541_U60 );
nand NAND2_21051 ( P3_ADD_541_U140 , P3_ADD_541_U121 , P3_ADD_541_U61 );
nand NAND2_21052 ( P3_ADD_541_U141 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_541_U4 );
nand NAND2_21053 ( P3_ADD_541_U142 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_541_U5 );
nand NAND2_21054 ( P3_ADD_541_U143 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_541_U58 );
nand NAND2_21055 ( P3_ADD_541_U144 , P3_ADD_541_U120 , P3_ADD_541_U59 );
nand NAND2_21056 ( P3_ADD_541_U145 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_541_U56 );
nand NAND2_21057 ( P3_ADD_541_U146 , P3_ADD_541_U119 , P3_ADD_541_U57 );
nand NAND2_21058 ( P3_ADD_541_U147 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_541_U54 );
nand NAND2_21059 ( P3_ADD_541_U148 , P3_ADD_541_U118 , P3_ADD_541_U55 );
nand NAND2_21060 ( P3_ADD_541_U149 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_541_U52 );
nand NAND2_21061 ( P3_ADD_541_U150 , P3_ADD_541_U117 , P3_ADD_541_U53 );
nand NAND2_21062 ( P3_ADD_541_U151 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_541_U50 );
nand NAND2_21063 ( P3_ADD_541_U152 , P3_ADD_541_U116 , P3_ADD_541_U51 );
nand NAND2_21064 ( P3_ADD_541_U153 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_541_U48 );
nand NAND2_21065 ( P3_ADD_541_U154 , P3_ADD_541_U115 , P3_ADD_541_U49 );
nand NAND2_21066 ( P3_ADD_541_U155 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_541_U46 );
nand NAND2_21067 ( P3_ADD_541_U156 , P3_ADD_541_U114 , P3_ADD_541_U47 );
nand NAND2_21068 ( P3_ADD_541_U157 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_541_U44 );
nand NAND2_21069 ( P3_ADD_541_U158 , P3_ADD_541_U113 , P3_ADD_541_U45 );
nand NAND2_21070 ( P3_ADD_541_U159 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_541_U42 );
nand NAND2_21071 ( P3_ADD_541_U160 , P3_ADD_541_U112 , P3_ADD_541_U43 );
nand NAND2_21072 ( P3_ADD_541_U161 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_541_U40 );
nand NAND2_21073 ( P3_ADD_541_U162 , P3_ADD_541_U111 , P3_ADD_541_U41 );
nand NAND2_21074 ( P3_ADD_541_U163 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_541_U38 );
nand NAND2_21075 ( P3_ADD_541_U164 , P3_ADD_541_U110 , P3_ADD_541_U39 );
nand NAND2_21076 ( P3_ADD_541_U165 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_541_U36 );
nand NAND2_21077 ( P3_ADD_541_U166 , P3_ADD_541_U109 , P3_ADD_541_U37 );
nand NAND2_21078 ( P3_ADD_541_U167 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_541_U34 );
nand NAND2_21079 ( P3_ADD_541_U168 , P3_ADD_541_U108 , P3_ADD_541_U35 );
nand NAND2_21080 ( P3_ADD_541_U169 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_541_U32 );
nand NAND2_21081 ( P3_ADD_541_U170 , P3_ADD_541_U107 , P3_ADD_541_U33 );
nand NAND2_21082 ( P3_ADD_541_U171 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_541_U30 );
nand NAND2_21083 ( P3_ADD_541_U172 , P3_ADD_541_U106 , P3_ADD_541_U31 );
nand NAND2_21084 ( P3_ADD_541_U173 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_541_U28 );
nand NAND2_21085 ( P3_ADD_541_U174 , P3_ADD_541_U105 , P3_ADD_541_U29 );
nand NAND2_21086 ( P3_ADD_541_U175 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_541_U26 );
nand NAND2_21087 ( P3_ADD_541_U176 , P3_ADD_541_U104 , P3_ADD_541_U27 );
nand NAND2_21088 ( P3_ADD_541_U177 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_541_U24 );
nand NAND2_21089 ( P3_ADD_541_U178 , P3_ADD_541_U103 , P3_ADD_541_U25 );
nand NAND2_21090 ( P3_ADD_541_U179 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_541_U22 );
nand NAND2_21091 ( P3_ADD_541_U180 , P3_ADD_541_U102 , P3_ADD_541_U23 );
nand NAND2_21092 ( P3_ADD_541_U181 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_541_U20 );
nand NAND2_21093 ( P3_ADD_541_U182 , P3_ADD_541_U101 , P3_ADD_541_U21 );
nand NAND2_21094 ( P3_SUB_355_U6 , P3_SUB_355_U45 , P3_SUB_355_U44 );
nand NAND2_21095 ( P3_SUB_355_U7 , P3_SUB_355_U9 , P3_SUB_355_U46 );
not NOT1_21096 ( P3_SUB_355_U8 , P3_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_21097 ( P3_SUB_355_U9 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_SUB_355_U18 );
not NOT1_21098 ( P3_SUB_355_U10 , P3_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_21099 ( P3_SUB_355_U11 , P3_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_21100 ( P3_SUB_355_U12 , P3_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_21101 ( P3_SUB_355_U13 , P3_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_21102 ( P3_SUB_355_U14 , P3_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_21103 ( P3_SUB_355_U15 , P3_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_21104 ( P3_SUB_355_U16 , P3_SUB_355_U41 , P3_SUB_355_U40 );
not NOT1_21105 ( P3_SUB_355_U17 , P3_INSTQUEUERD_ADDR_REG_4_ );
not NOT1_21106 ( P3_SUB_355_U18 , P3_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_21107 ( P3_SUB_355_U19 , P3_SUB_355_U51 , P3_SUB_355_U50 );
nand NAND2_21108 ( P3_SUB_355_U20 , P3_SUB_355_U56 , P3_SUB_355_U55 );
nand NAND2_21109 ( P3_SUB_355_U21 , P3_SUB_355_U61 , P3_SUB_355_U60 );
nand NAND2_21110 ( P3_SUB_355_U22 , P3_SUB_355_U66 , P3_SUB_355_U65 );
nand NAND2_21111 ( P3_SUB_355_U23 , P3_SUB_355_U48 , P3_SUB_355_U47 );
nand NAND2_21112 ( P3_SUB_355_U24 , P3_SUB_355_U53 , P3_SUB_355_U52 );
nand NAND2_21113 ( P3_SUB_355_U25 , P3_SUB_355_U58 , P3_SUB_355_U57 );
nand NAND2_21114 ( P3_SUB_355_U26 , P3_SUB_355_U63 , P3_SUB_355_U62 );
nand NAND2_21115 ( P3_SUB_355_U27 , P3_SUB_355_U37 , P3_SUB_355_U36 );
nand NAND2_21116 ( P3_SUB_355_U28 , P3_SUB_355_U33 , P3_SUB_355_U32 );
not NOT1_21117 ( P3_SUB_355_U29 , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_21118 ( P3_SUB_355_U30 , P3_SUB_355_U9 );
nand NAND2_21119 ( P3_SUB_355_U31 , P3_SUB_355_U30 , P3_SUB_355_U10 );
nand NAND2_21120 ( P3_SUB_355_U32 , P3_SUB_355_U31 , P3_SUB_355_U29 );
nand NAND2_21121 ( P3_SUB_355_U33 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_355_U9 );
not NOT1_21122 ( P3_SUB_355_U34 , P3_SUB_355_U28 );
nand NAND2_21123 ( P3_SUB_355_U35 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_355_U12 );
nand NAND2_21124 ( P3_SUB_355_U36 , P3_SUB_355_U35 , P3_SUB_355_U28 );
nand NAND2_21125 ( P3_SUB_355_U37 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_355_U11 );
not NOT1_21126 ( P3_SUB_355_U38 , P3_SUB_355_U27 );
nand NAND2_21127 ( P3_SUB_355_U39 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_355_U14 );
nand NAND2_21128 ( P3_SUB_355_U40 , P3_SUB_355_U39 , P3_SUB_355_U27 );
nand NAND2_21129 ( P3_SUB_355_U41 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_355_U13 );
not NOT1_21130 ( P3_SUB_355_U42 , P3_SUB_355_U16 );
nand NAND2_21131 ( P3_SUB_355_U43 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_355_U17 );
nand NAND2_21132 ( P3_SUB_355_U44 , P3_SUB_355_U42 , P3_SUB_355_U43 );
nand NAND2_21133 ( P3_SUB_355_U45 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_355_U15 );
nand NAND2_21134 ( P3_SUB_355_U46 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_SUB_355_U8 );
nand NAND2_21135 ( P3_SUB_355_U47 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_355_U15 );
nand NAND2_21136 ( P3_SUB_355_U48 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_355_U17 );
not NOT1_21137 ( P3_SUB_355_U49 , P3_SUB_355_U23 );
nand NAND2_21138 ( P3_SUB_355_U50 , P3_SUB_355_U49 , P3_SUB_355_U42 );
nand NAND2_21139 ( P3_SUB_355_U51 , P3_SUB_355_U23 , P3_SUB_355_U16 );
nand NAND2_21140 ( P3_SUB_355_U52 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_355_U14 );
nand NAND2_21141 ( P3_SUB_355_U53 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_355_U13 );
not NOT1_21142 ( P3_SUB_355_U54 , P3_SUB_355_U24 );
nand NAND2_21143 ( P3_SUB_355_U55 , P3_SUB_355_U38 , P3_SUB_355_U54 );
nand NAND2_21144 ( P3_SUB_355_U56 , P3_SUB_355_U24 , P3_SUB_355_U27 );
nand NAND2_21145 ( P3_SUB_355_U57 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_355_U12 );
nand NAND2_21146 ( P3_SUB_355_U58 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_355_U11 );
not NOT1_21147 ( P3_SUB_355_U59 , P3_SUB_355_U25 );
nand NAND2_21148 ( P3_SUB_355_U60 , P3_SUB_355_U34 , P3_SUB_355_U59 );
nand NAND2_21149 ( P3_SUB_355_U61 , P3_SUB_355_U25 , P3_SUB_355_U28 );
nand NAND2_21150 ( P3_SUB_355_U62 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_SUB_355_U10 );
nand NAND2_21151 ( P3_SUB_355_U63 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_355_U29 );
not NOT1_21152 ( P3_SUB_355_U64 , P3_SUB_355_U26 );
nand NAND2_21153 ( P3_SUB_355_U65 , P3_SUB_355_U64 , P3_SUB_355_U30 );
nand NAND2_21154 ( P3_SUB_355_U66 , P3_SUB_355_U26 , P3_SUB_355_U9 );
nand NAND2_21155 ( P3_SUB_450_U6 , P3_SUB_450_U43 , P3_SUB_450_U42 );
nand NAND2_21156 ( P3_SUB_450_U7 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_SUB_450_U27 );
not NOT1_21157 ( P3_SUB_450_U8 , P3_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_21158 ( P3_SUB_450_U9 , P3_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_21159 ( P3_SUB_450_U10 , P3_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_21160 ( P3_SUB_450_U11 , P3_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_21161 ( P3_SUB_450_U12 , P3_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_21162 ( P3_SUB_450_U13 , P3_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_21163 ( P3_SUB_450_U14 , P3_SUB_450_U39 , P3_SUB_450_U38 );
not NOT1_21164 ( P3_SUB_450_U15 , P3_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_21165 ( P3_SUB_450_U16 , P3_SUB_450_U48 , P3_SUB_450_U47 );
nand NAND2_21166 ( P3_SUB_450_U17 , P3_SUB_450_U53 , P3_SUB_450_U52 );
nand NAND2_21167 ( P3_SUB_450_U18 , P3_SUB_450_U58 , P3_SUB_450_U57 );
nand NAND2_21168 ( P3_SUB_450_U19 , P3_SUB_450_U63 , P3_SUB_450_U62 );
nand NAND2_21169 ( P3_SUB_450_U20 , P3_SUB_450_U45 , P3_SUB_450_U44 );
nand NAND2_21170 ( P3_SUB_450_U21 , P3_SUB_450_U50 , P3_SUB_450_U49 );
nand NAND2_21171 ( P3_SUB_450_U22 , P3_SUB_450_U55 , P3_SUB_450_U54 );
nand NAND2_21172 ( P3_SUB_450_U23 , P3_SUB_450_U60 , P3_SUB_450_U59 );
nand NAND2_21173 ( P3_SUB_450_U24 , P3_SUB_450_U35 , P3_SUB_450_U34 );
nand NAND2_21174 ( P3_SUB_450_U25 , P3_SUB_450_U31 , P3_SUB_450_U30 );
not NOT1_21175 ( P3_SUB_450_U26 , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_21176 ( P3_SUB_450_U27 , P3_INSTQUEUEWR_ADDR_REG_0_ );
not NOT1_21177 ( P3_SUB_450_U28 , P3_SUB_450_U7 );
nand NAND2_21178 ( P3_SUB_450_U29 , P3_SUB_450_U28 , P3_SUB_450_U8 );
nand NAND2_21179 ( P3_SUB_450_U30 , P3_SUB_450_U29 , P3_SUB_450_U26 );
nand NAND2_21180 ( P3_SUB_450_U31 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_450_U7 );
not NOT1_21181 ( P3_SUB_450_U32 , P3_SUB_450_U25 );
nand NAND2_21182 ( P3_SUB_450_U33 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_450_U10 );
nand NAND2_21183 ( P3_SUB_450_U34 , P3_SUB_450_U33 , P3_SUB_450_U25 );
nand NAND2_21184 ( P3_SUB_450_U35 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_450_U9 );
not NOT1_21185 ( P3_SUB_450_U36 , P3_SUB_450_U24 );
nand NAND2_21186 ( P3_SUB_450_U37 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_450_U12 );
nand NAND2_21187 ( P3_SUB_450_U38 , P3_SUB_450_U37 , P3_SUB_450_U24 );
nand NAND2_21188 ( P3_SUB_450_U39 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_450_U11 );
not NOT1_21189 ( P3_SUB_450_U40 , P3_SUB_450_U14 );
nand NAND2_21190 ( P3_SUB_450_U41 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_450_U15 );
nand NAND2_21191 ( P3_SUB_450_U42 , P3_SUB_450_U40 , P3_SUB_450_U41 );
nand NAND2_21192 ( P3_SUB_450_U43 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_450_U13 );
nand NAND2_21193 ( P3_SUB_450_U44 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_450_U13 );
nand NAND2_21194 ( P3_SUB_450_U45 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_450_U15 );
not NOT1_21195 ( P3_SUB_450_U46 , P3_SUB_450_U20 );
nand NAND2_21196 ( P3_SUB_450_U47 , P3_SUB_450_U46 , P3_SUB_450_U40 );
nand NAND2_21197 ( P3_SUB_450_U48 , P3_SUB_450_U20 , P3_SUB_450_U14 );
nand NAND2_21198 ( P3_SUB_450_U49 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_450_U12 );
nand NAND2_21199 ( P3_SUB_450_U50 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_450_U11 );
not NOT1_21200 ( P3_SUB_450_U51 , P3_SUB_450_U21 );
nand NAND2_21201 ( P3_SUB_450_U52 , P3_SUB_450_U36 , P3_SUB_450_U51 );
nand NAND2_21202 ( P3_SUB_450_U53 , P3_SUB_450_U21 , P3_SUB_450_U24 );
nand NAND2_21203 ( P3_SUB_450_U54 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_450_U10 );
nand NAND2_21204 ( P3_SUB_450_U55 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_450_U9 );
not NOT1_21205 ( P3_SUB_450_U56 , P3_SUB_450_U22 );
nand NAND2_21206 ( P3_SUB_450_U57 , P3_SUB_450_U32 , P3_SUB_450_U56 );
nand NAND2_21207 ( P3_SUB_450_U58 , P3_SUB_450_U22 , P3_SUB_450_U25 );
nand NAND2_21208 ( P3_SUB_450_U59 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_SUB_450_U8 );
nand NAND2_21209 ( P3_SUB_450_U60 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_450_U26 );
not NOT1_21210 ( P3_SUB_450_U61 , P3_SUB_450_U23 );
nand NAND2_21211 ( P3_SUB_450_U62 , P3_SUB_450_U61 , P3_SUB_450_U28 );
nand NAND2_21212 ( P3_SUB_450_U63 , P3_SUB_450_U23 , P3_SUB_450_U7 );
and AND2_21213 ( P3_SUB_357_1258_U4 , P3_INSTADDRPOINTER_REG_27_ , P3_INSTADDRPOINTER_REG_28_ );
and AND2_21214 ( P3_SUB_357_1258_U5 , P3_SUB_357_1258_U188 , P3_SUB_357_1258_U186 );
and AND2_21215 ( P3_SUB_357_1258_U6 , P3_SUB_357_1258_U187 , P3_SUB_357_1258_U178 );
and AND2_21216 ( P3_SUB_357_1258_U7 , P3_SUB_357_1258_U6 , P3_SUB_357_1258_U189 );
and AND2_21217 ( P3_SUB_357_1258_U8 , P3_SUB_357_1258_U5 , P3_SUB_357_1258_U190 );
and AND2_21218 ( P3_SUB_357_1258_U9 , P3_SUB_357_1258_U209 , P3_SUB_357_1258_U204 );
and AND4_21219 ( P3_SUB_357_1258_U10 , P3_SUB_357_1258_U210 , P3_SUB_357_1258_U205 , P3_SUB_357_1258_U206 , P3_SUB_357_1258_U156 );
and AND2_21220 ( P3_SUB_357_1258_U11 , P3_SUB_357_1258_U9 , P3_SUB_357_1258_U211 );
and AND2_21221 ( P3_SUB_357_1258_U12 , P3_SUB_357_1258_U10 , P3_SUB_357_1258_U212 );
and AND2_21222 ( P3_SUB_357_1258_U13 , P3_SUB_357_1258_U11 , P3_SUB_357_1258_U213 );
and AND2_21223 ( P3_SUB_357_1258_U14 , P3_SUB_357_1258_U12 , P3_SUB_357_1258_U214 );
and AND2_21224 ( P3_SUB_357_1258_U15 , P3_SUB_357_1258_U255 , P3_SUB_357_1258_U252 );
and AND2_21225 ( P3_SUB_357_1258_U16 , P3_SUB_357_1258_U249 , P3_SUB_357_1258_U248 );
and AND2_21226 ( P3_SUB_357_1258_U17 , P3_SUB_357_1258_U244 , P3_SUB_357_1258_U241 );
and AND2_21227 ( P3_SUB_357_1258_U18 , P3_SUB_357_1258_U233 , P3_SUB_357_1258_U230 );
and AND2_21228 ( P3_SUB_357_1258_U19 , P3_SUB_357_1258_U227 , P3_SUB_357_1258_U303 );
and AND2_21229 ( P3_SUB_357_1258_U20 , P3_SUB_357_1258_U225 , P3_SUB_357_1258_U296 );
nand NAND3_21230 ( P3_SUB_357_1258_U21 , P3_SUB_357_1258_U426 , P3_SUB_357_1258_U425 , P3_SUB_357_1258_U307 );
not NOT1_21231 ( P3_SUB_357_1258_U22 , P3_ADD_357_U9 );
not NOT1_21232 ( P3_SUB_357_1258_U23 , P3_INSTADDRPOINTER_REG_7_ );
not NOT1_21233 ( P3_SUB_357_1258_U24 , P3_ADD_357_U8 );
not NOT1_21234 ( P3_SUB_357_1258_U25 , P3_INSTADDRPOINTER_REG_5_ );
not NOT1_21235 ( P3_SUB_357_1258_U26 , P3_ADD_357_U19 );
not NOT1_21236 ( P3_SUB_357_1258_U27 , P3_INSTADDRPOINTER_REG_4_ );
not NOT1_21237 ( P3_SUB_357_1258_U28 , P3_ADD_357_U10 );
not NOT1_21238 ( P3_SUB_357_1258_U29 , P3_INSTADDRPOINTER_REG_0_ );
nand NAND2_21239 ( P3_SUB_357_1258_U30 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_357_U10 );
not NOT1_21240 ( P3_SUB_357_1258_U31 , P3_SUB_357_U7 );
not NOT1_21241 ( P3_SUB_357_1258_U32 , P3_ADD_357_U13 );
not NOT1_21242 ( P3_SUB_357_1258_U33 , P3_INSTADDRPOINTER_REG_2_ );
not NOT1_21243 ( P3_SUB_357_1258_U34 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_21244 ( P3_SUB_357_1258_U35 , P3_ADD_357_U7 );
not NOT1_21245 ( P3_SUB_357_1258_U36 , P3_INSTADDRPOINTER_REG_3_ );
not NOT1_21246 ( P3_SUB_357_1258_U37 , P3_ADD_357_U17 );
not NOT1_21247 ( P3_SUB_357_1258_U38 , P3_INSTADDRPOINTER_REG_6_ );
not NOT1_21248 ( P3_SUB_357_1258_U39 , P3_ADD_357_U6 );
not NOT1_21249 ( P3_SUB_357_1258_U40 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_21250 ( P3_SUB_357_1258_U41 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_21251 ( P3_SUB_357_1258_U42 , P3_INSTADDRPOINTER_REG_25_ );
not NOT1_21252 ( P3_SUB_357_1258_U43 , P3_INSTADDRPOINTER_REG_26_ );
not NOT1_21253 ( P3_SUB_357_1258_U44 , P3_INSTADDRPOINTER_REG_24_ );
not NOT1_21254 ( P3_SUB_357_1258_U45 , P3_INSTADDRPOINTER_REG_23_ );
not NOT1_21255 ( P3_SUB_357_1258_U46 , P3_INSTADDRPOINTER_REG_22_ );
not NOT1_21256 ( P3_SUB_357_1258_U47 , P3_INSTADDRPOINTER_REG_19_ );
not NOT1_21257 ( P3_SUB_357_1258_U48 , P3_INSTADDRPOINTER_REG_21_ );
not NOT1_21258 ( P3_SUB_357_1258_U49 , P3_INSTADDRPOINTER_REG_18_ );
not NOT1_21259 ( P3_SUB_357_1258_U50 , P3_INSTADDRPOINTER_REG_12_ );
not NOT1_21260 ( P3_SUB_357_1258_U51 , P3_INSTADDRPOINTER_REG_13_ );
not NOT1_21261 ( P3_SUB_357_1258_U52 , P3_INSTADDRPOINTER_REG_11_ );
not NOT1_21262 ( P3_SUB_357_1258_U53 , P3_INSTADDRPOINTER_REG_10_ );
not NOT1_21263 ( P3_SUB_357_1258_U54 , P3_INSTADDRPOINTER_REG_14_ );
not NOT1_21264 ( P3_SUB_357_1258_U55 , P3_INSTADDRPOINTER_REG_15_ );
not NOT1_21265 ( P3_SUB_357_1258_U56 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_21266 ( P3_SUB_357_1258_U57 , P3_INSTADDRPOINTER_REG_19_ , P3_INSTADDRPOINTER_REG_20_ );
not NOT1_21267 ( P3_SUB_357_1258_U58 , P3_INSTADDRPOINTER_REG_27_ );
not NOT1_21268 ( P3_SUB_357_1258_U59 , P3_INSTADDRPOINTER_REG_29_ );
not NOT1_21269 ( P3_SUB_357_1258_U60 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND3_21270 ( P3_SUB_357_1258_U61 , P3_SUB_357_1258_U222 , P3_SUB_357_1258_U151 , P3_SUB_357_1258_U269 );
nand NAND2_21271 ( P3_SUB_357_1258_U62 , P3_SUB_357_1258_U105 , P3_SUB_357_1258_U218 );
nand NAND2_21272 ( P3_SUB_357_1258_U63 , P3_SUB_357_1258_U104 , P3_SUB_357_1258_U284 );
nand NAND2_21273 ( P3_SUB_357_1258_U64 , P3_SUB_357_1258_U276 , P3_SUB_357_1258_U205 );
nand NAND2_21274 ( P3_SUB_357_1258_U65 , P3_SUB_357_1258_U277 , P3_SUB_357_1258_U47 );
nand NAND2_21275 ( P3_SUB_357_1258_U66 , P3_SUB_357_U7 , P3_SUB_357_1258_U161 );
nand NAND2_21276 ( P3_SUB_357_1258_U67 , P3_SUB_357_1258_U102 , P3_SUB_357_1258_U198 );
nand NAND2_21277 ( P3_SUB_357_1258_U68 , P3_SUB_357_1258_U290 , P3_SUB_357_1258_U8 );
nand NAND2_21278 ( P3_SUB_357_1258_U69 , P3_SUB_357_1258_U484 , P3_SUB_357_1258_U483 );
nand NAND2_21279 ( P3_SUB_357_1258_U70 , P3_SUB_357_1258_U312 , P3_SUB_357_1258_U311 );
nand NAND2_21280 ( P3_SUB_357_1258_U71 , P3_SUB_357_1258_U319 , P3_SUB_357_1258_U318 );
nand NAND2_21281 ( P3_SUB_357_1258_U72 , P3_SUB_357_1258_U326 , P3_SUB_357_1258_U325 );
nand NAND2_21282 ( P3_SUB_357_1258_U73 , P3_SUB_357_1258_U333 , P3_SUB_357_1258_U332 );
nand NAND2_21283 ( P3_SUB_357_1258_U74 , P3_SUB_357_1258_U340 , P3_SUB_357_1258_U339 );
nand NAND2_21284 ( P3_SUB_357_1258_U75 , P3_SUB_357_1258_U345 , P3_SUB_357_1258_U344 );
nand NAND2_21285 ( P3_SUB_357_1258_U76 , P3_SUB_357_1258_U350 , P3_SUB_357_1258_U349 );
nand NAND2_21286 ( P3_SUB_357_1258_U77 , P3_SUB_357_1258_U361 , P3_SUB_357_1258_U360 );
nand NAND2_21287 ( P3_SUB_357_1258_U78 , P3_SUB_357_1258_U366 , P3_SUB_357_1258_U365 );
nand NAND2_21288 ( P3_SUB_357_1258_U79 , P3_SUB_357_1258_U373 , P3_SUB_357_1258_U372 );
nand NAND2_21289 ( P3_SUB_357_1258_U80 , P3_SUB_357_1258_U384 , P3_SUB_357_1258_U383 );
nand NAND2_21290 ( P3_SUB_357_1258_U81 , P3_SUB_357_1258_U391 , P3_SUB_357_1258_U390 );
nand NAND2_21291 ( P3_SUB_357_1258_U82 , P3_SUB_357_1258_U398 , P3_SUB_357_1258_U397 );
nand NAND2_21292 ( P3_SUB_357_1258_U83 , P3_SUB_357_1258_U405 , P3_SUB_357_1258_U404 );
nand NAND2_21293 ( P3_SUB_357_1258_U84 , P3_SUB_357_1258_U412 , P3_SUB_357_1258_U411 );
nand NAND2_21294 ( P3_SUB_357_1258_U85 , P3_SUB_357_1258_U419 , P3_SUB_357_1258_U418 );
nand NAND2_21295 ( P3_SUB_357_1258_U86 , P3_SUB_357_1258_U431 , P3_SUB_357_1258_U430 );
nand NAND2_21296 ( P3_SUB_357_1258_U87 , P3_SUB_357_1258_U438 , P3_SUB_357_1258_U437 );
nand NAND2_21297 ( P3_SUB_357_1258_U88 , P3_SUB_357_1258_U449 , P3_SUB_357_1258_U448 );
nand NAND2_21298 ( P3_SUB_357_1258_U89 , P3_SUB_357_1258_U456 , P3_SUB_357_1258_U455 );
nand NAND2_21299 ( P3_SUB_357_1258_U90 , P3_SUB_357_1258_U463 , P3_SUB_357_1258_U462 );
nand NAND2_21300 ( P3_SUB_357_1258_U91 , P3_SUB_357_1258_U470 , P3_SUB_357_1258_U469 );
nand NAND2_21301 ( P3_SUB_357_1258_U92 , P3_SUB_357_1258_U477 , P3_SUB_357_1258_U476 );
nand NAND2_21302 ( P3_SUB_357_1258_U93 , P3_SUB_357_1258_U482 , P3_SUB_357_1258_U481 );
and AND3_21303 ( P3_SUB_357_1258_U94 , P3_SUB_357_1258_U163 , P3_SUB_357_1258_U164 , P3_SUB_357_1258_U160 );
and AND2_21304 ( P3_SUB_357_1258_U95 , P3_ADD_357_U7 , P3_INSTADDRPOINTER_REG_3_ );
and AND2_21305 ( P3_SUB_357_1258_U96 , P3_SUB_357_1258_U168 , P3_SUB_357_1258_U162 );
and AND2_21306 ( P3_SUB_357_1258_U97 , P3_SUB_357_1258_U164 , P3_SUB_357_1258_U163 );
and AND2_21307 ( P3_SUB_357_1258_U98 , P3_SUB_357_1258_U7 , P3_SUB_357_1258_U154 );
and AND2_21308 ( P3_SUB_357_1258_U99 , P3_SUB_357_1258_U192 , P3_SUB_357_1258_U155 );
and AND2_21309 ( P3_SUB_357_1258_U100 , P3_SUB_357_1258_U99 , P3_SUB_357_1258_U8 );
and AND2_21310 ( P3_SUB_357_1258_U101 , P3_INSTADDRPOINTER_REG_17_ , P3_INSTADDRPOINTER_REG_16_ );
and AND2_21311 ( P3_SUB_357_1258_U102 , P3_SUB_357_1258_U199 , P3_SUB_357_1258_U56 );
and AND2_21312 ( P3_SUB_357_1258_U103 , P3_SUB_357_1258_U215 , P3_SUB_357_1258_U13 );
and AND2_21313 ( P3_SUB_357_1258_U104 , P3_SUB_357_1258_U14 , P3_SUB_357_1258_U216 );
and AND3_21314 ( P3_SUB_357_1258_U105 , P3_SUB_357_1258_U157 , P3_SUB_357_1258_U58 , P3_SUB_357_1258_U219 );
and AND2_21315 ( P3_SUB_357_1258_U106 , P3_SUB_357_1258_U219 , P3_SUB_357_1258_U157 );
and AND3_21316 ( P3_SUB_357_1258_U107 , P3_INSTADDRPOINTER_REG_31_ , P3_SUB_357_1258_U60 , P3_SUB_357_1258_U269 );
and AND2_21317 ( P3_SUB_357_1258_U108 , P3_INSTADDRPOINTER_REG_30_ , P3_INSTADDRPOINTER_REG_31_ );
and AND3_21318 ( P3_SUB_357_1258_U109 , P3_SUB_357_1258_U386 , P3_SUB_357_1258_U385 , P3_SUB_357_1258_U157 );
and AND2_21319 ( P3_SUB_357_1258_U110 , P3_SUB_357_1258_U232 , P3_SUB_357_1258_U153 );
and AND2_21320 ( P3_SUB_357_1258_U111 , P3_SUB_357_1258_U237 , P3_SUB_357_1258_U156 );
and AND2_21321 ( P3_SUB_357_1258_U112 , P3_SUB_357_1258_U243 , P3_SUB_357_1258_U156 );
and AND3_21322 ( P3_SUB_357_1258_U113 , P3_SUB_357_1258_U465 , P3_SUB_357_1258_U464 , P3_SUB_357_1258_U155 );
and AND2_21323 ( P3_SUB_357_1258_U114 , P3_SUB_357_1258_U254 , P3_SUB_357_1258_U154 );
nand NAND3_21324 ( P3_SUB_357_1258_U115 , P3_SUB_357_1258_U176 , P3_SUB_357_1258_U152 , P3_SUB_357_1258_U268 );
and AND2_21325 ( P3_SUB_357_1258_U116 , P3_SUB_357_1258_U314 , P3_SUB_357_1258_U313 );
nand NAND2_21326 ( P3_SUB_357_1258_U117 , P3_SUB_357_1258_U300 , P3_SUB_357_1258_U267 );
and AND2_21327 ( P3_SUB_357_1258_U118 , P3_SUB_357_1258_U321 , P3_SUB_357_1258_U320 );
nand NAND2_21328 ( P3_SUB_357_1258_U119 , P3_SUB_357_1258_U173 , P3_SUB_357_1258_U172 );
and AND2_21329 ( P3_SUB_357_1258_U120 , P3_SUB_357_1258_U328 , P3_SUB_357_1258_U327 );
nand NAND2_21330 ( P3_SUB_357_1258_U121 , P3_SUB_357_1258_U298 , P3_SUB_357_1258_U266 );
and AND2_21331 ( P3_SUB_357_1258_U122 , P3_SUB_357_1258_U335 , P3_SUB_357_1258_U334 );
nand NAND2_21332 ( P3_SUB_357_1258_U123 , P3_SUB_357_1258_U96 , P3_SUB_357_1258_U167 );
nand NAND2_21333 ( P3_SUB_357_1258_U124 , P3_SUB_357_1258_U181 , P3_SUB_357_1258_U180 );
nand NAND2_21334 ( P3_SUB_357_1258_U125 , P3_SUB_357_1258_U159 , P3_SUB_357_1258_U183 );
and AND2_21335 ( P3_SUB_357_1258_U126 , P3_SUB_357_1258_U356 , P3_SUB_357_1258_U355 );
nand NAND3_21336 ( P3_SUB_357_1258_U127 , P3_SUB_357_1258_U270 , P3_SUB_357_1258_U66 , P3_SUB_357_1258_U271 );
and AND2_21337 ( P3_SUB_357_1258_U128 , P3_SUB_357_1258_U368 , P3_SUB_357_1258_U367 );
nand NAND3_21338 ( P3_SUB_357_1258_U129 , P3_SUB_357_1258_U275 , P3_SUB_357_1258_U274 , P3_SUB_357_1258_U304 );
and AND2_21339 ( P3_SUB_357_1258_U130 , P3_SUB_357_1258_U379 , P3_SUB_357_1258_U378 );
nand NAND2_21340 ( P3_SUB_357_1258_U131 , P3_SUB_357_1258_U106 , P3_SUB_357_1258_U218 );
and AND2_21341 ( P3_SUB_357_1258_U132 , P3_SUB_357_1258_U393 , P3_SUB_357_1258_U392 );
nand NAND2_21342 ( P3_SUB_357_1258_U133 , P3_SUB_357_1258_U282 , P3_SUB_357_1258_U14 );
and AND2_21343 ( P3_SUB_357_1258_U134 , P3_SUB_357_1258_U400 , P3_SUB_357_1258_U399 );
nand NAND2_21344 ( P3_SUB_357_1258_U135 , P3_SUB_357_1258_U280 , P3_SUB_357_1258_U12 );
and AND2_21345 ( P3_SUB_357_1258_U136 , P3_SUB_357_1258_U407 , P3_SUB_357_1258_U406 );
nand NAND2_21346 ( P3_SUB_357_1258_U137 , P3_SUB_357_1258_U278 , P3_SUB_357_1258_U10 );
and AND2_21347 ( P3_SUB_357_1258_U138 , P3_SUB_357_1258_U414 , P3_SUB_357_1258_U413 );
nand NAND2_21348 ( P3_SUB_357_1258_U139 , P3_SUB_357_1258_U111 , P3_SUB_357_1258_U236 );
and AND2_21349 ( P3_SUB_357_1258_U140 , P3_SUB_357_1258_U433 , P3_SUB_357_1258_U432 );
nand NAND3_21350 ( P3_SUB_357_1258_U141 , P3_SUB_357_1258_U272 , P3_SUB_357_1258_U201 , P3_SUB_357_1258_U273 );
and AND2_21351 ( P3_SUB_357_1258_U142 , P3_SUB_357_1258_U444 , P3_SUB_357_1258_U443 );
nand NAND2_21352 ( P3_SUB_357_1258_U143 , P3_SUB_357_1258_U199 , P3_SUB_357_1258_U198 );
and AND2_21353 ( P3_SUB_357_1258_U144 , P3_SUB_357_1258_U451 , P3_SUB_357_1258_U450 );
nand NAND2_21354 ( P3_SUB_357_1258_U145 , P3_SUB_357_1258_U195 , P3_SUB_357_1258_U194 );
and AND2_21355 ( P3_SUB_357_1258_U146 , P3_SUB_357_1258_U458 , P3_SUB_357_1258_U457 );
nand NAND2_21356 ( P3_SUB_357_1258_U147 , P3_SUB_357_1258_U100 , P3_SUB_357_1258_U292 );
and AND2_21357 ( P3_SUB_357_1258_U148 , P3_SUB_357_1258_U472 , P3_SUB_357_1258_U471 );
nand NAND2_21358 ( P3_SUB_357_1258_U149 , P3_SUB_357_1258_U288 , P3_SUB_357_1258_U5 );
nand NAND2_21359 ( P3_SUB_357_1258_U150 , P3_SUB_357_1258_U286 , P3_SUB_357_1258_U186 );
nand NAND2_21360 ( P3_SUB_357_1258_U151 , P3_ADD_357_U6 , P3_SUB_357_1258_U129 );
nand NAND2_21361 ( P3_SUB_357_1258_U152 , P3_ADD_357_U6 , P3_SUB_357_1258_U117 );
nand NAND2_21362 ( P3_SUB_357_1258_U153 , P3_SUB_357_1258_U217 , P3_SUB_357_1258_U39 );
nand NAND2_21363 ( P3_SUB_357_1258_U154 , P3_SUB_357_1258_U191 , P3_SUB_357_1258_U39 );
nand NAND2_21364 ( P3_SUB_357_1258_U155 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_357_U6 );
nand NAND2_21365 ( P3_SUB_357_1258_U156 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_357_U6 );
nand NAND2_21366 ( P3_SUB_357_1258_U157 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_357_U6 );
not NOT1_21367 ( P3_SUB_357_1258_U158 , P3_SUB_357_1258_U66 );
nand NAND2_21368 ( P3_SUB_357_1258_U159 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_357_U13 );
or OR2_21369 ( P3_SUB_357_1258_U160 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_357_U19 );
not NOT1_21370 ( P3_SUB_357_1258_U161 , P3_SUB_357_1258_U30 );
nand NAND2_21371 ( P3_SUB_357_1258_U162 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_357_U19 );
or OR2_21372 ( P3_SUB_357_1258_U163 , P3_ADD_357_U7 , P3_INSTADDRPOINTER_REG_3_ );
or OR2_21373 ( P3_SUB_357_1258_U164 , P3_ADD_357_U13 , P3_INSTADDRPOINTER_REG_2_ );
not NOT1_21374 ( P3_SUB_357_1258_U165 , P3_SUB_357_1258_U127 );
nand NAND4_21375 ( P3_SUB_357_1258_U166 , P3_SUB_357_1258_U271 , P3_SUB_357_1258_U270 , P3_SUB_357_1258_U159 , P3_SUB_357_1258_U66 );
nand NAND2_21376 ( P3_SUB_357_1258_U167 , P3_SUB_357_1258_U94 , P3_SUB_357_1258_U166 );
nand NAND2_21377 ( P3_SUB_357_1258_U168 , P3_SUB_357_1258_U95 , P3_SUB_357_1258_U160 );
not NOT1_21378 ( P3_SUB_357_1258_U169 , P3_SUB_357_1258_U123 );
or OR2_21379 ( P3_SUB_357_1258_U170 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_357_U8 );
or OR2_21380 ( P3_SUB_357_1258_U171 , P3_ADD_357_U17 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_21381 ( P3_SUB_357_1258_U172 , P3_SUB_357_1258_U171 , P3_SUB_357_1258_U121 );
nand NAND2_21382 ( P3_SUB_357_1258_U173 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_357_U17 );
not NOT1_21383 ( P3_SUB_357_1258_U174 , P3_SUB_357_1258_U119 );
or OR2_21384 ( P3_SUB_357_1258_U175 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_357_U9 );
nand NAND2_21385 ( P3_SUB_357_1258_U176 , P3_INSTADDRPOINTER_REG_8_ , P3_SUB_357_1258_U117 );
not NOT1_21386 ( P3_SUB_357_1258_U177 , P3_SUB_357_1258_U115 );
or OR2_21387 ( P3_SUB_357_1258_U178 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_357_U6 );
nand NAND2_21388 ( P3_SUB_357_1258_U179 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_357_U6 );
nand NAND2_21389 ( P3_SUB_357_1258_U180 , P3_SUB_357_1258_U97 , P3_SUB_357_1258_U166 );
nand NAND2_21390 ( P3_SUB_357_1258_U181 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_357_U7 );
not NOT1_21391 ( P3_SUB_357_1258_U182 , P3_SUB_357_1258_U124 );
nand NAND2_21392 ( P3_SUB_357_1258_U183 , P3_SUB_357_1258_U127 , P3_SUB_357_1258_U164 );
not NOT1_21393 ( P3_SUB_357_1258_U184 , P3_SUB_357_1258_U125 );
nand NAND2_21394 ( P3_SUB_357_1258_U185 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_357_U7 );
nand NAND2_21395 ( P3_SUB_357_1258_U186 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_357_U6 );
or OR2_21396 ( P3_SUB_357_1258_U187 , P3_ADD_357_U6 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_21397 ( P3_SUB_357_1258_U188 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_357_U6 );
or OR2_21398 ( P3_SUB_357_1258_U189 , P3_ADD_357_U6 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_21399 ( P3_SUB_357_1258_U190 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_357_U6 );
nand NAND2_21400 ( P3_SUB_357_1258_U191 , P3_INSTADDRPOINTER_REG_13_ , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_21401 ( P3_SUB_357_1258_U192 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_357_U6 );
or OR2_21402 ( P3_SUB_357_1258_U193 , P3_ADD_357_U6 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_21403 ( P3_SUB_357_1258_U194 , P3_SUB_357_1258_U193 , P3_SUB_357_1258_U147 );
nand NAND2_21404 ( P3_SUB_357_1258_U195 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_357_U6 );
not NOT1_21405 ( P3_SUB_357_1258_U196 , P3_SUB_357_1258_U145 );
or OR2_21406 ( P3_SUB_357_1258_U197 , P3_ADD_357_U6 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_21407 ( P3_SUB_357_1258_U198 , P3_SUB_357_1258_U197 , P3_SUB_357_1258_U145 );
nand NAND2_21408 ( P3_SUB_357_1258_U199 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_357_U6 );
not NOT1_21409 ( P3_SUB_357_1258_U200 , P3_SUB_357_1258_U143 );
nand NAND2_21410 ( P3_SUB_357_1258_U201 , P3_SUB_357_1258_U101 , P3_SUB_357_1258_U143 );
not NOT1_21411 ( P3_SUB_357_1258_U202 , P3_SUB_357_1258_U67 );
not NOT1_21412 ( P3_SUB_357_1258_U203 , P3_SUB_357_1258_U141 );
or OR2_21413 ( P3_SUB_357_1258_U204 , P3_ADD_357_U6 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_21414 ( P3_SUB_357_1258_U205 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_357_U6 );
nand NAND2_21415 ( P3_SUB_357_1258_U206 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_357_U6 );
not NOT1_21416 ( P3_SUB_357_1258_U207 , P3_SUB_357_1258_U57 );
nand NAND2_21417 ( P3_SUB_357_1258_U208 , P3_SUB_357_1258_U207 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_21418 ( P3_SUB_357_1258_U209 , P3_SUB_357_1258_U39 , P3_SUB_357_1258_U208 );
nand NAND2_21419 ( P3_SUB_357_1258_U210 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_357_U6 );
or OR2_21420 ( P3_SUB_357_1258_U211 , P3_ADD_357_U6 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_21421 ( P3_SUB_357_1258_U212 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_357_U6 );
or OR2_21422 ( P3_SUB_357_1258_U213 , P3_ADD_357_U6 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_21423 ( P3_SUB_357_1258_U214 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_357_U6 );
or OR2_21424 ( P3_SUB_357_1258_U215 , P3_ADD_357_U6 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_21425 ( P3_SUB_357_1258_U216 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_357_U6 );
nand NAND2_21426 ( P3_SUB_357_1258_U217 , P3_INSTADDRPOINTER_REG_26_ , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_21427 ( P3_SUB_357_1258_U218 , P3_SUB_357_1258_U63 , P3_SUB_357_1258_U153 );
nand NAND2_21428 ( P3_SUB_357_1258_U219 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_357_U6 );
not NOT1_21429 ( P3_SUB_357_1258_U220 , P3_SUB_357_1258_U131 );
not NOT1_21430 ( P3_SUB_357_1258_U221 , P3_SUB_357_1258_U62 );
nand NAND2_21431 ( P3_SUB_357_1258_U222 , P3_INSTADDRPOINTER_REG_29_ , P3_SUB_357_1258_U129 );
not NOT1_21432 ( P3_SUB_357_1258_U223 , P3_SUB_357_1258_U61 );
nand NAND2_21433 ( P3_SUB_357_1258_U224 , P3_SUB_357_1258_U151 , P3_SUB_357_1258_U107 );
nand NAND3_21434 ( P3_SUB_357_1258_U225 , P3_SUB_357_1258_U354 , P3_SUB_357_1258_U353 , P3_SUB_357_1258_U294 );
nand NAND2_21435 ( P3_SUB_357_1258_U226 , P3_SUB_357_1258_U221 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND3_21436 ( P3_SUB_357_1258_U227 , P3_SUB_357_1258_U377 , P3_SUB_357_1258_U376 , P3_SUB_357_1258_U62 );
or OR2_21437 ( P3_SUB_357_1258_U228 , P3_ADD_357_U6 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_21438 ( P3_SUB_357_1258_U229 , P3_SUB_357_1258_U228 , P3_SUB_357_1258_U63 );
nand NAND2_21439 ( P3_SUB_357_1258_U230 , P3_SUB_357_1258_U109 , P3_SUB_357_1258_U229 );
nand NAND2_21440 ( P3_SUB_357_1258_U231 , P3_SUB_357_1258_U285 , P3_SUB_357_1258_U157 );
nand NAND2_21441 ( P3_SUB_357_1258_U232 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_357_U6 );
nand NAND2_21442 ( P3_SUB_357_1258_U233 , P3_SUB_357_1258_U110 , P3_SUB_357_1258_U231 );
or OR2_21443 ( P3_SUB_357_1258_U234 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_357_U6 );
not NOT1_21444 ( P3_SUB_357_1258_U235 , P3_SUB_357_1258_U65 );
nand NAND2_21445 ( P3_SUB_357_1258_U236 , P3_ADD_357_U6 , P3_SUB_357_1258_U65 );
nand NAND2_21446 ( P3_SUB_357_1258_U237 , P3_SUB_357_1258_U207 , P3_SUB_357_1258_U64 );
not NOT1_21447 ( P3_SUB_357_1258_U238 , P3_SUB_357_1258_U139 );
nand NAND2_21448 ( P3_SUB_357_1258_U239 , P3_SUB_357_1258_U235 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_21449 ( P3_SUB_357_1258_U240 , P3_INSTADDRPOINTER_REG_19_ , P3_SUB_357_1258_U64 );
nand NAND3_21450 ( P3_SUB_357_1258_U241 , P3_SUB_357_1258_U421 , P3_SUB_357_1258_U420 , P3_SUB_357_1258_U240 );
nand NAND2_21451 ( P3_SUB_357_1258_U242 , P3_SUB_357_1258_U277 , P3_SUB_357_1258_U206 );
nand NAND2_21452 ( P3_SUB_357_1258_U243 , P3_SUB_357_1258_U57 , P3_SUB_357_1258_U39 );
nand NAND2_21453 ( P3_SUB_357_1258_U244 , P3_SUB_357_1258_U112 , P3_SUB_357_1258_U242 );
or OR2_21454 ( P3_SUB_357_1258_U245 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_357_U6 );
nand NAND2_21455 ( P3_SUB_357_1258_U246 , P3_SUB_357_1258_U202 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_21456 ( P3_SUB_357_1258_U247 , P3_INSTADDRPOINTER_REG_16_ , P3_SUB_357_1258_U143 );
nand NAND3_21457 ( P3_SUB_357_1258_U248 , P3_SUB_357_1258_U440 , P3_SUB_357_1258_U439 , P3_SUB_357_1258_U247 );
nand NAND3_21458 ( P3_SUB_357_1258_U249 , P3_SUB_357_1258_U442 , P3_SUB_357_1258_U441 , P3_SUB_357_1258_U67 );
or OR2_21459 ( P3_SUB_357_1258_U250 , P3_ADD_357_U6 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_21460 ( P3_SUB_357_1258_U251 , P3_SUB_357_1258_U250 , P3_SUB_357_1258_U68 );
nand NAND2_21461 ( P3_SUB_357_1258_U252 , P3_SUB_357_1258_U113 , P3_SUB_357_1258_U251 );
nand NAND2_21462 ( P3_SUB_357_1258_U253 , P3_SUB_357_1258_U291 , P3_SUB_357_1258_U155 );
nand NAND2_21463 ( P3_SUB_357_1258_U254 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_357_U6 );
nand NAND2_21464 ( P3_SUB_357_1258_U255 , P3_SUB_357_1258_U114 , P3_SUB_357_1258_U253 );
or OR2_21465 ( P3_SUB_357_1258_U256 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_357_U6 );
nand NAND2_21466 ( P3_SUB_357_1258_U257 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_357_U6 );
nand NAND2_21467 ( P3_SUB_357_1258_U258 , P3_SUB_357_1258_U179 , P3_SUB_357_1258_U178 );
nand NAND2_21468 ( P3_SUB_357_1258_U259 , P3_SUB_357_1258_U162 , P3_SUB_357_1258_U160 );
nand NAND2_21469 ( P3_SUB_357_1258_U260 , P3_SUB_357_1258_U185 , P3_SUB_357_1258_U163 );
nand NAND2_21470 ( P3_SUB_357_1258_U261 , P3_SUB_357_1258_U164 , P3_SUB_357_1258_U159 );
nand NAND2_21471 ( P3_SUB_357_1258_U262 , P3_SUB_357_1258_U234 , P3_SUB_357_1258_U157 );
nand NAND2_21472 ( P3_SUB_357_1258_U263 , P3_SUB_357_1258_U245 , P3_SUB_357_1258_U206 );
nand NAND2_21473 ( P3_SUB_357_1258_U264 , P3_SUB_357_1258_U256 , P3_SUB_357_1258_U155 );
nand NAND2_21474 ( P3_SUB_357_1258_U265 , P3_SUB_357_1258_U257 , P3_SUB_357_1258_U187 );
nand NAND2_21475 ( P3_SUB_357_1258_U266 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_357_U8 );
nand NAND2_21476 ( P3_SUB_357_1258_U267 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_357_U9 );
nand NAND2_21477 ( P3_SUB_357_1258_U268 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_357_U6 );
nand NAND2_21478 ( P3_SUB_357_1258_U269 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_357_U6 );
nand NAND2_21479 ( P3_SUB_357_1258_U270 , P3_INSTADDRPOINTER_REG_1_ , P3_SUB_357_1258_U161 );
nand NAND2_21480 ( P3_SUB_357_1258_U271 , P3_INSTADDRPOINTER_REG_1_ , P3_SUB_357_U7 );
nand NAND2_21481 ( P3_SUB_357_1258_U272 , P3_ADD_357_U6 , P3_SUB_357_1258_U67 );
nand NAND2_21482 ( P3_SUB_357_1258_U273 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_357_U6 );
nand NAND2_21483 ( P3_SUB_357_1258_U274 , P3_ADD_357_U6 , P3_SUB_357_1258_U62 );
nand NAND2_21484 ( P3_SUB_357_1258_U275 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_357_U6 );
nand NAND2_21485 ( P3_SUB_357_1258_U276 , P3_SUB_357_1258_U204 , P3_SUB_357_1258_U141 );
not NOT1_21486 ( P3_SUB_357_1258_U277 , P3_SUB_357_1258_U64 );
nand NAND2_21487 ( P3_SUB_357_1258_U278 , P3_SUB_357_1258_U9 , P3_SUB_357_1258_U141 );
not NOT1_21488 ( P3_SUB_357_1258_U279 , P3_SUB_357_1258_U137 );
nand NAND2_21489 ( P3_SUB_357_1258_U280 , P3_SUB_357_1258_U11 , P3_SUB_357_1258_U141 );
not NOT1_21490 ( P3_SUB_357_1258_U281 , P3_SUB_357_1258_U135 );
nand NAND2_21491 ( P3_SUB_357_1258_U282 , P3_SUB_357_1258_U13 , P3_SUB_357_1258_U141 );
not NOT1_21492 ( P3_SUB_357_1258_U283 , P3_SUB_357_1258_U133 );
nand NAND2_21493 ( P3_SUB_357_1258_U284 , P3_SUB_357_1258_U103 , P3_SUB_357_1258_U141 );
not NOT1_21494 ( P3_SUB_357_1258_U285 , P3_SUB_357_1258_U63 );
nand NAND2_21495 ( P3_SUB_357_1258_U286 , P3_SUB_357_1258_U178 , P3_SUB_357_1258_U115 );
not NOT1_21496 ( P3_SUB_357_1258_U287 , P3_SUB_357_1258_U150 );
nand NAND2_21497 ( P3_SUB_357_1258_U288 , P3_SUB_357_1258_U6 , P3_SUB_357_1258_U115 );
not NOT1_21498 ( P3_SUB_357_1258_U289 , P3_SUB_357_1258_U149 );
nand NAND2_21499 ( P3_SUB_357_1258_U290 , P3_SUB_357_1258_U7 , P3_SUB_357_1258_U115 );
not NOT1_21500 ( P3_SUB_357_1258_U291 , P3_SUB_357_1258_U68 );
nand NAND2_21501 ( P3_SUB_357_1258_U292 , P3_SUB_357_1258_U98 , P3_SUB_357_1258_U115 );
not NOT1_21502 ( P3_SUB_357_1258_U293 , P3_SUB_357_1258_U147 );
nand NAND2_21503 ( P3_SUB_357_1258_U294 , P3_SUB_357_1258_U223 , P3_SUB_357_1258_U60 );
nand NAND2_21504 ( P3_SUB_357_1258_U295 , P3_INSTADDRPOINTER_REG_30_ , P3_SUB_357_1258_U61 );
nand NAND3_21505 ( P3_SUB_357_1258_U296 , P3_SUB_357_1258_U352 , P3_SUB_357_1258_U351 , P3_SUB_357_1258_U295 );
nand NAND2_21506 ( P3_SUB_357_1258_U297 , P3_SUB_357_1258_U108 , P3_SUB_357_1258_U61 );
nand NAND2_21507 ( P3_SUB_357_1258_U298 , P3_SUB_357_1258_U170 , P3_SUB_357_1258_U123 );
not NOT1_21508 ( P3_SUB_357_1258_U299 , P3_SUB_357_1258_U121 );
nand NAND2_21509 ( P3_SUB_357_1258_U300 , P3_SUB_357_1258_U175 , P3_SUB_357_1258_U119 );
not NOT1_21510 ( P3_SUB_357_1258_U301 , P3_SUB_357_1258_U117 );
nand NAND2_21511 ( P3_SUB_357_1258_U302 , P3_INSTADDRPOINTER_REG_27_ , P3_SUB_357_1258_U131 );
nand NAND3_21512 ( P3_SUB_357_1258_U303 , P3_SUB_357_1258_U375 , P3_SUB_357_1258_U374 , P3_SUB_357_1258_U302 );
nand NAND2_21513 ( P3_SUB_357_1258_U304 , P3_SUB_357_1258_U4 , P3_SUB_357_1258_U131 );
not NOT1_21514 ( P3_SUB_357_1258_U305 , P3_SUB_357_1258_U129 );
nand NAND2_21515 ( P3_SUB_357_1258_U306 , P3_SUB_357_1258_U4 , P3_SUB_357_1258_U131 );
nand NAND2_21516 ( P3_SUB_357_1258_U307 , P3_SUB_357_1258_U158 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_21517 ( P3_SUB_357_1258_U308 , P3_ADD_357_U6 , P3_SUB_357_1258_U41 );
nand NAND2_21518 ( P3_SUB_357_1258_U309 , P3_INSTADDRPOINTER_REG_9_ , P3_SUB_357_1258_U39 );
nand NAND2_21519 ( P3_SUB_357_1258_U310 , P3_SUB_357_1258_U309 , P3_SUB_357_1258_U308 );
nand NAND2_21520 ( P3_SUB_357_1258_U311 , P3_SUB_357_1258_U258 , P3_SUB_357_1258_U115 );
nand NAND2_21521 ( P3_SUB_357_1258_U312 , P3_SUB_357_1258_U177 , P3_SUB_357_1258_U310 );
nand NAND2_21522 ( P3_SUB_357_1258_U313 , P3_ADD_357_U6 , P3_SUB_357_1258_U40 );
nand NAND2_21523 ( P3_SUB_357_1258_U314 , P3_INSTADDRPOINTER_REG_8_ , P3_SUB_357_1258_U39 );
nand NAND2_21524 ( P3_SUB_357_1258_U315 , P3_ADD_357_U6 , P3_SUB_357_1258_U40 );
nand NAND2_21525 ( P3_SUB_357_1258_U316 , P3_INSTADDRPOINTER_REG_8_ , P3_SUB_357_1258_U39 );
nand NAND2_21526 ( P3_SUB_357_1258_U317 , P3_SUB_357_1258_U316 , P3_SUB_357_1258_U315 );
nand NAND2_21527 ( P3_SUB_357_1258_U318 , P3_SUB_357_1258_U116 , P3_SUB_357_1258_U117 );
nand NAND2_21528 ( P3_SUB_357_1258_U319 , P3_SUB_357_1258_U301 , P3_SUB_357_1258_U317 );
nand NAND2_21529 ( P3_SUB_357_1258_U320 , P3_INSTADDRPOINTER_REG_7_ , P3_SUB_357_1258_U22 );
nand NAND2_21530 ( P3_SUB_357_1258_U321 , P3_ADD_357_U9 , P3_SUB_357_1258_U23 );
nand NAND2_21531 ( P3_SUB_357_1258_U322 , P3_INSTADDRPOINTER_REG_7_ , P3_SUB_357_1258_U22 );
nand NAND2_21532 ( P3_SUB_357_1258_U323 , P3_ADD_357_U9 , P3_SUB_357_1258_U23 );
nand NAND2_21533 ( P3_SUB_357_1258_U324 , P3_SUB_357_1258_U323 , P3_SUB_357_1258_U322 );
nand NAND2_21534 ( P3_SUB_357_1258_U325 , P3_SUB_357_1258_U118 , P3_SUB_357_1258_U119 );
nand NAND2_21535 ( P3_SUB_357_1258_U326 , P3_SUB_357_1258_U174 , P3_SUB_357_1258_U324 );
nand NAND2_21536 ( P3_SUB_357_1258_U327 , P3_INSTADDRPOINTER_REG_6_ , P3_SUB_357_1258_U37 );
nand NAND2_21537 ( P3_SUB_357_1258_U328 , P3_ADD_357_U17 , P3_SUB_357_1258_U38 );
nand NAND2_21538 ( P3_SUB_357_1258_U329 , P3_INSTADDRPOINTER_REG_6_ , P3_SUB_357_1258_U37 );
nand NAND2_21539 ( P3_SUB_357_1258_U330 , P3_ADD_357_U17 , P3_SUB_357_1258_U38 );
nand NAND2_21540 ( P3_SUB_357_1258_U331 , P3_SUB_357_1258_U330 , P3_SUB_357_1258_U329 );
nand NAND2_21541 ( P3_SUB_357_1258_U332 , P3_SUB_357_1258_U120 , P3_SUB_357_1258_U121 );
nand NAND2_21542 ( P3_SUB_357_1258_U333 , P3_SUB_357_1258_U299 , P3_SUB_357_1258_U331 );
nand NAND2_21543 ( P3_SUB_357_1258_U334 , P3_INSTADDRPOINTER_REG_5_ , P3_SUB_357_1258_U24 );
nand NAND2_21544 ( P3_SUB_357_1258_U335 , P3_ADD_357_U8 , P3_SUB_357_1258_U25 );
nand NAND2_21545 ( P3_SUB_357_1258_U336 , P3_INSTADDRPOINTER_REG_5_ , P3_SUB_357_1258_U24 );
nand NAND2_21546 ( P3_SUB_357_1258_U337 , P3_ADD_357_U8 , P3_SUB_357_1258_U25 );
nand NAND2_21547 ( P3_SUB_357_1258_U338 , P3_SUB_357_1258_U337 , P3_SUB_357_1258_U336 );
nand NAND2_21548 ( P3_SUB_357_1258_U339 , P3_SUB_357_1258_U122 , P3_SUB_357_1258_U123 );
nand NAND2_21549 ( P3_SUB_357_1258_U340 , P3_SUB_357_1258_U169 , P3_SUB_357_1258_U338 );
nand NAND2_21550 ( P3_SUB_357_1258_U341 , P3_INSTADDRPOINTER_REG_4_ , P3_SUB_357_1258_U26 );
nand NAND2_21551 ( P3_SUB_357_1258_U342 , P3_ADD_357_U19 , P3_SUB_357_1258_U27 );
nand NAND2_21552 ( P3_SUB_357_1258_U343 , P3_SUB_357_1258_U342 , P3_SUB_357_1258_U341 );
nand NAND2_21553 ( P3_SUB_357_1258_U344 , P3_SUB_357_1258_U259 , P3_SUB_357_1258_U124 );
nand NAND2_21554 ( P3_SUB_357_1258_U345 , P3_SUB_357_1258_U182 , P3_SUB_357_1258_U343 );
nand NAND2_21555 ( P3_SUB_357_1258_U346 , P3_INSTADDRPOINTER_REG_3_ , P3_SUB_357_1258_U35 );
nand NAND2_21556 ( P3_SUB_357_1258_U347 , P3_ADD_357_U7 , P3_SUB_357_1258_U36 );
nand NAND2_21557 ( P3_SUB_357_1258_U348 , P3_SUB_357_1258_U347 , P3_SUB_357_1258_U346 );
nand NAND2_21558 ( P3_SUB_357_1258_U349 , P3_SUB_357_1258_U260 , P3_SUB_357_1258_U125 );
nand NAND2_21559 ( P3_SUB_357_1258_U350 , P3_SUB_357_1258_U184 , P3_SUB_357_1258_U348 );
nand NAND2_21560 ( P3_SUB_357_1258_U351 , P3_INSTADDRPOINTER_REG_31_ , P3_SUB_357_1258_U39 );
nand NAND2_21561 ( P3_SUB_357_1258_U352 , P3_ADD_357_U6 , P3_SUB_357_1258_U224 );
nand NAND2_21562 ( P3_SUB_357_1258_U353 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_357_U6 );
nand NAND2_21563 ( P3_SUB_357_1258_U354 , P3_SUB_357_1258_U297 , P3_SUB_357_1258_U39 );
nand NAND2_21564 ( P3_SUB_357_1258_U355 , P3_ADD_357_U6 , P3_SUB_357_1258_U60 );
nand NAND2_21565 ( P3_SUB_357_1258_U356 , P3_INSTADDRPOINTER_REG_30_ , P3_SUB_357_1258_U39 );
nand NAND2_21566 ( P3_SUB_357_1258_U357 , P3_ADD_357_U6 , P3_SUB_357_1258_U60 );
nand NAND2_21567 ( P3_SUB_357_1258_U358 , P3_INSTADDRPOINTER_REG_30_ , P3_SUB_357_1258_U39 );
nand NAND2_21568 ( P3_SUB_357_1258_U359 , P3_SUB_357_1258_U358 , P3_SUB_357_1258_U357 );
nand NAND2_21569 ( P3_SUB_357_1258_U360 , P3_SUB_357_1258_U126 , P3_SUB_357_1258_U61 );
nand NAND2_21570 ( P3_SUB_357_1258_U361 , P3_SUB_357_1258_U359 , P3_SUB_357_1258_U223 );
nand NAND2_21571 ( P3_SUB_357_1258_U362 , P3_INSTADDRPOINTER_REG_2_ , P3_SUB_357_1258_U32 );
nand NAND2_21572 ( P3_SUB_357_1258_U363 , P3_ADD_357_U13 , P3_SUB_357_1258_U33 );
nand NAND2_21573 ( P3_SUB_357_1258_U364 , P3_SUB_357_1258_U363 , P3_SUB_357_1258_U362 );
nand NAND2_21574 ( P3_SUB_357_1258_U365 , P3_SUB_357_1258_U261 , P3_SUB_357_1258_U127 );
nand NAND2_21575 ( P3_SUB_357_1258_U366 , P3_SUB_357_1258_U165 , P3_SUB_357_1258_U364 );
nand NAND2_21576 ( P3_SUB_357_1258_U367 , P3_ADD_357_U6 , P3_SUB_357_1258_U59 );
nand NAND2_21577 ( P3_SUB_357_1258_U368 , P3_INSTADDRPOINTER_REG_29_ , P3_SUB_357_1258_U39 );
nand NAND2_21578 ( P3_SUB_357_1258_U369 , P3_ADD_357_U6 , P3_SUB_357_1258_U59 );
nand NAND2_21579 ( P3_SUB_357_1258_U370 , P3_INSTADDRPOINTER_REG_29_ , P3_SUB_357_1258_U39 );
nand NAND2_21580 ( P3_SUB_357_1258_U371 , P3_SUB_357_1258_U370 , P3_SUB_357_1258_U369 );
nand NAND2_21581 ( P3_SUB_357_1258_U372 , P3_SUB_357_1258_U128 , P3_SUB_357_1258_U129 );
nand NAND2_21582 ( P3_SUB_357_1258_U373 , P3_SUB_357_1258_U305 , P3_SUB_357_1258_U371 );
nand NAND2_21583 ( P3_SUB_357_1258_U374 , P3_INSTADDRPOINTER_REG_28_ , P3_SUB_357_1258_U39 );
nand NAND2_21584 ( P3_SUB_357_1258_U375 , P3_ADD_357_U6 , P3_SUB_357_1258_U226 );
nand NAND2_21585 ( P3_SUB_357_1258_U376 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_357_U6 );
nand NAND2_21586 ( P3_SUB_357_1258_U377 , P3_SUB_357_1258_U306 , P3_SUB_357_1258_U39 );
nand NAND2_21587 ( P3_SUB_357_1258_U378 , P3_INSTADDRPOINTER_REG_27_ , P3_SUB_357_1258_U39 );
nand NAND2_21588 ( P3_SUB_357_1258_U379 , P3_ADD_357_U6 , P3_SUB_357_1258_U58 );
nand NAND2_21589 ( P3_SUB_357_1258_U380 , P3_INSTADDRPOINTER_REG_27_ , P3_SUB_357_1258_U39 );
nand NAND2_21590 ( P3_SUB_357_1258_U381 , P3_ADD_357_U6 , P3_SUB_357_1258_U58 );
nand NAND2_21591 ( P3_SUB_357_1258_U382 , P3_SUB_357_1258_U381 , P3_SUB_357_1258_U380 );
nand NAND2_21592 ( P3_SUB_357_1258_U383 , P3_SUB_357_1258_U130 , P3_SUB_357_1258_U131 );
nand NAND2_21593 ( P3_SUB_357_1258_U384 , P3_SUB_357_1258_U220 , P3_SUB_357_1258_U382 );
nand NAND2_21594 ( P3_SUB_357_1258_U385 , P3_INSTADDRPOINTER_REG_26_ , P3_SUB_357_1258_U39 );
nand NAND2_21595 ( P3_SUB_357_1258_U386 , P3_ADD_357_U6 , P3_SUB_357_1258_U43 );
nand NAND2_21596 ( P3_SUB_357_1258_U387 , P3_INSTADDRPOINTER_REG_25_ , P3_SUB_357_1258_U39 );
nand NAND2_21597 ( P3_SUB_357_1258_U388 , P3_ADD_357_U6 , P3_SUB_357_1258_U42 );
nand NAND2_21598 ( P3_SUB_357_1258_U389 , P3_SUB_357_1258_U388 , P3_SUB_357_1258_U387 );
nand NAND2_21599 ( P3_SUB_357_1258_U390 , P3_SUB_357_1258_U63 , P3_SUB_357_1258_U262 );
nand NAND2_21600 ( P3_SUB_357_1258_U391 , P3_SUB_357_1258_U389 , P3_SUB_357_1258_U285 );
nand NAND2_21601 ( P3_SUB_357_1258_U392 , P3_INSTADDRPOINTER_REG_24_ , P3_SUB_357_1258_U39 );
nand NAND2_21602 ( P3_SUB_357_1258_U393 , P3_ADD_357_U6 , P3_SUB_357_1258_U44 );
nand NAND2_21603 ( P3_SUB_357_1258_U394 , P3_INSTADDRPOINTER_REG_24_ , P3_SUB_357_1258_U39 );
nand NAND2_21604 ( P3_SUB_357_1258_U395 , P3_ADD_357_U6 , P3_SUB_357_1258_U44 );
nand NAND2_21605 ( P3_SUB_357_1258_U396 , P3_SUB_357_1258_U395 , P3_SUB_357_1258_U394 );
nand NAND2_21606 ( P3_SUB_357_1258_U397 , P3_SUB_357_1258_U132 , P3_SUB_357_1258_U133 );
nand NAND2_21607 ( P3_SUB_357_1258_U398 , P3_SUB_357_1258_U283 , P3_SUB_357_1258_U396 );
nand NAND2_21608 ( P3_SUB_357_1258_U399 , P3_INSTADDRPOINTER_REG_23_ , P3_SUB_357_1258_U39 );
nand NAND2_21609 ( P3_SUB_357_1258_U400 , P3_ADD_357_U6 , P3_SUB_357_1258_U45 );
nand NAND2_21610 ( P3_SUB_357_1258_U401 , P3_INSTADDRPOINTER_REG_23_ , P3_SUB_357_1258_U39 );
nand NAND2_21611 ( P3_SUB_357_1258_U402 , P3_ADD_357_U6 , P3_SUB_357_1258_U45 );
nand NAND2_21612 ( P3_SUB_357_1258_U403 , P3_SUB_357_1258_U402 , P3_SUB_357_1258_U401 );
nand NAND2_21613 ( P3_SUB_357_1258_U404 , P3_SUB_357_1258_U134 , P3_SUB_357_1258_U135 );
nand NAND2_21614 ( P3_SUB_357_1258_U405 , P3_SUB_357_1258_U281 , P3_SUB_357_1258_U403 );
nand NAND2_21615 ( P3_SUB_357_1258_U406 , P3_INSTADDRPOINTER_REG_22_ , P3_SUB_357_1258_U39 );
nand NAND2_21616 ( P3_SUB_357_1258_U407 , P3_ADD_357_U6 , P3_SUB_357_1258_U46 );
nand NAND2_21617 ( P3_SUB_357_1258_U408 , P3_INSTADDRPOINTER_REG_22_ , P3_SUB_357_1258_U39 );
nand NAND2_21618 ( P3_SUB_357_1258_U409 , P3_ADD_357_U6 , P3_SUB_357_1258_U46 );
nand NAND2_21619 ( P3_SUB_357_1258_U410 , P3_SUB_357_1258_U409 , P3_SUB_357_1258_U408 );
nand NAND2_21620 ( P3_SUB_357_1258_U411 , P3_SUB_357_1258_U136 , P3_SUB_357_1258_U137 );
nand NAND2_21621 ( P3_SUB_357_1258_U412 , P3_SUB_357_1258_U279 , P3_SUB_357_1258_U410 );
nand NAND2_21622 ( P3_SUB_357_1258_U413 , P3_INSTADDRPOINTER_REG_21_ , P3_SUB_357_1258_U39 );
nand NAND2_21623 ( P3_SUB_357_1258_U414 , P3_ADD_357_U6 , P3_SUB_357_1258_U48 );
nand NAND2_21624 ( P3_SUB_357_1258_U415 , P3_INSTADDRPOINTER_REG_21_ , P3_SUB_357_1258_U39 );
nand NAND2_21625 ( P3_SUB_357_1258_U416 , P3_ADD_357_U6 , P3_SUB_357_1258_U48 );
nand NAND2_21626 ( P3_SUB_357_1258_U417 , P3_SUB_357_1258_U416 , P3_SUB_357_1258_U415 );
nand NAND2_21627 ( P3_SUB_357_1258_U418 , P3_SUB_357_1258_U138 , P3_SUB_357_1258_U139 );
nand NAND2_21628 ( P3_SUB_357_1258_U419 , P3_SUB_357_1258_U238 , P3_SUB_357_1258_U417 );
nand NAND2_21629 ( P3_SUB_357_1258_U420 , P3_INSTADDRPOINTER_REG_20_ , P3_SUB_357_1258_U39 );
nand NAND2_21630 ( P3_SUB_357_1258_U421 , P3_ADD_357_U6 , P3_SUB_357_1258_U239 );
nand NAND2_21631 ( P3_SUB_357_1258_U422 , P3_INSTADDRPOINTER_REG_1_ , P3_SUB_357_1258_U30 );
nand NAND2_21632 ( P3_SUB_357_1258_U423 , P3_SUB_357_1258_U161 , P3_SUB_357_1258_U34 );
nand NAND2_21633 ( P3_SUB_357_1258_U424 , P3_SUB_357_1258_U423 , P3_SUB_357_1258_U422 );
nand NAND3_21634 ( P3_SUB_357_1258_U425 , P3_SUB_357_1258_U30 , P3_SUB_357_1258_U34 , P3_SUB_357_U7 );
nand NAND2_21635 ( P3_SUB_357_1258_U426 , P3_SUB_357_1258_U424 , P3_SUB_357_1258_U31 );
nand NAND2_21636 ( P3_SUB_357_1258_U427 , P3_INSTADDRPOINTER_REG_19_ , P3_SUB_357_1258_U39 );
nand NAND2_21637 ( P3_SUB_357_1258_U428 , P3_ADD_357_U6 , P3_SUB_357_1258_U47 );
nand NAND2_21638 ( P3_SUB_357_1258_U429 , P3_SUB_357_1258_U428 , P3_SUB_357_1258_U427 );
nand NAND2_21639 ( P3_SUB_357_1258_U430 , P3_SUB_357_1258_U64 , P3_SUB_357_1258_U263 );
nand NAND2_21640 ( P3_SUB_357_1258_U431 , P3_SUB_357_1258_U429 , P3_SUB_357_1258_U277 );
nand NAND2_21641 ( P3_SUB_357_1258_U432 , P3_INSTADDRPOINTER_REG_18_ , P3_SUB_357_1258_U39 );
nand NAND2_21642 ( P3_SUB_357_1258_U433 , P3_ADD_357_U6 , P3_SUB_357_1258_U49 );
nand NAND2_21643 ( P3_SUB_357_1258_U434 , P3_INSTADDRPOINTER_REG_18_ , P3_SUB_357_1258_U39 );
nand NAND2_21644 ( P3_SUB_357_1258_U435 , P3_ADD_357_U6 , P3_SUB_357_1258_U49 );
nand NAND2_21645 ( P3_SUB_357_1258_U436 , P3_SUB_357_1258_U435 , P3_SUB_357_1258_U434 );
nand NAND2_21646 ( P3_SUB_357_1258_U437 , P3_SUB_357_1258_U140 , P3_SUB_357_1258_U141 );
nand NAND2_21647 ( P3_SUB_357_1258_U438 , P3_SUB_357_1258_U203 , P3_SUB_357_1258_U436 );
nand NAND2_21648 ( P3_SUB_357_1258_U439 , P3_INSTADDRPOINTER_REG_17_ , P3_SUB_357_1258_U39 );
nand NAND2_21649 ( P3_SUB_357_1258_U440 , P3_ADD_357_U6 , P3_SUB_357_1258_U246 );
nand NAND2_21650 ( P3_SUB_357_1258_U441 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_357_U6 );
nand NAND2_21651 ( P3_SUB_357_1258_U442 , P3_SUB_357_1258_U201 , P3_SUB_357_1258_U39 );
nand NAND2_21652 ( P3_SUB_357_1258_U443 , P3_INSTADDRPOINTER_REG_16_ , P3_SUB_357_1258_U39 );
nand NAND2_21653 ( P3_SUB_357_1258_U444 , P3_ADD_357_U6 , P3_SUB_357_1258_U56 );
nand NAND2_21654 ( P3_SUB_357_1258_U445 , P3_INSTADDRPOINTER_REG_16_ , P3_SUB_357_1258_U39 );
nand NAND2_21655 ( P3_SUB_357_1258_U446 , P3_ADD_357_U6 , P3_SUB_357_1258_U56 );
nand NAND2_21656 ( P3_SUB_357_1258_U447 , P3_SUB_357_1258_U446 , P3_SUB_357_1258_U445 );
nand NAND2_21657 ( P3_SUB_357_1258_U448 , P3_SUB_357_1258_U142 , P3_SUB_357_1258_U143 );
nand NAND2_21658 ( P3_SUB_357_1258_U449 , P3_SUB_357_1258_U200 , P3_SUB_357_1258_U447 );
nand NAND2_21659 ( P3_SUB_357_1258_U450 , P3_INSTADDRPOINTER_REG_15_ , P3_SUB_357_1258_U39 );
nand NAND2_21660 ( P3_SUB_357_1258_U451 , P3_ADD_357_U6 , P3_SUB_357_1258_U55 );
nand NAND2_21661 ( P3_SUB_357_1258_U452 , P3_INSTADDRPOINTER_REG_15_ , P3_SUB_357_1258_U39 );
nand NAND2_21662 ( P3_SUB_357_1258_U453 , P3_ADD_357_U6 , P3_SUB_357_1258_U55 );
nand NAND2_21663 ( P3_SUB_357_1258_U454 , P3_SUB_357_1258_U453 , P3_SUB_357_1258_U452 );
nand NAND2_21664 ( P3_SUB_357_1258_U455 , P3_SUB_357_1258_U144 , P3_SUB_357_1258_U145 );
nand NAND2_21665 ( P3_SUB_357_1258_U456 , P3_SUB_357_1258_U196 , P3_SUB_357_1258_U454 );
nand NAND2_21666 ( P3_SUB_357_1258_U457 , P3_INSTADDRPOINTER_REG_14_ , P3_SUB_357_1258_U39 );
nand NAND2_21667 ( P3_SUB_357_1258_U458 , P3_ADD_357_U6 , P3_SUB_357_1258_U54 );
nand NAND2_21668 ( P3_SUB_357_1258_U459 , P3_INSTADDRPOINTER_REG_14_ , P3_SUB_357_1258_U39 );
nand NAND2_21669 ( P3_SUB_357_1258_U460 , P3_ADD_357_U6 , P3_SUB_357_1258_U54 );
nand NAND2_21670 ( P3_SUB_357_1258_U461 , P3_SUB_357_1258_U460 , P3_SUB_357_1258_U459 );
nand NAND2_21671 ( P3_SUB_357_1258_U462 , P3_SUB_357_1258_U146 , P3_SUB_357_1258_U147 );
nand NAND2_21672 ( P3_SUB_357_1258_U463 , P3_SUB_357_1258_U293 , P3_SUB_357_1258_U461 );
nand NAND2_21673 ( P3_SUB_357_1258_U464 , P3_INSTADDRPOINTER_REG_13_ , P3_SUB_357_1258_U39 );
nand NAND2_21674 ( P3_SUB_357_1258_U465 , P3_ADD_357_U6 , P3_SUB_357_1258_U51 );
nand NAND2_21675 ( P3_SUB_357_1258_U466 , P3_INSTADDRPOINTER_REG_12_ , P3_SUB_357_1258_U39 );
nand NAND2_21676 ( P3_SUB_357_1258_U467 , P3_ADD_357_U6 , P3_SUB_357_1258_U50 );
nand NAND2_21677 ( P3_SUB_357_1258_U468 , P3_SUB_357_1258_U467 , P3_SUB_357_1258_U466 );
nand NAND2_21678 ( P3_SUB_357_1258_U469 , P3_SUB_357_1258_U68 , P3_SUB_357_1258_U264 );
nand NAND2_21679 ( P3_SUB_357_1258_U470 , P3_SUB_357_1258_U468 , P3_SUB_357_1258_U291 );
nand NAND2_21680 ( P3_SUB_357_1258_U471 , P3_INSTADDRPOINTER_REG_11_ , P3_SUB_357_1258_U39 );
nand NAND2_21681 ( P3_SUB_357_1258_U472 , P3_ADD_357_U6 , P3_SUB_357_1258_U52 );
nand NAND2_21682 ( P3_SUB_357_1258_U473 , P3_INSTADDRPOINTER_REG_11_ , P3_SUB_357_1258_U39 );
nand NAND2_21683 ( P3_SUB_357_1258_U474 , P3_ADD_357_U6 , P3_SUB_357_1258_U52 );
nand NAND2_21684 ( P3_SUB_357_1258_U475 , P3_SUB_357_1258_U474 , P3_SUB_357_1258_U473 );
nand NAND2_21685 ( P3_SUB_357_1258_U476 , P3_SUB_357_1258_U148 , P3_SUB_357_1258_U149 );
nand NAND2_21686 ( P3_SUB_357_1258_U477 , P3_SUB_357_1258_U289 , P3_SUB_357_1258_U475 );
nand NAND2_21687 ( P3_SUB_357_1258_U478 , P3_INSTADDRPOINTER_REG_10_ , P3_SUB_357_1258_U39 );
nand NAND2_21688 ( P3_SUB_357_1258_U479 , P3_ADD_357_U6 , P3_SUB_357_1258_U53 );
nand NAND2_21689 ( P3_SUB_357_1258_U480 , P3_SUB_357_1258_U479 , P3_SUB_357_1258_U478 );
nand NAND2_21690 ( P3_SUB_357_1258_U481 , P3_SUB_357_1258_U150 , P3_SUB_357_1258_U265 );
nand NAND2_21691 ( P3_SUB_357_1258_U482 , P3_SUB_357_1258_U287 , P3_SUB_357_1258_U480 );
nand NAND2_21692 ( P3_SUB_357_1258_U483 , P3_INSTADDRPOINTER_REG_0_ , P3_SUB_357_1258_U28 );
nand NAND2_21693 ( P3_SUB_357_1258_U484 , P3_ADD_357_U10 , P3_SUB_357_1258_U29 );
not NOT1_21694 ( P3_ADD_486_U5 , P3_INSTQUEUERD_ADDR_REG_0_ );
and AND2_21695 ( P3_ADD_486_U6 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_ADD_486_U20 );
not NOT1_21696 ( P3_ADD_486_U7 , P3_INSTQUEUERD_ADDR_REG_1_ );
nand NAND2_21697 ( P3_ADD_486_U8 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_INSTQUEUERD_ADDR_REG_0_ );
not NOT1_21698 ( P3_ADD_486_U9 , P3_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_21699 ( P3_ADD_486_U10 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_ADD_486_U18 );
not NOT1_21700 ( P3_ADD_486_U11 , P3_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_21701 ( P3_ADD_486_U12 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_ADD_486_U19 );
not NOT1_21702 ( P3_ADD_486_U13 , P3_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_21703 ( P3_ADD_486_U14 , P3_ADD_486_U22 , P3_ADD_486_U21 );
nand NAND2_21704 ( P3_ADD_486_U15 , P3_ADD_486_U24 , P3_ADD_486_U23 );
nand NAND2_21705 ( P3_ADD_486_U16 , P3_ADD_486_U26 , P3_ADD_486_U25 );
nand NAND2_21706 ( P3_ADD_486_U17 , P3_ADD_486_U28 , P3_ADD_486_U27 );
not NOT1_21707 ( P3_ADD_486_U18 , P3_ADD_486_U8 );
not NOT1_21708 ( P3_ADD_486_U19 , P3_ADD_486_U10 );
not NOT1_21709 ( P3_ADD_486_U20 , P3_ADD_486_U12 );
nand NAND2_21710 ( P3_ADD_486_U21 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_ADD_486_U12 );
nand NAND2_21711 ( P3_ADD_486_U22 , P3_ADD_486_U20 , P3_ADD_486_U13 );
nand NAND2_21712 ( P3_ADD_486_U23 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_ADD_486_U10 );
nand NAND2_21713 ( P3_ADD_486_U24 , P3_ADD_486_U19 , P3_ADD_486_U11 );
nand NAND2_21714 ( P3_ADD_486_U25 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_ADD_486_U8 );
nand NAND2_21715 ( P3_ADD_486_U26 , P3_ADD_486_U18 , P3_ADD_486_U9 );
nand NAND2_21716 ( P3_ADD_486_U27 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_ADD_486_U5 );
nand NAND2_21717 ( P3_ADD_486_U28 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_ADD_486_U7 );
nand NAND2_21718 ( P3_SUB_485_U6 , P3_SUB_485_U43 , P3_SUB_485_U42 );
nand NAND2_21719 ( P3_SUB_485_U7 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_SUB_485_U27 );
not NOT1_21720 ( P3_SUB_485_U8 , P3_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_21721 ( P3_SUB_485_U9 , P3_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_21722 ( P3_SUB_485_U10 , P3_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_21723 ( P3_SUB_485_U11 , P3_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_21724 ( P3_SUB_485_U12 , P3_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_21725 ( P3_SUB_485_U13 , P3_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_21726 ( P3_SUB_485_U14 , P3_SUB_485_U39 , P3_SUB_485_U38 );
not NOT1_21727 ( P3_SUB_485_U15 , P3_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_21728 ( P3_SUB_485_U16 , P3_SUB_485_U48 , P3_SUB_485_U47 );
nand NAND2_21729 ( P3_SUB_485_U17 , P3_SUB_485_U53 , P3_SUB_485_U52 );
nand NAND2_21730 ( P3_SUB_485_U18 , P3_SUB_485_U58 , P3_SUB_485_U57 );
nand NAND2_21731 ( P3_SUB_485_U19 , P3_SUB_485_U63 , P3_SUB_485_U62 );
nand NAND2_21732 ( P3_SUB_485_U20 , P3_SUB_485_U45 , P3_SUB_485_U44 );
nand NAND2_21733 ( P3_SUB_485_U21 , P3_SUB_485_U50 , P3_SUB_485_U49 );
nand NAND2_21734 ( P3_SUB_485_U22 , P3_SUB_485_U55 , P3_SUB_485_U54 );
nand NAND2_21735 ( P3_SUB_485_U23 , P3_SUB_485_U60 , P3_SUB_485_U59 );
nand NAND2_21736 ( P3_SUB_485_U24 , P3_SUB_485_U35 , P3_SUB_485_U34 );
nand NAND2_21737 ( P3_SUB_485_U25 , P3_SUB_485_U31 , P3_SUB_485_U30 );
not NOT1_21738 ( P3_SUB_485_U26 , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_21739 ( P3_SUB_485_U27 , P3_INSTQUEUEWR_ADDR_REG_0_ );
not NOT1_21740 ( P3_SUB_485_U28 , P3_SUB_485_U7 );
nand NAND2_21741 ( P3_SUB_485_U29 , P3_SUB_485_U28 , P3_SUB_485_U8 );
nand NAND2_21742 ( P3_SUB_485_U30 , P3_SUB_485_U29 , P3_SUB_485_U26 );
nand NAND2_21743 ( P3_SUB_485_U31 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_485_U7 );
not NOT1_21744 ( P3_SUB_485_U32 , P3_SUB_485_U25 );
nand NAND2_21745 ( P3_SUB_485_U33 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_485_U10 );
nand NAND2_21746 ( P3_SUB_485_U34 , P3_SUB_485_U33 , P3_SUB_485_U25 );
nand NAND2_21747 ( P3_SUB_485_U35 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_485_U9 );
not NOT1_21748 ( P3_SUB_485_U36 , P3_SUB_485_U24 );
nand NAND2_21749 ( P3_SUB_485_U37 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_485_U12 );
nand NAND2_21750 ( P3_SUB_485_U38 , P3_SUB_485_U37 , P3_SUB_485_U24 );
nand NAND2_21751 ( P3_SUB_485_U39 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_485_U11 );
not NOT1_21752 ( P3_SUB_485_U40 , P3_SUB_485_U14 );
nand NAND2_21753 ( P3_SUB_485_U41 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_485_U15 );
nand NAND2_21754 ( P3_SUB_485_U42 , P3_SUB_485_U40 , P3_SUB_485_U41 );
nand NAND2_21755 ( P3_SUB_485_U43 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_485_U13 );
nand NAND2_21756 ( P3_SUB_485_U44 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_485_U13 );
nand NAND2_21757 ( P3_SUB_485_U45 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_485_U15 );
not NOT1_21758 ( P3_SUB_485_U46 , P3_SUB_485_U20 );
nand NAND2_21759 ( P3_SUB_485_U47 , P3_SUB_485_U46 , P3_SUB_485_U40 );
nand NAND2_21760 ( P3_SUB_485_U48 , P3_SUB_485_U20 , P3_SUB_485_U14 );
nand NAND2_21761 ( P3_SUB_485_U49 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_485_U12 );
nand NAND2_21762 ( P3_SUB_485_U50 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_485_U11 );
not NOT1_21763 ( P3_SUB_485_U51 , P3_SUB_485_U21 );
nand NAND2_21764 ( P3_SUB_485_U52 , P3_SUB_485_U36 , P3_SUB_485_U51 );
nand NAND2_21765 ( P3_SUB_485_U53 , P3_SUB_485_U21 , P3_SUB_485_U24 );
nand NAND2_21766 ( P3_SUB_485_U54 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_485_U10 );
nand NAND2_21767 ( P3_SUB_485_U55 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_485_U9 );
not NOT1_21768 ( P3_SUB_485_U56 , P3_SUB_485_U22 );
nand NAND2_21769 ( P3_SUB_485_U57 , P3_SUB_485_U32 , P3_SUB_485_U56 );
nand NAND2_21770 ( P3_SUB_485_U58 , P3_SUB_485_U22 , P3_SUB_485_U25 );
nand NAND2_21771 ( P3_SUB_485_U59 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_SUB_485_U8 );
nand NAND2_21772 ( P3_SUB_485_U60 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_485_U26 );
not NOT1_21773 ( P3_SUB_485_U61 , P3_SUB_485_U23 );
nand NAND2_21774 ( P3_SUB_485_U62 , P3_SUB_485_U61 , P3_SUB_485_U28 );
nand NAND2_21775 ( P3_SUB_485_U63 , P3_SUB_485_U23 , P3_SUB_485_U7 );
not NOT1_21776 ( P3_SUB_563_U6 , P3_U3305 );
not NOT1_21777 ( P3_SUB_563_U7 , P3_U3306 );
not NOT1_21778 ( P3_ADD_515_U4 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_21779 ( P3_ADD_515_U5 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_21780 ( P3_ADD_515_U6 , P3_INSTADDRPOINTER_REG_2_ , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_21781 ( P3_ADD_515_U7 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_21782 ( P3_ADD_515_U8 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_515_U94 );
not NOT1_21783 ( P3_ADD_515_U9 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_21784 ( P3_ADD_515_U10 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_515_U95 );
not NOT1_21785 ( P3_ADD_515_U11 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_21786 ( P3_ADD_515_U12 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_515_U96 );
not NOT1_21787 ( P3_ADD_515_U13 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_21788 ( P3_ADD_515_U14 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_515_U97 );
not NOT1_21789 ( P3_ADD_515_U15 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_21790 ( P3_ADD_515_U16 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_515_U98 );
not NOT1_21791 ( P3_ADD_515_U17 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_21792 ( P3_ADD_515_U18 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_21793 ( P3_ADD_515_U19 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_515_U99 );
nand NAND2_21794 ( P3_ADD_515_U20 , P3_ADD_515_U100 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_21795 ( P3_ADD_515_U21 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_21796 ( P3_ADD_515_U22 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_515_U101 );
not NOT1_21797 ( P3_ADD_515_U23 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_21798 ( P3_ADD_515_U24 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_515_U102 );
not NOT1_21799 ( P3_ADD_515_U25 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_21800 ( P3_ADD_515_U26 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_515_U103 );
not NOT1_21801 ( P3_ADD_515_U27 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_21802 ( P3_ADD_515_U28 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_515_U104 );
not NOT1_21803 ( P3_ADD_515_U29 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_21804 ( P3_ADD_515_U30 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_515_U105 );
not NOT1_21805 ( P3_ADD_515_U31 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_21806 ( P3_ADD_515_U32 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_515_U106 );
not NOT1_21807 ( P3_ADD_515_U33 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_21808 ( P3_ADD_515_U34 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_515_U107 );
not NOT1_21809 ( P3_ADD_515_U35 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_21810 ( P3_ADD_515_U36 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_515_U108 );
not NOT1_21811 ( P3_ADD_515_U37 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_21812 ( P3_ADD_515_U38 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_515_U109 );
not NOT1_21813 ( P3_ADD_515_U39 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_21814 ( P3_ADD_515_U40 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_515_U110 );
not NOT1_21815 ( P3_ADD_515_U41 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_21816 ( P3_ADD_515_U42 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_515_U111 );
not NOT1_21817 ( P3_ADD_515_U43 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_21818 ( P3_ADD_515_U44 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_515_U112 );
not NOT1_21819 ( P3_ADD_515_U45 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_21820 ( P3_ADD_515_U46 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_515_U113 );
not NOT1_21821 ( P3_ADD_515_U47 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_21822 ( P3_ADD_515_U48 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_515_U114 );
not NOT1_21823 ( P3_ADD_515_U49 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_21824 ( P3_ADD_515_U50 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_515_U115 );
not NOT1_21825 ( P3_ADD_515_U51 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_21826 ( P3_ADD_515_U52 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_515_U116 );
not NOT1_21827 ( P3_ADD_515_U53 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_21828 ( P3_ADD_515_U54 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_515_U117 );
not NOT1_21829 ( P3_ADD_515_U55 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_21830 ( P3_ADD_515_U56 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_515_U118 );
not NOT1_21831 ( P3_ADD_515_U57 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_21832 ( P3_ADD_515_U58 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_515_U119 );
not NOT1_21833 ( P3_ADD_515_U59 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_21834 ( P3_ADD_515_U60 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_515_U120 );
not NOT1_21835 ( P3_ADD_515_U61 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_21836 ( P3_ADD_515_U62 , P3_ADD_515_U124 , P3_ADD_515_U123 );
nand NAND2_21837 ( P3_ADD_515_U63 , P3_ADD_515_U126 , P3_ADD_515_U125 );
nand NAND2_21838 ( P3_ADD_515_U64 , P3_ADD_515_U128 , P3_ADD_515_U127 );
nand NAND2_21839 ( P3_ADD_515_U65 , P3_ADD_515_U130 , P3_ADD_515_U129 );
nand NAND2_21840 ( P3_ADD_515_U66 , P3_ADD_515_U132 , P3_ADD_515_U131 );
nand NAND2_21841 ( P3_ADD_515_U67 , P3_ADD_515_U134 , P3_ADD_515_U133 );
nand NAND2_21842 ( P3_ADD_515_U68 , P3_ADD_515_U136 , P3_ADD_515_U135 );
nand NAND2_21843 ( P3_ADD_515_U69 , P3_ADD_515_U138 , P3_ADD_515_U137 );
nand NAND2_21844 ( P3_ADD_515_U70 , P3_ADD_515_U140 , P3_ADD_515_U139 );
nand NAND2_21845 ( P3_ADD_515_U71 , P3_ADD_515_U142 , P3_ADD_515_U141 );
nand NAND2_21846 ( P3_ADD_515_U72 , P3_ADD_515_U144 , P3_ADD_515_U143 );
nand NAND2_21847 ( P3_ADD_515_U73 , P3_ADD_515_U146 , P3_ADD_515_U145 );
nand NAND2_21848 ( P3_ADD_515_U74 , P3_ADD_515_U148 , P3_ADD_515_U147 );
nand NAND2_21849 ( P3_ADD_515_U75 , P3_ADD_515_U150 , P3_ADD_515_U149 );
nand NAND2_21850 ( P3_ADD_515_U76 , P3_ADD_515_U152 , P3_ADD_515_U151 );
nand NAND2_21851 ( P3_ADD_515_U77 , P3_ADD_515_U154 , P3_ADD_515_U153 );
nand NAND2_21852 ( P3_ADD_515_U78 , P3_ADD_515_U156 , P3_ADD_515_U155 );
nand NAND2_21853 ( P3_ADD_515_U79 , P3_ADD_515_U158 , P3_ADD_515_U157 );
nand NAND2_21854 ( P3_ADD_515_U80 , P3_ADD_515_U160 , P3_ADD_515_U159 );
nand NAND2_21855 ( P3_ADD_515_U81 , P3_ADD_515_U162 , P3_ADD_515_U161 );
nand NAND2_21856 ( P3_ADD_515_U82 , P3_ADD_515_U164 , P3_ADD_515_U163 );
nand NAND2_21857 ( P3_ADD_515_U83 , P3_ADD_515_U166 , P3_ADD_515_U165 );
nand NAND2_21858 ( P3_ADD_515_U84 , P3_ADD_515_U168 , P3_ADD_515_U167 );
nand NAND2_21859 ( P3_ADD_515_U85 , P3_ADD_515_U170 , P3_ADD_515_U169 );
nand NAND2_21860 ( P3_ADD_515_U86 , P3_ADD_515_U172 , P3_ADD_515_U171 );
nand NAND2_21861 ( P3_ADD_515_U87 , P3_ADD_515_U174 , P3_ADD_515_U173 );
nand NAND2_21862 ( P3_ADD_515_U88 , P3_ADD_515_U176 , P3_ADD_515_U175 );
nand NAND2_21863 ( P3_ADD_515_U89 , P3_ADD_515_U178 , P3_ADD_515_U177 );
nand NAND2_21864 ( P3_ADD_515_U90 , P3_ADD_515_U180 , P3_ADD_515_U179 );
nand NAND2_21865 ( P3_ADD_515_U91 , P3_ADD_515_U182 , P3_ADD_515_U181 );
not NOT1_21866 ( P3_ADD_515_U92 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_21867 ( P3_ADD_515_U93 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_515_U121 );
not NOT1_21868 ( P3_ADD_515_U94 , P3_ADD_515_U6 );
not NOT1_21869 ( P3_ADD_515_U95 , P3_ADD_515_U8 );
not NOT1_21870 ( P3_ADD_515_U96 , P3_ADD_515_U10 );
not NOT1_21871 ( P3_ADD_515_U97 , P3_ADD_515_U12 );
not NOT1_21872 ( P3_ADD_515_U98 , P3_ADD_515_U14 );
not NOT1_21873 ( P3_ADD_515_U99 , P3_ADD_515_U16 );
not NOT1_21874 ( P3_ADD_515_U100 , P3_ADD_515_U19 );
not NOT1_21875 ( P3_ADD_515_U101 , P3_ADD_515_U20 );
not NOT1_21876 ( P3_ADD_515_U102 , P3_ADD_515_U22 );
not NOT1_21877 ( P3_ADD_515_U103 , P3_ADD_515_U24 );
not NOT1_21878 ( P3_ADD_515_U104 , P3_ADD_515_U26 );
not NOT1_21879 ( P3_ADD_515_U105 , P3_ADD_515_U28 );
not NOT1_21880 ( P3_ADD_515_U106 , P3_ADD_515_U30 );
not NOT1_21881 ( P3_ADD_515_U107 , P3_ADD_515_U32 );
not NOT1_21882 ( P3_ADD_515_U108 , P3_ADD_515_U34 );
not NOT1_21883 ( P3_ADD_515_U109 , P3_ADD_515_U36 );
not NOT1_21884 ( P3_ADD_515_U110 , P3_ADD_515_U38 );
not NOT1_21885 ( P3_ADD_515_U111 , P3_ADD_515_U40 );
not NOT1_21886 ( P3_ADD_515_U112 , P3_ADD_515_U42 );
not NOT1_21887 ( P3_ADD_515_U113 , P3_ADD_515_U44 );
not NOT1_21888 ( P3_ADD_515_U114 , P3_ADD_515_U46 );
not NOT1_21889 ( P3_ADD_515_U115 , P3_ADD_515_U48 );
not NOT1_21890 ( P3_ADD_515_U116 , P3_ADD_515_U50 );
not NOT1_21891 ( P3_ADD_515_U117 , P3_ADD_515_U52 );
not NOT1_21892 ( P3_ADD_515_U118 , P3_ADD_515_U54 );
not NOT1_21893 ( P3_ADD_515_U119 , P3_ADD_515_U56 );
not NOT1_21894 ( P3_ADD_515_U120 , P3_ADD_515_U58 );
not NOT1_21895 ( P3_ADD_515_U121 , P3_ADD_515_U60 );
not NOT1_21896 ( P3_ADD_515_U122 , P3_ADD_515_U93 );
nand NAND2_21897 ( P3_ADD_515_U123 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_515_U19 );
nand NAND2_21898 ( P3_ADD_515_U124 , P3_ADD_515_U100 , P3_ADD_515_U18 );
nand NAND2_21899 ( P3_ADD_515_U125 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_515_U16 );
nand NAND2_21900 ( P3_ADD_515_U126 , P3_ADD_515_U99 , P3_ADD_515_U17 );
nand NAND2_21901 ( P3_ADD_515_U127 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_515_U14 );
nand NAND2_21902 ( P3_ADD_515_U128 , P3_ADD_515_U98 , P3_ADD_515_U15 );
nand NAND2_21903 ( P3_ADD_515_U129 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_515_U12 );
nand NAND2_21904 ( P3_ADD_515_U130 , P3_ADD_515_U97 , P3_ADD_515_U13 );
nand NAND2_21905 ( P3_ADD_515_U131 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_515_U10 );
nand NAND2_21906 ( P3_ADD_515_U132 , P3_ADD_515_U96 , P3_ADD_515_U11 );
nand NAND2_21907 ( P3_ADD_515_U133 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_515_U8 );
nand NAND2_21908 ( P3_ADD_515_U134 , P3_ADD_515_U95 , P3_ADD_515_U9 );
nand NAND2_21909 ( P3_ADD_515_U135 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_515_U6 );
nand NAND2_21910 ( P3_ADD_515_U136 , P3_ADD_515_U94 , P3_ADD_515_U7 );
nand NAND2_21911 ( P3_ADD_515_U137 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_515_U93 );
nand NAND2_21912 ( P3_ADD_515_U138 , P3_ADD_515_U122 , P3_ADD_515_U92 );
nand NAND2_21913 ( P3_ADD_515_U139 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_515_U60 );
nand NAND2_21914 ( P3_ADD_515_U140 , P3_ADD_515_U121 , P3_ADD_515_U61 );
nand NAND2_21915 ( P3_ADD_515_U141 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_515_U4 );
nand NAND2_21916 ( P3_ADD_515_U142 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_515_U5 );
nand NAND2_21917 ( P3_ADD_515_U143 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_515_U58 );
nand NAND2_21918 ( P3_ADD_515_U144 , P3_ADD_515_U120 , P3_ADD_515_U59 );
nand NAND2_21919 ( P3_ADD_515_U145 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_515_U56 );
nand NAND2_21920 ( P3_ADD_515_U146 , P3_ADD_515_U119 , P3_ADD_515_U57 );
nand NAND2_21921 ( P3_ADD_515_U147 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_515_U54 );
nand NAND2_21922 ( P3_ADD_515_U148 , P3_ADD_515_U118 , P3_ADD_515_U55 );
nand NAND2_21923 ( P3_ADD_515_U149 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_515_U52 );
nand NAND2_21924 ( P3_ADD_515_U150 , P3_ADD_515_U117 , P3_ADD_515_U53 );
nand NAND2_21925 ( P3_ADD_515_U151 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_515_U50 );
nand NAND2_21926 ( P3_ADD_515_U152 , P3_ADD_515_U116 , P3_ADD_515_U51 );
nand NAND2_21927 ( P3_ADD_515_U153 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_515_U48 );
nand NAND2_21928 ( P3_ADD_515_U154 , P3_ADD_515_U115 , P3_ADD_515_U49 );
nand NAND2_21929 ( P3_ADD_515_U155 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_515_U46 );
nand NAND2_21930 ( P3_ADD_515_U156 , P3_ADD_515_U114 , P3_ADD_515_U47 );
nand NAND2_21931 ( P3_ADD_515_U157 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_515_U44 );
nand NAND2_21932 ( P3_ADD_515_U158 , P3_ADD_515_U113 , P3_ADD_515_U45 );
nand NAND2_21933 ( P3_ADD_515_U159 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_515_U42 );
nand NAND2_21934 ( P3_ADD_515_U160 , P3_ADD_515_U112 , P3_ADD_515_U43 );
nand NAND2_21935 ( P3_ADD_515_U161 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_515_U40 );
nand NAND2_21936 ( P3_ADD_515_U162 , P3_ADD_515_U111 , P3_ADD_515_U41 );
nand NAND2_21937 ( P3_ADD_515_U163 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_515_U38 );
nand NAND2_21938 ( P3_ADD_515_U164 , P3_ADD_515_U110 , P3_ADD_515_U39 );
nand NAND2_21939 ( P3_ADD_515_U165 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_515_U36 );
nand NAND2_21940 ( P3_ADD_515_U166 , P3_ADD_515_U109 , P3_ADD_515_U37 );
nand NAND2_21941 ( P3_ADD_515_U167 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_515_U34 );
nand NAND2_21942 ( P3_ADD_515_U168 , P3_ADD_515_U108 , P3_ADD_515_U35 );
nand NAND2_21943 ( P3_ADD_515_U169 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_515_U32 );
nand NAND2_21944 ( P3_ADD_515_U170 , P3_ADD_515_U107 , P3_ADD_515_U33 );
nand NAND2_21945 ( P3_ADD_515_U171 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_515_U30 );
nand NAND2_21946 ( P3_ADD_515_U172 , P3_ADD_515_U106 , P3_ADD_515_U31 );
nand NAND2_21947 ( P3_ADD_515_U173 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_515_U28 );
nand NAND2_21948 ( P3_ADD_515_U174 , P3_ADD_515_U105 , P3_ADD_515_U29 );
nand NAND2_21949 ( P3_ADD_515_U175 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_515_U26 );
nand NAND2_21950 ( P3_ADD_515_U176 , P3_ADD_515_U104 , P3_ADD_515_U27 );
nand NAND2_21951 ( P3_ADD_515_U177 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_515_U24 );
nand NAND2_21952 ( P3_ADD_515_U178 , P3_ADD_515_U103 , P3_ADD_515_U25 );
nand NAND2_21953 ( P3_ADD_515_U179 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_515_U22 );
nand NAND2_21954 ( P3_ADD_515_U180 , P3_ADD_515_U102 , P3_ADD_515_U23 );
nand NAND2_21955 ( P3_ADD_515_U181 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_515_U20 );
nand NAND2_21956 ( P3_ADD_515_U182 , P3_ADD_515_U101 , P3_ADD_515_U21 );
not NOT1_21957 ( P3_ADD_394_U4 , P3_INSTADDRPOINTER_REG_0_ );
nand NAND2_21958 ( P3_ADD_394_U5 , P3_ADD_394_U92 , P3_ADD_394_U126 );
not NOT1_21959 ( P3_ADD_394_U6 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_21960 ( P3_ADD_394_U7 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_21961 ( P3_ADD_394_U8 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_394_U92 );
not NOT1_21962 ( P3_ADD_394_U9 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_21963 ( P3_ADD_394_U10 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_394_U98 );
not NOT1_21964 ( P3_ADD_394_U11 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_21965 ( P3_ADD_394_U12 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_394_U99 );
not NOT1_21966 ( P3_ADD_394_U13 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_21967 ( P3_ADD_394_U14 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_394_U100 );
not NOT1_21968 ( P3_ADD_394_U15 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_21969 ( P3_ADD_394_U16 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_394_U101 );
not NOT1_21970 ( P3_ADD_394_U17 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_21971 ( P3_ADD_394_U18 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_21972 ( P3_ADD_394_U19 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_394_U102 );
nand NAND2_21973 ( P3_ADD_394_U20 , P3_ADD_394_U103 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_21974 ( P3_ADD_394_U21 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_21975 ( P3_ADD_394_U22 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_394_U104 );
not NOT1_21976 ( P3_ADD_394_U23 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_21977 ( P3_ADD_394_U24 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_394_U105 );
not NOT1_21978 ( P3_ADD_394_U25 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_21979 ( P3_ADD_394_U26 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_394_U106 );
not NOT1_21980 ( P3_ADD_394_U27 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_21981 ( P3_ADD_394_U28 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_394_U107 );
not NOT1_21982 ( P3_ADD_394_U29 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_21983 ( P3_ADD_394_U30 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_394_U108 );
not NOT1_21984 ( P3_ADD_394_U31 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_21985 ( P3_ADD_394_U32 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_394_U109 );
not NOT1_21986 ( P3_ADD_394_U33 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_21987 ( P3_ADD_394_U34 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_394_U110 );
not NOT1_21988 ( P3_ADD_394_U35 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_21989 ( P3_ADD_394_U36 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_394_U111 );
not NOT1_21990 ( P3_ADD_394_U37 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_21991 ( P3_ADD_394_U38 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_394_U112 );
not NOT1_21992 ( P3_ADD_394_U39 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_21993 ( P3_ADD_394_U40 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_394_U113 );
not NOT1_21994 ( P3_ADD_394_U41 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_21995 ( P3_ADD_394_U42 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_394_U114 );
not NOT1_21996 ( P3_ADD_394_U43 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_21997 ( P3_ADD_394_U44 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_394_U115 );
not NOT1_21998 ( P3_ADD_394_U45 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_21999 ( P3_ADD_394_U46 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_394_U116 );
not NOT1_22000 ( P3_ADD_394_U47 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_22001 ( P3_ADD_394_U48 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_394_U117 );
not NOT1_22002 ( P3_ADD_394_U49 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_22003 ( P3_ADD_394_U50 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_394_U118 );
not NOT1_22004 ( P3_ADD_394_U51 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_22005 ( P3_ADD_394_U52 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_394_U119 );
not NOT1_22006 ( P3_ADD_394_U53 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_22007 ( P3_ADD_394_U54 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_394_U120 );
not NOT1_22008 ( P3_ADD_394_U55 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_22009 ( P3_ADD_394_U56 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_394_U121 );
not NOT1_22010 ( P3_ADD_394_U57 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_22011 ( P3_ADD_394_U58 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_394_U122 );
not NOT1_22012 ( P3_ADD_394_U59 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_22013 ( P3_ADD_394_U60 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_394_U123 );
not NOT1_22014 ( P3_ADD_394_U61 , P3_INSTADDRPOINTER_REG_30_ );
not NOT1_22015 ( P3_ADD_394_U62 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_22016 ( P3_ADD_394_U63 , P3_ADD_394_U128 , P3_ADD_394_U127 );
nand NAND2_22017 ( P3_ADD_394_U64 , P3_ADD_394_U130 , P3_ADD_394_U129 );
nand NAND2_22018 ( P3_ADD_394_U65 , P3_ADD_394_U132 , P3_ADD_394_U131 );
nand NAND2_22019 ( P3_ADD_394_U66 , P3_ADD_394_U134 , P3_ADD_394_U133 );
nand NAND2_22020 ( P3_ADD_394_U67 , P3_ADD_394_U136 , P3_ADD_394_U135 );
nand NAND2_22021 ( P3_ADD_394_U68 , P3_ADD_394_U138 , P3_ADD_394_U137 );
nand NAND2_22022 ( P3_ADD_394_U69 , P3_ADD_394_U142 , P3_ADD_394_U141 );
nand NAND2_22023 ( P3_ADD_394_U70 , P3_ADD_394_U144 , P3_ADD_394_U143 );
nand NAND2_22024 ( P3_ADD_394_U71 , P3_ADD_394_U146 , P3_ADD_394_U145 );
nand NAND2_22025 ( P3_ADD_394_U72 , P3_ADD_394_U148 , P3_ADD_394_U147 );
nand NAND2_22026 ( P3_ADD_394_U73 , P3_ADD_394_U150 , P3_ADD_394_U149 );
nand NAND2_22027 ( P3_ADD_394_U74 , P3_ADD_394_U152 , P3_ADD_394_U151 );
nand NAND2_22028 ( P3_ADD_394_U75 , P3_ADD_394_U154 , P3_ADD_394_U153 );
nand NAND2_22029 ( P3_ADD_394_U76 , P3_ADD_394_U156 , P3_ADD_394_U155 );
nand NAND2_22030 ( P3_ADD_394_U77 , P3_ADD_394_U158 , P3_ADD_394_U157 );
nand NAND2_22031 ( P3_ADD_394_U78 , P3_ADD_394_U160 , P3_ADD_394_U159 );
nand NAND2_22032 ( P3_ADD_394_U79 , P3_ADD_394_U162 , P3_ADD_394_U161 );
nand NAND2_22033 ( P3_ADD_394_U80 , P3_ADD_394_U164 , P3_ADD_394_U163 );
nand NAND2_22034 ( P3_ADD_394_U81 , P3_ADD_394_U166 , P3_ADD_394_U165 );
nand NAND2_22035 ( P3_ADD_394_U82 , P3_ADD_394_U168 , P3_ADD_394_U167 );
nand NAND2_22036 ( P3_ADD_394_U83 , P3_ADD_394_U170 , P3_ADD_394_U169 );
nand NAND2_22037 ( P3_ADD_394_U84 , P3_ADD_394_U172 , P3_ADD_394_U171 );
nand NAND2_22038 ( P3_ADD_394_U85 , P3_ADD_394_U174 , P3_ADD_394_U173 );
nand NAND2_22039 ( P3_ADD_394_U86 , P3_ADD_394_U176 , P3_ADD_394_U175 );
nand NAND2_22040 ( P3_ADD_394_U87 , P3_ADD_394_U178 , P3_ADD_394_U177 );
nand NAND2_22041 ( P3_ADD_394_U88 , P3_ADD_394_U180 , P3_ADD_394_U179 );
nand NAND2_22042 ( P3_ADD_394_U89 , P3_ADD_394_U182 , P3_ADD_394_U181 );
nand NAND2_22043 ( P3_ADD_394_U90 , P3_ADD_394_U184 , P3_ADD_394_U183 );
nand NAND2_22044 ( P3_ADD_394_U91 , P3_ADD_394_U186 , P3_ADD_394_U185 );
nand NAND2_22045 ( P3_ADD_394_U92 , P3_ADD_394_U62 , P3_ADD_394_U96 );
and AND2_22046 ( P3_ADD_394_U93 , P3_ADD_394_U140 , P3_ADD_394_U139 );
not NOT1_22047 ( P3_ADD_394_U94 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_22048 ( P3_ADD_394_U95 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_394_U124 );
nand NAND2_22049 ( P3_ADD_394_U96 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_22050 ( P3_ADD_394_U97 , P3_ADD_394_U92 );
not NOT1_22051 ( P3_ADD_394_U98 , P3_ADD_394_U8 );
not NOT1_22052 ( P3_ADD_394_U99 , P3_ADD_394_U10 );
not NOT1_22053 ( P3_ADD_394_U100 , P3_ADD_394_U12 );
not NOT1_22054 ( P3_ADD_394_U101 , P3_ADD_394_U14 );
not NOT1_22055 ( P3_ADD_394_U102 , P3_ADD_394_U16 );
not NOT1_22056 ( P3_ADD_394_U103 , P3_ADD_394_U19 );
not NOT1_22057 ( P3_ADD_394_U104 , P3_ADD_394_U20 );
not NOT1_22058 ( P3_ADD_394_U105 , P3_ADD_394_U22 );
not NOT1_22059 ( P3_ADD_394_U106 , P3_ADD_394_U24 );
not NOT1_22060 ( P3_ADD_394_U107 , P3_ADD_394_U26 );
not NOT1_22061 ( P3_ADD_394_U108 , P3_ADD_394_U28 );
not NOT1_22062 ( P3_ADD_394_U109 , P3_ADD_394_U30 );
not NOT1_22063 ( P3_ADD_394_U110 , P3_ADD_394_U32 );
not NOT1_22064 ( P3_ADD_394_U111 , P3_ADD_394_U34 );
not NOT1_22065 ( P3_ADD_394_U112 , P3_ADD_394_U36 );
not NOT1_22066 ( P3_ADD_394_U113 , P3_ADD_394_U38 );
not NOT1_22067 ( P3_ADD_394_U114 , P3_ADD_394_U40 );
not NOT1_22068 ( P3_ADD_394_U115 , P3_ADD_394_U42 );
not NOT1_22069 ( P3_ADD_394_U116 , P3_ADD_394_U44 );
not NOT1_22070 ( P3_ADD_394_U117 , P3_ADD_394_U46 );
not NOT1_22071 ( P3_ADD_394_U118 , P3_ADD_394_U48 );
not NOT1_22072 ( P3_ADD_394_U119 , P3_ADD_394_U50 );
not NOT1_22073 ( P3_ADD_394_U120 , P3_ADD_394_U52 );
not NOT1_22074 ( P3_ADD_394_U121 , P3_ADD_394_U54 );
not NOT1_22075 ( P3_ADD_394_U122 , P3_ADD_394_U56 );
not NOT1_22076 ( P3_ADD_394_U123 , P3_ADD_394_U58 );
not NOT1_22077 ( P3_ADD_394_U124 , P3_ADD_394_U60 );
not NOT1_22078 ( P3_ADD_394_U125 , P3_ADD_394_U95 );
nand NAND3_22079 ( P3_ADD_394_U126 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_22080 ( P3_ADD_394_U127 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_394_U19 );
nand NAND2_22081 ( P3_ADD_394_U128 , P3_ADD_394_U103 , P3_ADD_394_U18 );
nand NAND2_22082 ( P3_ADD_394_U129 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_394_U16 );
nand NAND2_22083 ( P3_ADD_394_U130 , P3_ADD_394_U102 , P3_ADD_394_U17 );
nand NAND2_22084 ( P3_ADD_394_U131 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_394_U14 );
nand NAND2_22085 ( P3_ADD_394_U132 , P3_ADD_394_U101 , P3_ADD_394_U15 );
nand NAND2_22086 ( P3_ADD_394_U133 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_394_U12 );
nand NAND2_22087 ( P3_ADD_394_U134 , P3_ADD_394_U100 , P3_ADD_394_U13 );
nand NAND2_22088 ( P3_ADD_394_U135 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_394_U10 );
nand NAND2_22089 ( P3_ADD_394_U136 , P3_ADD_394_U99 , P3_ADD_394_U11 );
nand NAND2_22090 ( P3_ADD_394_U137 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_394_U8 );
nand NAND2_22091 ( P3_ADD_394_U138 , P3_ADD_394_U98 , P3_ADD_394_U9 );
nand NAND2_22092 ( P3_ADD_394_U139 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_394_U92 );
nand NAND2_22093 ( P3_ADD_394_U140 , P3_ADD_394_U97 , P3_ADD_394_U7 );
nand NAND2_22094 ( P3_ADD_394_U141 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_394_U95 );
nand NAND2_22095 ( P3_ADD_394_U142 , P3_ADD_394_U125 , P3_ADD_394_U94 );
nand NAND2_22096 ( P3_ADD_394_U143 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_394_U60 );
nand NAND2_22097 ( P3_ADD_394_U144 , P3_ADD_394_U124 , P3_ADD_394_U61 );
nand NAND2_22098 ( P3_ADD_394_U145 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_394_U58 );
nand NAND2_22099 ( P3_ADD_394_U146 , P3_ADD_394_U123 , P3_ADD_394_U59 );
nand NAND2_22100 ( P3_ADD_394_U147 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_394_U56 );
nand NAND2_22101 ( P3_ADD_394_U148 , P3_ADD_394_U122 , P3_ADD_394_U57 );
nand NAND2_22102 ( P3_ADD_394_U149 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_394_U54 );
nand NAND2_22103 ( P3_ADD_394_U150 , P3_ADD_394_U121 , P3_ADD_394_U55 );
nand NAND2_22104 ( P3_ADD_394_U151 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_394_U52 );
nand NAND2_22105 ( P3_ADD_394_U152 , P3_ADD_394_U120 , P3_ADD_394_U53 );
nand NAND2_22106 ( P3_ADD_394_U153 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_394_U50 );
nand NAND2_22107 ( P3_ADD_394_U154 , P3_ADD_394_U119 , P3_ADD_394_U51 );
nand NAND2_22108 ( P3_ADD_394_U155 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_394_U48 );
nand NAND2_22109 ( P3_ADD_394_U156 , P3_ADD_394_U118 , P3_ADD_394_U49 );
nand NAND2_22110 ( P3_ADD_394_U157 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_394_U46 );
nand NAND2_22111 ( P3_ADD_394_U158 , P3_ADD_394_U117 , P3_ADD_394_U47 );
nand NAND2_22112 ( P3_ADD_394_U159 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_394_U44 );
nand NAND2_22113 ( P3_ADD_394_U160 , P3_ADD_394_U116 , P3_ADD_394_U45 );
nand NAND2_22114 ( P3_ADD_394_U161 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_394_U42 );
nand NAND2_22115 ( P3_ADD_394_U162 , P3_ADD_394_U115 , P3_ADD_394_U43 );
nand NAND2_22116 ( P3_ADD_394_U163 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_394_U40 );
nand NAND2_22117 ( P3_ADD_394_U164 , P3_ADD_394_U114 , P3_ADD_394_U41 );
nand NAND2_22118 ( P3_ADD_394_U165 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_394_U4 );
nand NAND2_22119 ( P3_ADD_394_U166 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_394_U6 );
nand NAND2_22120 ( P3_ADD_394_U167 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_394_U38 );
nand NAND2_22121 ( P3_ADD_394_U168 , P3_ADD_394_U113 , P3_ADD_394_U39 );
nand NAND2_22122 ( P3_ADD_394_U169 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_394_U36 );
nand NAND2_22123 ( P3_ADD_394_U170 , P3_ADD_394_U112 , P3_ADD_394_U37 );
nand NAND2_22124 ( P3_ADD_394_U171 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_394_U34 );
nand NAND2_22125 ( P3_ADD_394_U172 , P3_ADD_394_U111 , P3_ADD_394_U35 );
nand NAND2_22126 ( P3_ADD_394_U173 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_394_U32 );
nand NAND2_22127 ( P3_ADD_394_U174 , P3_ADD_394_U110 , P3_ADD_394_U33 );
nand NAND2_22128 ( P3_ADD_394_U175 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_394_U30 );
nand NAND2_22129 ( P3_ADD_394_U176 , P3_ADD_394_U109 , P3_ADD_394_U31 );
nand NAND2_22130 ( P3_ADD_394_U177 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_394_U28 );
nand NAND2_22131 ( P3_ADD_394_U178 , P3_ADD_394_U108 , P3_ADD_394_U29 );
nand NAND2_22132 ( P3_ADD_394_U179 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_394_U26 );
nand NAND2_22133 ( P3_ADD_394_U180 , P3_ADD_394_U107 , P3_ADD_394_U27 );
nand NAND2_22134 ( P3_ADD_394_U181 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_394_U24 );
nand NAND2_22135 ( P3_ADD_394_U182 , P3_ADD_394_U106 , P3_ADD_394_U25 );
nand NAND2_22136 ( P3_ADD_394_U183 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_394_U22 );
nand NAND2_22137 ( P3_ADD_394_U184 , P3_ADD_394_U105 , P3_ADD_394_U23 );
nand NAND2_22138 ( P3_ADD_394_U185 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_394_U20 );
nand NAND2_22139 ( P3_ADD_394_U186 , P3_ADD_394_U104 , P3_ADD_394_U21 );
nor nor_22140 ( P3_GTE_450_U6 , P3_SUB_450_U6 , P3_GTE_450_U7 );
nor nor_22141 ( P3_GTE_450_U7 , P3_SUB_450_U16 , P3_SUB_450_U17 , P3_SUB_450_U19 , P3_SUB_450_U18 );
and AND2_22142 ( P3_SUB_414_U6 , P3_SUB_414_U126 , P3_SUB_414_U28 );
and AND2_22143 ( P3_SUB_414_U7 , P3_SUB_414_U124 , P3_SUB_414_U29 );
and AND2_22144 ( P3_SUB_414_U8 , P3_SUB_414_U122 , P3_SUB_414_U30 );
and AND2_22145 ( P3_SUB_414_U9 , P3_SUB_414_U120 , P3_SUB_414_U31 );
and AND2_22146 ( P3_SUB_414_U10 , P3_SUB_414_U118 , P3_SUB_414_U32 );
and AND2_22147 ( P3_SUB_414_U11 , P3_SUB_414_U116 , P3_SUB_414_U33 );
and AND2_22148 ( P3_SUB_414_U12 , P3_SUB_414_U114 , P3_SUB_414_U34 );
and AND2_22149 ( P3_SUB_414_U13 , P3_SUB_414_U112 , P3_SUB_414_U35 );
and AND2_22150 ( P3_SUB_414_U14 , P3_SUB_414_U110 , P3_SUB_414_U36 );
and AND2_22151 ( P3_SUB_414_U15 , P3_SUB_414_U108 , P3_SUB_414_U37 );
and AND2_22152 ( P3_SUB_414_U16 , P3_SUB_414_U106 , P3_SUB_414_U38 );
and AND2_22153 ( P3_SUB_414_U17 , P3_SUB_414_U105 , P3_SUB_414_U21 );
and AND2_22154 ( P3_SUB_414_U18 , P3_SUB_414_U92 , P3_SUB_414_U22 );
and AND2_22155 ( P3_SUB_414_U19 , P3_SUB_414_U90 , P3_SUB_414_U23 );
and AND2_22156 ( P3_SUB_414_U20 , P3_SUB_414_U88 , P3_SUB_414_U24 );
or OR3_22157 ( P3_SUB_414_U21 , P3_EBX_REG_1_ , P3_EBX_REG_0_ , P3_EBX_REG_2_ );
nand NAND3_22158 ( P3_SUB_414_U22 , P3_SUB_414_U27 , P3_SUB_414_U58 , P3_SUB_414_U83 );
nand NAND3_22159 ( P3_SUB_414_U23 , P3_SUB_414_U26 , P3_SUB_414_U56 , P3_SUB_414_U84 );
nand NAND3_22160 ( P3_SUB_414_U24 , P3_SUB_414_U25 , P3_SUB_414_U54 , P3_SUB_414_U85 );
not NOT1_22161 ( P3_SUB_414_U25 , P3_EBX_REG_8_ );
not NOT1_22162 ( P3_SUB_414_U26 , P3_EBX_REG_6_ );
not NOT1_22163 ( P3_SUB_414_U27 , P3_EBX_REG_4_ );
nand NAND3_22164 ( P3_SUB_414_U28 , P3_SUB_414_U52 , P3_SUB_414_U49 , P3_SUB_414_U86 );
nand NAND3_22165 ( P3_SUB_414_U29 , P3_SUB_414_U48 , P3_SUB_414_U81 , P3_SUB_414_U93 );
nand NAND3_22166 ( P3_SUB_414_U30 , P3_SUB_414_U47 , P3_SUB_414_U79 , P3_SUB_414_U94 );
nand NAND3_22167 ( P3_SUB_414_U31 , P3_SUB_414_U46 , P3_SUB_414_U77 , P3_SUB_414_U95 );
nand NAND3_22168 ( P3_SUB_414_U32 , P3_SUB_414_U45 , P3_SUB_414_U75 , P3_SUB_414_U96 );
nand NAND3_22169 ( P3_SUB_414_U33 , P3_SUB_414_U44 , P3_SUB_414_U73 , P3_SUB_414_U97 );
nand NAND3_22170 ( P3_SUB_414_U34 , P3_SUB_414_U43 , P3_SUB_414_U69 , P3_SUB_414_U98 );
nand NAND3_22171 ( P3_SUB_414_U35 , P3_SUB_414_U42 , P3_SUB_414_U67 , P3_SUB_414_U99 );
nand NAND3_22172 ( P3_SUB_414_U36 , P3_SUB_414_U41 , P3_SUB_414_U65 , P3_SUB_414_U100 );
nand NAND3_22173 ( P3_SUB_414_U37 , P3_SUB_414_U40 , P3_SUB_414_U63 , P3_SUB_414_U101 );
nand NAND2_22174 ( P3_SUB_414_U38 , P3_SUB_414_U102 , P3_SUB_414_U39 );
not NOT1_22175 ( P3_SUB_414_U39 , P3_EBX_REG_29_ );
not NOT1_22176 ( P3_SUB_414_U40 , P3_EBX_REG_28_ );
not NOT1_22177 ( P3_SUB_414_U41 , P3_EBX_REG_26_ );
not NOT1_22178 ( P3_SUB_414_U42 , P3_EBX_REG_24_ );
not NOT1_22179 ( P3_SUB_414_U43 , P3_EBX_REG_22_ );
not NOT1_22180 ( P3_SUB_414_U44 , P3_EBX_REG_20_ );
not NOT1_22181 ( P3_SUB_414_U45 , P3_EBX_REG_18_ );
not NOT1_22182 ( P3_SUB_414_U46 , P3_EBX_REG_16_ );
not NOT1_22183 ( P3_SUB_414_U47 , P3_EBX_REG_14_ );
not NOT1_22184 ( P3_SUB_414_U48 , P3_EBX_REG_12_ );
not NOT1_22185 ( P3_SUB_414_U49 , P3_EBX_REG_10_ );
nand NAND2_22186 ( P3_SUB_414_U50 , P3_SUB_414_U149 , P3_SUB_414_U148 );
nand NAND2_22187 ( P3_SUB_414_U51 , P3_SUB_414_U137 , P3_SUB_414_U136 );
not NOT1_22188 ( P3_SUB_414_U52 , P3_EBX_REG_9_ );
and AND2_22189 ( P3_SUB_414_U53 , P3_SUB_414_U129 , P3_SUB_414_U128 );
not NOT1_22190 ( P3_SUB_414_U54 , P3_EBX_REG_7_ );
and AND2_22191 ( P3_SUB_414_U55 , P3_SUB_414_U131 , P3_SUB_414_U130 );
not NOT1_22192 ( P3_SUB_414_U56 , P3_EBX_REG_5_ );
and AND2_22193 ( P3_SUB_414_U57 , P3_SUB_414_U133 , P3_SUB_414_U132 );
not NOT1_22194 ( P3_SUB_414_U58 , P3_EBX_REG_3_ );
and AND2_22195 ( P3_SUB_414_U59 , P3_SUB_414_U135 , P3_SUB_414_U134 );
not NOT1_22196 ( P3_SUB_414_U60 , P3_EBX_REG_31_ );
not NOT1_22197 ( P3_SUB_414_U61 , P3_EBX_REG_30_ );
and AND2_22198 ( P3_SUB_414_U62 , P3_SUB_414_U139 , P3_SUB_414_U138 );
not NOT1_22199 ( P3_SUB_414_U63 , P3_EBX_REG_27_ );
and AND2_22200 ( P3_SUB_414_U64 , P3_SUB_414_U141 , P3_SUB_414_U140 );
not NOT1_22201 ( P3_SUB_414_U65 , P3_EBX_REG_25_ );
and AND2_22202 ( P3_SUB_414_U66 , P3_SUB_414_U143 , P3_SUB_414_U142 );
not NOT1_22203 ( P3_SUB_414_U67 , P3_EBX_REG_23_ );
and AND2_22204 ( P3_SUB_414_U68 , P3_SUB_414_U145 , P3_SUB_414_U144 );
not NOT1_22205 ( P3_SUB_414_U69 , P3_EBX_REG_21_ );
and AND2_22206 ( P3_SUB_414_U70 , P3_SUB_414_U147 , P3_SUB_414_U146 );
not NOT1_22207 ( P3_SUB_414_U71 , P3_EBX_REG_1_ );
not NOT1_22208 ( P3_SUB_414_U72 , P3_EBX_REG_0_ );
not NOT1_22209 ( P3_SUB_414_U73 , P3_EBX_REG_19_ );
and AND2_22210 ( P3_SUB_414_U74 , P3_SUB_414_U151 , P3_SUB_414_U150 );
not NOT1_22211 ( P3_SUB_414_U75 , P3_EBX_REG_17_ );
and AND2_22212 ( P3_SUB_414_U76 , P3_SUB_414_U153 , P3_SUB_414_U152 );
not NOT1_22213 ( P3_SUB_414_U77 , P3_EBX_REG_15_ );
and AND2_22214 ( P3_SUB_414_U78 , P3_SUB_414_U155 , P3_SUB_414_U154 );
not NOT1_22215 ( P3_SUB_414_U79 , P3_EBX_REG_13_ );
and AND2_22216 ( P3_SUB_414_U80 , P3_SUB_414_U157 , P3_SUB_414_U156 );
not NOT1_22217 ( P3_SUB_414_U81 , P3_EBX_REG_11_ );
and AND2_22218 ( P3_SUB_414_U82 , P3_SUB_414_U159 , P3_SUB_414_U158 );
not NOT1_22219 ( P3_SUB_414_U83 , P3_SUB_414_U21 );
not NOT1_22220 ( P3_SUB_414_U84 , P3_SUB_414_U22 );
not NOT1_22221 ( P3_SUB_414_U85 , P3_SUB_414_U23 );
not NOT1_22222 ( P3_SUB_414_U86 , P3_SUB_414_U24 );
nand NAND2_22223 ( P3_SUB_414_U87 , P3_SUB_414_U85 , P3_SUB_414_U54 );
nand NAND2_22224 ( P3_SUB_414_U88 , P3_EBX_REG_8_ , P3_SUB_414_U87 );
nand NAND2_22225 ( P3_SUB_414_U89 , P3_SUB_414_U84 , P3_SUB_414_U56 );
nand NAND2_22226 ( P3_SUB_414_U90 , P3_EBX_REG_6_ , P3_SUB_414_U89 );
nand NAND2_22227 ( P3_SUB_414_U91 , P3_SUB_414_U83 , P3_SUB_414_U58 );
nand NAND2_22228 ( P3_SUB_414_U92 , P3_EBX_REG_4_ , P3_SUB_414_U91 );
not NOT1_22229 ( P3_SUB_414_U93 , P3_SUB_414_U28 );
not NOT1_22230 ( P3_SUB_414_U94 , P3_SUB_414_U29 );
not NOT1_22231 ( P3_SUB_414_U95 , P3_SUB_414_U30 );
not NOT1_22232 ( P3_SUB_414_U96 , P3_SUB_414_U31 );
not NOT1_22233 ( P3_SUB_414_U97 , P3_SUB_414_U32 );
not NOT1_22234 ( P3_SUB_414_U98 , P3_SUB_414_U33 );
not NOT1_22235 ( P3_SUB_414_U99 , P3_SUB_414_U34 );
not NOT1_22236 ( P3_SUB_414_U100 , P3_SUB_414_U35 );
not NOT1_22237 ( P3_SUB_414_U101 , P3_SUB_414_U36 );
not NOT1_22238 ( P3_SUB_414_U102 , P3_SUB_414_U37 );
not NOT1_22239 ( P3_SUB_414_U103 , P3_SUB_414_U38 );
or OR2_22240 ( P3_SUB_414_U104 , P3_EBX_REG_1_ , P3_EBX_REG_0_ );
nand NAND2_22241 ( P3_SUB_414_U105 , P3_EBX_REG_2_ , P3_SUB_414_U104 );
nand NAND2_22242 ( P3_SUB_414_U106 , P3_EBX_REG_29_ , P3_SUB_414_U37 );
nand NAND2_22243 ( P3_SUB_414_U107 , P3_SUB_414_U101 , P3_SUB_414_U63 );
nand NAND2_22244 ( P3_SUB_414_U108 , P3_EBX_REG_28_ , P3_SUB_414_U107 );
nand NAND2_22245 ( P3_SUB_414_U109 , P3_SUB_414_U100 , P3_SUB_414_U65 );
nand NAND2_22246 ( P3_SUB_414_U110 , P3_EBX_REG_26_ , P3_SUB_414_U109 );
nand NAND2_22247 ( P3_SUB_414_U111 , P3_SUB_414_U99 , P3_SUB_414_U67 );
nand NAND2_22248 ( P3_SUB_414_U112 , P3_EBX_REG_24_ , P3_SUB_414_U111 );
nand NAND2_22249 ( P3_SUB_414_U113 , P3_SUB_414_U98 , P3_SUB_414_U69 );
nand NAND2_22250 ( P3_SUB_414_U114 , P3_EBX_REG_22_ , P3_SUB_414_U113 );
nand NAND2_22251 ( P3_SUB_414_U115 , P3_SUB_414_U97 , P3_SUB_414_U73 );
nand NAND2_22252 ( P3_SUB_414_U116 , P3_EBX_REG_20_ , P3_SUB_414_U115 );
nand NAND2_22253 ( P3_SUB_414_U117 , P3_SUB_414_U96 , P3_SUB_414_U75 );
nand NAND2_22254 ( P3_SUB_414_U118 , P3_EBX_REG_18_ , P3_SUB_414_U117 );
nand NAND2_22255 ( P3_SUB_414_U119 , P3_SUB_414_U95 , P3_SUB_414_U77 );
nand NAND2_22256 ( P3_SUB_414_U120 , P3_EBX_REG_16_ , P3_SUB_414_U119 );
nand NAND2_22257 ( P3_SUB_414_U121 , P3_SUB_414_U94 , P3_SUB_414_U79 );
nand NAND2_22258 ( P3_SUB_414_U122 , P3_EBX_REG_14_ , P3_SUB_414_U121 );
nand NAND2_22259 ( P3_SUB_414_U123 , P3_SUB_414_U93 , P3_SUB_414_U81 );
nand NAND2_22260 ( P3_SUB_414_U124 , P3_EBX_REG_12_ , P3_SUB_414_U123 );
nand NAND2_22261 ( P3_SUB_414_U125 , P3_SUB_414_U86 , P3_SUB_414_U52 );
nand NAND2_22262 ( P3_SUB_414_U126 , P3_EBX_REG_10_ , P3_SUB_414_U125 );
nand NAND2_22263 ( P3_SUB_414_U127 , P3_SUB_414_U103 , P3_SUB_414_U61 );
nand NAND2_22264 ( P3_SUB_414_U128 , P3_EBX_REG_9_ , P3_SUB_414_U24 );
nand NAND2_22265 ( P3_SUB_414_U129 , P3_SUB_414_U86 , P3_SUB_414_U52 );
nand NAND2_22266 ( P3_SUB_414_U130 , P3_EBX_REG_7_ , P3_SUB_414_U23 );
nand NAND2_22267 ( P3_SUB_414_U131 , P3_SUB_414_U85 , P3_SUB_414_U54 );
nand NAND2_22268 ( P3_SUB_414_U132 , P3_EBX_REG_5_ , P3_SUB_414_U22 );
nand NAND2_22269 ( P3_SUB_414_U133 , P3_SUB_414_U84 , P3_SUB_414_U56 );
nand NAND2_22270 ( P3_SUB_414_U134 , P3_EBX_REG_3_ , P3_SUB_414_U21 );
nand NAND2_22271 ( P3_SUB_414_U135 , P3_SUB_414_U83 , P3_SUB_414_U58 );
nand NAND2_22272 ( P3_SUB_414_U136 , P3_SUB_414_U127 , P3_SUB_414_U60 );
nand NAND3_22273 ( P3_SUB_414_U137 , P3_SUB_414_U103 , P3_SUB_414_U61 , P3_EBX_REG_31_ );
nand NAND2_22274 ( P3_SUB_414_U138 , P3_EBX_REG_30_ , P3_SUB_414_U38 );
nand NAND2_22275 ( P3_SUB_414_U139 , P3_SUB_414_U103 , P3_SUB_414_U61 );
nand NAND2_22276 ( P3_SUB_414_U140 , P3_EBX_REG_27_ , P3_SUB_414_U36 );
nand NAND2_22277 ( P3_SUB_414_U141 , P3_SUB_414_U101 , P3_SUB_414_U63 );
nand NAND2_22278 ( P3_SUB_414_U142 , P3_EBX_REG_25_ , P3_SUB_414_U35 );
nand NAND2_22279 ( P3_SUB_414_U143 , P3_SUB_414_U100 , P3_SUB_414_U65 );
nand NAND2_22280 ( P3_SUB_414_U144 , P3_EBX_REG_23_ , P3_SUB_414_U34 );
nand NAND2_22281 ( P3_SUB_414_U145 , P3_SUB_414_U99 , P3_SUB_414_U67 );
nand NAND2_22282 ( P3_SUB_414_U146 , P3_EBX_REG_21_ , P3_SUB_414_U33 );
nand NAND2_22283 ( P3_SUB_414_U147 , P3_SUB_414_U98 , P3_SUB_414_U69 );
nand NAND2_22284 ( P3_SUB_414_U148 , P3_EBX_REG_1_ , P3_SUB_414_U72 );
nand NAND2_22285 ( P3_SUB_414_U149 , P3_EBX_REG_0_ , P3_SUB_414_U71 );
nand NAND2_22286 ( P3_SUB_414_U150 , P3_EBX_REG_19_ , P3_SUB_414_U32 );
nand NAND2_22287 ( P3_SUB_414_U151 , P3_SUB_414_U97 , P3_SUB_414_U73 );
nand NAND2_22288 ( P3_SUB_414_U152 , P3_EBX_REG_17_ , P3_SUB_414_U31 );
nand NAND2_22289 ( P3_SUB_414_U153 , P3_SUB_414_U96 , P3_SUB_414_U75 );
nand NAND2_22290 ( P3_SUB_414_U154 , P3_EBX_REG_15_ , P3_SUB_414_U30 );
nand NAND2_22291 ( P3_SUB_414_U155 , P3_SUB_414_U95 , P3_SUB_414_U77 );
nand NAND2_22292 ( P3_SUB_414_U156 , P3_EBX_REG_13_ , P3_SUB_414_U29 );
nand NAND2_22293 ( P3_SUB_414_U157 , P3_SUB_414_U94 , P3_SUB_414_U79 );
nand NAND2_22294 ( P3_SUB_414_U158 , P3_EBX_REG_11_ , P3_SUB_414_U28 );
nand NAND2_22295 ( P3_SUB_414_U159 , P3_SUB_414_U93 , P3_SUB_414_U81 );
not NOT1_22296 ( P3_ADD_441_U4 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_22297 ( P3_ADD_441_U5 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_22298 ( P3_ADD_441_U6 , P3_INSTADDRPOINTER_REG_2_ , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_22299 ( P3_ADD_441_U7 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_22300 ( P3_ADD_441_U8 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_441_U94 );
not NOT1_22301 ( P3_ADD_441_U9 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_22302 ( P3_ADD_441_U10 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_441_U95 );
not NOT1_22303 ( P3_ADD_441_U11 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_22304 ( P3_ADD_441_U12 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_441_U96 );
not NOT1_22305 ( P3_ADD_441_U13 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_22306 ( P3_ADD_441_U14 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_441_U97 );
not NOT1_22307 ( P3_ADD_441_U15 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_22308 ( P3_ADD_441_U16 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_441_U98 );
not NOT1_22309 ( P3_ADD_441_U17 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_22310 ( P3_ADD_441_U18 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_22311 ( P3_ADD_441_U19 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_441_U99 );
nand NAND2_22312 ( P3_ADD_441_U20 , P3_ADD_441_U100 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_22313 ( P3_ADD_441_U21 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_22314 ( P3_ADD_441_U22 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_441_U101 );
not NOT1_22315 ( P3_ADD_441_U23 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_22316 ( P3_ADD_441_U24 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_441_U102 );
not NOT1_22317 ( P3_ADD_441_U25 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_22318 ( P3_ADD_441_U26 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_441_U103 );
not NOT1_22319 ( P3_ADD_441_U27 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_22320 ( P3_ADD_441_U28 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_441_U104 );
not NOT1_22321 ( P3_ADD_441_U29 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_22322 ( P3_ADD_441_U30 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_441_U105 );
not NOT1_22323 ( P3_ADD_441_U31 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_22324 ( P3_ADD_441_U32 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_441_U106 );
not NOT1_22325 ( P3_ADD_441_U33 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_22326 ( P3_ADD_441_U34 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_441_U107 );
not NOT1_22327 ( P3_ADD_441_U35 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_22328 ( P3_ADD_441_U36 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_441_U108 );
not NOT1_22329 ( P3_ADD_441_U37 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_22330 ( P3_ADD_441_U38 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_441_U109 );
not NOT1_22331 ( P3_ADD_441_U39 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_22332 ( P3_ADD_441_U40 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_441_U110 );
not NOT1_22333 ( P3_ADD_441_U41 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_22334 ( P3_ADD_441_U42 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_441_U111 );
not NOT1_22335 ( P3_ADD_441_U43 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_22336 ( P3_ADD_441_U44 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_441_U112 );
not NOT1_22337 ( P3_ADD_441_U45 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_22338 ( P3_ADD_441_U46 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_441_U113 );
not NOT1_22339 ( P3_ADD_441_U47 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_22340 ( P3_ADD_441_U48 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_441_U114 );
not NOT1_22341 ( P3_ADD_441_U49 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_22342 ( P3_ADD_441_U50 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_441_U115 );
not NOT1_22343 ( P3_ADD_441_U51 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_22344 ( P3_ADD_441_U52 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_441_U116 );
not NOT1_22345 ( P3_ADD_441_U53 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_22346 ( P3_ADD_441_U54 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_441_U117 );
not NOT1_22347 ( P3_ADD_441_U55 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_22348 ( P3_ADD_441_U56 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_441_U118 );
not NOT1_22349 ( P3_ADD_441_U57 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_22350 ( P3_ADD_441_U58 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_441_U119 );
not NOT1_22351 ( P3_ADD_441_U59 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_22352 ( P3_ADD_441_U60 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_441_U120 );
not NOT1_22353 ( P3_ADD_441_U61 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_22354 ( P3_ADD_441_U62 , P3_ADD_441_U124 , P3_ADD_441_U123 );
nand NAND2_22355 ( P3_ADD_441_U63 , P3_ADD_441_U126 , P3_ADD_441_U125 );
nand NAND2_22356 ( P3_ADD_441_U64 , P3_ADD_441_U128 , P3_ADD_441_U127 );
nand NAND2_22357 ( P3_ADD_441_U65 , P3_ADD_441_U130 , P3_ADD_441_U129 );
nand NAND2_22358 ( P3_ADD_441_U66 , P3_ADD_441_U132 , P3_ADD_441_U131 );
nand NAND2_22359 ( P3_ADD_441_U67 , P3_ADD_441_U134 , P3_ADD_441_U133 );
nand NAND2_22360 ( P3_ADD_441_U68 , P3_ADD_441_U136 , P3_ADD_441_U135 );
nand NAND2_22361 ( P3_ADD_441_U69 , P3_ADD_441_U138 , P3_ADD_441_U137 );
nand NAND2_22362 ( P3_ADD_441_U70 , P3_ADD_441_U140 , P3_ADD_441_U139 );
nand NAND2_22363 ( P3_ADD_441_U71 , P3_ADD_441_U142 , P3_ADD_441_U141 );
nand NAND2_22364 ( P3_ADD_441_U72 , P3_ADD_441_U144 , P3_ADD_441_U143 );
nand NAND2_22365 ( P3_ADD_441_U73 , P3_ADD_441_U146 , P3_ADD_441_U145 );
nand NAND2_22366 ( P3_ADD_441_U74 , P3_ADD_441_U148 , P3_ADD_441_U147 );
nand NAND2_22367 ( P3_ADD_441_U75 , P3_ADD_441_U150 , P3_ADD_441_U149 );
nand NAND2_22368 ( P3_ADD_441_U76 , P3_ADD_441_U152 , P3_ADD_441_U151 );
nand NAND2_22369 ( P3_ADD_441_U77 , P3_ADD_441_U154 , P3_ADD_441_U153 );
nand NAND2_22370 ( P3_ADD_441_U78 , P3_ADD_441_U156 , P3_ADD_441_U155 );
nand NAND2_22371 ( P3_ADD_441_U79 , P3_ADD_441_U158 , P3_ADD_441_U157 );
nand NAND2_22372 ( P3_ADD_441_U80 , P3_ADD_441_U160 , P3_ADD_441_U159 );
nand NAND2_22373 ( P3_ADD_441_U81 , P3_ADD_441_U162 , P3_ADD_441_U161 );
nand NAND2_22374 ( P3_ADD_441_U82 , P3_ADD_441_U164 , P3_ADD_441_U163 );
nand NAND2_22375 ( P3_ADD_441_U83 , P3_ADD_441_U166 , P3_ADD_441_U165 );
nand NAND2_22376 ( P3_ADD_441_U84 , P3_ADD_441_U168 , P3_ADD_441_U167 );
nand NAND2_22377 ( P3_ADD_441_U85 , P3_ADD_441_U170 , P3_ADD_441_U169 );
nand NAND2_22378 ( P3_ADD_441_U86 , P3_ADD_441_U172 , P3_ADD_441_U171 );
nand NAND2_22379 ( P3_ADD_441_U87 , P3_ADD_441_U174 , P3_ADD_441_U173 );
nand NAND2_22380 ( P3_ADD_441_U88 , P3_ADD_441_U176 , P3_ADD_441_U175 );
nand NAND2_22381 ( P3_ADD_441_U89 , P3_ADD_441_U178 , P3_ADD_441_U177 );
nand NAND2_22382 ( P3_ADD_441_U90 , P3_ADD_441_U180 , P3_ADD_441_U179 );
nand NAND2_22383 ( P3_ADD_441_U91 , P3_ADD_441_U182 , P3_ADD_441_U181 );
not NOT1_22384 ( P3_ADD_441_U92 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_22385 ( P3_ADD_441_U93 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_441_U121 );
not NOT1_22386 ( P3_ADD_441_U94 , P3_ADD_441_U6 );
not NOT1_22387 ( P3_ADD_441_U95 , P3_ADD_441_U8 );
not NOT1_22388 ( P3_ADD_441_U96 , P3_ADD_441_U10 );
not NOT1_22389 ( P3_ADD_441_U97 , P3_ADD_441_U12 );
not NOT1_22390 ( P3_ADD_441_U98 , P3_ADD_441_U14 );
not NOT1_22391 ( P3_ADD_441_U99 , P3_ADD_441_U16 );
not NOT1_22392 ( P3_ADD_441_U100 , P3_ADD_441_U19 );
not NOT1_22393 ( P3_ADD_441_U101 , P3_ADD_441_U20 );
not NOT1_22394 ( P3_ADD_441_U102 , P3_ADD_441_U22 );
not NOT1_22395 ( P3_ADD_441_U103 , P3_ADD_441_U24 );
not NOT1_22396 ( P3_ADD_441_U104 , P3_ADD_441_U26 );
not NOT1_22397 ( P3_ADD_441_U105 , P3_ADD_441_U28 );
not NOT1_22398 ( P3_ADD_441_U106 , P3_ADD_441_U30 );
not NOT1_22399 ( P3_ADD_441_U107 , P3_ADD_441_U32 );
not NOT1_22400 ( P3_ADD_441_U108 , P3_ADD_441_U34 );
not NOT1_22401 ( P3_ADD_441_U109 , P3_ADD_441_U36 );
not NOT1_22402 ( P3_ADD_441_U110 , P3_ADD_441_U38 );
not NOT1_22403 ( P3_ADD_441_U111 , P3_ADD_441_U40 );
not NOT1_22404 ( P3_ADD_441_U112 , P3_ADD_441_U42 );
not NOT1_22405 ( P3_ADD_441_U113 , P3_ADD_441_U44 );
not NOT1_22406 ( P3_ADD_441_U114 , P3_ADD_441_U46 );
not NOT1_22407 ( P3_ADD_441_U115 , P3_ADD_441_U48 );
not NOT1_22408 ( P3_ADD_441_U116 , P3_ADD_441_U50 );
not NOT1_22409 ( P3_ADD_441_U117 , P3_ADD_441_U52 );
not NOT1_22410 ( P3_ADD_441_U118 , P3_ADD_441_U54 );
not NOT1_22411 ( P3_ADD_441_U119 , P3_ADD_441_U56 );
not NOT1_22412 ( P3_ADD_441_U120 , P3_ADD_441_U58 );
not NOT1_22413 ( P3_ADD_441_U121 , P3_ADD_441_U60 );
not NOT1_22414 ( P3_ADD_441_U122 , P3_ADD_441_U93 );
nand NAND2_22415 ( P3_ADD_441_U123 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_441_U19 );
nand NAND2_22416 ( P3_ADD_441_U124 , P3_ADD_441_U100 , P3_ADD_441_U18 );
nand NAND2_22417 ( P3_ADD_441_U125 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_441_U16 );
nand NAND2_22418 ( P3_ADD_441_U126 , P3_ADD_441_U99 , P3_ADD_441_U17 );
nand NAND2_22419 ( P3_ADD_441_U127 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_441_U14 );
nand NAND2_22420 ( P3_ADD_441_U128 , P3_ADD_441_U98 , P3_ADD_441_U15 );
nand NAND2_22421 ( P3_ADD_441_U129 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_441_U12 );
nand NAND2_22422 ( P3_ADD_441_U130 , P3_ADD_441_U97 , P3_ADD_441_U13 );
nand NAND2_22423 ( P3_ADD_441_U131 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_441_U10 );
nand NAND2_22424 ( P3_ADD_441_U132 , P3_ADD_441_U96 , P3_ADD_441_U11 );
nand NAND2_22425 ( P3_ADD_441_U133 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_441_U8 );
nand NAND2_22426 ( P3_ADD_441_U134 , P3_ADD_441_U95 , P3_ADD_441_U9 );
nand NAND2_22427 ( P3_ADD_441_U135 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_441_U6 );
nand NAND2_22428 ( P3_ADD_441_U136 , P3_ADD_441_U94 , P3_ADD_441_U7 );
nand NAND2_22429 ( P3_ADD_441_U137 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_441_U93 );
nand NAND2_22430 ( P3_ADD_441_U138 , P3_ADD_441_U122 , P3_ADD_441_U92 );
nand NAND2_22431 ( P3_ADD_441_U139 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_441_U60 );
nand NAND2_22432 ( P3_ADD_441_U140 , P3_ADD_441_U121 , P3_ADD_441_U61 );
nand NAND2_22433 ( P3_ADD_441_U141 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_441_U4 );
nand NAND2_22434 ( P3_ADD_441_U142 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_441_U5 );
nand NAND2_22435 ( P3_ADD_441_U143 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_441_U58 );
nand NAND2_22436 ( P3_ADD_441_U144 , P3_ADD_441_U120 , P3_ADD_441_U59 );
nand NAND2_22437 ( P3_ADD_441_U145 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_441_U56 );
nand NAND2_22438 ( P3_ADD_441_U146 , P3_ADD_441_U119 , P3_ADD_441_U57 );
nand NAND2_22439 ( P3_ADD_441_U147 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_441_U54 );
nand NAND2_22440 ( P3_ADD_441_U148 , P3_ADD_441_U118 , P3_ADD_441_U55 );
nand NAND2_22441 ( P3_ADD_441_U149 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_441_U52 );
nand NAND2_22442 ( P3_ADD_441_U150 , P3_ADD_441_U117 , P3_ADD_441_U53 );
nand NAND2_22443 ( P3_ADD_441_U151 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_441_U50 );
nand NAND2_22444 ( P3_ADD_441_U152 , P3_ADD_441_U116 , P3_ADD_441_U51 );
nand NAND2_22445 ( P3_ADD_441_U153 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_441_U48 );
nand NAND2_22446 ( P3_ADD_441_U154 , P3_ADD_441_U115 , P3_ADD_441_U49 );
nand NAND2_22447 ( P3_ADD_441_U155 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_441_U46 );
nand NAND2_22448 ( P3_ADD_441_U156 , P3_ADD_441_U114 , P3_ADD_441_U47 );
nand NAND2_22449 ( P3_ADD_441_U157 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_441_U44 );
nand NAND2_22450 ( P3_ADD_441_U158 , P3_ADD_441_U113 , P3_ADD_441_U45 );
nand NAND2_22451 ( P3_ADD_441_U159 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_441_U42 );
nand NAND2_22452 ( P3_ADD_441_U160 , P3_ADD_441_U112 , P3_ADD_441_U43 );
nand NAND2_22453 ( P3_ADD_441_U161 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_441_U40 );
nand NAND2_22454 ( P3_ADD_441_U162 , P3_ADD_441_U111 , P3_ADD_441_U41 );
nand NAND2_22455 ( P3_ADD_441_U163 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_441_U38 );
nand NAND2_22456 ( P3_ADD_441_U164 , P3_ADD_441_U110 , P3_ADD_441_U39 );
nand NAND2_22457 ( P3_ADD_441_U165 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_441_U36 );
nand NAND2_22458 ( P3_ADD_441_U166 , P3_ADD_441_U109 , P3_ADD_441_U37 );
nand NAND2_22459 ( P3_ADD_441_U167 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_441_U34 );
nand NAND2_22460 ( P3_ADD_441_U168 , P3_ADD_441_U108 , P3_ADD_441_U35 );
nand NAND2_22461 ( P3_ADD_441_U169 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_441_U32 );
nand NAND2_22462 ( P3_ADD_441_U170 , P3_ADD_441_U107 , P3_ADD_441_U33 );
nand NAND2_22463 ( P3_ADD_441_U171 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_441_U30 );
nand NAND2_22464 ( P3_ADD_441_U172 , P3_ADD_441_U106 , P3_ADD_441_U31 );
nand NAND2_22465 ( P3_ADD_441_U173 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_441_U28 );
nand NAND2_22466 ( P3_ADD_441_U174 , P3_ADD_441_U105 , P3_ADD_441_U29 );
nand NAND2_22467 ( P3_ADD_441_U175 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_441_U26 );
nand NAND2_22468 ( P3_ADD_441_U176 , P3_ADD_441_U104 , P3_ADD_441_U27 );
nand NAND2_22469 ( P3_ADD_441_U177 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_441_U24 );
nand NAND2_22470 ( P3_ADD_441_U178 , P3_ADD_441_U103 , P3_ADD_441_U25 );
nand NAND2_22471 ( P3_ADD_441_U179 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_441_U22 );
nand NAND2_22472 ( P3_ADD_441_U180 , P3_ADD_441_U102 , P3_ADD_441_U23 );
nand NAND2_22473 ( P3_ADD_441_U181 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_441_U20 );
nand NAND2_22474 ( P3_ADD_441_U182 , P3_ADD_441_U101 , P3_ADD_441_U21 );
not NOT1_22475 ( P3_ADD_349_U5 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_22476 ( P3_ADD_349_U6 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_22477 ( P3_ADD_349_U7 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_22478 ( P3_ADD_349_U8 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_22479 ( P3_ADD_349_U9 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_349_U98 );
not NOT1_22480 ( P3_ADD_349_U10 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_22481 ( P3_ADD_349_U11 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_349_U99 );
not NOT1_22482 ( P3_ADD_349_U12 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_22483 ( P3_ADD_349_U13 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_349_U100 );
not NOT1_22484 ( P3_ADD_349_U14 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_22485 ( P3_ADD_349_U15 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_349_U101 );
not NOT1_22486 ( P3_ADD_349_U16 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_22487 ( P3_ADD_349_U17 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_349_U102 );
not NOT1_22488 ( P3_ADD_349_U18 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_22489 ( P3_ADD_349_U19 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_349_U103 );
not NOT1_22490 ( P3_ADD_349_U20 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_22491 ( P3_ADD_349_U21 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_22492 ( P3_ADD_349_U22 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_349_U104 );
nand NAND2_22493 ( P3_ADD_349_U23 , P3_ADD_349_U105 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_22494 ( P3_ADD_349_U24 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_22495 ( P3_ADD_349_U25 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_349_U106 );
not NOT1_22496 ( P3_ADD_349_U26 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_22497 ( P3_ADD_349_U27 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_349_U107 );
not NOT1_22498 ( P3_ADD_349_U28 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_22499 ( P3_ADD_349_U29 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_349_U108 );
not NOT1_22500 ( P3_ADD_349_U30 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_22501 ( P3_ADD_349_U31 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_349_U109 );
not NOT1_22502 ( P3_ADD_349_U32 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_22503 ( P3_ADD_349_U33 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_349_U110 );
not NOT1_22504 ( P3_ADD_349_U34 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_22505 ( P3_ADD_349_U35 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_349_U111 );
not NOT1_22506 ( P3_ADD_349_U36 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_22507 ( P3_ADD_349_U37 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_349_U112 );
not NOT1_22508 ( P3_ADD_349_U38 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_22509 ( P3_ADD_349_U39 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_349_U113 );
not NOT1_22510 ( P3_ADD_349_U40 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_22511 ( P3_ADD_349_U41 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_349_U114 );
not NOT1_22512 ( P3_ADD_349_U42 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_22513 ( P3_ADD_349_U43 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_349_U115 );
not NOT1_22514 ( P3_ADD_349_U44 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_22515 ( P3_ADD_349_U45 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_349_U116 );
not NOT1_22516 ( P3_ADD_349_U46 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_22517 ( P3_ADD_349_U47 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_349_U117 );
not NOT1_22518 ( P3_ADD_349_U48 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_22519 ( P3_ADD_349_U49 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_349_U118 );
not NOT1_22520 ( P3_ADD_349_U50 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_22521 ( P3_ADD_349_U51 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_349_U119 );
not NOT1_22522 ( P3_ADD_349_U52 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_22523 ( P3_ADD_349_U53 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_349_U120 );
not NOT1_22524 ( P3_ADD_349_U54 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_22525 ( P3_ADD_349_U55 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_349_U121 );
not NOT1_22526 ( P3_ADD_349_U56 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_22527 ( P3_ADD_349_U57 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_349_U122 );
not NOT1_22528 ( P3_ADD_349_U58 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_22529 ( P3_ADD_349_U59 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_349_U123 );
not NOT1_22530 ( P3_ADD_349_U60 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_22531 ( P3_ADD_349_U61 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_349_U124 );
not NOT1_22532 ( P3_ADD_349_U62 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_22533 ( P3_ADD_349_U63 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_349_U125 );
not NOT1_22534 ( P3_ADD_349_U64 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_22535 ( P3_ADD_349_U65 , P3_ADD_349_U129 , P3_ADD_349_U128 );
nand NAND2_22536 ( P3_ADD_349_U66 , P3_ADD_349_U131 , P3_ADD_349_U130 );
nand NAND2_22537 ( P3_ADD_349_U67 , P3_ADD_349_U133 , P3_ADD_349_U132 );
nand NAND2_22538 ( P3_ADD_349_U68 , P3_ADD_349_U135 , P3_ADD_349_U134 );
nand NAND2_22539 ( P3_ADD_349_U69 , P3_ADD_349_U137 , P3_ADD_349_U136 );
nand NAND2_22540 ( P3_ADD_349_U70 , P3_ADD_349_U139 , P3_ADD_349_U138 );
nand NAND2_22541 ( P3_ADD_349_U71 , P3_ADD_349_U141 , P3_ADD_349_U140 );
nand NAND2_22542 ( P3_ADD_349_U72 , P3_ADD_349_U143 , P3_ADD_349_U142 );
nand NAND2_22543 ( P3_ADD_349_U73 , P3_ADD_349_U145 , P3_ADD_349_U144 );
nand NAND2_22544 ( P3_ADD_349_U74 , P3_ADD_349_U147 , P3_ADD_349_U146 );
nand NAND2_22545 ( P3_ADD_349_U75 , P3_ADD_349_U149 , P3_ADD_349_U148 );
nand NAND2_22546 ( P3_ADD_349_U76 , P3_ADD_349_U151 , P3_ADD_349_U150 );
nand NAND2_22547 ( P3_ADD_349_U77 , P3_ADD_349_U153 , P3_ADD_349_U152 );
nand NAND2_22548 ( P3_ADD_349_U78 , P3_ADD_349_U155 , P3_ADD_349_U154 );
nand NAND2_22549 ( P3_ADD_349_U79 , P3_ADD_349_U157 , P3_ADD_349_U156 );
nand NAND2_22550 ( P3_ADD_349_U80 , P3_ADD_349_U159 , P3_ADD_349_U158 );
nand NAND2_22551 ( P3_ADD_349_U81 , P3_ADD_349_U161 , P3_ADD_349_U160 );
nand NAND2_22552 ( P3_ADD_349_U82 , P3_ADD_349_U163 , P3_ADD_349_U162 );
nand NAND2_22553 ( P3_ADD_349_U83 , P3_ADD_349_U165 , P3_ADD_349_U164 );
nand NAND2_22554 ( P3_ADD_349_U84 , P3_ADD_349_U167 , P3_ADD_349_U166 );
nand NAND2_22555 ( P3_ADD_349_U85 , P3_ADD_349_U169 , P3_ADD_349_U168 );
nand NAND2_22556 ( P3_ADD_349_U86 , P3_ADD_349_U171 , P3_ADD_349_U170 );
nand NAND2_22557 ( P3_ADD_349_U87 , P3_ADD_349_U173 , P3_ADD_349_U172 );
nand NAND2_22558 ( P3_ADD_349_U88 , P3_ADD_349_U175 , P3_ADD_349_U174 );
nand NAND2_22559 ( P3_ADD_349_U89 , P3_ADD_349_U177 , P3_ADD_349_U176 );
nand NAND2_22560 ( P3_ADD_349_U90 , P3_ADD_349_U179 , P3_ADD_349_U178 );
nand NAND2_22561 ( P3_ADD_349_U91 , P3_ADD_349_U181 , P3_ADD_349_U180 );
nand NAND2_22562 ( P3_ADD_349_U92 , P3_ADD_349_U183 , P3_ADD_349_U182 );
nand NAND2_22563 ( P3_ADD_349_U93 , P3_ADD_349_U185 , P3_ADD_349_U184 );
nand NAND2_22564 ( P3_ADD_349_U94 , P3_ADD_349_U187 , P3_ADD_349_U186 );
nand NAND2_22565 ( P3_ADD_349_U95 , P3_ADD_349_U189 , P3_ADD_349_U188 );
not NOT1_22566 ( P3_ADD_349_U96 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_22567 ( P3_ADD_349_U97 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_349_U126 );
not NOT1_22568 ( P3_ADD_349_U98 , P3_ADD_349_U7 );
not NOT1_22569 ( P3_ADD_349_U99 , P3_ADD_349_U9 );
not NOT1_22570 ( P3_ADD_349_U100 , P3_ADD_349_U11 );
not NOT1_22571 ( P3_ADD_349_U101 , P3_ADD_349_U13 );
not NOT1_22572 ( P3_ADD_349_U102 , P3_ADD_349_U15 );
not NOT1_22573 ( P3_ADD_349_U103 , P3_ADD_349_U17 );
not NOT1_22574 ( P3_ADD_349_U104 , P3_ADD_349_U19 );
not NOT1_22575 ( P3_ADD_349_U105 , P3_ADD_349_U22 );
not NOT1_22576 ( P3_ADD_349_U106 , P3_ADD_349_U23 );
not NOT1_22577 ( P3_ADD_349_U107 , P3_ADD_349_U25 );
not NOT1_22578 ( P3_ADD_349_U108 , P3_ADD_349_U27 );
not NOT1_22579 ( P3_ADD_349_U109 , P3_ADD_349_U29 );
not NOT1_22580 ( P3_ADD_349_U110 , P3_ADD_349_U31 );
not NOT1_22581 ( P3_ADD_349_U111 , P3_ADD_349_U33 );
not NOT1_22582 ( P3_ADD_349_U112 , P3_ADD_349_U35 );
not NOT1_22583 ( P3_ADD_349_U113 , P3_ADD_349_U37 );
not NOT1_22584 ( P3_ADD_349_U114 , P3_ADD_349_U39 );
not NOT1_22585 ( P3_ADD_349_U115 , P3_ADD_349_U41 );
not NOT1_22586 ( P3_ADD_349_U116 , P3_ADD_349_U43 );
not NOT1_22587 ( P3_ADD_349_U117 , P3_ADD_349_U45 );
not NOT1_22588 ( P3_ADD_349_U118 , P3_ADD_349_U47 );
not NOT1_22589 ( P3_ADD_349_U119 , P3_ADD_349_U49 );
not NOT1_22590 ( P3_ADD_349_U120 , P3_ADD_349_U51 );
not NOT1_22591 ( P3_ADD_349_U121 , P3_ADD_349_U53 );
not NOT1_22592 ( P3_ADD_349_U122 , P3_ADD_349_U55 );
not NOT1_22593 ( P3_ADD_349_U123 , P3_ADD_349_U57 );
not NOT1_22594 ( P3_ADD_349_U124 , P3_ADD_349_U59 );
not NOT1_22595 ( P3_ADD_349_U125 , P3_ADD_349_U61 );
not NOT1_22596 ( P3_ADD_349_U126 , P3_ADD_349_U63 );
not NOT1_22597 ( P3_ADD_349_U127 , P3_ADD_349_U97 );
nand NAND2_22598 ( P3_ADD_349_U128 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_349_U22 );
nand NAND2_22599 ( P3_ADD_349_U129 , P3_ADD_349_U105 , P3_ADD_349_U21 );
nand NAND2_22600 ( P3_ADD_349_U130 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_349_U19 );
nand NAND2_22601 ( P3_ADD_349_U131 , P3_ADD_349_U104 , P3_ADD_349_U20 );
nand NAND2_22602 ( P3_ADD_349_U132 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_349_U17 );
nand NAND2_22603 ( P3_ADD_349_U133 , P3_ADD_349_U103 , P3_ADD_349_U18 );
nand NAND2_22604 ( P3_ADD_349_U134 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_349_U15 );
nand NAND2_22605 ( P3_ADD_349_U135 , P3_ADD_349_U102 , P3_ADD_349_U16 );
nand NAND2_22606 ( P3_ADD_349_U136 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_349_U13 );
nand NAND2_22607 ( P3_ADD_349_U137 , P3_ADD_349_U101 , P3_ADD_349_U14 );
nand NAND2_22608 ( P3_ADD_349_U138 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_349_U11 );
nand NAND2_22609 ( P3_ADD_349_U139 , P3_ADD_349_U100 , P3_ADD_349_U12 );
nand NAND2_22610 ( P3_ADD_349_U140 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_349_U9 );
nand NAND2_22611 ( P3_ADD_349_U141 , P3_ADD_349_U99 , P3_ADD_349_U10 );
nand NAND2_22612 ( P3_ADD_349_U142 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_349_U97 );
nand NAND2_22613 ( P3_ADD_349_U143 , P3_ADD_349_U127 , P3_ADD_349_U96 );
nand NAND2_22614 ( P3_ADD_349_U144 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_349_U63 );
nand NAND2_22615 ( P3_ADD_349_U145 , P3_ADD_349_U126 , P3_ADD_349_U64 );
nand NAND2_22616 ( P3_ADD_349_U146 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_349_U7 );
nand NAND2_22617 ( P3_ADD_349_U147 , P3_ADD_349_U98 , P3_ADD_349_U8 );
nand NAND2_22618 ( P3_ADD_349_U148 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_349_U61 );
nand NAND2_22619 ( P3_ADD_349_U149 , P3_ADD_349_U125 , P3_ADD_349_U62 );
nand NAND2_22620 ( P3_ADD_349_U150 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_349_U59 );
nand NAND2_22621 ( P3_ADD_349_U151 , P3_ADD_349_U124 , P3_ADD_349_U60 );
nand NAND2_22622 ( P3_ADD_349_U152 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_349_U57 );
nand NAND2_22623 ( P3_ADD_349_U153 , P3_ADD_349_U123 , P3_ADD_349_U58 );
nand NAND2_22624 ( P3_ADD_349_U154 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_349_U55 );
nand NAND2_22625 ( P3_ADD_349_U155 , P3_ADD_349_U122 , P3_ADD_349_U56 );
nand NAND2_22626 ( P3_ADD_349_U156 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_349_U53 );
nand NAND2_22627 ( P3_ADD_349_U157 , P3_ADD_349_U121 , P3_ADD_349_U54 );
nand NAND2_22628 ( P3_ADD_349_U158 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_349_U51 );
nand NAND2_22629 ( P3_ADD_349_U159 , P3_ADD_349_U120 , P3_ADD_349_U52 );
nand NAND2_22630 ( P3_ADD_349_U160 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_349_U49 );
nand NAND2_22631 ( P3_ADD_349_U161 , P3_ADD_349_U119 , P3_ADD_349_U50 );
nand NAND2_22632 ( P3_ADD_349_U162 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_349_U47 );
nand NAND2_22633 ( P3_ADD_349_U163 , P3_ADD_349_U118 , P3_ADD_349_U48 );
nand NAND2_22634 ( P3_ADD_349_U164 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_349_U45 );
nand NAND2_22635 ( P3_ADD_349_U165 , P3_ADD_349_U117 , P3_ADD_349_U46 );
nand NAND2_22636 ( P3_ADD_349_U166 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_349_U43 );
nand NAND2_22637 ( P3_ADD_349_U167 , P3_ADD_349_U116 , P3_ADD_349_U44 );
nand NAND2_22638 ( P3_ADD_349_U168 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_349_U5 );
nand NAND2_22639 ( P3_ADD_349_U169 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_349_U6 );
nand NAND2_22640 ( P3_ADD_349_U170 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_349_U41 );
nand NAND2_22641 ( P3_ADD_349_U171 , P3_ADD_349_U115 , P3_ADD_349_U42 );
nand NAND2_22642 ( P3_ADD_349_U172 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_349_U39 );
nand NAND2_22643 ( P3_ADD_349_U173 , P3_ADD_349_U114 , P3_ADD_349_U40 );
nand NAND2_22644 ( P3_ADD_349_U174 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_349_U37 );
nand NAND2_22645 ( P3_ADD_349_U175 , P3_ADD_349_U113 , P3_ADD_349_U38 );
nand NAND2_22646 ( P3_ADD_349_U176 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_349_U35 );
nand NAND2_22647 ( P3_ADD_349_U177 , P3_ADD_349_U112 , P3_ADD_349_U36 );
nand NAND2_22648 ( P3_ADD_349_U178 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_349_U33 );
nand NAND2_22649 ( P3_ADD_349_U179 , P3_ADD_349_U111 , P3_ADD_349_U34 );
nand NAND2_22650 ( P3_ADD_349_U180 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_349_U31 );
nand NAND2_22651 ( P3_ADD_349_U181 , P3_ADD_349_U110 , P3_ADD_349_U32 );
nand NAND2_22652 ( P3_ADD_349_U182 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_349_U29 );
nand NAND2_22653 ( P3_ADD_349_U183 , P3_ADD_349_U109 , P3_ADD_349_U30 );
nand NAND2_22654 ( P3_ADD_349_U184 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_349_U27 );
nand NAND2_22655 ( P3_ADD_349_U185 , P3_ADD_349_U108 , P3_ADD_349_U28 );
nand NAND2_22656 ( P3_ADD_349_U186 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_349_U25 );
nand NAND2_22657 ( P3_ADD_349_U187 , P3_ADD_349_U107 , P3_ADD_349_U26 );
nand NAND2_22658 ( P3_ADD_349_U188 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_349_U23 );
nand NAND2_22659 ( P3_ADD_349_U189 , P3_ADD_349_U106 , P3_ADD_349_U24 );
not NOT1_22660 ( P3_ADD_405_U4 , P3_INSTADDRPOINTER_REG_0_ );
nand NAND2_22661 ( P3_ADD_405_U5 , P3_ADD_405_U92 , P3_ADD_405_U126 );
not NOT1_22662 ( P3_ADD_405_U6 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_22663 ( P3_ADD_405_U7 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_22664 ( P3_ADD_405_U8 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_405_U92 );
not NOT1_22665 ( P3_ADD_405_U9 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_22666 ( P3_ADD_405_U10 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_405_U98 );
not NOT1_22667 ( P3_ADD_405_U11 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_22668 ( P3_ADD_405_U12 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_405_U99 );
not NOT1_22669 ( P3_ADD_405_U13 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_22670 ( P3_ADD_405_U14 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_405_U100 );
not NOT1_22671 ( P3_ADD_405_U15 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_22672 ( P3_ADD_405_U16 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_405_U101 );
not NOT1_22673 ( P3_ADD_405_U17 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_22674 ( P3_ADD_405_U18 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_22675 ( P3_ADD_405_U19 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_405_U102 );
nand NAND2_22676 ( P3_ADD_405_U20 , P3_ADD_405_U103 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_22677 ( P3_ADD_405_U21 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_22678 ( P3_ADD_405_U22 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_405_U104 );
not NOT1_22679 ( P3_ADD_405_U23 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_22680 ( P3_ADD_405_U24 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_405_U105 );
not NOT1_22681 ( P3_ADD_405_U25 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_22682 ( P3_ADD_405_U26 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_405_U106 );
not NOT1_22683 ( P3_ADD_405_U27 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_22684 ( P3_ADD_405_U28 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_405_U107 );
not NOT1_22685 ( P3_ADD_405_U29 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_22686 ( P3_ADD_405_U30 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_405_U108 );
not NOT1_22687 ( P3_ADD_405_U31 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_22688 ( P3_ADD_405_U32 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_405_U109 );
not NOT1_22689 ( P3_ADD_405_U33 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_22690 ( P3_ADD_405_U34 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_405_U110 );
not NOT1_22691 ( P3_ADD_405_U35 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_22692 ( P3_ADD_405_U36 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_405_U111 );
not NOT1_22693 ( P3_ADD_405_U37 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_22694 ( P3_ADD_405_U38 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_405_U112 );
not NOT1_22695 ( P3_ADD_405_U39 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_22696 ( P3_ADD_405_U40 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_405_U113 );
not NOT1_22697 ( P3_ADD_405_U41 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_22698 ( P3_ADD_405_U42 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_405_U114 );
not NOT1_22699 ( P3_ADD_405_U43 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_22700 ( P3_ADD_405_U44 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_405_U115 );
not NOT1_22701 ( P3_ADD_405_U45 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_22702 ( P3_ADD_405_U46 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_405_U116 );
not NOT1_22703 ( P3_ADD_405_U47 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_22704 ( P3_ADD_405_U48 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_405_U117 );
not NOT1_22705 ( P3_ADD_405_U49 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_22706 ( P3_ADD_405_U50 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_405_U118 );
not NOT1_22707 ( P3_ADD_405_U51 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_22708 ( P3_ADD_405_U52 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_405_U119 );
not NOT1_22709 ( P3_ADD_405_U53 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_22710 ( P3_ADD_405_U54 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_405_U120 );
not NOT1_22711 ( P3_ADD_405_U55 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_22712 ( P3_ADD_405_U56 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_405_U121 );
not NOT1_22713 ( P3_ADD_405_U57 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_22714 ( P3_ADD_405_U58 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_405_U122 );
not NOT1_22715 ( P3_ADD_405_U59 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_22716 ( P3_ADD_405_U60 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_405_U123 );
not NOT1_22717 ( P3_ADD_405_U61 , P3_INSTADDRPOINTER_REG_30_ );
not NOT1_22718 ( P3_ADD_405_U62 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_22719 ( P3_ADD_405_U63 , P3_ADD_405_U128 , P3_ADD_405_U127 );
nand NAND2_22720 ( P3_ADD_405_U64 , P3_ADD_405_U130 , P3_ADD_405_U129 );
nand NAND2_22721 ( P3_ADD_405_U65 , P3_ADD_405_U132 , P3_ADD_405_U131 );
nand NAND2_22722 ( P3_ADD_405_U66 , P3_ADD_405_U134 , P3_ADD_405_U133 );
nand NAND2_22723 ( P3_ADD_405_U67 , P3_ADD_405_U136 , P3_ADD_405_U135 );
nand NAND2_22724 ( P3_ADD_405_U68 , P3_ADD_405_U138 , P3_ADD_405_U137 );
nand NAND2_22725 ( P3_ADD_405_U69 , P3_ADD_405_U142 , P3_ADD_405_U141 );
nand NAND2_22726 ( P3_ADD_405_U70 , P3_ADD_405_U144 , P3_ADD_405_U143 );
nand NAND2_22727 ( P3_ADD_405_U71 , P3_ADD_405_U146 , P3_ADD_405_U145 );
nand NAND2_22728 ( P3_ADD_405_U72 , P3_ADD_405_U148 , P3_ADD_405_U147 );
nand NAND2_22729 ( P3_ADD_405_U73 , P3_ADD_405_U150 , P3_ADD_405_U149 );
nand NAND2_22730 ( P3_ADD_405_U74 , P3_ADD_405_U152 , P3_ADD_405_U151 );
nand NAND2_22731 ( P3_ADD_405_U75 , P3_ADD_405_U154 , P3_ADD_405_U153 );
nand NAND2_22732 ( P3_ADD_405_U76 , P3_ADD_405_U156 , P3_ADD_405_U155 );
nand NAND2_22733 ( P3_ADD_405_U77 , P3_ADD_405_U158 , P3_ADD_405_U157 );
nand NAND2_22734 ( P3_ADD_405_U78 , P3_ADD_405_U160 , P3_ADD_405_U159 );
nand NAND2_22735 ( P3_ADD_405_U79 , P3_ADD_405_U162 , P3_ADD_405_U161 );
nand NAND2_22736 ( P3_ADD_405_U80 , P3_ADD_405_U164 , P3_ADD_405_U163 );
nand NAND2_22737 ( P3_ADD_405_U81 , P3_ADD_405_U166 , P3_ADD_405_U165 );
nand NAND2_22738 ( P3_ADD_405_U82 , P3_ADD_405_U168 , P3_ADD_405_U167 );
nand NAND2_22739 ( P3_ADD_405_U83 , P3_ADD_405_U170 , P3_ADD_405_U169 );
nand NAND2_22740 ( P3_ADD_405_U84 , P3_ADD_405_U172 , P3_ADD_405_U171 );
nand NAND2_22741 ( P3_ADD_405_U85 , P3_ADD_405_U174 , P3_ADD_405_U173 );
nand NAND2_22742 ( P3_ADD_405_U86 , P3_ADD_405_U176 , P3_ADD_405_U175 );
nand NAND2_22743 ( P3_ADD_405_U87 , P3_ADD_405_U178 , P3_ADD_405_U177 );
nand NAND2_22744 ( P3_ADD_405_U88 , P3_ADD_405_U180 , P3_ADD_405_U179 );
nand NAND2_22745 ( P3_ADD_405_U89 , P3_ADD_405_U182 , P3_ADD_405_U181 );
nand NAND2_22746 ( P3_ADD_405_U90 , P3_ADD_405_U184 , P3_ADD_405_U183 );
nand NAND2_22747 ( P3_ADD_405_U91 , P3_ADD_405_U186 , P3_ADD_405_U185 );
nand NAND2_22748 ( P3_ADD_405_U92 , P3_ADD_405_U62 , P3_ADD_405_U96 );
and AND2_22749 ( P3_ADD_405_U93 , P3_ADD_405_U140 , P3_ADD_405_U139 );
not NOT1_22750 ( P3_ADD_405_U94 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_22751 ( P3_ADD_405_U95 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_405_U124 );
nand NAND2_22752 ( P3_ADD_405_U96 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_22753 ( P3_ADD_405_U97 , P3_ADD_405_U92 );
not NOT1_22754 ( P3_ADD_405_U98 , P3_ADD_405_U8 );
not NOT1_22755 ( P3_ADD_405_U99 , P3_ADD_405_U10 );
not NOT1_22756 ( P3_ADD_405_U100 , P3_ADD_405_U12 );
not NOT1_22757 ( P3_ADD_405_U101 , P3_ADD_405_U14 );
not NOT1_22758 ( P3_ADD_405_U102 , P3_ADD_405_U16 );
not NOT1_22759 ( P3_ADD_405_U103 , P3_ADD_405_U19 );
not NOT1_22760 ( P3_ADD_405_U104 , P3_ADD_405_U20 );
not NOT1_22761 ( P3_ADD_405_U105 , P3_ADD_405_U22 );
not NOT1_22762 ( P3_ADD_405_U106 , P3_ADD_405_U24 );
not NOT1_22763 ( P3_ADD_405_U107 , P3_ADD_405_U26 );
not NOT1_22764 ( P3_ADD_405_U108 , P3_ADD_405_U28 );
not NOT1_22765 ( P3_ADD_405_U109 , P3_ADD_405_U30 );
not NOT1_22766 ( P3_ADD_405_U110 , P3_ADD_405_U32 );
not NOT1_22767 ( P3_ADD_405_U111 , P3_ADD_405_U34 );
not NOT1_22768 ( P3_ADD_405_U112 , P3_ADD_405_U36 );
not NOT1_22769 ( P3_ADD_405_U113 , P3_ADD_405_U38 );
not NOT1_22770 ( P3_ADD_405_U114 , P3_ADD_405_U40 );
not NOT1_22771 ( P3_ADD_405_U115 , P3_ADD_405_U42 );
not NOT1_22772 ( P3_ADD_405_U116 , P3_ADD_405_U44 );
not NOT1_22773 ( P3_ADD_405_U117 , P3_ADD_405_U46 );
not NOT1_22774 ( P3_ADD_405_U118 , P3_ADD_405_U48 );
not NOT1_22775 ( P3_ADD_405_U119 , P3_ADD_405_U50 );
not NOT1_22776 ( P3_ADD_405_U120 , P3_ADD_405_U52 );
not NOT1_22777 ( P3_ADD_405_U121 , P3_ADD_405_U54 );
not NOT1_22778 ( P3_ADD_405_U122 , P3_ADD_405_U56 );
not NOT1_22779 ( P3_ADD_405_U123 , P3_ADD_405_U58 );
not NOT1_22780 ( P3_ADD_405_U124 , P3_ADD_405_U60 );
not NOT1_22781 ( P3_ADD_405_U125 , P3_ADD_405_U95 );
nand NAND3_22782 ( P3_ADD_405_U126 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_22783 ( P3_ADD_405_U127 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_405_U19 );
nand NAND2_22784 ( P3_ADD_405_U128 , P3_ADD_405_U103 , P3_ADD_405_U18 );
nand NAND2_22785 ( P3_ADD_405_U129 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_405_U16 );
nand NAND2_22786 ( P3_ADD_405_U130 , P3_ADD_405_U102 , P3_ADD_405_U17 );
nand NAND2_22787 ( P3_ADD_405_U131 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_405_U14 );
nand NAND2_22788 ( P3_ADD_405_U132 , P3_ADD_405_U101 , P3_ADD_405_U15 );
nand NAND2_22789 ( P3_ADD_405_U133 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_405_U12 );
nand NAND2_22790 ( P3_ADD_405_U134 , P3_ADD_405_U100 , P3_ADD_405_U13 );
nand NAND2_22791 ( P3_ADD_405_U135 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_405_U10 );
nand NAND2_22792 ( P3_ADD_405_U136 , P3_ADD_405_U99 , P3_ADD_405_U11 );
nand NAND2_22793 ( P3_ADD_405_U137 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_405_U8 );
nand NAND2_22794 ( P3_ADD_405_U138 , P3_ADD_405_U98 , P3_ADD_405_U9 );
nand NAND2_22795 ( P3_ADD_405_U139 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_405_U92 );
nand NAND2_22796 ( P3_ADD_405_U140 , P3_ADD_405_U97 , P3_ADD_405_U7 );
nand NAND2_22797 ( P3_ADD_405_U141 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_405_U95 );
nand NAND2_22798 ( P3_ADD_405_U142 , P3_ADD_405_U125 , P3_ADD_405_U94 );
nand NAND2_22799 ( P3_ADD_405_U143 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_405_U60 );
nand NAND2_22800 ( P3_ADD_405_U144 , P3_ADD_405_U124 , P3_ADD_405_U61 );
nand NAND2_22801 ( P3_ADD_405_U145 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_405_U58 );
nand NAND2_22802 ( P3_ADD_405_U146 , P3_ADD_405_U123 , P3_ADD_405_U59 );
nand NAND2_22803 ( P3_ADD_405_U147 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_405_U56 );
nand NAND2_22804 ( P3_ADD_405_U148 , P3_ADD_405_U122 , P3_ADD_405_U57 );
nand NAND2_22805 ( P3_ADD_405_U149 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_405_U54 );
nand NAND2_22806 ( P3_ADD_405_U150 , P3_ADD_405_U121 , P3_ADD_405_U55 );
nand NAND2_22807 ( P3_ADD_405_U151 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_405_U52 );
nand NAND2_22808 ( P3_ADD_405_U152 , P3_ADD_405_U120 , P3_ADD_405_U53 );
nand NAND2_22809 ( P3_ADD_405_U153 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_405_U50 );
nand NAND2_22810 ( P3_ADD_405_U154 , P3_ADD_405_U119 , P3_ADD_405_U51 );
nand NAND2_22811 ( P3_ADD_405_U155 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_405_U48 );
nand NAND2_22812 ( P3_ADD_405_U156 , P3_ADD_405_U118 , P3_ADD_405_U49 );
nand NAND2_22813 ( P3_ADD_405_U157 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_405_U46 );
nand NAND2_22814 ( P3_ADD_405_U158 , P3_ADD_405_U117 , P3_ADD_405_U47 );
nand NAND2_22815 ( P3_ADD_405_U159 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_405_U44 );
nand NAND2_22816 ( P3_ADD_405_U160 , P3_ADD_405_U116 , P3_ADD_405_U45 );
nand NAND2_22817 ( P3_ADD_405_U161 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_405_U42 );
nand NAND2_22818 ( P3_ADD_405_U162 , P3_ADD_405_U115 , P3_ADD_405_U43 );
nand NAND2_22819 ( P3_ADD_405_U163 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_405_U40 );
nand NAND2_22820 ( P3_ADD_405_U164 , P3_ADD_405_U114 , P3_ADD_405_U41 );
nand NAND2_22821 ( P3_ADD_405_U165 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_405_U4 );
nand NAND2_22822 ( P3_ADD_405_U166 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_405_U6 );
nand NAND2_22823 ( P3_ADD_405_U167 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_405_U38 );
nand NAND2_22824 ( P3_ADD_405_U168 , P3_ADD_405_U113 , P3_ADD_405_U39 );
nand NAND2_22825 ( P3_ADD_405_U169 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_405_U36 );
nand NAND2_22826 ( P3_ADD_405_U170 , P3_ADD_405_U112 , P3_ADD_405_U37 );
nand NAND2_22827 ( P3_ADD_405_U171 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_405_U34 );
nand NAND2_22828 ( P3_ADD_405_U172 , P3_ADD_405_U111 , P3_ADD_405_U35 );
nand NAND2_22829 ( P3_ADD_405_U173 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_405_U32 );
nand NAND2_22830 ( P3_ADD_405_U174 , P3_ADD_405_U110 , P3_ADD_405_U33 );
nand NAND2_22831 ( P3_ADD_405_U175 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_405_U30 );
nand NAND2_22832 ( P3_ADD_405_U176 , P3_ADD_405_U109 , P3_ADD_405_U31 );
nand NAND2_22833 ( P3_ADD_405_U177 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_405_U28 );
nand NAND2_22834 ( P3_ADD_405_U178 , P3_ADD_405_U108 , P3_ADD_405_U29 );
nand NAND2_22835 ( P3_ADD_405_U179 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_405_U26 );
nand NAND2_22836 ( P3_ADD_405_U180 , P3_ADD_405_U107 , P3_ADD_405_U27 );
nand NAND2_22837 ( P3_ADD_405_U181 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_405_U24 );
nand NAND2_22838 ( P3_ADD_405_U182 , P3_ADD_405_U106 , P3_ADD_405_U25 );
nand NAND2_22839 ( P3_ADD_405_U183 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_405_U22 );
nand NAND2_22840 ( P3_ADD_405_U184 , P3_ADD_405_U105 , P3_ADD_405_U23 );
nand NAND2_22841 ( P3_ADD_405_U185 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_405_U20 );
nand NAND2_22842 ( P3_ADD_405_U186 , P3_ADD_405_U104 , P3_ADD_405_U21 );
not NOT1_22843 ( P3_ADD_553_U5 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_22844 ( P3_ADD_553_U6 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_22845 ( P3_ADD_553_U7 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_22846 ( P3_ADD_553_U8 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_22847 ( P3_ADD_553_U9 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_553_U98 );
not NOT1_22848 ( P3_ADD_553_U10 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_22849 ( P3_ADD_553_U11 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_553_U99 );
not NOT1_22850 ( P3_ADD_553_U12 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_22851 ( P3_ADD_553_U13 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_553_U100 );
not NOT1_22852 ( P3_ADD_553_U14 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_22853 ( P3_ADD_553_U15 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_553_U101 );
not NOT1_22854 ( P3_ADD_553_U16 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_22855 ( P3_ADD_553_U17 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_553_U102 );
not NOT1_22856 ( P3_ADD_553_U18 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_22857 ( P3_ADD_553_U19 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_553_U103 );
not NOT1_22858 ( P3_ADD_553_U20 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_22859 ( P3_ADD_553_U21 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_22860 ( P3_ADD_553_U22 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_553_U104 );
nand NAND2_22861 ( P3_ADD_553_U23 , P3_ADD_553_U105 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_22862 ( P3_ADD_553_U24 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_22863 ( P3_ADD_553_U25 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_553_U106 );
not NOT1_22864 ( P3_ADD_553_U26 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_22865 ( P3_ADD_553_U27 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_553_U107 );
not NOT1_22866 ( P3_ADD_553_U28 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_22867 ( P3_ADD_553_U29 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_553_U108 );
not NOT1_22868 ( P3_ADD_553_U30 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_22869 ( P3_ADD_553_U31 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_553_U109 );
not NOT1_22870 ( P3_ADD_553_U32 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_22871 ( P3_ADD_553_U33 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_553_U110 );
not NOT1_22872 ( P3_ADD_553_U34 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_22873 ( P3_ADD_553_U35 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_553_U111 );
not NOT1_22874 ( P3_ADD_553_U36 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_22875 ( P3_ADD_553_U37 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_553_U112 );
not NOT1_22876 ( P3_ADD_553_U38 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_22877 ( P3_ADD_553_U39 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_553_U113 );
not NOT1_22878 ( P3_ADD_553_U40 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_22879 ( P3_ADD_553_U41 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_553_U114 );
not NOT1_22880 ( P3_ADD_553_U42 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_22881 ( P3_ADD_553_U43 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_553_U115 );
not NOT1_22882 ( P3_ADD_553_U44 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_22883 ( P3_ADD_553_U45 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_553_U116 );
not NOT1_22884 ( P3_ADD_553_U46 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_22885 ( P3_ADD_553_U47 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_553_U117 );
not NOT1_22886 ( P3_ADD_553_U48 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_22887 ( P3_ADD_553_U49 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_553_U118 );
not NOT1_22888 ( P3_ADD_553_U50 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_22889 ( P3_ADD_553_U51 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_553_U119 );
not NOT1_22890 ( P3_ADD_553_U52 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_22891 ( P3_ADD_553_U53 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_553_U120 );
not NOT1_22892 ( P3_ADD_553_U54 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_22893 ( P3_ADD_553_U55 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_553_U121 );
not NOT1_22894 ( P3_ADD_553_U56 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_22895 ( P3_ADD_553_U57 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_553_U122 );
not NOT1_22896 ( P3_ADD_553_U58 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_22897 ( P3_ADD_553_U59 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_553_U123 );
not NOT1_22898 ( P3_ADD_553_U60 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_22899 ( P3_ADD_553_U61 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_553_U124 );
not NOT1_22900 ( P3_ADD_553_U62 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_22901 ( P3_ADD_553_U63 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_553_U125 );
not NOT1_22902 ( P3_ADD_553_U64 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_22903 ( P3_ADD_553_U65 , P3_ADD_553_U129 , P3_ADD_553_U128 );
nand NAND2_22904 ( P3_ADD_553_U66 , P3_ADD_553_U131 , P3_ADD_553_U130 );
nand NAND2_22905 ( P3_ADD_553_U67 , P3_ADD_553_U133 , P3_ADD_553_U132 );
nand NAND2_22906 ( P3_ADD_553_U68 , P3_ADD_553_U135 , P3_ADD_553_U134 );
nand NAND2_22907 ( P3_ADD_553_U69 , P3_ADD_553_U137 , P3_ADD_553_U136 );
nand NAND2_22908 ( P3_ADD_553_U70 , P3_ADD_553_U139 , P3_ADD_553_U138 );
nand NAND2_22909 ( P3_ADD_553_U71 , P3_ADD_553_U141 , P3_ADD_553_U140 );
nand NAND2_22910 ( P3_ADD_553_U72 , P3_ADD_553_U143 , P3_ADD_553_U142 );
nand NAND2_22911 ( P3_ADD_553_U73 , P3_ADD_553_U145 , P3_ADD_553_U144 );
nand NAND2_22912 ( P3_ADD_553_U74 , P3_ADD_553_U147 , P3_ADD_553_U146 );
nand NAND2_22913 ( P3_ADD_553_U75 , P3_ADD_553_U149 , P3_ADD_553_U148 );
nand NAND2_22914 ( P3_ADD_553_U76 , P3_ADD_553_U151 , P3_ADD_553_U150 );
nand NAND2_22915 ( P3_ADD_553_U77 , P3_ADD_553_U153 , P3_ADD_553_U152 );
nand NAND2_22916 ( P3_ADD_553_U78 , P3_ADD_553_U155 , P3_ADD_553_U154 );
nand NAND2_22917 ( P3_ADD_553_U79 , P3_ADD_553_U157 , P3_ADD_553_U156 );
nand NAND2_22918 ( P3_ADD_553_U80 , P3_ADD_553_U159 , P3_ADD_553_U158 );
nand NAND2_22919 ( P3_ADD_553_U81 , P3_ADD_553_U161 , P3_ADD_553_U160 );
nand NAND2_22920 ( P3_ADD_553_U82 , P3_ADD_553_U163 , P3_ADD_553_U162 );
nand NAND2_22921 ( P3_ADD_553_U83 , P3_ADD_553_U165 , P3_ADD_553_U164 );
nand NAND2_22922 ( P3_ADD_553_U84 , P3_ADD_553_U167 , P3_ADD_553_U166 );
nand NAND2_22923 ( P3_ADD_553_U85 , P3_ADD_553_U169 , P3_ADD_553_U168 );
nand NAND2_22924 ( P3_ADD_553_U86 , P3_ADD_553_U171 , P3_ADD_553_U170 );
nand NAND2_22925 ( P3_ADD_553_U87 , P3_ADD_553_U173 , P3_ADD_553_U172 );
nand NAND2_22926 ( P3_ADD_553_U88 , P3_ADD_553_U175 , P3_ADD_553_U174 );
nand NAND2_22927 ( P3_ADD_553_U89 , P3_ADD_553_U177 , P3_ADD_553_U176 );
nand NAND2_22928 ( P3_ADD_553_U90 , P3_ADD_553_U179 , P3_ADD_553_U178 );
nand NAND2_22929 ( P3_ADD_553_U91 , P3_ADD_553_U181 , P3_ADD_553_U180 );
nand NAND2_22930 ( P3_ADD_553_U92 , P3_ADD_553_U183 , P3_ADD_553_U182 );
nand NAND2_22931 ( P3_ADD_553_U93 , P3_ADD_553_U185 , P3_ADD_553_U184 );
nand NAND2_22932 ( P3_ADD_553_U94 , P3_ADD_553_U187 , P3_ADD_553_U186 );
nand NAND2_22933 ( P3_ADD_553_U95 , P3_ADD_553_U189 , P3_ADD_553_U188 );
not NOT1_22934 ( P3_ADD_553_U96 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_22935 ( P3_ADD_553_U97 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_553_U126 );
not NOT1_22936 ( P3_ADD_553_U98 , P3_ADD_553_U7 );
not NOT1_22937 ( P3_ADD_553_U99 , P3_ADD_553_U9 );
not NOT1_22938 ( P3_ADD_553_U100 , P3_ADD_553_U11 );
not NOT1_22939 ( P3_ADD_553_U101 , P3_ADD_553_U13 );
not NOT1_22940 ( P3_ADD_553_U102 , P3_ADD_553_U15 );
not NOT1_22941 ( P3_ADD_553_U103 , P3_ADD_553_U17 );
not NOT1_22942 ( P3_ADD_553_U104 , P3_ADD_553_U19 );
not NOT1_22943 ( P3_ADD_553_U105 , P3_ADD_553_U22 );
not NOT1_22944 ( P3_ADD_553_U106 , P3_ADD_553_U23 );
not NOT1_22945 ( P3_ADD_553_U107 , P3_ADD_553_U25 );
not NOT1_22946 ( P3_ADD_553_U108 , P3_ADD_553_U27 );
not NOT1_22947 ( P3_ADD_553_U109 , P3_ADD_553_U29 );
not NOT1_22948 ( P3_ADD_553_U110 , P3_ADD_553_U31 );
not NOT1_22949 ( P3_ADD_553_U111 , P3_ADD_553_U33 );
not NOT1_22950 ( P3_ADD_553_U112 , P3_ADD_553_U35 );
not NOT1_22951 ( P3_ADD_553_U113 , P3_ADD_553_U37 );
not NOT1_22952 ( P3_ADD_553_U114 , P3_ADD_553_U39 );
not NOT1_22953 ( P3_ADD_553_U115 , P3_ADD_553_U41 );
not NOT1_22954 ( P3_ADD_553_U116 , P3_ADD_553_U43 );
not NOT1_22955 ( P3_ADD_553_U117 , P3_ADD_553_U45 );
not NOT1_22956 ( P3_ADD_553_U118 , P3_ADD_553_U47 );
not NOT1_22957 ( P3_ADD_553_U119 , P3_ADD_553_U49 );
not NOT1_22958 ( P3_ADD_553_U120 , P3_ADD_553_U51 );
not NOT1_22959 ( P3_ADD_553_U121 , P3_ADD_553_U53 );
not NOT1_22960 ( P3_ADD_553_U122 , P3_ADD_553_U55 );
not NOT1_22961 ( P3_ADD_553_U123 , P3_ADD_553_U57 );
not NOT1_22962 ( P3_ADD_553_U124 , P3_ADD_553_U59 );
not NOT1_22963 ( P3_ADD_553_U125 , P3_ADD_553_U61 );
not NOT1_22964 ( P3_ADD_553_U126 , P3_ADD_553_U63 );
not NOT1_22965 ( P3_ADD_553_U127 , P3_ADD_553_U97 );
nand NAND2_22966 ( P3_ADD_553_U128 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_553_U22 );
nand NAND2_22967 ( P3_ADD_553_U129 , P3_ADD_553_U105 , P3_ADD_553_U21 );
nand NAND2_22968 ( P3_ADD_553_U130 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_553_U19 );
nand NAND2_22969 ( P3_ADD_553_U131 , P3_ADD_553_U104 , P3_ADD_553_U20 );
nand NAND2_22970 ( P3_ADD_553_U132 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_553_U17 );
nand NAND2_22971 ( P3_ADD_553_U133 , P3_ADD_553_U103 , P3_ADD_553_U18 );
nand NAND2_22972 ( P3_ADD_553_U134 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_553_U15 );
nand NAND2_22973 ( P3_ADD_553_U135 , P3_ADD_553_U102 , P3_ADD_553_U16 );
nand NAND2_22974 ( P3_ADD_553_U136 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_553_U13 );
nand NAND2_22975 ( P3_ADD_553_U137 , P3_ADD_553_U101 , P3_ADD_553_U14 );
nand NAND2_22976 ( P3_ADD_553_U138 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_553_U11 );
nand NAND2_22977 ( P3_ADD_553_U139 , P3_ADD_553_U100 , P3_ADD_553_U12 );
nand NAND2_22978 ( P3_ADD_553_U140 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_553_U9 );
nand NAND2_22979 ( P3_ADD_553_U141 , P3_ADD_553_U99 , P3_ADD_553_U10 );
nand NAND2_22980 ( P3_ADD_553_U142 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_553_U97 );
nand NAND2_22981 ( P3_ADD_553_U143 , P3_ADD_553_U127 , P3_ADD_553_U96 );
nand NAND2_22982 ( P3_ADD_553_U144 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_553_U63 );
nand NAND2_22983 ( P3_ADD_553_U145 , P3_ADD_553_U126 , P3_ADD_553_U64 );
nand NAND2_22984 ( P3_ADD_553_U146 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_553_U7 );
nand NAND2_22985 ( P3_ADD_553_U147 , P3_ADD_553_U98 , P3_ADD_553_U8 );
nand NAND2_22986 ( P3_ADD_553_U148 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_553_U61 );
nand NAND2_22987 ( P3_ADD_553_U149 , P3_ADD_553_U125 , P3_ADD_553_U62 );
nand NAND2_22988 ( P3_ADD_553_U150 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_553_U59 );
nand NAND2_22989 ( P3_ADD_553_U151 , P3_ADD_553_U124 , P3_ADD_553_U60 );
nand NAND2_22990 ( P3_ADD_553_U152 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_553_U57 );
nand NAND2_22991 ( P3_ADD_553_U153 , P3_ADD_553_U123 , P3_ADD_553_U58 );
nand NAND2_22992 ( P3_ADD_553_U154 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_553_U55 );
nand NAND2_22993 ( P3_ADD_553_U155 , P3_ADD_553_U122 , P3_ADD_553_U56 );
nand NAND2_22994 ( P3_ADD_553_U156 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_553_U53 );
nand NAND2_22995 ( P3_ADD_553_U157 , P3_ADD_553_U121 , P3_ADD_553_U54 );
nand NAND2_22996 ( P3_ADD_553_U158 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_553_U51 );
nand NAND2_22997 ( P3_ADD_553_U159 , P3_ADD_553_U120 , P3_ADD_553_U52 );
nand NAND2_22998 ( P3_ADD_553_U160 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_553_U49 );
nand NAND2_22999 ( P3_ADD_553_U161 , P3_ADD_553_U119 , P3_ADD_553_U50 );
nand NAND2_23000 ( P3_ADD_553_U162 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_553_U47 );
nand NAND2_23001 ( P3_ADD_553_U163 , P3_ADD_553_U118 , P3_ADD_553_U48 );
nand NAND2_23002 ( P3_ADD_553_U164 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_553_U45 );
nand NAND2_23003 ( P3_ADD_553_U165 , P3_ADD_553_U117 , P3_ADD_553_U46 );
nand NAND2_23004 ( P3_ADD_553_U166 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_553_U43 );
nand NAND2_23005 ( P3_ADD_553_U167 , P3_ADD_553_U116 , P3_ADD_553_U44 );
nand NAND2_23006 ( P3_ADD_553_U168 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_553_U5 );
nand NAND2_23007 ( P3_ADD_553_U169 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_553_U6 );
nand NAND2_23008 ( P3_ADD_553_U170 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_553_U41 );
nand NAND2_23009 ( P3_ADD_553_U171 , P3_ADD_553_U115 , P3_ADD_553_U42 );
nand NAND2_23010 ( P3_ADD_553_U172 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_553_U39 );
nand NAND2_23011 ( P3_ADD_553_U173 , P3_ADD_553_U114 , P3_ADD_553_U40 );
nand NAND2_23012 ( P3_ADD_553_U174 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_553_U37 );
nand NAND2_23013 ( P3_ADD_553_U175 , P3_ADD_553_U113 , P3_ADD_553_U38 );
nand NAND2_23014 ( P3_ADD_553_U176 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_553_U35 );
nand NAND2_23015 ( P3_ADD_553_U177 , P3_ADD_553_U112 , P3_ADD_553_U36 );
nand NAND2_23016 ( P3_ADD_553_U178 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_553_U33 );
nand NAND2_23017 ( P3_ADD_553_U179 , P3_ADD_553_U111 , P3_ADD_553_U34 );
nand NAND2_23018 ( P3_ADD_553_U180 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_553_U31 );
nand NAND2_23019 ( P3_ADD_553_U181 , P3_ADD_553_U110 , P3_ADD_553_U32 );
nand NAND2_23020 ( P3_ADD_553_U182 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_553_U29 );
nand NAND2_23021 ( P3_ADD_553_U183 , P3_ADD_553_U109 , P3_ADD_553_U30 );
nand NAND2_23022 ( P3_ADD_553_U184 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_553_U27 );
nand NAND2_23023 ( P3_ADD_553_U185 , P3_ADD_553_U108 , P3_ADD_553_U28 );
nand NAND2_23024 ( P3_ADD_553_U186 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_553_U25 );
nand NAND2_23025 ( P3_ADD_553_U187 , P3_ADD_553_U107 , P3_ADD_553_U26 );
nand NAND2_23026 ( P3_ADD_553_U188 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_553_U23 );
nand NAND2_23027 ( P3_ADD_553_U189 , P3_ADD_553_U106 , P3_ADD_553_U24 );
not NOT1_23028 ( P3_ADD_558_U5 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_23029 ( P3_ADD_558_U6 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_23030 ( P3_ADD_558_U7 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_23031 ( P3_ADD_558_U8 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_23032 ( P3_ADD_558_U9 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_558_U98 );
not NOT1_23033 ( P3_ADD_558_U10 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_23034 ( P3_ADD_558_U11 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_558_U99 );
not NOT1_23035 ( P3_ADD_558_U12 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_23036 ( P3_ADD_558_U13 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_558_U100 );
not NOT1_23037 ( P3_ADD_558_U14 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_23038 ( P3_ADD_558_U15 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_558_U101 );
not NOT1_23039 ( P3_ADD_558_U16 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_23040 ( P3_ADD_558_U17 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_558_U102 );
not NOT1_23041 ( P3_ADD_558_U18 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_23042 ( P3_ADD_558_U19 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_558_U103 );
not NOT1_23043 ( P3_ADD_558_U20 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_23044 ( P3_ADD_558_U21 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_23045 ( P3_ADD_558_U22 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_558_U104 );
nand NAND2_23046 ( P3_ADD_558_U23 , P3_ADD_558_U105 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_23047 ( P3_ADD_558_U24 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_23048 ( P3_ADD_558_U25 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_558_U106 );
not NOT1_23049 ( P3_ADD_558_U26 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_23050 ( P3_ADD_558_U27 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_558_U107 );
not NOT1_23051 ( P3_ADD_558_U28 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_23052 ( P3_ADD_558_U29 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_558_U108 );
not NOT1_23053 ( P3_ADD_558_U30 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_23054 ( P3_ADD_558_U31 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_558_U109 );
not NOT1_23055 ( P3_ADD_558_U32 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_23056 ( P3_ADD_558_U33 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_558_U110 );
not NOT1_23057 ( P3_ADD_558_U34 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_23058 ( P3_ADD_558_U35 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_558_U111 );
not NOT1_23059 ( P3_ADD_558_U36 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_23060 ( P3_ADD_558_U37 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_558_U112 );
not NOT1_23061 ( P3_ADD_558_U38 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_23062 ( P3_ADD_558_U39 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_558_U113 );
not NOT1_23063 ( P3_ADD_558_U40 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_23064 ( P3_ADD_558_U41 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_558_U114 );
not NOT1_23065 ( P3_ADD_558_U42 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_23066 ( P3_ADD_558_U43 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_558_U115 );
not NOT1_23067 ( P3_ADD_558_U44 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_23068 ( P3_ADD_558_U45 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_558_U116 );
not NOT1_23069 ( P3_ADD_558_U46 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_23070 ( P3_ADD_558_U47 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_558_U117 );
not NOT1_23071 ( P3_ADD_558_U48 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_23072 ( P3_ADD_558_U49 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_558_U118 );
not NOT1_23073 ( P3_ADD_558_U50 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_23074 ( P3_ADD_558_U51 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_558_U119 );
not NOT1_23075 ( P3_ADD_558_U52 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_23076 ( P3_ADD_558_U53 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_558_U120 );
not NOT1_23077 ( P3_ADD_558_U54 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_23078 ( P3_ADD_558_U55 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_558_U121 );
not NOT1_23079 ( P3_ADD_558_U56 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_23080 ( P3_ADD_558_U57 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_558_U122 );
not NOT1_23081 ( P3_ADD_558_U58 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_23082 ( P3_ADD_558_U59 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_558_U123 );
not NOT1_23083 ( P3_ADD_558_U60 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_23084 ( P3_ADD_558_U61 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_558_U124 );
not NOT1_23085 ( P3_ADD_558_U62 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_23086 ( P3_ADD_558_U63 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_558_U125 );
not NOT1_23087 ( P3_ADD_558_U64 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_23088 ( P3_ADD_558_U65 , P3_ADD_558_U129 , P3_ADD_558_U128 );
nand NAND2_23089 ( P3_ADD_558_U66 , P3_ADD_558_U131 , P3_ADD_558_U130 );
nand NAND2_23090 ( P3_ADD_558_U67 , P3_ADD_558_U133 , P3_ADD_558_U132 );
nand NAND2_23091 ( P3_ADD_558_U68 , P3_ADD_558_U135 , P3_ADD_558_U134 );
nand NAND2_23092 ( P3_ADD_558_U69 , P3_ADD_558_U137 , P3_ADD_558_U136 );
nand NAND2_23093 ( P3_ADD_558_U70 , P3_ADD_558_U139 , P3_ADD_558_U138 );
nand NAND2_23094 ( P3_ADD_558_U71 , P3_ADD_558_U141 , P3_ADD_558_U140 );
nand NAND2_23095 ( P3_ADD_558_U72 , P3_ADD_558_U143 , P3_ADD_558_U142 );
nand NAND2_23096 ( P3_ADD_558_U73 , P3_ADD_558_U145 , P3_ADD_558_U144 );
nand NAND2_23097 ( P3_ADD_558_U74 , P3_ADD_558_U147 , P3_ADD_558_U146 );
nand NAND2_23098 ( P3_ADD_558_U75 , P3_ADD_558_U149 , P3_ADD_558_U148 );
nand NAND2_23099 ( P3_ADD_558_U76 , P3_ADD_558_U151 , P3_ADD_558_U150 );
nand NAND2_23100 ( P3_ADD_558_U77 , P3_ADD_558_U153 , P3_ADD_558_U152 );
nand NAND2_23101 ( P3_ADD_558_U78 , P3_ADD_558_U155 , P3_ADD_558_U154 );
nand NAND2_23102 ( P3_ADD_558_U79 , P3_ADD_558_U157 , P3_ADD_558_U156 );
nand NAND2_23103 ( P3_ADD_558_U80 , P3_ADD_558_U159 , P3_ADD_558_U158 );
nand NAND2_23104 ( P3_ADD_558_U81 , P3_ADD_558_U161 , P3_ADD_558_U160 );
nand NAND2_23105 ( P3_ADD_558_U82 , P3_ADD_558_U163 , P3_ADD_558_U162 );
nand NAND2_23106 ( P3_ADD_558_U83 , P3_ADD_558_U165 , P3_ADD_558_U164 );
nand NAND2_23107 ( P3_ADD_558_U84 , P3_ADD_558_U167 , P3_ADD_558_U166 );
nand NAND2_23108 ( P3_ADD_558_U85 , P3_ADD_558_U169 , P3_ADD_558_U168 );
nand NAND2_23109 ( P3_ADD_558_U86 , P3_ADD_558_U171 , P3_ADD_558_U170 );
nand NAND2_23110 ( P3_ADD_558_U87 , P3_ADD_558_U173 , P3_ADD_558_U172 );
nand NAND2_23111 ( P3_ADD_558_U88 , P3_ADD_558_U175 , P3_ADD_558_U174 );
nand NAND2_23112 ( P3_ADD_558_U89 , P3_ADD_558_U177 , P3_ADD_558_U176 );
nand NAND2_23113 ( P3_ADD_558_U90 , P3_ADD_558_U179 , P3_ADD_558_U178 );
nand NAND2_23114 ( P3_ADD_558_U91 , P3_ADD_558_U181 , P3_ADD_558_U180 );
nand NAND2_23115 ( P3_ADD_558_U92 , P3_ADD_558_U183 , P3_ADD_558_U182 );
nand NAND2_23116 ( P3_ADD_558_U93 , P3_ADD_558_U185 , P3_ADD_558_U184 );
nand NAND2_23117 ( P3_ADD_558_U94 , P3_ADD_558_U187 , P3_ADD_558_U186 );
nand NAND2_23118 ( P3_ADD_558_U95 , P3_ADD_558_U189 , P3_ADD_558_U188 );
not NOT1_23119 ( P3_ADD_558_U96 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_23120 ( P3_ADD_558_U97 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_558_U126 );
not NOT1_23121 ( P3_ADD_558_U98 , P3_ADD_558_U7 );
not NOT1_23122 ( P3_ADD_558_U99 , P3_ADD_558_U9 );
not NOT1_23123 ( P3_ADD_558_U100 , P3_ADD_558_U11 );
not NOT1_23124 ( P3_ADD_558_U101 , P3_ADD_558_U13 );
not NOT1_23125 ( P3_ADD_558_U102 , P3_ADD_558_U15 );
not NOT1_23126 ( P3_ADD_558_U103 , P3_ADD_558_U17 );
not NOT1_23127 ( P3_ADD_558_U104 , P3_ADD_558_U19 );
not NOT1_23128 ( P3_ADD_558_U105 , P3_ADD_558_U22 );
not NOT1_23129 ( P3_ADD_558_U106 , P3_ADD_558_U23 );
not NOT1_23130 ( P3_ADD_558_U107 , P3_ADD_558_U25 );
not NOT1_23131 ( P3_ADD_558_U108 , P3_ADD_558_U27 );
not NOT1_23132 ( P3_ADD_558_U109 , P3_ADD_558_U29 );
not NOT1_23133 ( P3_ADD_558_U110 , P3_ADD_558_U31 );
not NOT1_23134 ( P3_ADD_558_U111 , P3_ADD_558_U33 );
not NOT1_23135 ( P3_ADD_558_U112 , P3_ADD_558_U35 );
not NOT1_23136 ( P3_ADD_558_U113 , P3_ADD_558_U37 );
not NOT1_23137 ( P3_ADD_558_U114 , P3_ADD_558_U39 );
not NOT1_23138 ( P3_ADD_558_U115 , P3_ADD_558_U41 );
not NOT1_23139 ( P3_ADD_558_U116 , P3_ADD_558_U43 );
not NOT1_23140 ( P3_ADD_558_U117 , P3_ADD_558_U45 );
not NOT1_23141 ( P3_ADD_558_U118 , P3_ADD_558_U47 );
not NOT1_23142 ( P3_ADD_558_U119 , P3_ADD_558_U49 );
not NOT1_23143 ( P3_ADD_558_U120 , P3_ADD_558_U51 );
not NOT1_23144 ( P3_ADD_558_U121 , P3_ADD_558_U53 );
not NOT1_23145 ( P3_ADD_558_U122 , P3_ADD_558_U55 );
not NOT1_23146 ( P3_ADD_558_U123 , P3_ADD_558_U57 );
not NOT1_23147 ( P3_ADD_558_U124 , P3_ADD_558_U59 );
not NOT1_23148 ( P3_ADD_558_U125 , P3_ADD_558_U61 );
not NOT1_23149 ( P3_ADD_558_U126 , P3_ADD_558_U63 );
not NOT1_23150 ( P3_ADD_558_U127 , P3_ADD_558_U97 );
nand NAND2_23151 ( P3_ADD_558_U128 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_558_U22 );
nand NAND2_23152 ( P3_ADD_558_U129 , P3_ADD_558_U105 , P3_ADD_558_U21 );
nand NAND2_23153 ( P3_ADD_558_U130 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_558_U19 );
nand NAND2_23154 ( P3_ADD_558_U131 , P3_ADD_558_U104 , P3_ADD_558_U20 );
nand NAND2_23155 ( P3_ADD_558_U132 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_558_U17 );
nand NAND2_23156 ( P3_ADD_558_U133 , P3_ADD_558_U103 , P3_ADD_558_U18 );
nand NAND2_23157 ( P3_ADD_558_U134 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_558_U15 );
nand NAND2_23158 ( P3_ADD_558_U135 , P3_ADD_558_U102 , P3_ADD_558_U16 );
nand NAND2_23159 ( P3_ADD_558_U136 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_558_U13 );
nand NAND2_23160 ( P3_ADD_558_U137 , P3_ADD_558_U101 , P3_ADD_558_U14 );
nand NAND2_23161 ( P3_ADD_558_U138 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_558_U11 );
nand NAND2_23162 ( P3_ADD_558_U139 , P3_ADD_558_U100 , P3_ADD_558_U12 );
nand NAND2_23163 ( P3_ADD_558_U140 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_558_U9 );
nand NAND2_23164 ( P3_ADD_558_U141 , P3_ADD_558_U99 , P3_ADD_558_U10 );
nand NAND2_23165 ( P3_ADD_558_U142 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_558_U97 );
nand NAND2_23166 ( P3_ADD_558_U143 , P3_ADD_558_U127 , P3_ADD_558_U96 );
nand NAND2_23167 ( P3_ADD_558_U144 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_558_U63 );
nand NAND2_23168 ( P3_ADD_558_U145 , P3_ADD_558_U126 , P3_ADD_558_U64 );
nand NAND2_23169 ( P3_ADD_558_U146 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_558_U7 );
nand NAND2_23170 ( P3_ADD_558_U147 , P3_ADD_558_U98 , P3_ADD_558_U8 );
nand NAND2_23171 ( P3_ADD_558_U148 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_558_U61 );
nand NAND2_23172 ( P3_ADD_558_U149 , P3_ADD_558_U125 , P3_ADD_558_U62 );
nand NAND2_23173 ( P3_ADD_558_U150 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_558_U59 );
nand NAND2_23174 ( P3_ADD_558_U151 , P3_ADD_558_U124 , P3_ADD_558_U60 );
nand NAND2_23175 ( P3_ADD_558_U152 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_558_U57 );
nand NAND2_23176 ( P3_ADD_558_U153 , P3_ADD_558_U123 , P3_ADD_558_U58 );
nand NAND2_23177 ( P3_ADD_558_U154 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_558_U55 );
nand NAND2_23178 ( P3_ADD_558_U155 , P3_ADD_558_U122 , P3_ADD_558_U56 );
nand NAND2_23179 ( P3_ADD_558_U156 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_558_U53 );
nand NAND2_23180 ( P3_ADD_558_U157 , P3_ADD_558_U121 , P3_ADD_558_U54 );
nand NAND2_23181 ( P3_ADD_558_U158 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_558_U51 );
nand NAND2_23182 ( P3_ADD_558_U159 , P3_ADD_558_U120 , P3_ADD_558_U52 );
nand NAND2_23183 ( P3_ADD_558_U160 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_558_U49 );
nand NAND2_23184 ( P3_ADD_558_U161 , P3_ADD_558_U119 , P3_ADD_558_U50 );
nand NAND2_23185 ( P3_ADD_558_U162 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_558_U47 );
nand NAND2_23186 ( P3_ADD_558_U163 , P3_ADD_558_U118 , P3_ADD_558_U48 );
nand NAND2_23187 ( P3_ADD_558_U164 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_558_U45 );
nand NAND2_23188 ( P3_ADD_558_U165 , P3_ADD_558_U117 , P3_ADD_558_U46 );
nand NAND2_23189 ( P3_ADD_558_U166 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_558_U43 );
nand NAND2_23190 ( P3_ADD_558_U167 , P3_ADD_558_U116 , P3_ADD_558_U44 );
nand NAND2_23191 ( P3_ADD_558_U168 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_558_U5 );
nand NAND2_23192 ( P3_ADD_558_U169 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_558_U6 );
nand NAND2_23193 ( P3_ADD_558_U170 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_558_U41 );
nand NAND2_23194 ( P3_ADD_558_U171 , P3_ADD_558_U115 , P3_ADD_558_U42 );
nand NAND2_23195 ( P3_ADD_558_U172 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_558_U39 );
nand NAND2_23196 ( P3_ADD_558_U173 , P3_ADD_558_U114 , P3_ADD_558_U40 );
nand NAND2_23197 ( P3_ADD_558_U174 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_558_U37 );
nand NAND2_23198 ( P3_ADD_558_U175 , P3_ADD_558_U113 , P3_ADD_558_U38 );
nand NAND2_23199 ( P3_ADD_558_U176 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_558_U35 );
nand NAND2_23200 ( P3_ADD_558_U177 , P3_ADD_558_U112 , P3_ADD_558_U36 );
nand NAND2_23201 ( P3_ADD_558_U178 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_558_U33 );
nand NAND2_23202 ( P3_ADD_558_U179 , P3_ADD_558_U111 , P3_ADD_558_U34 );
nand NAND2_23203 ( P3_ADD_558_U180 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_558_U31 );
nand NAND2_23204 ( P3_ADD_558_U181 , P3_ADD_558_U110 , P3_ADD_558_U32 );
nand NAND2_23205 ( P3_ADD_558_U182 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_558_U29 );
nand NAND2_23206 ( P3_ADD_558_U183 , P3_ADD_558_U109 , P3_ADD_558_U30 );
nand NAND2_23207 ( P3_ADD_558_U184 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_558_U27 );
nand NAND2_23208 ( P3_ADD_558_U185 , P3_ADD_558_U108 , P3_ADD_558_U28 );
nand NAND2_23209 ( P3_ADD_558_U186 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_558_U25 );
nand NAND2_23210 ( P3_ADD_558_U187 , P3_ADD_558_U107 , P3_ADD_558_U26 );
nand NAND2_23211 ( P3_ADD_558_U188 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_558_U23 );
nand NAND2_23212 ( P3_ADD_558_U189 , P3_ADD_558_U106 , P3_ADD_558_U24 );
not NOT1_23213 ( P3_ADD_385_U5 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_23214 ( P3_ADD_385_U6 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_23215 ( P3_ADD_385_U7 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_23216 ( P3_ADD_385_U8 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_23217 ( P3_ADD_385_U9 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_385_U98 );
not NOT1_23218 ( P3_ADD_385_U10 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_23219 ( P3_ADD_385_U11 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_385_U99 );
not NOT1_23220 ( P3_ADD_385_U12 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_23221 ( P3_ADD_385_U13 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_385_U100 );
not NOT1_23222 ( P3_ADD_385_U14 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_23223 ( P3_ADD_385_U15 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_385_U101 );
not NOT1_23224 ( P3_ADD_385_U16 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_23225 ( P3_ADD_385_U17 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_385_U102 );
not NOT1_23226 ( P3_ADD_385_U18 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_23227 ( P3_ADD_385_U19 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_385_U103 );
not NOT1_23228 ( P3_ADD_385_U20 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_23229 ( P3_ADD_385_U21 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_23230 ( P3_ADD_385_U22 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_385_U104 );
nand NAND2_23231 ( P3_ADD_385_U23 , P3_ADD_385_U105 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_23232 ( P3_ADD_385_U24 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_23233 ( P3_ADD_385_U25 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_385_U106 );
not NOT1_23234 ( P3_ADD_385_U26 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_23235 ( P3_ADD_385_U27 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_385_U107 );
not NOT1_23236 ( P3_ADD_385_U28 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_23237 ( P3_ADD_385_U29 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_385_U108 );
not NOT1_23238 ( P3_ADD_385_U30 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_23239 ( P3_ADD_385_U31 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_385_U109 );
not NOT1_23240 ( P3_ADD_385_U32 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_23241 ( P3_ADD_385_U33 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_385_U110 );
not NOT1_23242 ( P3_ADD_385_U34 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_23243 ( P3_ADD_385_U35 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_385_U111 );
not NOT1_23244 ( P3_ADD_385_U36 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_23245 ( P3_ADD_385_U37 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_385_U112 );
not NOT1_23246 ( P3_ADD_385_U38 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_23247 ( P3_ADD_385_U39 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_385_U113 );
not NOT1_23248 ( P3_ADD_385_U40 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_23249 ( P3_ADD_385_U41 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_385_U114 );
not NOT1_23250 ( P3_ADD_385_U42 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_23251 ( P3_ADD_385_U43 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_385_U115 );
not NOT1_23252 ( P3_ADD_385_U44 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_23253 ( P3_ADD_385_U45 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_385_U116 );
not NOT1_23254 ( P3_ADD_385_U46 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_23255 ( P3_ADD_385_U47 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_385_U117 );
not NOT1_23256 ( P3_ADD_385_U48 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_23257 ( P3_ADD_385_U49 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_385_U118 );
not NOT1_23258 ( P3_ADD_385_U50 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_23259 ( P3_ADD_385_U51 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_385_U119 );
not NOT1_23260 ( P3_ADD_385_U52 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_23261 ( P3_ADD_385_U53 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_385_U120 );
not NOT1_23262 ( P3_ADD_385_U54 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_23263 ( P3_ADD_385_U55 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_385_U121 );
not NOT1_23264 ( P3_ADD_385_U56 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_23265 ( P3_ADD_385_U57 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_385_U122 );
not NOT1_23266 ( P3_ADD_385_U58 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_23267 ( P3_ADD_385_U59 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_385_U123 );
not NOT1_23268 ( P3_ADD_385_U60 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_23269 ( P3_ADD_385_U61 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_385_U124 );
not NOT1_23270 ( P3_ADD_385_U62 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_23271 ( P3_ADD_385_U63 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_385_U125 );
not NOT1_23272 ( P3_ADD_385_U64 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_23273 ( P3_ADD_385_U65 , P3_ADD_385_U129 , P3_ADD_385_U128 );
nand NAND2_23274 ( P3_ADD_385_U66 , P3_ADD_385_U131 , P3_ADD_385_U130 );
nand NAND2_23275 ( P3_ADD_385_U67 , P3_ADD_385_U133 , P3_ADD_385_U132 );
nand NAND2_23276 ( P3_ADD_385_U68 , P3_ADD_385_U135 , P3_ADD_385_U134 );
nand NAND2_23277 ( P3_ADD_385_U69 , P3_ADD_385_U137 , P3_ADD_385_U136 );
nand NAND2_23278 ( P3_ADD_385_U70 , P3_ADD_385_U139 , P3_ADD_385_U138 );
nand NAND2_23279 ( P3_ADD_385_U71 , P3_ADD_385_U141 , P3_ADD_385_U140 );
nand NAND2_23280 ( P3_ADD_385_U72 , P3_ADD_385_U143 , P3_ADD_385_U142 );
nand NAND2_23281 ( P3_ADD_385_U73 , P3_ADD_385_U145 , P3_ADD_385_U144 );
nand NAND2_23282 ( P3_ADD_385_U74 , P3_ADD_385_U147 , P3_ADD_385_U146 );
nand NAND2_23283 ( P3_ADD_385_U75 , P3_ADD_385_U149 , P3_ADD_385_U148 );
nand NAND2_23284 ( P3_ADD_385_U76 , P3_ADD_385_U151 , P3_ADD_385_U150 );
nand NAND2_23285 ( P3_ADD_385_U77 , P3_ADD_385_U153 , P3_ADD_385_U152 );
nand NAND2_23286 ( P3_ADD_385_U78 , P3_ADD_385_U155 , P3_ADD_385_U154 );
nand NAND2_23287 ( P3_ADD_385_U79 , P3_ADD_385_U157 , P3_ADD_385_U156 );
nand NAND2_23288 ( P3_ADD_385_U80 , P3_ADD_385_U159 , P3_ADD_385_U158 );
nand NAND2_23289 ( P3_ADD_385_U81 , P3_ADD_385_U161 , P3_ADD_385_U160 );
nand NAND2_23290 ( P3_ADD_385_U82 , P3_ADD_385_U163 , P3_ADD_385_U162 );
nand NAND2_23291 ( P3_ADD_385_U83 , P3_ADD_385_U165 , P3_ADD_385_U164 );
nand NAND2_23292 ( P3_ADD_385_U84 , P3_ADD_385_U167 , P3_ADD_385_U166 );
nand NAND2_23293 ( P3_ADD_385_U85 , P3_ADD_385_U169 , P3_ADD_385_U168 );
nand NAND2_23294 ( P3_ADD_385_U86 , P3_ADD_385_U171 , P3_ADD_385_U170 );
nand NAND2_23295 ( P3_ADD_385_U87 , P3_ADD_385_U173 , P3_ADD_385_U172 );
nand NAND2_23296 ( P3_ADD_385_U88 , P3_ADD_385_U175 , P3_ADD_385_U174 );
nand NAND2_23297 ( P3_ADD_385_U89 , P3_ADD_385_U177 , P3_ADD_385_U176 );
nand NAND2_23298 ( P3_ADD_385_U90 , P3_ADD_385_U179 , P3_ADD_385_U178 );
nand NAND2_23299 ( P3_ADD_385_U91 , P3_ADD_385_U181 , P3_ADD_385_U180 );
nand NAND2_23300 ( P3_ADD_385_U92 , P3_ADD_385_U183 , P3_ADD_385_U182 );
nand NAND2_23301 ( P3_ADD_385_U93 , P3_ADD_385_U185 , P3_ADD_385_U184 );
nand NAND2_23302 ( P3_ADD_385_U94 , P3_ADD_385_U187 , P3_ADD_385_U186 );
nand NAND2_23303 ( P3_ADD_385_U95 , P3_ADD_385_U189 , P3_ADD_385_U188 );
not NOT1_23304 ( P3_ADD_385_U96 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_23305 ( P3_ADD_385_U97 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_385_U126 );
not NOT1_23306 ( P3_ADD_385_U98 , P3_ADD_385_U7 );
not NOT1_23307 ( P3_ADD_385_U99 , P3_ADD_385_U9 );
not NOT1_23308 ( P3_ADD_385_U100 , P3_ADD_385_U11 );
not NOT1_23309 ( P3_ADD_385_U101 , P3_ADD_385_U13 );
not NOT1_23310 ( P3_ADD_385_U102 , P3_ADD_385_U15 );
not NOT1_23311 ( P3_ADD_385_U103 , P3_ADD_385_U17 );
not NOT1_23312 ( P3_ADD_385_U104 , P3_ADD_385_U19 );
not NOT1_23313 ( P3_ADD_385_U105 , P3_ADD_385_U22 );
not NOT1_23314 ( P3_ADD_385_U106 , P3_ADD_385_U23 );
not NOT1_23315 ( P3_ADD_385_U107 , P3_ADD_385_U25 );
not NOT1_23316 ( P3_ADD_385_U108 , P3_ADD_385_U27 );
not NOT1_23317 ( P3_ADD_385_U109 , P3_ADD_385_U29 );
not NOT1_23318 ( P3_ADD_385_U110 , P3_ADD_385_U31 );
not NOT1_23319 ( P3_ADD_385_U111 , P3_ADD_385_U33 );
not NOT1_23320 ( P3_ADD_385_U112 , P3_ADD_385_U35 );
not NOT1_23321 ( P3_ADD_385_U113 , P3_ADD_385_U37 );
not NOT1_23322 ( P3_ADD_385_U114 , P3_ADD_385_U39 );
not NOT1_23323 ( P3_ADD_385_U115 , P3_ADD_385_U41 );
not NOT1_23324 ( P3_ADD_385_U116 , P3_ADD_385_U43 );
not NOT1_23325 ( P3_ADD_385_U117 , P3_ADD_385_U45 );
not NOT1_23326 ( P3_ADD_385_U118 , P3_ADD_385_U47 );
not NOT1_23327 ( P3_ADD_385_U119 , P3_ADD_385_U49 );
not NOT1_23328 ( P3_ADD_385_U120 , P3_ADD_385_U51 );
not NOT1_23329 ( P3_ADD_385_U121 , P3_ADD_385_U53 );
not NOT1_23330 ( P3_ADD_385_U122 , P3_ADD_385_U55 );
not NOT1_23331 ( P3_ADD_385_U123 , P3_ADD_385_U57 );
not NOT1_23332 ( P3_ADD_385_U124 , P3_ADD_385_U59 );
not NOT1_23333 ( P3_ADD_385_U125 , P3_ADD_385_U61 );
not NOT1_23334 ( P3_ADD_385_U126 , P3_ADD_385_U63 );
not NOT1_23335 ( P3_ADD_385_U127 , P3_ADD_385_U97 );
nand NAND2_23336 ( P3_ADD_385_U128 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_385_U22 );
nand NAND2_23337 ( P3_ADD_385_U129 , P3_ADD_385_U105 , P3_ADD_385_U21 );
nand NAND2_23338 ( P3_ADD_385_U130 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_385_U19 );
nand NAND2_23339 ( P3_ADD_385_U131 , P3_ADD_385_U104 , P3_ADD_385_U20 );
nand NAND2_23340 ( P3_ADD_385_U132 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_385_U17 );
nand NAND2_23341 ( P3_ADD_385_U133 , P3_ADD_385_U103 , P3_ADD_385_U18 );
nand NAND2_23342 ( P3_ADD_385_U134 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_385_U15 );
nand NAND2_23343 ( P3_ADD_385_U135 , P3_ADD_385_U102 , P3_ADD_385_U16 );
nand NAND2_23344 ( P3_ADD_385_U136 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_385_U13 );
nand NAND2_23345 ( P3_ADD_385_U137 , P3_ADD_385_U101 , P3_ADD_385_U14 );
nand NAND2_23346 ( P3_ADD_385_U138 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_385_U11 );
nand NAND2_23347 ( P3_ADD_385_U139 , P3_ADD_385_U100 , P3_ADD_385_U12 );
nand NAND2_23348 ( P3_ADD_385_U140 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_385_U9 );
nand NAND2_23349 ( P3_ADD_385_U141 , P3_ADD_385_U99 , P3_ADD_385_U10 );
nand NAND2_23350 ( P3_ADD_385_U142 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_385_U97 );
nand NAND2_23351 ( P3_ADD_385_U143 , P3_ADD_385_U127 , P3_ADD_385_U96 );
nand NAND2_23352 ( P3_ADD_385_U144 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_385_U63 );
nand NAND2_23353 ( P3_ADD_385_U145 , P3_ADD_385_U126 , P3_ADD_385_U64 );
nand NAND2_23354 ( P3_ADD_385_U146 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_385_U7 );
nand NAND2_23355 ( P3_ADD_385_U147 , P3_ADD_385_U98 , P3_ADD_385_U8 );
nand NAND2_23356 ( P3_ADD_385_U148 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_385_U61 );
nand NAND2_23357 ( P3_ADD_385_U149 , P3_ADD_385_U125 , P3_ADD_385_U62 );
nand NAND2_23358 ( P3_ADD_385_U150 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_385_U59 );
nand NAND2_23359 ( P3_ADD_385_U151 , P3_ADD_385_U124 , P3_ADD_385_U60 );
nand NAND2_23360 ( P3_ADD_385_U152 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_385_U57 );
nand NAND2_23361 ( P3_ADD_385_U153 , P3_ADD_385_U123 , P3_ADD_385_U58 );
nand NAND2_23362 ( P3_ADD_385_U154 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_385_U55 );
nand NAND2_23363 ( P3_ADD_385_U155 , P3_ADD_385_U122 , P3_ADD_385_U56 );
nand NAND2_23364 ( P3_ADD_385_U156 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_385_U53 );
nand NAND2_23365 ( P3_ADD_385_U157 , P3_ADD_385_U121 , P3_ADD_385_U54 );
nand NAND2_23366 ( P3_ADD_385_U158 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_385_U51 );
nand NAND2_23367 ( P3_ADD_385_U159 , P3_ADD_385_U120 , P3_ADD_385_U52 );
nand NAND2_23368 ( P3_ADD_385_U160 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_385_U49 );
nand NAND2_23369 ( P3_ADD_385_U161 , P3_ADD_385_U119 , P3_ADD_385_U50 );
nand NAND2_23370 ( P3_ADD_385_U162 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_385_U47 );
nand NAND2_23371 ( P3_ADD_385_U163 , P3_ADD_385_U118 , P3_ADD_385_U48 );
nand NAND2_23372 ( P3_ADD_385_U164 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_385_U45 );
nand NAND2_23373 ( P3_ADD_385_U165 , P3_ADD_385_U117 , P3_ADD_385_U46 );
nand NAND2_23374 ( P3_ADD_385_U166 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_385_U43 );
nand NAND2_23375 ( P3_ADD_385_U167 , P3_ADD_385_U116 , P3_ADD_385_U44 );
nand NAND2_23376 ( P3_ADD_385_U168 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_385_U5 );
nand NAND2_23377 ( P3_ADD_385_U169 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_385_U6 );
nand NAND2_23378 ( P3_ADD_385_U170 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_385_U41 );
nand NAND2_23379 ( P3_ADD_385_U171 , P3_ADD_385_U115 , P3_ADD_385_U42 );
nand NAND2_23380 ( P3_ADD_385_U172 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_385_U39 );
nand NAND2_23381 ( P3_ADD_385_U173 , P3_ADD_385_U114 , P3_ADD_385_U40 );
nand NAND2_23382 ( P3_ADD_385_U174 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_385_U37 );
nand NAND2_23383 ( P3_ADD_385_U175 , P3_ADD_385_U113 , P3_ADD_385_U38 );
nand NAND2_23384 ( P3_ADD_385_U176 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_385_U35 );
nand NAND2_23385 ( P3_ADD_385_U177 , P3_ADD_385_U112 , P3_ADD_385_U36 );
nand NAND2_23386 ( P3_ADD_385_U178 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_385_U33 );
nand NAND2_23387 ( P3_ADD_385_U179 , P3_ADD_385_U111 , P3_ADD_385_U34 );
nand NAND2_23388 ( P3_ADD_385_U180 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_385_U31 );
nand NAND2_23389 ( P3_ADD_385_U181 , P3_ADD_385_U110 , P3_ADD_385_U32 );
nand NAND2_23390 ( P3_ADD_385_U182 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_385_U29 );
nand NAND2_23391 ( P3_ADD_385_U183 , P3_ADD_385_U109 , P3_ADD_385_U30 );
nand NAND2_23392 ( P3_ADD_385_U184 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_385_U27 );
nand NAND2_23393 ( P3_ADD_385_U185 , P3_ADD_385_U108 , P3_ADD_385_U28 );
nand NAND2_23394 ( P3_ADD_385_U186 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_385_U25 );
nand NAND2_23395 ( P3_ADD_385_U187 , P3_ADD_385_U107 , P3_ADD_385_U26 );
nand NAND2_23396 ( P3_ADD_385_U188 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_385_U23 );
nand NAND2_23397 ( P3_ADD_385_U189 , P3_ADD_385_U106 , P3_ADD_385_U24 );
nand NAND2_23398 ( P3_ADD_357_U6 , P3_ADD_357_U15 , P3_ADD_357_U23 );
and AND2_23399 ( P3_ADD_357_U7 , P3_ADD_357_U29 , P3_ADD_357_U11 );
and AND2_23400 ( P3_ADD_357_U8 , P3_ADD_357_U27 , P3_ADD_357_U12 );
and AND2_23401 ( P3_ADD_357_U9 , P3_ADD_357_U25 , P3_ADD_357_U6 );
not NOT1_23402 ( P3_ADD_357_U10 , P3_SUB_357_U10 );
or OR3_23403 ( P3_ADD_357_U11 , P3_SUB_357_U7 , P3_SUB_357_U12 , P3_SUB_357_U11 );
nand NAND2_23404 ( P3_ADD_357_U12 , P3_ADD_357_U14 , P3_ADD_357_U22 );
nand NAND2_23405 ( P3_ADD_357_U13 , P3_ADD_357_U35 , P3_ADD_357_U34 );
nor nor_23406 ( P3_ADD_357_U14 , P3_SUB_357_U13 , P3_SUB_357_U9 );
nor nor_23407 ( P3_ADD_357_U15 , P3_SUB_357_U6 , P3_SUB_357_U8 );
not NOT1_23408 ( P3_ADD_357_U16 , P3_SUB_357_U6 );
and AND2_23409 ( P3_ADD_357_U17 , P3_ADD_357_U31 , P3_ADD_357_U30 );
not NOT1_23410 ( P3_ADD_357_U18 , P3_SUB_357_U13 );
and AND2_23411 ( P3_ADD_357_U19 , P3_ADD_357_U33 , P3_ADD_357_U32 );
not NOT1_23412 ( P3_ADD_357_U20 , P3_SUB_357_U7 );
not NOT1_23413 ( P3_ADD_357_U21 , P3_SUB_357_U12 );
not NOT1_23414 ( P3_ADD_357_U22 , P3_ADD_357_U11 );
not NOT1_23415 ( P3_ADD_357_U23 , P3_ADD_357_U12 );
nand NAND2_23416 ( P3_ADD_357_U24 , P3_ADD_357_U23 , P3_ADD_357_U16 );
nand NAND2_23417 ( P3_ADD_357_U25 , P3_SUB_357_U8 , P3_ADD_357_U24 );
nand NAND2_23418 ( P3_ADD_357_U26 , P3_ADD_357_U22 , P3_ADD_357_U18 );
nand NAND2_23419 ( P3_ADD_357_U27 , P3_SUB_357_U9 , P3_ADD_357_U26 );
or OR2_23420 ( P3_ADD_357_U28 , P3_SUB_357_U7 , P3_SUB_357_U12 );
nand NAND2_23421 ( P3_ADD_357_U29 , P3_SUB_357_U11 , P3_ADD_357_U28 );
nand NAND2_23422 ( P3_ADD_357_U30 , P3_SUB_357_U6 , P3_ADD_357_U12 );
nand NAND2_23423 ( P3_ADD_357_U31 , P3_ADD_357_U23 , P3_ADD_357_U16 );
nand NAND2_23424 ( P3_ADD_357_U32 , P3_SUB_357_U13 , P3_ADD_357_U11 );
nand NAND2_23425 ( P3_ADD_357_U33 , P3_ADD_357_U22 , P3_ADD_357_U18 );
nand NAND2_23426 ( P3_ADD_357_U34 , P3_SUB_357_U7 , P3_ADD_357_U21 );
nand NAND2_23427 ( P3_ADD_357_U35 , P3_SUB_357_U12 , P3_ADD_357_U20 );
not NOT1_23428 ( P3_ADD_547_U5 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_23429 ( P3_ADD_547_U6 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_23430 ( P3_ADD_547_U7 , P3_INSTADDRPOINTER_REG_1_ , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_23431 ( P3_ADD_547_U8 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_23432 ( P3_ADD_547_U9 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_547_U98 );
not NOT1_23433 ( P3_ADD_547_U10 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_23434 ( P3_ADD_547_U11 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_547_U99 );
not NOT1_23435 ( P3_ADD_547_U12 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_23436 ( P3_ADD_547_U13 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_547_U100 );
not NOT1_23437 ( P3_ADD_547_U14 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_23438 ( P3_ADD_547_U15 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_547_U101 );
not NOT1_23439 ( P3_ADD_547_U16 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_23440 ( P3_ADD_547_U17 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_547_U102 );
not NOT1_23441 ( P3_ADD_547_U18 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_23442 ( P3_ADD_547_U19 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_547_U103 );
not NOT1_23443 ( P3_ADD_547_U20 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_23444 ( P3_ADD_547_U21 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_23445 ( P3_ADD_547_U22 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_547_U104 );
nand NAND2_23446 ( P3_ADD_547_U23 , P3_ADD_547_U105 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_23447 ( P3_ADD_547_U24 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_23448 ( P3_ADD_547_U25 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_547_U106 );
not NOT1_23449 ( P3_ADD_547_U26 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_23450 ( P3_ADD_547_U27 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_547_U107 );
not NOT1_23451 ( P3_ADD_547_U28 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_23452 ( P3_ADD_547_U29 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_547_U108 );
not NOT1_23453 ( P3_ADD_547_U30 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_23454 ( P3_ADD_547_U31 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_547_U109 );
not NOT1_23455 ( P3_ADD_547_U32 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_23456 ( P3_ADD_547_U33 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_547_U110 );
not NOT1_23457 ( P3_ADD_547_U34 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_23458 ( P3_ADD_547_U35 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_547_U111 );
not NOT1_23459 ( P3_ADD_547_U36 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_23460 ( P3_ADD_547_U37 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_547_U112 );
not NOT1_23461 ( P3_ADD_547_U38 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_23462 ( P3_ADD_547_U39 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_547_U113 );
not NOT1_23463 ( P3_ADD_547_U40 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_23464 ( P3_ADD_547_U41 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_547_U114 );
not NOT1_23465 ( P3_ADD_547_U42 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_23466 ( P3_ADD_547_U43 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_547_U115 );
not NOT1_23467 ( P3_ADD_547_U44 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_23468 ( P3_ADD_547_U45 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_547_U116 );
not NOT1_23469 ( P3_ADD_547_U46 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_23470 ( P3_ADD_547_U47 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_547_U117 );
not NOT1_23471 ( P3_ADD_547_U48 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_23472 ( P3_ADD_547_U49 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_547_U118 );
not NOT1_23473 ( P3_ADD_547_U50 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_23474 ( P3_ADD_547_U51 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_547_U119 );
not NOT1_23475 ( P3_ADD_547_U52 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_23476 ( P3_ADD_547_U53 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_547_U120 );
not NOT1_23477 ( P3_ADD_547_U54 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_23478 ( P3_ADD_547_U55 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_547_U121 );
not NOT1_23479 ( P3_ADD_547_U56 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_23480 ( P3_ADD_547_U57 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_547_U122 );
not NOT1_23481 ( P3_ADD_547_U58 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_23482 ( P3_ADD_547_U59 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_547_U123 );
not NOT1_23483 ( P3_ADD_547_U60 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_23484 ( P3_ADD_547_U61 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_547_U124 );
not NOT1_23485 ( P3_ADD_547_U62 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_23486 ( P3_ADD_547_U63 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_547_U125 );
not NOT1_23487 ( P3_ADD_547_U64 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_23488 ( P3_ADD_547_U65 , P3_ADD_547_U129 , P3_ADD_547_U128 );
nand NAND2_23489 ( P3_ADD_547_U66 , P3_ADD_547_U131 , P3_ADD_547_U130 );
nand NAND2_23490 ( P3_ADD_547_U67 , P3_ADD_547_U133 , P3_ADD_547_U132 );
nand NAND2_23491 ( P3_ADD_547_U68 , P3_ADD_547_U135 , P3_ADD_547_U134 );
nand NAND2_23492 ( P3_ADD_547_U69 , P3_ADD_547_U137 , P3_ADD_547_U136 );
nand NAND2_23493 ( P3_ADD_547_U70 , P3_ADD_547_U139 , P3_ADD_547_U138 );
nand NAND2_23494 ( P3_ADD_547_U71 , P3_ADD_547_U141 , P3_ADD_547_U140 );
nand NAND2_23495 ( P3_ADD_547_U72 , P3_ADD_547_U143 , P3_ADD_547_U142 );
nand NAND2_23496 ( P3_ADD_547_U73 , P3_ADD_547_U145 , P3_ADD_547_U144 );
nand NAND2_23497 ( P3_ADD_547_U74 , P3_ADD_547_U147 , P3_ADD_547_U146 );
nand NAND2_23498 ( P3_ADD_547_U75 , P3_ADD_547_U149 , P3_ADD_547_U148 );
nand NAND2_23499 ( P3_ADD_547_U76 , P3_ADD_547_U151 , P3_ADD_547_U150 );
nand NAND2_23500 ( P3_ADD_547_U77 , P3_ADD_547_U153 , P3_ADD_547_U152 );
nand NAND2_23501 ( P3_ADD_547_U78 , P3_ADD_547_U155 , P3_ADD_547_U154 );
nand NAND2_23502 ( P3_ADD_547_U79 , P3_ADD_547_U157 , P3_ADD_547_U156 );
nand NAND2_23503 ( P3_ADD_547_U80 , P3_ADD_547_U159 , P3_ADD_547_U158 );
nand NAND2_23504 ( P3_ADD_547_U81 , P3_ADD_547_U161 , P3_ADD_547_U160 );
nand NAND2_23505 ( P3_ADD_547_U82 , P3_ADD_547_U163 , P3_ADD_547_U162 );
nand NAND2_23506 ( P3_ADD_547_U83 , P3_ADD_547_U165 , P3_ADD_547_U164 );
nand NAND2_23507 ( P3_ADD_547_U84 , P3_ADD_547_U167 , P3_ADD_547_U166 );
nand NAND2_23508 ( P3_ADD_547_U85 , P3_ADD_547_U169 , P3_ADD_547_U168 );
nand NAND2_23509 ( P3_ADD_547_U86 , P3_ADD_547_U171 , P3_ADD_547_U170 );
nand NAND2_23510 ( P3_ADD_547_U87 , P3_ADD_547_U173 , P3_ADD_547_U172 );
nand NAND2_23511 ( P3_ADD_547_U88 , P3_ADD_547_U175 , P3_ADD_547_U174 );
nand NAND2_23512 ( P3_ADD_547_U89 , P3_ADD_547_U177 , P3_ADD_547_U176 );
nand NAND2_23513 ( P3_ADD_547_U90 , P3_ADD_547_U179 , P3_ADD_547_U178 );
nand NAND2_23514 ( P3_ADD_547_U91 , P3_ADD_547_U181 , P3_ADD_547_U180 );
nand NAND2_23515 ( P3_ADD_547_U92 , P3_ADD_547_U183 , P3_ADD_547_U182 );
nand NAND2_23516 ( P3_ADD_547_U93 , P3_ADD_547_U185 , P3_ADD_547_U184 );
nand NAND2_23517 ( P3_ADD_547_U94 , P3_ADD_547_U187 , P3_ADD_547_U186 );
nand NAND2_23518 ( P3_ADD_547_U95 , P3_ADD_547_U189 , P3_ADD_547_U188 );
not NOT1_23519 ( P3_ADD_547_U96 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_23520 ( P3_ADD_547_U97 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_547_U126 );
not NOT1_23521 ( P3_ADD_547_U98 , P3_ADD_547_U7 );
not NOT1_23522 ( P3_ADD_547_U99 , P3_ADD_547_U9 );
not NOT1_23523 ( P3_ADD_547_U100 , P3_ADD_547_U11 );
not NOT1_23524 ( P3_ADD_547_U101 , P3_ADD_547_U13 );
not NOT1_23525 ( P3_ADD_547_U102 , P3_ADD_547_U15 );
not NOT1_23526 ( P3_ADD_547_U103 , P3_ADD_547_U17 );
not NOT1_23527 ( P3_ADD_547_U104 , P3_ADD_547_U19 );
not NOT1_23528 ( P3_ADD_547_U105 , P3_ADD_547_U22 );
not NOT1_23529 ( P3_ADD_547_U106 , P3_ADD_547_U23 );
not NOT1_23530 ( P3_ADD_547_U107 , P3_ADD_547_U25 );
not NOT1_23531 ( P3_ADD_547_U108 , P3_ADD_547_U27 );
not NOT1_23532 ( P3_ADD_547_U109 , P3_ADD_547_U29 );
not NOT1_23533 ( P3_ADD_547_U110 , P3_ADD_547_U31 );
not NOT1_23534 ( P3_ADD_547_U111 , P3_ADD_547_U33 );
not NOT1_23535 ( P3_ADD_547_U112 , P3_ADD_547_U35 );
not NOT1_23536 ( P3_ADD_547_U113 , P3_ADD_547_U37 );
not NOT1_23537 ( P3_ADD_547_U114 , P3_ADD_547_U39 );
not NOT1_23538 ( P3_ADD_547_U115 , P3_ADD_547_U41 );
not NOT1_23539 ( P3_ADD_547_U116 , P3_ADD_547_U43 );
not NOT1_23540 ( P3_ADD_547_U117 , P3_ADD_547_U45 );
not NOT1_23541 ( P3_ADD_547_U118 , P3_ADD_547_U47 );
not NOT1_23542 ( P3_ADD_547_U119 , P3_ADD_547_U49 );
not NOT1_23543 ( P3_ADD_547_U120 , P3_ADD_547_U51 );
not NOT1_23544 ( P3_ADD_547_U121 , P3_ADD_547_U53 );
not NOT1_23545 ( P3_ADD_547_U122 , P3_ADD_547_U55 );
not NOT1_23546 ( P3_ADD_547_U123 , P3_ADD_547_U57 );
not NOT1_23547 ( P3_ADD_547_U124 , P3_ADD_547_U59 );
not NOT1_23548 ( P3_ADD_547_U125 , P3_ADD_547_U61 );
not NOT1_23549 ( P3_ADD_547_U126 , P3_ADD_547_U63 );
not NOT1_23550 ( P3_ADD_547_U127 , P3_ADD_547_U97 );
nand NAND2_23551 ( P3_ADD_547_U128 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_547_U22 );
nand NAND2_23552 ( P3_ADD_547_U129 , P3_ADD_547_U105 , P3_ADD_547_U21 );
nand NAND2_23553 ( P3_ADD_547_U130 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_547_U19 );
nand NAND2_23554 ( P3_ADD_547_U131 , P3_ADD_547_U104 , P3_ADD_547_U20 );
nand NAND2_23555 ( P3_ADD_547_U132 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_547_U17 );
nand NAND2_23556 ( P3_ADD_547_U133 , P3_ADD_547_U103 , P3_ADD_547_U18 );
nand NAND2_23557 ( P3_ADD_547_U134 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_547_U15 );
nand NAND2_23558 ( P3_ADD_547_U135 , P3_ADD_547_U102 , P3_ADD_547_U16 );
nand NAND2_23559 ( P3_ADD_547_U136 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_547_U13 );
nand NAND2_23560 ( P3_ADD_547_U137 , P3_ADD_547_U101 , P3_ADD_547_U14 );
nand NAND2_23561 ( P3_ADD_547_U138 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_547_U11 );
nand NAND2_23562 ( P3_ADD_547_U139 , P3_ADD_547_U100 , P3_ADD_547_U12 );
nand NAND2_23563 ( P3_ADD_547_U140 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_547_U9 );
nand NAND2_23564 ( P3_ADD_547_U141 , P3_ADD_547_U99 , P3_ADD_547_U10 );
nand NAND2_23565 ( P3_ADD_547_U142 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_547_U97 );
nand NAND2_23566 ( P3_ADD_547_U143 , P3_ADD_547_U127 , P3_ADD_547_U96 );
nand NAND2_23567 ( P3_ADD_547_U144 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_547_U63 );
nand NAND2_23568 ( P3_ADD_547_U145 , P3_ADD_547_U126 , P3_ADD_547_U64 );
nand NAND2_23569 ( P3_ADD_547_U146 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_547_U7 );
nand NAND2_23570 ( P3_ADD_547_U147 , P3_ADD_547_U98 , P3_ADD_547_U8 );
nand NAND2_23571 ( P3_ADD_547_U148 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_547_U61 );
nand NAND2_23572 ( P3_ADD_547_U149 , P3_ADD_547_U125 , P3_ADD_547_U62 );
nand NAND2_23573 ( P3_ADD_547_U150 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_547_U59 );
nand NAND2_23574 ( P3_ADD_547_U151 , P3_ADD_547_U124 , P3_ADD_547_U60 );
nand NAND2_23575 ( P3_ADD_547_U152 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_547_U57 );
nand NAND2_23576 ( P3_ADD_547_U153 , P3_ADD_547_U123 , P3_ADD_547_U58 );
nand NAND2_23577 ( P3_ADD_547_U154 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_547_U55 );
nand NAND2_23578 ( P3_ADD_547_U155 , P3_ADD_547_U122 , P3_ADD_547_U56 );
nand NAND2_23579 ( P3_ADD_547_U156 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_547_U53 );
nand NAND2_23580 ( P3_ADD_547_U157 , P3_ADD_547_U121 , P3_ADD_547_U54 );
nand NAND2_23581 ( P3_ADD_547_U158 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_547_U51 );
nand NAND2_23582 ( P3_ADD_547_U159 , P3_ADD_547_U120 , P3_ADD_547_U52 );
nand NAND2_23583 ( P3_ADD_547_U160 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_547_U49 );
nand NAND2_23584 ( P3_ADD_547_U161 , P3_ADD_547_U119 , P3_ADD_547_U50 );
nand NAND2_23585 ( P3_ADD_547_U162 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_547_U47 );
nand NAND2_23586 ( P3_ADD_547_U163 , P3_ADD_547_U118 , P3_ADD_547_U48 );
nand NAND2_23587 ( P3_ADD_547_U164 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_547_U45 );
nand NAND2_23588 ( P3_ADD_547_U165 , P3_ADD_547_U117 , P3_ADD_547_U46 );
nand NAND2_23589 ( P3_ADD_547_U166 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_547_U43 );
nand NAND2_23590 ( P3_ADD_547_U167 , P3_ADD_547_U116 , P3_ADD_547_U44 );
nand NAND2_23591 ( P3_ADD_547_U168 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_547_U5 );
nand NAND2_23592 ( P3_ADD_547_U169 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_547_U6 );
nand NAND2_23593 ( P3_ADD_547_U170 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_547_U41 );
nand NAND2_23594 ( P3_ADD_547_U171 , P3_ADD_547_U115 , P3_ADD_547_U42 );
nand NAND2_23595 ( P3_ADD_547_U172 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_547_U39 );
nand NAND2_23596 ( P3_ADD_547_U173 , P3_ADD_547_U114 , P3_ADD_547_U40 );
nand NAND2_23597 ( P3_ADD_547_U174 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_547_U37 );
nand NAND2_23598 ( P3_ADD_547_U175 , P3_ADD_547_U113 , P3_ADD_547_U38 );
nand NAND2_23599 ( P3_ADD_547_U176 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_547_U35 );
nand NAND2_23600 ( P3_ADD_547_U177 , P3_ADD_547_U112 , P3_ADD_547_U36 );
nand NAND2_23601 ( P3_ADD_547_U178 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_547_U33 );
nand NAND2_23602 ( P3_ADD_547_U179 , P3_ADD_547_U111 , P3_ADD_547_U34 );
nand NAND2_23603 ( P3_ADD_547_U180 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_547_U31 );
nand NAND2_23604 ( P3_ADD_547_U181 , P3_ADD_547_U110 , P3_ADD_547_U32 );
nand NAND2_23605 ( P3_ADD_547_U182 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_547_U29 );
nand NAND2_23606 ( P3_ADD_547_U183 , P3_ADD_547_U109 , P3_ADD_547_U30 );
nand NAND2_23607 ( P3_ADD_547_U184 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_547_U27 );
nand NAND2_23608 ( P3_ADD_547_U185 , P3_ADD_547_U108 , P3_ADD_547_U28 );
nand NAND2_23609 ( P3_ADD_547_U186 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_547_U25 );
nand NAND2_23610 ( P3_ADD_547_U187 , P3_ADD_547_U107 , P3_ADD_547_U26 );
nand NAND2_23611 ( P3_ADD_547_U188 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_547_U23 );
nand NAND2_23612 ( P3_ADD_547_U189 , P3_ADD_547_U106 , P3_ADD_547_U24 );
nand NAND2_23613 ( P3_SUB_412_U6 , P3_SUB_412_U43 , P3_SUB_412_U42 );
nand NAND2_23614 ( P3_SUB_412_U7 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_SUB_412_U27 );
not NOT1_23615 ( P3_SUB_412_U8 , P3_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_23616 ( P3_SUB_412_U9 , P3_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_23617 ( P3_SUB_412_U10 , P3_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_23618 ( P3_SUB_412_U11 , P3_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_23619 ( P3_SUB_412_U12 , P3_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_23620 ( P3_SUB_412_U13 , P3_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_23621 ( P3_SUB_412_U14 , P3_SUB_412_U39 , P3_SUB_412_U38 );
not NOT1_23622 ( P3_SUB_412_U15 , P3_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_23623 ( P3_SUB_412_U16 , P3_SUB_412_U48 , P3_SUB_412_U47 );
nand NAND2_23624 ( P3_SUB_412_U17 , P3_SUB_412_U53 , P3_SUB_412_U52 );
nand NAND2_23625 ( P3_SUB_412_U18 , P3_SUB_412_U58 , P3_SUB_412_U57 );
nand NAND2_23626 ( P3_SUB_412_U19 , P3_SUB_412_U63 , P3_SUB_412_U62 );
nand NAND2_23627 ( P3_SUB_412_U20 , P3_SUB_412_U45 , P3_SUB_412_U44 );
nand NAND2_23628 ( P3_SUB_412_U21 , P3_SUB_412_U50 , P3_SUB_412_U49 );
nand NAND2_23629 ( P3_SUB_412_U22 , P3_SUB_412_U55 , P3_SUB_412_U54 );
nand NAND2_23630 ( P3_SUB_412_U23 , P3_SUB_412_U60 , P3_SUB_412_U59 );
nand NAND2_23631 ( P3_SUB_412_U24 , P3_SUB_412_U35 , P3_SUB_412_U34 );
nand NAND2_23632 ( P3_SUB_412_U25 , P3_SUB_412_U31 , P3_SUB_412_U30 );
not NOT1_23633 ( P3_SUB_412_U26 , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_23634 ( P3_SUB_412_U27 , P3_INSTQUEUEWR_ADDR_REG_0_ );
not NOT1_23635 ( P3_SUB_412_U28 , P3_SUB_412_U7 );
nand NAND2_23636 ( P3_SUB_412_U29 , P3_SUB_412_U28 , P3_SUB_412_U8 );
nand NAND2_23637 ( P3_SUB_412_U30 , P3_SUB_412_U29 , P3_SUB_412_U26 );
nand NAND2_23638 ( P3_SUB_412_U31 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_412_U7 );
not NOT1_23639 ( P3_SUB_412_U32 , P3_SUB_412_U25 );
nand NAND2_23640 ( P3_SUB_412_U33 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_412_U10 );
nand NAND2_23641 ( P3_SUB_412_U34 , P3_SUB_412_U33 , P3_SUB_412_U25 );
nand NAND2_23642 ( P3_SUB_412_U35 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_412_U9 );
not NOT1_23643 ( P3_SUB_412_U36 , P3_SUB_412_U24 );
nand NAND2_23644 ( P3_SUB_412_U37 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_412_U12 );
nand NAND2_23645 ( P3_SUB_412_U38 , P3_SUB_412_U37 , P3_SUB_412_U24 );
nand NAND2_23646 ( P3_SUB_412_U39 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_412_U11 );
not NOT1_23647 ( P3_SUB_412_U40 , P3_SUB_412_U14 );
nand NAND2_23648 ( P3_SUB_412_U41 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_412_U15 );
nand NAND2_23649 ( P3_SUB_412_U42 , P3_SUB_412_U40 , P3_SUB_412_U41 );
nand NAND2_23650 ( P3_SUB_412_U43 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_412_U13 );
nand NAND2_23651 ( P3_SUB_412_U44 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_412_U13 );
nand NAND2_23652 ( P3_SUB_412_U45 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_412_U15 );
not NOT1_23653 ( P3_SUB_412_U46 , P3_SUB_412_U20 );
nand NAND2_23654 ( P3_SUB_412_U47 , P3_SUB_412_U46 , P3_SUB_412_U40 );
nand NAND2_23655 ( P3_SUB_412_U48 , P3_SUB_412_U20 , P3_SUB_412_U14 );
nand NAND2_23656 ( P3_SUB_412_U49 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_412_U12 );
nand NAND2_23657 ( P3_SUB_412_U50 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_412_U11 );
not NOT1_23658 ( P3_SUB_412_U51 , P3_SUB_412_U21 );
nand NAND2_23659 ( P3_SUB_412_U52 , P3_SUB_412_U36 , P3_SUB_412_U51 );
nand NAND2_23660 ( P3_SUB_412_U53 , P3_SUB_412_U21 , P3_SUB_412_U24 );
nand NAND2_23661 ( P3_SUB_412_U54 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_412_U10 );
nand NAND2_23662 ( P3_SUB_412_U55 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_412_U9 );
not NOT1_23663 ( P3_SUB_412_U56 , P3_SUB_412_U22 );
nand NAND2_23664 ( P3_SUB_412_U57 , P3_SUB_412_U32 , P3_SUB_412_U56 );
nand NAND2_23665 ( P3_SUB_412_U58 , P3_SUB_412_U22 , P3_SUB_412_U25 );
nand NAND2_23666 ( P3_SUB_412_U59 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_SUB_412_U8 );
nand NAND2_23667 ( P3_SUB_412_U60 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_412_U26 );
not NOT1_23668 ( P3_SUB_412_U61 , P3_SUB_412_U23 );
nand NAND2_23669 ( P3_SUB_412_U62 , P3_SUB_412_U61 , P3_SUB_412_U28 );
nand NAND2_23670 ( P3_SUB_412_U63 , P3_SUB_412_U23 , P3_SUB_412_U7 );
and AND2_23671 ( P3_ADD_371_1212_U4 , P3_ADD_371_1212_U133 , P3_ADD_371_1212_U132 );
and AND2_23672 ( P3_ADD_371_1212_U5 , P3_ADD_371_1212_U196 , P3_ADD_371_1212_U48 );
and AND2_23673 ( P3_ADD_371_1212_U6 , P3_ADD_371_1212_U194 , P3_ADD_371_1212_U49 );
and AND2_23674 ( P3_ADD_371_1212_U7 , P3_ADD_371_1212_U192 , P3_ADD_371_1212_U78 );
and AND2_23675 ( P3_ADD_371_1212_U8 , P3_ADD_371_1212_U191 , P3_ADD_371_1212_U53 );
and AND2_23676 ( P3_ADD_371_1212_U9 , P3_ADD_371_1212_U189 , P3_ADD_371_1212_U56 );
and AND2_23677 ( P3_ADD_371_1212_U10 , P3_ADD_371_1212_U187 , P3_ADD_371_1212_U59 );
and AND2_23678 ( P3_ADD_371_1212_U11 , P3_ADD_371_1212_U185 , P3_ADD_371_1212_U168 );
and AND2_23679 ( P3_ADD_371_1212_U12 , P3_ADD_371_1212_U184 , P3_ADD_371_1212_U62 );
and AND2_23680 ( P3_ADD_371_1212_U13 , P3_ADD_371_1212_U183 , P3_ADD_371_1212_U65 );
and AND2_23681 ( P3_ADD_371_1212_U14 , P3_ADD_371_1212_U181 , P3_ADD_371_1212_U68 );
and AND2_23682 ( P3_ADD_371_1212_U15 , P3_ADD_371_1212_U179 , P3_ADD_371_1212_U70 );
and AND2_23683 ( P3_ADD_371_1212_U16 , P3_ADD_371_1212_U178 , P3_ADD_371_1212_U73 );
and AND2_23684 ( P3_ADD_371_1212_U17 , P3_ADD_371_1212_U176 , P3_ADD_371_1212_U75 );
and AND2_23685 ( P3_ADD_371_1212_U18 , P3_ADD_371_1212_U162 , P3_ADD_371_1212_U159 );
and AND2_23686 ( P3_ADD_371_1212_U19 , P3_ADD_371_1212_U155 , P3_ADD_371_1212_U152 );
nand NAND3_23687 ( P3_ADD_371_1212_U20 , P3_ADD_371_1212_U255 , P3_ADD_371_1212_U254 , P3_ADD_371_1212_U203 );
not NOT1_23688 ( P3_ADD_371_1212_U21 , P3_ADD_371_U20 );
not NOT1_23689 ( P3_ADD_371_1212_U22 , P3_INSTADDRPOINTER_REG_4_ );
not NOT1_23690 ( P3_ADD_371_1212_U23 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_23691 ( P3_ADD_371_1212_U24 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_371_U20 );
not NOT1_23692 ( P3_ADD_371_1212_U25 , P3_ADD_371_U19 );
not NOT1_23693 ( P3_ADD_371_1212_U26 , P3_ADD_371_U5 );
not NOT1_23694 ( P3_ADD_371_1212_U27 , P3_INSTADDRPOINTER_REG_2_ );
not NOT1_23695 ( P3_ADD_371_1212_U28 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_23696 ( P3_ADD_371_1212_U29 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_371_U5 );
not NOT1_23697 ( P3_ADD_371_1212_U30 , P3_ADD_371_U25 );
not NOT1_23698 ( P3_ADD_371_1212_U31 , P3_ADD_371_U4 );
not NOT1_23699 ( P3_ADD_371_1212_U32 , P3_INSTADDRPOINTER_REG_0_ );
not NOT1_23700 ( P3_ADD_371_1212_U33 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_23701 ( P3_ADD_371_1212_U34 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_371_U4 );
not NOT1_23702 ( P3_ADD_371_1212_U35 , P3_ADD_371_U21 );
not NOT1_23703 ( P3_ADD_371_1212_U36 , P3_ADD_371_U18 );
not NOT1_23704 ( P3_ADD_371_1212_U37 , P3_INSTADDRPOINTER_REG_6_ );
not NOT1_23705 ( P3_ADD_371_1212_U38 , P3_INSTADDRPOINTER_REG_7_ );
not NOT1_23706 ( P3_ADD_371_1212_U39 , P3_ADD_371_U17 );
not NOT1_23707 ( P3_ADD_371_1212_U40 , P3_ADD_371_U6 );
not NOT1_23708 ( P3_ADD_371_1212_U41 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_23709 ( P3_ADD_371_1212_U42 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_23710 ( P3_ADD_371_1212_U43 , P3_ADD_371_1212_U94 , P3_ADD_371_1212_U130 );
nand NAND2_23711 ( P3_ADD_371_1212_U44 , P3_ADD_371_1212_U77 , P3_ADD_371_1212_U123 );
not NOT1_23712 ( P3_ADD_371_1212_U45 , P3_INSTADDRPOINTER_REG_10_ );
not NOT1_23713 ( P3_ADD_371_1212_U46 , P3_INSTADDRPOINTER_REG_11_ );
not NOT1_23714 ( P3_ADD_371_1212_U47 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_23715 ( P3_ADD_371_1212_U48 , P3_ADD_371_1212_U99 , P3_ADD_371_1212_U108 );
nand NAND2_23716 ( P3_ADD_371_1212_U49 , P3_ADD_371_1212_U100 , P3_ADD_371_1212_U117 );
not NOT1_23717 ( P3_ADD_371_1212_U50 , P3_INSTADDRPOINTER_REG_13_ );
not NOT1_23718 ( P3_ADD_371_1212_U51 , P3_INSTADDRPOINTER_REG_15_ );
not NOT1_23719 ( P3_ADD_371_1212_U52 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_23720 ( P3_ADD_371_1212_U53 , P3_ADD_371_1212_U163 , P3_ADD_371_1212_U101 );
not NOT1_23721 ( P3_ADD_371_1212_U54 , P3_INSTADDRPOINTER_REG_17_ );
not NOT1_23722 ( P3_ADD_371_1212_U55 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_23723 ( P3_ADD_371_1212_U56 , P3_ADD_371_1212_U102 , P3_ADD_371_1212_U165 );
not NOT1_23724 ( P3_ADD_371_1212_U57 , P3_INSTADDRPOINTER_REG_18_ );
not NOT1_23725 ( P3_ADD_371_1212_U58 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_23726 ( P3_ADD_371_1212_U59 , P3_ADD_371_1212_U103 , P3_ADD_371_1212_U166 );
not NOT1_23727 ( P3_ADD_371_1212_U60 , P3_INSTADDRPOINTER_REG_20_ );
not NOT1_23728 ( P3_ADD_371_1212_U61 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_23729 ( P3_ADD_371_1212_U62 , P3_ADD_371_1212_U104 , P3_ADD_371_1212_U167 );
not NOT1_23730 ( P3_ADD_371_1212_U63 , P3_INSTADDRPOINTER_REG_23_ );
not NOT1_23731 ( P3_ADD_371_1212_U64 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_23732 ( P3_ADD_371_1212_U65 , P3_ADD_371_1212_U105 , P3_ADD_371_1212_U169 );
not NOT1_23733 ( P3_ADD_371_1212_U66 , P3_INSTADDRPOINTER_REG_25_ );
not NOT1_23734 ( P3_ADD_371_1212_U67 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_23735 ( P3_ADD_371_1212_U68 , P3_ADD_371_1212_U106 , P3_ADD_371_1212_U170 );
not NOT1_23736 ( P3_ADD_371_1212_U69 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_23737 ( P3_ADD_371_1212_U70 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_371_1212_U171 );
not NOT1_23738 ( P3_ADD_371_1212_U71 , P3_INSTADDRPOINTER_REG_28_ );
not NOT1_23739 ( P3_ADD_371_1212_U72 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_23740 ( P3_ADD_371_1212_U73 , P3_ADD_371_1212_U107 , P3_ADD_371_1212_U172 );
not NOT1_23741 ( P3_ADD_371_1212_U74 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_23742 ( P3_ADD_371_1212_U75 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_371_1212_U173 );
not NOT1_23743 ( P3_ADD_371_1212_U76 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_23744 ( P3_ADD_371_1212_U77 , P3_ADD_371_U21 , P3_ADD_371_1212_U121 );
nand NAND2_23745 ( P3_ADD_371_1212_U78 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_371_1212_U163 );
nand NAND2_23746 ( P3_ADD_371_1212_U79 , P3_ADD_371_1212_U239 , P3_ADD_371_1212_U238 );
nand NAND2_23747 ( P3_ADD_371_1212_U80 , P3_ADD_371_1212_U246 , P3_ADD_371_1212_U245 );
nand NAND2_23748 ( P3_ADD_371_1212_U81 , P3_ADD_371_1212_U248 , P3_ADD_371_1212_U247 );
nand NAND2_23749 ( P3_ADD_371_1212_U82 , P3_ADD_371_1212_U250 , P3_ADD_371_1212_U249 );
nand NAND2_23750 ( P3_ADD_371_1212_U83 , P3_ADD_371_1212_U257 , P3_ADD_371_1212_U256 );
nand NAND2_23751 ( P3_ADD_371_1212_U84 , P3_ADD_371_1212_U259 , P3_ADD_371_1212_U258 );
nand NAND2_23752 ( P3_ADD_371_1212_U85 , P3_ADD_371_1212_U261 , P3_ADD_371_1212_U260 );
nand NAND2_23753 ( P3_ADD_371_1212_U86 , P3_ADD_371_1212_U263 , P3_ADD_371_1212_U262 );
nand NAND2_23754 ( P3_ADD_371_1212_U87 , P3_ADD_371_1212_U265 , P3_ADD_371_1212_U264 );
nand NAND2_23755 ( P3_ADD_371_1212_U88 , P3_ADD_371_1212_U212 , P3_ADD_371_1212_U211 );
nand NAND2_23756 ( P3_ADD_371_1212_U89 , P3_ADD_371_1212_U219 , P3_ADD_371_1212_U218 );
nand NAND2_23757 ( P3_ADD_371_1212_U90 , P3_ADD_371_1212_U226 , P3_ADD_371_1212_U225 );
nand NAND2_23758 ( P3_ADD_371_1212_U91 , P3_ADD_371_1212_U233 , P3_ADD_371_1212_U232 );
nand NAND2_23759 ( P3_ADD_371_1212_U92 , P3_ADD_371_1212_U237 , P3_ADD_371_1212_U236 );
nand NAND2_23760 ( P3_ADD_371_1212_U93 , P3_ADD_371_1212_U244 , P3_ADD_371_1212_U243 );
and AND2_23761 ( P3_ADD_371_1212_U94 , P3_ADD_371_1212_U129 , P3_ADD_371_1212_U128 );
and AND2_23762 ( P3_ADD_371_1212_U95 , P3_ADD_371_1212_U137 , P3_ADD_371_1212_U136 );
and AND3_23763 ( P3_ADD_371_1212_U96 , P3_ADD_371_1212_U228 , P3_ADD_371_1212_U227 , P3_ADD_371_1212_U24 );
and AND2_23764 ( P3_ADD_371_1212_U97 , P3_ADD_371_1212_U154 , P3_ADD_371_1212_U4 );
and AND3_23765 ( P3_ADD_371_1212_U98 , P3_ADD_371_1212_U235 , P3_ADD_371_1212_U234 , P3_ADD_371_1212_U29 );
and AND2_23766 ( P3_ADD_371_1212_U99 , P3_INSTADDRPOINTER_REG_9_ , P3_INSTADDRPOINTER_REG_10_ );
and AND2_23767 ( P3_ADD_371_1212_U100 , P3_INSTADDRPOINTER_REG_12_ , P3_INSTADDRPOINTER_REG_11_ );
and AND3_23768 ( P3_ADD_371_1212_U101 , P3_INSTADDRPOINTER_REG_14_ , P3_INSTADDRPOINTER_REG_15_ , P3_INSTADDRPOINTER_REG_13_ );
and AND2_23769 ( P3_ADD_371_1212_U102 , P3_INSTADDRPOINTER_REG_17_ , P3_INSTADDRPOINTER_REG_16_ );
and AND2_23770 ( P3_ADD_371_1212_U103 , P3_INSTADDRPOINTER_REG_18_ , P3_INSTADDRPOINTER_REG_19_ );
and AND2_23771 ( P3_ADD_371_1212_U104 , P3_INSTADDRPOINTER_REG_20_ , P3_INSTADDRPOINTER_REG_21_ );
and AND2_23772 ( P3_ADD_371_1212_U105 , P3_INSTADDRPOINTER_REG_23_ , P3_INSTADDRPOINTER_REG_22_ );
and AND2_23773 ( P3_ADD_371_1212_U106 , P3_INSTADDRPOINTER_REG_25_ , P3_INSTADDRPOINTER_REG_24_ );
and AND2_23774 ( P3_ADD_371_1212_U107 , P3_INSTADDRPOINTER_REG_28_ , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_23775 ( P3_ADD_371_1212_U108 , P3_ADD_371_1212_U148 , P3_ADD_371_1212_U147 );
and AND2_23776 ( P3_ADD_371_1212_U109 , P3_ADD_371_1212_U205 , P3_ADD_371_1212_U204 );
and AND2_23777 ( P3_ADD_371_1212_U110 , P3_ADD_371_1212_U207 , P3_ADD_371_1212_U206 );
nand NAND3_23778 ( P3_ADD_371_1212_U111 , P3_ADD_371_1212_U144 , P3_ADD_371_1212_U118 , P3_ADD_371_1212_U200 );
and AND2_23779 ( P3_ADD_371_1212_U112 , P3_ADD_371_1212_U214 , P3_ADD_371_1212_U213 );
nand NAND2_23780 ( P3_ADD_371_1212_U113 , P3_ADD_371_1212_U142 , P3_ADD_371_1212_U141 );
and AND2_23781 ( P3_ADD_371_1212_U114 , P3_ADD_371_1212_U221 , P3_ADD_371_1212_U220 );
nand NAND2_23782 ( P3_ADD_371_1212_U115 , P3_ADD_371_1212_U95 , P3_ADD_371_1212_U138 );
not NOT1_23783 ( P3_ADD_371_1212_U116 , P3_INSTADDRPOINTER_REG_31_ );
not NOT1_23784 ( P3_ADD_371_1212_U117 , P3_ADD_371_1212_U48 );
nand NAND2_23785 ( P3_ADD_371_1212_U118 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_371_1212_U113 );
nand NAND2_23786 ( P3_ADD_371_1212_U119 , P3_ADD_371_1212_U202 , P3_ADD_371_1212_U201 );
not NOT1_23787 ( P3_ADD_371_1212_U120 , P3_ADD_371_1212_U77 );
not NOT1_23788 ( P3_ADD_371_1212_U121 , P3_ADD_371_1212_U34 );
nand NAND2_23789 ( P3_ADD_371_1212_U122 , P3_ADD_371_1212_U35 , P3_ADD_371_1212_U34 );
nand NAND2_23790 ( P3_ADD_371_1212_U123 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_371_1212_U122 );
not NOT1_23791 ( P3_ADD_371_1212_U124 , P3_ADD_371_1212_U44 );
or OR2_23792 ( P3_ADD_371_1212_U125 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_371_U5 );
not NOT1_23793 ( P3_ADD_371_1212_U126 , P3_ADD_371_1212_U29 );
nand NAND2_23794 ( P3_ADD_371_1212_U127 , P3_ADD_371_1212_U30 , P3_ADD_371_1212_U29 );
nand NAND2_23795 ( P3_ADD_371_1212_U128 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_371_1212_U127 );
nand NAND2_23796 ( P3_ADD_371_1212_U129 , P3_ADD_371_U25 , P3_ADD_371_1212_U126 );
nand NAND2_23797 ( P3_ADD_371_1212_U130 , P3_ADD_371_1212_U44 , P3_ADD_371_1212_U119 );
not NOT1_23798 ( P3_ADD_371_1212_U131 , P3_ADD_371_1212_U43 );
or OR2_23799 ( P3_ADD_371_1212_U132 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_371_U19 );
or OR2_23800 ( P3_ADD_371_1212_U133 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_371_U20 );
not NOT1_23801 ( P3_ADD_371_1212_U134 , P3_ADD_371_1212_U24 );
nand NAND2_23802 ( P3_ADD_371_1212_U135 , P3_ADD_371_1212_U25 , P3_ADD_371_1212_U24 );
nand NAND2_23803 ( P3_ADD_371_1212_U136 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_371_1212_U135 );
nand NAND2_23804 ( P3_ADD_371_1212_U137 , P3_ADD_371_U19 , P3_ADD_371_1212_U134 );
nand NAND2_23805 ( P3_ADD_371_1212_U138 , P3_ADD_371_1212_U4 , P3_ADD_371_1212_U43 );
not NOT1_23806 ( P3_ADD_371_1212_U139 , P3_ADD_371_1212_U115 );
or OR2_23807 ( P3_ADD_371_1212_U140 , P3_ADD_371_U18 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_23808 ( P3_ADD_371_1212_U141 , P3_ADD_371_1212_U140 , P3_ADD_371_1212_U115 );
nand NAND2_23809 ( P3_ADD_371_1212_U142 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_371_U18 );
not NOT1_23810 ( P3_ADD_371_1212_U143 , P3_ADD_371_1212_U113 );
nand NAND2_23811 ( P3_ADD_371_1212_U144 , P3_ADD_371_U17 , P3_ADD_371_1212_U113 );
not NOT1_23812 ( P3_ADD_371_1212_U145 , P3_ADD_371_1212_U111 );
or OR2_23813 ( P3_ADD_371_1212_U146 , P3_ADD_371_U6 , P3_INSTADDRPOINTER_REG_8_ );
nand NAND2_23814 ( P3_ADD_371_1212_U147 , P3_ADD_371_1212_U146 , P3_ADD_371_1212_U111 );
nand NAND2_23815 ( P3_ADD_371_1212_U148 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_371_U6 );
not NOT1_23816 ( P3_ADD_371_1212_U149 , P3_ADD_371_1212_U108 );
or OR2_23817 ( P3_ADD_371_1212_U150 , P3_ADD_371_U20 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_23818 ( P3_ADD_371_1212_U151 , P3_ADD_371_1212_U150 , P3_ADD_371_1212_U43 );
nand NAND2_23819 ( P3_ADD_371_1212_U152 , P3_ADD_371_1212_U96 , P3_ADD_371_1212_U151 );
nand NAND2_23820 ( P3_ADD_371_1212_U153 , P3_ADD_371_1212_U131 , P3_ADD_371_1212_U24 );
nand NAND2_23821 ( P3_ADD_371_1212_U154 , P3_ADD_371_U19 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_23822 ( P3_ADD_371_1212_U155 , P3_ADD_371_1212_U97 , P3_ADD_371_1212_U153 );
or OR2_23823 ( P3_ADD_371_1212_U156 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_371_U20 );
or OR2_23824 ( P3_ADD_371_1212_U157 , P3_ADD_371_U5 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_23825 ( P3_ADD_371_1212_U158 , P3_ADD_371_1212_U157 , P3_ADD_371_1212_U44 );
nand NAND2_23826 ( P3_ADD_371_1212_U159 , P3_ADD_371_1212_U98 , P3_ADD_371_1212_U158 );
nand NAND2_23827 ( P3_ADD_371_1212_U160 , P3_ADD_371_1212_U124 , P3_ADD_371_1212_U29 );
nand NAND2_23828 ( P3_ADD_371_1212_U161 , P3_ADD_371_U25 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND3_23829 ( P3_ADD_371_1212_U162 , P3_ADD_371_1212_U160 , P3_ADD_371_1212_U161 , P3_ADD_371_1212_U119 );
not NOT1_23830 ( P3_ADD_371_1212_U163 , P3_ADD_371_1212_U49 );
not NOT1_23831 ( P3_ADD_371_1212_U164 , P3_ADD_371_1212_U78 );
not NOT1_23832 ( P3_ADD_371_1212_U165 , P3_ADD_371_1212_U53 );
not NOT1_23833 ( P3_ADD_371_1212_U166 , P3_ADD_371_1212_U56 );
not NOT1_23834 ( P3_ADD_371_1212_U167 , P3_ADD_371_1212_U59 );
nand NAND2_23835 ( P3_ADD_371_1212_U168 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_371_1212_U167 );
not NOT1_23836 ( P3_ADD_371_1212_U169 , P3_ADD_371_1212_U62 );
not NOT1_23837 ( P3_ADD_371_1212_U170 , P3_ADD_371_1212_U65 );
not NOT1_23838 ( P3_ADD_371_1212_U171 , P3_ADD_371_1212_U68 );
not NOT1_23839 ( P3_ADD_371_1212_U172 , P3_ADD_371_1212_U70 );
not NOT1_23840 ( P3_ADD_371_1212_U173 , P3_ADD_371_1212_U73 );
not NOT1_23841 ( P3_ADD_371_1212_U174 , P3_ADD_371_1212_U75 );
or OR2_23842 ( P3_ADD_371_1212_U175 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_371_U5 );
nand NAND2_23843 ( P3_ADD_371_1212_U176 , P3_ADD_371_1212_U74 , P3_ADD_371_1212_U73 );
nand NAND2_23844 ( P3_ADD_371_1212_U177 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_371_1212_U172 );
nand NAND2_23845 ( P3_ADD_371_1212_U178 , P3_ADD_371_1212_U71 , P3_ADD_371_1212_U177 );
nand NAND2_23846 ( P3_ADD_371_1212_U179 , P3_ADD_371_1212_U69 , P3_ADD_371_1212_U68 );
nand NAND2_23847 ( P3_ADD_371_1212_U180 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_371_1212_U170 );
nand NAND2_23848 ( P3_ADD_371_1212_U181 , P3_ADD_371_1212_U66 , P3_ADD_371_1212_U180 );
nand NAND2_23849 ( P3_ADD_371_1212_U182 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_371_1212_U169 );
nand NAND2_23850 ( P3_ADD_371_1212_U183 , P3_ADD_371_1212_U63 , P3_ADD_371_1212_U182 );
nand NAND2_23851 ( P3_ADD_371_1212_U184 , P3_ADD_371_1212_U61 , P3_ADD_371_1212_U168 );
nand NAND2_23852 ( P3_ADD_371_1212_U185 , P3_ADD_371_1212_U60 , P3_ADD_371_1212_U59 );
nand NAND2_23853 ( P3_ADD_371_1212_U186 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_371_1212_U166 );
nand NAND2_23854 ( P3_ADD_371_1212_U187 , P3_ADD_371_1212_U58 , P3_ADD_371_1212_U186 );
nand NAND2_23855 ( P3_ADD_371_1212_U188 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_371_1212_U165 );
nand NAND2_23856 ( P3_ADD_371_1212_U189 , P3_ADD_371_1212_U54 , P3_ADD_371_1212_U188 );
nand NAND2_23857 ( P3_ADD_371_1212_U190 , P3_ADD_371_1212_U164 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_23858 ( P3_ADD_371_1212_U191 , P3_ADD_371_1212_U51 , P3_ADD_371_1212_U190 );
nand NAND2_23859 ( P3_ADD_371_1212_U192 , P3_ADD_371_1212_U50 , P3_ADD_371_1212_U49 );
nand NAND2_23860 ( P3_ADD_371_1212_U193 , P3_ADD_371_1212_U117 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_23861 ( P3_ADD_371_1212_U194 , P3_ADD_371_1212_U47 , P3_ADD_371_1212_U193 );
nand NAND2_23862 ( P3_ADD_371_1212_U195 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_371_1212_U108 );
nand NAND2_23863 ( P3_ADD_371_1212_U196 , P3_ADD_371_1212_U45 , P3_ADD_371_1212_U195 );
nand NAND2_23864 ( P3_ADD_371_1212_U197 , P3_ADD_371_1212_U156 , P3_ADD_371_1212_U24 );
nand NAND2_23865 ( P3_ADD_371_1212_U198 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_371_1212_U174 );
nand NAND2_23866 ( P3_ADD_371_1212_U199 , P3_ADD_371_1212_U175 , P3_ADD_371_1212_U29 );
nand NAND2_23867 ( P3_ADD_371_1212_U200 , P3_ADD_371_U17 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_23868 ( P3_ADD_371_1212_U201 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_371_1212_U125 );
nand NAND2_23869 ( P3_ADD_371_1212_U202 , P3_ADD_371_U25 , P3_ADD_371_1212_U125 );
nand NAND2_23870 ( P3_ADD_371_1212_U203 , P3_ADD_371_1212_U120 , P3_INSTADDRPOINTER_REG_1_ );
nand NAND2_23871 ( P3_ADD_371_1212_U204 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_371_1212_U108 );
nand NAND2_23872 ( P3_ADD_371_1212_U205 , P3_ADD_371_1212_U149 , P3_ADD_371_1212_U42 );
nand NAND2_23873 ( P3_ADD_371_1212_U206 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_371_1212_U40 );
nand NAND2_23874 ( P3_ADD_371_1212_U207 , P3_ADD_371_U6 , P3_ADD_371_1212_U41 );
nand NAND2_23875 ( P3_ADD_371_1212_U208 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_371_1212_U40 );
nand NAND2_23876 ( P3_ADD_371_1212_U209 , P3_ADD_371_U6 , P3_ADD_371_1212_U41 );
nand NAND2_23877 ( P3_ADD_371_1212_U210 , P3_ADD_371_1212_U209 , P3_ADD_371_1212_U208 );
nand NAND2_23878 ( P3_ADD_371_1212_U211 , P3_ADD_371_1212_U110 , P3_ADD_371_1212_U111 );
nand NAND2_23879 ( P3_ADD_371_1212_U212 , P3_ADD_371_1212_U145 , P3_ADD_371_1212_U210 );
nand NAND2_23880 ( P3_ADD_371_1212_U213 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_371_1212_U39 );
nand NAND2_23881 ( P3_ADD_371_1212_U214 , P3_ADD_371_U17 , P3_ADD_371_1212_U38 );
nand NAND2_23882 ( P3_ADD_371_1212_U215 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_371_1212_U39 );
nand NAND2_23883 ( P3_ADD_371_1212_U216 , P3_ADD_371_U17 , P3_ADD_371_1212_U38 );
nand NAND2_23884 ( P3_ADD_371_1212_U217 , P3_ADD_371_1212_U216 , P3_ADD_371_1212_U215 );
nand NAND2_23885 ( P3_ADD_371_1212_U218 , P3_ADD_371_1212_U112 , P3_ADD_371_1212_U113 );
nand NAND2_23886 ( P3_ADD_371_1212_U219 , P3_ADD_371_1212_U143 , P3_ADD_371_1212_U217 );
nand NAND2_23887 ( P3_ADD_371_1212_U220 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_371_1212_U36 );
nand NAND2_23888 ( P3_ADD_371_1212_U221 , P3_ADD_371_U18 , P3_ADD_371_1212_U37 );
nand NAND2_23889 ( P3_ADD_371_1212_U222 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_371_1212_U36 );
nand NAND2_23890 ( P3_ADD_371_1212_U223 , P3_ADD_371_U18 , P3_ADD_371_1212_U37 );
nand NAND2_23891 ( P3_ADD_371_1212_U224 , P3_ADD_371_1212_U223 , P3_ADD_371_1212_U222 );
nand NAND2_23892 ( P3_ADD_371_1212_U225 , P3_ADD_371_1212_U114 , P3_ADD_371_1212_U115 );
nand NAND2_23893 ( P3_ADD_371_1212_U226 , P3_ADD_371_1212_U139 , P3_ADD_371_1212_U224 );
nand NAND2_23894 ( P3_ADD_371_1212_U227 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_371_1212_U25 );
nand NAND2_23895 ( P3_ADD_371_1212_U228 , P3_ADD_371_U19 , P3_ADD_371_1212_U23 );
nand NAND2_23896 ( P3_ADD_371_1212_U229 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_371_1212_U21 );
nand NAND2_23897 ( P3_ADD_371_1212_U230 , P3_ADD_371_U20 , P3_ADD_371_1212_U22 );
nand NAND2_23898 ( P3_ADD_371_1212_U231 , P3_ADD_371_1212_U230 , P3_ADD_371_1212_U229 );
nand NAND2_23899 ( P3_ADD_371_1212_U232 , P3_ADD_371_1212_U197 , P3_ADD_371_1212_U43 );
nand NAND2_23900 ( P3_ADD_371_1212_U233 , P3_ADD_371_1212_U231 , P3_ADD_371_1212_U131 );
nand NAND2_23901 ( P3_ADD_371_1212_U234 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_371_1212_U30 );
nand NAND2_23902 ( P3_ADD_371_1212_U235 , P3_ADD_371_U25 , P3_ADD_371_1212_U28 );
nand NAND2_23903 ( P3_ADD_371_1212_U236 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_371_1212_U198 );
nand NAND3_23904 ( P3_ADD_371_1212_U237 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_371_1212_U174 , P3_ADD_371_1212_U116 );
nand NAND2_23905 ( P3_ADD_371_1212_U238 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_371_1212_U75 );
nand NAND2_23906 ( P3_ADD_371_1212_U239 , P3_ADD_371_1212_U174 , P3_ADD_371_1212_U76 );
nand NAND2_23907 ( P3_ADD_371_1212_U240 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_371_1212_U26 );
nand NAND2_23908 ( P3_ADD_371_1212_U241 , P3_ADD_371_U5 , P3_ADD_371_1212_U27 );
nand NAND2_23909 ( P3_ADD_371_1212_U242 , P3_ADD_371_1212_U241 , P3_ADD_371_1212_U240 );
nand NAND2_23910 ( P3_ADD_371_1212_U243 , P3_ADD_371_1212_U199 , P3_ADD_371_1212_U44 );
nand NAND2_23911 ( P3_ADD_371_1212_U244 , P3_ADD_371_1212_U242 , P3_ADD_371_1212_U124 );
nand NAND2_23912 ( P3_ADD_371_1212_U245 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_371_1212_U70 );
nand NAND2_23913 ( P3_ADD_371_1212_U246 , P3_ADD_371_1212_U172 , P3_ADD_371_1212_U72 );
nand NAND2_23914 ( P3_ADD_371_1212_U247 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_371_1212_U65 );
nand NAND2_23915 ( P3_ADD_371_1212_U248 , P3_ADD_371_1212_U170 , P3_ADD_371_1212_U67 );
nand NAND2_23916 ( P3_ADD_371_1212_U249 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_371_1212_U62 );
nand NAND2_23917 ( P3_ADD_371_1212_U250 , P3_ADD_371_1212_U169 , P3_ADD_371_1212_U64 );
nand NAND2_23918 ( P3_ADD_371_1212_U251 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_371_1212_U34 );
nand NAND2_23919 ( P3_ADD_371_1212_U252 , P3_ADD_371_1212_U121 , P3_ADD_371_1212_U33 );
nand NAND2_23920 ( P3_ADD_371_1212_U253 , P3_ADD_371_1212_U252 , P3_ADD_371_1212_U251 );
nand NAND3_23921 ( P3_ADD_371_1212_U254 , P3_ADD_371_1212_U34 , P3_ADD_371_1212_U33 , P3_ADD_371_U21 );
nand NAND2_23922 ( P3_ADD_371_1212_U255 , P3_ADD_371_1212_U253 , P3_ADD_371_1212_U35 );
nand NAND2_23923 ( P3_ADD_371_1212_U256 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_371_1212_U56 );
nand NAND2_23924 ( P3_ADD_371_1212_U257 , P3_ADD_371_1212_U166 , P3_ADD_371_1212_U57 );
nand NAND2_23925 ( P3_ADD_371_1212_U258 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_371_1212_U53 );
nand NAND2_23926 ( P3_ADD_371_1212_U259 , P3_ADD_371_1212_U165 , P3_ADD_371_1212_U55 );
nand NAND2_23927 ( P3_ADD_371_1212_U260 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_371_1212_U78 );
nand NAND2_23928 ( P3_ADD_371_1212_U261 , P3_ADD_371_1212_U164 , P3_ADD_371_1212_U52 );
nand NAND2_23929 ( P3_ADD_371_1212_U262 , P3_ADD_371_1212_U117 , P3_ADD_371_1212_U46 );
nand NAND2_23930 ( P3_ADD_371_1212_U263 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_371_1212_U48 );
nand NAND2_23931 ( P3_ADD_371_1212_U264 , P3_INSTADDRPOINTER_REG_0_ , P3_ADD_371_1212_U31 );
nand NAND2_23932 ( P3_ADD_371_1212_U265 , P3_ADD_371_U4 , P3_ADD_371_1212_U32 );
nand NAND2_23933 ( P3_SUB_504_U6 , P3_SUB_504_U43 , P3_SUB_504_U42 );
nand NAND2_23934 ( P3_SUB_504_U7 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_SUB_504_U27 );
not NOT1_23935 ( P3_SUB_504_U8 , P3_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_23936 ( P3_SUB_504_U9 , P3_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_23937 ( P3_SUB_504_U10 , P3_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_23938 ( P3_SUB_504_U11 , P3_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_23939 ( P3_SUB_504_U12 , P3_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_23940 ( P3_SUB_504_U13 , P3_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_23941 ( P3_SUB_504_U14 , P3_SUB_504_U39 , P3_SUB_504_U38 );
not NOT1_23942 ( P3_SUB_504_U15 , P3_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_23943 ( P3_SUB_504_U16 , P3_SUB_504_U48 , P3_SUB_504_U47 );
nand NAND2_23944 ( P3_SUB_504_U17 , P3_SUB_504_U53 , P3_SUB_504_U52 );
nand NAND2_23945 ( P3_SUB_504_U18 , P3_SUB_504_U58 , P3_SUB_504_U57 );
nand NAND2_23946 ( P3_SUB_504_U19 , P3_SUB_504_U63 , P3_SUB_504_U62 );
nand NAND2_23947 ( P3_SUB_504_U20 , P3_SUB_504_U45 , P3_SUB_504_U44 );
nand NAND2_23948 ( P3_SUB_504_U21 , P3_SUB_504_U50 , P3_SUB_504_U49 );
nand NAND2_23949 ( P3_SUB_504_U22 , P3_SUB_504_U55 , P3_SUB_504_U54 );
nand NAND2_23950 ( P3_SUB_504_U23 , P3_SUB_504_U60 , P3_SUB_504_U59 );
nand NAND2_23951 ( P3_SUB_504_U24 , P3_SUB_504_U35 , P3_SUB_504_U34 );
nand NAND2_23952 ( P3_SUB_504_U25 , P3_SUB_504_U31 , P3_SUB_504_U30 );
not NOT1_23953 ( P3_SUB_504_U26 , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_23954 ( P3_SUB_504_U27 , P3_INSTQUEUEWR_ADDR_REG_0_ );
not NOT1_23955 ( P3_SUB_504_U28 , P3_SUB_504_U7 );
nand NAND2_23956 ( P3_SUB_504_U29 , P3_SUB_504_U28 , P3_SUB_504_U8 );
nand NAND2_23957 ( P3_SUB_504_U30 , P3_SUB_504_U29 , P3_SUB_504_U26 );
nand NAND2_23958 ( P3_SUB_504_U31 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_504_U7 );
not NOT1_23959 ( P3_SUB_504_U32 , P3_SUB_504_U25 );
nand NAND2_23960 ( P3_SUB_504_U33 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_504_U10 );
nand NAND2_23961 ( P3_SUB_504_U34 , P3_SUB_504_U33 , P3_SUB_504_U25 );
nand NAND2_23962 ( P3_SUB_504_U35 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_504_U9 );
not NOT1_23963 ( P3_SUB_504_U36 , P3_SUB_504_U24 );
nand NAND2_23964 ( P3_SUB_504_U37 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_504_U12 );
nand NAND2_23965 ( P3_SUB_504_U38 , P3_SUB_504_U37 , P3_SUB_504_U24 );
nand NAND2_23966 ( P3_SUB_504_U39 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_504_U11 );
not NOT1_23967 ( P3_SUB_504_U40 , P3_SUB_504_U14 );
nand NAND2_23968 ( P3_SUB_504_U41 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_504_U15 );
nand NAND2_23969 ( P3_SUB_504_U42 , P3_SUB_504_U40 , P3_SUB_504_U41 );
nand NAND2_23970 ( P3_SUB_504_U43 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_504_U13 );
nand NAND2_23971 ( P3_SUB_504_U44 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_504_U13 );
nand NAND2_23972 ( P3_SUB_504_U45 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_504_U15 );
not NOT1_23973 ( P3_SUB_504_U46 , P3_SUB_504_U20 );
nand NAND2_23974 ( P3_SUB_504_U47 , P3_SUB_504_U46 , P3_SUB_504_U40 );
nand NAND2_23975 ( P3_SUB_504_U48 , P3_SUB_504_U20 , P3_SUB_504_U14 );
nand NAND2_23976 ( P3_SUB_504_U49 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_504_U12 );
nand NAND2_23977 ( P3_SUB_504_U50 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_504_U11 );
not NOT1_23978 ( P3_SUB_504_U51 , P3_SUB_504_U21 );
nand NAND2_23979 ( P3_SUB_504_U52 , P3_SUB_504_U36 , P3_SUB_504_U51 );
nand NAND2_23980 ( P3_SUB_504_U53 , P3_SUB_504_U21 , P3_SUB_504_U24 );
nand NAND2_23981 ( P3_SUB_504_U54 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_504_U10 );
nand NAND2_23982 ( P3_SUB_504_U55 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_504_U9 );
not NOT1_23983 ( P3_SUB_504_U56 , P3_SUB_504_U22 );
nand NAND2_23984 ( P3_SUB_504_U57 , P3_SUB_504_U32 , P3_SUB_504_U56 );
nand NAND2_23985 ( P3_SUB_504_U58 , P3_SUB_504_U22 , P3_SUB_504_U25 );
nand NAND2_23986 ( P3_SUB_504_U59 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_SUB_504_U8 );
nand NAND2_23987 ( P3_SUB_504_U60 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_504_U26 );
not NOT1_23988 ( P3_SUB_504_U61 , P3_SUB_504_U23 );
nand NAND2_23989 ( P3_SUB_504_U62 , P3_SUB_504_U61 , P3_SUB_504_U28 );
nand NAND2_23990 ( P3_SUB_504_U63 , P3_SUB_504_U23 , P3_SUB_504_U7 );
nand NAND2_23991 ( P3_SUB_401_U6 , P3_SUB_401_U45 , P3_SUB_401_U44 );
nand NAND2_23992 ( P3_SUB_401_U7 , P3_SUB_401_U9 , P3_SUB_401_U46 );
not NOT1_23993 ( P3_SUB_401_U8 , P3_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_23994 ( P3_SUB_401_U9 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_SUB_401_U18 );
not NOT1_23995 ( P3_SUB_401_U10 , P3_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_23996 ( P3_SUB_401_U11 , P3_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_23997 ( P3_SUB_401_U12 , P3_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_23998 ( P3_SUB_401_U13 , P3_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_23999 ( P3_SUB_401_U14 , P3_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_24000 ( P3_SUB_401_U15 , P3_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_24001 ( P3_SUB_401_U16 , P3_SUB_401_U41 , P3_SUB_401_U40 );
not NOT1_24002 ( P3_SUB_401_U17 , P3_INSTQUEUERD_ADDR_REG_4_ );
not NOT1_24003 ( P3_SUB_401_U18 , P3_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_24004 ( P3_SUB_401_U19 , P3_SUB_401_U51 , P3_SUB_401_U50 );
nand NAND2_24005 ( P3_SUB_401_U20 , P3_SUB_401_U56 , P3_SUB_401_U55 );
nand NAND2_24006 ( P3_SUB_401_U21 , P3_SUB_401_U61 , P3_SUB_401_U60 );
nand NAND2_24007 ( P3_SUB_401_U22 , P3_SUB_401_U66 , P3_SUB_401_U65 );
nand NAND2_24008 ( P3_SUB_401_U23 , P3_SUB_401_U48 , P3_SUB_401_U47 );
nand NAND2_24009 ( P3_SUB_401_U24 , P3_SUB_401_U53 , P3_SUB_401_U52 );
nand NAND2_24010 ( P3_SUB_401_U25 , P3_SUB_401_U58 , P3_SUB_401_U57 );
nand NAND2_24011 ( P3_SUB_401_U26 , P3_SUB_401_U63 , P3_SUB_401_U62 );
nand NAND2_24012 ( P3_SUB_401_U27 , P3_SUB_401_U37 , P3_SUB_401_U36 );
nand NAND2_24013 ( P3_SUB_401_U28 , P3_SUB_401_U33 , P3_SUB_401_U32 );
not NOT1_24014 ( P3_SUB_401_U29 , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_24015 ( P3_SUB_401_U30 , P3_SUB_401_U9 );
nand NAND2_24016 ( P3_SUB_401_U31 , P3_SUB_401_U30 , P3_SUB_401_U10 );
nand NAND2_24017 ( P3_SUB_401_U32 , P3_SUB_401_U31 , P3_SUB_401_U29 );
nand NAND2_24018 ( P3_SUB_401_U33 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_401_U9 );
not NOT1_24019 ( P3_SUB_401_U34 , P3_SUB_401_U28 );
nand NAND2_24020 ( P3_SUB_401_U35 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_401_U12 );
nand NAND2_24021 ( P3_SUB_401_U36 , P3_SUB_401_U35 , P3_SUB_401_U28 );
nand NAND2_24022 ( P3_SUB_401_U37 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_401_U11 );
not NOT1_24023 ( P3_SUB_401_U38 , P3_SUB_401_U27 );
nand NAND2_24024 ( P3_SUB_401_U39 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_401_U14 );
nand NAND2_24025 ( P3_SUB_401_U40 , P3_SUB_401_U39 , P3_SUB_401_U27 );
nand NAND2_24026 ( P3_SUB_401_U41 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_401_U13 );
not NOT1_24027 ( P3_SUB_401_U42 , P3_SUB_401_U16 );
nand NAND2_24028 ( P3_SUB_401_U43 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_401_U17 );
nand NAND2_24029 ( P3_SUB_401_U44 , P3_SUB_401_U42 , P3_SUB_401_U43 );
nand NAND2_24030 ( P3_SUB_401_U45 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_401_U15 );
nand NAND2_24031 ( P3_SUB_401_U46 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_SUB_401_U8 );
nand NAND2_24032 ( P3_SUB_401_U47 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_401_U15 );
nand NAND2_24033 ( P3_SUB_401_U48 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_401_U17 );
not NOT1_24034 ( P3_SUB_401_U49 , P3_SUB_401_U23 );
nand NAND2_24035 ( P3_SUB_401_U50 , P3_SUB_401_U49 , P3_SUB_401_U42 );
nand NAND2_24036 ( P3_SUB_401_U51 , P3_SUB_401_U23 , P3_SUB_401_U16 );
nand NAND2_24037 ( P3_SUB_401_U52 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_401_U14 );
nand NAND2_24038 ( P3_SUB_401_U53 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_401_U13 );
not NOT1_24039 ( P3_SUB_401_U54 , P3_SUB_401_U24 );
nand NAND2_24040 ( P3_SUB_401_U55 , P3_SUB_401_U38 , P3_SUB_401_U54 );
nand NAND2_24041 ( P3_SUB_401_U56 , P3_SUB_401_U24 , P3_SUB_401_U27 );
nand NAND2_24042 ( P3_SUB_401_U57 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_401_U12 );
nand NAND2_24043 ( P3_SUB_401_U58 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_401_U11 );
not NOT1_24044 ( P3_SUB_401_U59 , P3_SUB_401_U25 );
nand NAND2_24045 ( P3_SUB_401_U60 , P3_SUB_401_U34 , P3_SUB_401_U59 );
nand NAND2_24046 ( P3_SUB_401_U61 , P3_SUB_401_U25 , P3_SUB_401_U28 );
nand NAND2_24047 ( P3_SUB_401_U62 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_SUB_401_U10 );
nand NAND2_24048 ( P3_SUB_401_U63 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_401_U29 );
not NOT1_24049 ( P3_SUB_401_U64 , P3_SUB_401_U26 );
nand NAND2_24050 ( P3_SUB_401_U65 , P3_SUB_401_U64 , P3_SUB_401_U30 );
nand NAND2_24051 ( P3_SUB_401_U66 , P3_SUB_401_U26 , P3_SUB_401_U9 );
not NOT1_24052 ( P3_ADD_371_U4 , P3_U2621 );
nand NAND2_24053 ( P3_ADD_371_U5 , P3_ADD_371_U24 , P3_ADD_371_U32 );
and AND2_24054 ( P3_ADD_371_U6 , P3_ADD_371_U22 , P3_ADD_371_U30 );
not NOT1_24055 ( P3_ADD_371_U7 , P3_U2622 );
not NOT1_24056 ( P3_ADD_371_U8 , P3_U2624 );
nand NAND2_24057 ( P3_ADD_371_U9 , P3_U2624 , P3_ADD_371_U24 );
not NOT1_24058 ( P3_ADD_371_U10 , P3_U2625 );
nand NAND2_24059 ( P3_ADD_371_U11 , P3_U2625 , P3_ADD_371_U28 );
not NOT1_24060 ( P3_ADD_371_U12 , P3_U2626 );
nand NAND2_24061 ( P3_ADD_371_U13 , P3_U2626 , P3_ADD_371_U29 );
not NOT1_24062 ( P3_ADD_371_U14 , P3_U2628 );
not NOT1_24063 ( P3_ADD_371_U15 , P3_U2627 );
not NOT1_24064 ( P3_ADD_371_U16 , P3_U2623 );
nand NAND2_24065 ( P3_ADD_371_U17 , P3_ADD_371_U34 , P3_ADD_371_U33 );
nand NAND2_24066 ( P3_ADD_371_U18 , P3_ADD_371_U36 , P3_ADD_371_U35 );
nand NAND2_24067 ( P3_ADD_371_U19 , P3_ADD_371_U38 , P3_ADD_371_U37 );
nand NAND2_24068 ( P3_ADD_371_U20 , P3_ADD_371_U40 , P3_ADD_371_U39 );
nand NAND2_24069 ( P3_ADD_371_U21 , P3_ADD_371_U44 , P3_ADD_371_U43 );
and AND2_24070 ( P3_ADD_371_U22 , P3_U2628 , P3_U2627 );
nand NAND2_24071 ( P3_ADD_371_U23 , P3_U2627 , P3_ADD_371_U30 );
nand NAND2_24072 ( P3_ADD_371_U24 , P3_ADD_371_U16 , P3_ADD_371_U26 );
and AND2_24073 ( P3_ADD_371_U25 , P3_ADD_371_U42 , P3_ADD_371_U41 );
nand NAND2_24074 ( P3_ADD_371_U26 , P3_U2622 , P3_U2621 );
not NOT1_24075 ( P3_ADD_371_U27 , P3_ADD_371_U24 );
not NOT1_24076 ( P3_ADD_371_U28 , P3_ADD_371_U9 );
not NOT1_24077 ( P3_ADD_371_U29 , P3_ADD_371_U11 );
not NOT1_24078 ( P3_ADD_371_U30 , P3_ADD_371_U13 );
not NOT1_24079 ( P3_ADD_371_U31 , P3_ADD_371_U23 );
nand NAND3_24080 ( P3_ADD_371_U32 , P3_U2622 , P3_U2621 , P3_U2623 );
nand NAND2_24081 ( P3_ADD_371_U33 , P3_U2628 , P3_ADD_371_U23 );
nand NAND2_24082 ( P3_ADD_371_U34 , P3_ADD_371_U31 , P3_ADD_371_U14 );
nand NAND2_24083 ( P3_ADD_371_U35 , P3_U2627 , P3_ADD_371_U13 );
nand NAND2_24084 ( P3_ADD_371_U36 , P3_ADD_371_U30 , P3_ADD_371_U15 );
nand NAND2_24085 ( P3_ADD_371_U37 , P3_U2626 , P3_ADD_371_U11 );
nand NAND2_24086 ( P3_ADD_371_U38 , P3_ADD_371_U29 , P3_ADD_371_U12 );
nand NAND2_24087 ( P3_ADD_371_U39 , P3_U2625 , P3_ADD_371_U9 );
nand NAND2_24088 ( P3_ADD_371_U40 , P3_ADD_371_U28 , P3_ADD_371_U10 );
nand NAND2_24089 ( P3_ADD_371_U41 , P3_U2624 , P3_ADD_371_U24 );
nand NAND2_24090 ( P3_ADD_371_U42 , P3_ADD_371_U27 , P3_ADD_371_U8 );
nand NAND2_24091 ( P3_ADD_371_U43 , P3_U2622 , P3_ADD_371_U4 );
nand NAND2_24092 ( P3_ADD_371_U44 , P3_U2621 , P3_ADD_371_U7 );
nand NAND2_24093 ( P3_SUB_390_U6 , P3_SUB_390_U45 , P3_SUB_390_U44 );
nand NAND2_24094 ( P3_SUB_390_U7 , P3_SUB_390_U9 , P3_SUB_390_U46 );
not NOT1_24095 ( P3_SUB_390_U8 , P3_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_24096 ( P3_SUB_390_U9 , P3_INSTQUEUERD_ADDR_REG_0_ , P3_SUB_390_U18 );
not NOT1_24097 ( P3_SUB_390_U10 , P3_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_24098 ( P3_SUB_390_U11 , P3_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_24099 ( P3_SUB_390_U12 , P3_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_24100 ( P3_SUB_390_U13 , P3_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_24101 ( P3_SUB_390_U14 , P3_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_24102 ( P3_SUB_390_U15 , P3_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_24103 ( P3_SUB_390_U16 , P3_SUB_390_U41 , P3_SUB_390_U40 );
not NOT1_24104 ( P3_SUB_390_U17 , P3_INSTQUEUERD_ADDR_REG_4_ );
not NOT1_24105 ( P3_SUB_390_U18 , P3_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_24106 ( P3_SUB_390_U19 , P3_SUB_390_U51 , P3_SUB_390_U50 );
nand NAND2_24107 ( P3_SUB_390_U20 , P3_SUB_390_U56 , P3_SUB_390_U55 );
nand NAND2_24108 ( P3_SUB_390_U21 , P3_SUB_390_U61 , P3_SUB_390_U60 );
nand NAND2_24109 ( P3_SUB_390_U22 , P3_SUB_390_U66 , P3_SUB_390_U65 );
nand NAND2_24110 ( P3_SUB_390_U23 , P3_SUB_390_U48 , P3_SUB_390_U47 );
nand NAND2_24111 ( P3_SUB_390_U24 , P3_SUB_390_U53 , P3_SUB_390_U52 );
nand NAND2_24112 ( P3_SUB_390_U25 , P3_SUB_390_U58 , P3_SUB_390_U57 );
nand NAND2_24113 ( P3_SUB_390_U26 , P3_SUB_390_U63 , P3_SUB_390_U62 );
nand NAND2_24114 ( P3_SUB_390_U27 , P3_SUB_390_U37 , P3_SUB_390_U36 );
nand NAND2_24115 ( P3_SUB_390_U28 , P3_SUB_390_U33 , P3_SUB_390_U32 );
not NOT1_24116 ( P3_SUB_390_U29 , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_24117 ( P3_SUB_390_U30 , P3_SUB_390_U9 );
nand NAND2_24118 ( P3_SUB_390_U31 , P3_SUB_390_U30 , P3_SUB_390_U10 );
nand NAND2_24119 ( P3_SUB_390_U32 , P3_SUB_390_U31 , P3_SUB_390_U29 );
nand NAND2_24120 ( P3_SUB_390_U33 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_390_U9 );
not NOT1_24121 ( P3_SUB_390_U34 , P3_SUB_390_U28 );
nand NAND2_24122 ( P3_SUB_390_U35 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_390_U12 );
nand NAND2_24123 ( P3_SUB_390_U36 , P3_SUB_390_U35 , P3_SUB_390_U28 );
nand NAND2_24124 ( P3_SUB_390_U37 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_390_U11 );
not NOT1_24125 ( P3_SUB_390_U38 , P3_SUB_390_U27 );
nand NAND2_24126 ( P3_SUB_390_U39 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_390_U14 );
nand NAND2_24127 ( P3_SUB_390_U40 , P3_SUB_390_U39 , P3_SUB_390_U27 );
nand NAND2_24128 ( P3_SUB_390_U41 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_390_U13 );
not NOT1_24129 ( P3_SUB_390_U42 , P3_SUB_390_U16 );
nand NAND2_24130 ( P3_SUB_390_U43 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_390_U17 );
nand NAND2_24131 ( P3_SUB_390_U44 , P3_SUB_390_U42 , P3_SUB_390_U43 );
nand NAND2_24132 ( P3_SUB_390_U45 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_390_U15 );
nand NAND2_24133 ( P3_SUB_390_U46 , P3_INSTQUEUEWR_ADDR_REG_0_ , P3_SUB_390_U8 );
nand NAND2_24134 ( P3_SUB_390_U47 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_SUB_390_U15 );
nand NAND2_24135 ( P3_SUB_390_U48 , P3_INSTQUEUEWR_ADDR_REG_4_ , P3_SUB_390_U17 );
not NOT1_24136 ( P3_SUB_390_U49 , P3_SUB_390_U23 );
nand NAND2_24137 ( P3_SUB_390_U50 , P3_SUB_390_U49 , P3_SUB_390_U42 );
nand NAND2_24138 ( P3_SUB_390_U51 , P3_SUB_390_U23 , P3_SUB_390_U16 );
nand NAND2_24139 ( P3_SUB_390_U52 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_SUB_390_U14 );
nand NAND2_24140 ( P3_SUB_390_U53 , P3_INSTQUEUEWR_ADDR_REG_3_ , P3_SUB_390_U13 );
not NOT1_24141 ( P3_SUB_390_U54 , P3_SUB_390_U24 );
nand NAND2_24142 ( P3_SUB_390_U55 , P3_SUB_390_U38 , P3_SUB_390_U54 );
nand NAND2_24143 ( P3_SUB_390_U56 , P3_SUB_390_U24 , P3_SUB_390_U27 );
nand NAND2_24144 ( P3_SUB_390_U57 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_SUB_390_U12 );
nand NAND2_24145 ( P3_SUB_390_U58 , P3_INSTQUEUEWR_ADDR_REG_2_ , P3_SUB_390_U11 );
not NOT1_24146 ( P3_SUB_390_U59 , P3_SUB_390_U25 );
nand NAND2_24147 ( P3_SUB_390_U60 , P3_SUB_390_U34 , P3_SUB_390_U59 );
nand NAND2_24148 ( P3_SUB_390_U61 , P3_SUB_390_U25 , P3_SUB_390_U28 );
nand NAND2_24149 ( P3_SUB_390_U62 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_SUB_390_U10 );
nand NAND2_24150 ( P3_SUB_390_U63 , P3_INSTQUEUEWR_ADDR_REG_1_ , P3_SUB_390_U29 );
not NOT1_24151 ( P3_SUB_390_U64 , P3_SUB_390_U26 );
nand NAND2_24152 ( P3_SUB_390_U65 , P3_SUB_390_U64 , P3_SUB_390_U30 );
nand NAND2_24153 ( P3_SUB_390_U66 , P3_SUB_390_U26 , P3_SUB_390_U9 );
not NOT1_24154 ( P3_SUB_357_U6 , P3_U2627 );
not NOT1_24155 ( P3_SUB_357_U7 , P3_U2622 );
not NOT1_24156 ( P3_SUB_357_U8 , P3_U2628 );
not NOT1_24157 ( P3_SUB_357_U9 , P3_U2626 );
not NOT1_24158 ( P3_SUB_357_U10 , P3_U2621 );
not NOT1_24159 ( P3_SUB_357_U11 , P3_U2624 );
not NOT1_24160 ( P3_SUB_357_U12 , P3_U2623 );
not NOT1_24161 ( P3_SUB_357_U13 , P3_U2625 );
not NOT1_24162 ( P3_ADD_495_U4 , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_24163 ( P3_ADD_495_U5 , P3_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_24164 ( P3_ADD_495_U6 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_24165 ( P3_ADD_495_U7 , P3_INSTQUEUERD_ADDR_REG_3_ );
nand NAND2_24166 ( P3_ADD_495_U8 , P3_ADD_495_U16 , P3_ADD_495_U15 );
nand NAND2_24167 ( P3_ADD_495_U9 , P3_ADD_495_U18 , P3_ADD_495_U17 );
nand NAND2_24168 ( P3_ADD_495_U10 , P3_ADD_495_U20 , P3_ADD_495_U19 );
not NOT1_24169 ( P3_ADD_495_U11 , P3_INSTQUEUERD_ADDR_REG_4_ );
nand NAND2_24170 ( P3_ADD_495_U12 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_ADD_495_U13 );
not NOT1_24171 ( P3_ADD_495_U13 , P3_ADD_495_U6 );
not NOT1_24172 ( P3_ADD_495_U14 , P3_ADD_495_U12 );
nand NAND2_24173 ( P3_ADD_495_U15 , P3_INSTQUEUERD_ADDR_REG_4_ , P3_ADD_495_U12 );
nand NAND2_24174 ( P3_ADD_495_U16 , P3_ADD_495_U14 , P3_ADD_495_U11 );
nand NAND2_24175 ( P3_ADD_495_U17 , P3_INSTQUEUERD_ADDR_REG_3_ , P3_ADD_495_U6 );
nand NAND2_24176 ( P3_ADD_495_U18 , P3_ADD_495_U13 , P3_ADD_495_U7 );
nand NAND2_24177 ( P3_ADD_495_U19 , P3_INSTQUEUERD_ADDR_REG_2_ , P3_ADD_495_U4 );
nand NAND2_24178 ( P3_ADD_495_U20 , P3_INSTQUEUERD_ADDR_REG_1_ , P3_ADD_495_U5 );
nor nor_24179 ( P3_GTE_412_U6 , P3_SUB_412_U6 , P3_GTE_412_U7 );
nor nor_24180 ( P3_GTE_412_U7 , P3_SUB_412_U16 , P3_SUB_412_U17 , P3_SUB_412_U19 , P3_SUB_412_U18 );
nor nor_24181 ( P3_GTE_504_U6 , P3_SUB_504_U6 , P3_GTE_504_U7 );
nor nor_24182 ( P3_GTE_504_U7 , P3_SUB_504_U16 , P3_SUB_504_U17 , P3_SUB_504_U19 , P3_SUB_504_U18 );
not NOT1_24183 ( P3_ADD_494_U4 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_24184 ( P3_ADD_494_U5 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_24185 ( P3_ADD_494_U6 , P3_INSTADDRPOINTER_REG_2_ , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_24186 ( P3_ADD_494_U7 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_24187 ( P3_ADD_494_U8 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_494_U94 );
not NOT1_24188 ( P3_ADD_494_U9 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_24189 ( P3_ADD_494_U10 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_494_U95 );
not NOT1_24190 ( P3_ADD_494_U11 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_24191 ( P3_ADD_494_U12 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_494_U96 );
not NOT1_24192 ( P3_ADD_494_U13 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_24193 ( P3_ADD_494_U14 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_494_U97 );
not NOT1_24194 ( P3_ADD_494_U15 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_24195 ( P3_ADD_494_U16 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_494_U98 );
not NOT1_24196 ( P3_ADD_494_U17 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_24197 ( P3_ADD_494_U18 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_24198 ( P3_ADD_494_U19 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_494_U99 );
nand NAND2_24199 ( P3_ADD_494_U20 , P3_ADD_494_U100 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_24200 ( P3_ADD_494_U21 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_24201 ( P3_ADD_494_U22 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_494_U101 );
not NOT1_24202 ( P3_ADD_494_U23 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_24203 ( P3_ADD_494_U24 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_494_U102 );
not NOT1_24204 ( P3_ADD_494_U25 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_24205 ( P3_ADD_494_U26 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_494_U103 );
not NOT1_24206 ( P3_ADD_494_U27 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_24207 ( P3_ADD_494_U28 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_494_U104 );
not NOT1_24208 ( P3_ADD_494_U29 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_24209 ( P3_ADD_494_U30 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_494_U105 );
not NOT1_24210 ( P3_ADD_494_U31 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_24211 ( P3_ADD_494_U32 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_494_U106 );
not NOT1_24212 ( P3_ADD_494_U33 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_24213 ( P3_ADD_494_U34 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_494_U107 );
not NOT1_24214 ( P3_ADD_494_U35 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_24215 ( P3_ADD_494_U36 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_494_U108 );
not NOT1_24216 ( P3_ADD_494_U37 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_24217 ( P3_ADD_494_U38 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_494_U109 );
not NOT1_24218 ( P3_ADD_494_U39 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_24219 ( P3_ADD_494_U40 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_494_U110 );
not NOT1_24220 ( P3_ADD_494_U41 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_24221 ( P3_ADD_494_U42 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_494_U111 );
not NOT1_24222 ( P3_ADD_494_U43 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_24223 ( P3_ADD_494_U44 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_494_U112 );
not NOT1_24224 ( P3_ADD_494_U45 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_24225 ( P3_ADD_494_U46 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_494_U113 );
not NOT1_24226 ( P3_ADD_494_U47 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_24227 ( P3_ADD_494_U48 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_494_U114 );
not NOT1_24228 ( P3_ADD_494_U49 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_24229 ( P3_ADD_494_U50 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_494_U115 );
not NOT1_24230 ( P3_ADD_494_U51 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_24231 ( P3_ADD_494_U52 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_494_U116 );
not NOT1_24232 ( P3_ADD_494_U53 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_24233 ( P3_ADD_494_U54 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_494_U117 );
not NOT1_24234 ( P3_ADD_494_U55 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_24235 ( P3_ADD_494_U56 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_494_U118 );
not NOT1_24236 ( P3_ADD_494_U57 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_24237 ( P3_ADD_494_U58 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_494_U119 );
not NOT1_24238 ( P3_ADD_494_U59 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_24239 ( P3_ADD_494_U60 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_494_U120 );
not NOT1_24240 ( P3_ADD_494_U61 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_24241 ( P3_ADD_494_U62 , P3_ADD_494_U124 , P3_ADD_494_U123 );
nand NAND2_24242 ( P3_ADD_494_U63 , P3_ADD_494_U126 , P3_ADD_494_U125 );
nand NAND2_24243 ( P3_ADD_494_U64 , P3_ADD_494_U128 , P3_ADD_494_U127 );
nand NAND2_24244 ( P3_ADD_494_U65 , P3_ADD_494_U130 , P3_ADD_494_U129 );
nand NAND2_24245 ( P3_ADD_494_U66 , P3_ADD_494_U132 , P3_ADD_494_U131 );
nand NAND2_24246 ( P3_ADD_494_U67 , P3_ADD_494_U134 , P3_ADD_494_U133 );
nand NAND2_24247 ( P3_ADD_494_U68 , P3_ADD_494_U136 , P3_ADD_494_U135 );
nand NAND2_24248 ( P3_ADD_494_U69 , P3_ADD_494_U138 , P3_ADD_494_U137 );
nand NAND2_24249 ( P3_ADD_494_U70 , P3_ADD_494_U140 , P3_ADD_494_U139 );
nand NAND2_24250 ( P3_ADD_494_U71 , P3_ADD_494_U142 , P3_ADD_494_U141 );
nand NAND2_24251 ( P3_ADD_494_U72 , P3_ADD_494_U144 , P3_ADD_494_U143 );
nand NAND2_24252 ( P3_ADD_494_U73 , P3_ADD_494_U146 , P3_ADD_494_U145 );
nand NAND2_24253 ( P3_ADD_494_U74 , P3_ADD_494_U148 , P3_ADD_494_U147 );
nand NAND2_24254 ( P3_ADD_494_U75 , P3_ADD_494_U150 , P3_ADD_494_U149 );
nand NAND2_24255 ( P3_ADD_494_U76 , P3_ADD_494_U152 , P3_ADD_494_U151 );
nand NAND2_24256 ( P3_ADD_494_U77 , P3_ADD_494_U154 , P3_ADD_494_U153 );
nand NAND2_24257 ( P3_ADD_494_U78 , P3_ADD_494_U156 , P3_ADD_494_U155 );
nand NAND2_24258 ( P3_ADD_494_U79 , P3_ADD_494_U158 , P3_ADD_494_U157 );
nand NAND2_24259 ( P3_ADD_494_U80 , P3_ADD_494_U160 , P3_ADD_494_U159 );
nand NAND2_24260 ( P3_ADD_494_U81 , P3_ADD_494_U162 , P3_ADD_494_U161 );
nand NAND2_24261 ( P3_ADD_494_U82 , P3_ADD_494_U164 , P3_ADD_494_U163 );
nand NAND2_24262 ( P3_ADD_494_U83 , P3_ADD_494_U166 , P3_ADD_494_U165 );
nand NAND2_24263 ( P3_ADD_494_U84 , P3_ADD_494_U168 , P3_ADD_494_U167 );
nand NAND2_24264 ( P3_ADD_494_U85 , P3_ADD_494_U170 , P3_ADD_494_U169 );
nand NAND2_24265 ( P3_ADD_494_U86 , P3_ADD_494_U172 , P3_ADD_494_U171 );
nand NAND2_24266 ( P3_ADD_494_U87 , P3_ADD_494_U174 , P3_ADD_494_U173 );
nand NAND2_24267 ( P3_ADD_494_U88 , P3_ADD_494_U176 , P3_ADD_494_U175 );
nand NAND2_24268 ( P3_ADD_494_U89 , P3_ADD_494_U178 , P3_ADD_494_U177 );
nand NAND2_24269 ( P3_ADD_494_U90 , P3_ADD_494_U180 , P3_ADD_494_U179 );
nand NAND2_24270 ( P3_ADD_494_U91 , P3_ADD_494_U182 , P3_ADD_494_U181 );
not NOT1_24271 ( P3_ADD_494_U92 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_24272 ( P3_ADD_494_U93 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_494_U121 );
not NOT1_24273 ( P3_ADD_494_U94 , P3_ADD_494_U6 );
not NOT1_24274 ( P3_ADD_494_U95 , P3_ADD_494_U8 );
not NOT1_24275 ( P3_ADD_494_U96 , P3_ADD_494_U10 );
not NOT1_24276 ( P3_ADD_494_U97 , P3_ADD_494_U12 );
not NOT1_24277 ( P3_ADD_494_U98 , P3_ADD_494_U14 );
not NOT1_24278 ( P3_ADD_494_U99 , P3_ADD_494_U16 );
not NOT1_24279 ( P3_ADD_494_U100 , P3_ADD_494_U19 );
not NOT1_24280 ( P3_ADD_494_U101 , P3_ADD_494_U20 );
not NOT1_24281 ( P3_ADD_494_U102 , P3_ADD_494_U22 );
not NOT1_24282 ( P3_ADD_494_U103 , P3_ADD_494_U24 );
not NOT1_24283 ( P3_ADD_494_U104 , P3_ADD_494_U26 );
not NOT1_24284 ( P3_ADD_494_U105 , P3_ADD_494_U28 );
not NOT1_24285 ( P3_ADD_494_U106 , P3_ADD_494_U30 );
not NOT1_24286 ( P3_ADD_494_U107 , P3_ADD_494_U32 );
not NOT1_24287 ( P3_ADD_494_U108 , P3_ADD_494_U34 );
not NOT1_24288 ( P3_ADD_494_U109 , P3_ADD_494_U36 );
not NOT1_24289 ( P3_ADD_494_U110 , P3_ADD_494_U38 );
not NOT1_24290 ( P3_ADD_494_U111 , P3_ADD_494_U40 );
not NOT1_24291 ( P3_ADD_494_U112 , P3_ADD_494_U42 );
not NOT1_24292 ( P3_ADD_494_U113 , P3_ADD_494_U44 );
not NOT1_24293 ( P3_ADD_494_U114 , P3_ADD_494_U46 );
not NOT1_24294 ( P3_ADD_494_U115 , P3_ADD_494_U48 );
not NOT1_24295 ( P3_ADD_494_U116 , P3_ADD_494_U50 );
not NOT1_24296 ( P3_ADD_494_U117 , P3_ADD_494_U52 );
not NOT1_24297 ( P3_ADD_494_U118 , P3_ADD_494_U54 );
not NOT1_24298 ( P3_ADD_494_U119 , P3_ADD_494_U56 );
not NOT1_24299 ( P3_ADD_494_U120 , P3_ADD_494_U58 );
not NOT1_24300 ( P3_ADD_494_U121 , P3_ADD_494_U60 );
not NOT1_24301 ( P3_ADD_494_U122 , P3_ADD_494_U93 );
nand NAND2_24302 ( P3_ADD_494_U123 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_494_U19 );
nand NAND2_24303 ( P3_ADD_494_U124 , P3_ADD_494_U100 , P3_ADD_494_U18 );
nand NAND2_24304 ( P3_ADD_494_U125 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_494_U16 );
nand NAND2_24305 ( P3_ADD_494_U126 , P3_ADD_494_U99 , P3_ADD_494_U17 );
nand NAND2_24306 ( P3_ADD_494_U127 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_494_U14 );
nand NAND2_24307 ( P3_ADD_494_U128 , P3_ADD_494_U98 , P3_ADD_494_U15 );
nand NAND2_24308 ( P3_ADD_494_U129 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_494_U12 );
nand NAND2_24309 ( P3_ADD_494_U130 , P3_ADD_494_U97 , P3_ADD_494_U13 );
nand NAND2_24310 ( P3_ADD_494_U131 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_494_U10 );
nand NAND2_24311 ( P3_ADD_494_U132 , P3_ADD_494_U96 , P3_ADD_494_U11 );
nand NAND2_24312 ( P3_ADD_494_U133 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_494_U8 );
nand NAND2_24313 ( P3_ADD_494_U134 , P3_ADD_494_U95 , P3_ADD_494_U9 );
nand NAND2_24314 ( P3_ADD_494_U135 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_494_U6 );
nand NAND2_24315 ( P3_ADD_494_U136 , P3_ADD_494_U94 , P3_ADD_494_U7 );
nand NAND2_24316 ( P3_ADD_494_U137 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_494_U93 );
nand NAND2_24317 ( P3_ADD_494_U138 , P3_ADD_494_U122 , P3_ADD_494_U92 );
nand NAND2_24318 ( P3_ADD_494_U139 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_494_U60 );
nand NAND2_24319 ( P3_ADD_494_U140 , P3_ADD_494_U121 , P3_ADD_494_U61 );
nand NAND2_24320 ( P3_ADD_494_U141 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_494_U4 );
nand NAND2_24321 ( P3_ADD_494_U142 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_494_U5 );
nand NAND2_24322 ( P3_ADD_494_U143 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_494_U58 );
nand NAND2_24323 ( P3_ADD_494_U144 , P3_ADD_494_U120 , P3_ADD_494_U59 );
nand NAND2_24324 ( P3_ADD_494_U145 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_494_U56 );
nand NAND2_24325 ( P3_ADD_494_U146 , P3_ADD_494_U119 , P3_ADD_494_U57 );
nand NAND2_24326 ( P3_ADD_494_U147 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_494_U54 );
nand NAND2_24327 ( P3_ADD_494_U148 , P3_ADD_494_U118 , P3_ADD_494_U55 );
nand NAND2_24328 ( P3_ADD_494_U149 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_494_U52 );
nand NAND2_24329 ( P3_ADD_494_U150 , P3_ADD_494_U117 , P3_ADD_494_U53 );
nand NAND2_24330 ( P3_ADD_494_U151 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_494_U50 );
nand NAND2_24331 ( P3_ADD_494_U152 , P3_ADD_494_U116 , P3_ADD_494_U51 );
nand NAND2_24332 ( P3_ADD_494_U153 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_494_U48 );
nand NAND2_24333 ( P3_ADD_494_U154 , P3_ADD_494_U115 , P3_ADD_494_U49 );
nand NAND2_24334 ( P3_ADD_494_U155 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_494_U46 );
nand NAND2_24335 ( P3_ADD_494_U156 , P3_ADD_494_U114 , P3_ADD_494_U47 );
nand NAND2_24336 ( P3_ADD_494_U157 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_494_U44 );
nand NAND2_24337 ( P3_ADD_494_U158 , P3_ADD_494_U113 , P3_ADD_494_U45 );
nand NAND2_24338 ( P3_ADD_494_U159 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_494_U42 );
nand NAND2_24339 ( P3_ADD_494_U160 , P3_ADD_494_U112 , P3_ADD_494_U43 );
nand NAND2_24340 ( P3_ADD_494_U161 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_494_U40 );
nand NAND2_24341 ( P3_ADD_494_U162 , P3_ADD_494_U111 , P3_ADD_494_U41 );
nand NAND2_24342 ( P3_ADD_494_U163 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_494_U38 );
nand NAND2_24343 ( P3_ADD_494_U164 , P3_ADD_494_U110 , P3_ADD_494_U39 );
nand NAND2_24344 ( P3_ADD_494_U165 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_494_U36 );
nand NAND2_24345 ( P3_ADD_494_U166 , P3_ADD_494_U109 , P3_ADD_494_U37 );
nand NAND2_24346 ( P3_ADD_494_U167 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_494_U34 );
nand NAND2_24347 ( P3_ADD_494_U168 , P3_ADD_494_U108 , P3_ADD_494_U35 );
nand NAND2_24348 ( P3_ADD_494_U169 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_494_U32 );
nand NAND2_24349 ( P3_ADD_494_U170 , P3_ADD_494_U107 , P3_ADD_494_U33 );
nand NAND2_24350 ( P3_ADD_494_U171 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_494_U30 );
nand NAND2_24351 ( P3_ADD_494_U172 , P3_ADD_494_U106 , P3_ADD_494_U31 );
nand NAND2_24352 ( P3_ADD_494_U173 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_494_U28 );
nand NAND2_24353 ( P3_ADD_494_U174 , P3_ADD_494_U105 , P3_ADD_494_U29 );
nand NAND2_24354 ( P3_ADD_494_U175 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_494_U26 );
nand NAND2_24355 ( P3_ADD_494_U176 , P3_ADD_494_U104 , P3_ADD_494_U27 );
nand NAND2_24356 ( P3_ADD_494_U177 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_494_U24 );
nand NAND2_24357 ( P3_ADD_494_U178 , P3_ADD_494_U103 , P3_ADD_494_U25 );
nand NAND2_24358 ( P3_ADD_494_U179 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_494_U22 );
nand NAND2_24359 ( P3_ADD_494_U180 , P3_ADD_494_U102 , P3_ADD_494_U23 );
nand NAND2_24360 ( P3_ADD_494_U181 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_494_U20 );
nand NAND2_24361 ( P3_ADD_494_U182 , P3_ADD_494_U101 , P3_ADD_494_U21 );
not NOT1_24362 ( P3_ADD_536_U4 , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_24363 ( P3_ADD_536_U5 , P3_INSTADDRPOINTER_REG_2_ );
nand NAND2_24364 ( P3_ADD_536_U6 , P3_INSTADDRPOINTER_REG_2_ , P3_INSTADDRPOINTER_REG_1_ );
not NOT1_24365 ( P3_ADD_536_U7 , P3_INSTADDRPOINTER_REG_3_ );
nand NAND2_24366 ( P3_ADD_536_U8 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_536_U94 );
not NOT1_24367 ( P3_ADD_536_U9 , P3_INSTADDRPOINTER_REG_4_ );
nand NAND2_24368 ( P3_ADD_536_U10 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_536_U95 );
not NOT1_24369 ( P3_ADD_536_U11 , P3_INSTADDRPOINTER_REG_5_ );
nand NAND2_24370 ( P3_ADD_536_U12 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_536_U96 );
not NOT1_24371 ( P3_ADD_536_U13 , P3_INSTADDRPOINTER_REG_6_ );
nand NAND2_24372 ( P3_ADD_536_U14 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_536_U97 );
not NOT1_24373 ( P3_ADD_536_U15 , P3_INSTADDRPOINTER_REG_7_ );
nand NAND2_24374 ( P3_ADD_536_U16 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_536_U98 );
not NOT1_24375 ( P3_ADD_536_U17 , P3_INSTADDRPOINTER_REG_8_ );
not NOT1_24376 ( P3_ADD_536_U18 , P3_INSTADDRPOINTER_REG_9_ );
nand NAND2_24377 ( P3_ADD_536_U19 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_536_U99 );
nand NAND2_24378 ( P3_ADD_536_U20 , P3_ADD_536_U100 , P3_INSTADDRPOINTER_REG_9_ );
not NOT1_24379 ( P3_ADD_536_U21 , P3_INSTADDRPOINTER_REG_10_ );
nand NAND2_24380 ( P3_ADD_536_U22 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_536_U101 );
not NOT1_24381 ( P3_ADD_536_U23 , P3_INSTADDRPOINTER_REG_11_ );
nand NAND2_24382 ( P3_ADD_536_U24 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_536_U102 );
not NOT1_24383 ( P3_ADD_536_U25 , P3_INSTADDRPOINTER_REG_12_ );
nand NAND2_24384 ( P3_ADD_536_U26 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_536_U103 );
not NOT1_24385 ( P3_ADD_536_U27 , P3_INSTADDRPOINTER_REG_13_ );
nand NAND2_24386 ( P3_ADD_536_U28 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_536_U104 );
not NOT1_24387 ( P3_ADD_536_U29 , P3_INSTADDRPOINTER_REG_14_ );
nand NAND2_24388 ( P3_ADD_536_U30 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_536_U105 );
not NOT1_24389 ( P3_ADD_536_U31 , P3_INSTADDRPOINTER_REG_15_ );
nand NAND2_24390 ( P3_ADD_536_U32 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_536_U106 );
not NOT1_24391 ( P3_ADD_536_U33 , P3_INSTADDRPOINTER_REG_16_ );
nand NAND2_24392 ( P3_ADD_536_U34 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_536_U107 );
not NOT1_24393 ( P3_ADD_536_U35 , P3_INSTADDRPOINTER_REG_17_ );
nand NAND2_24394 ( P3_ADD_536_U36 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_536_U108 );
not NOT1_24395 ( P3_ADD_536_U37 , P3_INSTADDRPOINTER_REG_18_ );
nand NAND2_24396 ( P3_ADD_536_U38 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_536_U109 );
not NOT1_24397 ( P3_ADD_536_U39 , P3_INSTADDRPOINTER_REG_19_ );
nand NAND2_24398 ( P3_ADD_536_U40 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_536_U110 );
not NOT1_24399 ( P3_ADD_536_U41 , P3_INSTADDRPOINTER_REG_20_ );
nand NAND2_24400 ( P3_ADD_536_U42 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_536_U111 );
not NOT1_24401 ( P3_ADD_536_U43 , P3_INSTADDRPOINTER_REG_21_ );
nand NAND2_24402 ( P3_ADD_536_U44 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_536_U112 );
not NOT1_24403 ( P3_ADD_536_U45 , P3_INSTADDRPOINTER_REG_22_ );
nand NAND2_24404 ( P3_ADD_536_U46 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_536_U113 );
not NOT1_24405 ( P3_ADD_536_U47 , P3_INSTADDRPOINTER_REG_23_ );
nand NAND2_24406 ( P3_ADD_536_U48 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_536_U114 );
not NOT1_24407 ( P3_ADD_536_U49 , P3_INSTADDRPOINTER_REG_24_ );
nand NAND2_24408 ( P3_ADD_536_U50 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_536_U115 );
not NOT1_24409 ( P3_ADD_536_U51 , P3_INSTADDRPOINTER_REG_25_ );
nand NAND2_24410 ( P3_ADD_536_U52 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_536_U116 );
not NOT1_24411 ( P3_ADD_536_U53 , P3_INSTADDRPOINTER_REG_26_ );
nand NAND2_24412 ( P3_ADD_536_U54 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_536_U117 );
not NOT1_24413 ( P3_ADD_536_U55 , P3_INSTADDRPOINTER_REG_27_ );
nand NAND2_24414 ( P3_ADD_536_U56 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_536_U118 );
not NOT1_24415 ( P3_ADD_536_U57 , P3_INSTADDRPOINTER_REG_28_ );
nand NAND2_24416 ( P3_ADD_536_U58 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_536_U119 );
not NOT1_24417 ( P3_ADD_536_U59 , P3_INSTADDRPOINTER_REG_29_ );
nand NAND2_24418 ( P3_ADD_536_U60 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_536_U120 );
not NOT1_24419 ( P3_ADD_536_U61 , P3_INSTADDRPOINTER_REG_30_ );
nand NAND2_24420 ( P3_ADD_536_U62 , P3_ADD_536_U124 , P3_ADD_536_U123 );
nand NAND2_24421 ( P3_ADD_536_U63 , P3_ADD_536_U126 , P3_ADD_536_U125 );
nand NAND2_24422 ( P3_ADD_536_U64 , P3_ADD_536_U128 , P3_ADD_536_U127 );
nand NAND2_24423 ( P3_ADD_536_U65 , P3_ADD_536_U130 , P3_ADD_536_U129 );
nand NAND2_24424 ( P3_ADD_536_U66 , P3_ADD_536_U132 , P3_ADD_536_U131 );
nand NAND2_24425 ( P3_ADD_536_U67 , P3_ADD_536_U134 , P3_ADD_536_U133 );
nand NAND2_24426 ( P3_ADD_536_U68 , P3_ADD_536_U136 , P3_ADD_536_U135 );
nand NAND2_24427 ( P3_ADD_536_U69 , P3_ADD_536_U138 , P3_ADD_536_U137 );
nand NAND2_24428 ( P3_ADD_536_U70 , P3_ADD_536_U140 , P3_ADD_536_U139 );
nand NAND2_24429 ( P3_ADD_536_U71 , P3_ADD_536_U142 , P3_ADD_536_U141 );
nand NAND2_24430 ( P3_ADD_536_U72 , P3_ADD_536_U144 , P3_ADD_536_U143 );
nand NAND2_24431 ( P3_ADD_536_U73 , P3_ADD_536_U146 , P3_ADD_536_U145 );
nand NAND2_24432 ( P3_ADD_536_U74 , P3_ADD_536_U148 , P3_ADD_536_U147 );
nand NAND2_24433 ( P3_ADD_536_U75 , P3_ADD_536_U150 , P3_ADD_536_U149 );
nand NAND2_24434 ( P3_ADD_536_U76 , P3_ADD_536_U152 , P3_ADD_536_U151 );
nand NAND2_24435 ( P3_ADD_536_U77 , P3_ADD_536_U154 , P3_ADD_536_U153 );
nand NAND2_24436 ( P3_ADD_536_U78 , P3_ADD_536_U156 , P3_ADD_536_U155 );
nand NAND2_24437 ( P3_ADD_536_U79 , P3_ADD_536_U158 , P3_ADD_536_U157 );
nand NAND2_24438 ( P3_ADD_536_U80 , P3_ADD_536_U160 , P3_ADD_536_U159 );
nand NAND2_24439 ( P3_ADD_536_U81 , P3_ADD_536_U162 , P3_ADD_536_U161 );
nand NAND2_24440 ( P3_ADD_536_U82 , P3_ADD_536_U164 , P3_ADD_536_U163 );
nand NAND2_24441 ( P3_ADD_536_U83 , P3_ADD_536_U166 , P3_ADD_536_U165 );
nand NAND2_24442 ( P3_ADD_536_U84 , P3_ADD_536_U168 , P3_ADD_536_U167 );
nand NAND2_24443 ( P3_ADD_536_U85 , P3_ADD_536_U170 , P3_ADD_536_U169 );
nand NAND2_24444 ( P3_ADD_536_U86 , P3_ADD_536_U172 , P3_ADD_536_U171 );
nand NAND2_24445 ( P3_ADD_536_U87 , P3_ADD_536_U174 , P3_ADD_536_U173 );
nand NAND2_24446 ( P3_ADD_536_U88 , P3_ADD_536_U176 , P3_ADD_536_U175 );
nand NAND2_24447 ( P3_ADD_536_U89 , P3_ADD_536_U178 , P3_ADD_536_U177 );
nand NAND2_24448 ( P3_ADD_536_U90 , P3_ADD_536_U180 , P3_ADD_536_U179 );
nand NAND2_24449 ( P3_ADD_536_U91 , P3_ADD_536_U182 , P3_ADD_536_U181 );
not NOT1_24450 ( P3_ADD_536_U92 , P3_INSTADDRPOINTER_REG_31_ );
nand NAND2_24451 ( P3_ADD_536_U93 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_536_U121 );
not NOT1_24452 ( P3_ADD_536_U94 , P3_ADD_536_U6 );
not NOT1_24453 ( P3_ADD_536_U95 , P3_ADD_536_U8 );
not NOT1_24454 ( P3_ADD_536_U96 , P3_ADD_536_U10 );
not NOT1_24455 ( P3_ADD_536_U97 , P3_ADD_536_U12 );
not NOT1_24456 ( P3_ADD_536_U98 , P3_ADD_536_U14 );
not NOT1_24457 ( P3_ADD_536_U99 , P3_ADD_536_U16 );
not NOT1_24458 ( P3_ADD_536_U100 , P3_ADD_536_U19 );
not NOT1_24459 ( P3_ADD_536_U101 , P3_ADD_536_U20 );
not NOT1_24460 ( P3_ADD_536_U102 , P3_ADD_536_U22 );
not NOT1_24461 ( P3_ADD_536_U103 , P3_ADD_536_U24 );
not NOT1_24462 ( P3_ADD_536_U104 , P3_ADD_536_U26 );
not NOT1_24463 ( P3_ADD_536_U105 , P3_ADD_536_U28 );
not NOT1_24464 ( P3_ADD_536_U106 , P3_ADD_536_U30 );
not NOT1_24465 ( P3_ADD_536_U107 , P3_ADD_536_U32 );
not NOT1_24466 ( P3_ADD_536_U108 , P3_ADD_536_U34 );
not NOT1_24467 ( P3_ADD_536_U109 , P3_ADD_536_U36 );
not NOT1_24468 ( P3_ADD_536_U110 , P3_ADD_536_U38 );
not NOT1_24469 ( P3_ADD_536_U111 , P3_ADD_536_U40 );
not NOT1_24470 ( P3_ADD_536_U112 , P3_ADD_536_U42 );
not NOT1_24471 ( P3_ADD_536_U113 , P3_ADD_536_U44 );
not NOT1_24472 ( P3_ADD_536_U114 , P3_ADD_536_U46 );
not NOT1_24473 ( P3_ADD_536_U115 , P3_ADD_536_U48 );
not NOT1_24474 ( P3_ADD_536_U116 , P3_ADD_536_U50 );
not NOT1_24475 ( P3_ADD_536_U117 , P3_ADD_536_U52 );
not NOT1_24476 ( P3_ADD_536_U118 , P3_ADD_536_U54 );
not NOT1_24477 ( P3_ADD_536_U119 , P3_ADD_536_U56 );
not NOT1_24478 ( P3_ADD_536_U120 , P3_ADD_536_U58 );
not NOT1_24479 ( P3_ADD_536_U121 , P3_ADD_536_U60 );
not NOT1_24480 ( P3_ADD_536_U122 , P3_ADD_536_U93 );
nand NAND2_24481 ( P3_ADD_536_U123 , P3_INSTADDRPOINTER_REG_9_ , P3_ADD_536_U19 );
nand NAND2_24482 ( P3_ADD_536_U124 , P3_ADD_536_U100 , P3_ADD_536_U18 );
nand NAND2_24483 ( P3_ADD_536_U125 , P3_INSTADDRPOINTER_REG_8_ , P3_ADD_536_U16 );
nand NAND2_24484 ( P3_ADD_536_U126 , P3_ADD_536_U99 , P3_ADD_536_U17 );
nand NAND2_24485 ( P3_ADD_536_U127 , P3_INSTADDRPOINTER_REG_7_ , P3_ADD_536_U14 );
nand NAND2_24486 ( P3_ADD_536_U128 , P3_ADD_536_U98 , P3_ADD_536_U15 );
nand NAND2_24487 ( P3_ADD_536_U129 , P3_INSTADDRPOINTER_REG_6_ , P3_ADD_536_U12 );
nand NAND2_24488 ( P3_ADD_536_U130 , P3_ADD_536_U97 , P3_ADD_536_U13 );
nand NAND2_24489 ( P3_ADD_536_U131 , P3_INSTADDRPOINTER_REG_5_ , P3_ADD_536_U10 );
nand NAND2_24490 ( P3_ADD_536_U132 , P3_ADD_536_U96 , P3_ADD_536_U11 );
nand NAND2_24491 ( P3_ADD_536_U133 , P3_INSTADDRPOINTER_REG_4_ , P3_ADD_536_U8 );
nand NAND2_24492 ( P3_ADD_536_U134 , P3_ADD_536_U95 , P3_ADD_536_U9 );
nand NAND2_24493 ( P3_ADD_536_U135 , P3_INSTADDRPOINTER_REG_3_ , P3_ADD_536_U6 );
nand NAND2_24494 ( P3_ADD_536_U136 , P3_ADD_536_U94 , P3_ADD_536_U7 );
nand NAND2_24495 ( P3_ADD_536_U137 , P3_INSTADDRPOINTER_REG_31_ , P3_ADD_536_U93 );
nand NAND2_24496 ( P3_ADD_536_U138 , P3_ADD_536_U122 , P3_ADD_536_U92 );
nand NAND2_24497 ( P3_ADD_536_U139 , P3_INSTADDRPOINTER_REG_30_ , P3_ADD_536_U60 );
nand NAND2_24498 ( P3_ADD_536_U140 , P3_ADD_536_U121 , P3_ADD_536_U61 );
nand NAND2_24499 ( P3_ADD_536_U141 , P3_INSTADDRPOINTER_REG_2_ , P3_ADD_536_U4 );
nand NAND2_24500 ( P3_ADD_536_U142 , P3_INSTADDRPOINTER_REG_1_ , P3_ADD_536_U5 );
nand NAND2_24501 ( P3_ADD_536_U143 , P3_INSTADDRPOINTER_REG_29_ , P3_ADD_536_U58 );
nand NAND2_24502 ( P3_ADD_536_U144 , P3_ADD_536_U120 , P3_ADD_536_U59 );
nand NAND2_24503 ( P3_ADD_536_U145 , P3_INSTADDRPOINTER_REG_28_ , P3_ADD_536_U56 );
nand NAND2_24504 ( P3_ADD_536_U146 , P3_ADD_536_U119 , P3_ADD_536_U57 );
nand NAND2_24505 ( P3_ADD_536_U147 , P3_INSTADDRPOINTER_REG_27_ , P3_ADD_536_U54 );
nand NAND2_24506 ( P3_ADD_536_U148 , P3_ADD_536_U118 , P3_ADD_536_U55 );
nand NAND2_24507 ( P3_ADD_536_U149 , P3_INSTADDRPOINTER_REG_26_ , P3_ADD_536_U52 );
nand NAND2_24508 ( P3_ADD_536_U150 , P3_ADD_536_U117 , P3_ADD_536_U53 );
nand NAND2_24509 ( P3_ADD_536_U151 , P3_INSTADDRPOINTER_REG_25_ , P3_ADD_536_U50 );
nand NAND2_24510 ( P3_ADD_536_U152 , P3_ADD_536_U116 , P3_ADD_536_U51 );
nand NAND2_24511 ( P3_ADD_536_U153 , P3_INSTADDRPOINTER_REG_24_ , P3_ADD_536_U48 );
nand NAND2_24512 ( P3_ADD_536_U154 , P3_ADD_536_U115 , P3_ADD_536_U49 );
nand NAND2_24513 ( P3_ADD_536_U155 , P3_INSTADDRPOINTER_REG_23_ , P3_ADD_536_U46 );
nand NAND2_24514 ( P3_ADD_536_U156 , P3_ADD_536_U114 , P3_ADD_536_U47 );
nand NAND2_24515 ( P3_ADD_536_U157 , P3_INSTADDRPOINTER_REG_22_ , P3_ADD_536_U44 );
nand NAND2_24516 ( P3_ADD_536_U158 , P3_ADD_536_U113 , P3_ADD_536_U45 );
nand NAND2_24517 ( P3_ADD_536_U159 , P3_INSTADDRPOINTER_REG_21_ , P3_ADD_536_U42 );
nand NAND2_24518 ( P3_ADD_536_U160 , P3_ADD_536_U112 , P3_ADD_536_U43 );
nand NAND2_24519 ( P3_ADD_536_U161 , P3_INSTADDRPOINTER_REG_20_ , P3_ADD_536_U40 );
nand NAND2_24520 ( P3_ADD_536_U162 , P3_ADD_536_U111 , P3_ADD_536_U41 );
nand NAND2_24521 ( P3_ADD_536_U163 , P3_INSTADDRPOINTER_REG_19_ , P3_ADD_536_U38 );
nand NAND2_24522 ( P3_ADD_536_U164 , P3_ADD_536_U110 , P3_ADD_536_U39 );
nand NAND2_24523 ( P3_ADD_536_U165 , P3_INSTADDRPOINTER_REG_18_ , P3_ADD_536_U36 );
nand NAND2_24524 ( P3_ADD_536_U166 , P3_ADD_536_U109 , P3_ADD_536_U37 );
nand NAND2_24525 ( P3_ADD_536_U167 , P3_INSTADDRPOINTER_REG_17_ , P3_ADD_536_U34 );
nand NAND2_24526 ( P3_ADD_536_U168 , P3_ADD_536_U108 , P3_ADD_536_U35 );
nand NAND2_24527 ( P3_ADD_536_U169 , P3_INSTADDRPOINTER_REG_16_ , P3_ADD_536_U32 );
nand NAND2_24528 ( P3_ADD_536_U170 , P3_ADD_536_U107 , P3_ADD_536_U33 );
nand NAND2_24529 ( P3_ADD_536_U171 , P3_INSTADDRPOINTER_REG_15_ , P3_ADD_536_U30 );
nand NAND2_24530 ( P3_ADD_536_U172 , P3_ADD_536_U106 , P3_ADD_536_U31 );
nand NAND2_24531 ( P3_ADD_536_U173 , P3_INSTADDRPOINTER_REG_14_ , P3_ADD_536_U28 );
nand NAND2_24532 ( P3_ADD_536_U174 , P3_ADD_536_U105 , P3_ADD_536_U29 );
nand NAND2_24533 ( P3_ADD_536_U175 , P3_INSTADDRPOINTER_REG_13_ , P3_ADD_536_U26 );
nand NAND2_24534 ( P3_ADD_536_U176 , P3_ADD_536_U104 , P3_ADD_536_U27 );
nand NAND2_24535 ( P3_ADD_536_U177 , P3_INSTADDRPOINTER_REG_12_ , P3_ADD_536_U24 );
nand NAND2_24536 ( P3_ADD_536_U178 , P3_ADD_536_U103 , P3_ADD_536_U25 );
nand NAND2_24537 ( P3_ADD_536_U179 , P3_INSTADDRPOINTER_REG_11_ , P3_ADD_536_U22 );
nand NAND2_24538 ( P3_ADD_536_U180 , P3_ADD_536_U102 , P3_ADD_536_U23 );
nand NAND2_24539 ( P3_ADD_536_U181 , P3_INSTADDRPOINTER_REG_10_ , P3_ADD_536_U20 );
nand NAND2_24540 ( P3_ADD_536_U182 , P3_ADD_536_U101 , P3_ADD_536_U21 );
not NOT1_24541 ( P3_ADD_402_1132_U4 , P3_U2613 );
not NOT1_24542 ( P3_ADD_402_1132_U5 , P3_U3069 );
nand NAND2_24543 ( P3_ADD_402_1132_U6 , P3_U3069 , P3_U2613 );
not NOT1_24544 ( P3_ADD_402_1132_U7 , P3_U2614 );
nand NAND2_24545 ( P3_ADD_402_1132_U8 , P3_U2614 , P3_ADD_402_1132_U28 );
not NOT1_24546 ( P3_ADD_402_1132_U9 , P3_U2615 );
nand NAND2_24547 ( P3_ADD_402_1132_U10 , P3_U2615 , P3_ADD_402_1132_U29 );
not NOT1_24548 ( P3_ADD_402_1132_U11 , P3_U2616 );
nand NAND2_24549 ( P3_ADD_402_1132_U12 , P3_U2616 , P3_ADD_402_1132_U30 );
not NOT1_24550 ( P3_ADD_402_1132_U13 , P3_U2617 );
nand NAND2_24551 ( P3_ADD_402_1132_U14 , P3_U2617 , P3_ADD_402_1132_U31 );
not NOT1_24552 ( P3_ADD_402_1132_U15 , P3_U2618 );
nand NAND2_24553 ( P3_ADD_402_1132_U16 , P3_U2618 , P3_ADD_402_1132_U32 );
not NOT1_24554 ( P3_ADD_402_1132_U17 , P3_U2619 );
nand NAND2_24555 ( P3_ADD_402_1132_U18 , P3_ADD_402_1132_U36 , P3_ADD_402_1132_U35 );
nand NAND2_24556 ( P3_ADD_402_1132_U19 , P3_ADD_402_1132_U38 , P3_ADD_402_1132_U37 );
nand NAND2_24557 ( P3_ADD_402_1132_U20 , P3_ADD_402_1132_U40 , P3_ADD_402_1132_U39 );
nand NAND2_24558 ( P3_ADD_402_1132_U21 , P3_ADD_402_1132_U42 , P3_ADD_402_1132_U41 );
nand NAND2_24559 ( P3_ADD_402_1132_U22 , P3_ADD_402_1132_U44 , P3_ADD_402_1132_U43 );
nand NAND2_24560 ( P3_ADD_402_1132_U23 , P3_ADD_402_1132_U46 , P3_ADD_402_1132_U45 );
nand NAND2_24561 ( P3_ADD_402_1132_U24 , P3_ADD_402_1132_U48 , P3_ADD_402_1132_U47 );
nand NAND2_24562 ( P3_ADD_402_1132_U25 , P3_ADD_402_1132_U50 , P3_ADD_402_1132_U49 );
not NOT1_24563 ( P3_ADD_402_1132_U26 , P3_U2620 );
nand NAND2_24564 ( P3_ADD_402_1132_U27 , P3_U2619 , P3_ADD_402_1132_U33 );
not NOT1_24565 ( P3_ADD_402_1132_U28 , P3_ADD_402_1132_U6 );
not NOT1_24566 ( P3_ADD_402_1132_U29 , P3_ADD_402_1132_U8 );
not NOT1_24567 ( P3_ADD_402_1132_U30 , P3_ADD_402_1132_U10 );
not NOT1_24568 ( P3_ADD_402_1132_U31 , P3_ADD_402_1132_U12 );
not NOT1_24569 ( P3_ADD_402_1132_U32 , P3_ADD_402_1132_U14 );
not NOT1_24570 ( P3_ADD_402_1132_U33 , P3_ADD_402_1132_U16 );
not NOT1_24571 ( P3_ADD_402_1132_U34 , P3_ADD_402_1132_U27 );
nand NAND2_24572 ( P3_ADD_402_1132_U35 , P3_U2620 , P3_ADD_402_1132_U27 );
nand NAND2_24573 ( P3_ADD_402_1132_U36 , P3_ADD_402_1132_U34 , P3_ADD_402_1132_U26 );
nand NAND2_24574 ( P3_ADD_402_1132_U37 , P3_U2619 , P3_ADD_402_1132_U16 );
nand NAND2_24575 ( P3_ADD_402_1132_U38 , P3_ADD_402_1132_U33 , P3_ADD_402_1132_U17 );
nand NAND2_24576 ( P3_ADD_402_1132_U39 , P3_U2618 , P3_ADD_402_1132_U14 );
nand NAND2_24577 ( P3_ADD_402_1132_U40 , P3_ADD_402_1132_U32 , P3_ADD_402_1132_U15 );
nand NAND2_24578 ( P3_ADD_402_1132_U41 , P3_U2617 , P3_ADD_402_1132_U12 );
nand NAND2_24579 ( P3_ADD_402_1132_U42 , P3_ADD_402_1132_U31 , P3_ADD_402_1132_U13 );
nand NAND2_24580 ( P3_ADD_402_1132_U43 , P3_U2616 , P3_ADD_402_1132_U10 );
nand NAND2_24581 ( P3_ADD_402_1132_U44 , P3_ADD_402_1132_U30 , P3_ADD_402_1132_U11 );
nand NAND2_24582 ( P3_ADD_402_1132_U45 , P3_U2615 , P3_ADD_402_1132_U8 );
nand NAND2_24583 ( P3_ADD_402_1132_U46 , P3_ADD_402_1132_U29 , P3_ADD_402_1132_U9 );
nand NAND2_24584 ( P3_ADD_402_1132_U47 , P3_U2614 , P3_ADD_402_1132_U6 );
nand NAND2_24585 ( P3_ADD_402_1132_U48 , P3_ADD_402_1132_U28 , P3_ADD_402_1132_U7 );
nand NAND2_24586 ( P3_ADD_402_1132_U49 , P3_U3069 , P3_ADD_402_1132_U4 );
nand NAND2_24587 ( P3_ADD_402_1132_U50 , P3_U2613 , P3_ADD_402_1132_U5 );
nand NAND2_24588 ( P2_R2099_U5 , P2_R2099_U107 , P2_R2099_U148 );
not NOT1_24589 ( P2_R2099_U6 , P2_U2747 );
not NOT1_24590 ( P2_R2099_U7 , P2_U2751 );
not NOT1_24591 ( P2_R2099_U8 , P2_U2750 );
not NOT1_24592 ( P2_R2099_U9 , P2_U2746 );
not NOT1_24593 ( P2_R2099_U10 , P2_U2749 );
not NOT1_24594 ( P2_R2099_U11 , P2_U2745 );
not NOT1_24595 ( P2_R2099_U12 , P2_U2748 );
not NOT1_24596 ( P2_R2099_U13 , P2_U2744 );
not NOT1_24597 ( P2_R2099_U14 , P2_U2743 );
nand NAND2_24598 ( P2_R2099_U15 , P2_U2743 , P2_R2099_U97 );
not NOT1_24599 ( P2_R2099_U16 , P2_U2742 );
nand NAND2_24600 ( P2_R2099_U17 , P2_U2742 , P2_R2099_U120 );
not NOT1_24601 ( P2_R2099_U18 , P2_U2741 );
nand NAND2_24602 ( P2_R2099_U19 , P2_U2741 , P2_R2099_U121 );
not NOT1_24603 ( P2_R2099_U20 , P2_U2740 );
nand NAND2_24604 ( P2_R2099_U21 , P2_U2740 , P2_R2099_U122 );
not NOT1_24605 ( P2_R2099_U22 , P2_U2739 );
not NOT1_24606 ( P2_R2099_U23 , P2_U2738 );
nand NAND2_24607 ( P2_R2099_U24 , P2_U2739 , P2_R2099_U123 );
nand NAND2_24608 ( P2_R2099_U25 , P2_R2099_U124 , P2_U2738 );
not NOT1_24609 ( P2_R2099_U26 , P2_U2737 );
nand NAND2_24610 ( P2_R2099_U27 , P2_U2737 , P2_R2099_U125 );
not NOT1_24611 ( P2_R2099_U28 , P2_U2736 );
nand NAND2_24612 ( P2_R2099_U29 , P2_U2736 , P2_R2099_U126 );
not NOT1_24613 ( P2_R2099_U30 , P2_U2735 );
nand NAND2_24614 ( P2_R2099_U31 , P2_U2735 , P2_R2099_U127 );
not NOT1_24615 ( P2_R2099_U32 , P2_U2734 );
nand NAND2_24616 ( P2_R2099_U33 , P2_U2734 , P2_R2099_U128 );
not NOT1_24617 ( P2_R2099_U34 , P2_U2733 );
nand NAND2_24618 ( P2_R2099_U35 , P2_U2733 , P2_R2099_U129 );
not NOT1_24619 ( P2_R2099_U36 , P2_U2732 );
nand NAND2_24620 ( P2_R2099_U37 , P2_U2732 , P2_R2099_U130 );
not NOT1_24621 ( P2_R2099_U38 , P2_U2731 );
nand NAND2_24622 ( P2_R2099_U39 , P2_U2731 , P2_R2099_U131 );
not NOT1_24623 ( P2_R2099_U40 , P2_U2730 );
nand NAND2_24624 ( P2_R2099_U41 , P2_U2730 , P2_R2099_U132 );
not NOT1_24625 ( P2_R2099_U42 , P2_U2729 );
nand NAND2_24626 ( P2_R2099_U43 , P2_U2729 , P2_R2099_U133 );
not NOT1_24627 ( P2_R2099_U44 , P2_U2728 );
nand NAND2_24628 ( P2_R2099_U45 , P2_U2728 , P2_R2099_U134 );
not NOT1_24629 ( P2_R2099_U46 , P2_U2727 );
nand NAND2_24630 ( P2_R2099_U47 , P2_U2727 , P2_R2099_U135 );
not NOT1_24631 ( P2_R2099_U48 , P2_U2726 );
nand NAND2_24632 ( P2_R2099_U49 , P2_U2726 , P2_R2099_U136 );
not NOT1_24633 ( P2_R2099_U50 , P2_U2725 );
nand NAND2_24634 ( P2_R2099_U51 , P2_U2725 , P2_R2099_U137 );
not NOT1_24635 ( P2_R2099_U52 , P2_U2724 );
nand NAND2_24636 ( P2_R2099_U53 , P2_U2724 , P2_R2099_U138 );
not NOT1_24637 ( P2_R2099_U54 , P2_U2723 );
nand NAND2_24638 ( P2_R2099_U55 , P2_U2723 , P2_R2099_U139 );
not NOT1_24639 ( P2_R2099_U56 , P2_U2722 );
nand NAND2_24640 ( P2_R2099_U57 , P2_U2722 , P2_R2099_U140 );
not NOT1_24641 ( P2_R2099_U58 , P2_U2721 );
nand NAND2_24642 ( P2_R2099_U59 , P2_U2721 , P2_R2099_U141 );
not NOT1_24643 ( P2_R2099_U60 , P2_U2720 );
nand NAND2_24644 ( P2_R2099_U61 , P2_U2720 , P2_R2099_U142 );
not NOT1_24645 ( P2_R2099_U62 , P2_U2719 );
nand NAND2_24646 ( P2_R2099_U63 , P2_U2719 , P2_R2099_U143 );
not NOT1_24647 ( P2_R2099_U64 , P2_U2718 );
nand NAND2_24648 ( P2_R2099_U65 , P2_U2718 , P2_R2099_U144 );
not NOT1_24649 ( P2_R2099_U66 , P2_U2717 );
nand NAND2_24650 ( P2_R2099_U67 , P2_R2099_U150 , P2_R2099_U149 );
nand NAND2_24651 ( P2_R2099_U68 , P2_R2099_U152 , P2_R2099_U151 );
nand NAND2_24652 ( P2_R2099_U69 , P2_R2099_U154 , P2_R2099_U153 );
nand NAND2_24653 ( P2_R2099_U70 , P2_R2099_U156 , P2_R2099_U155 );
nand NAND2_24654 ( P2_R2099_U71 , P2_R2099_U158 , P2_R2099_U157 );
nand NAND2_24655 ( P2_R2099_U72 , P2_R2099_U169 , P2_R2099_U168 );
nand NAND2_24656 ( P2_R2099_U73 , P2_R2099_U171 , P2_R2099_U170 );
nand NAND2_24657 ( P2_R2099_U74 , P2_R2099_U180 , P2_R2099_U179 );
nand NAND2_24658 ( P2_R2099_U75 , P2_R2099_U182 , P2_R2099_U181 );
nand NAND2_24659 ( P2_R2099_U76 , P2_R2099_U184 , P2_R2099_U183 );
nand NAND2_24660 ( P2_R2099_U77 , P2_R2099_U186 , P2_R2099_U185 );
nand NAND2_24661 ( P2_R2099_U78 , P2_R2099_U188 , P2_R2099_U187 );
nand NAND2_24662 ( P2_R2099_U79 , P2_R2099_U190 , P2_R2099_U189 );
nand NAND2_24663 ( P2_R2099_U80 , P2_R2099_U192 , P2_R2099_U191 );
nand NAND2_24664 ( P2_R2099_U81 , P2_R2099_U194 , P2_R2099_U193 );
nand NAND2_24665 ( P2_R2099_U82 , P2_R2099_U196 , P2_R2099_U195 );
nand NAND2_24666 ( P2_R2099_U83 , P2_R2099_U198 , P2_R2099_U197 );
nand NAND2_24667 ( P2_R2099_U84 , P2_R2099_U205 , P2_R2099_U204 );
nand NAND2_24668 ( P2_R2099_U85 , P2_R2099_U207 , P2_R2099_U206 );
nand NAND2_24669 ( P2_R2099_U86 , P2_R2099_U209 , P2_R2099_U208 );
nand NAND2_24670 ( P2_R2099_U87 , P2_R2099_U211 , P2_R2099_U210 );
nand NAND2_24671 ( P2_R2099_U88 , P2_R2099_U213 , P2_R2099_U212 );
nand NAND2_24672 ( P2_R2099_U89 , P2_R2099_U215 , P2_R2099_U214 );
nand NAND2_24673 ( P2_R2099_U90 , P2_R2099_U217 , P2_R2099_U216 );
nand NAND2_24674 ( P2_R2099_U91 , P2_R2099_U219 , P2_R2099_U218 );
nand NAND2_24675 ( P2_R2099_U92 , P2_R2099_U221 , P2_R2099_U220 );
nand NAND2_24676 ( P2_R2099_U93 , P2_R2099_U223 , P2_R2099_U222 );
nand NAND2_24677 ( P2_R2099_U94 , P2_R2099_U225 , P2_R2099_U224 );
nand NAND2_24678 ( P2_R2099_U95 , P2_R2099_U167 , P2_R2099_U166 );
nand NAND2_24679 ( P2_R2099_U96 , P2_R2099_U178 , P2_R2099_U177 );
nand NAND2_24680 ( P2_R2099_U97 , P2_R2099_U118 , P2_R2099_U117 );
and AND2_24681 ( P2_R2099_U98 , P2_R2099_U160 , P2_R2099_U159 );
and AND2_24682 ( P2_R2099_U99 , P2_R2099_U162 , P2_R2099_U161 );
nand NAND2_24683 ( P2_R2099_U100 , P2_R2099_U114 , P2_R2099_U113 );
not NOT1_24684 ( P2_R2099_U101 , P2_U2716 );
nand NAND2_24685 ( P2_R2099_U102 , P2_U2717 , P2_R2099_U145 );
and AND2_24686 ( P2_R2099_U103 , P2_R2099_U173 , P2_R2099_U172 );
nand NAND2_24687 ( P2_R2099_U104 , P2_R2099_U106 , P2_R2099_U110 );
nand NAND2_24688 ( P2_R2099_U105 , P2_U2751 , P2_U2747 );
nand NAND3_24689 ( P2_R2099_U106 , P2_U2746 , P2_U2747 , P2_U2751 );
and AND2_24690 ( P2_R2099_U107 , P2_R2099_U203 , P2_R2099_U202 );
not NOT1_24691 ( P2_R2099_U108 , P2_R2099_U106 );
nand NAND2_24692 ( P2_R2099_U109 , P2_R2099_U9 , P2_R2099_U105 );
nand NAND2_24693 ( P2_R2099_U110 , P2_U2750 , P2_R2099_U109 );
not NOT1_24694 ( P2_R2099_U111 , P2_R2099_U104 );
or OR2_24695 ( P2_R2099_U112 , P2_U2749 , P2_U2745 );
nand NAND2_24696 ( P2_R2099_U113 , P2_R2099_U112 , P2_R2099_U104 );
nand NAND2_24697 ( P2_R2099_U114 , P2_U2745 , P2_U2749 );
not NOT1_24698 ( P2_R2099_U115 , P2_R2099_U100 );
or OR2_24699 ( P2_R2099_U116 , P2_U2748 , P2_U2744 );
nand NAND2_24700 ( P2_R2099_U117 , P2_R2099_U116 , P2_R2099_U100 );
nand NAND2_24701 ( P2_R2099_U118 , P2_U2744 , P2_U2748 );
not NOT1_24702 ( P2_R2099_U119 , P2_R2099_U97 );
not NOT1_24703 ( P2_R2099_U120 , P2_R2099_U15 );
not NOT1_24704 ( P2_R2099_U121 , P2_R2099_U17 );
not NOT1_24705 ( P2_R2099_U122 , P2_R2099_U19 );
not NOT1_24706 ( P2_R2099_U123 , P2_R2099_U21 );
not NOT1_24707 ( P2_R2099_U124 , P2_R2099_U24 );
not NOT1_24708 ( P2_R2099_U125 , P2_R2099_U25 );
not NOT1_24709 ( P2_R2099_U126 , P2_R2099_U27 );
not NOT1_24710 ( P2_R2099_U127 , P2_R2099_U29 );
not NOT1_24711 ( P2_R2099_U128 , P2_R2099_U31 );
not NOT1_24712 ( P2_R2099_U129 , P2_R2099_U33 );
not NOT1_24713 ( P2_R2099_U130 , P2_R2099_U35 );
not NOT1_24714 ( P2_R2099_U131 , P2_R2099_U37 );
not NOT1_24715 ( P2_R2099_U132 , P2_R2099_U39 );
not NOT1_24716 ( P2_R2099_U133 , P2_R2099_U41 );
not NOT1_24717 ( P2_R2099_U134 , P2_R2099_U43 );
not NOT1_24718 ( P2_R2099_U135 , P2_R2099_U45 );
not NOT1_24719 ( P2_R2099_U136 , P2_R2099_U47 );
not NOT1_24720 ( P2_R2099_U137 , P2_R2099_U49 );
not NOT1_24721 ( P2_R2099_U138 , P2_R2099_U51 );
not NOT1_24722 ( P2_R2099_U139 , P2_R2099_U53 );
not NOT1_24723 ( P2_R2099_U140 , P2_R2099_U55 );
not NOT1_24724 ( P2_R2099_U141 , P2_R2099_U57 );
not NOT1_24725 ( P2_R2099_U142 , P2_R2099_U59 );
not NOT1_24726 ( P2_R2099_U143 , P2_R2099_U61 );
not NOT1_24727 ( P2_R2099_U144 , P2_R2099_U63 );
not NOT1_24728 ( P2_R2099_U145 , P2_R2099_U65 );
not NOT1_24729 ( P2_R2099_U146 , P2_R2099_U102 );
not NOT1_24730 ( P2_R2099_U147 , P2_R2099_U105 );
nand NAND2_24731 ( P2_R2099_U148 , P2_R2099_U201 , P2_R2099_U9 );
nand NAND2_24732 ( P2_R2099_U149 , P2_U2738 , P2_R2099_U24 );
nand NAND2_24733 ( P2_R2099_U150 , P2_R2099_U124 , P2_R2099_U23 );
nand NAND2_24734 ( P2_R2099_U151 , P2_U2739 , P2_R2099_U21 );
nand NAND2_24735 ( P2_R2099_U152 , P2_R2099_U123 , P2_R2099_U22 );
nand NAND2_24736 ( P2_R2099_U153 , P2_U2740 , P2_R2099_U19 );
nand NAND2_24737 ( P2_R2099_U154 , P2_R2099_U122 , P2_R2099_U20 );
nand NAND2_24738 ( P2_R2099_U155 , P2_U2741 , P2_R2099_U17 );
nand NAND2_24739 ( P2_R2099_U156 , P2_R2099_U121 , P2_R2099_U18 );
nand NAND2_24740 ( P2_R2099_U157 , P2_U2742 , P2_R2099_U15 );
nand NAND2_24741 ( P2_R2099_U158 , P2_R2099_U120 , P2_R2099_U16 );
nand NAND2_24742 ( P2_R2099_U159 , P2_U2743 , P2_R2099_U97 );
nand NAND2_24743 ( P2_R2099_U160 , P2_R2099_U119 , P2_R2099_U14 );
nand NAND2_24744 ( P2_R2099_U161 , P2_U2744 , P2_R2099_U12 );
nand NAND2_24745 ( P2_R2099_U162 , P2_U2748 , P2_R2099_U13 );
nand NAND2_24746 ( P2_R2099_U163 , P2_U2744 , P2_R2099_U12 );
nand NAND2_24747 ( P2_R2099_U164 , P2_U2748 , P2_R2099_U13 );
nand NAND2_24748 ( P2_R2099_U165 , P2_R2099_U164 , P2_R2099_U163 );
nand NAND2_24749 ( P2_R2099_U166 , P2_R2099_U99 , P2_R2099_U100 );
nand NAND2_24750 ( P2_R2099_U167 , P2_R2099_U115 , P2_R2099_U165 );
nand NAND2_24751 ( P2_R2099_U168 , P2_U2716 , P2_R2099_U102 );
nand NAND2_24752 ( P2_R2099_U169 , P2_R2099_U146 , P2_R2099_U101 );
nand NAND2_24753 ( P2_R2099_U170 , P2_U2717 , P2_R2099_U65 );
nand NAND2_24754 ( P2_R2099_U171 , P2_R2099_U145 , P2_R2099_U66 );
nand NAND2_24755 ( P2_R2099_U172 , P2_U2745 , P2_R2099_U10 );
nand NAND2_24756 ( P2_R2099_U173 , P2_U2749 , P2_R2099_U11 );
nand NAND2_24757 ( P2_R2099_U174 , P2_U2745 , P2_R2099_U10 );
nand NAND2_24758 ( P2_R2099_U175 , P2_U2749 , P2_R2099_U11 );
nand NAND2_24759 ( P2_R2099_U176 , P2_R2099_U175 , P2_R2099_U174 );
nand NAND2_24760 ( P2_R2099_U177 , P2_R2099_U103 , P2_R2099_U104 );
nand NAND2_24761 ( P2_R2099_U178 , P2_R2099_U111 , P2_R2099_U176 );
nand NAND2_24762 ( P2_R2099_U179 , P2_U2718 , P2_R2099_U63 );
nand NAND2_24763 ( P2_R2099_U180 , P2_R2099_U144 , P2_R2099_U64 );
nand NAND2_24764 ( P2_R2099_U181 , P2_U2719 , P2_R2099_U61 );
nand NAND2_24765 ( P2_R2099_U182 , P2_R2099_U143 , P2_R2099_U62 );
nand NAND2_24766 ( P2_R2099_U183 , P2_U2720 , P2_R2099_U59 );
nand NAND2_24767 ( P2_R2099_U184 , P2_R2099_U142 , P2_R2099_U60 );
nand NAND2_24768 ( P2_R2099_U185 , P2_U2721 , P2_R2099_U57 );
nand NAND2_24769 ( P2_R2099_U186 , P2_R2099_U141 , P2_R2099_U58 );
nand NAND2_24770 ( P2_R2099_U187 , P2_U2722 , P2_R2099_U55 );
nand NAND2_24771 ( P2_R2099_U188 , P2_R2099_U140 , P2_R2099_U56 );
nand NAND2_24772 ( P2_R2099_U189 , P2_U2723 , P2_R2099_U53 );
nand NAND2_24773 ( P2_R2099_U190 , P2_R2099_U139 , P2_R2099_U54 );
nand NAND2_24774 ( P2_R2099_U191 , P2_U2724 , P2_R2099_U51 );
nand NAND2_24775 ( P2_R2099_U192 , P2_R2099_U138 , P2_R2099_U52 );
nand NAND2_24776 ( P2_R2099_U193 , P2_U2725 , P2_R2099_U49 );
nand NAND2_24777 ( P2_R2099_U194 , P2_R2099_U137 , P2_R2099_U50 );
nand NAND2_24778 ( P2_R2099_U195 , P2_U2726 , P2_R2099_U47 );
nand NAND2_24779 ( P2_R2099_U196 , P2_R2099_U136 , P2_R2099_U48 );
nand NAND2_24780 ( P2_R2099_U197 , P2_U2727 , P2_R2099_U45 );
nand NAND2_24781 ( P2_R2099_U198 , P2_R2099_U135 , P2_R2099_U46 );
nand NAND2_24782 ( P2_R2099_U199 , P2_U2750 , P2_R2099_U105 );
nand NAND2_24783 ( P2_R2099_U200 , P2_R2099_U147 , P2_R2099_U8 );
nand NAND2_24784 ( P2_R2099_U201 , P2_R2099_U200 , P2_R2099_U199 );
nand NAND3_24785 ( P2_R2099_U202 , P2_U2746 , P2_R2099_U105 , P2_R2099_U8 );
nand NAND2_24786 ( P2_R2099_U203 , P2_R2099_U108 , P2_U2750 );
nand NAND2_24787 ( P2_R2099_U204 , P2_U2728 , P2_R2099_U43 );
nand NAND2_24788 ( P2_R2099_U205 , P2_R2099_U134 , P2_R2099_U44 );
nand NAND2_24789 ( P2_R2099_U206 , P2_U2729 , P2_R2099_U41 );
nand NAND2_24790 ( P2_R2099_U207 , P2_R2099_U133 , P2_R2099_U42 );
nand NAND2_24791 ( P2_R2099_U208 , P2_U2730 , P2_R2099_U39 );
nand NAND2_24792 ( P2_R2099_U209 , P2_R2099_U132 , P2_R2099_U40 );
nand NAND2_24793 ( P2_R2099_U210 , P2_U2731 , P2_R2099_U37 );
nand NAND2_24794 ( P2_R2099_U211 , P2_R2099_U131 , P2_R2099_U38 );
nand NAND2_24795 ( P2_R2099_U212 , P2_U2732 , P2_R2099_U35 );
nand NAND2_24796 ( P2_R2099_U213 , P2_R2099_U130 , P2_R2099_U36 );
nand NAND2_24797 ( P2_R2099_U214 , P2_U2733 , P2_R2099_U33 );
nand NAND2_24798 ( P2_R2099_U215 , P2_R2099_U129 , P2_R2099_U34 );
nand NAND2_24799 ( P2_R2099_U216 , P2_U2734 , P2_R2099_U31 );
nand NAND2_24800 ( P2_R2099_U217 , P2_R2099_U128 , P2_R2099_U32 );
nand NAND2_24801 ( P2_R2099_U218 , P2_U2735 , P2_R2099_U29 );
nand NAND2_24802 ( P2_R2099_U219 , P2_R2099_U127 , P2_R2099_U30 );
nand NAND2_24803 ( P2_R2099_U220 , P2_U2736 , P2_R2099_U27 );
nand NAND2_24804 ( P2_R2099_U221 , P2_R2099_U126 , P2_R2099_U28 );
nand NAND2_24805 ( P2_R2099_U222 , P2_U2737 , P2_R2099_U25 );
nand NAND2_24806 ( P2_R2099_U223 , P2_R2099_U125 , P2_R2099_U26 );
nand NAND2_24807 ( P2_R2099_U224 , P2_U2751 , P2_R2099_U6 );
nand NAND2_24808 ( P2_R2099_U225 , P2_U2747 , P2_R2099_U7 );
and AND2_24809 ( P2_ADD_391_1196_U5 , P2_ADD_391_1196_U301 , P2_ADD_391_1196_U299 );
and AND2_24810 ( P2_ADD_391_1196_U6 , P2_ADD_391_1196_U296 , P2_ADD_391_1196_U294 );
and AND2_24811 ( P2_ADD_391_1196_U7 , P2_ADD_391_1196_U292 , P2_ADD_391_1196_U290 );
and AND2_24812 ( P2_ADD_391_1196_U8 , P2_ADD_391_1196_U287 , P2_ADD_391_1196_U283 );
and AND2_24813 ( P2_ADD_391_1196_U9 , P2_ADD_391_1196_U205 , P2_ADD_391_1196_U203 );
and AND2_24814 ( P2_ADD_391_1196_U10 , P2_ADD_391_1196_U201 , P2_ADD_391_1196_U199 );
and AND2_24815 ( P2_ADD_391_1196_U11 , P2_ADD_391_1196_U196 , P2_ADD_391_1196_U192 );
nand NAND2_24816 ( P2_ADD_391_1196_U12 , P2_ADD_391_1196_U144 , P2_ADD_391_1196_U306 );
not NOT1_24817 ( P2_ADD_391_1196_U13 , P2_R2182_U72 );
not NOT1_24818 ( P2_ADD_391_1196_U14 , P2_R2096_U71 );
not NOT1_24819 ( P2_ADD_391_1196_U15 , P2_R2182_U73 );
not NOT1_24820 ( P2_ADD_391_1196_U16 , P2_R2096_U72 );
not NOT1_24821 ( P2_ADD_391_1196_U17 , P2_R2182_U74 );
not NOT1_24822 ( P2_ADD_391_1196_U18 , P2_R2096_U73 );
not NOT1_24823 ( P2_ADD_391_1196_U19 , P2_R2096_U68 );
not NOT1_24824 ( P2_ADD_391_1196_U20 , P2_R2182_U69 );
not NOT1_24825 ( P2_ADD_391_1196_U21 , P2_R2182_U68 );
nand NAND2_24826 ( P2_ADD_391_1196_U22 , P2_R2182_U69 , P2_R2096_U68 );
not NOT1_24827 ( P2_ADD_391_1196_U23 , P2_R2096_U51 );
not NOT1_24828 ( P2_ADD_391_1196_U24 , P2_R2182_U40 );
not NOT1_24829 ( P2_ADD_391_1196_U25 , P2_R2096_U77 );
not NOT1_24830 ( P2_ADD_391_1196_U26 , P2_R2182_U76 );
not NOT1_24831 ( P2_ADD_391_1196_U27 , P2_R2096_U75 );
not NOT1_24832 ( P2_ADD_391_1196_U28 , P2_R2182_U75 );
not NOT1_24833 ( P2_ADD_391_1196_U29 , P2_R2096_U74 );
nand NAND2_24834 ( P2_ADD_391_1196_U30 , P2_ADD_391_1196_U39 , P2_ADD_391_1196_U180 );
not NOT1_24835 ( P2_ADD_391_1196_U31 , P2_R2182_U71 );
not NOT1_24836 ( P2_ADD_391_1196_U32 , P2_R2096_U70 );
not NOT1_24837 ( P2_ADD_391_1196_U33 , P2_R2096_U69 );
not NOT1_24838 ( P2_ADD_391_1196_U34 , P2_R2182_U70 );
nand NAND2_24839 ( P2_ADD_391_1196_U35 , P2_ADD_391_1196_U190 , P2_ADD_391_1196_U189 );
nand NAND2_24840 ( P2_ADD_391_1196_U36 , P2_ADD_391_1196_U35 , P2_ADD_391_1196_U193 );
nand NAND3_24841 ( P2_ADD_391_1196_U37 , P2_ADD_391_1196_U184 , P2_ADD_391_1196_U182 , P2_ADD_391_1196_U183 );
nand NAND2_24842 ( P2_ADD_391_1196_U38 , P2_ADD_391_1196_U176 , P2_ADD_391_1196_U175 );
nand NAND2_24843 ( P2_ADD_391_1196_U39 , P2_ADD_391_1196_U38 , P2_ADD_391_1196_U178 );
not NOT1_24844 ( P2_ADD_391_1196_U40 , P2_R2182_U91 );
not NOT1_24845 ( P2_ADD_391_1196_U41 , P2_R2096_U92 );
not NOT1_24846 ( P2_ADD_391_1196_U42 , P2_R2182_U92 );
not NOT1_24847 ( P2_ADD_391_1196_U43 , P2_R2096_U93 );
not NOT1_24848 ( P2_ADD_391_1196_U44 , P2_R2182_U93 );
not NOT1_24849 ( P2_ADD_391_1196_U45 , P2_R2096_U94 );
not NOT1_24850 ( P2_ADD_391_1196_U46 , P2_R2182_U95 );
not NOT1_24851 ( P2_ADD_391_1196_U47 , P2_R2096_U96 );
not NOT1_24852 ( P2_ADD_391_1196_U48 , P2_R2182_U96 );
not NOT1_24853 ( P2_ADD_391_1196_U49 , P2_R2096_U97 );
nand NAND2_24854 ( P2_ADD_391_1196_U50 , P2_ADD_391_1196_U36 , P2_ADD_391_1196_U206 );
not NOT1_24855 ( P2_ADD_391_1196_U51 , P2_R2182_U94 );
not NOT1_24856 ( P2_ADD_391_1196_U52 , P2_R2096_U95 );
nand NAND2_24857 ( P2_ADD_391_1196_U53 , P2_ADD_391_1196_U85 , P2_ADD_391_1196_U220 );
not NOT1_24858 ( P2_ADD_391_1196_U54 , P2_R2182_U90 );
not NOT1_24859 ( P2_ADD_391_1196_U55 , P2_R2096_U91 );
not NOT1_24860 ( P2_ADD_391_1196_U56 , P2_R2182_U89 );
not NOT1_24861 ( P2_ADD_391_1196_U57 , P2_R2096_U90 );
not NOT1_24862 ( P2_ADD_391_1196_U58 , P2_R2182_U88 );
not NOT1_24863 ( P2_ADD_391_1196_U59 , P2_R2096_U89 );
not NOT1_24864 ( P2_ADD_391_1196_U60 , P2_R2182_U87 );
not NOT1_24865 ( P2_ADD_391_1196_U61 , P2_R2096_U88 );
not NOT1_24866 ( P2_ADD_391_1196_U62 , P2_R2182_U86 );
not NOT1_24867 ( P2_ADD_391_1196_U63 , P2_R2096_U87 );
not NOT1_24868 ( P2_ADD_391_1196_U64 , P2_R2182_U85 );
not NOT1_24869 ( P2_ADD_391_1196_U65 , P2_R2096_U86 );
not NOT1_24870 ( P2_ADD_391_1196_U66 , P2_R2182_U84 );
not NOT1_24871 ( P2_ADD_391_1196_U67 , P2_R2096_U85 );
not NOT1_24872 ( P2_ADD_391_1196_U68 , P2_R2182_U83 );
not NOT1_24873 ( P2_ADD_391_1196_U69 , P2_R2096_U84 );
not NOT1_24874 ( P2_ADD_391_1196_U70 , P2_R2182_U82 );
not NOT1_24875 ( P2_ADD_391_1196_U71 , P2_R2096_U83 );
not NOT1_24876 ( P2_ADD_391_1196_U72 , P2_R2182_U81 );
not NOT1_24877 ( P2_ADD_391_1196_U73 , P2_R2096_U82 );
not NOT1_24878 ( P2_ADD_391_1196_U74 , P2_R2182_U80 );
not NOT1_24879 ( P2_ADD_391_1196_U75 , P2_R2096_U81 );
not NOT1_24880 ( P2_ADD_391_1196_U76 , P2_R2182_U79 );
not NOT1_24881 ( P2_ADD_391_1196_U77 , P2_R2096_U80 );
not NOT1_24882 ( P2_ADD_391_1196_U78 , P2_R2096_U79 );
not NOT1_24883 ( P2_ADD_391_1196_U79 , P2_R2182_U78 );
not NOT1_24884 ( P2_ADD_391_1196_U80 , P2_R2096_U78 );
not NOT1_24885 ( P2_ADD_391_1196_U81 , P2_R2182_U77 );
nand NAND2_24886 ( P2_ADD_391_1196_U82 , P2_ADD_391_1196_U278 , P2_ADD_391_1196_U277 );
nand NAND3_24887 ( P2_ADD_391_1196_U83 , P2_ADD_391_1196_U224 , P2_ADD_391_1196_U222 , P2_ADD_391_1196_U223 );
nand NAND2_24888 ( P2_ADD_391_1196_U84 , P2_ADD_391_1196_U216 , P2_ADD_391_1196_U215 );
nand NAND2_24889 ( P2_ADD_391_1196_U85 , P2_ADD_391_1196_U84 , P2_ADD_391_1196_U218 );
nand NAND3_24890 ( P2_ADD_391_1196_U86 , P2_ADD_391_1196_U210 , P2_ADD_391_1196_U208 , P2_ADD_391_1196_U209 );
nand NAND2_24891 ( P2_ADD_391_1196_U87 , P2_ADD_391_1196_U478 , P2_ADD_391_1196_U477 );
nand NAND2_24892 ( P2_ADD_391_1196_U88 , P2_ADD_391_1196_U315 , P2_ADD_391_1196_U314 );
nand NAND2_24893 ( P2_ADD_391_1196_U89 , P2_ADD_391_1196_U322 , P2_ADD_391_1196_U321 );
nand NAND2_24894 ( P2_ADD_391_1196_U90 , P2_ADD_391_1196_U331 , P2_ADD_391_1196_U330 );
nand NAND2_24895 ( P2_ADD_391_1196_U91 , P2_ADD_391_1196_U338 , P2_ADD_391_1196_U337 );
nand NAND2_24896 ( P2_ADD_391_1196_U92 , P2_ADD_391_1196_U350 , P2_ADD_391_1196_U349 );
nand NAND2_24897 ( P2_ADD_391_1196_U93 , P2_ADD_391_1196_U357 , P2_ADD_391_1196_U356 );
nand NAND2_24898 ( P2_ADD_391_1196_U94 , P2_ADD_391_1196_U364 , P2_ADD_391_1196_U363 );
nand NAND2_24899 ( P2_ADD_391_1196_U95 , P2_ADD_391_1196_U371 , P2_ADD_391_1196_U370 );
nand NAND2_24900 ( P2_ADD_391_1196_U96 , P2_ADD_391_1196_U378 , P2_ADD_391_1196_U377 );
nand NAND2_24901 ( P2_ADD_391_1196_U97 , P2_ADD_391_1196_U385 , P2_ADD_391_1196_U384 );
nand NAND2_24902 ( P2_ADD_391_1196_U98 , P2_ADD_391_1196_U392 , P2_ADD_391_1196_U391 );
nand NAND2_24903 ( P2_ADD_391_1196_U99 , P2_ADD_391_1196_U399 , P2_ADD_391_1196_U398 );
nand NAND2_24904 ( P2_ADD_391_1196_U100 , P2_ADD_391_1196_U406 , P2_ADD_391_1196_U405 );
nand NAND2_24905 ( P2_ADD_391_1196_U101 , P2_ADD_391_1196_U413 , P2_ADD_391_1196_U412 );
nand NAND2_24906 ( P2_ADD_391_1196_U102 , P2_ADD_391_1196_U420 , P2_ADD_391_1196_U419 );
nand NAND2_24907 ( P2_ADD_391_1196_U103 , P2_ADD_391_1196_U432 , P2_ADD_391_1196_U431 );
nand NAND2_24908 ( P2_ADD_391_1196_U104 , P2_ADD_391_1196_U439 , P2_ADD_391_1196_U438 );
nand NAND2_24909 ( P2_ADD_391_1196_U105 , P2_ADD_391_1196_U446 , P2_ADD_391_1196_U445 );
nand NAND2_24910 ( P2_ADD_391_1196_U106 , P2_ADD_391_1196_U453 , P2_ADD_391_1196_U452 );
nand NAND2_24911 ( P2_ADD_391_1196_U107 , P2_ADD_391_1196_U460 , P2_ADD_391_1196_U459 );
nand NAND2_24912 ( P2_ADD_391_1196_U108 , P2_ADD_391_1196_U469 , P2_ADD_391_1196_U468 );
nand NAND2_24913 ( P2_ADD_391_1196_U109 , P2_ADD_391_1196_U476 , P2_ADD_391_1196_U475 );
and AND2_24914 ( P2_ADD_391_1196_U110 , P2_ADD_391_1196_U308 , P2_ADD_391_1196_U307 );
and AND2_24915 ( P2_ADD_391_1196_U111 , P2_ADD_391_1196_U310 , P2_ADD_391_1196_U309 );
nand NAND2_24916 ( P2_ADD_391_1196_U112 , P2_ADD_391_1196_U37 , P2_ADD_391_1196_U186 );
and AND2_24917 ( P2_ADD_391_1196_U113 , P2_ADD_391_1196_U317 , P2_ADD_391_1196_U316 );
and AND2_24918 ( P2_ADD_391_1196_U114 , P2_ADD_391_1196_U324 , P2_ADD_391_1196_U323 );
and AND2_24919 ( P2_ADD_391_1196_U115 , P2_ADD_391_1196_U326 , P2_ADD_391_1196_U325 );
nand NAND2_24920 ( P2_ADD_391_1196_U116 , P2_ADD_391_1196_U172 , P2_ADD_391_1196_U171 );
and AND2_24921 ( P2_ADD_391_1196_U117 , P2_ADD_391_1196_U333 , P2_ADD_391_1196_U332 );
nand NAND2_24922 ( P2_ADD_391_1196_U118 , P2_ADD_391_1196_U168 , P2_ADD_391_1196_U167 );
not NOT1_24923 ( P2_ADD_391_1196_U119 , P2_R2182_U41 );
not NOT1_24924 ( P2_ADD_391_1196_U120 , P2_R2096_U76 );
and AND2_24925 ( P2_ADD_391_1196_U121 , P2_ADD_391_1196_U340 , P2_ADD_391_1196_U339 );
and AND2_24926 ( P2_ADD_391_1196_U122 , P2_ADD_391_1196_U345 , P2_ADD_391_1196_U344 );
nand NAND2_24927 ( P2_ADD_391_1196_U123 , P2_ADD_391_1196_U143 , P2_ADD_391_1196_U164 );
and AND2_24928 ( P2_ADD_391_1196_U124 , P2_ADD_391_1196_U352 , P2_ADD_391_1196_U351 );
and AND2_24929 ( P2_ADD_391_1196_U125 , P2_ADD_391_1196_U359 , P2_ADD_391_1196_U358 );
nand NAND2_24930 ( P2_ADD_391_1196_U126 , P2_ADD_391_1196_U274 , P2_ADD_391_1196_U273 );
and AND2_24931 ( P2_ADD_391_1196_U127 , P2_ADD_391_1196_U366 , P2_ADD_391_1196_U365 );
nand NAND2_24932 ( P2_ADD_391_1196_U128 , P2_ADD_391_1196_U270 , P2_ADD_391_1196_U269 );
and AND2_24933 ( P2_ADD_391_1196_U129 , P2_ADD_391_1196_U373 , P2_ADD_391_1196_U372 );
nand NAND2_24934 ( P2_ADD_391_1196_U130 , P2_ADD_391_1196_U266 , P2_ADD_391_1196_U265 );
and AND2_24935 ( P2_ADD_391_1196_U131 , P2_ADD_391_1196_U380 , P2_ADD_391_1196_U379 );
nand NAND2_24936 ( P2_ADD_391_1196_U132 , P2_ADD_391_1196_U262 , P2_ADD_391_1196_U261 );
and AND2_24937 ( P2_ADD_391_1196_U133 , P2_ADD_391_1196_U387 , P2_ADD_391_1196_U386 );
nand NAND2_24938 ( P2_ADD_391_1196_U134 , P2_ADD_391_1196_U258 , P2_ADD_391_1196_U257 );
and AND2_24939 ( P2_ADD_391_1196_U135 , P2_ADD_391_1196_U394 , P2_ADD_391_1196_U393 );
nand NAND2_24940 ( P2_ADD_391_1196_U136 , P2_ADD_391_1196_U254 , P2_ADD_391_1196_U253 );
and AND2_24941 ( P2_ADD_391_1196_U137 , P2_ADD_391_1196_U401 , P2_ADD_391_1196_U400 );
nand NAND2_24942 ( P2_ADD_391_1196_U138 , P2_ADD_391_1196_U250 , P2_ADD_391_1196_U249 );
and AND2_24943 ( P2_ADD_391_1196_U139 , P2_ADD_391_1196_U408 , P2_ADD_391_1196_U407 );
nand NAND2_24944 ( P2_ADD_391_1196_U140 , P2_ADD_391_1196_U246 , P2_ADD_391_1196_U245 );
and AND2_24945 ( P2_ADD_391_1196_U141 , P2_ADD_391_1196_U415 , P2_ADD_391_1196_U414 );
nand NAND2_24946 ( P2_ADD_391_1196_U142 , P2_ADD_391_1196_U242 , P2_ADD_391_1196_U241 );
nand NAND2_24947 ( P2_ADD_391_1196_U143 , P2_R2096_U51 , P2_ADD_391_1196_U162 );
and AND2_24948 ( P2_ADD_391_1196_U144 , P2_ADD_391_1196_U425 , P2_ADD_391_1196_U424 );
and AND2_24949 ( P2_ADD_391_1196_U145 , P2_ADD_391_1196_U427 , P2_ADD_391_1196_U426 );
nand NAND2_24950 ( P2_ADD_391_1196_U146 , P2_ADD_391_1196_U238 , P2_ADD_391_1196_U237 );
and AND2_24951 ( P2_ADD_391_1196_U147 , P2_ADD_391_1196_U434 , P2_ADD_391_1196_U433 );
nand NAND2_24952 ( P2_ADD_391_1196_U148 , P2_ADD_391_1196_U234 , P2_ADD_391_1196_U233 );
and AND2_24953 ( P2_ADD_391_1196_U149 , P2_ADD_391_1196_U441 , P2_ADD_391_1196_U440 );
nand NAND2_24954 ( P2_ADD_391_1196_U150 , P2_ADD_391_1196_U230 , P2_ADD_391_1196_U229 );
and AND2_24955 ( P2_ADD_391_1196_U151 , P2_ADD_391_1196_U448 , P2_ADD_391_1196_U447 );
nand NAND2_24956 ( P2_ADD_391_1196_U152 , P2_ADD_391_1196_U83 , P2_ADD_391_1196_U226 );
and AND2_24957 ( P2_ADD_391_1196_U153 , P2_ADD_391_1196_U455 , P2_ADD_391_1196_U454 );
and AND2_24958 ( P2_ADD_391_1196_U154 , P2_ADD_391_1196_U462 , P2_ADD_391_1196_U461 );
and AND2_24959 ( P2_ADD_391_1196_U155 , P2_ADD_391_1196_U464 , P2_ADD_391_1196_U463 );
nand NAND2_24960 ( P2_ADD_391_1196_U156 , P2_ADD_391_1196_U86 , P2_ADD_391_1196_U212 );
and AND2_24961 ( P2_ADD_391_1196_U157 , P2_ADD_391_1196_U471 , P2_ADD_391_1196_U470 );
nand NAND2_24962 ( P2_ADD_391_1196_U158 , P2_R2096_U97 , P2_R2182_U96 );
nand NAND2_24963 ( P2_ADD_391_1196_U159 , P2_R2096_U93 , P2_R2182_U92 );
not NOT1_24964 ( P2_ADD_391_1196_U160 , P2_ADD_391_1196_U143 );
nand NAND2_24965 ( P2_ADD_391_1196_U161 , P2_R2096_U72 , P2_R2182_U73 );
not NOT1_24966 ( P2_ADD_391_1196_U162 , P2_ADD_391_1196_U22 );
nand NAND2_24967 ( P2_ADD_391_1196_U163 , P2_ADD_391_1196_U23 , P2_ADD_391_1196_U22 );
nand NAND2_24968 ( P2_ADD_391_1196_U164 , P2_R2182_U68 , P2_ADD_391_1196_U163 );
not NOT1_24969 ( P2_ADD_391_1196_U165 , P2_ADD_391_1196_U123 );
or OR2_24970 ( P2_ADD_391_1196_U166 , P2_R2182_U40 , P2_R2096_U77 );
nand NAND2_24971 ( P2_ADD_391_1196_U167 , P2_ADD_391_1196_U166 , P2_ADD_391_1196_U123 );
nand NAND2_24972 ( P2_ADD_391_1196_U168 , P2_R2096_U77 , P2_R2182_U40 );
not NOT1_24973 ( P2_ADD_391_1196_U169 , P2_ADD_391_1196_U118 );
or OR2_24974 ( P2_ADD_391_1196_U170 , P2_R2182_U76 , P2_R2096_U75 );
nand NAND2_24975 ( P2_ADD_391_1196_U171 , P2_ADD_391_1196_U170 , P2_ADD_391_1196_U118 );
nand NAND2_24976 ( P2_ADD_391_1196_U172 , P2_R2096_U75 , P2_R2182_U76 );
not NOT1_24977 ( P2_ADD_391_1196_U173 , P2_ADD_391_1196_U116 );
or OR2_24978 ( P2_ADD_391_1196_U174 , P2_R2182_U75 , P2_R2096_U74 );
nand NAND2_24979 ( P2_ADD_391_1196_U175 , P2_ADD_391_1196_U174 , P2_ADD_391_1196_U116 );
nand NAND2_24980 ( P2_ADD_391_1196_U176 , P2_R2096_U74 , P2_R2182_U75 );
not NOT1_24981 ( P2_ADD_391_1196_U177 , P2_ADD_391_1196_U38 );
or OR2_24982 ( P2_ADD_391_1196_U178 , P2_R2096_U73 , P2_R2182_U74 );
not NOT1_24983 ( P2_ADD_391_1196_U179 , P2_ADD_391_1196_U39 );
nand NAND2_24984 ( P2_ADD_391_1196_U180 , P2_R2096_U73 , P2_R2182_U74 );
not NOT1_24985 ( P2_ADD_391_1196_U181 , P2_ADD_391_1196_U30 );
nand NAND2_24986 ( P2_ADD_391_1196_U182 , P2_ADD_391_1196_U181 , P2_ADD_391_1196_U161 );
or OR2_24987 ( P2_ADD_391_1196_U183 , P2_R2096_U71 , P2_R2182_U72 );
or OR2_24988 ( P2_ADD_391_1196_U184 , P2_R2096_U72 , P2_R2182_U73 );
not NOT1_24989 ( P2_ADD_391_1196_U185 , P2_ADD_391_1196_U37 );
nand NAND2_24990 ( P2_ADD_391_1196_U186 , P2_R2096_U71 , P2_R2182_U72 );
not NOT1_24991 ( P2_ADD_391_1196_U187 , P2_ADD_391_1196_U112 );
or OR2_24992 ( P2_ADD_391_1196_U188 , P2_R2182_U71 , P2_R2096_U70 );
nand NAND2_24993 ( P2_ADD_391_1196_U189 , P2_ADD_391_1196_U188 , P2_ADD_391_1196_U112 );
nand NAND2_24994 ( P2_ADD_391_1196_U190 , P2_R2096_U70 , P2_R2182_U71 );
not NOT1_24995 ( P2_ADD_391_1196_U191 , P2_ADD_391_1196_U35 );
nand NAND2_24996 ( P2_ADD_391_1196_U192 , P2_ADD_391_1196_U110 , P2_ADD_391_1196_U191 );
or OR2_24997 ( P2_ADD_391_1196_U193 , P2_R2096_U69 , P2_R2182_U70 );
not NOT1_24998 ( P2_ADD_391_1196_U194 , P2_ADD_391_1196_U36 );
nand NAND2_24999 ( P2_ADD_391_1196_U195 , P2_R2182_U70 , P2_R2096_U69 );
nand NAND2_25000 ( P2_ADD_391_1196_U196 , P2_ADD_391_1196_U194 , P2_ADD_391_1196_U195 );
or OR2_25001 ( P2_ADD_391_1196_U197 , P2_R2182_U73 , P2_R2096_U72 );
nand NAND2_25002 ( P2_ADD_391_1196_U198 , P2_ADD_391_1196_U197 , P2_ADD_391_1196_U30 );
nand NAND3_25003 ( P2_ADD_391_1196_U199 , P2_ADD_391_1196_U198 , P2_ADD_391_1196_U161 , P2_ADD_391_1196_U113 );
nand NAND2_25004 ( P2_ADD_391_1196_U200 , P2_R2096_U71 , P2_R2182_U72 );
nand NAND2_25005 ( P2_ADD_391_1196_U201 , P2_ADD_391_1196_U185 , P2_ADD_391_1196_U200 );
or OR2_25006 ( P2_ADD_391_1196_U202 , P2_R2096_U72 , P2_R2182_U73 );
nand NAND2_25007 ( P2_ADD_391_1196_U203 , P2_ADD_391_1196_U114 , P2_ADD_391_1196_U177 );
nand NAND2_25008 ( P2_ADD_391_1196_U204 , P2_R2096_U73 , P2_R2182_U74 );
nand NAND2_25009 ( P2_ADD_391_1196_U205 , P2_ADD_391_1196_U179 , P2_ADD_391_1196_U204 );
nand NAND2_25010 ( P2_ADD_391_1196_U206 , P2_R2182_U70 , P2_R2096_U69 );
not NOT1_25011 ( P2_ADD_391_1196_U207 , P2_ADD_391_1196_U50 );
nand NAND2_25012 ( P2_ADD_391_1196_U208 , P2_ADD_391_1196_U207 , P2_ADD_391_1196_U158 );
or OR2_25013 ( P2_ADD_391_1196_U209 , P2_R2096_U96 , P2_R2182_U95 );
or OR2_25014 ( P2_ADD_391_1196_U210 , P2_R2096_U97 , P2_R2182_U96 );
not NOT1_25015 ( P2_ADD_391_1196_U211 , P2_ADD_391_1196_U86 );
nand NAND2_25016 ( P2_ADD_391_1196_U212 , P2_R2096_U96 , P2_R2182_U95 );
not NOT1_25017 ( P2_ADD_391_1196_U213 , P2_ADD_391_1196_U156 );
or OR2_25018 ( P2_ADD_391_1196_U214 , P2_R2182_U94 , P2_R2096_U95 );
nand NAND2_25019 ( P2_ADD_391_1196_U215 , P2_ADD_391_1196_U214 , P2_ADD_391_1196_U156 );
nand NAND2_25020 ( P2_ADD_391_1196_U216 , P2_R2096_U95 , P2_R2182_U94 );
not NOT1_25021 ( P2_ADD_391_1196_U217 , P2_ADD_391_1196_U84 );
or OR2_25022 ( P2_ADD_391_1196_U218 , P2_R2096_U94 , P2_R2182_U93 );
not NOT1_25023 ( P2_ADD_391_1196_U219 , P2_ADD_391_1196_U85 );
nand NAND2_25024 ( P2_ADD_391_1196_U220 , P2_R2096_U94 , P2_R2182_U93 );
not NOT1_25025 ( P2_ADD_391_1196_U221 , P2_ADD_391_1196_U53 );
nand NAND2_25026 ( P2_ADD_391_1196_U222 , P2_ADD_391_1196_U221 , P2_ADD_391_1196_U159 );
or OR2_25027 ( P2_ADD_391_1196_U223 , P2_R2096_U92 , P2_R2182_U91 );
or OR2_25028 ( P2_ADD_391_1196_U224 , P2_R2096_U93 , P2_R2182_U92 );
not NOT1_25029 ( P2_ADD_391_1196_U225 , P2_ADD_391_1196_U83 );
nand NAND2_25030 ( P2_ADD_391_1196_U226 , P2_R2096_U92 , P2_R2182_U91 );
not NOT1_25031 ( P2_ADD_391_1196_U227 , P2_ADD_391_1196_U152 );
or OR2_25032 ( P2_ADD_391_1196_U228 , P2_R2182_U90 , P2_R2096_U91 );
nand NAND2_25033 ( P2_ADD_391_1196_U229 , P2_ADD_391_1196_U228 , P2_ADD_391_1196_U152 );
nand NAND2_25034 ( P2_ADD_391_1196_U230 , P2_R2096_U91 , P2_R2182_U90 );
not NOT1_25035 ( P2_ADD_391_1196_U231 , P2_ADD_391_1196_U150 );
or OR2_25036 ( P2_ADD_391_1196_U232 , P2_R2182_U89 , P2_R2096_U90 );
nand NAND2_25037 ( P2_ADD_391_1196_U233 , P2_ADD_391_1196_U232 , P2_ADD_391_1196_U150 );
nand NAND2_25038 ( P2_ADD_391_1196_U234 , P2_R2096_U90 , P2_R2182_U89 );
not NOT1_25039 ( P2_ADD_391_1196_U235 , P2_ADD_391_1196_U148 );
or OR2_25040 ( P2_ADD_391_1196_U236 , P2_R2182_U88 , P2_R2096_U89 );
nand NAND2_25041 ( P2_ADD_391_1196_U237 , P2_ADD_391_1196_U236 , P2_ADD_391_1196_U148 );
nand NAND2_25042 ( P2_ADD_391_1196_U238 , P2_R2096_U89 , P2_R2182_U88 );
not NOT1_25043 ( P2_ADD_391_1196_U239 , P2_ADD_391_1196_U146 );
or OR2_25044 ( P2_ADD_391_1196_U240 , P2_R2182_U87 , P2_R2096_U88 );
nand NAND2_25045 ( P2_ADD_391_1196_U241 , P2_ADD_391_1196_U240 , P2_ADD_391_1196_U146 );
nand NAND2_25046 ( P2_ADD_391_1196_U242 , P2_R2096_U88 , P2_R2182_U87 );
not NOT1_25047 ( P2_ADD_391_1196_U243 , P2_ADD_391_1196_U142 );
or OR2_25048 ( P2_ADD_391_1196_U244 , P2_R2182_U86 , P2_R2096_U87 );
nand NAND2_25049 ( P2_ADD_391_1196_U245 , P2_ADD_391_1196_U244 , P2_ADD_391_1196_U142 );
nand NAND2_25050 ( P2_ADD_391_1196_U246 , P2_R2096_U87 , P2_R2182_U86 );
not NOT1_25051 ( P2_ADD_391_1196_U247 , P2_ADD_391_1196_U140 );
or OR2_25052 ( P2_ADD_391_1196_U248 , P2_R2182_U85 , P2_R2096_U86 );
nand NAND2_25053 ( P2_ADD_391_1196_U249 , P2_ADD_391_1196_U248 , P2_ADD_391_1196_U140 );
nand NAND2_25054 ( P2_ADD_391_1196_U250 , P2_R2096_U86 , P2_R2182_U85 );
not NOT1_25055 ( P2_ADD_391_1196_U251 , P2_ADD_391_1196_U138 );
or OR2_25056 ( P2_ADD_391_1196_U252 , P2_R2182_U84 , P2_R2096_U85 );
nand NAND2_25057 ( P2_ADD_391_1196_U253 , P2_ADD_391_1196_U252 , P2_ADD_391_1196_U138 );
nand NAND2_25058 ( P2_ADD_391_1196_U254 , P2_R2096_U85 , P2_R2182_U84 );
not NOT1_25059 ( P2_ADD_391_1196_U255 , P2_ADD_391_1196_U136 );
or OR2_25060 ( P2_ADD_391_1196_U256 , P2_R2182_U83 , P2_R2096_U84 );
nand NAND2_25061 ( P2_ADD_391_1196_U257 , P2_ADD_391_1196_U256 , P2_ADD_391_1196_U136 );
nand NAND2_25062 ( P2_ADD_391_1196_U258 , P2_R2096_U84 , P2_R2182_U83 );
not NOT1_25063 ( P2_ADD_391_1196_U259 , P2_ADD_391_1196_U134 );
or OR2_25064 ( P2_ADD_391_1196_U260 , P2_R2182_U82 , P2_R2096_U83 );
nand NAND2_25065 ( P2_ADD_391_1196_U261 , P2_ADD_391_1196_U260 , P2_ADD_391_1196_U134 );
nand NAND2_25066 ( P2_ADD_391_1196_U262 , P2_R2096_U83 , P2_R2182_U82 );
not NOT1_25067 ( P2_ADD_391_1196_U263 , P2_ADD_391_1196_U132 );
or OR2_25068 ( P2_ADD_391_1196_U264 , P2_R2182_U81 , P2_R2096_U82 );
nand NAND2_25069 ( P2_ADD_391_1196_U265 , P2_ADD_391_1196_U264 , P2_ADD_391_1196_U132 );
nand NAND2_25070 ( P2_ADD_391_1196_U266 , P2_R2096_U82 , P2_R2182_U81 );
not NOT1_25071 ( P2_ADD_391_1196_U267 , P2_ADD_391_1196_U130 );
or OR2_25072 ( P2_ADD_391_1196_U268 , P2_R2182_U80 , P2_R2096_U81 );
nand NAND2_25073 ( P2_ADD_391_1196_U269 , P2_ADD_391_1196_U268 , P2_ADD_391_1196_U130 );
nand NAND2_25074 ( P2_ADD_391_1196_U270 , P2_R2096_U81 , P2_R2182_U80 );
not NOT1_25075 ( P2_ADD_391_1196_U271 , P2_ADD_391_1196_U128 );
or OR2_25076 ( P2_ADD_391_1196_U272 , P2_R2182_U79 , P2_R2096_U80 );
nand NAND2_25077 ( P2_ADD_391_1196_U273 , P2_ADD_391_1196_U272 , P2_ADD_391_1196_U128 );
nand NAND2_25078 ( P2_ADD_391_1196_U274 , P2_R2096_U80 , P2_R2182_U79 );
not NOT1_25079 ( P2_ADD_391_1196_U275 , P2_ADD_391_1196_U126 );
or OR2_25080 ( P2_ADD_391_1196_U276 , P2_R2096_U79 , P2_R2182_U78 );
nand NAND2_25081 ( P2_ADD_391_1196_U277 , P2_ADD_391_1196_U276 , P2_ADD_391_1196_U126 );
nand NAND2_25082 ( P2_ADD_391_1196_U278 , P2_R2182_U78 , P2_R2096_U79 );
not NOT1_25083 ( P2_ADD_391_1196_U279 , P2_ADD_391_1196_U82 );
or OR2_25084 ( P2_ADD_391_1196_U280 , P2_R2096_U78 , P2_R2182_U77 );
nand NAND2_25085 ( P2_ADD_391_1196_U281 , P2_ADD_391_1196_U280 , P2_ADD_391_1196_U82 );
nand NAND2_25086 ( P2_ADD_391_1196_U282 , P2_R2182_U77 , P2_R2096_U78 );
nand NAND3_25087 ( P2_ADD_391_1196_U283 , P2_ADD_391_1196_U282 , P2_ADD_391_1196_U281 , P2_ADD_391_1196_U121 );
nand NAND2_25088 ( P2_ADD_391_1196_U284 , P2_R2182_U77 , P2_R2096_U78 );
nand NAND2_25089 ( P2_ADD_391_1196_U285 , P2_ADD_391_1196_U279 , P2_ADD_391_1196_U284 );
or OR2_25090 ( P2_ADD_391_1196_U286 , P2_R2182_U77 , P2_R2096_U78 );
nand NAND3_25091 ( P2_ADD_391_1196_U287 , P2_ADD_391_1196_U286 , P2_ADD_391_1196_U285 , P2_ADD_391_1196_U343 );
or OR2_25092 ( P2_ADD_391_1196_U288 , P2_R2182_U92 , P2_R2096_U93 );
nand NAND2_25093 ( P2_ADD_391_1196_U289 , P2_ADD_391_1196_U288 , P2_ADD_391_1196_U53 );
nand NAND3_25094 ( P2_ADD_391_1196_U290 , P2_ADD_391_1196_U289 , P2_ADD_391_1196_U159 , P2_ADD_391_1196_U153 );
nand NAND2_25095 ( P2_ADD_391_1196_U291 , P2_R2096_U92 , P2_R2182_U91 );
nand NAND2_25096 ( P2_ADD_391_1196_U292 , P2_ADD_391_1196_U225 , P2_ADD_391_1196_U291 );
or OR2_25097 ( P2_ADD_391_1196_U293 , P2_R2096_U93 , P2_R2182_U92 );
nand NAND2_25098 ( P2_ADD_391_1196_U294 , P2_ADD_391_1196_U154 , P2_ADD_391_1196_U217 );
nand NAND2_25099 ( P2_ADD_391_1196_U295 , P2_R2096_U94 , P2_R2182_U93 );
nand NAND2_25100 ( P2_ADD_391_1196_U296 , P2_ADD_391_1196_U219 , P2_ADD_391_1196_U295 );
or OR2_25101 ( P2_ADD_391_1196_U297 , P2_R2182_U96 , P2_R2096_U97 );
nand NAND2_25102 ( P2_ADD_391_1196_U298 , P2_ADD_391_1196_U297 , P2_ADD_391_1196_U50 );
nand NAND3_25103 ( P2_ADD_391_1196_U299 , P2_ADD_391_1196_U298 , P2_ADD_391_1196_U158 , P2_ADD_391_1196_U157 );
nand NAND2_25104 ( P2_ADD_391_1196_U300 , P2_R2096_U96 , P2_R2182_U95 );
nand NAND2_25105 ( P2_ADD_391_1196_U301 , P2_ADD_391_1196_U211 , P2_ADD_391_1196_U300 );
or OR2_25106 ( P2_ADD_391_1196_U302 , P2_R2096_U97 , P2_R2182_U96 );
nand NAND2_25107 ( P2_ADD_391_1196_U303 , P2_ADD_391_1196_U202 , P2_ADD_391_1196_U161 );
nand NAND2_25108 ( P2_ADD_391_1196_U304 , P2_ADD_391_1196_U293 , P2_ADD_391_1196_U159 );
nand NAND2_25109 ( P2_ADD_391_1196_U305 , P2_ADD_391_1196_U302 , P2_ADD_391_1196_U158 );
nand NAND2_25110 ( P2_ADD_391_1196_U306 , P2_ADD_391_1196_U423 , P2_ADD_391_1196_U23 );
nand NAND2_25111 ( P2_ADD_391_1196_U307 , P2_R2096_U69 , P2_ADD_391_1196_U34 );
nand NAND2_25112 ( P2_ADD_391_1196_U308 , P2_R2182_U70 , P2_ADD_391_1196_U33 );
nand NAND2_25113 ( P2_ADD_391_1196_U309 , P2_R2096_U70 , P2_ADD_391_1196_U31 );
nand NAND2_25114 ( P2_ADD_391_1196_U310 , P2_R2182_U71 , P2_ADD_391_1196_U32 );
nand NAND2_25115 ( P2_ADD_391_1196_U311 , P2_R2096_U70 , P2_ADD_391_1196_U31 );
nand NAND2_25116 ( P2_ADD_391_1196_U312 , P2_R2182_U71 , P2_ADD_391_1196_U32 );
nand NAND2_25117 ( P2_ADD_391_1196_U313 , P2_ADD_391_1196_U312 , P2_ADD_391_1196_U311 );
nand NAND2_25118 ( P2_ADD_391_1196_U314 , P2_ADD_391_1196_U111 , P2_ADD_391_1196_U112 );
nand NAND2_25119 ( P2_ADD_391_1196_U315 , P2_ADD_391_1196_U187 , P2_ADD_391_1196_U313 );
nand NAND2_25120 ( P2_ADD_391_1196_U316 , P2_R2096_U71 , P2_ADD_391_1196_U13 );
nand NAND2_25121 ( P2_ADD_391_1196_U317 , P2_R2182_U72 , P2_ADD_391_1196_U14 );
nand NAND2_25122 ( P2_ADD_391_1196_U318 , P2_R2096_U72 , P2_ADD_391_1196_U15 );
nand NAND2_25123 ( P2_ADD_391_1196_U319 , P2_R2182_U73 , P2_ADD_391_1196_U16 );
nand NAND2_25124 ( P2_ADD_391_1196_U320 , P2_ADD_391_1196_U319 , P2_ADD_391_1196_U318 );
nand NAND2_25125 ( P2_ADD_391_1196_U321 , P2_ADD_391_1196_U303 , P2_ADD_391_1196_U30 );
nand NAND2_25126 ( P2_ADD_391_1196_U322 , P2_ADD_391_1196_U320 , P2_ADD_391_1196_U181 );
nand NAND2_25127 ( P2_ADD_391_1196_U323 , P2_R2096_U73 , P2_ADD_391_1196_U17 );
nand NAND2_25128 ( P2_ADD_391_1196_U324 , P2_R2182_U74 , P2_ADD_391_1196_U18 );
nand NAND2_25129 ( P2_ADD_391_1196_U325 , P2_R2096_U74 , P2_ADD_391_1196_U28 );
nand NAND2_25130 ( P2_ADD_391_1196_U326 , P2_R2182_U75 , P2_ADD_391_1196_U29 );
nand NAND2_25131 ( P2_ADD_391_1196_U327 , P2_R2096_U74 , P2_ADD_391_1196_U28 );
nand NAND2_25132 ( P2_ADD_391_1196_U328 , P2_R2182_U75 , P2_ADD_391_1196_U29 );
nand NAND2_25133 ( P2_ADD_391_1196_U329 , P2_ADD_391_1196_U328 , P2_ADD_391_1196_U327 );
nand NAND2_25134 ( P2_ADD_391_1196_U330 , P2_ADD_391_1196_U115 , P2_ADD_391_1196_U116 );
nand NAND2_25135 ( P2_ADD_391_1196_U331 , P2_ADD_391_1196_U173 , P2_ADD_391_1196_U329 );
nand NAND2_25136 ( P2_ADD_391_1196_U332 , P2_R2096_U75 , P2_ADD_391_1196_U26 );
nand NAND2_25137 ( P2_ADD_391_1196_U333 , P2_R2182_U76 , P2_ADD_391_1196_U27 );
nand NAND2_25138 ( P2_ADD_391_1196_U334 , P2_R2096_U75 , P2_ADD_391_1196_U26 );
nand NAND2_25139 ( P2_ADD_391_1196_U335 , P2_R2182_U76 , P2_ADD_391_1196_U27 );
nand NAND2_25140 ( P2_ADD_391_1196_U336 , P2_ADD_391_1196_U335 , P2_ADD_391_1196_U334 );
nand NAND2_25141 ( P2_ADD_391_1196_U337 , P2_ADD_391_1196_U117 , P2_ADD_391_1196_U118 );
nand NAND2_25142 ( P2_ADD_391_1196_U338 , P2_ADD_391_1196_U169 , P2_ADD_391_1196_U336 );
nand NAND2_25143 ( P2_ADD_391_1196_U339 , P2_R2182_U41 , P2_ADD_391_1196_U120 );
nand NAND2_25144 ( P2_ADD_391_1196_U340 , P2_R2096_U76 , P2_ADD_391_1196_U119 );
nand NAND2_25145 ( P2_ADD_391_1196_U341 , P2_R2182_U41 , P2_ADD_391_1196_U120 );
nand NAND2_25146 ( P2_ADD_391_1196_U342 , P2_R2096_U76 , P2_ADD_391_1196_U119 );
nand NAND2_25147 ( P2_ADD_391_1196_U343 , P2_ADD_391_1196_U342 , P2_ADD_391_1196_U341 );
nand NAND2_25148 ( P2_ADD_391_1196_U344 , P2_R2096_U77 , P2_ADD_391_1196_U24 );
nand NAND2_25149 ( P2_ADD_391_1196_U345 , P2_R2182_U40 , P2_ADD_391_1196_U25 );
nand NAND2_25150 ( P2_ADD_391_1196_U346 , P2_R2096_U77 , P2_ADD_391_1196_U24 );
nand NAND2_25151 ( P2_ADD_391_1196_U347 , P2_R2182_U40 , P2_ADD_391_1196_U25 );
nand NAND2_25152 ( P2_ADD_391_1196_U348 , P2_ADD_391_1196_U347 , P2_ADD_391_1196_U346 );
nand NAND2_25153 ( P2_ADD_391_1196_U349 , P2_ADD_391_1196_U122 , P2_ADD_391_1196_U123 );
nand NAND2_25154 ( P2_ADD_391_1196_U350 , P2_ADD_391_1196_U165 , P2_ADD_391_1196_U348 );
nand NAND2_25155 ( P2_ADD_391_1196_U351 , P2_R2182_U77 , P2_ADD_391_1196_U80 );
nand NAND2_25156 ( P2_ADD_391_1196_U352 , P2_R2096_U78 , P2_ADD_391_1196_U81 );
nand NAND2_25157 ( P2_ADD_391_1196_U353 , P2_R2182_U77 , P2_ADD_391_1196_U80 );
nand NAND2_25158 ( P2_ADD_391_1196_U354 , P2_R2096_U78 , P2_ADD_391_1196_U81 );
nand NAND2_25159 ( P2_ADD_391_1196_U355 , P2_ADD_391_1196_U354 , P2_ADD_391_1196_U353 );
nand NAND2_25160 ( P2_ADD_391_1196_U356 , P2_ADD_391_1196_U124 , P2_ADD_391_1196_U82 );
nand NAND2_25161 ( P2_ADD_391_1196_U357 , P2_ADD_391_1196_U355 , P2_ADD_391_1196_U279 );
nand NAND2_25162 ( P2_ADD_391_1196_U358 , P2_R2182_U78 , P2_ADD_391_1196_U78 );
nand NAND2_25163 ( P2_ADD_391_1196_U359 , P2_R2096_U79 , P2_ADD_391_1196_U79 );
nand NAND2_25164 ( P2_ADD_391_1196_U360 , P2_R2182_U78 , P2_ADD_391_1196_U78 );
nand NAND2_25165 ( P2_ADD_391_1196_U361 , P2_R2096_U79 , P2_ADD_391_1196_U79 );
nand NAND2_25166 ( P2_ADD_391_1196_U362 , P2_ADD_391_1196_U361 , P2_ADD_391_1196_U360 );
nand NAND2_25167 ( P2_ADD_391_1196_U363 , P2_ADD_391_1196_U125 , P2_ADD_391_1196_U126 );
nand NAND2_25168 ( P2_ADD_391_1196_U364 , P2_ADD_391_1196_U275 , P2_ADD_391_1196_U362 );
nand NAND2_25169 ( P2_ADD_391_1196_U365 , P2_R2096_U80 , P2_ADD_391_1196_U76 );
nand NAND2_25170 ( P2_ADD_391_1196_U366 , P2_R2182_U79 , P2_ADD_391_1196_U77 );
nand NAND2_25171 ( P2_ADD_391_1196_U367 , P2_R2096_U80 , P2_ADD_391_1196_U76 );
nand NAND2_25172 ( P2_ADD_391_1196_U368 , P2_R2182_U79 , P2_ADD_391_1196_U77 );
nand NAND2_25173 ( P2_ADD_391_1196_U369 , P2_ADD_391_1196_U368 , P2_ADD_391_1196_U367 );
nand NAND2_25174 ( P2_ADD_391_1196_U370 , P2_ADD_391_1196_U127 , P2_ADD_391_1196_U128 );
nand NAND2_25175 ( P2_ADD_391_1196_U371 , P2_ADD_391_1196_U271 , P2_ADD_391_1196_U369 );
nand NAND2_25176 ( P2_ADD_391_1196_U372 , P2_R2096_U81 , P2_ADD_391_1196_U74 );
nand NAND2_25177 ( P2_ADD_391_1196_U373 , P2_R2182_U80 , P2_ADD_391_1196_U75 );
nand NAND2_25178 ( P2_ADD_391_1196_U374 , P2_R2096_U81 , P2_ADD_391_1196_U74 );
nand NAND2_25179 ( P2_ADD_391_1196_U375 , P2_R2182_U80 , P2_ADD_391_1196_U75 );
nand NAND2_25180 ( P2_ADD_391_1196_U376 , P2_ADD_391_1196_U375 , P2_ADD_391_1196_U374 );
nand NAND2_25181 ( P2_ADD_391_1196_U377 , P2_ADD_391_1196_U129 , P2_ADD_391_1196_U130 );
nand NAND2_25182 ( P2_ADD_391_1196_U378 , P2_ADD_391_1196_U267 , P2_ADD_391_1196_U376 );
nand NAND2_25183 ( P2_ADD_391_1196_U379 , P2_R2096_U82 , P2_ADD_391_1196_U72 );
nand NAND2_25184 ( P2_ADD_391_1196_U380 , P2_R2182_U81 , P2_ADD_391_1196_U73 );
nand NAND2_25185 ( P2_ADD_391_1196_U381 , P2_R2096_U82 , P2_ADD_391_1196_U72 );
nand NAND2_25186 ( P2_ADD_391_1196_U382 , P2_R2182_U81 , P2_ADD_391_1196_U73 );
nand NAND2_25187 ( P2_ADD_391_1196_U383 , P2_ADD_391_1196_U382 , P2_ADD_391_1196_U381 );
nand NAND2_25188 ( P2_ADD_391_1196_U384 , P2_ADD_391_1196_U131 , P2_ADD_391_1196_U132 );
nand NAND2_25189 ( P2_ADD_391_1196_U385 , P2_ADD_391_1196_U263 , P2_ADD_391_1196_U383 );
nand NAND2_25190 ( P2_ADD_391_1196_U386 , P2_R2096_U83 , P2_ADD_391_1196_U70 );
nand NAND2_25191 ( P2_ADD_391_1196_U387 , P2_R2182_U82 , P2_ADD_391_1196_U71 );
nand NAND2_25192 ( P2_ADD_391_1196_U388 , P2_R2096_U83 , P2_ADD_391_1196_U70 );
nand NAND2_25193 ( P2_ADD_391_1196_U389 , P2_R2182_U82 , P2_ADD_391_1196_U71 );
nand NAND2_25194 ( P2_ADD_391_1196_U390 , P2_ADD_391_1196_U389 , P2_ADD_391_1196_U388 );
nand NAND2_25195 ( P2_ADD_391_1196_U391 , P2_ADD_391_1196_U133 , P2_ADD_391_1196_U134 );
nand NAND2_25196 ( P2_ADD_391_1196_U392 , P2_ADD_391_1196_U259 , P2_ADD_391_1196_U390 );
nand NAND2_25197 ( P2_ADD_391_1196_U393 , P2_R2096_U84 , P2_ADD_391_1196_U68 );
nand NAND2_25198 ( P2_ADD_391_1196_U394 , P2_R2182_U83 , P2_ADD_391_1196_U69 );
nand NAND2_25199 ( P2_ADD_391_1196_U395 , P2_R2096_U84 , P2_ADD_391_1196_U68 );
nand NAND2_25200 ( P2_ADD_391_1196_U396 , P2_R2182_U83 , P2_ADD_391_1196_U69 );
nand NAND2_25201 ( P2_ADD_391_1196_U397 , P2_ADD_391_1196_U396 , P2_ADD_391_1196_U395 );
nand NAND2_25202 ( P2_ADD_391_1196_U398 , P2_ADD_391_1196_U135 , P2_ADD_391_1196_U136 );
nand NAND2_25203 ( P2_ADD_391_1196_U399 , P2_ADD_391_1196_U255 , P2_ADD_391_1196_U397 );
nand NAND2_25204 ( P2_ADD_391_1196_U400 , P2_R2096_U85 , P2_ADD_391_1196_U66 );
nand NAND2_25205 ( P2_ADD_391_1196_U401 , P2_R2182_U84 , P2_ADD_391_1196_U67 );
nand NAND2_25206 ( P2_ADD_391_1196_U402 , P2_R2096_U85 , P2_ADD_391_1196_U66 );
nand NAND2_25207 ( P2_ADD_391_1196_U403 , P2_R2182_U84 , P2_ADD_391_1196_U67 );
nand NAND2_25208 ( P2_ADD_391_1196_U404 , P2_ADD_391_1196_U403 , P2_ADD_391_1196_U402 );
nand NAND2_25209 ( P2_ADD_391_1196_U405 , P2_ADD_391_1196_U137 , P2_ADD_391_1196_U138 );
nand NAND2_25210 ( P2_ADD_391_1196_U406 , P2_ADD_391_1196_U251 , P2_ADD_391_1196_U404 );
nand NAND2_25211 ( P2_ADD_391_1196_U407 , P2_R2096_U86 , P2_ADD_391_1196_U64 );
nand NAND2_25212 ( P2_ADD_391_1196_U408 , P2_R2182_U85 , P2_ADD_391_1196_U65 );
nand NAND2_25213 ( P2_ADD_391_1196_U409 , P2_R2096_U86 , P2_ADD_391_1196_U64 );
nand NAND2_25214 ( P2_ADD_391_1196_U410 , P2_R2182_U85 , P2_ADD_391_1196_U65 );
nand NAND2_25215 ( P2_ADD_391_1196_U411 , P2_ADD_391_1196_U410 , P2_ADD_391_1196_U409 );
nand NAND2_25216 ( P2_ADD_391_1196_U412 , P2_ADD_391_1196_U139 , P2_ADD_391_1196_U140 );
nand NAND2_25217 ( P2_ADD_391_1196_U413 , P2_ADD_391_1196_U247 , P2_ADD_391_1196_U411 );
nand NAND2_25218 ( P2_ADD_391_1196_U414 , P2_R2096_U87 , P2_ADD_391_1196_U62 );
nand NAND2_25219 ( P2_ADD_391_1196_U415 , P2_R2182_U86 , P2_ADD_391_1196_U63 );
nand NAND2_25220 ( P2_ADD_391_1196_U416 , P2_R2096_U87 , P2_ADD_391_1196_U62 );
nand NAND2_25221 ( P2_ADD_391_1196_U417 , P2_R2182_U86 , P2_ADD_391_1196_U63 );
nand NAND2_25222 ( P2_ADD_391_1196_U418 , P2_ADD_391_1196_U417 , P2_ADD_391_1196_U416 );
nand NAND2_25223 ( P2_ADD_391_1196_U419 , P2_ADD_391_1196_U141 , P2_ADD_391_1196_U142 );
nand NAND2_25224 ( P2_ADD_391_1196_U420 , P2_ADD_391_1196_U243 , P2_ADD_391_1196_U418 );
nand NAND2_25225 ( P2_ADD_391_1196_U421 , P2_R2182_U68 , P2_ADD_391_1196_U22 );
nand NAND2_25226 ( P2_ADD_391_1196_U422 , P2_ADD_391_1196_U162 , P2_ADD_391_1196_U21 );
nand NAND2_25227 ( P2_ADD_391_1196_U423 , P2_ADD_391_1196_U422 , P2_ADD_391_1196_U421 );
nand NAND3_25228 ( P2_ADD_391_1196_U424 , P2_R2096_U51 , P2_ADD_391_1196_U22 , P2_ADD_391_1196_U21 );
nand NAND2_25229 ( P2_ADD_391_1196_U425 , P2_ADD_391_1196_U160 , P2_R2182_U68 );
nand NAND2_25230 ( P2_ADD_391_1196_U426 , P2_R2096_U88 , P2_ADD_391_1196_U60 );
nand NAND2_25231 ( P2_ADD_391_1196_U427 , P2_R2182_U87 , P2_ADD_391_1196_U61 );
nand NAND2_25232 ( P2_ADD_391_1196_U428 , P2_R2096_U88 , P2_ADD_391_1196_U60 );
nand NAND2_25233 ( P2_ADD_391_1196_U429 , P2_R2182_U87 , P2_ADD_391_1196_U61 );
nand NAND2_25234 ( P2_ADD_391_1196_U430 , P2_ADD_391_1196_U429 , P2_ADD_391_1196_U428 );
nand NAND2_25235 ( P2_ADD_391_1196_U431 , P2_ADD_391_1196_U145 , P2_ADD_391_1196_U146 );
nand NAND2_25236 ( P2_ADD_391_1196_U432 , P2_ADD_391_1196_U239 , P2_ADD_391_1196_U430 );
nand NAND2_25237 ( P2_ADD_391_1196_U433 , P2_R2096_U89 , P2_ADD_391_1196_U58 );
nand NAND2_25238 ( P2_ADD_391_1196_U434 , P2_R2182_U88 , P2_ADD_391_1196_U59 );
nand NAND2_25239 ( P2_ADD_391_1196_U435 , P2_R2096_U89 , P2_ADD_391_1196_U58 );
nand NAND2_25240 ( P2_ADD_391_1196_U436 , P2_R2182_U88 , P2_ADD_391_1196_U59 );
nand NAND2_25241 ( P2_ADD_391_1196_U437 , P2_ADD_391_1196_U436 , P2_ADD_391_1196_U435 );
nand NAND2_25242 ( P2_ADD_391_1196_U438 , P2_ADD_391_1196_U147 , P2_ADD_391_1196_U148 );
nand NAND2_25243 ( P2_ADD_391_1196_U439 , P2_ADD_391_1196_U235 , P2_ADD_391_1196_U437 );
nand NAND2_25244 ( P2_ADD_391_1196_U440 , P2_R2096_U90 , P2_ADD_391_1196_U56 );
nand NAND2_25245 ( P2_ADD_391_1196_U441 , P2_R2182_U89 , P2_ADD_391_1196_U57 );
nand NAND2_25246 ( P2_ADD_391_1196_U442 , P2_R2096_U90 , P2_ADD_391_1196_U56 );
nand NAND2_25247 ( P2_ADD_391_1196_U443 , P2_R2182_U89 , P2_ADD_391_1196_U57 );
nand NAND2_25248 ( P2_ADD_391_1196_U444 , P2_ADD_391_1196_U443 , P2_ADD_391_1196_U442 );
nand NAND2_25249 ( P2_ADD_391_1196_U445 , P2_ADD_391_1196_U149 , P2_ADD_391_1196_U150 );
nand NAND2_25250 ( P2_ADD_391_1196_U446 , P2_ADD_391_1196_U231 , P2_ADD_391_1196_U444 );
nand NAND2_25251 ( P2_ADD_391_1196_U447 , P2_R2096_U91 , P2_ADD_391_1196_U54 );
nand NAND2_25252 ( P2_ADD_391_1196_U448 , P2_R2182_U90 , P2_ADD_391_1196_U55 );
nand NAND2_25253 ( P2_ADD_391_1196_U449 , P2_R2096_U91 , P2_ADD_391_1196_U54 );
nand NAND2_25254 ( P2_ADD_391_1196_U450 , P2_R2182_U90 , P2_ADD_391_1196_U55 );
nand NAND2_25255 ( P2_ADD_391_1196_U451 , P2_ADD_391_1196_U450 , P2_ADD_391_1196_U449 );
nand NAND2_25256 ( P2_ADD_391_1196_U452 , P2_ADD_391_1196_U151 , P2_ADD_391_1196_U152 );
nand NAND2_25257 ( P2_ADD_391_1196_U453 , P2_ADD_391_1196_U227 , P2_ADD_391_1196_U451 );
nand NAND2_25258 ( P2_ADD_391_1196_U454 , P2_R2096_U92 , P2_ADD_391_1196_U40 );
nand NAND2_25259 ( P2_ADD_391_1196_U455 , P2_R2182_U91 , P2_ADD_391_1196_U41 );
nand NAND2_25260 ( P2_ADD_391_1196_U456 , P2_R2096_U93 , P2_ADD_391_1196_U42 );
nand NAND2_25261 ( P2_ADD_391_1196_U457 , P2_R2182_U92 , P2_ADD_391_1196_U43 );
nand NAND2_25262 ( P2_ADD_391_1196_U458 , P2_ADD_391_1196_U457 , P2_ADD_391_1196_U456 );
nand NAND2_25263 ( P2_ADD_391_1196_U459 , P2_ADD_391_1196_U304 , P2_ADD_391_1196_U53 );
nand NAND2_25264 ( P2_ADD_391_1196_U460 , P2_ADD_391_1196_U458 , P2_ADD_391_1196_U221 );
nand NAND2_25265 ( P2_ADD_391_1196_U461 , P2_R2096_U94 , P2_ADD_391_1196_U44 );
nand NAND2_25266 ( P2_ADD_391_1196_U462 , P2_R2182_U93 , P2_ADD_391_1196_U45 );
nand NAND2_25267 ( P2_ADD_391_1196_U463 , P2_R2096_U95 , P2_ADD_391_1196_U51 );
nand NAND2_25268 ( P2_ADD_391_1196_U464 , P2_R2182_U94 , P2_ADD_391_1196_U52 );
nand NAND2_25269 ( P2_ADD_391_1196_U465 , P2_R2096_U95 , P2_ADD_391_1196_U51 );
nand NAND2_25270 ( P2_ADD_391_1196_U466 , P2_R2182_U94 , P2_ADD_391_1196_U52 );
nand NAND2_25271 ( P2_ADD_391_1196_U467 , P2_ADD_391_1196_U466 , P2_ADD_391_1196_U465 );
nand NAND2_25272 ( P2_ADD_391_1196_U468 , P2_ADD_391_1196_U155 , P2_ADD_391_1196_U156 );
nand NAND2_25273 ( P2_ADD_391_1196_U469 , P2_ADD_391_1196_U213 , P2_ADD_391_1196_U467 );
nand NAND2_25274 ( P2_ADD_391_1196_U470 , P2_R2096_U96 , P2_ADD_391_1196_U46 );
nand NAND2_25275 ( P2_ADD_391_1196_U471 , P2_R2182_U95 , P2_ADD_391_1196_U47 );
nand NAND2_25276 ( P2_ADD_391_1196_U472 , P2_R2096_U97 , P2_ADD_391_1196_U48 );
nand NAND2_25277 ( P2_ADD_391_1196_U473 , P2_R2182_U96 , P2_ADD_391_1196_U49 );
nand NAND2_25278 ( P2_ADD_391_1196_U474 , P2_ADD_391_1196_U473 , P2_ADD_391_1196_U472 );
nand NAND2_25279 ( P2_ADD_391_1196_U475 , P2_ADD_391_1196_U305 , P2_ADD_391_1196_U50 );
nand NAND2_25280 ( P2_ADD_391_1196_U476 , P2_ADD_391_1196_U474 , P2_ADD_391_1196_U207 );
nand NAND2_25281 ( P2_ADD_391_1196_U477 , P2_R2182_U69 , P2_ADD_391_1196_U19 );
nand NAND2_25282 ( P2_ADD_391_1196_U478 , P2_R2096_U68 , P2_ADD_391_1196_U20 );
not NOT1_25283 ( P2_ADD_402_1132_U4 , P2_U2606 );
not NOT1_25284 ( P2_ADD_402_1132_U5 , P2_U2591 );
nand NAND2_25285 ( P2_ADD_402_1132_U6 , P2_U2591 , P2_U2606 );
not NOT1_25286 ( P2_ADD_402_1132_U7 , P2_U2592 );
nand NAND2_25287 ( P2_ADD_402_1132_U8 , P2_U2592 , P2_ADD_402_1132_U28 );
not NOT1_25288 ( P2_ADD_402_1132_U9 , P2_U2593 );
nand NAND2_25289 ( P2_ADD_402_1132_U10 , P2_U2593 , P2_ADD_402_1132_U29 );
not NOT1_25290 ( P2_ADD_402_1132_U11 , P2_U2594 );
nand NAND2_25291 ( P2_ADD_402_1132_U12 , P2_U2594 , P2_ADD_402_1132_U30 );
not NOT1_25292 ( P2_ADD_402_1132_U13 , P2_U2595 );
nand NAND2_25293 ( P2_ADD_402_1132_U14 , P2_U2595 , P2_ADD_402_1132_U31 );
not NOT1_25294 ( P2_ADD_402_1132_U15 , P2_U2596 );
nand NAND2_25295 ( P2_ADD_402_1132_U16 , P2_U2596 , P2_ADD_402_1132_U32 );
not NOT1_25296 ( P2_ADD_402_1132_U17 , P2_U2597 );
nand NAND2_25297 ( P2_ADD_402_1132_U18 , P2_ADD_402_1132_U36 , P2_ADD_402_1132_U35 );
nand NAND2_25298 ( P2_ADD_402_1132_U19 , P2_ADD_402_1132_U38 , P2_ADD_402_1132_U37 );
nand NAND2_25299 ( P2_ADD_402_1132_U20 , P2_ADD_402_1132_U40 , P2_ADD_402_1132_U39 );
nand NAND2_25300 ( P2_ADD_402_1132_U21 , P2_ADD_402_1132_U42 , P2_ADD_402_1132_U41 );
nand NAND2_25301 ( P2_ADD_402_1132_U22 , P2_ADD_402_1132_U44 , P2_ADD_402_1132_U43 );
nand NAND2_25302 ( P2_ADD_402_1132_U23 , P2_ADD_402_1132_U46 , P2_ADD_402_1132_U45 );
nand NAND2_25303 ( P2_ADD_402_1132_U24 , P2_ADD_402_1132_U48 , P2_ADD_402_1132_U47 );
nand NAND2_25304 ( P2_ADD_402_1132_U25 , P2_ADD_402_1132_U50 , P2_ADD_402_1132_U49 );
not NOT1_25305 ( P2_ADD_402_1132_U26 , P2_U2598 );
nand NAND2_25306 ( P2_ADD_402_1132_U27 , P2_U2597 , P2_ADD_402_1132_U33 );
not NOT1_25307 ( P2_ADD_402_1132_U28 , P2_ADD_402_1132_U6 );
not NOT1_25308 ( P2_ADD_402_1132_U29 , P2_ADD_402_1132_U8 );
not NOT1_25309 ( P2_ADD_402_1132_U30 , P2_ADD_402_1132_U10 );
not NOT1_25310 ( P2_ADD_402_1132_U31 , P2_ADD_402_1132_U12 );
not NOT1_25311 ( P2_ADD_402_1132_U32 , P2_ADD_402_1132_U14 );
not NOT1_25312 ( P2_ADD_402_1132_U33 , P2_ADD_402_1132_U16 );
not NOT1_25313 ( P2_ADD_402_1132_U34 , P2_ADD_402_1132_U27 );
nand NAND2_25314 ( P2_ADD_402_1132_U35 , P2_U2598 , P2_ADD_402_1132_U27 );
nand NAND2_25315 ( P2_ADD_402_1132_U36 , P2_ADD_402_1132_U34 , P2_ADD_402_1132_U26 );
nand NAND2_25316 ( P2_ADD_402_1132_U37 , P2_U2597 , P2_ADD_402_1132_U16 );
nand NAND2_25317 ( P2_ADD_402_1132_U38 , P2_ADD_402_1132_U33 , P2_ADD_402_1132_U17 );
nand NAND2_25318 ( P2_ADD_402_1132_U39 , P2_U2592 , P2_ADD_402_1132_U6 );
nand NAND2_25319 ( P2_ADD_402_1132_U40 , P2_ADD_402_1132_U28 , P2_ADD_402_1132_U7 );
nand NAND2_25320 ( P2_ADD_402_1132_U41 , P2_U2594 , P2_ADD_402_1132_U10 );
nand NAND2_25321 ( P2_ADD_402_1132_U42 , P2_ADD_402_1132_U30 , P2_ADD_402_1132_U11 );
nand NAND2_25322 ( P2_ADD_402_1132_U43 , P2_U2595 , P2_ADD_402_1132_U12 );
nand NAND2_25323 ( P2_ADD_402_1132_U44 , P2_ADD_402_1132_U31 , P2_ADD_402_1132_U13 );
nand NAND2_25324 ( P2_ADD_402_1132_U45 , P2_U2591 , P2_ADD_402_1132_U4 );
nand NAND2_25325 ( P2_ADD_402_1132_U46 , P2_U2606 , P2_ADD_402_1132_U5 );
nand NAND2_25326 ( P2_ADD_402_1132_U47 , P2_U2596 , P2_ADD_402_1132_U14 );
nand NAND2_25327 ( P2_ADD_402_1132_U48 , P2_ADD_402_1132_U32 , P2_ADD_402_1132_U15 );
nand NAND2_25328 ( P2_ADD_402_1132_U49 , P2_U2593 , P2_ADD_402_1132_U8 );
nand NAND2_25329 ( P2_ADD_402_1132_U50 , P2_ADD_402_1132_U29 , P2_ADD_402_1132_U9 );
not NOT1_25330 ( P2_SUB_563_U6 , P2_U3618 );
not NOT1_25331 ( P2_SUB_563_U7 , P2_U3619 );
and AND2_25332 ( P2_R2182_U4 , P2_U2671 , P2_R2182_U20 );
and AND2_25333 ( P2_R2182_U5 , P2_U2670 , P2_R2182_U4 );
and AND2_25334 ( P2_R2182_U6 , P2_U2669 , P2_R2182_U5 );
and AND2_25335 ( P2_R2182_U7 , P2_U2690 , P2_R2182_U8 );
and AND2_25336 ( P2_R2182_U8 , P2_U2691 , P2_R2182_U11 );
and AND2_25337 ( P2_R2182_U9 , P2_U2675 , P2_R2182_U21 );
and AND2_25338 ( P2_R2182_U10 , P2_U2674 , P2_R2182_U9 );
and AND2_25339 ( P2_R2182_U11 , P2_U2692 , P2_R2182_U13 );
and AND2_25340 ( P2_R2182_U12 , P2_U2694 , P2_R2182_U18 );
and AND2_25341 ( P2_R2182_U13 , P2_U2693 , P2_R2182_U12 );
and AND2_25342 ( P2_R2182_U14 , P2_U2668 , P2_R2182_U6 );
and AND2_25343 ( P2_R2182_U15 , P2_U2667 , P2_R2182_U14 );
and AND2_25344 ( P2_R2182_U16 , P2_U2666 , P2_R2182_U15 );
and AND2_25345 ( P2_R2182_U17 , P2_U2696 , P2_R2182_U16 );
and AND2_25346 ( P2_R2182_U18 , P2_U2695 , P2_R2182_U17 );
and AND2_25347 ( P2_R2182_U19 , P2_U2673 , P2_R2182_U10 );
and AND2_25348 ( P2_R2182_U20 , P2_U2672 , P2_R2182_U19 );
and AND2_25349 ( P2_R2182_U21 , P2_U2676 , P2_R2182_U102 );
not NOT1_25350 ( P2_R2182_U22 , P2_U2675 );
not NOT1_25351 ( P2_R2182_U23 , P2_U2671 );
not NOT1_25352 ( P2_R2182_U24 , P2_U2676 );
not NOT1_25353 ( P2_R2182_U25 , P2_U2666 );
not NOT1_25354 ( P2_R2182_U26 , P2_U2667 );
not NOT1_25355 ( P2_R2182_U27 , P2_U2696 );
not NOT1_25356 ( P2_R2182_U28 , P2_U2695 );
not NOT1_25357 ( P2_R2182_U29 , P2_U2694 );
not NOT1_25358 ( P2_R2182_U30 , P2_U2693 );
not NOT1_25359 ( P2_R2182_U31 , P2_U2692 );
not NOT1_25360 ( P2_R2182_U32 , P2_U2691 );
not NOT1_25361 ( P2_R2182_U33 , P2_U2670 );
not NOT1_25362 ( P2_R2182_U34 , P2_U2672 );
not NOT1_25363 ( P2_R2182_U35 , P2_U2674 );
not NOT1_25364 ( P2_R2182_U36 , P2_U2673 );
not NOT1_25365 ( P2_R2182_U37 , P2_U2690 );
not NOT1_25366 ( P2_R2182_U38 , P2_U2668 );
not NOT1_25367 ( P2_R2182_U39 , P2_U2669 );
and AND2_25368 ( P2_R2182_U40 , P2_R2182_U192 , P2_R2182_U190 );
and AND2_25369 ( P2_R2182_U41 , P2_R2182_U186 , P2_R2182_U182 );
not NOT1_25370 ( P2_R2182_U42 , P2_U2700 );
not NOT1_25371 ( P2_R2182_U43 , P2_U2679 );
not NOT1_25372 ( P2_R2182_U44 , P2_U2702 );
not NOT1_25373 ( P2_R2182_U45 , P2_U2681 );
nand NAND2_25374 ( P2_R2182_U46 , P2_U2681 , P2_U2702 );
not NOT1_25375 ( P2_R2182_U47 , P2_U2680 );
not NOT1_25376 ( P2_R2182_U48 , P2_U2699 );
not NOT1_25377 ( P2_R2182_U49 , P2_U2678 );
not NOT1_25378 ( P2_R2182_U50 , P2_U2698 );
not NOT1_25379 ( P2_R2182_U51 , P2_U2677 );
not NOT1_25380 ( P2_R2182_U52 , P2_U2689 );
not NOT1_25381 ( P2_R2182_U53 , P2_U2665 );
not NOT1_25382 ( P2_R2182_U54 , P2_U2688 );
not NOT1_25383 ( P2_R2182_U55 , P2_U2664 );
not NOT1_25384 ( P2_R2182_U56 , P2_U2687 );
not NOT1_25385 ( P2_R2182_U57 , P2_U2663 );
not NOT1_25386 ( P2_R2182_U58 , P2_U2686 );
not NOT1_25387 ( P2_R2182_U59 , P2_U2662 );
not NOT1_25388 ( P2_R2182_U60 , P2_U2685 );
not NOT1_25389 ( P2_R2182_U61 , P2_U2661 );
not NOT1_25390 ( P2_R2182_U62 , P2_U2684 );
not NOT1_25391 ( P2_R2182_U63 , P2_U2660 );
not NOT1_25392 ( P2_R2182_U64 , P2_U2683 );
not NOT1_25393 ( P2_R2182_U65 , P2_U2659 );
nand NAND2_25394 ( P2_R2182_U66 , P2_R2182_U177 , P2_R2182_U176 );
not NOT1_25395 ( P2_R2182_U67 , P2_U2701 );
nand NAND2_25396 ( P2_R2182_U68 , P2_R2182_U283 , P2_R2182_U282 );
nand NAND2_25397 ( P2_R2182_U69 , P2_R2182_U305 , P2_R2182_U304 );
nand NAND2_25398 ( P2_R2182_U70 , P2_R2182_U194 , P2_R2182_U193 );
nand NAND2_25399 ( P2_R2182_U71 , P2_R2182_U196 , P2_R2182_U195 );
nand NAND2_25400 ( P2_R2182_U72 , P2_R2182_U198 , P2_R2182_U197 );
nand NAND2_25401 ( P2_R2182_U73 , P2_R2182_U200 , P2_R2182_U199 );
nand NAND2_25402 ( P2_R2182_U74 , P2_R2182_U202 , P2_R2182_U201 );
nand NAND2_25403 ( P2_R2182_U75 , P2_R2182_U209 , P2_R2182_U208 );
nand NAND2_25404 ( P2_R2182_U76 , P2_R2182_U216 , P2_R2182_U215 );
nand NAND2_25405 ( P2_R2182_U77 , P2_R2182_U230 , P2_R2182_U229 );
nand NAND2_25406 ( P2_R2182_U78 , P2_R2182_U237 , P2_R2182_U236 );
nand NAND2_25407 ( P2_R2182_U79 , P2_R2182_U244 , P2_R2182_U243 );
nand NAND2_25408 ( P2_R2182_U80 , P2_R2182_U251 , P2_R2182_U250 );
nand NAND2_25409 ( P2_R2182_U81 , P2_R2182_U258 , P2_R2182_U257 );
nand NAND2_25410 ( P2_R2182_U82 , P2_R2182_U265 , P2_R2182_U264 );
nand NAND2_25411 ( P2_R2182_U83 , P2_R2182_U272 , P2_R2182_U271 );
nand NAND2_25412 ( P2_R2182_U84 , P2_R2182_U274 , P2_R2182_U273 );
nand NAND2_25413 ( P2_R2182_U85 , P2_R2182_U276 , P2_R2182_U275 );
nand NAND2_25414 ( P2_R2182_U86 , P2_R2182_U278 , P2_R2182_U277 );
nand NAND2_25415 ( P2_R2182_U87 , P2_R2182_U285 , P2_R2182_U284 );
nand NAND2_25416 ( P2_R2182_U88 , P2_R2182_U287 , P2_R2182_U286 );
nand NAND2_25417 ( P2_R2182_U89 , P2_R2182_U289 , P2_R2182_U288 );
nand NAND2_25418 ( P2_R2182_U90 , P2_R2182_U291 , P2_R2182_U290 );
nand NAND2_25419 ( P2_R2182_U91 , P2_R2182_U293 , P2_R2182_U292 );
nand NAND2_25420 ( P2_R2182_U92 , P2_R2182_U295 , P2_R2182_U294 );
nand NAND2_25421 ( P2_R2182_U93 , P2_R2182_U297 , P2_R2182_U296 );
nand NAND2_25422 ( P2_R2182_U94 , P2_R2182_U299 , P2_R2182_U298 );
nand NAND2_25423 ( P2_R2182_U95 , P2_R2182_U301 , P2_R2182_U300 );
nand NAND2_25424 ( P2_R2182_U96 , P2_R2182_U303 , P2_R2182_U302 );
and AND3_25425 ( P2_R2182_U97 , P2_R2182_U218 , P2_R2182_U217 , P2_R2182_U181 );
and AND2_25426 ( P2_R2182_U98 , P2_R2182_U185 , P2_R2182_U221 );
and AND3_25427 ( P2_R2182_U99 , P2_R2182_U223 , P2_R2182_U222 , P2_R2182_U189 );
and AND2_25428 ( P2_R2182_U100 , P2_R2182_U191 , P2_R2182_U125 );
nand NAND2_25429 ( P2_R2182_U101 , P2_R2182_U280 , P2_R2182_U279 );
nand NAND2_25430 ( P2_R2182_U102 , P2_R2182_U135 , P2_R2182_U134 );
and AND2_25431 ( P2_R2182_U103 , P2_R2182_U204 , P2_R2182_U203 );
nand NAND2_25432 ( P2_R2182_U104 , P2_R2182_U131 , P2_R2182_U130 );
and AND2_25433 ( P2_R2182_U105 , P2_R2182_U211 , P2_R2182_U210 );
nand NAND2_25434 ( P2_R2182_U106 , P2_R2182_U126 , P2_R2182_U127 );
not NOT1_25435 ( P2_R2182_U107 , P2_U2658 );
not NOT1_25436 ( P2_R2182_U108 , P2_U2682 );
and AND2_25437 ( P2_R2182_U109 , P2_R2182_U225 , P2_R2182_U224 );
and AND2_25438 ( P2_R2182_U110 , P2_R2182_U232 , P2_R2182_U231 );
nand NAND2_25439 ( P2_R2182_U111 , P2_R2182_U173 , P2_R2182_U172 );
and AND2_25440 ( P2_R2182_U112 , P2_R2182_U239 , P2_R2182_U238 );
nand NAND2_25441 ( P2_R2182_U113 , P2_R2182_U169 , P2_R2182_U168 );
and AND2_25442 ( P2_R2182_U114 , P2_R2182_U246 , P2_R2182_U245 );
nand NAND2_25443 ( P2_R2182_U115 , P2_R2182_U165 , P2_R2182_U164 );
and AND2_25444 ( P2_R2182_U116 , P2_R2182_U253 , P2_R2182_U252 );
nand NAND2_25445 ( P2_R2182_U117 , P2_R2182_U161 , P2_R2182_U160 );
and AND2_25446 ( P2_R2182_U118 , P2_R2182_U260 , P2_R2182_U259 );
nand NAND2_25447 ( P2_R2182_U119 , P2_R2182_U157 , P2_R2182_U156 );
and AND2_25448 ( P2_R2182_U120 , P2_R2182_U267 , P2_R2182_U266 );
not NOT1_25449 ( P2_R2182_U121 , P2_R2182_U46 );
nand NAND2_25450 ( P2_R2182_U122 , P2_U2680 , P2_R2182_U121 );
nand NAND2_25451 ( P2_R2182_U123 , P2_R2182_U122 , P2_R2182_U67 );
or OR2_25452 ( P2_R2182_U124 , P2_U2679 , P2_U2700 );
nand NAND2_25453 ( P2_R2182_U125 , P2_R2182_U46 , P2_R2182_U47 );
nand NAND3_25454 ( P2_R2182_U126 , P2_R2182_U125 , P2_R2182_U123 , P2_R2182_U124 );
nand NAND2_25455 ( P2_R2182_U127 , P2_U2679 , P2_U2700 );
not NOT1_25456 ( P2_R2182_U128 , P2_R2182_U106 );
or OR2_25457 ( P2_R2182_U129 , P2_U2699 , P2_U2678 );
nand NAND2_25458 ( P2_R2182_U130 , P2_R2182_U129 , P2_R2182_U106 );
nand NAND2_25459 ( P2_R2182_U131 , P2_U2678 , P2_U2699 );
not NOT1_25460 ( P2_R2182_U132 , P2_R2182_U104 );
or OR2_25461 ( P2_R2182_U133 , P2_U2698 , P2_U2677 );
nand NAND2_25462 ( P2_R2182_U134 , P2_R2182_U133 , P2_R2182_U104 );
nand NAND2_25463 ( P2_R2182_U135 , P2_U2677 , P2_U2698 );
not NOT1_25464 ( P2_R2182_U136 , P2_R2182_U102 );
not NOT1_25465 ( P2_R2182_U137 , P2_R2182_U21 );
not NOT1_25466 ( P2_R2182_U138 , P2_R2182_U9 );
not NOT1_25467 ( P2_R2182_U139 , P2_R2182_U10 );
not NOT1_25468 ( P2_R2182_U140 , P2_R2182_U19 );
not NOT1_25469 ( P2_R2182_U141 , P2_R2182_U20 );
not NOT1_25470 ( P2_R2182_U142 , P2_R2182_U4 );
not NOT1_25471 ( P2_R2182_U143 , P2_R2182_U5 );
not NOT1_25472 ( P2_R2182_U144 , P2_R2182_U6 );
not NOT1_25473 ( P2_R2182_U145 , P2_R2182_U14 );
not NOT1_25474 ( P2_R2182_U146 , P2_R2182_U15 );
not NOT1_25475 ( P2_R2182_U147 , P2_R2182_U16 );
not NOT1_25476 ( P2_R2182_U148 , P2_R2182_U17 );
not NOT1_25477 ( P2_R2182_U149 , P2_R2182_U18 );
not NOT1_25478 ( P2_R2182_U150 , P2_R2182_U12 );
not NOT1_25479 ( P2_R2182_U151 , P2_R2182_U13 );
not NOT1_25480 ( P2_R2182_U152 , P2_R2182_U11 );
not NOT1_25481 ( P2_R2182_U153 , P2_R2182_U8 );
not NOT1_25482 ( P2_R2182_U154 , P2_R2182_U7 );
or OR2_25483 ( P2_R2182_U155 , P2_U2689 , P2_U2665 );
nand NAND2_25484 ( P2_R2182_U156 , P2_R2182_U155 , P2_R2182_U7 );
nand NAND2_25485 ( P2_R2182_U157 , P2_U2665 , P2_U2689 );
not NOT1_25486 ( P2_R2182_U158 , P2_R2182_U119 );
or OR2_25487 ( P2_R2182_U159 , P2_U2688 , P2_U2664 );
nand NAND2_25488 ( P2_R2182_U160 , P2_R2182_U159 , P2_R2182_U119 );
nand NAND2_25489 ( P2_R2182_U161 , P2_U2664 , P2_U2688 );
not NOT1_25490 ( P2_R2182_U162 , P2_R2182_U117 );
or OR2_25491 ( P2_R2182_U163 , P2_U2687 , P2_U2663 );
nand NAND2_25492 ( P2_R2182_U164 , P2_R2182_U163 , P2_R2182_U117 );
nand NAND2_25493 ( P2_R2182_U165 , P2_U2663 , P2_U2687 );
not NOT1_25494 ( P2_R2182_U166 , P2_R2182_U115 );
or OR2_25495 ( P2_R2182_U167 , P2_U2686 , P2_U2662 );
nand NAND2_25496 ( P2_R2182_U168 , P2_R2182_U167 , P2_R2182_U115 );
nand NAND2_25497 ( P2_R2182_U169 , P2_U2662 , P2_U2686 );
not NOT1_25498 ( P2_R2182_U170 , P2_R2182_U113 );
or OR2_25499 ( P2_R2182_U171 , P2_U2685 , P2_U2661 );
nand NAND2_25500 ( P2_R2182_U172 , P2_R2182_U171 , P2_R2182_U113 );
nand NAND2_25501 ( P2_R2182_U173 , P2_U2661 , P2_U2685 );
not NOT1_25502 ( P2_R2182_U174 , P2_R2182_U111 );
or OR2_25503 ( P2_R2182_U175 , P2_U2684 , P2_U2660 );
nand NAND2_25504 ( P2_R2182_U176 , P2_R2182_U175 , P2_R2182_U111 );
nand NAND2_25505 ( P2_R2182_U177 , P2_U2660 , P2_U2684 );
not NOT1_25506 ( P2_R2182_U178 , P2_R2182_U66 );
or OR2_25507 ( P2_R2182_U179 , P2_U2683 , P2_U2659 );
nand NAND2_25508 ( P2_R2182_U180 , P2_R2182_U179 , P2_R2182_U66 );
nand NAND2_25509 ( P2_R2182_U181 , P2_U2659 , P2_U2683 );
nand NAND2_25510 ( P2_R2182_U182 , P2_R2182_U97 , P2_R2182_U180 );
nand NAND2_25511 ( P2_R2182_U183 , P2_U2659 , P2_U2683 );
nand NAND2_25512 ( P2_R2182_U184 , P2_R2182_U178 , P2_R2182_U183 );
or OR2_25513 ( P2_R2182_U185 , P2_U2659 , P2_U2683 );
nand NAND2_25514 ( P2_R2182_U186 , P2_R2182_U98 , P2_R2182_U184 );
nand NAND2_25515 ( P2_R2182_U187 , P2_R2182_U47 , P2_R2182_U46 );
nand NAND2_25516 ( P2_R2182_U188 , P2_U2701 , P2_R2182_U187 );
nand NAND2_25517 ( P2_R2182_U189 , P2_U2680 , P2_R2182_U121 );
nand NAND2_25518 ( P2_R2182_U190 , P2_R2182_U99 , P2_R2182_U188 );
nand NAND2_25519 ( P2_R2182_U191 , P2_U2679 , P2_U2700 );
nand NAND3_25520 ( P2_R2182_U192 , P2_R2182_U124 , P2_R2182_U123 , P2_R2182_U100 );
nand NAND2_25521 ( P2_R2182_U193 , P2_R2182_U34 , P2_R2182_U19 );
nand NAND2_25522 ( P2_R2182_U194 , P2_R2182_U140 , P2_U2672 );
nand NAND2_25523 ( P2_R2182_U195 , P2_R2182_U36 , P2_R2182_U10 );
nand NAND2_25524 ( P2_R2182_U196 , P2_R2182_U139 , P2_U2673 );
nand NAND2_25525 ( P2_R2182_U197 , P2_R2182_U35 , P2_R2182_U9 );
nand NAND2_25526 ( P2_R2182_U198 , P2_R2182_U138 , P2_U2674 );
nand NAND2_25527 ( P2_R2182_U199 , P2_R2182_U22 , P2_R2182_U21 );
nand NAND2_25528 ( P2_R2182_U200 , P2_R2182_U137 , P2_U2675 );
nand NAND2_25529 ( P2_R2182_U201 , P2_R2182_U24 , P2_R2182_U102 );
nand NAND2_25530 ( P2_R2182_U202 , P2_R2182_U136 , P2_U2676 );
nand NAND2_25531 ( P2_R2182_U203 , P2_U2677 , P2_R2182_U50 );
nand NAND2_25532 ( P2_R2182_U204 , P2_U2698 , P2_R2182_U51 );
nand NAND2_25533 ( P2_R2182_U205 , P2_U2677 , P2_R2182_U50 );
nand NAND2_25534 ( P2_R2182_U206 , P2_U2698 , P2_R2182_U51 );
nand NAND2_25535 ( P2_R2182_U207 , P2_R2182_U206 , P2_R2182_U205 );
nand NAND2_25536 ( P2_R2182_U208 , P2_R2182_U103 , P2_R2182_U104 );
nand NAND2_25537 ( P2_R2182_U209 , P2_R2182_U132 , P2_R2182_U207 );
nand NAND2_25538 ( P2_R2182_U210 , P2_U2678 , P2_R2182_U48 );
nand NAND2_25539 ( P2_R2182_U211 , P2_U2699 , P2_R2182_U49 );
nand NAND2_25540 ( P2_R2182_U212 , P2_U2678 , P2_R2182_U48 );
nand NAND2_25541 ( P2_R2182_U213 , P2_U2699 , P2_R2182_U49 );
nand NAND2_25542 ( P2_R2182_U214 , P2_R2182_U213 , P2_R2182_U212 );
nand NAND2_25543 ( P2_R2182_U215 , P2_R2182_U105 , P2_R2182_U106 );
nand NAND2_25544 ( P2_R2182_U216 , P2_R2182_U128 , P2_R2182_U214 );
nand NAND2_25545 ( P2_R2182_U217 , P2_U2658 , P2_R2182_U108 );
nand NAND2_25546 ( P2_R2182_U218 , P2_U2682 , P2_R2182_U107 );
nand NAND2_25547 ( P2_R2182_U219 , P2_U2658 , P2_R2182_U108 );
nand NAND2_25548 ( P2_R2182_U220 , P2_U2682 , P2_R2182_U107 );
nand NAND2_25549 ( P2_R2182_U221 , P2_R2182_U220 , P2_R2182_U219 );
nand NAND2_25550 ( P2_R2182_U222 , P2_U2679 , P2_R2182_U42 );
nand NAND2_25551 ( P2_R2182_U223 , P2_U2700 , P2_R2182_U43 );
nand NAND2_25552 ( P2_R2182_U224 , P2_U2659 , P2_R2182_U64 );
nand NAND2_25553 ( P2_R2182_U225 , P2_U2683 , P2_R2182_U65 );
nand NAND2_25554 ( P2_R2182_U226 , P2_U2659 , P2_R2182_U64 );
nand NAND2_25555 ( P2_R2182_U227 , P2_U2683 , P2_R2182_U65 );
nand NAND2_25556 ( P2_R2182_U228 , P2_R2182_U227 , P2_R2182_U226 );
nand NAND2_25557 ( P2_R2182_U229 , P2_R2182_U109 , P2_R2182_U66 );
nand NAND2_25558 ( P2_R2182_U230 , P2_R2182_U228 , P2_R2182_U178 );
nand NAND2_25559 ( P2_R2182_U231 , P2_U2660 , P2_R2182_U62 );
nand NAND2_25560 ( P2_R2182_U232 , P2_U2684 , P2_R2182_U63 );
nand NAND2_25561 ( P2_R2182_U233 , P2_U2660 , P2_R2182_U62 );
nand NAND2_25562 ( P2_R2182_U234 , P2_U2684 , P2_R2182_U63 );
nand NAND2_25563 ( P2_R2182_U235 , P2_R2182_U234 , P2_R2182_U233 );
nand NAND2_25564 ( P2_R2182_U236 , P2_R2182_U110 , P2_R2182_U111 );
nand NAND2_25565 ( P2_R2182_U237 , P2_R2182_U174 , P2_R2182_U235 );
nand NAND2_25566 ( P2_R2182_U238 , P2_U2661 , P2_R2182_U60 );
nand NAND2_25567 ( P2_R2182_U239 , P2_U2685 , P2_R2182_U61 );
nand NAND2_25568 ( P2_R2182_U240 , P2_U2661 , P2_R2182_U60 );
nand NAND2_25569 ( P2_R2182_U241 , P2_U2685 , P2_R2182_U61 );
nand NAND2_25570 ( P2_R2182_U242 , P2_R2182_U241 , P2_R2182_U240 );
nand NAND2_25571 ( P2_R2182_U243 , P2_R2182_U112 , P2_R2182_U113 );
nand NAND2_25572 ( P2_R2182_U244 , P2_R2182_U170 , P2_R2182_U242 );
nand NAND2_25573 ( P2_R2182_U245 , P2_U2662 , P2_R2182_U58 );
nand NAND2_25574 ( P2_R2182_U246 , P2_U2686 , P2_R2182_U59 );
nand NAND2_25575 ( P2_R2182_U247 , P2_U2662 , P2_R2182_U58 );
nand NAND2_25576 ( P2_R2182_U248 , P2_U2686 , P2_R2182_U59 );
nand NAND2_25577 ( P2_R2182_U249 , P2_R2182_U248 , P2_R2182_U247 );
nand NAND2_25578 ( P2_R2182_U250 , P2_R2182_U114 , P2_R2182_U115 );
nand NAND2_25579 ( P2_R2182_U251 , P2_R2182_U166 , P2_R2182_U249 );
nand NAND2_25580 ( P2_R2182_U252 , P2_U2663 , P2_R2182_U56 );
nand NAND2_25581 ( P2_R2182_U253 , P2_U2687 , P2_R2182_U57 );
nand NAND2_25582 ( P2_R2182_U254 , P2_U2663 , P2_R2182_U56 );
nand NAND2_25583 ( P2_R2182_U255 , P2_U2687 , P2_R2182_U57 );
nand NAND2_25584 ( P2_R2182_U256 , P2_R2182_U255 , P2_R2182_U254 );
nand NAND2_25585 ( P2_R2182_U257 , P2_R2182_U116 , P2_R2182_U117 );
nand NAND2_25586 ( P2_R2182_U258 , P2_R2182_U162 , P2_R2182_U256 );
nand NAND2_25587 ( P2_R2182_U259 , P2_U2664 , P2_R2182_U54 );
nand NAND2_25588 ( P2_R2182_U260 , P2_U2688 , P2_R2182_U55 );
nand NAND2_25589 ( P2_R2182_U261 , P2_U2664 , P2_R2182_U54 );
nand NAND2_25590 ( P2_R2182_U262 , P2_U2688 , P2_R2182_U55 );
nand NAND2_25591 ( P2_R2182_U263 , P2_R2182_U262 , P2_R2182_U261 );
nand NAND2_25592 ( P2_R2182_U264 , P2_R2182_U118 , P2_R2182_U119 );
nand NAND2_25593 ( P2_R2182_U265 , P2_R2182_U158 , P2_R2182_U263 );
nand NAND2_25594 ( P2_R2182_U266 , P2_U2665 , P2_R2182_U52 );
nand NAND2_25595 ( P2_R2182_U267 , P2_U2689 , P2_R2182_U53 );
nand NAND2_25596 ( P2_R2182_U268 , P2_U2665 , P2_R2182_U52 );
nand NAND2_25597 ( P2_R2182_U269 , P2_U2689 , P2_R2182_U53 );
nand NAND2_25598 ( P2_R2182_U270 , P2_R2182_U269 , P2_R2182_U268 );
nand NAND2_25599 ( P2_R2182_U271 , P2_R2182_U120 , P2_R2182_U7 );
nand NAND2_25600 ( P2_R2182_U272 , P2_R2182_U154 , P2_R2182_U270 );
nand NAND2_25601 ( P2_R2182_U273 , P2_R2182_U37 , P2_R2182_U8 );
nand NAND2_25602 ( P2_R2182_U274 , P2_R2182_U153 , P2_U2690 );
nand NAND2_25603 ( P2_R2182_U275 , P2_R2182_U32 , P2_R2182_U11 );
nand NAND2_25604 ( P2_R2182_U276 , P2_R2182_U152 , P2_U2691 );
nand NAND2_25605 ( P2_R2182_U277 , P2_R2182_U31 , P2_R2182_U13 );
nand NAND2_25606 ( P2_R2182_U278 , P2_R2182_U151 , P2_U2692 );
nand NAND2_25607 ( P2_R2182_U279 , P2_R2182_U121 , P2_R2182_U47 );
nand NAND2_25608 ( P2_R2182_U280 , P2_U2680 , P2_R2182_U46 );
not NOT1_25609 ( P2_R2182_U281 , P2_R2182_U101 );
nand NAND2_25610 ( P2_R2182_U282 , P2_R2182_U281 , P2_U2701 );
nand NAND2_25611 ( P2_R2182_U283 , P2_R2182_U101 , P2_R2182_U67 );
nand NAND2_25612 ( P2_R2182_U284 , P2_R2182_U30 , P2_R2182_U12 );
nand NAND2_25613 ( P2_R2182_U285 , P2_R2182_U150 , P2_U2693 );
nand NAND2_25614 ( P2_R2182_U286 , P2_R2182_U29 , P2_R2182_U18 );
nand NAND2_25615 ( P2_R2182_U287 , P2_R2182_U149 , P2_U2694 );
nand NAND2_25616 ( P2_R2182_U288 , P2_R2182_U28 , P2_R2182_U17 );
nand NAND2_25617 ( P2_R2182_U289 , P2_R2182_U148 , P2_U2695 );
nand NAND2_25618 ( P2_R2182_U290 , P2_R2182_U27 , P2_R2182_U16 );
nand NAND2_25619 ( P2_R2182_U291 , P2_R2182_U147 , P2_U2696 );
nand NAND2_25620 ( P2_R2182_U292 , P2_R2182_U25 , P2_R2182_U15 );
nand NAND2_25621 ( P2_R2182_U293 , P2_R2182_U146 , P2_U2666 );
nand NAND2_25622 ( P2_R2182_U294 , P2_R2182_U26 , P2_R2182_U14 );
nand NAND2_25623 ( P2_R2182_U295 , P2_R2182_U145 , P2_U2667 );
nand NAND2_25624 ( P2_R2182_U296 , P2_R2182_U38 , P2_R2182_U6 );
nand NAND2_25625 ( P2_R2182_U297 , P2_R2182_U144 , P2_U2668 );
nand NAND2_25626 ( P2_R2182_U298 , P2_R2182_U39 , P2_R2182_U5 );
nand NAND2_25627 ( P2_R2182_U299 , P2_R2182_U143 , P2_U2669 );
nand NAND2_25628 ( P2_R2182_U300 , P2_R2182_U33 , P2_R2182_U4 );
nand NAND2_25629 ( P2_R2182_U301 , P2_R2182_U142 , P2_U2670 );
nand NAND2_25630 ( P2_R2182_U302 , P2_R2182_U23 , P2_R2182_U20 );
nand NAND2_25631 ( P2_R2182_U303 , P2_R2182_U141 , P2_U2671 );
nand NAND2_25632 ( P2_R2182_U304 , P2_U2681 , P2_R2182_U44 );
nand NAND2_25633 ( P2_R2182_U305 , P2_U2702 , P2_R2182_U45 );
nand NAND3_25634 ( P2_R2167_U6 , P2_R2167_U42 , P2_R2167_U41 , P2_R2167_U38 );
not NOT1_25635 ( P2_R2167_U7 , P2_U2706 );
not NOT1_25636 ( P2_R2167_U8 , P2_U2713 );
not NOT1_25637 ( P2_R2167_U9 , P2_U2712 );
not NOT1_25638 ( P2_R2167_U10 , P2_U2705 );
not NOT1_25639 ( P2_R2167_U11 , P2_U2704 );
not NOT1_25640 ( P2_R2167_U12 , P2_U2711 );
not NOT1_25641 ( P2_R2167_U13 , P2_U2710 );
not NOT1_25642 ( P2_R2167_U14 , P2_U2703 );
not NOT1_25643 ( P2_R2167_U15 , P2_U2361 );
not NOT1_25644 ( P2_R2167_U16 , P2_U2709 );
not NOT1_25645 ( P2_R2167_U17 , P2_STATE2_REG_0_ );
not NOT1_25646 ( P2_R2167_U18 , P2_U2708 );
nand NAND2_25647 ( P2_R2167_U19 , P2_U2714 , P2_U2715 );
nand NAND2_25648 ( P2_R2167_U20 , P2_U2707 , P2_R2167_U19 );
or OR2_25649 ( P2_R2167_U21 , P2_U2714 , P2_U2715 );
nand NAND2_25650 ( P2_R2167_U22 , P2_U2706 , P2_R2167_U8 );
nand NAND3_25651 ( P2_R2167_U23 , P2_R2167_U21 , P2_R2167_U20 , P2_R2167_U22 );
nand NAND2_25652 ( P2_R2167_U24 , P2_U2713 , P2_R2167_U7 );
nand NAND2_25653 ( P2_R2167_U25 , P2_U2712 , P2_R2167_U10 );
nand NAND3_25654 ( P2_R2167_U26 , P2_R2167_U24 , P2_R2167_U25 , P2_R2167_U23 );
nand NAND2_25655 ( P2_R2167_U27 , P2_U2705 , P2_R2167_U9 );
nand NAND2_25656 ( P2_R2167_U28 , P2_U2704 , P2_R2167_U12 );
nand NAND3_25657 ( P2_R2167_U29 , P2_R2167_U27 , P2_R2167_U28 , P2_R2167_U26 );
nand NAND2_25658 ( P2_R2167_U30 , P2_U2711 , P2_R2167_U11 );
nand NAND2_25659 ( P2_R2167_U31 , P2_U2710 , P2_R2167_U14 );
nand NAND3_25660 ( P2_R2167_U32 , P2_R2167_U30 , P2_R2167_U29 , P2_R2167_U31 );
nand NAND2_25661 ( P2_R2167_U33 , P2_U2703 , P2_R2167_U13 );
nand NAND2_25662 ( P2_R2167_U34 , P2_U2361 , P2_R2167_U16 );
nand NAND3_25663 ( P2_R2167_U35 , P2_R2167_U33 , P2_R2167_U32 , P2_R2167_U34 );
nand NAND2_25664 ( P2_R2167_U36 , P2_U2709 , P2_R2167_U15 );
nand NAND2_25665 ( P2_R2167_U37 , P2_R2167_U36 , P2_R2167_U35 );
nand NAND3_25666 ( P2_R2167_U38 , P2_R2167_U40 , P2_R2167_U39 , P2_R2167_U37 );
nand NAND2_25667 ( P2_R2167_U39 , P2_U2361 , P2_R2167_U18 );
nand NAND2_25668 ( P2_R2167_U40 , P2_U2708 , P2_R2167_U15 );
nand NAND3_25669 ( P2_R2167_U41 , P2_STATE2_REG_0_ , P2_U2361 , P2_R2167_U18 );
nand NAND3_25670 ( P2_R2167_U42 , P2_R2167_U17 , P2_R2167_U15 , P2_U2708 );
not NOT1_25671 ( P2_R2027_U5 , P2_INSTADDRPOINTER_REG_0_ );
not NOT1_25672 ( P2_R2027_U6 , P2_INSTADDRPOINTER_REG_1_ );
nand NAND2_25673 ( P2_R2027_U7 , P2_INSTADDRPOINTER_REG_1_ , P2_INSTADDRPOINTER_REG_0_ );
not NOT1_25674 ( P2_R2027_U8 , P2_INSTADDRPOINTER_REG_2_ );
nand NAND2_25675 ( P2_R2027_U9 , P2_INSTADDRPOINTER_REG_2_ , P2_R2027_U98 );
not NOT1_25676 ( P2_R2027_U10 , P2_INSTADDRPOINTER_REG_3_ );
nand NAND2_25677 ( P2_R2027_U11 , P2_INSTADDRPOINTER_REG_3_ , P2_R2027_U99 );
not NOT1_25678 ( P2_R2027_U12 , P2_INSTADDRPOINTER_REG_4_ );
nand NAND2_25679 ( P2_R2027_U13 , P2_INSTADDRPOINTER_REG_4_ , P2_R2027_U100 );
not NOT1_25680 ( P2_R2027_U14 , P2_INSTADDRPOINTER_REG_5_ );
nand NAND2_25681 ( P2_R2027_U15 , P2_INSTADDRPOINTER_REG_5_ , P2_R2027_U101 );
not NOT1_25682 ( P2_R2027_U16 , P2_INSTADDRPOINTER_REG_6_ );
nand NAND2_25683 ( P2_R2027_U17 , P2_INSTADDRPOINTER_REG_6_ , P2_R2027_U102 );
not NOT1_25684 ( P2_R2027_U18 , P2_INSTADDRPOINTER_REG_7_ );
nand NAND2_25685 ( P2_R2027_U19 , P2_INSTADDRPOINTER_REG_7_ , P2_R2027_U103 );
not NOT1_25686 ( P2_R2027_U20 , P2_INSTADDRPOINTER_REG_8_ );
not NOT1_25687 ( P2_R2027_U21 , P2_INSTADDRPOINTER_REG_9_ );
nand NAND2_25688 ( P2_R2027_U22 , P2_INSTADDRPOINTER_REG_8_ , P2_R2027_U104 );
nand NAND2_25689 ( P2_R2027_U23 , P2_R2027_U105 , P2_INSTADDRPOINTER_REG_9_ );
not NOT1_25690 ( P2_R2027_U24 , P2_INSTADDRPOINTER_REG_10_ );
nand NAND2_25691 ( P2_R2027_U25 , P2_INSTADDRPOINTER_REG_10_ , P2_R2027_U106 );
not NOT1_25692 ( P2_R2027_U26 , P2_INSTADDRPOINTER_REG_11_ );
nand NAND2_25693 ( P2_R2027_U27 , P2_INSTADDRPOINTER_REG_11_ , P2_R2027_U107 );
not NOT1_25694 ( P2_R2027_U28 , P2_INSTADDRPOINTER_REG_12_ );
nand NAND2_25695 ( P2_R2027_U29 , P2_INSTADDRPOINTER_REG_12_ , P2_R2027_U108 );
not NOT1_25696 ( P2_R2027_U30 , P2_INSTADDRPOINTER_REG_13_ );
nand NAND2_25697 ( P2_R2027_U31 , P2_INSTADDRPOINTER_REG_13_ , P2_R2027_U109 );
not NOT1_25698 ( P2_R2027_U32 , P2_INSTADDRPOINTER_REG_14_ );
nand NAND2_25699 ( P2_R2027_U33 , P2_INSTADDRPOINTER_REG_14_ , P2_R2027_U110 );
not NOT1_25700 ( P2_R2027_U34 , P2_INSTADDRPOINTER_REG_15_ );
nand NAND2_25701 ( P2_R2027_U35 , P2_INSTADDRPOINTER_REG_15_ , P2_R2027_U111 );
not NOT1_25702 ( P2_R2027_U36 , P2_INSTADDRPOINTER_REG_16_ );
nand NAND2_25703 ( P2_R2027_U37 , P2_INSTADDRPOINTER_REG_16_ , P2_R2027_U112 );
not NOT1_25704 ( P2_R2027_U38 , P2_INSTADDRPOINTER_REG_17_ );
nand NAND2_25705 ( P2_R2027_U39 , P2_INSTADDRPOINTER_REG_17_ , P2_R2027_U113 );
not NOT1_25706 ( P2_R2027_U40 , P2_INSTADDRPOINTER_REG_18_ );
nand NAND2_25707 ( P2_R2027_U41 , P2_INSTADDRPOINTER_REG_18_ , P2_R2027_U114 );
not NOT1_25708 ( P2_R2027_U42 , P2_INSTADDRPOINTER_REG_19_ );
nand NAND2_25709 ( P2_R2027_U43 , P2_INSTADDRPOINTER_REG_19_ , P2_R2027_U115 );
not NOT1_25710 ( P2_R2027_U44 , P2_INSTADDRPOINTER_REG_20_ );
nand NAND2_25711 ( P2_R2027_U45 , P2_INSTADDRPOINTER_REG_20_ , P2_R2027_U116 );
not NOT1_25712 ( P2_R2027_U46 , P2_INSTADDRPOINTER_REG_21_ );
nand NAND2_25713 ( P2_R2027_U47 , P2_INSTADDRPOINTER_REG_21_ , P2_R2027_U117 );
not NOT1_25714 ( P2_R2027_U48 , P2_INSTADDRPOINTER_REG_22_ );
nand NAND2_25715 ( P2_R2027_U49 , P2_INSTADDRPOINTER_REG_22_ , P2_R2027_U118 );
not NOT1_25716 ( P2_R2027_U50 , P2_INSTADDRPOINTER_REG_23_ );
nand NAND2_25717 ( P2_R2027_U51 , P2_INSTADDRPOINTER_REG_23_ , P2_R2027_U119 );
not NOT1_25718 ( P2_R2027_U52 , P2_INSTADDRPOINTER_REG_24_ );
nand NAND2_25719 ( P2_R2027_U53 , P2_INSTADDRPOINTER_REG_24_ , P2_R2027_U120 );
not NOT1_25720 ( P2_R2027_U54 , P2_INSTADDRPOINTER_REG_25_ );
nand NAND2_25721 ( P2_R2027_U55 , P2_INSTADDRPOINTER_REG_25_ , P2_R2027_U121 );
not NOT1_25722 ( P2_R2027_U56 , P2_INSTADDRPOINTER_REG_26_ );
nand NAND2_25723 ( P2_R2027_U57 , P2_INSTADDRPOINTER_REG_26_ , P2_R2027_U122 );
not NOT1_25724 ( P2_R2027_U58 , P2_INSTADDRPOINTER_REG_27_ );
nand NAND2_25725 ( P2_R2027_U59 , P2_INSTADDRPOINTER_REG_27_ , P2_R2027_U123 );
not NOT1_25726 ( P2_R2027_U60 , P2_INSTADDRPOINTER_REG_28_ );
nand NAND2_25727 ( P2_R2027_U61 , P2_INSTADDRPOINTER_REG_28_ , P2_R2027_U124 );
not NOT1_25728 ( P2_R2027_U62 , P2_INSTADDRPOINTER_REG_29_ );
nand NAND2_25729 ( P2_R2027_U63 , P2_INSTADDRPOINTER_REG_29_ , P2_R2027_U125 );
not NOT1_25730 ( P2_R2027_U64 , P2_INSTADDRPOINTER_REG_30_ );
nand NAND2_25731 ( P2_R2027_U65 , P2_R2027_U129 , P2_R2027_U128 );
nand NAND2_25732 ( P2_R2027_U66 , P2_R2027_U131 , P2_R2027_U130 );
nand NAND2_25733 ( P2_R2027_U67 , P2_R2027_U133 , P2_R2027_U132 );
nand NAND2_25734 ( P2_R2027_U68 , P2_R2027_U135 , P2_R2027_U134 );
nand NAND2_25735 ( P2_R2027_U69 , P2_R2027_U137 , P2_R2027_U136 );
nand NAND2_25736 ( P2_R2027_U70 , P2_R2027_U139 , P2_R2027_U138 );
nand NAND2_25737 ( P2_R2027_U71 , P2_R2027_U141 , P2_R2027_U140 );
nand NAND2_25738 ( P2_R2027_U72 , P2_R2027_U143 , P2_R2027_U142 );
nand NAND2_25739 ( P2_R2027_U73 , P2_R2027_U145 , P2_R2027_U144 );
nand NAND2_25740 ( P2_R2027_U74 , P2_R2027_U147 , P2_R2027_U146 );
nand NAND2_25741 ( P2_R2027_U75 , P2_R2027_U149 , P2_R2027_U148 );
nand NAND2_25742 ( P2_R2027_U76 , P2_R2027_U151 , P2_R2027_U150 );
nand NAND2_25743 ( P2_R2027_U77 , P2_R2027_U153 , P2_R2027_U152 );
nand NAND2_25744 ( P2_R2027_U78 , P2_R2027_U155 , P2_R2027_U154 );
nand NAND2_25745 ( P2_R2027_U79 , P2_R2027_U157 , P2_R2027_U156 );
nand NAND2_25746 ( P2_R2027_U80 , P2_R2027_U159 , P2_R2027_U158 );
nand NAND2_25747 ( P2_R2027_U81 , P2_R2027_U161 , P2_R2027_U160 );
nand NAND2_25748 ( P2_R2027_U82 , P2_R2027_U163 , P2_R2027_U162 );
nand NAND2_25749 ( P2_R2027_U83 , P2_R2027_U165 , P2_R2027_U164 );
nand NAND2_25750 ( P2_R2027_U84 , P2_R2027_U167 , P2_R2027_U166 );
nand NAND2_25751 ( P2_R2027_U85 , P2_R2027_U169 , P2_R2027_U168 );
nand NAND2_25752 ( P2_R2027_U86 , P2_R2027_U171 , P2_R2027_U170 );
nand NAND2_25753 ( P2_R2027_U87 , P2_R2027_U173 , P2_R2027_U172 );
nand NAND2_25754 ( P2_R2027_U88 , P2_R2027_U175 , P2_R2027_U174 );
nand NAND2_25755 ( P2_R2027_U89 , P2_R2027_U177 , P2_R2027_U176 );
nand NAND2_25756 ( P2_R2027_U90 , P2_R2027_U179 , P2_R2027_U178 );
nand NAND2_25757 ( P2_R2027_U91 , P2_R2027_U181 , P2_R2027_U180 );
nand NAND2_25758 ( P2_R2027_U92 , P2_R2027_U183 , P2_R2027_U182 );
nand NAND2_25759 ( P2_R2027_U93 , P2_R2027_U185 , P2_R2027_U184 );
nand NAND2_25760 ( P2_R2027_U94 , P2_R2027_U187 , P2_R2027_U186 );
nand NAND2_25761 ( P2_R2027_U95 , P2_R2027_U189 , P2_R2027_U188 );
not NOT1_25762 ( P2_R2027_U96 , P2_INSTADDRPOINTER_REG_31_ );
nand NAND2_25763 ( P2_R2027_U97 , P2_INSTADDRPOINTER_REG_30_ , P2_R2027_U126 );
not NOT1_25764 ( P2_R2027_U98 , P2_R2027_U7 );
not NOT1_25765 ( P2_R2027_U99 , P2_R2027_U9 );
not NOT1_25766 ( P2_R2027_U100 , P2_R2027_U11 );
not NOT1_25767 ( P2_R2027_U101 , P2_R2027_U13 );
not NOT1_25768 ( P2_R2027_U102 , P2_R2027_U15 );
not NOT1_25769 ( P2_R2027_U103 , P2_R2027_U17 );
not NOT1_25770 ( P2_R2027_U104 , P2_R2027_U19 );
not NOT1_25771 ( P2_R2027_U105 , P2_R2027_U22 );
not NOT1_25772 ( P2_R2027_U106 , P2_R2027_U23 );
not NOT1_25773 ( P2_R2027_U107 , P2_R2027_U25 );
not NOT1_25774 ( P2_R2027_U108 , P2_R2027_U27 );
not NOT1_25775 ( P2_R2027_U109 , P2_R2027_U29 );
not NOT1_25776 ( P2_R2027_U110 , P2_R2027_U31 );
not NOT1_25777 ( P2_R2027_U111 , P2_R2027_U33 );
not NOT1_25778 ( P2_R2027_U112 , P2_R2027_U35 );
not NOT1_25779 ( P2_R2027_U113 , P2_R2027_U37 );
not NOT1_25780 ( P2_R2027_U114 , P2_R2027_U39 );
not NOT1_25781 ( P2_R2027_U115 , P2_R2027_U41 );
not NOT1_25782 ( P2_R2027_U116 , P2_R2027_U43 );
not NOT1_25783 ( P2_R2027_U117 , P2_R2027_U45 );
not NOT1_25784 ( P2_R2027_U118 , P2_R2027_U47 );
not NOT1_25785 ( P2_R2027_U119 , P2_R2027_U49 );
not NOT1_25786 ( P2_R2027_U120 , P2_R2027_U51 );
not NOT1_25787 ( P2_R2027_U121 , P2_R2027_U53 );
not NOT1_25788 ( P2_R2027_U122 , P2_R2027_U55 );
not NOT1_25789 ( P2_R2027_U123 , P2_R2027_U57 );
not NOT1_25790 ( P2_R2027_U124 , P2_R2027_U59 );
not NOT1_25791 ( P2_R2027_U125 , P2_R2027_U61 );
not NOT1_25792 ( P2_R2027_U126 , P2_R2027_U63 );
not NOT1_25793 ( P2_R2027_U127 , P2_R2027_U97 );
nand NAND2_25794 ( P2_R2027_U128 , P2_INSTADDRPOINTER_REG_9_ , P2_R2027_U22 );
nand NAND2_25795 ( P2_R2027_U129 , P2_R2027_U105 , P2_R2027_U21 );
nand NAND2_25796 ( P2_R2027_U130 , P2_INSTADDRPOINTER_REG_8_ , P2_R2027_U19 );
nand NAND2_25797 ( P2_R2027_U131 , P2_R2027_U104 , P2_R2027_U20 );
nand NAND2_25798 ( P2_R2027_U132 , P2_INSTADDRPOINTER_REG_7_ , P2_R2027_U17 );
nand NAND2_25799 ( P2_R2027_U133 , P2_R2027_U103 , P2_R2027_U18 );
nand NAND2_25800 ( P2_R2027_U134 , P2_INSTADDRPOINTER_REG_6_ , P2_R2027_U15 );
nand NAND2_25801 ( P2_R2027_U135 , P2_R2027_U102 , P2_R2027_U16 );
nand NAND2_25802 ( P2_R2027_U136 , P2_INSTADDRPOINTER_REG_5_ , P2_R2027_U13 );
nand NAND2_25803 ( P2_R2027_U137 , P2_R2027_U101 , P2_R2027_U14 );
nand NAND2_25804 ( P2_R2027_U138 , P2_INSTADDRPOINTER_REG_4_ , P2_R2027_U11 );
nand NAND2_25805 ( P2_R2027_U139 , P2_R2027_U100 , P2_R2027_U12 );
nand NAND2_25806 ( P2_R2027_U140 , P2_INSTADDRPOINTER_REG_3_ , P2_R2027_U9 );
nand NAND2_25807 ( P2_R2027_U141 , P2_R2027_U99 , P2_R2027_U10 );
nand NAND2_25808 ( P2_R2027_U142 , P2_INSTADDRPOINTER_REG_31_ , P2_R2027_U97 );
nand NAND2_25809 ( P2_R2027_U143 , P2_R2027_U127 , P2_R2027_U96 );
nand NAND2_25810 ( P2_R2027_U144 , P2_INSTADDRPOINTER_REG_30_ , P2_R2027_U63 );
nand NAND2_25811 ( P2_R2027_U145 , P2_R2027_U126 , P2_R2027_U64 );
nand NAND2_25812 ( P2_R2027_U146 , P2_INSTADDRPOINTER_REG_2_ , P2_R2027_U7 );
nand NAND2_25813 ( P2_R2027_U147 , P2_R2027_U98 , P2_R2027_U8 );
nand NAND2_25814 ( P2_R2027_U148 , P2_INSTADDRPOINTER_REG_29_ , P2_R2027_U61 );
nand NAND2_25815 ( P2_R2027_U149 , P2_R2027_U125 , P2_R2027_U62 );
nand NAND2_25816 ( P2_R2027_U150 , P2_INSTADDRPOINTER_REG_28_ , P2_R2027_U59 );
nand NAND2_25817 ( P2_R2027_U151 , P2_R2027_U124 , P2_R2027_U60 );
nand NAND2_25818 ( P2_R2027_U152 , P2_INSTADDRPOINTER_REG_27_ , P2_R2027_U57 );
nand NAND2_25819 ( P2_R2027_U153 , P2_R2027_U123 , P2_R2027_U58 );
nand NAND2_25820 ( P2_R2027_U154 , P2_INSTADDRPOINTER_REG_26_ , P2_R2027_U55 );
nand NAND2_25821 ( P2_R2027_U155 , P2_R2027_U122 , P2_R2027_U56 );
nand NAND2_25822 ( P2_R2027_U156 , P2_INSTADDRPOINTER_REG_25_ , P2_R2027_U53 );
nand NAND2_25823 ( P2_R2027_U157 , P2_R2027_U121 , P2_R2027_U54 );
nand NAND2_25824 ( P2_R2027_U158 , P2_INSTADDRPOINTER_REG_24_ , P2_R2027_U51 );
nand NAND2_25825 ( P2_R2027_U159 , P2_R2027_U120 , P2_R2027_U52 );
nand NAND2_25826 ( P2_R2027_U160 , P2_INSTADDRPOINTER_REG_23_ , P2_R2027_U49 );
nand NAND2_25827 ( P2_R2027_U161 , P2_R2027_U119 , P2_R2027_U50 );
nand NAND2_25828 ( P2_R2027_U162 , P2_INSTADDRPOINTER_REG_22_ , P2_R2027_U47 );
nand NAND2_25829 ( P2_R2027_U163 , P2_R2027_U118 , P2_R2027_U48 );
nand NAND2_25830 ( P2_R2027_U164 , P2_INSTADDRPOINTER_REG_21_ , P2_R2027_U45 );
nand NAND2_25831 ( P2_R2027_U165 , P2_R2027_U117 , P2_R2027_U46 );
nand NAND2_25832 ( P2_R2027_U166 , P2_INSTADDRPOINTER_REG_20_ , P2_R2027_U43 );
nand NAND2_25833 ( P2_R2027_U167 , P2_R2027_U116 , P2_R2027_U44 );
nand NAND2_25834 ( P2_R2027_U168 , P2_INSTADDRPOINTER_REG_1_ , P2_R2027_U5 );
nand NAND2_25835 ( P2_R2027_U169 , P2_INSTADDRPOINTER_REG_0_ , P2_R2027_U6 );
nand NAND2_25836 ( P2_R2027_U170 , P2_INSTADDRPOINTER_REG_19_ , P2_R2027_U41 );
nand NAND2_25837 ( P2_R2027_U171 , P2_R2027_U115 , P2_R2027_U42 );
nand NAND2_25838 ( P2_R2027_U172 , P2_INSTADDRPOINTER_REG_18_ , P2_R2027_U39 );
nand NAND2_25839 ( P2_R2027_U173 , P2_R2027_U114 , P2_R2027_U40 );
nand NAND2_25840 ( P2_R2027_U174 , P2_INSTADDRPOINTER_REG_17_ , P2_R2027_U37 );
nand NAND2_25841 ( P2_R2027_U175 , P2_R2027_U113 , P2_R2027_U38 );
nand NAND2_25842 ( P2_R2027_U176 , P2_INSTADDRPOINTER_REG_16_ , P2_R2027_U35 );
nand NAND2_25843 ( P2_R2027_U177 , P2_R2027_U112 , P2_R2027_U36 );
nand NAND2_25844 ( P2_R2027_U178 , P2_INSTADDRPOINTER_REG_15_ , P2_R2027_U33 );
nand NAND2_25845 ( P2_R2027_U179 , P2_R2027_U111 , P2_R2027_U34 );
nand NAND2_25846 ( P2_R2027_U180 , P2_INSTADDRPOINTER_REG_14_ , P2_R2027_U31 );
nand NAND2_25847 ( P2_R2027_U181 , P2_R2027_U110 , P2_R2027_U32 );
nand NAND2_25848 ( P2_R2027_U182 , P2_INSTADDRPOINTER_REG_13_ , P2_R2027_U29 );
nand NAND2_25849 ( P2_R2027_U183 , P2_R2027_U109 , P2_R2027_U30 );
nand NAND2_25850 ( P2_R2027_U184 , P2_INSTADDRPOINTER_REG_12_ , P2_R2027_U27 );
nand NAND2_25851 ( P2_R2027_U185 , P2_R2027_U108 , P2_R2027_U28 );
nand NAND2_25852 ( P2_R2027_U186 , P2_INSTADDRPOINTER_REG_11_ , P2_R2027_U25 );
nand NAND2_25853 ( P2_R2027_U187 , P2_R2027_U107 , P2_R2027_U26 );
nand NAND2_25854 ( P2_R2027_U188 , P2_INSTADDRPOINTER_REG_10_ , P2_R2027_U23 );
nand NAND2_25855 ( P2_R2027_U189 , P2_R2027_U106 , P2_R2027_U24 );
or OR2_25856 ( P2_LT_563_1260_U6 , P2_LT_563_1260_U7 , P2_U3617 );
nor nor_25857 ( P2_LT_563_1260_U7 , P2_SUB_563_U6 , P2_SUB_563_U7 );
not NOT1_25858 ( P2_R2337_U4 , P2_PHYADDRPOINTER_REG_1_ );
not NOT1_25859 ( P2_R2337_U5 , P2_PHYADDRPOINTER_REG_3_ );
not NOT1_25860 ( P2_R2337_U6 , P2_PHYADDRPOINTER_REG_2_ );
nand NAND3_25861 ( P2_R2337_U7 , P2_PHYADDRPOINTER_REG_3_ , P2_PHYADDRPOINTER_REG_1_ , P2_PHYADDRPOINTER_REG_2_ );
not NOT1_25862 ( P2_R2337_U8 , P2_PHYADDRPOINTER_REG_4_ );
nand NAND2_25863 ( P2_R2337_U9 , P2_PHYADDRPOINTER_REG_4_ , P2_R2337_U95 );
not NOT1_25864 ( P2_R2337_U10 , P2_PHYADDRPOINTER_REG_5_ );
nand NAND2_25865 ( P2_R2337_U11 , P2_PHYADDRPOINTER_REG_5_ , P2_R2337_U96 );
not NOT1_25866 ( P2_R2337_U12 , P2_PHYADDRPOINTER_REG_6_ );
nand NAND2_25867 ( P2_R2337_U13 , P2_PHYADDRPOINTER_REG_6_ , P2_R2337_U97 );
not NOT1_25868 ( P2_R2337_U14 , P2_PHYADDRPOINTER_REG_7_ );
nand NAND2_25869 ( P2_R2337_U15 , P2_PHYADDRPOINTER_REG_7_ , P2_R2337_U98 );
not NOT1_25870 ( P2_R2337_U16 , P2_PHYADDRPOINTER_REG_8_ );
not NOT1_25871 ( P2_R2337_U17 , P2_PHYADDRPOINTER_REG_9_ );
nand NAND2_25872 ( P2_R2337_U18 , P2_PHYADDRPOINTER_REG_8_ , P2_R2337_U99 );
nand NAND2_25873 ( P2_R2337_U19 , P2_R2337_U100 , P2_PHYADDRPOINTER_REG_9_ );
not NOT1_25874 ( P2_R2337_U20 , P2_PHYADDRPOINTER_REG_10_ );
nand NAND2_25875 ( P2_R2337_U21 , P2_PHYADDRPOINTER_REG_10_ , P2_R2337_U101 );
not NOT1_25876 ( P2_R2337_U22 , P2_PHYADDRPOINTER_REG_11_ );
nand NAND2_25877 ( P2_R2337_U23 , P2_PHYADDRPOINTER_REG_11_ , P2_R2337_U102 );
not NOT1_25878 ( P2_R2337_U24 , P2_PHYADDRPOINTER_REG_12_ );
nand NAND2_25879 ( P2_R2337_U25 , P2_PHYADDRPOINTER_REG_12_ , P2_R2337_U103 );
not NOT1_25880 ( P2_R2337_U26 , P2_PHYADDRPOINTER_REG_13_ );
nand NAND2_25881 ( P2_R2337_U27 , P2_PHYADDRPOINTER_REG_13_ , P2_R2337_U104 );
not NOT1_25882 ( P2_R2337_U28 , P2_PHYADDRPOINTER_REG_14_ );
nand NAND2_25883 ( P2_R2337_U29 , P2_PHYADDRPOINTER_REG_14_ , P2_R2337_U105 );
not NOT1_25884 ( P2_R2337_U30 , P2_PHYADDRPOINTER_REG_15_ );
nand NAND2_25885 ( P2_R2337_U31 , P2_PHYADDRPOINTER_REG_15_ , P2_R2337_U106 );
not NOT1_25886 ( P2_R2337_U32 , P2_PHYADDRPOINTER_REG_16_ );
nand NAND2_25887 ( P2_R2337_U33 , P2_PHYADDRPOINTER_REG_16_ , P2_R2337_U107 );
not NOT1_25888 ( P2_R2337_U34 , P2_PHYADDRPOINTER_REG_17_ );
nand NAND2_25889 ( P2_R2337_U35 , P2_PHYADDRPOINTER_REG_17_ , P2_R2337_U108 );
not NOT1_25890 ( P2_R2337_U36 , P2_PHYADDRPOINTER_REG_18_ );
nand NAND2_25891 ( P2_R2337_U37 , P2_PHYADDRPOINTER_REG_18_ , P2_R2337_U109 );
not NOT1_25892 ( P2_R2337_U38 , P2_PHYADDRPOINTER_REG_19_ );
nand NAND2_25893 ( P2_R2337_U39 , P2_PHYADDRPOINTER_REG_19_ , P2_R2337_U110 );
not NOT1_25894 ( P2_R2337_U40 , P2_PHYADDRPOINTER_REG_20_ );
nand NAND2_25895 ( P2_R2337_U41 , P2_PHYADDRPOINTER_REG_20_ , P2_R2337_U111 );
not NOT1_25896 ( P2_R2337_U42 , P2_PHYADDRPOINTER_REG_21_ );
nand NAND2_25897 ( P2_R2337_U43 , P2_PHYADDRPOINTER_REG_21_ , P2_R2337_U112 );
not NOT1_25898 ( P2_R2337_U44 , P2_PHYADDRPOINTER_REG_22_ );
nand NAND2_25899 ( P2_R2337_U45 , P2_PHYADDRPOINTER_REG_22_ , P2_R2337_U113 );
not NOT1_25900 ( P2_R2337_U46 , P2_PHYADDRPOINTER_REG_23_ );
nand NAND2_25901 ( P2_R2337_U47 , P2_PHYADDRPOINTER_REG_23_ , P2_R2337_U114 );
not NOT1_25902 ( P2_R2337_U48 , P2_PHYADDRPOINTER_REG_24_ );
nand NAND2_25903 ( P2_R2337_U49 , P2_PHYADDRPOINTER_REG_24_ , P2_R2337_U115 );
not NOT1_25904 ( P2_R2337_U50 , P2_PHYADDRPOINTER_REG_25_ );
nand NAND2_25905 ( P2_R2337_U51 , P2_PHYADDRPOINTER_REG_25_ , P2_R2337_U116 );
not NOT1_25906 ( P2_R2337_U52 , P2_PHYADDRPOINTER_REG_26_ );
nand NAND2_25907 ( P2_R2337_U53 , P2_PHYADDRPOINTER_REG_26_ , P2_R2337_U117 );
not NOT1_25908 ( P2_R2337_U54 , P2_PHYADDRPOINTER_REG_27_ );
nand NAND2_25909 ( P2_R2337_U55 , P2_PHYADDRPOINTER_REG_27_ , P2_R2337_U118 );
not NOT1_25910 ( P2_R2337_U56 , P2_PHYADDRPOINTER_REG_28_ );
nand NAND2_25911 ( P2_R2337_U57 , P2_PHYADDRPOINTER_REG_28_ , P2_R2337_U119 );
not NOT1_25912 ( P2_R2337_U58 , P2_PHYADDRPOINTER_REG_29_ );
nand NAND2_25913 ( P2_R2337_U59 , P2_PHYADDRPOINTER_REG_29_ , P2_R2337_U120 );
not NOT1_25914 ( P2_R2337_U60 , P2_PHYADDRPOINTER_REG_30_ );
nand NAND2_25915 ( P2_R2337_U61 , P2_R2337_U124 , P2_R2337_U123 );
nand NAND2_25916 ( P2_R2337_U62 , P2_R2337_U126 , P2_R2337_U125 );
nand NAND2_25917 ( P2_R2337_U63 , P2_R2337_U128 , P2_R2337_U127 );
nand NAND2_25918 ( P2_R2337_U64 , P2_R2337_U130 , P2_R2337_U129 );
nand NAND2_25919 ( P2_R2337_U65 , P2_R2337_U132 , P2_R2337_U131 );
nand NAND2_25920 ( P2_R2337_U66 , P2_R2337_U134 , P2_R2337_U133 );
nand NAND2_25921 ( P2_R2337_U67 , P2_R2337_U136 , P2_R2337_U135 );
nand NAND2_25922 ( P2_R2337_U68 , P2_R2337_U138 , P2_R2337_U137 );
nand NAND2_25923 ( P2_R2337_U69 , P2_R2337_U140 , P2_R2337_U139 );
nand NAND2_25924 ( P2_R2337_U70 , P2_R2337_U142 , P2_R2337_U141 );
nand NAND2_25925 ( P2_R2337_U71 , P2_R2337_U144 , P2_R2337_U143 );
nand NAND2_25926 ( P2_R2337_U72 , P2_R2337_U146 , P2_R2337_U145 );
nand NAND2_25927 ( P2_R2337_U73 , P2_R2337_U148 , P2_R2337_U147 );
nand NAND2_25928 ( P2_R2337_U74 , P2_R2337_U150 , P2_R2337_U149 );
nand NAND2_25929 ( P2_R2337_U75 , P2_R2337_U152 , P2_R2337_U151 );
nand NAND2_25930 ( P2_R2337_U76 , P2_R2337_U154 , P2_R2337_U153 );
nand NAND2_25931 ( P2_R2337_U77 , P2_R2337_U156 , P2_R2337_U155 );
nand NAND2_25932 ( P2_R2337_U78 , P2_R2337_U158 , P2_R2337_U157 );
nand NAND2_25933 ( P2_R2337_U79 , P2_R2337_U160 , P2_R2337_U159 );
nand NAND2_25934 ( P2_R2337_U80 , P2_R2337_U162 , P2_R2337_U161 );
nand NAND2_25935 ( P2_R2337_U81 , P2_R2337_U164 , P2_R2337_U163 );
nand NAND2_25936 ( P2_R2337_U82 , P2_R2337_U166 , P2_R2337_U165 );
nand NAND2_25937 ( P2_R2337_U83 , P2_R2337_U168 , P2_R2337_U167 );
nand NAND2_25938 ( P2_R2337_U84 , P2_R2337_U170 , P2_R2337_U169 );
nand NAND2_25939 ( P2_R2337_U85 , P2_R2337_U172 , P2_R2337_U171 );
nand NAND2_25940 ( P2_R2337_U86 , P2_R2337_U174 , P2_R2337_U173 );
nand NAND2_25941 ( P2_R2337_U87 , P2_R2337_U176 , P2_R2337_U175 );
nand NAND2_25942 ( P2_R2337_U88 , P2_R2337_U178 , P2_R2337_U177 );
nand NAND2_25943 ( P2_R2337_U89 , P2_R2337_U180 , P2_R2337_U179 );
nand NAND2_25944 ( P2_R2337_U90 , P2_R2337_U182 , P2_R2337_U181 );
nand NAND2_25945 ( P2_R2337_U91 , P2_PHYADDRPOINTER_REG_2_ , P2_PHYADDRPOINTER_REG_1_ );
not NOT1_25946 ( P2_R2337_U92 , P2_PHYADDRPOINTER_REG_31_ );
nand NAND2_25947 ( P2_R2337_U93 , P2_PHYADDRPOINTER_REG_30_ , P2_R2337_U121 );
not NOT1_25948 ( P2_R2337_U94 , P2_R2337_U91 );
not NOT1_25949 ( P2_R2337_U95 , P2_R2337_U7 );
not NOT1_25950 ( P2_R2337_U96 , P2_R2337_U9 );
not NOT1_25951 ( P2_R2337_U97 , P2_R2337_U11 );
not NOT1_25952 ( P2_R2337_U98 , P2_R2337_U13 );
not NOT1_25953 ( P2_R2337_U99 , P2_R2337_U15 );
not NOT1_25954 ( P2_R2337_U100 , P2_R2337_U18 );
not NOT1_25955 ( P2_R2337_U101 , P2_R2337_U19 );
not NOT1_25956 ( P2_R2337_U102 , P2_R2337_U21 );
not NOT1_25957 ( P2_R2337_U103 , P2_R2337_U23 );
not NOT1_25958 ( P2_R2337_U104 , P2_R2337_U25 );
not NOT1_25959 ( P2_R2337_U105 , P2_R2337_U27 );
not NOT1_25960 ( P2_R2337_U106 , P2_R2337_U29 );
not NOT1_25961 ( P2_R2337_U107 , P2_R2337_U31 );
not NOT1_25962 ( P2_R2337_U108 , P2_R2337_U33 );
not NOT1_25963 ( P2_R2337_U109 , P2_R2337_U35 );
not NOT1_25964 ( P2_R2337_U110 , P2_R2337_U37 );
not NOT1_25965 ( P2_R2337_U111 , P2_R2337_U39 );
not NOT1_25966 ( P2_R2337_U112 , P2_R2337_U41 );
not NOT1_25967 ( P2_R2337_U113 , P2_R2337_U43 );
not NOT1_25968 ( P2_R2337_U114 , P2_R2337_U45 );
not NOT1_25969 ( P2_R2337_U115 , P2_R2337_U47 );
not NOT1_25970 ( P2_R2337_U116 , P2_R2337_U49 );
not NOT1_25971 ( P2_R2337_U117 , P2_R2337_U51 );
not NOT1_25972 ( P2_R2337_U118 , P2_R2337_U53 );
not NOT1_25973 ( P2_R2337_U119 , P2_R2337_U55 );
not NOT1_25974 ( P2_R2337_U120 , P2_R2337_U57 );
not NOT1_25975 ( P2_R2337_U121 , P2_R2337_U59 );
not NOT1_25976 ( P2_R2337_U122 , P2_R2337_U93 );
nand NAND2_25977 ( P2_R2337_U123 , P2_PHYADDRPOINTER_REG_9_ , P2_R2337_U18 );
nand NAND2_25978 ( P2_R2337_U124 , P2_R2337_U100 , P2_R2337_U17 );
nand NAND2_25979 ( P2_R2337_U125 , P2_PHYADDRPOINTER_REG_8_ , P2_R2337_U15 );
nand NAND2_25980 ( P2_R2337_U126 , P2_R2337_U99 , P2_R2337_U16 );
nand NAND2_25981 ( P2_R2337_U127 , P2_PHYADDRPOINTER_REG_7_ , P2_R2337_U13 );
nand NAND2_25982 ( P2_R2337_U128 , P2_R2337_U98 , P2_R2337_U14 );
nand NAND2_25983 ( P2_R2337_U129 , P2_PHYADDRPOINTER_REG_6_ , P2_R2337_U11 );
nand NAND2_25984 ( P2_R2337_U130 , P2_R2337_U97 , P2_R2337_U12 );
nand NAND2_25985 ( P2_R2337_U131 , P2_PHYADDRPOINTER_REG_5_ , P2_R2337_U9 );
nand NAND2_25986 ( P2_R2337_U132 , P2_R2337_U96 , P2_R2337_U10 );
nand NAND2_25987 ( P2_R2337_U133 , P2_PHYADDRPOINTER_REG_4_ , P2_R2337_U7 );
nand NAND2_25988 ( P2_R2337_U134 , P2_R2337_U95 , P2_R2337_U8 );
nand NAND2_25989 ( P2_R2337_U135 , P2_PHYADDRPOINTER_REG_3_ , P2_R2337_U91 );
nand NAND2_25990 ( P2_R2337_U136 , P2_R2337_U94 , P2_R2337_U5 );
nand NAND2_25991 ( P2_R2337_U137 , P2_PHYADDRPOINTER_REG_31_ , P2_R2337_U93 );
nand NAND2_25992 ( P2_R2337_U138 , P2_R2337_U122 , P2_R2337_U92 );
nand NAND2_25993 ( P2_R2337_U139 , P2_PHYADDRPOINTER_REG_30_ , P2_R2337_U59 );
nand NAND2_25994 ( P2_R2337_U140 , P2_R2337_U121 , P2_R2337_U60 );
nand NAND2_25995 ( P2_R2337_U141 , P2_PHYADDRPOINTER_REG_2_ , P2_R2337_U4 );
nand NAND2_25996 ( P2_R2337_U142 , P2_PHYADDRPOINTER_REG_1_ , P2_R2337_U6 );
nand NAND2_25997 ( P2_R2337_U143 , P2_PHYADDRPOINTER_REG_29_ , P2_R2337_U57 );
nand NAND2_25998 ( P2_R2337_U144 , P2_R2337_U120 , P2_R2337_U58 );
nand NAND2_25999 ( P2_R2337_U145 , P2_PHYADDRPOINTER_REG_28_ , P2_R2337_U55 );
nand NAND2_26000 ( P2_R2337_U146 , P2_R2337_U119 , P2_R2337_U56 );
nand NAND2_26001 ( P2_R2337_U147 , P2_PHYADDRPOINTER_REG_27_ , P2_R2337_U53 );
nand NAND2_26002 ( P2_R2337_U148 , P2_R2337_U118 , P2_R2337_U54 );
nand NAND2_26003 ( P2_R2337_U149 , P2_PHYADDRPOINTER_REG_26_ , P2_R2337_U51 );
nand NAND2_26004 ( P2_R2337_U150 , P2_R2337_U117 , P2_R2337_U52 );
nand NAND2_26005 ( P2_R2337_U151 , P2_PHYADDRPOINTER_REG_25_ , P2_R2337_U49 );
nand NAND2_26006 ( P2_R2337_U152 , P2_R2337_U116 , P2_R2337_U50 );
nand NAND2_26007 ( P2_R2337_U153 , P2_PHYADDRPOINTER_REG_24_ , P2_R2337_U47 );
nand NAND2_26008 ( P2_R2337_U154 , P2_R2337_U115 , P2_R2337_U48 );
nand NAND2_26009 ( P2_R2337_U155 , P2_PHYADDRPOINTER_REG_23_ , P2_R2337_U45 );
nand NAND2_26010 ( P2_R2337_U156 , P2_R2337_U114 , P2_R2337_U46 );
nand NAND2_26011 ( P2_R2337_U157 , P2_PHYADDRPOINTER_REG_22_ , P2_R2337_U43 );
nand NAND2_26012 ( P2_R2337_U158 , P2_R2337_U113 , P2_R2337_U44 );
nand NAND2_26013 ( P2_R2337_U159 , P2_PHYADDRPOINTER_REG_21_ , P2_R2337_U41 );
nand NAND2_26014 ( P2_R2337_U160 , P2_R2337_U112 , P2_R2337_U42 );
nand NAND2_26015 ( P2_R2337_U161 , P2_PHYADDRPOINTER_REG_20_ , P2_R2337_U39 );
nand NAND2_26016 ( P2_R2337_U162 , P2_R2337_U111 , P2_R2337_U40 );
nand NAND2_26017 ( P2_R2337_U163 , P2_PHYADDRPOINTER_REG_19_ , P2_R2337_U37 );
nand NAND2_26018 ( P2_R2337_U164 , P2_R2337_U110 , P2_R2337_U38 );
nand NAND2_26019 ( P2_R2337_U165 , P2_PHYADDRPOINTER_REG_18_ , P2_R2337_U35 );
nand NAND2_26020 ( P2_R2337_U166 , P2_R2337_U109 , P2_R2337_U36 );
nand NAND2_26021 ( P2_R2337_U167 , P2_PHYADDRPOINTER_REG_17_ , P2_R2337_U33 );
nand NAND2_26022 ( P2_R2337_U168 , P2_R2337_U108 , P2_R2337_U34 );
nand NAND2_26023 ( P2_R2337_U169 , P2_PHYADDRPOINTER_REG_16_ , P2_R2337_U31 );
nand NAND2_26024 ( P2_R2337_U170 , P2_R2337_U107 , P2_R2337_U32 );
nand NAND2_26025 ( P2_R2337_U171 , P2_PHYADDRPOINTER_REG_15_ , P2_R2337_U29 );
nand NAND2_26026 ( P2_R2337_U172 , P2_R2337_U106 , P2_R2337_U30 );
nand NAND2_26027 ( P2_R2337_U173 , P2_PHYADDRPOINTER_REG_14_ , P2_R2337_U27 );
nand NAND2_26028 ( P2_R2337_U174 , P2_R2337_U105 , P2_R2337_U28 );
nand NAND2_26029 ( P2_R2337_U175 , P2_PHYADDRPOINTER_REG_13_ , P2_R2337_U25 );
nand NAND2_26030 ( P2_R2337_U176 , P2_R2337_U104 , P2_R2337_U26 );
nand NAND2_26031 ( P2_R2337_U177 , P2_PHYADDRPOINTER_REG_12_ , P2_R2337_U23 );
nand NAND2_26032 ( P2_R2337_U178 , P2_R2337_U103 , P2_R2337_U24 );
nand NAND2_26033 ( P2_R2337_U179 , P2_PHYADDRPOINTER_REG_11_ , P2_R2337_U21 );
nand NAND2_26034 ( P2_R2337_U180 , P2_R2337_U102 , P2_R2337_U22 );
nand NAND2_26035 ( P2_R2337_U181 , P2_PHYADDRPOINTER_REG_10_ , P2_R2337_U19 );
nand NAND2_26036 ( P2_R2337_U182 , P2_R2337_U101 , P2_R2337_U20 );
not NOT1_26037 ( P2_R2147_U4 , P2_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_26038 ( P2_R2147_U5 , P2_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_26039 ( P2_R2147_U6 , P2_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_26040 ( P2_R2147_U7 , P2_R2147_U16 , P2_R2147_U15 );
nand NAND2_26041 ( P2_R2147_U8 , P2_R2147_U18 , P2_R2147_U17 );
nand NAND2_26042 ( P2_R2147_U9 , P2_R2147_U20 , P2_R2147_U19 );
not NOT1_26043 ( P2_R2147_U10 , P2_U2752 );
nand NAND3_26044 ( P2_R2147_U11 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_INSTQUEUERD_ADDR_REG_1_ , P2_INSTQUEUERD_ADDR_REG_2_ );
nand NAND2_26045 ( P2_R2147_U12 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_26046 ( P2_R2147_U13 , P2_R2147_U11 );
not NOT1_26047 ( P2_R2147_U14 , P2_R2147_U12 );
nand NAND2_26048 ( P2_R2147_U15 , P2_U2752 , P2_R2147_U11 );
nand NAND2_26049 ( P2_R2147_U16 , P2_R2147_U13 , P2_R2147_U10 );
nand NAND2_26050 ( P2_R2147_U17 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_R2147_U12 );
nand NAND2_26051 ( P2_R2147_U18 , P2_R2147_U14 , P2_R2147_U5 );
nand NAND2_26052 ( P2_R2147_U19 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_R2147_U4 );
nand NAND2_26053 ( P2_R2147_U20 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_R2147_U6 );
and AND2_26054 ( P2_R2219_U6 , P2_R2219_U52 , P2_R2219_U48 );
and AND2_26055 ( P2_R2219_U7 , P2_R2219_U68 , P2_R2219_U66 );
nand NAND2_26056 ( P2_R2219_U8 , P2_R2219_U45 , P2_R2219_U69 );
not NOT1_26057 ( P2_R2219_U9 , P2_U4428 );
not NOT1_26058 ( P2_R2219_U10 , P2_U2753 );
not NOT1_26059 ( P2_R2219_U11 , P2_U2761 );
not NOT1_26060 ( P2_R2219_U12 , P2_U2763 );
not NOT1_26061 ( P2_R2219_U13 , P2_U2762 );
not NOT1_26062 ( P2_R2219_U14 , P2_U2756 );
not NOT1_26063 ( P2_R2219_U15 , P2_U2765 );
not NOT1_26064 ( P2_R2219_U16 , P2_U2764 );
not NOT1_26065 ( P2_R2219_U17 , P2_U2755 );
not NOT1_26066 ( P2_R2219_U18 , P2_U2754 );
nand NAND2_26067 ( P2_R2219_U19 , P2_R2219_U72 , P2_R2219_U76 );
not NOT1_26068 ( P2_R2219_U20 , P2_U2760 );
not NOT1_26069 ( P2_R2219_U21 , P2_U2759 );
not NOT1_26070 ( P2_R2219_U22 , P2_U2758 );
not NOT1_26071 ( P2_R2219_U23 , P2_U2757 );
nand NAND2_26072 ( P2_R2219_U24 , P2_R2219_U86 , P2_R2219_U85 );
nand NAND2_26073 ( P2_R2219_U25 , P2_R2219_U91 , P2_R2219_U90 );
nand NAND2_26074 ( P2_R2219_U26 , P2_R2219_U96 , P2_R2219_U95 );
nand NAND2_26075 ( P2_R2219_U27 , P2_R2219_U101 , P2_R2219_U100 );
nand NAND2_26076 ( P2_R2219_U28 , P2_R2219_U106 , P2_R2219_U105 );
nand NAND2_26077 ( P2_R2219_U29 , P2_R2219_U111 , P2_R2219_U110 );
nand NAND2_26078 ( P2_R2219_U30 , P2_R2219_U116 , P2_R2219_U115 );
and AND2_26079 ( P2_R2219_U31 , P2_R2219_U6 , P2_R2219_U55 );
nand NAND2_26080 ( P2_R2219_U32 , P2_R2219_U83 , P2_R2219_U82 );
nand NAND2_26081 ( P2_R2219_U33 , P2_R2219_U88 , P2_R2219_U87 );
nand NAND2_26082 ( P2_R2219_U34 , P2_R2219_U93 , P2_R2219_U92 );
nand NAND2_26083 ( P2_R2219_U35 , P2_R2219_U98 , P2_R2219_U97 );
nand NAND2_26084 ( P2_R2219_U36 , P2_R2219_U103 , P2_R2219_U102 );
nand NAND2_26085 ( P2_R2219_U37 , P2_R2219_U108 , P2_R2219_U107 );
nand NAND2_26086 ( P2_R2219_U38 , P2_R2219_U113 , P2_R2219_U112 );
nand NAND2_26087 ( P2_R2219_U39 , P2_R2219_U64 , P2_R2219_U63 );
nand NAND2_26088 ( P2_R2219_U40 , P2_R2219_U60 , P2_R2219_U59 );
nand NAND3_26089 ( P2_R2219_U41 , P2_R2219_U75 , P2_R2219_U56 , P2_R2219_U74 );
nand NAND2_26090 ( P2_R2219_U42 , P2_R2219_U19 , P2_R2219_U71 );
nand NAND2_26091 ( P2_R2219_U43 , P2_R2219_U50 , P2_R2219_U49 );
nand NAND2_26092 ( P2_R2219_U44 , P2_R2219_U78 , P2_R2219_U70 );
nand NAND2_26093 ( P2_R2219_U45 , P2_U2765 , P2_R2219_U23 );
not NOT1_26094 ( P2_R2219_U46 , P2_R2219_U45 );
nand NAND2_26095 ( P2_R2219_U47 , P2_U2764 , P2_R2219_U14 );
nand NAND2_26096 ( P2_R2219_U48 , P2_U2763 , P2_R2219_U17 );
nand NAND2_26097 ( P2_R2219_U49 , P2_R2219_U48 , P2_R2219_U81 );
nand NAND2_26098 ( P2_R2219_U50 , P2_U2755 , P2_R2219_U12 );
not NOT1_26099 ( P2_R2219_U51 , P2_R2219_U43 );
nand NAND2_26100 ( P2_R2219_U52 , P2_U2762 , P2_R2219_U18 );
nand NAND2_26101 ( P2_R2219_U53 , P2_U2754 , P2_R2219_U13 );
not NOT1_26102 ( P2_R2219_U54 , P2_R2219_U42 );
nand NAND2_26103 ( P2_R2219_U55 , P2_U2761 , P2_R2219_U10 );
nand NAND2_26104 ( P2_R2219_U56 , P2_U2753 , P2_R2219_U11 );
not NOT1_26105 ( P2_R2219_U57 , P2_R2219_U41 );
nand NAND2_26106 ( P2_R2219_U58 , P2_U2760 , P2_R2219_U9 );
nand NAND2_26107 ( P2_R2219_U59 , P2_R2219_U58 , P2_R2219_U41 );
nand NAND2_26108 ( P2_R2219_U60 , P2_U4428 , P2_R2219_U20 );
not NOT1_26109 ( P2_R2219_U61 , P2_R2219_U40 );
nand NAND2_26110 ( P2_R2219_U62 , P2_U2759 , P2_R2219_U9 );
nand NAND2_26111 ( P2_R2219_U63 , P2_R2219_U62 , P2_R2219_U40 );
nand NAND2_26112 ( P2_R2219_U64 , P2_U4428 , P2_R2219_U21 );
not NOT1_26113 ( P2_R2219_U65 , P2_R2219_U39 );
nand NAND2_26114 ( P2_R2219_U66 , P2_U4428 , P2_R2219_U22 );
nand NAND2_26115 ( P2_R2219_U67 , P2_U2758 , P2_R2219_U9 );
nand NAND2_26116 ( P2_R2219_U68 , P2_R2219_U67 , P2_R2219_U39 );
nand NAND2_26117 ( P2_R2219_U69 , P2_U2757 , P2_R2219_U15 );
nand NAND2_26118 ( P2_R2219_U70 , P2_U2756 , P2_R2219_U16 );
nand NAND2_26119 ( P2_R2219_U71 , P2_R2219_U6 , P2_R2219_U44 );
nand NAND2_26120 ( P2_R2219_U72 , P2_R2219_U53 , P2_R2219_U50 );
not NOT1_26121 ( P2_R2219_U73 , P2_R2219_U19 );
nand NAND2_26122 ( P2_R2219_U74 , P2_R2219_U31 , P2_R2219_U44 );
nand NAND2_26123 ( P2_R2219_U75 , P2_R2219_U73 , P2_R2219_U55 );
nand NAND2_26124 ( P2_R2219_U76 , P2_U2762 , P2_R2219_U18 );
nand NAND2_26125 ( P2_R2219_U77 , P2_U2764 , P2_R2219_U14 );
nand NAND2_26126 ( P2_R2219_U78 , P2_R2219_U47 , P2_R2219_U45 );
not NOT1_26127 ( P2_R2219_U79 , P2_R2219_U44 );
nand NAND2_26128 ( P2_R2219_U80 , P2_R2219_U77 , P2_R2219_U45 );
nand NAND2_26129 ( P2_R2219_U81 , P2_R2219_U80 , P2_R2219_U70 );
nand NAND2_26130 ( P2_R2219_U82 , P2_U2758 , P2_R2219_U9 );
nand NAND2_26131 ( P2_R2219_U83 , P2_U4428 , P2_R2219_U22 );
not NOT1_26132 ( P2_R2219_U84 , P2_R2219_U32 );
nand NAND2_26133 ( P2_R2219_U85 , P2_R2219_U65 , P2_R2219_U84 );
nand NAND2_26134 ( P2_R2219_U86 , P2_R2219_U32 , P2_R2219_U39 );
nand NAND2_26135 ( P2_R2219_U87 , P2_U2759 , P2_R2219_U9 );
nand NAND2_26136 ( P2_R2219_U88 , P2_U4428 , P2_R2219_U21 );
not NOT1_26137 ( P2_R2219_U89 , P2_R2219_U33 );
nand NAND2_26138 ( P2_R2219_U90 , P2_R2219_U61 , P2_R2219_U89 );
nand NAND2_26139 ( P2_R2219_U91 , P2_R2219_U33 , P2_R2219_U40 );
nand NAND2_26140 ( P2_R2219_U92 , P2_U2760 , P2_R2219_U9 );
nand NAND2_26141 ( P2_R2219_U93 , P2_U4428 , P2_R2219_U20 );
not NOT1_26142 ( P2_R2219_U94 , P2_R2219_U34 );
nand NAND2_26143 ( P2_R2219_U95 , P2_R2219_U57 , P2_R2219_U94 );
nand NAND2_26144 ( P2_R2219_U96 , P2_R2219_U34 , P2_R2219_U41 );
nand NAND2_26145 ( P2_R2219_U97 , P2_U2761 , P2_R2219_U10 );
nand NAND2_26146 ( P2_R2219_U98 , P2_U2753 , P2_R2219_U11 );
not NOT1_26147 ( P2_R2219_U99 , P2_R2219_U35 );
nand NAND2_26148 ( P2_R2219_U100 , P2_R2219_U54 , P2_R2219_U99 );
nand NAND2_26149 ( P2_R2219_U101 , P2_R2219_U35 , P2_R2219_U42 );
nand NAND2_26150 ( P2_R2219_U102 , P2_U2762 , P2_R2219_U18 );
nand NAND2_26151 ( P2_R2219_U103 , P2_U2754 , P2_R2219_U13 );
not NOT1_26152 ( P2_R2219_U104 , P2_R2219_U36 );
nand NAND2_26153 ( P2_R2219_U105 , P2_R2219_U51 , P2_R2219_U104 );
nand NAND2_26154 ( P2_R2219_U106 , P2_R2219_U36 , P2_R2219_U43 );
nand NAND2_26155 ( P2_R2219_U107 , P2_U2763 , P2_R2219_U17 );
nand NAND2_26156 ( P2_R2219_U108 , P2_U2755 , P2_R2219_U12 );
not NOT1_26157 ( P2_R2219_U109 , P2_R2219_U37 );
nand NAND2_26158 ( P2_R2219_U110 , P2_R2219_U79 , P2_R2219_U109 );
nand NAND2_26159 ( P2_R2219_U111 , P2_R2219_U37 , P2_R2219_U44 );
nand NAND2_26160 ( P2_R2219_U112 , P2_U2764 , P2_R2219_U14 );
nand NAND2_26161 ( P2_R2219_U113 , P2_U2756 , P2_R2219_U16 );
not NOT1_26162 ( P2_R2219_U114 , P2_R2219_U38 );
nand NAND2_26163 ( P2_R2219_U115 , P2_R2219_U46 , P2_R2219_U114 );
nand NAND2_26164 ( P2_R2219_U116 , P2_R2219_U38 , P2_R2219_U45 );
nor nor_26165 ( P2_R2243_U6 , P2_U3686 , P2_U3685 , P2_U3684 , P2_U3687 );
nor nor_26166 ( P2_R2243_U7 , P2_U3684 , P2_R2243_U9 );
nand NAND2_26167 ( P2_R2243_U8 , P2_R2243_U7 , P2_R2243_U11 );
nor nor_26168 ( P2_R2243_U9 , P2_U3689 , P2_U3687 , P2_U3684 , P2_U3686 , P2_U3685 );
not NOT1_26169 ( P2_R2243_U10 , P2_U3688 );
nand NAND2_26170 ( P2_R2243_U11 , P2_R2243_U6 , P2_R2243_U10 );
not NOT1_26171 ( P2_SUB_589_U6 , P2_U3614 );
not NOT1_26172 ( P2_SUB_589_U7 , P2_U3615 );
not NOT1_26173 ( P2_SUB_589_U8 , P2_U2813 );
not NOT1_26174 ( P2_SUB_589_U9 , P2_U3613 );
and AND2_26175 ( P2_R2096_U4 , P2_U2640 , P2_R2096_U23 );
and AND2_26176 ( P2_R2096_U5 , P2_U2633 , P2_R2096_U18 );
and AND2_26177 ( P2_R2096_U6 , P2_U2631 , P2_R2096_U25 );
and AND2_26178 ( P2_R2096_U7 , P2_U2629 , P2_R2096_U16 );
and AND2_26179 ( P2_R2096_U8 , P2_U2628 , P2_R2096_U7 );
and AND2_26180 ( P2_R2096_U9 , P2_U2627 , P2_R2096_U8 );
and AND2_26181 ( P2_R2096_U10 , P2_U2626 , P2_R2096_U9 );
and AND2_26182 ( P2_R2096_U11 , P2_U2625 , P2_R2096_U10 );
and AND2_26183 ( P2_R2096_U12 , P2_U2624 , P2_R2096_U11 );
and AND2_26184 ( P2_R2096_U13 , P2_U2622 , P2_R2096_U15 );
and AND2_26185 ( P2_R2096_U14 , P2_U2621 , P2_R2096_U13 );
and AND2_26186 ( P2_R2096_U15 , P2_U2623 , P2_R2096_U12 );
and AND2_26187 ( P2_R2096_U16 , P2_U2630 , P2_R2096_U6 );
and AND2_26188 ( P2_R2096_U17 , P2_U2635 , P2_R2096_U21 );
and AND2_26189 ( P2_R2096_U18 , P2_U2634 , P2_R2096_U17 );
and AND2_26190 ( P2_R2096_U19 , P2_U2638 , P2_R2096_U24 );
and AND2_26191 ( P2_R2096_U20 , P2_U2637 , P2_R2096_U19 );
and AND2_26192 ( P2_R2096_U21 , P2_U2636 , P2_R2096_U20 );
and AND2_26193 ( P2_R2096_U22 , P2_U2620 , P2_R2096_U14 );
and AND2_26194 ( P2_R2096_U23 , P2_U2641 , P2_R2096_U99 );
and AND2_26195 ( P2_R2096_U24 , P2_U2639 , P2_R2096_U4 );
and AND2_26196 ( P2_R2096_U25 , P2_U2632 , P2_R2096_U5 );
not NOT1_26197 ( P2_R2096_U26 , P2_U2631 );
not NOT1_26198 ( P2_R2096_U27 , P2_U2638 );
not NOT1_26199 ( P2_R2096_U28 , P2_U2640 );
not NOT1_26200 ( P2_R2096_U29 , P2_U2618 );
not NOT1_26201 ( P2_R2096_U30 , P2_U2619 );
not NOT1_26202 ( P2_R2096_U31 , P2_U2635 );
not NOT1_26203 ( P2_R2096_U32 , P2_U2636 );
not NOT1_26204 ( P2_R2096_U33 , P2_U2637 );
not NOT1_26205 ( P2_R2096_U34 , P2_U2633 );
not NOT1_26206 ( P2_R2096_U35 , P2_U2634 );
not NOT1_26207 ( P2_R2096_U36 , P2_U2629 );
not NOT1_26208 ( P2_R2096_U37 , P2_U2641 );
not NOT1_26209 ( P2_R2096_U38 , P2_U2622 );
not NOT1_26210 ( P2_R2096_U39 , P2_U2627 );
not NOT1_26211 ( P2_R2096_U40 , P2_U2620 );
not NOT1_26212 ( P2_R2096_U41 , P2_U2621 );
not NOT1_26213 ( P2_R2096_U42 , P2_U2623 );
not NOT1_26214 ( P2_R2096_U43 , P2_U2624 );
not NOT1_26215 ( P2_R2096_U44 , P2_U2625 );
not NOT1_26216 ( P2_R2096_U45 , P2_U2626 );
not NOT1_26217 ( P2_R2096_U46 , P2_U2628 );
not NOT1_26218 ( P2_R2096_U47 , P2_U2630 );
not NOT1_26219 ( P2_R2096_U48 , P2_U2632 );
not NOT1_26220 ( P2_R2096_U49 , P2_U2639 );
and AND2_26221 ( P2_R2096_U50 , P2_R2096_U168 , P2_R2096_U167 );
nand NAND2_26222 ( P2_R2096_U51 , P2_R2096_U114 , P2_R2096_U170 );
not NOT1_26223 ( P2_R2096_U52 , P2_U2657 );
not NOT1_26224 ( P2_R2096_U53 , P2_U2649 );
not NOT1_26225 ( P2_R2096_U54 , P2_U2648 );
not NOT1_26226 ( P2_R2096_U55 , P2_U2656 );
not NOT1_26227 ( P2_R2096_U56 , P2_U2655 );
not NOT1_26228 ( P2_R2096_U57 , P2_U2647 );
not NOT1_26229 ( P2_R2096_U58 , P2_U2654 );
not NOT1_26230 ( P2_R2096_U59 , P2_U2646 );
not NOT1_26231 ( P2_R2096_U60 , P2_U2653 );
not NOT1_26232 ( P2_R2096_U61 , P2_U2645 );
not NOT1_26233 ( P2_R2096_U62 , P2_U2652 );
not NOT1_26234 ( P2_R2096_U63 , P2_U2644 );
not NOT1_26235 ( P2_R2096_U64 , P2_U2651 );
not NOT1_26236 ( P2_R2096_U65 , P2_U2643 );
not NOT1_26237 ( P2_R2096_U66 , P2_U2650 );
not NOT1_26238 ( P2_R2096_U67 , P2_U2642 );
nand NAND2_26239 ( P2_R2096_U68 , P2_R2096_U265 , P2_R2096_U264 );
nand NAND2_26240 ( P2_R2096_U69 , P2_R2096_U172 , P2_R2096_U171 );
nand NAND2_26241 ( P2_R2096_U70 , P2_R2096_U174 , P2_R2096_U173 );
nand NAND2_26242 ( P2_R2096_U71 , P2_R2096_U181 , P2_R2096_U180 );
nand NAND2_26243 ( P2_R2096_U72 , P2_R2096_U188 , P2_R2096_U187 );
nand NAND2_26244 ( P2_R2096_U73 , P2_R2096_U195 , P2_R2096_U194 );
nand NAND2_26245 ( P2_R2096_U74 , P2_R2096_U202 , P2_R2096_U201 );
nand NAND2_26246 ( P2_R2096_U75 , P2_R2096_U209 , P2_R2096_U208 );
nand NAND2_26247 ( P2_R2096_U76 , P2_R2096_U211 , P2_R2096_U210 );
nand NAND2_26248 ( P2_R2096_U77 , P2_R2096_U218 , P2_R2096_U217 );
nand NAND2_26249 ( P2_R2096_U78 , P2_R2096_U220 , P2_R2096_U219 );
nand NAND2_26250 ( P2_R2096_U79 , P2_R2096_U222 , P2_R2096_U221 );
nand NAND2_26251 ( P2_R2096_U80 , P2_R2096_U224 , P2_R2096_U223 );
nand NAND2_26252 ( P2_R2096_U81 , P2_R2096_U226 , P2_R2096_U225 );
nand NAND2_26253 ( P2_R2096_U82 , P2_R2096_U228 , P2_R2096_U227 );
nand NAND2_26254 ( P2_R2096_U83 , P2_R2096_U230 , P2_R2096_U229 );
nand NAND2_26255 ( P2_R2096_U84 , P2_R2096_U232 , P2_R2096_U231 );
nand NAND2_26256 ( P2_R2096_U85 , P2_R2096_U234 , P2_R2096_U233 );
nand NAND2_26257 ( P2_R2096_U86 , P2_R2096_U236 , P2_R2096_U235 );
nand NAND2_26258 ( P2_R2096_U87 , P2_R2096_U238 , P2_R2096_U237 );
nand NAND2_26259 ( P2_R2096_U88 , P2_R2096_U245 , P2_R2096_U244 );
nand NAND2_26260 ( P2_R2096_U89 , P2_R2096_U247 , P2_R2096_U246 );
nand NAND2_26261 ( P2_R2096_U90 , P2_R2096_U249 , P2_R2096_U248 );
nand NAND2_26262 ( P2_R2096_U91 , P2_R2096_U251 , P2_R2096_U250 );
nand NAND2_26263 ( P2_R2096_U92 , P2_R2096_U253 , P2_R2096_U252 );
nand NAND2_26264 ( P2_R2096_U93 , P2_R2096_U255 , P2_R2096_U254 );
nand NAND2_26265 ( P2_R2096_U94 , P2_R2096_U257 , P2_R2096_U256 );
nand NAND2_26266 ( P2_R2096_U95 , P2_R2096_U259 , P2_R2096_U258 );
nand NAND2_26267 ( P2_R2096_U96 , P2_R2096_U261 , P2_R2096_U260 );
nand NAND2_26268 ( P2_R2096_U97 , P2_R2096_U263 , P2_R2096_U262 );
and AND2_26269 ( P2_R2096_U98 , P2_U2619 , P2_U2618 );
nand NAND2_26270 ( P2_R2096_U99 , P2_R2096_U142 , P2_R2096_U141 );
and AND2_26271 ( P2_R2096_U100 , P2_R2096_U176 , P2_R2096_U175 );
nand NAND2_26272 ( P2_R2096_U101 , P2_R2096_U138 , P2_R2096_U137 );
and AND2_26273 ( P2_R2096_U102 , P2_R2096_U183 , P2_R2096_U182 );
nand NAND2_26274 ( P2_R2096_U103 , P2_R2096_U134 , P2_R2096_U133 );
and AND2_26275 ( P2_R2096_U104 , P2_R2096_U190 , P2_R2096_U189 );
nand NAND2_26276 ( P2_R2096_U105 , P2_R2096_U130 , P2_R2096_U129 );
and AND2_26277 ( P2_R2096_U106 , P2_R2096_U197 , P2_R2096_U196 );
nand NAND2_26278 ( P2_R2096_U107 , P2_R2096_U126 , P2_R2096_U125 );
and AND2_26279 ( P2_R2096_U108 , P2_R2096_U204 , P2_R2096_U203 );
nand NAND2_26280 ( P2_R2096_U109 , P2_R2096_U122 , P2_R2096_U121 );
and AND2_26281 ( P2_R2096_U110 , P2_R2096_U213 , P2_R2096_U212 );
nand NAND2_26282 ( P2_R2096_U111 , P2_R2096_U113 , P2_R2096_U118 );
nand NAND2_26283 ( P2_R2096_U112 , P2_U2649 , P2_U2657 );
nand NAND3_26284 ( P2_R2096_U113 , P2_U2649 , P2_U2657 , P2_U2656 );
and AND2_26285 ( P2_R2096_U114 , P2_R2096_U243 , P2_R2096_U242 );
not NOT1_26286 ( P2_R2096_U115 , P2_R2096_U113 );
nand NAND2_26287 ( P2_R2096_U116 , P2_U2649 , P2_U2657 );
nand NAND2_26288 ( P2_R2096_U117 , P2_R2096_U55 , P2_R2096_U116 );
nand NAND2_26289 ( P2_R2096_U118 , P2_U2648 , P2_R2096_U117 );
not NOT1_26290 ( P2_R2096_U119 , P2_R2096_U111 );
or OR2_26291 ( P2_R2096_U120 , P2_U2655 , P2_U2647 );
nand NAND2_26292 ( P2_R2096_U121 , P2_R2096_U120 , P2_R2096_U111 );
nand NAND2_26293 ( P2_R2096_U122 , P2_U2647 , P2_U2655 );
not NOT1_26294 ( P2_R2096_U123 , P2_R2096_U109 );
or OR2_26295 ( P2_R2096_U124 , P2_U2654 , P2_U2646 );
nand NAND2_26296 ( P2_R2096_U125 , P2_R2096_U124 , P2_R2096_U109 );
nand NAND2_26297 ( P2_R2096_U126 , P2_U2646 , P2_U2654 );
not NOT1_26298 ( P2_R2096_U127 , P2_R2096_U107 );
or OR2_26299 ( P2_R2096_U128 , P2_U2653 , P2_U2645 );
nand NAND2_26300 ( P2_R2096_U129 , P2_R2096_U128 , P2_R2096_U107 );
nand NAND2_26301 ( P2_R2096_U130 , P2_U2645 , P2_U2653 );
not NOT1_26302 ( P2_R2096_U131 , P2_R2096_U105 );
or OR2_26303 ( P2_R2096_U132 , P2_U2652 , P2_U2644 );
nand NAND2_26304 ( P2_R2096_U133 , P2_R2096_U132 , P2_R2096_U105 );
nand NAND2_26305 ( P2_R2096_U134 , P2_U2644 , P2_U2652 );
not NOT1_26306 ( P2_R2096_U135 , P2_R2096_U103 );
or OR2_26307 ( P2_R2096_U136 , P2_U2651 , P2_U2643 );
nand NAND2_26308 ( P2_R2096_U137 , P2_R2096_U136 , P2_R2096_U103 );
nand NAND2_26309 ( P2_R2096_U138 , P2_U2643 , P2_U2651 );
not NOT1_26310 ( P2_R2096_U139 , P2_R2096_U101 );
or OR2_26311 ( P2_R2096_U140 , P2_U2650 , P2_U2642 );
nand NAND2_26312 ( P2_R2096_U141 , P2_R2096_U140 , P2_R2096_U101 );
nand NAND2_26313 ( P2_R2096_U142 , P2_U2642 , P2_U2650 );
not NOT1_26314 ( P2_R2096_U143 , P2_R2096_U99 );
not NOT1_26315 ( P2_R2096_U144 , P2_R2096_U23 );
not NOT1_26316 ( P2_R2096_U145 , P2_R2096_U4 );
not NOT1_26317 ( P2_R2096_U146 , P2_R2096_U24 );
not NOT1_26318 ( P2_R2096_U147 , P2_R2096_U19 );
not NOT1_26319 ( P2_R2096_U148 , P2_R2096_U20 );
not NOT1_26320 ( P2_R2096_U149 , P2_R2096_U21 );
not NOT1_26321 ( P2_R2096_U150 , P2_R2096_U17 );
not NOT1_26322 ( P2_R2096_U151 , P2_R2096_U18 );
not NOT1_26323 ( P2_R2096_U152 , P2_R2096_U5 );
not NOT1_26324 ( P2_R2096_U153 , P2_R2096_U25 );
not NOT1_26325 ( P2_R2096_U154 , P2_R2096_U6 );
not NOT1_26326 ( P2_R2096_U155 , P2_R2096_U16 );
not NOT1_26327 ( P2_R2096_U156 , P2_R2096_U7 );
not NOT1_26328 ( P2_R2096_U157 , P2_R2096_U8 );
not NOT1_26329 ( P2_R2096_U158 , P2_R2096_U9 );
not NOT1_26330 ( P2_R2096_U159 , P2_R2096_U10 );
not NOT1_26331 ( P2_R2096_U160 , P2_R2096_U11 );
not NOT1_26332 ( P2_R2096_U161 , P2_R2096_U12 );
not NOT1_26333 ( P2_R2096_U162 , P2_R2096_U15 );
not NOT1_26334 ( P2_R2096_U163 , P2_R2096_U13 );
not NOT1_26335 ( P2_R2096_U164 , P2_R2096_U14 );
not NOT1_26336 ( P2_R2096_U165 , P2_R2096_U22 );
nand NAND2_26337 ( P2_R2096_U166 , P2_U2619 , P2_R2096_U22 );
nand NAND2_26338 ( P2_R2096_U167 , P2_R2096_U29 , P2_R2096_U166 );
nand NAND2_26339 ( P2_R2096_U168 , P2_R2096_U98 , P2_R2096_U22 );
not NOT1_26340 ( P2_R2096_U169 , P2_R2096_U112 );
nand NAND2_26341 ( P2_R2096_U170 , P2_R2096_U241 , P2_R2096_U55 );
nand NAND2_26342 ( P2_R2096_U171 , P2_R2096_U28 , P2_R2096_U23 );
nand NAND2_26343 ( P2_R2096_U172 , P2_R2096_U144 , P2_U2640 );
nand NAND2_26344 ( P2_R2096_U173 , P2_R2096_U37 , P2_R2096_U99 );
nand NAND2_26345 ( P2_R2096_U174 , P2_R2096_U143 , P2_U2641 );
nand NAND2_26346 ( P2_R2096_U175 , P2_U2642 , P2_R2096_U66 );
nand NAND2_26347 ( P2_R2096_U176 , P2_U2650 , P2_R2096_U67 );
nand NAND2_26348 ( P2_R2096_U177 , P2_U2642 , P2_R2096_U66 );
nand NAND2_26349 ( P2_R2096_U178 , P2_U2650 , P2_R2096_U67 );
nand NAND2_26350 ( P2_R2096_U179 , P2_R2096_U178 , P2_R2096_U177 );
nand NAND2_26351 ( P2_R2096_U180 , P2_R2096_U100 , P2_R2096_U101 );
nand NAND2_26352 ( P2_R2096_U181 , P2_R2096_U139 , P2_R2096_U179 );
nand NAND2_26353 ( P2_R2096_U182 , P2_U2643 , P2_R2096_U64 );
nand NAND2_26354 ( P2_R2096_U183 , P2_U2651 , P2_R2096_U65 );
nand NAND2_26355 ( P2_R2096_U184 , P2_U2643 , P2_R2096_U64 );
nand NAND2_26356 ( P2_R2096_U185 , P2_U2651 , P2_R2096_U65 );
nand NAND2_26357 ( P2_R2096_U186 , P2_R2096_U185 , P2_R2096_U184 );
nand NAND2_26358 ( P2_R2096_U187 , P2_R2096_U102 , P2_R2096_U103 );
nand NAND2_26359 ( P2_R2096_U188 , P2_R2096_U135 , P2_R2096_U186 );
nand NAND2_26360 ( P2_R2096_U189 , P2_U2644 , P2_R2096_U62 );
nand NAND2_26361 ( P2_R2096_U190 , P2_U2652 , P2_R2096_U63 );
nand NAND2_26362 ( P2_R2096_U191 , P2_U2644 , P2_R2096_U62 );
nand NAND2_26363 ( P2_R2096_U192 , P2_U2652 , P2_R2096_U63 );
nand NAND2_26364 ( P2_R2096_U193 , P2_R2096_U192 , P2_R2096_U191 );
nand NAND2_26365 ( P2_R2096_U194 , P2_R2096_U104 , P2_R2096_U105 );
nand NAND2_26366 ( P2_R2096_U195 , P2_R2096_U131 , P2_R2096_U193 );
nand NAND2_26367 ( P2_R2096_U196 , P2_U2645 , P2_R2096_U60 );
nand NAND2_26368 ( P2_R2096_U197 , P2_U2653 , P2_R2096_U61 );
nand NAND2_26369 ( P2_R2096_U198 , P2_U2645 , P2_R2096_U60 );
nand NAND2_26370 ( P2_R2096_U199 , P2_U2653 , P2_R2096_U61 );
nand NAND2_26371 ( P2_R2096_U200 , P2_R2096_U199 , P2_R2096_U198 );
nand NAND2_26372 ( P2_R2096_U201 , P2_R2096_U106 , P2_R2096_U107 );
nand NAND2_26373 ( P2_R2096_U202 , P2_R2096_U127 , P2_R2096_U200 );
nand NAND2_26374 ( P2_R2096_U203 , P2_U2646 , P2_R2096_U58 );
nand NAND2_26375 ( P2_R2096_U204 , P2_U2654 , P2_R2096_U59 );
nand NAND2_26376 ( P2_R2096_U205 , P2_U2646 , P2_R2096_U58 );
nand NAND2_26377 ( P2_R2096_U206 , P2_U2654 , P2_R2096_U59 );
nand NAND2_26378 ( P2_R2096_U207 , P2_R2096_U206 , P2_R2096_U205 );
nand NAND2_26379 ( P2_R2096_U208 , P2_R2096_U108 , P2_R2096_U109 );
nand NAND2_26380 ( P2_R2096_U209 , P2_R2096_U123 , P2_R2096_U207 );
nand NAND2_26381 ( P2_R2096_U210 , P2_R2096_U30 , P2_R2096_U22 );
nand NAND2_26382 ( P2_R2096_U211 , P2_U2619 , P2_R2096_U165 );
nand NAND2_26383 ( P2_R2096_U212 , P2_U2647 , P2_R2096_U56 );
nand NAND2_26384 ( P2_R2096_U213 , P2_U2655 , P2_R2096_U57 );
nand NAND2_26385 ( P2_R2096_U214 , P2_U2647 , P2_R2096_U56 );
nand NAND2_26386 ( P2_R2096_U215 , P2_U2655 , P2_R2096_U57 );
nand NAND2_26387 ( P2_R2096_U216 , P2_R2096_U215 , P2_R2096_U214 );
nand NAND2_26388 ( P2_R2096_U217 , P2_R2096_U110 , P2_R2096_U111 );
nand NAND2_26389 ( P2_R2096_U218 , P2_R2096_U119 , P2_R2096_U216 );
nand NAND2_26390 ( P2_R2096_U219 , P2_R2096_U40 , P2_R2096_U14 );
nand NAND2_26391 ( P2_R2096_U220 , P2_R2096_U164 , P2_U2620 );
nand NAND2_26392 ( P2_R2096_U221 , P2_R2096_U41 , P2_R2096_U13 );
nand NAND2_26393 ( P2_R2096_U222 , P2_R2096_U163 , P2_U2621 );
nand NAND2_26394 ( P2_R2096_U223 , P2_R2096_U38 , P2_R2096_U15 );
nand NAND2_26395 ( P2_R2096_U224 , P2_R2096_U162 , P2_U2622 );
nand NAND2_26396 ( P2_R2096_U225 , P2_R2096_U42 , P2_R2096_U12 );
nand NAND2_26397 ( P2_R2096_U226 , P2_R2096_U161 , P2_U2623 );
nand NAND2_26398 ( P2_R2096_U227 , P2_R2096_U43 , P2_R2096_U11 );
nand NAND2_26399 ( P2_R2096_U228 , P2_R2096_U160 , P2_U2624 );
nand NAND2_26400 ( P2_R2096_U229 , P2_R2096_U44 , P2_R2096_U10 );
nand NAND2_26401 ( P2_R2096_U230 , P2_R2096_U159 , P2_U2625 );
nand NAND2_26402 ( P2_R2096_U231 , P2_R2096_U45 , P2_R2096_U9 );
nand NAND2_26403 ( P2_R2096_U232 , P2_R2096_U158 , P2_U2626 );
nand NAND2_26404 ( P2_R2096_U233 , P2_R2096_U39 , P2_R2096_U8 );
nand NAND2_26405 ( P2_R2096_U234 , P2_R2096_U157 , P2_U2627 );
nand NAND2_26406 ( P2_R2096_U235 , P2_R2096_U46 , P2_R2096_U7 );
nand NAND2_26407 ( P2_R2096_U236 , P2_R2096_U156 , P2_U2628 );
nand NAND2_26408 ( P2_R2096_U237 , P2_R2096_U36 , P2_R2096_U16 );
nand NAND2_26409 ( P2_R2096_U238 , P2_R2096_U155 , P2_U2629 );
nand NAND2_26410 ( P2_R2096_U239 , P2_U2648 , P2_R2096_U112 );
nand NAND2_26411 ( P2_R2096_U240 , P2_R2096_U169 , P2_R2096_U54 );
nand NAND2_26412 ( P2_R2096_U241 , P2_R2096_U240 , P2_R2096_U239 );
nand NAND3_26413 ( P2_R2096_U242 , P2_U2656 , P2_R2096_U116 , P2_R2096_U54 );
nand NAND2_26414 ( P2_R2096_U243 , P2_R2096_U115 , P2_U2648 );
nand NAND2_26415 ( P2_R2096_U244 , P2_R2096_U47 , P2_R2096_U6 );
nand NAND2_26416 ( P2_R2096_U245 , P2_R2096_U154 , P2_U2630 );
nand NAND2_26417 ( P2_R2096_U246 , P2_R2096_U26 , P2_R2096_U25 );
nand NAND2_26418 ( P2_R2096_U247 , P2_R2096_U153 , P2_U2631 );
nand NAND2_26419 ( P2_R2096_U248 , P2_R2096_U48 , P2_R2096_U5 );
nand NAND2_26420 ( P2_R2096_U249 , P2_R2096_U152 , P2_U2632 );
nand NAND2_26421 ( P2_R2096_U250 , P2_R2096_U34 , P2_R2096_U18 );
nand NAND2_26422 ( P2_R2096_U251 , P2_R2096_U151 , P2_U2633 );
nand NAND2_26423 ( P2_R2096_U252 , P2_R2096_U35 , P2_R2096_U17 );
nand NAND2_26424 ( P2_R2096_U253 , P2_R2096_U150 , P2_U2634 );
nand NAND2_26425 ( P2_R2096_U254 , P2_R2096_U31 , P2_R2096_U21 );
nand NAND2_26426 ( P2_R2096_U255 , P2_R2096_U149 , P2_U2635 );
nand NAND2_26427 ( P2_R2096_U256 , P2_R2096_U32 , P2_R2096_U20 );
nand NAND2_26428 ( P2_R2096_U257 , P2_R2096_U148 , P2_U2636 );
nand NAND2_26429 ( P2_R2096_U258 , P2_R2096_U33 , P2_R2096_U19 );
nand NAND2_26430 ( P2_R2096_U259 , P2_R2096_U147 , P2_U2637 );
nand NAND2_26431 ( P2_R2096_U260 , P2_R2096_U27 , P2_R2096_U24 );
nand NAND2_26432 ( P2_R2096_U261 , P2_R2096_U146 , P2_U2638 );
nand NAND2_26433 ( P2_R2096_U262 , P2_R2096_U49 , P2_R2096_U4 );
nand NAND2_26434 ( P2_R2096_U263 , P2_R2096_U145 , P2_U2639 );
nand NAND2_26435 ( P2_R2096_U264 , P2_U2649 , P2_R2096_U52 );
nand NAND2_26436 ( P2_R2096_U265 , P2_U2657 , P2_R2096_U53 );
nor nor_26437 ( P2_GTE_370_U6 , P2_R2219_U25 , P2_GTE_370_U8 );
and AND2_26438 ( P2_GTE_370_U7 , P2_R2219_U29 , P2_GTE_370_U9 );
nor nor_26439 ( P2_GTE_370_U8 , P2_R2219_U26 , P2_R2219_U27 , P2_R2219_U28 , P2_GTE_370_U7 );
or OR2_26440 ( P2_GTE_370_U9 , P2_R2219_U8 , P2_R2219_U30 );
and AND2_26441 ( P2_LT_563_U6 , P2_LT_563_U27 , P2_LT_563_U26 );
not NOT1_26442 ( P2_LT_563_U7 , P2_U3620 );
not NOT1_26443 ( P2_LT_563_U8 , P2_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_26444 ( P2_LT_563_U9 , P2_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_26445 ( P2_LT_563_U10 , P2_U3619 );
not NOT1_26446 ( P2_LT_563_U11 , P2_U3618 );
not NOT1_26447 ( P2_LT_563_U12 , P2_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_26448 ( P2_LT_563_U13 , P2_INSTQUEUEWR_ADDR_REG_4_ );
not NOT1_26449 ( P2_LT_563_U14 , P2_U3617 );
not NOT1_26450 ( P2_LT_563_U15 , P2_U3621 );
nand NAND2_26451 ( P2_LT_563_U16 , P2_U3620 , P2_LT_563_U8 );
nand NAND3_26452 ( P2_LT_563_U17 , P2_INSTQUEUEWR_ADDR_REG_0_ , P2_LT_563_U15 , P2_LT_563_U16 );
nand NAND2_26453 ( P2_LT_563_U18 , P2_INSTQUEUEWR_ADDR_REG_1_ , P2_LT_563_U7 );
nand NAND2_26454 ( P2_LT_563_U19 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_LT_563_U10 );
nand NAND3_26455 ( P2_LT_563_U20 , P2_LT_563_U18 , P2_LT_563_U19 , P2_LT_563_U17 );
nand NAND2_26456 ( P2_LT_563_U21 , P2_U3619 , P2_LT_563_U9 );
nand NAND2_26457 ( P2_LT_563_U22 , P2_U3618 , P2_LT_563_U12 );
nand NAND3_26458 ( P2_LT_563_U23 , P2_LT_563_U21 , P2_LT_563_U22 , P2_LT_563_U20 );
nand NAND2_26459 ( P2_LT_563_U24 , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_LT_563_U11 );
nand NAND2_26460 ( P2_LT_563_U25 , P2_INSTQUEUEWR_ADDR_REG_4_ , P2_LT_563_U14 );
nand NAND3_26461 ( P2_LT_563_U26 , P2_LT_563_U24 , P2_LT_563_U25 , P2_LT_563_U23 );
nand NAND2_26462 ( P2_LT_563_U27 , P2_U3617 , P2_LT_563_U13 );
nand NAND2_26463 ( P2_R2256_U4 , P2_R2256_U31 , P2_R2256_U46 );
and AND2_26464 ( P2_R2256_U5 , P2_R2256_U23 , P2_R2256_U43 );
not NOT1_26465 ( P2_R2256_U6 , P2_U3629 );
not NOT1_26466 ( P2_R2256_U7 , P2_U3628 );
not NOT1_26467 ( P2_R2256_U8 , P2_U3627 );
not NOT1_26468 ( P2_R2256_U9 , P2_U3626 );
nand NAND2_26469 ( P2_R2256_U10 , P2_U3626 , P2_R2256_U25 );
not NOT1_26470 ( P2_R2256_U11 , P2_U3625 );
nand NAND2_26471 ( P2_R2256_U12 , P2_U3625 , P2_R2256_U41 );
not NOT1_26472 ( P2_R2256_U13 , P2_U3624 );
nand NAND2_26473 ( P2_R2256_U14 , P2_U3624 , P2_R2256_U42 );
not NOT1_26474 ( P2_R2256_U15 , P2_U3622 );
not NOT1_26475 ( P2_R2256_U16 , P2_U3623 );
nand NAND2_26476 ( P2_R2256_U17 , P2_R2256_U48 , P2_R2256_U47 );
nand NAND2_26477 ( P2_R2256_U18 , P2_R2256_U50 , P2_R2256_U49 );
nand NAND2_26478 ( P2_R2256_U19 , P2_R2256_U52 , P2_R2256_U51 );
nand NAND2_26479 ( P2_R2256_U20 , P2_R2256_U54 , P2_R2256_U53 );
nand NAND2_26480 ( P2_R2256_U21 , P2_R2256_U70 , P2_R2256_U69 );
nand NAND2_26481 ( P2_R2256_U22 , P2_R2256_U63 , P2_R2256_U62 );
and AND2_26482 ( P2_R2256_U23 , P2_U3622 , P2_U3623 );
nand NAND2_26483 ( P2_R2256_U24 , P2_U3623 , P2_R2256_U43 );
nand NAND2_26484 ( P2_R2256_U25 , P2_R2256_U39 , P2_R2256_U38 );
and AND2_26485 ( P2_R2256_U26 , P2_R2256_U56 , P2_R2256_U55 );
and AND2_26486 ( P2_R2256_U27 , P2_R2256_U58 , P2_R2256_U57 );
nand NAND2_26487 ( P2_R2256_U28 , P2_R2256_U30 , P2_R2256_U35 );
nand NAND2_26488 ( P2_R2256_U29 , P2_U7873 , P2_U3629 );
nand NAND3_26489 ( P2_R2256_U30 , P2_U7873 , P2_U3629 , P2_U3628 );
and AND2_26490 ( P2_R2256_U31 , P2_R2256_U68 , P2_R2256_U67 );
not NOT1_26491 ( P2_R2256_U32 , P2_R2256_U30 );
nand NAND2_26492 ( P2_R2256_U33 , P2_U7873 , P2_U3629 );
nand NAND2_26493 ( P2_R2256_U34 , P2_R2256_U7 , P2_R2256_U33 );
nand NAND2_26494 ( P2_R2256_U35 , P2_U2616 , P2_R2256_U34 );
not NOT1_26495 ( P2_R2256_U36 , P2_R2256_U28 );
or OR2_26496 ( P2_R2256_U37 , P2_U3627 , P2_U7873 );
nand NAND2_26497 ( P2_R2256_U38 , P2_R2256_U37 , P2_R2256_U28 );
nand NAND2_26498 ( P2_R2256_U39 , P2_U7873 , P2_U3627 );
not NOT1_26499 ( P2_R2256_U40 , P2_R2256_U25 );
not NOT1_26500 ( P2_R2256_U41 , P2_R2256_U10 );
not NOT1_26501 ( P2_R2256_U42 , P2_R2256_U12 );
not NOT1_26502 ( P2_R2256_U43 , P2_R2256_U14 );
not NOT1_26503 ( P2_R2256_U44 , P2_R2256_U24 );
not NOT1_26504 ( P2_R2256_U45 , P2_R2256_U29 );
nand NAND2_26505 ( P2_R2256_U46 , P2_R2256_U66 , P2_R2256_U7 );
nand NAND2_26506 ( P2_R2256_U47 , P2_U3622 , P2_R2256_U24 );
nand NAND2_26507 ( P2_R2256_U48 , P2_R2256_U44 , P2_R2256_U15 );
nand NAND2_26508 ( P2_R2256_U49 , P2_U3623 , P2_R2256_U14 );
nand NAND2_26509 ( P2_R2256_U50 , P2_R2256_U43 , P2_R2256_U16 );
nand NAND2_26510 ( P2_R2256_U51 , P2_U3624 , P2_R2256_U12 );
nand NAND2_26511 ( P2_R2256_U52 , P2_R2256_U42 , P2_R2256_U13 );
nand NAND2_26512 ( P2_R2256_U53 , P2_U3625 , P2_R2256_U10 );
nand NAND2_26513 ( P2_R2256_U54 , P2_R2256_U41 , P2_R2256_U11 );
nand NAND2_26514 ( P2_R2256_U55 , P2_U3626 , P2_R2256_U25 );
nand NAND2_26515 ( P2_R2256_U56 , P2_R2256_U40 , P2_R2256_U9 );
nand NAND2_26516 ( P2_R2256_U57 , P2_U7873 , P2_R2256_U8 );
nand NAND2_26517 ( P2_R2256_U58 , P2_U3627 , P2_U2616 );
nand NAND2_26518 ( P2_R2256_U59 , P2_U7873 , P2_R2256_U8 );
nand NAND2_26519 ( P2_R2256_U60 , P2_U3627 , P2_U2616 );
nand NAND2_26520 ( P2_R2256_U61 , P2_R2256_U60 , P2_R2256_U59 );
nand NAND2_26521 ( P2_R2256_U62 , P2_R2256_U27 , P2_R2256_U28 );
nand NAND2_26522 ( P2_R2256_U63 , P2_R2256_U36 , P2_R2256_U61 );
nand NAND2_26523 ( P2_R2256_U64 , P2_U2616 , P2_R2256_U29 );
nand NAND2_26524 ( P2_R2256_U65 , P2_R2256_U45 , P2_U7873 );
nand NAND2_26525 ( P2_R2256_U66 , P2_R2256_U65 , P2_R2256_U64 );
nand NAND3_26526 ( P2_R2256_U67 , P2_U3628 , P2_R2256_U33 , P2_U7873 );
nand NAND2_26527 ( P2_R2256_U68 , P2_R2256_U32 , P2_U2616 );
nand NAND2_26528 ( P2_R2256_U69 , P2_U7873 , P2_R2256_U6 );
nand NAND2_26529 ( P2_R2256_U70 , P2_U3629 , P2_U2616 );
nand NAND2_26530 ( P2_R2238_U6 , P2_R2238_U45 , P2_R2238_U44 );
nand NAND2_26531 ( P2_R2238_U7 , P2_R2238_U9 , P2_R2238_U46 );
not NOT1_26532 ( P2_R2238_U8 , P2_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_26533 ( P2_R2238_U9 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_R2238_U18 );
not NOT1_26534 ( P2_R2238_U10 , P2_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_26535 ( P2_R2238_U11 , P2_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_26536 ( P2_R2238_U12 , P2_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_26537 ( P2_R2238_U13 , P2_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_26538 ( P2_R2238_U14 , P2_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_26539 ( P2_R2238_U15 , P2_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_26540 ( P2_R2238_U16 , P2_R2238_U41 , P2_R2238_U40 );
not NOT1_26541 ( P2_R2238_U17 , P2_INSTQUEUERD_ADDR_REG_4_ );
not NOT1_26542 ( P2_R2238_U18 , P2_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_26543 ( P2_R2238_U19 , P2_R2238_U51 , P2_R2238_U50 );
nand NAND2_26544 ( P2_R2238_U20 , P2_R2238_U56 , P2_R2238_U55 );
nand NAND2_26545 ( P2_R2238_U21 , P2_R2238_U61 , P2_R2238_U60 );
nand NAND2_26546 ( P2_R2238_U22 , P2_R2238_U66 , P2_R2238_U65 );
nand NAND2_26547 ( P2_R2238_U23 , P2_R2238_U48 , P2_R2238_U47 );
nand NAND2_26548 ( P2_R2238_U24 , P2_R2238_U53 , P2_R2238_U52 );
nand NAND2_26549 ( P2_R2238_U25 , P2_R2238_U58 , P2_R2238_U57 );
nand NAND2_26550 ( P2_R2238_U26 , P2_R2238_U63 , P2_R2238_U62 );
nand NAND2_26551 ( P2_R2238_U27 , P2_R2238_U37 , P2_R2238_U36 );
nand NAND2_26552 ( P2_R2238_U28 , P2_R2238_U33 , P2_R2238_U32 );
not NOT1_26553 ( P2_R2238_U29 , P2_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_26554 ( P2_R2238_U30 , P2_R2238_U9 );
nand NAND2_26555 ( P2_R2238_U31 , P2_R2238_U30 , P2_R2238_U10 );
nand NAND2_26556 ( P2_R2238_U32 , P2_R2238_U31 , P2_R2238_U29 );
nand NAND2_26557 ( P2_R2238_U33 , P2_INSTQUEUEWR_ADDR_REG_1_ , P2_R2238_U9 );
not NOT1_26558 ( P2_R2238_U34 , P2_R2238_U28 );
nand NAND2_26559 ( P2_R2238_U35 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_R2238_U12 );
nand NAND2_26560 ( P2_R2238_U36 , P2_R2238_U35 , P2_R2238_U28 );
nand NAND2_26561 ( P2_R2238_U37 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_R2238_U11 );
not NOT1_26562 ( P2_R2238_U38 , P2_R2238_U27 );
nand NAND2_26563 ( P2_R2238_U39 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_R2238_U14 );
nand NAND2_26564 ( P2_R2238_U40 , P2_R2238_U39 , P2_R2238_U27 );
nand NAND2_26565 ( P2_R2238_U41 , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_R2238_U13 );
not NOT1_26566 ( P2_R2238_U42 , P2_R2238_U16 );
nand NAND2_26567 ( P2_R2238_U43 , P2_INSTQUEUEWR_ADDR_REG_4_ , P2_R2238_U17 );
nand NAND2_26568 ( P2_R2238_U44 , P2_R2238_U42 , P2_R2238_U43 );
nand NAND2_26569 ( P2_R2238_U45 , P2_INSTQUEUERD_ADDR_REG_4_ , P2_R2238_U15 );
nand NAND2_26570 ( P2_R2238_U46 , P2_INSTQUEUEWR_ADDR_REG_0_ , P2_R2238_U8 );
nand NAND2_26571 ( P2_R2238_U47 , P2_INSTQUEUERD_ADDR_REG_4_ , P2_R2238_U15 );
nand NAND2_26572 ( P2_R2238_U48 , P2_INSTQUEUEWR_ADDR_REG_4_ , P2_R2238_U17 );
not NOT1_26573 ( P2_R2238_U49 , P2_R2238_U23 );
nand NAND2_26574 ( P2_R2238_U50 , P2_R2238_U49 , P2_R2238_U42 );
nand NAND2_26575 ( P2_R2238_U51 , P2_R2238_U23 , P2_R2238_U16 );
nand NAND2_26576 ( P2_R2238_U52 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_R2238_U14 );
nand NAND2_26577 ( P2_R2238_U53 , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_R2238_U13 );
not NOT1_26578 ( P2_R2238_U54 , P2_R2238_U24 );
nand NAND2_26579 ( P2_R2238_U55 , P2_R2238_U38 , P2_R2238_U54 );
nand NAND2_26580 ( P2_R2238_U56 , P2_R2238_U24 , P2_R2238_U27 );
nand NAND2_26581 ( P2_R2238_U57 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_R2238_U12 );
nand NAND2_26582 ( P2_R2238_U58 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_R2238_U11 );
not NOT1_26583 ( P2_R2238_U59 , P2_R2238_U25 );
nand NAND2_26584 ( P2_R2238_U60 , P2_R2238_U34 , P2_R2238_U59 );
nand NAND2_26585 ( P2_R2238_U61 , P2_R2238_U25 , P2_R2238_U28 );
nand NAND2_26586 ( P2_R2238_U62 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_R2238_U10 );
nand NAND2_26587 ( P2_R2238_U63 , P2_INSTQUEUEWR_ADDR_REG_1_ , P2_R2238_U29 );
not NOT1_26588 ( P2_R2238_U64 , P2_R2238_U26 );
nand NAND2_26589 ( P2_R2238_U65 , P2_R2238_U64 , P2_R2238_U30 );
nand NAND2_26590 ( P2_R2238_U66 , P2_R2238_U26 , P2_R2238_U9 );
and AND2_26591 ( P2_R1957_U6 , P2_R1957_U126 , P2_R1957_U27 );
and AND2_26592 ( P2_R1957_U7 , P2_R1957_U124 , P2_R1957_U28 );
and AND2_26593 ( P2_R1957_U8 , P2_R1957_U122 , P2_R1957_U29 );
and AND2_26594 ( P2_R1957_U9 , P2_R1957_U120 , P2_R1957_U30 );
and AND2_26595 ( P2_R1957_U10 , P2_R1957_U118 , P2_R1957_U31 );
and AND2_26596 ( P2_R1957_U11 , P2_R1957_U116 , P2_R1957_U32 );
and AND2_26597 ( P2_R1957_U12 , P2_R1957_U114 , P2_R1957_U33 );
and AND2_26598 ( P2_R1957_U13 , P2_R1957_U112 , P2_R1957_U34 );
and AND2_26599 ( P2_R1957_U14 , P2_R1957_U110 , P2_R1957_U35 );
and AND2_26600 ( P2_R1957_U15 , P2_R1957_U108 , P2_R1957_U36 );
and AND2_26601 ( P2_R1957_U16 , P2_R1957_U106 , P2_R1957_U37 );
and AND2_26602 ( P2_R1957_U17 , P2_R1957_U105 , P2_R1957_U21 );
and AND2_26603 ( P2_R1957_U18 , P2_R1957_U92 , P2_R1957_U22 );
and AND2_26604 ( P2_R1957_U19 , P2_R1957_U90 , P2_R1957_U23 );
and AND2_26605 ( P2_R1957_U20 , P2_R1957_U88 , P2_R1957_U24 );
or OR3_26606 ( P2_R1957_U21 , P2_U3682 , P2_U3683 , P2_U3671 );
nand NAND2_26607 ( P2_R1957_U22 , P2_R1957_U51 , P2_R1957_U83 );
nand NAND3_26608 ( P2_R1957_U23 , P2_R1957_U84 , P2_R1957_U56 , P2_R1957_U26 );
nand NAND3_26609 ( P2_R1957_U24 , P2_R1957_U85 , P2_R1957_U54 , P2_R1957_U25 );
not NOT1_26610 ( P2_R1957_U25 , P2_U3654 );
not NOT1_26611 ( P2_R1957_U26 , P2_U3656 );
nand NAND3_26612 ( P2_R1957_U27 , P2_R1957_U52 , P2_R1957_U86 , P2_R1957_U48 );
nand NAND3_26613 ( P2_R1957_U28 , P2_R1957_U93 , P2_R1957_U81 , P2_R1957_U47 );
nand NAND3_26614 ( P2_R1957_U29 , P2_R1957_U94 , P2_R1957_U79 , P2_R1957_U46 );
nand NAND3_26615 ( P2_R1957_U30 , P2_R1957_U95 , P2_R1957_U77 , P2_R1957_U45 );
nand NAND3_26616 ( P2_R1957_U31 , P2_R1957_U96 , P2_R1957_U75 , P2_R1957_U44 );
nand NAND3_26617 ( P2_R1957_U32 , P2_R1957_U97 , P2_R1957_U73 , P2_R1957_U43 );
nand NAND3_26618 ( P2_R1957_U33 , P2_R1957_U98 , P2_R1957_U69 , P2_R1957_U42 );
nand NAND3_26619 ( P2_R1957_U34 , P2_R1957_U99 , P2_R1957_U67 , P2_R1957_U41 );
nand NAND3_26620 ( P2_R1957_U35 , P2_R1957_U100 , P2_R1957_U65 , P2_R1957_U40 );
nand NAND3_26621 ( P2_R1957_U36 , P2_R1957_U101 , P2_R1957_U63 , P2_R1957_U39 );
nand NAND2_26622 ( P2_R1957_U37 , P2_R1957_U102 , P2_R1957_U38 );
not NOT1_26623 ( P2_R1957_U38 , P2_U3661 );
not NOT1_26624 ( P2_R1957_U39 , P2_U3662 );
not NOT1_26625 ( P2_R1957_U40 , P2_U3664 );
not NOT1_26626 ( P2_R1957_U41 , P2_U3666 );
not NOT1_26627 ( P2_R1957_U42 , P2_U3668 );
not NOT1_26628 ( P2_R1957_U43 , P2_U3670 );
not NOT1_26629 ( P2_R1957_U44 , P2_U3673 );
not NOT1_26630 ( P2_R1957_U45 , P2_U3675 );
not NOT1_26631 ( P2_R1957_U46 , P2_U3677 );
not NOT1_26632 ( P2_R1957_U47 , P2_U3679 );
not NOT1_26633 ( P2_R1957_U48 , P2_U3681 );
nand NAND2_26634 ( P2_R1957_U49 , P2_R1957_U149 , P2_R1957_U148 );
nand NAND2_26635 ( P2_R1957_U50 , P2_R1957_U137 , P2_R1957_U136 );
nor nor_26636 ( P2_R1957_U51 , P2_U3660 , P2_U3658 );
not NOT1_26637 ( P2_R1957_U52 , P2_U3653 );
and AND2_26638 ( P2_R1957_U53 , P2_R1957_U129 , P2_R1957_U128 );
not NOT1_26639 ( P2_R1957_U54 , P2_U3655 );
and AND2_26640 ( P2_R1957_U55 , P2_R1957_U131 , P2_R1957_U130 );
not NOT1_26641 ( P2_R1957_U56 , P2_U3657 );
and AND2_26642 ( P2_R1957_U57 , P2_R1957_U133 , P2_R1957_U132 );
not NOT1_26643 ( P2_R1957_U58 , P2_U3660 );
and AND2_26644 ( P2_R1957_U59 , P2_R1957_U135 , P2_R1957_U134 );
not NOT1_26645 ( P2_R1957_U60 , P2_U3647 );
not NOT1_26646 ( P2_R1957_U61 , P2_U3659 );
and AND2_26647 ( P2_R1957_U62 , P2_R1957_U139 , P2_R1957_U138 );
not NOT1_26648 ( P2_R1957_U63 , P2_U3663 );
and AND2_26649 ( P2_R1957_U64 , P2_R1957_U141 , P2_R1957_U140 );
not NOT1_26650 ( P2_R1957_U65 , P2_U3665 );
and AND2_26651 ( P2_R1957_U66 , P2_R1957_U143 , P2_R1957_U142 );
not NOT1_26652 ( P2_R1957_U67 , P2_U3667 );
and AND2_26653 ( P2_R1957_U68 , P2_R1957_U145 , P2_R1957_U144 );
not NOT1_26654 ( P2_R1957_U69 , P2_U3669 );
and AND2_26655 ( P2_R1957_U70 , P2_R1957_U147 , P2_R1957_U146 );
not NOT1_26656 ( P2_R1957_U71 , P2_U3682 );
not NOT1_26657 ( P2_R1957_U72 , P2_U3683 );
not NOT1_26658 ( P2_R1957_U73 , P2_U3672 );
and AND2_26659 ( P2_R1957_U74 , P2_R1957_U151 , P2_R1957_U150 );
not NOT1_26660 ( P2_R1957_U75 , P2_U3674 );
and AND2_26661 ( P2_R1957_U76 , P2_R1957_U153 , P2_R1957_U152 );
not NOT1_26662 ( P2_R1957_U77 , P2_U3676 );
and AND2_26663 ( P2_R1957_U78 , P2_R1957_U155 , P2_R1957_U154 );
not NOT1_26664 ( P2_R1957_U79 , P2_U3678 );
and AND2_26665 ( P2_R1957_U80 , P2_R1957_U157 , P2_R1957_U156 );
not NOT1_26666 ( P2_R1957_U81 , P2_U3680 );
and AND2_26667 ( P2_R1957_U82 , P2_R1957_U159 , P2_R1957_U158 );
not NOT1_26668 ( P2_R1957_U83 , P2_R1957_U21 );
not NOT1_26669 ( P2_R1957_U84 , P2_R1957_U22 );
not NOT1_26670 ( P2_R1957_U85 , P2_R1957_U23 );
not NOT1_26671 ( P2_R1957_U86 , P2_R1957_U24 );
nand NAND2_26672 ( P2_R1957_U87 , P2_R1957_U85 , P2_R1957_U54 );
nand NAND2_26673 ( P2_R1957_U88 , P2_U3654 , P2_R1957_U87 );
nand NAND2_26674 ( P2_R1957_U89 , P2_R1957_U84 , P2_R1957_U56 );
nand NAND2_26675 ( P2_R1957_U90 , P2_U3656 , P2_R1957_U89 );
nand NAND2_26676 ( P2_R1957_U91 , P2_R1957_U83 , P2_R1957_U58 );
nand NAND2_26677 ( P2_R1957_U92 , P2_U3658 , P2_R1957_U91 );
not NOT1_26678 ( P2_R1957_U93 , P2_R1957_U27 );
not NOT1_26679 ( P2_R1957_U94 , P2_R1957_U28 );
not NOT1_26680 ( P2_R1957_U95 , P2_R1957_U29 );
not NOT1_26681 ( P2_R1957_U96 , P2_R1957_U30 );
not NOT1_26682 ( P2_R1957_U97 , P2_R1957_U31 );
not NOT1_26683 ( P2_R1957_U98 , P2_R1957_U32 );
not NOT1_26684 ( P2_R1957_U99 , P2_R1957_U33 );
not NOT1_26685 ( P2_R1957_U100 , P2_R1957_U34 );
not NOT1_26686 ( P2_R1957_U101 , P2_R1957_U35 );
not NOT1_26687 ( P2_R1957_U102 , P2_R1957_U36 );
not NOT1_26688 ( P2_R1957_U103 , P2_R1957_U37 );
or OR2_26689 ( P2_R1957_U104 , P2_U3682 , P2_U3683 );
nand NAND2_26690 ( P2_R1957_U105 , P2_U3671 , P2_R1957_U104 );
nand NAND2_26691 ( P2_R1957_U106 , P2_U3661 , P2_R1957_U36 );
nand NAND2_26692 ( P2_R1957_U107 , P2_R1957_U101 , P2_R1957_U63 );
nand NAND2_26693 ( P2_R1957_U108 , P2_U3662 , P2_R1957_U107 );
nand NAND2_26694 ( P2_R1957_U109 , P2_R1957_U100 , P2_R1957_U65 );
nand NAND2_26695 ( P2_R1957_U110 , P2_U3664 , P2_R1957_U109 );
nand NAND2_26696 ( P2_R1957_U111 , P2_R1957_U99 , P2_R1957_U67 );
nand NAND2_26697 ( P2_R1957_U112 , P2_U3666 , P2_R1957_U111 );
nand NAND2_26698 ( P2_R1957_U113 , P2_R1957_U98 , P2_R1957_U69 );
nand NAND2_26699 ( P2_R1957_U114 , P2_U3668 , P2_R1957_U113 );
nand NAND2_26700 ( P2_R1957_U115 , P2_R1957_U97 , P2_R1957_U73 );
nand NAND2_26701 ( P2_R1957_U116 , P2_U3670 , P2_R1957_U115 );
nand NAND2_26702 ( P2_R1957_U117 , P2_R1957_U96 , P2_R1957_U75 );
nand NAND2_26703 ( P2_R1957_U118 , P2_U3673 , P2_R1957_U117 );
nand NAND2_26704 ( P2_R1957_U119 , P2_R1957_U95 , P2_R1957_U77 );
nand NAND2_26705 ( P2_R1957_U120 , P2_U3675 , P2_R1957_U119 );
nand NAND2_26706 ( P2_R1957_U121 , P2_R1957_U94 , P2_R1957_U79 );
nand NAND2_26707 ( P2_R1957_U122 , P2_U3677 , P2_R1957_U121 );
nand NAND2_26708 ( P2_R1957_U123 , P2_R1957_U93 , P2_R1957_U81 );
nand NAND2_26709 ( P2_R1957_U124 , P2_U3679 , P2_R1957_U123 );
nand NAND2_26710 ( P2_R1957_U125 , P2_R1957_U86 , P2_R1957_U52 );
nand NAND2_26711 ( P2_R1957_U126 , P2_U3681 , P2_R1957_U125 );
nand NAND2_26712 ( P2_R1957_U127 , P2_R1957_U103 , P2_R1957_U61 );
nand NAND2_26713 ( P2_R1957_U128 , P2_U3653 , P2_R1957_U24 );
nand NAND2_26714 ( P2_R1957_U129 , P2_R1957_U86 , P2_R1957_U52 );
nand NAND2_26715 ( P2_R1957_U130 , P2_U3655 , P2_R1957_U23 );
nand NAND2_26716 ( P2_R1957_U131 , P2_R1957_U85 , P2_R1957_U54 );
nand NAND2_26717 ( P2_R1957_U132 , P2_U3657 , P2_R1957_U22 );
nand NAND2_26718 ( P2_R1957_U133 , P2_R1957_U84 , P2_R1957_U56 );
nand NAND2_26719 ( P2_R1957_U134 , P2_U3660 , P2_R1957_U21 );
nand NAND2_26720 ( P2_R1957_U135 , P2_R1957_U83 , P2_R1957_U58 );
nand NAND2_26721 ( P2_R1957_U136 , P2_R1957_U127 , P2_R1957_U60 );
nand NAND3_26722 ( P2_R1957_U137 , P2_R1957_U103 , P2_R1957_U61 , P2_U3647 );
nand NAND2_26723 ( P2_R1957_U138 , P2_U3659 , P2_R1957_U37 );
nand NAND2_26724 ( P2_R1957_U139 , P2_R1957_U103 , P2_R1957_U61 );
nand NAND2_26725 ( P2_R1957_U140 , P2_U3663 , P2_R1957_U35 );
nand NAND2_26726 ( P2_R1957_U141 , P2_R1957_U101 , P2_R1957_U63 );
nand NAND2_26727 ( P2_R1957_U142 , P2_U3665 , P2_R1957_U34 );
nand NAND2_26728 ( P2_R1957_U143 , P2_R1957_U100 , P2_R1957_U65 );
nand NAND2_26729 ( P2_R1957_U144 , P2_U3667 , P2_R1957_U33 );
nand NAND2_26730 ( P2_R1957_U145 , P2_R1957_U99 , P2_R1957_U67 );
nand NAND2_26731 ( P2_R1957_U146 , P2_U3669 , P2_R1957_U32 );
nand NAND2_26732 ( P2_R1957_U147 , P2_R1957_U98 , P2_R1957_U69 );
nand NAND2_26733 ( P2_R1957_U148 , P2_U3682 , P2_R1957_U72 );
nand NAND2_26734 ( P2_R1957_U149 , P2_U3683 , P2_R1957_U71 );
nand NAND2_26735 ( P2_R1957_U150 , P2_U3672 , P2_R1957_U31 );
nand NAND2_26736 ( P2_R1957_U151 , P2_R1957_U97 , P2_R1957_U73 );
nand NAND2_26737 ( P2_R1957_U152 , P2_U3674 , P2_R1957_U30 );
nand NAND2_26738 ( P2_R1957_U153 , P2_R1957_U96 , P2_R1957_U75 );
nand NAND2_26739 ( P2_R1957_U154 , P2_U3676 , P2_R1957_U29 );
nand NAND2_26740 ( P2_R1957_U155 , P2_R1957_U95 , P2_R1957_U77 );
nand NAND2_26741 ( P2_R1957_U156 , P2_U3678 , P2_R1957_U28 );
nand NAND2_26742 ( P2_R1957_U157 , P2_R1957_U94 , P2_R1957_U79 );
nand NAND2_26743 ( P2_R1957_U158 , P2_U3680 , P2_R1957_U27 );
nand NAND2_26744 ( P2_R1957_U159 , P2_R1957_U93 , P2_R1957_U81 );
and AND2_26745 ( P2_R2278_U4 , P2_R2278_U399 , P2_R2278_U398 );
and AND3_26746 ( P2_R2278_U5 , P2_R2278_U161 , P2_R2278_U309 , P2_R2278_U206 );
nand NAND3_26747 ( P2_R2278_U6 , P2_R2278_U490 , P2_R2278_U489 , P2_R2278_U345 );
not NOT1_26748 ( P2_R2278_U7 , P2_U3631 );
not NOT1_26749 ( P2_R2278_U8 , P2_INSTADDRPOINTER_REG_7_ );
not NOT1_26750 ( P2_R2278_U9 , P2_U3633 );
not NOT1_26751 ( P2_R2278_U10 , P2_INSTADDRPOINTER_REG_5_ );
not NOT1_26752 ( P2_R2278_U11 , P2_U3635 );
not NOT1_26753 ( P2_R2278_U12 , P2_INSTADDRPOINTER_REG_3_ );
not NOT1_26754 ( P2_R2278_U13 , P2_U3638 );
not NOT1_26755 ( P2_R2278_U14 , P2_INSTADDRPOINTER_REG_0_ );
nand NAND2_26756 ( P2_R2278_U15 , P2_INSTADDRPOINTER_REG_0_ , P2_U3638 );
not NOT1_26757 ( P2_R2278_U16 , P2_U3637 );
not NOT1_26758 ( P2_R2278_U17 , P2_INSTADDRPOINTER_REG_1_ );
not NOT1_26759 ( P2_R2278_U18 , P2_U3636 );
not NOT1_26760 ( P2_R2278_U19 , P2_INSTADDRPOINTER_REG_2_ );
nand NAND2_26761 ( P2_R2278_U20 , P2_INSTADDRPOINTER_REG_2_ , P2_U3636 );
not NOT1_26762 ( P2_R2278_U21 , P2_U3634 );
not NOT1_26763 ( P2_R2278_U22 , P2_INSTADDRPOINTER_REG_4_ );
nand NAND2_26764 ( P2_R2278_U23 , P2_INSTADDRPOINTER_REG_4_ , P2_U3634 );
not NOT1_26765 ( P2_R2278_U24 , P2_U3632 );
not NOT1_26766 ( P2_R2278_U25 , P2_INSTADDRPOINTER_REG_6_ );
nand NAND2_26767 ( P2_R2278_U26 , P2_INSTADDRPOINTER_REG_6_ , P2_U3632 );
not NOT1_26768 ( P2_R2278_U27 , P2_U3630 );
not NOT1_26769 ( P2_R2278_U28 , P2_INSTADDRPOINTER_REG_8_ );
not NOT1_26770 ( P2_R2278_U29 , P2_INSTADDRPOINTER_REG_9_ );
not NOT1_26771 ( P2_R2278_U30 , P2_U2812 );
not NOT1_26772 ( P2_R2278_U31 , P2_U2793 );
not NOT1_26773 ( P2_R2278_U32 , P2_INSTADDRPOINTER_REG_28_ );
not NOT1_26774 ( P2_R2278_U33 , P2_U2792 );
not NOT1_26775 ( P2_R2278_U34 , P2_INSTADDRPOINTER_REG_29_ );
not NOT1_26776 ( P2_R2278_U35 , P2_U2797 );
not NOT1_26777 ( P2_R2278_U36 , P2_INSTADDRPOINTER_REG_24_ );
not NOT1_26778 ( P2_R2278_U37 , P2_U2799 );
not NOT1_26779 ( P2_R2278_U38 , P2_INSTADDRPOINTER_REG_22_ );
not NOT1_26780 ( P2_R2278_U39 , P2_U2801 );
not NOT1_26781 ( P2_R2278_U40 , P2_INSTADDRPOINTER_REG_20_ );
not NOT1_26782 ( P2_R2278_U41 , P2_U2804 );
not NOT1_26783 ( P2_R2278_U42 , P2_INSTADDRPOINTER_REG_17_ );
not NOT1_26784 ( P2_R2278_U43 , P2_U2806 );
not NOT1_26785 ( P2_R2278_U44 , P2_INSTADDRPOINTER_REG_15_ );
not NOT1_26786 ( P2_R2278_U45 , P2_U2808 );
not NOT1_26787 ( P2_R2278_U46 , P2_INSTADDRPOINTER_REG_13_ );
not NOT1_26788 ( P2_R2278_U47 , P2_U2810 );
not NOT1_26789 ( P2_R2278_U48 , P2_INSTADDRPOINTER_REG_11_ );
nand NAND2_26790 ( P2_R2278_U49 , P2_INSTADDRPOINTER_REG_8_ , P2_U3630 );
not NOT1_26791 ( P2_R2278_U50 , P2_U2811 );
not NOT1_26792 ( P2_R2278_U51 , P2_INSTADDRPOINTER_REG_10_ );
nand NAND2_26793 ( P2_R2278_U52 , P2_INSTADDRPOINTER_REG_10_ , P2_U2811 );
not NOT1_26794 ( P2_R2278_U53 , P2_U2809 );
not NOT1_26795 ( P2_R2278_U54 , P2_INSTADDRPOINTER_REG_12_ );
nand NAND2_26796 ( P2_R2278_U55 , P2_INSTADDRPOINTER_REG_12_ , P2_U2809 );
not NOT1_26797 ( P2_R2278_U56 , P2_U2807 );
not NOT1_26798 ( P2_R2278_U57 , P2_INSTADDRPOINTER_REG_14_ );
nand NAND2_26799 ( P2_R2278_U58 , P2_INSTADDRPOINTER_REG_14_ , P2_U2807 );
not NOT1_26800 ( P2_R2278_U59 , P2_U2805 );
not NOT1_26801 ( P2_R2278_U60 , P2_INSTADDRPOINTER_REG_16_ );
nand NAND2_26802 ( P2_R2278_U61 , P2_INSTADDRPOINTER_REG_16_ , P2_U2805 );
not NOT1_26803 ( P2_R2278_U62 , P2_U2802 );
not NOT1_26804 ( P2_R2278_U63 , P2_INSTADDRPOINTER_REG_19_ );
not NOT1_26805 ( P2_R2278_U64 , P2_U2803 );
not NOT1_26806 ( P2_R2278_U65 , P2_INSTADDRPOINTER_REG_18_ );
not NOT1_26807 ( P2_R2278_U66 , P2_U2800 );
not NOT1_26808 ( P2_R2278_U67 , P2_INSTADDRPOINTER_REG_21_ );
nand NAND2_26809 ( P2_R2278_U68 , P2_INSTADDRPOINTER_REG_21_ , P2_U2800 );
not NOT1_26810 ( P2_R2278_U69 , P2_U2798 );
not NOT1_26811 ( P2_R2278_U70 , P2_INSTADDRPOINTER_REG_23_ );
nand NAND2_26812 ( P2_R2278_U71 , P2_INSTADDRPOINTER_REG_23_ , P2_U2798 );
not NOT1_26813 ( P2_R2278_U72 , P2_U2796 );
not NOT1_26814 ( P2_R2278_U73 , P2_INSTADDRPOINTER_REG_25_ );
not NOT1_26815 ( P2_R2278_U74 , P2_U2794 );
not NOT1_26816 ( P2_R2278_U75 , P2_INSTADDRPOINTER_REG_27_ );
not NOT1_26817 ( P2_R2278_U76 , P2_U2795 );
not NOT1_26818 ( P2_R2278_U77 , P2_INSTADDRPOINTER_REG_26_ );
nand NAND2_26819 ( P2_R2278_U78 , P2_INSTADDRPOINTER_REG_26_ , P2_U2795 );
not NOT1_26820 ( P2_R2278_U79 , P2_U2791 );
not NOT1_26821 ( P2_R2278_U80 , P2_INSTADDRPOINTER_REG_30_ );
nand NAND2_26822 ( P2_R2278_U81 , P2_R2278_U340 , P2_R2278_U297 );
nand NAND2_26823 ( P2_R2278_U82 , P2_U3637 , P2_R2278_U208 );
nand NAND2_26824 ( P2_R2278_U83 , P2_R2278_U562 , P2_R2278_U561 );
nand NAND2_26825 ( P2_R2278_U84 , P2_R2278_U352 , P2_R2278_U351 );
nand NAND2_26826 ( P2_R2278_U85 , P2_R2278_U359 , P2_R2278_U358 );
nand NAND2_26827 ( P2_R2278_U86 , P2_R2278_U366 , P2_R2278_U365 );
nand NAND2_26828 ( P2_R2278_U87 , P2_R2278_U373 , P2_R2278_U372 );
nand NAND2_26829 ( P2_R2278_U88 , P2_R2278_U380 , P2_R2278_U379 );
nand NAND2_26830 ( P2_R2278_U89 , P2_R2278_U387 , P2_R2278_U386 );
nand NAND2_26831 ( P2_R2278_U90 , P2_R2278_U394 , P2_R2278_U393 );
nand NAND2_26832 ( P2_R2278_U91 , P2_R2278_U408 , P2_R2278_U407 );
nand NAND2_26833 ( P2_R2278_U92 , P2_R2278_U415 , P2_R2278_U414 );
nand NAND2_26834 ( P2_R2278_U93 , P2_R2278_U422 , P2_R2278_U421 );
nand NAND2_26835 ( P2_R2278_U94 , P2_R2278_U429 , P2_R2278_U428 );
nand NAND2_26836 ( P2_R2278_U95 , P2_R2278_U436 , P2_R2278_U435 );
nand NAND2_26837 ( P2_R2278_U96 , P2_R2278_U443 , P2_R2278_U442 );
nand NAND2_26838 ( P2_R2278_U97 , P2_R2278_U450 , P2_R2278_U449 );
nand NAND2_26839 ( P2_R2278_U98 , P2_R2278_U457 , P2_R2278_U456 );
nand NAND2_26840 ( P2_R2278_U99 , P2_R2278_U464 , P2_R2278_U463 );
nand NAND2_26841 ( P2_R2278_U100 , P2_R2278_U471 , P2_R2278_U470 );
nand NAND2_26842 ( P2_R2278_U101 , P2_R2278_U478 , P2_R2278_U477 );
nand NAND2_26843 ( P2_R2278_U102 , P2_R2278_U485 , P2_R2278_U484 );
nand NAND2_26844 ( P2_R2278_U103 , P2_R2278_U497 , P2_R2278_U496 );
nand NAND2_26845 ( P2_R2278_U104 , P2_R2278_U504 , P2_R2278_U503 );
nand NAND2_26846 ( P2_R2278_U105 , P2_R2278_U511 , P2_R2278_U510 );
nand NAND2_26847 ( P2_R2278_U106 , P2_R2278_U518 , P2_R2278_U517 );
nand NAND2_26848 ( P2_R2278_U107 , P2_R2278_U525 , P2_R2278_U524 );
nand NAND2_26849 ( P2_R2278_U108 , P2_R2278_U532 , P2_R2278_U531 );
nand NAND2_26850 ( P2_R2278_U109 , P2_R2278_U539 , P2_R2278_U538 );
nand NAND2_26851 ( P2_R2278_U110 , P2_R2278_U546 , P2_R2278_U545 );
nand NAND2_26852 ( P2_R2278_U111 , P2_R2278_U553 , P2_R2278_U552 );
nand NAND2_26853 ( P2_R2278_U112 , P2_R2278_U560 , P2_R2278_U559 );
and AND2_26854 ( P2_R2278_U113 , P2_R2278_U210 , P2_R2278_U314 );
and AND2_26855 ( P2_R2278_U114 , P2_R2278_U313 , P2_R2278_U215 );
and AND2_26856 ( P2_R2278_U115 , P2_R2278_U217 , P2_R2278_U221 );
and AND2_26857 ( P2_R2278_U116 , P2_R2278_U316 , P2_R2278_U222 );
and AND2_26858 ( P2_R2278_U117 , P2_R2278_U224 , P2_R2278_U228 );
and AND2_26859 ( P2_R2278_U118 , P2_R2278_U318 , P2_R2278_U229 );
and AND2_26860 ( P2_R2278_U119 , P2_R2278_U231 , P2_R2278_U235 );
and AND2_26861 ( P2_R2278_U120 , P2_R2278_U320 , P2_R2278_U236 );
and AND2_26862 ( P2_R2278_U121 , P2_R2278_U238 , P2_R2278_U242 );
and AND2_26863 ( P2_R2278_U122 , P2_R2278_U322 , P2_R2278_U243 );
and AND2_26864 ( P2_R2278_U123 , P2_R2278_U245 , P2_R2278_U249 );
and AND2_26865 ( P2_R2278_U124 , P2_R2278_U324 , P2_R2278_U250 );
and AND2_26866 ( P2_R2278_U125 , P2_R2278_U252 , P2_R2278_U256 );
and AND2_26867 ( P2_R2278_U126 , P2_R2278_U326 , P2_R2278_U257 );
and AND2_26868 ( P2_R2278_U127 , P2_R2278_U259 , P2_R2278_U263 );
and AND2_26869 ( P2_R2278_U128 , P2_R2278_U328 , P2_R2278_U264 );
and AND2_26870 ( P2_R2278_U129 , P2_R2278_U273 , P2_R2278_U270 );
and AND2_26871 ( P2_R2278_U130 , P2_R2278_U331 , P2_R2278_U273 );
and AND2_26872 ( P2_R2278_U131 , P2_R2278_U334 , P2_R2278_U274 );
and AND2_26873 ( P2_R2278_U132 , P2_R2278_U276 , P2_R2278_U280 );
and AND2_26874 ( P2_R2278_U133 , P2_R2278_U336 , P2_R2278_U281 );
and AND2_26875 ( P2_R2278_U134 , P2_R2278_U283 , P2_R2278_U287 );
and AND2_26876 ( P2_R2278_U135 , P2_R2278_U338 , P2_R2278_U288 );
and AND3_26877 ( P2_R2278_U136 , P2_R2278_U299 , P2_R2278_U296 , P2_R2278_U292 );
and AND2_26878 ( P2_R2278_U137 , P2_R2278_U304 , P2_R2278_U300 );
and AND2_26879 ( P2_R2278_U138 , P2_R2278_U307 , P2_R2278_U302 );
and AND2_26880 ( P2_R2278_U139 , P2_R2278_U397 , P2_R2278_U138 );
and AND2_26881 ( P2_R2278_U140 , P2_R2278_U343 , P2_R2278_U300 );
and AND2_26882 ( P2_R2278_U141 , P2_R2278_U4 , P2_R2278_U142 );
and AND2_26883 ( P2_R2278_U142 , P2_R2278_U304 , P2_R2278_U306 );
and AND2_26884 ( P2_R2278_U143 , P2_R2278_U292 , P2_R2278_U296 );
and AND2_26885 ( P2_R2278_U144 , P2_R2278_U266 , P2_R2278_U270 );
and AND2_26886 ( P2_R2278_U145 , P2_R2278_U347 , P2_R2278_U346 );
nand NAND2_26887 ( P2_R2278_U146 , P2_R2278_U49 , P2_R2278_U232 );
and AND2_26888 ( P2_R2278_U147 , P2_R2278_U354 , P2_R2278_U353 );
nand NAND2_26889 ( P2_R2278_U148 , P2_R2278_U118 , P2_R2278_U317 );
and AND2_26890 ( P2_R2278_U149 , P2_R2278_U361 , P2_R2278_U360 );
nand NAND2_26891 ( P2_R2278_U150 , P2_R2278_U26 , P2_R2278_U225 );
and AND2_26892 ( P2_R2278_U151 , P2_R2278_U368 , P2_R2278_U367 );
nand NAND2_26893 ( P2_R2278_U152 , P2_R2278_U116 , P2_R2278_U315 );
and AND2_26894 ( P2_R2278_U153 , P2_R2278_U375 , P2_R2278_U374 );
nand NAND2_26895 ( P2_R2278_U154 , P2_R2278_U23 , P2_R2278_U218 );
and AND2_26896 ( P2_R2278_U155 , P2_R2278_U382 , P2_R2278_U381 );
nand NAND2_26897 ( P2_R2278_U156 , P2_R2278_U114 , P2_R2278_U312 );
and AND2_26898 ( P2_R2278_U157 , P2_R2278_U389 , P2_R2278_U388 );
nand NAND2_26899 ( P2_R2278_U158 , P2_R2278_U20 , P2_R2278_U211 );
not NOT1_26900 ( P2_R2278_U159 , P2_INSTADDRPOINTER_REG_31_ );
not NOT1_26901 ( P2_R2278_U160 , P2_U2790 );
and AND2_26902 ( P2_R2278_U161 , P2_R2278_U401 , P2_R2278_U400 );
and AND2_26903 ( P2_R2278_U162 , P2_R2278_U403 , P2_R2278_U402 );
nand NAND2_26904 ( P2_R2278_U163 , P2_R2278_U304 , P2_R2278_U303 );
and AND2_26905 ( P2_R2278_U164 , P2_R2278_U410 , P2_R2278_U409 );
nand NAND3_26906 ( P2_R2278_U165 , P2_R2278_U310 , P2_R2278_U82 , P2_R2278_U311 );
and AND2_26907 ( P2_R2278_U166 , P2_R2278_U417 , P2_R2278_U416 );
nand NAND2_26908 ( P2_R2278_U167 , P2_R2278_U140 , P2_R2278_U342 );
and AND2_26909 ( P2_R2278_U168 , P2_R2278_U424 , P2_R2278_U423 );
nand NAND2_26910 ( P2_R2278_U169 , P2_R2278_U341 , P2_R2278_U339 );
and AND2_26911 ( P2_R2278_U170 , P2_R2278_U431 , P2_R2278_U430 );
nand NAND2_26912 ( P2_R2278_U171 , P2_R2278_U78 , P2_R2278_U293 );
and AND2_26913 ( P2_R2278_U172 , P2_R2278_U438 , P2_R2278_U437 );
nand NAND3_26914 ( P2_R2278_U173 , P2_R2278_U290 , P2_R2278_U205 , P2_R2278_U308 );
nand NAND2_26915 ( P2_R2278_U174 , P2_R2278_U135 , P2_R2278_U337 );
and AND2_26916 ( P2_R2278_U175 , P2_R2278_U452 , P2_R2278_U451 );
nand NAND2_26917 ( P2_R2278_U176 , P2_R2278_U71 , P2_R2278_U284 );
and AND2_26918 ( P2_R2278_U177 , P2_R2278_U459 , P2_R2278_U458 );
nand NAND2_26919 ( P2_R2278_U178 , P2_R2278_U133 , P2_R2278_U335 );
and AND2_26920 ( P2_R2278_U179 , P2_R2278_U466 , P2_R2278_U465 );
nand NAND2_26921 ( P2_R2278_U180 , P2_R2278_U68 , P2_R2278_U277 );
and AND2_26922 ( P2_R2278_U181 , P2_R2278_U473 , P2_R2278_U472 );
nand NAND2_26923 ( P2_R2278_U182 , P2_R2278_U131 , P2_R2278_U333 );
and AND2_26924 ( P2_R2278_U183 , P2_R2278_U480 , P2_R2278_U479 );
nand NAND2_26925 ( P2_R2278_U184 , P2_R2278_U330 , P2_R2278_U329 );
and AND2_26926 ( P2_R2278_U185 , P2_R2278_U492 , P2_R2278_U491 );
nand NAND2_26927 ( P2_R2278_U186 , P2_R2278_U268 , P2_R2278_U267 );
and AND2_26928 ( P2_R2278_U187 , P2_R2278_U499 , P2_R2278_U498 );
nand NAND2_26929 ( P2_R2278_U188 , P2_R2278_U128 , P2_R2278_U327 );
and AND2_26930 ( P2_R2278_U189 , P2_R2278_U506 , P2_R2278_U505 );
nand NAND2_26931 ( P2_R2278_U190 , P2_R2278_U61 , P2_R2278_U260 );
and AND2_26932 ( P2_R2278_U191 , P2_R2278_U513 , P2_R2278_U512 );
nand NAND2_26933 ( P2_R2278_U192 , P2_R2278_U126 , P2_R2278_U325 );
and AND2_26934 ( P2_R2278_U193 , P2_R2278_U520 , P2_R2278_U519 );
nand NAND2_26935 ( P2_R2278_U194 , P2_R2278_U58 , P2_R2278_U253 );
and AND2_26936 ( P2_R2278_U195 , P2_R2278_U527 , P2_R2278_U526 );
nand NAND2_26937 ( P2_R2278_U196 , P2_R2278_U124 , P2_R2278_U323 );
and AND2_26938 ( P2_R2278_U197 , P2_R2278_U534 , P2_R2278_U533 );
nand NAND2_26939 ( P2_R2278_U198 , P2_R2278_U55 , P2_R2278_U246 );
and AND2_26940 ( P2_R2278_U199 , P2_R2278_U541 , P2_R2278_U540 );
nand NAND2_26941 ( P2_R2278_U200 , P2_R2278_U122 , P2_R2278_U321 );
and AND2_26942 ( P2_R2278_U201 , P2_R2278_U548 , P2_R2278_U547 );
nand NAND2_26943 ( P2_R2278_U202 , P2_R2278_U52 , P2_R2278_U239 );
and AND2_26944 ( P2_R2278_U203 , P2_R2278_U555 , P2_R2278_U554 );
nand NAND2_26945 ( P2_R2278_U204 , P2_R2278_U120 , P2_R2278_U319 );
nand NAND2_26946 ( P2_R2278_U205 , P2_U2796 , P2_R2278_U174 );
nand NAND2_26947 ( P2_R2278_U206 , P2_R2278_U139 , P2_R2278_U344 );
not NOT1_26948 ( P2_R2278_U207 , P2_R2278_U82 );
not NOT1_26949 ( P2_R2278_U208 , P2_R2278_U15 );
not NOT1_26950 ( P2_R2278_U209 , P2_R2278_U165 );
or OR2_26951 ( P2_R2278_U210 , P2_U3636 , P2_INSTADDRPOINTER_REG_2_ );
nand NAND2_26952 ( P2_R2278_U211 , P2_R2278_U210 , P2_R2278_U165 );
not NOT1_26953 ( P2_R2278_U212 , P2_R2278_U20 );
not NOT1_26954 ( P2_R2278_U213 , P2_R2278_U158 );
or OR2_26955 ( P2_R2278_U214 , P2_U3635 , P2_INSTADDRPOINTER_REG_3_ );
nand NAND2_26956 ( P2_R2278_U215 , P2_INSTADDRPOINTER_REG_3_ , P2_U3635 );
not NOT1_26957 ( P2_R2278_U216 , P2_R2278_U156 );
or OR2_26958 ( P2_R2278_U217 , P2_U3634 , P2_INSTADDRPOINTER_REG_4_ );
nand NAND2_26959 ( P2_R2278_U218 , P2_R2278_U217 , P2_R2278_U156 );
not NOT1_26960 ( P2_R2278_U219 , P2_R2278_U23 );
not NOT1_26961 ( P2_R2278_U220 , P2_R2278_U154 );
or OR2_26962 ( P2_R2278_U221 , P2_U3633 , P2_INSTADDRPOINTER_REG_5_ );
nand NAND2_26963 ( P2_R2278_U222 , P2_INSTADDRPOINTER_REG_5_ , P2_U3633 );
not NOT1_26964 ( P2_R2278_U223 , P2_R2278_U152 );
or OR2_26965 ( P2_R2278_U224 , P2_U3632 , P2_INSTADDRPOINTER_REG_6_ );
nand NAND2_26966 ( P2_R2278_U225 , P2_R2278_U224 , P2_R2278_U152 );
not NOT1_26967 ( P2_R2278_U226 , P2_R2278_U26 );
not NOT1_26968 ( P2_R2278_U227 , P2_R2278_U150 );
or OR2_26969 ( P2_R2278_U228 , P2_U3631 , P2_INSTADDRPOINTER_REG_7_ );
nand NAND2_26970 ( P2_R2278_U229 , P2_INSTADDRPOINTER_REG_7_ , P2_U3631 );
not NOT1_26971 ( P2_R2278_U230 , P2_R2278_U148 );
or OR2_26972 ( P2_R2278_U231 , P2_U3630 , P2_INSTADDRPOINTER_REG_8_ );
nand NAND2_26973 ( P2_R2278_U232 , P2_R2278_U231 , P2_R2278_U148 );
not NOT1_26974 ( P2_R2278_U233 , P2_R2278_U49 );
not NOT1_26975 ( P2_R2278_U234 , P2_R2278_U146 );
or OR2_26976 ( P2_R2278_U235 , P2_U2812 , P2_INSTADDRPOINTER_REG_9_ );
nand NAND2_26977 ( P2_R2278_U236 , P2_U2812 , P2_INSTADDRPOINTER_REG_9_ );
not NOT1_26978 ( P2_R2278_U237 , P2_R2278_U204 );
or OR2_26979 ( P2_R2278_U238 , P2_U2811 , P2_INSTADDRPOINTER_REG_10_ );
nand NAND2_26980 ( P2_R2278_U239 , P2_R2278_U238 , P2_R2278_U204 );
not NOT1_26981 ( P2_R2278_U240 , P2_R2278_U52 );
not NOT1_26982 ( P2_R2278_U241 , P2_R2278_U202 );
or OR2_26983 ( P2_R2278_U242 , P2_U2810 , P2_INSTADDRPOINTER_REG_11_ );
nand NAND2_26984 ( P2_R2278_U243 , P2_INSTADDRPOINTER_REG_11_ , P2_U2810 );
not NOT1_26985 ( P2_R2278_U244 , P2_R2278_U200 );
or OR2_26986 ( P2_R2278_U245 , P2_U2809 , P2_INSTADDRPOINTER_REG_12_ );
nand NAND2_26987 ( P2_R2278_U246 , P2_R2278_U245 , P2_R2278_U200 );
not NOT1_26988 ( P2_R2278_U247 , P2_R2278_U55 );
not NOT1_26989 ( P2_R2278_U248 , P2_R2278_U198 );
or OR2_26990 ( P2_R2278_U249 , P2_U2808 , P2_INSTADDRPOINTER_REG_13_ );
nand NAND2_26991 ( P2_R2278_U250 , P2_INSTADDRPOINTER_REG_13_ , P2_U2808 );
not NOT1_26992 ( P2_R2278_U251 , P2_R2278_U196 );
or OR2_26993 ( P2_R2278_U252 , P2_U2807 , P2_INSTADDRPOINTER_REG_14_ );
nand NAND2_26994 ( P2_R2278_U253 , P2_R2278_U252 , P2_R2278_U196 );
not NOT1_26995 ( P2_R2278_U254 , P2_R2278_U58 );
not NOT1_26996 ( P2_R2278_U255 , P2_R2278_U194 );
or OR2_26997 ( P2_R2278_U256 , P2_U2806 , P2_INSTADDRPOINTER_REG_15_ );
nand NAND2_26998 ( P2_R2278_U257 , P2_INSTADDRPOINTER_REG_15_ , P2_U2806 );
not NOT1_26999 ( P2_R2278_U258 , P2_R2278_U192 );
or OR2_27000 ( P2_R2278_U259 , P2_U2805 , P2_INSTADDRPOINTER_REG_16_ );
nand NAND2_27001 ( P2_R2278_U260 , P2_R2278_U259 , P2_R2278_U192 );
not NOT1_27002 ( P2_R2278_U261 , P2_R2278_U61 );
not NOT1_27003 ( P2_R2278_U262 , P2_R2278_U190 );
or OR2_27004 ( P2_R2278_U263 , P2_U2804 , P2_INSTADDRPOINTER_REG_17_ );
nand NAND2_27005 ( P2_R2278_U264 , P2_INSTADDRPOINTER_REG_17_ , P2_U2804 );
not NOT1_27006 ( P2_R2278_U265 , P2_R2278_U188 );
or OR2_27007 ( P2_R2278_U266 , P2_U2803 , P2_INSTADDRPOINTER_REG_18_ );
nand NAND2_27008 ( P2_R2278_U267 , P2_R2278_U266 , P2_R2278_U188 );
nand NAND2_27009 ( P2_R2278_U268 , P2_INSTADDRPOINTER_REG_18_ , P2_U2803 );
not NOT1_27010 ( P2_R2278_U269 , P2_R2278_U186 );
or OR2_27011 ( P2_R2278_U270 , P2_U2802 , P2_INSTADDRPOINTER_REG_19_ );
nand NAND2_27012 ( P2_R2278_U271 , P2_INSTADDRPOINTER_REG_19_ , P2_U2802 );
not NOT1_27013 ( P2_R2278_U272 , P2_R2278_U184 );
or OR2_27014 ( P2_R2278_U273 , P2_U2801 , P2_INSTADDRPOINTER_REG_20_ );
nand NAND2_27015 ( P2_R2278_U274 , P2_INSTADDRPOINTER_REG_20_ , P2_U2801 );
not NOT1_27016 ( P2_R2278_U275 , P2_R2278_U182 );
or OR2_27017 ( P2_R2278_U276 , P2_U2800 , P2_INSTADDRPOINTER_REG_21_ );
nand NAND2_27018 ( P2_R2278_U277 , P2_R2278_U276 , P2_R2278_U182 );
not NOT1_27019 ( P2_R2278_U278 , P2_R2278_U68 );
not NOT1_27020 ( P2_R2278_U279 , P2_R2278_U180 );
or OR2_27021 ( P2_R2278_U280 , P2_U2799 , P2_INSTADDRPOINTER_REG_22_ );
nand NAND2_27022 ( P2_R2278_U281 , P2_INSTADDRPOINTER_REG_22_ , P2_U2799 );
not NOT1_27023 ( P2_R2278_U282 , P2_R2278_U178 );
or OR2_27024 ( P2_R2278_U283 , P2_U2798 , P2_INSTADDRPOINTER_REG_23_ );
nand NAND2_27025 ( P2_R2278_U284 , P2_R2278_U283 , P2_R2278_U178 );
not NOT1_27026 ( P2_R2278_U285 , P2_R2278_U71 );
not NOT1_27027 ( P2_R2278_U286 , P2_R2278_U176 );
or OR2_27028 ( P2_R2278_U287 , P2_U2797 , P2_INSTADDRPOINTER_REG_24_ );
nand NAND2_27029 ( P2_R2278_U288 , P2_INSTADDRPOINTER_REG_24_ , P2_U2797 );
not NOT1_27030 ( P2_R2278_U289 , P2_R2278_U174 );
nand NAND2_27031 ( P2_R2278_U290 , P2_INSTADDRPOINTER_REG_25_ , P2_R2278_U174 );
not NOT1_27032 ( P2_R2278_U291 , P2_R2278_U173 );
or OR2_27033 ( P2_R2278_U292 , P2_U2795 , P2_INSTADDRPOINTER_REG_26_ );
nand NAND2_27034 ( P2_R2278_U293 , P2_R2278_U292 , P2_R2278_U173 );
not NOT1_27035 ( P2_R2278_U294 , P2_R2278_U78 );
not NOT1_27036 ( P2_R2278_U295 , P2_R2278_U171 );
or OR2_27037 ( P2_R2278_U296 , P2_U2794 , P2_INSTADDRPOINTER_REG_27_ );
nand NAND2_27038 ( P2_R2278_U297 , P2_INSTADDRPOINTER_REG_27_ , P2_U2794 );
not NOT1_27039 ( P2_R2278_U298 , P2_R2278_U169 );
or OR2_27040 ( P2_R2278_U299 , P2_U2793 , P2_INSTADDRPOINTER_REG_28_ );
nand NAND2_27041 ( P2_R2278_U300 , P2_INSTADDRPOINTER_REG_28_ , P2_U2793 );
not NOT1_27042 ( P2_R2278_U301 , P2_R2278_U167 );
or OR2_27043 ( P2_R2278_U302 , P2_U2792 , P2_INSTADDRPOINTER_REG_29_ );
nand NAND2_27044 ( P2_R2278_U303 , P2_R2278_U302 , P2_R2278_U167 );
nand NAND2_27045 ( P2_R2278_U304 , P2_INSTADDRPOINTER_REG_29_ , P2_U2792 );
not NOT1_27046 ( P2_R2278_U305 , P2_R2278_U163 );
nand NAND2_27047 ( P2_R2278_U306 , P2_INSTADDRPOINTER_REG_30_ , P2_U2791 );
or OR2_27048 ( P2_R2278_U307 , P2_INSTADDRPOINTER_REG_30_ , P2_U2791 );
nand NAND2_27049 ( P2_R2278_U308 , P2_INSTADDRPOINTER_REG_25_ , P2_U2796 );
nand NAND2_27050 ( P2_R2278_U309 , P2_R2278_U303 , P2_R2278_U141 );
nand NAND2_27051 ( P2_R2278_U310 , P2_INSTADDRPOINTER_REG_1_ , P2_R2278_U208 );
nand NAND2_27052 ( P2_R2278_U311 , P2_INSTADDRPOINTER_REG_1_ , P2_U3637 );
nand NAND2_27053 ( P2_R2278_U312 , P2_R2278_U113 , P2_R2278_U165 );
nand NAND2_27054 ( P2_R2278_U313 , P2_R2278_U212 , P2_R2278_U214 );
or OR2_27055 ( P2_R2278_U314 , P2_U3635 , P2_INSTADDRPOINTER_REG_3_ );
nand NAND2_27056 ( P2_R2278_U315 , P2_R2278_U115 , P2_R2278_U156 );
nand NAND2_27057 ( P2_R2278_U316 , P2_R2278_U219 , P2_R2278_U221 );
nand NAND2_27058 ( P2_R2278_U317 , P2_R2278_U117 , P2_R2278_U152 );
nand NAND2_27059 ( P2_R2278_U318 , P2_R2278_U226 , P2_R2278_U228 );
nand NAND2_27060 ( P2_R2278_U319 , P2_R2278_U119 , P2_R2278_U148 );
nand NAND2_27061 ( P2_R2278_U320 , P2_R2278_U233 , P2_R2278_U235 );
nand NAND2_27062 ( P2_R2278_U321 , P2_R2278_U121 , P2_R2278_U204 );
nand NAND2_27063 ( P2_R2278_U322 , P2_R2278_U240 , P2_R2278_U242 );
nand NAND2_27064 ( P2_R2278_U323 , P2_R2278_U123 , P2_R2278_U200 );
nand NAND2_27065 ( P2_R2278_U324 , P2_R2278_U247 , P2_R2278_U249 );
nand NAND2_27066 ( P2_R2278_U325 , P2_R2278_U125 , P2_R2278_U196 );
nand NAND2_27067 ( P2_R2278_U326 , P2_R2278_U254 , P2_R2278_U256 );
nand NAND2_27068 ( P2_R2278_U327 , P2_R2278_U127 , P2_R2278_U192 );
nand NAND2_27069 ( P2_R2278_U328 , P2_R2278_U261 , P2_R2278_U263 );
nand NAND2_27070 ( P2_R2278_U329 , P2_R2278_U144 , P2_R2278_U188 );
nand NAND2_27071 ( P2_R2278_U330 , P2_R2278_U331 , P2_R2278_U332 );
or OR2_27072 ( P2_R2278_U331 , P2_U2802 , P2_INSTADDRPOINTER_REG_19_ );
nand NAND2_27073 ( P2_R2278_U332 , P2_R2278_U268 , P2_R2278_U271 );
nand NAND3_27074 ( P2_R2278_U333 , P2_R2278_U266 , P2_R2278_U188 , P2_R2278_U129 );
nand NAND2_27075 ( P2_R2278_U334 , P2_R2278_U130 , P2_R2278_U332 );
nand NAND2_27076 ( P2_R2278_U335 , P2_R2278_U132 , P2_R2278_U182 );
nand NAND2_27077 ( P2_R2278_U336 , P2_R2278_U278 , P2_R2278_U280 );
nand NAND2_27078 ( P2_R2278_U337 , P2_R2278_U134 , P2_R2278_U178 );
nand NAND2_27079 ( P2_R2278_U338 , P2_R2278_U285 , P2_R2278_U287 );
nand NAND2_27080 ( P2_R2278_U339 , P2_R2278_U143 , P2_R2278_U173 );
nand NAND2_27081 ( P2_R2278_U340 , P2_R2278_U294 , P2_R2278_U296 );
not NOT1_27082 ( P2_R2278_U341 , P2_R2278_U81 );
nand NAND2_27083 ( P2_R2278_U342 , P2_R2278_U173 , P2_R2278_U136 );
nand NAND2_27084 ( P2_R2278_U343 , P2_R2278_U81 , P2_R2278_U299 );
nand NAND3_27085 ( P2_R2278_U344 , P2_R2278_U343 , P2_R2278_U342 , P2_R2278_U137 );
nand NAND2_27086 ( P2_R2278_U345 , P2_R2278_U207 , P2_INSTADDRPOINTER_REG_1_ );
nand NAND2_27087 ( P2_R2278_U346 , P2_INSTADDRPOINTER_REG_9_ , P2_R2278_U30 );
nand NAND2_27088 ( P2_R2278_U347 , P2_U2812 , P2_R2278_U29 );
nand NAND2_27089 ( P2_R2278_U348 , P2_INSTADDRPOINTER_REG_9_ , P2_R2278_U30 );
nand NAND2_27090 ( P2_R2278_U349 , P2_U2812 , P2_R2278_U29 );
nand NAND2_27091 ( P2_R2278_U350 , P2_R2278_U349 , P2_R2278_U348 );
nand NAND2_27092 ( P2_R2278_U351 , P2_R2278_U145 , P2_R2278_U146 );
nand NAND2_27093 ( P2_R2278_U352 , P2_R2278_U234 , P2_R2278_U350 );
nand NAND2_27094 ( P2_R2278_U353 , P2_INSTADDRPOINTER_REG_8_ , P2_R2278_U27 );
nand NAND2_27095 ( P2_R2278_U354 , P2_U3630 , P2_R2278_U28 );
nand NAND2_27096 ( P2_R2278_U355 , P2_INSTADDRPOINTER_REG_8_ , P2_R2278_U27 );
nand NAND2_27097 ( P2_R2278_U356 , P2_U3630 , P2_R2278_U28 );
nand NAND2_27098 ( P2_R2278_U357 , P2_R2278_U356 , P2_R2278_U355 );
nand NAND2_27099 ( P2_R2278_U358 , P2_R2278_U147 , P2_R2278_U148 );
nand NAND2_27100 ( P2_R2278_U359 , P2_R2278_U230 , P2_R2278_U357 );
nand NAND2_27101 ( P2_R2278_U360 , P2_INSTADDRPOINTER_REG_7_ , P2_R2278_U7 );
nand NAND2_27102 ( P2_R2278_U361 , P2_U3631 , P2_R2278_U8 );
nand NAND2_27103 ( P2_R2278_U362 , P2_INSTADDRPOINTER_REG_7_ , P2_R2278_U7 );
nand NAND2_27104 ( P2_R2278_U363 , P2_U3631 , P2_R2278_U8 );
nand NAND2_27105 ( P2_R2278_U364 , P2_R2278_U363 , P2_R2278_U362 );
nand NAND2_27106 ( P2_R2278_U365 , P2_R2278_U149 , P2_R2278_U150 );
nand NAND2_27107 ( P2_R2278_U366 , P2_R2278_U227 , P2_R2278_U364 );
nand NAND2_27108 ( P2_R2278_U367 , P2_INSTADDRPOINTER_REG_6_ , P2_R2278_U24 );
nand NAND2_27109 ( P2_R2278_U368 , P2_U3632 , P2_R2278_U25 );
nand NAND2_27110 ( P2_R2278_U369 , P2_INSTADDRPOINTER_REG_6_ , P2_R2278_U24 );
nand NAND2_27111 ( P2_R2278_U370 , P2_U3632 , P2_R2278_U25 );
nand NAND2_27112 ( P2_R2278_U371 , P2_R2278_U370 , P2_R2278_U369 );
nand NAND2_27113 ( P2_R2278_U372 , P2_R2278_U151 , P2_R2278_U152 );
nand NAND2_27114 ( P2_R2278_U373 , P2_R2278_U223 , P2_R2278_U371 );
nand NAND2_27115 ( P2_R2278_U374 , P2_INSTADDRPOINTER_REG_5_ , P2_R2278_U9 );
nand NAND2_27116 ( P2_R2278_U375 , P2_U3633 , P2_R2278_U10 );
nand NAND2_27117 ( P2_R2278_U376 , P2_INSTADDRPOINTER_REG_5_ , P2_R2278_U9 );
nand NAND2_27118 ( P2_R2278_U377 , P2_U3633 , P2_R2278_U10 );
nand NAND2_27119 ( P2_R2278_U378 , P2_R2278_U377 , P2_R2278_U376 );
nand NAND2_27120 ( P2_R2278_U379 , P2_R2278_U153 , P2_R2278_U154 );
nand NAND2_27121 ( P2_R2278_U380 , P2_R2278_U220 , P2_R2278_U378 );
nand NAND2_27122 ( P2_R2278_U381 , P2_INSTADDRPOINTER_REG_4_ , P2_R2278_U21 );
nand NAND2_27123 ( P2_R2278_U382 , P2_U3634 , P2_R2278_U22 );
nand NAND2_27124 ( P2_R2278_U383 , P2_INSTADDRPOINTER_REG_4_ , P2_R2278_U21 );
nand NAND2_27125 ( P2_R2278_U384 , P2_U3634 , P2_R2278_U22 );
nand NAND2_27126 ( P2_R2278_U385 , P2_R2278_U384 , P2_R2278_U383 );
nand NAND2_27127 ( P2_R2278_U386 , P2_R2278_U155 , P2_R2278_U156 );
nand NAND2_27128 ( P2_R2278_U387 , P2_R2278_U216 , P2_R2278_U385 );
nand NAND2_27129 ( P2_R2278_U388 , P2_INSTADDRPOINTER_REG_3_ , P2_R2278_U11 );
nand NAND2_27130 ( P2_R2278_U389 , P2_U3635 , P2_R2278_U12 );
nand NAND2_27131 ( P2_R2278_U390 , P2_INSTADDRPOINTER_REG_3_ , P2_R2278_U11 );
nand NAND2_27132 ( P2_R2278_U391 , P2_U3635 , P2_R2278_U12 );
nand NAND2_27133 ( P2_R2278_U392 , P2_R2278_U391 , P2_R2278_U390 );
nand NAND2_27134 ( P2_R2278_U393 , P2_R2278_U157 , P2_R2278_U158 );
nand NAND2_27135 ( P2_R2278_U394 , P2_R2278_U213 , P2_R2278_U392 );
nand NAND2_27136 ( P2_R2278_U395 , P2_INSTADDRPOINTER_REG_31_ , P2_R2278_U160 );
nand NAND2_27137 ( P2_R2278_U396 , P2_U2790 , P2_R2278_U159 );
nand NAND2_27138 ( P2_R2278_U397 , P2_R2278_U396 , P2_R2278_U395 );
nand NAND2_27139 ( P2_R2278_U398 , P2_INSTADDRPOINTER_REG_31_ , P2_R2278_U160 );
nand NAND2_27140 ( P2_R2278_U399 , P2_U2790 , P2_R2278_U159 );
nand NAND3_27141 ( P2_R2278_U400 , P2_R2278_U4 , P2_R2278_U79 , P2_R2278_U80 );
nand NAND3_27142 ( P2_R2278_U401 , P2_U2791 , P2_R2278_U397 , P2_INSTADDRPOINTER_REG_30_ );
nand NAND2_27143 ( P2_R2278_U402 , P2_INSTADDRPOINTER_REG_30_ , P2_R2278_U79 );
nand NAND2_27144 ( P2_R2278_U403 , P2_U2791 , P2_R2278_U80 );
nand NAND2_27145 ( P2_R2278_U404 , P2_INSTADDRPOINTER_REG_30_ , P2_R2278_U79 );
nand NAND2_27146 ( P2_R2278_U405 , P2_U2791 , P2_R2278_U80 );
nand NAND2_27147 ( P2_R2278_U406 , P2_R2278_U405 , P2_R2278_U404 );
nand NAND2_27148 ( P2_R2278_U407 , P2_R2278_U162 , P2_R2278_U163 );
nand NAND2_27149 ( P2_R2278_U408 , P2_R2278_U305 , P2_R2278_U406 );
nand NAND2_27150 ( P2_R2278_U409 , P2_INSTADDRPOINTER_REG_2_ , P2_R2278_U18 );
nand NAND2_27151 ( P2_R2278_U410 , P2_U3636 , P2_R2278_U19 );
nand NAND2_27152 ( P2_R2278_U411 , P2_INSTADDRPOINTER_REG_2_ , P2_R2278_U18 );
nand NAND2_27153 ( P2_R2278_U412 , P2_U3636 , P2_R2278_U19 );
nand NAND2_27154 ( P2_R2278_U413 , P2_R2278_U412 , P2_R2278_U411 );
nand NAND2_27155 ( P2_R2278_U414 , P2_R2278_U164 , P2_R2278_U165 );
nand NAND2_27156 ( P2_R2278_U415 , P2_R2278_U209 , P2_R2278_U413 );
nand NAND2_27157 ( P2_R2278_U416 , P2_INSTADDRPOINTER_REG_29_ , P2_R2278_U33 );
nand NAND2_27158 ( P2_R2278_U417 , P2_U2792 , P2_R2278_U34 );
nand NAND2_27159 ( P2_R2278_U418 , P2_INSTADDRPOINTER_REG_29_ , P2_R2278_U33 );
nand NAND2_27160 ( P2_R2278_U419 , P2_U2792 , P2_R2278_U34 );
nand NAND2_27161 ( P2_R2278_U420 , P2_R2278_U419 , P2_R2278_U418 );
nand NAND2_27162 ( P2_R2278_U421 , P2_R2278_U166 , P2_R2278_U167 );
nand NAND2_27163 ( P2_R2278_U422 , P2_R2278_U301 , P2_R2278_U420 );
nand NAND2_27164 ( P2_R2278_U423 , P2_INSTADDRPOINTER_REG_28_ , P2_R2278_U31 );
nand NAND2_27165 ( P2_R2278_U424 , P2_U2793 , P2_R2278_U32 );
nand NAND2_27166 ( P2_R2278_U425 , P2_INSTADDRPOINTER_REG_28_ , P2_R2278_U31 );
nand NAND2_27167 ( P2_R2278_U426 , P2_U2793 , P2_R2278_U32 );
nand NAND2_27168 ( P2_R2278_U427 , P2_R2278_U426 , P2_R2278_U425 );
nand NAND2_27169 ( P2_R2278_U428 , P2_R2278_U168 , P2_R2278_U169 );
nand NAND2_27170 ( P2_R2278_U429 , P2_R2278_U298 , P2_R2278_U427 );
nand NAND2_27171 ( P2_R2278_U430 , P2_INSTADDRPOINTER_REG_27_ , P2_R2278_U74 );
nand NAND2_27172 ( P2_R2278_U431 , P2_U2794 , P2_R2278_U75 );
nand NAND2_27173 ( P2_R2278_U432 , P2_INSTADDRPOINTER_REG_27_ , P2_R2278_U74 );
nand NAND2_27174 ( P2_R2278_U433 , P2_U2794 , P2_R2278_U75 );
nand NAND2_27175 ( P2_R2278_U434 , P2_R2278_U433 , P2_R2278_U432 );
nand NAND2_27176 ( P2_R2278_U435 , P2_R2278_U170 , P2_R2278_U171 );
nand NAND2_27177 ( P2_R2278_U436 , P2_R2278_U295 , P2_R2278_U434 );
nand NAND2_27178 ( P2_R2278_U437 , P2_INSTADDRPOINTER_REG_26_ , P2_R2278_U76 );
nand NAND2_27179 ( P2_R2278_U438 , P2_U2795 , P2_R2278_U77 );
nand NAND2_27180 ( P2_R2278_U439 , P2_INSTADDRPOINTER_REG_26_ , P2_R2278_U76 );
nand NAND2_27181 ( P2_R2278_U440 , P2_U2795 , P2_R2278_U77 );
nand NAND2_27182 ( P2_R2278_U441 , P2_R2278_U440 , P2_R2278_U439 );
nand NAND2_27183 ( P2_R2278_U442 , P2_R2278_U172 , P2_R2278_U173 );
nand NAND2_27184 ( P2_R2278_U443 , P2_R2278_U291 , P2_R2278_U441 );
nand NAND2_27185 ( P2_R2278_U444 , P2_INSTADDRPOINTER_REG_25_ , P2_R2278_U174 );
nand NAND2_27186 ( P2_R2278_U445 , P2_R2278_U289 , P2_R2278_U73 );
nand NAND2_27187 ( P2_R2278_U446 , P2_INSTADDRPOINTER_REG_25_ , P2_R2278_U174 );
nand NAND2_27188 ( P2_R2278_U447 , P2_R2278_U289 , P2_R2278_U73 );
nand NAND2_27189 ( P2_R2278_U448 , P2_R2278_U447 , P2_R2278_U446 );
nand NAND3_27190 ( P2_R2278_U449 , P2_R2278_U445 , P2_R2278_U444 , P2_R2278_U72 );
nand NAND2_27191 ( P2_R2278_U450 , P2_R2278_U448 , P2_U2796 );
nand NAND2_27192 ( P2_R2278_U451 , P2_INSTADDRPOINTER_REG_24_ , P2_R2278_U35 );
nand NAND2_27193 ( P2_R2278_U452 , P2_U2797 , P2_R2278_U36 );
nand NAND2_27194 ( P2_R2278_U453 , P2_INSTADDRPOINTER_REG_24_ , P2_R2278_U35 );
nand NAND2_27195 ( P2_R2278_U454 , P2_U2797 , P2_R2278_U36 );
nand NAND2_27196 ( P2_R2278_U455 , P2_R2278_U454 , P2_R2278_U453 );
nand NAND2_27197 ( P2_R2278_U456 , P2_R2278_U175 , P2_R2278_U176 );
nand NAND2_27198 ( P2_R2278_U457 , P2_R2278_U286 , P2_R2278_U455 );
nand NAND2_27199 ( P2_R2278_U458 , P2_INSTADDRPOINTER_REG_23_ , P2_R2278_U69 );
nand NAND2_27200 ( P2_R2278_U459 , P2_U2798 , P2_R2278_U70 );
nand NAND2_27201 ( P2_R2278_U460 , P2_INSTADDRPOINTER_REG_23_ , P2_R2278_U69 );
nand NAND2_27202 ( P2_R2278_U461 , P2_U2798 , P2_R2278_U70 );
nand NAND2_27203 ( P2_R2278_U462 , P2_R2278_U461 , P2_R2278_U460 );
nand NAND2_27204 ( P2_R2278_U463 , P2_R2278_U177 , P2_R2278_U178 );
nand NAND2_27205 ( P2_R2278_U464 , P2_R2278_U282 , P2_R2278_U462 );
nand NAND2_27206 ( P2_R2278_U465 , P2_INSTADDRPOINTER_REG_22_ , P2_R2278_U37 );
nand NAND2_27207 ( P2_R2278_U466 , P2_U2799 , P2_R2278_U38 );
nand NAND2_27208 ( P2_R2278_U467 , P2_INSTADDRPOINTER_REG_22_ , P2_R2278_U37 );
nand NAND2_27209 ( P2_R2278_U468 , P2_U2799 , P2_R2278_U38 );
nand NAND2_27210 ( P2_R2278_U469 , P2_R2278_U468 , P2_R2278_U467 );
nand NAND2_27211 ( P2_R2278_U470 , P2_R2278_U179 , P2_R2278_U180 );
nand NAND2_27212 ( P2_R2278_U471 , P2_R2278_U279 , P2_R2278_U469 );
nand NAND2_27213 ( P2_R2278_U472 , P2_INSTADDRPOINTER_REG_21_ , P2_R2278_U66 );
nand NAND2_27214 ( P2_R2278_U473 , P2_U2800 , P2_R2278_U67 );
nand NAND2_27215 ( P2_R2278_U474 , P2_INSTADDRPOINTER_REG_21_ , P2_R2278_U66 );
nand NAND2_27216 ( P2_R2278_U475 , P2_U2800 , P2_R2278_U67 );
nand NAND2_27217 ( P2_R2278_U476 , P2_R2278_U475 , P2_R2278_U474 );
nand NAND2_27218 ( P2_R2278_U477 , P2_R2278_U181 , P2_R2278_U182 );
nand NAND2_27219 ( P2_R2278_U478 , P2_R2278_U275 , P2_R2278_U476 );
nand NAND2_27220 ( P2_R2278_U479 , P2_INSTADDRPOINTER_REG_20_ , P2_R2278_U39 );
nand NAND2_27221 ( P2_R2278_U480 , P2_U2801 , P2_R2278_U40 );
nand NAND2_27222 ( P2_R2278_U481 , P2_INSTADDRPOINTER_REG_20_ , P2_R2278_U39 );
nand NAND2_27223 ( P2_R2278_U482 , P2_U2801 , P2_R2278_U40 );
nand NAND2_27224 ( P2_R2278_U483 , P2_R2278_U482 , P2_R2278_U481 );
nand NAND2_27225 ( P2_R2278_U484 , P2_R2278_U183 , P2_R2278_U184 );
nand NAND2_27226 ( P2_R2278_U485 , P2_R2278_U272 , P2_R2278_U483 );
nand NAND2_27227 ( P2_R2278_U486 , P2_INSTADDRPOINTER_REG_1_ , P2_R2278_U15 );
nand NAND2_27228 ( P2_R2278_U487 , P2_R2278_U208 , P2_R2278_U17 );
nand NAND2_27229 ( P2_R2278_U488 , P2_R2278_U487 , P2_R2278_U486 );
nand NAND3_27230 ( P2_R2278_U489 , P2_R2278_U15 , P2_R2278_U17 , P2_U3637 );
nand NAND2_27231 ( P2_R2278_U490 , P2_R2278_U488 , P2_R2278_U16 );
nand NAND2_27232 ( P2_R2278_U491 , P2_INSTADDRPOINTER_REG_19_ , P2_R2278_U62 );
nand NAND2_27233 ( P2_R2278_U492 , P2_U2802 , P2_R2278_U63 );
nand NAND2_27234 ( P2_R2278_U493 , P2_INSTADDRPOINTER_REG_19_ , P2_R2278_U62 );
nand NAND2_27235 ( P2_R2278_U494 , P2_U2802 , P2_R2278_U63 );
nand NAND2_27236 ( P2_R2278_U495 , P2_R2278_U494 , P2_R2278_U493 );
nand NAND2_27237 ( P2_R2278_U496 , P2_R2278_U185 , P2_R2278_U186 );
nand NAND2_27238 ( P2_R2278_U497 , P2_R2278_U269 , P2_R2278_U495 );
nand NAND2_27239 ( P2_R2278_U498 , P2_INSTADDRPOINTER_REG_18_ , P2_R2278_U64 );
nand NAND2_27240 ( P2_R2278_U499 , P2_U2803 , P2_R2278_U65 );
nand NAND2_27241 ( P2_R2278_U500 , P2_INSTADDRPOINTER_REG_18_ , P2_R2278_U64 );
nand NAND2_27242 ( P2_R2278_U501 , P2_U2803 , P2_R2278_U65 );
nand NAND2_27243 ( P2_R2278_U502 , P2_R2278_U501 , P2_R2278_U500 );
nand NAND2_27244 ( P2_R2278_U503 , P2_R2278_U187 , P2_R2278_U188 );
nand NAND2_27245 ( P2_R2278_U504 , P2_R2278_U265 , P2_R2278_U502 );
nand NAND2_27246 ( P2_R2278_U505 , P2_INSTADDRPOINTER_REG_17_ , P2_R2278_U41 );
nand NAND2_27247 ( P2_R2278_U506 , P2_U2804 , P2_R2278_U42 );
nand NAND2_27248 ( P2_R2278_U507 , P2_INSTADDRPOINTER_REG_17_ , P2_R2278_U41 );
nand NAND2_27249 ( P2_R2278_U508 , P2_U2804 , P2_R2278_U42 );
nand NAND2_27250 ( P2_R2278_U509 , P2_R2278_U508 , P2_R2278_U507 );
nand NAND2_27251 ( P2_R2278_U510 , P2_R2278_U189 , P2_R2278_U190 );
nand NAND2_27252 ( P2_R2278_U511 , P2_R2278_U262 , P2_R2278_U509 );
nand NAND2_27253 ( P2_R2278_U512 , P2_INSTADDRPOINTER_REG_16_ , P2_R2278_U59 );
nand NAND2_27254 ( P2_R2278_U513 , P2_U2805 , P2_R2278_U60 );
nand NAND2_27255 ( P2_R2278_U514 , P2_INSTADDRPOINTER_REG_16_ , P2_R2278_U59 );
nand NAND2_27256 ( P2_R2278_U515 , P2_U2805 , P2_R2278_U60 );
nand NAND2_27257 ( P2_R2278_U516 , P2_R2278_U515 , P2_R2278_U514 );
nand NAND2_27258 ( P2_R2278_U517 , P2_R2278_U191 , P2_R2278_U192 );
nand NAND2_27259 ( P2_R2278_U518 , P2_R2278_U258 , P2_R2278_U516 );
nand NAND2_27260 ( P2_R2278_U519 , P2_INSTADDRPOINTER_REG_15_ , P2_R2278_U43 );
nand NAND2_27261 ( P2_R2278_U520 , P2_U2806 , P2_R2278_U44 );
nand NAND2_27262 ( P2_R2278_U521 , P2_INSTADDRPOINTER_REG_15_ , P2_R2278_U43 );
nand NAND2_27263 ( P2_R2278_U522 , P2_U2806 , P2_R2278_U44 );
nand NAND2_27264 ( P2_R2278_U523 , P2_R2278_U522 , P2_R2278_U521 );
nand NAND2_27265 ( P2_R2278_U524 , P2_R2278_U193 , P2_R2278_U194 );
nand NAND2_27266 ( P2_R2278_U525 , P2_R2278_U255 , P2_R2278_U523 );
nand NAND2_27267 ( P2_R2278_U526 , P2_INSTADDRPOINTER_REG_14_ , P2_R2278_U56 );
nand NAND2_27268 ( P2_R2278_U527 , P2_U2807 , P2_R2278_U57 );
nand NAND2_27269 ( P2_R2278_U528 , P2_INSTADDRPOINTER_REG_14_ , P2_R2278_U56 );
nand NAND2_27270 ( P2_R2278_U529 , P2_U2807 , P2_R2278_U57 );
nand NAND2_27271 ( P2_R2278_U530 , P2_R2278_U529 , P2_R2278_U528 );
nand NAND2_27272 ( P2_R2278_U531 , P2_R2278_U195 , P2_R2278_U196 );
nand NAND2_27273 ( P2_R2278_U532 , P2_R2278_U251 , P2_R2278_U530 );
nand NAND2_27274 ( P2_R2278_U533 , P2_INSTADDRPOINTER_REG_13_ , P2_R2278_U45 );
nand NAND2_27275 ( P2_R2278_U534 , P2_U2808 , P2_R2278_U46 );
nand NAND2_27276 ( P2_R2278_U535 , P2_INSTADDRPOINTER_REG_13_ , P2_R2278_U45 );
nand NAND2_27277 ( P2_R2278_U536 , P2_U2808 , P2_R2278_U46 );
nand NAND2_27278 ( P2_R2278_U537 , P2_R2278_U536 , P2_R2278_U535 );
nand NAND2_27279 ( P2_R2278_U538 , P2_R2278_U197 , P2_R2278_U198 );
nand NAND2_27280 ( P2_R2278_U539 , P2_R2278_U248 , P2_R2278_U537 );
nand NAND2_27281 ( P2_R2278_U540 , P2_INSTADDRPOINTER_REG_12_ , P2_R2278_U53 );
nand NAND2_27282 ( P2_R2278_U541 , P2_U2809 , P2_R2278_U54 );
nand NAND2_27283 ( P2_R2278_U542 , P2_INSTADDRPOINTER_REG_12_ , P2_R2278_U53 );
nand NAND2_27284 ( P2_R2278_U543 , P2_U2809 , P2_R2278_U54 );
nand NAND2_27285 ( P2_R2278_U544 , P2_R2278_U543 , P2_R2278_U542 );
nand NAND2_27286 ( P2_R2278_U545 , P2_R2278_U199 , P2_R2278_U200 );
nand NAND2_27287 ( P2_R2278_U546 , P2_R2278_U244 , P2_R2278_U544 );
nand NAND2_27288 ( P2_R2278_U547 , P2_INSTADDRPOINTER_REG_11_ , P2_R2278_U47 );
nand NAND2_27289 ( P2_R2278_U548 , P2_U2810 , P2_R2278_U48 );
nand NAND2_27290 ( P2_R2278_U549 , P2_INSTADDRPOINTER_REG_11_ , P2_R2278_U47 );
nand NAND2_27291 ( P2_R2278_U550 , P2_U2810 , P2_R2278_U48 );
nand NAND2_27292 ( P2_R2278_U551 , P2_R2278_U550 , P2_R2278_U549 );
nand NAND2_27293 ( P2_R2278_U552 , P2_R2278_U201 , P2_R2278_U202 );
nand NAND2_27294 ( P2_R2278_U553 , P2_R2278_U241 , P2_R2278_U551 );
nand NAND2_27295 ( P2_R2278_U554 , P2_INSTADDRPOINTER_REG_10_ , P2_R2278_U50 );
nand NAND2_27296 ( P2_R2278_U555 , P2_U2811 , P2_R2278_U51 );
nand NAND2_27297 ( P2_R2278_U556 , P2_INSTADDRPOINTER_REG_10_ , P2_R2278_U50 );
nand NAND2_27298 ( P2_R2278_U557 , P2_U2811 , P2_R2278_U51 );
nand NAND2_27299 ( P2_R2278_U558 , P2_R2278_U557 , P2_R2278_U556 );
nand NAND2_27300 ( P2_R2278_U559 , P2_R2278_U203 , P2_R2278_U204 );
nand NAND2_27301 ( P2_R2278_U560 , P2_R2278_U237 , P2_R2278_U558 );
nand NAND2_27302 ( P2_R2278_U561 , P2_INSTADDRPOINTER_REG_0_ , P2_R2278_U13 );
nand NAND2_27303 ( P2_R2278_U562 , P2_U3638 , P2_R2278_U14 );
nand NAND2_27304 ( P2_SUB_450_U6 , P2_SUB_450_U43 , P2_SUB_450_U42 );
nand NAND2_27305 ( P2_SUB_450_U7 , P2_INSTQUEUERD_ADDR_REG_0_ , P2_SUB_450_U16 );
not NOT1_27306 ( P2_SUB_450_U8 , P2_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_27307 ( P2_SUB_450_U9 , P2_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_27308 ( P2_SUB_450_U10 , P2_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_27309 ( P2_SUB_450_U11 , P2_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_27310 ( P2_SUB_450_U12 , P2_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_27311 ( P2_SUB_450_U13 , P2_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_27312 ( P2_SUB_450_U14 , P2_SUB_450_U39 , P2_SUB_450_U38 );
not NOT1_27313 ( P2_SUB_450_U15 , P2_INSTQUEUERD_ADDR_REG_4_ );
not NOT1_27314 ( P2_SUB_450_U16 , P2_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_27315 ( P2_SUB_450_U17 , P2_SUB_450_U48 , P2_SUB_450_U47 );
nand NAND2_27316 ( P2_SUB_450_U18 , P2_SUB_450_U53 , P2_SUB_450_U52 );
nand NAND2_27317 ( P2_SUB_450_U19 , P2_SUB_450_U58 , P2_SUB_450_U57 );
nand NAND2_27318 ( P2_SUB_450_U20 , P2_SUB_450_U63 , P2_SUB_450_U62 );
nand NAND2_27319 ( P2_SUB_450_U21 , P2_SUB_450_U45 , P2_SUB_450_U44 );
nand NAND2_27320 ( P2_SUB_450_U22 , P2_SUB_450_U50 , P2_SUB_450_U49 );
nand NAND2_27321 ( P2_SUB_450_U23 , P2_SUB_450_U55 , P2_SUB_450_U54 );
nand NAND2_27322 ( P2_SUB_450_U24 , P2_SUB_450_U60 , P2_SUB_450_U59 );
nand NAND2_27323 ( P2_SUB_450_U25 , P2_SUB_450_U35 , P2_SUB_450_U34 );
nand NAND2_27324 ( P2_SUB_450_U26 , P2_SUB_450_U31 , P2_SUB_450_U30 );
not NOT1_27325 ( P2_SUB_450_U27 , P2_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_27326 ( P2_SUB_450_U28 , P2_SUB_450_U7 );
nand NAND2_27327 ( P2_SUB_450_U29 , P2_SUB_450_U28 , P2_SUB_450_U8 );
nand NAND2_27328 ( P2_SUB_450_U30 , P2_SUB_450_U29 , P2_SUB_450_U27 );
nand NAND2_27329 ( P2_SUB_450_U31 , P2_INSTQUEUEWR_ADDR_REG_1_ , P2_SUB_450_U7 );
not NOT1_27330 ( P2_SUB_450_U32 , P2_SUB_450_U26 );
nand NAND2_27331 ( P2_SUB_450_U33 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_SUB_450_U10 );
nand NAND2_27332 ( P2_SUB_450_U34 , P2_SUB_450_U33 , P2_SUB_450_U26 );
nand NAND2_27333 ( P2_SUB_450_U35 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_SUB_450_U9 );
not NOT1_27334 ( P2_SUB_450_U36 , P2_SUB_450_U25 );
nand NAND2_27335 ( P2_SUB_450_U37 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_SUB_450_U12 );
nand NAND2_27336 ( P2_SUB_450_U38 , P2_SUB_450_U37 , P2_SUB_450_U25 );
nand NAND2_27337 ( P2_SUB_450_U39 , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_SUB_450_U11 );
not NOT1_27338 ( P2_SUB_450_U40 , P2_SUB_450_U14 );
nand NAND2_27339 ( P2_SUB_450_U41 , P2_INSTQUEUEWR_ADDR_REG_4_ , P2_SUB_450_U15 );
nand NAND2_27340 ( P2_SUB_450_U42 , P2_SUB_450_U40 , P2_SUB_450_U41 );
nand NAND2_27341 ( P2_SUB_450_U43 , P2_INSTQUEUERD_ADDR_REG_4_ , P2_SUB_450_U13 );
nand NAND2_27342 ( P2_SUB_450_U44 , P2_INSTQUEUERD_ADDR_REG_4_ , P2_SUB_450_U13 );
nand NAND2_27343 ( P2_SUB_450_U45 , P2_INSTQUEUEWR_ADDR_REG_4_ , P2_SUB_450_U15 );
not NOT1_27344 ( P2_SUB_450_U46 , P2_SUB_450_U21 );
nand NAND2_27345 ( P2_SUB_450_U47 , P2_SUB_450_U46 , P2_SUB_450_U40 );
nand NAND2_27346 ( P2_SUB_450_U48 , P2_SUB_450_U21 , P2_SUB_450_U14 );
nand NAND2_27347 ( P2_SUB_450_U49 , P2_INSTQUEUERD_ADDR_REG_3_ , P2_SUB_450_U12 );
nand NAND2_27348 ( P2_SUB_450_U50 , P2_INSTQUEUEWR_ADDR_REG_3_ , P2_SUB_450_U11 );
not NOT1_27349 ( P2_SUB_450_U51 , P2_SUB_450_U22 );
nand NAND2_27350 ( P2_SUB_450_U52 , P2_SUB_450_U36 , P2_SUB_450_U51 );
nand NAND2_27351 ( P2_SUB_450_U53 , P2_SUB_450_U22 , P2_SUB_450_U25 );
nand NAND2_27352 ( P2_SUB_450_U54 , P2_INSTQUEUERD_ADDR_REG_2_ , P2_SUB_450_U10 );
nand NAND2_27353 ( P2_SUB_450_U55 , P2_INSTQUEUEWR_ADDR_REG_2_ , P2_SUB_450_U9 );
not NOT1_27354 ( P2_SUB_450_U56 , P2_SUB_450_U23 );
nand NAND2_27355 ( P2_SUB_450_U57 , P2_SUB_450_U32 , P2_SUB_450_U56 );
nand NAND2_27356 ( P2_SUB_450_U58 , P2_SUB_450_U23 , P2_SUB_450_U26 );
nand NAND2_27357 ( P2_SUB_450_U59 , P2_INSTQUEUERD_ADDR_REG_1_ , P2_SUB_450_U8 );
nand NAND2_27358 ( P2_SUB_450_U60 , P2_INSTQUEUEWR_ADDR_REG_1_ , P2_SUB_450_U27 );
not NOT1_27359 ( P2_SUB_450_U61 , P2_SUB_450_U24 );
nand NAND2_27360 ( P2_SUB_450_U62 , P2_SUB_450_U61 , P2_SUB_450_U28 );
nand NAND2_27361 ( P2_SUB_450_U63 , P2_SUB_450_U24 , P2_SUB_450_U7 );
nor nor_27362 ( P2_R2088_U6 , P2_U3648 , P2_R2088_U7 );
nor nor_27363 ( P2_R2088_U7 , P2_U3648 , P2_U3649 , P2_U3650 , P2_U3652 , P2_U3651 );
not NOT1_27364 ( P2_ADD_394_U4 , P2_INSTADDRPOINTER_REG_0_ );
nand NAND2_27365 ( P2_ADD_394_U5 , P2_ADD_394_U94 , P2_ADD_394_U125 );
not NOT1_27366 ( P2_ADD_394_U6 , P2_INSTADDRPOINTER_REG_1_ );
not NOT1_27367 ( P2_ADD_394_U7 , P2_INSTADDRPOINTER_REG_3_ );
nand NAND2_27368 ( P2_ADD_394_U8 , P2_INSTADDRPOINTER_REG_3_ , P2_ADD_394_U94 );
not NOT1_27369 ( P2_ADD_394_U9 , P2_INSTADDRPOINTER_REG_4_ );
nand NAND2_27370 ( P2_ADD_394_U10 , P2_INSTADDRPOINTER_REG_4_ , P2_ADD_394_U98 );
not NOT1_27371 ( P2_ADD_394_U11 , P2_INSTADDRPOINTER_REG_5_ );
not NOT1_27372 ( P2_ADD_394_U12 , P2_INSTADDRPOINTER_REG_6_ );
nand NAND2_27373 ( P2_ADD_394_U13 , P2_INSTADDRPOINTER_REG_5_ , P2_ADD_394_U99 );
nand NAND2_27374 ( P2_ADD_394_U14 , P2_ADD_394_U100 , P2_INSTADDRPOINTER_REG_6_ );
not NOT1_27375 ( P2_ADD_394_U15 , P2_INSTADDRPOINTER_REG_7_ );
nand NAND2_27376 ( P2_ADD_394_U16 , P2_INSTADDRPOINTER_REG_7_ , P2_ADD_394_U101 );
not NOT1_27377 ( P2_ADD_394_U17 , P2_INSTADDRPOINTER_REG_8_ );
nand NAND2_27378 ( P2_ADD_394_U18 , P2_INSTADDRPOINTER_REG_8_ , P2_ADD_394_U102 );
not NOT1_27379 ( P2_ADD_394_U19 , P2_INSTADDRPOINTER_REG_9_ );
nand NAND2_27380 ( P2_ADD_394_U20 , P2_INSTADDRPOINTER_REG_9_ , P2_ADD_394_U103 );
not NOT1_27381 ( P2_ADD_394_U21 , P2_INSTADDRPOINTER_REG_10_ );
nand NAND2_27382 ( P2_ADD_394_U22 , P2_INSTADDRPOINTER_REG_10_ , P2_ADD_394_U104 );
not NOT1_27383 ( P2_ADD_394_U23 , P2_INSTADDRPOINTER_REG_11_ );
nand NAND2_27384 ( P2_ADD_394_U24 , P2_INSTADDRPOINTER_REG_11_ , P2_ADD_394_U105 );
not NOT1_27385 ( P2_ADD_394_U25 , P2_INSTADDRPOINTER_REG_12_ );
nand NAND2_27386 ( P2_ADD_394_U26 , P2_INSTADDRPOINTER_REG_12_ , P2_ADD_394_U106 );
not NOT1_27387 ( P2_ADD_394_U27 , P2_INSTADDRPOINTER_REG_13_ );
nand NAND2_27388 ( P2_ADD_394_U28 , P2_INSTADDRPOINTER_REG_13_ , P2_ADD_394_U107 );
not NOT1_27389 ( P2_ADD_394_U29 , P2_INSTADDRPOINTER_REG_14_ );
nand NAND2_27390 ( P2_ADD_394_U30 , P2_INSTADDRPOINTER_REG_14_ , P2_ADD_394_U108 );
not NOT1_27391 ( P2_ADD_394_U31 , P2_INSTADDRPOINTER_REG_15_ );
nand NAND2_27392 ( P2_ADD_394_U32 , P2_INSTADDRPOINTER_REG_15_ , P2_ADD_394_U109 );
not NOT1_27393 ( P2_ADD_394_U33 , P2_INSTADDRPOINTER_REG_16_ );
nand NAND2_27394 ( P2_ADD_394_U34 , P2_INSTADDRPOINTER_REG_16_ , P2_ADD_394_U110 );
not NOT1_27395 ( P2_ADD_394_U35 , P2_INSTADDRPOINTER_REG_17_ );
nand NAND2_27396 ( P2_ADD_394_U36 , P2_INSTADDRPOINTER_REG_17_ , P2_ADD_394_U111 );
not NOT1_27397 ( P2_ADD_394_U37 , P2_INSTADDRPOINTER_REG_18_ );
nand NAND2_27398 ( P2_ADD_394_U38 , P2_INSTADDRPOINTER_REG_18_ , P2_ADD_394_U112 );
not NOT1_27399 ( P2_ADD_394_U39 , P2_INSTADDRPOINTER_REG_19_ );
nand NAND2_27400 ( P2_ADD_394_U40 , P2_INSTADDRPOINTER_REG_19_ , P2_ADD_394_U113 );
not NOT1_27401 ( P2_ADD_394_U41 , P2_INSTADDRPOINTER_REG_20_ );
nand NAND2_27402 ( P2_ADD_394_U42 , P2_INSTADDRPOINTER_REG_20_ , P2_ADD_394_U114 );
not NOT1_27403 ( P2_ADD_394_U43 , P2_INSTADDRPOINTER_REG_21_ );
nand NAND2_27404 ( P2_ADD_394_U44 , P2_INSTADDRPOINTER_REG_21_ , P2_ADD_394_U115 );
not NOT1_27405 ( P2_ADD_394_U45 , P2_INSTADDRPOINTER_REG_22_ );
nand NAND2_27406 ( P2_ADD_394_U46 , P2_INSTADDRPOINTER_REG_22_ , P2_ADD_394_U116 );
not NOT1_27407 ( P2_ADD_394_U47 , P2_INSTADDRPOINTER_REG_23_ );
nand NAND2_27408 ( P2_ADD_394_U48 , P2_INSTADDRPOINTER_REG_23_ , P2_ADD_394_U117 );
not NOT1_27409 ( P2_ADD_394_U49 , P2_INSTADDRPOINTER_REG_24_ );
nand NAND2_27410 ( P2_ADD_394_U50 , P2_INSTADDRPOINTER_REG_24_ , P2_ADD_394_U118 );
not NOT1_27411 ( P2_ADD_394_U51 , P2_INSTADDRPOINTER_REG_25_ );
nand NAND2_27412 ( P2_ADD_394_U52 , P2_INSTADDRPOINTER_REG_25_ , P2_ADD_394_U119 );
not NOT1_27413 ( P2_ADD_394_U53 , P2_INSTADDRPOINTER_REG_26_ );
nand NAND2_27414 ( P2_ADD_394_U54 , P2_INSTADDRPOINTER_REG_26_ , P2_ADD_394_U120 );
not NOT1_27415 ( P2_ADD_394_U55 , P2_INSTADDRPOINTER_REG_27_ );
nand NAND2_27416 ( P2_ADD_394_U56 , P2_INSTADDRPOINTER_REG_27_ , P2_ADD_394_U121 );
not NOT1_27417 ( P2_ADD_394_U57 , P2_INSTADDRPOINTER_REG_28_ );
nand NAND2_27418 ( P2_ADD_394_U58 , P2_INSTADDRPOINTER_REG_28_ , P2_ADD_394_U122 );
not NOT1_27419 ( P2_ADD_394_U59 , P2_INSTADDRPOINTER_REG_29_ );
not NOT1_27420 ( P2_ADD_394_U60 , P2_INSTADDRPOINTER_REG_30_ );
nand NAND2_27421 ( P2_ADD_394_U61 , P2_INSTADDRPOINTER_REG_29_ , P2_ADD_394_U123 );
not NOT1_27422 ( P2_ADD_394_U62 , P2_INSTADDRPOINTER_REG_2_ );
nand NAND2_27423 ( P2_ADD_394_U63 , P2_ADD_394_U128 , P2_ADD_394_U127 );
nand NAND2_27424 ( P2_ADD_394_U64 , P2_ADD_394_U130 , P2_ADD_394_U129 );
nand NAND2_27425 ( P2_ADD_394_U65 , P2_ADD_394_U132 , P2_ADD_394_U131 );
nand NAND2_27426 ( P2_ADD_394_U66 , P2_ADD_394_U134 , P2_ADD_394_U133 );
nand NAND2_27427 ( P2_ADD_394_U67 , P2_ADD_394_U136 , P2_ADD_394_U135 );
nand NAND2_27428 ( P2_ADD_394_U68 , P2_ADD_394_U138 , P2_ADD_394_U137 );
nand NAND2_27429 ( P2_ADD_394_U69 , P2_ADD_394_U140 , P2_ADD_394_U139 );
nand NAND2_27430 ( P2_ADD_394_U70 , P2_ADD_394_U142 , P2_ADD_394_U141 );
nand NAND2_27431 ( P2_ADD_394_U71 , P2_ADD_394_U144 , P2_ADD_394_U143 );
nand NAND2_27432 ( P2_ADD_394_U72 , P2_ADD_394_U146 , P2_ADD_394_U145 );
nand NAND2_27433 ( P2_ADD_394_U73 , P2_ADD_394_U148 , P2_ADD_394_U147 );
nand NAND2_27434 ( P2_ADD_394_U74 , P2_ADD_394_U150 , P2_ADD_394_U149 );
nand NAND2_27435 ( P2_ADD_394_U75 , P2_ADD_394_U152 , P2_ADD_394_U151 );
nand NAND2_27436 ( P2_ADD_394_U76 , P2_ADD_394_U154 , P2_ADD_394_U153 );
nand NAND2_27437 ( P2_ADD_394_U77 , P2_ADD_394_U156 , P2_ADD_394_U155 );
nand NAND2_27438 ( P2_ADD_394_U78 , P2_ADD_394_U158 , P2_ADD_394_U157 );
nand NAND2_27439 ( P2_ADD_394_U79 , P2_ADD_394_U160 , P2_ADD_394_U159 );
nand NAND2_27440 ( P2_ADD_394_U80 , P2_ADD_394_U162 , P2_ADD_394_U161 );
nand NAND2_27441 ( P2_ADD_394_U81 , P2_ADD_394_U164 , P2_ADD_394_U163 );
nand NAND2_27442 ( P2_ADD_394_U82 , P2_ADD_394_U166 , P2_ADD_394_U165 );
nand NAND2_27443 ( P2_ADD_394_U83 , P2_ADD_394_U168 , P2_ADD_394_U167 );
nand NAND2_27444 ( P2_ADD_394_U84 , P2_ADD_394_U170 , P2_ADD_394_U169 );
nand NAND2_27445 ( P2_ADD_394_U85 , P2_ADD_394_U174 , P2_ADD_394_U173 );
nand NAND2_27446 ( P2_ADD_394_U86 , P2_ADD_394_U176 , P2_ADD_394_U175 );
nand NAND2_27447 ( P2_ADD_394_U87 , P2_ADD_394_U178 , P2_ADD_394_U177 );
nand NAND2_27448 ( P2_ADD_394_U88 , P2_ADD_394_U180 , P2_ADD_394_U179 );
nand NAND2_27449 ( P2_ADD_394_U89 , P2_ADD_394_U182 , P2_ADD_394_U181 );
nand NAND2_27450 ( P2_ADD_394_U90 , P2_ADD_394_U184 , P2_ADD_394_U183 );
nand NAND2_27451 ( P2_ADD_394_U91 , P2_ADD_394_U186 , P2_ADD_394_U185 );
not NOT1_27452 ( P2_ADD_394_U92 , P2_INSTADDRPOINTER_REG_31_ );
nand NAND2_27453 ( P2_ADD_394_U93 , P2_ADD_394_U124 , P2_INSTADDRPOINTER_REG_30_ );
nand NAND2_27454 ( P2_ADD_394_U94 , P2_ADD_394_U62 , P2_ADD_394_U96 );
and AND2_27455 ( P2_ADD_394_U95 , P2_ADD_394_U172 , P2_ADD_394_U171 );
nand NAND2_27456 ( P2_ADD_394_U96 , P2_INSTADDRPOINTER_REG_1_ , P2_INSTADDRPOINTER_REG_0_ );
not NOT1_27457 ( P2_ADD_394_U97 , P2_ADD_394_U94 );
not NOT1_27458 ( P2_ADD_394_U98 , P2_ADD_394_U8 );
not NOT1_27459 ( P2_ADD_394_U99 , P2_ADD_394_U10 );
not NOT1_27460 ( P2_ADD_394_U100 , P2_ADD_394_U13 );
not NOT1_27461 ( P2_ADD_394_U101 , P2_ADD_394_U14 );
not NOT1_27462 ( P2_ADD_394_U102 , P2_ADD_394_U16 );
not NOT1_27463 ( P2_ADD_394_U103 , P2_ADD_394_U18 );
not NOT1_27464 ( P2_ADD_394_U104 , P2_ADD_394_U20 );
not NOT1_27465 ( P2_ADD_394_U105 , P2_ADD_394_U22 );
not NOT1_27466 ( P2_ADD_394_U106 , P2_ADD_394_U24 );
not NOT1_27467 ( P2_ADD_394_U107 , P2_ADD_394_U26 );
not NOT1_27468 ( P2_ADD_394_U108 , P2_ADD_394_U28 );
not NOT1_27469 ( P2_ADD_394_U109 , P2_ADD_394_U30 );
not NOT1_27470 ( P2_ADD_394_U110 , P2_ADD_394_U32 );
not NOT1_27471 ( P2_ADD_394_U111 , P2_ADD_394_U34 );
not NOT1_27472 ( P2_ADD_394_U112 , P2_ADD_394_U36 );
not NOT1_27473 ( P2_ADD_394_U113 , P2_ADD_394_U38 );
not NOT1_27474 ( P2_ADD_394_U114 , P2_ADD_394_U40 );
not NOT1_27475 ( P2_ADD_394_U115 , P2_ADD_394_U42 );
not NOT1_27476 ( P2_ADD_394_U116 , P2_ADD_394_U44 );
not NOT1_27477 ( P2_ADD_394_U117 , P2_ADD_394_U46 );
not NOT1_27478 ( P2_ADD_394_U118 , P2_ADD_394_U48 );
not NOT1_27479 ( P2_ADD_394_U119 , P2_ADD_394_U50 );
not NOT1_27480 ( P2_ADD_394_U120 , P2_ADD_394_U52 );
not NOT1_27481 ( P2_ADD_394_U121 , P2_ADD_394_U54 );
not NOT1_27482 ( P2_ADD_394_U122 , P2_ADD_394_U56 );
not NOT1_27483 ( P2_ADD_394_U123 , P2_ADD_394_U58 );
not NOT1_27484 ( P2_ADD_394_U124 , P2_ADD_394_U61 );
nand NAND3_27485 ( P2_ADD_394_U125 , P2_INSTADDRPOINTER_REG_1_ , P2_INSTADDRPOINTER_REG_0_ , P2_INSTADDRPOINTER_REG_2_ );
not NOT1_27486 ( P2_ADD_394_U126 , P2_ADD_394_U93 );
nand NAND2_27487 ( P2_ADD_394_U127 , P2_INSTADDRPOINTER_REG_6_ , P2_ADD_394_U13 );
nand NAND2_27488 ( P2_ADD_394_U128 , P2_ADD_394_U100 , P2_ADD_394_U12 );
nand NAND2_27489 ( P2_ADD_394_U129 , P2_INSTADDRPOINTER_REG_30_ , P2_ADD_394_U61 );
nand NAND2_27490 ( P2_ADD_394_U130 , P2_ADD_394_U124 , P2_ADD_394_U60 );
nand NAND2_27491 ( P2_ADD_394_U131 , P2_INSTADDRPOINTER_REG_29_ , P2_ADD_394_U58 );
nand NAND2_27492 ( P2_ADD_394_U132 , P2_ADD_394_U123 , P2_ADD_394_U59 );
nand NAND2_27493 ( P2_ADD_394_U133 , P2_INSTADDRPOINTER_REG_24_ , P2_ADD_394_U48 );
nand NAND2_27494 ( P2_ADD_394_U134 , P2_ADD_394_U118 , P2_ADD_394_U49 );
nand NAND2_27495 ( P2_ADD_394_U135 , P2_INSTADDRPOINTER_REG_17_ , P2_ADD_394_U34 );
nand NAND2_27496 ( P2_ADD_394_U136 , P2_ADD_394_U111 , P2_ADD_394_U35 );
nand NAND2_27497 ( P2_ADD_394_U137 , P2_INSTADDRPOINTER_REG_20_ , P2_ADD_394_U40 );
nand NAND2_27498 ( P2_ADD_394_U138 , P2_ADD_394_U114 , P2_ADD_394_U41 );
nand NAND2_27499 ( P2_ADD_394_U139 , P2_INSTADDRPOINTER_REG_13_ , P2_ADD_394_U26 );
nand NAND2_27500 ( P2_ADD_394_U140 , P2_ADD_394_U107 , P2_ADD_394_U27 );
nand NAND2_27501 ( P2_ADD_394_U141 , P2_INSTADDRPOINTER_REG_9_ , P2_ADD_394_U18 );
nand NAND2_27502 ( P2_ADD_394_U142 , P2_ADD_394_U103 , P2_ADD_394_U19 );
nand NAND2_27503 ( P2_ADD_394_U143 , P2_INSTADDRPOINTER_REG_22_ , P2_ADD_394_U44 );
nand NAND2_27504 ( P2_ADD_394_U144 , P2_ADD_394_U116 , P2_ADD_394_U45 );
nand NAND2_27505 ( P2_ADD_394_U145 , P2_INSTADDRPOINTER_REG_18_ , P2_ADD_394_U36 );
nand NAND2_27506 ( P2_ADD_394_U146 , P2_ADD_394_U112 , P2_ADD_394_U37 );
nand NAND2_27507 ( P2_ADD_394_U147 , P2_INSTADDRPOINTER_REG_11_ , P2_ADD_394_U22 );
nand NAND2_27508 ( P2_ADD_394_U148 , P2_ADD_394_U105 , P2_ADD_394_U23 );
nand NAND2_27509 ( P2_ADD_394_U149 , P2_INSTADDRPOINTER_REG_26_ , P2_ADD_394_U52 );
nand NAND2_27510 ( P2_ADD_394_U150 , P2_ADD_394_U120 , P2_ADD_394_U53 );
nand NAND2_27511 ( P2_ADD_394_U151 , P2_INSTADDRPOINTER_REG_15_ , P2_ADD_394_U30 );
nand NAND2_27512 ( P2_ADD_394_U152 , P2_ADD_394_U109 , P2_ADD_394_U31 );
nand NAND2_27513 ( P2_ADD_394_U153 , P2_INSTADDRPOINTER_REG_4_ , P2_ADD_394_U8 );
nand NAND2_27514 ( P2_ADD_394_U154 , P2_ADD_394_U98 , P2_ADD_394_U9 );
nand NAND2_27515 ( P2_ADD_394_U155 , P2_INSTADDRPOINTER_REG_27_ , P2_ADD_394_U54 );
nand NAND2_27516 ( P2_ADD_394_U156 , P2_ADD_394_U121 , P2_ADD_394_U55 );
nand NAND2_27517 ( P2_ADD_394_U157 , P2_INSTADDRPOINTER_REG_14_ , P2_ADD_394_U28 );
nand NAND2_27518 ( P2_ADD_394_U158 , P2_ADD_394_U108 , P2_ADD_394_U29 );
nand NAND2_27519 ( P2_ADD_394_U159 , P2_INSTADDRPOINTER_REG_5_ , P2_ADD_394_U10 );
nand NAND2_27520 ( P2_ADD_394_U160 , P2_ADD_394_U99 , P2_ADD_394_U11 );
nand NAND2_27521 ( P2_ADD_394_U161 , P2_INSTADDRPOINTER_REG_8_ , P2_ADD_394_U16 );
nand NAND2_27522 ( P2_ADD_394_U162 , P2_ADD_394_U102 , P2_ADD_394_U17 );
nand NAND2_27523 ( P2_ADD_394_U163 , P2_INSTADDRPOINTER_REG_23_ , P2_ADD_394_U46 );
nand NAND2_27524 ( P2_ADD_394_U164 , P2_ADD_394_U117 , P2_ADD_394_U47 );
nand NAND2_27525 ( P2_ADD_394_U165 , P2_INSTADDRPOINTER_REG_19_ , P2_ADD_394_U38 );
nand NAND2_27526 ( P2_ADD_394_U166 , P2_ADD_394_U113 , P2_ADD_394_U39 );
nand NAND2_27527 ( P2_ADD_394_U167 , P2_INSTADDRPOINTER_REG_10_ , P2_ADD_394_U20 );
nand NAND2_27528 ( P2_ADD_394_U168 , P2_ADD_394_U104 , P2_ADD_394_U21 );
nand NAND2_27529 ( P2_ADD_394_U169 , P2_INSTADDRPOINTER_REG_31_ , P2_ADD_394_U93 );
nand NAND2_27530 ( P2_ADD_394_U170 , P2_ADD_394_U126 , P2_ADD_394_U92 );
nand NAND2_27531 ( P2_ADD_394_U171 , P2_INSTADDRPOINTER_REG_3_ , P2_ADD_394_U94 );
nand NAND2_27532 ( P2_ADD_394_U172 , P2_ADD_394_U97 , P2_ADD_394_U7 );
nand NAND2_27533 ( P2_ADD_394_U173 , P2_INSTADDRPOINTER_REG_1_ , P2_ADD_394_U4 );
nand NAND2_27534 ( P2_ADD_394_U174 , P2_INSTADDRPOINTER_REG_0_ , P2_ADD_394_U6 );
nand NAND2_27535 ( P2_ADD_394_U175 , P2_INSTADDRPOINTER_REG_28_ , P2_ADD_394_U56 );
nand NAND2_27536 ( P2_ADD_394_U176 , P2_ADD_394_U122 , P2_ADD_394_U57 );
nand NAND2_27537 ( P2_ADD_394_U177 , P2_INSTADDRPOINTER_REG_21_ , P2_ADD_394_U42 );
nand NAND2_27538 ( P2_ADD_394_U178 , P2_ADD_394_U115 , P2_ADD_394_U43 );
nand NAND2_27539 ( P2_ADD_394_U179 , P2_INSTADDRPOINTER_REG_12_ , P2_ADD_394_U24 );
nand NAND2_27540 ( P2_ADD_394_U180 , P2_ADD_394_U106 , P2_ADD_394_U25 );
nand NAND2_27541 ( P2_ADD_394_U181 , P2_INSTADDRPOINTER_REG_7_ , P2_ADD_394_U14 );
nand NAND2_27542 ( P2_ADD_394_U182 , P2_ADD_394_U101 , P2_ADD_394_U15 );
nand NAND2_27543 ( P2_ADD_394_U183 , P2_INSTADDRPOINTER_REG_25_ , P2_ADD_394_U50 );
nand NAND2_27544 ( P2_ADD_394_U184 , P2_ADD_394_U119 , P2_ADD_394_U51 );
nand NAND2_27545 ( P2_ADD_394_U185 , P2_INSTADDRPOINTER_REG_16_ , P2_ADD_394_U32 );
nand NAND2_27546 ( P2_ADD_394_U186 , P2_ADD_394_U110 , P2_ADD_394_U33 );
and AND2_27547 ( P2_R2267_U6 , P2_R2267_U133 , P2_R2267_U31 );
and AND2_27548 ( P2_R2267_U7 , P2_R2267_U131 , P2_R2267_U32 );
and AND2_27549 ( P2_R2267_U8 , P2_R2267_U129 , P2_R2267_U33 );
and AND2_27550 ( P2_R2267_U9 , P2_R2267_U127 , P2_R2267_U34 );
and AND2_27551 ( P2_R2267_U10 , P2_R2267_U125 , P2_R2267_U35 );
and AND2_27552 ( P2_R2267_U11 , P2_R2267_U123 , P2_R2267_U36 );
and AND2_27553 ( P2_R2267_U12 , P2_R2267_U121 , P2_R2267_U37 );
and AND2_27554 ( P2_R2267_U13 , P2_R2267_U119 , P2_R2267_U38 );
and AND2_27555 ( P2_R2267_U14 , P2_R2267_U117 , P2_R2267_U39 );
and AND2_27556 ( P2_R2267_U15 , P2_R2267_U115 , P2_R2267_U40 );
and AND2_27557 ( P2_R2267_U16 , P2_R2267_U113 , P2_R2267_U62 );
and AND2_27558 ( P2_R2267_U17 , P2_R2267_U101 , P2_R2267_U24 );
and AND2_27559 ( P2_R2267_U18 , P2_R2267_U99 , P2_R2267_U25 );
and AND2_27560 ( P2_R2267_U19 , P2_R2267_U97 , P2_R2267_U26 );
and AND2_27561 ( P2_R2267_U20 , P2_R2267_U95 , P2_R2267_U30 );
nand NAND2_27562 ( P2_R2267_U21 , P2_R2267_U77 , P2_R2267_U134 );
not NOT1_27563 ( P2_R2267_U22 , P2_U3646 );
nand NAND2_27564 ( P2_R2267_U23 , P2_R2267_U76 , P2_R2267_U77 );
nand NAND3_27565 ( P2_R2267_U24 , P2_R2267_U89 , P2_R2267_U64 , P2_R2267_U29 );
nand NAND3_27566 ( P2_R2267_U25 , P2_R2267_U90 , P2_R2267_U59 , P2_R2267_U28 );
nand NAND3_27567 ( P2_R2267_U26 , P2_R2267_U91 , P2_R2267_U57 , P2_R2267_U27 );
not NOT1_27568 ( P2_R2267_U27 , P2_U3639 );
not NOT1_27569 ( P2_R2267_U28 , P2_U3641 );
not NOT1_27570 ( P2_R2267_U29 , P2_U3643 );
nand NAND2_27571 ( P2_R2267_U30 , P2_R2267_U44 , P2_R2267_U92 );
nand NAND2_27572 ( P2_R2267_U31 , P2_R2267_U45 , P2_R2267_U93 );
nand NAND2_27573 ( P2_R2267_U32 , P2_R2267_U46 , P2_R2267_U102 );
nand NAND2_27574 ( P2_R2267_U33 , P2_R2267_U47 , P2_R2267_U103 );
nand NAND2_27575 ( P2_R2267_U34 , P2_R2267_U48 , P2_R2267_U104 );
nand NAND2_27576 ( P2_R2267_U35 , P2_R2267_U49 , P2_R2267_U105 );
nand NAND2_27577 ( P2_R2267_U36 , P2_R2267_U50 , P2_R2267_U106 );
nand NAND2_27578 ( P2_R2267_U37 , P2_R2267_U51 , P2_R2267_U107 );
nand NAND2_27579 ( P2_R2267_U38 , P2_R2267_U52 , P2_R2267_U108 );
nand NAND2_27580 ( P2_R2267_U39 , P2_R2267_U53 , P2_R2267_U109 );
nand NAND2_27581 ( P2_R2267_U40 , P2_R2267_U54 , P2_R2267_U110 );
not NOT1_27582 ( P2_R2267_U41 , P2_U2767 );
not NOT1_27583 ( P2_R2267_U42 , P2_U2617 );
nand NAND2_27584 ( P2_R2267_U43 , P2_R2267_U156 , P2_R2267_U155 );
nor nor_27585 ( P2_R2267_U44 , P2_U2789 , P2_U2788 );
nor nor_27586 ( P2_R2267_U45 , P2_U2787 , P2_U2786 );
nor nor_27587 ( P2_R2267_U46 , P2_U2785 , P2_U2784 );
nor nor_27588 ( P2_R2267_U47 , P2_U2783 , P2_U2782 );
nor nor_27589 ( P2_R2267_U48 , P2_U2781 , P2_U2780 );
nor nor_27590 ( P2_R2267_U49 , P2_U2779 , P2_U2778 );
nor nor_27591 ( P2_R2267_U50 , P2_U2777 , P2_U2776 );
nor nor_27592 ( P2_R2267_U51 , P2_U2775 , P2_U2774 );
nor nor_27593 ( P2_R2267_U52 , P2_U2773 , P2_U2772 );
nor nor_27594 ( P2_R2267_U53 , P2_U2771 , P2_U2770 );
nor nor_27595 ( P2_R2267_U54 , P2_U2769 , P2_U2768 );
not NOT1_27596 ( P2_R2267_U55 , P2_U2789 );
and AND2_27597 ( P2_R2267_U56 , P2_R2267_U136 , P2_R2267_U135 );
not NOT1_27598 ( P2_R2267_U57 , P2_U3640 );
and AND2_27599 ( P2_R2267_U58 , P2_R2267_U138 , P2_R2267_U137 );
not NOT1_27600 ( P2_R2267_U59 , P2_U3642 );
and AND2_27601 ( P2_R2267_U60 , P2_R2267_U140 , P2_R2267_U139 );
not NOT1_27602 ( P2_R2267_U61 , P2_U2766 );
nand NAND2_27603 ( P2_R2267_U62 , P2_R2267_U111 , P2_R2267_U41 );
and AND2_27604 ( P2_R2267_U63 , P2_R2267_U142 , P2_R2267_U141 );
not NOT1_27605 ( P2_R2267_U64 , P2_U3644 );
and AND2_27606 ( P2_R2267_U65 , P2_R2267_U144 , P2_R2267_U143 );
not NOT1_27607 ( P2_R2267_U66 , P2_U2769 );
and AND2_27608 ( P2_R2267_U67 , P2_R2267_U146 , P2_R2267_U145 );
not NOT1_27609 ( P2_R2267_U68 , P2_U2771 );
and AND2_27610 ( P2_R2267_U69 , P2_R2267_U148 , P2_R2267_U147 );
not NOT1_27611 ( P2_R2267_U70 , P2_U2773 );
and AND2_27612 ( P2_R2267_U71 , P2_R2267_U150 , P2_R2267_U149 );
not NOT1_27613 ( P2_R2267_U72 , P2_U2775 );
and AND2_27614 ( P2_R2267_U73 , P2_R2267_U152 , P2_R2267_U151 );
not NOT1_27615 ( P2_R2267_U74 , P2_U2777 );
and AND2_27616 ( P2_R2267_U75 , P2_R2267_U154 , P2_R2267_U153 );
not NOT1_27617 ( P2_R2267_U76 , P2_U3645 );
nand NAND2_27618 ( P2_R2267_U77 , P2_U3646 , P2_R2267_U42 );
not NOT1_27619 ( P2_R2267_U78 , P2_U2779 );
and AND2_27620 ( P2_R2267_U79 , P2_R2267_U158 , P2_R2267_U157 );
not NOT1_27621 ( P2_R2267_U80 , P2_U2781 );
and AND2_27622 ( P2_R2267_U81 , P2_R2267_U160 , P2_R2267_U159 );
not NOT1_27623 ( P2_R2267_U82 , P2_U2783 );
and AND2_27624 ( P2_R2267_U83 , P2_R2267_U162 , P2_R2267_U161 );
not NOT1_27625 ( P2_R2267_U84 , P2_U2785 );
and AND2_27626 ( P2_R2267_U85 , P2_R2267_U164 , P2_R2267_U163 );
not NOT1_27627 ( P2_R2267_U86 , P2_U2787 );
and AND2_27628 ( P2_R2267_U87 , P2_R2267_U166 , P2_R2267_U165 );
not NOT1_27629 ( P2_R2267_U88 , P2_R2267_U77 );
not NOT1_27630 ( P2_R2267_U89 , P2_R2267_U23 );
not NOT1_27631 ( P2_R2267_U90 , P2_R2267_U24 );
not NOT1_27632 ( P2_R2267_U91 , P2_R2267_U25 );
not NOT1_27633 ( P2_R2267_U92 , P2_R2267_U26 );
not NOT1_27634 ( P2_R2267_U93 , P2_R2267_U30 );
nand NAND2_27635 ( P2_R2267_U94 , P2_R2267_U92 , P2_R2267_U55 );
nand NAND2_27636 ( P2_R2267_U95 , P2_U2788 , P2_R2267_U94 );
nand NAND2_27637 ( P2_R2267_U96 , P2_R2267_U91 , P2_R2267_U57 );
nand NAND2_27638 ( P2_R2267_U97 , P2_U3639 , P2_R2267_U96 );
nand NAND2_27639 ( P2_R2267_U98 , P2_R2267_U90 , P2_R2267_U59 );
nand NAND2_27640 ( P2_R2267_U99 , P2_U3641 , P2_R2267_U98 );
nand NAND2_27641 ( P2_R2267_U100 , P2_R2267_U89 , P2_R2267_U64 );
nand NAND2_27642 ( P2_R2267_U101 , P2_U3643 , P2_R2267_U100 );
not NOT1_27643 ( P2_R2267_U102 , P2_R2267_U31 );
not NOT1_27644 ( P2_R2267_U103 , P2_R2267_U32 );
not NOT1_27645 ( P2_R2267_U104 , P2_R2267_U33 );
not NOT1_27646 ( P2_R2267_U105 , P2_R2267_U34 );
not NOT1_27647 ( P2_R2267_U106 , P2_R2267_U35 );
not NOT1_27648 ( P2_R2267_U107 , P2_R2267_U36 );
not NOT1_27649 ( P2_R2267_U108 , P2_R2267_U37 );
not NOT1_27650 ( P2_R2267_U109 , P2_R2267_U38 );
not NOT1_27651 ( P2_R2267_U110 , P2_R2267_U39 );
not NOT1_27652 ( P2_R2267_U111 , P2_R2267_U40 );
not NOT1_27653 ( P2_R2267_U112 , P2_R2267_U62 );
nand NAND2_27654 ( P2_R2267_U113 , P2_U2767 , P2_R2267_U40 );
nand NAND2_27655 ( P2_R2267_U114 , P2_R2267_U110 , P2_R2267_U66 );
nand NAND2_27656 ( P2_R2267_U115 , P2_U2768 , P2_R2267_U114 );
nand NAND2_27657 ( P2_R2267_U116 , P2_R2267_U109 , P2_R2267_U68 );
nand NAND2_27658 ( P2_R2267_U117 , P2_U2770 , P2_R2267_U116 );
nand NAND2_27659 ( P2_R2267_U118 , P2_R2267_U108 , P2_R2267_U70 );
nand NAND2_27660 ( P2_R2267_U119 , P2_U2772 , P2_R2267_U118 );
nand NAND2_27661 ( P2_R2267_U120 , P2_R2267_U107 , P2_R2267_U72 );
nand NAND2_27662 ( P2_R2267_U121 , P2_U2774 , P2_R2267_U120 );
nand NAND2_27663 ( P2_R2267_U122 , P2_R2267_U106 , P2_R2267_U74 );
nand NAND2_27664 ( P2_R2267_U123 , P2_U2776 , P2_R2267_U122 );
nand NAND2_27665 ( P2_R2267_U124 , P2_R2267_U105 , P2_R2267_U78 );
nand NAND2_27666 ( P2_R2267_U125 , P2_U2778 , P2_R2267_U124 );
nand NAND2_27667 ( P2_R2267_U126 , P2_R2267_U104 , P2_R2267_U80 );
nand NAND2_27668 ( P2_R2267_U127 , P2_U2780 , P2_R2267_U126 );
nand NAND2_27669 ( P2_R2267_U128 , P2_R2267_U103 , P2_R2267_U82 );
nand NAND2_27670 ( P2_R2267_U129 , P2_U2782 , P2_R2267_U128 );
nand NAND2_27671 ( P2_R2267_U130 , P2_R2267_U102 , P2_R2267_U84 );
nand NAND2_27672 ( P2_R2267_U131 , P2_U2784 , P2_R2267_U130 );
nand NAND2_27673 ( P2_R2267_U132 , P2_R2267_U93 , P2_R2267_U86 );
nand NAND2_27674 ( P2_R2267_U133 , P2_U2786 , P2_R2267_U132 );
nand NAND2_27675 ( P2_R2267_U134 , P2_U2617 , P2_R2267_U22 );
nand NAND2_27676 ( P2_R2267_U135 , P2_U2789 , P2_R2267_U26 );
nand NAND2_27677 ( P2_R2267_U136 , P2_R2267_U92 , P2_R2267_U55 );
nand NAND2_27678 ( P2_R2267_U137 , P2_U3640 , P2_R2267_U25 );
nand NAND2_27679 ( P2_R2267_U138 , P2_R2267_U91 , P2_R2267_U57 );
nand NAND2_27680 ( P2_R2267_U139 , P2_U3642 , P2_R2267_U24 );
nand NAND2_27681 ( P2_R2267_U140 , P2_R2267_U90 , P2_R2267_U59 );
nand NAND2_27682 ( P2_R2267_U141 , P2_U2766 , P2_R2267_U62 );
nand NAND2_27683 ( P2_R2267_U142 , P2_R2267_U112 , P2_R2267_U61 );
nand NAND2_27684 ( P2_R2267_U143 , P2_U3644 , P2_R2267_U23 );
nand NAND2_27685 ( P2_R2267_U144 , P2_R2267_U89 , P2_R2267_U64 );
nand NAND2_27686 ( P2_R2267_U145 , P2_U2769 , P2_R2267_U39 );
nand NAND2_27687 ( P2_R2267_U146 , P2_R2267_U110 , P2_R2267_U66 );
nand NAND2_27688 ( P2_R2267_U147 , P2_U2771 , P2_R2267_U38 );
nand NAND2_27689 ( P2_R2267_U148 , P2_R2267_U109 , P2_R2267_U68 );
nand NAND2_27690 ( P2_R2267_U149 , P2_U2773 , P2_R2267_U37 );
nand NAND2_27691 ( P2_R2267_U150 , P2_R2267_U108 , P2_R2267_U70 );
nand NAND2_27692 ( P2_R2267_U151 , P2_U2775 , P2_R2267_U36 );
nand NAND2_27693 ( P2_R2267_U152 , P2_R2267_U107 , P2_R2267_U72 );
nand NAND2_27694 ( P2_R2267_U153 , P2_U2777 , P2_R2267_U35 );
nand NAND2_27695 ( P2_R2267_U154 , P2_R2267_U106 , P2_R2267_U74 );
nand NAND2_27696 ( P2_R2267_U155 , P2_U3645 , P2_R2267_U77 );
nand NAND2_27697 ( P2_R2267_U156 , P2_R2267_U88 , P2_R2267_U76 );
nand NAND2_27698 ( P2_R2267_U157 , P2_U2779 , P2_R2267_U34 );
nand NAND2_27699 ( P2_R2267_U158 , P2_R2267_U105 , P2_R2267_U78 );
nand NAND2_27700 ( P2_R2267_U159 , P2_U2781 , P2_R2267_U33 );
nand NAND2_27701 ( P2_R2267_U160 , P2_R2267_U104 , P2_R2267_U80 );
nand NAND2_27702 ( P2_R2267_U161 , P2_U2783 , P2_R2267_U32 );
nand NAND2_27703 ( P2_R2267_U162 , P2_R2267_U103 , P2_R2267_U82 );
nand NAND2_27704 ( P2_R2267_U163 , P2_U2785 , P2_R2267_U31 );
nand NAND2_27705 ( P2_R2267_U164 , P2_R2267_U102 , P2_R2267_U84 );
nand NAND2_27706 ( P2_R2267_U165 , P2_U2787 , P2_R2267_U30 );
nand NAND2_27707 ( P2_R2267_U166 , P2_R2267_U93 , P2_R2267_U86 );
and AND2_27708 ( P2_ADD_371_1212_U4 , P2_INSTADDRPOINTER_REG_13_ , P2_ADD_371_1212_U10 );
and AND2_27709 ( P2_ADD_371_1212_U5 , P2_INSTADDRPOINTER_REG_10_ , P2_INSTADDRPOINTER_REG_9_ );
and AND2_27710 ( P2_ADD_371_1212_U6 , P2_ADD_371_1212_U89 , P2_ADD_371_1212_U11 );
and AND2_27711 ( P2_ADD_371_1212_U7 , P2_ADD_371_1212_U10 , P2_ADD_371_1212_U87 );
and AND2_27712 ( P2_ADD_371_1212_U8 , P2_ADD_371_1212_U9 , P2_ADD_371_1212_U91 );
and AND2_27713 ( P2_ADD_371_1212_U9 , P2_ADD_371_1212_U6 , P2_ADD_371_1212_U90 );
and AND4_27714 ( P2_ADD_371_1212_U10 , P2_INSTADDRPOINTER_REG_12_ , P2_INSTADDRPOINTER_REG_11_ , P2_INSTADDRPOINTER_REG_10_ , P2_INSTADDRPOINTER_REG_9_ );
and AND2_27715 ( P2_ADD_371_1212_U11 , P2_ADD_371_1212_U7 , P2_ADD_371_1212_U88 );
and AND2_27716 ( P2_ADD_371_1212_U12 , P2_ADD_371_1212_U8 , P2_ADD_371_1212_U92 );
and AND2_27717 ( P2_ADD_371_1212_U13 , P2_ADD_371_1212_U196 , P2_ADD_371_1212_U168 );
and AND2_27718 ( P2_ADD_371_1212_U14 , P2_ADD_371_1212_U188 , P2_ADD_371_1212_U132 );
and AND2_27719 ( P2_ADD_371_1212_U15 , P2_ADD_371_1212_U185 , P2_ADD_371_1212_U170 );
and AND2_27720 ( P2_ADD_371_1212_U16 , P2_ADD_371_1212_U191 , P2_ADD_371_1212_U120 );
and AND2_27721 ( P2_ADD_371_1212_U17 , P2_ADD_371_1212_U200 , P2_ADD_371_1212_U114 );
and AND2_27722 ( P2_ADD_371_1212_U18 , P2_ADD_371_1212_U194 , P2_ADD_371_1212_U174 );
and AND2_27723 ( P2_ADD_371_1212_U19 , P2_ADD_371_1212_U183 , P2_ADD_371_1212_U131 );
and AND2_27724 ( P2_ADD_371_1212_U20 , P2_ADD_371_1212_U187 , P2_ADD_371_1212_U176 );
and AND2_27725 ( P2_ADD_371_1212_U21 , P2_ADD_371_1212_U192 , P2_ADD_371_1212_U113 );
and AND2_27726 ( P2_ADD_371_1212_U22 , P2_ADD_371_1212_U190 , P2_ADD_371_1212_U123 );
and AND2_27727 ( P2_ADD_371_1212_U23 , P2_ADD_371_1212_U198 , P2_ADD_371_1212_U180 );
and AND2_27728 ( P2_ADD_371_1212_U24 , P2_ADD_371_1212_U182 , P2_ADD_371_1212_U112 );
nand NAND3_27729 ( P2_ADD_371_1212_U25 , P2_ADD_371_1212_U269 , P2_ADD_371_1212_U268 , P2_ADD_371_1212_U204 );
not NOT1_27730 ( P2_ADD_371_1212_U26 , P2_INSTADDRPOINTER_REG_0_ );
not NOT1_27731 ( P2_ADD_371_1212_U27 , P2_R2256_U21 );
not NOT1_27732 ( P2_ADD_371_1212_U28 , P2_INSTADDRPOINTER_REG_1_ );
nand NAND2_27733 ( P2_ADD_371_1212_U29 , P2_R2256_U21 , P2_INSTADDRPOINTER_REG_0_ );
not NOT1_27734 ( P2_ADD_371_1212_U30 , P2_R2256_U4 );
not NOT1_27735 ( P2_ADD_371_1212_U31 , P2_R2256_U22 );
not NOT1_27736 ( P2_ADD_371_1212_U32 , P2_INSTADDRPOINTER_REG_2_ );
not NOT1_27737 ( P2_ADD_371_1212_U33 , P2_R2256_U26 );
not NOT1_27738 ( P2_ADD_371_1212_U34 , P2_INSTADDRPOINTER_REG_3_ );
not NOT1_27739 ( P2_ADD_371_1212_U35 , P2_R2256_U20 );
not NOT1_27740 ( P2_ADD_371_1212_U36 , P2_INSTADDRPOINTER_REG_4_ );
not NOT1_27741 ( P2_ADD_371_1212_U37 , P2_R2256_U19 );
not NOT1_27742 ( P2_ADD_371_1212_U38 , P2_INSTADDRPOINTER_REG_5_ );
not NOT1_27743 ( P2_ADD_371_1212_U39 , P2_INSTADDRPOINTER_REG_6_ );
not NOT1_27744 ( P2_ADD_371_1212_U40 , P2_R2256_U18 );
not NOT1_27745 ( P2_ADD_371_1212_U41 , P2_R2256_U5 );
not NOT1_27746 ( P2_ADD_371_1212_U42 , P2_INSTADDRPOINTER_REG_8_ );
not NOT1_27747 ( P2_ADD_371_1212_U43 , P2_R2256_U17 );
not NOT1_27748 ( P2_ADD_371_1212_U44 , P2_INSTADDRPOINTER_REG_7_ );
not NOT1_27749 ( P2_ADD_371_1212_U45 , P2_INSTADDRPOINTER_REG_9_ );
not NOT1_27750 ( P2_ADD_371_1212_U46 , P2_INSTADDRPOINTER_REG_10_ );
not NOT1_27751 ( P2_ADD_371_1212_U47 , P2_INSTADDRPOINTER_REG_11_ );
not NOT1_27752 ( P2_ADD_371_1212_U48 , P2_INSTADDRPOINTER_REG_12_ );
not NOT1_27753 ( P2_ADD_371_1212_U49 , P2_INSTADDRPOINTER_REG_13_ );
not NOT1_27754 ( P2_ADD_371_1212_U50 , P2_INSTADDRPOINTER_REG_14_ );
not NOT1_27755 ( P2_ADD_371_1212_U51 , P2_INSTADDRPOINTER_REG_15_ );
not NOT1_27756 ( P2_ADD_371_1212_U52 , P2_INSTADDRPOINTER_REG_16_ );
not NOT1_27757 ( P2_ADD_371_1212_U53 , P2_INSTADDRPOINTER_REG_18_ );
not NOT1_27758 ( P2_ADD_371_1212_U54 , P2_INSTADDRPOINTER_REG_17_ );
not NOT1_27759 ( P2_ADD_371_1212_U55 , P2_INSTADDRPOINTER_REG_19_ );
not NOT1_27760 ( P2_ADD_371_1212_U56 , P2_INSTADDRPOINTER_REG_20_ );
not NOT1_27761 ( P2_ADD_371_1212_U57 , P2_INSTADDRPOINTER_REG_21_ );
not NOT1_27762 ( P2_ADD_371_1212_U58 , P2_INSTADDRPOINTER_REG_22_ );
not NOT1_27763 ( P2_ADD_371_1212_U59 , P2_INSTADDRPOINTER_REG_23_ );
not NOT1_27764 ( P2_ADD_371_1212_U60 , P2_INSTADDRPOINTER_REG_24_ );
not NOT1_27765 ( P2_ADD_371_1212_U61 , P2_INSTADDRPOINTER_REG_26_ );
not NOT1_27766 ( P2_ADD_371_1212_U62 , P2_INSTADDRPOINTER_REG_25_ );
not NOT1_27767 ( P2_ADD_371_1212_U63 , P2_INSTADDRPOINTER_REG_27_ );
not NOT1_27768 ( P2_ADD_371_1212_U64 , P2_INSTADDRPOINTER_REG_28_ );
not NOT1_27769 ( P2_ADD_371_1212_U65 , P2_INSTADDRPOINTER_REG_29_ );
not NOT1_27770 ( P2_ADD_371_1212_U66 , P2_INSTADDRPOINTER_REG_30_ );
nand NAND2_27771 ( P2_ADD_371_1212_U67 , P2_R2256_U4 , P2_ADD_371_1212_U137 );
nand NAND2_27772 ( P2_ADD_371_1212_U68 , P2_ADD_371_1212_U206 , P2_ADD_371_1212_U205 );
nand NAND2_27773 ( P2_ADD_371_1212_U69 , P2_ADD_371_1212_U215 , P2_ADD_371_1212_U214 );
nand NAND2_27774 ( P2_ADD_371_1212_U70 , P2_ADD_371_1212_U217 , P2_ADD_371_1212_U216 );
nand NAND2_27775 ( P2_ADD_371_1212_U71 , P2_ADD_371_1212_U219 , P2_ADD_371_1212_U218 );
nand NAND2_27776 ( P2_ADD_371_1212_U72 , P2_ADD_371_1212_U230 , P2_ADD_371_1212_U229 );
nand NAND2_27777 ( P2_ADD_371_1212_U73 , P2_ADD_371_1212_U232 , P2_ADD_371_1212_U231 );
nand NAND2_27778 ( P2_ADD_371_1212_U74 , P2_ADD_371_1212_U241 , P2_ADD_371_1212_U240 );
nand NAND2_27779 ( P2_ADD_371_1212_U75 , P2_ADD_371_1212_U271 , P2_ADD_371_1212_U270 );
nand NAND2_27780 ( P2_ADD_371_1212_U76 , P2_ADD_371_1212_U273 , P2_ADD_371_1212_U272 );
nand NAND2_27781 ( P2_ADD_371_1212_U77 , P2_ADD_371_1212_U282 , P2_ADD_371_1212_U281 );
nand NAND2_27782 ( P2_ADD_371_1212_U78 , P2_ADD_371_1212_U213 , P2_ADD_371_1212_U212 );
nand NAND2_27783 ( P2_ADD_371_1212_U79 , P2_ADD_371_1212_U226 , P2_ADD_371_1212_U225 );
nand NAND2_27784 ( P2_ADD_371_1212_U80 , P2_ADD_371_1212_U239 , P2_ADD_371_1212_U238 );
nand NAND2_27785 ( P2_ADD_371_1212_U81 , P2_ADD_371_1212_U248 , P2_ADD_371_1212_U247 );
nand NAND2_27786 ( P2_ADD_371_1212_U82 , P2_ADD_371_1212_U255 , P2_ADD_371_1212_U254 );
nand NAND2_27787 ( P2_ADD_371_1212_U83 , P2_ADD_371_1212_U257 , P2_ADD_371_1212_U256 );
nand NAND2_27788 ( P2_ADD_371_1212_U84 , P2_ADD_371_1212_U264 , P2_ADD_371_1212_U263 );
nand NAND2_27789 ( P2_ADD_371_1212_U85 , P2_ADD_371_1212_U280 , P2_ADD_371_1212_U279 );
and AND2_27790 ( P2_ADD_371_1212_U86 , P2_ADD_371_1212_U203 , P2_ADD_371_1212_U166 );
and AND3_27791 ( P2_ADD_371_1212_U87 , P2_INSTADDRPOINTER_REG_15_ , P2_INSTADDRPOINTER_REG_14_ , P2_INSTADDRPOINTER_REG_13_ );
and AND3_27792 ( P2_ADD_371_1212_U88 , P2_INSTADDRPOINTER_REG_17_ , P2_INSTADDRPOINTER_REG_18_ , P2_INSTADDRPOINTER_REG_16_ );
and AND2_27793 ( P2_ADD_371_1212_U89 , P2_INSTADDRPOINTER_REG_19_ , P2_INSTADDRPOINTER_REG_20_ );
and AND3_27794 ( P2_ADD_371_1212_U90 , P2_INSTADDRPOINTER_REG_23_ , P2_INSTADDRPOINTER_REG_22_ , P2_INSTADDRPOINTER_REG_21_ );
and AND3_27795 ( P2_ADD_371_1212_U91 , P2_INSTADDRPOINTER_REG_25_ , P2_INSTADDRPOINTER_REG_26_ , P2_INSTADDRPOINTER_REG_24_ );
and AND3_27796 ( P2_ADD_371_1212_U92 , P2_INSTADDRPOINTER_REG_29_ , P2_INSTADDRPOINTER_REG_28_ , P2_INSTADDRPOINTER_REG_27_ );
and AND2_27797 ( P2_ADD_371_1212_U93 , P2_ADD_371_1212_U8 , P2_ADD_371_1212_U94 );
and AND2_27798 ( P2_ADD_371_1212_U94 , P2_INSTADDRPOINTER_REG_28_ , P2_INSTADDRPOINTER_REG_27_ );
and AND2_27799 ( P2_ADD_371_1212_U95 , P2_ADD_371_1212_U7 , P2_INSTADDRPOINTER_REG_16_ );
and AND2_27800 ( P2_ADD_371_1212_U96 , P2_ADD_371_1212_U11 , P2_INSTADDRPOINTER_REG_19_ );
and AND2_27801 ( P2_ADD_371_1212_U97 , P2_ADD_371_1212_U6 , P2_ADD_371_1212_U98 );
and AND2_27802 ( P2_ADD_371_1212_U98 , P2_INSTADDRPOINTER_REG_22_ , P2_INSTADDRPOINTER_REG_21_ );
and AND2_27803 ( P2_ADD_371_1212_U99 , P2_ADD_371_1212_U6 , P2_INSTADDRPOINTER_REG_21_ );
and AND2_27804 ( P2_ADD_371_1212_U100 , P2_ADD_371_1212_U7 , P2_ADD_371_1212_U101 );
and AND2_27805 ( P2_ADD_371_1212_U101 , P2_INSTADDRPOINTER_REG_17_ , P2_INSTADDRPOINTER_REG_16_ );
and AND2_27806 ( P2_ADD_371_1212_U102 , P2_INSTADDRPOINTER_REG_11_ , P2_ADD_371_1212_U5 );
and AND2_27807 ( P2_ADD_371_1212_U103 , P2_ADD_371_1212_U9 , P2_ADD_371_1212_U104 );
and AND2_27808 ( P2_ADD_371_1212_U104 , P2_INSTADDRPOINTER_REG_25_ , P2_INSTADDRPOINTER_REG_24_ );
and AND2_27809 ( P2_ADD_371_1212_U105 , P2_INSTADDRPOINTER_REG_14_ , P2_ADD_371_1212_U4 );
and AND2_27810 ( P2_ADD_371_1212_U106 , P2_ADD_371_1212_U12 , P2_INSTADDRPOINTER_REG_30_ );
and AND2_27811 ( P2_ADD_371_1212_U107 , P2_ADD_371_1212_U12 , P2_INSTADDRPOINTER_REG_30_ );
and AND2_27812 ( P2_ADD_371_1212_U108 , P2_ADD_371_1212_U8 , P2_INSTADDRPOINTER_REG_27_ );
and AND2_27813 ( P2_ADD_371_1212_U109 , P2_ADD_371_1212_U9 , P2_INSTADDRPOINTER_REG_24_ );
and AND2_27814 ( P2_ADD_371_1212_U110 , P2_ADD_371_1212_U208 , P2_ADD_371_1212_U207 );
nand NAND2_27815 ( P2_ADD_371_1212_U111 , P2_ADD_371_1212_U155 , P2_ADD_371_1212_U154 );
nand NAND2_27816 ( P2_ADD_371_1212_U112 , P2_ADD_371_1212_U12 , P2_ADD_371_1212_U117 );
nand NAND2_27817 ( P2_ADD_371_1212_U113 , P2_ADD_371_1212_U9 , P2_ADD_371_1212_U117 );
nand NAND2_27818 ( P2_ADD_371_1212_U114 , P2_ADD_371_1212_U95 , P2_ADD_371_1212_U117 );
and AND2_27819 ( P2_ADD_371_1212_U115 , P2_ADD_371_1212_U221 , P2_ADD_371_1212_U220 );
nand NAND2_27820 ( P2_ADD_371_1212_U116 , P2_ADD_371_1212_U67 , P2_ADD_371_1212_U139 );
nand NAND2_27821 ( P2_ADD_371_1212_U117 , P2_ADD_371_1212_U86 , P2_ADD_371_1212_U202 );
and AND2_27822 ( P2_ADD_371_1212_U118 , P2_ADD_371_1212_U228 , P2_ADD_371_1212_U227 );
nand NAND2_27823 ( P2_ADD_371_1212_U119 , P2_ADD_371_1212_U117 , P2_ADD_371_1212_U100 );
nand NAND2_27824 ( P2_ADD_371_1212_U120 , P2_ADD_371_1212_U105 , P2_ADD_371_1212_U117 );
and AND2_27825 ( P2_ADD_371_1212_U121 , P2_ADD_371_1212_U234 , P2_ADD_371_1212_U233 );
nand NAND2_27826 ( P2_ADD_371_1212_U122 , P2_ADD_371_1212_U147 , P2_ADD_371_1212_U146 );
nand NAND2_27827 ( P2_ADD_371_1212_U123 , P2_ADD_371_1212_U8 , P2_ADD_371_1212_U117 );
and AND2_27828 ( P2_ADD_371_1212_U124 , P2_ADD_371_1212_U243 , P2_ADD_371_1212_U242 );
nand NAND2_27829 ( P2_ADD_371_1212_U125 , P2_ADD_371_1212_U151 , P2_ADD_371_1212_U150 );
and AND2_27830 ( P2_ADD_371_1212_U126 , P2_ADD_371_1212_U250 , P2_ADD_371_1212_U249 );
nand NAND2_27831 ( P2_ADD_371_1212_U127 , P2_ADD_371_1212_U163 , P2_ADD_371_1212_U162 );
not NOT1_27832 ( P2_ADD_371_1212_U128 , P2_INSTADDRPOINTER_REG_31_ );
and AND2_27833 ( P2_ADD_371_1212_U129 , P2_ADD_371_1212_U259 , P2_ADD_371_1212_U258 );
nand NAND2_27834 ( P2_ADD_371_1212_U130 , P2_ADD_371_1212_U143 , P2_ADD_371_1212_U142 );
nand NAND2_27835 ( P2_ADD_371_1212_U131 , P2_ADD_371_1212_U6 , P2_ADD_371_1212_U117 );
nand NAND2_27836 ( P2_ADD_371_1212_U132 , P2_ADD_371_1212_U102 , P2_ADD_371_1212_U117 );
and AND2_27837 ( P2_ADD_371_1212_U133 , P2_ADD_371_1212_U275 , P2_ADD_371_1212_U274 );
nand NAND2_27838 ( P2_ADD_371_1212_U134 , P2_ADD_371_1212_U159 , P2_ADD_371_1212_U158 );
nand NAND2_27839 ( P2_ADD_371_1212_U135 , P2_ADD_371_1212_U109 , P2_ADD_371_1212_U117 );
not NOT1_27840 ( P2_ADD_371_1212_U136 , P2_ADD_371_1212_U67 );
not NOT1_27841 ( P2_ADD_371_1212_U137 , P2_ADD_371_1212_U29 );
nand NAND2_27842 ( P2_ADD_371_1212_U138 , P2_ADD_371_1212_U30 , P2_ADD_371_1212_U29 );
nand NAND2_27843 ( P2_ADD_371_1212_U139 , P2_INSTADDRPOINTER_REG_1_ , P2_ADD_371_1212_U138 );
not NOT1_27844 ( P2_ADD_371_1212_U140 , P2_ADD_371_1212_U116 );
or OR2_27845 ( P2_ADD_371_1212_U141 , P2_R2256_U22 , P2_INSTADDRPOINTER_REG_2_ );
nand NAND2_27846 ( P2_ADD_371_1212_U142 , P2_ADD_371_1212_U141 , P2_ADD_371_1212_U116 );
nand NAND2_27847 ( P2_ADD_371_1212_U143 , P2_INSTADDRPOINTER_REG_2_ , P2_R2256_U22 );
not NOT1_27848 ( P2_ADD_371_1212_U144 , P2_ADD_371_1212_U130 );
or OR2_27849 ( P2_ADD_371_1212_U145 , P2_R2256_U26 , P2_INSTADDRPOINTER_REG_3_ );
nand NAND2_27850 ( P2_ADD_371_1212_U146 , P2_ADD_371_1212_U145 , P2_ADD_371_1212_U130 );
nand NAND2_27851 ( P2_ADD_371_1212_U147 , P2_INSTADDRPOINTER_REG_3_ , P2_R2256_U26 );
not NOT1_27852 ( P2_ADD_371_1212_U148 , P2_ADD_371_1212_U122 );
or OR2_27853 ( P2_ADD_371_1212_U149 , P2_R2256_U20 , P2_INSTADDRPOINTER_REG_4_ );
nand NAND2_27854 ( P2_ADD_371_1212_U150 , P2_ADD_371_1212_U149 , P2_ADD_371_1212_U122 );
nand NAND2_27855 ( P2_ADD_371_1212_U151 , P2_INSTADDRPOINTER_REG_4_ , P2_R2256_U20 );
not NOT1_27856 ( P2_ADD_371_1212_U152 , P2_ADD_371_1212_U125 );
or OR2_27857 ( P2_ADD_371_1212_U153 , P2_R2256_U19 , P2_INSTADDRPOINTER_REG_5_ );
nand NAND2_27858 ( P2_ADD_371_1212_U154 , P2_ADD_371_1212_U153 , P2_ADD_371_1212_U125 );
nand NAND2_27859 ( P2_ADD_371_1212_U155 , P2_INSTADDRPOINTER_REG_5_ , P2_R2256_U19 );
not NOT1_27860 ( P2_ADD_371_1212_U156 , P2_ADD_371_1212_U111 );
or OR2_27861 ( P2_ADD_371_1212_U157 , P2_R2256_U18 , P2_INSTADDRPOINTER_REG_6_ );
nand NAND2_27862 ( P2_ADD_371_1212_U158 , P2_ADD_371_1212_U157 , P2_ADD_371_1212_U111 );
nand NAND2_27863 ( P2_ADD_371_1212_U159 , P2_R2256_U18 , P2_INSTADDRPOINTER_REG_6_ );
not NOT1_27864 ( P2_ADD_371_1212_U160 , P2_ADD_371_1212_U134 );
or OR2_27865 ( P2_ADD_371_1212_U161 , P2_R2256_U17 , P2_INSTADDRPOINTER_REG_7_ );
nand NAND2_27866 ( P2_ADD_371_1212_U162 , P2_ADD_371_1212_U161 , P2_ADD_371_1212_U134 );
nand NAND2_27867 ( P2_ADD_371_1212_U163 , P2_INSTADDRPOINTER_REG_7_ , P2_R2256_U17 );
not NOT1_27868 ( P2_ADD_371_1212_U164 , P2_ADD_371_1212_U127 );
or OR2_27869 ( P2_ADD_371_1212_U165 , P2_R2256_U5 , P2_INSTADDRPOINTER_REG_8_ );
nand NAND2_27870 ( P2_ADD_371_1212_U166 , P2_INSTADDRPOINTER_REG_8_ , P2_R2256_U5 );
not NOT1_27871 ( P2_ADD_371_1212_U167 , P2_ADD_371_1212_U117 );
nand NAND2_27872 ( P2_ADD_371_1212_U168 , P2_ADD_371_1212_U5 , P2_ADD_371_1212_U117 );
not NOT1_27873 ( P2_ADD_371_1212_U169 , P2_ADD_371_1212_U132 );
nand NAND2_27874 ( P2_ADD_371_1212_U170 , P2_ADD_371_1212_U4 , P2_ADD_371_1212_U117 );
not NOT1_27875 ( P2_ADD_371_1212_U171 , P2_ADD_371_1212_U120 );
not NOT1_27876 ( P2_ADD_371_1212_U172 , P2_ADD_371_1212_U114 );
not NOT1_27877 ( P2_ADD_371_1212_U173 , P2_ADD_371_1212_U119 );
nand NAND2_27878 ( P2_ADD_371_1212_U174 , P2_ADD_371_1212_U96 , P2_ADD_371_1212_U117 );
not NOT1_27879 ( P2_ADD_371_1212_U175 , P2_ADD_371_1212_U131 );
nand NAND2_27880 ( P2_ADD_371_1212_U176 , P2_ADD_371_1212_U117 , P2_ADD_371_1212_U97 );
not NOT1_27881 ( P2_ADD_371_1212_U177 , P2_ADD_371_1212_U113 );
not NOT1_27882 ( P2_ADD_371_1212_U178 , P2_ADD_371_1212_U135 );
not NOT1_27883 ( P2_ADD_371_1212_U179 , P2_ADD_371_1212_U123 );
nand NAND2_27884 ( P2_ADD_371_1212_U180 , P2_ADD_371_1212_U117 , P2_ADD_371_1212_U93 );
not NOT1_27885 ( P2_ADD_371_1212_U181 , P2_ADD_371_1212_U112 );
nand NAND2_27886 ( P2_ADD_371_1212_U182 , P2_ADD_371_1212_U65 , P2_ADD_371_1212_U180 );
nand NAND2_27887 ( P2_ADD_371_1212_U183 , P2_ADD_371_1212_U56 , P2_ADD_371_1212_U174 );
nand NAND2_27888 ( P2_ADD_371_1212_U184 , P2_ADD_371_1212_U10 , P2_ADD_371_1212_U117 );
nand NAND2_27889 ( P2_ADD_371_1212_U185 , P2_ADD_371_1212_U49 , P2_ADD_371_1212_U184 );
nand NAND2_27890 ( P2_ADD_371_1212_U186 , P2_ADD_371_1212_U99 , P2_ADD_371_1212_U117 );
nand NAND2_27891 ( P2_ADD_371_1212_U187 , P2_ADD_371_1212_U58 , P2_ADD_371_1212_U186 );
nand NAND2_27892 ( P2_ADD_371_1212_U188 , P2_ADD_371_1212_U47 , P2_ADD_371_1212_U168 );
nand NAND2_27893 ( P2_ADD_371_1212_U189 , P2_ADD_371_1212_U117 , P2_ADD_371_1212_U103 );
nand NAND2_27894 ( P2_ADD_371_1212_U190 , P2_ADD_371_1212_U61 , P2_ADD_371_1212_U189 );
nand NAND2_27895 ( P2_ADD_371_1212_U191 , P2_ADD_371_1212_U50 , P2_ADD_371_1212_U170 );
nand NAND2_27896 ( P2_ADD_371_1212_U192 , P2_ADD_371_1212_U59 , P2_ADD_371_1212_U176 );
nand NAND2_27897 ( P2_ADD_371_1212_U193 , P2_ADD_371_1212_U11 , P2_ADD_371_1212_U117 );
nand NAND2_27898 ( P2_ADD_371_1212_U194 , P2_ADD_371_1212_U55 , P2_ADD_371_1212_U193 );
nand NAND2_27899 ( P2_ADD_371_1212_U195 , P2_INSTADDRPOINTER_REG_9_ , P2_ADD_371_1212_U117 );
nand NAND2_27900 ( P2_ADD_371_1212_U196 , P2_ADD_371_1212_U46 , P2_ADD_371_1212_U195 );
nand NAND2_27901 ( P2_ADD_371_1212_U197 , P2_ADD_371_1212_U108 , P2_ADD_371_1212_U117 );
nand NAND2_27902 ( P2_ADD_371_1212_U198 , P2_ADD_371_1212_U64 , P2_ADD_371_1212_U197 );
nand NAND2_27903 ( P2_ADD_371_1212_U199 , P2_ADD_371_1212_U7 , P2_ADD_371_1212_U117 );
nand NAND2_27904 ( P2_ADD_371_1212_U200 , P2_ADD_371_1212_U52 , P2_ADD_371_1212_U199 );
nand NAND2_27905 ( P2_ADD_371_1212_U201 , P2_ADD_371_1212_U107 , P2_ADD_371_1212_U117 );
nand NAND3_27906 ( P2_ADD_371_1212_U202 , P2_ADD_371_1212_U165 , P2_ADD_371_1212_U134 , P2_ADD_371_1212_U161 );
nand NAND3_27907 ( P2_ADD_371_1212_U203 , P2_INSTADDRPOINTER_REG_7_ , P2_ADD_371_1212_U165 , P2_R2256_U17 );
nand NAND2_27908 ( P2_ADD_371_1212_U204 , P2_ADD_371_1212_U136 , P2_INSTADDRPOINTER_REG_1_ );
nand NAND2_27909 ( P2_ADD_371_1212_U205 , P2_INSTADDRPOINTER_REG_0_ , P2_ADD_371_1212_U27 );
nand NAND2_27910 ( P2_ADD_371_1212_U206 , P2_R2256_U21 , P2_ADD_371_1212_U26 );
nand NAND2_27911 ( P2_ADD_371_1212_U207 , P2_INSTADDRPOINTER_REG_6_ , P2_ADD_371_1212_U40 );
nand NAND2_27912 ( P2_ADD_371_1212_U208 , P2_R2256_U18 , P2_ADD_371_1212_U39 );
nand NAND2_27913 ( P2_ADD_371_1212_U209 , P2_INSTADDRPOINTER_REG_6_ , P2_ADD_371_1212_U40 );
nand NAND2_27914 ( P2_ADD_371_1212_U210 , P2_R2256_U18 , P2_ADD_371_1212_U39 );
nand NAND2_27915 ( P2_ADD_371_1212_U211 , P2_ADD_371_1212_U210 , P2_ADD_371_1212_U209 );
nand NAND2_27916 ( P2_ADD_371_1212_U212 , P2_ADD_371_1212_U110 , P2_ADD_371_1212_U111 );
nand NAND2_27917 ( P2_ADD_371_1212_U213 , P2_ADD_371_1212_U156 , P2_ADD_371_1212_U211 );
nand NAND2_27918 ( P2_ADD_371_1212_U214 , P2_INSTADDRPOINTER_REG_30_ , P2_ADD_371_1212_U112 );
nand NAND2_27919 ( P2_ADD_371_1212_U215 , P2_ADD_371_1212_U181 , P2_ADD_371_1212_U66 );
nand NAND2_27920 ( P2_ADD_371_1212_U216 , P2_INSTADDRPOINTER_REG_24_ , P2_ADD_371_1212_U113 );
nand NAND2_27921 ( P2_ADD_371_1212_U217 , P2_ADD_371_1212_U177 , P2_ADD_371_1212_U60 );
nand NAND2_27922 ( P2_ADD_371_1212_U218 , P2_INSTADDRPOINTER_REG_17_ , P2_ADD_371_1212_U114 );
nand NAND2_27923 ( P2_ADD_371_1212_U219 , P2_ADD_371_1212_U172 , P2_ADD_371_1212_U54 );
nand NAND2_27924 ( P2_ADD_371_1212_U220 , P2_INSTADDRPOINTER_REG_2_ , P2_ADD_371_1212_U31 );
nand NAND2_27925 ( P2_ADD_371_1212_U221 , P2_R2256_U22 , P2_ADD_371_1212_U32 );
nand NAND2_27926 ( P2_ADD_371_1212_U222 , P2_INSTADDRPOINTER_REG_2_ , P2_ADD_371_1212_U31 );
nand NAND2_27927 ( P2_ADD_371_1212_U223 , P2_R2256_U22 , P2_ADD_371_1212_U32 );
nand NAND2_27928 ( P2_ADD_371_1212_U224 , P2_ADD_371_1212_U223 , P2_ADD_371_1212_U222 );
nand NAND2_27929 ( P2_ADD_371_1212_U225 , P2_ADD_371_1212_U115 , P2_ADD_371_1212_U116 );
nand NAND2_27930 ( P2_ADD_371_1212_U226 , P2_ADD_371_1212_U140 , P2_ADD_371_1212_U224 );
nand NAND2_27931 ( P2_ADD_371_1212_U227 , P2_INSTADDRPOINTER_REG_9_ , P2_ADD_371_1212_U117 );
nand NAND2_27932 ( P2_ADD_371_1212_U228 , P2_ADD_371_1212_U167 , P2_ADD_371_1212_U45 );
nand NAND2_27933 ( P2_ADD_371_1212_U229 , P2_INSTADDRPOINTER_REG_18_ , P2_ADD_371_1212_U119 );
nand NAND2_27934 ( P2_ADD_371_1212_U230 , P2_ADD_371_1212_U173 , P2_ADD_371_1212_U53 );
nand NAND2_27935 ( P2_ADD_371_1212_U231 , P2_INSTADDRPOINTER_REG_15_ , P2_ADD_371_1212_U120 );
nand NAND2_27936 ( P2_ADD_371_1212_U232 , P2_ADD_371_1212_U171 , P2_ADD_371_1212_U51 );
nand NAND2_27937 ( P2_ADD_371_1212_U233 , P2_INSTADDRPOINTER_REG_4_ , P2_ADD_371_1212_U35 );
nand NAND2_27938 ( P2_ADD_371_1212_U234 , P2_R2256_U20 , P2_ADD_371_1212_U36 );
nand NAND2_27939 ( P2_ADD_371_1212_U235 , P2_INSTADDRPOINTER_REG_4_ , P2_ADD_371_1212_U35 );
nand NAND2_27940 ( P2_ADD_371_1212_U236 , P2_R2256_U20 , P2_ADD_371_1212_U36 );
nand NAND2_27941 ( P2_ADD_371_1212_U237 , P2_ADD_371_1212_U236 , P2_ADD_371_1212_U235 );
nand NAND2_27942 ( P2_ADD_371_1212_U238 , P2_ADD_371_1212_U121 , P2_ADD_371_1212_U122 );
nand NAND2_27943 ( P2_ADD_371_1212_U239 , P2_ADD_371_1212_U148 , P2_ADD_371_1212_U237 );
nand NAND2_27944 ( P2_ADD_371_1212_U240 , P2_INSTADDRPOINTER_REG_27_ , P2_ADD_371_1212_U123 );
nand NAND2_27945 ( P2_ADD_371_1212_U241 , P2_ADD_371_1212_U179 , P2_ADD_371_1212_U63 );
nand NAND2_27946 ( P2_ADD_371_1212_U242 , P2_INSTADDRPOINTER_REG_5_ , P2_ADD_371_1212_U37 );
nand NAND2_27947 ( P2_ADD_371_1212_U243 , P2_R2256_U19 , P2_ADD_371_1212_U38 );
nand NAND2_27948 ( P2_ADD_371_1212_U244 , P2_INSTADDRPOINTER_REG_5_ , P2_ADD_371_1212_U37 );
nand NAND2_27949 ( P2_ADD_371_1212_U245 , P2_R2256_U19 , P2_ADD_371_1212_U38 );
nand NAND2_27950 ( P2_ADD_371_1212_U246 , P2_ADD_371_1212_U245 , P2_ADD_371_1212_U244 );
nand NAND2_27951 ( P2_ADD_371_1212_U247 , P2_ADD_371_1212_U124 , P2_ADD_371_1212_U125 );
nand NAND2_27952 ( P2_ADD_371_1212_U248 , P2_ADD_371_1212_U152 , P2_ADD_371_1212_U246 );
nand NAND2_27953 ( P2_ADD_371_1212_U249 , P2_INSTADDRPOINTER_REG_8_ , P2_ADD_371_1212_U41 );
nand NAND2_27954 ( P2_ADD_371_1212_U250 , P2_R2256_U5 , P2_ADD_371_1212_U42 );
nand NAND2_27955 ( P2_ADD_371_1212_U251 , P2_INSTADDRPOINTER_REG_8_ , P2_ADD_371_1212_U41 );
nand NAND2_27956 ( P2_ADD_371_1212_U252 , P2_R2256_U5 , P2_ADD_371_1212_U42 );
nand NAND2_27957 ( P2_ADD_371_1212_U253 , P2_ADD_371_1212_U252 , P2_ADD_371_1212_U251 );
nand NAND2_27958 ( P2_ADD_371_1212_U254 , P2_ADD_371_1212_U126 , P2_ADD_371_1212_U127 );
nand NAND2_27959 ( P2_ADD_371_1212_U255 , P2_ADD_371_1212_U164 , P2_ADD_371_1212_U253 );
nand NAND2_27960 ( P2_ADD_371_1212_U256 , P2_INSTADDRPOINTER_REG_31_ , P2_ADD_371_1212_U201 );
nand NAND3_27961 ( P2_ADD_371_1212_U257 , P2_ADD_371_1212_U106 , P2_ADD_371_1212_U117 , P2_ADD_371_1212_U128 );
nand NAND2_27962 ( P2_ADD_371_1212_U258 , P2_INSTADDRPOINTER_REG_3_ , P2_ADD_371_1212_U33 );
nand NAND2_27963 ( P2_ADD_371_1212_U259 , P2_R2256_U26 , P2_ADD_371_1212_U34 );
nand NAND2_27964 ( P2_ADD_371_1212_U260 , P2_INSTADDRPOINTER_REG_3_ , P2_ADD_371_1212_U33 );
nand NAND2_27965 ( P2_ADD_371_1212_U261 , P2_R2256_U26 , P2_ADD_371_1212_U34 );
nand NAND2_27966 ( P2_ADD_371_1212_U262 , P2_ADD_371_1212_U261 , P2_ADD_371_1212_U260 );
nand NAND2_27967 ( P2_ADD_371_1212_U263 , P2_ADD_371_1212_U129 , P2_ADD_371_1212_U130 );
nand NAND2_27968 ( P2_ADD_371_1212_U264 , P2_ADD_371_1212_U144 , P2_ADD_371_1212_U262 );
nand NAND2_27969 ( P2_ADD_371_1212_U265 , P2_INSTADDRPOINTER_REG_1_ , P2_ADD_371_1212_U29 );
nand NAND2_27970 ( P2_ADD_371_1212_U266 , P2_ADD_371_1212_U137 , P2_ADD_371_1212_U28 );
nand NAND2_27971 ( P2_ADD_371_1212_U267 , P2_ADD_371_1212_U266 , P2_ADD_371_1212_U265 );
nand NAND3_27972 ( P2_ADD_371_1212_U268 , P2_ADD_371_1212_U29 , P2_ADD_371_1212_U28 , P2_R2256_U4 );
nand NAND2_27973 ( P2_ADD_371_1212_U269 , P2_ADD_371_1212_U267 , P2_ADD_371_1212_U30 );
nand NAND2_27974 ( P2_ADD_371_1212_U270 , P2_INSTADDRPOINTER_REG_21_ , P2_ADD_371_1212_U131 );
nand NAND2_27975 ( P2_ADD_371_1212_U271 , P2_ADD_371_1212_U175 , P2_ADD_371_1212_U57 );
nand NAND2_27976 ( P2_ADD_371_1212_U272 , P2_INSTADDRPOINTER_REG_12_ , P2_ADD_371_1212_U132 );
nand NAND2_27977 ( P2_ADD_371_1212_U273 , P2_ADD_371_1212_U169 , P2_ADD_371_1212_U48 );
nand NAND2_27978 ( P2_ADD_371_1212_U274 , P2_INSTADDRPOINTER_REG_7_ , P2_ADD_371_1212_U43 );
nand NAND2_27979 ( P2_ADD_371_1212_U275 , P2_R2256_U17 , P2_ADD_371_1212_U44 );
nand NAND2_27980 ( P2_ADD_371_1212_U276 , P2_INSTADDRPOINTER_REG_7_ , P2_ADD_371_1212_U43 );
nand NAND2_27981 ( P2_ADD_371_1212_U277 , P2_R2256_U17 , P2_ADD_371_1212_U44 );
nand NAND2_27982 ( P2_ADD_371_1212_U278 , P2_ADD_371_1212_U277 , P2_ADD_371_1212_U276 );
nand NAND2_27983 ( P2_ADD_371_1212_U279 , P2_ADD_371_1212_U133 , P2_ADD_371_1212_U134 );
nand NAND2_27984 ( P2_ADD_371_1212_U280 , P2_ADD_371_1212_U160 , P2_ADD_371_1212_U278 );
nand NAND2_27985 ( P2_ADD_371_1212_U281 , P2_INSTADDRPOINTER_REG_25_ , P2_ADD_371_1212_U135 );
nand NAND2_27986 ( P2_ADD_371_1212_U282 , P2_ADD_371_1212_U178 , P2_ADD_371_1212_U62 );
not NOT1_27987 ( P1_R2027_U5 , P1_INSTADDRPOINTER_REG_0_ );
not NOT1_27988 ( P1_R2027_U6 , P1_INSTADDRPOINTER_REG_2_ );
not NOT1_27989 ( P1_R2027_U7 , P1_INSTADDRPOINTER_REG_1_ );
not NOT1_27990 ( P1_R2027_U8 , P1_INSTADDRPOINTER_REG_4_ );
not NOT1_27991 ( P1_R2027_U9 , P1_INSTADDRPOINTER_REG_3_ );
nand NAND3_27992 ( P1_R2027_U10 , P1_INSTADDRPOINTER_REG_2_ , P1_INSTADDRPOINTER_REG_0_ , P1_INSTADDRPOINTER_REG_1_ );
not NOT1_27993 ( P1_R2027_U11 , P1_INSTADDRPOINTER_REG_6_ );
not NOT1_27994 ( P1_R2027_U12 , P1_INSTADDRPOINTER_REG_5_ );
nand NAND2_27995 ( P1_R2027_U13 , P1_R2027_U82 , P1_R2027_U111 );
not NOT1_27996 ( P1_R2027_U14 , P1_INSTADDRPOINTER_REG_8_ );
not NOT1_27997 ( P1_R2027_U15 , P1_INSTADDRPOINTER_REG_7_ );
nand NAND2_27998 ( P1_R2027_U16 , P1_R2027_U83 , P1_R2027_U112 );
nand NAND2_27999 ( P1_R2027_U17 , P1_R2027_U84 , P1_R2027_U118 );
not NOT1_28000 ( P1_R2027_U18 , P1_INSTADDRPOINTER_REG_9_ );
not NOT1_28001 ( P1_R2027_U19 , P1_INSTADDRPOINTER_REG_10_ );
not NOT1_28002 ( P1_R2027_U20 , P1_INSTADDRPOINTER_REG_12_ );
not NOT1_28003 ( P1_R2027_U21 , P1_INSTADDRPOINTER_REG_11_ );
nand NAND2_28004 ( P1_R2027_U22 , P1_R2027_U85 , P1_R2027_U120 );
not NOT1_28005 ( P1_R2027_U23 , P1_INSTADDRPOINTER_REG_14_ );
not NOT1_28006 ( P1_R2027_U24 , P1_INSTADDRPOINTER_REG_13_ );
nand NAND2_28007 ( P1_R2027_U25 , P1_R2027_U86 , P1_R2027_U113 );
not NOT1_28008 ( P1_R2027_U26 , P1_INSTADDRPOINTER_REG_15_ );
nand NAND2_28009 ( P1_R2027_U27 , P1_R2027_U87 , P1_R2027_U119 );
not NOT1_28010 ( P1_R2027_U28 , P1_INSTADDRPOINTER_REG_16_ );
not NOT1_28011 ( P1_R2027_U29 , P1_INSTADDRPOINTER_REG_18_ );
not NOT1_28012 ( P1_R2027_U30 , P1_INSTADDRPOINTER_REG_17_ );
nand NAND2_28013 ( P1_R2027_U31 , P1_R2027_U88 , P1_R2027_U124 );
not NOT1_28014 ( P1_R2027_U32 , P1_INSTADDRPOINTER_REG_20_ );
not NOT1_28015 ( P1_R2027_U33 , P1_INSTADDRPOINTER_REG_19_ );
nand NAND2_28016 ( P1_R2027_U34 , P1_R2027_U89 , P1_R2027_U117 );
not NOT1_28017 ( P1_R2027_U35 , P1_INSTADDRPOINTER_REG_21_ );
nand NAND2_28018 ( P1_R2027_U36 , P1_R2027_U90 , P1_R2027_U114 );
not NOT1_28019 ( P1_R2027_U37 , P1_INSTADDRPOINTER_REG_22_ );
not NOT1_28020 ( P1_R2027_U38 , P1_INSTADDRPOINTER_REG_24_ );
not NOT1_28021 ( P1_R2027_U39 , P1_INSTADDRPOINTER_REG_23_ );
nand NAND2_28022 ( P1_R2027_U40 , P1_R2027_U91 , P1_R2027_U121 );
not NOT1_28023 ( P1_R2027_U41 , P1_INSTADDRPOINTER_REG_26_ );
not NOT1_28024 ( P1_R2027_U42 , P1_INSTADDRPOINTER_REG_25_ );
nand NAND2_28025 ( P1_R2027_U43 , P1_R2027_U92 , P1_R2027_U115 );
not NOT1_28026 ( P1_R2027_U44 , P1_INSTADDRPOINTER_REG_27_ );
not NOT1_28027 ( P1_R2027_U45 , P1_INSTADDRPOINTER_REG_28_ );
nand NAND2_28028 ( P1_R2027_U46 , P1_R2027_U93 , P1_R2027_U116 );
not NOT1_28029 ( P1_R2027_U47 , P1_INSTADDRPOINTER_REG_29_ );
nand NAND2_28030 ( P1_R2027_U48 , P1_R2027_U94 , P1_R2027_U122 );
nand NAND2_28031 ( P1_R2027_U49 , P1_R2027_U123 , P1_INSTADDRPOINTER_REG_29_ );
not NOT1_28032 ( P1_R2027_U50 , P1_INSTADDRPOINTER_REG_30_ );
nand NAND2_28033 ( P1_R2027_U51 , P1_R2027_U142 , P1_R2027_U141 );
nand NAND2_28034 ( P1_R2027_U52 , P1_R2027_U144 , P1_R2027_U143 );
nand NAND2_28035 ( P1_R2027_U53 , P1_R2027_U146 , P1_R2027_U145 );
nand NAND2_28036 ( P1_R2027_U54 , P1_R2027_U148 , P1_R2027_U147 );
nand NAND2_28037 ( P1_R2027_U55 , P1_R2027_U150 , P1_R2027_U149 );
nand NAND2_28038 ( P1_R2027_U56 , P1_R2027_U152 , P1_R2027_U151 );
nand NAND2_28039 ( P1_R2027_U57 , P1_R2027_U154 , P1_R2027_U153 );
nand NAND2_28040 ( P1_R2027_U58 , P1_R2027_U156 , P1_R2027_U155 );
nand NAND2_28041 ( P1_R2027_U59 , P1_R2027_U158 , P1_R2027_U157 );
nand NAND2_28042 ( P1_R2027_U60 , P1_R2027_U160 , P1_R2027_U159 );
nand NAND2_28043 ( P1_R2027_U61 , P1_R2027_U162 , P1_R2027_U161 );
nand NAND2_28044 ( P1_R2027_U62 , P1_R2027_U164 , P1_R2027_U163 );
nand NAND2_28045 ( P1_R2027_U63 , P1_R2027_U166 , P1_R2027_U165 );
nand NAND2_28046 ( P1_R2027_U64 , P1_R2027_U168 , P1_R2027_U167 );
nand NAND2_28047 ( P1_R2027_U65 , P1_R2027_U170 , P1_R2027_U169 );
nand NAND2_28048 ( P1_R2027_U66 , P1_R2027_U172 , P1_R2027_U171 );
nand NAND2_28049 ( P1_R2027_U67 , P1_R2027_U174 , P1_R2027_U173 );
nand NAND2_28050 ( P1_R2027_U68 , P1_R2027_U176 , P1_R2027_U175 );
nand NAND2_28051 ( P1_R2027_U69 , P1_R2027_U178 , P1_R2027_U177 );
nand NAND2_28052 ( P1_R2027_U70 , P1_R2027_U180 , P1_R2027_U179 );
nand NAND2_28053 ( P1_R2027_U71 , P1_R2027_U182 , P1_R2027_U181 );
nand NAND2_28054 ( P1_R2027_U72 , P1_R2027_U184 , P1_R2027_U183 );
nand NAND2_28055 ( P1_R2027_U73 , P1_R2027_U186 , P1_R2027_U185 );
nand NAND2_28056 ( P1_R2027_U74 , P1_R2027_U188 , P1_R2027_U187 );
nand NAND2_28057 ( P1_R2027_U75 , P1_R2027_U190 , P1_R2027_U189 );
nand NAND2_28058 ( P1_R2027_U76 , P1_R2027_U192 , P1_R2027_U191 );
nand NAND2_28059 ( P1_R2027_U77 , P1_R2027_U194 , P1_R2027_U193 );
nand NAND2_28060 ( P1_R2027_U78 , P1_R2027_U196 , P1_R2027_U195 );
nand NAND2_28061 ( P1_R2027_U79 , P1_R2027_U198 , P1_R2027_U197 );
nand NAND2_28062 ( P1_R2027_U80 , P1_R2027_U200 , P1_R2027_U199 );
nand NAND2_28063 ( P1_R2027_U81 , P1_R2027_U202 , P1_R2027_U201 );
and AND2_28064 ( P1_R2027_U82 , P1_INSTADDRPOINTER_REG_3_ , P1_INSTADDRPOINTER_REG_4_ );
and AND2_28065 ( P1_R2027_U83 , P1_INSTADDRPOINTER_REG_5_ , P1_INSTADDRPOINTER_REG_6_ );
and AND2_28066 ( P1_R2027_U84 , P1_INSTADDRPOINTER_REG_7_ , P1_INSTADDRPOINTER_REG_8_ );
and AND2_28067 ( P1_R2027_U85 , P1_INSTADDRPOINTER_REG_9_ , P1_INSTADDRPOINTER_REG_10_ );
and AND2_28068 ( P1_R2027_U86 , P1_INSTADDRPOINTER_REG_11_ , P1_INSTADDRPOINTER_REG_12_ );
and AND2_28069 ( P1_R2027_U87 , P1_INSTADDRPOINTER_REG_13_ , P1_INSTADDRPOINTER_REG_14_ );
and AND2_28070 ( P1_R2027_U88 , P1_INSTADDRPOINTER_REG_16_ , P1_INSTADDRPOINTER_REG_15_ );
and AND2_28071 ( P1_R2027_U89 , P1_INSTADDRPOINTER_REG_17_ , P1_INSTADDRPOINTER_REG_18_ );
and AND2_28072 ( P1_R2027_U90 , P1_INSTADDRPOINTER_REG_19_ , P1_INSTADDRPOINTER_REG_20_ );
and AND2_28073 ( P1_R2027_U91 , P1_INSTADDRPOINTER_REG_22_ , P1_INSTADDRPOINTER_REG_21_ );
and AND2_28074 ( P1_R2027_U92 , P1_INSTADDRPOINTER_REG_23_ , P1_INSTADDRPOINTER_REG_24_ );
and AND2_28075 ( P1_R2027_U93 , P1_INSTADDRPOINTER_REG_25_ , P1_INSTADDRPOINTER_REG_26_ );
and AND2_28076 ( P1_R2027_U94 , P1_INSTADDRPOINTER_REG_28_ , P1_INSTADDRPOINTER_REG_27_ );
nand NAND2_28077 ( P1_R2027_U95 , P1_R2027_U118 , P1_INSTADDRPOINTER_REG_7_ );
nand NAND2_28078 ( P1_R2027_U96 , P1_R2027_U112 , P1_INSTADDRPOINTER_REG_5_ );
nand NAND2_28079 ( P1_R2027_U97 , P1_R2027_U111 , P1_INSTADDRPOINTER_REG_3_ );
not NOT1_28080 ( P1_R2027_U98 , P1_INSTADDRPOINTER_REG_31_ );
nand NAND2_28081 ( P1_R2027_U99 , P1_INSTADDRPOINTER_REG_30_ , P1_R2027_U128 );
nand NAND2_28082 ( P1_R2027_U100 , P1_INSTADDRPOINTER_REG_1_ , P1_INSTADDRPOINTER_REG_0_ );
nand NAND2_28083 ( P1_R2027_U101 , P1_R2027_U122 , P1_INSTADDRPOINTER_REG_27_ );
nand NAND2_28084 ( P1_R2027_U102 , P1_R2027_U116 , P1_INSTADDRPOINTER_REG_25_ );
nand NAND2_28085 ( P1_R2027_U103 , P1_R2027_U115 , P1_INSTADDRPOINTER_REG_23_ );
nand NAND2_28086 ( P1_R2027_U104 , P1_R2027_U121 , P1_INSTADDRPOINTER_REG_21_ );
nand NAND2_28087 ( P1_R2027_U105 , P1_R2027_U114 , P1_INSTADDRPOINTER_REG_19_ );
nand NAND2_28088 ( P1_R2027_U106 , P1_R2027_U117 , P1_INSTADDRPOINTER_REG_17_ );
nand NAND2_28089 ( P1_R2027_U107 , P1_R2027_U124 , P1_INSTADDRPOINTER_REG_15_ );
nand NAND2_28090 ( P1_R2027_U108 , P1_R2027_U119 , P1_INSTADDRPOINTER_REG_13_ );
nand NAND2_28091 ( P1_R2027_U109 , P1_R2027_U113 , P1_INSTADDRPOINTER_REG_11_ );
nand NAND2_28092 ( P1_R2027_U110 , P1_INSTADDRPOINTER_REG_9_ , P1_R2027_U120 );
not NOT1_28093 ( P1_R2027_U111 , P1_R2027_U10 );
not NOT1_28094 ( P1_R2027_U112 , P1_R2027_U13 );
not NOT1_28095 ( P1_R2027_U113 , P1_R2027_U22 );
not NOT1_28096 ( P1_R2027_U114 , P1_R2027_U34 );
not NOT1_28097 ( P1_R2027_U115 , P1_R2027_U40 );
not NOT1_28098 ( P1_R2027_U116 , P1_R2027_U43 );
not NOT1_28099 ( P1_R2027_U117 , P1_R2027_U31 );
not NOT1_28100 ( P1_R2027_U118 , P1_R2027_U16 );
not NOT1_28101 ( P1_R2027_U119 , P1_R2027_U25 );
not NOT1_28102 ( P1_R2027_U120 , P1_R2027_U17 );
not NOT1_28103 ( P1_R2027_U121 , P1_R2027_U36 );
not NOT1_28104 ( P1_R2027_U122 , P1_R2027_U46 );
not NOT1_28105 ( P1_R2027_U123 , P1_R2027_U48 );
not NOT1_28106 ( P1_R2027_U124 , P1_R2027_U27 );
not NOT1_28107 ( P1_R2027_U125 , P1_R2027_U95 );
not NOT1_28108 ( P1_R2027_U126 , P1_R2027_U96 );
not NOT1_28109 ( P1_R2027_U127 , P1_R2027_U97 );
not NOT1_28110 ( P1_R2027_U128 , P1_R2027_U49 );
not NOT1_28111 ( P1_R2027_U129 , P1_R2027_U99 );
not NOT1_28112 ( P1_R2027_U130 , P1_R2027_U100 );
not NOT1_28113 ( P1_R2027_U131 , P1_R2027_U101 );
not NOT1_28114 ( P1_R2027_U132 , P1_R2027_U102 );
not NOT1_28115 ( P1_R2027_U133 , P1_R2027_U103 );
not NOT1_28116 ( P1_R2027_U134 , P1_R2027_U104 );
not NOT1_28117 ( P1_R2027_U135 , P1_R2027_U105 );
not NOT1_28118 ( P1_R2027_U136 , P1_R2027_U106 );
not NOT1_28119 ( P1_R2027_U137 , P1_R2027_U107 );
not NOT1_28120 ( P1_R2027_U138 , P1_R2027_U108 );
not NOT1_28121 ( P1_R2027_U139 , P1_R2027_U109 );
not NOT1_28122 ( P1_R2027_U140 , P1_R2027_U110 );
nand NAND2_28123 ( P1_R2027_U141 , P1_R2027_U120 , P1_R2027_U18 );
nand NAND2_28124 ( P1_R2027_U142 , P1_INSTADDRPOINTER_REG_9_ , P1_R2027_U17 );
nand NAND2_28125 ( P1_R2027_U143 , P1_INSTADDRPOINTER_REG_8_ , P1_R2027_U95 );
nand NAND2_28126 ( P1_R2027_U144 , P1_R2027_U125 , P1_R2027_U14 );
nand NAND2_28127 ( P1_R2027_U145 , P1_R2027_U118 , P1_R2027_U15 );
nand NAND2_28128 ( P1_R2027_U146 , P1_INSTADDRPOINTER_REG_7_ , P1_R2027_U16 );
nand NAND2_28129 ( P1_R2027_U147 , P1_INSTADDRPOINTER_REG_6_ , P1_R2027_U96 );
nand NAND2_28130 ( P1_R2027_U148 , P1_R2027_U126 , P1_R2027_U11 );
nand NAND2_28131 ( P1_R2027_U149 , P1_R2027_U112 , P1_R2027_U12 );
nand NAND2_28132 ( P1_R2027_U150 , P1_INSTADDRPOINTER_REG_5_ , P1_R2027_U13 );
nand NAND2_28133 ( P1_R2027_U151 , P1_INSTADDRPOINTER_REG_4_ , P1_R2027_U97 );
nand NAND2_28134 ( P1_R2027_U152 , P1_R2027_U127 , P1_R2027_U8 );
nand NAND2_28135 ( P1_R2027_U153 , P1_R2027_U111 , P1_R2027_U9 );
nand NAND2_28136 ( P1_R2027_U154 , P1_INSTADDRPOINTER_REG_3_ , P1_R2027_U10 );
nand NAND2_28137 ( P1_R2027_U155 , P1_INSTADDRPOINTER_REG_31_ , P1_R2027_U99 );
nand NAND2_28138 ( P1_R2027_U156 , P1_R2027_U129 , P1_R2027_U98 );
nand NAND2_28139 ( P1_R2027_U157 , P1_INSTADDRPOINTER_REG_30_ , P1_R2027_U49 );
nand NAND2_28140 ( P1_R2027_U158 , P1_R2027_U128 , P1_R2027_U50 );
nand NAND2_28141 ( P1_R2027_U159 , P1_INSTADDRPOINTER_REG_2_ , P1_R2027_U100 );
nand NAND2_28142 ( P1_R2027_U160 , P1_R2027_U130 , P1_R2027_U6 );
nand NAND2_28143 ( P1_R2027_U161 , P1_R2027_U123 , P1_R2027_U47 );
nand NAND2_28144 ( P1_R2027_U162 , P1_INSTADDRPOINTER_REG_29_ , P1_R2027_U48 );
nand NAND2_28145 ( P1_R2027_U163 , P1_INSTADDRPOINTER_REG_28_ , P1_R2027_U101 );
nand NAND2_28146 ( P1_R2027_U164 , P1_R2027_U131 , P1_R2027_U45 );
nand NAND2_28147 ( P1_R2027_U165 , P1_R2027_U122 , P1_R2027_U44 );
nand NAND2_28148 ( P1_R2027_U166 , P1_INSTADDRPOINTER_REG_27_ , P1_R2027_U46 );
nand NAND2_28149 ( P1_R2027_U167 , P1_INSTADDRPOINTER_REG_26_ , P1_R2027_U102 );
nand NAND2_28150 ( P1_R2027_U168 , P1_R2027_U132 , P1_R2027_U41 );
nand NAND2_28151 ( P1_R2027_U169 , P1_R2027_U116 , P1_R2027_U42 );
nand NAND2_28152 ( P1_R2027_U170 , P1_INSTADDRPOINTER_REG_25_ , P1_R2027_U43 );
nand NAND2_28153 ( P1_R2027_U171 , P1_INSTADDRPOINTER_REG_24_ , P1_R2027_U103 );
nand NAND2_28154 ( P1_R2027_U172 , P1_R2027_U133 , P1_R2027_U38 );
nand NAND2_28155 ( P1_R2027_U173 , P1_R2027_U115 , P1_R2027_U39 );
nand NAND2_28156 ( P1_R2027_U174 , P1_INSTADDRPOINTER_REG_23_ , P1_R2027_U40 );
nand NAND2_28157 ( P1_R2027_U175 , P1_INSTADDRPOINTER_REG_22_ , P1_R2027_U104 );
nand NAND2_28158 ( P1_R2027_U176 , P1_R2027_U134 , P1_R2027_U37 );
nand NAND2_28159 ( P1_R2027_U177 , P1_R2027_U121 , P1_R2027_U35 );
nand NAND2_28160 ( P1_R2027_U178 , P1_INSTADDRPOINTER_REG_21_ , P1_R2027_U36 );
nand NAND2_28161 ( P1_R2027_U179 , P1_INSTADDRPOINTER_REG_20_ , P1_R2027_U105 );
nand NAND2_28162 ( P1_R2027_U180 , P1_R2027_U135 , P1_R2027_U32 );
nand NAND2_28163 ( P1_R2027_U181 , P1_INSTADDRPOINTER_REG_0_ , P1_R2027_U7 );
nand NAND2_28164 ( P1_R2027_U182 , P1_INSTADDRPOINTER_REG_1_ , P1_R2027_U5 );
nand NAND2_28165 ( P1_R2027_U183 , P1_R2027_U114 , P1_R2027_U33 );
nand NAND2_28166 ( P1_R2027_U184 , P1_INSTADDRPOINTER_REG_19_ , P1_R2027_U34 );
nand NAND2_28167 ( P1_R2027_U185 , P1_INSTADDRPOINTER_REG_18_ , P1_R2027_U106 );
nand NAND2_28168 ( P1_R2027_U186 , P1_R2027_U136 , P1_R2027_U29 );
nand NAND2_28169 ( P1_R2027_U187 , P1_R2027_U117 , P1_R2027_U30 );
nand NAND2_28170 ( P1_R2027_U188 , P1_INSTADDRPOINTER_REG_17_ , P1_R2027_U31 );
nand NAND2_28171 ( P1_R2027_U189 , P1_INSTADDRPOINTER_REG_16_ , P1_R2027_U107 );
nand NAND2_28172 ( P1_R2027_U190 , P1_R2027_U137 , P1_R2027_U28 );
nand NAND2_28173 ( P1_R2027_U191 , P1_R2027_U124 , P1_R2027_U26 );
nand NAND2_28174 ( P1_R2027_U192 , P1_INSTADDRPOINTER_REG_15_ , P1_R2027_U27 );
nand NAND2_28175 ( P1_R2027_U193 , P1_INSTADDRPOINTER_REG_14_ , P1_R2027_U108 );
nand NAND2_28176 ( P1_R2027_U194 , P1_R2027_U138 , P1_R2027_U23 );
nand NAND2_28177 ( P1_R2027_U195 , P1_R2027_U119 , P1_R2027_U24 );
nand NAND2_28178 ( P1_R2027_U196 , P1_INSTADDRPOINTER_REG_13_ , P1_R2027_U25 );
nand NAND2_28179 ( P1_R2027_U197 , P1_INSTADDRPOINTER_REG_12_ , P1_R2027_U109 );
nand NAND2_28180 ( P1_R2027_U198 , P1_R2027_U139 , P1_R2027_U20 );
nand NAND2_28181 ( P1_R2027_U199 , P1_R2027_U113 , P1_R2027_U21 );
nand NAND2_28182 ( P1_R2027_U200 , P1_INSTADDRPOINTER_REG_11_ , P1_R2027_U22 );
nand NAND2_28183 ( P1_R2027_U201 , P1_INSTADDRPOINTER_REG_10_ , P1_R2027_U110 );
nand NAND2_28184 ( P1_R2027_U202 , P1_R2027_U140 , P1_R2027_U19 );
and AND2_28185 ( P1_R2182_U5 , P1_R2182_U47 , P1_U2740 );
and AND2_28186 ( P1_R2182_U6 , P1_R2182_U60 , P1_R2182_U16 );
not NOT1_28187 ( P1_R2182_U7 , P1_U2744 );
not NOT1_28188 ( P1_R2182_U8 , P1_U3246 );
nand NAND2_28189 ( P1_R2182_U9 , P1_U3246 , P1_U2744 );
not NOT1_28190 ( P1_R2182_U10 , P1_U2742 );
not NOT1_28191 ( P1_R2182_U11 , P1_U2741 );
not NOT1_28192 ( P1_R2182_U12 , P1_U2740 );
nand NAND2_28193 ( P1_R2182_U13 , P1_R2182_U35 , P1_R2182_U41 );
not NOT1_28194 ( P1_R2182_U14 , P1_U2737 );
not NOT1_28195 ( P1_R2182_U15 , P1_U2738 );
nand NAND2_28196 ( P1_R2182_U16 , P1_U2723 , P1_U2739 );
not NOT1_28197 ( P1_R2182_U17 , P1_U2736 );
not NOT1_28198 ( P1_R2182_U18 , P1_U2735 );
nand NAND2_28199 ( P1_R2182_U19 , P1_R2182_U36 , P1_R2182_U49 );
not NOT1_28200 ( P1_R2182_U20 , P1_U2734 );
nand NAND2_28201 ( P1_R2182_U21 , P1_R2182_U37 , P1_R2182_U46 );
nand NAND2_28202 ( P1_R2182_U22 , P1_R2182_U48 , P1_U2734 );
not NOT1_28203 ( P1_R2182_U23 , P1_U2733 );
nand NAND2_28204 ( P1_R2182_U24 , P1_R2182_U64 , P1_R2182_U63 );
nand NAND2_28205 ( P1_R2182_U25 , P1_R2182_U66 , P1_R2182_U65 );
nand NAND2_28206 ( P1_R2182_U26 , P1_R2182_U68 , P1_R2182_U67 );
nand NAND2_28207 ( P1_R2182_U27 , P1_R2182_U72 , P1_R2182_U71 );
nand NAND2_28208 ( P1_R2182_U28 , P1_R2182_U74 , P1_R2182_U73 );
nand NAND2_28209 ( P1_R2182_U29 , P1_R2182_U76 , P1_R2182_U75 );
nand NAND2_28210 ( P1_R2182_U30 , P1_R2182_U78 , P1_R2182_U77 );
nand NAND2_28211 ( P1_R2182_U31 , P1_R2182_U80 , P1_R2182_U79 );
nand NAND2_28212 ( P1_R2182_U32 , P1_R2182_U82 , P1_R2182_U81 );
nand NAND2_28213 ( P1_R2182_U33 , P1_R2182_U84 , P1_R2182_U83 );
nand NAND2_28214 ( P1_R2182_U34 , P1_R2182_U86 , P1_R2182_U85 );
and AND2_28215 ( P1_R2182_U35 , P1_U2742 , P1_U2741 );
and AND2_28216 ( P1_R2182_U36 , P1_U2738 , P1_U2737 );
and AND2_28217 ( P1_R2182_U37 , P1_U2735 , P1_U2736 );
nand NAND2_28218 ( P1_R2182_U38 , P1_U2742 , P1_R2182_U41 );
not NOT1_28219 ( P1_R2182_U39 , P1_U2732 );
nand NAND2_28220 ( P1_R2182_U40 , P1_U2733 , P1_R2182_U56 );
nand NAND2_28221 ( P1_R2182_U41 , P1_R2182_U52 , P1_R2182_U53 );
and AND2_28222 ( P1_R2182_U42 , P1_R2182_U70 , P1_R2182_U69 );
nand NAND2_28223 ( P1_R2182_U43 , P1_R2182_U46 , P1_U2736 );
nand NAND2_28224 ( P1_R2182_U44 , P1_R2182_U49 , P1_U2738 );
nand NAND2_28225 ( P1_R2182_U45 , P1_R2182_U51 , P1_R2182_U62 );
not NOT1_28226 ( P1_R2182_U46 , P1_R2182_U19 );
not NOT1_28227 ( P1_R2182_U47 , P1_R2182_U13 );
not NOT1_28228 ( P1_R2182_U48 , P1_R2182_U21 );
not NOT1_28229 ( P1_R2182_U49 , P1_R2182_U16 );
not NOT1_28230 ( P1_R2182_U50 , P1_R2182_U9 );
or OR2_28231 ( P1_R2182_U51 , P1_U2743 , P1_U2731 );
nand NAND2_28232 ( P1_R2182_U52 , P1_U2731 , P1_U2743 );
nand NAND2_28233 ( P1_R2182_U53 , P1_R2182_U50 , P1_R2182_U51 );
not NOT1_28234 ( P1_R2182_U54 , P1_R2182_U41 );
not NOT1_28235 ( P1_R2182_U55 , P1_R2182_U38 );
not NOT1_28236 ( P1_R2182_U56 , P1_R2182_U22 );
not NOT1_28237 ( P1_R2182_U57 , P1_R2182_U40 );
not NOT1_28238 ( P1_R2182_U58 , P1_R2182_U43 );
not NOT1_28239 ( P1_R2182_U59 , P1_R2182_U44 );
or OR2_28240 ( P1_R2182_U60 , P1_U2739 , P1_U2723 );
not NOT1_28241 ( P1_R2182_U61 , P1_R2182_U45 );
nand NAND2_28242 ( P1_R2182_U62 , P1_U2731 , P1_U2743 );
nand NAND2_28243 ( P1_R2182_U63 , P1_R2182_U47 , P1_R2182_U12 );
nand NAND2_28244 ( P1_R2182_U64 , P1_U2740 , P1_R2182_U13 );
nand NAND2_28245 ( P1_R2182_U65 , P1_U2741 , P1_R2182_U38 );
nand NAND2_28246 ( P1_R2182_U66 , P1_R2182_U55 , P1_R2182_U11 );
nand NAND2_28247 ( P1_R2182_U67 , P1_U2732 , P1_R2182_U40 );
nand NAND2_28248 ( P1_R2182_U68 , P1_R2182_U57 , P1_R2182_U39 );
nand NAND2_28249 ( P1_R2182_U69 , P1_U2742 , P1_R2182_U41 );
nand NAND2_28250 ( P1_R2182_U70 , P1_R2182_U54 , P1_R2182_U10 );
nand NAND2_28251 ( P1_R2182_U71 , P1_U2733 , P1_R2182_U22 );
nand NAND2_28252 ( P1_R2182_U72 , P1_R2182_U56 , P1_R2182_U23 );
nand NAND2_28253 ( P1_R2182_U73 , P1_R2182_U48 , P1_R2182_U20 );
nand NAND2_28254 ( P1_R2182_U74 , P1_U2734 , P1_R2182_U21 );
nand NAND2_28255 ( P1_R2182_U75 , P1_U2735 , P1_R2182_U43 );
nand NAND2_28256 ( P1_R2182_U76 , P1_R2182_U58 , P1_R2182_U18 );
nand NAND2_28257 ( P1_R2182_U77 , P1_R2182_U46 , P1_R2182_U17 );
nand NAND2_28258 ( P1_R2182_U78 , P1_U2736 , P1_R2182_U19 );
nand NAND2_28259 ( P1_R2182_U79 , P1_U2737 , P1_R2182_U44 );
nand NAND2_28260 ( P1_R2182_U80 , P1_R2182_U59 , P1_R2182_U14 );
nand NAND2_28261 ( P1_R2182_U81 , P1_R2182_U49 , P1_R2182_U15 );
nand NAND2_28262 ( P1_R2182_U82 , P1_U2738 , P1_R2182_U16 );
nand NAND2_28263 ( P1_R2182_U83 , P1_R2182_U50 , P1_R2182_U45 );
nand NAND2_28264 ( P1_R2182_U84 , P1_R2182_U61 , P1_R2182_U9 );
nand NAND2_28265 ( P1_R2182_U85 , P1_U3246 , P1_R2182_U7 );
nand NAND2_28266 ( P1_R2182_U86 , P1_U2744 , P1_R2182_U8 );
and AND2_28267 ( P1_R2144_U5 , P1_R2144_U104 , P1_R2144_U103 );
and AND4_28268 ( P1_R2144_U6 , P1_R2144_U36 , P1_R2144_U35 , P1_R2144_U27 , P1_R2144_U29 );
and AND2_28269 ( P1_R2144_U7 , P1_R2144_U104 , P1_R2144_U81 );
and AND2_28270 ( P1_R2144_U8 , P1_R2144_U138 , P1_R2144_U136 );
and AND2_28271 ( P1_R2144_U9 , P1_R2144_U128 , P1_R2144_U127 );
and AND3_28272 ( P1_R2144_U10 , P1_R2144_U213 , P1_R2144_U212 , P1_R2144_U82 );
nand NAND2_28273 ( P1_R2144_U11 , P1_R2144_U144 , P1_R2144_U146 );
not NOT1_28274 ( P1_R2144_U12 , P1_U2355 );
not NOT1_28275 ( P1_R2144_U13 , P1_U2750 );
not NOT1_28276 ( P1_R2144_U14 , P1_U2751 );
not NOT1_28277 ( P1_R2144_U15 , P1_U2752 );
not NOT1_28278 ( P1_R2144_U16 , P1_U2749 );
not NOT1_28279 ( P1_R2144_U17 , P1_U2745 );
not NOT1_28280 ( P1_R2144_U18 , P1_U2748 );
nand NAND2_28281 ( P1_R2144_U19 , P1_U2748 , P1_R2144_U178 );
not NOT1_28282 ( P1_R2144_U20 , P1_U2747 );
nand NAND2_28283 ( P1_R2144_U21 , P1_U2747 , P1_R2144_U170 );
not NOT1_28284 ( P1_R2144_U22 , P1_U2746 );
nand NAND2_28285 ( P1_R2144_U23 , P1_U2746 , P1_R2144_U173 );
nand NAND2_28286 ( P1_R2144_U24 , P1_R2144_U79 , P1_R2144_U63 );
nand NAND2_28287 ( P1_R2144_U25 , P1_R2144_U6 , P1_R2144_U79 );
nand NAND2_28288 ( P1_R2144_U26 , P1_R2144_U65 , P1_R2144_U141 );
nand NAND2_28289 ( P1_R2144_U27 , P1_R2144_U206 , P1_R2144_U205 );
nand NAND2_28290 ( P1_R2144_U28 , P1_R2144_U186 , P1_R2144_U185 );
nand NAND2_28291 ( P1_R2144_U29 , P1_R2144_U203 , P1_R2144_U202 );
nand NAND2_28292 ( P1_R2144_U30 , P1_R2144_U209 , P1_R2144_U208 );
nand NAND2_28293 ( P1_R2144_U31 , P1_R2144_U224 , P1_R2144_U223 );
nand NAND2_28294 ( P1_R2144_U32 , P1_R2144_U221 , P1_R2144_U220 );
nand NAND2_28295 ( P1_R2144_U33 , P1_R2144_U227 , P1_R2144_U226 );
nand NAND2_28296 ( P1_R2144_U34 , P1_R2144_U230 , P1_R2144_U229 );
nand NAND2_28297 ( P1_R2144_U35 , P1_R2144_U233 , P1_R2144_U232 );
nand NAND2_28298 ( P1_R2144_U36 , P1_R2144_U236 , P1_R2144_U235 );
nand NAND2_28299 ( P1_R2144_U37 , P1_R2144_U248 , P1_R2144_U247 );
nand NAND2_28300 ( P1_R2144_U38 , P1_R2144_U250 , P1_R2144_U249 );
nand NAND2_28301 ( P1_R2144_U39 , P1_R2144_U252 , P1_R2144_U251 );
nand NAND2_28302 ( P1_R2144_U40 , P1_R2144_U254 , P1_R2144_U253 );
nand NAND2_28303 ( P1_R2144_U41 , P1_R2144_U256 , P1_R2144_U255 );
nand NAND2_28304 ( P1_R2144_U42 , P1_R2144_U258 , P1_R2144_U257 );
nand NAND2_28305 ( P1_R2144_U43 , P1_R2144_U260 , P1_R2144_U259 );
and AND2_28306 ( P1_R2144_U44 , P1_R2144_U21 , P1_R2144_U105 );
nand NAND2_28307 ( P1_R2144_U45 , P1_R2144_U217 , P1_R2144_U216 );
and AND2_28308 ( P1_R2144_U46 , P1_R2144_U19 , P1_R2144_U106 );
nand NAND2_28309 ( P1_R2144_U47 , P1_R2144_U219 , P1_R2144_U218 );
and AND2_28310 ( P1_R2144_U48 , P1_R2144_U162 , P1_R2144_U109 );
nand NAND2_28311 ( P1_R2144_U49 , P1_R2144_U239 , P1_R2144_U238 );
nand NAND2_28312 ( P1_R2144_U50 , P1_R2144_U246 , P1_R2144_U245 );
and AND2_28313 ( P1_R2144_U51 , P1_R2144_U110 , P1_R2144_U109 );
and AND2_28314 ( P1_R2144_U52 , P1_R2144_U106 , P1_R2144_U105 );
and AND2_28315 ( P1_R2144_U53 , P1_R2144_U7 , P1_R2144_U52 );
and AND4_28316 ( P1_R2144_U54 , P1_R2144_U103 , P1_R2144_U151 , P1_R2144_U153 , P1_R2144_U152 );
and AND2_28317 ( P1_R2144_U55 , P1_R2144_U109 , P1_R2144_U106 );
and AND2_28318 ( P1_R2144_U56 , P1_R2144_U159 , P1_R2144_U19 );
and AND2_28319 ( P1_R2144_U57 , P1_R2144_U156 , P1_R2144_U21 );
and AND3_28320 ( P1_R2144_U58 , P1_R2144_U19 , P1_R2144_U21 , P1_R2144_U159 );
and AND2_28321 ( P1_R2144_U59 , P1_R2144_U5 , P1_R2144_U105 );
and AND2_28322 ( P1_R2144_U60 , P1_R2144_U126 , P1_R2144_U21 );
and AND2_28323 ( P1_R2144_U61 , P1_R2144_U23 , P1_R2144_U81 );
and AND2_28324 ( P1_R2144_U62 , P1_R2144_U111 , P1_R2144_U110 );
and AND2_28325 ( P1_R2144_U63 , P1_R2144_U6 , P1_R2144_U64 );
and AND4_28326 ( P1_R2144_U64 , P1_R2144_U34 , P1_R2144_U33 , P1_R2144_U31 , P1_R2144_U32 );
and AND2_28327 ( P1_R2144_U65 , P1_R2144_U34 , P1_R2144_U33 );
and AND3_28328 ( P1_R2144_U66 , P1_R2144_U36 , P1_R2144_U27 , P1_R2144_U29 );
and AND2_28329 ( P1_R2144_U67 , P1_R2144_U29 , P1_R2144_U27 );
not NOT1_28330 ( P1_R2144_U68 , P1_U2762 );
not NOT1_28331 ( P1_R2144_U69 , P1_U2761 );
not NOT1_28332 ( P1_R2144_U70 , P1_U2763 );
not NOT1_28333 ( P1_R2144_U71 , P1_U2764 );
not NOT1_28334 ( P1_R2144_U72 , P1_U2766 );
not NOT1_28335 ( P1_R2144_U73 , P1_U2767 );
not NOT1_28336 ( P1_R2144_U74 , P1_U2768 );
not NOT1_28337 ( P1_R2144_U75 , P1_U2765 );
not NOT1_28338 ( P1_R2144_U76 , P1_U2760 );
not NOT1_28339 ( P1_R2144_U77 , P1_U2759 );
nand NAND2_28340 ( P1_R2144_U78 , P1_R2144_U29 , P1_R2144_U79 );
nand NAND2_28341 ( P1_R2144_U79 , P1_R2144_U99 , P1_R2144_U54 );
and AND2_28342 ( P1_R2144_U80 , P1_R2144_U211 , P1_R2144_U210 );
nand NAND3_28343 ( P1_R2144_U81 , P1_R2144_U165 , P1_R2144_U164 , P1_R2144_U22 );
and AND2_28344 ( P1_R2144_U82 , P1_R2144_U215 , P1_R2144_U214 );
nand NAND2_28345 ( P1_R2144_U83 , P1_R2144_U56 , P1_R2144_U158 );
nand NAND2_28346 ( P1_R2144_U84 , P1_R2144_U111 , P1_R2144_U118 );
not NOT1_28347 ( P1_R2144_U85 , P1_U2754 );
not NOT1_28348 ( P1_R2144_U86 , P1_U2753 );
not NOT1_28349 ( P1_R2144_U87 , P1_U2755 );
not NOT1_28350 ( P1_R2144_U88 , P1_U2756 );
not NOT1_28351 ( P1_R2144_U89 , P1_U2757 );
not NOT1_28352 ( P1_R2144_U90 , P1_U2758 );
nand NAND2_28353 ( P1_R2144_U91 , P1_R2144_U100 , P1_R2144_U132 );
and AND2_28354 ( P1_R2144_U92 , P1_R2144_U241 , P1_R2144_U240 );
nand NAND2_28355 ( P1_R2144_U93 , P1_R2144_U129 , P1_R2144_U113 );
nand NAND2_28356 ( P1_R2144_U94 , P1_R2144_U143 , P1_R2144_U32 );
nand NAND2_28357 ( P1_R2144_U95 , P1_R2144_U141 , P1_R2144_U34 );
nand NAND2_28358 ( P1_R2144_U96 , P1_R2144_U79 , P1_R2144_U66 );
nand NAND2_28359 ( P1_R2144_U97 , P1_R2144_U67 , P1_R2144_U79 );
nand NAND2_28360 ( P1_R2144_U98 , P1_R2144_U113 , P1_R2144_U112 );
nand NAND2_28361 ( P1_R2144_U99 , P1_R2144_U53 , P1_R2144_U84 );
nand NAND2_28362 ( P1_R2144_U100 , P1_U2751 , P1_R2144_U28 );
not NOT1_28363 ( P1_R2144_U101 , P1_R2144_U24 );
not NOT1_28364 ( P1_R2144_U102 , P1_R2144_U81 );
nand NAND2_28365 ( P1_R2144_U103 , P1_U2745 , P1_R2144_U181 );
nand NAND3_28366 ( P1_R2144_U104 , P1_R2144_U167 , P1_R2144_U166 , P1_R2144_U17 );
nand NAND3_28367 ( P1_R2144_U105 , P1_R2144_U175 , P1_R2144_U174 , P1_R2144_U20 );
nand NAND3_28368 ( P1_R2144_U106 , P1_R2144_U201 , P1_R2144_U200 , P1_R2144_U18 );
not NOT1_28369 ( P1_R2144_U107 , P1_R2144_U21 );
not NOT1_28370 ( P1_R2144_U108 , P1_R2144_U23 );
nand NAND3_28371 ( P1_R2144_U109 , P1_R2144_U194 , P1_R2144_U193 , P1_R2144_U13 );
nand NAND3_28372 ( P1_R2144_U110 , P1_R2144_U196 , P1_R2144_U195 , P1_R2144_U16 );
nand NAND2_28373 ( P1_R2144_U111 , P1_U2749 , P1_R2144_U199 );
nand NAND3_28374 ( P1_R2144_U112 , P1_R2144_U189 , P1_R2144_U188 , P1_R2144_U15 );
nand NAND2_28375 ( P1_R2144_U113 , P1_U2752 , P1_R2144_U192 );
nand NAND2_28376 ( P1_R2144_U114 , P1_R2144_U187 , P1_R2144_U14 );
nand NAND2_28377 ( P1_R2144_U115 , P1_U2355 , P1_R2144_U112 );
nand NAND2_28378 ( P1_R2144_U116 , P1_U2750 , P1_R2144_U184 );
nand NAND2_28379 ( P1_R2144_U117 , P1_R2144_U155 , P1_R2144_U157 );
nand NAND2_28380 ( P1_R2144_U118 , P1_R2144_U51 , P1_R2144_U117 );
not NOT1_28381 ( P1_R2144_U119 , P1_R2144_U84 );
not NOT1_28382 ( P1_R2144_U120 , P1_R2144_U19 );
not NOT1_28383 ( P1_R2144_U121 , P1_R2144_U79 );
not NOT1_28384 ( P1_R2144_U122 , P1_R2144_U78 );
not NOT1_28385 ( P1_R2144_U123 , P1_R2144_U83 );
nand NAND2_28386 ( P1_R2144_U124 , P1_R2144_U83 , P1_R2144_U105 );
nand NAND2_28387 ( P1_R2144_U125 , P1_R2144_U21 , P1_R2144_U124 );
nand NAND2_28388 ( P1_R2144_U126 , P1_R2144_U23 , P1_R2144_U81 );
nand NAND2_28389 ( P1_R2144_U127 , P1_R2144_U60 , P1_R2144_U124 );
nand NAND2_28390 ( P1_R2144_U128 , P1_R2144_U61 , P1_R2144_U125 );
nand NAND2_28391 ( P1_R2144_U129 , P1_U2355 , P1_R2144_U112 );
not NOT1_28392 ( P1_R2144_U130 , P1_R2144_U93 );
nand NAND2_28393 ( P1_R2144_U131 , P1_R2144_U187 , P1_R2144_U14 );
nand NAND2_28394 ( P1_R2144_U132 , P1_R2144_U131 , P1_R2144_U93 );
not NOT1_28395 ( P1_R2144_U133 , P1_R2144_U91 );
nand NAND2_28396 ( P1_R2144_U134 , P1_R2144_U91 , P1_R2144_U109 );
nand NAND2_28397 ( P1_R2144_U135 , P1_R2144_U134 , P1_R2144_U116 );
nand NAND2_28398 ( P1_R2144_U136 , P1_R2144_U62 , P1_R2144_U135 );
nand NAND2_28399 ( P1_R2144_U137 , P1_R2144_U161 , P1_R2144_U110 );
nand NAND3_28400 ( P1_R2144_U138 , P1_R2144_U134 , P1_R2144_U116 , P1_R2144_U137 );
not NOT1_28401 ( P1_R2144_U139 , P1_R2144_U97 );
not NOT1_28402 ( P1_R2144_U140 , P1_R2144_U96 );
not NOT1_28403 ( P1_R2144_U141 , P1_R2144_U25 );
not NOT1_28404 ( P1_R2144_U142 , P1_R2144_U95 );
not NOT1_28405 ( P1_R2144_U143 , P1_R2144_U26 );
nand NAND2_28406 ( P1_R2144_U144 , P1_U2355 , P1_R2144_U24 );
not NOT1_28407 ( P1_R2144_U145 , P1_R2144_U144 );
nand NAND2_28408 ( P1_R2144_U146 , P1_R2144_U101 , P1_R2144_U12 );
not NOT1_28409 ( P1_R2144_U147 , P1_R2144_U94 );
not NOT1_28410 ( P1_R2144_U148 , P1_R2144_U98 );
nand NAND2_28411 ( P1_R2144_U149 , P1_R2144_U21 , P1_R2144_U105 );
nand NAND2_28412 ( P1_R2144_U150 , P1_R2144_U19 , P1_R2144_U106 );
nand NAND3_28413 ( P1_R2144_U151 , P1_R2144_U120 , P1_R2144_U105 , P1_R2144_U7 );
nand NAND2_28414 ( P1_R2144_U152 , P1_R2144_U107 , P1_R2144_U7 );
nand NAND2_28415 ( P1_R2144_U153 , P1_R2144_U108 , P1_R2144_U7 );
nand NAND3_28416 ( P1_R2144_U154 , P1_R2144_U113 , P1_R2144_U115 , P1_R2144_U100 );
nand NAND2_28417 ( P1_R2144_U155 , P1_R2144_U154 , P1_R2144_U114 );
nand NAND2_28418 ( P1_R2144_U156 , P1_R2144_U104 , P1_R2144_U103 );
nand NAND2_28419 ( P1_R2144_U157 , P1_U2750 , P1_R2144_U184 );
nand NAND3_28420 ( P1_R2144_U158 , P1_R2144_U117 , P1_R2144_U110 , P1_R2144_U55 );
nand NAND3_28421 ( P1_R2144_U159 , P1_U2749 , P1_R2144_U106 , P1_R2144_U199 );
nand NAND2_28422 ( P1_R2144_U160 , P1_R2144_U58 , P1_R2144_U158 );
nand NAND2_28423 ( P1_R2144_U161 , P1_U2749 , P1_R2144_U199 );
nand NAND2_28424 ( P1_R2144_U162 , P1_U2750 , P1_R2144_U184 );
nand NAND2_28425 ( P1_R2144_U163 , P1_R2144_U116 , P1_R2144_U109 );
nand NAND2_28426 ( P1_R2144_U164 , P1_U2355 , P1_R2144_U68 );
nand NAND2_28427 ( P1_R2144_U165 , P1_U2762 , P1_R2144_U12 );
nand NAND2_28428 ( P1_R2144_U166 , P1_U2355 , P1_R2144_U69 );
nand NAND2_28429 ( P1_R2144_U167 , P1_U2761 , P1_R2144_U12 );
nand NAND2_28430 ( P1_R2144_U168 , P1_U2355 , P1_R2144_U70 );
nand NAND2_28431 ( P1_R2144_U169 , P1_U2763 , P1_R2144_U12 );
nand NAND2_28432 ( P1_R2144_U170 , P1_R2144_U169 , P1_R2144_U168 );
nand NAND2_28433 ( P1_R2144_U171 , P1_U2355 , P1_R2144_U68 );
nand NAND2_28434 ( P1_R2144_U172 , P1_U2762 , P1_R2144_U12 );
nand NAND2_28435 ( P1_R2144_U173 , P1_R2144_U172 , P1_R2144_U171 );
nand NAND2_28436 ( P1_R2144_U174 , P1_U2355 , P1_R2144_U70 );
nand NAND2_28437 ( P1_R2144_U175 , P1_U2763 , P1_R2144_U12 );
nand NAND2_28438 ( P1_R2144_U176 , P1_U2355 , P1_R2144_U71 );
nand NAND2_28439 ( P1_R2144_U177 , P1_U2764 , P1_R2144_U12 );
nand NAND2_28440 ( P1_R2144_U178 , P1_R2144_U177 , P1_R2144_U176 );
nand NAND2_28441 ( P1_R2144_U179 , P1_U2355 , P1_R2144_U69 );
nand NAND2_28442 ( P1_R2144_U180 , P1_U2761 , P1_R2144_U12 );
nand NAND2_28443 ( P1_R2144_U181 , P1_R2144_U180 , P1_R2144_U179 );
nand NAND2_28444 ( P1_R2144_U182 , P1_U2355 , P1_R2144_U72 );
nand NAND2_28445 ( P1_R2144_U183 , P1_U2766 , P1_R2144_U12 );
nand NAND2_28446 ( P1_R2144_U184 , P1_R2144_U183 , P1_R2144_U182 );
nand NAND2_28447 ( P1_R2144_U185 , P1_U2355 , P1_R2144_U73 );
nand NAND2_28448 ( P1_R2144_U186 , P1_U2767 , P1_R2144_U12 );
not NOT1_28449 ( P1_R2144_U187 , P1_R2144_U28 );
nand NAND2_28450 ( P1_R2144_U188 , P1_U2355 , P1_R2144_U74 );
nand NAND2_28451 ( P1_R2144_U189 , P1_U2768 , P1_R2144_U12 );
nand NAND2_28452 ( P1_R2144_U190 , P1_U2355 , P1_R2144_U74 );
nand NAND2_28453 ( P1_R2144_U191 , P1_U2768 , P1_R2144_U12 );
nand NAND2_28454 ( P1_R2144_U192 , P1_R2144_U191 , P1_R2144_U190 );
nand NAND2_28455 ( P1_R2144_U193 , P1_U2355 , P1_R2144_U72 );
nand NAND2_28456 ( P1_R2144_U194 , P1_U2766 , P1_R2144_U12 );
nand NAND2_28457 ( P1_R2144_U195 , P1_U2355 , P1_R2144_U75 );
nand NAND2_28458 ( P1_R2144_U196 , P1_U2765 , P1_R2144_U12 );
nand NAND2_28459 ( P1_R2144_U197 , P1_U2355 , P1_R2144_U75 );
nand NAND2_28460 ( P1_R2144_U198 , P1_U2765 , P1_R2144_U12 );
nand NAND2_28461 ( P1_R2144_U199 , P1_R2144_U198 , P1_R2144_U197 );
nand NAND2_28462 ( P1_R2144_U200 , P1_U2355 , P1_R2144_U71 );
nand NAND2_28463 ( P1_R2144_U201 , P1_U2764 , P1_R2144_U12 );
nand NAND2_28464 ( P1_R2144_U202 , P1_U2355 , P1_R2144_U76 );
nand NAND2_28465 ( P1_R2144_U203 , P1_U2760 , P1_R2144_U12 );
not NOT1_28466 ( P1_R2144_U204 , P1_R2144_U29 );
nand NAND2_28467 ( P1_R2144_U205 , P1_U2355 , P1_R2144_U77 );
nand NAND2_28468 ( P1_R2144_U206 , P1_U2759 , P1_R2144_U12 );
not NOT1_28469 ( P1_R2144_U207 , P1_R2144_U27 );
nand NAND2_28470 ( P1_R2144_U208 , P1_R2144_U122 , P1_R2144_U207 );
nand NAND2_28471 ( P1_R2144_U209 , P1_R2144_U27 , P1_R2144_U78 );
nand NAND2_28472 ( P1_R2144_U210 , P1_R2144_U121 , P1_R2144_U204 );
nand NAND2_28473 ( P1_R2144_U211 , P1_R2144_U29 , P1_R2144_U79 );
nand NAND3_28474 ( P1_R2144_U212 , P1_R2144_U57 , P1_R2144_U124 , P1_R2144_U23 );
nand NAND2_28475 ( P1_R2144_U213 , P1_R2144_U5 , P1_R2144_U108 );
nand NAND2_28476 ( P1_R2144_U214 , P1_R2144_U102 , P1_R2144_U156 );
nand NAND3_28477 ( P1_R2144_U215 , P1_R2144_U59 , P1_R2144_U160 , P1_R2144_U81 );
nand NAND2_28478 ( P1_R2144_U216 , P1_R2144_U149 , P1_R2144_U83 );
nand NAND2_28479 ( P1_R2144_U217 , P1_R2144_U44 , P1_R2144_U123 );
nand NAND2_28480 ( P1_R2144_U218 , P1_R2144_U150 , P1_R2144_U84 );
nand NAND2_28481 ( P1_R2144_U219 , P1_R2144_U46 , P1_R2144_U119 );
nand NAND2_28482 ( P1_R2144_U220 , P1_U2355 , P1_R2144_U85 );
nand NAND2_28483 ( P1_R2144_U221 , P1_U2754 , P1_R2144_U12 );
not NOT1_28484 ( P1_R2144_U222 , P1_R2144_U32 );
nand NAND2_28485 ( P1_R2144_U223 , P1_U2355 , P1_R2144_U86 );
nand NAND2_28486 ( P1_R2144_U224 , P1_U2753 , P1_R2144_U12 );
not NOT1_28487 ( P1_R2144_U225 , P1_R2144_U31 );
nand NAND2_28488 ( P1_R2144_U226 , P1_U2355 , P1_R2144_U87 );
nand NAND2_28489 ( P1_R2144_U227 , P1_U2755 , P1_R2144_U12 );
not NOT1_28490 ( P1_R2144_U228 , P1_R2144_U33 );
nand NAND2_28491 ( P1_R2144_U229 , P1_U2355 , P1_R2144_U88 );
nand NAND2_28492 ( P1_R2144_U230 , P1_U2756 , P1_R2144_U12 );
not NOT1_28493 ( P1_R2144_U231 , P1_R2144_U34 );
nand NAND2_28494 ( P1_R2144_U232 , P1_U2355 , P1_R2144_U89 );
nand NAND2_28495 ( P1_R2144_U233 , P1_U2757 , P1_R2144_U12 );
not NOT1_28496 ( P1_R2144_U234 , P1_R2144_U35 );
nand NAND2_28497 ( P1_R2144_U235 , P1_U2355 , P1_R2144_U90 );
nand NAND2_28498 ( P1_R2144_U236 , P1_U2758 , P1_R2144_U12 );
not NOT1_28499 ( P1_R2144_U237 , P1_R2144_U36 );
nand NAND2_28500 ( P1_R2144_U238 , P1_R2144_U163 , P1_R2144_U91 );
nand NAND2_28501 ( P1_R2144_U239 , P1_R2144_U48 , P1_R2144_U133 );
nand NAND2_28502 ( P1_R2144_U240 , P1_R2144_U187 , P1_U2751 );
nand NAND2_28503 ( P1_R2144_U241 , P1_R2144_U28 , P1_R2144_U14 );
nand NAND2_28504 ( P1_R2144_U242 , P1_R2144_U187 , P1_U2751 );
nand NAND2_28505 ( P1_R2144_U243 , P1_R2144_U28 , P1_R2144_U14 );
nand NAND2_28506 ( P1_R2144_U244 , P1_R2144_U243 , P1_R2144_U242 );
nand NAND2_28507 ( P1_R2144_U245 , P1_R2144_U92 , P1_R2144_U93 );
nand NAND2_28508 ( P1_R2144_U246 , P1_R2144_U130 , P1_R2144_U244 );
nand NAND2_28509 ( P1_R2144_U247 , P1_R2144_U147 , P1_R2144_U225 );
nand NAND2_28510 ( P1_R2144_U248 , P1_R2144_U31 , P1_R2144_U94 );
nand NAND2_28511 ( P1_R2144_U249 , P1_R2144_U222 , P1_R2144_U143 );
nand NAND2_28512 ( P1_R2144_U250 , P1_R2144_U32 , P1_R2144_U26 );
nand NAND2_28513 ( P1_R2144_U251 , P1_R2144_U142 , P1_R2144_U228 );
nand NAND2_28514 ( P1_R2144_U252 , P1_R2144_U33 , P1_R2144_U95 );
nand NAND2_28515 ( P1_R2144_U253 , P1_R2144_U231 , P1_R2144_U141 );
nand NAND2_28516 ( P1_R2144_U254 , P1_R2144_U34 , P1_R2144_U25 );
nand NAND2_28517 ( P1_R2144_U255 , P1_R2144_U140 , P1_R2144_U234 );
nand NAND2_28518 ( P1_R2144_U256 , P1_R2144_U35 , P1_R2144_U96 );
nand NAND2_28519 ( P1_R2144_U257 , P1_R2144_U139 , P1_R2144_U237 );
nand NAND2_28520 ( P1_R2144_U258 , P1_R2144_U36 , P1_R2144_U97 );
nand NAND2_28521 ( P1_R2144_U259 , P1_U2355 , P1_R2144_U98 );
nand NAND2_28522 ( P1_R2144_U260 , P1_R2144_U148 , P1_R2144_U12 );
and AND2_28523 ( P1_R2278_U5 , P1_R2278_U466 , P1_R2278_U327 );
and AND2_28524 ( P1_R2278_U6 , P1_R2278_U292 , P1_R2278_U288 );
and AND2_28525 ( P1_R2278_U7 , P1_R2278_U6 , P1_R2278_U295 );
and AND3_28526 ( P1_R2278_U8 , P1_R2278_U302 , P1_R2278_U298 , P1_R2278_U305 );
and AND2_28527 ( P1_R2278_U9 , P1_R2278_U8 , P1_R2278_U308 );
and AND3_28528 ( P1_R2278_U10 , P1_R2278_U313 , P1_R2278_U311 , P1_R2278_U315 );
and AND2_28529 ( P1_R2278_U11 , P1_R2278_U134 , P1_R2278_U10 );
and AND2_28530 ( P1_R2278_U12 , P1_R2278_U295 , P1_R2278_U292 );
and AND2_28531 ( P1_R2278_U13 , P1_R2278_U9 , P1_R2278_U321 );
and AND2_28532 ( P1_R2278_U14 , P1_R2278_U463 , P1_R2278_U462 );
and AND2_28533 ( P1_R2278_U15 , P1_R2278_U344 , P1_R2278_U342 );
and AND4_28534 ( P1_R2278_U16 , P1_R2278_U188 , P1_R2278_U375 , P1_R2278_U468 , P1_R2278_U467 );
and AND2_28535 ( P1_R2278_U17 , P1_R2278_U272 , P1_R2278_U270 );
and AND2_28536 ( P1_R2278_U18 , P1_R2278_U268 , P1_R2278_U266 );
nand NAND2_28537 ( P1_R2278_U19 , P1_R2278_U214 , P1_R2278_U429 );
and AND2_28538 ( P1_R2278_U20 , P1_R2278_U414 , P1_R2278_U335 );
not NOT1_28539 ( P1_R2278_U21 , P1_INSTADDRPOINTER_REG_8_ );
not NOT1_28540 ( P1_R2278_U22 , P1_U2792 );
not NOT1_28541 ( P1_R2278_U23 , P1_INSTADDRPOINTER_REG_7_ );
not NOT1_28542 ( P1_R2278_U24 , P1_U2793 );
not NOT1_28543 ( P1_R2278_U25 , P1_INSTADDRPOINTER_REG_6_ );
not NOT1_28544 ( P1_R2278_U26 , P1_U2794 );
not NOT1_28545 ( P1_R2278_U27 , P1_INSTADDRPOINTER_REG_5_ );
not NOT1_28546 ( P1_R2278_U28 , P1_U2795 );
not NOT1_28547 ( P1_R2278_U29 , P1_U2800 );
not NOT1_28548 ( P1_R2278_U30 , P1_INSTADDRPOINTER_REG_0_ );
not NOT1_28549 ( P1_R2278_U31 , P1_INSTADDRPOINTER_REG_1_ );
nand NAND2_28550 ( P1_R2278_U32 , P1_INSTADDRPOINTER_REG_0_ , P1_U2800 );
not NOT1_28551 ( P1_R2278_U33 , P1_U2799 );
not NOT1_28552 ( P1_R2278_U34 , P1_INSTADDRPOINTER_REG_2_ );
not NOT1_28553 ( P1_R2278_U35 , P1_U2798 );
not NOT1_28554 ( P1_R2278_U36 , P1_INSTADDRPOINTER_REG_3_ );
not NOT1_28555 ( P1_R2278_U37 , P1_U2797 );
not NOT1_28556 ( P1_R2278_U38 , P1_INSTADDRPOINTER_REG_4_ );
not NOT1_28557 ( P1_R2278_U39 , P1_U2796 );
nand NAND2_28558 ( P1_R2278_U40 , P1_R2278_U43 , P1_R2278_U250 );
nand NAND3_28559 ( P1_R2278_U41 , P1_R2278_U254 , P1_R2278_U252 , P1_R2278_U253 );
nand NAND2_28560 ( P1_R2278_U42 , P1_R2278_U246 , P1_R2278_U245 );
nand NAND2_28561 ( P1_R2278_U43 , P1_R2278_U42 , P1_R2278_U248 );
not NOT1_28562 ( P1_R2278_U44 , P1_INSTADDRPOINTER_REG_25_ );
not NOT1_28563 ( P1_R2278_U45 , P1_U2775 );
not NOT1_28564 ( P1_R2278_U46 , P1_INSTADDRPOINTER_REG_26_ );
not NOT1_28565 ( P1_R2278_U47 , P1_U2774 );
not NOT1_28566 ( P1_R2278_U48 , P1_INSTADDRPOINTER_REG_24_ );
not NOT1_28567 ( P1_R2278_U49 , P1_U2776 );
not NOT1_28568 ( P1_R2278_U50 , P1_INSTADDRPOINTER_REG_23_ );
not NOT1_28569 ( P1_R2278_U51 , P1_U2777 );
not NOT1_28570 ( P1_R2278_U52 , P1_INSTADDRPOINTER_REG_21_ );
not NOT1_28571 ( P1_R2278_U53 , P1_U2779 );
not NOT1_28572 ( P1_R2278_U54 , P1_INSTADDRPOINTER_REG_20_ );
not NOT1_28573 ( P1_R2278_U55 , P1_U2780 );
not NOT1_28574 ( P1_R2278_U56 , P1_INSTADDRPOINTER_REG_19_ );
not NOT1_28575 ( P1_R2278_U57 , P1_U2781 );
not NOT1_28576 ( P1_R2278_U58 , P1_INSTADDRPOINTER_REG_11_ );
not NOT1_28577 ( P1_R2278_U59 , P1_U2789 );
not NOT1_28578 ( P1_R2278_U60 , P1_INSTADDRPOINTER_REG_10_ );
not NOT1_28579 ( P1_R2278_U61 , P1_U2790 );
not NOT1_28580 ( P1_R2278_U62 , P1_INSTADDRPOINTER_REG_15_ );
not NOT1_28581 ( P1_R2278_U63 , P1_U2785 );
not NOT1_28582 ( P1_R2278_U64 , P1_INSTADDRPOINTER_REG_13_ );
not NOT1_28583 ( P1_R2278_U65 , P1_U2787 );
not NOT1_28584 ( P1_R2278_U66 , P1_INSTADDRPOINTER_REG_14_ );
not NOT1_28585 ( P1_R2278_U67 , P1_U2786 );
nand NAND2_28586 ( P1_R2278_U68 , P1_U2788 , P1_INSTADDRPOINTER_REG_12_ );
not NOT1_28587 ( P1_R2278_U69 , P1_INSTADDRPOINTER_REG_16_ );
not NOT1_28588 ( P1_R2278_U70 , P1_U2784 );
not NOT1_28589 ( P1_R2278_U71 , P1_INSTADDRPOINTER_REG_17_ );
not NOT1_28590 ( P1_R2278_U72 , P1_U2783 );
nand NAND4_28591 ( P1_R2278_U73 , P1_R2278_U12 , P1_R2278_U8 , P1_R2278_U359 , P1_R2278_U308 );
not NOT1_28592 ( P1_R2278_U74 , P1_INSTADDRPOINTER_REG_22_ );
not NOT1_28593 ( P1_R2278_U75 , P1_U2778 );
nand NAND2_28594 ( P1_R2278_U76 , P1_U2778 , P1_INSTADDRPOINTER_REG_22_ );
not NOT1_28595 ( P1_R2278_U77 , P1_INSTADDRPOINTER_REG_18_ );
not NOT1_28596 ( P1_R2278_U78 , P1_U2782 );
nand NAND2_28597 ( P1_R2278_U79 , P1_U2782 , P1_INSTADDRPOINTER_REG_18_ );
nand NAND2_28598 ( P1_R2278_U80 , P1_R2278_U144 , P1_R2278_U8 );
not NOT1_28599 ( P1_R2278_U81 , P1_U2772 );
not NOT1_28600 ( P1_R2278_U82 , P1_INSTADDRPOINTER_REG_28_ );
not NOT1_28601 ( P1_R2278_U83 , P1_INSTADDRPOINTER_REG_27_ );
not NOT1_28602 ( P1_R2278_U84 , P1_U2773 );
nand NAND2_28603 ( P1_R2278_U85 , P1_U2773 , P1_INSTADDRPOINTER_REG_27_ );
nand NAND2_28604 ( P1_R2278_U86 , P1_R2278_U379 , P1_R2278_U322 );
nand NAND3_28605 ( P1_R2278_U87 , P1_R2278_U392 , P1_R2278_U92 , P1_R2278_U93 );
not NOT1_28606 ( P1_R2278_U88 , P1_U2770 );
not NOT1_28607 ( P1_R2278_U89 , P1_INSTADDRPOINTER_REG_30_ );
not NOT1_28608 ( P1_R2278_U90 , P1_U2771 );
not NOT1_28609 ( P1_R2278_U91 , P1_INSTADDRPOINTER_REG_29_ );
nand NAND2_28610 ( P1_R2278_U92 , P1_R2278_U143 , P1_R2278_U11 );
nand NAND3_28611 ( P1_R2278_U93 , P1_R2278_U11 , P1_R2278_U321 , P1_R2278_U377 );
nand NAND2_28612 ( P1_R2278_U94 , P1_R2278_U132 , P1_R2278_U372 );
nand NAND2_28613 ( P1_R2278_U95 , P1_R2278_U136 , P1_R2278_U368 );
nand NAND3_28614 ( P1_R2278_U96 , P1_R2278_U11 , P1_R2278_U321 , P1_R2278_U378 );
nand NAND2_28615 ( P1_R2278_U97 , P1_R2278_U229 , P1_R2278_U331 );
nand NAND2_28616 ( P1_R2278_U98 , P1_R2278_U138 , P1_R2278_U354 );
nand NAND2_28617 ( P1_R2278_U99 , P1_R2278_U610 , P1_R2278_U609 );
and AND2_28618 ( P1_R2278_U100 , P1_R2278_U262 , P1_R2278_U261 );
nand NAND2_28619 ( P1_R2278_U101 , P1_R2278_U431 , P1_R2278_U430 );
nand NAND2_28620 ( P1_R2278_U102 , P1_R2278_U438 , P1_R2278_U437 );
nand NAND2_28621 ( P1_R2278_U103 , P1_R2278_U445 , P1_R2278_U444 );
nand NAND2_28622 ( P1_R2278_U104 , P1_R2278_U454 , P1_R2278_U453 );
nand NAND2_28623 ( P1_R2278_U105 , P1_R2278_U461 , P1_R2278_U460 );
nand NAND2_28624 ( P1_R2278_U106 , P1_R2278_U477 , P1_R2278_U476 );
nand NAND2_28625 ( P1_R2278_U107 , P1_R2278_U484 , P1_R2278_U483 );
nand NAND2_28626 ( P1_R2278_U108 , P1_R2278_U491 , P1_R2278_U490 );
nand NAND2_28627 ( P1_R2278_U109 , P1_R2278_U498 , P1_R2278_U497 );
nand NAND2_28628 ( P1_R2278_U110 , P1_R2278_U505 , P1_R2278_U504 );
nand NAND2_28629 ( P1_R2278_U111 , P1_R2278_U512 , P1_R2278_U511 );
nand NAND2_28630 ( P1_R2278_U112 , P1_R2278_U519 , P1_R2278_U518 );
nand NAND2_28631 ( P1_R2278_U113 , P1_R2278_U526 , P1_R2278_U525 );
nand NAND2_28632 ( P1_R2278_U114 , P1_R2278_U533 , P1_R2278_U532 );
nand NAND2_28633 ( P1_R2278_U115 , P1_R2278_U540 , P1_R2278_U539 );
nand NAND2_28634 ( P1_R2278_U116 , P1_R2278_U547 , P1_R2278_U546 );
nand NAND2_28635 ( P1_R2278_U117 , P1_R2278_U554 , P1_R2278_U553 );
nand NAND2_28636 ( P1_R2278_U118 , P1_R2278_U566 , P1_R2278_U565 );
nand NAND2_28637 ( P1_R2278_U119 , P1_R2278_U573 , P1_R2278_U572 );
nand NAND2_28638 ( P1_R2278_U120 , P1_R2278_U580 , P1_R2278_U579 );
nand NAND2_28639 ( P1_R2278_U121 , P1_R2278_U587 , P1_R2278_U586 );
nand NAND2_28640 ( P1_R2278_U122 , P1_R2278_U594 , P1_R2278_U593 );
nand NAND2_28641 ( P1_R2278_U123 , P1_R2278_U599 , P1_R2278_U598 );
and AND2_28642 ( P1_R2278_U124 , P1_R2278_U68 , P1_R2278_U281 );
nand NAND2_28643 ( P1_R2278_U125 , P1_R2278_U601 , P1_R2278_U600 );
nand NAND2_28644 ( P1_R2278_U126 , P1_R2278_U608 , P1_R2278_U607 );
and AND2_28645 ( P1_R2278_U127 , P1_INSTADDRPOINTER_REG_7_ , P1_U2793 );
and AND2_28646 ( P1_R2278_U128 , P1_R2278_U258 , P1_R2278_U254 );
and AND2_28647 ( P1_R2278_U129 , P1_R2278_U352 , P1_R2278_U259 );
and AND2_28648 ( P1_R2278_U130 , P1_INSTADDRPOINTER_REG_23_ , P1_U2777 );
and AND2_28649 ( P1_R2278_U131 , P1_R2278_U318 , P1_R2278_U316 );
and AND3_28650 ( P1_R2278_U132 , P1_R2278_U319 , P1_R2278_U317 , P1_R2278_U321 );
and AND2_28651 ( P1_R2278_U133 , P1_INSTADDRPOINTER_REG_19_ , P1_U2781 );
and AND2_28652 ( P1_R2278_U134 , P1_R2278_U319 , P1_R2278_U317 );
and AND2_28653 ( P1_R2278_U135 , P1_R2278_U321 , P1_R2278_U308 );
and AND2_28654 ( P1_R2278_U136 , P1_R2278_U11 , P1_R2278_U135 );
and AND3_28655 ( P1_R2278_U137 , P1_R2278_U259 , P1_R2278_U228 , P1_R2278_U273 );
and AND2_28656 ( P1_R2278_U138 , P1_R2278_U389 , P1_R2278_U276 );
and AND2_28657 ( P1_R2278_U139 , P1_R2278_U357 , P1_R2278_U140 );
and AND3_28658 ( P1_R2278_U140 , P1_R2278_U281 , P1_R2278_U283 , P1_R2278_U284 );
and AND2_28659 ( P1_R2278_U141 , P1_R2278_U286 , P1_R2278_U410 );
and AND2_28660 ( P1_R2278_U142 , P1_R2278_U7 , P1_R2278_U13 );
and AND2_28661 ( P1_R2278_U143 , P1_R2278_U309 , P1_R2278_U321 );
and AND2_28662 ( P1_R2278_U144 , P1_R2278_U296 , P1_R2278_U308 );
and AND2_28663 ( P1_R2278_U145 , P1_R2278_U95 , P1_R2278_U94 );
and AND2_28664 ( P1_R2278_U146 , P1_R2278_U401 , P1_R2278_U96 );
and AND2_28665 ( P1_R2278_U147 , P1_R2278_U324 , P1_R2278_U5 );
and AND4_28666 ( P1_R2278_U148 , P1_R2278_U324 , P1_R2278_U321 , P1_R2278_U319 , P1_R2278_U317 );
and AND3_28667 ( P1_R2278_U149 , P1_R2278_U321 , P1_R2278_U308 , P1_R2278_U324 );
and AND2_28668 ( P1_R2278_U150 , P1_R2278_U11 , P1_R2278_U149 );
and AND2_28669 ( P1_R2278_U151 , P1_R2278_U286 , P1_R2278_U412 );
and AND2_28670 ( P1_R2278_U152 , P1_R2278_U11 , P1_R2278_U324 );
and AND2_28671 ( P1_R2278_U153 , P1_R2278_U7 , P1_R2278_U13 );
and AND2_28672 ( P1_R2278_U154 , P1_R2278_U324 , P1_R2278_U321 );
and AND5_28673 ( P1_R2278_U155 , P1_R2278_U394 , P1_R2278_U393 , P1_R2278_U395 , P1_R2278_U398 , P1_R2278_U156 );
and AND3_28674 ( P1_R2278_U156 , P1_R2278_U14 , P1_R2278_U400 , P1_R2278_U399 );
and AND2_28675 ( P1_R2278_U157 , P1_R2278_U11 , P1_R2278_U324 );
and AND2_28676 ( P1_R2278_U158 , P1_R2278_U7 , P1_R2278_U13 );
and AND3_28677 ( P1_R2278_U159 , P1_R2278_U403 , P1_R2278_U187 , P1_R2278_U404 );
and AND2_28678 ( P1_R2278_U160 , P1_R2278_U286 , P1_R2278_U417 );
and AND2_28679 ( P1_R2278_U161 , P1_R2278_U9 , P1_R2278_U7 );
and AND2_28680 ( P1_R2278_U162 , P1_R2278_U369 , P1_R2278_U76 );
and AND2_28681 ( P1_R2278_U163 , P1_R2278_U73 , P1_R2278_U80 );
and AND2_28682 ( P1_R2278_U164 , P1_R2278_U317 , P1_R2278_U10 );
and AND2_28683 ( P1_R2278_U165 , P1_R2278_U371 , P1_R2278_U316 );
and AND2_28684 ( P1_R2278_U166 , P1_R2278_U311 , P1_R2278_U313 );
and AND2_28685 ( P1_R2278_U167 , P1_R2278_U370 , P1_R2278_U314 );
and AND2_28686 ( P1_R2278_U168 , P1_R2278_U286 , P1_R2278_U415 );
and AND2_28687 ( P1_R2278_U169 , P1_R2278_U362 , P1_R2278_U79 );
and AND2_28688 ( P1_R2278_U170 , P1_R2278_U367 , P1_R2278_U306 );
and AND2_28689 ( P1_R2278_U171 , P1_R2278_U298 , P1_R2278_U302 );
and AND2_28690 ( P1_R2278_U172 , P1_R2278_U364 , P1_R2278_U303 );
and AND3_28691 ( P1_R2278_U173 , P1_R2278_U589 , P1_R2278_U588 , P1_R2278_U285 );
and AND2_28692 ( P1_R2278_U174 , P1_R2278_U337 , P1_R2278_U227 );
and AND3_28693 ( P1_R2278_U175 , P1_R2278_U603 , P1_R2278_U602 , P1_R2278_U228 );
nand NAND2_28694 ( P1_R2278_U176 , P1_R2278_U129 , P1_R2278_U353 );
and AND2_28695 ( P1_R2278_U177 , P1_R2278_U433 , P1_R2278_U432 );
nand NAND2_28696 ( P1_R2278_U178 , P1_R2278_U41 , P1_R2278_U256 );
and AND2_28697 ( P1_R2278_U179 , P1_R2278_U440 , P1_R2278_U439 );
and AND2_28698 ( P1_R2278_U180 , P1_R2278_U447 , P1_R2278_U446 );
and AND2_28699 ( P1_R2278_U181 , P1_R2278_U449 , P1_R2278_U448 );
nand NAND2_28700 ( P1_R2278_U182 , P1_R2278_U242 , P1_R2278_U241 );
and AND2_28701 ( P1_R2278_U183 , P1_R2278_U456 , P1_R2278_U455 );
nand NAND2_28702 ( P1_R2278_U184 , P1_R2278_U238 , P1_R2278_U237 );
not NOT1_28703 ( P1_R2278_U185 , P1_INSTADDRPOINTER_REG_31_ );
not NOT1_28704 ( P1_R2278_U186 , P1_U2769 );
nand NAND2_28705 ( P1_R2278_U187 , P1_INSTADDRPOINTER_REG_29_ , P1_U2771 );
and AND2_28706 ( P1_R2278_U188 , P1_R2278_U470 , P1_R2278_U469 );
and AND2_28707 ( P1_R2278_U189 , P1_R2278_U472 , P1_R2278_U471 );
nand NAND4_28708 ( P1_R2278_U190 , P1_R2278_U406 , P1_R2278_U405 , P1_R2278_U407 , P1_R2278_U159 );
and AND2_28709 ( P1_R2278_U191 , P1_R2278_U479 , P1_R2278_U478 );
nand NAND2_28710 ( P1_R2278_U192 , P1_R2278_U213 , P1_R2278_U234 );
and AND2_28711 ( P1_R2278_U193 , P1_R2278_U486 , P1_R2278_U485 );
nand NAND3_28712 ( P1_R2278_U194 , P1_R2278_U145 , P1_R2278_U385 , P1_R2278_U146 );
and AND2_28713 ( P1_R2278_U195 , P1_R2278_U493 , P1_R2278_U492 );
nand NAND2_28714 ( P1_R2278_U196 , P1_R2278_U419 , P1_R2278_U409 );
and AND2_28715 ( P1_R2278_U197 , P1_R2278_U500 , P1_R2278_U499 );
nand NAND2_28716 ( P1_R2278_U198 , P1_R2278_U425 , P1_R2278_U373 );
and AND2_28717 ( P1_R2278_U199 , P1_R2278_U507 , P1_R2278_U506 );
nand NAND2_28718 ( P1_R2278_U200 , P1_R2278_U165 , P1_R2278_U423 );
and AND2_28719 ( P1_R2278_U201 , P1_R2278_U514 , P1_R2278_U513 );
nand NAND2_28720 ( P1_R2278_U202 , P1_R2278_U167 , P1_R2278_U427 );
and AND2_28721 ( P1_R2278_U203 , P1_R2278_U521 , P1_R2278_U520 );
nand NAND2_28722 ( P1_R2278_U204 , P1_R2278_U421 , P1_R2278_U312 );
and AND2_28723 ( P1_R2278_U205 , P1_R2278_U528 , P1_R2278_U527 );
nand NAND3_28724 ( P1_R2278_U206 , P1_R2278_U163 , P1_R2278_U376 , P1_R2278_U162 );
and AND2_28725 ( P1_R2278_U207 , P1_R2278_U535 , P1_R2278_U534 );
nand NAND2_28726 ( P1_R2278_U208 , P1_R2278_U170 , P1_R2278_U365 );
and AND2_28727 ( P1_R2278_U209 , P1_R2278_U542 , P1_R2278_U541 );
nand NAND2_28728 ( P1_R2278_U210 , P1_R2278_U172 , P1_R2278_U363 );
and AND2_28729 ( P1_R2278_U211 , P1_R2278_U549 , P1_R2278_U548 );
nand NAND2_28730 ( P1_R2278_U212 , P1_R2278_U300 , P1_R2278_U299 );
nand NAND2_28731 ( P1_R2278_U213 , P1_U2799 , P1_R2278_U232 );
and AND2_28732 ( P1_R2278_U214 , P1_R2278_U559 , P1_R2278_U558 );
and AND2_28733 ( P1_R2278_U215 , P1_R2278_U561 , P1_R2278_U560 );
nand NAND2_28734 ( P1_R2278_U216 , P1_R2278_U169 , P1_R2278_U361 );
and AND2_28735 ( P1_R2278_U217 , P1_R2278_U568 , P1_R2278_U567 );
nand NAND2_28736 ( P1_R2278_U218 , P1_R2278_U360 , P1_R2278_U358 );
and AND2_28737 ( P1_R2278_U219 , P1_R2278_U575 , P1_R2278_U574 );
nand NAND2_28738 ( P1_R2278_U220 , P1_R2278_U290 , P1_R2278_U289 );
and AND2_28739 ( P1_R2278_U221 , P1_R2278_U582 , P1_R2278_U581 );
nand NAND2_28740 ( P1_R2278_U222 , P1_R2278_U168 , P1_R2278_U226 );
nand NAND2_28741 ( P1_R2278_U223 , P1_R2278_U68 , P1_R2278_U328 );
nand NAND2_28742 ( P1_R2278_U224 , P1_R2278_U98 , P1_R2278_U279 );
nand NAND2_28743 ( P1_R2278_U225 , P1_R2278_U274 , P1_R2278_U273 );
nand NAND2_28744 ( P1_R2278_U226 , P1_R2278_U224 , P1_R2278_U139 );
nand NAND2_28745 ( P1_R2278_U227 , P1_R2278_U356 , P1_R2278_U355 );
nand NAND2_28746 ( P1_R2278_U228 , P1_U2790 , P1_INSTADDRPOINTER_REG_10_ );
nand NAND2_28747 ( P1_R2278_U229 , P1_U2787 , P1_INSTADDRPOINTER_REG_13_ );
not NOT1_28748 ( P1_R2278_U230 , P1_R2278_U213 );
nand NAND2_28749 ( P1_R2278_U231 , P1_U2794 , P1_INSTADDRPOINTER_REG_6_ );
not NOT1_28750 ( P1_R2278_U232 , P1_R2278_U32 );
nand NAND2_28751 ( P1_R2278_U233 , P1_R2278_U33 , P1_R2278_U32 );
nand NAND2_28752 ( P1_R2278_U234 , P1_INSTADDRPOINTER_REG_1_ , P1_R2278_U233 );
not NOT1_28753 ( P1_R2278_U235 , P1_R2278_U192 );
or OR2_28754 ( P1_R2278_U236 , P1_INSTADDRPOINTER_REG_2_ , P1_U2798 );
nand NAND2_28755 ( P1_R2278_U237 , P1_R2278_U236 , P1_R2278_U192 );
nand NAND2_28756 ( P1_R2278_U238 , P1_U2798 , P1_INSTADDRPOINTER_REG_2_ );
not NOT1_28757 ( P1_R2278_U239 , P1_R2278_U184 );
or OR2_28758 ( P1_R2278_U240 , P1_INSTADDRPOINTER_REG_3_ , P1_U2797 );
nand NAND2_28759 ( P1_R2278_U241 , P1_R2278_U240 , P1_R2278_U184 );
nand NAND2_28760 ( P1_R2278_U242 , P1_U2797 , P1_INSTADDRPOINTER_REG_3_ );
not NOT1_28761 ( P1_R2278_U243 , P1_R2278_U182 );
or OR2_28762 ( P1_R2278_U244 , P1_INSTADDRPOINTER_REG_4_ , P1_U2796 );
nand NAND2_28763 ( P1_R2278_U245 , P1_R2278_U244 , P1_R2278_U182 );
nand NAND2_28764 ( P1_R2278_U246 , P1_U2796 , P1_INSTADDRPOINTER_REG_4_ );
not NOT1_28765 ( P1_R2278_U247 , P1_R2278_U42 );
or OR2_28766 ( P1_R2278_U248 , P1_U2795 , P1_INSTADDRPOINTER_REG_5_ );
not NOT1_28767 ( P1_R2278_U249 , P1_R2278_U43 );
nand NAND2_28768 ( P1_R2278_U250 , P1_U2795 , P1_INSTADDRPOINTER_REG_5_ );
not NOT1_28769 ( P1_R2278_U251 , P1_R2278_U40 );
nand NAND2_28770 ( P1_R2278_U252 , P1_R2278_U251 , P1_R2278_U231 );
or OR2_28771 ( P1_R2278_U253 , P1_U2793 , P1_INSTADDRPOINTER_REG_7_ );
or OR2_28772 ( P1_R2278_U254 , P1_U2794 , P1_INSTADDRPOINTER_REG_6_ );
not NOT1_28773 ( P1_R2278_U255 , P1_R2278_U41 );
nand NAND2_28774 ( P1_R2278_U256 , P1_U2793 , P1_INSTADDRPOINTER_REG_7_ );
not NOT1_28775 ( P1_R2278_U257 , P1_R2278_U178 );
or OR2_28776 ( P1_R2278_U258 , P1_INSTADDRPOINTER_REG_8_ , P1_U2792 );
nand NAND2_28777 ( P1_R2278_U259 , P1_U2792 , P1_INSTADDRPOINTER_REG_8_ );
not NOT1_28778 ( P1_R2278_U260 , P1_R2278_U176 );
or OR2_28779 ( P1_R2278_U261 , P1_INSTADDRPOINTER_REG_9_ , P1_U2791 );
nand NAND2_28780 ( P1_R2278_U262 , P1_U2791 , P1_INSTADDRPOINTER_REG_9_ );
nand NAND2_28781 ( P1_R2278_U263 , P1_U2791 , P1_INSTADDRPOINTER_REG_9_ );
or OR2_28782 ( P1_R2278_U264 , P1_INSTADDRPOINTER_REG_6_ , P1_U2794 );
nand NAND2_28783 ( P1_R2278_U265 , P1_R2278_U264 , P1_R2278_U40 );
nand NAND3_28784 ( P1_R2278_U266 , P1_R2278_U265 , P1_R2278_U231 , P1_R2278_U179 );
nand NAND2_28785 ( P1_R2278_U267 , P1_U2793 , P1_INSTADDRPOINTER_REG_7_ );
nand NAND2_28786 ( P1_R2278_U268 , P1_R2278_U255 , P1_R2278_U267 );
or OR2_28787 ( P1_R2278_U269 , P1_U2794 , P1_INSTADDRPOINTER_REG_6_ );
nand NAND2_28788 ( P1_R2278_U270 , P1_R2278_U180 , P1_R2278_U247 );
nand NAND2_28789 ( P1_R2278_U271 , P1_U2795 , P1_INSTADDRPOINTER_REG_5_ );
nand NAND2_28790 ( P1_R2278_U272 , P1_R2278_U249 , P1_R2278_U271 );
nand NAND2_28791 ( P1_R2278_U273 , P1_U2791 , P1_INSTADDRPOINTER_REG_9_ );
nand NAND2_28792 ( P1_R2278_U274 , P1_R2278_U261 , P1_R2278_U176 );
not NOT1_28793 ( P1_R2278_U275 , P1_R2278_U225 );
or OR2_28794 ( P1_R2278_U276 , P1_U2789 , P1_INSTADDRPOINTER_REG_11_ );
or OR2_28795 ( P1_R2278_U277 , P1_U2790 , P1_INSTADDRPOINTER_REG_10_ );
not NOT1_28796 ( P1_R2278_U278 , P1_R2278_U98 );
nand NAND2_28797 ( P1_R2278_U279 , P1_U2789 , P1_INSTADDRPOINTER_REG_11_ );
not NOT1_28798 ( P1_R2278_U280 , P1_R2278_U224 );
or OR2_28799 ( P1_R2278_U281 , P1_INSTADDRPOINTER_REG_12_ , P1_U2788 );
not NOT1_28800 ( P1_R2278_U282 , P1_R2278_U68 );
or OR2_28801 ( P1_R2278_U283 , P1_U2787 , P1_INSTADDRPOINTER_REG_13_ );
or OR2_28802 ( P1_R2278_U284 , P1_U2786 , P1_INSTADDRPOINTER_REG_14_ );
nand NAND2_28803 ( P1_R2278_U285 , P1_U2786 , P1_INSTADDRPOINTER_REG_14_ );
nand NAND2_28804 ( P1_R2278_U286 , P1_U2785 , P1_INSTADDRPOINTER_REG_15_ );
nand NAND3_28805 ( P1_R2278_U287 , P1_R2278_U391 , P1_R2278_U229 , P1_R2278_U285 );
or OR2_28806 ( P1_R2278_U288 , P1_INSTADDRPOINTER_REG_16_ , P1_U2784 );
nand NAND2_28807 ( P1_R2278_U289 , P1_R2278_U288 , P1_R2278_U222 );
nand NAND2_28808 ( P1_R2278_U290 , P1_U2784 , P1_INSTADDRPOINTER_REG_16_ );
not NOT1_28809 ( P1_R2278_U291 , P1_R2278_U220 );
or OR2_28810 ( P1_R2278_U292 , P1_INSTADDRPOINTER_REG_17_ , P1_U2783 );
nand NAND2_28811 ( P1_R2278_U293 , P1_U2783 , P1_INSTADDRPOINTER_REG_17_ );
not NOT1_28812 ( P1_R2278_U294 , P1_R2278_U218 );
or OR2_28813 ( P1_R2278_U295 , P1_INSTADDRPOINTER_REG_18_ , P1_U2782 );
not NOT1_28814 ( P1_R2278_U296 , P1_R2278_U79 );
not NOT1_28815 ( P1_R2278_U297 , P1_R2278_U216 );
or OR2_28816 ( P1_R2278_U298 , P1_INSTADDRPOINTER_REG_19_ , P1_U2781 );
nand NAND2_28817 ( P1_R2278_U299 , P1_R2278_U298 , P1_R2278_U216 );
nand NAND2_28818 ( P1_R2278_U300 , P1_U2781 , P1_INSTADDRPOINTER_REG_19_ );
not NOT1_28819 ( P1_R2278_U301 , P1_R2278_U212 );
or OR2_28820 ( P1_R2278_U302 , P1_INSTADDRPOINTER_REG_20_ , P1_U2780 );
nand NAND2_28821 ( P1_R2278_U303 , P1_U2780 , P1_INSTADDRPOINTER_REG_20_ );
not NOT1_28822 ( P1_R2278_U304 , P1_R2278_U210 );
or OR2_28823 ( P1_R2278_U305 , P1_INSTADDRPOINTER_REG_21_ , P1_U2779 );
nand NAND2_28824 ( P1_R2278_U306 , P1_U2779 , P1_INSTADDRPOINTER_REG_21_ );
not NOT1_28825 ( P1_R2278_U307 , P1_R2278_U208 );
or OR2_28826 ( P1_R2278_U308 , P1_INSTADDRPOINTER_REG_22_ , P1_U2778 );
not NOT1_28827 ( P1_R2278_U309 , P1_R2278_U76 );
not NOT1_28828 ( P1_R2278_U310 , P1_R2278_U206 );
or OR2_28829 ( P1_R2278_U311 , P1_INSTADDRPOINTER_REG_23_ , P1_U2777 );
nand NAND2_28830 ( P1_R2278_U312 , P1_U2777 , P1_INSTADDRPOINTER_REG_23_ );
or OR2_28831 ( P1_R2278_U313 , P1_INSTADDRPOINTER_REG_24_ , P1_U2776 );
nand NAND2_28832 ( P1_R2278_U314 , P1_U2776 , P1_INSTADDRPOINTER_REG_24_ );
or OR2_28833 ( P1_R2278_U315 , P1_INSTADDRPOINTER_REG_25_ , P1_U2775 );
nand NAND2_28834 ( P1_R2278_U316 , P1_U2775 , P1_INSTADDRPOINTER_REG_25_ );
or OR2_28835 ( P1_R2278_U317 , P1_INSTADDRPOINTER_REG_26_ , P1_U2774 );
nand NAND2_28836 ( P1_R2278_U318 , P1_U2774 , P1_INSTADDRPOINTER_REG_26_ );
or OR2_28837 ( P1_R2278_U319 , P1_INSTADDRPOINTER_REG_27_ , P1_U2773 );
not NOT1_28838 ( P1_R2278_U320 , P1_R2278_U85 );
or OR2_28839 ( P1_R2278_U321 , P1_U2772 , P1_INSTADDRPOINTER_REG_28_ );
nand NAND2_28840 ( P1_R2278_U322 , P1_INSTADDRPOINTER_REG_28_ , P1_U2772 );
not NOT1_28841 ( P1_R2278_U323 , P1_R2278_U194 );
or OR2_28842 ( P1_R2278_U324 , P1_U2771 , P1_INSTADDRPOINTER_REG_29_ );
not NOT1_28843 ( P1_R2278_U325 , P1_R2278_U187 );
not NOT1_28844 ( P1_R2278_U326 , P1_R2278_U190 );
or OR2_28845 ( P1_R2278_U327 , P1_INSTADDRPOINTER_REG_30_ , P1_U2770 );
nand NAND2_28846 ( P1_R2278_U328 , P1_R2278_U281 , P1_R2278_U224 );
not NOT1_28847 ( P1_R2278_U329 , P1_R2278_U223 );
or OR2_28848 ( P1_R2278_U330 , P1_INSTADDRPOINTER_REG_13_ , P1_U2787 );
nand NAND2_28849 ( P1_R2278_U331 , P1_R2278_U330 , P1_R2278_U223 );
not NOT1_28850 ( P1_R2278_U332 , P1_R2278_U97 );
or OR2_28851 ( P1_R2278_U333 , P1_INSTADDRPOINTER_REG_14_ , P1_U2786 );
nand NAND2_28852 ( P1_R2278_U334 , P1_R2278_U333 , P1_R2278_U97 );
nand NAND2_28853 ( P1_R2278_U335 , P1_R2278_U173 , P1_R2278_U334 );
nand NAND2_28854 ( P1_R2278_U336 , P1_R2278_U332 , P1_R2278_U285 );
nand NAND2_28855 ( P1_R2278_U337 , P1_U2785 , P1_INSTADDRPOINTER_REG_15_ );
or OR2_28856 ( P1_R2278_U338 , P1_U2786 , P1_INSTADDRPOINTER_REG_14_ );
or OR2_28857 ( P1_R2278_U339 , P1_U2787 , P1_INSTADDRPOINTER_REG_13_ );
or OR2_28858 ( P1_R2278_U340 , P1_INSTADDRPOINTER_REG_10_ , P1_U2790 );
nand NAND2_28859 ( P1_R2278_U341 , P1_R2278_U340 , P1_R2278_U225 );
nand NAND2_28860 ( P1_R2278_U342 , P1_R2278_U175 , P1_R2278_U341 );
nand NAND2_28861 ( P1_R2278_U343 , P1_U2789 , P1_INSTADDRPOINTER_REG_11_ );
nand NAND2_28862 ( P1_R2278_U344 , P1_R2278_U278 , P1_R2278_U343 );
or OR2_28863 ( P1_R2278_U345 , P1_U2790 , P1_INSTADDRPOINTER_REG_10_ );
nand NAND2_28864 ( P1_R2278_U346 , P1_R2278_U263 , P1_R2278_U261 );
nand NAND2_28865 ( P1_R2278_U347 , P1_R2278_U269 , P1_R2278_U231 );
nand NAND2_28866 ( P1_R2278_U348 , P1_R2278_U338 , P1_R2278_U285 );
nand NAND2_28867 ( P1_R2278_U349 , P1_R2278_U339 , P1_R2278_U229 );
nand NAND2_28868 ( P1_R2278_U350 , P1_R2278_U68 , P1_R2278_U281 );
nand NAND2_28869 ( P1_R2278_U351 , P1_R2278_U345 , P1_R2278_U228 );
nand NAND2_28870 ( P1_R2278_U352 , P1_R2278_U127 , P1_R2278_U258 );
nand NAND3_28871 ( P1_R2278_U353 , P1_R2278_U253 , P1_R2278_U252 , P1_R2278_U128 );
nand NAND3_28872 ( P1_R2278_U354 , P1_R2278_U353 , P1_R2278_U352 , P1_R2278_U137 );
nand NAND2_28873 ( P1_R2278_U355 , P1_U2785 , P1_R2278_U284 );
nand NAND2_28874 ( P1_R2278_U356 , P1_INSTADDRPOINTER_REG_15_ , P1_R2278_U284 );
nand NAND2_28875 ( P1_R2278_U357 , P1_R2278_U356 , P1_R2278_U63 );
nand NAND2_28876 ( P1_R2278_U358 , P1_R2278_U6 , P1_R2278_U222 );
nand NAND2_28877 ( P1_R2278_U359 , P1_R2278_U293 , P1_R2278_U290 );
nand NAND2_28878 ( P1_R2278_U360 , P1_R2278_U359 , P1_R2278_U292 );
nand NAND2_28879 ( P1_R2278_U361 , P1_R2278_U7 , P1_R2278_U222 );
nand NAND2_28880 ( P1_R2278_U362 , P1_R2278_U12 , P1_R2278_U359 );
nand NAND2_28881 ( P1_R2278_U363 , P1_R2278_U171 , P1_R2278_U216 );
nand NAND2_28882 ( P1_R2278_U364 , P1_R2278_U133 , P1_R2278_U302 );
nand NAND2_28883 ( P1_R2278_U365 , P1_R2278_U8 , P1_R2278_U216 );
nand NAND2_28884 ( P1_R2278_U366 , P1_R2278_U364 , P1_R2278_U303 );
nand NAND2_28885 ( P1_R2278_U367 , P1_R2278_U366 , P1_R2278_U305 );
nand NAND2_28886 ( P1_R2278_U368 , P1_R2278_U367 , P1_R2278_U306 );
nand NAND2_28887 ( P1_R2278_U369 , P1_R2278_U368 , P1_R2278_U308 );
nand NAND2_28888 ( P1_R2278_U370 , P1_R2278_U130 , P1_R2278_U313 );
nand NAND2_28889 ( P1_R2278_U371 , P1_R2278_U381 , P1_R2278_U315 );
nand NAND2_28890 ( P1_R2278_U372 , P1_R2278_U131 , P1_R2278_U371 );
nand NAND2_28891 ( P1_R2278_U373 , P1_R2278_U372 , P1_R2278_U317 );
nand NAND2_28892 ( P1_R2278_U374 , P1_R2278_U372 , P1_R2278_U317 );
nand NAND2_28893 ( P1_R2278_U375 , P1_R2278_U147 , P1_R2278_U194 );
nand NAND2_28894 ( P1_R2278_U376 , P1_R2278_U161 , P1_R2278_U418 );
not NOT1_28895 ( P1_R2278_U377 , P1_R2278_U80 );
not NOT1_28896 ( P1_R2278_U378 , P1_R2278_U73 );
nand NAND2_28897 ( P1_R2278_U379 , P1_R2278_U320 , P1_R2278_U321 );
not NOT1_28898 ( P1_R2278_U380 , P1_R2278_U94 );
nand NAND2_28899 ( P1_R2278_U381 , P1_R2278_U370 , P1_R2278_U314 );
nand NAND3_28900 ( P1_R2278_U382 , P1_R2278_U391 , P1_R2278_U229 , P1_R2278_U285 );
not NOT1_28901 ( P1_R2278_U383 , P1_R2278_U92 );
not NOT1_28902 ( P1_R2278_U384 , P1_R2278_U95 );
nand NAND3_28903 ( P1_R2278_U385 , P1_R2278_U11 , P1_R2278_U411 , P1_R2278_U142 );
not NOT1_28904 ( P1_R2278_U386 , P1_R2278_U93 );
not NOT1_28905 ( P1_R2278_U387 , P1_R2278_U96 );
nand NAND2_28906 ( P1_R2278_U388 , P1_R2278_U277 , P1_R2278_U261 );
nand NAND2_28907 ( P1_R2278_U389 , P1_R2278_U388 , P1_R2278_U228 );
nand NAND3_28908 ( P1_R2278_U390 , P1_R2278_U391 , P1_R2278_U229 , P1_R2278_U285 );
nand NAND2_28909 ( P1_R2278_U391 , P1_R2278_U282 , P1_R2278_U283 );
not NOT1_28910 ( P1_R2278_U392 , P1_R2278_U86 );
nand NAND2_28911 ( P1_R2278_U393 , P1_INSTADDRPOINTER_REG_30_ , P1_U2770 );
nand NAND2_28912 ( P1_R2278_U394 , P1_R2278_U148 , P1_R2278_U372 );
nand NAND2_28913 ( P1_R2278_U395 , P1_R2278_U383 , P1_R2278_U324 );
nand NAND2_28914 ( P1_R2278_U396 , P1_R2278_U150 , P1_R2278_U368 );
nand NAND3_28915 ( P1_R2278_U397 , P1_R2278_U152 , P1_R2278_U413 , P1_R2278_U153 );
nand NAND2_28916 ( P1_R2278_U398 , P1_R2278_U386 , P1_R2278_U324 );
nand NAND3_28917 ( P1_R2278_U399 , P1_R2278_U154 , P1_R2278_U11 , P1_R2278_U378 );
nand NAND2_28918 ( P1_R2278_U400 , P1_R2278_U86 , P1_R2278_U324 );
not NOT1_28919 ( P1_R2278_U401 , P1_R2278_U87 );
nand NAND3_28920 ( P1_R2278_U402 , P1_R2278_U391 , P1_R2278_U229 , P1_R2278_U285 );
nand NAND2_28921 ( P1_R2278_U403 , P1_R2278_U380 , P1_R2278_U324 );
nand NAND2_28922 ( P1_R2278_U404 , P1_R2278_U384 , P1_R2278_U324 );
nand NAND3_28923 ( P1_R2278_U405 , P1_R2278_U157 , P1_R2278_U411 , P1_R2278_U158 );
nand NAND2_28924 ( P1_R2278_U406 , P1_R2278_U387 , P1_R2278_U324 );
nand NAND2_28925 ( P1_R2278_U407 , P1_R2278_U87 , P1_R2278_U324 );
nand NAND2_28926 ( P1_R2278_U408 , P1_R2278_U374 , P1_R2278_U85 );
nand NAND2_28927 ( P1_R2278_U409 , P1_R2278_U408 , P1_R2278_U319 );
nand NAND2_28928 ( P1_R2278_U410 , P1_R2278_U402 , P1_R2278_U227 );
nand NAND2_28929 ( P1_R2278_U411 , P1_R2278_U141 , P1_R2278_U226 );
nand NAND2_28930 ( P1_R2278_U412 , P1_R2278_U390 , P1_R2278_U227 );
nand NAND2_28931 ( P1_R2278_U413 , P1_R2278_U151 , P1_R2278_U226 );
nand NAND2_28932 ( P1_R2278_U414 , P1_R2278_U174 , P1_R2278_U336 );
nand NAND2_28933 ( P1_R2278_U415 , P1_R2278_U287 , P1_R2278_U227 );
not NOT1_28934 ( P1_R2278_U416 , P1_R2278_U222 );
nand NAND2_28935 ( P1_R2278_U417 , P1_R2278_U382 , P1_R2278_U227 );
nand NAND2_28936 ( P1_R2278_U418 , P1_R2278_U160 , P1_R2278_U226 );
nand NAND2_28937 ( P1_R2278_U419 , P1_R2278_U11 , P1_R2278_U206 );
not NOT1_28938 ( P1_R2278_U420 , P1_R2278_U196 );
nand NAND2_28939 ( P1_R2278_U421 , P1_R2278_U311 , P1_R2278_U206 );
not NOT1_28940 ( P1_R2278_U422 , P1_R2278_U204 );
nand NAND2_28941 ( P1_R2278_U423 , P1_R2278_U10 , P1_R2278_U206 );
not NOT1_28942 ( P1_R2278_U424 , P1_R2278_U200 );
nand NAND2_28943 ( P1_R2278_U425 , P1_R2278_U164 , P1_R2278_U206 );
not NOT1_28944 ( P1_R2278_U426 , P1_R2278_U198 );
nand NAND2_28945 ( P1_R2278_U427 , P1_R2278_U166 , P1_R2278_U206 );
not NOT1_28946 ( P1_R2278_U428 , P1_R2278_U202 );
nand NAND2_28947 ( P1_R2278_U429 , P1_R2278_U557 , P1_R2278_U33 );
nand NAND2_28948 ( P1_R2278_U430 , P1_R2278_U346 , P1_R2278_U176 );
nand NAND2_28949 ( P1_R2278_U431 , P1_R2278_U100 , P1_R2278_U260 );
nand NAND2_28950 ( P1_R2278_U432 , P1_U2792 , P1_R2278_U21 );
nand NAND2_28951 ( P1_R2278_U433 , P1_INSTADDRPOINTER_REG_8_ , P1_R2278_U22 );
nand NAND2_28952 ( P1_R2278_U434 , P1_U2792 , P1_R2278_U21 );
nand NAND2_28953 ( P1_R2278_U435 , P1_INSTADDRPOINTER_REG_8_ , P1_R2278_U22 );
nand NAND2_28954 ( P1_R2278_U436 , P1_R2278_U435 , P1_R2278_U434 );
nand NAND2_28955 ( P1_R2278_U437 , P1_R2278_U177 , P1_R2278_U178 );
nand NAND2_28956 ( P1_R2278_U438 , P1_R2278_U257 , P1_R2278_U436 );
nand NAND2_28957 ( P1_R2278_U439 , P1_U2793 , P1_R2278_U23 );
nand NAND2_28958 ( P1_R2278_U440 , P1_INSTADDRPOINTER_REG_7_ , P1_R2278_U24 );
nand NAND2_28959 ( P1_R2278_U441 , P1_U2794 , P1_R2278_U25 );
nand NAND2_28960 ( P1_R2278_U442 , P1_INSTADDRPOINTER_REG_6_ , P1_R2278_U26 );
nand NAND2_28961 ( P1_R2278_U443 , P1_R2278_U442 , P1_R2278_U441 );
nand NAND2_28962 ( P1_R2278_U444 , P1_R2278_U347 , P1_R2278_U40 );
nand NAND2_28963 ( P1_R2278_U445 , P1_R2278_U443 , P1_R2278_U251 );
nand NAND2_28964 ( P1_R2278_U446 , P1_U2795 , P1_R2278_U27 );
nand NAND2_28965 ( P1_R2278_U447 , P1_INSTADDRPOINTER_REG_5_ , P1_R2278_U28 );
nand NAND2_28966 ( P1_R2278_U448 , P1_U2796 , P1_R2278_U38 );
nand NAND2_28967 ( P1_R2278_U449 , P1_INSTADDRPOINTER_REG_4_ , P1_R2278_U39 );
nand NAND2_28968 ( P1_R2278_U450 , P1_U2796 , P1_R2278_U38 );
nand NAND2_28969 ( P1_R2278_U451 , P1_INSTADDRPOINTER_REG_4_ , P1_R2278_U39 );
nand NAND2_28970 ( P1_R2278_U452 , P1_R2278_U451 , P1_R2278_U450 );
nand NAND2_28971 ( P1_R2278_U453 , P1_R2278_U181 , P1_R2278_U182 );
nand NAND2_28972 ( P1_R2278_U454 , P1_R2278_U243 , P1_R2278_U452 );
nand NAND2_28973 ( P1_R2278_U455 , P1_U2797 , P1_R2278_U36 );
nand NAND2_28974 ( P1_R2278_U456 , P1_INSTADDRPOINTER_REG_3_ , P1_R2278_U37 );
nand NAND2_28975 ( P1_R2278_U457 , P1_U2797 , P1_R2278_U36 );
nand NAND2_28976 ( P1_R2278_U458 , P1_INSTADDRPOINTER_REG_3_ , P1_R2278_U37 );
nand NAND2_28977 ( P1_R2278_U459 , P1_R2278_U458 , P1_R2278_U457 );
nand NAND2_28978 ( P1_R2278_U460 , P1_R2278_U183 , P1_R2278_U184 );
nand NAND2_28979 ( P1_R2278_U461 , P1_R2278_U239 , P1_R2278_U459 );
nand NAND2_28980 ( P1_R2278_U462 , P1_INSTADDRPOINTER_REG_31_ , P1_R2278_U186 );
nand NAND2_28981 ( P1_R2278_U463 , P1_U2769 , P1_R2278_U185 );
nand NAND2_28982 ( P1_R2278_U464 , P1_INSTADDRPOINTER_REG_31_ , P1_R2278_U186 );
nand NAND2_28983 ( P1_R2278_U465 , P1_U2769 , P1_R2278_U185 );
nand NAND2_28984 ( P1_R2278_U466 , P1_R2278_U465 , P1_R2278_U464 );
nand NAND4_28985 ( P1_R2278_U467 , P1_R2278_U397 , P1_R2278_U396 , P1_R2278_U155 , P1_R2278_U187 );
nand NAND2_28986 ( P1_R2278_U468 , P1_R2278_U325 , P1_R2278_U5 );
nand NAND3_28987 ( P1_R2278_U469 , P1_R2278_U14 , P1_R2278_U88 , P1_R2278_U89 );
nand NAND3_28988 ( P1_R2278_U470 , P1_U2770 , P1_R2278_U466 , P1_INSTADDRPOINTER_REG_30_ );
nand NAND2_28989 ( P1_R2278_U471 , P1_INSTADDRPOINTER_REG_30_ , P1_R2278_U88 );
nand NAND2_28990 ( P1_R2278_U472 , P1_U2770 , P1_R2278_U89 );
nand NAND2_28991 ( P1_R2278_U473 , P1_INSTADDRPOINTER_REG_30_ , P1_R2278_U88 );
nand NAND2_28992 ( P1_R2278_U474 , P1_U2770 , P1_R2278_U89 );
nand NAND2_28993 ( P1_R2278_U475 , P1_R2278_U474 , P1_R2278_U473 );
nand NAND2_28994 ( P1_R2278_U476 , P1_R2278_U189 , P1_R2278_U190 );
nand NAND2_28995 ( P1_R2278_U477 , P1_R2278_U326 , P1_R2278_U475 );
nand NAND2_28996 ( P1_R2278_U478 , P1_U2798 , P1_R2278_U34 );
nand NAND2_28997 ( P1_R2278_U479 , P1_INSTADDRPOINTER_REG_2_ , P1_R2278_U35 );
nand NAND2_28998 ( P1_R2278_U480 , P1_U2798 , P1_R2278_U34 );
nand NAND2_28999 ( P1_R2278_U481 , P1_INSTADDRPOINTER_REG_2_ , P1_R2278_U35 );
nand NAND2_29000 ( P1_R2278_U482 , P1_R2278_U481 , P1_R2278_U480 );
nand NAND2_29001 ( P1_R2278_U483 , P1_R2278_U191 , P1_R2278_U192 );
nand NAND2_29002 ( P1_R2278_U484 , P1_R2278_U235 , P1_R2278_U482 );
nand NAND2_29003 ( P1_R2278_U485 , P1_INSTADDRPOINTER_REG_29_ , P1_R2278_U90 );
nand NAND2_29004 ( P1_R2278_U486 , P1_U2771 , P1_R2278_U91 );
nand NAND2_29005 ( P1_R2278_U487 , P1_INSTADDRPOINTER_REG_29_ , P1_R2278_U90 );
nand NAND2_29006 ( P1_R2278_U488 , P1_U2771 , P1_R2278_U91 );
nand NAND2_29007 ( P1_R2278_U489 , P1_R2278_U488 , P1_R2278_U487 );
nand NAND2_29008 ( P1_R2278_U490 , P1_R2278_U193 , P1_R2278_U194 );
nand NAND2_29009 ( P1_R2278_U491 , P1_R2278_U323 , P1_R2278_U489 );
nand NAND2_29010 ( P1_R2278_U492 , P1_INSTADDRPOINTER_REG_28_ , P1_R2278_U81 );
nand NAND2_29011 ( P1_R2278_U493 , P1_U2772 , P1_R2278_U82 );
nand NAND2_29012 ( P1_R2278_U494 , P1_INSTADDRPOINTER_REG_28_ , P1_R2278_U81 );
nand NAND2_29013 ( P1_R2278_U495 , P1_U2772 , P1_R2278_U82 );
nand NAND2_29014 ( P1_R2278_U496 , P1_R2278_U495 , P1_R2278_U494 );
nand NAND2_29015 ( P1_R2278_U497 , P1_R2278_U195 , P1_R2278_U196 );
nand NAND2_29016 ( P1_R2278_U498 , P1_R2278_U420 , P1_R2278_U496 );
nand NAND2_29017 ( P1_R2278_U499 , P1_U2773 , P1_R2278_U83 );
nand NAND2_29018 ( P1_R2278_U500 , P1_INSTADDRPOINTER_REG_27_ , P1_R2278_U84 );
nand NAND2_29019 ( P1_R2278_U501 , P1_U2773 , P1_R2278_U83 );
nand NAND2_29020 ( P1_R2278_U502 , P1_INSTADDRPOINTER_REG_27_ , P1_R2278_U84 );
nand NAND2_29021 ( P1_R2278_U503 , P1_R2278_U502 , P1_R2278_U501 );
nand NAND2_29022 ( P1_R2278_U504 , P1_R2278_U197 , P1_R2278_U198 );
nand NAND2_29023 ( P1_R2278_U505 , P1_R2278_U426 , P1_R2278_U503 );
nand NAND2_29024 ( P1_R2278_U506 , P1_U2774 , P1_R2278_U46 );
nand NAND2_29025 ( P1_R2278_U507 , P1_INSTADDRPOINTER_REG_26_ , P1_R2278_U47 );
nand NAND2_29026 ( P1_R2278_U508 , P1_U2774 , P1_R2278_U46 );
nand NAND2_29027 ( P1_R2278_U509 , P1_INSTADDRPOINTER_REG_26_ , P1_R2278_U47 );
nand NAND2_29028 ( P1_R2278_U510 , P1_R2278_U509 , P1_R2278_U508 );
nand NAND2_29029 ( P1_R2278_U511 , P1_R2278_U199 , P1_R2278_U200 );
nand NAND2_29030 ( P1_R2278_U512 , P1_R2278_U424 , P1_R2278_U510 );
nand NAND2_29031 ( P1_R2278_U513 , P1_U2775 , P1_R2278_U44 );
nand NAND2_29032 ( P1_R2278_U514 , P1_INSTADDRPOINTER_REG_25_ , P1_R2278_U45 );
nand NAND2_29033 ( P1_R2278_U515 , P1_U2775 , P1_R2278_U44 );
nand NAND2_29034 ( P1_R2278_U516 , P1_INSTADDRPOINTER_REG_25_ , P1_R2278_U45 );
nand NAND2_29035 ( P1_R2278_U517 , P1_R2278_U516 , P1_R2278_U515 );
nand NAND2_29036 ( P1_R2278_U518 , P1_R2278_U201 , P1_R2278_U202 );
nand NAND2_29037 ( P1_R2278_U519 , P1_R2278_U428 , P1_R2278_U517 );
nand NAND2_29038 ( P1_R2278_U520 , P1_U2776 , P1_R2278_U48 );
nand NAND2_29039 ( P1_R2278_U521 , P1_INSTADDRPOINTER_REG_24_ , P1_R2278_U49 );
nand NAND2_29040 ( P1_R2278_U522 , P1_U2776 , P1_R2278_U48 );
nand NAND2_29041 ( P1_R2278_U523 , P1_INSTADDRPOINTER_REG_24_ , P1_R2278_U49 );
nand NAND2_29042 ( P1_R2278_U524 , P1_R2278_U523 , P1_R2278_U522 );
nand NAND2_29043 ( P1_R2278_U525 , P1_R2278_U203 , P1_R2278_U204 );
nand NAND2_29044 ( P1_R2278_U526 , P1_R2278_U422 , P1_R2278_U524 );
nand NAND2_29045 ( P1_R2278_U527 , P1_U2777 , P1_R2278_U50 );
nand NAND2_29046 ( P1_R2278_U528 , P1_INSTADDRPOINTER_REG_23_ , P1_R2278_U51 );
nand NAND2_29047 ( P1_R2278_U529 , P1_U2777 , P1_R2278_U50 );
nand NAND2_29048 ( P1_R2278_U530 , P1_INSTADDRPOINTER_REG_23_ , P1_R2278_U51 );
nand NAND2_29049 ( P1_R2278_U531 , P1_R2278_U530 , P1_R2278_U529 );
nand NAND2_29050 ( P1_R2278_U532 , P1_R2278_U205 , P1_R2278_U206 );
nand NAND2_29051 ( P1_R2278_U533 , P1_R2278_U310 , P1_R2278_U531 );
nand NAND2_29052 ( P1_R2278_U534 , P1_U2778 , P1_R2278_U74 );
nand NAND2_29053 ( P1_R2278_U535 , P1_INSTADDRPOINTER_REG_22_ , P1_R2278_U75 );
nand NAND2_29054 ( P1_R2278_U536 , P1_U2778 , P1_R2278_U74 );
nand NAND2_29055 ( P1_R2278_U537 , P1_INSTADDRPOINTER_REG_22_ , P1_R2278_U75 );
nand NAND2_29056 ( P1_R2278_U538 , P1_R2278_U537 , P1_R2278_U536 );
nand NAND2_29057 ( P1_R2278_U539 , P1_R2278_U207 , P1_R2278_U208 );
nand NAND2_29058 ( P1_R2278_U540 , P1_R2278_U307 , P1_R2278_U538 );
nand NAND2_29059 ( P1_R2278_U541 , P1_U2779 , P1_R2278_U52 );
nand NAND2_29060 ( P1_R2278_U542 , P1_INSTADDRPOINTER_REG_21_ , P1_R2278_U53 );
nand NAND2_29061 ( P1_R2278_U543 , P1_U2779 , P1_R2278_U52 );
nand NAND2_29062 ( P1_R2278_U544 , P1_INSTADDRPOINTER_REG_21_ , P1_R2278_U53 );
nand NAND2_29063 ( P1_R2278_U545 , P1_R2278_U544 , P1_R2278_U543 );
nand NAND2_29064 ( P1_R2278_U546 , P1_R2278_U209 , P1_R2278_U210 );
nand NAND2_29065 ( P1_R2278_U547 , P1_R2278_U304 , P1_R2278_U545 );
nand NAND2_29066 ( P1_R2278_U548 , P1_U2780 , P1_R2278_U54 );
nand NAND2_29067 ( P1_R2278_U549 , P1_INSTADDRPOINTER_REG_20_ , P1_R2278_U55 );
nand NAND2_29068 ( P1_R2278_U550 , P1_U2780 , P1_R2278_U54 );
nand NAND2_29069 ( P1_R2278_U551 , P1_INSTADDRPOINTER_REG_20_ , P1_R2278_U55 );
nand NAND2_29070 ( P1_R2278_U552 , P1_R2278_U551 , P1_R2278_U550 );
nand NAND2_29071 ( P1_R2278_U553 , P1_R2278_U211 , P1_R2278_U212 );
nand NAND2_29072 ( P1_R2278_U554 , P1_R2278_U301 , P1_R2278_U552 );
nand NAND2_29073 ( P1_R2278_U555 , P1_INSTADDRPOINTER_REG_1_ , P1_R2278_U32 );
nand NAND2_29074 ( P1_R2278_U556 , P1_R2278_U232 , P1_R2278_U31 );
nand NAND2_29075 ( P1_R2278_U557 , P1_R2278_U556 , P1_R2278_U555 );
nand NAND3_29076 ( P1_R2278_U558 , P1_U2799 , P1_R2278_U32 , P1_R2278_U31 );
nand NAND2_29077 ( P1_R2278_U559 , P1_R2278_U230 , P1_INSTADDRPOINTER_REG_1_ );
nand NAND2_29078 ( P1_R2278_U560 , P1_U2781 , P1_R2278_U56 );
nand NAND2_29079 ( P1_R2278_U561 , P1_INSTADDRPOINTER_REG_19_ , P1_R2278_U57 );
nand NAND2_29080 ( P1_R2278_U562 , P1_U2781 , P1_R2278_U56 );
nand NAND2_29081 ( P1_R2278_U563 , P1_INSTADDRPOINTER_REG_19_ , P1_R2278_U57 );
nand NAND2_29082 ( P1_R2278_U564 , P1_R2278_U563 , P1_R2278_U562 );
nand NAND2_29083 ( P1_R2278_U565 , P1_R2278_U215 , P1_R2278_U216 );
nand NAND2_29084 ( P1_R2278_U566 , P1_R2278_U297 , P1_R2278_U564 );
nand NAND2_29085 ( P1_R2278_U567 , P1_U2782 , P1_R2278_U77 );
nand NAND2_29086 ( P1_R2278_U568 , P1_INSTADDRPOINTER_REG_18_ , P1_R2278_U78 );
nand NAND2_29087 ( P1_R2278_U569 , P1_U2782 , P1_R2278_U77 );
nand NAND2_29088 ( P1_R2278_U570 , P1_INSTADDRPOINTER_REG_18_ , P1_R2278_U78 );
nand NAND2_29089 ( P1_R2278_U571 , P1_R2278_U570 , P1_R2278_U569 );
nand NAND2_29090 ( P1_R2278_U572 , P1_R2278_U217 , P1_R2278_U218 );
nand NAND2_29091 ( P1_R2278_U573 , P1_R2278_U294 , P1_R2278_U571 );
nand NAND2_29092 ( P1_R2278_U574 , P1_U2783 , P1_R2278_U71 );
nand NAND2_29093 ( P1_R2278_U575 , P1_INSTADDRPOINTER_REG_17_ , P1_R2278_U72 );
nand NAND2_29094 ( P1_R2278_U576 , P1_U2783 , P1_R2278_U71 );
nand NAND2_29095 ( P1_R2278_U577 , P1_INSTADDRPOINTER_REG_17_ , P1_R2278_U72 );
nand NAND2_29096 ( P1_R2278_U578 , P1_R2278_U577 , P1_R2278_U576 );
nand NAND2_29097 ( P1_R2278_U579 , P1_R2278_U219 , P1_R2278_U220 );
nand NAND2_29098 ( P1_R2278_U580 , P1_R2278_U291 , P1_R2278_U578 );
nand NAND2_29099 ( P1_R2278_U581 , P1_U2784 , P1_R2278_U69 );
nand NAND2_29100 ( P1_R2278_U582 , P1_INSTADDRPOINTER_REG_16_ , P1_R2278_U70 );
nand NAND2_29101 ( P1_R2278_U583 , P1_U2784 , P1_R2278_U69 );
nand NAND2_29102 ( P1_R2278_U584 , P1_INSTADDRPOINTER_REG_16_ , P1_R2278_U70 );
nand NAND2_29103 ( P1_R2278_U585 , P1_R2278_U584 , P1_R2278_U583 );
nand NAND2_29104 ( P1_R2278_U586 , P1_R2278_U221 , P1_R2278_U222 );
nand NAND2_29105 ( P1_R2278_U587 , P1_R2278_U416 , P1_R2278_U585 );
nand NAND2_29106 ( P1_R2278_U588 , P1_U2785 , P1_R2278_U62 );
nand NAND2_29107 ( P1_R2278_U589 , P1_INSTADDRPOINTER_REG_15_ , P1_R2278_U63 );
nand NAND2_29108 ( P1_R2278_U590 , P1_U2786 , P1_R2278_U66 );
nand NAND2_29109 ( P1_R2278_U591 , P1_INSTADDRPOINTER_REG_14_ , P1_R2278_U67 );
nand NAND2_29110 ( P1_R2278_U592 , P1_R2278_U591 , P1_R2278_U590 );
nand NAND2_29111 ( P1_R2278_U593 , P1_R2278_U348 , P1_R2278_U97 );
nand NAND2_29112 ( P1_R2278_U594 , P1_R2278_U592 , P1_R2278_U332 );
nand NAND2_29113 ( P1_R2278_U595 , P1_U2787 , P1_R2278_U64 );
nand NAND2_29114 ( P1_R2278_U596 , P1_INSTADDRPOINTER_REG_13_ , P1_R2278_U65 );
nand NAND2_29115 ( P1_R2278_U597 , P1_R2278_U596 , P1_R2278_U595 );
nand NAND2_29116 ( P1_R2278_U598 , P1_R2278_U349 , P1_R2278_U223 );
nand NAND2_29117 ( P1_R2278_U599 , P1_R2278_U329 , P1_R2278_U597 );
nand NAND2_29118 ( P1_R2278_U600 , P1_R2278_U350 , P1_R2278_U224 );
nand NAND2_29119 ( P1_R2278_U601 , P1_R2278_U124 , P1_R2278_U280 );
nand NAND2_29120 ( P1_R2278_U602 , P1_U2789 , P1_R2278_U58 );
nand NAND2_29121 ( P1_R2278_U603 , P1_INSTADDRPOINTER_REG_11_ , P1_R2278_U59 );
nand NAND2_29122 ( P1_R2278_U604 , P1_U2790 , P1_R2278_U60 );
nand NAND2_29123 ( P1_R2278_U605 , P1_INSTADDRPOINTER_REG_10_ , P1_R2278_U61 );
nand NAND2_29124 ( P1_R2278_U606 , P1_R2278_U605 , P1_R2278_U604 );
nand NAND2_29125 ( P1_R2278_U607 , P1_R2278_U351 , P1_R2278_U225 );
nand NAND2_29126 ( P1_R2278_U608 , P1_R2278_U275 , P1_R2278_U606 );
nand NAND2_29127 ( P1_R2278_U609 , P1_INSTADDRPOINTER_REG_0_ , P1_R2278_U29 );
nand NAND2_29128 ( P1_R2278_U610 , P1_U2800 , P1_R2278_U30 );
and AND2_29129 ( P1_R2358_U5 , P1_R2358_U274 , P1_R2358_U272 );
and AND2_29130 ( P1_R2358_U6 , P1_R2358_U280 , P1_R2358_U278 );
and AND2_29131 ( P1_R2358_U7 , P1_R2358_U6 , P1_R2358_U282 );
and AND2_29132 ( P1_R2358_U8 , P1_R2358_U288 , P1_R2358_U286 );
and AND2_29133 ( P1_R2358_U9 , P1_R2358_U8 , P1_R2358_U290 );
and AND2_29134 ( P1_R2358_U10 , P1_R2358_U9 , P1_R2358_U292 );
and AND2_29135 ( P1_R2358_U11 , P1_R2358_U458 , P1_R2358_U457 );
and AND2_29136 ( P1_R2358_U12 , P1_R2358_U481 , P1_R2358_U480 );
and AND2_29137 ( P1_R2358_U13 , P1_R2358_U555 , P1_R2358_U554 );
and AND2_29138 ( P1_R2358_U14 , P1_R2358_U330 , P1_R2358_U329 );
and AND2_29139 ( P1_R2358_U15 , P1_R2358_U327 , P1_R2358_U325 );
and AND2_29140 ( P1_R2358_U16 , P1_R2358_U320 , P1_R2358_U319 );
and AND2_29141 ( P1_R2358_U17 , P1_R2358_U317 , P1_R2358_U315 );
and AND2_29142 ( P1_R2358_U18 , P1_R2358_U308 , P1_R2358_U307 );
and AND2_29143 ( P1_R2358_U19 , P1_R2358_U254 , P1_R2358_U252 );
and AND2_29144 ( P1_R2358_U20 , P1_R2358_U245 , P1_R2358_U244 );
and AND2_29145 ( P1_R2358_U21 , P1_R2358_U242 , P1_R2358_U240 );
and AND3_29146 ( P1_R2358_U22 , P1_R2358_U566 , P1_R2358_U565 , P1_R2358_U136 );
not NOT1_29147 ( P1_R2358_U23 , P1_U2352 );
not NOT1_29148 ( P1_R2358_U24 , P1_U2643 );
not NOT1_29149 ( P1_R2358_U25 , P1_U2644 );
not NOT1_29150 ( P1_R2358_U26 , P1_U2645 );
not NOT1_29151 ( P1_R2358_U27 , P1_U2646 );
nand NAND2_29152 ( P1_R2358_U28 , P1_U2646 , P1_R2358_U413 );
not NOT1_29153 ( P1_R2358_U29 , P1_U2649 );
not NOT1_29154 ( P1_R2358_U30 , P1_U2648 );
not NOT1_29155 ( P1_R2358_U31 , P1_U2650 );
not NOT1_29156 ( P1_R2358_U32 , P1_U2647 );
not NOT1_29157 ( P1_R2358_U33 , P1_U2642 );
not NOT1_29158 ( P1_R2358_U34 , P1_U2641 );
nand NAND2_29159 ( P1_R2358_U35 , P1_R2358_U236 , P1_R2358_U220 );
nand NAND2_29160 ( P1_R2358_U36 , P1_R2358_U35 , P1_R2358_U218 );
not NOT1_29161 ( P1_R2358_U37 , P1_U2623 );
not NOT1_29162 ( P1_R2358_U38 , P1_U2624 );
not NOT1_29163 ( P1_R2358_U39 , P1_U2625 );
not NOT1_29164 ( P1_R2358_U40 , P1_U2626 );
not NOT1_29165 ( P1_R2358_U41 , P1_U2627 );
nand NAND2_29166 ( P1_R2358_U42 , P1_U2627 , P1_R2358_U546 );
not NOT1_29167 ( P1_R2358_U43 , P1_U2628 );
not NOT1_29168 ( P1_R2358_U44 , P1_U2629 );
not NOT1_29169 ( P1_R2358_U45 , P1_U2630 );
not NOT1_29170 ( P1_R2358_U46 , P1_U2631 );
nand NAND2_29171 ( P1_R2358_U47 , P1_U2631 , P1_R2358_U521 );
not NOT1_29172 ( P1_R2358_U48 , P1_U2632 );
not NOT1_29173 ( P1_R2358_U49 , P1_U2633 );
not NOT1_29174 ( P1_R2358_U50 , P1_U2634 );
nand NAND2_29175 ( P1_R2358_U51 , P1_U2634 , P1_R2358_U501 );
not NOT1_29176 ( P1_R2358_U52 , P1_U2639 );
not NOT1_29177 ( P1_R2358_U53 , P1_U2640 );
nand NAND3_29178 ( P1_R2358_U54 , P1_R2358_U400 , P1_R2358_U399 , P1_R2358_U34 );
not NOT1_29179 ( P1_R2358_U55 , P1_U2635 );
not NOT1_29180 ( P1_R2358_U56 , P1_U2638 );
nand NAND2_29181 ( P1_R2358_U57 , P1_U2638 , P1_R2358_U471 );
not NOT1_29182 ( P1_R2358_U58 , P1_U2637 );
nand NAND2_29183 ( P1_R2358_U59 , P1_U2637 , P1_R2358_U463 );
not NOT1_29184 ( P1_R2358_U60 , P1_U2636 );
nand NAND2_29185 ( P1_R2358_U61 , P1_U2636 , P1_R2358_U466 );
not NOT1_29186 ( P1_R2358_U62 , P1_U2622 );
not NOT1_29187 ( P1_R2358_U63 , P1_U2620 );
not NOT1_29188 ( P1_R2358_U64 , P1_U2621 );
nand NAND2_29189 ( P1_R2358_U65 , P1_R2358_U206 , P1_R2358_U248 );
nand NAND2_29190 ( P1_R2358_U66 , P1_R2358_U65 , P1_R2358_U202 );
nand NAND2_29191 ( P1_R2358_U67 , P1_R2358_U371 , P1_R2358_U293 );
nand NAND2_29192 ( P1_R2358_U68 , P1_R2358_U369 , P1_R2358_U291 );
nand NAND2_29193 ( P1_R2358_U69 , P1_R2358_U364 , P1_R2358_U283 );
nand NAND2_29194 ( P1_R2358_U70 , P1_R2358_U358 , P1_R2358_U275 );
nand NAND2_29195 ( P1_R2358_U71 , P1_R2358_U59 , P1_R2358_U311 );
nand NAND2_29196 ( P1_R2358_U72 , P1_R2358_U71 , P1_R2358_U255 );
nand NAND2_29197 ( P1_R2358_U73 , P1_R2358_U233 , P1_R2358_U321 );
nand NAND2_29198 ( P1_R2358_U74 , P1_R2358_U73 , P1_R2358_U262 );
nand NAND2_29199 ( P1_R2358_U75 , P1_R2358_U557 , P1_R2358_U556 );
nand NAND2_29200 ( P1_R2358_U76 , P1_R2358_U611 , P1_R2358_U610 );
and AND2_29201 ( P1_R2358_U77 , P1_R2358_U233 , P1_R2358_U54 );
nand NAND2_29202 ( P1_R2358_U78 , P1_R2358_U450 , P1_R2358_U449 );
and AND2_29203 ( P1_R2358_U79 , P1_R2358_U229 , P1_R2358_U228 );
nand NAND2_29204 ( P1_R2358_U80 , P1_R2358_U452 , P1_R2358_U451 );
and AND2_29205 ( P1_R2358_U81 , P1_R2358_U220 , P1_R2358_U219 );
nand NAND2_29206 ( P1_R2358_U82 , P1_R2358_U454 , P1_R2358_U453 );
and AND2_29207 ( P1_R2358_U83 , P1_R2358_U225 , P1_R2358_U28 );
nand NAND2_29208 ( P1_R2358_U84 , P1_R2358_U456 , P1_R2358_U455 );
nand NAND2_29209 ( P1_R2358_U85 , P1_R2358_U575 , P1_R2358_U574 );
and AND2_29210 ( P1_R2358_U86 , P1_R2358_U179 , P1_R2358_U300 );
nand NAND2_29211 ( P1_R2358_U87 , P1_R2358_U577 , P1_R2358_U576 );
and AND2_29212 ( P1_R2358_U88 , P1_R2358_U297 , P1_R2358_U296 );
nand NAND2_29213 ( P1_R2358_U89 , P1_R2358_U579 , P1_R2358_U578 );
and AND2_29214 ( P1_R2358_U90 , P1_R2358_U295 , P1_R2358_U294 );
nand NAND2_29215 ( P1_R2358_U91 , P1_R2358_U581 , P1_R2358_U580 );
and AND2_29216 ( P1_R2358_U92 , P1_R2358_U293 , P1_R2358_U292 );
nand NAND2_29217 ( P1_R2358_U93 , P1_R2358_U583 , P1_R2358_U582 );
and AND2_29218 ( P1_R2358_U94 , P1_R2358_U291 , P1_R2358_U290 );
nand NAND2_29219 ( P1_R2358_U95 , P1_R2358_U585 , P1_R2358_U584 );
and AND2_29220 ( P1_R2358_U96 , P1_R2358_U289 , P1_R2358_U288 );
nand NAND2_29221 ( P1_R2358_U97 , P1_R2358_U587 , P1_R2358_U586 );
and AND2_29222 ( P1_R2358_U98 , P1_R2358_U42 , P1_R2358_U286 );
nand NAND2_29223 ( P1_R2358_U99 , P1_R2358_U589 , P1_R2358_U588 );
and AND2_29224 ( P1_R2358_U100 , P1_R2358_U285 , P1_R2358_U284 );
nand NAND2_29225 ( P1_R2358_U101 , P1_R2358_U591 , P1_R2358_U590 );
and AND2_29226 ( P1_R2358_U102 , P1_R2358_U283 , P1_R2358_U282 );
nand NAND2_29227 ( P1_R2358_U103 , P1_R2358_U593 , P1_R2358_U592 );
and AND2_29228 ( P1_R2358_U104 , P1_R2358_U281 , P1_R2358_U280 );
nand NAND2_29229 ( P1_R2358_U105 , P1_R2358_U595 , P1_R2358_U594 );
and AND2_29230 ( P1_R2358_U106 , P1_R2358_U206 , P1_R2358_U205 );
nand NAND2_29231 ( P1_R2358_U107 , P1_R2358_U597 , P1_R2358_U596 );
and AND2_29232 ( P1_R2358_U108 , P1_R2358_U47 , P1_R2358_U278 );
nand NAND2_29233 ( P1_R2358_U109 , P1_R2358_U599 , P1_R2358_U598 );
and AND2_29234 ( P1_R2358_U110 , P1_R2358_U277 , P1_R2358_U276 );
nand NAND2_29235 ( P1_R2358_U111 , P1_R2358_U601 , P1_R2358_U600 );
and AND2_29236 ( P1_R2358_U112 , P1_R2358_U275 , P1_R2358_U274 );
nand NAND2_29237 ( P1_R2358_U113 , P1_R2358_U603 , P1_R2358_U602 );
and AND2_29238 ( P1_R2358_U114 , P1_R2358_U51 , P1_R2358_U272 );
nand NAND2_29239 ( P1_R2358_U115 , P1_R2358_U605 , P1_R2358_U604 );
and AND2_29240 ( P1_R2358_U116 , P1_R2358_U59 , P1_R2358_U258 );
nand NAND2_29241 ( P1_R2358_U117 , P1_R2358_U607 , P1_R2358_U606 );
and AND2_29242 ( P1_R2358_U118 , P1_R2358_U57 , P1_R2358_U259 );
nand NAND2_29243 ( P1_R2358_U119 , P1_R2358_U609 , P1_R2358_U608 );
and AND2_29244 ( P1_R2358_U120 , P1_R2358_U208 , P1_R2358_U205 );
and AND2_29245 ( P1_R2358_U121 , P1_R2358_U204 , P1_R2358_U202 );
and AND2_29246 ( P1_R2358_U122 , P1_R2358_U217 , P1_R2358_U216 );
and AND2_29247 ( P1_R2358_U123 , P1_R2358_U204 , P1_R2358_U203 );
and AND2_29248 ( P1_R2358_U124 , P1_R2358_U229 , P1_R2358_U54 );
and AND2_29249 ( P1_R2358_U125 , P1_R2358_U265 , P1_R2358_U262 );
and AND4_29250 ( P1_R2358_U126 , P1_R2358_U258 , P1_R2358_U259 , P1_R2358_U255 , P1_R2358_U356 );
and AND4_29251 ( P1_R2358_U127 , P1_R2358_U256 , P1_R2358_U353 , P1_R2358_U355 , P1_R2358_U354 );
and AND2_29252 ( P1_R2358_U128 , P1_R2358_U276 , P1_R2358_U5 );
and AND2_29253 ( P1_R2358_U129 , P1_R2358_U361 , P1_R2358_U277 );
and AND2_29254 ( P1_R2358_U130 , P1_R2358_U7 , P1_R2358_U284 );
and AND2_29255 ( P1_R2358_U131 , P1_R2358_U366 , P1_R2358_U285 );
and AND2_29256 ( P1_R2358_U132 , P1_R2358_U10 , P1_R2358_U294 );
and AND2_29257 ( P1_R2358_U133 , P1_R2358_U373 , P1_R2358_U295 );
and AND2_29258 ( P1_R2358_U134 , P1_R2358_U561 , P1_R2358_U305 );
and AND2_29259 ( P1_R2358_U135 , P1_R2358_U304 , P1_R2358_U13 );
and AND2_29260 ( P1_R2358_U136 , P1_R2358_U180 , P1_R2358_U374 );
and AND2_29261 ( P1_R2358_U137 , P1_R2358_U367 , P1_R2358_U289 );
and AND2_29262 ( P1_R2358_U138 , P1_R2358_U362 , P1_R2358_U281 );
and AND2_29263 ( P1_R2358_U139 , P1_R2358_U257 , P1_R2358_U256 );
and AND2_29264 ( P1_R2358_U140 , P1_R2358_U316 , P1_R2358_U61 );
and AND2_29265 ( P1_R2358_U141 , P1_R2358_U265 , P1_R2358_U264 );
and AND2_29266 ( P1_R2358_U142 , P1_R2358_U326 , P1_R2358_U263 );
not NOT1_29267 ( P1_R2358_U143 , P1_U2618 );
not NOT1_29268 ( P1_R2358_U144 , P1_U2615 );
not NOT1_29269 ( P1_R2358_U145 , P1_U2614 );
not NOT1_29270 ( P1_R2358_U146 , P1_U2667 );
not NOT1_29271 ( P1_R2358_U147 , P1_U2668 );
not NOT1_29272 ( P1_R2358_U148 , P1_U2670 );
not NOT1_29273 ( P1_R2358_U149 , P1_U2671 );
not NOT1_29274 ( P1_R2358_U150 , P1_U2672 );
not NOT1_29275 ( P1_R2358_U151 , P1_U2669 );
not NOT1_29276 ( P1_R2358_U152 , P1_U2617 );
nand NAND2_29277 ( P1_R2358_U153 , P1_R2358_U228 , P1_R2358_U230 );
nand NAND3_29278 ( P1_R2358_U154 , P1_R2358_U226 , P1_R2358_U216 , P1_R2358_U224 );
nand NAND2_29279 ( P1_R2358_U155 , P1_R2358_U28 , P1_R2358_U234 );
nand NAND2_29280 ( P1_R2358_U156 , P1_R2358_U203 , P1_R2358_U213 );
not NOT1_29281 ( P1_R2358_U157 , P1_U2611 );
not NOT1_29282 ( P1_R2358_U158 , P1_U2612 );
not NOT1_29283 ( P1_R2358_U159 , P1_U2613 );
not NOT1_29284 ( P1_R2358_U160 , P1_U2616 );
not NOT1_29285 ( P1_R2358_U161 , P1_U2610 );
not NOT1_29286 ( P1_R2358_U162 , P1_U2609 );
not NOT1_29287 ( P1_R2358_U163 , P1_U2666 );
not NOT1_29288 ( P1_R2358_U164 , P1_U2665 );
not NOT1_29289 ( P1_R2358_U165 , P1_U2664 );
not NOT1_29290 ( P1_R2358_U166 , P1_U2660 );
not NOT1_29291 ( P1_R2358_U167 , P1_U2661 );
not NOT1_29292 ( P1_R2358_U168 , P1_U2663 );
not NOT1_29293 ( P1_R2358_U169 , P1_U2662 );
not NOT1_29294 ( P1_R2358_U170 , P1_U2655 );
not NOT1_29295 ( P1_R2358_U171 , P1_U2656 );
not NOT1_29296 ( P1_R2358_U172 , P1_U2657 );
not NOT1_29297 ( P1_R2358_U173 , P1_U2659 );
not NOT1_29298 ( P1_R2358_U174 , P1_U2658 );
not NOT1_29299 ( P1_R2358_U175 , P1_U2654 );
not NOT1_29300 ( P1_R2358_U176 , P1_U2653 );
not NOT1_29301 ( P1_R2358_U177 , P1_U2651 );
not NOT1_29302 ( P1_R2358_U178 , P1_U2652 );
nand NAND2_29303 ( P1_R2358_U179 , P1_U2621 , P1_R2358_U564 );
and AND2_29304 ( P1_R2358_U180 , P1_R2358_U568 , P1_R2358_U567 );
and AND2_29305 ( P1_R2358_U181 , P1_R2358_U570 , P1_R2358_U569 );
nand NAND2_29306 ( P1_R2358_U182 , P1_R2358_U179 , P1_R2358_U302 );
nand NAND2_29307 ( P1_R2358_U183 , P1_R2358_U297 , P1_R2358_U298 );
nand NAND2_29308 ( P1_R2358_U184 , P1_R2358_U133 , P1_R2358_U383 );
nand NAND2_29309 ( P1_R2358_U185 , P1_R2358_U372 , P1_R2358_U381 );
nand NAND2_29310 ( P1_R2358_U186 , P1_R2358_U370 , P1_R2358_U379 );
nand NAND2_29311 ( P1_R2358_U187 , P1_R2358_U137 , P1_R2358_U377 );
nand NAND2_29312 ( P1_R2358_U188 , P1_R2358_U375 , P1_R2358_U42 );
nand NAND2_29313 ( P1_R2358_U189 , P1_R2358_U131 , P1_R2358_U385 );
nand NAND2_29314 ( P1_R2358_U190 , P1_R2358_U365 , P1_R2358_U387 );
nand NAND2_29315 ( P1_R2358_U191 , P1_R2358_U138 , P1_R2358_U389 );
nand NAND2_29316 ( P1_R2358_U192 , P1_R2358_U391 , P1_R2358_U47 );
nand NAND2_29317 ( P1_R2358_U193 , P1_R2358_U209 , P1_R2358_U246 );
nand NAND2_29318 ( P1_R2358_U194 , P1_R2358_U129 , P1_R2358_U393 );
nand NAND2_29319 ( P1_R2358_U195 , P1_R2358_U359 , P1_R2358_U395 );
nand NAND2_29320 ( P1_R2358_U196 , P1_R2358_U397 , P1_R2358_U51 );
nand NAND2_29321 ( P1_R2358_U197 , P1_R2358_U201 , P1_R2358_U127 );
nand NAND2_29322 ( P1_R2358_U198 , P1_R2358_U57 , P1_R2358_U309 );
nand NAND3_29323 ( P1_R2358_U199 , P1_R2358_U268 , P1_R2358_U264 , P1_R2358_U267 );
nand NAND2_29324 ( P1_R2358_U200 , P1_R2358_U209 , P1_R2358_U208 );
nand NAND2_29325 ( P1_R2358_U201 , P1_R2358_U126 , P1_R2358_U199 );
nand NAND3_29326 ( P1_R2358_U202 , P1_R2358_U436 , P1_R2358_U435 , P1_R2358_U30 );
nand NAND2_29327 ( P1_R2358_U203 , P1_U2647 , P1_R2358_U441 );
nand NAND3_29328 ( P1_R2358_U204 , P1_R2358_U438 , P1_R2358_U437 , P1_R2358_U32 );
nand NAND3_29329 ( P1_R2358_U205 , P1_R2358_U432 , P1_R2358_U431 , P1_R2358_U29 );
nand NAND2_29330 ( P1_R2358_U206 , P1_U2649 , P1_R2358_U427 );
nand NAND2_29331 ( P1_R2358_U207 , P1_U2648 , P1_R2358_U424 );
nand NAND3_29332 ( P1_R2358_U208 , P1_R2358_U434 , P1_R2358_U433 , P1_R2358_U31 );
nand NAND2_29333 ( P1_R2358_U209 , P1_U2650 , P1_R2358_U430 );
nand NAND2_29334 ( P1_R2358_U210 , P1_R2358_U209 , P1_R2358_U23 );
nand NAND2_29335 ( P1_R2358_U211 , P1_R2358_U120 , P1_R2358_U210 );
nand NAND3_29336 ( P1_R2358_U212 , P1_R2358_U211 , P1_R2358_U206 , P1_R2358_U207 );
nand NAND2_29337 ( P1_R2358_U213 , P1_R2358_U121 , P1_R2358_U212 );
not NOT1_29338 ( P1_R2358_U214 , P1_R2358_U156 );
nand NAND2_29339 ( P1_R2358_U215 , P1_U2644 , P1_R2358_U408 );
nand NAND2_29340 ( P1_R2358_U216 , P1_U2643 , P1_R2358_U421 );
nand NAND3_29341 ( P1_R2358_U217 , P1_R2358_U405 , P1_R2358_U404 , P1_R2358_U24 );
nand NAND3_29342 ( P1_R2358_U218 , P1_R2358_U418 , P1_R2358_U417 , P1_R2358_U25 );
nand NAND3_29343 ( P1_R2358_U219 , P1_R2358_U410 , P1_R2358_U409 , P1_R2358_U26 );
nand NAND2_29344 ( P1_R2358_U220 , P1_U2645 , P1_R2358_U416 );
not NOT1_29345 ( P1_R2358_U221 , P1_R2358_U28 );
nand NAND2_29346 ( P1_R2358_U222 , P1_R2358_U221 , P1_R2358_U219 );
nand NAND3_29347 ( P1_R2358_U223 , P1_R2358_U220 , P1_R2358_U222 , P1_R2358_U215 );
nand NAND3_29348 ( P1_R2358_U224 , P1_R2358_U218 , P1_R2358_U223 , P1_R2358_U217 );
nand NAND3_29349 ( P1_R2358_U225 , P1_R2358_U443 , P1_R2358_U442 , P1_R2358_U27 );
nand NAND5_29350 ( P1_R2358_U226 , P1_R2358_U225 , P1_R2358_U156 , P1_R2358_U219 , P1_R2358_U218 , P1_R2358_U217 );
not NOT1_29351 ( P1_R2358_U227 , P1_R2358_U154 );
nand NAND2_29352 ( P1_R2358_U228 , P1_U2642 , P1_R2358_U448 );
nand NAND3_29353 ( P1_R2358_U229 , P1_R2358_U445 , P1_R2358_U444 , P1_R2358_U33 );
nand NAND2_29354 ( P1_R2358_U230 , P1_R2358_U229 , P1_R2358_U154 );
not NOT1_29355 ( P1_R2358_U231 , P1_R2358_U153 );
not NOT1_29356 ( P1_R2358_U232 , P1_R2358_U54 );
nand NAND2_29357 ( P1_R2358_U233 , P1_U2641 , P1_R2358_U403 );
nand NAND2_29358 ( P1_R2358_U234 , P1_R2358_U225 , P1_R2358_U156 );
not NOT1_29359 ( P1_R2358_U235 , P1_R2358_U155 );
nand NAND2_29360 ( P1_R2358_U236 , P1_R2358_U155 , P1_R2358_U219 );
not NOT1_29361 ( P1_R2358_U237 , P1_R2358_U35 );
not NOT1_29362 ( P1_R2358_U238 , P1_R2358_U36 );
nand NAND2_29363 ( P1_R2358_U239 , P1_R2358_U36 , P1_R2358_U215 );
nand NAND2_29364 ( P1_R2358_U240 , P1_R2358_U122 , P1_R2358_U239 );
nand NAND2_29365 ( P1_R2358_U241 , P1_R2358_U217 , P1_R2358_U216 );
nand NAND3_29366 ( P1_R2358_U242 , P1_R2358_U36 , P1_R2358_U215 , P1_R2358_U241 );
nand NAND2_29367 ( P1_R2358_U243 , P1_R2358_U218 , P1_R2358_U215 );
nand NAND2_29368 ( P1_R2358_U244 , P1_R2358_U237 , P1_R2358_U243 );
nand NAND2_29369 ( P1_R2358_U245 , P1_R2358_U238 , P1_R2358_U215 );
nand NAND2_29370 ( P1_R2358_U246 , P1_U2352 , P1_R2358_U208 );
not NOT1_29371 ( P1_R2358_U247 , P1_R2358_U193 );
nand NAND2_29372 ( P1_R2358_U248 , P1_R2358_U193 , P1_R2358_U205 );
not NOT1_29373 ( P1_R2358_U249 , P1_R2358_U65 );
not NOT1_29374 ( P1_R2358_U250 , P1_R2358_U66 );
nand NAND2_29375 ( P1_R2358_U251 , P1_R2358_U66 , P1_R2358_U207 );
nand NAND2_29376 ( P1_R2358_U252 , P1_R2358_U123 , P1_R2358_U251 );
nand NAND2_29377 ( P1_R2358_U253 , P1_R2358_U204 , P1_R2358_U203 );
nand NAND3_29378 ( P1_R2358_U254 , P1_R2358_U66 , P1_R2358_U207 , P1_R2358_U253 );
nand NAND3_29379 ( P1_R2358_U255 , P1_R2358_U460 , P1_R2358_U459 , P1_R2358_U60 );
nand NAND2_29380 ( P1_R2358_U256 , P1_U2635 , P1_R2358_U474 );
nand NAND2_29381 ( P1_R2358_U257 , P1_R2358_U11 , P1_R2358_U55 );
nand NAND3_29382 ( P1_R2358_U258 , P1_R2358_U468 , P1_R2358_U467 , P1_R2358_U58 );
nand NAND3_29383 ( P1_R2358_U259 , P1_R2358_U486 , P1_R2358_U485 , P1_R2358_U56 );
not NOT1_29384 ( P1_R2358_U260 , P1_R2358_U59 );
not NOT1_29385 ( P1_R2358_U261 , P1_R2358_U61 );
nand NAND3_29386 ( P1_R2358_U262 , P1_R2358_U476 , P1_R2358_U475 , P1_R2358_U53 );
nand NAND2_29387 ( P1_R2358_U263 , P1_U2640 , P1_R2358_U479 );
nand NAND2_29388 ( P1_R2358_U264 , P1_U2639 , P1_R2358_U484 );
nand NAND2_29389 ( P1_R2358_U265 , P1_R2358_U12 , P1_R2358_U52 );
nand NAND3_29390 ( P1_R2358_U266 , P1_R2358_U233 , P1_R2358_U228 , P1_R2358_U263 );
nand NAND4_29391 ( P1_R2358_U267 , P1_R2358_U360 , P1_R2358_U357 , P1_R2358_U266 , P1_R2358_U262 );
nand NAND3_29392 ( P1_R2358_U268 , P1_R2358_U124 , P1_R2358_U154 , P1_R2358_U125 );
not NOT1_29393 ( P1_R2358_U269 , P1_R2358_U199 );
not NOT1_29394 ( P1_R2358_U270 , P1_R2358_U57 );
not NOT1_29395 ( P1_R2358_U271 , P1_R2358_U197 );
nand NAND3_29396 ( P1_R2358_U272 , P1_R2358_U488 , P1_R2358_U487 , P1_R2358_U50 );
not NOT1_29397 ( P1_R2358_U273 , P1_R2358_U51 );
nand NAND3_29398 ( P1_R2358_U274 , P1_R2358_U490 , P1_R2358_U489 , P1_R2358_U49 );
nand NAND2_29399 ( P1_R2358_U275 , P1_U2633 , P1_R2358_U498 );
nand NAND3_29400 ( P1_R2358_U276 , P1_R2358_U492 , P1_R2358_U491 , P1_R2358_U48 );
nand NAND2_29401 ( P1_R2358_U277 , P1_U2632 , P1_R2358_U495 );
nand NAND3_29402 ( P1_R2358_U278 , P1_R2358_U507 , P1_R2358_U506 , P1_R2358_U46 );
not NOT1_29403 ( P1_R2358_U279 , P1_R2358_U47 );
nand NAND3_29404 ( P1_R2358_U280 , P1_R2358_U509 , P1_R2358_U508 , P1_R2358_U45 );
nand NAND2_29405 ( P1_R2358_U281 , P1_U2630 , P1_R2358_U518 );
nand NAND3_29406 ( P1_R2358_U282 , P1_R2358_U505 , P1_R2358_U504 , P1_R2358_U44 );
nand NAND2_29407 ( P1_R2358_U283 , P1_U2629 , P1_R2358_U515 );
nand NAND3_29408 ( P1_R2358_U284 , P1_R2358_U503 , P1_R2358_U502 , P1_R2358_U43 );
nand NAND2_29409 ( P1_R2358_U285 , P1_U2628 , P1_R2358_U512 );
nand NAND3_29410 ( P1_R2358_U286 , P1_R2358_U529 , P1_R2358_U528 , P1_R2358_U41 );
not NOT1_29411 ( P1_R2358_U287 , P1_R2358_U42 );
nand NAND3_29412 ( P1_R2358_U288 , P1_R2358_U531 , P1_R2358_U530 , P1_R2358_U40 );
nand NAND2_29413 ( P1_R2358_U289 , P1_U2626 , P1_R2358_U543 );
nand NAND3_29414 ( P1_R2358_U290 , P1_R2358_U527 , P1_R2358_U526 , P1_R2358_U39 );
nand NAND2_29415 ( P1_R2358_U291 , P1_U2625 , P1_R2358_U540 );
nand NAND3_29416 ( P1_R2358_U292 , P1_R2358_U525 , P1_R2358_U524 , P1_R2358_U38 );
nand NAND2_29417 ( P1_R2358_U293 , P1_U2624 , P1_R2358_U537 );
nand NAND3_29418 ( P1_R2358_U294 , P1_R2358_U523 , P1_R2358_U522 , P1_R2358_U37 );
nand NAND2_29419 ( P1_R2358_U295 , P1_U2623 , P1_R2358_U534 );
nand NAND3_29420 ( P1_R2358_U296 , P1_R2358_U548 , P1_R2358_U547 , P1_R2358_U62 );
nand NAND2_29421 ( P1_R2358_U297 , P1_U2622 , P1_R2358_U551 );
nand NAND2_29422 ( P1_R2358_U298 , P1_R2358_U296 , P1_R2358_U184 );
not NOT1_29423 ( P1_R2358_U299 , P1_R2358_U183 );
nand NAND3_29424 ( P1_R2358_U300 , P1_R2358_U553 , P1_R2358_U552 , P1_R2358_U64 );
not NOT1_29425 ( P1_R2358_U301 , P1_R2358_U179 );
nand NAND2_29426 ( P1_R2358_U302 , P1_R2358_U300 , P1_R2358_U183 );
not NOT1_29427 ( P1_R2358_U303 , P1_R2358_U182 );
nand NAND2_29428 ( P1_R2358_U304 , P1_U2620 , P1_R2358_U75 );
nand NAND2_29429 ( P1_R2358_U305 , P1_R2358_U558 , P1_R2358_U63 );
nand NAND2_29430 ( P1_R2358_U306 , P1_R2358_U207 , P1_R2358_U202 );
nand NAND2_29431 ( P1_R2358_U307 , P1_R2358_U249 , P1_R2358_U306 );
nand NAND2_29432 ( P1_R2358_U308 , P1_R2358_U250 , P1_R2358_U207 );
nand NAND2_29433 ( P1_R2358_U309 , P1_R2358_U199 , P1_R2358_U259 );
not NOT1_29434 ( P1_R2358_U310 , P1_R2358_U198 );
nand NAND2_29435 ( P1_R2358_U311 , P1_R2358_U198 , P1_R2358_U258 );
not NOT1_29436 ( P1_R2358_U312 , P1_R2358_U71 );
not NOT1_29437 ( P1_R2358_U313 , P1_R2358_U72 );
nand NAND2_29438 ( P1_R2358_U314 , P1_R2358_U72 , P1_R2358_U61 );
nand NAND2_29439 ( P1_R2358_U315 , P1_R2358_U139 , P1_R2358_U314 );
nand NAND2_29440 ( P1_R2358_U316 , P1_R2358_U257 , P1_R2358_U256 );
nand NAND2_29441 ( P1_R2358_U317 , P1_R2358_U140 , P1_R2358_U72 );
nand NAND2_29442 ( P1_R2358_U318 , P1_R2358_U61 , P1_R2358_U255 );
nand NAND2_29443 ( P1_R2358_U319 , P1_R2358_U312 , P1_R2358_U318 );
nand NAND2_29444 ( P1_R2358_U320 , P1_R2358_U313 , P1_R2358_U61 );
nand NAND2_29445 ( P1_R2358_U321 , P1_R2358_U54 , P1_R2358_U153 );
not NOT1_29446 ( P1_R2358_U322 , P1_R2358_U73 );
not NOT1_29447 ( P1_R2358_U323 , P1_R2358_U74 );
nand NAND2_29448 ( P1_R2358_U324 , P1_R2358_U74 , P1_R2358_U263 );
nand NAND2_29449 ( P1_R2358_U325 , P1_R2358_U141 , P1_R2358_U324 );
nand NAND2_29450 ( P1_R2358_U326 , P1_R2358_U265 , P1_R2358_U264 );
nand NAND2_29451 ( P1_R2358_U327 , P1_R2358_U142 , P1_R2358_U74 );
nand NAND2_29452 ( P1_R2358_U328 , P1_R2358_U263 , P1_R2358_U262 );
nand NAND2_29453 ( P1_R2358_U329 , P1_R2358_U322 , P1_R2358_U328 );
nand NAND2_29454 ( P1_R2358_U330 , P1_R2358_U323 , P1_R2358_U263 );
not NOT1_29455 ( P1_R2358_U331 , P1_R2358_U200 );
nand NAND2_29456 ( P1_R2358_U332 , P1_R2358_U233 , P1_R2358_U54 );
nand NAND2_29457 ( P1_R2358_U333 , P1_R2358_U229 , P1_R2358_U228 );
nand NAND2_29458 ( P1_R2358_U334 , P1_R2358_U220 , P1_R2358_U219 );
nand NAND2_29459 ( P1_R2358_U335 , P1_R2358_U225 , P1_R2358_U28 );
nand NAND2_29460 ( P1_R2358_U336 , P1_R2358_U179 , P1_R2358_U300 );
nand NAND2_29461 ( P1_R2358_U337 , P1_R2358_U297 , P1_R2358_U296 );
nand NAND2_29462 ( P1_R2358_U338 , P1_R2358_U295 , P1_R2358_U294 );
nand NAND2_29463 ( P1_R2358_U339 , P1_R2358_U293 , P1_R2358_U292 );
nand NAND2_29464 ( P1_R2358_U340 , P1_R2358_U291 , P1_R2358_U290 );
nand NAND2_29465 ( P1_R2358_U341 , P1_R2358_U289 , P1_R2358_U288 );
nand NAND2_29466 ( P1_R2358_U342 , P1_R2358_U42 , P1_R2358_U286 );
nand NAND2_29467 ( P1_R2358_U343 , P1_R2358_U285 , P1_R2358_U284 );
nand NAND2_29468 ( P1_R2358_U344 , P1_R2358_U283 , P1_R2358_U282 );
nand NAND2_29469 ( P1_R2358_U345 , P1_R2358_U281 , P1_R2358_U280 );
nand NAND2_29470 ( P1_R2358_U346 , P1_R2358_U206 , P1_R2358_U205 );
nand NAND2_29471 ( P1_R2358_U347 , P1_R2358_U47 , P1_R2358_U278 );
nand NAND2_29472 ( P1_R2358_U348 , P1_R2358_U277 , P1_R2358_U276 );
nand NAND2_29473 ( P1_R2358_U349 , P1_R2358_U275 , P1_R2358_U274 );
nand NAND2_29474 ( P1_R2358_U350 , P1_R2358_U51 , P1_R2358_U272 );
nand NAND2_29475 ( P1_R2358_U351 , P1_R2358_U59 , P1_R2358_U258 );
nand NAND2_29476 ( P1_R2358_U352 , P1_R2358_U57 , P1_R2358_U259 );
nand NAND4_29477 ( P1_R2358_U353 , P1_R2358_U270 , P1_R2358_U258 , P1_R2358_U255 , P1_R2358_U257 );
nand NAND3_29478 ( P1_R2358_U354 , P1_R2358_U260 , P1_R2358_U255 , P1_R2358_U257 );
nand NAND2_29479 ( P1_R2358_U355 , P1_R2358_U261 , P1_R2358_U257 );
nand NAND2_29480 ( P1_R2358_U356 , P1_R2358_U11 , P1_R2358_U55 );
nand NAND2_29481 ( P1_R2358_U357 , P1_R2358_U232 , P1_R2358_U263 );
nand NAND2_29482 ( P1_R2358_U358 , P1_R2358_U273 , P1_R2358_U274 );
not NOT1_29483 ( P1_R2358_U359 , P1_R2358_U70 );
nand NAND2_29484 ( P1_R2358_U360 , P1_R2358_U12 , P1_R2358_U52 );
nand NAND2_29485 ( P1_R2358_U361 , P1_R2358_U70 , P1_R2358_U276 );
nand NAND2_29486 ( P1_R2358_U362 , P1_R2358_U279 , P1_R2358_U280 );
nand NAND2_29487 ( P1_R2358_U363 , P1_R2358_U362 , P1_R2358_U281 );
nand NAND2_29488 ( P1_R2358_U364 , P1_R2358_U363 , P1_R2358_U282 );
not NOT1_29489 ( P1_R2358_U365 , P1_R2358_U69 );
nand NAND2_29490 ( P1_R2358_U366 , P1_R2358_U69 , P1_R2358_U284 );
nand NAND2_29491 ( P1_R2358_U367 , P1_R2358_U287 , P1_R2358_U288 );
nand NAND2_29492 ( P1_R2358_U368 , P1_R2358_U367 , P1_R2358_U289 );
nand NAND2_29493 ( P1_R2358_U369 , P1_R2358_U368 , P1_R2358_U290 );
not NOT1_29494 ( P1_R2358_U370 , P1_R2358_U68 );
nand NAND2_29495 ( P1_R2358_U371 , P1_R2358_U68 , P1_R2358_U292 );
not NOT1_29496 ( P1_R2358_U372 , P1_R2358_U67 );
nand NAND2_29497 ( P1_R2358_U373 , P1_R2358_U67 , P1_R2358_U294 );
nand NAND3_29498 ( P1_R2358_U374 , P1_R2358_U300 , P1_R2358_U183 , P1_R2358_U134 );
nand NAND2_29499 ( P1_R2358_U375 , P1_R2358_U286 , P1_R2358_U189 );
not NOT1_29500 ( P1_R2358_U376 , P1_R2358_U188 );
nand NAND2_29501 ( P1_R2358_U377 , P1_R2358_U8 , P1_R2358_U189 );
not NOT1_29502 ( P1_R2358_U378 , P1_R2358_U187 );
nand NAND2_29503 ( P1_R2358_U379 , P1_R2358_U9 , P1_R2358_U189 );
not NOT1_29504 ( P1_R2358_U380 , P1_R2358_U186 );
nand NAND2_29505 ( P1_R2358_U381 , P1_R2358_U10 , P1_R2358_U189 );
not NOT1_29506 ( P1_R2358_U382 , P1_R2358_U185 );
nand NAND2_29507 ( P1_R2358_U383 , P1_R2358_U132 , P1_R2358_U189 );
not NOT1_29508 ( P1_R2358_U384 , P1_R2358_U184 );
nand NAND2_29509 ( P1_R2358_U385 , P1_R2358_U130 , P1_R2358_U194 );
not NOT1_29510 ( P1_R2358_U386 , P1_R2358_U189 );
nand NAND2_29511 ( P1_R2358_U387 , P1_R2358_U7 , P1_R2358_U194 );
not NOT1_29512 ( P1_R2358_U388 , P1_R2358_U190 );
nand NAND2_29513 ( P1_R2358_U389 , P1_R2358_U6 , P1_R2358_U194 );
not NOT1_29514 ( P1_R2358_U390 , P1_R2358_U191 );
nand NAND2_29515 ( P1_R2358_U391 , P1_R2358_U278 , P1_R2358_U194 );
not NOT1_29516 ( P1_R2358_U392 , P1_R2358_U192 );
nand NAND2_29517 ( P1_R2358_U393 , P1_R2358_U128 , P1_R2358_U197 );
not NOT1_29518 ( P1_R2358_U394 , P1_R2358_U194 );
nand NAND2_29519 ( P1_R2358_U395 , P1_R2358_U5 , P1_R2358_U197 );
not NOT1_29520 ( P1_R2358_U396 , P1_R2358_U195 );
nand NAND2_29521 ( P1_R2358_U397 , P1_R2358_U272 , P1_R2358_U197 );
not NOT1_29522 ( P1_R2358_U398 , P1_R2358_U196 );
nand NAND2_29523 ( P1_R2358_U399 , P1_U2352 , P1_R2358_U143 );
nand NAND2_29524 ( P1_R2358_U400 , P1_U2618 , P1_R2358_U23 );
nand NAND2_29525 ( P1_R2358_U401 , P1_U2352 , P1_R2358_U143 );
nand NAND2_29526 ( P1_R2358_U402 , P1_U2618 , P1_R2358_U23 );
nand NAND2_29527 ( P1_R2358_U403 , P1_R2358_U402 , P1_R2358_U401 );
nand NAND2_29528 ( P1_R2358_U404 , P1_U2352 , P1_R2358_U144 );
nand NAND2_29529 ( P1_R2358_U405 , P1_U2615 , P1_R2358_U23 );
nand NAND2_29530 ( P1_R2358_U406 , P1_U2352 , P1_R2358_U145 );
nand NAND2_29531 ( P1_R2358_U407 , P1_U2614 , P1_R2358_U23 );
nand NAND2_29532 ( P1_R2358_U408 , P1_R2358_U407 , P1_R2358_U406 );
nand NAND2_29533 ( P1_R2358_U409 , P1_U2352 , P1_R2358_U146 );
nand NAND2_29534 ( P1_R2358_U410 , P1_U2667 , P1_R2358_U23 );
nand NAND2_29535 ( P1_R2358_U411 , P1_U2352 , P1_R2358_U147 );
nand NAND2_29536 ( P1_R2358_U412 , P1_U2668 , P1_R2358_U23 );
nand NAND2_29537 ( P1_R2358_U413 , P1_R2358_U412 , P1_R2358_U411 );
nand NAND2_29538 ( P1_R2358_U414 , P1_U2352 , P1_R2358_U146 );
nand NAND2_29539 ( P1_R2358_U415 , P1_U2667 , P1_R2358_U23 );
nand NAND2_29540 ( P1_R2358_U416 , P1_R2358_U415 , P1_R2358_U414 );
nand NAND2_29541 ( P1_R2358_U417 , P1_U2352 , P1_R2358_U145 );
nand NAND2_29542 ( P1_R2358_U418 , P1_U2614 , P1_R2358_U23 );
nand NAND2_29543 ( P1_R2358_U419 , P1_U2352 , P1_R2358_U144 );
nand NAND2_29544 ( P1_R2358_U420 , P1_U2615 , P1_R2358_U23 );
nand NAND2_29545 ( P1_R2358_U421 , P1_R2358_U420 , P1_R2358_U419 );
nand NAND2_29546 ( P1_R2358_U422 , P1_U2352 , P1_R2358_U148 );
nand NAND2_29547 ( P1_R2358_U423 , P1_U2670 , P1_R2358_U23 );
nand NAND2_29548 ( P1_R2358_U424 , P1_R2358_U423 , P1_R2358_U422 );
nand NAND2_29549 ( P1_R2358_U425 , P1_U2352 , P1_R2358_U149 );
nand NAND2_29550 ( P1_R2358_U426 , P1_U2671 , P1_R2358_U23 );
nand NAND2_29551 ( P1_R2358_U427 , P1_R2358_U426 , P1_R2358_U425 );
nand NAND2_29552 ( P1_R2358_U428 , P1_U2352 , P1_R2358_U150 );
nand NAND2_29553 ( P1_R2358_U429 , P1_U2672 , P1_R2358_U23 );
nand NAND2_29554 ( P1_R2358_U430 , P1_R2358_U429 , P1_R2358_U428 );
nand NAND2_29555 ( P1_R2358_U431 , P1_U2352 , P1_R2358_U149 );
nand NAND2_29556 ( P1_R2358_U432 , P1_U2671 , P1_R2358_U23 );
nand NAND2_29557 ( P1_R2358_U433 , P1_U2352 , P1_R2358_U150 );
nand NAND2_29558 ( P1_R2358_U434 , P1_U2672 , P1_R2358_U23 );
nand NAND2_29559 ( P1_R2358_U435 , P1_U2352 , P1_R2358_U148 );
nand NAND2_29560 ( P1_R2358_U436 , P1_U2670 , P1_R2358_U23 );
nand NAND2_29561 ( P1_R2358_U437 , P1_U2352 , P1_R2358_U151 );
nand NAND2_29562 ( P1_R2358_U438 , P1_U2669 , P1_R2358_U23 );
nand NAND2_29563 ( P1_R2358_U439 , P1_U2352 , P1_R2358_U151 );
nand NAND2_29564 ( P1_R2358_U440 , P1_U2669 , P1_R2358_U23 );
nand NAND2_29565 ( P1_R2358_U441 , P1_R2358_U440 , P1_R2358_U439 );
nand NAND2_29566 ( P1_R2358_U442 , P1_U2352 , P1_R2358_U147 );
nand NAND2_29567 ( P1_R2358_U443 , P1_U2668 , P1_R2358_U23 );
nand NAND2_29568 ( P1_R2358_U444 , P1_U2352 , P1_R2358_U152 );
nand NAND2_29569 ( P1_R2358_U445 , P1_U2617 , P1_R2358_U23 );
nand NAND2_29570 ( P1_R2358_U446 , P1_U2352 , P1_R2358_U152 );
nand NAND2_29571 ( P1_R2358_U447 , P1_U2617 , P1_R2358_U23 );
nand NAND2_29572 ( P1_R2358_U448 , P1_R2358_U447 , P1_R2358_U446 );
nand NAND2_29573 ( P1_R2358_U449 , P1_R2358_U332 , P1_R2358_U153 );
nand NAND2_29574 ( P1_R2358_U450 , P1_R2358_U77 , P1_R2358_U231 );
nand NAND2_29575 ( P1_R2358_U451 , P1_R2358_U333 , P1_R2358_U154 );
nand NAND2_29576 ( P1_R2358_U452 , P1_R2358_U79 , P1_R2358_U227 );
nand NAND2_29577 ( P1_R2358_U453 , P1_R2358_U334 , P1_R2358_U155 );
nand NAND2_29578 ( P1_R2358_U454 , P1_R2358_U81 , P1_R2358_U235 );
nand NAND2_29579 ( P1_R2358_U455 , P1_R2358_U335 , P1_R2358_U156 );
nand NAND2_29580 ( P1_R2358_U456 , P1_R2358_U83 , P1_R2358_U214 );
nand NAND2_29581 ( P1_R2358_U457 , P1_U2352 , P1_R2358_U157 );
nand NAND2_29582 ( P1_R2358_U458 , P1_U2611 , P1_R2358_U23 );
nand NAND2_29583 ( P1_R2358_U459 , P1_U2352 , P1_R2358_U158 );
nand NAND2_29584 ( P1_R2358_U460 , P1_U2612 , P1_R2358_U23 );
nand NAND2_29585 ( P1_R2358_U461 , P1_U2352 , P1_R2358_U159 );
nand NAND2_29586 ( P1_R2358_U462 , P1_U2613 , P1_R2358_U23 );
nand NAND2_29587 ( P1_R2358_U463 , P1_R2358_U462 , P1_R2358_U461 );
nand NAND2_29588 ( P1_R2358_U464 , P1_U2352 , P1_R2358_U158 );
nand NAND2_29589 ( P1_R2358_U465 , P1_U2612 , P1_R2358_U23 );
nand NAND2_29590 ( P1_R2358_U466 , P1_R2358_U465 , P1_R2358_U464 );
nand NAND2_29591 ( P1_R2358_U467 , P1_U2352 , P1_R2358_U159 );
nand NAND2_29592 ( P1_R2358_U468 , P1_U2613 , P1_R2358_U23 );
nand NAND2_29593 ( P1_R2358_U469 , P1_U2352 , P1_R2358_U160 );
nand NAND2_29594 ( P1_R2358_U470 , P1_U2616 , P1_R2358_U23 );
nand NAND2_29595 ( P1_R2358_U471 , P1_R2358_U470 , P1_R2358_U469 );
nand NAND2_29596 ( P1_R2358_U472 , P1_U2352 , P1_R2358_U157 );
nand NAND2_29597 ( P1_R2358_U473 , P1_U2611 , P1_R2358_U23 );
nand NAND2_29598 ( P1_R2358_U474 , P1_R2358_U473 , P1_R2358_U472 );
nand NAND2_29599 ( P1_R2358_U475 , P1_U2352 , P1_R2358_U161 );
nand NAND2_29600 ( P1_R2358_U476 , P1_U2610 , P1_R2358_U23 );
nand NAND2_29601 ( P1_R2358_U477 , P1_U2352 , P1_R2358_U161 );
nand NAND2_29602 ( P1_R2358_U478 , P1_U2610 , P1_R2358_U23 );
nand NAND2_29603 ( P1_R2358_U479 , P1_R2358_U478 , P1_R2358_U477 );
nand NAND2_29604 ( P1_R2358_U480 , P1_U2352 , P1_R2358_U162 );
nand NAND2_29605 ( P1_R2358_U481 , P1_U2609 , P1_R2358_U23 );
nand NAND2_29606 ( P1_R2358_U482 , P1_U2352 , P1_R2358_U162 );
nand NAND2_29607 ( P1_R2358_U483 , P1_U2609 , P1_R2358_U23 );
nand NAND2_29608 ( P1_R2358_U484 , P1_R2358_U483 , P1_R2358_U482 );
nand NAND2_29609 ( P1_R2358_U485 , P1_U2352 , P1_R2358_U160 );
nand NAND2_29610 ( P1_R2358_U486 , P1_U2616 , P1_R2358_U23 );
nand NAND2_29611 ( P1_R2358_U487 , P1_U2352 , P1_R2358_U163 );
nand NAND2_29612 ( P1_R2358_U488 , P1_U2666 , P1_R2358_U23 );
nand NAND2_29613 ( P1_R2358_U489 , P1_U2352 , P1_R2358_U164 );
nand NAND2_29614 ( P1_R2358_U490 , P1_U2665 , P1_R2358_U23 );
nand NAND2_29615 ( P1_R2358_U491 , P1_U2352 , P1_R2358_U165 );
nand NAND2_29616 ( P1_R2358_U492 , P1_U2664 , P1_R2358_U23 );
nand NAND2_29617 ( P1_R2358_U493 , P1_U2352 , P1_R2358_U165 );
nand NAND2_29618 ( P1_R2358_U494 , P1_U2664 , P1_R2358_U23 );
nand NAND2_29619 ( P1_R2358_U495 , P1_R2358_U494 , P1_R2358_U493 );
nand NAND2_29620 ( P1_R2358_U496 , P1_U2352 , P1_R2358_U164 );
nand NAND2_29621 ( P1_R2358_U497 , P1_U2665 , P1_R2358_U23 );
nand NAND2_29622 ( P1_R2358_U498 , P1_R2358_U497 , P1_R2358_U496 );
nand NAND2_29623 ( P1_R2358_U499 , P1_U2352 , P1_R2358_U163 );
nand NAND2_29624 ( P1_R2358_U500 , P1_U2666 , P1_R2358_U23 );
nand NAND2_29625 ( P1_R2358_U501 , P1_R2358_U500 , P1_R2358_U499 );
nand NAND2_29626 ( P1_R2358_U502 , P1_U2352 , P1_R2358_U166 );
nand NAND2_29627 ( P1_R2358_U503 , P1_U2660 , P1_R2358_U23 );
nand NAND2_29628 ( P1_R2358_U504 , P1_U2352 , P1_R2358_U167 );
nand NAND2_29629 ( P1_R2358_U505 , P1_U2661 , P1_R2358_U23 );
nand NAND2_29630 ( P1_R2358_U506 , P1_U2352 , P1_R2358_U168 );
nand NAND2_29631 ( P1_R2358_U507 , P1_U2663 , P1_R2358_U23 );
nand NAND2_29632 ( P1_R2358_U508 , P1_U2352 , P1_R2358_U169 );
nand NAND2_29633 ( P1_R2358_U509 , P1_U2662 , P1_R2358_U23 );
nand NAND2_29634 ( P1_R2358_U510 , P1_U2352 , P1_R2358_U166 );
nand NAND2_29635 ( P1_R2358_U511 , P1_U2660 , P1_R2358_U23 );
nand NAND2_29636 ( P1_R2358_U512 , P1_R2358_U511 , P1_R2358_U510 );
nand NAND2_29637 ( P1_R2358_U513 , P1_U2352 , P1_R2358_U167 );
nand NAND2_29638 ( P1_R2358_U514 , P1_U2661 , P1_R2358_U23 );
nand NAND2_29639 ( P1_R2358_U515 , P1_R2358_U514 , P1_R2358_U513 );
nand NAND2_29640 ( P1_R2358_U516 , P1_U2352 , P1_R2358_U169 );
nand NAND2_29641 ( P1_R2358_U517 , P1_U2662 , P1_R2358_U23 );
nand NAND2_29642 ( P1_R2358_U518 , P1_R2358_U517 , P1_R2358_U516 );
nand NAND2_29643 ( P1_R2358_U519 , P1_U2352 , P1_R2358_U168 );
nand NAND2_29644 ( P1_R2358_U520 , P1_U2663 , P1_R2358_U23 );
nand NAND2_29645 ( P1_R2358_U521 , P1_R2358_U520 , P1_R2358_U519 );
nand NAND2_29646 ( P1_R2358_U522 , P1_U2352 , P1_R2358_U170 );
nand NAND2_29647 ( P1_R2358_U523 , P1_U2655 , P1_R2358_U23 );
nand NAND2_29648 ( P1_R2358_U524 , P1_U2352 , P1_R2358_U171 );
nand NAND2_29649 ( P1_R2358_U525 , P1_U2656 , P1_R2358_U23 );
nand NAND2_29650 ( P1_R2358_U526 , P1_U2352 , P1_R2358_U172 );
nand NAND2_29651 ( P1_R2358_U527 , P1_U2657 , P1_R2358_U23 );
nand NAND2_29652 ( P1_R2358_U528 , P1_U2352 , P1_R2358_U173 );
nand NAND2_29653 ( P1_R2358_U529 , P1_U2659 , P1_R2358_U23 );
nand NAND2_29654 ( P1_R2358_U530 , P1_U2352 , P1_R2358_U174 );
nand NAND2_29655 ( P1_R2358_U531 , P1_U2658 , P1_R2358_U23 );
nand NAND2_29656 ( P1_R2358_U532 , P1_U2352 , P1_R2358_U170 );
nand NAND2_29657 ( P1_R2358_U533 , P1_U2655 , P1_R2358_U23 );
nand NAND2_29658 ( P1_R2358_U534 , P1_R2358_U533 , P1_R2358_U532 );
nand NAND2_29659 ( P1_R2358_U535 , P1_U2352 , P1_R2358_U171 );
nand NAND2_29660 ( P1_R2358_U536 , P1_U2656 , P1_R2358_U23 );
nand NAND2_29661 ( P1_R2358_U537 , P1_R2358_U536 , P1_R2358_U535 );
nand NAND2_29662 ( P1_R2358_U538 , P1_U2352 , P1_R2358_U172 );
nand NAND2_29663 ( P1_R2358_U539 , P1_U2657 , P1_R2358_U23 );
nand NAND2_29664 ( P1_R2358_U540 , P1_R2358_U539 , P1_R2358_U538 );
nand NAND2_29665 ( P1_R2358_U541 , P1_U2352 , P1_R2358_U174 );
nand NAND2_29666 ( P1_R2358_U542 , P1_U2658 , P1_R2358_U23 );
nand NAND2_29667 ( P1_R2358_U543 , P1_R2358_U542 , P1_R2358_U541 );
nand NAND2_29668 ( P1_R2358_U544 , P1_U2352 , P1_R2358_U173 );
nand NAND2_29669 ( P1_R2358_U545 , P1_U2659 , P1_R2358_U23 );
nand NAND2_29670 ( P1_R2358_U546 , P1_R2358_U545 , P1_R2358_U544 );
nand NAND2_29671 ( P1_R2358_U547 , P1_U2352 , P1_R2358_U175 );
nand NAND2_29672 ( P1_R2358_U548 , P1_U2654 , P1_R2358_U23 );
nand NAND2_29673 ( P1_R2358_U549 , P1_U2352 , P1_R2358_U175 );
nand NAND2_29674 ( P1_R2358_U550 , P1_U2654 , P1_R2358_U23 );
nand NAND2_29675 ( P1_R2358_U551 , P1_R2358_U550 , P1_R2358_U549 );
nand NAND2_29676 ( P1_R2358_U552 , P1_U2352 , P1_R2358_U176 );
nand NAND2_29677 ( P1_R2358_U553 , P1_U2653 , P1_R2358_U23 );
nand NAND2_29678 ( P1_R2358_U554 , P1_U2352 , P1_R2358_U177 );
nand NAND2_29679 ( P1_R2358_U555 , P1_U2651 , P1_R2358_U23 );
nand NAND2_29680 ( P1_R2358_U556 , P1_U2352 , P1_R2358_U178 );
nand NAND2_29681 ( P1_R2358_U557 , P1_U2652 , P1_R2358_U23 );
not NOT1_29682 ( P1_R2358_U558 , P1_R2358_U75 );
nand NAND2_29683 ( P1_R2358_U559 , P1_U2352 , P1_R2358_U177 );
nand NAND2_29684 ( P1_R2358_U560 , P1_U2651 , P1_R2358_U23 );
nand NAND2_29685 ( P1_R2358_U561 , P1_R2358_U560 , P1_R2358_U559 );
nand NAND2_29686 ( P1_R2358_U562 , P1_U2352 , P1_R2358_U176 );
nand NAND2_29687 ( P1_R2358_U563 , P1_U2653 , P1_R2358_U23 );
nand NAND2_29688 ( P1_R2358_U564 , P1_R2358_U563 , P1_R2358_U562 );
nand NAND3_29689 ( P1_R2358_U565 , P1_R2358_U135 , P1_R2358_U302 , P1_R2358_U179 );
nand NAND3_29690 ( P1_R2358_U566 , P1_R2358_U561 , P1_R2358_U305 , P1_R2358_U301 );
nand NAND3_29691 ( P1_R2358_U567 , P1_R2358_U13 , P1_R2358_U558 , P1_R2358_U63 );
nand NAND3_29692 ( P1_R2358_U568 , P1_R2358_U561 , P1_R2358_U75 , P1_U2620 );
nand NAND2_29693 ( P1_R2358_U569 , P1_R2358_U558 , P1_U2620 );
nand NAND2_29694 ( P1_R2358_U570 , P1_R2358_U75 , P1_R2358_U63 );
nand NAND2_29695 ( P1_R2358_U571 , P1_R2358_U558 , P1_U2620 );
nand NAND2_29696 ( P1_R2358_U572 , P1_R2358_U75 , P1_R2358_U63 );
nand NAND2_29697 ( P1_R2358_U573 , P1_R2358_U572 , P1_R2358_U571 );
nand NAND2_29698 ( P1_R2358_U574 , P1_R2358_U181 , P1_R2358_U182 );
nand NAND2_29699 ( P1_R2358_U575 , P1_R2358_U303 , P1_R2358_U573 );
nand NAND2_29700 ( P1_R2358_U576 , P1_R2358_U336 , P1_R2358_U183 );
nand NAND2_29701 ( P1_R2358_U577 , P1_R2358_U86 , P1_R2358_U299 );
nand NAND2_29702 ( P1_R2358_U578 , P1_R2358_U184 , P1_R2358_U337 );
nand NAND2_29703 ( P1_R2358_U579 , P1_R2358_U88 , P1_R2358_U384 );
nand NAND2_29704 ( P1_R2358_U580 , P1_R2358_U185 , P1_R2358_U338 );
nand NAND2_29705 ( P1_R2358_U581 , P1_R2358_U90 , P1_R2358_U382 );
nand NAND2_29706 ( P1_R2358_U582 , P1_R2358_U186 , P1_R2358_U339 );
nand NAND2_29707 ( P1_R2358_U583 , P1_R2358_U92 , P1_R2358_U380 );
nand NAND2_29708 ( P1_R2358_U584 , P1_R2358_U187 , P1_R2358_U340 );
nand NAND2_29709 ( P1_R2358_U585 , P1_R2358_U94 , P1_R2358_U378 );
nand NAND2_29710 ( P1_R2358_U586 , P1_R2358_U188 , P1_R2358_U341 );
nand NAND2_29711 ( P1_R2358_U587 , P1_R2358_U96 , P1_R2358_U376 );
nand NAND2_29712 ( P1_R2358_U588 , P1_R2358_U189 , P1_R2358_U342 );
nand NAND2_29713 ( P1_R2358_U589 , P1_R2358_U98 , P1_R2358_U386 );
nand NAND2_29714 ( P1_R2358_U590 , P1_R2358_U190 , P1_R2358_U343 );
nand NAND2_29715 ( P1_R2358_U591 , P1_R2358_U100 , P1_R2358_U388 );
nand NAND2_29716 ( P1_R2358_U592 , P1_R2358_U191 , P1_R2358_U344 );
nand NAND2_29717 ( P1_R2358_U593 , P1_R2358_U102 , P1_R2358_U390 );
nand NAND2_29718 ( P1_R2358_U594 , P1_R2358_U192 , P1_R2358_U345 );
nand NAND2_29719 ( P1_R2358_U595 , P1_R2358_U104 , P1_R2358_U392 );
nand NAND2_29720 ( P1_R2358_U596 , P1_R2358_U346 , P1_R2358_U193 );
nand NAND2_29721 ( P1_R2358_U597 , P1_R2358_U106 , P1_R2358_U247 );
nand NAND2_29722 ( P1_R2358_U598 , P1_R2358_U194 , P1_R2358_U347 );
nand NAND2_29723 ( P1_R2358_U599 , P1_R2358_U108 , P1_R2358_U394 );
nand NAND2_29724 ( P1_R2358_U600 , P1_R2358_U195 , P1_R2358_U348 );
nand NAND2_29725 ( P1_R2358_U601 , P1_R2358_U110 , P1_R2358_U396 );
nand NAND2_29726 ( P1_R2358_U602 , P1_R2358_U196 , P1_R2358_U349 );
nand NAND2_29727 ( P1_R2358_U603 , P1_R2358_U112 , P1_R2358_U398 );
nand NAND2_29728 ( P1_R2358_U604 , P1_R2358_U350 , P1_R2358_U197 );
nand NAND2_29729 ( P1_R2358_U605 , P1_R2358_U114 , P1_R2358_U271 );
nand NAND2_29730 ( P1_R2358_U606 , P1_R2358_U351 , P1_R2358_U198 );
nand NAND2_29731 ( P1_R2358_U607 , P1_R2358_U116 , P1_R2358_U310 );
nand NAND2_29732 ( P1_R2358_U608 , P1_R2358_U352 , P1_R2358_U199 );
nand NAND2_29733 ( P1_R2358_U609 , P1_R2358_U118 , P1_R2358_U269 );
nand NAND2_29734 ( P1_R2358_U610 , P1_U2352 , P1_R2358_U200 );
nand NAND2_29735 ( P1_R2358_U611 , P1_R2358_U331 , P1_R2358_U23 );
or OR2_29736 ( P1_LT_589_U6 , P1_LT_589_U8 , P1_U2673 );
and AND2_29737 ( P1_LT_589_U7 , P1_R584_U7 , P1_R584_U6 );
nor nor_29738 ( P1_LT_589_U8 , P1_LT_589_U7 , P1_R584_U9 , P1_R584_U8 );
not NOT1_29739 ( P1_R584_U6 , P1_U2676 );
not NOT1_29740 ( P1_R584_U7 , P1_U2677 );
not NOT1_29741 ( P1_R584_U8 , P1_U2674 );
not NOT1_29742 ( P1_R584_U9 , P1_U2675 );
not NOT1_29743 ( P1_R2099_U4 , P1_U4190 );
not NOT1_29744 ( P1_R2099_U5 , P1_U4189 );
not NOT1_29745 ( P1_R2099_U6 , P1_U2678 );
nand NAND2_29746 ( P1_R2099_U7 , P1_R2099_U88 , P1_R2099_U137 );
nand NAND2_29747 ( P1_R2099_U8 , P1_R2099_U89 , P1_R2099_U155 );
nand NAND2_29748 ( P1_R2099_U9 , P1_R2099_U90 , P1_R2099_U157 );
nand NAND2_29749 ( P1_R2099_U10 , P1_R2099_U91 , P1_R2099_U159 );
nand NAND2_29750 ( P1_R2099_U11 , P1_R2099_U92 , P1_R2099_U161 );
nand NAND2_29751 ( P1_R2099_U12 , P1_R2099_U93 , P1_R2099_U163 );
nand NAND2_29752 ( P1_R2099_U13 , P1_R2099_U94 , P1_R2099_U165 );
nand NAND2_29753 ( P1_R2099_U14 , P1_R2099_U95 , P1_R2099_U167 );
nand NAND2_29754 ( P1_R2099_U15 , P1_R2099_U169 , P1_R2099_U55 );
nand NAND2_29755 ( P1_R2099_U16 , P1_R2099_U170 , P1_R2099_U54 );
nand NAND2_29756 ( P1_R2099_U17 , P1_R2099_U171 , P1_R2099_U53 );
nand NAND2_29757 ( P1_R2099_U18 , P1_R2099_U172 , P1_R2099_U52 );
nand NAND2_29758 ( P1_R2099_U19 , P1_R2099_U173 , P1_R2099_U51 );
nand NAND2_29759 ( P1_R2099_U20 , P1_R2099_U174 , P1_R2099_U50 );
nand NAND2_29760 ( P1_R2099_U21 , P1_R2099_U175 , P1_R2099_U49 );
nand NAND2_29761 ( P1_R2099_U22 , P1_R2099_U176 , P1_R2099_U48 );
nand NAND2_29762 ( P1_R2099_U23 , P1_R2099_U177 , P1_R2099_U47 );
nand NAND2_29763 ( P1_R2099_U24 , P1_R2099_U178 , P1_R2099_U46 );
nand NAND2_29764 ( P1_R2099_U25 , P1_R2099_U179 , P1_R2099_U45 );
nand NAND2_29765 ( P1_R2099_U26 , P1_R2099_U210 , P1_R2099_U209 );
nand NAND2_29766 ( P1_R2099_U27 , P1_R2099_U183 , P1_R2099_U182 );
nand NAND2_29767 ( P1_R2099_U28 , P1_R2099_U204 , P1_R2099_U203 );
nand NAND2_29768 ( P1_R2099_U29 , P1_R2099_U207 , P1_R2099_U206 );
nand NAND2_29769 ( P1_R2099_U30 , P1_R2099_U198 , P1_R2099_U197 );
nand NAND2_29770 ( P1_R2099_U31 , P1_R2099_U201 , P1_R2099_U200 );
nand NAND2_29771 ( P1_R2099_U32 , P1_R2099_U186 , P1_R2099_U185 );
nand NAND2_29772 ( P1_R2099_U33 , P1_R2099_U189 , P1_R2099_U188 );
nand NAND2_29773 ( P1_R2099_U34 , P1_R2099_U195 , P1_R2099_U194 );
nand NAND2_29774 ( P1_R2099_U35 , P1_R2099_U192 , P1_R2099_U191 );
nand NAND2_29775 ( P1_R2099_U36 , P1_R2099_U213 , P1_R2099_U212 );
nand NAND2_29776 ( P1_R2099_U37 , P1_R2099_U215 , P1_R2099_U214 );
nand NAND2_29777 ( P1_R2099_U38 , P1_R2099_U217 , P1_R2099_U216 );
nand NAND2_29778 ( P1_R2099_U39 , P1_R2099_U219 , P1_R2099_U218 );
nand NAND2_29779 ( P1_R2099_U40 , P1_R2099_U221 , P1_R2099_U220 );
nand NAND2_29780 ( P1_R2099_U41 , P1_R2099_U223 , P1_R2099_U222 );
nand NAND2_29781 ( P1_R2099_U42 , P1_R2099_U225 , P1_R2099_U224 );
nand NAND2_29782 ( P1_R2099_U43 , P1_R2099_U284 , P1_R2099_U283 );
nand NAND2_29783 ( P1_R2099_U44 , P1_R2099_U287 , P1_R2099_U286 );
nand NAND2_29784 ( P1_R2099_U45 , P1_R2099_U227 , P1_R2099_U226 );
nand NAND2_29785 ( P1_R2099_U46 , P1_R2099_U230 , P1_R2099_U229 );
nand NAND2_29786 ( P1_R2099_U47 , P1_R2099_U233 , P1_R2099_U232 );
nand NAND2_29787 ( P1_R2099_U48 , P1_R2099_U236 , P1_R2099_U235 );
nand NAND2_29788 ( P1_R2099_U49 , P1_R2099_U239 , P1_R2099_U238 );
nand NAND2_29789 ( P1_R2099_U50 , P1_R2099_U242 , P1_R2099_U241 );
nand NAND2_29790 ( P1_R2099_U51 , P1_R2099_U245 , P1_R2099_U244 );
nand NAND2_29791 ( P1_R2099_U52 , P1_R2099_U248 , P1_R2099_U247 );
nand NAND2_29792 ( P1_R2099_U53 , P1_R2099_U251 , P1_R2099_U250 );
nand NAND2_29793 ( P1_R2099_U54 , P1_R2099_U254 , P1_R2099_U253 );
nand NAND2_29794 ( P1_R2099_U55 , P1_R2099_U257 , P1_R2099_U256 );
nand NAND2_29795 ( P1_R2099_U56 , P1_R2099_U278 , P1_R2099_U277 );
nand NAND2_29796 ( P1_R2099_U57 , P1_R2099_U281 , P1_R2099_U280 );
nand NAND2_29797 ( P1_R2099_U58 , P1_R2099_U272 , P1_R2099_U271 );
nand NAND2_29798 ( P1_R2099_U59 , P1_R2099_U275 , P1_R2099_U274 );
nand NAND2_29799 ( P1_R2099_U60 , P1_R2099_U266 , P1_R2099_U265 );
nand NAND2_29800 ( P1_R2099_U61 , P1_R2099_U269 , P1_R2099_U268 );
nand NAND2_29801 ( P1_R2099_U62 , P1_R2099_U260 , P1_R2099_U259 );
nand NAND2_29802 ( P1_R2099_U63 , P1_R2099_U263 , P1_R2099_U262 );
nand NAND2_29803 ( P1_R2099_U64 , P1_R2099_U293 , P1_R2099_U292 );
nand NAND2_29804 ( P1_R2099_U65 , P1_R2099_U295 , P1_R2099_U294 );
nand NAND2_29805 ( P1_R2099_U66 , P1_R2099_U299 , P1_R2099_U298 );
nand NAND2_29806 ( P1_R2099_U67 , P1_R2099_U301 , P1_R2099_U300 );
nand NAND2_29807 ( P1_R2099_U68 , P1_R2099_U303 , P1_R2099_U302 );
nand NAND2_29808 ( P1_R2099_U69 , P1_R2099_U305 , P1_R2099_U304 );
nand NAND2_29809 ( P1_R2099_U70 , P1_R2099_U307 , P1_R2099_U306 );
nand NAND2_29810 ( P1_R2099_U71 , P1_R2099_U309 , P1_R2099_U308 );
nand NAND2_29811 ( P1_R2099_U72 , P1_R2099_U311 , P1_R2099_U310 );
nand NAND2_29812 ( P1_R2099_U73 , P1_R2099_U313 , P1_R2099_U312 );
nand NAND2_29813 ( P1_R2099_U74 , P1_R2099_U315 , P1_R2099_U314 );
nand NAND2_29814 ( P1_R2099_U75 , P1_R2099_U317 , P1_R2099_U316 );
nand NAND2_29815 ( P1_R2099_U76 , P1_R2099_U326 , P1_R2099_U325 );
nand NAND2_29816 ( P1_R2099_U77 , P1_R2099_U328 , P1_R2099_U327 );
nand NAND2_29817 ( P1_R2099_U78 , P1_R2099_U330 , P1_R2099_U329 );
nand NAND2_29818 ( P1_R2099_U79 , P1_R2099_U332 , P1_R2099_U331 );
nand NAND2_29819 ( P1_R2099_U80 , P1_R2099_U334 , P1_R2099_U333 );
nand NAND2_29820 ( P1_R2099_U81 , P1_R2099_U336 , P1_R2099_U335 );
nand NAND2_29821 ( P1_R2099_U82 , P1_R2099_U338 , P1_R2099_U337 );
nand NAND2_29822 ( P1_R2099_U83 , P1_R2099_U340 , P1_R2099_U339 );
nand NAND2_29823 ( P1_R2099_U84 , P1_R2099_U342 , P1_R2099_U341 );
nand NAND2_29824 ( P1_R2099_U85 , P1_R2099_U344 , P1_R2099_U343 );
nand NAND2_29825 ( P1_R2099_U86 , P1_R2099_U349 , P1_R2099_U348 );
nand NAND2_29826 ( P1_R2099_U87 , P1_R2099_U324 , P1_R2099_U323 );
and AND2_29827 ( P1_R2099_U88 , P1_R2099_U34 , P1_R2099_U35 );
and AND2_29828 ( P1_R2099_U89 , P1_R2099_U31 , P1_R2099_U30 );
and AND2_29829 ( P1_R2099_U90 , P1_R2099_U29 , P1_R2099_U28 );
and AND2_29830 ( P1_R2099_U91 , P1_R2099_U26 , P1_R2099_U27 );
and AND2_29831 ( P1_R2099_U92 , P1_R2099_U63 , P1_R2099_U62 );
and AND2_29832 ( P1_R2099_U93 , P1_R2099_U61 , P1_R2099_U60 );
and AND2_29833 ( P1_R2099_U94 , P1_R2099_U59 , P1_R2099_U58 );
and AND2_29834 ( P1_R2099_U95 , P1_R2099_U57 , P1_R2099_U56 );
and AND2_29835 ( P1_R2099_U96 , P1_R2099_U44 , P1_R2099_U43 );
nand NAND2_29836 ( P1_R2099_U97 , P1_R2099_U290 , P1_R2099_U289 );
nand NAND2_29837 ( P1_R2099_U98 , P1_R2099_U346 , P1_R2099_U345 );
not NOT1_29838 ( P1_R2099_U99 , P1_U2702 );
not NOT1_29839 ( P1_R2099_U100 , P1_U2710 );
not NOT1_29840 ( P1_R2099_U101 , P1_U2709 );
not NOT1_29841 ( P1_R2099_U102 , P1_U2708 );
not NOT1_29842 ( P1_R2099_U103 , P1_U2707 );
not NOT1_29843 ( P1_R2099_U104 , P1_U2706 );
not NOT1_29844 ( P1_R2099_U105 , P1_U2705 );
not NOT1_29845 ( P1_R2099_U106 , P1_U2704 );
not NOT1_29846 ( P1_R2099_U107 , P1_U2703 );
not NOT1_29847 ( P1_R2099_U108 , P1_U2701 );
nand NAND2_29848 ( P1_R2099_U109 , P1_R2099_U159 , P1_R2099_U27 );
nand NAND2_29849 ( P1_R2099_U110 , P1_R2099_U157 , P1_R2099_U28 );
nand NAND2_29850 ( P1_R2099_U111 , P1_R2099_U155 , P1_R2099_U30 );
nand NAND2_29851 ( P1_R2099_U112 , P1_R2099_U35 , P1_R2099_U137 );
not NOT1_29852 ( P1_R2099_U113 , P1_U2682 );
not NOT1_29853 ( P1_R2099_U114 , P1_U2683 );
not NOT1_29854 ( P1_R2099_U115 , P1_U2684 );
not NOT1_29855 ( P1_R2099_U116 , P1_U2685 );
not NOT1_29856 ( P1_R2099_U117 , P1_U2686 );
not NOT1_29857 ( P1_R2099_U118 , P1_U2687 );
not NOT1_29858 ( P1_R2099_U119 , P1_U2688 );
not NOT1_29859 ( P1_R2099_U120 , P1_U2689 );
not NOT1_29860 ( P1_R2099_U121 , P1_U2690 );
not NOT1_29861 ( P1_R2099_U122 , P1_U2691 );
not NOT1_29862 ( P1_R2099_U123 , P1_U2692 );
not NOT1_29863 ( P1_R2099_U124 , P1_U2700 );
not NOT1_29864 ( P1_R2099_U125 , P1_U2699 );
not NOT1_29865 ( P1_R2099_U126 , P1_U2698 );
not NOT1_29866 ( P1_R2099_U127 , P1_U2697 );
not NOT1_29867 ( P1_R2099_U128 , P1_U2696 );
not NOT1_29868 ( P1_R2099_U129 , P1_U2695 );
not NOT1_29869 ( P1_R2099_U130 , P1_U2694 );
not NOT1_29870 ( P1_R2099_U131 , P1_U2693 );
not NOT1_29871 ( P1_R2099_U132 , P1_U2680 );
not NOT1_29872 ( P1_R2099_U133 , P1_U2681 );
not NOT1_29873 ( P1_R2099_U134 , P1_U2679 );
nand NAND2_29874 ( P1_R2099_U135 , P1_R2099_U96 , P1_R2099_U180 );
nand NAND2_29875 ( P1_R2099_U136 , P1_R2099_U180 , P1_R2099_U44 );
nand NAND2_29876 ( P1_R2099_U137 , P1_R2099_U152 , P1_R2099_U151 );
and AND2_29877 ( P1_R2099_U138 , P1_R2099_U297 , P1_R2099_U296 );
and AND2_29878 ( P1_R2099_U139 , P1_R2099_U319 , P1_R2099_U318 );
nand NAND2_29879 ( P1_R2099_U140 , P1_R2099_U148 , P1_R2099_U147 );
nand NAND2_29880 ( P1_R2099_U141 , P1_R2099_U167 , P1_R2099_U56 );
nand NAND2_29881 ( P1_R2099_U142 , P1_R2099_U165 , P1_R2099_U58 );
nand NAND2_29882 ( P1_R2099_U143 , P1_R2099_U163 , P1_R2099_U60 );
nand NAND2_29883 ( P1_R2099_U144 , P1_R2099_U161 , P1_R2099_U62 );
not NOT1_29884 ( P1_R2099_U145 , P1_R2099_U135 );
or OR2_29885 ( P1_R2099_U146 , P1_U4190 , P1_U4189 );
nand NAND2_29886 ( P1_R2099_U147 , P1_R2099_U32 , P1_R2099_U146 );
nand NAND2_29887 ( P1_R2099_U148 , P1_U4189 , P1_U4190 );
not NOT1_29888 ( P1_R2099_U149 , P1_R2099_U140 );
nand NAND2_29889 ( P1_R2099_U150 , P1_R2099_U190 , P1_R2099_U6 );
nand NAND2_29890 ( P1_R2099_U151 , P1_R2099_U150 , P1_R2099_U140 );
nand NAND2_29891 ( P1_R2099_U152 , P1_U2678 , P1_R2099_U33 );
not NOT1_29892 ( P1_R2099_U153 , P1_R2099_U137 );
not NOT1_29893 ( P1_R2099_U154 , P1_R2099_U112 );
not NOT1_29894 ( P1_R2099_U155 , P1_R2099_U7 );
not NOT1_29895 ( P1_R2099_U156 , P1_R2099_U111 );
not NOT1_29896 ( P1_R2099_U157 , P1_R2099_U8 );
not NOT1_29897 ( P1_R2099_U158 , P1_R2099_U110 );
not NOT1_29898 ( P1_R2099_U159 , P1_R2099_U9 );
not NOT1_29899 ( P1_R2099_U160 , P1_R2099_U109 );
not NOT1_29900 ( P1_R2099_U161 , P1_R2099_U10 );
not NOT1_29901 ( P1_R2099_U162 , P1_R2099_U144 );
not NOT1_29902 ( P1_R2099_U163 , P1_R2099_U11 );
not NOT1_29903 ( P1_R2099_U164 , P1_R2099_U143 );
not NOT1_29904 ( P1_R2099_U165 , P1_R2099_U12 );
not NOT1_29905 ( P1_R2099_U166 , P1_R2099_U142 );
not NOT1_29906 ( P1_R2099_U167 , P1_R2099_U13 );
not NOT1_29907 ( P1_R2099_U168 , P1_R2099_U141 );
not NOT1_29908 ( P1_R2099_U169 , P1_R2099_U14 );
not NOT1_29909 ( P1_R2099_U170 , P1_R2099_U15 );
not NOT1_29910 ( P1_R2099_U171 , P1_R2099_U16 );
not NOT1_29911 ( P1_R2099_U172 , P1_R2099_U17 );
not NOT1_29912 ( P1_R2099_U173 , P1_R2099_U18 );
not NOT1_29913 ( P1_R2099_U174 , P1_R2099_U19 );
not NOT1_29914 ( P1_R2099_U175 , P1_R2099_U20 );
not NOT1_29915 ( P1_R2099_U176 , P1_R2099_U21 );
not NOT1_29916 ( P1_R2099_U177 , P1_R2099_U22 );
not NOT1_29917 ( P1_R2099_U178 , P1_R2099_U23 );
not NOT1_29918 ( P1_R2099_U179 , P1_R2099_U24 );
not NOT1_29919 ( P1_R2099_U180 , P1_R2099_U25 );
not NOT1_29920 ( P1_R2099_U181 , P1_R2099_U136 );
nand NAND2_29921 ( P1_R2099_U182 , P1_U4190 , P1_R2099_U99 );
nand NAND2_29922 ( P1_R2099_U183 , P1_U2702 , P1_R2099_U4 );
not NOT1_29923 ( P1_R2099_U184 , P1_R2099_U27 );
nand NAND2_29924 ( P1_R2099_U185 , P1_U4190 , P1_R2099_U100 );
nand NAND2_29925 ( P1_R2099_U186 , P1_U2710 , P1_R2099_U4 );
not NOT1_29926 ( P1_R2099_U187 , P1_R2099_U32 );
nand NAND2_29927 ( P1_R2099_U188 , P1_U4190 , P1_R2099_U101 );
nand NAND2_29928 ( P1_R2099_U189 , P1_U2709 , P1_R2099_U4 );
not NOT1_29929 ( P1_R2099_U190 , P1_R2099_U33 );
nand NAND2_29930 ( P1_R2099_U191 , P1_U4190 , P1_R2099_U102 );
nand NAND2_29931 ( P1_R2099_U192 , P1_U2708 , P1_R2099_U4 );
not NOT1_29932 ( P1_R2099_U193 , P1_R2099_U35 );
nand NAND2_29933 ( P1_R2099_U194 , P1_U4190 , P1_R2099_U103 );
nand NAND2_29934 ( P1_R2099_U195 , P1_U2707 , P1_R2099_U4 );
not NOT1_29935 ( P1_R2099_U196 , P1_R2099_U34 );
nand NAND2_29936 ( P1_R2099_U197 , P1_U4190 , P1_R2099_U104 );
nand NAND2_29937 ( P1_R2099_U198 , P1_U2706 , P1_R2099_U4 );
not NOT1_29938 ( P1_R2099_U199 , P1_R2099_U30 );
nand NAND2_29939 ( P1_R2099_U200 , P1_U4190 , P1_R2099_U105 );
nand NAND2_29940 ( P1_R2099_U201 , P1_U2705 , P1_R2099_U4 );
not NOT1_29941 ( P1_R2099_U202 , P1_R2099_U31 );
nand NAND2_29942 ( P1_R2099_U203 , P1_U4190 , P1_R2099_U106 );
nand NAND2_29943 ( P1_R2099_U204 , P1_U2704 , P1_R2099_U4 );
not NOT1_29944 ( P1_R2099_U205 , P1_R2099_U28 );
nand NAND2_29945 ( P1_R2099_U206 , P1_U4190 , P1_R2099_U107 );
nand NAND2_29946 ( P1_R2099_U207 , P1_U2703 , P1_R2099_U4 );
not NOT1_29947 ( P1_R2099_U208 , P1_R2099_U29 );
nand NAND2_29948 ( P1_R2099_U209 , P1_U4190 , P1_R2099_U108 );
nand NAND2_29949 ( P1_R2099_U210 , P1_U2701 , P1_R2099_U4 );
not NOT1_29950 ( P1_R2099_U211 , P1_R2099_U26 );
nand NAND2_29951 ( P1_R2099_U212 , P1_R2099_U160 , P1_R2099_U211 );
nand NAND2_29952 ( P1_R2099_U213 , P1_R2099_U26 , P1_R2099_U109 );
nand NAND2_29953 ( P1_R2099_U214 , P1_R2099_U184 , P1_R2099_U159 );
nand NAND2_29954 ( P1_R2099_U215 , P1_R2099_U27 , P1_R2099_U9 );
nand NAND2_29955 ( P1_R2099_U216 , P1_R2099_U158 , P1_R2099_U208 );
nand NAND2_29956 ( P1_R2099_U217 , P1_R2099_U29 , P1_R2099_U110 );
nand NAND2_29957 ( P1_R2099_U218 , P1_R2099_U205 , P1_R2099_U157 );
nand NAND2_29958 ( P1_R2099_U219 , P1_R2099_U28 , P1_R2099_U8 );
nand NAND2_29959 ( P1_R2099_U220 , P1_R2099_U156 , P1_R2099_U202 );
nand NAND2_29960 ( P1_R2099_U221 , P1_R2099_U31 , P1_R2099_U111 );
nand NAND2_29961 ( P1_R2099_U222 , P1_R2099_U199 , P1_R2099_U155 );
nand NAND2_29962 ( P1_R2099_U223 , P1_R2099_U30 , P1_R2099_U7 );
nand NAND2_29963 ( P1_R2099_U224 , P1_R2099_U154 , P1_R2099_U196 );
nand NAND2_29964 ( P1_R2099_U225 , P1_R2099_U34 , P1_R2099_U112 );
nand NAND2_29965 ( P1_R2099_U226 , P1_U4190 , P1_R2099_U113 );
nand NAND2_29966 ( P1_R2099_U227 , P1_U2682 , P1_R2099_U4 );
not NOT1_29967 ( P1_R2099_U228 , P1_R2099_U45 );
nand NAND2_29968 ( P1_R2099_U229 , P1_U4190 , P1_R2099_U114 );
nand NAND2_29969 ( P1_R2099_U230 , P1_U2683 , P1_R2099_U4 );
not NOT1_29970 ( P1_R2099_U231 , P1_R2099_U46 );
nand NAND2_29971 ( P1_R2099_U232 , P1_U4190 , P1_R2099_U115 );
nand NAND2_29972 ( P1_R2099_U233 , P1_U2684 , P1_R2099_U4 );
not NOT1_29973 ( P1_R2099_U234 , P1_R2099_U47 );
nand NAND2_29974 ( P1_R2099_U235 , P1_U4190 , P1_R2099_U116 );
nand NAND2_29975 ( P1_R2099_U236 , P1_U2685 , P1_R2099_U4 );
not NOT1_29976 ( P1_R2099_U237 , P1_R2099_U48 );
nand NAND2_29977 ( P1_R2099_U238 , P1_U4190 , P1_R2099_U117 );
nand NAND2_29978 ( P1_R2099_U239 , P1_U2686 , P1_R2099_U4 );
not NOT1_29979 ( P1_R2099_U240 , P1_R2099_U49 );
nand NAND2_29980 ( P1_R2099_U241 , P1_U4190 , P1_R2099_U118 );
nand NAND2_29981 ( P1_R2099_U242 , P1_U2687 , P1_R2099_U4 );
not NOT1_29982 ( P1_R2099_U243 , P1_R2099_U50 );
nand NAND2_29983 ( P1_R2099_U244 , P1_U4190 , P1_R2099_U119 );
nand NAND2_29984 ( P1_R2099_U245 , P1_U2688 , P1_R2099_U4 );
not NOT1_29985 ( P1_R2099_U246 , P1_R2099_U51 );
nand NAND2_29986 ( P1_R2099_U247 , P1_U4190 , P1_R2099_U120 );
nand NAND2_29987 ( P1_R2099_U248 , P1_U2689 , P1_R2099_U4 );
not NOT1_29988 ( P1_R2099_U249 , P1_R2099_U52 );
nand NAND2_29989 ( P1_R2099_U250 , P1_U4190 , P1_R2099_U121 );
nand NAND2_29990 ( P1_R2099_U251 , P1_U2690 , P1_R2099_U4 );
not NOT1_29991 ( P1_R2099_U252 , P1_R2099_U53 );
nand NAND2_29992 ( P1_R2099_U253 , P1_U4190 , P1_R2099_U122 );
nand NAND2_29993 ( P1_R2099_U254 , P1_U2691 , P1_R2099_U4 );
not NOT1_29994 ( P1_R2099_U255 , P1_R2099_U54 );
nand NAND2_29995 ( P1_R2099_U256 , P1_U4190 , P1_R2099_U123 );
nand NAND2_29996 ( P1_R2099_U257 , P1_U2692 , P1_R2099_U4 );
not NOT1_29997 ( P1_R2099_U258 , P1_R2099_U55 );
nand NAND2_29998 ( P1_R2099_U259 , P1_U4190 , P1_R2099_U124 );
nand NAND2_29999 ( P1_R2099_U260 , P1_U2700 , P1_R2099_U4 );
not NOT1_30000 ( P1_R2099_U261 , P1_R2099_U62 );
nand NAND2_30001 ( P1_R2099_U262 , P1_U4190 , P1_R2099_U125 );
nand NAND2_30002 ( P1_R2099_U263 , P1_U2699 , P1_R2099_U4 );
not NOT1_30003 ( P1_R2099_U264 , P1_R2099_U63 );
nand NAND2_30004 ( P1_R2099_U265 , P1_U4190 , P1_R2099_U126 );
nand NAND2_30005 ( P1_R2099_U266 , P1_U2698 , P1_R2099_U4 );
not NOT1_30006 ( P1_R2099_U267 , P1_R2099_U60 );
nand NAND2_30007 ( P1_R2099_U268 , P1_U4190 , P1_R2099_U127 );
nand NAND2_30008 ( P1_R2099_U269 , P1_U2697 , P1_R2099_U4 );
not NOT1_30009 ( P1_R2099_U270 , P1_R2099_U61 );
nand NAND2_30010 ( P1_R2099_U271 , P1_U4190 , P1_R2099_U128 );
nand NAND2_30011 ( P1_R2099_U272 , P1_U2696 , P1_R2099_U4 );
not NOT1_30012 ( P1_R2099_U273 , P1_R2099_U58 );
nand NAND2_30013 ( P1_R2099_U274 , P1_U4190 , P1_R2099_U129 );
nand NAND2_30014 ( P1_R2099_U275 , P1_U2695 , P1_R2099_U4 );
not NOT1_30015 ( P1_R2099_U276 , P1_R2099_U59 );
nand NAND2_30016 ( P1_R2099_U277 , P1_U4190 , P1_R2099_U130 );
nand NAND2_30017 ( P1_R2099_U278 , P1_U2694 , P1_R2099_U4 );
not NOT1_30018 ( P1_R2099_U279 , P1_R2099_U56 );
nand NAND2_30019 ( P1_R2099_U280 , P1_U4190 , P1_R2099_U131 );
nand NAND2_30020 ( P1_R2099_U281 , P1_U2693 , P1_R2099_U4 );
not NOT1_30021 ( P1_R2099_U282 , P1_R2099_U57 );
nand NAND2_30022 ( P1_R2099_U283 , P1_U4190 , P1_R2099_U132 );
nand NAND2_30023 ( P1_R2099_U284 , P1_U2680 , P1_R2099_U4 );
not NOT1_30024 ( P1_R2099_U285 , P1_R2099_U43 );
nand NAND2_30025 ( P1_R2099_U286 , P1_U4190 , P1_R2099_U133 );
nand NAND2_30026 ( P1_R2099_U287 , P1_U2681 , P1_R2099_U4 );
not NOT1_30027 ( P1_R2099_U288 , P1_R2099_U44 );
nand NAND2_30028 ( P1_R2099_U289 , P1_U4190 , P1_R2099_U134 );
nand NAND2_30029 ( P1_R2099_U290 , P1_U2679 , P1_R2099_U4 );
not NOT1_30030 ( P1_R2099_U291 , P1_R2099_U97 );
nand NAND2_30031 ( P1_R2099_U292 , P1_R2099_U145 , P1_R2099_U291 );
nand NAND2_30032 ( P1_R2099_U293 , P1_R2099_U97 , P1_R2099_U135 );
nand NAND2_30033 ( P1_R2099_U294 , P1_R2099_U181 , P1_R2099_U285 );
nand NAND2_30034 ( P1_R2099_U295 , P1_R2099_U43 , P1_R2099_U136 );
nand NAND2_30035 ( P1_R2099_U296 , P1_R2099_U153 , P1_R2099_U193 );
nand NAND2_30036 ( P1_R2099_U297 , P1_R2099_U35 , P1_R2099_U137 );
nand NAND2_30037 ( P1_R2099_U298 , P1_R2099_U288 , P1_R2099_U180 );
nand NAND2_30038 ( P1_R2099_U299 , P1_R2099_U44 , P1_R2099_U25 );
nand NAND2_30039 ( P1_R2099_U300 , P1_R2099_U228 , P1_R2099_U179 );
nand NAND2_30040 ( P1_R2099_U301 , P1_R2099_U45 , P1_R2099_U24 );
nand NAND2_30041 ( P1_R2099_U302 , P1_R2099_U231 , P1_R2099_U178 );
nand NAND2_30042 ( P1_R2099_U303 , P1_R2099_U46 , P1_R2099_U23 );
nand NAND2_30043 ( P1_R2099_U304 , P1_R2099_U234 , P1_R2099_U177 );
nand NAND2_30044 ( P1_R2099_U305 , P1_R2099_U47 , P1_R2099_U22 );
nand NAND2_30045 ( P1_R2099_U306 , P1_R2099_U237 , P1_R2099_U176 );
nand NAND2_30046 ( P1_R2099_U307 , P1_R2099_U48 , P1_R2099_U21 );
nand NAND2_30047 ( P1_R2099_U308 , P1_R2099_U240 , P1_R2099_U175 );
nand NAND2_30048 ( P1_R2099_U309 , P1_R2099_U49 , P1_R2099_U20 );
nand NAND2_30049 ( P1_R2099_U310 , P1_R2099_U243 , P1_R2099_U174 );
nand NAND2_30050 ( P1_R2099_U311 , P1_R2099_U50 , P1_R2099_U19 );
nand NAND2_30051 ( P1_R2099_U312 , P1_R2099_U246 , P1_R2099_U173 );
nand NAND2_30052 ( P1_R2099_U313 , P1_R2099_U51 , P1_R2099_U18 );
nand NAND2_30053 ( P1_R2099_U314 , P1_R2099_U249 , P1_R2099_U172 );
nand NAND2_30054 ( P1_R2099_U315 , P1_R2099_U52 , P1_R2099_U17 );
nand NAND2_30055 ( P1_R2099_U316 , P1_R2099_U252 , P1_R2099_U171 );
nand NAND2_30056 ( P1_R2099_U317 , P1_R2099_U53 , P1_R2099_U16 );
nand NAND2_30057 ( P1_R2099_U318 , P1_R2099_U190 , P1_U2678 );
nand NAND2_30058 ( P1_R2099_U319 , P1_R2099_U33 , P1_R2099_U6 );
nand NAND2_30059 ( P1_R2099_U320 , P1_R2099_U190 , P1_U2678 );
nand NAND2_30060 ( P1_R2099_U321 , P1_R2099_U33 , P1_R2099_U6 );
nand NAND2_30061 ( P1_R2099_U322 , P1_R2099_U321 , P1_R2099_U320 );
nand NAND2_30062 ( P1_R2099_U323 , P1_R2099_U139 , P1_R2099_U140 );
nand NAND2_30063 ( P1_R2099_U324 , P1_R2099_U149 , P1_R2099_U322 );
nand NAND2_30064 ( P1_R2099_U325 , P1_R2099_U255 , P1_R2099_U170 );
nand NAND2_30065 ( P1_R2099_U326 , P1_R2099_U54 , P1_R2099_U15 );
nand NAND2_30066 ( P1_R2099_U327 , P1_R2099_U258 , P1_R2099_U169 );
nand NAND2_30067 ( P1_R2099_U328 , P1_R2099_U55 , P1_R2099_U14 );
nand NAND2_30068 ( P1_R2099_U329 , P1_R2099_U168 , P1_R2099_U282 );
nand NAND2_30069 ( P1_R2099_U330 , P1_R2099_U57 , P1_R2099_U141 );
nand NAND2_30070 ( P1_R2099_U331 , P1_R2099_U279 , P1_R2099_U167 );
nand NAND2_30071 ( P1_R2099_U332 , P1_R2099_U56 , P1_R2099_U13 );
nand NAND2_30072 ( P1_R2099_U333 , P1_R2099_U166 , P1_R2099_U276 );
nand NAND2_30073 ( P1_R2099_U334 , P1_R2099_U59 , P1_R2099_U142 );
nand NAND2_30074 ( P1_R2099_U335 , P1_R2099_U273 , P1_R2099_U165 );
nand NAND2_30075 ( P1_R2099_U336 , P1_R2099_U58 , P1_R2099_U12 );
nand NAND2_30076 ( P1_R2099_U337 , P1_R2099_U164 , P1_R2099_U270 );
nand NAND2_30077 ( P1_R2099_U338 , P1_R2099_U61 , P1_R2099_U143 );
nand NAND2_30078 ( P1_R2099_U339 , P1_R2099_U267 , P1_R2099_U163 );
nand NAND2_30079 ( P1_R2099_U340 , P1_R2099_U60 , P1_R2099_U11 );
nand NAND2_30080 ( P1_R2099_U341 , P1_R2099_U162 , P1_R2099_U264 );
nand NAND2_30081 ( P1_R2099_U342 , P1_R2099_U63 , P1_R2099_U144 );
nand NAND2_30082 ( P1_R2099_U343 , P1_R2099_U261 , P1_R2099_U161 );
nand NAND2_30083 ( P1_R2099_U344 , P1_R2099_U62 , P1_R2099_U10 );
nand NAND2_30084 ( P1_R2099_U345 , P1_U4189 , P1_R2099_U4 );
nand NAND2_30085 ( P1_R2099_U346 , P1_U4190 , P1_R2099_U5 );
not NOT1_30086 ( P1_R2099_U347 , P1_R2099_U98 );
nand NAND2_30087 ( P1_R2099_U348 , P1_R2099_U32 , P1_R2099_U347 );
nand NAND2_30088 ( P1_R2099_U349 , P1_R2099_U98 , P1_R2099_U187 );
not NOT1_30089 ( P1_R2167_U6 , P1_U2716 );
not NOT1_30090 ( P1_R2167_U7 , P1_U2714 );
not NOT1_30091 ( P1_R2167_U8 , P1_U2720 );
not NOT1_30092 ( P1_R2167_U9 , P1_U2719 );
not NOT1_30093 ( P1_R2167_U10 , P1_U2713 );
not NOT1_30094 ( P1_R2167_U11 , P1_U2712 );
not NOT1_30095 ( P1_R2167_U12 , P1_U2718 );
not NOT1_30096 ( P1_R2167_U13 , P1_U2717 );
not NOT1_30097 ( P1_R2167_U14 , P1_U2711 );
not NOT1_30098 ( P1_R2167_U15 , P1_U2356 );
not NOT1_30099 ( P1_R2167_U16 , P1_STATE2_REG_0_ );
nand NAND2_30100 ( P1_R2167_U17 , P1_R2167_U50 , P1_R2167_U49 );
and AND2_30101 ( P1_R2167_U18 , P1_R2167_U29 , P1_R2167_U30 );
and AND2_30102 ( P1_R2167_U19 , P1_R2167_U32 , P1_R2167_U33 );
and AND2_30103 ( P1_R2167_U20 , P1_R2167_U35 , P1_R2167_U36 );
and AND2_30104 ( P1_R2167_U21 , P1_R2167_U38 , P1_R2167_U39 );
not NOT1_30105 ( P1_R2167_U22 , P1_U2721 );
not NOT1_30106 ( P1_R2167_U23 , P1_U2722 );
nand NAND2_30107 ( P1_R2167_U24 , P1_U2715 , P1_R2167_U23 );
nand NAND2_30108 ( P1_R2167_U25 , P1_U2715 , P1_R2167_U22 );
or OR2_30109 ( P1_R2167_U26 , P1_U2721 , P1_U2722 );
nand NAND2_30110 ( P1_R2167_U27 , P1_U2714 , P1_R2167_U8 );
nand NAND4_30111 ( P1_R2167_U28 , P1_R2167_U27 , P1_R2167_U26 , P1_R2167_U25 , P1_R2167_U24 );
nand NAND2_30112 ( P1_R2167_U29 , P1_U2720 , P1_R2167_U7 );
nand NAND2_30113 ( P1_R2167_U30 , P1_U2719 , P1_R2167_U10 );
nand NAND2_30114 ( P1_R2167_U31 , P1_R2167_U18 , P1_R2167_U28 );
nand NAND2_30115 ( P1_R2167_U32 , P1_U2713 , P1_R2167_U9 );
nand NAND2_30116 ( P1_R2167_U33 , P1_U2712 , P1_R2167_U12 );
nand NAND2_30117 ( P1_R2167_U34 , P1_R2167_U19 , P1_R2167_U31 );
nand NAND2_30118 ( P1_R2167_U35 , P1_U2718 , P1_R2167_U11 );
nand NAND2_30119 ( P1_R2167_U36 , P1_U2717 , P1_R2167_U14 );
nand NAND2_30120 ( P1_R2167_U37 , P1_R2167_U20 , P1_R2167_U34 );
nand NAND2_30121 ( P1_R2167_U38 , P1_U2711 , P1_R2167_U13 );
nand NAND2_30122 ( P1_R2167_U39 , P1_U2356 , P1_R2167_U6 );
nand NAND2_30123 ( P1_R2167_U40 , P1_R2167_U21 , P1_R2167_U37 );
nand NAND2_30124 ( P1_R2167_U41 , P1_U2716 , P1_R2167_U15 );
nand NAND2_30125 ( P1_R2167_U42 , P1_R2167_U40 , P1_R2167_U41 );
nand NAND2_30126 ( P1_R2167_U43 , P1_U2716 , P1_R2167_U16 );
nand NAND2_30127 ( P1_R2167_U44 , P1_R2167_U42 , P1_R2167_U6 );
nand NAND2_30128 ( P1_R2167_U45 , P1_R2167_U44 , P1_R2167_U43 );
nand NAND2_30129 ( P1_R2167_U46 , P1_STATE2_REG_0_ , P1_R2167_U6 );
nand NAND2_30130 ( P1_R2167_U47 , P1_U2716 , P1_R2167_U42 );
nand NAND2_30131 ( P1_R2167_U48 , P1_R2167_U47 , P1_R2167_U46 );
nand NAND2_30132 ( P1_R2167_U49 , P1_R2167_U45 , P1_R2167_U15 );
nand NAND2_30133 ( P1_R2167_U50 , P1_U2356 , P1_R2167_U48 );
not NOT1_30134 ( P1_R2337_U4 , P1_PHYADDRPOINTER_REG_1_ );
not NOT1_30135 ( P1_R2337_U5 , P1_PHYADDRPOINTER_REG_2_ );
nand NAND2_30136 ( P1_R2337_U6 , P1_PHYADDRPOINTER_REG_2_ , P1_PHYADDRPOINTER_REG_1_ );
not NOT1_30137 ( P1_R2337_U7 , P1_PHYADDRPOINTER_REG_3_ );
nand NAND2_30138 ( P1_R2337_U8 , P1_PHYADDRPOINTER_REG_3_ , P1_R2337_U94 );
not NOT1_30139 ( P1_R2337_U9 , P1_PHYADDRPOINTER_REG_4_ );
nand NAND2_30140 ( P1_R2337_U10 , P1_PHYADDRPOINTER_REG_4_ , P1_R2337_U95 );
not NOT1_30141 ( P1_R2337_U11 , P1_PHYADDRPOINTER_REG_5_ );
nand NAND2_30142 ( P1_R2337_U12 , P1_PHYADDRPOINTER_REG_5_ , P1_R2337_U96 );
not NOT1_30143 ( P1_R2337_U13 , P1_PHYADDRPOINTER_REG_6_ );
nand NAND2_30144 ( P1_R2337_U14 , P1_PHYADDRPOINTER_REG_6_ , P1_R2337_U97 );
not NOT1_30145 ( P1_R2337_U15 , P1_PHYADDRPOINTER_REG_7_ );
nand NAND2_30146 ( P1_R2337_U16 , P1_PHYADDRPOINTER_REG_7_ , P1_R2337_U98 );
not NOT1_30147 ( P1_R2337_U17 , P1_PHYADDRPOINTER_REG_8_ );
not NOT1_30148 ( P1_R2337_U18 , P1_PHYADDRPOINTER_REG_9_ );
nand NAND2_30149 ( P1_R2337_U19 , P1_PHYADDRPOINTER_REG_8_ , P1_R2337_U99 );
nand NAND2_30150 ( P1_R2337_U20 , P1_R2337_U100 , P1_PHYADDRPOINTER_REG_9_ );
not NOT1_30151 ( P1_R2337_U21 , P1_PHYADDRPOINTER_REG_10_ );
nand NAND2_30152 ( P1_R2337_U22 , P1_PHYADDRPOINTER_REG_10_ , P1_R2337_U101 );
not NOT1_30153 ( P1_R2337_U23 , P1_PHYADDRPOINTER_REG_11_ );
nand NAND2_30154 ( P1_R2337_U24 , P1_PHYADDRPOINTER_REG_11_ , P1_R2337_U102 );
not NOT1_30155 ( P1_R2337_U25 , P1_PHYADDRPOINTER_REG_12_ );
nand NAND2_30156 ( P1_R2337_U26 , P1_PHYADDRPOINTER_REG_12_ , P1_R2337_U103 );
not NOT1_30157 ( P1_R2337_U27 , P1_PHYADDRPOINTER_REG_13_ );
nand NAND2_30158 ( P1_R2337_U28 , P1_PHYADDRPOINTER_REG_13_ , P1_R2337_U104 );
not NOT1_30159 ( P1_R2337_U29 , P1_PHYADDRPOINTER_REG_14_ );
nand NAND2_30160 ( P1_R2337_U30 , P1_PHYADDRPOINTER_REG_14_ , P1_R2337_U105 );
not NOT1_30161 ( P1_R2337_U31 , P1_PHYADDRPOINTER_REG_15_ );
nand NAND2_30162 ( P1_R2337_U32 , P1_PHYADDRPOINTER_REG_15_ , P1_R2337_U106 );
not NOT1_30163 ( P1_R2337_U33 , P1_PHYADDRPOINTER_REG_16_ );
nand NAND2_30164 ( P1_R2337_U34 , P1_PHYADDRPOINTER_REG_16_ , P1_R2337_U107 );
not NOT1_30165 ( P1_R2337_U35 , P1_PHYADDRPOINTER_REG_17_ );
nand NAND2_30166 ( P1_R2337_U36 , P1_PHYADDRPOINTER_REG_17_ , P1_R2337_U108 );
not NOT1_30167 ( P1_R2337_U37 , P1_PHYADDRPOINTER_REG_18_ );
nand NAND2_30168 ( P1_R2337_U38 , P1_PHYADDRPOINTER_REG_18_ , P1_R2337_U109 );
not NOT1_30169 ( P1_R2337_U39 , P1_PHYADDRPOINTER_REG_19_ );
nand NAND2_30170 ( P1_R2337_U40 , P1_PHYADDRPOINTER_REG_19_ , P1_R2337_U110 );
not NOT1_30171 ( P1_R2337_U41 , P1_PHYADDRPOINTER_REG_20_ );
nand NAND2_30172 ( P1_R2337_U42 , P1_PHYADDRPOINTER_REG_20_ , P1_R2337_U111 );
not NOT1_30173 ( P1_R2337_U43 , P1_PHYADDRPOINTER_REG_21_ );
nand NAND2_30174 ( P1_R2337_U44 , P1_PHYADDRPOINTER_REG_21_ , P1_R2337_U112 );
not NOT1_30175 ( P1_R2337_U45 , P1_PHYADDRPOINTER_REG_22_ );
nand NAND2_30176 ( P1_R2337_U46 , P1_PHYADDRPOINTER_REG_22_ , P1_R2337_U113 );
not NOT1_30177 ( P1_R2337_U47 , P1_PHYADDRPOINTER_REG_23_ );
nand NAND2_30178 ( P1_R2337_U48 , P1_PHYADDRPOINTER_REG_23_ , P1_R2337_U114 );
not NOT1_30179 ( P1_R2337_U49 , P1_PHYADDRPOINTER_REG_24_ );
nand NAND2_30180 ( P1_R2337_U50 , P1_PHYADDRPOINTER_REG_24_ , P1_R2337_U115 );
not NOT1_30181 ( P1_R2337_U51 , P1_PHYADDRPOINTER_REG_25_ );
nand NAND2_30182 ( P1_R2337_U52 , P1_PHYADDRPOINTER_REG_25_ , P1_R2337_U116 );
not NOT1_30183 ( P1_R2337_U53 , P1_PHYADDRPOINTER_REG_26_ );
nand NAND2_30184 ( P1_R2337_U54 , P1_PHYADDRPOINTER_REG_26_ , P1_R2337_U117 );
not NOT1_30185 ( P1_R2337_U55 , P1_PHYADDRPOINTER_REG_27_ );
nand NAND2_30186 ( P1_R2337_U56 , P1_PHYADDRPOINTER_REG_27_ , P1_R2337_U118 );
not NOT1_30187 ( P1_R2337_U57 , P1_PHYADDRPOINTER_REG_28_ );
nand NAND2_30188 ( P1_R2337_U58 , P1_PHYADDRPOINTER_REG_28_ , P1_R2337_U119 );
not NOT1_30189 ( P1_R2337_U59 , P1_PHYADDRPOINTER_REG_29_ );
nand NAND2_30190 ( P1_R2337_U60 , P1_PHYADDRPOINTER_REG_29_ , P1_R2337_U120 );
not NOT1_30191 ( P1_R2337_U61 , P1_PHYADDRPOINTER_REG_30_ );
nand NAND2_30192 ( P1_R2337_U62 , P1_R2337_U124 , P1_R2337_U123 );
nand NAND2_30193 ( P1_R2337_U63 , P1_R2337_U126 , P1_R2337_U125 );
nand NAND2_30194 ( P1_R2337_U64 , P1_R2337_U128 , P1_R2337_U127 );
nand NAND2_30195 ( P1_R2337_U65 , P1_R2337_U130 , P1_R2337_U129 );
nand NAND2_30196 ( P1_R2337_U66 , P1_R2337_U132 , P1_R2337_U131 );
nand NAND2_30197 ( P1_R2337_U67 , P1_R2337_U134 , P1_R2337_U133 );
nand NAND2_30198 ( P1_R2337_U68 , P1_R2337_U136 , P1_R2337_U135 );
nand NAND2_30199 ( P1_R2337_U69 , P1_R2337_U138 , P1_R2337_U137 );
nand NAND2_30200 ( P1_R2337_U70 , P1_R2337_U140 , P1_R2337_U139 );
nand NAND2_30201 ( P1_R2337_U71 , P1_R2337_U142 , P1_R2337_U141 );
nand NAND2_30202 ( P1_R2337_U72 , P1_R2337_U144 , P1_R2337_U143 );
nand NAND2_30203 ( P1_R2337_U73 , P1_R2337_U146 , P1_R2337_U145 );
nand NAND2_30204 ( P1_R2337_U74 , P1_R2337_U148 , P1_R2337_U147 );
nand NAND2_30205 ( P1_R2337_U75 , P1_R2337_U150 , P1_R2337_U149 );
nand NAND2_30206 ( P1_R2337_U76 , P1_R2337_U152 , P1_R2337_U151 );
nand NAND2_30207 ( P1_R2337_U77 , P1_R2337_U154 , P1_R2337_U153 );
nand NAND2_30208 ( P1_R2337_U78 , P1_R2337_U156 , P1_R2337_U155 );
nand NAND2_30209 ( P1_R2337_U79 , P1_R2337_U158 , P1_R2337_U157 );
nand NAND2_30210 ( P1_R2337_U80 , P1_R2337_U160 , P1_R2337_U159 );
nand NAND2_30211 ( P1_R2337_U81 , P1_R2337_U162 , P1_R2337_U161 );
nand NAND2_30212 ( P1_R2337_U82 , P1_R2337_U164 , P1_R2337_U163 );
nand NAND2_30213 ( P1_R2337_U83 , P1_R2337_U166 , P1_R2337_U165 );
nand NAND2_30214 ( P1_R2337_U84 , P1_R2337_U168 , P1_R2337_U167 );
nand NAND2_30215 ( P1_R2337_U85 , P1_R2337_U170 , P1_R2337_U169 );
nand NAND2_30216 ( P1_R2337_U86 , P1_R2337_U172 , P1_R2337_U171 );
nand NAND2_30217 ( P1_R2337_U87 , P1_R2337_U174 , P1_R2337_U173 );
nand NAND2_30218 ( P1_R2337_U88 , P1_R2337_U176 , P1_R2337_U175 );
nand NAND2_30219 ( P1_R2337_U89 , P1_R2337_U178 , P1_R2337_U177 );
nand NAND2_30220 ( P1_R2337_U90 , P1_R2337_U180 , P1_R2337_U179 );
nand NAND2_30221 ( P1_R2337_U91 , P1_R2337_U182 , P1_R2337_U181 );
not NOT1_30222 ( P1_R2337_U92 , P1_PHYADDRPOINTER_REG_31_ );
nand NAND2_30223 ( P1_R2337_U93 , P1_PHYADDRPOINTER_REG_30_ , P1_R2337_U121 );
not NOT1_30224 ( P1_R2337_U94 , P1_R2337_U6 );
not NOT1_30225 ( P1_R2337_U95 , P1_R2337_U8 );
not NOT1_30226 ( P1_R2337_U96 , P1_R2337_U10 );
not NOT1_30227 ( P1_R2337_U97 , P1_R2337_U12 );
not NOT1_30228 ( P1_R2337_U98 , P1_R2337_U14 );
not NOT1_30229 ( P1_R2337_U99 , P1_R2337_U16 );
not NOT1_30230 ( P1_R2337_U100 , P1_R2337_U19 );
not NOT1_30231 ( P1_R2337_U101 , P1_R2337_U20 );
not NOT1_30232 ( P1_R2337_U102 , P1_R2337_U22 );
not NOT1_30233 ( P1_R2337_U103 , P1_R2337_U24 );
not NOT1_30234 ( P1_R2337_U104 , P1_R2337_U26 );
not NOT1_30235 ( P1_R2337_U105 , P1_R2337_U28 );
not NOT1_30236 ( P1_R2337_U106 , P1_R2337_U30 );
not NOT1_30237 ( P1_R2337_U107 , P1_R2337_U32 );
not NOT1_30238 ( P1_R2337_U108 , P1_R2337_U34 );
not NOT1_30239 ( P1_R2337_U109 , P1_R2337_U36 );
not NOT1_30240 ( P1_R2337_U110 , P1_R2337_U38 );
not NOT1_30241 ( P1_R2337_U111 , P1_R2337_U40 );
not NOT1_30242 ( P1_R2337_U112 , P1_R2337_U42 );
not NOT1_30243 ( P1_R2337_U113 , P1_R2337_U44 );
not NOT1_30244 ( P1_R2337_U114 , P1_R2337_U46 );
not NOT1_30245 ( P1_R2337_U115 , P1_R2337_U48 );
not NOT1_30246 ( P1_R2337_U116 , P1_R2337_U50 );
not NOT1_30247 ( P1_R2337_U117 , P1_R2337_U52 );
not NOT1_30248 ( P1_R2337_U118 , P1_R2337_U54 );
not NOT1_30249 ( P1_R2337_U119 , P1_R2337_U56 );
not NOT1_30250 ( P1_R2337_U120 , P1_R2337_U58 );
not NOT1_30251 ( P1_R2337_U121 , P1_R2337_U60 );
not NOT1_30252 ( P1_R2337_U122 , P1_R2337_U93 );
nand NAND2_30253 ( P1_R2337_U123 , P1_PHYADDRPOINTER_REG_9_ , P1_R2337_U19 );
nand NAND2_30254 ( P1_R2337_U124 , P1_R2337_U100 , P1_R2337_U18 );
nand NAND2_30255 ( P1_R2337_U125 , P1_PHYADDRPOINTER_REG_8_ , P1_R2337_U16 );
nand NAND2_30256 ( P1_R2337_U126 , P1_R2337_U99 , P1_R2337_U17 );
nand NAND2_30257 ( P1_R2337_U127 , P1_PHYADDRPOINTER_REG_7_ , P1_R2337_U14 );
nand NAND2_30258 ( P1_R2337_U128 , P1_R2337_U98 , P1_R2337_U15 );
nand NAND2_30259 ( P1_R2337_U129 , P1_PHYADDRPOINTER_REG_6_ , P1_R2337_U12 );
nand NAND2_30260 ( P1_R2337_U130 , P1_R2337_U97 , P1_R2337_U13 );
nand NAND2_30261 ( P1_R2337_U131 , P1_PHYADDRPOINTER_REG_5_ , P1_R2337_U10 );
nand NAND2_30262 ( P1_R2337_U132 , P1_R2337_U96 , P1_R2337_U11 );
nand NAND2_30263 ( P1_R2337_U133 , P1_PHYADDRPOINTER_REG_4_ , P1_R2337_U8 );
nand NAND2_30264 ( P1_R2337_U134 , P1_R2337_U95 , P1_R2337_U9 );
nand NAND2_30265 ( P1_R2337_U135 , P1_PHYADDRPOINTER_REG_3_ , P1_R2337_U6 );
nand NAND2_30266 ( P1_R2337_U136 , P1_R2337_U94 , P1_R2337_U7 );
nand NAND2_30267 ( P1_R2337_U137 , P1_PHYADDRPOINTER_REG_31_ , P1_R2337_U93 );
nand NAND2_30268 ( P1_R2337_U138 , P1_R2337_U122 , P1_R2337_U92 );
nand NAND2_30269 ( P1_R2337_U139 , P1_PHYADDRPOINTER_REG_30_ , P1_R2337_U60 );
nand NAND2_30270 ( P1_R2337_U140 , P1_R2337_U121 , P1_R2337_U61 );
nand NAND2_30271 ( P1_R2337_U141 , P1_PHYADDRPOINTER_REG_2_ , P1_R2337_U4 );
nand NAND2_30272 ( P1_R2337_U142 , P1_PHYADDRPOINTER_REG_1_ , P1_R2337_U5 );
nand NAND2_30273 ( P1_R2337_U143 , P1_PHYADDRPOINTER_REG_29_ , P1_R2337_U58 );
nand NAND2_30274 ( P1_R2337_U144 , P1_R2337_U120 , P1_R2337_U59 );
nand NAND2_30275 ( P1_R2337_U145 , P1_PHYADDRPOINTER_REG_28_ , P1_R2337_U56 );
nand NAND2_30276 ( P1_R2337_U146 , P1_R2337_U119 , P1_R2337_U57 );
nand NAND2_30277 ( P1_R2337_U147 , P1_PHYADDRPOINTER_REG_27_ , P1_R2337_U54 );
nand NAND2_30278 ( P1_R2337_U148 , P1_R2337_U118 , P1_R2337_U55 );
nand NAND2_30279 ( P1_R2337_U149 , P1_PHYADDRPOINTER_REG_26_ , P1_R2337_U52 );
nand NAND2_30280 ( P1_R2337_U150 , P1_R2337_U117 , P1_R2337_U53 );
nand NAND2_30281 ( P1_R2337_U151 , P1_PHYADDRPOINTER_REG_25_ , P1_R2337_U50 );
nand NAND2_30282 ( P1_R2337_U152 , P1_R2337_U116 , P1_R2337_U51 );
nand NAND2_30283 ( P1_R2337_U153 , P1_PHYADDRPOINTER_REG_24_ , P1_R2337_U48 );
nand NAND2_30284 ( P1_R2337_U154 , P1_R2337_U115 , P1_R2337_U49 );
nand NAND2_30285 ( P1_R2337_U155 , P1_PHYADDRPOINTER_REG_23_ , P1_R2337_U46 );
nand NAND2_30286 ( P1_R2337_U156 , P1_R2337_U114 , P1_R2337_U47 );
nand NAND2_30287 ( P1_R2337_U157 , P1_PHYADDRPOINTER_REG_22_ , P1_R2337_U44 );
nand NAND2_30288 ( P1_R2337_U158 , P1_R2337_U113 , P1_R2337_U45 );
nand NAND2_30289 ( P1_R2337_U159 , P1_PHYADDRPOINTER_REG_21_ , P1_R2337_U42 );
nand NAND2_30290 ( P1_R2337_U160 , P1_R2337_U112 , P1_R2337_U43 );
nand NAND2_30291 ( P1_R2337_U161 , P1_PHYADDRPOINTER_REG_20_ , P1_R2337_U40 );
nand NAND2_30292 ( P1_R2337_U162 , P1_R2337_U111 , P1_R2337_U41 );
nand NAND2_30293 ( P1_R2337_U163 , P1_PHYADDRPOINTER_REG_19_ , P1_R2337_U38 );
nand NAND2_30294 ( P1_R2337_U164 , P1_R2337_U110 , P1_R2337_U39 );
nand NAND2_30295 ( P1_R2337_U165 , P1_PHYADDRPOINTER_REG_18_ , P1_R2337_U36 );
nand NAND2_30296 ( P1_R2337_U166 , P1_R2337_U109 , P1_R2337_U37 );
nand NAND2_30297 ( P1_R2337_U167 , P1_PHYADDRPOINTER_REG_17_ , P1_R2337_U34 );
nand NAND2_30298 ( P1_R2337_U168 , P1_R2337_U108 , P1_R2337_U35 );
nand NAND2_30299 ( P1_R2337_U169 , P1_PHYADDRPOINTER_REG_16_ , P1_R2337_U32 );
nand NAND2_30300 ( P1_R2337_U170 , P1_R2337_U107 , P1_R2337_U33 );
nand NAND2_30301 ( P1_R2337_U171 , P1_PHYADDRPOINTER_REG_15_ , P1_R2337_U30 );
nand NAND2_30302 ( P1_R2337_U172 , P1_R2337_U106 , P1_R2337_U31 );
nand NAND2_30303 ( P1_R2337_U173 , P1_PHYADDRPOINTER_REG_14_ , P1_R2337_U28 );
nand NAND2_30304 ( P1_R2337_U174 , P1_R2337_U105 , P1_R2337_U29 );
nand NAND2_30305 ( P1_R2337_U175 , P1_PHYADDRPOINTER_REG_13_ , P1_R2337_U26 );
nand NAND2_30306 ( P1_R2337_U176 , P1_R2337_U104 , P1_R2337_U27 );
nand NAND2_30307 ( P1_R2337_U177 , P1_PHYADDRPOINTER_REG_12_ , P1_R2337_U24 );
nand NAND2_30308 ( P1_R2337_U178 , P1_R2337_U103 , P1_R2337_U25 );
nand NAND2_30309 ( P1_R2337_U179 , P1_PHYADDRPOINTER_REG_11_ , P1_R2337_U22 );
nand NAND2_30310 ( P1_R2337_U180 , P1_R2337_U102 , P1_R2337_U23 );
nand NAND2_30311 ( P1_R2337_U181 , P1_PHYADDRPOINTER_REG_10_ , P1_R2337_U20 );
nand NAND2_30312 ( P1_R2337_U182 , P1_R2337_U101 , P1_R2337_U21 );
not NOT1_30313 ( P1_SUB_357_U6 , P1_U3233 );
not NOT1_30314 ( P1_SUB_357_U7 , P1_U3228 );
not NOT1_30315 ( P1_SUB_357_U8 , P1_U3234 );
not NOT1_30316 ( P1_SUB_357_U9 , P1_U3232 );
not NOT1_30317 ( P1_SUB_357_U10 , P1_U3227 );
not NOT1_30318 ( P1_SUB_357_U11 , P1_U3230 );
not NOT1_30319 ( P1_SUB_357_U12 , P1_U3229 );
not NOT1_30320 ( P1_SUB_357_U13 , P1_U3231 );
and AND2_30321 ( P1_LT_563_1260_U6 , P1_LT_563_1260_U9 , P1_LT_563_1260_U8 );
not NOT1_30322 ( P1_LT_563_1260_U7 , P1_U2673 );
nand NAND2_30323 ( P1_LT_563_1260_U8 , P1_R584_U8 , P1_LT_563_1260_U7 );
nand NAND2_30324 ( P1_LT_563_1260_U9 , P1_R584_U9 , P1_LT_563_1260_U7 );
nand NAND2_30325 ( P1_SUB_580_U6 , P1_SUB_580_U10 , P1_SUB_580_U9 );
not NOT1_30326 ( P1_SUB_580_U7 , P1_INSTADDRPOINTER_REG_1_ );
not NOT1_30327 ( P1_SUB_580_U8 , P1_INSTADDRPOINTER_REG_0_ );
nand NAND2_30328 ( P1_SUB_580_U9 , P1_INSTADDRPOINTER_REG_1_ , P1_SUB_580_U8 );
nand NAND2_30329 ( P1_SUB_580_U10 , P1_INSTADDRPOINTER_REG_0_ , P1_SUB_580_U7 );
not NOT1_30330 ( P1_R2096_U4 , P1_REIP_REG_1_ );
not NOT1_30331 ( P1_R2096_U5 , P1_REIP_REG_2_ );
nand NAND2_30332 ( P1_R2096_U6 , P1_REIP_REG_2_ , P1_REIP_REG_1_ );
not NOT1_30333 ( P1_R2096_U7 , P1_REIP_REG_3_ );
nand NAND2_30334 ( P1_R2096_U8 , P1_REIP_REG_3_ , P1_R2096_U94 );
not NOT1_30335 ( P1_R2096_U9 , P1_REIP_REG_4_ );
nand NAND2_30336 ( P1_R2096_U10 , P1_REIP_REG_4_ , P1_R2096_U95 );
not NOT1_30337 ( P1_R2096_U11 , P1_REIP_REG_5_ );
nand NAND2_30338 ( P1_R2096_U12 , P1_REIP_REG_5_ , P1_R2096_U96 );
not NOT1_30339 ( P1_R2096_U13 , P1_REIP_REG_6_ );
nand NAND2_30340 ( P1_R2096_U14 , P1_REIP_REG_6_ , P1_R2096_U97 );
not NOT1_30341 ( P1_R2096_U15 , P1_REIP_REG_7_ );
nand NAND2_30342 ( P1_R2096_U16 , P1_REIP_REG_7_ , P1_R2096_U98 );
not NOT1_30343 ( P1_R2096_U17 , P1_REIP_REG_8_ );
not NOT1_30344 ( P1_R2096_U18 , P1_REIP_REG_9_ );
nand NAND2_30345 ( P1_R2096_U19 , P1_REIP_REG_8_ , P1_R2096_U99 );
nand NAND2_30346 ( P1_R2096_U20 , P1_R2096_U100 , P1_REIP_REG_9_ );
not NOT1_30347 ( P1_R2096_U21 , P1_REIP_REG_10_ );
nand NAND2_30348 ( P1_R2096_U22 , P1_REIP_REG_10_ , P1_R2096_U101 );
not NOT1_30349 ( P1_R2096_U23 , P1_REIP_REG_11_ );
nand NAND2_30350 ( P1_R2096_U24 , P1_REIP_REG_11_ , P1_R2096_U102 );
not NOT1_30351 ( P1_R2096_U25 , P1_REIP_REG_12_ );
nand NAND2_30352 ( P1_R2096_U26 , P1_REIP_REG_12_ , P1_R2096_U103 );
not NOT1_30353 ( P1_R2096_U27 , P1_REIP_REG_13_ );
nand NAND2_30354 ( P1_R2096_U28 , P1_REIP_REG_13_ , P1_R2096_U104 );
not NOT1_30355 ( P1_R2096_U29 , P1_REIP_REG_14_ );
nand NAND2_30356 ( P1_R2096_U30 , P1_REIP_REG_14_ , P1_R2096_U105 );
not NOT1_30357 ( P1_R2096_U31 , P1_REIP_REG_15_ );
nand NAND2_30358 ( P1_R2096_U32 , P1_REIP_REG_15_ , P1_R2096_U106 );
not NOT1_30359 ( P1_R2096_U33 , P1_REIP_REG_16_ );
nand NAND2_30360 ( P1_R2096_U34 , P1_REIP_REG_16_ , P1_R2096_U107 );
not NOT1_30361 ( P1_R2096_U35 , P1_REIP_REG_17_ );
nand NAND2_30362 ( P1_R2096_U36 , P1_REIP_REG_17_ , P1_R2096_U108 );
not NOT1_30363 ( P1_R2096_U37 , P1_REIP_REG_18_ );
nand NAND2_30364 ( P1_R2096_U38 , P1_REIP_REG_18_ , P1_R2096_U109 );
not NOT1_30365 ( P1_R2096_U39 , P1_REIP_REG_19_ );
nand NAND2_30366 ( P1_R2096_U40 , P1_REIP_REG_19_ , P1_R2096_U110 );
not NOT1_30367 ( P1_R2096_U41 , P1_REIP_REG_20_ );
nand NAND2_30368 ( P1_R2096_U42 , P1_REIP_REG_20_ , P1_R2096_U111 );
not NOT1_30369 ( P1_R2096_U43 , P1_REIP_REG_21_ );
nand NAND2_30370 ( P1_R2096_U44 , P1_REIP_REG_21_ , P1_R2096_U112 );
not NOT1_30371 ( P1_R2096_U45 , P1_REIP_REG_22_ );
nand NAND2_30372 ( P1_R2096_U46 , P1_REIP_REG_22_ , P1_R2096_U113 );
not NOT1_30373 ( P1_R2096_U47 , P1_REIP_REG_23_ );
nand NAND2_30374 ( P1_R2096_U48 , P1_REIP_REG_23_ , P1_R2096_U114 );
not NOT1_30375 ( P1_R2096_U49 , P1_REIP_REG_24_ );
nand NAND2_30376 ( P1_R2096_U50 , P1_REIP_REG_24_ , P1_R2096_U115 );
not NOT1_30377 ( P1_R2096_U51 , P1_REIP_REG_25_ );
nand NAND2_30378 ( P1_R2096_U52 , P1_REIP_REG_25_ , P1_R2096_U116 );
not NOT1_30379 ( P1_R2096_U53 , P1_REIP_REG_26_ );
nand NAND2_30380 ( P1_R2096_U54 , P1_REIP_REG_26_ , P1_R2096_U117 );
not NOT1_30381 ( P1_R2096_U55 , P1_REIP_REG_27_ );
nand NAND2_30382 ( P1_R2096_U56 , P1_REIP_REG_27_ , P1_R2096_U118 );
not NOT1_30383 ( P1_R2096_U57 , P1_REIP_REG_28_ );
nand NAND2_30384 ( P1_R2096_U58 , P1_REIP_REG_28_ , P1_R2096_U119 );
not NOT1_30385 ( P1_R2096_U59 , P1_REIP_REG_29_ );
nand NAND2_30386 ( P1_R2096_U60 , P1_REIP_REG_29_ , P1_R2096_U120 );
not NOT1_30387 ( P1_R2096_U61 , P1_REIP_REG_30_ );
nand NAND2_30388 ( P1_R2096_U62 , P1_R2096_U124 , P1_R2096_U123 );
nand NAND2_30389 ( P1_R2096_U63 , P1_R2096_U126 , P1_R2096_U125 );
nand NAND2_30390 ( P1_R2096_U64 , P1_R2096_U128 , P1_R2096_U127 );
nand NAND2_30391 ( P1_R2096_U65 , P1_R2096_U130 , P1_R2096_U129 );
nand NAND2_30392 ( P1_R2096_U66 , P1_R2096_U132 , P1_R2096_U131 );
nand NAND2_30393 ( P1_R2096_U67 , P1_R2096_U134 , P1_R2096_U133 );
nand NAND2_30394 ( P1_R2096_U68 , P1_R2096_U136 , P1_R2096_U135 );
nand NAND2_30395 ( P1_R2096_U69 , P1_R2096_U138 , P1_R2096_U137 );
nand NAND2_30396 ( P1_R2096_U70 , P1_R2096_U140 , P1_R2096_U139 );
nand NAND2_30397 ( P1_R2096_U71 , P1_R2096_U142 , P1_R2096_U141 );
nand NAND2_30398 ( P1_R2096_U72 , P1_R2096_U144 , P1_R2096_U143 );
nand NAND2_30399 ( P1_R2096_U73 , P1_R2096_U146 , P1_R2096_U145 );
nand NAND2_30400 ( P1_R2096_U74 , P1_R2096_U148 , P1_R2096_U147 );
nand NAND2_30401 ( P1_R2096_U75 , P1_R2096_U150 , P1_R2096_U149 );
nand NAND2_30402 ( P1_R2096_U76 , P1_R2096_U152 , P1_R2096_U151 );
nand NAND2_30403 ( P1_R2096_U77 , P1_R2096_U154 , P1_R2096_U153 );
nand NAND2_30404 ( P1_R2096_U78 , P1_R2096_U156 , P1_R2096_U155 );
nand NAND2_30405 ( P1_R2096_U79 , P1_R2096_U158 , P1_R2096_U157 );
nand NAND2_30406 ( P1_R2096_U80 , P1_R2096_U160 , P1_R2096_U159 );
nand NAND2_30407 ( P1_R2096_U81 , P1_R2096_U162 , P1_R2096_U161 );
nand NAND2_30408 ( P1_R2096_U82 , P1_R2096_U164 , P1_R2096_U163 );
nand NAND2_30409 ( P1_R2096_U83 , P1_R2096_U166 , P1_R2096_U165 );
nand NAND2_30410 ( P1_R2096_U84 , P1_R2096_U168 , P1_R2096_U167 );
nand NAND2_30411 ( P1_R2096_U85 , P1_R2096_U170 , P1_R2096_U169 );
nand NAND2_30412 ( P1_R2096_U86 , P1_R2096_U172 , P1_R2096_U171 );
nand NAND2_30413 ( P1_R2096_U87 , P1_R2096_U174 , P1_R2096_U173 );
nand NAND2_30414 ( P1_R2096_U88 , P1_R2096_U176 , P1_R2096_U175 );
nand NAND2_30415 ( P1_R2096_U89 , P1_R2096_U178 , P1_R2096_U177 );
nand NAND2_30416 ( P1_R2096_U90 , P1_R2096_U180 , P1_R2096_U179 );
nand NAND2_30417 ( P1_R2096_U91 , P1_R2096_U182 , P1_R2096_U181 );
not NOT1_30418 ( P1_R2096_U92 , P1_REIP_REG_31_ );
nand NAND2_30419 ( P1_R2096_U93 , P1_REIP_REG_30_ , P1_R2096_U121 );
not NOT1_30420 ( P1_R2096_U94 , P1_R2096_U6 );
not NOT1_30421 ( P1_R2096_U95 , P1_R2096_U8 );
not NOT1_30422 ( P1_R2096_U96 , P1_R2096_U10 );
not NOT1_30423 ( P1_R2096_U97 , P1_R2096_U12 );
not NOT1_30424 ( P1_R2096_U98 , P1_R2096_U14 );
not NOT1_30425 ( P1_R2096_U99 , P1_R2096_U16 );
not NOT1_30426 ( P1_R2096_U100 , P1_R2096_U19 );
not NOT1_30427 ( P1_R2096_U101 , P1_R2096_U20 );
not NOT1_30428 ( P1_R2096_U102 , P1_R2096_U22 );
not NOT1_30429 ( P1_R2096_U103 , P1_R2096_U24 );
not NOT1_30430 ( P1_R2096_U104 , P1_R2096_U26 );
not NOT1_30431 ( P1_R2096_U105 , P1_R2096_U28 );
not NOT1_30432 ( P1_R2096_U106 , P1_R2096_U30 );
not NOT1_30433 ( P1_R2096_U107 , P1_R2096_U32 );
not NOT1_30434 ( P1_R2096_U108 , P1_R2096_U34 );
not NOT1_30435 ( P1_R2096_U109 , P1_R2096_U36 );
not NOT1_30436 ( P1_R2096_U110 , P1_R2096_U38 );
not NOT1_30437 ( P1_R2096_U111 , P1_R2096_U40 );
not NOT1_30438 ( P1_R2096_U112 , P1_R2096_U42 );
not NOT1_30439 ( P1_R2096_U113 , P1_R2096_U44 );
not NOT1_30440 ( P1_R2096_U114 , P1_R2096_U46 );
not NOT1_30441 ( P1_R2096_U115 , P1_R2096_U48 );
not NOT1_30442 ( P1_R2096_U116 , P1_R2096_U50 );
not NOT1_30443 ( P1_R2096_U117 , P1_R2096_U52 );
not NOT1_30444 ( P1_R2096_U118 , P1_R2096_U54 );
not NOT1_30445 ( P1_R2096_U119 , P1_R2096_U56 );
not NOT1_30446 ( P1_R2096_U120 , P1_R2096_U58 );
not NOT1_30447 ( P1_R2096_U121 , P1_R2096_U60 );
not NOT1_30448 ( P1_R2096_U122 , P1_R2096_U93 );
nand NAND2_30449 ( P1_R2096_U123 , P1_REIP_REG_9_ , P1_R2096_U19 );
nand NAND2_30450 ( P1_R2096_U124 , P1_R2096_U100 , P1_R2096_U18 );
nand NAND2_30451 ( P1_R2096_U125 , P1_REIP_REG_8_ , P1_R2096_U16 );
nand NAND2_30452 ( P1_R2096_U126 , P1_R2096_U99 , P1_R2096_U17 );
nand NAND2_30453 ( P1_R2096_U127 , P1_REIP_REG_7_ , P1_R2096_U14 );
nand NAND2_30454 ( P1_R2096_U128 , P1_R2096_U98 , P1_R2096_U15 );
nand NAND2_30455 ( P1_R2096_U129 , P1_REIP_REG_6_ , P1_R2096_U12 );
nand NAND2_30456 ( P1_R2096_U130 , P1_R2096_U97 , P1_R2096_U13 );
nand NAND2_30457 ( P1_R2096_U131 , P1_REIP_REG_5_ , P1_R2096_U10 );
nand NAND2_30458 ( P1_R2096_U132 , P1_R2096_U96 , P1_R2096_U11 );
nand NAND2_30459 ( P1_R2096_U133 , P1_REIP_REG_4_ , P1_R2096_U8 );
nand NAND2_30460 ( P1_R2096_U134 , P1_R2096_U95 , P1_R2096_U9 );
nand NAND2_30461 ( P1_R2096_U135 , P1_REIP_REG_3_ , P1_R2096_U6 );
nand NAND2_30462 ( P1_R2096_U136 , P1_R2096_U94 , P1_R2096_U7 );
nand NAND2_30463 ( P1_R2096_U137 , P1_REIP_REG_31_ , P1_R2096_U93 );
nand NAND2_30464 ( P1_R2096_U138 , P1_R2096_U122 , P1_R2096_U92 );
nand NAND2_30465 ( P1_R2096_U139 , P1_REIP_REG_30_ , P1_R2096_U60 );
nand NAND2_30466 ( P1_R2096_U140 , P1_R2096_U121 , P1_R2096_U61 );
nand NAND2_30467 ( P1_R2096_U141 , P1_REIP_REG_2_ , P1_R2096_U4 );
nand NAND2_30468 ( P1_R2096_U142 , P1_REIP_REG_1_ , P1_R2096_U5 );
nand NAND2_30469 ( P1_R2096_U143 , P1_REIP_REG_29_ , P1_R2096_U58 );
nand NAND2_30470 ( P1_R2096_U144 , P1_R2096_U120 , P1_R2096_U59 );
nand NAND2_30471 ( P1_R2096_U145 , P1_REIP_REG_28_ , P1_R2096_U56 );
nand NAND2_30472 ( P1_R2096_U146 , P1_R2096_U119 , P1_R2096_U57 );
nand NAND2_30473 ( P1_R2096_U147 , P1_REIP_REG_27_ , P1_R2096_U54 );
nand NAND2_30474 ( P1_R2096_U148 , P1_R2096_U118 , P1_R2096_U55 );
nand NAND2_30475 ( P1_R2096_U149 , P1_REIP_REG_26_ , P1_R2096_U52 );
nand NAND2_30476 ( P1_R2096_U150 , P1_R2096_U117 , P1_R2096_U53 );
nand NAND2_30477 ( P1_R2096_U151 , P1_REIP_REG_25_ , P1_R2096_U50 );
nand NAND2_30478 ( P1_R2096_U152 , P1_R2096_U116 , P1_R2096_U51 );
nand NAND2_30479 ( P1_R2096_U153 , P1_REIP_REG_24_ , P1_R2096_U48 );
nand NAND2_30480 ( P1_R2096_U154 , P1_R2096_U115 , P1_R2096_U49 );
nand NAND2_30481 ( P1_R2096_U155 , P1_REIP_REG_23_ , P1_R2096_U46 );
nand NAND2_30482 ( P1_R2096_U156 , P1_R2096_U114 , P1_R2096_U47 );
nand NAND2_30483 ( P1_R2096_U157 , P1_REIP_REG_22_ , P1_R2096_U44 );
nand NAND2_30484 ( P1_R2096_U158 , P1_R2096_U113 , P1_R2096_U45 );
nand NAND2_30485 ( P1_R2096_U159 , P1_REIP_REG_21_ , P1_R2096_U42 );
nand NAND2_30486 ( P1_R2096_U160 , P1_R2096_U112 , P1_R2096_U43 );
nand NAND2_30487 ( P1_R2096_U161 , P1_REIP_REG_20_ , P1_R2096_U40 );
nand NAND2_30488 ( P1_R2096_U162 , P1_R2096_U111 , P1_R2096_U41 );
nand NAND2_30489 ( P1_R2096_U163 , P1_REIP_REG_19_ , P1_R2096_U38 );
nand NAND2_30490 ( P1_R2096_U164 , P1_R2096_U110 , P1_R2096_U39 );
nand NAND2_30491 ( P1_R2096_U165 , P1_REIP_REG_18_ , P1_R2096_U36 );
nand NAND2_30492 ( P1_R2096_U166 , P1_R2096_U109 , P1_R2096_U37 );
nand NAND2_30493 ( P1_R2096_U167 , P1_REIP_REG_17_ , P1_R2096_U34 );
nand NAND2_30494 ( P1_R2096_U168 , P1_R2096_U108 , P1_R2096_U35 );
nand NAND2_30495 ( P1_R2096_U169 , P1_REIP_REG_16_ , P1_R2096_U32 );
nand NAND2_30496 ( P1_R2096_U170 , P1_R2096_U107 , P1_R2096_U33 );
nand NAND2_30497 ( P1_R2096_U171 , P1_REIP_REG_15_ , P1_R2096_U30 );
nand NAND2_30498 ( P1_R2096_U172 , P1_R2096_U106 , P1_R2096_U31 );
nand NAND2_30499 ( P1_R2096_U173 , P1_REIP_REG_14_ , P1_R2096_U28 );
nand NAND2_30500 ( P1_R2096_U174 , P1_R2096_U105 , P1_R2096_U29 );
nand NAND2_30501 ( P1_R2096_U175 , P1_REIP_REG_13_ , P1_R2096_U26 );
nand NAND2_30502 ( P1_R2096_U176 , P1_R2096_U104 , P1_R2096_U27 );
nand NAND2_30503 ( P1_R2096_U177 , P1_REIP_REG_12_ , P1_R2096_U24 );
nand NAND2_30504 ( P1_R2096_U178 , P1_R2096_U103 , P1_R2096_U25 );
nand NAND2_30505 ( P1_R2096_U179 , P1_REIP_REG_11_ , P1_R2096_U22 );
nand NAND2_30506 ( P1_R2096_U180 , P1_R2096_U102 , P1_R2096_U23 );
nand NAND2_30507 ( P1_R2096_U181 , P1_REIP_REG_10_ , P1_R2096_U20 );
nand NAND2_30508 ( P1_R2096_U182 , P1_R2096_U101 , P1_R2096_U21 );
and AND2_30509 ( P1_LT_563_U6 , P1_LT_563_U27 , P1_LT_563_U26 );
not NOT1_30510 ( P1_LT_563_U7 , P1_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_30511 ( P1_LT_563_U8 , P1_U3491 );
not NOT1_30512 ( P1_LT_563_U9 , P1_U3490 );
not NOT1_30513 ( P1_LT_563_U10 , P1_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_30514 ( P1_LT_563_U11 , P1_INSTQUEUEWR_ADDR_REG_4_ );
not NOT1_30515 ( P1_LT_563_U12 , P1_U3489 );
and AND2_30516 ( P1_LT_563_U13 , P1_LT_563_U21 , P1_LT_563_U22 );
and AND2_30517 ( P1_LT_563_U14 , P1_LT_563_U24 , P1_LT_563_U25 );
not NOT1_30518 ( P1_LT_563_U15 , P1_U3492 );
not NOT1_30519 ( P1_LT_563_U16 , P1_U3493 );
nand NAND3_30520 ( P1_LT_563_U17 , P1_LT_563_U16 , P1_LT_563_U15 , P1_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_30521 ( P1_LT_563_U18 , P1_INSTQUEUEWR_ADDR_REG_1_ , P1_LT_563_U15 );
nand NAND2_30522 ( P1_LT_563_U19 , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_LT_563_U8 );
nand NAND4_30523 ( P1_LT_563_U20 , P1_LT_563_U28 , P1_LT_563_U19 , P1_LT_563_U18 , P1_LT_563_U17 );
nand NAND2_30524 ( P1_LT_563_U21 , P1_U3491 , P1_LT_563_U7 );
nand NAND2_30525 ( P1_LT_563_U22 , P1_U3490 , P1_LT_563_U10 );
nand NAND2_30526 ( P1_LT_563_U23 , P1_LT_563_U13 , P1_LT_563_U20 );
nand NAND2_30527 ( P1_LT_563_U24 , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_LT_563_U9 );
nand NAND2_30528 ( P1_LT_563_U25 , P1_INSTQUEUEWR_ADDR_REG_4_ , P1_LT_563_U12 );
nand NAND2_30529 ( P1_LT_563_U26 , P1_LT_563_U14 , P1_LT_563_U23 );
nand NAND2_30530 ( P1_LT_563_U27 , P1_U3489 , P1_LT_563_U11 );
nand NAND3_30531 ( P1_LT_563_U28 , P1_INSTQUEUEWR_ADDR_REG_0_ , P1_INSTQUEUEWR_ADDR_REG_1_ , P1_LT_563_U16 );
nand NAND2_30532 ( P1_R2238_U6 , P1_R2238_U45 , P1_R2238_U44 );
nand NAND2_30533 ( P1_R2238_U7 , P1_R2238_U9 , P1_R2238_U46 );
not NOT1_30534 ( P1_R2238_U8 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_30535 ( P1_R2238_U9 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_R2238_U18 );
not NOT1_30536 ( P1_R2238_U10 , P1_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_30537 ( P1_R2238_U11 , P1_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_30538 ( P1_R2238_U12 , P1_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_30539 ( P1_R2238_U13 , P1_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_30540 ( P1_R2238_U14 , P1_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_30541 ( P1_R2238_U15 , P1_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_30542 ( P1_R2238_U16 , P1_R2238_U41 , P1_R2238_U40 );
not NOT1_30543 ( P1_R2238_U17 , P1_INSTQUEUERD_ADDR_REG_4_ );
not NOT1_30544 ( P1_R2238_U18 , P1_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_30545 ( P1_R2238_U19 , P1_R2238_U51 , P1_R2238_U50 );
nand NAND2_30546 ( P1_R2238_U20 , P1_R2238_U56 , P1_R2238_U55 );
nand NAND2_30547 ( P1_R2238_U21 , P1_R2238_U61 , P1_R2238_U60 );
nand NAND2_30548 ( P1_R2238_U22 , P1_R2238_U66 , P1_R2238_U65 );
nand NAND2_30549 ( P1_R2238_U23 , P1_R2238_U48 , P1_R2238_U47 );
nand NAND2_30550 ( P1_R2238_U24 , P1_R2238_U53 , P1_R2238_U52 );
nand NAND2_30551 ( P1_R2238_U25 , P1_R2238_U58 , P1_R2238_U57 );
nand NAND2_30552 ( P1_R2238_U26 , P1_R2238_U63 , P1_R2238_U62 );
nand NAND2_30553 ( P1_R2238_U27 , P1_R2238_U37 , P1_R2238_U36 );
nand NAND2_30554 ( P1_R2238_U28 , P1_R2238_U33 , P1_R2238_U32 );
not NOT1_30555 ( P1_R2238_U29 , P1_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_30556 ( P1_R2238_U30 , P1_R2238_U9 );
nand NAND2_30557 ( P1_R2238_U31 , P1_R2238_U30 , P1_R2238_U10 );
nand NAND2_30558 ( P1_R2238_U32 , P1_R2238_U31 , P1_R2238_U29 );
nand NAND2_30559 ( P1_R2238_U33 , P1_INSTQUEUEWR_ADDR_REG_1_ , P1_R2238_U9 );
not NOT1_30560 ( P1_R2238_U34 , P1_R2238_U28 );
nand NAND2_30561 ( P1_R2238_U35 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_R2238_U12 );
nand NAND2_30562 ( P1_R2238_U36 , P1_R2238_U35 , P1_R2238_U28 );
nand NAND2_30563 ( P1_R2238_U37 , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_R2238_U11 );
not NOT1_30564 ( P1_R2238_U38 , P1_R2238_U27 );
nand NAND2_30565 ( P1_R2238_U39 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_R2238_U14 );
nand NAND2_30566 ( P1_R2238_U40 , P1_R2238_U39 , P1_R2238_U27 );
nand NAND2_30567 ( P1_R2238_U41 , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_R2238_U13 );
not NOT1_30568 ( P1_R2238_U42 , P1_R2238_U16 );
nand NAND2_30569 ( P1_R2238_U43 , P1_INSTQUEUEWR_ADDR_REG_4_ , P1_R2238_U17 );
nand NAND2_30570 ( P1_R2238_U44 , P1_R2238_U42 , P1_R2238_U43 );
nand NAND2_30571 ( P1_R2238_U45 , P1_INSTQUEUERD_ADDR_REG_4_ , P1_R2238_U15 );
nand NAND2_30572 ( P1_R2238_U46 , P1_INSTQUEUEWR_ADDR_REG_0_ , P1_R2238_U8 );
nand NAND2_30573 ( P1_R2238_U47 , P1_INSTQUEUERD_ADDR_REG_4_ , P1_R2238_U15 );
nand NAND2_30574 ( P1_R2238_U48 , P1_INSTQUEUEWR_ADDR_REG_4_ , P1_R2238_U17 );
not NOT1_30575 ( P1_R2238_U49 , P1_R2238_U23 );
nand NAND2_30576 ( P1_R2238_U50 , P1_R2238_U49 , P1_R2238_U42 );
nand NAND2_30577 ( P1_R2238_U51 , P1_R2238_U23 , P1_R2238_U16 );
nand NAND2_30578 ( P1_R2238_U52 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_R2238_U14 );
nand NAND2_30579 ( P1_R2238_U53 , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_R2238_U13 );
not NOT1_30580 ( P1_R2238_U54 , P1_R2238_U24 );
nand NAND2_30581 ( P1_R2238_U55 , P1_R2238_U38 , P1_R2238_U54 );
nand NAND2_30582 ( P1_R2238_U56 , P1_R2238_U24 , P1_R2238_U27 );
nand NAND2_30583 ( P1_R2238_U57 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_R2238_U12 );
nand NAND2_30584 ( P1_R2238_U58 , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_R2238_U11 );
not NOT1_30585 ( P1_R2238_U59 , P1_R2238_U25 );
nand NAND2_30586 ( P1_R2238_U60 , P1_R2238_U34 , P1_R2238_U59 );
nand NAND2_30587 ( P1_R2238_U61 , P1_R2238_U25 , P1_R2238_U28 );
nand NAND2_30588 ( P1_R2238_U62 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_R2238_U10 );
nand NAND2_30589 ( P1_R2238_U63 , P1_INSTQUEUEWR_ADDR_REG_1_ , P1_R2238_U29 );
not NOT1_30590 ( P1_R2238_U64 , P1_R2238_U26 );
nand NAND2_30591 ( P1_R2238_U65 , P1_R2238_U64 , P1_R2238_U30 );
nand NAND2_30592 ( P1_R2238_U66 , P1_R2238_U26 , P1_R2238_U9 );
nand NAND2_30593 ( P1_SUB_450_U6 , P1_SUB_450_U45 , P1_SUB_450_U44 );
nand NAND2_30594 ( P1_SUB_450_U7 , P1_SUB_450_U9 , P1_SUB_450_U46 );
not NOT1_30595 ( P1_SUB_450_U8 , P1_INSTQUEUERD_ADDR_REG_0_ );
nand NAND2_30596 ( P1_SUB_450_U9 , P1_INSTQUEUERD_ADDR_REG_0_ , P1_SUB_450_U18 );
not NOT1_30597 ( P1_SUB_450_U10 , P1_INSTQUEUEWR_ADDR_REG_1_ );
not NOT1_30598 ( P1_SUB_450_U11 , P1_INSTQUEUERD_ADDR_REG_2_ );
not NOT1_30599 ( P1_SUB_450_U12 , P1_INSTQUEUEWR_ADDR_REG_2_ );
not NOT1_30600 ( P1_SUB_450_U13 , P1_INSTQUEUERD_ADDR_REG_3_ );
not NOT1_30601 ( P1_SUB_450_U14 , P1_INSTQUEUEWR_ADDR_REG_3_ );
not NOT1_30602 ( P1_SUB_450_U15 , P1_INSTQUEUEWR_ADDR_REG_4_ );
nand NAND2_30603 ( P1_SUB_450_U16 , P1_SUB_450_U41 , P1_SUB_450_U40 );
not NOT1_30604 ( P1_SUB_450_U17 , P1_INSTQUEUERD_ADDR_REG_4_ );
not NOT1_30605 ( P1_SUB_450_U18 , P1_INSTQUEUEWR_ADDR_REG_0_ );
nand NAND2_30606 ( P1_SUB_450_U19 , P1_SUB_450_U51 , P1_SUB_450_U50 );
nand NAND2_30607 ( P1_SUB_450_U20 , P1_SUB_450_U56 , P1_SUB_450_U55 );
nand NAND2_30608 ( P1_SUB_450_U21 , P1_SUB_450_U61 , P1_SUB_450_U60 );
nand NAND2_30609 ( P1_SUB_450_U22 , P1_SUB_450_U66 , P1_SUB_450_U65 );
nand NAND2_30610 ( P1_SUB_450_U23 , P1_SUB_450_U48 , P1_SUB_450_U47 );
nand NAND2_30611 ( P1_SUB_450_U24 , P1_SUB_450_U53 , P1_SUB_450_U52 );
nand NAND2_30612 ( P1_SUB_450_U25 , P1_SUB_450_U58 , P1_SUB_450_U57 );
nand NAND2_30613 ( P1_SUB_450_U26 , P1_SUB_450_U63 , P1_SUB_450_U62 );
nand NAND2_30614 ( P1_SUB_450_U27 , P1_SUB_450_U37 , P1_SUB_450_U36 );
nand NAND2_30615 ( P1_SUB_450_U28 , P1_SUB_450_U33 , P1_SUB_450_U32 );
not NOT1_30616 ( P1_SUB_450_U29 , P1_INSTQUEUERD_ADDR_REG_1_ );
not NOT1_30617 ( P1_SUB_450_U30 , P1_SUB_450_U9 );
nand NAND2_30618 ( P1_SUB_450_U31 , P1_SUB_450_U30 , P1_SUB_450_U10 );
nand NAND2_30619 ( P1_SUB_450_U32 , P1_SUB_450_U31 , P1_SUB_450_U29 );
nand NAND2_30620 ( P1_SUB_450_U33 , P1_INSTQUEUEWR_ADDR_REG_1_ , P1_SUB_450_U9 );
not NOT1_30621 ( P1_SUB_450_U34 , P1_SUB_450_U28 );
nand NAND2_30622 ( P1_SUB_450_U35 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_SUB_450_U12 );
nand NAND2_30623 ( P1_SUB_450_U36 , P1_SUB_450_U35 , P1_SUB_450_U28 );
nand NAND2_30624 ( P1_SUB_450_U37 , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_SUB_450_U11 );
not NOT1_30625 ( P1_SUB_450_U38 , P1_SUB_450_U27 );
nand NAND2_30626 ( P1_SUB_450_U39 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_SUB_450_U14 );
nand NAND2_30627 ( P1_SUB_450_U40 , P1_SUB_450_U39 , P1_SUB_450_U27 );
nand NAND2_30628 ( P1_SUB_450_U41 , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_SUB_450_U13 );
not NOT1_30629 ( P1_SUB_450_U42 , P1_SUB_450_U16 );
nand NAND2_30630 ( P1_SUB_450_U43 , P1_INSTQUEUEWR_ADDR_REG_4_ , P1_SUB_450_U17 );
nand NAND2_30631 ( P1_SUB_450_U44 , P1_SUB_450_U42 , P1_SUB_450_U43 );
nand NAND2_30632 ( P1_SUB_450_U45 , P1_INSTQUEUERD_ADDR_REG_4_ , P1_SUB_450_U15 );
nand NAND2_30633 ( P1_SUB_450_U46 , P1_INSTQUEUEWR_ADDR_REG_0_ , P1_SUB_450_U8 );
nand NAND2_30634 ( P1_SUB_450_U47 , P1_INSTQUEUERD_ADDR_REG_4_ , P1_SUB_450_U15 );
nand NAND2_30635 ( P1_SUB_450_U48 , P1_INSTQUEUEWR_ADDR_REG_4_ , P1_SUB_450_U17 );
not NOT1_30636 ( P1_SUB_450_U49 , P1_SUB_450_U23 );
nand NAND2_30637 ( P1_SUB_450_U50 , P1_SUB_450_U49 , P1_SUB_450_U42 );
nand NAND2_30638 ( P1_SUB_450_U51 , P1_SUB_450_U23 , P1_SUB_450_U16 );
nand NAND2_30639 ( P1_SUB_450_U52 , P1_INSTQUEUERD_ADDR_REG_3_ , P1_SUB_450_U14 );
nand NAND2_30640 ( P1_SUB_450_U53 , P1_INSTQUEUEWR_ADDR_REG_3_ , P1_SUB_450_U13 );
not NOT1_30641 ( P1_SUB_450_U54 , P1_SUB_450_U24 );
nand NAND2_30642 ( P1_SUB_450_U55 , P1_SUB_450_U38 , P1_SUB_450_U54 );
nand NAND2_30643 ( P1_SUB_450_U56 , P1_SUB_450_U24 , P1_SUB_450_U27 );
nand NAND2_30644 ( P1_SUB_450_U57 , P1_INSTQUEUERD_ADDR_REG_2_ , P1_SUB_450_U12 );
nand NAND2_30645 ( P1_SUB_450_U58 , P1_INSTQUEUEWR_ADDR_REG_2_ , P1_SUB_450_U11 );
not NOT1_30646 ( P1_SUB_450_U59 , P1_SUB_450_U25 );
nand NAND2_30647 ( P1_SUB_450_U60 , P1_SUB_450_U34 , P1_SUB_450_U59 );
nand NAND2_30648 ( P1_SUB_450_U61 , P1_SUB_450_U25 , P1_SUB_450_U28 );
nand NAND2_30649 ( P1_SUB_450_U62 , P1_INSTQUEUERD_ADDR_REG_1_ , P1_SUB_450_U10 );
nand NAND2_30650 ( P1_SUB_450_U63 , P1_INSTQUEUEWR_ADDR_REG_1_ , P1_SUB_450_U29 );
not NOT1_30651 ( P1_SUB_450_U64 , P1_SUB_450_U26 );
nand NAND2_30652 ( P1_SUB_450_U65 , P1_SUB_450_U64 , P1_SUB_450_U30 );
nand NAND2_30653 ( P1_SUB_450_U66 , P1_SUB_450_U26 , P1_SUB_450_U9 );
not NOT1_30654 ( P1_ADD_371_U4 , P1_U3227 );
nand NAND2_30655 ( P1_ADD_371_U5 , P1_ADD_371_U23 , P1_ADD_371_U31 );
and AND2_30656 ( P1_ADD_371_U6 , P1_ADD_371_U22 , P1_ADD_371_U30 );
not NOT1_30657 ( P1_ADD_371_U7 , P1_U3228 );
not NOT1_30658 ( P1_ADD_371_U8 , P1_U3230 );
nand NAND2_30659 ( P1_ADD_371_U9 , P1_U3230 , P1_ADD_371_U23 );
not NOT1_30660 ( P1_ADD_371_U10 , P1_U3231 );
nand NAND2_30661 ( P1_ADD_371_U11 , P1_U3231 , P1_ADD_371_U28 );
not NOT1_30662 ( P1_ADD_371_U12 , P1_U3232 );
not NOT1_30663 ( P1_ADD_371_U13 , P1_U3233 );
nand NAND2_30664 ( P1_ADD_371_U14 , P1_U3232 , P1_ADD_371_U29 );
not NOT1_30665 ( P1_ADD_371_U15 , P1_U3229 );
not NOT1_30666 ( P1_ADD_371_U16 , P1_U3234 );
nand NAND2_30667 ( P1_ADD_371_U17 , P1_ADD_371_U34 , P1_ADD_371_U33 );
nand NAND2_30668 ( P1_ADD_371_U18 , P1_ADD_371_U36 , P1_ADD_371_U35 );
nand NAND2_30669 ( P1_ADD_371_U19 , P1_ADD_371_U38 , P1_ADD_371_U37 );
nand NAND2_30670 ( P1_ADD_371_U20 , P1_ADD_371_U42 , P1_ADD_371_U41 );
nand NAND2_30671 ( P1_ADD_371_U21 , P1_ADD_371_U44 , P1_ADD_371_U43 );
and AND2_30672 ( P1_ADD_371_U22 , P1_U3234 , P1_U3233 );
nand NAND2_30673 ( P1_ADD_371_U23 , P1_ADD_371_U15 , P1_ADD_371_U26 );
and AND2_30674 ( P1_ADD_371_U24 , P1_ADD_371_U40 , P1_ADD_371_U39 );
nand NAND2_30675 ( P1_ADD_371_U25 , P1_ADD_371_U30 , P1_U3233 );
nand NAND2_30676 ( P1_ADD_371_U26 , P1_U3228 , P1_U3227 );
not NOT1_30677 ( P1_ADD_371_U27 , P1_ADD_371_U23 );
not NOT1_30678 ( P1_ADD_371_U28 , P1_ADD_371_U9 );
not NOT1_30679 ( P1_ADD_371_U29 , P1_ADD_371_U11 );
not NOT1_30680 ( P1_ADD_371_U30 , P1_ADD_371_U14 );
nand NAND3_30681 ( P1_ADD_371_U31 , P1_U3228 , P1_U3227 , P1_U3229 );
not NOT1_30682 ( P1_ADD_371_U32 , P1_ADD_371_U25 );
nand NAND2_30683 ( P1_ADD_371_U33 , P1_U3233 , P1_ADD_371_U14 );
nand NAND2_30684 ( P1_ADD_371_U34 , P1_ADD_371_U30 , P1_ADD_371_U13 );
nand NAND2_30685 ( P1_ADD_371_U35 , P1_U3231 , P1_ADD_371_U9 );
nand NAND2_30686 ( P1_ADD_371_U36 , P1_ADD_371_U28 , P1_ADD_371_U10 );
nand NAND2_30687 ( P1_ADD_371_U37 , P1_U3232 , P1_ADD_371_U11 );
nand NAND2_30688 ( P1_ADD_371_U38 , P1_ADD_371_U29 , P1_ADD_371_U12 );
nand NAND2_30689 ( P1_ADD_371_U39 , P1_U3230 , P1_ADD_371_U23 );
nand NAND2_30690 ( P1_ADD_371_U40 , P1_ADD_371_U27 , P1_ADD_371_U8 );
nand NAND2_30691 ( P1_ADD_371_U41 , P1_U3228 , P1_ADD_371_U4 );
nand NAND2_30692 ( P1_ADD_371_U42 , P1_U3227 , P1_ADD_371_U7 );
nand NAND2_30693 ( P1_ADD_371_U43 , P1_U3234 , P1_ADD_371_U25 );
nand NAND2_30694 ( P1_ADD_371_U44 , P1_ADD_371_U32 , P1_ADD_371_U16 );
not NOT1_30695 ( P1_ADD_405_U4 , P1_INSTADDRPOINTER_REG_0_ );
nand NAND2_30696 ( P1_ADD_405_U5 , P1_ADD_405_U94 , P1_ADD_405_U125 );
not NOT1_30697 ( P1_ADD_405_U6 , P1_INSTADDRPOINTER_REG_1_ );
not NOT1_30698 ( P1_ADD_405_U7 , P1_INSTADDRPOINTER_REG_3_ );
nand NAND2_30699 ( P1_ADD_405_U8 , P1_INSTADDRPOINTER_REG_3_ , P1_ADD_405_U94 );
not NOT1_30700 ( P1_ADD_405_U9 , P1_INSTADDRPOINTER_REG_4_ );
nand NAND2_30701 ( P1_ADD_405_U10 , P1_INSTADDRPOINTER_REG_4_ , P1_ADD_405_U98 );
not NOT1_30702 ( P1_ADD_405_U11 , P1_INSTADDRPOINTER_REG_5_ );
not NOT1_30703 ( P1_ADD_405_U12 , P1_INSTADDRPOINTER_REG_6_ );
nand NAND2_30704 ( P1_ADD_405_U13 , P1_INSTADDRPOINTER_REG_5_ , P1_ADD_405_U99 );
nand NAND2_30705 ( P1_ADD_405_U14 , P1_ADD_405_U100 , P1_INSTADDRPOINTER_REG_6_ );
not NOT1_30706 ( P1_ADD_405_U15 , P1_INSTADDRPOINTER_REG_7_ );
nand NAND2_30707 ( P1_ADD_405_U16 , P1_INSTADDRPOINTER_REG_7_ , P1_ADD_405_U101 );
not NOT1_30708 ( P1_ADD_405_U17 , P1_INSTADDRPOINTER_REG_8_ );
nand NAND2_30709 ( P1_ADD_405_U18 , P1_INSTADDRPOINTER_REG_8_ , P1_ADD_405_U102 );
not NOT1_30710 ( P1_ADD_405_U19 , P1_INSTADDRPOINTER_REG_9_ );
nand NAND2_30711 ( P1_ADD_405_U20 , P1_INSTADDRPOINTER_REG_9_ , P1_ADD_405_U103 );
not NOT1_30712 ( P1_ADD_405_U21 , P1_INSTADDRPOINTER_REG_10_ );
nand NAND2_30713 ( P1_ADD_405_U22 , P1_INSTADDRPOINTER_REG_10_ , P1_ADD_405_U104 );
not NOT1_30714 ( P1_ADD_405_U23 , P1_INSTADDRPOINTER_REG_11_ );
nand NAND2_30715 ( P1_ADD_405_U24 , P1_INSTADDRPOINTER_REG_11_ , P1_ADD_405_U105 );
not NOT1_30716 ( P1_ADD_405_U25 , P1_INSTADDRPOINTER_REG_12_ );
nand NAND2_30717 ( P1_ADD_405_U26 , P1_INSTADDRPOINTER_REG_12_ , P1_ADD_405_U106 );
not NOT1_30718 ( P1_ADD_405_U27 , P1_INSTADDRPOINTER_REG_13_ );
nand NAND2_30719 ( P1_ADD_405_U28 , P1_INSTADDRPOINTER_REG_13_ , P1_ADD_405_U107 );
not NOT1_30720 ( P1_ADD_405_U29 , P1_INSTADDRPOINTER_REG_14_ );
nand NAND2_30721 ( P1_ADD_405_U30 , P1_INSTADDRPOINTER_REG_14_ , P1_ADD_405_U108 );
not NOT1_30722 ( P1_ADD_405_U31 , P1_INSTADDRPOINTER_REG_15_ );
nand NAND2_30723 ( P1_ADD_405_U32 , P1_INSTADDRPOINTER_REG_15_ , P1_ADD_405_U109 );
not NOT1_30724 ( P1_ADD_405_U33 , P1_INSTADDRPOINTER_REG_16_ );
nand NAND2_30725 ( P1_ADD_405_U34 , P1_INSTADDRPOINTER_REG_16_ , P1_ADD_405_U110 );
not NOT1_30726 ( P1_ADD_405_U35 , P1_INSTADDRPOINTER_REG_17_ );
nand NAND2_30727 ( P1_ADD_405_U36 , P1_INSTADDRPOINTER_REG_17_ , P1_ADD_405_U111 );
not NOT1_30728 ( P1_ADD_405_U37 , P1_INSTADDRPOINTER_REG_18_ );
nand NAND2_30729 ( P1_ADD_405_U38 , P1_INSTADDRPOINTER_REG_18_ , P1_ADD_405_U112 );
not NOT1_30730 ( P1_ADD_405_U39 , P1_INSTADDRPOINTER_REG_19_ );
nand NAND2_30731 ( P1_ADD_405_U40 , P1_INSTADDRPOINTER_REG_19_ , P1_ADD_405_U113 );
not NOT1_30732 ( P1_ADD_405_U41 , P1_INSTADDRPOINTER_REG_20_ );
nand NAND2_30733 ( P1_ADD_405_U42 , P1_INSTADDRPOINTER_REG_20_ , P1_ADD_405_U114 );
not NOT1_30734 ( P1_ADD_405_U43 , P1_INSTADDRPOINTER_REG_21_ );
nand NAND2_30735 ( P1_ADD_405_U44 , P1_INSTADDRPOINTER_REG_21_ , P1_ADD_405_U115 );
not NOT1_30736 ( P1_ADD_405_U45 , P1_INSTADDRPOINTER_REG_22_ );
nand NAND2_30737 ( P1_ADD_405_U46 , P1_INSTADDRPOINTER_REG_22_ , P1_ADD_405_U116 );
not NOT1_30738 ( P1_ADD_405_U47 , P1_INSTADDRPOINTER_REG_23_ );
nand NAND2_30739 ( P1_ADD_405_U48 , P1_INSTADDRPOINTER_REG_23_ , P1_ADD_405_U117 );
not NOT1_30740 ( P1_ADD_405_U49 , P1_INSTADDRPOINTER_REG_24_ );
nand NAND2_30741 ( P1_ADD_405_U50 , P1_INSTADDRPOINTER_REG_24_ , P1_ADD_405_U118 );
not NOT1_30742 ( P1_ADD_405_U51 , P1_INSTADDRPOINTER_REG_25_ );
nand NAND2_30743 ( P1_ADD_405_U52 , P1_INSTADDRPOINTER_REG_25_ , P1_ADD_405_U119 );
not NOT1_30744 ( P1_ADD_405_U53 , P1_INSTADDRPOINTER_REG_26_ );
nand NAND2_30745 ( P1_ADD_405_U54 , P1_INSTADDRPOINTER_REG_26_ , P1_ADD_405_U120 );
not NOT1_30746 ( P1_ADD_405_U55 , P1_INSTADDRPOINTER_REG_27_ );
nand NAND2_30747 ( P1_ADD_405_U56 , P1_INSTADDRPOINTER_REG_27_ , P1_ADD_405_U121 );
not NOT1_30748 ( P1_ADD_405_U57 , P1_INSTADDRPOINTER_REG_28_ );
nand NAND2_30749 ( P1_ADD_405_U58 , P1_INSTADDRPOINTER_REG_28_ , P1_ADD_405_U122 );
not NOT1_30750 ( P1_ADD_405_U59 , P1_INSTADDRPOINTER_REG_29_ );
not NOT1_30751 ( P1_ADD_405_U60 , P1_INSTADDRPOINTER_REG_30_ );
nand NAND2_30752 ( P1_ADD_405_U61 , P1_INSTADDRPOINTER_REG_29_ , P1_ADD_405_U123 );
not NOT1_30753 ( P1_ADD_405_U62 , P1_INSTADDRPOINTER_REG_2_ );
nand NAND2_30754 ( P1_ADD_405_U63 , P1_ADD_405_U128 , P1_ADD_405_U127 );
nand NAND2_30755 ( P1_ADD_405_U64 , P1_ADD_405_U130 , P1_ADD_405_U129 );
nand NAND2_30756 ( P1_ADD_405_U65 , P1_ADD_405_U132 , P1_ADD_405_U131 );
nand NAND2_30757 ( P1_ADD_405_U66 , P1_ADD_405_U134 , P1_ADD_405_U133 );
nand NAND2_30758 ( P1_ADD_405_U67 , P1_ADD_405_U136 , P1_ADD_405_U135 );
nand NAND2_30759 ( P1_ADD_405_U68 , P1_ADD_405_U138 , P1_ADD_405_U137 );
nand NAND2_30760 ( P1_ADD_405_U69 , P1_ADD_405_U140 , P1_ADD_405_U139 );
nand NAND2_30761 ( P1_ADD_405_U70 , P1_ADD_405_U142 , P1_ADD_405_U141 );
nand NAND2_30762 ( P1_ADD_405_U71 , P1_ADD_405_U144 , P1_ADD_405_U143 );
nand NAND2_30763 ( P1_ADD_405_U72 , P1_ADD_405_U146 , P1_ADD_405_U145 );
nand NAND2_30764 ( P1_ADD_405_U73 , P1_ADD_405_U148 , P1_ADD_405_U147 );
nand NAND2_30765 ( P1_ADD_405_U74 , P1_ADD_405_U150 , P1_ADD_405_U149 );
nand NAND2_30766 ( P1_ADD_405_U75 , P1_ADD_405_U152 , P1_ADD_405_U151 );
nand NAND2_30767 ( P1_ADD_405_U76 , P1_ADD_405_U154 , P1_ADD_405_U153 );
nand NAND2_30768 ( P1_ADD_405_U77 , P1_ADD_405_U156 , P1_ADD_405_U155 );
nand NAND2_30769 ( P1_ADD_405_U78 , P1_ADD_405_U158 , P1_ADD_405_U157 );
nand NAND2_30770 ( P1_ADD_405_U79 , P1_ADD_405_U160 , P1_ADD_405_U159 );
nand NAND2_30771 ( P1_ADD_405_U80 , P1_ADD_405_U162 , P1_ADD_405_U161 );
nand NAND2_30772 ( P1_ADD_405_U81 , P1_ADD_405_U164 , P1_ADD_405_U163 );
nand NAND2_30773 ( P1_ADD_405_U82 , P1_ADD_405_U166 , P1_ADD_405_U165 );
nand NAND2_30774 ( P1_ADD_405_U83 , P1_ADD_405_U168 , P1_ADD_405_U167 );
nand NAND2_30775 ( P1_ADD_405_U84 , P1_ADD_405_U170 , P1_ADD_405_U169 );
nand NAND2_30776 ( P1_ADD_405_U85 , P1_ADD_405_U174 , P1_ADD_405_U173 );
nand NAND2_30777 ( P1_ADD_405_U86 , P1_ADD_405_U176 , P1_ADD_405_U175 );

// 67 Additional buffers.
buf add_BUF1_1 ( P3_DATAO_REG_0_ , P3_DATAO_REG_0__EXTRA );
buf add_BUF1_2 ( P3_DATAO_REG_1_ , P3_DATAO_REG_1__EXTRA );
buf add_BUF1_3 ( P3_DATAO_REG_2_ , P3_DATAO_REG_2__EXTRA );
buf add_BUF1_4 ( P3_DATAO_REG_3_ , P3_DATAO_REG_3__EXTRA );
buf add_BUF1_5 ( P3_DATAO_REG_4_ , P3_DATAO_REG_4__EXTRA );
buf add_BUF1_6 ( P3_DATAO_REG_5_ , P3_DATAO_REG_5__EXTRA );
buf add_BUF1_7 ( P3_DATAO_REG_6_ , P3_DATAO_REG_6__EXTRA );
buf add_BUF1_8 ( P3_DATAO_REG_7_ , P3_DATAO_REG_7__EXTRA );
buf add_BUF1_9 ( P3_DATAO_REG_8_ , P3_DATAO_REG_8__EXTRA );
buf add_BUF1_10 ( P3_DATAO_REG_9_ , P3_DATAO_REG_9__EXTRA );
buf add_BUF1_11 ( P3_DATAO_REG_10_ , P3_DATAO_REG_10__EXTRA );
buf add_BUF1_12 ( P3_DATAO_REG_11_ , P3_DATAO_REG_11__EXTRA );
buf add_BUF1_13 ( P3_DATAO_REG_12_ , P3_DATAO_REG_12__EXTRA );
buf add_BUF1_14 ( P3_DATAO_REG_13_ , P3_DATAO_REG_13__EXTRA );
buf add_BUF1_15 ( P3_DATAO_REG_14_ , P3_DATAO_REG_14__EXTRA );
buf add_BUF1_16 ( P3_DATAO_REG_15_ , P3_DATAO_REG_15__EXTRA );
buf add_BUF1_17 ( P3_DATAO_REG_16_ , P3_DATAO_REG_16__EXTRA );
buf add_BUF1_18 ( P3_DATAO_REG_17_ , P3_DATAO_REG_17__EXTRA );
buf add_BUF1_19 ( P3_DATAO_REG_18_ , P3_DATAO_REG_18__EXTRA );
buf add_BUF1_20 ( P3_DATAO_REG_19_ , P3_DATAO_REG_19__EXTRA );
buf add_BUF1_21 ( P3_DATAO_REG_20_ , P3_DATAO_REG_20__EXTRA );
buf add_BUF1_22 ( P3_DATAO_REG_21_ , P3_DATAO_REG_21__EXTRA );
buf add_BUF1_23 ( P3_DATAO_REG_22_ , P3_DATAO_REG_22__EXTRA );
buf add_BUF1_24 ( P3_DATAO_REG_23_ , P3_DATAO_REG_23__EXTRA );
buf add_BUF1_25 ( P3_DATAO_REG_24_ , P3_DATAO_REG_24__EXTRA );
buf add_BUF1_26 ( P3_DATAO_REG_25_ , P3_DATAO_REG_25__EXTRA );
buf add_BUF1_27 ( P3_DATAO_REG_26_ , P3_DATAO_REG_26__EXTRA );
buf add_BUF1_28 ( P3_DATAO_REG_27_ , P3_DATAO_REG_27__EXTRA );
buf add_BUF1_29 ( P3_DATAO_REG_28_ , P3_DATAO_REG_28__EXTRA );
buf add_BUF1_30 ( P3_DATAO_REG_29_ , P3_DATAO_REG_29__EXTRA );
buf add_BUF1_31 ( P3_DATAO_REG_30_ , P3_DATAO_REG_30__EXTRA );
buf add_BUF1_32 ( P3_DATAO_REG_31_ , P3_DATAO_REG_31__EXTRA );
buf add_BUF1_33 ( P3_W_R_N_REG , P3_W_R_N_REG_EXTRA );
buf add_BUF1_34 ( P3_D_C_N_REG , P3_D_C_N_REG_EXTRA );
buf add_BUF1_35 ( P3_M_IO_N_REG , P3_M_IO_N_REG_EXTRA );
buf add_BUF1_36 ( P3_ADS_N_REG , P3_ADS_N_REG_EXTRA );
buf add_BUF1_37 ( P1_ADDRESS_REG_29_ , P1_ADDRESS_REG_29__EXTRA );
buf add_BUF1_38 ( P1_ADDRESS_REG_28_ , P1_ADDRESS_REG_28__EXTRA );
buf add_BUF1_39 ( P1_ADDRESS_REG_27_ , P1_ADDRESS_REG_27__EXTRA );
buf add_BUF1_40 ( P1_ADDRESS_REG_26_ , P1_ADDRESS_REG_26__EXTRA );
buf add_BUF1_41 ( P1_ADDRESS_REG_25_ , P1_ADDRESS_REG_25__EXTRA );
buf add_BUF1_42 ( P1_ADDRESS_REG_24_ , P1_ADDRESS_REG_24__EXTRA );
buf add_BUF1_43 ( P1_ADDRESS_REG_23_ , P1_ADDRESS_REG_23__EXTRA );
buf add_BUF1_44 ( P1_ADDRESS_REG_22_ , P1_ADDRESS_REG_22__EXTRA );
buf add_BUF1_45 ( P1_ADDRESS_REG_21_ , P1_ADDRESS_REG_21__EXTRA );
buf add_BUF1_46 ( P1_ADDRESS_REG_20_ , P1_ADDRESS_REG_20__EXTRA );
buf add_BUF1_47 ( P1_ADDRESS_REG_19_ , P1_ADDRESS_REG_19__EXTRA );
buf add_BUF1_48 ( P1_ADDRESS_REG_18_ , P1_ADDRESS_REG_18__EXTRA );
buf add_BUF1_49 ( P1_ADDRESS_REG_17_ , P1_ADDRESS_REG_17__EXTRA );
buf add_BUF1_50 ( P1_ADDRESS_REG_16_ , P1_ADDRESS_REG_16__EXTRA );
buf add_BUF1_51 ( P1_ADDRESS_REG_15_ , P1_ADDRESS_REG_15__EXTRA );
buf add_BUF1_52 ( P1_ADDRESS_REG_14_ , P1_ADDRESS_REG_14__EXTRA );
buf add_BUF1_53 ( P1_ADDRESS_REG_13_ , P1_ADDRESS_REG_13__EXTRA );
buf add_BUF1_54 ( P1_ADDRESS_REG_12_ , P1_ADDRESS_REG_12__EXTRA );
buf add_BUF1_55 ( P1_ADDRESS_REG_11_ , P1_ADDRESS_REG_11__EXTRA );
buf add_BUF1_56 ( P1_ADDRESS_REG_10_ , P1_ADDRESS_REG_10__EXTRA );
buf add_BUF1_57 ( P1_ADDRESS_REG_9_ , P1_ADDRESS_REG_9__EXTRA );
buf add_BUF1_58 ( P1_ADDRESS_REG_8_ , P1_ADDRESS_REG_8__EXTRA );
buf add_BUF1_59 ( P1_ADDRESS_REG_7_ , P1_ADDRESS_REG_7__EXTRA );
buf add_BUF1_60 ( P1_ADDRESS_REG_6_ , P1_ADDRESS_REG_6__EXTRA );
buf add_BUF1_61 ( P1_ADDRESS_REG_5_ , P1_ADDRESS_REG_5__EXTRA );
buf add_BUF1_62 ( P1_ADDRESS_REG_4_ , P1_ADDRESS_REG_4__EXTRA );
buf add_BUF1_63 ( P1_ADDRESS_REG_3_ , P1_ADDRESS_REG_3__EXTRA );
buf add_BUF1_64 ( P1_ADDRESS_REG_2_ , P1_ADDRESS_REG_2__EXTRA );
buf add_BUF1_65 ( P1_ADDRESS_REG_1_ , P1_ADDRESS_REG_1__EXTRA );
buf add_BUF1_66 ( P1_ADDRESS_REG_0_ , P1_ADDRESS_REG_0__EXTRA );
buf add_BUF1_67 ( P1_ADS_N_REG , P1_ADS_N_REG_EXTRA );

endmodule
